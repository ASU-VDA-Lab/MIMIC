module fake_ariane_42_n_2116 (n_83, n_8, n_56, n_60, n_170, n_190, n_160, n_64, n_179, n_180, n_119, n_124, n_167, n_90, n_195, n_38, n_47, n_110, n_153, n_18, n_197, n_86, n_75, n_89, n_67, n_176, n_149, n_34, n_158, n_172, n_69, n_95, n_175, n_92, n_143, n_183, n_203, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_181, n_152, n_120, n_169, n_106, n_12, n_53, n_173, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_156, n_49, n_20, n_174, n_100, n_17, n_50, n_187, n_132, n_62, n_147, n_204, n_200, n_51, n_166, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_199, n_91, n_159, n_107, n_189, n_72, n_105, n_128, n_44, n_30, n_82, n_178, n_31, n_42, n_57, n_131, n_201, n_70, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_188, n_185, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_198, n_148, n_164, n_52, n_157, n_184, n_177, n_135, n_73, n_77, n_171, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_182, n_196, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_191, n_151, n_136, n_192, n_28, n_80, n_146, n_194, n_97, n_154, n_142, n_161, n_14, n_163, n_88, n_186, n_141, n_68, n_116, n_104, n_202, n_145, n_78, n_193, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_2116);

input n_83;
input n_8;
input n_56;
input n_60;
input n_170;
input n_190;
input n_160;
input n_64;
input n_179;
input n_180;
input n_119;
input n_124;
input n_167;
input n_90;
input n_195;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_197;
input n_86;
input n_75;
input n_89;
input n_67;
input n_176;
input n_149;
input n_34;
input n_158;
input n_172;
input n_69;
input n_95;
input n_175;
input n_92;
input n_143;
input n_183;
input n_203;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_181;
input n_152;
input n_120;
input n_169;
input n_106;
input n_12;
input n_53;
input n_173;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_156;
input n_49;
input n_20;
input n_174;
input n_100;
input n_17;
input n_50;
input n_187;
input n_132;
input n_62;
input n_147;
input n_204;
input n_200;
input n_51;
input n_166;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_199;
input n_91;
input n_159;
input n_107;
input n_189;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_178;
input n_31;
input n_42;
input n_57;
input n_131;
input n_201;
input n_70;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_188;
input n_185;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_198;
input n_148;
input n_164;
input n_52;
input n_157;
input n_184;
input n_177;
input n_135;
input n_73;
input n_77;
input n_171;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_182;
input n_196;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_191;
input n_151;
input n_136;
input n_192;
input n_28;
input n_80;
input n_146;
input n_194;
input n_97;
input n_154;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_186;
input n_141;
input n_68;
input n_116;
input n_104;
input n_202;
input n_145;
input n_78;
input n_193;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_2116;

wire n_913;
wire n_1681;
wire n_1486;
wire n_1507;
wire n_1938;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_1250;
wire n_2030;
wire n_1169;
wire n_789;
wire n_850;
wire n_1916;
wire n_610;
wire n_245;
wire n_1713;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_2002;
wire n_1463;
wire n_1238;
wire n_2011;
wire n_1515;
wire n_817;
wire n_1837;
wire n_924;
wire n_781;
wire n_2013;
wire n_1566;
wire n_717;
wire n_2006;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_1706;
wire n_524;
wire n_1214;
wire n_634;
wire n_1839;
wire n_1246;
wire n_1138;
wire n_214;
wire n_2042;
wire n_1853;
wire n_764;
wire n_1503;
wire n_462;
wire n_1196;
wire n_1181;
wire n_1999;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1745;
wire n_1366;
wire n_232;
wire n_2084;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1835;
wire n_1457;
wire n_377;
wire n_1682;
wire n_1836;
wire n_520;
wire n_870;
wire n_1453;
wire n_279;
wire n_958;
wire n_945;
wire n_813;
wire n_419;
wire n_1985;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1909;
wire n_1184;
wire n_1961;
wire n_1535;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_1979;
wire n_1277;
wire n_2107;
wire n_1746;
wire n_829;
wire n_1761;
wire n_1062;
wire n_339;
wire n_738;
wire n_1690;
wire n_672;
wire n_740;
wire n_1283;
wire n_1974;
wire n_1736;
wire n_1018;
wire n_259;
wire n_953;
wire n_1364;
wire n_1888;
wire n_1224;
wire n_2109;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_1688;
wire n_989;
wire n_645;
wire n_242;
wire n_1944;
wire n_331;
wire n_559;
wire n_267;
wire n_495;
wire n_1988;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_1936;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_2078;
wire n_1145;
wire n_971;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_2049;
wire n_1522;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_1404;
wire n_868;
wire n_1847;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1851;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_1676;
wire n_1085;
wire n_277;
wire n_1636;
wire n_432;
wire n_293;
wire n_823;
wire n_1900;
wire n_620;
wire n_1074;
wire n_859;
wire n_1765;
wire n_1889;
wire n_587;
wire n_1977;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_206;
wire n_352;
wire n_899;
wire n_1703;
wire n_611;
wire n_1295;
wire n_2060;
wire n_1850;
wire n_365;
wire n_238;
wire n_2004;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_334;
wire n_661;
wire n_2098;
wire n_1751;
wire n_300;
wire n_533;
wire n_1917;
wire n_1924;
wire n_438;
wire n_1654;
wire n_1560;
wire n_1548;
wire n_1811;
wire n_2045;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_1840;
wire n_376;
wire n_512;
wire n_1597;
wire n_1771;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_2061;
wire n_2094;
wire n_1354;
wire n_1790;
wire n_1213;
wire n_237;
wire n_2043;
wire n_780;
wire n_1918;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1949;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_2077;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_209;
wire n_490;
wire n_1461;
wire n_1391;
wire n_1947;
wire n_225;
wire n_1599;
wire n_1876;
wire n_1006;
wire n_1830;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_2038;
wire n_1838;
wire n_1594;
wire n_680;
wire n_1935;
wire n_287;
wire n_1716;
wire n_302;
wire n_1872;
wire n_380;
wire n_1585;
wire n_1432;
wire n_249;
wire n_1108;
wire n_355;
wire n_212;
wire n_851;
wire n_444;
wire n_1590;
wire n_1351;
wire n_1274;
wire n_257;
wire n_652;
wire n_1819;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_1833;
wire n_407;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_1884;
wire n_460;
wire n_1555;
wire n_1842;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_966;
wire n_992;
wire n_955;
wire n_1182;
wire n_794;
wire n_1692;
wire n_1562;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_288;
wire n_1292;
wire n_1178;
wire n_1972;
wire n_2015;
wire n_1435;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_2072;
wire n_306;
wire n_436;
wire n_324;
wire n_2087;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_437;
wire n_967;
wire n_274;
wire n_337;
wire n_1083;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1787;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_1717;
wire n_1812;
wire n_824;
wire n_428;
wire n_892;
wire n_1880;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_1855;
wire n_2100;
wire n_990;
wire n_1623;
wire n_1903;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_1932;
wire n_1780;
wire n_1970;
wire n_1920;
wire n_2083;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1911;
wire n_1825;
wire n_1908;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1832;
wire n_1841;
wire n_1680;
wire n_2066;
wire n_964;
wire n_1627;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_1731;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_1914;
wire n_934;
wire n_1447;
wire n_1220;
wire n_356;
wire n_2019;
wire n_698;
wire n_1674;
wire n_2021;
wire n_2025;
wire n_1992;
wire n_307;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_1633;
wire n_404;
wire n_1913;
wire n_2069;
wire n_1058;
wire n_347;
wire n_1042;
wire n_1234;
wire n_479;
wire n_1578;
wire n_1455;
wire n_299;
wire n_836;
wire n_1279;
wire n_564;
wire n_205;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_1689;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_1728;
wire n_370;
wire n_706;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_2041;
wire n_2113;
wire n_1933;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_1817;
wire n_552;
wire n_348;
wire n_670;
wire n_1826;
wire n_379;
wire n_264;
wire n_441;
wire n_1951;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_1618;
wire n_1869;
wire n_1743;
wire n_905;
wire n_207;
wire n_720;
wire n_926;
wire n_1943;
wire n_1802;
wire n_2112;
wire n_1163;
wire n_1795;
wire n_1384;
wire n_1868;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_2099;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1879;
wire n_1886;
wire n_1648;
wire n_1413;
wire n_855;
wire n_808;
wire n_1365;
wire n_553;
wire n_2059;
wire n_1439;
wire n_814;
wire n_578;
wire n_2074;
wire n_1665;
wire n_1287;
wire n_405;
wire n_1611;
wire n_320;
wire n_1414;
wire n_1134;
wire n_2067;
wire n_1484;
wire n_1901;
wire n_647;
wire n_2055;
wire n_2027;
wire n_1423;
wire n_600;
wire n_481;
wire n_1053;
wire n_1609;
wire n_1939;
wire n_1906;
wire n_529;
wire n_1899;
wire n_502;
wire n_218;
wire n_1467;
wire n_247;
wire n_1828;
wire n_1798;
wire n_1304;
wire n_1608;
wire n_1744;
wire n_1105;
wire n_547;
wire n_439;
wire n_604;
wire n_677;
wire n_478;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_2102;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_2023;
wire n_1278;
wire n_707;
wire n_983;
wire n_590;
wire n_699;
wire n_727;
wire n_301;
wire n_1726;
wire n_2075;
wire n_1945;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_2031;
wire n_325;
wire n_1740;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_1963;
wire n_729;
wire n_887;
wire n_2057;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_1693;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1823;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_2033;
wire n_233;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_221;
wire n_321;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1863;
wire n_1763;
wire n_1666;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_281;
wire n_1859;
wire n_262;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_1883;
wire n_1969;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_1667;
wire n_845;
wire n_888;
wire n_1649;
wire n_1677;
wire n_1927;
wire n_1297;
wire n_551;
wire n_417;
wire n_1708;
wire n_343;
wire n_1222;
wire n_1844;
wire n_582;
wire n_1957;
wire n_1953;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_1919;
wire n_534;
wire n_1791;
wire n_1894;
wire n_1460;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_1898;
wire n_451;
wire n_745;
wire n_1741;
wire n_1572;
wire n_1907;
wire n_1793;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1975;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_769;
wire n_1797;
wire n_1753;
wire n_1990;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_1895;
wire n_982;
wire n_1800;
wire n_915;
wire n_215;
wire n_1075;
wire n_2008;
wire n_454;
wire n_298;
wire n_1331;
wire n_1890;
wire n_1529;
wire n_1227;
wire n_655;
wire n_1734;
wire n_1860;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_1700;
wire n_659;
wire n_1332;
wire n_509;
wire n_1854;
wire n_666;
wire n_1747;
wire n_2071;
wire n_430;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_2082;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1766;
wire n_1338;
wire n_1342;
wire n_456;
wire n_1867;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_521;
wire n_873;
wire n_1301;
wire n_1748;
wire n_1966;
wire n_1243;
wire n_1400;
wire n_342;
wire n_2035;
wire n_1466;
wire n_1513;
wire n_1527;
wire n_358;
wire n_1783;
wire n_608;
wire n_1538;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1993;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1954;
wire n_1668;
wire n_1878;
wire n_1605;
wire n_1078;
wire n_266;
wire n_1897;
wire n_1161;
wire n_811;
wire n_624;
wire n_876;
wire n_791;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_687;
wire n_797;
wire n_2026;
wire n_1786;
wire n_480;
wire n_1327;
wire n_1475;
wire n_211;
wire n_642;
wire n_1804;
wire n_2106;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_1757;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_2091;
wire n_393;
wire n_1632;
wire n_1769;
wire n_474;
wire n_1929;
wire n_1950;
wire n_805;
wire n_2032;
wire n_2090;
wire n_295;
wire n_1658;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_730;
wire n_386;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1997;
wire n_1137;
wire n_1873;
wire n_1258;
wire n_640;
wire n_463;
wire n_1524;
wire n_1476;
wire n_1733;
wire n_1856;
wire n_2016;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1874;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_1807;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_1784;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_283;
wire n_806;
wire n_1984;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_1824;
wire n_643;
wire n_1492;
wire n_226;
wire n_1441;
wire n_1822;
wire n_682;
wire n_1616;
wire n_819;
wire n_1971;
wire n_586;
wire n_1324;
wire n_1429;
wire n_2064;
wire n_1778;
wire n_1776;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1759;
wire n_1829;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_2022;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_1815;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_1864;
wire n_1887;
wire n_1208;
wire n_1987;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1577;
wire n_1448;
wire n_1009;
wire n_230;
wire n_1133;
wire n_883;
wire n_473;
wire n_1852;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_594;
wire n_1995;
wire n_1877;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_1849;
wire n_2076;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_2001;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_1201;
wire n_1288;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_2070;
wire n_426;
wire n_433;
wire n_398;
wire n_210;
wire n_1090;
wire n_1367;
wire n_2044;
wire n_253;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_224;
wire n_894;
wire n_1380;
wire n_1624;
wire n_1801;
wire n_420;
wire n_1291;
wire n_562;
wire n_2020;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1882;
wire n_1976;
wire n_1023;
wire n_1881;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_1958;
wire n_467;
wire n_1511;
wire n_1422;
wire n_1965;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_1641;
wire n_538;
wire n_1517;
wire n_2036;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_2003;
wire n_1307;
wire n_1128;
wire n_2053;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1921;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1955;
wire n_2110;
wire n_1773;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_1948;
wire n_810;
wire n_1290;
wire n_1959;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_236;
wire n_683;
wire n_601;
wire n_565;
wire n_628;
wire n_1300;
wire n_1960;
wire n_2068;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_1968;
wire n_1885;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_1978;
wire n_414;
wire n_571;
wire n_1521;
wire n_1694;
wire n_1940;
wire n_284;
wire n_593;
wire n_1695;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_1774;
wire n_409;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_2007;
wire n_526;
wire n_1994;
wire n_1767;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1973;
wire n_1444;
wire n_1803;
wire n_820;
wire n_1749;
wire n_872;
wire n_1653;
wire n_254;
wire n_1157;
wire n_1584;
wire n_234;
wire n_848;
wire n_1664;
wire n_280;
wire n_629;
wire n_1739;
wire n_1814;
wire n_532;
wire n_1789;
wire n_763;
wire n_1986;
wire n_540;
wire n_216;
wire n_692;
wire n_2054;
wire n_1857;
wire n_984;
wire n_1687;
wire n_2073;
wire n_223;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_2046;
wire n_1816;
wire n_1910;
wire n_1756;
wire n_1606;
wire n_395;
wire n_621;
wire n_1587;
wire n_213;
wire n_2093;
wire n_2018;
wire n_1772;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_2040;
wire n_493;
wire n_1311;
wire n_1956;
wire n_1589;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_697;
wire n_622;
wire n_1626;
wire n_1962;
wire n_1335;
wire n_1715;
wire n_296;
wire n_880;
wire n_793;
wire n_2114;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_1785;
wire n_792;
wire n_1262;
wire n_1942;
wire n_580;
wire n_1579;
wire n_494;
wire n_434;
wire n_2014;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1893;
wire n_1183;
wire n_1326;
wire n_1805;
wire n_981;
wire n_1110;
wire n_1758;
wire n_243;
wire n_1407;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_2010;
wire n_1054;
wire n_508;
wire n_1679;
wire n_1952;
wire n_1858;
wire n_353;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_1834;
wire n_1011;
wire n_978;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_1721;
wire n_653;
wire n_1445;
wire n_1317;
wire n_2050;
wire n_783;
wire n_556;
wire n_1127;
wire n_1536;
wire n_1471;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_1980;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_1998;
wire n_541;
wire n_499;
wire n_1775;
wire n_788;
wire n_908;
wire n_1036;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_2028;
wire n_919;
wire n_1663;
wire n_2092;
wire n_1625;
wire n_2086;
wire n_1926;
wire n_318;
wire n_1458;
wire n_244;
wire n_679;
wire n_1630;
wire n_220;
wire n_663;
wire n_1720;
wire n_443;
wire n_1412;
wire n_1738;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_1922;
wire n_1735;
wire n_1788;
wire n_391;
wire n_940;
wire n_1537;
wire n_2065;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_1930;
wire n_765;
wire n_1809;
wire n_1843;
wire n_1904;
wire n_2000;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_2096;
wire n_1530;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_898;
wire n_857;
wire n_363;
wire n_1067;
wire n_968;
wire n_1235;
wire n_1323;
wire n_1462;
wire n_2012;
wire n_1937;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_2039;
wire n_1755;
wire n_1285;
wire n_761;
wire n_733;
wire n_731;
wire n_336;
wire n_1813;
wire n_315;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_2111;
wire n_1996;
wire n_1106;
wire n_2009;
wire n_648;
wire n_784;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_2024;
wire n_1348;
wire n_753;
wire n_1770;
wire n_701;
wire n_1003;
wire n_1125;
wire n_2103;
wire n_1710;
wire n_1865;
wire n_309;
wire n_1344;
wire n_1390;
wire n_401;
wire n_485;
wire n_1792;
wire n_504;
wire n_2062;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_291;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1510;
wire n_1099;
wire n_839;
wire n_1754;
wire n_759;
wire n_567;
wire n_240;
wire n_369;
wire n_1727;
wire n_1991;
wire n_1575;
wire n_1848;
wire n_1892;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_323;
wire n_550;
wire n_1315;
wire n_1660;
wire n_1902;
wire n_997;
wire n_635;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_248;
wire n_1152;
wire n_2034;
wire n_1845;
wire n_1934;
wire n_2101;
wire n_921;
wire n_1615;
wire n_1236;
wire n_228;
wire n_2104;
wire n_1265;
wire n_1576;
wire n_2105;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1806;
wire n_1409;
wire n_1148;
wire n_1684;
wire n_1588;
wire n_1673;
wire n_1334;
wire n_654;
wire n_2088;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_2005;
wire n_2048;
wire n_1696;
wire n_498;
wire n_1875;
wire n_1059;
wire n_684;
wire n_2108;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1831;
wire n_1497;
wire n_1866;
wire n_2056;
wire n_459;
wire n_1136;
wire n_1782;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_838;
wire n_383;
wire n_1558;
wire n_1941;
wire n_1316;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_1915;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_1781;
wire n_709;
wire n_809;
wire n_2085;
wire n_1686;
wire n_1964;
wire n_235;
wire n_881;
wire n_1019;
wire n_1477;
wire n_1777;
wire n_1982;
wire n_2097;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_217;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_708;
wire n_308;
wire n_1223;
wire n_1768;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1983;
wire n_1041;
wire n_2115;
wire n_993;
wire n_1862;
wire n_948;
wire n_2017;
wire n_922;
wire n_1004;
wire n_1810;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_1923;
wire n_1764;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_1337;
wire n_774;
wire n_1946;
wire n_933;
wire n_1779;
wire n_596;
wire n_954;
wire n_2051;
wire n_1168;
wire n_1821;
wire n_219;
wire n_1310;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_252;
wire n_664;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_1896;
wire n_1732;
wire n_415;
wire n_1967;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_2052;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1724;
wire n_1670;
wire n_1707;
wire n_1799;
wire n_2080;
wire n_2058;
wire n_1126;
wire n_2029;
wire n_1846;
wire n_1912;
wire n_938;
wire n_1891;
wire n_1328;
wire n_895;
wire n_304;
wire n_1639;
wire n_583;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_1928;
wire n_946;
wire n_757;
wire n_2047;
wire n_375;
wire n_1655;
wire n_1818;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_472;
wire n_937;
wire n_1474;
wire n_2081;
wire n_265;
wire n_1583;
wire n_1604;
wire n_208;
wire n_1631;
wire n_1702;
wire n_275;
wire n_1794;
wire n_1375;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_496;
wire n_1827;
wire n_866;
wire n_246;
wire n_925;
wire n_1752;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_1129;
wire n_1252;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_1871;
wire n_329;
wire n_718;
wire n_1434;
wire n_340;
wire n_1905;
wire n_1569;
wire n_548;
wire n_289;
wire n_523;
wire n_1662;
wire n_457;
wire n_1299;
wire n_1870;
wire n_2063;
wire n_1925;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1861;
wire n_2079;
wire n_1228;
wire n_1931;
wire n_1244;
wire n_1796;
wire n_411;
wire n_484;
wire n_849;
wire n_2095;
wire n_1820;
wire n_357;
wire n_412;
wire n_1251;
wire n_1989;
wire n_447;
wire n_1421;
wire n_1762;
wire n_1233;
wire n_1808;
wire n_1574;
wire n_1672;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_1981;
wire n_2037;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_2089;
wire n_1487;
wire n_675;

BUFx10_ASAP7_75t_L g205 ( 
.A(n_36),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_45),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_67),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_61),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_24),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_188),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_87),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_25),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_119),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_166),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_33),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_140),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_60),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_40),
.Y(n_218)
);

BUFx2_ASAP7_75t_L g219 ( 
.A(n_186),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_163),
.Y(n_220)
);

HB1xp67_ASAP7_75t_L g221 ( 
.A(n_66),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_152),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_192),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_167),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_68),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_133),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_23),
.Y(n_227)
);

CKINVDCx16_ASAP7_75t_R g228 ( 
.A(n_31),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_193),
.Y(n_229)
);

INVx1_ASAP7_75t_SL g230 ( 
.A(n_29),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_195),
.Y(n_231)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_122),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_43),
.Y(n_233)
);

CKINVDCx16_ASAP7_75t_R g234 ( 
.A(n_41),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_2),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_61),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_107),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_79),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_124),
.Y(n_239)
);

BUFx3_ASAP7_75t_L g240 ( 
.A(n_58),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_39),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_178),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_132),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_157),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_96),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_191),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_118),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_71),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_103),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_33),
.Y(n_250)
);

BUFx3_ASAP7_75t_L g251 ( 
.A(n_104),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_204),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_16),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_100),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_187),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_137),
.Y(n_256)
);

INVxp67_ASAP7_75t_SL g257 ( 
.A(n_161),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_128),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_37),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_169),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_171),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_183),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_149),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_69),
.Y(n_264)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_82),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_185),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_44),
.Y(n_267)
);

CKINVDCx16_ASAP7_75t_R g268 ( 
.A(n_83),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_46),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_45),
.Y(n_270)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_111),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_184),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_30),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_6),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_139),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_32),
.Y(n_276)
);

BUFx6f_ASAP7_75t_L g277 ( 
.A(n_141),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_115),
.Y(n_278)
);

CKINVDCx16_ASAP7_75t_R g279 ( 
.A(n_92),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_42),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_14),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_73),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_190),
.Y(n_283)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_198),
.Y(n_284)
);

INVx1_ASAP7_75t_SL g285 ( 
.A(n_32),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_131),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_26),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_41),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_196),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_42),
.Y(n_290)
);

INVx2_ASAP7_75t_L g291 ( 
.A(n_75),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_75),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_176),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_199),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_159),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_5),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_43),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_76),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_136),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_180),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_39),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_181),
.Y(n_302)
);

INVx2_ASAP7_75t_L g303 ( 
.A(n_123),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_13),
.Y(n_304)
);

BUFx3_ASAP7_75t_L g305 ( 
.A(n_86),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g306 ( 
.A(n_135),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_168),
.Y(n_307)
);

BUFx10_ASAP7_75t_L g308 ( 
.A(n_162),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_71),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_63),
.Y(n_310)
);

BUFx2_ASAP7_75t_L g311 ( 
.A(n_114),
.Y(n_311)
);

BUFx10_ASAP7_75t_L g312 ( 
.A(n_34),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_35),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_194),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_37),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_47),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_30),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_101),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_138),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_155),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_72),
.Y(n_321)
);

INVx2_ASAP7_75t_L g322 ( 
.A(n_81),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g323 ( 
.A(n_94),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_27),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_203),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_1),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_51),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_179),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_27),
.Y(n_329)
);

INVx2_ASAP7_75t_L g330 ( 
.A(n_134),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_154),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_44),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_95),
.Y(n_333)
);

INVx2_ASAP7_75t_SL g334 ( 
.A(n_12),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_19),
.Y(n_335)
);

BUFx5_ASAP7_75t_L g336 ( 
.A(n_52),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_150),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_127),
.Y(n_338)
);

BUFx3_ASAP7_75t_L g339 ( 
.A(n_102),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_10),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_18),
.Y(n_341)
);

CKINVDCx16_ASAP7_75t_R g342 ( 
.A(n_91),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_130),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_197),
.Y(n_344)
);

INVx2_ASAP7_75t_SL g345 ( 
.A(n_54),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_36),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_108),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_170),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_19),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_49),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_174),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_54),
.Y(n_352)
);

CKINVDCx20_ASAP7_75t_R g353 ( 
.A(n_15),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_17),
.Y(n_354)
);

CKINVDCx20_ASAP7_75t_R g355 ( 
.A(n_144),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_89),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_125),
.Y(n_357)
);

CKINVDCx20_ASAP7_75t_R g358 ( 
.A(n_34),
.Y(n_358)
);

CKINVDCx20_ASAP7_75t_R g359 ( 
.A(n_25),
.Y(n_359)
);

CKINVDCx20_ASAP7_75t_R g360 ( 
.A(n_67),
.Y(n_360)
);

BUFx6f_ASAP7_75t_L g361 ( 
.A(n_189),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_151),
.Y(n_362)
);

BUFx10_ASAP7_75t_L g363 ( 
.A(n_2),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_200),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_76),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_49),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_53),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_60),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_120),
.Y(n_369)
);

CKINVDCx20_ASAP7_75t_R g370 ( 
.A(n_110),
.Y(n_370)
);

BUFx6f_ASAP7_75t_L g371 ( 
.A(n_7),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_97),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_77),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_143),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_16),
.Y(n_375)
);

CKINVDCx16_ASAP7_75t_R g376 ( 
.A(n_17),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_175),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_23),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_126),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_202),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_56),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_22),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_172),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_6),
.Y(n_384)
);

INVx2_ASAP7_75t_L g385 ( 
.A(n_77),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_173),
.Y(n_386)
);

CKINVDCx14_ASAP7_75t_R g387 ( 
.A(n_160),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_112),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_56),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_55),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_51),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_58),
.Y(n_392)
);

INVxp67_ASAP7_75t_SL g393 ( 
.A(n_11),
.Y(n_393)
);

BUFx6f_ASAP7_75t_L g394 ( 
.A(n_148),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_50),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_22),
.Y(n_396)
);

BUFx3_ASAP7_75t_L g397 ( 
.A(n_121),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_85),
.Y(n_398)
);

BUFx3_ASAP7_75t_L g399 ( 
.A(n_73),
.Y(n_399)
);

CKINVDCx20_ASAP7_75t_R g400 ( 
.A(n_5),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_78),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_12),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_106),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_145),
.Y(n_404)
);

BUFx2_ASAP7_75t_L g405 ( 
.A(n_113),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_74),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_31),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_336),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_336),
.Y(n_409)
);

BUFx2_ASAP7_75t_L g410 ( 
.A(n_221),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_336),
.Y(n_411)
);

BUFx2_ASAP7_75t_L g412 ( 
.A(n_240),
.Y(n_412)
);

CKINVDCx16_ASAP7_75t_R g413 ( 
.A(n_228),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_336),
.Y(n_414)
);

INVx2_ASAP7_75t_L g415 ( 
.A(n_336),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_336),
.Y(n_416)
);

CKINVDCx20_ASAP7_75t_R g417 ( 
.A(n_220),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_336),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_336),
.Y(n_419)
);

INVx2_ASAP7_75t_L g420 ( 
.A(n_371),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_371),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_371),
.Y(n_422)
);

INVxp67_ASAP7_75t_L g423 ( 
.A(n_334),
.Y(n_423)
);

INVxp67_ASAP7_75t_L g424 ( 
.A(n_334),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_371),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_371),
.Y(n_426)
);

HB1xp67_ASAP7_75t_L g427 ( 
.A(n_234),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_291),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_291),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_385),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_385),
.Y(n_431)
);

INVx2_ASAP7_75t_L g432 ( 
.A(n_251),
.Y(n_432)
);

INVx2_ASAP7_75t_L g433 ( 
.A(n_251),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_376),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_232),
.Y(n_435)
);

CKINVDCx5p33_ASAP7_75t_R g436 ( 
.A(n_263),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_232),
.Y(n_437)
);

CKINVDCx16_ASAP7_75t_R g438 ( 
.A(n_268),
.Y(n_438)
);

HB1xp67_ASAP7_75t_L g439 ( 
.A(n_208),
.Y(n_439)
);

CKINVDCx5p33_ASAP7_75t_R g440 ( 
.A(n_306),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_265),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_265),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_271),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_271),
.Y(n_444)
);

INVxp67_ASAP7_75t_SL g445 ( 
.A(n_240),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_284),
.Y(n_446)
);

HB1xp67_ASAP7_75t_L g447 ( 
.A(n_208),
.Y(n_447)
);

CKINVDCx20_ASAP7_75t_R g448 ( 
.A(n_323),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_284),
.Y(n_449)
);

INVxp33_ASAP7_75t_SL g450 ( 
.A(n_407),
.Y(n_450)
);

HB1xp67_ASAP7_75t_L g451 ( 
.A(n_209),
.Y(n_451)
);

CKINVDCx5p33_ASAP7_75t_R g452 ( 
.A(n_355),
.Y(n_452)
);

CKINVDCx16_ASAP7_75t_R g453 ( 
.A(n_279),
.Y(n_453)
);

CKINVDCx20_ASAP7_75t_R g454 ( 
.A(n_370),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_303),
.Y(n_455)
);

CKINVDCx20_ASAP7_75t_R g456 ( 
.A(n_225),
.Y(n_456)
);

BUFx3_ASAP7_75t_L g457 ( 
.A(n_305),
.Y(n_457)
);

CKINVDCx16_ASAP7_75t_R g458 ( 
.A(n_342),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_303),
.Y(n_459)
);

CKINVDCx16_ASAP7_75t_R g460 ( 
.A(n_387),
.Y(n_460)
);

INVxp67_ASAP7_75t_SL g461 ( 
.A(n_399),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_322),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_322),
.Y(n_463)
);

CKINVDCx20_ASAP7_75t_R g464 ( 
.A(n_233),
.Y(n_464)
);

CKINVDCx5p33_ASAP7_75t_R g465 ( 
.A(n_264),
.Y(n_465)
);

INVxp67_ASAP7_75t_SL g466 ( 
.A(n_399),
.Y(n_466)
);

INVxp67_ASAP7_75t_SL g467 ( 
.A(n_206),
.Y(n_467)
);

CKINVDCx5p33_ASAP7_75t_R g468 ( 
.A(n_267),
.Y(n_468)
);

CKINVDCx16_ASAP7_75t_R g469 ( 
.A(n_205),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_330),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_330),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_207),
.Y(n_472)
);

CKINVDCx20_ASAP7_75t_R g473 ( 
.A(n_241),
.Y(n_473)
);

CKINVDCx5p33_ASAP7_75t_R g474 ( 
.A(n_270),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_215),
.Y(n_475)
);

INVx2_ASAP7_75t_L g476 ( 
.A(n_305),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_217),
.Y(n_477)
);

CKINVDCx5p33_ASAP7_75t_R g478 ( 
.A(n_273),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_218),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_253),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_259),
.Y(n_481)
);

CKINVDCx5p33_ASAP7_75t_R g482 ( 
.A(n_274),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_280),
.Y(n_483)
);

INVxp33_ASAP7_75t_SL g484 ( 
.A(n_209),
.Y(n_484)
);

INVxp67_ASAP7_75t_L g485 ( 
.A(n_345),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_281),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_282),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_288),
.Y(n_488)
);

CKINVDCx5p33_ASAP7_75t_R g489 ( 
.A(n_276),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_297),
.Y(n_490)
);

CKINVDCx20_ASAP7_75t_R g491 ( 
.A(n_269),
.Y(n_491)
);

CKINVDCx20_ASAP7_75t_R g492 ( 
.A(n_353),
.Y(n_492)
);

CKINVDCx16_ASAP7_75t_R g493 ( 
.A(n_205),
.Y(n_493)
);

CKINVDCx20_ASAP7_75t_R g494 ( 
.A(n_358),
.Y(n_494)
);

INVx2_ASAP7_75t_L g495 ( 
.A(n_339),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_298),
.Y(n_496)
);

CKINVDCx5p33_ASAP7_75t_R g497 ( 
.A(n_287),
.Y(n_497)
);

INVxp33_ASAP7_75t_L g498 ( 
.A(n_304),
.Y(n_498)
);

CKINVDCx5p33_ASAP7_75t_R g499 ( 
.A(n_290),
.Y(n_499)
);

CKINVDCx20_ASAP7_75t_R g500 ( 
.A(n_359),
.Y(n_500)
);

CKINVDCx5p33_ASAP7_75t_R g501 ( 
.A(n_292),
.Y(n_501)
);

INVxp33_ASAP7_75t_L g502 ( 
.A(n_309),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_321),
.Y(n_503)
);

HB1xp67_ASAP7_75t_L g504 ( 
.A(n_212),
.Y(n_504)
);

INVxp33_ASAP7_75t_SL g505 ( 
.A(n_212),
.Y(n_505)
);

CKINVDCx5p33_ASAP7_75t_R g506 ( 
.A(n_301),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_349),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_350),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_352),
.Y(n_509)
);

INVxp33_ASAP7_75t_SL g510 ( 
.A(n_407),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_365),
.Y(n_511)
);

CKINVDCx5p33_ASAP7_75t_R g512 ( 
.A(n_310),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_366),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_368),
.Y(n_514)
);

INVxp33_ASAP7_75t_SL g515 ( 
.A(n_227),
.Y(n_515)
);

AND2x4_ASAP7_75t_L g516 ( 
.A(n_457),
.B(n_219),
.Y(n_516)
);

INVx2_ASAP7_75t_L g517 ( 
.A(n_420),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_408),
.Y(n_518)
);

BUFx6f_ASAP7_75t_L g519 ( 
.A(n_420),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_408),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_409),
.Y(n_521)
);

CKINVDCx5p33_ASAP7_75t_R g522 ( 
.A(n_436),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_L g523 ( 
.A(n_445),
.B(n_311),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_409),
.Y(n_524)
);

CKINVDCx5p33_ASAP7_75t_R g525 ( 
.A(n_440),
.Y(n_525)
);

CKINVDCx5p33_ASAP7_75t_R g526 ( 
.A(n_452),
.Y(n_526)
);

BUFx6f_ASAP7_75t_L g527 ( 
.A(n_415),
.Y(n_527)
);

CKINVDCx5p33_ASAP7_75t_R g528 ( 
.A(n_417),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_411),
.Y(n_529)
);

INVxp67_ASAP7_75t_L g530 ( 
.A(n_427),
.Y(n_530)
);

BUFx6f_ASAP7_75t_L g531 ( 
.A(n_415),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_L g532 ( 
.A(n_461),
.B(n_405),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_L g533 ( 
.A(n_466),
.B(n_211),
.Y(n_533)
);

INVx2_ASAP7_75t_L g534 ( 
.A(n_411),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_L g535 ( 
.A(n_457),
.B(n_213),
.Y(n_535)
);

CKINVDCx6p67_ASAP7_75t_R g536 ( 
.A(n_460),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_414),
.Y(n_537)
);

AND2x4_ASAP7_75t_L g538 ( 
.A(n_432),
.B(n_339),
.Y(n_538)
);

NAND2xp33_ASAP7_75t_R g539 ( 
.A(n_434),
.B(n_227),
.Y(n_539)
);

INVx2_ASAP7_75t_L g540 ( 
.A(n_414),
.Y(n_540)
);

INVx2_ASAP7_75t_L g541 ( 
.A(n_421),
.Y(n_541)
);

AND2x2_ASAP7_75t_L g542 ( 
.A(n_412),
.B(n_205),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_416),
.Y(n_543)
);

OAI22xp5_ASAP7_75t_SL g544 ( 
.A1(n_456),
.A2(n_400),
.B1(n_360),
.B2(n_235),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_416),
.Y(n_545)
);

BUFx6f_ASAP7_75t_L g546 ( 
.A(n_421),
.Y(n_546)
);

AND2x2_ASAP7_75t_L g547 ( 
.A(n_412),
.B(n_312),
.Y(n_547)
);

BUFx3_ASAP7_75t_L g548 ( 
.A(n_432),
.Y(n_548)
);

HB1xp67_ASAP7_75t_L g549 ( 
.A(n_413),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_418),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_L g551 ( 
.A(n_460),
.B(n_224),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_418),
.Y(n_552)
);

INVx2_ASAP7_75t_L g553 ( 
.A(n_419),
.Y(n_553)
);

AND2x2_ASAP7_75t_L g554 ( 
.A(n_498),
.B(n_312),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_419),
.Y(n_555)
);

AND2x4_ASAP7_75t_L g556 ( 
.A(n_433),
.B(n_397),
.Y(n_556)
);

NOR2xp33_ASAP7_75t_L g557 ( 
.A(n_450),
.B(n_484),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_L g558 ( 
.A(n_433),
.B(n_226),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_422),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_L g560 ( 
.A(n_476),
.B(n_231),
.Y(n_560)
);

INVxp67_ASAP7_75t_L g561 ( 
.A(n_439),
.Y(n_561)
);

BUFx6f_ASAP7_75t_L g562 ( 
.A(n_422),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_425),
.Y(n_563)
);

OAI22xp5_ASAP7_75t_L g564 ( 
.A1(n_438),
.A2(n_230),
.B1(n_285),
.B2(n_401),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_425),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_L g566 ( 
.A(n_476),
.B(n_238),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_426),
.Y(n_567)
);

CKINVDCx20_ASAP7_75t_R g568 ( 
.A(n_464),
.Y(n_568)
);

CKINVDCx5p33_ASAP7_75t_R g569 ( 
.A(n_448),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_426),
.Y(n_570)
);

HB1xp67_ASAP7_75t_L g571 ( 
.A(n_465),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_435),
.Y(n_572)
);

BUFx2_ASAP7_75t_L g573 ( 
.A(n_468),
.Y(n_573)
);

NOR2xp33_ASAP7_75t_L g574 ( 
.A(n_505),
.B(n_244),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_435),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_L g576 ( 
.A(n_495),
.B(n_247),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_437),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_437),
.Y(n_578)
);

INVx2_ASAP7_75t_L g579 ( 
.A(n_441),
.Y(n_579)
);

AND2x4_ASAP7_75t_L g580 ( 
.A(n_495),
.B(n_397),
.Y(n_580)
);

AND2x2_ASAP7_75t_L g581 ( 
.A(n_502),
.B(n_312),
.Y(n_581)
);

BUFx6f_ASAP7_75t_L g582 ( 
.A(n_441),
.Y(n_582)
);

CKINVDCx5p33_ASAP7_75t_R g583 ( 
.A(n_454),
.Y(n_583)
);

XNOR2xp5_ASAP7_75t_L g584 ( 
.A(n_473),
.B(n_235),
.Y(n_584)
);

INVx2_ASAP7_75t_L g585 ( 
.A(n_442),
.Y(n_585)
);

OAI22xp5_ASAP7_75t_SL g586 ( 
.A1(n_491),
.A2(n_332),
.B1(n_236),
.B2(n_248),
.Y(n_586)
);

OA21x2_ASAP7_75t_L g587 ( 
.A1(n_442),
.A2(n_252),
.B(n_249),
.Y(n_587)
);

INVx2_ASAP7_75t_SL g588 ( 
.A(n_474),
.Y(n_588)
);

BUFx2_ASAP7_75t_L g589 ( 
.A(n_478),
.Y(n_589)
);

BUFx3_ASAP7_75t_L g590 ( 
.A(n_443),
.Y(n_590)
);

NOR2xp33_ASAP7_75t_R g591 ( 
.A(n_482),
.B(n_261),
.Y(n_591)
);

INVx4_ASAP7_75t_L g592 ( 
.A(n_443),
.Y(n_592)
);

CKINVDCx5p33_ASAP7_75t_R g593 ( 
.A(n_489),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_444),
.Y(n_594)
);

INVx2_ASAP7_75t_L g595 ( 
.A(n_444),
.Y(n_595)
);

HB1xp67_ASAP7_75t_L g596 ( 
.A(n_497),
.Y(n_596)
);

NAND2xp33_ASAP7_75t_R g597 ( 
.A(n_499),
.B(n_236),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_446),
.Y(n_598)
);

CKINVDCx5p33_ASAP7_75t_R g599 ( 
.A(n_501),
.Y(n_599)
);

INVx3_ASAP7_75t_L g600 ( 
.A(n_446),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_534),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_534),
.Y(n_602)
);

INVx2_ASAP7_75t_L g603 ( 
.A(n_534),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_L g604 ( 
.A(n_574),
.B(n_438),
.Y(n_604)
);

INVx2_ASAP7_75t_SL g605 ( 
.A(n_554),
.Y(n_605)
);

NAND2xp33_ASAP7_75t_L g606 ( 
.A(n_588),
.B(n_506),
.Y(n_606)
);

INVx2_ASAP7_75t_L g607 ( 
.A(n_540),
.Y(n_607)
);

INVx2_ASAP7_75t_L g608 ( 
.A(n_540),
.Y(n_608)
);

AOI22xp33_ASAP7_75t_SL g609 ( 
.A1(n_586),
.A2(n_458),
.B1(n_453),
.B2(n_469),
.Y(n_609)
);

AOI21x1_ASAP7_75t_L g610 ( 
.A1(n_518),
.A2(n_455),
.B(n_449),
.Y(n_610)
);

OAI22xp5_ASAP7_75t_SL g611 ( 
.A1(n_544),
.A2(n_494),
.B1(n_500),
.B2(n_492),
.Y(n_611)
);

INVx2_ASAP7_75t_L g612 ( 
.A(n_540),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_L g613 ( 
.A(n_548),
.B(n_458),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_553),
.Y(n_614)
);

AOI22xp5_ASAP7_75t_L g615 ( 
.A1(n_586),
.A2(n_393),
.B1(n_250),
.B2(n_296),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_SL g616 ( 
.A(n_591),
.B(n_512),
.Y(n_616)
);

CKINVDCx5p33_ASAP7_75t_R g617 ( 
.A(n_593),
.Y(n_617)
);

INVx2_ASAP7_75t_L g618 ( 
.A(n_553),
.Y(n_618)
);

AND2x2_ASAP7_75t_L g619 ( 
.A(n_554),
.B(n_467),
.Y(n_619)
);

INVx2_ASAP7_75t_L g620 ( 
.A(n_553),
.Y(n_620)
);

INVx2_ASAP7_75t_L g621 ( 
.A(n_518),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_559),
.Y(n_622)
);

NOR2xp33_ASAP7_75t_L g623 ( 
.A(n_551),
.B(n_510),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_559),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_563),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_L g626 ( 
.A(n_548),
.B(n_455),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_563),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_L g628 ( 
.A(n_516),
.B(n_459),
.Y(n_628)
);

INVx2_ASAP7_75t_L g629 ( 
.A(n_520),
.Y(n_629)
);

OAI22xp5_ASAP7_75t_L g630 ( 
.A1(n_557),
.A2(n_515),
.B1(n_250),
.B2(n_296),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_SL g631 ( 
.A(n_588),
.B(n_599),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_SL g632 ( 
.A(n_573),
.B(n_493),
.Y(n_632)
);

OR2x2_ASAP7_75t_L g633 ( 
.A(n_581),
.B(n_410),
.Y(n_633)
);

AOI22xp5_ASAP7_75t_L g634 ( 
.A1(n_564),
.A2(n_597),
.B1(n_581),
.B2(n_547),
.Y(n_634)
);

CKINVDCx5p33_ASAP7_75t_R g635 ( 
.A(n_522),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_565),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_SL g637 ( 
.A(n_573),
.B(n_447),
.Y(n_637)
);

AOI22xp5_ASAP7_75t_SL g638 ( 
.A1(n_584),
.A2(n_410),
.B1(n_424),
.B2(n_423),
.Y(n_638)
);

AOI22xp33_ASAP7_75t_SL g639 ( 
.A1(n_544),
.A2(n_363),
.B1(n_504),
.B2(n_451),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_565),
.Y(n_640)
);

INVx2_ASAP7_75t_L g641 ( 
.A(n_520),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_L g642 ( 
.A(n_516),
.B(n_459),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_567),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_567),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_L g645 ( 
.A(n_516),
.B(n_462),
.Y(n_645)
);

INVx2_ASAP7_75t_L g646 ( 
.A(n_521),
.Y(n_646)
);

NAND3xp33_ASAP7_75t_SL g647 ( 
.A(n_589),
.B(n_316),
.C(n_248),
.Y(n_647)
);

AND2x2_ASAP7_75t_L g648 ( 
.A(n_590),
.B(n_472),
.Y(n_648)
);

BUFx4f_ASAP7_75t_L g649 ( 
.A(n_587),
.Y(n_649)
);

INVx1_ASAP7_75t_SL g650 ( 
.A(n_568),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_L g651 ( 
.A(n_516),
.B(n_462),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_SL g652 ( 
.A(n_589),
.B(n_210),
.Y(n_652)
);

INVx8_ASAP7_75t_L g653 ( 
.A(n_538),
.Y(n_653)
);

INVx2_ASAP7_75t_SL g654 ( 
.A(n_542),
.Y(n_654)
);

INVx2_ASAP7_75t_L g655 ( 
.A(n_521),
.Y(n_655)
);

INVx4_ASAP7_75t_L g656 ( 
.A(n_527),
.Y(n_656)
);

INVx1_ASAP7_75t_SL g657 ( 
.A(n_528),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_SL g658 ( 
.A(n_542),
.B(n_210),
.Y(n_658)
);

INVx2_ASAP7_75t_L g659 ( 
.A(n_524),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_570),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_570),
.Y(n_661)
);

INVx3_ASAP7_75t_L g662 ( 
.A(n_527),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_524),
.Y(n_663)
);

OAI22xp5_ASAP7_75t_SL g664 ( 
.A1(n_584),
.A2(n_317),
.B1(n_324),
.B2(n_316),
.Y(n_664)
);

OAI22xp5_ASAP7_75t_SL g665 ( 
.A1(n_569),
.A2(n_324),
.B1(n_326),
.B2(n_317),
.Y(n_665)
);

NAND3xp33_ASAP7_75t_L g666 ( 
.A(n_529),
.B(n_470),
.C(n_463),
.Y(n_666)
);

INVx2_ASAP7_75t_L g667 ( 
.A(n_529),
.Y(n_667)
);

BUFx2_ASAP7_75t_L g668 ( 
.A(n_530),
.Y(n_668)
);

NAND2xp33_ASAP7_75t_R g669 ( 
.A(n_525),
.B(n_475),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_L g670 ( 
.A(n_537),
.B(n_463),
.Y(n_670)
);

HB1xp67_ASAP7_75t_L g671 ( 
.A(n_549),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_537),
.Y(n_672)
);

INVx2_ASAP7_75t_SL g673 ( 
.A(n_547),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_543),
.Y(n_674)
);

INVx2_ASAP7_75t_L g675 ( 
.A(n_543),
.Y(n_675)
);

INVxp33_ASAP7_75t_SL g676 ( 
.A(n_526),
.Y(n_676)
);

NAND2xp33_ASAP7_75t_L g677 ( 
.A(n_571),
.B(n_214),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_SL g678 ( 
.A(n_523),
.B(n_214),
.Y(n_678)
);

BUFx2_ASAP7_75t_L g679 ( 
.A(n_561),
.Y(n_679)
);

AND2x2_ASAP7_75t_SL g680 ( 
.A(n_587),
.B(n_277),
.Y(n_680)
);

BUFx3_ASAP7_75t_L g681 ( 
.A(n_545),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_L g682 ( 
.A(n_550),
.B(n_470),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_550),
.Y(n_683)
);

INVx2_ASAP7_75t_L g684 ( 
.A(n_552),
.Y(n_684)
);

BUFx6f_ASAP7_75t_L g685 ( 
.A(n_527),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_552),
.Y(n_686)
);

CKINVDCx5p33_ASAP7_75t_R g687 ( 
.A(n_583),
.Y(n_687)
);

INVx2_ASAP7_75t_L g688 ( 
.A(n_555),
.Y(n_688)
);

INVx2_ASAP7_75t_L g689 ( 
.A(n_527),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_582),
.Y(n_690)
);

BUFx6f_ASAP7_75t_L g691 ( 
.A(n_527),
.Y(n_691)
);

AOI21x1_ASAP7_75t_L g692 ( 
.A1(n_587),
.A2(n_471),
.B(n_255),
.Y(n_692)
);

AOI22xp5_ASAP7_75t_L g693 ( 
.A1(n_539),
.A2(n_367),
.B1(n_326),
.B2(n_354),
.Y(n_693)
);

INVx2_ASAP7_75t_L g694 ( 
.A(n_527),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_582),
.Y(n_695)
);

INVx3_ASAP7_75t_L g696 ( 
.A(n_531),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_SL g697 ( 
.A(n_532),
.B(n_216),
.Y(n_697)
);

AO21x2_ASAP7_75t_L g698 ( 
.A1(n_533),
.A2(n_258),
.B(n_254),
.Y(n_698)
);

INVx2_ASAP7_75t_L g699 ( 
.A(n_531),
.Y(n_699)
);

INVx2_ASAP7_75t_L g700 ( 
.A(n_531),
.Y(n_700)
);

INVx2_ASAP7_75t_L g701 ( 
.A(n_531),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_582),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_582),
.Y(n_703)
);

BUFx10_ASAP7_75t_L g704 ( 
.A(n_596),
.Y(n_704)
);

INVx2_ASAP7_75t_L g705 ( 
.A(n_531),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_SL g706 ( 
.A(n_592),
.B(n_216),
.Y(n_706)
);

INVx2_ASAP7_75t_L g707 ( 
.A(n_531),
.Y(n_707)
);

CKINVDCx20_ASAP7_75t_R g708 ( 
.A(n_536),
.Y(n_708)
);

NOR2xp33_ASAP7_75t_SL g709 ( 
.A(n_536),
.B(n_308),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_582),
.Y(n_710)
);

AO21x2_ASAP7_75t_L g711 ( 
.A1(n_535),
.A2(n_278),
.B(n_260),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_582),
.Y(n_712)
);

INVx2_ASAP7_75t_L g713 ( 
.A(n_541),
.Y(n_713)
);

INVx2_ASAP7_75t_L g714 ( 
.A(n_541),
.Y(n_714)
);

AND2x2_ASAP7_75t_L g715 ( 
.A(n_590),
.B(n_475),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_579),
.Y(n_716)
);

INVx2_ASAP7_75t_L g717 ( 
.A(n_517),
.Y(n_717)
);

INVx2_ASAP7_75t_L g718 ( 
.A(n_517),
.Y(n_718)
);

INVx2_ASAP7_75t_L g719 ( 
.A(n_546),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_579),
.Y(n_720)
);

NAND2xp33_ASAP7_75t_SL g721 ( 
.A(n_592),
.B(n_327),
.Y(n_721)
);

INVx2_ASAP7_75t_L g722 ( 
.A(n_546),
.Y(n_722)
);

INVx3_ASAP7_75t_L g723 ( 
.A(n_546),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_579),
.Y(n_724)
);

INVx3_ASAP7_75t_L g725 ( 
.A(n_546),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_585),
.Y(n_726)
);

INVx2_ASAP7_75t_L g727 ( 
.A(n_546),
.Y(n_727)
);

INVx3_ASAP7_75t_L g728 ( 
.A(n_546),
.Y(n_728)
);

INVxp67_ASAP7_75t_L g729 ( 
.A(n_558),
.Y(n_729)
);

INVx2_ASAP7_75t_L g730 ( 
.A(n_562),
.Y(n_730)
);

AND2x2_ASAP7_75t_L g731 ( 
.A(n_592),
.B(n_477),
.Y(n_731)
);

INVx2_ASAP7_75t_L g732 ( 
.A(n_562),
.Y(n_732)
);

INVx2_ASAP7_75t_L g733 ( 
.A(n_562),
.Y(n_733)
);

BUFx2_ASAP7_75t_L g734 ( 
.A(n_538),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_L g735 ( 
.A(n_538),
.B(n_479),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_585),
.Y(n_736)
);

INVx4_ASAP7_75t_L g737 ( 
.A(n_587),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_585),
.Y(n_738)
);

INVx2_ASAP7_75t_L g739 ( 
.A(n_562),
.Y(n_739)
);

INVx2_ASAP7_75t_L g740 ( 
.A(n_562),
.Y(n_740)
);

INVx2_ASAP7_75t_L g741 ( 
.A(n_562),
.Y(n_741)
);

INVxp67_ASAP7_75t_L g742 ( 
.A(n_560),
.Y(n_742)
);

BUFx6f_ASAP7_75t_SL g743 ( 
.A(n_556),
.Y(n_743)
);

NAND3xp33_ASAP7_75t_L g744 ( 
.A(n_572),
.B(n_378),
.C(n_375),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_SL g745 ( 
.A(n_556),
.B(n_222),
.Y(n_745)
);

INVx2_ASAP7_75t_L g746 ( 
.A(n_519),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_SL g747 ( 
.A(n_681),
.B(n_600),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_L g748 ( 
.A(n_729),
.B(n_556),
.Y(n_748)
);

INVx2_ASAP7_75t_L g749 ( 
.A(n_603),
.Y(n_749)
);

NOR2xp33_ASAP7_75t_L g750 ( 
.A(n_623),
.B(n_566),
.Y(n_750)
);

AOI22xp5_ASAP7_75t_L g751 ( 
.A1(n_605),
.A2(n_257),
.B1(n_600),
.B2(n_575),
.Y(n_751)
);

INVx2_ASAP7_75t_L g752 ( 
.A(n_603),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_SL g753 ( 
.A(n_681),
.B(n_600),
.Y(n_753)
);

INVx2_ASAP7_75t_L g754 ( 
.A(n_603),
.Y(n_754)
);

NOR2xp33_ASAP7_75t_L g755 ( 
.A(n_605),
.B(n_576),
.Y(n_755)
);

INVx2_ASAP7_75t_L g756 ( 
.A(n_655),
.Y(n_756)
);

BUFx6f_ASAP7_75t_L g757 ( 
.A(n_685),
.Y(n_757)
);

CKINVDCx5p33_ASAP7_75t_R g758 ( 
.A(n_617),
.Y(n_758)
);

INVx2_ASAP7_75t_SL g759 ( 
.A(n_668),
.Y(n_759)
);

BUFx3_ASAP7_75t_L g760 ( 
.A(n_653),
.Y(n_760)
);

INVxp67_ASAP7_75t_L g761 ( 
.A(n_668),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_L g762 ( 
.A(n_742),
.B(n_556),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_L g763 ( 
.A(n_619),
.B(n_580),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_L g764 ( 
.A(n_731),
.B(n_580),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_622),
.Y(n_765)
);

AOI22xp5_ASAP7_75t_L g766 ( 
.A1(n_654),
.A2(n_572),
.B1(n_594),
.B2(n_578),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_SL g767 ( 
.A(n_681),
.B(n_222),
.Y(n_767)
);

INVxp33_ASAP7_75t_L g768 ( 
.A(n_679),
.Y(n_768)
);

BUFx6f_ASAP7_75t_L g769 ( 
.A(n_685),
.Y(n_769)
);

NAND2xp33_ASAP7_75t_L g770 ( 
.A(n_655),
.B(n_223),
.Y(n_770)
);

OR2x2_ASAP7_75t_L g771 ( 
.A(n_633),
.B(n_485),
.Y(n_771)
);

INVx2_ASAP7_75t_L g772 ( 
.A(n_607),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_L g773 ( 
.A(n_648),
.B(n_577),
.Y(n_773)
);

INVxp67_ASAP7_75t_L g774 ( 
.A(n_679),
.Y(n_774)
);

INVx2_ASAP7_75t_L g775 ( 
.A(n_607),
.Y(n_775)
);

BUFx6f_ASAP7_75t_L g776 ( 
.A(n_685),
.Y(n_776)
);

INVx2_ASAP7_75t_L g777 ( 
.A(n_607),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_L g778 ( 
.A(n_648),
.B(n_577),
.Y(n_778)
);

INVx2_ASAP7_75t_SL g779 ( 
.A(n_671),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_SL g780 ( 
.A(n_663),
.B(n_223),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_SL g781 ( 
.A(n_663),
.B(n_229),
.Y(n_781)
);

BUFx6f_ASAP7_75t_L g782 ( 
.A(n_685),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_L g783 ( 
.A(n_715),
.B(n_578),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_L g784 ( 
.A(n_715),
.B(n_594),
.Y(n_784)
);

NAND2xp33_ASAP7_75t_L g785 ( 
.A(n_655),
.B(n_229),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_L g786 ( 
.A(n_654),
.B(n_598),
.Y(n_786)
);

AOI22xp5_ASAP7_75t_L g787 ( 
.A1(n_673),
.A2(n_295),
.B1(n_404),
.B2(n_403),
.Y(n_787)
);

NOR3xp33_ASAP7_75t_L g788 ( 
.A(n_665),
.B(n_604),
.C(n_630),
.Y(n_788)
);

INVx2_ASAP7_75t_L g789 ( 
.A(n_659),
.Y(n_789)
);

INVx2_ASAP7_75t_SL g790 ( 
.A(n_704),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_SL g791 ( 
.A(n_672),
.B(n_237),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_L g792 ( 
.A(n_673),
.B(n_595),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_L g793 ( 
.A(n_628),
.B(n_595),
.Y(n_793)
);

NOR2xp33_ASAP7_75t_L g794 ( 
.A(n_613),
.B(n_595),
.Y(n_794)
);

OAI22xp33_ASAP7_75t_L g795 ( 
.A1(n_615),
.A2(n_384),
.B1(n_389),
.B2(n_395),
.Y(n_795)
);

NOR2xp33_ASAP7_75t_L g796 ( 
.A(n_658),
.B(n_313),
.Y(n_796)
);

INVx2_ASAP7_75t_L g797 ( 
.A(n_659),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_SL g798 ( 
.A(n_672),
.B(n_237),
.Y(n_798)
);

NAND2x1p5_ASAP7_75t_L g799 ( 
.A(n_734),
.B(n_283),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_L g800 ( 
.A(n_642),
.B(n_239),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_L g801 ( 
.A(n_645),
.B(n_239),
.Y(n_801)
);

OR2x2_ASAP7_75t_L g802 ( 
.A(n_633),
.B(n_650),
.Y(n_802)
);

AND2x4_ASAP7_75t_L g803 ( 
.A(n_734),
.B(n_479),
.Y(n_803)
);

AND2x2_ASAP7_75t_L g804 ( 
.A(n_638),
.B(n_480),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_L g805 ( 
.A(n_651),
.B(n_242),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_SL g806 ( 
.A(n_674),
.B(n_242),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_624),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_625),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_SL g809 ( 
.A(n_674),
.B(n_243),
.Y(n_809)
);

INVx4_ASAP7_75t_L g810 ( 
.A(n_653),
.Y(n_810)
);

NOR2xp33_ASAP7_75t_L g811 ( 
.A(n_634),
.B(n_315),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_625),
.Y(n_812)
);

INVxp67_ASAP7_75t_L g813 ( 
.A(n_669),
.Y(n_813)
);

NOR2xp33_ASAP7_75t_L g814 ( 
.A(n_634),
.B(n_381),
.Y(n_814)
);

NAND2xp33_ASAP7_75t_L g815 ( 
.A(n_659),
.B(n_667),
.Y(n_815)
);

NAND2xp33_ASAP7_75t_SL g816 ( 
.A(n_635),
.B(n_327),
.Y(n_816)
);

INVx2_ASAP7_75t_L g817 ( 
.A(n_667),
.Y(n_817)
);

NAND2xp33_ASAP7_75t_L g818 ( 
.A(n_667),
.B(n_243),
.Y(n_818)
);

INVx3_ASAP7_75t_L g819 ( 
.A(n_653),
.Y(n_819)
);

INVx2_ASAP7_75t_L g820 ( 
.A(n_608),
.Y(n_820)
);

INVx1_ASAP7_75t_L g821 ( 
.A(n_627),
.Y(n_821)
);

AND2x6_ASAP7_75t_SL g822 ( 
.A(n_676),
.B(n_396),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_627),
.Y(n_823)
);

AOI22xp33_ASAP7_75t_L g824 ( 
.A1(n_664),
.A2(n_406),
.B1(n_308),
.B2(n_363),
.Y(n_824)
);

NOR2xp33_ASAP7_75t_L g825 ( 
.A(n_678),
.B(n_382),
.Y(n_825)
);

OAI22xp5_ASAP7_75t_L g826 ( 
.A1(n_683),
.A2(n_373),
.B1(n_367),
.B2(n_340),
.Y(n_826)
);

AOI21xp5_ASAP7_75t_L g827 ( 
.A1(n_683),
.A2(n_294),
.B(n_289),
.Y(n_827)
);

NOR2xp67_ASAP7_75t_SL g828 ( 
.A(n_616),
.B(n_329),
.Y(n_828)
);

NOR2xp33_ASAP7_75t_L g829 ( 
.A(n_697),
.B(n_390),
.Y(n_829)
);

AND2x2_ASAP7_75t_L g830 ( 
.A(n_638),
.B(n_480),
.Y(n_830)
);

OR2x6_ASAP7_75t_L g831 ( 
.A(n_653),
.B(n_611),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_636),
.Y(n_832)
);

INVx2_ASAP7_75t_L g833 ( 
.A(n_608),
.Y(n_833)
);

NOR2xp33_ASAP7_75t_L g834 ( 
.A(n_745),
.B(n_329),
.Y(n_834)
);

BUFx6f_ASAP7_75t_SL g835 ( 
.A(n_704),
.Y(n_835)
);

INVx2_ASAP7_75t_L g836 ( 
.A(n_608),
.Y(n_836)
);

O2A1O1Ixp33_ASAP7_75t_L g837 ( 
.A1(n_686),
.A2(n_486),
.B(n_514),
.C(n_513),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_SL g838 ( 
.A(n_685),
.B(n_245),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_L g839 ( 
.A(n_735),
.B(n_245),
.Y(n_839)
);

AOI22xp5_ASAP7_75t_L g840 ( 
.A1(n_677),
.A2(n_295),
.B1(n_256),
.B2(n_246),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_L g841 ( 
.A(n_698),
.B(n_246),
.Y(n_841)
);

NOR2xp33_ASAP7_75t_L g842 ( 
.A(n_652),
.B(n_332),
.Y(n_842)
);

INVx2_ASAP7_75t_L g843 ( 
.A(n_612),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_SL g844 ( 
.A(n_685),
.B(n_256),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_SL g845 ( 
.A(n_691),
.B(n_649),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_L g846 ( 
.A(n_698),
.B(n_320),
.Y(n_846)
);

INVx2_ASAP7_75t_L g847 ( 
.A(n_612),
.Y(n_847)
);

NAND2xp33_ASAP7_75t_L g848 ( 
.A(n_621),
.B(n_320),
.Y(n_848)
);

INVx2_ASAP7_75t_L g849 ( 
.A(n_612),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_636),
.Y(n_850)
);

NOR2xp33_ASAP7_75t_L g851 ( 
.A(n_706),
.B(n_335),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_L g852 ( 
.A(n_698),
.B(n_325),
.Y(n_852)
);

NAND2xp33_ASAP7_75t_SL g853 ( 
.A(n_631),
.B(n_335),
.Y(n_853)
);

OR2x6_ASAP7_75t_L g854 ( 
.A(n_653),
.B(n_481),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_640),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_640),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_L g857 ( 
.A(n_621),
.B(n_325),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_L g858 ( 
.A(n_629),
.B(n_328),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_643),
.Y(n_859)
);

NAND3xp33_ASAP7_75t_L g860 ( 
.A(n_693),
.B(n_341),
.C(n_340),
.Y(n_860)
);

INVxp67_ASAP7_75t_L g861 ( 
.A(n_657),
.Y(n_861)
);

AND2x2_ASAP7_75t_L g862 ( 
.A(n_704),
.B(n_483),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_L g863 ( 
.A(n_641),
.B(n_331),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_643),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_L g865 ( 
.A(n_646),
.B(n_333),
.Y(n_865)
);

A2O1A1Ixp33_ASAP7_75t_L g866 ( 
.A1(n_615),
.A2(n_486),
.B(n_514),
.C(n_513),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_L g867 ( 
.A(n_646),
.B(n_333),
.Y(n_867)
);

INVx3_ASAP7_75t_L g868 ( 
.A(n_610),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_L g869 ( 
.A(n_675),
.B(n_338),
.Y(n_869)
);

NAND3xp33_ASAP7_75t_L g870 ( 
.A(n_606),
.B(n_346),
.C(n_341),
.Y(n_870)
);

INVx4_ASAP7_75t_L g871 ( 
.A(n_743),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_SL g872 ( 
.A(n_691),
.B(n_344),
.Y(n_872)
);

INVx1_ASAP7_75t_L g873 ( 
.A(n_644),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_644),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_L g875 ( 
.A(n_684),
.B(n_344),
.Y(n_875)
);

AND2x2_ASAP7_75t_SL g876 ( 
.A(n_709),
.B(n_314),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_660),
.Y(n_877)
);

NOR2xp33_ASAP7_75t_L g878 ( 
.A(n_743),
.B(n_346),
.Y(n_878)
);

INVx2_ASAP7_75t_L g879 ( 
.A(n_618),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_660),
.Y(n_880)
);

BUFx6f_ASAP7_75t_SL g881 ( 
.A(n_704),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_L g882 ( 
.A(n_684),
.B(n_351),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_661),
.Y(n_883)
);

CKINVDCx5p33_ASAP7_75t_R g884 ( 
.A(n_687),
.Y(n_884)
);

NOR2xp33_ASAP7_75t_SL g885 ( 
.A(n_708),
.B(n_308),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_L g886 ( 
.A(n_688),
.B(n_351),
.Y(n_886)
);

INVx2_ASAP7_75t_L g887 ( 
.A(n_618),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_SL g888 ( 
.A(n_691),
.B(n_357),
.Y(n_888)
);

INVx2_ASAP7_75t_L g889 ( 
.A(n_618),
.Y(n_889)
);

OR2x2_ASAP7_75t_L g890 ( 
.A(n_632),
.B(n_483),
.Y(n_890)
);

INVx2_ASAP7_75t_SL g891 ( 
.A(n_637),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_SL g892 ( 
.A(n_691),
.B(n_357),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_L g893 ( 
.A(n_688),
.B(n_369),
.Y(n_893)
);

NOR2xp67_ASAP7_75t_L g894 ( 
.A(n_647),
.B(n_487),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_SL g895 ( 
.A(n_691),
.B(n_369),
.Y(n_895)
);

INVx1_ASAP7_75t_L g896 ( 
.A(n_661),
.Y(n_896)
);

INVx8_ASAP7_75t_L g897 ( 
.A(n_743),
.Y(n_897)
);

BUFx2_ASAP7_75t_L g898 ( 
.A(n_665),
.Y(n_898)
);

NAND2xp5_ASAP7_75t_L g899 ( 
.A(n_601),
.B(n_372),
.Y(n_899)
);

OR2x2_ASAP7_75t_L g900 ( 
.A(n_664),
.B(n_487),
.Y(n_900)
);

AO221x1_ASAP7_75t_L g901 ( 
.A1(n_611),
.A2(n_277),
.B1(n_361),
.B2(n_394),
.C(n_343),
.Y(n_901)
);

CKINVDCx6p67_ASAP7_75t_R g902 ( 
.A(n_743),
.Y(n_902)
);

AND2x4_ASAP7_75t_L g903 ( 
.A(n_810),
.B(n_716),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_SL g904 ( 
.A(n_810),
.B(n_691),
.Y(n_904)
);

INVxp67_ASAP7_75t_L g905 ( 
.A(n_759),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_765),
.Y(n_906)
);

INVx2_ASAP7_75t_L g907 ( 
.A(n_749),
.Y(n_907)
);

BUFx3_ASAP7_75t_L g908 ( 
.A(n_897),
.Y(n_908)
);

NOR2xp33_ASAP7_75t_L g909 ( 
.A(n_750),
.B(n_721),
.Y(n_909)
);

INVx2_ASAP7_75t_L g910 ( 
.A(n_749),
.Y(n_910)
);

NAND2xp5_ASAP7_75t_L g911 ( 
.A(n_750),
.B(n_601),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_L g912 ( 
.A(n_755),
.B(n_602),
.Y(n_912)
);

BUFx2_ASAP7_75t_L g913 ( 
.A(n_761),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_L g914 ( 
.A(n_755),
.B(n_602),
.Y(n_914)
);

AND2x6_ASAP7_75t_SL g915 ( 
.A(n_811),
.B(n_488),
.Y(n_915)
);

AND2x4_ASAP7_75t_L g916 ( 
.A(n_760),
.B(n_716),
.Y(n_916)
);

NOR3xp33_ASAP7_75t_SL g917 ( 
.A(n_758),
.B(n_373),
.C(n_354),
.Y(n_917)
);

INVx2_ASAP7_75t_L g918 ( 
.A(n_752),
.Y(n_918)
);

NAND2xp5_ASAP7_75t_SL g919 ( 
.A(n_819),
.B(n_656),
.Y(n_919)
);

INVx3_ASAP7_75t_L g920 ( 
.A(n_760),
.Y(n_920)
);

AOI21xp5_ASAP7_75t_L g921 ( 
.A1(n_815),
.A2(n_696),
.B(n_662),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_L g922 ( 
.A(n_763),
.B(n_614),
.Y(n_922)
);

NAND2xp5_ASAP7_75t_SL g923 ( 
.A(n_819),
.B(n_656),
.Y(n_923)
);

HB1xp67_ASAP7_75t_L g924 ( 
.A(n_774),
.Y(n_924)
);

BUFx6f_ASAP7_75t_L g925 ( 
.A(n_897),
.Y(n_925)
);

INVx2_ASAP7_75t_L g926 ( 
.A(n_752),
.Y(n_926)
);

AND2x6_ASAP7_75t_SL g927 ( 
.A(n_811),
.B(n_488),
.Y(n_927)
);

AOI21xp33_ASAP7_75t_L g928 ( 
.A1(n_814),
.A2(n_609),
.B(n_649),
.Y(n_928)
);

AND2x2_ASAP7_75t_L g929 ( 
.A(n_804),
.B(n_639),
.Y(n_929)
);

INVx3_ASAP7_75t_L g930 ( 
.A(n_871),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_807),
.Y(n_931)
);

INVx1_ASAP7_75t_L g932 ( 
.A(n_808),
.Y(n_932)
);

INVx1_ASAP7_75t_L g933 ( 
.A(n_812),
.Y(n_933)
);

NOR2xp33_ASAP7_75t_R g934 ( 
.A(n_884),
.B(n_649),
.Y(n_934)
);

BUFx6f_ASAP7_75t_L g935 ( 
.A(n_897),
.Y(n_935)
);

NOR3xp33_ASAP7_75t_SL g936 ( 
.A(n_816),
.B(n_392),
.C(n_391),
.Y(n_936)
);

INVx1_ASAP7_75t_L g937 ( 
.A(n_821),
.Y(n_937)
);

AND2x2_ASAP7_75t_L g938 ( 
.A(n_830),
.B(n_490),
.Y(n_938)
);

NOR2xp33_ASAP7_75t_L g939 ( 
.A(n_813),
.B(n_656),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_L g940 ( 
.A(n_794),
.B(n_720),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_L g941 ( 
.A(n_862),
.B(n_720),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_SL g942 ( 
.A(n_757),
.B(n_656),
.Y(n_942)
);

INVx1_ASAP7_75t_L g943 ( 
.A(n_823),
.Y(n_943)
);

AND2x2_ASAP7_75t_L g944 ( 
.A(n_768),
.B(n_771),
.Y(n_944)
);

INVx2_ASAP7_75t_L g945 ( 
.A(n_754),
.Y(n_945)
);

INVx1_ASAP7_75t_L g946 ( 
.A(n_832),
.Y(n_946)
);

AND2x4_ASAP7_75t_L g947 ( 
.A(n_871),
.B(n_724),
.Y(n_947)
);

BUFx3_ASAP7_75t_L g948 ( 
.A(n_902),
.Y(n_948)
);

INVx1_ASAP7_75t_L g949 ( 
.A(n_850),
.Y(n_949)
);

NOR2xp33_ASAP7_75t_SL g950 ( 
.A(n_876),
.B(n_744),
.Y(n_950)
);

CKINVDCx11_ASAP7_75t_R g951 ( 
.A(n_822),
.Y(n_951)
);

NAND2xp5_ASAP7_75t_L g952 ( 
.A(n_803),
.B(n_724),
.Y(n_952)
);

INVx2_ASAP7_75t_L g953 ( 
.A(n_754),
.Y(n_953)
);

AND2x4_ASAP7_75t_L g954 ( 
.A(n_854),
.B(n_726),
.Y(n_954)
);

NOR3xp33_ASAP7_75t_SL g955 ( 
.A(n_853),
.B(n_392),
.C(n_391),
.Y(n_955)
);

INVx3_ASAP7_75t_L g956 ( 
.A(n_757),
.Y(n_956)
);

INVx2_ASAP7_75t_L g957 ( 
.A(n_772),
.Y(n_957)
);

INVx1_ASAP7_75t_L g958 ( 
.A(n_855),
.Y(n_958)
);

NOR3xp33_ASAP7_75t_L g959 ( 
.A(n_898),
.B(n_402),
.C(n_401),
.Y(n_959)
);

NAND2xp5_ASAP7_75t_SL g960 ( 
.A(n_757),
.B(n_662),
.Y(n_960)
);

AND2x4_ASAP7_75t_L g961 ( 
.A(n_854),
.B(n_736),
.Y(n_961)
);

BUFx6f_ASAP7_75t_L g962 ( 
.A(n_769),
.Y(n_962)
);

INVx4_ASAP7_75t_L g963 ( 
.A(n_854),
.Y(n_963)
);

NOR2xp33_ASAP7_75t_L g964 ( 
.A(n_814),
.B(n_662),
.Y(n_964)
);

INVx2_ASAP7_75t_L g965 ( 
.A(n_772),
.Y(n_965)
);

INVx1_ASAP7_75t_L g966 ( 
.A(n_856),
.Y(n_966)
);

NAND2xp5_ASAP7_75t_SL g967 ( 
.A(n_769),
.B(n_662),
.Y(n_967)
);

INVx1_ASAP7_75t_L g968 ( 
.A(n_859),
.Y(n_968)
);

NAND2x1p5_ASAP7_75t_L g969 ( 
.A(n_864),
.B(n_696),
.Y(n_969)
);

AOI22xp33_ASAP7_75t_L g970 ( 
.A1(n_900),
.A2(n_795),
.B1(n_824),
.B2(n_788),
.Y(n_970)
);

HB1xp67_ASAP7_75t_L g971 ( 
.A(n_779),
.Y(n_971)
);

INVx2_ASAP7_75t_L g972 ( 
.A(n_775),
.Y(n_972)
);

INVx1_ASAP7_75t_L g973 ( 
.A(n_873),
.Y(n_973)
);

AND2x2_ASAP7_75t_L g974 ( 
.A(n_802),
.B(n_490),
.Y(n_974)
);

AOI22xp5_ASAP7_75t_L g975 ( 
.A1(n_876),
.A2(n_738),
.B1(n_710),
.B2(n_703),
.Y(n_975)
);

NOR3xp33_ASAP7_75t_SL g976 ( 
.A(n_870),
.B(n_402),
.C(n_744),
.Y(n_976)
);

NAND2xp5_ASAP7_75t_L g977 ( 
.A(n_748),
.B(n_738),
.Y(n_977)
);

INVx2_ASAP7_75t_L g978 ( 
.A(n_775),
.Y(n_978)
);

BUFx3_ASAP7_75t_L g979 ( 
.A(n_769),
.Y(n_979)
);

INVx1_ASAP7_75t_L g980 ( 
.A(n_874),
.Y(n_980)
);

INVx1_ASAP7_75t_L g981 ( 
.A(n_877),
.Y(n_981)
);

AOI22xp33_ASAP7_75t_L g982 ( 
.A1(n_795),
.A2(n_711),
.B1(n_680),
.B2(n_737),
.Y(n_982)
);

INVx1_ASAP7_75t_L g983 ( 
.A(n_880),
.Y(n_983)
);

NAND2xp5_ASAP7_75t_SL g984 ( 
.A(n_776),
.B(n_696),
.Y(n_984)
);

NAND2xp5_ASAP7_75t_SL g985 ( 
.A(n_776),
.B(n_620),
.Y(n_985)
);

INVx1_ASAP7_75t_L g986 ( 
.A(n_883),
.Y(n_986)
);

NOR2xp33_ASAP7_75t_L g987 ( 
.A(n_762),
.B(n_737),
.Y(n_987)
);

NAND2xp5_ASAP7_75t_SL g988 ( 
.A(n_776),
.B(n_782),
.Y(n_988)
);

AND2x4_ASAP7_75t_L g989 ( 
.A(n_831),
.B(n_737),
.Y(n_989)
);

INVx1_ASAP7_75t_L g990 ( 
.A(n_896),
.Y(n_990)
);

AO22x1_ASAP7_75t_L g991 ( 
.A1(n_861),
.A2(n_503),
.B1(n_511),
.B2(n_509),
.Y(n_991)
);

NAND2xp5_ASAP7_75t_L g992 ( 
.A(n_764),
.B(n_626),
.Y(n_992)
);

NAND2xp5_ASAP7_75t_L g993 ( 
.A(n_786),
.B(n_620),
.Y(n_993)
);

BUFx6f_ASAP7_75t_L g994 ( 
.A(n_782),
.Y(n_994)
);

AOI22xp5_ASAP7_75t_L g995 ( 
.A1(n_851),
.A2(n_842),
.B1(n_878),
.B2(n_829),
.Y(n_995)
);

INVx1_ASAP7_75t_L g996 ( 
.A(n_792),
.Y(n_996)
);

NAND2xp5_ASAP7_75t_SL g997 ( 
.A(n_782),
.B(n_723),
.Y(n_997)
);

AND2x6_ASAP7_75t_L g998 ( 
.A(n_782),
.B(n_701),
.Y(n_998)
);

HB1xp67_ASAP7_75t_L g999 ( 
.A(n_799),
.Y(n_999)
);

NAND2xp5_ASAP7_75t_SL g1000 ( 
.A(n_756),
.B(n_723),
.Y(n_1000)
);

BUFx3_ASAP7_75t_L g1001 ( 
.A(n_799),
.Y(n_1001)
);

INVx2_ASAP7_75t_SL g1002 ( 
.A(n_890),
.Y(n_1002)
);

INVx1_ASAP7_75t_L g1003 ( 
.A(n_773),
.Y(n_1003)
);

AND2x2_ASAP7_75t_L g1004 ( 
.A(n_891),
.B(n_496),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_L g1005 ( 
.A(n_778),
.B(n_711),
.Y(n_1005)
);

NOR3xp33_ASAP7_75t_SL g1006 ( 
.A(n_826),
.B(n_398),
.C(n_372),
.Y(n_1006)
);

CKINVDCx5p33_ASAP7_75t_R g1007 ( 
.A(n_835),
.Y(n_1007)
);

INVx1_ASAP7_75t_L g1008 ( 
.A(n_783),
.Y(n_1008)
);

INVx1_ASAP7_75t_L g1009 ( 
.A(n_784),
.Y(n_1009)
);

INVx5_ASAP7_75t_L g1010 ( 
.A(n_868),
.Y(n_1010)
);

INVxp67_ASAP7_75t_L g1011 ( 
.A(n_894),
.Y(n_1011)
);

NAND2xp5_ASAP7_75t_L g1012 ( 
.A(n_766),
.B(n_711),
.Y(n_1012)
);

INVxp67_ASAP7_75t_L g1013 ( 
.A(n_885),
.Y(n_1013)
);

HB1xp67_ASAP7_75t_L g1014 ( 
.A(n_831),
.Y(n_1014)
);

AOI22xp33_ASAP7_75t_L g1015 ( 
.A1(n_824),
.A2(n_680),
.B1(n_737),
.B2(n_666),
.Y(n_1015)
);

HB1xp67_ASAP7_75t_L g1016 ( 
.A(n_831),
.Y(n_1016)
);

OR2x2_ASAP7_75t_L g1017 ( 
.A(n_860),
.B(n_670),
.Y(n_1017)
);

NOR2xp33_ASAP7_75t_L g1018 ( 
.A(n_842),
.B(n_701),
.Y(n_1018)
);

NAND2xp5_ASAP7_75t_SL g1019 ( 
.A(n_789),
.B(n_723),
.Y(n_1019)
);

OR2x2_ASAP7_75t_L g1020 ( 
.A(n_787),
.B(n_682),
.Y(n_1020)
);

NAND2xp5_ASAP7_75t_SL g1021 ( 
.A(n_797),
.B(n_723),
.Y(n_1021)
);

BUFx2_ASAP7_75t_L g1022 ( 
.A(n_790),
.Y(n_1022)
);

BUFx3_ASAP7_75t_L g1023 ( 
.A(n_817),
.Y(n_1023)
);

NOR2xp33_ASAP7_75t_L g1024 ( 
.A(n_780),
.B(n_781),
.Y(n_1024)
);

INVx5_ASAP7_75t_L g1025 ( 
.A(n_868),
.Y(n_1025)
);

AOI22xp5_ASAP7_75t_L g1026 ( 
.A1(n_851),
.A2(n_690),
.B1(n_695),
.B2(n_702),
.Y(n_1026)
);

INVx3_ASAP7_75t_L g1027 ( 
.A(n_777),
.Y(n_1027)
);

NOR2xp33_ASAP7_75t_R g1028 ( 
.A(n_835),
.B(n_610),
.Y(n_1028)
);

NAND2xp5_ASAP7_75t_L g1029 ( 
.A(n_878),
.B(n_680),
.Y(n_1029)
);

INVx2_ASAP7_75t_L g1030 ( 
.A(n_777),
.Y(n_1030)
);

CKINVDCx5p33_ASAP7_75t_R g1031 ( 
.A(n_881),
.Y(n_1031)
);

NOR3xp33_ASAP7_75t_SL g1032 ( 
.A(n_780),
.B(n_403),
.C(n_398),
.Y(n_1032)
);

NAND2xp5_ASAP7_75t_SL g1033 ( 
.A(n_845),
.B(n_725),
.Y(n_1033)
);

NAND2xp5_ASAP7_75t_L g1034 ( 
.A(n_866),
.B(n_713),
.Y(n_1034)
);

INVx1_ASAP7_75t_L g1035 ( 
.A(n_833),
.Y(n_1035)
);

INVx3_ASAP7_75t_L g1036 ( 
.A(n_833),
.Y(n_1036)
);

INVx2_ASAP7_75t_L g1037 ( 
.A(n_836),
.Y(n_1037)
);

NAND2xp5_ASAP7_75t_L g1038 ( 
.A(n_866),
.B(n_713),
.Y(n_1038)
);

NAND2x1p5_ASAP7_75t_L g1039 ( 
.A(n_747),
.B(n_725),
.Y(n_1039)
);

INVx1_ASAP7_75t_L g1040 ( 
.A(n_836),
.Y(n_1040)
);

BUFx6f_ASAP7_75t_L g1041 ( 
.A(n_843),
.Y(n_1041)
);

AOI22xp5_ASAP7_75t_L g1042 ( 
.A1(n_825),
.A2(n_690),
.B1(n_695),
.B2(n_702),
.Y(n_1042)
);

INVxp67_ASAP7_75t_L g1043 ( 
.A(n_834),
.Y(n_1043)
);

HB1xp67_ASAP7_75t_L g1044 ( 
.A(n_881),
.Y(n_1044)
);

AOI22xp33_ASAP7_75t_L g1045 ( 
.A1(n_901),
.A2(n_666),
.B1(n_714),
.B2(n_718),
.Y(n_1045)
);

INVx1_ASAP7_75t_L g1046 ( 
.A(n_843),
.Y(n_1046)
);

INVx2_ASAP7_75t_L g1047 ( 
.A(n_847),
.Y(n_1047)
);

O2A1O1Ixp33_ASAP7_75t_L g1048 ( 
.A1(n_747),
.A2(n_703),
.B(n_710),
.C(n_712),
.Y(n_1048)
);

NAND2x1p5_ASAP7_75t_L g1049 ( 
.A(n_753),
.B(n_725),
.Y(n_1049)
);

INVx1_ASAP7_75t_L g1050 ( 
.A(n_847),
.Y(n_1050)
);

OAI22xp5_ASAP7_75t_L g1051 ( 
.A1(n_753),
.A2(n_728),
.B1(n_712),
.B2(n_701),
.Y(n_1051)
);

BUFx3_ASAP7_75t_L g1052 ( 
.A(n_849),
.Y(n_1052)
);

AOI22xp5_ASAP7_75t_L g1053 ( 
.A1(n_825),
.A2(n_728),
.B1(n_700),
.B2(n_699),
.Y(n_1053)
);

XNOR2xp5_ASAP7_75t_L g1054 ( 
.A(n_840),
.B(n_692),
.Y(n_1054)
);

CKINVDCx5p33_ASAP7_75t_R g1055 ( 
.A(n_796),
.Y(n_1055)
);

NAND2xp5_ASAP7_75t_L g1056 ( 
.A(n_800),
.B(n_717),
.Y(n_1056)
);

INVx2_ASAP7_75t_SL g1057 ( 
.A(n_781),
.Y(n_1057)
);

INVx1_ASAP7_75t_SL g1058 ( 
.A(n_767),
.Y(n_1058)
);

INVx2_ASAP7_75t_L g1059 ( 
.A(n_849),
.Y(n_1059)
);

INVx5_ASAP7_75t_L g1060 ( 
.A(n_820),
.Y(n_1060)
);

INVx2_ASAP7_75t_L g1061 ( 
.A(n_879),
.Y(n_1061)
);

NAND2xp5_ASAP7_75t_SL g1062 ( 
.A(n_751),
.B(n_728),
.Y(n_1062)
);

INVx2_ASAP7_75t_L g1063 ( 
.A(n_887),
.Y(n_1063)
);

BUFx3_ASAP7_75t_L g1064 ( 
.A(n_889),
.Y(n_1064)
);

INVx2_ASAP7_75t_L g1065 ( 
.A(n_793),
.Y(n_1065)
);

INVx5_ASAP7_75t_L g1066 ( 
.A(n_828),
.Y(n_1066)
);

NAND2xp5_ASAP7_75t_SL g1067 ( 
.A(n_767),
.B(n_727),
.Y(n_1067)
);

BUFx2_ASAP7_75t_L g1068 ( 
.A(n_857),
.Y(n_1068)
);

NAND2xp5_ASAP7_75t_L g1069 ( 
.A(n_801),
.B(n_717),
.Y(n_1069)
);

AND2x2_ASAP7_75t_L g1070 ( 
.A(n_796),
.B(n_496),
.Y(n_1070)
);

NOR2x2_ASAP7_75t_L g1071 ( 
.A(n_834),
.B(n_727),
.Y(n_1071)
);

INVx2_ASAP7_75t_L g1072 ( 
.A(n_899),
.Y(n_1072)
);

INVx4_ASAP7_75t_L g1073 ( 
.A(n_770),
.Y(n_1073)
);

NOR2xp33_ASAP7_75t_L g1074 ( 
.A(n_791),
.B(n_689),
.Y(n_1074)
);

NAND2xp5_ASAP7_75t_L g1075 ( 
.A(n_805),
.B(n_718),
.Y(n_1075)
);

AND2x2_ASAP7_75t_SL g1076 ( 
.A(n_841),
.B(n_318),
.Y(n_1076)
);

NOR2xp33_ASAP7_75t_L g1077 ( 
.A(n_791),
.B(n_689),
.Y(n_1077)
);

NOR3xp33_ASAP7_75t_SL g1078 ( 
.A(n_798),
.B(n_404),
.C(n_509),
.Y(n_1078)
);

INVx1_ASAP7_75t_L g1079 ( 
.A(n_837),
.Y(n_1079)
);

NAND3xp33_ASAP7_75t_L g1080 ( 
.A(n_995),
.B(n_848),
.C(n_818),
.Y(n_1080)
);

NOR2xp33_ASAP7_75t_R g1081 ( 
.A(n_1007),
.B(n_785),
.Y(n_1081)
);

AOI21xp5_ASAP7_75t_L g1082 ( 
.A1(n_911),
.A2(n_844),
.B(n_838),
.Y(n_1082)
);

INVx1_ASAP7_75t_SL g1083 ( 
.A(n_913),
.Y(n_1083)
);

NOR2x1_ASAP7_75t_L g1084 ( 
.A(n_948),
.B(n_798),
.Y(n_1084)
);

NAND2x1p5_ASAP7_75t_L g1085 ( 
.A(n_925),
.B(n_806),
.Y(n_1085)
);

CKINVDCx5p33_ASAP7_75t_R g1086 ( 
.A(n_1031),
.Y(n_1086)
);

AOI21xp5_ASAP7_75t_L g1087 ( 
.A1(n_940),
.A2(n_888),
.B(n_872),
.Y(n_1087)
);

INVx1_ASAP7_75t_L g1088 ( 
.A(n_906),
.Y(n_1088)
);

NOR2xp33_ASAP7_75t_SL g1089 ( 
.A(n_1055),
.B(n_846),
.Y(n_1089)
);

O2A1O1Ixp33_ASAP7_75t_L g1090 ( 
.A1(n_909),
.A2(n_809),
.B(n_806),
.C(n_839),
.Y(n_1090)
);

BUFx12f_ASAP7_75t_L g1091 ( 
.A(n_951),
.Y(n_1091)
);

INVx2_ASAP7_75t_L g1092 ( 
.A(n_907),
.Y(n_1092)
);

NAND2xp5_ASAP7_75t_L g1093 ( 
.A(n_938),
.B(n_809),
.Y(n_1093)
);

NAND2xp5_ASAP7_75t_L g1094 ( 
.A(n_1003),
.B(n_858),
.Y(n_1094)
);

AOI22xp33_ASAP7_75t_L g1095 ( 
.A1(n_970),
.A2(n_852),
.B1(n_893),
.B2(n_867),
.Y(n_1095)
);

NAND2xp5_ASAP7_75t_L g1096 ( 
.A(n_1008),
.B(n_863),
.Y(n_1096)
);

AOI21xp5_ASAP7_75t_L g1097 ( 
.A1(n_912),
.A2(n_892),
.B(n_872),
.Y(n_1097)
);

BUFx3_ASAP7_75t_L g1098 ( 
.A(n_948),
.Y(n_1098)
);

AOI21xp5_ASAP7_75t_L g1099 ( 
.A1(n_914),
.A2(n_895),
.B(n_865),
.Y(n_1099)
);

AND2x2_ASAP7_75t_L g1100 ( 
.A(n_974),
.B(n_503),
.Y(n_1100)
);

O2A1O1Ixp33_ASAP7_75t_L g1101 ( 
.A1(n_1043),
.A2(n_886),
.B(n_882),
.C(n_875),
.Y(n_1101)
);

OR2x6_ASAP7_75t_L g1102 ( 
.A(n_963),
.B(n_827),
.Y(n_1102)
);

NAND2xp5_ASAP7_75t_L g1103 ( 
.A(n_1009),
.B(n_869),
.Y(n_1103)
);

BUFx2_ASAP7_75t_L g1104 ( 
.A(n_971),
.Y(n_1104)
);

NAND2xp5_ASAP7_75t_SL g1105 ( 
.A(n_964),
.B(n_1029),
.Y(n_1105)
);

NAND2xp5_ASAP7_75t_SL g1106 ( 
.A(n_964),
.B(n_694),
.Y(n_1106)
);

OAI21x1_ASAP7_75t_L g1107 ( 
.A1(n_921),
.A2(n_692),
.B(n_694),
.Y(n_1107)
);

AND2x2_ASAP7_75t_L g1108 ( 
.A(n_944),
.B(n_507),
.Y(n_1108)
);

CKINVDCx8_ASAP7_75t_R g1109 ( 
.A(n_915),
.Y(n_1109)
);

NOR2xp33_ASAP7_75t_L g1110 ( 
.A(n_970),
.B(n_705),
.Y(n_1110)
);

INVx2_ASAP7_75t_L g1111 ( 
.A(n_907),
.Y(n_1111)
);

A2O1A1Ixp33_ASAP7_75t_L g1112 ( 
.A1(n_1024),
.A2(n_928),
.B(n_1070),
.C(n_1018),
.Y(n_1112)
);

INVx1_ASAP7_75t_L g1113 ( 
.A(n_931),
.Y(n_1113)
);

AOI21xp5_ASAP7_75t_L g1114 ( 
.A1(n_987),
.A2(n_705),
.B(n_707),
.Y(n_1114)
);

O2A1O1Ixp33_ASAP7_75t_L g1115 ( 
.A1(n_1024),
.A2(n_511),
.B(n_507),
.C(n_508),
.Y(n_1115)
);

OAI21xp5_ASAP7_75t_L g1116 ( 
.A1(n_987),
.A2(n_707),
.B(n_741),
.Y(n_1116)
);

NAND2xp5_ASAP7_75t_SL g1117 ( 
.A(n_989),
.B(n_727),
.Y(n_1117)
);

BUFx2_ASAP7_75t_L g1118 ( 
.A(n_924),
.Y(n_1118)
);

INVx3_ASAP7_75t_L g1119 ( 
.A(n_925),
.Y(n_1119)
);

INVx1_ASAP7_75t_L g1120 ( 
.A(n_932),
.Y(n_1120)
);

INVx2_ASAP7_75t_L g1121 ( 
.A(n_910),
.Y(n_1121)
);

NAND2xp5_ASAP7_75t_SL g1122 ( 
.A(n_989),
.B(n_730),
.Y(n_1122)
);

HB1xp67_ASAP7_75t_L g1123 ( 
.A(n_954),
.Y(n_1123)
);

AO32x1_ASAP7_75t_L g1124 ( 
.A1(n_1054),
.A2(n_429),
.A3(n_428),
.B1(n_430),
.B2(n_431),
.Y(n_1124)
);

INVxp67_ASAP7_75t_SL g1125 ( 
.A(n_962),
.Y(n_1125)
);

OR2x2_ASAP7_75t_L g1126 ( 
.A(n_1002),
.B(n_508),
.Y(n_1126)
);

NAND2xp5_ASAP7_75t_SL g1127 ( 
.A(n_989),
.B(n_903),
.Y(n_1127)
);

AND2x4_ASAP7_75t_L g1128 ( 
.A(n_908),
.B(n_730),
.Y(n_1128)
);

INVx3_ASAP7_75t_L g1129 ( 
.A(n_925),
.Y(n_1129)
);

NOR2xp33_ASAP7_75t_L g1130 ( 
.A(n_927),
.B(n_719),
.Y(n_1130)
);

NAND2xp5_ASAP7_75t_SL g1131 ( 
.A(n_903),
.B(n_732),
.Y(n_1131)
);

INVx1_ASAP7_75t_L g1132 ( 
.A(n_933),
.Y(n_1132)
);

BUFx2_ASAP7_75t_L g1133 ( 
.A(n_905),
.Y(n_1133)
);

NAND2xp5_ASAP7_75t_L g1134 ( 
.A(n_1065),
.B(n_996),
.Y(n_1134)
);

OR2x6_ASAP7_75t_L g1135 ( 
.A(n_963),
.B(n_719),
.Y(n_1135)
);

NAND2xp5_ASAP7_75t_L g1136 ( 
.A(n_1004),
.B(n_952),
.Y(n_1136)
);

AND2x2_ASAP7_75t_L g1137 ( 
.A(n_929),
.B(n_363),
.Y(n_1137)
);

INVx4_ASAP7_75t_L g1138 ( 
.A(n_925),
.Y(n_1138)
);

NAND2xp5_ASAP7_75t_SL g1139 ( 
.A(n_903),
.B(n_732),
.Y(n_1139)
);

CKINVDCx14_ASAP7_75t_R g1140 ( 
.A(n_934),
.Y(n_1140)
);

BUFx8_ASAP7_75t_SL g1141 ( 
.A(n_1022),
.Y(n_1141)
);

CKINVDCx8_ASAP7_75t_R g1142 ( 
.A(n_935),
.Y(n_1142)
);

AOI21xp5_ASAP7_75t_L g1143 ( 
.A1(n_1033),
.A2(n_740),
.B(n_739),
.Y(n_1143)
);

AND2x2_ASAP7_75t_L g1144 ( 
.A(n_999),
.B(n_428),
.Y(n_1144)
);

A2O1A1Ixp33_ASAP7_75t_L g1145 ( 
.A1(n_1018),
.A2(n_356),
.B(n_364),
.C(n_362),
.Y(n_1145)
);

AND2x4_ASAP7_75t_L g1146 ( 
.A(n_908),
.B(n_733),
.Y(n_1146)
);

NAND2xp5_ASAP7_75t_L g1147 ( 
.A(n_1076),
.B(n_733),
.Y(n_1147)
);

INVxp67_ASAP7_75t_L g1148 ( 
.A(n_950),
.Y(n_1148)
);

NOR2xp33_ASAP7_75t_L g1149 ( 
.A(n_1058),
.B(n_722),
.Y(n_1149)
);

INVx1_ASAP7_75t_L g1150 ( 
.A(n_937),
.Y(n_1150)
);

INVx2_ASAP7_75t_SL g1151 ( 
.A(n_1044),
.Y(n_1151)
);

A2O1A1Ixp33_ASAP7_75t_L g1152 ( 
.A1(n_1079),
.A2(n_347),
.B(n_383),
.C(n_348),
.Y(n_1152)
);

AND2x4_ASAP7_75t_L g1153 ( 
.A(n_1001),
.B(n_739),
.Y(n_1153)
);

AOI21xp5_ASAP7_75t_L g1154 ( 
.A1(n_1033),
.A2(n_740),
.B(n_739),
.Y(n_1154)
);

NOR2xp33_ASAP7_75t_L g1155 ( 
.A(n_1068),
.B(n_722),
.Y(n_1155)
);

INVx1_ASAP7_75t_L g1156 ( 
.A(n_943),
.Y(n_1156)
);

NAND2xp5_ASAP7_75t_SL g1157 ( 
.A(n_954),
.B(n_961),
.Y(n_1157)
);

AND2x2_ASAP7_75t_L g1158 ( 
.A(n_1014),
.B(n_429),
.Y(n_1158)
);

BUFx6f_ASAP7_75t_L g1159 ( 
.A(n_935),
.Y(n_1159)
);

INVx2_ASAP7_75t_L g1160 ( 
.A(n_910),
.Y(n_1160)
);

NAND2xp5_ASAP7_75t_SL g1161 ( 
.A(n_954),
.B(n_746),
.Y(n_1161)
);

O2A1O1Ixp5_ASAP7_75t_SL g1162 ( 
.A1(n_1067),
.A2(n_988),
.B(n_985),
.C(n_967),
.Y(n_1162)
);

AND2x2_ASAP7_75t_L g1163 ( 
.A(n_1016),
.B(n_430),
.Y(n_1163)
);

INVx4_ASAP7_75t_L g1164 ( 
.A(n_935),
.Y(n_1164)
);

HB1xp67_ASAP7_75t_L g1165 ( 
.A(n_961),
.Y(n_1165)
);

AND2x4_ASAP7_75t_L g1166 ( 
.A(n_1001),
.B(n_746),
.Y(n_1166)
);

NAND3xp33_ASAP7_75t_SL g1167 ( 
.A(n_959),
.B(n_431),
.C(n_266),
.Y(n_1167)
);

O2A1O1Ixp33_ASAP7_75t_L g1168 ( 
.A1(n_1020),
.A2(n_319),
.B(n_337),
.C(n_374),
.Y(n_1168)
);

NOR3xp33_ASAP7_75t_SL g1169 ( 
.A(n_946),
.B(n_262),
.C(n_272),
.Y(n_1169)
);

AOI21xp5_ASAP7_75t_L g1170 ( 
.A1(n_977),
.A2(n_388),
.B(n_275),
.Y(n_1170)
);

INVx2_ASAP7_75t_L g1171 ( 
.A(n_918),
.Y(n_1171)
);

INVx1_ASAP7_75t_L g1172 ( 
.A(n_949),
.Y(n_1172)
);

NAND2xp5_ASAP7_75t_L g1173 ( 
.A(n_1076),
.B(n_0),
.Y(n_1173)
);

INVx3_ASAP7_75t_L g1174 ( 
.A(n_935),
.Y(n_1174)
);

AOI33xp33_ASAP7_75t_L g1175 ( 
.A1(n_958),
.A2(n_990),
.A3(n_986),
.B1(n_983),
.B2(n_981),
.B3(n_980),
.Y(n_1175)
);

O2A1O1Ixp33_ASAP7_75t_L g1176 ( 
.A1(n_1072),
.A2(n_0),
.B(n_3),
.C(n_4),
.Y(n_1176)
);

OAI22xp5_ASAP7_75t_L g1177 ( 
.A1(n_961),
.A2(n_307),
.B1(n_286),
.B2(n_386),
.Y(n_1177)
);

AOI22x1_ASAP7_75t_L g1178 ( 
.A1(n_969),
.A2(n_519),
.B1(n_293),
.B2(n_380),
.Y(n_1178)
);

OAI22xp5_ASAP7_75t_L g1179 ( 
.A1(n_1073),
.A2(n_299),
.B1(n_379),
.B2(n_377),
.Y(n_1179)
);

INVx3_ASAP7_75t_L g1180 ( 
.A(n_930),
.Y(n_1180)
);

AOI221xp5_ASAP7_75t_L g1181 ( 
.A1(n_991),
.A2(n_302),
.B1(n_300),
.B2(n_519),
.C(n_361),
.Y(n_1181)
);

INVx1_ASAP7_75t_L g1182 ( 
.A(n_966),
.Y(n_1182)
);

AOI21xp5_ASAP7_75t_L g1183 ( 
.A1(n_1010),
.A2(n_394),
.B(n_361),
.Y(n_1183)
);

NAND2xp5_ASAP7_75t_SL g1184 ( 
.A(n_962),
.B(n_519),
.Y(n_1184)
);

INVx1_ASAP7_75t_L g1185 ( 
.A(n_968),
.Y(n_1185)
);

INVx1_ASAP7_75t_L g1186 ( 
.A(n_973),
.Y(n_1186)
);

NAND2xp5_ASAP7_75t_L g1187 ( 
.A(n_941),
.B(n_3),
.Y(n_1187)
);

INVx1_ASAP7_75t_SL g1188 ( 
.A(n_934),
.Y(n_1188)
);

INVx2_ASAP7_75t_L g1189 ( 
.A(n_918),
.Y(n_1189)
);

HB1xp67_ASAP7_75t_L g1190 ( 
.A(n_1052),
.Y(n_1190)
);

INVx2_ASAP7_75t_L g1191 ( 
.A(n_926),
.Y(n_1191)
);

INVx1_ASAP7_75t_L g1192 ( 
.A(n_1035),
.Y(n_1192)
);

OR2x2_ASAP7_75t_L g1193 ( 
.A(n_1013),
.B(n_519),
.Y(n_1193)
);

NAND2xp5_ASAP7_75t_SL g1194 ( 
.A(n_962),
.B(n_519),
.Y(n_1194)
);

INVx2_ASAP7_75t_L g1195 ( 
.A(n_945),
.Y(n_1195)
);

INVx1_ASAP7_75t_L g1196 ( 
.A(n_1040),
.Y(n_1196)
);

A2O1A1Ixp33_ASAP7_75t_L g1197 ( 
.A1(n_1072),
.A2(n_394),
.B(n_277),
.C(n_8),
.Y(n_1197)
);

AO21x1_ASAP7_75t_L g1198 ( 
.A1(n_1005),
.A2(n_277),
.B(n_201),
.Y(n_1198)
);

OAI22xp5_ASAP7_75t_L g1199 ( 
.A1(n_1073),
.A2(n_277),
.B1(n_7),
.B2(n_8),
.Y(n_1199)
);

INVx2_ASAP7_75t_L g1200 ( 
.A(n_945),
.Y(n_1200)
);

NOR3xp33_ASAP7_75t_SL g1201 ( 
.A(n_919),
.B(n_923),
.C(n_997),
.Y(n_1201)
);

OAI22xp5_ASAP7_75t_L g1202 ( 
.A1(n_1057),
.A2(n_4),
.B1(n_9),
.B2(n_10),
.Y(n_1202)
);

AOI33xp33_ASAP7_75t_L g1203 ( 
.A1(n_1015),
.A2(n_9),
.A3(n_11),
.B1(n_13),
.B2(n_14),
.B3(n_15),
.Y(n_1203)
);

CKINVDCx16_ASAP7_75t_R g1204 ( 
.A(n_1028),
.Y(n_1204)
);

AOI22x1_ASAP7_75t_L g1205 ( 
.A1(n_969),
.A2(n_18),
.B1(n_20),
.B2(n_21),
.Y(n_1205)
);

NAND2xp5_ASAP7_75t_SL g1206 ( 
.A(n_962),
.B(n_21),
.Y(n_1206)
);

AND2x2_ASAP7_75t_L g1207 ( 
.A(n_917),
.B(n_24),
.Y(n_1207)
);

NAND2xp5_ASAP7_75t_SL g1208 ( 
.A(n_994),
.B(n_26),
.Y(n_1208)
);

NAND2xp5_ASAP7_75t_L g1209 ( 
.A(n_992),
.B(n_28),
.Y(n_1209)
);

INVx2_ASAP7_75t_L g1210 ( 
.A(n_953),
.Y(n_1210)
);

NOR2xp33_ASAP7_75t_R g1211 ( 
.A(n_920),
.B(n_182),
.Y(n_1211)
);

BUFx12f_ASAP7_75t_L g1212 ( 
.A(n_951),
.Y(n_1212)
);

AOI21xp5_ASAP7_75t_L g1213 ( 
.A1(n_1025),
.A2(n_922),
.B(n_942),
.Y(n_1213)
);

INVx2_ASAP7_75t_L g1214 ( 
.A(n_953),
.Y(n_1214)
);

OAI22xp5_ASAP7_75t_L g1215 ( 
.A1(n_1015),
.A2(n_916),
.B1(n_982),
.B2(n_1017),
.Y(n_1215)
);

NAND2xp5_ASAP7_75t_L g1216 ( 
.A(n_916),
.B(n_28),
.Y(n_1216)
);

BUFx2_ASAP7_75t_L g1217 ( 
.A(n_1028),
.Y(n_1217)
);

NAND2xp5_ASAP7_75t_L g1218 ( 
.A(n_916),
.B(n_29),
.Y(n_1218)
);

AOI22xp33_ASAP7_75t_L g1219 ( 
.A1(n_982),
.A2(n_35),
.B1(n_38),
.B2(n_40),
.Y(n_1219)
);

NAND3xp33_ASAP7_75t_L g1220 ( 
.A(n_1006),
.B(n_38),
.C(n_46),
.Y(n_1220)
);

NAND2xp5_ASAP7_75t_SL g1221 ( 
.A(n_994),
.B(n_47),
.Y(n_1221)
);

BUFx6f_ASAP7_75t_L g1222 ( 
.A(n_994),
.Y(n_1222)
);

OAI22xp5_ASAP7_75t_L g1223 ( 
.A1(n_975),
.A2(n_48),
.B1(n_50),
.B2(n_52),
.Y(n_1223)
);

INVx1_ASAP7_75t_L g1224 ( 
.A(n_1046),
.Y(n_1224)
);

BUFx3_ASAP7_75t_L g1225 ( 
.A(n_979),
.Y(n_1225)
);

OAI22xp5_ASAP7_75t_L g1226 ( 
.A1(n_920),
.A2(n_48),
.B1(n_53),
.B2(n_55),
.Y(n_1226)
);

BUFx12f_ASAP7_75t_L g1227 ( 
.A(n_1066),
.Y(n_1227)
);

NAND2xp5_ASAP7_75t_SL g1228 ( 
.A(n_1089),
.B(n_947),
.Y(n_1228)
);

INVx1_ASAP7_75t_SL g1229 ( 
.A(n_1083),
.Y(n_1229)
);

INVx1_ASAP7_75t_L g1230 ( 
.A(n_1088),
.Y(n_1230)
);

NAND2xp5_ASAP7_75t_L g1231 ( 
.A(n_1100),
.B(n_1078),
.Y(n_1231)
);

AND2x2_ASAP7_75t_L g1232 ( 
.A(n_1137),
.B(n_936),
.Y(n_1232)
);

OAI21x1_ASAP7_75t_L g1233 ( 
.A1(n_1107),
.A2(n_1162),
.B(n_1114),
.Y(n_1233)
);

AOI21xp5_ASAP7_75t_SL g1234 ( 
.A1(n_1112),
.A2(n_947),
.B(n_1012),
.Y(n_1234)
);

NAND2xp5_ASAP7_75t_L g1235 ( 
.A(n_1110),
.B(n_1052),
.Y(n_1235)
);

INVx1_ASAP7_75t_SL g1236 ( 
.A(n_1118),
.Y(n_1236)
);

A2O1A1Ixp33_ASAP7_75t_L g1237 ( 
.A1(n_1090),
.A2(n_976),
.B(n_939),
.C(n_1032),
.Y(n_1237)
);

OAI21x1_ASAP7_75t_L g1238 ( 
.A1(n_1213),
.A2(n_984),
.B(n_960),
.Y(n_1238)
);

CKINVDCx20_ASAP7_75t_R g1239 ( 
.A(n_1141),
.Y(n_1239)
);

NAND3xp33_ASAP7_75t_L g1240 ( 
.A(n_1080),
.B(n_1042),
.C(n_1026),
.Y(n_1240)
);

AND2x2_ASAP7_75t_L g1241 ( 
.A(n_1108),
.B(n_955),
.Y(n_1241)
);

NAND3xp33_ASAP7_75t_L g1242 ( 
.A(n_1219),
.B(n_1077),
.C(n_1074),
.Y(n_1242)
);

BUFx2_ASAP7_75t_L g1243 ( 
.A(n_1133),
.Y(n_1243)
);

AOI21xp5_ASAP7_75t_SL g1244 ( 
.A1(n_1112),
.A2(n_947),
.B(n_993),
.Y(n_1244)
);

AOI21xp5_ASAP7_75t_L g1245 ( 
.A1(n_1105),
.A2(n_904),
.B(n_919),
.Y(n_1245)
);

NOR2xp33_ASAP7_75t_L g1246 ( 
.A(n_1148),
.B(n_1011),
.Y(n_1246)
);

BUFx6f_ASAP7_75t_L g1247 ( 
.A(n_1142),
.Y(n_1247)
);

INVx1_ASAP7_75t_L g1248 ( 
.A(n_1113),
.Y(n_1248)
);

NAND2x1p5_ASAP7_75t_L g1249 ( 
.A(n_1157),
.B(n_930),
.Y(n_1249)
);

BUFx8_ASAP7_75t_SL g1250 ( 
.A(n_1091),
.Y(n_1250)
);

OA21x2_ASAP7_75t_L g1251 ( 
.A1(n_1198),
.A2(n_1034),
.B(n_1038),
.Y(n_1251)
);

AOI211x1_ASAP7_75t_L g1252 ( 
.A1(n_1173),
.A2(n_1067),
.B(n_1019),
.C(n_1000),
.Y(n_1252)
);

INVx4_ASAP7_75t_L g1253 ( 
.A(n_1086),
.Y(n_1253)
);

INVxp67_ASAP7_75t_L g1254 ( 
.A(n_1104),
.Y(n_1254)
);

AOI22xp5_ASAP7_75t_L g1255 ( 
.A1(n_1148),
.A2(n_939),
.B1(n_1062),
.B2(n_1077),
.Y(n_1255)
);

INVx1_ASAP7_75t_L g1256 ( 
.A(n_1120),
.Y(n_1256)
);

NAND2xp5_ASAP7_75t_L g1257 ( 
.A(n_1136),
.B(n_1023),
.Y(n_1257)
);

CKINVDCx8_ASAP7_75t_R g1258 ( 
.A(n_1204),
.Y(n_1258)
);

A2O1A1Ixp33_ASAP7_75t_L g1259 ( 
.A1(n_1168),
.A2(n_1074),
.B(n_1075),
.C(n_1069),
.Y(n_1259)
);

INVx2_ASAP7_75t_SL g1260 ( 
.A(n_1098),
.Y(n_1260)
);

OAI21x1_ASAP7_75t_SL g1261 ( 
.A1(n_1219),
.A2(n_1048),
.B(n_1053),
.Y(n_1261)
);

NAND2xp5_ASAP7_75t_L g1262 ( 
.A(n_1110),
.B(n_957),
.Y(n_1262)
);

INVx3_ASAP7_75t_L g1263 ( 
.A(n_1159),
.Y(n_1263)
);

NAND2xp5_ASAP7_75t_L g1264 ( 
.A(n_1134),
.B(n_957),
.Y(n_1264)
);

AOI21xp5_ASAP7_75t_L g1265 ( 
.A1(n_1106),
.A2(n_994),
.B(n_1019),
.Y(n_1265)
);

BUFx6f_ASAP7_75t_SL g1266 ( 
.A(n_1151),
.Y(n_1266)
);

INVx3_ASAP7_75t_L g1267 ( 
.A(n_1159),
.Y(n_1267)
);

AO31x2_ASAP7_75t_L g1268 ( 
.A1(n_1215),
.A2(n_1059),
.A3(n_965),
.B(n_972),
.Y(n_1268)
);

OAI22x1_ASAP7_75t_L g1269 ( 
.A1(n_1130),
.A2(n_1071),
.B1(n_1066),
.B2(n_1060),
.Y(n_1269)
);

AO22x2_ASAP7_75t_L g1270 ( 
.A1(n_1093),
.A2(n_1071),
.B1(n_1050),
.B2(n_1061),
.Y(n_1270)
);

OAI21x1_ASAP7_75t_L g1271 ( 
.A1(n_1143),
.A2(n_1047),
.B(n_972),
.Y(n_1271)
);

OAI21x1_ASAP7_75t_L g1272 ( 
.A1(n_1154),
.A2(n_1047),
.B(n_1030),
.Y(n_1272)
);

AOI21xp5_ASAP7_75t_L g1273 ( 
.A1(n_1099),
.A2(n_1116),
.B(n_1082),
.Y(n_1273)
);

AOI21xp5_ASAP7_75t_L g1274 ( 
.A1(n_1087),
.A2(n_1021),
.B(n_1056),
.Y(n_1274)
);

AOI21x1_ASAP7_75t_L g1275 ( 
.A1(n_1097),
.A2(n_1062),
.B(n_1051),
.Y(n_1275)
);

BUFx2_ASAP7_75t_L g1276 ( 
.A(n_1081),
.Y(n_1276)
);

AO31x2_ASAP7_75t_L g1277 ( 
.A1(n_1145),
.A2(n_978),
.A3(n_1037),
.B(n_965),
.Y(n_1277)
);

AND2x4_ASAP7_75t_L g1278 ( 
.A(n_1157),
.B(n_956),
.Y(n_1278)
);

NAND2x1_ASAP7_75t_L g1279 ( 
.A(n_1180),
.B(n_998),
.Y(n_1279)
);

AOI21x1_ASAP7_75t_L g1280 ( 
.A1(n_1184),
.A2(n_978),
.B(n_1059),
.Y(n_1280)
);

INVx3_ASAP7_75t_L g1281 ( 
.A(n_1159),
.Y(n_1281)
);

INVx2_ASAP7_75t_SL g1282 ( 
.A(n_1227),
.Y(n_1282)
);

INVx1_ASAP7_75t_L g1283 ( 
.A(n_1132),
.Y(n_1283)
);

OAI21x1_ASAP7_75t_L g1284 ( 
.A1(n_1184),
.A2(n_1039),
.B(n_1049),
.Y(n_1284)
);

AO32x2_ASAP7_75t_L g1285 ( 
.A1(n_1223),
.A2(n_1045),
.A3(n_1066),
.B1(n_1049),
.B2(n_1039),
.Y(n_1285)
);

AO31x2_ASAP7_75t_L g1286 ( 
.A1(n_1145),
.A2(n_1063),
.A3(n_1061),
.B(n_1045),
.Y(n_1286)
);

OR2x2_ASAP7_75t_L g1287 ( 
.A(n_1126),
.B(n_1023),
.Y(n_1287)
);

AOI21xp5_ASAP7_75t_L g1288 ( 
.A1(n_1209),
.A2(n_1127),
.B(n_1101),
.Y(n_1288)
);

AOI22xp5_ASAP7_75t_L g1289 ( 
.A1(n_1140),
.A2(n_998),
.B1(n_1066),
.B2(n_1036),
.Y(n_1289)
);

NAND2xp5_ASAP7_75t_L g1290 ( 
.A(n_1095),
.B(n_1036),
.Y(n_1290)
);

AOI21xp5_ASAP7_75t_L g1291 ( 
.A1(n_1125),
.A2(n_1041),
.B(n_1027),
.Y(n_1291)
);

OAI21x1_ASAP7_75t_L g1292 ( 
.A1(n_1194),
.A2(n_1027),
.B(n_1063),
.Y(n_1292)
);

NOR2xp67_ASAP7_75t_SL g1293 ( 
.A(n_1212),
.B(n_1041),
.Y(n_1293)
);

NAND2xp5_ASAP7_75t_SL g1294 ( 
.A(n_1217),
.B(n_1041),
.Y(n_1294)
);

AO31x2_ASAP7_75t_L g1295 ( 
.A1(n_1197),
.A2(n_1064),
.A3(n_998),
.B(n_99),
.Y(n_1295)
);

BUFx6f_ASAP7_75t_L g1296 ( 
.A(n_1225),
.Y(n_1296)
);

AOI22xp33_ASAP7_75t_L g1297 ( 
.A1(n_1130),
.A2(n_1064),
.B1(n_998),
.B2(n_62),
.Y(n_1297)
);

NAND3xp33_ASAP7_75t_L g1298 ( 
.A(n_1203),
.B(n_998),
.C(n_59),
.Y(n_1298)
);

NOR2xp33_ASAP7_75t_L g1299 ( 
.A(n_1109),
.B(n_57),
.Y(n_1299)
);

INVx3_ASAP7_75t_L g1300 ( 
.A(n_1159),
.Y(n_1300)
);

AOI221x1_ASAP7_75t_L g1301 ( 
.A1(n_1152),
.A2(n_57),
.B1(n_59),
.B2(n_62),
.C(n_63),
.Y(n_1301)
);

BUFx3_ASAP7_75t_L g1302 ( 
.A(n_1144),
.Y(n_1302)
);

INVx1_ASAP7_75t_L g1303 ( 
.A(n_1150),
.Y(n_1303)
);

CKINVDCx6p67_ASAP7_75t_R g1304 ( 
.A(n_1207),
.Y(n_1304)
);

INVx1_ASAP7_75t_SL g1305 ( 
.A(n_1123),
.Y(n_1305)
);

INVx1_ASAP7_75t_L g1306 ( 
.A(n_1156),
.Y(n_1306)
);

NAND2xp5_ASAP7_75t_L g1307 ( 
.A(n_1095),
.B(n_64),
.Y(n_1307)
);

INVx2_ASAP7_75t_L g1308 ( 
.A(n_1092),
.Y(n_1308)
);

OAI21xp33_ASAP7_75t_L g1309 ( 
.A1(n_1203),
.A2(n_64),
.B(n_65),
.Y(n_1309)
);

OAI21xp5_ASAP7_75t_L g1310 ( 
.A1(n_1152),
.A2(n_65),
.B(n_66),
.Y(n_1310)
);

NAND3xp33_ASAP7_75t_L g1311 ( 
.A(n_1197),
.B(n_68),
.C(n_69),
.Y(n_1311)
);

BUFx3_ASAP7_75t_L g1312 ( 
.A(n_1153),
.Y(n_1312)
);

INVxp67_ASAP7_75t_L g1313 ( 
.A(n_1155),
.Y(n_1313)
);

AOI221xp5_ASAP7_75t_SL g1314 ( 
.A1(n_1199),
.A2(n_70),
.B1(n_72),
.B2(n_74),
.C(n_78),
.Y(n_1314)
);

AOI21x1_ASAP7_75t_L g1315 ( 
.A1(n_1117),
.A2(n_129),
.B(n_80),
.Y(n_1315)
);

NAND3xp33_ASAP7_75t_L g1316 ( 
.A(n_1205),
.B(n_70),
.C(n_84),
.Y(n_1316)
);

AOI21xp5_ASAP7_75t_L g1317 ( 
.A1(n_1125),
.A2(n_88),
.B(n_90),
.Y(n_1317)
);

AO31x2_ASAP7_75t_L g1318 ( 
.A1(n_1111),
.A2(n_93),
.A3(n_98),
.B(n_105),
.Y(n_1318)
);

AO31x2_ASAP7_75t_L g1319 ( 
.A1(n_1121),
.A2(n_109),
.A3(n_116),
.B(n_117),
.Y(n_1319)
);

INVx3_ASAP7_75t_L g1320 ( 
.A(n_1138),
.Y(n_1320)
);

NOR3xp33_ASAP7_75t_L g1321 ( 
.A(n_1220),
.B(n_142),
.C(n_146),
.Y(n_1321)
);

INVx2_ASAP7_75t_L g1322 ( 
.A(n_1160),
.Y(n_1322)
);

BUFx12f_ASAP7_75t_L g1323 ( 
.A(n_1138),
.Y(n_1323)
);

NAND2xp5_ASAP7_75t_L g1324 ( 
.A(n_1175),
.B(n_147),
.Y(n_1324)
);

INVx8_ASAP7_75t_L g1325 ( 
.A(n_1135),
.Y(n_1325)
);

NAND2xp5_ASAP7_75t_L g1326 ( 
.A(n_1175),
.B(n_153),
.Y(n_1326)
);

OAI21x1_ASAP7_75t_L g1327 ( 
.A1(n_1183),
.A2(n_156),
.B(n_158),
.Y(n_1327)
);

AOI21xp33_ASAP7_75t_L g1328 ( 
.A1(n_1176),
.A2(n_164),
.B(n_165),
.Y(n_1328)
);

INVx5_ASAP7_75t_L g1329 ( 
.A(n_1135),
.Y(n_1329)
);

INVxp67_ASAP7_75t_L g1330 ( 
.A(n_1155),
.Y(n_1330)
);

AOI21x1_ASAP7_75t_L g1331 ( 
.A1(n_1117),
.A2(n_177),
.B(n_1122),
.Y(n_1331)
);

NAND2xp5_ASAP7_75t_L g1332 ( 
.A(n_1123),
.B(n_1165),
.Y(n_1332)
);

NAND2xp5_ASAP7_75t_L g1333 ( 
.A(n_1094),
.B(n_1096),
.Y(n_1333)
);

AOI21xp5_ASAP7_75t_L g1334 ( 
.A1(n_1103),
.A2(n_1187),
.B(n_1139),
.Y(n_1334)
);

NAND2xp5_ASAP7_75t_SL g1335 ( 
.A(n_1211),
.B(n_1153),
.Y(n_1335)
);

NOR2x1_ASAP7_75t_L g1336 ( 
.A(n_1188),
.B(n_1164),
.Y(n_1336)
);

NOR2x1_ASAP7_75t_SL g1337 ( 
.A(n_1135),
.B(n_1102),
.Y(n_1337)
);

OAI21xp33_ASAP7_75t_SL g1338 ( 
.A1(n_1206),
.A2(n_1208),
.B(n_1221),
.Y(n_1338)
);

AND2x4_ASAP7_75t_L g1339 ( 
.A(n_1165),
.B(n_1166),
.Y(n_1339)
);

OAI21xp5_ASAP7_75t_SL g1340 ( 
.A1(n_1202),
.A2(n_1226),
.B(n_1167),
.Y(n_1340)
);

HB1xp67_ASAP7_75t_L g1341 ( 
.A(n_1216),
.Y(n_1341)
);

NAND2xp5_ASAP7_75t_L g1342 ( 
.A(n_1190),
.B(n_1186),
.Y(n_1342)
);

NOR2xp33_ASAP7_75t_L g1343 ( 
.A(n_1140),
.B(n_1177),
.Y(n_1343)
);

NAND2xp5_ASAP7_75t_L g1344 ( 
.A(n_1190),
.B(n_1172),
.Y(n_1344)
);

OR2x6_ASAP7_75t_L g1345 ( 
.A(n_1102),
.B(n_1166),
.Y(n_1345)
);

OAI21x1_ASAP7_75t_L g1346 ( 
.A1(n_1122),
.A2(n_1178),
.B(n_1085),
.Y(n_1346)
);

A2O1A1Ixp33_ASAP7_75t_L g1347 ( 
.A1(n_1170),
.A2(n_1115),
.B(n_1181),
.C(n_1084),
.Y(n_1347)
);

INVx2_ASAP7_75t_L g1348 ( 
.A(n_1171),
.Y(n_1348)
);

NAND3xp33_ASAP7_75t_SL g1349 ( 
.A(n_1081),
.B(n_1169),
.C(n_1085),
.Y(n_1349)
);

OAI21x1_ASAP7_75t_L g1350 ( 
.A1(n_1224),
.A2(n_1192),
.B(n_1196),
.Y(n_1350)
);

BUFx2_ASAP7_75t_SL g1351 ( 
.A(n_1164),
.Y(n_1351)
);

AND2x4_ASAP7_75t_L g1352 ( 
.A(n_1128),
.B(n_1146),
.Y(n_1352)
);

O2A1O1Ixp33_ASAP7_75t_L g1353 ( 
.A1(n_1206),
.A2(n_1221),
.B(n_1208),
.C(n_1218),
.Y(n_1353)
);

BUFx3_ASAP7_75t_L g1354 ( 
.A(n_1119),
.Y(n_1354)
);

NAND2xp5_ASAP7_75t_L g1355 ( 
.A(n_1182),
.B(n_1185),
.Y(n_1355)
);

O2A1O1Ixp5_ASAP7_75t_L g1356 ( 
.A1(n_1131),
.A2(n_1161),
.B(n_1180),
.C(n_1179),
.Y(n_1356)
);

A2O1A1Ixp33_ASAP7_75t_L g1357 ( 
.A1(n_1149),
.A2(n_1169),
.B(n_1147),
.C(n_1201),
.Y(n_1357)
);

AOI21x1_ASAP7_75t_SL g1358 ( 
.A1(n_1128),
.A2(n_1146),
.B(n_1163),
.Y(n_1358)
);

BUFx2_ASAP7_75t_L g1359 ( 
.A(n_1211),
.Y(n_1359)
);

NOR2xp33_ASAP7_75t_R g1360 ( 
.A(n_1119),
.B(n_1129),
.Y(n_1360)
);

NAND2xp5_ASAP7_75t_L g1361 ( 
.A(n_1189),
.B(n_1191),
.Y(n_1361)
);

NOR2xp33_ASAP7_75t_L g1362 ( 
.A(n_1158),
.B(n_1174),
.Y(n_1362)
);

OAI21x1_ASAP7_75t_L g1363 ( 
.A1(n_1195),
.A2(n_1200),
.B(n_1214),
.Y(n_1363)
);

OAI21x1_ASAP7_75t_L g1364 ( 
.A1(n_1210),
.A2(n_1161),
.B(n_1174),
.Y(n_1364)
);

NAND2xp5_ASAP7_75t_L g1365 ( 
.A(n_1149),
.B(n_1201),
.Y(n_1365)
);

NOR2xp67_ASAP7_75t_L g1366 ( 
.A(n_1193),
.B(n_1222),
.Y(n_1366)
);

INVxp67_ASAP7_75t_SL g1367 ( 
.A(n_1222),
.Y(n_1367)
);

NAND2xp5_ASAP7_75t_L g1368 ( 
.A(n_1222),
.B(n_1124),
.Y(n_1368)
);

INVx1_ASAP7_75t_L g1369 ( 
.A(n_1222),
.Y(n_1369)
);

AOI211x1_ASAP7_75t_L g1370 ( 
.A1(n_1124),
.A2(n_795),
.B(n_860),
.C(n_1173),
.Y(n_1370)
);

OAI21xp5_ASAP7_75t_L g1371 ( 
.A1(n_1124),
.A2(n_909),
.B(n_1105),
.Y(n_1371)
);

INVx1_ASAP7_75t_L g1372 ( 
.A(n_1088),
.Y(n_1372)
);

INVx1_ASAP7_75t_L g1373 ( 
.A(n_1088),
.Y(n_1373)
);

NAND2xp5_ASAP7_75t_L g1374 ( 
.A(n_1100),
.B(n_974),
.Y(n_1374)
);

AND2x2_ASAP7_75t_L g1375 ( 
.A(n_1137),
.B(n_898),
.Y(n_1375)
);

OAI21x1_ASAP7_75t_L g1376 ( 
.A1(n_1107),
.A2(n_1162),
.B(n_1114),
.Y(n_1376)
);

OAI21x1_ASAP7_75t_L g1377 ( 
.A1(n_1107),
.A2(n_1162),
.B(n_1114),
.Y(n_1377)
);

A2O1A1Ixp33_ASAP7_75t_L g1378 ( 
.A1(n_1090),
.A2(n_995),
.B(n_909),
.C(n_1168),
.Y(n_1378)
);

AND2x2_ASAP7_75t_L g1379 ( 
.A(n_1137),
.B(n_898),
.Y(n_1379)
);

BUFx2_ASAP7_75t_L g1380 ( 
.A(n_1141),
.Y(n_1380)
);

BUFx2_ASAP7_75t_L g1381 ( 
.A(n_1141),
.Y(n_1381)
);

AO21x1_ASAP7_75t_L g1382 ( 
.A1(n_1215),
.A2(n_995),
.B(n_964),
.Y(n_1382)
);

A2O1A1Ixp33_ASAP7_75t_L g1383 ( 
.A1(n_1090),
.A2(n_995),
.B(n_909),
.C(n_1168),
.Y(n_1383)
);

INVx1_ASAP7_75t_L g1384 ( 
.A(n_1355),
.Y(n_1384)
);

INVx1_ASAP7_75t_L g1385 ( 
.A(n_1355),
.Y(n_1385)
);

CKINVDCx5p33_ASAP7_75t_R g1386 ( 
.A(n_1250),
.Y(n_1386)
);

AOI21x1_ASAP7_75t_L g1387 ( 
.A1(n_1275),
.A2(n_1273),
.B(n_1274),
.Y(n_1387)
);

OAI21x1_ASAP7_75t_L g1388 ( 
.A1(n_1233),
.A2(n_1377),
.B(n_1376),
.Y(n_1388)
);

NOR2x1_ASAP7_75t_R g1389 ( 
.A(n_1380),
.B(n_1381),
.Y(n_1389)
);

CKINVDCx20_ASAP7_75t_R g1390 ( 
.A(n_1239),
.Y(n_1390)
);

AO21x2_ASAP7_75t_L g1391 ( 
.A1(n_1371),
.A2(n_1280),
.B(n_1368),
.Y(n_1391)
);

AOI21xp5_ASAP7_75t_L g1392 ( 
.A1(n_1378),
.A2(n_1383),
.B(n_1244),
.Y(n_1392)
);

CKINVDCx14_ASAP7_75t_R g1393 ( 
.A(n_1276),
.Y(n_1393)
);

OAI21x1_ASAP7_75t_L g1394 ( 
.A1(n_1271),
.A2(n_1272),
.B(n_1238),
.Y(n_1394)
);

NAND2x1p5_ASAP7_75t_L g1395 ( 
.A(n_1329),
.B(n_1293),
.Y(n_1395)
);

INVx1_ASAP7_75t_L g1396 ( 
.A(n_1230),
.Y(n_1396)
);

OAI21xp5_ASAP7_75t_L g1397 ( 
.A1(n_1240),
.A2(n_1288),
.B(n_1311),
.Y(n_1397)
);

O2A1O1Ixp33_ASAP7_75t_L g1398 ( 
.A1(n_1340),
.A2(n_1310),
.B(n_1237),
.C(n_1307),
.Y(n_1398)
);

NAND3xp33_ASAP7_75t_L g1399 ( 
.A(n_1310),
.B(n_1314),
.C(n_1307),
.Y(n_1399)
);

INVx2_ASAP7_75t_SL g1400 ( 
.A(n_1296),
.Y(n_1400)
);

AOI22xp33_ASAP7_75t_L g1401 ( 
.A1(n_1382),
.A2(n_1309),
.B1(n_1298),
.B2(n_1311),
.Y(n_1401)
);

A2O1A1Ixp33_ASAP7_75t_L g1402 ( 
.A1(n_1298),
.A2(n_1240),
.B(n_1242),
.C(n_1340),
.Y(n_1402)
);

INVx2_ASAP7_75t_L g1403 ( 
.A(n_1350),
.Y(n_1403)
);

O2A1O1Ixp33_ASAP7_75t_L g1404 ( 
.A1(n_1347),
.A2(n_1357),
.B(n_1353),
.C(n_1231),
.Y(n_1404)
);

NAND2xp5_ASAP7_75t_L g1405 ( 
.A(n_1333),
.B(n_1374),
.Y(n_1405)
);

A2O1A1Ixp33_ASAP7_75t_L g1406 ( 
.A1(n_1242),
.A2(n_1371),
.B(n_1338),
.C(n_1255),
.Y(n_1406)
);

OAI21x1_ASAP7_75t_L g1407 ( 
.A1(n_1284),
.A2(n_1331),
.B(n_1265),
.Y(n_1407)
);

OAI21xp33_ASAP7_75t_SL g1408 ( 
.A1(n_1324),
.A2(n_1326),
.B(n_1365),
.Y(n_1408)
);

INVx1_ASAP7_75t_SL g1409 ( 
.A(n_1229),
.Y(n_1409)
);

INVx2_ASAP7_75t_L g1410 ( 
.A(n_1363),
.Y(n_1410)
);

AOI221xp5_ASAP7_75t_L g1411 ( 
.A1(n_1314),
.A2(n_1370),
.B1(n_1328),
.B2(n_1241),
.C(n_1299),
.Y(n_1411)
);

OAI22xp5_ASAP7_75t_L g1412 ( 
.A1(n_1236),
.A2(n_1365),
.B1(n_1297),
.B2(n_1313),
.Y(n_1412)
);

CKINVDCx16_ASAP7_75t_R g1413 ( 
.A(n_1375),
.Y(n_1413)
);

O2A1O1Ixp33_ASAP7_75t_L g1414 ( 
.A1(n_1328),
.A2(n_1261),
.B(n_1330),
.C(n_1326),
.Y(n_1414)
);

OAI21x1_ASAP7_75t_L g1415 ( 
.A1(n_1292),
.A2(n_1245),
.B(n_1346),
.Y(n_1415)
);

BUFx3_ASAP7_75t_L g1416 ( 
.A(n_1247),
.Y(n_1416)
);

AOI22xp33_ASAP7_75t_L g1417 ( 
.A1(n_1379),
.A2(n_1270),
.B1(n_1302),
.B2(n_1232),
.Y(n_1417)
);

INVx1_ASAP7_75t_SL g1418 ( 
.A(n_1229),
.Y(n_1418)
);

OAI221xp5_ASAP7_75t_L g1419 ( 
.A1(n_1343),
.A2(n_1316),
.B1(n_1246),
.B2(n_1321),
.C(n_1259),
.Y(n_1419)
);

CKINVDCx20_ASAP7_75t_R g1420 ( 
.A(n_1258),
.Y(n_1420)
);

OAI22xp5_ASAP7_75t_SL g1421 ( 
.A1(n_1253),
.A2(n_1359),
.B1(n_1236),
.B2(n_1316),
.Y(n_1421)
);

AOI22xp33_ASAP7_75t_L g1422 ( 
.A1(n_1270),
.A2(n_1341),
.B1(n_1287),
.B2(n_1257),
.Y(n_1422)
);

AND2x2_ASAP7_75t_L g1423 ( 
.A(n_1352),
.B(n_1243),
.Y(n_1423)
);

AND2x4_ASAP7_75t_L g1424 ( 
.A(n_1345),
.B(n_1339),
.Y(n_1424)
);

AND2x4_ASAP7_75t_L g1425 ( 
.A(n_1345),
.B(n_1339),
.Y(n_1425)
);

NAND2xp5_ASAP7_75t_L g1426 ( 
.A(n_1254),
.B(n_1342),
.Y(n_1426)
);

AND2x4_ASAP7_75t_L g1427 ( 
.A(n_1345),
.B(n_1337),
.Y(n_1427)
);

AND2x2_ASAP7_75t_L g1428 ( 
.A(n_1352),
.B(n_1362),
.Y(n_1428)
);

OR2x6_ASAP7_75t_L g1429 ( 
.A(n_1325),
.B(n_1234),
.Y(n_1429)
);

OR2x6_ASAP7_75t_SL g1430 ( 
.A(n_1235),
.B(n_1332),
.Y(n_1430)
);

BUFx2_ASAP7_75t_R g1431 ( 
.A(n_1335),
.Y(n_1431)
);

NAND2xp5_ASAP7_75t_L g1432 ( 
.A(n_1342),
.B(n_1344),
.Y(n_1432)
);

AO31x2_ASAP7_75t_L g1433 ( 
.A1(n_1368),
.A2(n_1262),
.A3(n_1290),
.B(n_1324),
.Y(n_1433)
);

AOI22xp33_ASAP7_75t_L g1434 ( 
.A1(n_1235),
.A2(n_1228),
.B1(n_1372),
.B2(n_1306),
.Y(n_1434)
);

OAI21x1_ASAP7_75t_L g1435 ( 
.A1(n_1315),
.A2(n_1251),
.B(n_1364),
.Y(n_1435)
);

BUFx4f_ASAP7_75t_L g1436 ( 
.A(n_1247),
.Y(n_1436)
);

AND2x2_ASAP7_75t_L g1437 ( 
.A(n_1296),
.B(n_1305),
.Y(n_1437)
);

NAND2xp5_ASAP7_75t_SL g1438 ( 
.A(n_1356),
.B(n_1334),
.Y(n_1438)
);

CKINVDCx16_ASAP7_75t_R g1439 ( 
.A(n_1253),
.Y(n_1439)
);

NAND2xp5_ASAP7_75t_L g1440 ( 
.A(n_1344),
.B(n_1332),
.Y(n_1440)
);

INVx2_ASAP7_75t_SL g1441 ( 
.A(n_1296),
.Y(n_1441)
);

INVx1_ASAP7_75t_L g1442 ( 
.A(n_1248),
.Y(n_1442)
);

OAI21x1_ASAP7_75t_L g1443 ( 
.A1(n_1251),
.A2(n_1327),
.B(n_1290),
.Y(n_1443)
);

AND2x2_ASAP7_75t_L g1444 ( 
.A(n_1305),
.B(n_1303),
.Y(n_1444)
);

INVx1_ASAP7_75t_L g1445 ( 
.A(n_1256),
.Y(n_1445)
);

OAI21x1_ASAP7_75t_L g1446 ( 
.A1(n_1291),
.A2(n_1279),
.B(n_1317),
.Y(n_1446)
);

CKINVDCx20_ASAP7_75t_R g1447 ( 
.A(n_1304),
.Y(n_1447)
);

INVx1_ASAP7_75t_L g1448 ( 
.A(n_1283),
.Y(n_1448)
);

INVx1_ASAP7_75t_SL g1449 ( 
.A(n_1260),
.Y(n_1449)
);

BUFx3_ASAP7_75t_L g1450 ( 
.A(n_1247),
.Y(n_1450)
);

BUFx2_ASAP7_75t_SL g1451 ( 
.A(n_1266),
.Y(n_1451)
);

INVx3_ASAP7_75t_L g1452 ( 
.A(n_1295),
.Y(n_1452)
);

AND2x2_ASAP7_75t_L g1453 ( 
.A(n_1373),
.B(n_1312),
.Y(n_1453)
);

AND2x4_ASAP7_75t_L g1454 ( 
.A(n_1278),
.B(n_1329),
.Y(n_1454)
);

AO21x2_ASAP7_75t_L g1455 ( 
.A1(n_1264),
.A2(n_1361),
.B(n_1366),
.Y(n_1455)
);

OR2x6_ASAP7_75t_L g1456 ( 
.A(n_1325),
.B(n_1252),
.Y(n_1456)
);

OR2x2_ASAP7_75t_L g1457 ( 
.A(n_1264),
.B(n_1361),
.Y(n_1457)
);

AND2x4_ASAP7_75t_L g1458 ( 
.A(n_1278),
.B(n_1329),
.Y(n_1458)
);

CKINVDCx11_ASAP7_75t_R g1459 ( 
.A(n_1323),
.Y(n_1459)
);

OAI21x1_ASAP7_75t_L g1460 ( 
.A1(n_1358),
.A2(n_1369),
.B(n_1249),
.Y(n_1460)
);

BUFx3_ASAP7_75t_L g1461 ( 
.A(n_1354),
.Y(n_1461)
);

INVx1_ASAP7_75t_L g1462 ( 
.A(n_1308),
.Y(n_1462)
);

OAI21x1_ASAP7_75t_L g1463 ( 
.A1(n_1249),
.A2(n_1289),
.B(n_1263),
.Y(n_1463)
);

OAI21x1_ASAP7_75t_L g1464 ( 
.A1(n_1263),
.A2(n_1300),
.B(n_1267),
.Y(n_1464)
);

INVx2_ASAP7_75t_L g1465 ( 
.A(n_1268),
.Y(n_1465)
);

BUFx2_ASAP7_75t_L g1466 ( 
.A(n_1360),
.Y(n_1466)
);

OR2x2_ASAP7_75t_L g1467 ( 
.A(n_1322),
.B(n_1348),
.Y(n_1467)
);

AO21x2_ASAP7_75t_L g1468 ( 
.A1(n_1294),
.A2(n_1367),
.B(n_1349),
.Y(n_1468)
);

OAI21x1_ASAP7_75t_L g1469 ( 
.A1(n_1267),
.A2(n_1300),
.B(n_1281),
.Y(n_1469)
);

BUFx3_ASAP7_75t_L g1470 ( 
.A(n_1325),
.Y(n_1470)
);

AOI22xp5_ASAP7_75t_L g1471 ( 
.A1(n_1269),
.A2(n_1266),
.B1(n_1282),
.B2(n_1336),
.Y(n_1471)
);

INVx6_ASAP7_75t_L g1472 ( 
.A(n_1329),
.Y(n_1472)
);

INVx2_ASAP7_75t_L g1473 ( 
.A(n_1277),
.Y(n_1473)
);

OAI21x1_ASAP7_75t_L g1474 ( 
.A1(n_1281),
.A2(n_1320),
.B(n_1301),
.Y(n_1474)
);

INVx4_ASAP7_75t_L g1475 ( 
.A(n_1351),
.Y(n_1475)
);

OAI21x1_ASAP7_75t_L g1476 ( 
.A1(n_1295),
.A2(n_1277),
.B(n_1285),
.Y(n_1476)
);

AND2x4_ASAP7_75t_L g1477 ( 
.A(n_1286),
.B(n_1295),
.Y(n_1477)
);

NAND3xp33_ASAP7_75t_L g1478 ( 
.A(n_1285),
.B(n_1318),
.C(n_1319),
.Y(n_1478)
);

CKINVDCx5p33_ASAP7_75t_R g1479 ( 
.A(n_1285),
.Y(n_1479)
);

INVx1_ASAP7_75t_L g1480 ( 
.A(n_1286),
.Y(n_1480)
);

OAI21x1_ASAP7_75t_L g1481 ( 
.A1(n_1318),
.A2(n_1376),
.B(n_1233),
.Y(n_1481)
);

AO21x2_ASAP7_75t_L g1482 ( 
.A1(n_1318),
.A2(n_1371),
.B(n_1280),
.Y(n_1482)
);

INVx2_ASAP7_75t_L g1483 ( 
.A(n_1319),
.Y(n_1483)
);

BUFx3_ASAP7_75t_L g1484 ( 
.A(n_1319),
.Y(n_1484)
);

INVx3_ASAP7_75t_L g1485 ( 
.A(n_1279),
.Y(n_1485)
);

OA21x2_ASAP7_75t_L g1486 ( 
.A1(n_1233),
.A2(n_1377),
.B(n_1376),
.Y(n_1486)
);

OAI21x1_ASAP7_75t_L g1487 ( 
.A1(n_1233),
.A2(n_1377),
.B(n_1376),
.Y(n_1487)
);

INVxp67_ASAP7_75t_L g1488 ( 
.A(n_1243),
.Y(n_1488)
);

INVx1_ASAP7_75t_L g1489 ( 
.A(n_1355),
.Y(n_1489)
);

INVx2_ASAP7_75t_L g1490 ( 
.A(n_1350),
.Y(n_1490)
);

OR2x2_ASAP7_75t_L g1491 ( 
.A(n_1342),
.B(n_1344),
.Y(n_1491)
);

AND2x4_ASAP7_75t_L g1492 ( 
.A(n_1345),
.B(n_1339),
.Y(n_1492)
);

OAI21xp5_ASAP7_75t_L g1493 ( 
.A1(n_1383),
.A2(n_909),
.B(n_995),
.Y(n_1493)
);

OAI21x1_ASAP7_75t_SL g1494 ( 
.A1(n_1310),
.A2(n_1382),
.B(n_1288),
.Y(n_1494)
);

OAI21x1_ASAP7_75t_L g1495 ( 
.A1(n_1233),
.A2(n_1377),
.B(n_1376),
.Y(n_1495)
);

INVx1_ASAP7_75t_L g1496 ( 
.A(n_1355),
.Y(n_1496)
);

OAI21x1_ASAP7_75t_L g1497 ( 
.A1(n_1233),
.A2(n_1377),
.B(n_1376),
.Y(n_1497)
);

HB1xp67_ASAP7_75t_L g1498 ( 
.A(n_1236),
.Y(n_1498)
);

OA21x2_ASAP7_75t_L g1499 ( 
.A1(n_1233),
.A2(n_1377),
.B(n_1376),
.Y(n_1499)
);

INVx2_ASAP7_75t_L g1500 ( 
.A(n_1350),
.Y(n_1500)
);

OAI21xp33_ASAP7_75t_L g1501 ( 
.A1(n_1309),
.A2(n_909),
.B(n_995),
.Y(n_1501)
);

CKINVDCx6p67_ASAP7_75t_R g1502 ( 
.A(n_1239),
.Y(n_1502)
);

OAI21x1_ASAP7_75t_L g1503 ( 
.A1(n_1233),
.A2(n_1377),
.B(n_1376),
.Y(n_1503)
);

OAI21xp5_ASAP7_75t_L g1504 ( 
.A1(n_1383),
.A2(n_909),
.B(n_995),
.Y(n_1504)
);

OR2x6_ASAP7_75t_L g1505 ( 
.A(n_1325),
.B(n_1234),
.Y(n_1505)
);

BUFx2_ASAP7_75t_L g1506 ( 
.A(n_1243),
.Y(n_1506)
);

OAI21x1_ASAP7_75t_L g1507 ( 
.A1(n_1233),
.A2(n_1377),
.B(n_1376),
.Y(n_1507)
);

INVx2_ASAP7_75t_L g1508 ( 
.A(n_1350),
.Y(n_1508)
);

OAI21x1_ASAP7_75t_L g1509 ( 
.A1(n_1233),
.A2(n_1377),
.B(n_1376),
.Y(n_1509)
);

NAND2xp5_ASAP7_75t_L g1510 ( 
.A(n_1333),
.B(n_1374),
.Y(n_1510)
);

OAI22xp5_ASAP7_75t_SL g1511 ( 
.A1(n_1299),
.A2(n_1055),
.B1(n_1109),
.B2(n_898),
.Y(n_1511)
);

AND2x2_ASAP7_75t_L g1512 ( 
.A(n_1375),
.B(n_1379),
.Y(n_1512)
);

HB1xp67_ASAP7_75t_L g1513 ( 
.A(n_1236),
.Y(n_1513)
);

OAI21x1_ASAP7_75t_L g1514 ( 
.A1(n_1233),
.A2(n_1377),
.B(n_1376),
.Y(n_1514)
);

NAND2xp5_ASAP7_75t_L g1515 ( 
.A(n_1333),
.B(n_1374),
.Y(n_1515)
);

AOI21xp5_ASAP7_75t_L g1516 ( 
.A1(n_1378),
.A2(n_1383),
.B(n_1105),
.Y(n_1516)
);

OA21x2_ASAP7_75t_L g1517 ( 
.A1(n_1233),
.A2(n_1377),
.B(n_1376),
.Y(n_1517)
);

INVx1_ASAP7_75t_SL g1518 ( 
.A(n_1229),
.Y(n_1518)
);

AOI21x1_ASAP7_75t_L g1519 ( 
.A1(n_1275),
.A2(n_1273),
.B(n_1274),
.Y(n_1519)
);

INVx6_ASAP7_75t_L g1520 ( 
.A(n_1247),
.Y(n_1520)
);

AO31x2_ASAP7_75t_L g1521 ( 
.A1(n_1382),
.A2(n_1198),
.A3(n_1368),
.B(n_1273),
.Y(n_1521)
);

INVx2_ASAP7_75t_L g1522 ( 
.A(n_1350),
.Y(n_1522)
);

OAI21xp5_ASAP7_75t_L g1523 ( 
.A1(n_1383),
.A2(n_909),
.B(n_995),
.Y(n_1523)
);

OAI22xp5_ASAP7_75t_L g1524 ( 
.A1(n_1378),
.A2(n_995),
.B1(n_970),
.B2(n_909),
.Y(n_1524)
);

OAI21xp5_ASAP7_75t_L g1525 ( 
.A1(n_1383),
.A2(n_909),
.B(n_995),
.Y(n_1525)
);

INVx2_ASAP7_75t_L g1526 ( 
.A(n_1350),
.Y(n_1526)
);

HB1xp67_ASAP7_75t_L g1527 ( 
.A(n_1236),
.Y(n_1527)
);

AND2x4_ASAP7_75t_L g1528 ( 
.A(n_1345),
.B(n_1339),
.Y(n_1528)
);

INVx1_ASAP7_75t_L g1529 ( 
.A(n_1355),
.Y(n_1529)
);

HB1xp67_ASAP7_75t_L g1530 ( 
.A(n_1236),
.Y(n_1530)
);

OA21x2_ASAP7_75t_L g1531 ( 
.A1(n_1233),
.A2(n_1377),
.B(n_1376),
.Y(n_1531)
);

OR2x6_ASAP7_75t_L g1532 ( 
.A(n_1325),
.B(n_1234),
.Y(n_1532)
);

AND2x4_ASAP7_75t_L g1533 ( 
.A(n_1345),
.B(n_1339),
.Y(n_1533)
);

AO31x2_ASAP7_75t_L g1534 ( 
.A1(n_1382),
.A2(n_1198),
.A3(n_1368),
.B(n_1273),
.Y(n_1534)
);

OAI21x1_ASAP7_75t_L g1535 ( 
.A1(n_1233),
.A2(n_1377),
.B(n_1376),
.Y(n_1535)
);

INVx2_ASAP7_75t_SL g1536 ( 
.A(n_1296),
.Y(n_1536)
);

OAI21x1_ASAP7_75t_L g1537 ( 
.A1(n_1233),
.A2(n_1377),
.B(n_1376),
.Y(n_1537)
);

CKINVDCx5p33_ASAP7_75t_R g1538 ( 
.A(n_1250),
.Y(n_1538)
);

NOR2x1_ASAP7_75t_SL g1539 ( 
.A(n_1345),
.B(n_1329),
.Y(n_1539)
);

INVx1_ASAP7_75t_L g1540 ( 
.A(n_1355),
.Y(n_1540)
);

INVx1_ASAP7_75t_L g1541 ( 
.A(n_1355),
.Y(n_1541)
);

OA21x2_ASAP7_75t_L g1542 ( 
.A1(n_1233),
.A2(n_1377),
.B(n_1376),
.Y(n_1542)
);

NAND2xp5_ASAP7_75t_L g1543 ( 
.A(n_1333),
.B(n_1374),
.Y(n_1543)
);

BUFx2_ASAP7_75t_L g1544 ( 
.A(n_1243),
.Y(n_1544)
);

INVx2_ASAP7_75t_L g1545 ( 
.A(n_1350),
.Y(n_1545)
);

NAND2xp5_ASAP7_75t_L g1546 ( 
.A(n_1333),
.B(n_1374),
.Y(n_1546)
);

OAI21xp5_ASAP7_75t_L g1547 ( 
.A1(n_1383),
.A2(n_909),
.B(n_995),
.Y(n_1547)
);

BUFx2_ASAP7_75t_L g1548 ( 
.A(n_1243),
.Y(n_1548)
);

OAI22xp5_ASAP7_75t_L g1549 ( 
.A1(n_1378),
.A2(n_995),
.B1(n_970),
.B2(n_909),
.Y(n_1549)
);

INVx1_ASAP7_75t_L g1550 ( 
.A(n_1355),
.Y(n_1550)
);

OAI21xp5_ASAP7_75t_L g1551 ( 
.A1(n_1383),
.A2(n_909),
.B(n_995),
.Y(n_1551)
);

OR2x2_ASAP7_75t_L g1552 ( 
.A(n_1342),
.B(n_1344),
.Y(n_1552)
);

OAI21x1_ASAP7_75t_L g1553 ( 
.A1(n_1233),
.A2(n_1377),
.B(n_1376),
.Y(n_1553)
);

AND2x4_ASAP7_75t_L g1554 ( 
.A(n_1345),
.B(n_1339),
.Y(n_1554)
);

INVx3_ASAP7_75t_L g1555 ( 
.A(n_1475),
.Y(n_1555)
);

A2O1A1Ixp33_ASAP7_75t_L g1556 ( 
.A1(n_1392),
.A2(n_1398),
.B(n_1501),
.C(n_1523),
.Y(n_1556)
);

AOI221x1_ASAP7_75t_SL g1557 ( 
.A1(n_1524),
.A2(n_1549),
.B1(n_1399),
.B2(n_1426),
.C(n_1405),
.Y(n_1557)
);

AOI21xp5_ASAP7_75t_SL g1558 ( 
.A1(n_1402),
.A2(n_1504),
.B(n_1493),
.Y(n_1558)
);

NAND2xp5_ASAP7_75t_L g1559 ( 
.A(n_1432),
.B(n_1440),
.Y(n_1559)
);

AND2x4_ASAP7_75t_L g1560 ( 
.A(n_1424),
.B(n_1425),
.Y(n_1560)
);

OAI22xp5_ASAP7_75t_L g1561 ( 
.A1(n_1402),
.A2(n_1547),
.B1(n_1551),
.B2(n_1525),
.Y(n_1561)
);

INVx2_ASAP7_75t_L g1562 ( 
.A(n_1467),
.Y(n_1562)
);

AOI21xp5_ASAP7_75t_L g1563 ( 
.A1(n_1397),
.A2(n_1516),
.B(n_1438),
.Y(n_1563)
);

CKINVDCx5p33_ASAP7_75t_R g1564 ( 
.A(n_1502),
.Y(n_1564)
);

AND2x2_ASAP7_75t_L g1565 ( 
.A(n_1428),
.B(n_1423),
.Y(n_1565)
);

OR2x2_ASAP7_75t_L g1566 ( 
.A(n_1491),
.B(n_1552),
.Y(n_1566)
);

AND2x2_ASAP7_75t_L g1567 ( 
.A(n_1512),
.B(n_1413),
.Y(n_1567)
);

OR2x2_ASAP7_75t_L g1568 ( 
.A(n_1498),
.B(n_1513),
.Y(n_1568)
);

CKINVDCx16_ASAP7_75t_R g1569 ( 
.A(n_1390),
.Y(n_1569)
);

AND2x2_ASAP7_75t_L g1570 ( 
.A(n_1437),
.B(n_1453),
.Y(n_1570)
);

OA21x2_ASAP7_75t_L g1571 ( 
.A1(n_1388),
.A2(n_1495),
.B(n_1487),
.Y(n_1571)
);

HB1xp67_ASAP7_75t_L g1572 ( 
.A(n_1391),
.Y(n_1572)
);

OA21x2_ASAP7_75t_L g1573 ( 
.A1(n_1388),
.A2(n_1495),
.B(n_1487),
.Y(n_1573)
);

INVx1_ASAP7_75t_SL g1574 ( 
.A(n_1420),
.Y(n_1574)
);

HB1xp67_ASAP7_75t_L g1575 ( 
.A(n_1391),
.Y(n_1575)
);

OR2x2_ASAP7_75t_L g1576 ( 
.A(n_1527),
.B(n_1530),
.Y(n_1576)
);

AND2x2_ASAP7_75t_L g1577 ( 
.A(n_1444),
.B(n_1506),
.Y(n_1577)
);

NAND2xp5_ASAP7_75t_L g1578 ( 
.A(n_1510),
.B(n_1515),
.Y(n_1578)
);

CKINVDCx5p33_ASAP7_75t_R g1579 ( 
.A(n_1502),
.Y(n_1579)
);

O2A1O1Ixp5_ASAP7_75t_L g1580 ( 
.A1(n_1406),
.A2(n_1452),
.B(n_1477),
.C(n_1519),
.Y(n_1580)
);

HB1xp67_ASAP7_75t_L g1581 ( 
.A(n_1433),
.Y(n_1581)
);

OR2x2_ASAP7_75t_L g1582 ( 
.A(n_1544),
.B(n_1548),
.Y(n_1582)
);

O2A1O1Ixp33_ASAP7_75t_L g1583 ( 
.A1(n_1419),
.A2(n_1404),
.B(n_1494),
.C(n_1414),
.Y(n_1583)
);

OAI22xp5_ASAP7_75t_L g1584 ( 
.A1(n_1401),
.A2(n_1411),
.B1(n_1393),
.B2(n_1412),
.Y(n_1584)
);

O2A1O1Ixp33_ASAP7_75t_L g1585 ( 
.A1(n_1401),
.A2(n_1408),
.B(n_1546),
.C(n_1543),
.Y(n_1585)
);

INVx1_ASAP7_75t_L g1586 ( 
.A(n_1442),
.Y(n_1586)
);

NAND2xp5_ASAP7_75t_L g1587 ( 
.A(n_1384),
.B(n_1385),
.Y(n_1587)
);

INVx1_ASAP7_75t_L g1588 ( 
.A(n_1445),
.Y(n_1588)
);

AND2x4_ASAP7_75t_L g1589 ( 
.A(n_1424),
.B(n_1425),
.Y(n_1589)
);

AND2x2_ASAP7_75t_L g1590 ( 
.A(n_1409),
.B(n_1418),
.Y(n_1590)
);

BUFx8_ASAP7_75t_SL g1591 ( 
.A(n_1390),
.Y(n_1591)
);

OR2x2_ASAP7_75t_L g1592 ( 
.A(n_1518),
.B(n_1489),
.Y(n_1592)
);

AOI22xp5_ASAP7_75t_L g1593 ( 
.A1(n_1511),
.A2(n_1417),
.B1(n_1421),
.B2(n_1434),
.Y(n_1593)
);

OAI22xp5_ASAP7_75t_L g1594 ( 
.A1(n_1393),
.A2(n_1488),
.B1(n_1417),
.B2(n_1447),
.Y(n_1594)
);

BUFx12f_ASAP7_75t_L g1595 ( 
.A(n_1386),
.Y(n_1595)
);

AOI21xp5_ASAP7_75t_SL g1596 ( 
.A1(n_1429),
.A2(n_1505),
.B(n_1532),
.Y(n_1596)
);

AOI21xp5_ASAP7_75t_SL g1597 ( 
.A1(n_1429),
.A2(n_1505),
.B(n_1532),
.Y(n_1597)
);

AOI221x1_ASAP7_75t_SL g1598 ( 
.A1(n_1448),
.A2(n_1529),
.B1(n_1550),
.B2(n_1496),
.C(n_1541),
.Y(n_1598)
);

OAI31xp33_ASAP7_75t_L g1599 ( 
.A1(n_1434),
.A2(n_1449),
.A3(n_1478),
.B(n_1422),
.Y(n_1599)
);

OA21x2_ASAP7_75t_L g1600 ( 
.A1(n_1497),
.A2(n_1503),
.B(n_1514),
.Y(n_1600)
);

CKINVDCx14_ASAP7_75t_R g1601 ( 
.A(n_1386),
.Y(n_1601)
);

O2A1O1Ixp5_ASAP7_75t_L g1602 ( 
.A1(n_1452),
.A2(n_1477),
.B(n_1387),
.C(n_1500),
.Y(n_1602)
);

NAND2xp5_ASAP7_75t_L g1603 ( 
.A(n_1540),
.B(n_1430),
.Y(n_1603)
);

OAI22xp5_ASAP7_75t_L g1604 ( 
.A1(n_1447),
.A2(n_1479),
.B1(n_1430),
.B2(n_1466),
.Y(n_1604)
);

AND2x2_ASAP7_75t_L g1605 ( 
.A(n_1492),
.B(n_1528),
.Y(n_1605)
);

BUFx6f_ASAP7_75t_L g1606 ( 
.A(n_1436),
.Y(n_1606)
);

AND2x2_ASAP7_75t_L g1607 ( 
.A(n_1533),
.B(n_1554),
.Y(n_1607)
);

AND2x4_ASAP7_75t_L g1608 ( 
.A(n_1533),
.B(n_1554),
.Y(n_1608)
);

INVx2_ASAP7_75t_L g1609 ( 
.A(n_1462),
.Y(n_1609)
);

AND2x2_ASAP7_75t_L g1610 ( 
.A(n_1461),
.B(n_1416),
.Y(n_1610)
);

AND2x4_ASAP7_75t_L g1611 ( 
.A(n_1427),
.B(n_1454),
.Y(n_1611)
);

AND2x2_ASAP7_75t_L g1612 ( 
.A(n_1450),
.B(n_1400),
.Y(n_1612)
);

NAND2xp5_ASAP7_75t_L g1613 ( 
.A(n_1457),
.B(n_1400),
.Y(n_1613)
);

BUFx6f_ASAP7_75t_L g1614 ( 
.A(n_1436),
.Y(n_1614)
);

CKINVDCx12_ASAP7_75t_R g1615 ( 
.A(n_1389),
.Y(n_1615)
);

CKINVDCx20_ASAP7_75t_R g1616 ( 
.A(n_1538),
.Y(n_1616)
);

NAND2xp5_ASAP7_75t_L g1617 ( 
.A(n_1441),
.B(n_1536),
.Y(n_1617)
);

OR2x2_ASAP7_75t_L g1618 ( 
.A(n_1433),
.B(n_1479),
.Y(n_1618)
);

O2A1O1Ixp5_ASAP7_75t_L g1619 ( 
.A1(n_1403),
.A2(n_1490),
.B(n_1545),
.C(n_1522),
.Y(n_1619)
);

NOR2x1_ASAP7_75t_L g1620 ( 
.A(n_1475),
.B(n_1451),
.Y(n_1620)
);

OR2x2_ASAP7_75t_L g1621 ( 
.A(n_1433),
.B(n_1450),
.Y(n_1621)
);

OA21x2_ASAP7_75t_L g1622 ( 
.A1(n_1497),
.A2(n_1553),
.B(n_1537),
.Y(n_1622)
);

AND2x2_ASAP7_75t_L g1623 ( 
.A(n_1441),
.B(n_1536),
.Y(n_1623)
);

OAI22xp5_ASAP7_75t_L g1624 ( 
.A1(n_1431),
.A2(n_1420),
.B1(n_1439),
.B2(n_1436),
.Y(n_1624)
);

OR2x2_ASAP7_75t_L g1625 ( 
.A(n_1433),
.B(n_1422),
.Y(n_1625)
);

NAND2xp5_ASAP7_75t_L g1626 ( 
.A(n_1520),
.B(n_1471),
.Y(n_1626)
);

AND2x4_ASAP7_75t_L g1627 ( 
.A(n_1427),
.B(n_1454),
.Y(n_1627)
);

INVx1_ASAP7_75t_L g1628 ( 
.A(n_1455),
.Y(n_1628)
);

NAND2xp5_ASAP7_75t_L g1629 ( 
.A(n_1520),
.B(n_1455),
.Y(n_1629)
);

AND2x4_ASAP7_75t_SL g1630 ( 
.A(n_1429),
.B(n_1505),
.Y(n_1630)
);

BUFx4f_ASAP7_75t_SL g1631 ( 
.A(n_1475),
.Y(n_1631)
);

AND2x4_ASAP7_75t_L g1632 ( 
.A(n_1427),
.B(n_1454),
.Y(n_1632)
);

OAI22xp5_ASAP7_75t_L g1633 ( 
.A1(n_1456),
.A2(n_1532),
.B1(n_1520),
.B2(n_1395),
.Y(n_1633)
);

INVx3_ASAP7_75t_SL g1634 ( 
.A(n_1538),
.Y(n_1634)
);

A2O1A1Ixp33_ASAP7_75t_L g1635 ( 
.A1(n_1476),
.A2(n_1484),
.B(n_1463),
.C(n_1443),
.Y(n_1635)
);

NOR2xp33_ASAP7_75t_L g1636 ( 
.A(n_1456),
.B(n_1468),
.Y(n_1636)
);

NAND2xp5_ASAP7_75t_L g1637 ( 
.A(n_1470),
.B(n_1468),
.Y(n_1637)
);

AND2x4_ASAP7_75t_L g1638 ( 
.A(n_1458),
.B(n_1470),
.Y(n_1638)
);

HB1xp67_ASAP7_75t_L g1639 ( 
.A(n_1403),
.Y(n_1639)
);

OAI22xp5_ASAP7_75t_L g1640 ( 
.A1(n_1456),
.A2(n_1395),
.B1(n_1485),
.B2(n_1458),
.Y(n_1640)
);

AND2x2_ASAP7_75t_L g1641 ( 
.A(n_1458),
.B(n_1469),
.Y(n_1641)
);

AND2x4_ASAP7_75t_L g1642 ( 
.A(n_1539),
.B(n_1463),
.Y(n_1642)
);

AND2x2_ASAP7_75t_L g1643 ( 
.A(n_1464),
.B(n_1469),
.Y(n_1643)
);

CKINVDCx20_ASAP7_75t_R g1644 ( 
.A(n_1459),
.Y(n_1644)
);

O2A1O1Ixp33_ASAP7_75t_L g1645 ( 
.A1(n_1490),
.A2(n_1500),
.B(n_1508),
.C(n_1522),
.Y(n_1645)
);

O2A1O1Ixp33_ASAP7_75t_L g1646 ( 
.A1(n_1508),
.A2(n_1526),
.B(n_1545),
.C(n_1485),
.Y(n_1646)
);

OAI22xp5_ASAP7_75t_L g1647 ( 
.A1(n_1485),
.A2(n_1472),
.B1(n_1484),
.B2(n_1480),
.Y(n_1647)
);

AND2x2_ASAP7_75t_L g1648 ( 
.A(n_1460),
.B(n_1474),
.Y(n_1648)
);

HB1xp67_ASAP7_75t_L g1649 ( 
.A(n_1521),
.Y(n_1649)
);

AND2x2_ASAP7_75t_L g1650 ( 
.A(n_1460),
.B(n_1521),
.Y(n_1650)
);

HB1xp67_ASAP7_75t_L g1651 ( 
.A(n_1521),
.Y(n_1651)
);

HB1xp67_ASAP7_75t_L g1652 ( 
.A(n_1521),
.Y(n_1652)
);

HB1xp67_ASAP7_75t_L g1653 ( 
.A(n_1534),
.Y(n_1653)
);

INVx3_ASAP7_75t_L g1654 ( 
.A(n_1472),
.Y(n_1654)
);

AND2x2_ASAP7_75t_L g1655 ( 
.A(n_1534),
.B(n_1459),
.Y(n_1655)
);

AND2x2_ASAP7_75t_L g1656 ( 
.A(n_1534),
.B(n_1482),
.Y(n_1656)
);

OR2x2_ASAP7_75t_L g1657 ( 
.A(n_1476),
.B(n_1473),
.Y(n_1657)
);

AND2x2_ASAP7_75t_L g1658 ( 
.A(n_1486),
.B(n_1499),
.Y(n_1658)
);

AND2x2_ASAP7_75t_L g1659 ( 
.A(n_1499),
.B(n_1517),
.Y(n_1659)
);

AND2x2_ASAP7_75t_L g1660 ( 
.A(n_1531),
.B(n_1542),
.Y(n_1660)
);

OAI22xp5_ASAP7_75t_L g1661 ( 
.A1(n_1483),
.A2(n_1531),
.B1(n_1542),
.B2(n_1465),
.Y(n_1661)
);

BUFx2_ASAP7_75t_R g1662 ( 
.A(n_1503),
.Y(n_1662)
);

O2A1O1Ixp33_ASAP7_75t_L g1663 ( 
.A1(n_1410),
.A2(n_1446),
.B(n_1407),
.C(n_1481),
.Y(n_1663)
);

AND2x4_ASAP7_75t_L g1664 ( 
.A(n_1410),
.B(n_1407),
.Y(n_1664)
);

CKINVDCx5p33_ASAP7_75t_R g1665 ( 
.A(n_1507),
.Y(n_1665)
);

NAND2xp5_ASAP7_75t_L g1666 ( 
.A(n_1415),
.B(n_1514),
.Y(n_1666)
);

HB1xp67_ASAP7_75t_L g1667 ( 
.A(n_1509),
.Y(n_1667)
);

OA21x2_ASAP7_75t_L g1668 ( 
.A1(n_1535),
.A2(n_1537),
.B(n_1553),
.Y(n_1668)
);

CKINVDCx6p67_ASAP7_75t_R g1669 ( 
.A(n_1435),
.Y(n_1669)
);

AND2x2_ASAP7_75t_L g1670 ( 
.A(n_1394),
.B(n_1428),
.Y(n_1670)
);

OAI22xp5_ASAP7_75t_L g1671 ( 
.A1(n_1394),
.A2(n_1402),
.B1(n_1549),
.B2(n_1524),
.Y(n_1671)
);

AND2x4_ASAP7_75t_L g1672 ( 
.A(n_1424),
.B(n_1425),
.Y(n_1672)
);

AOI21xp5_ASAP7_75t_SL g1673 ( 
.A1(n_1524),
.A2(n_1549),
.B(n_1402),
.Y(n_1673)
);

NOR2xp67_ASAP7_75t_L g1674 ( 
.A(n_1475),
.B(n_1471),
.Y(n_1674)
);

AND2x2_ASAP7_75t_L g1675 ( 
.A(n_1428),
.B(n_1423),
.Y(n_1675)
);

AOI21xp5_ASAP7_75t_SL g1676 ( 
.A1(n_1524),
.A2(n_1549),
.B(n_1402),
.Y(n_1676)
);

INVx4_ASAP7_75t_L g1677 ( 
.A(n_1475),
.Y(n_1677)
);

OAI22xp5_ASAP7_75t_L g1678 ( 
.A1(n_1402),
.A2(n_1524),
.B1(n_1549),
.B2(n_995),
.Y(n_1678)
);

NOR2xp67_ASAP7_75t_L g1679 ( 
.A(n_1475),
.B(n_1471),
.Y(n_1679)
);

CKINVDCx5p33_ASAP7_75t_R g1680 ( 
.A(n_1502),
.Y(n_1680)
);

INVx1_ASAP7_75t_L g1681 ( 
.A(n_1396),
.Y(n_1681)
);

AND2x4_ASAP7_75t_L g1682 ( 
.A(n_1424),
.B(n_1425),
.Y(n_1682)
);

O2A1O1Ixp33_ASAP7_75t_L g1683 ( 
.A1(n_1524),
.A2(n_1549),
.B(n_1504),
.C(n_1523),
.Y(n_1683)
);

NAND2xp5_ASAP7_75t_L g1684 ( 
.A(n_1432),
.B(n_1440),
.Y(n_1684)
);

HB1xp67_ASAP7_75t_L g1685 ( 
.A(n_1391),
.Y(n_1685)
);

NAND2xp5_ASAP7_75t_L g1686 ( 
.A(n_1432),
.B(n_1440),
.Y(n_1686)
);

AOI21x1_ASAP7_75t_SL g1687 ( 
.A1(n_1426),
.A2(n_1307),
.B(n_1368),
.Y(n_1687)
);

AOI21xp5_ASAP7_75t_L g1688 ( 
.A1(n_1392),
.A2(n_1504),
.B(n_1493),
.Y(n_1688)
);

AOI21x1_ASAP7_75t_SL g1689 ( 
.A1(n_1426),
.A2(n_1307),
.B(n_1368),
.Y(n_1689)
);

AND2x4_ASAP7_75t_L g1690 ( 
.A(n_1424),
.B(n_1425),
.Y(n_1690)
);

A2O1A1Ixp33_ASAP7_75t_L g1691 ( 
.A1(n_1392),
.A2(n_995),
.B(n_1398),
.C(n_811),
.Y(n_1691)
);

HB1xp67_ASAP7_75t_L g1692 ( 
.A(n_1568),
.Y(n_1692)
);

AOI22xp5_ASAP7_75t_L g1693 ( 
.A1(n_1678),
.A2(n_1561),
.B1(n_1691),
.B2(n_1584),
.Y(n_1693)
);

NAND2xp5_ASAP7_75t_L g1694 ( 
.A(n_1559),
.B(n_1684),
.Y(n_1694)
);

BUFx2_ASAP7_75t_L g1695 ( 
.A(n_1643),
.Y(n_1695)
);

AND2x2_ASAP7_75t_L g1696 ( 
.A(n_1670),
.B(n_1577),
.Y(n_1696)
);

NOR2xp33_ASAP7_75t_L g1697 ( 
.A(n_1569),
.B(n_1591),
.Y(n_1697)
);

HB1xp67_ASAP7_75t_L g1698 ( 
.A(n_1576),
.Y(n_1698)
);

BUFx6f_ASAP7_75t_L g1699 ( 
.A(n_1642),
.Y(n_1699)
);

CKINVDCx5p33_ASAP7_75t_R g1700 ( 
.A(n_1595),
.Y(n_1700)
);

BUFx2_ASAP7_75t_L g1701 ( 
.A(n_1665),
.Y(n_1701)
);

INVx1_ASAP7_75t_L g1702 ( 
.A(n_1586),
.Y(n_1702)
);

OAI22xp5_ASAP7_75t_L g1703 ( 
.A1(n_1673),
.A2(n_1676),
.B1(n_1558),
.B2(n_1556),
.Y(n_1703)
);

INVx1_ASAP7_75t_L g1704 ( 
.A(n_1588),
.Y(n_1704)
);

INVx1_ASAP7_75t_L g1705 ( 
.A(n_1681),
.Y(n_1705)
);

INVx1_ASAP7_75t_L g1706 ( 
.A(n_1587),
.Y(n_1706)
);

BUFx6f_ASAP7_75t_L g1707 ( 
.A(n_1642),
.Y(n_1707)
);

INVx3_ASAP7_75t_L g1708 ( 
.A(n_1669),
.Y(n_1708)
);

INVx1_ASAP7_75t_L g1709 ( 
.A(n_1639),
.Y(n_1709)
);

INVx1_ASAP7_75t_L g1710 ( 
.A(n_1629),
.Y(n_1710)
);

HB1xp67_ASAP7_75t_L g1711 ( 
.A(n_1603),
.Y(n_1711)
);

AO21x2_ASAP7_75t_L g1712 ( 
.A1(n_1628),
.A2(n_1661),
.B(n_1635),
.Y(n_1712)
);

AND2x2_ASAP7_75t_L g1713 ( 
.A(n_1650),
.B(n_1641),
.Y(n_1713)
);

OR2x2_ASAP7_75t_L g1714 ( 
.A(n_1618),
.B(n_1566),
.Y(n_1714)
);

OAI21xp5_ASAP7_75t_L g1715 ( 
.A1(n_1688),
.A2(n_1583),
.B(n_1683),
.Y(n_1715)
);

INVx1_ASAP7_75t_L g1716 ( 
.A(n_1621),
.Y(n_1716)
);

HB1xp67_ASAP7_75t_L g1717 ( 
.A(n_1582),
.Y(n_1717)
);

OR2x2_ASAP7_75t_L g1718 ( 
.A(n_1625),
.B(n_1592),
.Y(n_1718)
);

AND2x2_ASAP7_75t_L g1719 ( 
.A(n_1570),
.B(n_1655),
.Y(n_1719)
);

NOR2xp33_ASAP7_75t_L g1720 ( 
.A(n_1634),
.B(n_1574),
.Y(n_1720)
);

INVx1_ASAP7_75t_L g1721 ( 
.A(n_1609),
.Y(n_1721)
);

NAND4xp25_ASAP7_75t_L g1722 ( 
.A(n_1557),
.B(n_1563),
.C(n_1598),
.D(n_1671),
.Y(n_1722)
);

INVx1_ASAP7_75t_L g1723 ( 
.A(n_1581),
.Y(n_1723)
);

AND2x2_ASAP7_75t_L g1724 ( 
.A(n_1649),
.B(n_1651),
.Y(n_1724)
);

AOI21xp5_ASAP7_75t_SL g1725 ( 
.A1(n_1585),
.A2(n_1563),
.B(n_1633),
.Y(n_1725)
);

INVx2_ASAP7_75t_L g1726 ( 
.A(n_1657),
.Y(n_1726)
);

AND2x2_ASAP7_75t_L g1727 ( 
.A(n_1649),
.B(n_1651),
.Y(n_1727)
);

OA21x2_ASAP7_75t_L g1728 ( 
.A1(n_1580),
.A2(n_1602),
.B(n_1666),
.Y(n_1728)
);

INVx2_ASAP7_75t_L g1729 ( 
.A(n_1619),
.Y(n_1729)
);

INVx2_ASAP7_75t_L g1730 ( 
.A(n_1619),
.Y(n_1730)
);

INVx2_ASAP7_75t_L g1731 ( 
.A(n_1664),
.Y(n_1731)
);

INVx1_ASAP7_75t_L g1732 ( 
.A(n_1581),
.Y(n_1732)
);

INVx2_ASAP7_75t_L g1733 ( 
.A(n_1664),
.Y(n_1733)
);

NAND2xp5_ASAP7_75t_L g1734 ( 
.A(n_1686),
.B(n_1585),
.Y(n_1734)
);

INVx1_ASAP7_75t_L g1735 ( 
.A(n_1572),
.Y(n_1735)
);

BUFx2_ASAP7_75t_L g1736 ( 
.A(n_1648),
.Y(n_1736)
);

INVx1_ASAP7_75t_L g1737 ( 
.A(n_1575),
.Y(n_1737)
);

OR2x2_ASAP7_75t_L g1738 ( 
.A(n_1613),
.B(n_1604),
.Y(n_1738)
);

A2O1A1Ixp33_ASAP7_75t_L g1739 ( 
.A1(n_1593),
.A2(n_1599),
.B(n_1636),
.C(n_1594),
.Y(n_1739)
);

INVx1_ASAP7_75t_L g1740 ( 
.A(n_1575),
.Y(n_1740)
);

OR2x6_ASAP7_75t_L g1741 ( 
.A(n_1596),
.B(n_1597),
.Y(n_1741)
);

OR2x2_ASAP7_75t_L g1742 ( 
.A(n_1652),
.B(n_1653),
.Y(n_1742)
);

OR2x6_ASAP7_75t_L g1743 ( 
.A(n_1637),
.B(n_1636),
.Y(n_1743)
);

INVx1_ASAP7_75t_L g1744 ( 
.A(n_1685),
.Y(n_1744)
);

HB1xp67_ASAP7_75t_L g1745 ( 
.A(n_1590),
.Y(n_1745)
);

AND2x2_ASAP7_75t_L g1746 ( 
.A(n_1652),
.B(n_1653),
.Y(n_1746)
);

CKINVDCx5p33_ASAP7_75t_R g1747 ( 
.A(n_1564),
.Y(n_1747)
);

CKINVDCx5p33_ASAP7_75t_R g1748 ( 
.A(n_1579),
.Y(n_1748)
);

BUFx2_ASAP7_75t_L g1749 ( 
.A(n_1555),
.Y(n_1749)
);

INVx2_ASAP7_75t_L g1750 ( 
.A(n_1656),
.Y(n_1750)
);

INVx1_ASAP7_75t_L g1751 ( 
.A(n_1685),
.Y(n_1751)
);

HB1xp67_ASAP7_75t_L g1752 ( 
.A(n_1617),
.Y(n_1752)
);

OAI21xp5_ASAP7_75t_L g1753 ( 
.A1(n_1580),
.A2(n_1674),
.B(n_1679),
.Y(n_1753)
);

HB1xp67_ASAP7_75t_L g1754 ( 
.A(n_1623),
.Y(n_1754)
);

OAI211xp5_ASAP7_75t_L g1755 ( 
.A1(n_1620),
.A2(n_1567),
.B(n_1667),
.C(n_1626),
.Y(n_1755)
);

OR2x2_ASAP7_75t_L g1756 ( 
.A(n_1658),
.B(n_1659),
.Y(n_1756)
);

INVx1_ASAP7_75t_L g1757 ( 
.A(n_1645),
.Y(n_1757)
);

HB1xp67_ASAP7_75t_L g1758 ( 
.A(n_1612),
.Y(n_1758)
);

OR2x2_ASAP7_75t_L g1759 ( 
.A(n_1660),
.B(n_1562),
.Y(n_1759)
);

INVx2_ASAP7_75t_L g1760 ( 
.A(n_1602),
.Y(n_1760)
);

OR2x6_ASAP7_75t_L g1761 ( 
.A(n_1647),
.B(n_1640),
.Y(n_1761)
);

AND2x4_ASAP7_75t_L g1762 ( 
.A(n_1611),
.B(n_1632),
.Y(n_1762)
);

INVx1_ASAP7_75t_L g1763 ( 
.A(n_1645),
.Y(n_1763)
);

AND2x2_ASAP7_75t_L g1764 ( 
.A(n_1565),
.B(n_1675),
.Y(n_1764)
);

BUFx8_ASAP7_75t_L g1765 ( 
.A(n_1606),
.Y(n_1765)
);

INVx1_ASAP7_75t_L g1766 ( 
.A(n_1646),
.Y(n_1766)
);

INVx1_ASAP7_75t_L g1767 ( 
.A(n_1646),
.Y(n_1767)
);

INVx1_ASAP7_75t_L g1768 ( 
.A(n_1571),
.Y(n_1768)
);

INVx2_ASAP7_75t_L g1769 ( 
.A(n_1573),
.Y(n_1769)
);

HB1xp67_ASAP7_75t_SL g1770 ( 
.A(n_1680),
.Y(n_1770)
);

BUFx2_ASAP7_75t_L g1771 ( 
.A(n_1677),
.Y(n_1771)
);

BUFx3_ASAP7_75t_L g1772 ( 
.A(n_1610),
.Y(n_1772)
);

OAI221xp5_ASAP7_75t_L g1773 ( 
.A1(n_1693),
.A2(n_1624),
.B1(n_1578),
.B2(n_1654),
.C(n_1606),
.Y(n_1773)
);

AND2x2_ASAP7_75t_L g1774 ( 
.A(n_1696),
.B(n_1622),
.Y(n_1774)
);

NAND2xp5_ASAP7_75t_L g1775 ( 
.A(n_1734),
.B(n_1622),
.Y(n_1775)
);

NAND2xp5_ASAP7_75t_L g1776 ( 
.A(n_1706),
.B(n_1668),
.Y(n_1776)
);

INVx2_ASAP7_75t_L g1777 ( 
.A(n_1769),
.Y(n_1777)
);

NAND2x1_ASAP7_75t_L g1778 ( 
.A(n_1725),
.B(n_1677),
.Y(n_1778)
);

NOR2xp33_ASAP7_75t_L g1779 ( 
.A(n_1697),
.B(n_1634),
.Y(n_1779)
);

INVx2_ASAP7_75t_L g1780 ( 
.A(n_1768),
.Y(n_1780)
);

BUFx2_ASAP7_75t_L g1781 ( 
.A(n_1736),
.Y(n_1781)
);

AND2x2_ASAP7_75t_L g1782 ( 
.A(n_1756),
.B(n_1668),
.Y(n_1782)
);

AOI22xp5_ASAP7_75t_L g1783 ( 
.A1(n_1703),
.A2(n_1630),
.B1(n_1615),
.B2(n_1644),
.Y(n_1783)
);

NAND2xp5_ASAP7_75t_L g1784 ( 
.A(n_1706),
.B(n_1600),
.Y(n_1784)
);

AND2x2_ASAP7_75t_L g1785 ( 
.A(n_1756),
.B(n_1663),
.Y(n_1785)
);

INVx2_ASAP7_75t_L g1786 ( 
.A(n_1768),
.Y(n_1786)
);

OR2x2_ASAP7_75t_L g1787 ( 
.A(n_1759),
.B(n_1714),
.Y(n_1787)
);

AND2x2_ASAP7_75t_L g1788 ( 
.A(n_1695),
.B(n_1663),
.Y(n_1788)
);

INVx1_ASAP7_75t_L g1789 ( 
.A(n_1709),
.Y(n_1789)
);

HB1xp67_ASAP7_75t_L g1790 ( 
.A(n_1735),
.Y(n_1790)
);

INVx1_ASAP7_75t_L g1791 ( 
.A(n_1709),
.Y(n_1791)
);

AND2x2_ASAP7_75t_L g1792 ( 
.A(n_1696),
.B(n_1607),
.Y(n_1792)
);

AOI22xp33_ASAP7_75t_L g1793 ( 
.A1(n_1715),
.A2(n_1627),
.B1(n_1638),
.B2(n_1690),
.Y(n_1793)
);

NAND2xp33_ASAP7_75t_R g1794 ( 
.A(n_1700),
.B(n_1560),
.Y(n_1794)
);

BUFx2_ASAP7_75t_L g1795 ( 
.A(n_1736),
.Y(n_1795)
);

AND2x4_ASAP7_75t_L g1796 ( 
.A(n_1699),
.B(n_1560),
.Y(n_1796)
);

AND2x2_ASAP7_75t_L g1797 ( 
.A(n_1713),
.B(n_1695),
.Y(n_1797)
);

OAI21xp5_ASAP7_75t_SL g1798 ( 
.A1(n_1722),
.A2(n_1601),
.B(n_1606),
.Y(n_1798)
);

HB1xp67_ASAP7_75t_L g1799 ( 
.A(n_1735),
.Y(n_1799)
);

BUFx3_ASAP7_75t_L g1800 ( 
.A(n_1749),
.Y(n_1800)
);

INVxp67_ASAP7_75t_L g1801 ( 
.A(n_1711),
.Y(n_1801)
);

AOI221x1_ASAP7_75t_L g1802 ( 
.A1(n_1725),
.A2(n_1614),
.B1(n_1689),
.B2(n_1687),
.C(n_1589),
.Y(n_1802)
);

HB1xp67_ASAP7_75t_L g1803 ( 
.A(n_1737),
.Y(n_1803)
);

INVxp67_ASAP7_75t_L g1804 ( 
.A(n_1710),
.Y(n_1804)
);

INVxp67_ASAP7_75t_L g1805 ( 
.A(n_1710),
.Y(n_1805)
);

AND2x2_ASAP7_75t_L g1806 ( 
.A(n_1713),
.B(n_1605),
.Y(n_1806)
);

A2O1A1Ixp33_ASAP7_75t_L g1807 ( 
.A1(n_1739),
.A2(n_1662),
.B(n_1589),
.C(n_1608),
.Y(n_1807)
);

NOR2x1_ASAP7_75t_L g1808 ( 
.A(n_1755),
.B(n_1616),
.Y(n_1808)
);

BUFx3_ASAP7_75t_L g1809 ( 
.A(n_1749),
.Y(n_1809)
);

AND2x2_ASAP7_75t_L g1810 ( 
.A(n_1699),
.B(n_1707),
.Y(n_1810)
);

NAND3xp33_ASAP7_75t_L g1811 ( 
.A(n_1753),
.B(n_1614),
.C(n_1689),
.Y(n_1811)
);

AOI22xp33_ASAP7_75t_L g1812 ( 
.A1(n_1718),
.A2(n_1608),
.B1(n_1682),
.B2(n_1672),
.Y(n_1812)
);

AND2x2_ASAP7_75t_L g1813 ( 
.A(n_1719),
.B(n_1758),
.Y(n_1813)
);

AND2x2_ASAP7_75t_L g1814 ( 
.A(n_1707),
.B(n_1672),
.Y(n_1814)
);

AND2x4_ASAP7_75t_L g1815 ( 
.A(n_1707),
.B(n_1614),
.Y(n_1815)
);

OR2x2_ASAP7_75t_L g1816 ( 
.A(n_1775),
.B(n_1692),
.Y(n_1816)
);

INVxp67_ASAP7_75t_L g1817 ( 
.A(n_1808),
.Y(n_1817)
);

OAI22xp5_ASAP7_75t_L g1818 ( 
.A1(n_1808),
.A2(n_1738),
.B1(n_1761),
.B2(n_1631),
.Y(n_1818)
);

OAI321xp33_ASAP7_75t_L g1819 ( 
.A1(n_1773),
.A2(n_1807),
.A3(n_1775),
.B1(n_1811),
.B2(n_1788),
.C(n_1761),
.Y(n_1819)
);

AOI221xp5_ASAP7_75t_L g1820 ( 
.A1(n_1785),
.A2(n_1701),
.B1(n_1694),
.B2(n_1760),
.C(n_1702),
.Y(n_1820)
);

NOR2xp33_ASAP7_75t_R g1821 ( 
.A(n_1794),
.B(n_1747),
.Y(n_1821)
);

OAI31xp33_ASAP7_75t_L g1822 ( 
.A1(n_1773),
.A2(n_1701),
.A3(n_1738),
.B(n_1716),
.Y(n_1822)
);

AOI22xp33_ASAP7_75t_L g1823 ( 
.A1(n_1811),
.A2(n_1718),
.B1(n_1714),
.B2(n_1750),
.Y(n_1823)
);

BUFx2_ASAP7_75t_L g1824 ( 
.A(n_1781),
.Y(n_1824)
);

INVx1_ASAP7_75t_L g1825 ( 
.A(n_1790),
.Y(n_1825)
);

OAI33xp33_ASAP7_75t_L g1826 ( 
.A1(n_1801),
.A2(n_1705),
.A3(n_1704),
.B1(n_1716),
.B2(n_1742),
.B3(n_1732),
.Y(n_1826)
);

INVx1_ASAP7_75t_L g1827 ( 
.A(n_1790),
.Y(n_1827)
);

NOR2x1_ASAP7_75t_SL g1828 ( 
.A(n_1800),
.B(n_1741),
.Y(n_1828)
);

NOR2xp33_ASAP7_75t_L g1829 ( 
.A(n_1779),
.B(n_1770),
.Y(n_1829)
);

INVx2_ASAP7_75t_SL g1830 ( 
.A(n_1800),
.Y(n_1830)
);

OR2x2_ASAP7_75t_L g1831 ( 
.A(n_1781),
.B(n_1698),
.Y(n_1831)
);

NOR2xp33_ASAP7_75t_R g1832 ( 
.A(n_1795),
.B(n_1747),
.Y(n_1832)
);

BUFx6f_ASAP7_75t_L g1833 ( 
.A(n_1778),
.Y(n_1833)
);

BUFx12f_ASAP7_75t_L g1834 ( 
.A(n_1795),
.Y(n_1834)
);

INVx1_ASAP7_75t_L g1835 ( 
.A(n_1799),
.Y(n_1835)
);

AOI22xp33_ASAP7_75t_L g1836 ( 
.A1(n_1785),
.A2(n_1750),
.B1(n_1743),
.B2(n_1761),
.Y(n_1836)
);

BUFx3_ASAP7_75t_L g1837 ( 
.A(n_1815),
.Y(n_1837)
);

OAI21xp5_ASAP7_75t_L g1838 ( 
.A1(n_1802),
.A2(n_1752),
.B(n_1760),
.Y(n_1838)
);

NAND2xp5_ASAP7_75t_SL g1839 ( 
.A(n_1801),
.B(n_1708),
.Y(n_1839)
);

INVx1_ASAP7_75t_L g1840 ( 
.A(n_1799),
.Y(n_1840)
);

INVx1_ASAP7_75t_L g1841 ( 
.A(n_1803),
.Y(n_1841)
);

OAI21xp5_ASAP7_75t_L g1842 ( 
.A1(n_1802),
.A2(n_1745),
.B(n_1723),
.Y(n_1842)
);

INVx2_ASAP7_75t_L g1843 ( 
.A(n_1777),
.Y(n_1843)
);

HB1xp67_ASAP7_75t_L g1844 ( 
.A(n_1803),
.Y(n_1844)
);

INVx1_ASAP7_75t_L g1845 ( 
.A(n_1789),
.Y(n_1845)
);

BUFx2_ASAP7_75t_L g1846 ( 
.A(n_1809),
.Y(n_1846)
);

AOI211xp5_ASAP7_75t_L g1847 ( 
.A1(n_1798),
.A2(n_1746),
.B(n_1724),
.C(n_1727),
.Y(n_1847)
);

NAND3xp33_ASAP7_75t_SL g1848 ( 
.A(n_1783),
.B(n_1748),
.C(n_1720),
.Y(n_1848)
);

AOI33xp33_ASAP7_75t_L g1849 ( 
.A1(n_1785),
.A2(n_1704),
.A3(n_1705),
.B1(n_1764),
.B2(n_1740),
.B3(n_1744),
.Y(n_1849)
);

NAND2xp5_ASAP7_75t_L g1850 ( 
.A(n_1804),
.B(n_1717),
.Y(n_1850)
);

OAI221xp5_ASAP7_75t_L g1851 ( 
.A1(n_1783),
.A2(n_1743),
.B1(n_1708),
.B2(n_1731),
.C(n_1733),
.Y(n_1851)
);

AOI22xp33_ASAP7_75t_L g1852 ( 
.A1(n_1812),
.A2(n_1743),
.B1(n_1757),
.B2(n_1763),
.Y(n_1852)
);

INVx4_ASAP7_75t_L g1853 ( 
.A(n_1815),
.Y(n_1853)
);

AOI22xp33_ASAP7_75t_L g1854 ( 
.A1(n_1787),
.A2(n_1743),
.B1(n_1757),
.B2(n_1763),
.Y(n_1854)
);

OAI33xp33_ASAP7_75t_L g1855 ( 
.A1(n_1804),
.A2(n_1742),
.A3(n_1732),
.B1(n_1723),
.B2(n_1740),
.B3(n_1744),
.Y(n_1855)
);

NAND2xp33_ASAP7_75t_R g1856 ( 
.A(n_1788),
.B(n_1748),
.Y(n_1856)
);

INVx2_ASAP7_75t_L g1857 ( 
.A(n_1780),
.Y(n_1857)
);

INVx1_ASAP7_75t_L g1858 ( 
.A(n_1789),
.Y(n_1858)
);

AOI22xp33_ASAP7_75t_SL g1859 ( 
.A1(n_1788),
.A2(n_1712),
.B1(n_1767),
.B2(n_1766),
.Y(n_1859)
);

NAND2xp5_ASAP7_75t_L g1860 ( 
.A(n_1805),
.B(n_1764),
.Y(n_1860)
);

AND2x2_ASAP7_75t_L g1861 ( 
.A(n_1797),
.B(n_1754),
.Y(n_1861)
);

OAI221xp5_ASAP7_75t_L g1862 ( 
.A1(n_1793),
.A2(n_1708),
.B1(n_1733),
.B2(n_1731),
.C(n_1767),
.Y(n_1862)
);

HB1xp67_ASAP7_75t_L g1863 ( 
.A(n_1805),
.Y(n_1863)
);

OAI31xp33_ASAP7_75t_L g1864 ( 
.A1(n_1782),
.A2(n_1766),
.A3(n_1724),
.B(n_1727),
.Y(n_1864)
);

AOI221xp5_ASAP7_75t_L g1865 ( 
.A1(n_1782),
.A2(n_1746),
.B1(n_1751),
.B2(n_1712),
.C(n_1729),
.Y(n_1865)
);

AND2x2_ASAP7_75t_L g1866 ( 
.A(n_1797),
.B(n_1772),
.Y(n_1866)
);

AND2x4_ASAP7_75t_L g1867 ( 
.A(n_1796),
.B(n_1762),
.Y(n_1867)
);

NOR4xp25_ASAP7_75t_SL g1868 ( 
.A(n_1798),
.B(n_1700),
.C(n_1751),
.D(n_1771),
.Y(n_1868)
);

AOI211xp5_ASAP7_75t_L g1869 ( 
.A1(n_1782),
.A2(n_1707),
.B(n_1729),
.C(n_1730),
.Y(n_1869)
);

AOI22xp33_ASAP7_75t_L g1870 ( 
.A1(n_1787),
.A2(n_1712),
.B1(n_1726),
.B2(n_1721),
.Y(n_1870)
);

CKINVDCx16_ASAP7_75t_R g1871 ( 
.A(n_1821),
.Y(n_1871)
);

INVx2_ASAP7_75t_L g1872 ( 
.A(n_1857),
.Y(n_1872)
);

INVx3_ASAP7_75t_L g1873 ( 
.A(n_1833),
.Y(n_1873)
);

INVx1_ASAP7_75t_L g1874 ( 
.A(n_1845),
.Y(n_1874)
);

INVx1_ASAP7_75t_L g1875 ( 
.A(n_1845),
.Y(n_1875)
);

NAND3xp33_ASAP7_75t_SL g1876 ( 
.A(n_1868),
.B(n_1778),
.C(n_1813),
.Y(n_1876)
);

INVx3_ASAP7_75t_L g1877 ( 
.A(n_1833),
.Y(n_1877)
);

AND2x2_ASAP7_75t_L g1878 ( 
.A(n_1847),
.B(n_1774),
.Y(n_1878)
);

INVx1_ASAP7_75t_L g1879 ( 
.A(n_1858),
.Y(n_1879)
);

AND2x2_ASAP7_75t_L g1880 ( 
.A(n_1847),
.B(n_1774),
.Y(n_1880)
);

AND2x2_ASAP7_75t_L g1881 ( 
.A(n_1864),
.B(n_1792),
.Y(n_1881)
);

AND2x2_ASAP7_75t_L g1882 ( 
.A(n_1846),
.B(n_1792),
.Y(n_1882)
);

OR2x6_ASAP7_75t_L g1883 ( 
.A(n_1833),
.B(n_1741),
.Y(n_1883)
);

BUFx6f_ASAP7_75t_L g1884 ( 
.A(n_1833),
.Y(n_1884)
);

INVxp67_ASAP7_75t_SL g1885 ( 
.A(n_1863),
.Y(n_1885)
);

INVx1_ASAP7_75t_L g1886 ( 
.A(n_1858),
.Y(n_1886)
);

INVx1_ASAP7_75t_L g1887 ( 
.A(n_1825),
.Y(n_1887)
);

INVx1_ASAP7_75t_L g1888 ( 
.A(n_1825),
.Y(n_1888)
);

INVx4_ASAP7_75t_SL g1889 ( 
.A(n_1867),
.Y(n_1889)
);

INVx2_ASAP7_75t_L g1890 ( 
.A(n_1843),
.Y(n_1890)
);

BUFx6f_ASAP7_75t_L g1891 ( 
.A(n_1837),
.Y(n_1891)
);

OR2x2_ASAP7_75t_L g1892 ( 
.A(n_1816),
.B(n_1776),
.Y(n_1892)
);

NAND2xp5_ASAP7_75t_L g1893 ( 
.A(n_1865),
.B(n_1776),
.Y(n_1893)
);

NOR3xp33_ASAP7_75t_SL g1894 ( 
.A(n_1856),
.B(n_1784),
.C(n_1791),
.Y(n_1894)
);

INVx1_ASAP7_75t_L g1895 ( 
.A(n_1827),
.Y(n_1895)
);

AOI21xp5_ASAP7_75t_SL g1896 ( 
.A1(n_1828),
.A2(n_1728),
.B(n_1815),
.Y(n_1896)
);

OA21x2_ASAP7_75t_L g1897 ( 
.A1(n_1838),
.A2(n_1784),
.B(n_1786),
.Y(n_1897)
);

BUFx3_ASAP7_75t_L g1898 ( 
.A(n_1846),
.Y(n_1898)
);

INVx3_ASAP7_75t_L g1899 ( 
.A(n_1853),
.Y(n_1899)
);

INVx1_ASAP7_75t_L g1900 ( 
.A(n_1827),
.Y(n_1900)
);

INVx1_ASAP7_75t_L g1901 ( 
.A(n_1835),
.Y(n_1901)
);

INVx1_ASAP7_75t_L g1902 ( 
.A(n_1835),
.Y(n_1902)
);

AND2x2_ASAP7_75t_L g1903 ( 
.A(n_1866),
.B(n_1806),
.Y(n_1903)
);

OA21x2_ASAP7_75t_L g1904 ( 
.A1(n_1842),
.A2(n_1786),
.B(n_1780),
.Y(n_1904)
);

AND4x1_ASAP7_75t_L g1905 ( 
.A(n_1822),
.B(n_1810),
.C(n_1765),
.D(n_1814),
.Y(n_1905)
);

NOR2xp33_ASAP7_75t_L g1906 ( 
.A(n_1848),
.B(n_1806),
.Y(n_1906)
);

INVx1_ASAP7_75t_L g1907 ( 
.A(n_1840),
.Y(n_1907)
);

INVx1_ASAP7_75t_L g1908 ( 
.A(n_1874),
.Y(n_1908)
);

AND2x2_ASAP7_75t_L g1909 ( 
.A(n_1894),
.B(n_1824),
.Y(n_1909)
);

BUFx2_ASAP7_75t_L g1910 ( 
.A(n_1871),
.Y(n_1910)
);

OR2x2_ASAP7_75t_L g1911 ( 
.A(n_1893),
.B(n_1816),
.Y(n_1911)
);

INVx1_ASAP7_75t_L g1912 ( 
.A(n_1874),
.Y(n_1912)
);

INVx1_ASAP7_75t_L g1913 ( 
.A(n_1874),
.Y(n_1913)
);

INVx2_ASAP7_75t_L g1914 ( 
.A(n_1890),
.Y(n_1914)
);

INVx2_ASAP7_75t_L g1915 ( 
.A(n_1890),
.Y(n_1915)
);

AND2x4_ASAP7_75t_L g1916 ( 
.A(n_1889),
.B(n_1828),
.Y(n_1916)
);

AND2x4_ASAP7_75t_L g1917 ( 
.A(n_1889),
.B(n_1898),
.Y(n_1917)
);

INVx1_ASAP7_75t_L g1918 ( 
.A(n_1875),
.Y(n_1918)
);

NAND2xp5_ASAP7_75t_L g1919 ( 
.A(n_1885),
.B(n_1849),
.Y(n_1919)
);

NAND2xp33_ASAP7_75t_SL g1920 ( 
.A(n_1894),
.B(n_1832),
.Y(n_1920)
);

INVx2_ASAP7_75t_L g1921 ( 
.A(n_1890),
.Y(n_1921)
);

NAND4xp25_ASAP7_75t_L g1922 ( 
.A(n_1898),
.B(n_1820),
.C(n_1818),
.D(n_1839),
.Y(n_1922)
);

NAND2xp5_ASAP7_75t_L g1923 ( 
.A(n_1885),
.B(n_1860),
.Y(n_1923)
);

BUFx2_ASAP7_75t_SL g1924 ( 
.A(n_1884),
.Y(n_1924)
);

HB1xp67_ASAP7_75t_L g1925 ( 
.A(n_1887),
.Y(n_1925)
);

AOI22xp33_ASAP7_75t_L g1926 ( 
.A1(n_1893),
.A2(n_1859),
.B1(n_1897),
.B2(n_1904),
.Y(n_1926)
);

INVx1_ASAP7_75t_L g1927 ( 
.A(n_1875),
.Y(n_1927)
);

OAI31xp33_ASAP7_75t_L g1928 ( 
.A1(n_1893),
.A2(n_1817),
.A3(n_1862),
.B(n_1851),
.Y(n_1928)
);

INVx1_ASAP7_75t_L g1929 ( 
.A(n_1875),
.Y(n_1929)
);

AND2x2_ASAP7_75t_L g1930 ( 
.A(n_1889),
.B(n_1824),
.Y(n_1930)
);

OR2x2_ASAP7_75t_L g1931 ( 
.A(n_1892),
.B(n_1831),
.Y(n_1931)
);

INVx2_ASAP7_75t_L g1932 ( 
.A(n_1890),
.Y(n_1932)
);

NAND2xp5_ASAP7_75t_L g1933 ( 
.A(n_1882),
.B(n_1850),
.Y(n_1933)
);

AOI31xp33_ASAP7_75t_SL g1934 ( 
.A1(n_1906),
.A2(n_1829),
.A3(n_1869),
.B(n_1831),
.Y(n_1934)
);

INVx2_ASAP7_75t_L g1935 ( 
.A(n_1890),
.Y(n_1935)
);

INVx1_ASAP7_75t_L g1936 ( 
.A(n_1879),
.Y(n_1936)
);

INVx2_ASAP7_75t_L g1937 ( 
.A(n_1872),
.Y(n_1937)
);

NAND3xp33_ASAP7_75t_L g1938 ( 
.A(n_1897),
.B(n_1869),
.C(n_1854),
.Y(n_1938)
);

NAND2xp5_ASAP7_75t_L g1939 ( 
.A(n_1882),
.B(n_1844),
.Y(n_1939)
);

NOR2xp33_ASAP7_75t_R g1940 ( 
.A(n_1871),
.B(n_1834),
.Y(n_1940)
);

NOR2x1_ASAP7_75t_L g1941 ( 
.A(n_1898),
.B(n_1853),
.Y(n_1941)
);

INVx1_ASAP7_75t_L g1942 ( 
.A(n_1879),
.Y(n_1942)
);

AND2x2_ASAP7_75t_L g1943 ( 
.A(n_1889),
.B(n_1866),
.Y(n_1943)
);

OR2x2_ASAP7_75t_L g1944 ( 
.A(n_1892),
.B(n_1840),
.Y(n_1944)
);

NAND2xp5_ASAP7_75t_L g1945 ( 
.A(n_1882),
.B(n_1841),
.Y(n_1945)
);

INVx1_ASAP7_75t_L g1946 ( 
.A(n_1879),
.Y(n_1946)
);

OR2x2_ASAP7_75t_L g1947 ( 
.A(n_1892),
.B(n_1841),
.Y(n_1947)
);

INVx1_ASAP7_75t_L g1948 ( 
.A(n_1886),
.Y(n_1948)
);

NOR2xp33_ASAP7_75t_L g1949 ( 
.A(n_1871),
.B(n_1834),
.Y(n_1949)
);

OR2x2_ASAP7_75t_L g1950 ( 
.A(n_1892),
.B(n_1791),
.Y(n_1950)
);

HB1xp67_ASAP7_75t_L g1951 ( 
.A(n_1887),
.Y(n_1951)
);

INVx1_ASAP7_75t_L g1952 ( 
.A(n_1886),
.Y(n_1952)
);

NAND2xp5_ASAP7_75t_L g1953 ( 
.A(n_1882),
.B(n_1823),
.Y(n_1953)
);

NAND2xp5_ASAP7_75t_L g1954 ( 
.A(n_1903),
.B(n_1861),
.Y(n_1954)
);

NAND2x1p5_ASAP7_75t_L g1955 ( 
.A(n_1916),
.B(n_1905),
.Y(n_1955)
);

AOI22xp5_ASAP7_75t_L g1956 ( 
.A1(n_1926),
.A2(n_1897),
.B1(n_1904),
.B2(n_1878),
.Y(n_1956)
);

AND2x2_ASAP7_75t_L g1957 ( 
.A(n_1910),
.B(n_1878),
.Y(n_1957)
);

NAND2xp5_ASAP7_75t_L g1958 ( 
.A(n_1911),
.B(n_1881),
.Y(n_1958)
);

INVx1_ASAP7_75t_SL g1959 ( 
.A(n_1910),
.Y(n_1959)
);

INVx1_ASAP7_75t_L g1960 ( 
.A(n_1925),
.Y(n_1960)
);

INVx2_ASAP7_75t_L g1961 ( 
.A(n_1914),
.Y(n_1961)
);

INVx1_ASAP7_75t_L g1962 ( 
.A(n_1951),
.Y(n_1962)
);

OR2x2_ASAP7_75t_L g1963 ( 
.A(n_1911),
.B(n_1887),
.Y(n_1963)
);

OR2x2_ASAP7_75t_L g1964 ( 
.A(n_1931),
.B(n_1888),
.Y(n_1964)
);

OAI31xp33_ASAP7_75t_L g1965 ( 
.A1(n_1938),
.A2(n_1880),
.A3(n_1878),
.B(n_1906),
.Y(n_1965)
);

NAND2xp5_ASAP7_75t_L g1966 ( 
.A(n_1919),
.B(n_1881),
.Y(n_1966)
);

INVx1_ASAP7_75t_L g1967 ( 
.A(n_1908),
.Y(n_1967)
);

INVxp67_ASAP7_75t_L g1968 ( 
.A(n_1949),
.Y(n_1968)
);

NAND2xp5_ASAP7_75t_L g1969 ( 
.A(n_1954),
.B(n_1881),
.Y(n_1969)
);

INVx1_ASAP7_75t_L g1970 ( 
.A(n_1908),
.Y(n_1970)
);

INVx1_ASAP7_75t_L g1971 ( 
.A(n_1912),
.Y(n_1971)
);

AND2x2_ASAP7_75t_L g1972 ( 
.A(n_1917),
.B(n_1878),
.Y(n_1972)
);

INVx1_ASAP7_75t_L g1973 ( 
.A(n_1912),
.Y(n_1973)
);

OR2x2_ASAP7_75t_L g1974 ( 
.A(n_1931),
.B(n_1923),
.Y(n_1974)
);

NAND2xp5_ASAP7_75t_L g1975 ( 
.A(n_1933),
.B(n_1881),
.Y(n_1975)
);

OR2x2_ASAP7_75t_L g1976 ( 
.A(n_1953),
.B(n_1888),
.Y(n_1976)
);

AND2x2_ASAP7_75t_L g1977 ( 
.A(n_1917),
.B(n_1880),
.Y(n_1977)
);

AND2x2_ASAP7_75t_L g1978 ( 
.A(n_1917),
.B(n_1880),
.Y(n_1978)
);

NOR2xp33_ASAP7_75t_L g1979 ( 
.A(n_1922),
.B(n_1855),
.Y(n_1979)
);

O2A1O1Ixp5_ASAP7_75t_L g1980 ( 
.A1(n_1920),
.A2(n_1826),
.B(n_1880),
.C(n_1873),
.Y(n_1980)
);

INVx1_ASAP7_75t_L g1981 ( 
.A(n_1918),
.Y(n_1981)
);

OR2x2_ASAP7_75t_L g1982 ( 
.A(n_1945),
.B(n_1888),
.Y(n_1982)
);

OAI21xp33_ASAP7_75t_L g1983 ( 
.A1(n_1909),
.A2(n_1898),
.B(n_1876),
.Y(n_1983)
);

INVx2_ASAP7_75t_L g1984 ( 
.A(n_1914),
.Y(n_1984)
);

INVx1_ASAP7_75t_L g1985 ( 
.A(n_1918),
.Y(n_1985)
);

AOI22xp5_ASAP7_75t_L g1986 ( 
.A1(n_1920),
.A2(n_1897),
.B1(n_1904),
.B2(n_1852),
.Y(n_1986)
);

AOI21xp33_ASAP7_75t_L g1987 ( 
.A1(n_1928),
.A2(n_1819),
.B(n_1897),
.Y(n_1987)
);

AND2x2_ASAP7_75t_L g1988 ( 
.A(n_1943),
.B(n_1889),
.Y(n_1988)
);

OR2x2_ASAP7_75t_L g1989 ( 
.A(n_1939),
.B(n_1895),
.Y(n_1989)
);

NAND2xp5_ASAP7_75t_L g1990 ( 
.A(n_1950),
.B(n_1903),
.Y(n_1990)
);

AOI22xp5_ASAP7_75t_L g1991 ( 
.A1(n_1909),
.A2(n_1897),
.B1(n_1904),
.B2(n_1870),
.Y(n_1991)
);

OAI22xp5_ASAP7_75t_L g1992 ( 
.A1(n_1934),
.A2(n_1836),
.B1(n_1903),
.B2(n_1896),
.Y(n_1992)
);

AND2x2_ASAP7_75t_L g1993 ( 
.A(n_1943),
.B(n_1889),
.Y(n_1993)
);

INVx1_ASAP7_75t_L g1994 ( 
.A(n_1967),
.Y(n_1994)
);

NAND2xp5_ASAP7_75t_L g1995 ( 
.A(n_1979),
.B(n_1913),
.Y(n_1995)
);

INVx1_ASAP7_75t_SL g1996 ( 
.A(n_1959),
.Y(n_1996)
);

INVx2_ASAP7_75t_SL g1997 ( 
.A(n_1972),
.Y(n_1997)
);

NAND2xp5_ASAP7_75t_L g1998 ( 
.A(n_1979),
.B(n_1927),
.Y(n_1998)
);

INVx2_ASAP7_75t_L g1999 ( 
.A(n_1972),
.Y(n_1999)
);

OR2x2_ASAP7_75t_L g2000 ( 
.A(n_1958),
.B(n_1944),
.Y(n_2000)
);

OR2x2_ASAP7_75t_L g2001 ( 
.A(n_1974),
.B(n_1944),
.Y(n_2001)
);

INVx1_ASAP7_75t_L g2002 ( 
.A(n_1970),
.Y(n_2002)
);

AND2x4_ASAP7_75t_L g2003 ( 
.A(n_1968),
.B(n_1889),
.Y(n_2003)
);

OR2x6_ASAP7_75t_L g2004 ( 
.A(n_1968),
.B(n_1896),
.Y(n_2004)
);

INVx1_ASAP7_75t_SL g2005 ( 
.A(n_1957),
.Y(n_2005)
);

INVx1_ASAP7_75t_L g2006 ( 
.A(n_1971),
.Y(n_2006)
);

NAND2xp5_ASAP7_75t_L g2007 ( 
.A(n_1956),
.B(n_1929),
.Y(n_2007)
);

OR2x2_ASAP7_75t_L g2008 ( 
.A(n_1976),
.B(n_1947),
.Y(n_2008)
);

AND2x2_ASAP7_75t_L g2009 ( 
.A(n_1957),
.B(n_1940),
.Y(n_2009)
);

OR2x2_ASAP7_75t_L g2010 ( 
.A(n_1966),
.B(n_1947),
.Y(n_2010)
);

INVx1_ASAP7_75t_L g2011 ( 
.A(n_1973),
.Y(n_2011)
);

NAND2xp5_ASAP7_75t_SL g2012 ( 
.A(n_1980),
.B(n_1916),
.Y(n_2012)
);

INVx1_ASAP7_75t_SL g2013 ( 
.A(n_1960),
.Y(n_2013)
);

INVx1_ASAP7_75t_L g2014 ( 
.A(n_1981),
.Y(n_2014)
);

INVx1_ASAP7_75t_L g2015 ( 
.A(n_1985),
.Y(n_2015)
);

NOR2x1_ASAP7_75t_L g2016 ( 
.A(n_1962),
.B(n_1941),
.Y(n_2016)
);

OR2x2_ASAP7_75t_L g2017 ( 
.A(n_1975),
.B(n_1950),
.Y(n_2017)
);

NAND2xp33_ASAP7_75t_L g2018 ( 
.A(n_1983),
.B(n_1955),
.Y(n_2018)
);

INVx1_ASAP7_75t_L g2019 ( 
.A(n_1964),
.Y(n_2019)
);

OR2x2_ASAP7_75t_L g2020 ( 
.A(n_1990),
.B(n_1942),
.Y(n_2020)
);

INVx1_ASAP7_75t_L g2021 ( 
.A(n_1963),
.Y(n_2021)
);

INVx2_ASAP7_75t_L g2022 ( 
.A(n_1977),
.Y(n_2022)
);

NAND2xp5_ASAP7_75t_L g2023 ( 
.A(n_2005),
.B(n_1965),
.Y(n_2023)
);

AOI31xp33_ASAP7_75t_L g2024 ( 
.A1(n_1996),
.A2(n_1955),
.A3(n_1987),
.B(n_1977),
.Y(n_2024)
);

AND2x2_ASAP7_75t_L g2025 ( 
.A(n_2009),
.B(n_1978),
.Y(n_2025)
);

OR2x2_ASAP7_75t_L g2026 ( 
.A(n_2005),
.B(n_1969),
.Y(n_2026)
);

INVx1_ASAP7_75t_L g2027 ( 
.A(n_2001),
.Y(n_2027)
);

INVx1_ASAP7_75t_L g2028 ( 
.A(n_1994),
.Y(n_2028)
);

OAI221xp5_ASAP7_75t_L g2029 ( 
.A1(n_1995),
.A2(n_1991),
.B1(n_1986),
.B2(n_1980),
.C(n_1992),
.Y(n_2029)
);

OAI22xp33_ASAP7_75t_L g2030 ( 
.A1(n_2004),
.A2(n_1897),
.B1(n_1904),
.B2(n_1876),
.Y(n_2030)
);

NOR2x1_ASAP7_75t_L g2031 ( 
.A(n_1996),
.B(n_1898),
.Y(n_2031)
);

AOI21xp5_ASAP7_75t_L g2032 ( 
.A1(n_2012),
.A2(n_1876),
.B(n_1978),
.Y(n_2032)
);

NAND2xp5_ASAP7_75t_L g2033 ( 
.A(n_2013),
.B(n_1989),
.Y(n_2033)
);

INVx1_ASAP7_75t_L g2034 ( 
.A(n_2002),
.Y(n_2034)
);

NAND2xp5_ASAP7_75t_L g2035 ( 
.A(n_2013),
.B(n_1982),
.Y(n_2035)
);

AOI22xp33_ASAP7_75t_L g2036 ( 
.A1(n_1995),
.A2(n_1998),
.B1(n_2007),
.B2(n_2004),
.Y(n_2036)
);

INVx1_ASAP7_75t_SL g2037 ( 
.A(n_2018),
.Y(n_2037)
);

OAI22xp5_ASAP7_75t_L g2038 ( 
.A1(n_2004),
.A2(n_1993),
.B1(n_1988),
.B2(n_1916),
.Y(n_2038)
);

AOI211x1_ASAP7_75t_L g2039 ( 
.A1(n_1998),
.A2(n_1905),
.B(n_1930),
.C(n_1993),
.Y(n_2039)
);

INVx1_ASAP7_75t_L g2040 ( 
.A(n_2006),
.Y(n_2040)
);

NAND2xp5_ASAP7_75t_L g2041 ( 
.A(n_2021),
.B(n_1961),
.Y(n_2041)
);

OAI211xp5_ASAP7_75t_L g2042 ( 
.A1(n_2007),
.A2(n_1988),
.B(n_1930),
.C(n_1884),
.Y(n_2042)
);

AOI21xp33_ASAP7_75t_L g2043 ( 
.A1(n_2011),
.A2(n_1984),
.B(n_1961),
.Y(n_2043)
);

NAND2xp5_ASAP7_75t_L g2044 ( 
.A(n_2019),
.B(n_1984),
.Y(n_2044)
);

OAI21xp5_ASAP7_75t_L g2045 ( 
.A1(n_2016),
.A2(n_1904),
.B(n_1905),
.Y(n_2045)
);

NOR2xp33_ASAP7_75t_L g2046 ( 
.A(n_2037),
.B(n_1997),
.Y(n_2046)
);

AND2x2_ASAP7_75t_L g2047 ( 
.A(n_2025),
.B(n_1999),
.Y(n_2047)
);

NAND2xp5_ASAP7_75t_L g2048 ( 
.A(n_2031),
.B(n_2022),
.Y(n_2048)
);

NAND2xp5_ASAP7_75t_L g2049 ( 
.A(n_2036),
.B(n_2008),
.Y(n_2049)
);

NAND2xp5_ASAP7_75t_L g2050 ( 
.A(n_2036),
.B(n_2010),
.Y(n_2050)
);

INVx1_ASAP7_75t_L g2051 ( 
.A(n_2027),
.Y(n_2051)
);

HB1xp67_ASAP7_75t_L g2052 ( 
.A(n_2025),
.Y(n_2052)
);

NAND2xp5_ASAP7_75t_L g2053 ( 
.A(n_2033),
.B(n_2000),
.Y(n_2053)
);

NOR2x1p5_ASAP7_75t_L g2054 ( 
.A(n_2026),
.B(n_2035),
.Y(n_2054)
);

AND2x2_ASAP7_75t_L g2055 ( 
.A(n_2032),
.B(n_2003),
.Y(n_2055)
);

INVx1_ASAP7_75t_L g2056 ( 
.A(n_2041),
.Y(n_2056)
);

NAND2xp5_ASAP7_75t_L g2057 ( 
.A(n_2044),
.B(n_2017),
.Y(n_2057)
);

AND2x2_ASAP7_75t_L g2058 ( 
.A(n_2038),
.B(n_2003),
.Y(n_2058)
);

INVx1_ASAP7_75t_L g2059 ( 
.A(n_2028),
.Y(n_2059)
);

AND2x2_ASAP7_75t_L g2060 ( 
.A(n_2023),
.B(n_2020),
.Y(n_2060)
);

AND2x2_ASAP7_75t_L g2061 ( 
.A(n_2034),
.B(n_2014),
.Y(n_2061)
);

AOI221xp5_ASAP7_75t_L g2062 ( 
.A1(n_2049),
.A2(n_2029),
.B1(n_2024),
.B2(n_2030),
.C(n_2043),
.Y(n_2062)
);

OAI221xp5_ASAP7_75t_SL g2063 ( 
.A1(n_2050),
.A2(n_2030),
.B1(n_2042),
.B2(n_2040),
.C(n_2045),
.Y(n_2063)
);

NOR4xp25_ASAP7_75t_L g2064 ( 
.A(n_2051),
.B(n_2015),
.C(n_1915),
.D(n_1921),
.Y(n_2064)
);

NAND4xp25_ASAP7_75t_SL g2065 ( 
.A(n_2055),
.B(n_2047),
.C(n_2053),
.D(n_2057),
.Y(n_2065)
);

OR2x2_ASAP7_75t_L g2066 ( 
.A(n_2052),
.B(n_1946),
.Y(n_2066)
);

AOI32xp33_ASAP7_75t_L g2067 ( 
.A1(n_2060),
.A2(n_2039),
.A3(n_1915),
.B1(n_1921),
.B2(n_1932),
.Y(n_2067)
);

HB1xp67_ASAP7_75t_L g2068 ( 
.A(n_2047),
.Y(n_2068)
);

AOI322xp5_ASAP7_75t_L g2069 ( 
.A1(n_2060),
.A2(n_1935),
.A3(n_1932),
.B1(n_1937),
.B2(n_1936),
.C1(n_1952),
.C2(n_1948),
.Y(n_2069)
);

AOI221xp5_ASAP7_75t_L g2070 ( 
.A1(n_2056),
.A2(n_1935),
.B1(n_1937),
.B2(n_1952),
.C(n_1936),
.Y(n_2070)
);

NOR2xp67_ASAP7_75t_L g2071 ( 
.A(n_2046),
.B(n_1873),
.Y(n_2071)
);

AOI211xp5_ASAP7_75t_L g2072 ( 
.A1(n_2055),
.A2(n_1884),
.B(n_1948),
.C(n_1873),
.Y(n_2072)
);

AOI21xp33_ASAP7_75t_L g2073 ( 
.A1(n_2048),
.A2(n_1904),
.B(n_1924),
.Y(n_2073)
);

AOI22xp5_ASAP7_75t_L g2074 ( 
.A1(n_2054),
.A2(n_1884),
.B1(n_1924),
.B2(n_1873),
.Y(n_2074)
);

NOR3xp33_ASAP7_75t_L g2075 ( 
.A(n_2051),
.B(n_1873),
.C(n_1877),
.Y(n_2075)
);

INVx1_ASAP7_75t_L g2076 ( 
.A(n_2061),
.Y(n_2076)
);

AOI21xp33_ASAP7_75t_L g2077 ( 
.A1(n_2062),
.A2(n_2059),
.B(n_2061),
.Y(n_2077)
);

AOI211xp5_ASAP7_75t_L g2078 ( 
.A1(n_2063),
.A2(n_2058),
.B(n_1884),
.C(n_1873),
.Y(n_2078)
);

NAND3xp33_ASAP7_75t_L g2079 ( 
.A(n_2068),
.B(n_2076),
.C(n_2072),
.Y(n_2079)
);

INVx3_ASAP7_75t_L g2080 ( 
.A(n_2066),
.Y(n_2080)
);

INVxp67_ASAP7_75t_SL g2081 ( 
.A(n_2071),
.Y(n_2081)
);

INVx1_ASAP7_75t_L g2082 ( 
.A(n_2065),
.Y(n_2082)
);

INVx1_ASAP7_75t_L g2083 ( 
.A(n_2064),
.Y(n_2083)
);

AOI221xp5_ASAP7_75t_L g2084 ( 
.A1(n_2067),
.A2(n_2058),
.B1(n_1884),
.B2(n_1895),
.C(n_1901),
.Y(n_2084)
);

NOR2x1_ASAP7_75t_L g2085 ( 
.A(n_2083),
.B(n_1877),
.Y(n_2085)
);

NAND2xp5_ASAP7_75t_L g2086 ( 
.A(n_2080),
.B(n_2078),
.Y(n_2086)
);

OR2x2_ASAP7_75t_L g2087 ( 
.A(n_2080),
.B(n_2074),
.Y(n_2087)
);

OAI21xp33_ASAP7_75t_L g2088 ( 
.A1(n_2082),
.A2(n_2069),
.B(n_2075),
.Y(n_2088)
);

XNOR2xp5_ASAP7_75t_L g2089 ( 
.A(n_2079),
.B(n_2070),
.Y(n_2089)
);

NAND2xp5_ASAP7_75t_L g2090 ( 
.A(n_2081),
.B(n_2073),
.Y(n_2090)
);

INVx1_ASAP7_75t_L g2091 ( 
.A(n_2077),
.Y(n_2091)
);

AND2x2_ASAP7_75t_L g2092 ( 
.A(n_2084),
.B(n_1903),
.Y(n_2092)
);

AOI22xp33_ASAP7_75t_SL g2093 ( 
.A1(n_2091),
.A2(n_1884),
.B1(n_1877),
.B2(n_1891),
.Y(n_2093)
);

INVx1_ASAP7_75t_L g2094 ( 
.A(n_2086),
.Y(n_2094)
);

AOI22xp5_ASAP7_75t_L g2095 ( 
.A1(n_2090),
.A2(n_1884),
.B1(n_1877),
.B2(n_1891),
.Y(n_2095)
);

OAI22xp5_ASAP7_75t_L g2096 ( 
.A1(n_2089),
.A2(n_1884),
.B1(n_1877),
.B2(n_1891),
.Y(n_2096)
);

AOI21xp33_ASAP7_75t_L g2097 ( 
.A1(n_2085),
.A2(n_1884),
.B(n_1872),
.Y(n_2097)
);

OAI211xp5_ASAP7_75t_L g2098 ( 
.A1(n_2088),
.A2(n_1877),
.B(n_1899),
.C(n_1891),
.Y(n_2098)
);

NOR4xp25_ASAP7_75t_L g2099 ( 
.A(n_2094),
.B(n_2087),
.C(n_2092),
.D(n_1907),
.Y(n_2099)
);

NAND2xp5_ASAP7_75t_SL g2100 ( 
.A(n_2093),
.B(n_1891),
.Y(n_2100)
);

AND2x4_ASAP7_75t_L g2101 ( 
.A(n_2095),
.B(n_1899),
.Y(n_2101)
);

NAND4xp75_ASAP7_75t_L g2102 ( 
.A(n_2097),
.B(n_1907),
.C(n_1895),
.D(n_1900),
.Y(n_2102)
);

AND2x4_ASAP7_75t_L g2103 ( 
.A(n_2101),
.B(n_2100),
.Y(n_2103)
);

AOI322xp5_ASAP7_75t_L g2104 ( 
.A1(n_2103),
.A2(n_2099),
.A3(n_2098),
.B1(n_2102),
.B2(n_2096),
.C1(n_1907),
.C2(n_1900),
.Y(n_2104)
);

INVx2_ASAP7_75t_L g2105 ( 
.A(n_2104),
.Y(n_2105)
);

INVx3_ASAP7_75t_L g2106 ( 
.A(n_2104),
.Y(n_2106)
);

NAND2xp5_ASAP7_75t_L g2107 ( 
.A(n_2106),
.B(n_1872),
.Y(n_2107)
);

NAND2xp5_ASAP7_75t_SL g2108 ( 
.A(n_2106),
.B(n_1891),
.Y(n_2108)
);

INVx2_ASAP7_75t_L g2109 ( 
.A(n_2107),
.Y(n_2109)
);

CKINVDCx20_ASAP7_75t_R g2110 ( 
.A(n_2108),
.Y(n_2110)
);

OAI22xp5_ASAP7_75t_L g2111 ( 
.A1(n_2110),
.A2(n_2105),
.B1(n_1900),
.B2(n_1902),
.Y(n_2111)
);

AOI22xp5_ASAP7_75t_SL g2112 ( 
.A1(n_2111),
.A2(n_2109),
.B1(n_1891),
.B2(n_1899),
.Y(n_2112)
);

AOI22xp5_ASAP7_75t_L g2113 ( 
.A1(n_2112),
.A2(n_1902),
.B1(n_1901),
.B2(n_1891),
.Y(n_2113)
);

AO21x2_ASAP7_75t_L g2114 ( 
.A1(n_2113),
.A2(n_1902),
.B(n_1901),
.Y(n_2114)
);

OAI22xp33_ASAP7_75t_L g2115 ( 
.A1(n_2114),
.A2(n_1891),
.B1(n_1886),
.B2(n_1899),
.Y(n_2115)
);

OA22x2_ASAP7_75t_L g2116 ( 
.A1(n_2115),
.A2(n_1899),
.B1(n_1830),
.B2(n_1883),
.Y(n_2116)
);


endmodule