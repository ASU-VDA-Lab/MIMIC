module fake_ibex_1249_n_4896 (n_151, n_85, n_599, n_778, n_822, n_507, n_743, n_540, n_754, n_395, n_84, n_64, n_171, n_756, n_103, n_529, n_389, n_204, n_626, n_274, n_387, n_766, n_688, n_130, n_177, n_707, n_76, n_273, n_309, n_330, n_9, n_328, n_293, n_341, n_372, n_124, n_37, n_256, n_418, n_193, n_510, n_845, n_446, n_108, n_350, n_601, n_621, n_610, n_165, n_790, n_452, n_86, n_70, n_664, n_255, n_175, n_586, n_773, n_638, n_398, n_59, n_28, n_125, n_304, n_821, n_191, n_593, n_5, n_62, n_71, n_153, n_545, n_583, n_678, n_663, n_194, n_249, n_334, n_634, n_733, n_312, n_622, n_578, n_478, n_239, n_94, n_134, n_432, n_371, n_403, n_423, n_608, n_357, n_88, n_412, n_457, n_494, n_142, n_226, n_336, n_258, n_40, n_90, n_17, n_74, n_449, n_547, n_176, n_727, n_58, n_43, n_216, n_33, n_652, n_781, n_421, n_828, n_738, n_475, n_802, n_166, n_163, n_753, n_645, n_500, n_747, n_542, n_114, n_236, n_34, n_376, n_377, n_584, n_531, n_647, n_15, n_761, n_556, n_748, n_24, n_189, n_498, n_698, n_280, n_317, n_340, n_375, n_708, n_105, n_187, n_667, n_1, n_154, n_682, n_850, n_182, n_196, n_326, n_327, n_89, n_50, n_723, n_144, n_170, n_270, n_346, n_383, n_113, n_840, n_561, n_117, n_417, n_471, n_846, n_739, n_755, n_265, n_853, n_504, n_158, n_859, n_259, n_276, n_339, n_470, n_770, n_210, n_348, n_220, n_674, n_91, n_481, n_287, n_54, n_243, n_19, n_497, n_671, n_228, n_711, n_147, n_552, n_251, n_384, n_632, n_373, n_854, n_458, n_244, n_73, n_343, n_310, n_714, n_703, n_426, n_323, n_469, n_829, n_598, n_825, n_143, n_740, n_106, n_386, n_549, n_8, n_224, n_183, n_533, n_508, n_67, n_453, n_591, n_655, n_333, n_110, n_306, n_400, n_47, n_550, n_736, n_169, n_10, n_673, n_21, n_732, n_798, n_832, n_242, n_278, n_316, n_16, n_404, n_60, n_557, n_641, n_7, n_109, n_127, n_121, n_527, n_590, n_465, n_48, n_325, n_57, n_301, n_496, n_617, n_434, n_296, n_690, n_120, n_835, n_168, n_526, n_785, n_155, n_824, n_315, n_441, n_604, n_13, n_637, n_122, n_523, n_116, n_694, n_787, n_614, n_370, n_431, n_719, n_574, n_0, n_289, n_716, n_12, n_515, n_642, n_150, n_286, n_321, n_133, n_569, n_600, n_51, n_215, n_279, n_49, n_374, n_235, n_464, n_538, n_669, n_838, n_750, n_746, n_22, n_136, n_261, n_742, n_521, n_665, n_459, n_30, n_518, n_367, n_221, n_852, n_789, n_654, n_656, n_724, n_437, n_731, n_602, n_842, n_355, n_767, n_474, n_758, n_594, n_636, n_710, n_720, n_407, n_102, n_490, n_568, n_813, n_52, n_448, n_646, n_595, n_99, n_466, n_269, n_156, n_570, n_126, n_623, n_585, n_715, n_791, n_530, n_356, n_25, n_104, n_45, n_420, n_483, n_543, n_580, n_141, n_487, n_769, n_222, n_660, n_186, n_524, n_349, n_765, n_849, n_857, n_454, n_777, n_295, n_730, n_331, n_576, n_230, n_96, n_759, n_185, n_388, n_625, n_619, n_536, n_611, n_352, n_290, n_558, n_666, n_174, n_467, n_427, n_607, n_827, n_157, n_219, n_246, n_31, n_442, n_146, n_207, n_438, n_851, n_689, n_793, n_167, n_676, n_128, n_253, n_208, n_234, n_3, n_152, n_300, n_145, n_65, n_358, n_771, n_205, n_618, n_488, n_139, n_514, n_705, n_429, n_560, n_275, n_541, n_98, n_129, n_613, n_659, n_267, n_662, n_635, n_844, n_245, n_589, n_571, n_229, n_209, n_472, n_648, n_783, n_347, n_847, n_830, n_473, n_445, n_629, n_335, n_413, n_82, n_263, n_27, n_573, n_353, n_359, n_826, n_299, n_87, n_262, n_433, n_75, n_439, n_704, n_643, n_137, n_679, n_841, n_772, n_810, n_768, n_839, n_338, n_173, n_696, n_796, n_797, n_837, n_477, n_640, n_363, n_402, n_725, n_180, n_369, n_596, n_201, n_699, n_14, n_351, n_368, n_456, n_834, n_257, n_77, n_718, n_801, n_44, n_672, n_722, n_401, n_553, n_554, n_66, n_735, n_305, n_713, n_307, n_192, n_804, n_140, n_484, n_566, n_480, n_416, n_581, n_651, n_365, n_721, n_4, n_814, n_6, n_605, n_539, n_100, n_179, n_354, n_206, n_392, n_630, n_516, n_548, n_567, n_763, n_745, n_329, n_447, n_26, n_188, n_200, n_444, n_506, n_562, n_564, n_546, n_199, n_788, n_795, n_592, n_495, n_762, n_410, n_308, n_675, n_800, n_463, n_624, n_706, n_411, n_135, n_520, n_784, n_684, n_775, n_658, n_512, n_615, n_685, n_283, n_366, n_397, n_111, n_803, n_692, n_36, n_627, n_18, n_709, n_322, n_53, n_227, n_499, n_115, n_757, n_11, n_248, n_92, n_702, n_451, n_712, n_101, n_190, n_138, n_650, n_776, n_409, n_582, n_818, n_653, n_214, n_238, n_579, n_843, n_332, n_799, n_517, n_211, n_744, n_817, n_218, n_314, n_691, n_563, n_132, n_277, n_555, n_337, n_522, n_700, n_479, n_534, n_225, n_360, n_272, n_511, n_23, n_734, n_468, n_223, n_381, n_525, n_815, n_780, n_535, n_382, n_502, n_681, n_633, n_532, n_726, n_95, n_405, n_415, n_597, n_285, n_288, n_247, n_320, n_379, n_551, n_55, n_612, n_291, n_318, n_63, n_819, n_161, n_237, n_29, n_203, n_268, n_440, n_858, n_148, n_2, n_342, n_233, n_385, n_414, n_430, n_118, n_729, n_741, n_603, n_378, n_486, n_422, n_164, n_38, n_198, n_264, n_616, n_782, n_833, n_217, n_324, n_391, n_831, n_537, n_728, n_78, n_805, n_670, n_820, n_20, n_69, n_390, n_544, n_39, n_178, n_509, n_695, n_786, n_639, n_303, n_362, n_717, n_93, n_505, n_162, n_482, n_240, n_282, n_61, n_680, n_501, n_809, n_752, n_856, n_668, n_779, n_266, n_42, n_294, n_112, n_485, n_46, n_284, n_811, n_808, n_80, n_172, n_250, n_493, n_460, n_609, n_476, n_792, n_461, n_575, n_313, n_519, n_345, n_408, n_119, n_361, n_455, n_419, n_774, n_72, n_319, n_195, n_513, n_212, n_588, n_693, n_311, n_661, n_848, n_406, n_606, n_737, n_97, n_197, n_528, n_181, n_131, n_123, n_631, n_683, n_260, n_620, n_794, n_836, n_462, n_302, n_450, n_443, n_686, n_572, n_644, n_577, n_344, n_393, n_436, n_428, n_491, n_297, n_435, n_628, n_41, n_252, n_396, n_697, n_816, n_83, n_32, n_107, n_149, n_489, n_677, n_399, n_254, n_213, n_424, n_565, n_823, n_701, n_271, n_241, n_68, n_503, n_292, n_807, n_394, n_79, n_81, n_35, n_364, n_687, n_159, n_202, n_231, n_298, n_587, n_760, n_751, n_806, n_160, n_657, n_764, n_184, n_56, n_492, n_649, n_812, n_855, n_232, n_380, n_749, n_281, n_559, n_425, n_4896);

input n_151;
input n_85;
input n_599;
input n_778;
input n_822;
input n_507;
input n_743;
input n_540;
input n_754;
input n_395;
input n_84;
input n_64;
input n_171;
input n_756;
input n_103;
input n_529;
input n_389;
input n_204;
input n_626;
input n_274;
input n_387;
input n_766;
input n_688;
input n_130;
input n_177;
input n_707;
input n_76;
input n_273;
input n_309;
input n_330;
input n_9;
input n_328;
input n_293;
input n_341;
input n_372;
input n_124;
input n_37;
input n_256;
input n_418;
input n_193;
input n_510;
input n_845;
input n_446;
input n_108;
input n_350;
input n_601;
input n_621;
input n_610;
input n_165;
input n_790;
input n_452;
input n_86;
input n_70;
input n_664;
input n_255;
input n_175;
input n_586;
input n_773;
input n_638;
input n_398;
input n_59;
input n_28;
input n_125;
input n_304;
input n_821;
input n_191;
input n_593;
input n_5;
input n_62;
input n_71;
input n_153;
input n_545;
input n_583;
input n_678;
input n_663;
input n_194;
input n_249;
input n_334;
input n_634;
input n_733;
input n_312;
input n_622;
input n_578;
input n_478;
input n_239;
input n_94;
input n_134;
input n_432;
input n_371;
input n_403;
input n_423;
input n_608;
input n_357;
input n_88;
input n_412;
input n_457;
input n_494;
input n_142;
input n_226;
input n_336;
input n_258;
input n_40;
input n_90;
input n_17;
input n_74;
input n_449;
input n_547;
input n_176;
input n_727;
input n_58;
input n_43;
input n_216;
input n_33;
input n_652;
input n_781;
input n_421;
input n_828;
input n_738;
input n_475;
input n_802;
input n_166;
input n_163;
input n_753;
input n_645;
input n_500;
input n_747;
input n_542;
input n_114;
input n_236;
input n_34;
input n_376;
input n_377;
input n_584;
input n_531;
input n_647;
input n_15;
input n_761;
input n_556;
input n_748;
input n_24;
input n_189;
input n_498;
input n_698;
input n_280;
input n_317;
input n_340;
input n_375;
input n_708;
input n_105;
input n_187;
input n_667;
input n_1;
input n_154;
input n_682;
input n_850;
input n_182;
input n_196;
input n_326;
input n_327;
input n_89;
input n_50;
input n_723;
input n_144;
input n_170;
input n_270;
input n_346;
input n_383;
input n_113;
input n_840;
input n_561;
input n_117;
input n_417;
input n_471;
input n_846;
input n_739;
input n_755;
input n_265;
input n_853;
input n_504;
input n_158;
input n_859;
input n_259;
input n_276;
input n_339;
input n_470;
input n_770;
input n_210;
input n_348;
input n_220;
input n_674;
input n_91;
input n_481;
input n_287;
input n_54;
input n_243;
input n_19;
input n_497;
input n_671;
input n_228;
input n_711;
input n_147;
input n_552;
input n_251;
input n_384;
input n_632;
input n_373;
input n_854;
input n_458;
input n_244;
input n_73;
input n_343;
input n_310;
input n_714;
input n_703;
input n_426;
input n_323;
input n_469;
input n_829;
input n_598;
input n_825;
input n_143;
input n_740;
input n_106;
input n_386;
input n_549;
input n_8;
input n_224;
input n_183;
input n_533;
input n_508;
input n_67;
input n_453;
input n_591;
input n_655;
input n_333;
input n_110;
input n_306;
input n_400;
input n_47;
input n_550;
input n_736;
input n_169;
input n_10;
input n_673;
input n_21;
input n_732;
input n_798;
input n_832;
input n_242;
input n_278;
input n_316;
input n_16;
input n_404;
input n_60;
input n_557;
input n_641;
input n_7;
input n_109;
input n_127;
input n_121;
input n_527;
input n_590;
input n_465;
input n_48;
input n_325;
input n_57;
input n_301;
input n_496;
input n_617;
input n_434;
input n_296;
input n_690;
input n_120;
input n_835;
input n_168;
input n_526;
input n_785;
input n_155;
input n_824;
input n_315;
input n_441;
input n_604;
input n_13;
input n_637;
input n_122;
input n_523;
input n_116;
input n_694;
input n_787;
input n_614;
input n_370;
input n_431;
input n_719;
input n_574;
input n_0;
input n_289;
input n_716;
input n_12;
input n_515;
input n_642;
input n_150;
input n_286;
input n_321;
input n_133;
input n_569;
input n_600;
input n_51;
input n_215;
input n_279;
input n_49;
input n_374;
input n_235;
input n_464;
input n_538;
input n_669;
input n_838;
input n_750;
input n_746;
input n_22;
input n_136;
input n_261;
input n_742;
input n_521;
input n_665;
input n_459;
input n_30;
input n_518;
input n_367;
input n_221;
input n_852;
input n_789;
input n_654;
input n_656;
input n_724;
input n_437;
input n_731;
input n_602;
input n_842;
input n_355;
input n_767;
input n_474;
input n_758;
input n_594;
input n_636;
input n_710;
input n_720;
input n_407;
input n_102;
input n_490;
input n_568;
input n_813;
input n_52;
input n_448;
input n_646;
input n_595;
input n_99;
input n_466;
input n_269;
input n_156;
input n_570;
input n_126;
input n_623;
input n_585;
input n_715;
input n_791;
input n_530;
input n_356;
input n_25;
input n_104;
input n_45;
input n_420;
input n_483;
input n_543;
input n_580;
input n_141;
input n_487;
input n_769;
input n_222;
input n_660;
input n_186;
input n_524;
input n_349;
input n_765;
input n_849;
input n_857;
input n_454;
input n_777;
input n_295;
input n_730;
input n_331;
input n_576;
input n_230;
input n_96;
input n_759;
input n_185;
input n_388;
input n_625;
input n_619;
input n_536;
input n_611;
input n_352;
input n_290;
input n_558;
input n_666;
input n_174;
input n_467;
input n_427;
input n_607;
input n_827;
input n_157;
input n_219;
input n_246;
input n_31;
input n_442;
input n_146;
input n_207;
input n_438;
input n_851;
input n_689;
input n_793;
input n_167;
input n_676;
input n_128;
input n_253;
input n_208;
input n_234;
input n_3;
input n_152;
input n_300;
input n_145;
input n_65;
input n_358;
input n_771;
input n_205;
input n_618;
input n_488;
input n_139;
input n_514;
input n_705;
input n_429;
input n_560;
input n_275;
input n_541;
input n_98;
input n_129;
input n_613;
input n_659;
input n_267;
input n_662;
input n_635;
input n_844;
input n_245;
input n_589;
input n_571;
input n_229;
input n_209;
input n_472;
input n_648;
input n_783;
input n_347;
input n_847;
input n_830;
input n_473;
input n_445;
input n_629;
input n_335;
input n_413;
input n_82;
input n_263;
input n_27;
input n_573;
input n_353;
input n_359;
input n_826;
input n_299;
input n_87;
input n_262;
input n_433;
input n_75;
input n_439;
input n_704;
input n_643;
input n_137;
input n_679;
input n_841;
input n_772;
input n_810;
input n_768;
input n_839;
input n_338;
input n_173;
input n_696;
input n_796;
input n_797;
input n_837;
input n_477;
input n_640;
input n_363;
input n_402;
input n_725;
input n_180;
input n_369;
input n_596;
input n_201;
input n_699;
input n_14;
input n_351;
input n_368;
input n_456;
input n_834;
input n_257;
input n_77;
input n_718;
input n_801;
input n_44;
input n_672;
input n_722;
input n_401;
input n_553;
input n_554;
input n_66;
input n_735;
input n_305;
input n_713;
input n_307;
input n_192;
input n_804;
input n_140;
input n_484;
input n_566;
input n_480;
input n_416;
input n_581;
input n_651;
input n_365;
input n_721;
input n_4;
input n_814;
input n_6;
input n_605;
input n_539;
input n_100;
input n_179;
input n_354;
input n_206;
input n_392;
input n_630;
input n_516;
input n_548;
input n_567;
input n_763;
input n_745;
input n_329;
input n_447;
input n_26;
input n_188;
input n_200;
input n_444;
input n_506;
input n_562;
input n_564;
input n_546;
input n_199;
input n_788;
input n_795;
input n_592;
input n_495;
input n_762;
input n_410;
input n_308;
input n_675;
input n_800;
input n_463;
input n_624;
input n_706;
input n_411;
input n_135;
input n_520;
input n_784;
input n_684;
input n_775;
input n_658;
input n_512;
input n_615;
input n_685;
input n_283;
input n_366;
input n_397;
input n_111;
input n_803;
input n_692;
input n_36;
input n_627;
input n_18;
input n_709;
input n_322;
input n_53;
input n_227;
input n_499;
input n_115;
input n_757;
input n_11;
input n_248;
input n_92;
input n_702;
input n_451;
input n_712;
input n_101;
input n_190;
input n_138;
input n_650;
input n_776;
input n_409;
input n_582;
input n_818;
input n_653;
input n_214;
input n_238;
input n_579;
input n_843;
input n_332;
input n_799;
input n_517;
input n_211;
input n_744;
input n_817;
input n_218;
input n_314;
input n_691;
input n_563;
input n_132;
input n_277;
input n_555;
input n_337;
input n_522;
input n_700;
input n_479;
input n_534;
input n_225;
input n_360;
input n_272;
input n_511;
input n_23;
input n_734;
input n_468;
input n_223;
input n_381;
input n_525;
input n_815;
input n_780;
input n_535;
input n_382;
input n_502;
input n_681;
input n_633;
input n_532;
input n_726;
input n_95;
input n_405;
input n_415;
input n_597;
input n_285;
input n_288;
input n_247;
input n_320;
input n_379;
input n_551;
input n_55;
input n_612;
input n_291;
input n_318;
input n_63;
input n_819;
input n_161;
input n_237;
input n_29;
input n_203;
input n_268;
input n_440;
input n_858;
input n_148;
input n_2;
input n_342;
input n_233;
input n_385;
input n_414;
input n_430;
input n_118;
input n_729;
input n_741;
input n_603;
input n_378;
input n_486;
input n_422;
input n_164;
input n_38;
input n_198;
input n_264;
input n_616;
input n_782;
input n_833;
input n_217;
input n_324;
input n_391;
input n_831;
input n_537;
input n_728;
input n_78;
input n_805;
input n_670;
input n_820;
input n_20;
input n_69;
input n_390;
input n_544;
input n_39;
input n_178;
input n_509;
input n_695;
input n_786;
input n_639;
input n_303;
input n_362;
input n_717;
input n_93;
input n_505;
input n_162;
input n_482;
input n_240;
input n_282;
input n_61;
input n_680;
input n_501;
input n_809;
input n_752;
input n_856;
input n_668;
input n_779;
input n_266;
input n_42;
input n_294;
input n_112;
input n_485;
input n_46;
input n_284;
input n_811;
input n_808;
input n_80;
input n_172;
input n_250;
input n_493;
input n_460;
input n_609;
input n_476;
input n_792;
input n_461;
input n_575;
input n_313;
input n_519;
input n_345;
input n_408;
input n_119;
input n_361;
input n_455;
input n_419;
input n_774;
input n_72;
input n_319;
input n_195;
input n_513;
input n_212;
input n_588;
input n_693;
input n_311;
input n_661;
input n_848;
input n_406;
input n_606;
input n_737;
input n_97;
input n_197;
input n_528;
input n_181;
input n_131;
input n_123;
input n_631;
input n_683;
input n_260;
input n_620;
input n_794;
input n_836;
input n_462;
input n_302;
input n_450;
input n_443;
input n_686;
input n_572;
input n_644;
input n_577;
input n_344;
input n_393;
input n_436;
input n_428;
input n_491;
input n_297;
input n_435;
input n_628;
input n_41;
input n_252;
input n_396;
input n_697;
input n_816;
input n_83;
input n_32;
input n_107;
input n_149;
input n_489;
input n_677;
input n_399;
input n_254;
input n_213;
input n_424;
input n_565;
input n_823;
input n_701;
input n_271;
input n_241;
input n_68;
input n_503;
input n_292;
input n_807;
input n_394;
input n_79;
input n_81;
input n_35;
input n_364;
input n_687;
input n_159;
input n_202;
input n_231;
input n_298;
input n_587;
input n_760;
input n_751;
input n_806;
input n_160;
input n_657;
input n_764;
input n_184;
input n_56;
input n_492;
input n_649;
input n_812;
input n_855;
input n_232;
input n_380;
input n_749;
input n_281;
input n_559;
input n_425;

output n_4896;

wire n_1084;
wire n_4368;
wire n_2594;
wire n_1474;
wire n_1295;
wire n_1983;
wire n_2804;
wire n_4557;
wire n_3150;
wire n_992;
wire n_4773;
wire n_4798;
wire n_1582;
wire n_2201;
wire n_3853;
wire n_2512;
wire n_3590;
wire n_4449;
wire n_4056;
wire n_2960;
wire n_2175;
wire n_2071;
wire n_2796;
wire n_4688;
wire n_1110;
wire n_3610;
wire n_2607;
wire n_1382;
wire n_3548;
wire n_3911;
wire n_3144;
wire n_2569;
wire n_2949;
wire n_1998;
wire n_2840;
wire n_4234;
wire n_1596;
wire n_4883;
wire n_926;
wire n_3319;
wire n_1079;
wire n_3077;
wire n_4146;
wire n_2835;
wire n_4656;
wire n_3915;
wire n_1100;
wire n_3559;
wire n_4158;
wire n_4687;
wire n_4756;
wire n_4095;
wire n_2177;
wire n_1930;
wire n_2123;
wire n_4204;
wire n_4364;
wire n_1234;
wire n_3019;
wire n_4881;
wire n_2047;
wire n_1594;
wire n_1944;
wire n_2235;
wire n_1802;
wire n_2498;
wire n_3817;
wire n_3755;
wire n_2038;
wire n_2504;
wire n_1469;
wire n_4630;
wire n_3812;
wire n_2017;
wire n_873;
wire n_1227;
wire n_962;
wire n_4632;
wire n_1080;
wire n_909;
wire n_862;
wire n_2290;
wire n_4607;
wire n_3750;
wire n_4514;
wire n_957;
wire n_3838;
wire n_3255;
wire n_3272;
wire n_3674;
wire n_4249;
wire n_1652;
wire n_969;
wire n_1859;
wire n_1954;
wire n_2183;
wire n_4346;
wire n_2074;
wire n_2897;
wire n_4749;
wire n_1883;
wire n_1125;
wire n_4805;
wire n_2687;
wire n_3456;
wire n_2037;
wire n_4550;
wire n_4668;
wire n_1226;
wire n_1034;
wire n_2383;
wire n_3132;
wire n_1765;
wire n_4159;
wire n_872;
wire n_2392;
wire n_4651;
wire n_1873;
wire n_1619;
wire n_2640;
wire n_1666;
wire n_2682;
wire n_3605;
wire n_930;
wire n_4372;
wire n_1044;
wire n_3280;
wire n_3105;
wire n_3146;
wire n_4731;
wire n_1492;
wire n_1134;
wire n_4004;
wire n_1478;
wire n_1684;
wire n_4892;
wire n_1796;
wire n_3569;
wire n_4343;
wire n_1614;
wire n_2374;
wire n_3334;
wire n_3819;
wire n_2598;
wire n_4353;
wire n_4648;
wire n_1722;
wire n_4371;
wire n_3931;
wire n_911;
wire n_2023;
wire n_2720;
wire n_4421;
wire n_4601;
wire n_4179;
wire n_3870;
wire n_3340;
wire n_4142;
wire n_2335;
wire n_1233;
wire n_2322;
wire n_3025;
wire n_3411;
wire n_2955;
wire n_3458;
wire n_3653;
wire n_3519;
wire n_4360;
wire n_4785;
wire n_2276;
wire n_1045;
wire n_3235;
wire n_2989;
wire n_1856;
wire n_963;
wire n_1782;
wire n_2230;
wire n_2889;
wire n_3843;
wire n_2139;
wire n_2847;
wire n_3693;
wire n_3033;
wire n_4399;
wire n_1308;
wire n_1138;
wire n_2943;
wire n_1096;
wire n_2151;
wire n_2391;
wire n_1391;
wire n_3338;
wire n_4585;
wire n_3168;
wire n_884;
wire n_2396;
wire n_3135;
wire n_3440;
wire n_3904;
wire n_4378;
wire n_4239;
wire n_3175;
wire n_3729;
wire n_4169;
wire n_3484;
wire n_1971;
wire n_2485;
wire n_2479;
wire n_4477;
wire n_3570;
wire n_879;
wire n_2179;
wire n_4875;
wire n_1957;
wire n_4197;
wire n_2188;
wire n_1144;
wire n_2360;
wire n_2359;
wire n_4654;
wire n_2506;
wire n_3984;
wire n_4233;
wire n_4369;
wire n_4765;
wire n_1392;
wire n_2158;
wire n_1268;
wire n_2571;
wire n_3187;
wire n_3830;
wire n_3598;
wire n_2724;
wire n_3086;
wire n_2475;
wire n_3721;
wire n_4418;
wire n_948;
wire n_2799;
wire n_1752;
wire n_1829;
wire n_1338;
wire n_3726;
wire n_4708;
wire n_4592;
wire n_4172;
wire n_1730;
wire n_4277;
wire n_875;
wire n_1307;
wire n_4431;
wire n_1327;
wire n_2644;
wire n_4771;
wire n_4445;
wire n_876;
wire n_3211;
wire n_3479;
wire n_1840;
wire n_2837;
wire n_4652;
wire n_3751;
wire n_989;
wire n_3262;
wire n_3407;
wire n_3804;
wire n_1908;
wire n_4673;
wire n_3315;
wire n_3537;
wire n_4470;
wire n_4690;
wire n_1668;
wire n_3982;
wire n_2343;
wire n_2605;
wire n_2887;
wire n_1641;
wire n_2565;
wire n_4201;
wire n_1480;
wire n_1463;
wire n_1823;
wire n_3251;
wire n_4285;
wire n_1681;
wire n_2921;
wire n_4031;
wire n_4781;
wire n_3724;
wire n_1636;
wire n_939;
wire n_1687;
wire n_4120;
wire n_3192;
wire n_3753;
wire n_3533;
wire n_3896;
wire n_2192;
wire n_4423;
wire n_4584;
wire n_1766;
wire n_3184;
wire n_3566;
wire n_4065;
wire n_3469;
wire n_3170;
wire n_4155;
wire n_1922;
wire n_3890;
wire n_4578;
wire n_2032;
wire n_2820;
wire n_3323;
wire n_2311;
wire n_1937;
wire n_3392;
wire n_3347;
wire n_893;
wire n_3242;
wire n_3395;
wire n_3839;
wire n_1654;
wire n_4808;
wire n_4507;
wire n_3577;
wire n_2995;
wire n_4526;
wire n_4802;
wire n_4867;
wire n_3330;
wire n_1258;
wire n_1344;
wire n_2208;
wire n_2198;
wire n_1929;
wire n_2707;
wire n_3509;
wire n_3472;
wire n_1749;
wire n_4746;
wire n_1680;
wire n_1981;
wire n_1195;
wire n_2918;
wire n_3353;
wire n_3976;
wire n_4304;
wire n_4348;
wire n_4821;
wire n_1945;
wire n_2638;
wire n_4382;
wire n_3939;
wire n_4160;
wire n_2860;
wire n_2448;
wire n_3631;
wire n_4002;
wire n_2015;
wire n_3807;
wire n_4874;
wire n_2537;
wire n_1130;
wire n_4246;
wire n_2643;
wire n_4545;
wire n_1228;
wire n_2998;
wire n_2336;
wire n_3987;
wire n_3845;
wire n_3641;
wire n_2163;
wire n_4450;
wire n_3969;
wire n_4467;
wire n_1081;
wire n_4437;
wire n_4840;
wire n_4801;
wire n_4887;
wire n_2354;
wire n_3639;
wire n_3856;
wire n_1155;
wire n_1292;
wire n_3996;
wire n_4311;
wire n_2432;
wire n_3043;
wire n_2873;
wire n_1576;
wire n_1664;
wire n_4144;
wire n_2273;
wire n_3298;
wire n_1427;
wire n_4447;
wire n_4491;
wire n_4672;
wire n_1133;
wire n_3049;
wire n_2421;
wire n_1926;
wire n_3208;
wire n_4015;
wire n_904;
wire n_2363;
wire n_2814;
wire n_3237;
wire n_4211;
wire n_3264;
wire n_3204;
wire n_4119;
wire n_4569;
wire n_2003;
wire n_1970;
wire n_3671;
wire n_3946;
wire n_3727;
wire n_2621;
wire n_3620;
wire n_1778;
wire n_2558;
wire n_2953;
wire n_2922;
wire n_2347;
wire n_3881;
wire n_3949;
wire n_3507;
wire n_3884;
wire n_3103;
wire n_2839;
wire n_3926;
wire n_1030;
wire n_1698;
wire n_3688;
wire n_1094;
wire n_2462;
wire n_3770;
wire n_1496;
wire n_1910;
wire n_2333;
wire n_2436;
wire n_1663;
wire n_2705;
wire n_1214;
wire n_1274;
wire n_4591;
wire n_2527;
wire n_1606;
wire n_3711;
wire n_1595;
wire n_2164;
wire n_4267;
wire n_1509;
wire n_1648;
wire n_1618;
wire n_2944;
wire n_4349;
wire n_1886;
wire n_2269;
wire n_3748;
wire n_4723;
wire n_1841;
wire n_1070;
wire n_2472;
wire n_4389;
wire n_4510;
wire n_2685;
wire n_2846;
wire n_3197;
wire n_3699;
wire n_3668;
wire n_1955;
wire n_4312;
wire n_4567;
wire n_917;
wire n_4556;
wire n_2249;
wire n_2413;
wire n_2362;
wire n_968;
wire n_3148;
wire n_3022;
wire n_2822;
wire n_4014;
wire n_4779;
wire n_1253;
wire n_3707;
wire n_1306;
wire n_1484;
wire n_2686;
wire n_1493;
wire n_2597;
wire n_4217;
wire n_4214;
wire n_1313;
wire n_3973;
wire n_4430;
wire n_2774;
wire n_3151;
wire n_2090;
wire n_4223;
wire n_2260;
wire n_3977;
wire n_4724;
wire n_4769;
wire n_3125;
wire n_3722;
wire n_2812;
wire n_4889;
wire n_3802;
wire n_3681;
wire n_2753;
wire n_3603;
wire n_1638;
wire n_4221;
wire n_4721;
wire n_2215;
wire n_1449;
wire n_1071;
wire n_1723;
wire n_1960;
wire n_2663;
wire n_3882;
wire n_3129;
wire n_4806;
wire n_937;
wire n_2595;
wire n_2116;
wire n_3979;
wire n_3714;
wire n_3592;
wire n_4650;
wire n_1645;
wire n_3186;
wire n_4433;
wire n_973;
wire n_1038;
wire n_2280;
wire n_1943;
wire n_3541;
wire n_1863;
wire n_2844;
wire n_4428;
wire n_4784;
wire n_1269;
wire n_2393;
wire n_2773;
wire n_3565;
wire n_4766;
wire n_3883;
wire n_3097;
wire n_2906;
wire n_3030;
wire n_3943;
wire n_4563;
wire n_3809;
wire n_979;
wire n_4503;
wire n_1309;
wire n_1999;
wire n_3810;
wire n_3718;
wire n_1316;
wire n_1562;
wire n_3917;
wire n_1215;
wire n_3679;
wire n_4854;
wire n_3579;
wire n_2777;
wire n_2480;
wire n_3769;
wire n_1445;
wire n_2283;
wire n_2806;
wire n_3910;
wire n_2813;
wire n_2147;
wire n_4517;
wire n_4295;
wire n_1716;
wire n_4238;
wire n_1466;
wire n_1412;
wire n_3210;
wire n_3221;
wire n_3667;
wire n_1672;
wire n_4511;
wire n_1007;
wire n_2253;
wire n_4479;
wire n_1276;
wire n_3822;
wire n_4171;
wire n_1637;
wire n_3310;
wire n_2900;
wire n_4182;
wire n_3858;
wire n_1401;
wire n_4173;
wire n_3764;
wire n_3795;
wire n_4788;
wire n_4754;
wire n_1817;
wire n_2951;
wire n_2145;
wire n_2122;
wire n_1588;
wire n_3765;
wire n_2216;
wire n_1301;
wire n_2579;
wire n_4166;
wire n_2876;
wire n_2242;
wire n_869;
wire n_1620;
wire n_4259;
wire n_4845;
wire n_1561;
wire n_3301;
wire n_2370;
wire n_4600;
wire n_2025;
wire n_1078;
wire n_2247;
wire n_3451;
wire n_4422;
wire n_1219;
wire n_4513;
wire n_1865;
wire n_3177;
wire n_3518;
wire n_4188;
wire n_3399;
wire n_1252;
wire n_2022;
wire n_4786;
wire n_4842;
wire n_4850;
wire n_2730;
wire n_3967;
wire n_1170;
wire n_1927;
wire n_2373;
wire n_1869;
wire n_3842;
wire n_1853;
wire n_2275;
wire n_2980;
wire n_4735;
wire n_2189;
wire n_2482;
wire n_3799;
wire n_2767;
wire n_3676;
wire n_4667;
wire n_2899;
wire n_2826;
wire n_2112;
wire n_1753;
wire n_3351;
wire n_1322;
wire n_4457;
wire n_4060;
wire n_2008;
wire n_1305;
wire n_2088;
wire n_4610;
wire n_1248;
wire n_2762;
wire n_2171;
wire n_3307;
wire n_4774;
wire n_1388;
wire n_2859;
wire n_4711;
wire n_2564;
wire n_3780;
wire n_3023;
wire n_1653;
wire n_4067;
wire n_4799;
wire n_1375;
wire n_3224;
wire n_1356;
wire n_894;
wire n_1118;
wire n_2591;
wire n_4481;
wire n_1881;
wire n_3762;
wire n_3965;
wire n_1969;
wire n_3798;
wire n_4809;
wire n_1296;
wire n_3948;
wire n_3060;
wire n_4124;
wire n_4671;
wire n_971;
wire n_1326;
wire n_4444;
wire n_1350;
wire n_3627;
wire n_906;
wire n_4499;
wire n_2957;
wire n_4676;
wire n_2586;
wire n_3958;
wire n_1764;
wire n_1093;
wire n_2412;
wire n_2783;
wire n_4393;
wire n_978;
wire n_3777;
wire n_899;
wire n_1799;
wire n_3293;
wire n_1019;
wire n_902;
wire n_1689;
wire n_1250;
wire n_2550;
wire n_1190;
wire n_1304;
wire n_4595;
wire n_2541;
wire n_4598;
wire n_2987;
wire n_881;
wire n_4879;
wire n_3259;
wire n_1702;
wire n_3916;
wire n_4553;
wire n_3381;
wire n_3630;
wire n_1558;
wire n_2750;
wire n_1650;
wire n_1520;
wire n_1073;
wire n_1453;
wire n_3961;
wire n_1108;
wire n_2722;
wire n_4533;
wire n_2509;
wire n_2727;
wire n_3618;
wire n_4078;
wire n_4283;
wire n_1794;
wire n_1423;
wire n_3836;
wire n_4174;
wire n_1239;
wire n_4714;
wire n_4870;
wire n_2399;
wire n_1370;
wire n_2719;
wire n_1209;
wire n_1708;
wire n_2213;
wire n_3038;
wire n_3732;
wire n_3779;
wire n_3521;
wire n_3203;
wire n_3295;
wire n_3923;
wire n_4392;
wire n_2723;
wire n_1616;
wire n_3199;
wire n_3808;
wire n_4455;
wire n_4054;
wire n_3093;
wire n_1569;
wire n_2664;
wire n_4804;
wire n_1434;
wire n_3716;
wire n_1649;
wire n_2389;
wire n_3450;
wire n_4129;
wire n_4518;
wire n_4732;
wire n_4012;
wire n_1936;
wire n_2114;
wire n_1717;
wire n_3567;
wire n_2107;
wire n_1609;
wire n_2257;
wire n_3435;
wire n_4828;
wire n_4856;
wire n_4352;
wire n_3530;
wire n_4480;
wire n_1613;
wire n_1988;
wire n_1132;
wire n_892;
wire n_1467;
wire n_4548;
wire n_1803;
wire n_2401;
wire n_1787;
wire n_2782;
wire n_2511;
wire n_3217;
wire n_1281;
wire n_3094;
wire n_3874;
wire n_4258;
wire n_4535;
wire n_1447;
wire n_2166;
wire n_2451;
wire n_4665;
wire n_2150;
wire n_1549;
wire n_4290;
wire n_2631;
wire n_1867;
wire n_1531;
wire n_2919;
wire n_3909;
wire n_4252;
wire n_1332;
wire n_2660;
wire n_4505;
wire n_3971;
wire n_2661;
wire n_4079;
wire n_4219;
wire n_4577;
wire n_2292;
wire n_3573;
wire n_4604;
wire n_3563;
wire n_3510;
wire n_3560;
wire n_4248;
wire n_2334;
wire n_1424;
wire n_3467;
wire n_2444;
wire n_2350;
wire n_1742;
wire n_2625;
wire n_4240;
wire n_3652;
wire n_1818;
wire n_870;
wire n_2199;
wire n_1709;
wire n_1610;
wire n_2219;
wire n_4398;
wire n_3847;
wire n_1298;
wire n_1844;
wire n_4522;
wire n_1387;
wire n_2649;
wire n_1040;
wire n_2203;
wire n_4055;
wire n_2693;
wire n_3194;
wire n_3607;
wire n_3371;
wire n_4692;
wire n_4713;
wire n_1159;
wire n_1368;
wire n_2281;
wire n_4476;
wire n_1154;
wire n_3202;
wire n_2539;
wire n_2431;
wire n_1701;
wire n_2084;
wire n_1243;
wire n_3572;
wire n_2387;
wire n_2646;
wire n_3375;
wire n_2397;
wire n_1121;
wire n_2746;
wire n_3241;
wire n_4615;
wire n_4823;
wire n_2256;
wire n_3317;
wire n_3887;
wire n_3963;
wire n_3800;
wire n_3461;
wire n_2445;
wire n_2729;
wire n_1571;
wire n_1980;
wire n_3951;
wire n_3355;
wire n_2529;
wire n_4103;
wire n_3583;
wire n_2019;
wire n_4126;
wire n_4710;
wire n_1407;
wire n_3282;
wire n_4435;
wire n_4680;
wire n_1235;
wire n_1821;
wire n_3832;
wire n_3508;
wire n_1003;
wire n_4649;
wire n_4755;
wire n_889;
wire n_3827;
wire n_2708;
wire n_3156;
wire n_4303;
wire n_3457;
wire n_2748;
wire n_4757;
wire n_1058;
wire n_4803;
wire n_1835;
wire n_1862;
wire n_2224;
wire n_2697;
wire n_3531;
wire n_4693;
wire n_3415;
wire n_2470;
wire n_2355;
wire n_2890;
wire n_3698;
wire n_2731;
wire n_4451;
wire n_1543;
wire n_4653;
wire n_3466;
wire n_3386;
wire n_2233;
wire n_4400;
wire n_2499;
wire n_4568;
wire n_3370;
wire n_4359;
wire n_1504;
wire n_3814;
wire n_1519;
wire n_1425;
wire n_4812;
wire n_1781;
wire n_3888;
wire n_2069;
wire n_4331;
wire n_2602;
wire n_4090;
wire n_1441;
wire n_4105;
wire n_4549;
wire n_4573;
wire n_4206;
wire n_2028;
wire n_3309;
wire n_3678;
wire n_4136;
wire n_1924;
wire n_4216;
wire n_2856;
wire n_1921;
wire n_3024;
wire n_4767;
wire n_1156;
wire n_4358;
wire n_2857;
wire n_1293;
wire n_1360;
wire n_1555;
wire n_1394;
wire n_1347;
wire n_3968;
wire n_4825;
wire n_3950;
wire n_4177;
wire n_2070;
wire n_1042;
wire n_1888;
wire n_3471;
wire n_4098;
wire n_3117;
wire n_3320;
wire n_1786;
wire n_2033;
wire n_3039;
wire n_3900;
wire n_1319;
wire n_4376;
wire n_4050;
wire n_1553;
wire n_3478;
wire n_3701;
wire n_3542;
wire n_4623;
wire n_1041;
wire n_4700;
wire n_2766;
wire n_3756;
wire n_2828;
wire n_3754;
wire n_4411;
wire n_1964;
wire n_4523;
wire n_4156;
wire n_4408;
wire n_1090;
wire n_3720;
wire n_3374;
wire n_1196;
wire n_3704;
wire n_1182;
wire n_1271;
wire n_3811;
wire n_4074;
wire n_2416;
wire n_3633;
wire n_4878;
wire n_2786;
wire n_1731;
wire n_1905;
wire n_2962;
wire n_1031;
wire n_3416;
wire n_4355;
wire n_2879;
wire n_2958;
wire n_3147;
wire n_3694;
wire n_2052;
wire n_3690;
wire n_981;
wire n_3628;
wire n_3983;
wire n_2425;
wire n_2800;
wire n_4225;
wire n_3514;
wire n_3091;
wire n_4037;
wire n_4582;
wire n_3006;
wire n_3348;
wire n_2118;
wire n_2259;
wire n_3859;
wire n_2162;
wire n_4489;
wire n_2236;
wire n_3455;
wire n_4758;
wire n_4834;
wire n_3957;
wire n_3660;
wire n_2377;
wire n_2718;
wire n_2577;
wire n_4712;
wire n_1591;
wire n_3426;
wire n_3165;
wire n_4308;
wire n_2289;
wire n_2288;
wire n_2841;
wire n_4271;
wire n_3075;
wire n_1671;
wire n_1795;
wire n_1409;
wire n_1015;
wire n_3634;
wire n_3448;
wire n_2744;
wire n_2101;
wire n_2795;
wire n_3524;
wire n_3788;
wire n_1377;
wire n_2473;
wire n_4096;
wire n_4419;
wire n_1583;
wire n_3520;
wire n_4404;
wire n_1521;
wire n_2632;
wire n_1152;
wire n_2456;
wire n_3054;
wire n_2924;
wire n_2264;
wire n_2076;
wire n_2599;
wire n_974;
wire n_1036;
wire n_1831;
wire n_3626;
wire n_3733;
wire n_4853;
wire n_864;
wire n_1987;
wire n_4571;
wire n_959;
wire n_1106;
wire n_1312;
wire n_4655;
wire n_1129;
wire n_1244;
wire n_3171;
wire n_1733;
wire n_3365;
wire n_3684;
wire n_1634;
wire n_3986;
wire n_2853;
wire n_1932;
wire n_4725;
wire n_3775;
wire n_1452;
wire n_1552;
wire n_1318;
wire n_4006;
wire n_1508;
wire n_2217;
wire n_3741;
wire n_3854;
wire n_1217;
wire n_3594;
wire n_2866;
wire n_3970;
wire n_3153;
wire n_3291;
wire n_4570;
wire n_4658;
wire n_2655;
wire n_3487;
wire n_2454;
wire n_1715;
wire n_3966;
wire n_4293;
wire n_1189;
wire n_4008;
wire n_3300;
wire n_1713;
wire n_3621;
wire n_901;
wire n_1577;
wire n_2036;
wire n_1255;
wire n_2829;
wire n_2968;
wire n_4253;
wire n_4039;
wire n_2740;
wire n_4494;
wire n_3473;
wire n_1700;
wire n_2623;
wire n_4681;
wire n_4122;
wire n_4542;
wire n_2622;
wire n_3232;
wire n_4250;
wire n_2819;
wire n_1218;
wire n_2178;
wire n_4572;
wire n_1181;
wire n_3263;
wire n_3815;
wire n_4374;
wire n_1140;
wire n_1985;
wire n_4375;
wire n_4501;
wire n_4205;
wire n_1772;
wire n_4740;
wire n_2858;
wire n_3708;
wire n_4882;
wire n_1056;
wire n_2626;
wire n_1283;
wire n_3007;
wire n_3790;
wire n_1446;
wire n_2404;
wire n_1487;
wire n_3078;
wire n_2789;
wire n_2603;
wire n_4403;
wire n_1421;
wire n_1203;
wire n_3640;
wire n_3218;
wire n_2821;
wire n_2424;
wire n_1793;
wire n_2573;
wire n_1237;
wire n_2880;
wire n_2390;
wire n_4768;
wire n_2423;
wire n_4230;
wire n_3849;
wire n_965;
wire n_1109;
wire n_4402;
wire n_2741;
wire n_2793;
wire n_4333;
wire n_4813;
wire n_3098;
wire n_3490;
wire n_3055;
wire n_1633;
wire n_3299;
wire n_4469;
wire n_4070;
wire n_2580;
wire n_3222;
wire n_1711;
wire n_3529;
wire n_3069;
wire n_4558;
wire n_3107;
wire n_3352;
wire n_3436;
wire n_4134;
wire n_1051;
wire n_4180;
wire n_4131;
wire n_1008;
wire n_3065;
wire n_2964;
wire n_2375;
wire n_4062;
wire n_1498;
wire n_4460;
wire n_2312;
wire n_2572;
wire n_2946;
wire n_1053;
wire n_4330;
wire n_1656;
wire n_1207;
wire n_4040;
wire n_1735;
wire n_1076;
wire n_2063;
wire n_1032;
wire n_936;
wire n_3082;
wire n_1884;
wire n_2176;
wire n_3813;
wire n_1825;
wire n_2805;
wire n_4232;
wire n_1589;
wire n_2717;
wire n_4504;
wire n_4199;
wire n_2204;
wire n_2863;
wire n_2575;
wire n_1210;
wire n_2319;
wire n_4527;
wire n_4864;
wire n_3757;
wire n_2877;
wire n_1933;
wire n_2522;
wire n_3357;
wire n_3855;
wire n_4033;
wire n_4608;
wire n_4485;
wire n_1996;
wire n_1510;
wire n_1201;
wire n_1842;
wire n_2852;
wire n_2132;
wire n_3964;
wire n_3110;
wire n_1677;
wire n_1246;
wire n_3364;
wire n_1236;
wire n_4384;
wire n_2297;
wire n_3429;
wire n_3306;
wire n_3412;
wire n_4231;
wire n_3037;
wire n_3188;
wire n_2780;
wire n_3787;
wire n_1792;
wire n_1712;
wire n_3250;
wire n_1984;
wire n_1568;
wire n_2885;
wire n_4762;
wire n_1877;
wire n_4537;
wire n_3445;
wire n_1477;
wire n_1184;
wire n_2080;
wire n_2220;
wire n_2585;
wire n_4005;
wire n_1724;
wire n_2554;
wire n_3155;
wire n_2838;
wire n_1364;
wire n_3183;
wire n_1540;
wire n_1676;
wire n_1013;
wire n_3243;
wire n_4323;
wire n_4407;
wire n_4184;
wire n_2468;
wire n_929;
wire n_3248;
wire n_3214;
wire n_1890;
wire n_1136;
wire n_1075;
wire n_1249;
wire n_3128;
wire n_4073;
wire n_1918;
wire n_2606;
wire n_3642;
wire n_2549;
wire n_4325;
wire n_2461;
wire n_3468;
wire n_2006;
wire n_2440;
wire n_4113;
wire n_1229;
wire n_4337;
wire n_1440;
wire n_4826;
wire n_1490;
wire n_2152;
wire n_4646;
wire n_907;
wire n_1179;
wire n_1990;
wire n_4818;
wire n_3680;
wire n_4462;
wire n_1153;
wire n_3624;
wire n_1751;
wire n_2787;
wire n_3785;
wire n_2467;
wire n_2146;
wire n_2341;
wire n_4540;
wire n_3525;
wire n_1737;
wire n_4292;
wire n_4187;
wire n_3145;
wire n_4819;
wire n_2779;
wire n_1117;
wire n_1273;
wire n_3821;
wire n_2547;
wire n_2930;
wire n_2616;
wire n_1748;
wire n_4261;
wire n_2662;
wire n_4884;
wire n_1083;
wire n_3205;
wire n_3872;
wire n_1014;
wire n_4490;
wire n_3801;
wire n_2883;
wire n_938;
wire n_1178;
wire n_2935;
wire n_878;
wire n_2441;
wire n_3503;
wire n_2358;
wire n_2490;
wire n_3127;
wire n_3496;
wire n_2361;
wire n_4063;
wire n_1464;
wire n_1566;
wire n_4362;
wire n_3568;
wire n_944;
wire n_4876;
wire n_3312;
wire n_4128;
wire n_4092;
wire n_3003;
wire n_4244;
wire n_1848;
wire n_4009;
wire n_2062;
wire n_2277;
wire n_3841;
wire n_2650;
wire n_1982;
wire n_2252;
wire n_3932;
wire n_2888;
wire n_2339;
wire n_3614;
wire n_4626;
wire n_1334;
wire n_3879;
wire n_1963;
wire n_3394;
wire n_1695;
wire n_3331;
wire n_1418;
wire n_2999;
wire n_2402;
wire n_1137;
wire n_2552;
wire n_2910;
wire n_3119;
wire n_2590;
wire n_4414;
wire n_1977;
wire n_2294;
wire n_1200;
wire n_2295;
wire n_2530;
wire n_3345;
wire n_4706;
wire n_2379;
wire n_1120;
wire n_2300;
wire n_2792;
wire n_4747;
wire n_1602;
wire n_2965;
wire n_4114;
wire n_1776;
wire n_2372;
wire n_3341;
wire n_2382;
wire n_4347;
wire n_1852;
wire n_4191;
wire n_1522;
wire n_2523;
wire n_2557;
wire n_3544;
wire n_3868;
wire n_1279;
wire n_2505;
wire n_931;
wire n_4791;
wire n_3488;
wire n_4209;
wire n_3554;
wire n_2481;
wire n_3692;
wire n_1064;
wire n_4409;
wire n_1408;
wire n_2832;
wire n_3913;
wire n_1028;
wire n_1264;
wire n_3535;
wire n_3730;
wire n_2808;
wire n_2287;
wire n_3597;
wire n_4525;
wire n_3396;
wire n_4011;
wire n_4190;
wire n_2954;
wire n_4307;
wire n_3526;
wire n_2102;
wire n_4356;
wire n_1935;
wire n_2046;
wire n_3367;
wire n_3492;
wire n_1146;
wire n_2785;
wire n_2751;
wire n_3558;
wire n_2142;
wire n_1548;
wire n_4824;
wire n_3703;
wire n_2977;
wire n_4443;
wire n_1682;
wire n_4151;
wire n_4625;
wire n_1608;
wire n_3776;
wire n_3599;
wire n_4170;
wire n_1009;
wire n_4554;
wire n_1260;
wire n_1896;
wire n_1704;
wire n_2160;
wire n_2699;
wire n_2234;
wire n_2991;
wire n_4097;
wire n_4861;
wire n_1436;
wire n_3239;
wire n_4137;
wire n_2600;
wire n_1485;
wire n_1069;
wire n_4424;
wire n_2239;
wire n_4152;
wire n_1465;
wire n_3952;
wire n_1352;
wire n_1171;
wire n_1126;
wire n_3826;
wire n_4674;
wire n_4365;
wire n_1232;
wire n_1979;
wire n_2328;
wire n_2715;
wire n_3781;
wire n_4679;
wire n_4596;
wire n_4415;
wire n_1345;
wire n_4456;
wire n_4215;
wire n_4587;
wire n_4315;
wire n_2434;
wire n_1590;
wire n_2332;
wire n_2971;
wire n_954;
wire n_3578;
wire n_4734;
wire n_1628;
wire n_1773;
wire n_2133;
wire n_3553;
wire n_3072;
wire n_1545;
wire n_4492;
wire n_3249;
wire n_3580;
wire n_2369;
wire n_3470;
wire n_3584;
wire n_1471;
wire n_1738;
wire n_3441;
wire n_3797;
wire n_4559;
wire n_4500;
wire n_1395;
wire n_998;
wire n_1729;
wire n_1115;
wire n_2551;
wire n_4641;
wire n_3281;
wire n_2823;
wire n_3274;
wire n_4064;
wire n_4660;
wire n_4110;
wire n_2094;
wire n_2613;
wire n_1479;
wire n_3505;
wire n_4427;
wire n_4564;
wire n_2306;
wire n_1046;
wire n_2419;
wire n_4379;
wire n_3397;
wire n_2934;
wire n_4145;
wire n_2807;
wire n_4047;
wire n_882;
wire n_4157;
wire n_942;
wire n_1627;
wire n_1431;
wire n_3956;
wire n_3880;
wire n_4042;
wire n_2525;
wire n_4664;
wire n_3829;
wire n_4579;
wire n_1864;
wire n_4624;
wire n_943;
wire n_4317;
wire n_2568;
wire n_3087;
wire n_2629;
wire n_3587;
wire n_1523;
wire n_1086;
wire n_2197;
wire n_1756;
wire n_2010;
wire n_2097;
wire n_2733;
wire n_2241;
wire n_1470;
wire n_2098;
wire n_2109;
wire n_1761;
wire n_3796;
wire n_2648;
wire n_2458;
wire n_4041;
wire n_2398;
wire n_1836;
wire n_3032;
wire n_3401;
wire n_4753;
wire n_1593;
wire n_986;
wire n_1420;
wire n_2651;
wire n_1750;
wire n_1775;
wire n_2833;
wire n_4297;
wire n_1699;
wire n_3179;
wire n_4894;
wire n_927;
wire n_1563;
wire n_4115;
wire n_2905;
wire n_3460;
wire n_3954;
wire n_3978;
wire n_2570;
wire n_4051;
wire n_4321;
wire n_4709;
wire n_3123;
wire n_4025;
wire n_1875;
wire n_3379;
wire n_1615;
wire n_2184;
wire n_2418;
wire n_1087;
wire n_3390;
wire n_3719;
wire n_4425;
wire n_1599;
wire n_1400;
wire n_1539;
wire n_1806;
wire n_2842;
wire n_2711;
wire n_3070;
wire n_3646;
wire n_3477;
wire n_2635;
wire n_2469;
wire n_1575;
wire n_2209;
wire n_4416;
wire n_3074;
wire n_3897;
wire n_4077;
wire n_4640;
wire n_4024;
wire n_3020;
wire n_3142;
wire n_3975;
wire n_3164;
wire n_3475;
wire n_1448;
wire n_2077;
wire n_3136;
wire n_2520;
wire n_2193;
wire n_2612;
wire n_3034;
wire n_4010;
wire n_4255;
wire n_2095;
wire n_3108;
wire n_2486;
wire n_2628;
wire n_2395;
wire n_951;
wire n_2521;
wire n_2908;
wire n_4059;
wire n_4561;
wire n_4130;
wire n_2053;
wire n_2752;
wire n_1580;
wire n_2124;
wire n_3991;
wire n_4361;
wire n_3974;
wire n_1574;
wire n_2200;
wire n_4642;
wire n_4764;
wire n_1705;
wire n_3625;
wire n_2304;
wire n_4237;
wire n_4683;
wire n_1746;
wire n_2716;
wire n_1439;
wire n_2263;
wire n_2212;
wire n_2352;
wire n_4839;
wire n_3495;
wire n_863;
wire n_2185;
wire n_4141;
wire n_4614;
wire n_3169;
wire n_1832;
wire n_1128;
wire n_2476;
wire n_2376;
wire n_2979;
wire n_3398;
wire n_1266;
wire n_1300;
wire n_3759;
wire n_4035;
wire n_2781;
wire n_4291;
wire n_3419;
wire n_3629;
wire n_4800;
wire n_4880;
wire n_2460;
wire n_2170;
wire n_4694;
wire n_3600;
wire n_1785;
wire n_4109;
wire n_1870;
wire n_2484;
wire n_3999;
wire n_4117;
wire n_2721;
wire n_1405;
wire n_2884;
wire n_3383;
wire n_4087;
wire n_3167;
wire n_3687;
wire n_997;
wire n_4154;
wire n_3735;
wire n_2308;
wire n_3459;
wire n_3238;
wire n_2986;
wire n_3498;
wire n_4520;
wire n_1428;
wire n_2691;
wire n_4026;
wire n_4318;
wire n_2243;
wire n_2400;
wire n_3731;
wire n_3092;
wire n_3555;
wire n_4385;
wire n_2903;
wire n_891;
wire n_3659;
wire n_3254;
wire n_4496;
wire n_4717;
wire n_2507;
wire n_2759;
wire n_3682;
wire n_1528;
wire n_1495;
wire n_3131;
wire n_3434;
wire n_4052;
wire n_2463;
wire n_2654;
wire n_3840;
wire n_2975;
wire n_1357;
wire n_2503;
wire n_4072;
wire n_2478;
wire n_3178;
wire n_2794;
wire n_4566;
wire n_4245;
wire n_1512;
wire n_3672;
wire n_2496;
wire n_3378;
wire n_3481;
wire n_3885;
wire n_2974;
wire n_871;
wire n_2990;
wire n_2923;
wire n_1339;
wire n_1544;
wire n_1426;
wire n_2365;
wire n_3449;
wire n_4100;
wire n_4719;
wire n_3517;
wire n_3350;
wire n_2245;
wire n_4872;
wire n_1315;
wire n_1413;
wire n_2464;
wire n_3877;
wire n_4873;
wire n_945;
wire n_2925;
wire n_2270;
wire n_3260;
wire n_4647;
wire n_1706;
wire n_3936;
wire n_1560;
wire n_1592;
wire n_2776;
wire n_1461;
wire n_3166;
wire n_3953;
wire n_2695;
wire n_2630;
wire n_903;
wire n_1967;
wire n_2340;
wire n_3385;
wire n_2117;
wire n_1095;
wire n_1328;
wire n_1265;
wire n_3834;
wire n_2488;
wire n_1378;
wire n_2042;
wire n_3656;
wire n_4837;
wire n_3257;
wire n_1048;
wire n_2459;
wire n_3137;
wire n_3116;
wire n_4426;
wire n_1925;
wire n_2439;
wire n_3638;
wire n_2106;
wire n_1430;
wire n_2414;
wire n_1251;
wire n_3090;
wire n_1247;
wire n_3816;
wire n_2450;
wire n_4636;
wire n_4195;
wire n_1475;
wire n_3337;
wire n_2465;
wire n_1263;
wire n_3316;
wire n_3925;
wire n_4089;
wire n_4176;
wire n_1185;
wire n_1683;
wire n_4256;
wire n_3575;
wire n_4454;
wire n_4851;
wire n_4175;
wire n_1122;
wire n_2765;
wire n_3387;
wire n_890;
wire n_874;
wire n_4278;
wire n_4495;
wire n_1505;
wire n_3010;
wire n_2941;
wire n_1163;
wire n_4609;
wire n_1514;
wire n_964;
wire n_2728;
wire n_3772;
wire n_4685;
wire n_2948;
wire n_916;
wire n_4458;
wire n_4322;
wire n_3428;
wire n_2298;
wire n_2771;
wire n_4336;
wire n_4822;
wire n_3219;
wire n_2936;
wire n_895;
wire n_3955;
wire n_3867;
wire n_1035;
wire n_2427;
wire n_2045;
wire n_3158;
wire n_1535;
wire n_2985;
wire n_3106;
wire n_4227;
wire n_2190;
wire n_1127;
wire n_932;
wire n_3657;
wire n_4716;
wire n_1972;
wire n_3080;
wire n_4030;
wire n_2772;
wire n_2778;
wire n_947;
wire n_1004;
wire n_4276;
wire n_4612;
wire n_3929;
wire n_1898;
wire n_1254;
wire n_1148;
wire n_1667;
wire n_1845;
wire n_1104;
wire n_2205;
wire n_1011;
wire n_2875;
wire n_3284;
wire n_2684;
wire n_2524;
wire n_1437;
wire n_3835;
wire n_3723;
wire n_2747;
wire n_3389;
wire n_1707;
wire n_1941;
wire n_3902;
wire n_4185;
wire n_2422;
wire n_3927;
wire n_4203;
wire n_2064;
wire n_3088;
wire n_1679;
wire n_2342;
wire n_2755;
wire n_2301;
wire n_1497;
wire n_2002;
wire n_2055;
wire n_4866;
wire n_3564;
wire n_4815;
wire n_2385;
wire n_3095;
wire n_3864;
wire n_3026;
wire n_2545;
wire n_1578;
wire n_3294;
wire n_4831;
wire n_2050;
wire n_1143;
wire n_1783;
wire n_2712;
wire n_3695;
wire n_3279;
wire n_2584;
wire n_972;
wire n_1815;
wire n_2500;
wire n_3344;
wire n_4381;
wire n_1917;
wire n_4314;
wire n_1444;
wire n_4133;
wire n_920;
wire n_4316;
wire n_2442;
wire n_3985;
wire n_1067;
wire n_3328;
wire n_2763;
wire n_2788;
wire n_4441;
wire n_994;
wire n_2000;
wire n_4083;
wire n_2089;
wire n_1857;
wire n_2761;
wire n_4020;
wire n_1920;
wire n_2696;
wire n_3252;
wire n_887;
wire n_1162;
wire n_1997;
wire n_2578;
wire n_4306;
wire n_2745;
wire n_1894;
wire n_2110;
wire n_2904;
wire n_2896;
wire n_3064;
wire n_4228;
wire n_4699;
wire n_2997;
wire n_3314;
wire n_961;
wire n_991;
wire n_1331;
wire n_1349;
wire n_1223;
wire n_2127;
wire n_3891;
wire n_3747;
wire n_1323;
wire n_1739;
wire n_4704;
wire n_3130;
wire n_1777;
wire n_3228;
wire n_3028;
wire n_3710;
wire n_1353;
wire n_3409;
wire n_2386;
wire n_3706;
wire n_3324;
wire n_1429;
wire n_3073;
wire n_2029;
wire n_3209;
wire n_2026;
wire n_1546;
wire n_3588;
wire n_4003;
wire n_4254;
wire n_4775;
wire n_4536;
wire n_3420;
wire n_1432;
wire n_4192;
wire n_2103;
wire n_3322;
wire n_4633;
wire n_1950;
wire n_4497;
wire n_1320;
wire n_4247;
wire n_4071;
wire n_4388;
wire n_996;
wire n_4593;
wire n_3632;
wire n_3914;
wire n_915;
wire n_2238;
wire n_3289;
wire n_1174;
wire n_4512;
wire n_1874;
wire n_1834;
wire n_3372;
wire n_3499;
wire n_4483;
wire n_4138;
wire n_3552;
wire n_4121;
wire n_2862;
wire n_3850;
wire n_3100;
wire n_4488;
wire n_4116;
wire n_4164;
wire n_3405;
wire n_1727;
wire n_3377;
wire n_1286;
wire n_1657;
wire n_1741;
wire n_1294;
wire n_1601;
wire n_900;
wire n_3784;
wire n_3414;
wire n_1351;
wire n_2933;
wire n_4183;
wire n_4118;
wire n_2138;
wire n_1380;
wire n_1367;
wire n_3336;
wire n_3240;
wire n_3828;
wire n_1291;
wire n_2895;
wire n_3763;
wire n_4858;
wire n_1914;
wire n_3833;
wire n_4284;
wire n_4814;
wire n_1458;
wire n_1694;
wire n_4370;
wire n_1460;
wire n_2041;
wire n_3201;
wire n_2271;
wire n_4621;
wire n_2356;
wire n_3339;
wire n_1830;
wire n_2261;
wire n_3016;
wire n_1629;
wire n_3476;
wire n_3673;
wire n_4066;
wire n_3990;
wire n_2994;
wire n_2011;
wire n_2620;
wire n_4044;
wire n_1826;
wire n_1855;
wire n_4241;
wire n_1662;
wire n_2105;
wire n_2187;
wire n_3556;
wire n_1340;
wire n_2694;
wire n_3443;
wire n_2562;
wire n_2642;
wire n_3029;
wire n_3269;
wire n_3609;
wire n_4135;
wire n_3447;
wire n_4678;
wire n_3771;
wire n_2647;
wire n_1626;
wire n_3995;
wire n_4104;
wire n_2223;
wire n_1660;
wire n_1850;
wire n_1643;
wire n_1670;
wire n_1789;
wire n_2415;
wire n_3876;
wire n_3152;
wire n_4000;
wire n_3154;
wire n_4123;
wire n_2344;
wire n_3589;
wire n_2317;
wire n_2556;
wire n_1112;
wire n_1267;
wire n_2384;
wire n_2683;
wire n_1384;
wire n_1376;
wire n_1537;
wire n_1858;
wire n_3432;
wire n_3523;
wire n_2815;
wire n_1816;
wire n_2446;
wire n_3388;
wire n_1612;
wire n_4619;
wire n_4645;
wire n_2318;
wire n_1172;
wire n_2659;
wire n_3908;
wire n_3616;
wire n_1099;
wire n_2141;
wire n_3696;
wire n_3113;
wire n_4305;
wire n_2902;
wire n_4048;
wire n_4084;
wire n_2909;
wire n_1422;
wire n_1527;
wire n_3174;
wire n_3960;
wire n_4007;
wire n_4848;
wire n_3608;
wire n_4339;
wire n_4269;
wire n_4085;
wire n_3190;
wire n_1524;
wire n_1055;
wire n_3878;
wire n_4016;
wire n_2849;
wire n_4661;
wire n_2947;
wire n_4080;
wire n_4707;
wire n_1754;
wire n_4286;
wire n_4429;
wire n_3048;
wire n_3686;
wire n_1177;
wire n_1025;
wire n_1991;
wire n_2566;
wire n_2679;
wire n_3292;
wire n_4028;
wire n_2210;
wire n_1517;
wire n_3940;
wire n_2502;
wire n_1225;
wire n_1962;
wire n_4860;
wire n_2346;
wire n_4695;
wire n_982;
wire n_4438;
wire n_3670;
wire n_1624;
wire n_1952;
wire n_2180;
wire n_3002;
wire n_3376;
wire n_2087;
wire n_2920;
wire n_3290;
wire n_4795;
wire n_1598;
wire n_2952;
wire n_4289;
wire n_2617;
wire n_3585;
wire n_977;
wire n_2878;
wire n_1895;
wire n_2250;
wire n_1491;
wire n_1860;
wire n_4163;
wire n_2831;
wire n_1810;
wire n_1763;
wire n_923;
wire n_3912;
wire n_3778;
wire n_3818;
wire n_1607;
wire n_2865;
wire n_2075;
wire n_4816;
wire n_3047;
wire n_1625;
wire n_2959;
wire n_2610;
wire n_4638;
wire n_2380;
wire n_2420;
wire n_3335;
wire n_4498;
wire n_3265;
wire n_2240;
wire n_933;
wire n_2221;
wire n_1774;
wire n_4846;
wire n_1797;
wire n_4750;
wire n_2516;
wire n_3993;
wire n_2120;
wire n_1037;
wire n_1899;
wire n_2031;
wire n_3669;
wire n_3427;
wire n_4001;
wire n_1348;
wire n_1289;
wire n_2892;
wire n_1021;
wire n_1557;
wire n_1188;
wire n_1567;
wire n_2007;
wire n_1191;
wire n_2004;
wire n_3356;
wire n_4099;
wire n_4377;
wire n_3431;
wire n_3220;
wire n_2024;
wire n_3783;
wire n_2086;
wire n_1503;
wire n_3422;
wire n_1052;
wire n_4264;
wire n_1942;
wire n_4832;
wire n_4326;
wire n_3666;
wire n_3141;
wire n_2309;
wire n_2274;
wire n_2698;
wire n_3899;
wire n_1617;
wire n_1839;
wire n_3930;
wire n_4149;
wire n_1587;
wire n_2330;
wire n_2639;
wire n_2555;
wire n_1259;
wire n_2108;
wire n_3099;
wire n_3712;
wire n_4101;
wire n_2535;
wire n_1001;
wire n_2945;
wire n_4745;
wire n_3057;
wire n_2143;
wire n_4057;
wire n_2410;
wire n_3760;
wire n_4319;
wire n_4637;
wire n_1396;
wire n_4792;
wire n_2916;
wire n_1923;
wire n_1224;
wire n_3206;
wire n_3736;
wire n_2196;
wire n_2739;
wire n_2611;
wire n_4021;
wire n_1538;
wire n_2528;
wire n_3773;
wire n_4383;
wire n_2548;
wire n_3216;
wire n_2709;
wire n_3061;
wire n_3717;
wire n_2633;
wire n_1017;
wire n_2244;
wire n_2604;
wire n_3462;
wire n_3424;
wire n_3745;
wire n_4373;
wire n_2351;
wire n_2437;
wire n_3664;
wire n_2049;
wire n_1456;
wire n_3245;
wire n_1889;
wire n_3907;
wire n_2113;
wire n_2665;
wire n_1124;
wire n_4855;
wire n_1690;
wire n_3063;
wire n_4543;
wire n_4466;
wire n_2688;
wire n_2881;
wire n_4643;
wire n_3862;
wire n_3302;
wire n_1673;
wire n_4132;
wire n_3361;
wire n_2018;
wire n_3134;
wire n_4736;
wire n_922;
wire n_2817;
wire n_1790;
wire n_993;
wire n_4202;
wire n_3196;
wire n_2085;
wire n_3304;
wire n_4287;
wire n_2581;
wire n_1725;
wire n_2809;
wire n_2149;
wire n_4603;
wire n_2237;
wire n_2268;
wire n_2320;
wire n_1135;
wire n_2255;
wire n_2001;
wire n_1820;
wire n_4300;
wire n_3921;
wire n_1800;
wire n_3277;
wire n_3480;
wire n_2758;
wire n_3746;
wire n_4417;
wire n_1494;
wire n_1550;
wire n_3906;
wire n_2060;
wire n_1066;
wire n_2214;
wire n_3474;
wire n_1169;
wire n_1726;
wire n_1946;
wire n_3111;
wire n_1938;
wire n_3452;
wire n_4022;
wire n_4212;
wire n_1241;
wire n_3645;
wire n_4262;
wire n_2589;
wire n_1072;
wire n_2194;
wire n_4827;
wire n_1231;
wire n_1173;
wire n_4019;
wire n_2736;
wire n_4320;
wire n_1208;
wire n_1604;
wire n_1639;
wire n_2735;
wire n_2845;
wire n_3506;
wire n_1976;
wire n_2154;
wire n_2035;
wire n_1337;
wire n_2732;
wire n_2984;
wire n_3162;
wire n_4436;
wire n_4599;
wire n_1906;
wire n_3004;
wire n_4697;
wire n_3886;
wire n_4890;
wire n_1647;
wire n_1901;
wire n_4357;
wire n_4538;
wire n_3096;
wire n_3333;
wire n_4509;
wire n_3705;
wire n_4023;
wire n_3031;
wire n_4849;
wire n_4783;
wire n_1278;
wire n_2059;
wire n_3276;
wire n_4366;
wire n_1006;
wire n_2956;
wire n_4730;
wire n_1415;
wire n_1238;
wire n_4616;
wire n_3959;
wire n_3743;
wire n_4760;
wire n_976;
wire n_1710;
wire n_4139;
wire n_3021;
wire n_1063;
wire n_4068;
wire n_4288;
wire n_2153;
wire n_2452;
wire n_1270;
wire n_2891;
wire n_2457;
wire n_4340;
wire n_3825;
wire n_2144;
wire n_1476;
wire n_1603;
wire n_935;
wire n_4763;
wire n_925;
wire n_2592;
wire n_1054;
wire n_2027;
wire n_3404;
wire n_2072;
wire n_4434;
wire n_2737;
wire n_2012;
wire n_2251;
wire n_2963;
wire n_3512;
wire n_4720;
wire n_1644;
wire n_3892;
wire n_1406;
wire n_1489;
wire n_3591;
wire n_1880;
wire n_1993;
wire n_4586;
wire n_4859;
wire n_3860;
wire n_2137;
wire n_1455;
wire n_1642;
wire n_1871;
wire n_2182;
wire n_2868;
wire n_3044;
wire n_3493;
wire n_2447;
wire n_2818;
wire n_3358;
wire n_3115;
wire n_1057;
wire n_4583;
wire n_1473;
wire n_3140;
wire n_3486;
wire n_2125;
wire n_2426;
wire n_2894;
wire n_1403;
wire n_2181;
wire n_3253;
wire n_2587;
wire n_1149;
wire n_4034;
wire n_1176;
wire n_1502;
wire n_1605;
wire n_868;
wire n_2099;
wire n_3920;
wire n_1202;
wire n_3848;
wire n_1065;
wire n_1897;
wire n_2477;
wire n_1457;
wire n_3172;
wire n_905;
wire n_4082;
wire n_2159;
wire n_3410;
wire n_975;
wire n_934;
wire n_4622;
wire n_3273;
wire n_4367;
wire n_950;
wire n_2700;
wire n_3139;
wire n_1222;
wire n_4282;
wire n_4715;
wire n_4885;
wire n_1630;
wire n_3408;
wire n_4475;
wire n_2286;
wire n_4222;
wire n_3182;
wire n_1879;
wire n_1959;
wire n_2563;
wire n_1198;
wire n_2206;
wire n_3734;
wire n_3637;
wire n_4893;
wire n_1311;
wire n_3538;
wire n_1261;
wire n_2299;
wire n_3393;
wire n_2078;
wire n_3650;
wire n_3327;
wire n_4588;
wire n_2265;
wire n_1114;
wire n_3513;
wire n_3709;
wire n_3011;
wire n_1167;
wire n_3231;
wire n_2677;
wire n_2531;
wire n_2315;
wire n_3647;
wire n_3623;
wire n_3138;
wire n_2157;
wire n_3212;
wire n_1282;
wire n_4029;
wire n_2067;
wire n_2517;
wire n_1321;
wire n_1779;
wire n_3446;
wire n_3349;
wire n_3619;
wire n_3928;
wire n_4043;
wire n_2489;
wire n_1770;
wire n_1107;
wire n_4167;
wire n_3058;
wire n_3454;
wire n_4334;
wire n_1846;
wire n_2211;
wire n_1573;
wire n_2950;
wire n_919;
wire n_4143;
wire n_2272;
wire n_1956;
wire n_3574;
wire n_4410;
wire n_2608;
wire n_4270;
wire n_3384;
wire n_4698;
wire n_2983;
wire n_4273;
wire n_1718;
wire n_3229;
wire n_2225;
wire n_2546;
wire n_4741;
wire n_3739;
wire n_1411;
wire n_2825;
wire n_1139;
wire n_1018;
wire n_2345;
wire n_1324;
wire n_4338;
wire n_1669;
wire n_1501;
wire n_2742;
wire n_4440;
wire n_1885;
wire n_1740;
wire n_1989;
wire n_3604;
wire n_1838;
wire n_3540;
wire n_3649;
wire n_3824;
wire n_2680;
wire n_1343;
wire n_1801;
wire n_3439;
wire n_1371;
wire n_4198;
wire n_4739;
wire n_1513;
wire n_3740;
wire n_4397;
wire n_4529;
wire n_3001;
wire n_2861;
wire n_2976;
wire n_4181;
wire n_2161;
wire n_2191;
wire n_3611;
wire n_2329;
wire n_1788;
wire n_4186;
wire n_2093;
wire n_2348;
wire n_2675;
wire n_2417;
wire n_2576;
wire n_2043;
wire n_3601;
wire n_4344;
wire n_2366;
wire n_4229;
wire n_4294;
wire n_1621;
wire n_2338;
wire n_3571;
wire n_1919;
wire n_1342;
wire n_4351;
wire n_2756;
wire n_2893;
wire n_2009;
wire n_2248;
wire n_958;
wire n_1175;
wire n_3500;
wire n_1416;
wire n_1659;
wire n_4200;
wire n_4162;
wire n_4111;
wire n_2850;
wire n_3465;
wire n_1221;
wire n_3962;
wire n_4575;
wire n_3875;
wire n_4847;
wire n_1047;
wire n_1878;
wire n_1515;
wire n_1374;
wire n_3846;
wire n_4341;
wire n_4328;
wire n_2851;
wire n_4759;
wire n_2438;
wire n_1435;
wire n_4127;
wire n_1688;
wire n_2973;
wire n_3651;
wire n_4620;
wire n_1433;
wire n_1314;
wire n_2567;
wire n_3059;
wire n_3085;
wire n_1242;
wire n_1119;
wire n_2229;
wire n_2867;
wire n_2810;
wire n_4666;
wire n_4770;
wire n_3871;
wire n_1085;
wire n_3027;
wire n_4076;
wire n_4189;
wire n_2388;
wire n_2981;
wire n_3438;
wire n_2222;
wire n_4439;
wire n_3112;
wire n_1907;
wire n_3464;
wire n_4835;
wire n_4390;
wire n_885;
wire n_4722;
wire n_1530;
wire n_3215;
wire n_3413;
wire n_877;
wire n_4580;
wire n_3994;
wire n_2871;
wire n_2135;
wire n_4565;
wire n_1088;
wire n_896;
wire n_2764;
wire n_2624;
wire n_1813;
wire n_1451;
wire n_1005;
wire n_1102;
wire n_3234;
wire n_3648;
wire n_4663;
wire n_2471;
wire n_4581;
wire n_1288;
wire n_4058;
wire n_4618;
wire n_4487;
wire n_1275;
wire n_985;
wire n_1165;
wire n_4519;
wire n_4611;
wire n_897;
wire n_1622;
wire n_2757;
wire n_4148;
wire n_2714;
wire n_3066;
wire n_2669;
wire n_4081;
wire n_4391;
wire n_2869;
wire n_1105;
wire n_1459;
wire n_912;
wire n_4032;
wire n_4829;
wire n_2898;
wire n_2232;
wire n_3121;
wire n_2455;
wire n_2121;
wire n_4541;
wire n_4515;
wire n_1893;
wire n_2519;
wire n_1570;
wire n_2231;
wire n_4530;
wire n_2874;
wire n_995;
wire n_2278;
wire n_1000;
wire n_4463;
wire n_2284;
wire n_1931;
wire n_2433;
wire n_2816;
wire n_2803;
wire n_3402;
wire n_1256;
wire n_2798;
wire n_4670;
wire n_3425;
wire n_1303;
wire n_1994;
wire n_1771;
wire n_3308;
wire n_1526;
wire n_4268;
wire n_1507;
wire n_1809;
wire n_1206;
wire n_2367;
wire n_3236;
wire n_2658;
wire n_3491;
wire n_3109;
wire n_1961;
wire n_3576;
wire n_4838;
wire n_4844;
wire n_3271;
wire n_3013;
wire n_2553;
wire n_1050;
wire n_2218;
wire n_2667;
wire n_4524;
wire n_3062;
wire n_4265;
wire n_3806;
wire n_1769;
wire n_2130;
wire n_3256;
wire n_1060;
wire n_4862;
wire n_3126;
wire n_1372;
wire n_1847;
wire n_1565;
wire n_1257;
wire n_3805;
wire n_2325;
wire n_2406;
wire n_1632;
wire n_2864;
wire n_3346;
wire n_3104;
wire n_4260;
wire n_3391;
wire n_4628;
wire n_4017;
wire n_1542;
wire n_946;
wire n_1547;
wire n_1586;
wire n_1362;
wire n_3497;
wire n_4696;
wire n_4895;
wire n_4178;
wire n_4324;
wire n_1097;
wire n_3354;
wire n_4069;
wire n_3288;
wire n_3373;
wire n_3382;
wire n_3122;
wire n_2518;
wire n_2784;
wire n_4236;
wire n_3012;
wire n_4313;
wire n_4140;
wire n_3045;
wire n_1909;
wire n_2543;
wire n_3368;
wire n_2381;
wire n_2313;
wire n_3561;
wire n_956;
wire n_3586;
wire n_4125;
wire n_2495;
wire n_4531;
wire n_4597;
wire n_4778;
wire n_2992;
wire n_1541;
wire n_2703;
wire n_1812;
wire n_3014;
wire n_4789;
wire n_1951;
wire n_1330;
wire n_4574;
wire n_4659;
wire n_2574;
wire n_1697;
wire n_2128;
wire n_1872;
wire n_4242;
wire n_4748;
wire n_1940;
wire n_2690;
wire n_1747;
wire n_3767;
wire n_1887;
wire n_1212;
wire n_1199;
wire n_3400;
wire n_3942;
wire n_4852;
wire n_2020;
wire n_3504;
wire n_1978;
wire n_2508;
wire n_3511;
wire n_2540;
wire n_4243;
wire n_1767;
wire n_1939;
wire n_2428;
wire n_3820;
wire n_3159;
wire n_1768;
wire n_1443;
wire n_3697;
wire n_2068;
wire n_2636;
wire n_2672;
wire n_3360;
wire n_1585;
wire n_1861;
wire n_2316;
wire n_3101;
wire n_1564;
wire n_4053;
wire n_1995;
wire n_4677;
wire n_1631;
wire n_2593;
wire n_1623;
wire n_2911;
wire n_861;
wire n_1828;
wire n_4279;
wire n_3937;
wire n_2364;
wire n_1389;
wire n_3303;
wire n_1131;
wire n_2641;
wire n_4729;
wire n_1798;
wire n_4555;
wire n_1077;
wire n_3120;
wire n_1554;
wire n_4843;
wire n_4761;
wire n_3549;
wire n_4751;
wire n_4562;
wire n_1481;
wire n_1584;
wire n_2021;
wire n_1928;
wire n_2713;
wire n_3227;
wire n_2938;
wire n_4235;
wire n_1438;
wire n_3774;
wire n_3972;
wire n_3342;
wire n_1973;
wire n_2314;
wire n_2939;
wire n_2156;
wire n_2494;
wire n_4036;
wire n_2126;
wire n_1147;
wire n_3403;
wire n_1363;
wire n_3863;
wire n_2228;
wire n_1691;
wire n_4453;
wire n_1098;
wire n_4474;
wire n_1518;
wire n_1366;
wire n_4350;
wire n_4380;
wire n_1187;
wire n_1361;
wire n_2034;
wire n_1693;
wire n_2790;
wire n_2872;
wire n_3173;
wire n_3102;
wire n_4345;
wire n_4478;
wire n_4281;
wire n_2411;
wire n_4332;
wire n_2081;
wire n_1892;
wire n_1061;
wire n_3539;
wire n_2266;
wire n_2993;
wire n_4473;
wire n_3433;
wire n_2061;
wire n_3018;
wire n_1373;
wire n_3998;
wire n_4820;
wire n_2449;
wire n_1686;
wire n_2131;
wire n_4464;
wire n_3866;
wire n_3761;
wire n_2526;
wire n_4794;
wire n_2830;
wire n_1302;
wire n_3803;
wire n_3017;
wire n_4675;
wire n_3083;
wire n_2083;
wire n_886;
wire n_3989;
wire n_2119;
wire n_1010;
wire n_4605;
wire n_4737;
wire n_3844;
wire n_883;
wire n_2207;
wire n_4210;
wire n_4752;
wire n_4546;
wire n_2044;
wire n_4049;
wire n_2542;
wire n_2091;
wire n_3918;
wire n_2843;
wire n_3362;
wire n_3035;
wire n_4165;
wire n_3191;
wire n_1029;
wire n_4891;
wire n_3485;
wire n_2394;
wire n_3051;
wire n_3305;
wire n_1635;
wire n_1572;
wire n_4810;
wire n_3149;
wire n_2827;
wire n_941;
wire n_1245;
wire n_1317;
wire n_3643;
wire n_2615;
wire n_3278;
wire n_2487;
wire n_2701;
wire n_3163;
wire n_2929;
wire n_3343;
wire n_3752;
wire n_4310;
wire n_3786;
wire n_4061;
wire n_1329;
wire n_2409;
wire n_2637;
wire n_2337;
wire n_4045;
wire n_4432;
wire n_2405;
wire n_2601;
wire n_4871;
wire n_2513;
wire n_4405;
wire n_3118;
wire n_1369;
wire n_1912;
wire n_1297;
wire n_3143;
wire n_3655;
wire n_1734;
wire n_3543;
wire n_3791;
wire n_3742;
wire n_4552;
wire n_1876;
wire n_2666;
wire n_3050;
wire n_4461;
wire n_4091;
wire n_2323;
wire n_3532;
wire n_4257;
wire n_4790;
wire n_1811;
wire n_928;
wire n_898;
wire n_1285;
wire n_3042;
wire n_967;
wire n_2561;
wire n_4263;
wire n_3725;
wire n_4516;
wire n_2913;
wire n_2491;
wire n_4686;
wire n_1529;
wire n_1381;
wire n_1824;
wire n_2254;
wire n_1597;
wire n_1161;
wire n_1103;
wire n_3522;
wire n_4682;
wire n_4528;
wire n_1486;
wire n_1068;
wire n_4363;
wire n_4888;
wire n_4502;
wire n_1833;
wire n_2914;
wire n_3551;
wire n_4196;
wire n_4335;
wire n_2371;
wire n_914;
wire n_3992;
wire n_4147;
wire n_3444;
wire n_1986;
wire n_3898;
wire n_4218;
wire n_3366;
wire n_4705;
wire n_4811;
wire n_2882;
wire n_1024;
wire n_3009;
wire n_1141;
wire n_3453;
wire n_3297;
wire n_3176;
wire n_4301;
wire n_4107;
wire n_4471;
wire n_1949;
wire n_1197;
wire n_2493;
wire n_2429;
wire n_2408;
wire n_3326;
wire n_1168;
wire n_865;
wire n_3581;
wire n_3000;
wire n_2115;
wire n_2013;
wire n_2140;
wire n_2134;
wire n_2483;
wire n_2305;
wire n_1556;
wire n_3547;
wire n_3423;
wire n_1192;
wire n_1646;
wire n_1290;
wire n_3700;
wire n_4161;
wire n_2514;
wire n_2466;
wire n_3661;
wire n_4386;
wire n_4733;
wire n_1759;
wire n_2048;
wire n_2760;
wire n_987;
wire n_4547;
wire n_1299;
wire n_2942;
wire n_4420;
wire n_4684;
wire n_2096;
wire n_3663;
wire n_3947;
wire n_4836;
wire n_2129;
wire n_3230;
wire n_3545;
wire n_1101;
wire n_2532;
wire n_3665;
wire n_2079;
wire n_4193;
wire n_4807;
wire n_4886;
wire n_2296;
wire n_4342;
wire n_3782;
wire n_1720;
wire n_880;
wire n_2671;
wire n_1911;
wire n_2293;
wire n_3296;
wire n_3831;
wire n_1336;
wire n_3068;
wire n_3071;
wire n_3683;
wire n_3919;
wire n_2734;
wire n_2870;
wire n_1166;
wire n_4302;
wire n_1390;
wire n_2775;
wire n_1023;
wire n_4869;
wire n_1358;
wire n_2310;
wire n_3318;
wire n_3223;
wire n_4013;
wire n_1211;
wire n_1397;
wire n_2674;
wire n_1284;
wire n_2005;
wire n_4482;
wire n_3794;
wire n_1359;
wire n_1116;
wire n_2811;
wire n_1758;
wire n_3226;
wire n_3702;
wire n_3981;
wire n_1532;
wire n_4406;
wire n_2848;
wire n_1419;
wire n_2689;
wire n_1784;
wire n_1685;
wire n_1992;
wire n_1082;
wire n_3200;
wire n_3430;
wire n_4493;
wire n_4797;
wire n_4738;
wire n_1213;
wire n_2596;
wire n_2801;
wire n_980;
wire n_1488;
wire n_1193;
wire n_3067;
wire n_2928;
wire n_2227;
wire n_2652;
wire n_3225;
wire n_1074;
wire n_3380;
wire n_3557;
wire n_3207;
wire n_3596;
wire n_1379;
wire n_1721;
wire n_2972;
wire n_2627;
wire n_1827;
wire n_953;
wire n_1180;
wire n_1462;
wire n_4657;
wire n_3606;
wire n_3369;
wire n_3823;
wire n_4718;
wire n_4086;
wire n_3185;
wire n_2326;
wire n_3869;
wire n_1866;
wire n_3852;
wire n_1220;
wire n_1398;
wire n_2169;
wire n_2111;
wire n_1262;
wire n_1904;
wire n_2966;
wire n_3084;
wire n_3036;
wire n_4112;
wire n_4634;
wire n_4644;
wire n_1692;
wire n_2501;
wire n_2051;
wire n_1012;
wire n_1805;
wire n_4207;
wire n_960;
wire n_1022;
wire n_4412;
wire n_4796;
wire n_1760;
wire n_3737;
wire n_1240;
wire n_2173;
wire n_1183;
wire n_4560;
wire n_3285;
wire n_3160;
wire n_3483;
wire n_4266;
wire n_4744;
wire n_1204;
wire n_1151;
wire n_2824;
wire n_1814;
wire n_3124;
wire n_3286;
wire n_999;
wire n_2634;
wire n_2982;
wire n_4038;
wire n_1092;
wire n_4472;
wire n_4793;
wire n_1808;
wire n_2768;
wire n_2668;
wire n_1658;
wire n_1386;
wire n_2588;
wire n_3015;
wire n_2931;
wire n_3321;
wire n_2492;
wire n_3081;
wire n_4639;
wire n_3636;
wire n_910;
wire n_2291;
wire n_3837;
wire n_4102;
wire n_3612;
wire n_3046;
wire n_2172;
wire n_4841;
wire n_1728;
wire n_1020;
wire n_4787;
wire n_3076;
wire n_1385;
wire n_1142;
wire n_2927;
wire n_4274;
wire n_1062;
wire n_4395;
wire n_4635;
wire n_4521;
wire n_1230;
wire n_4459;
wire n_1516;
wire n_1027;
wire n_4551;
wire n_3893;
wire n_4484;
wire n_3622;
wire n_3857;
wire n_2533;
wire n_1499;
wire n_1500;
wire n_4272;
wire n_2155;
wire n_2706;
wire n_1868;
wire n_966;
wire n_2148;
wire n_2303;
wire n_949;
wire n_2104;
wire n_2357;
wire n_2618;
wire n_2855;
wire n_2653;
wire n_4448;
wire n_4354;
wire n_924;
wire n_3938;
wire n_2937;
wire n_3728;
wire n_3359;
wire n_4532;
wire n_4401;
wire n_4727;
wire n_3114;
wire n_2331;
wire n_4296;
wire n_3332;
wire n_3905;
wire n_1600;
wire n_1661;
wire n_2967;
wire n_4701;
wire n_1965;
wire n_3005;
wire n_4413;
wire n_1757;
wire n_4627;
wire n_4743;
wire n_4088;
wire n_2136;
wire n_4309;
wire n_4726;
wire n_3617;
wire n_4027;
wire n_3602;
wire n_4298;
wire n_2403;
wire n_918;
wire n_3053;
wire n_2056;
wire n_1913;
wire n_2702;
wire n_3922;
wire n_2054;
wire n_1039;
wire n_2226;
wire n_3894;
wire n_2407;
wire n_2791;
wire n_1043;
wire n_1402;
wire n_2267;
wire n_2302;
wire n_1450;
wire n_2082;
wire n_2453;
wire n_2560;
wire n_3056;
wire n_3267;
wire n_2092;
wire n_4208;
wire n_3008;
wire n_1472;
wire n_1365;
wire n_2802;
wire n_2443;
wire n_3189;
wire n_3052;
wire n_4544;
wire n_4728;
wire n_2797;
wire n_2279;
wire n_1089;
wire n_4865;
wire n_1536;
wire n_1049;
wire n_1719;
wire n_1974;
wire n_2066;
wire n_1158;
wire n_2988;
wire n_3945;
wire n_4275;
wire n_1882;
wire n_4046;
wire n_2770;
wire n_2996;
wire n_2704;
wire n_2961;
wire n_3924;
wire n_1915;
wire n_2836;
wire n_4589;
wire n_940;
wire n_1762;
wire n_2534;
wire n_1404;
wire n_3689;
wire n_3582;
wire n_4631;
wire n_4830;
wire n_3283;
wire n_4468;
wire n_1736;
wire n_4617;
wire n_4442;
wire n_3421;
wire n_2907;
wire n_3311;
wire n_1160;
wire n_1442;
wire n_1948;
wire n_2168;
wire n_1216;
wire n_2681;
wire n_1891;
wire n_1026;
wire n_3247;
wire n_2886;
wire n_1454;
wire n_1033;
wire n_4094;
wire n_4689;
wire n_4772;
wire n_4857;
wire n_3613;
wire n_1383;
wire n_990;
wire n_3675;
wire n_1968;
wire n_4108;
wire n_2057;
wire n_4594;
wire n_2609;
wire n_4018;
wire n_2378;
wire n_888;
wire n_2749;
wire n_3658;
wire n_1325;
wire n_4613;
wire n_3133;
wire n_2754;
wire n_3527;
wire n_4629;
wire n_2014;
wire n_3901;
wire n_3041;
wire n_1483;
wire n_1703;
wire n_4539;
wire n_1205;
wire n_1822;
wire n_1953;
wire n_3715;
wire n_4194;
wire n_1059;
wire n_2969;
wire n_3713;
wire n_2692;
wire n_3550;
wire n_3261;
wire n_1804;
wire n_1581;
wire n_3287;
wire n_3534;
wire n_1837;
wire n_3889;
wire n_4776;
wire n_3325;
wire n_4299;
wire n_1744;
wire n_1975;
wire n_3437;
wire n_3744;
wire n_1414;
wire n_2324;
wire n_2246;
wire n_2738;
wire n_3861;
wire n_3161;
wire n_1002;
wire n_1851;
wire n_1755;
wire n_2195;
wire n_2940;
wire n_4150;
wire n_1111;
wire n_1819;
wire n_3313;
wire n_4702;
wire n_1341;
wire n_1807;
wire n_2670;
wire n_2645;
wire n_2202;
wire n_1310;
wire n_3275;
wire n_4486;
wire n_4863;
wire n_1745;
wire n_1714;
wire n_3198;
wire n_3463;
wire n_3941;
wire n_1958;
wire n_1611;
wire n_2559;
wire n_3516;
wire n_2262;
wire n_3562;
wire n_3933;
wire n_955;
wire n_1916;
wire n_1333;
wire n_2619;
wire n_2726;
wire n_2917;
wire n_3873;
wire n_4506;
wire n_3738;
wire n_2073;
wire n_4093;
wire n_952;
wire n_1675;
wire n_1947;
wire n_2165;
wire n_1640;
wire n_2016;
wire n_3157;
wire n_4669;
wire n_4226;
wire n_1551;
wire n_4153;
wire n_3793;
wire n_1145;
wire n_1533;
wire n_2307;
wire n_2515;
wire n_3792;
wire n_3546;
wire n_1511;
wire n_4329;
wire n_1791;
wire n_1113;
wire n_3089;
wire n_1651;
wire n_4817;
wire n_1966;
wire n_2058;
wire n_2678;
wire n_3406;
wire n_1468;
wire n_3442;
wire n_2327;
wire n_3758;
wire n_3988;
wire n_4780;
wire n_4877;
wire n_4327;
wire n_2656;
wire n_913;
wire n_2353;
wire n_4106;
wire n_4251;
wire n_4168;
wire n_1164;
wire n_2258;
wire n_3944;
wire n_3662;
wire n_3595;
wire n_1732;
wire n_3749;
wire n_2167;
wire n_3079;
wire n_1354;
wire n_3329;
wire n_4396;
wire n_2039;
wire n_1696;
wire n_1277;
wire n_1016;
wire n_3233;
wire n_4465;
wire n_1355;
wire n_3691;
wire n_4452;
wire n_2544;
wire n_3193;
wire n_4534;
wire n_3501;
wire n_3635;
wire n_866;
wire n_2538;
wire n_3270;
wire n_2582;
wire n_1559;
wire n_2321;
wire n_4590;
wire n_2915;
wire n_1579;
wire n_4446;
wire n_1280;
wire n_4602;
wire n_2854;
wire n_2932;
wire n_3258;
wire n_1335;
wire n_3266;
wire n_4280;
wire n_2285;
wire n_3213;
wire n_3789;
wire n_1934;
wire n_4394;
wire n_1900;
wire n_2040;
wire n_2174;
wire n_3246;
wire n_1843;
wire n_2186;
wire n_2510;
wire n_2030;
wire n_2614;
wire n_3418;
wire n_2435;
wire n_3934;
wire n_1665;
wire n_4576;
wire n_2583;
wire n_3417;
wire n_1678;
wire n_1091;
wire n_1780;
wire n_2725;
wire n_3865;
wire n_1287;
wire n_2769;
wire n_4606;
wire n_1482;
wire n_4220;
wire n_4075;
wire n_4782;
wire n_860;
wire n_1525;
wire n_3244;
wire n_3195;
wire n_3997;
wire n_4742;
wire n_3593;
wire n_2100;
wire n_2349;
wire n_1902;
wire n_2536;
wire n_3903;
wire n_2474;
wire n_3895;
wire n_1150;
wire n_1194;
wire n_1399;
wire n_3685;
wire n_4777;
wire n_3851;
wire n_4508;
wire n_1903;
wire n_4833;
wire n_1674;
wire n_1849;
wire n_3768;
wire n_867;
wire n_983;
wire n_1417;
wire n_3482;
wire n_2282;
wire n_4224;
wire n_970;
wire n_3654;
wire n_4868;
wire n_3980;
wire n_2430;
wire n_2673;
wire n_921;
wire n_2676;
wire n_3515;
wire n_3489;
wire n_4213;
wire n_2926;
wire n_1534;
wire n_2912;
wire n_3181;
wire n_908;
wire n_3536;
wire n_1346;
wire n_2834;
wire n_3644;
wire n_3268;
wire n_1123;
wire n_2710;
wire n_1272;
wire n_4387;
wire n_4703;
wire n_2497;
wire n_1393;
wire n_2970;
wire n_984;
wire n_1655;
wire n_3040;
wire n_3494;
wire n_4691;
wire n_2978;
wire n_3615;
wire n_1410;
wire n_988;
wire n_2368;
wire n_3363;
wire n_3528;
wire n_1157;
wire n_3502;
wire n_3677;
wire n_3766;
wire n_2657;
wire n_3935;
wire n_1186;
wire n_2065;
wire n_2901;
wire n_3180;
wire n_1743;
wire n_2743;
wire n_1854;
wire n_1506;
wire n_4662;

CKINVDCx5p33_ASAP7_75t_R g860 ( 
.A(n_230),
.Y(n_860)
);

INVx1_ASAP7_75t_L g861 ( 
.A(n_144),
.Y(n_861)
);

INVx1_ASAP7_75t_L g862 ( 
.A(n_243),
.Y(n_862)
);

CKINVDCx20_ASAP7_75t_R g863 ( 
.A(n_828),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_616),
.Y(n_864)
);

CKINVDCx5p33_ASAP7_75t_R g865 ( 
.A(n_859),
.Y(n_865)
);

CKINVDCx5p33_ASAP7_75t_R g866 ( 
.A(n_735),
.Y(n_866)
);

CKINVDCx5p33_ASAP7_75t_R g867 ( 
.A(n_20),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_680),
.Y(n_868)
);

CKINVDCx5p33_ASAP7_75t_R g869 ( 
.A(n_96),
.Y(n_869)
);

CKINVDCx5p33_ASAP7_75t_R g870 ( 
.A(n_811),
.Y(n_870)
);

CKINVDCx5p33_ASAP7_75t_R g871 ( 
.A(n_747),
.Y(n_871)
);

BUFx10_ASAP7_75t_L g872 ( 
.A(n_278),
.Y(n_872)
);

INVx2_ASAP7_75t_SL g873 ( 
.A(n_613),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_401),
.Y(n_874)
);

CKINVDCx5p33_ASAP7_75t_R g875 ( 
.A(n_504),
.Y(n_875)
);

INVx1_ASAP7_75t_L g876 ( 
.A(n_682),
.Y(n_876)
);

INVx2_ASAP7_75t_L g877 ( 
.A(n_762),
.Y(n_877)
);

CKINVDCx5p33_ASAP7_75t_R g878 ( 
.A(n_449),
.Y(n_878)
);

CKINVDCx5p33_ASAP7_75t_R g879 ( 
.A(n_39),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_257),
.Y(n_880)
);

INVx2_ASAP7_75t_L g881 ( 
.A(n_42),
.Y(n_881)
);

INVx2_ASAP7_75t_L g882 ( 
.A(n_285),
.Y(n_882)
);

HB1xp67_ASAP7_75t_L g883 ( 
.A(n_744),
.Y(n_883)
);

CKINVDCx5p33_ASAP7_75t_R g884 ( 
.A(n_259),
.Y(n_884)
);

INVx1_ASAP7_75t_SL g885 ( 
.A(n_329),
.Y(n_885)
);

CKINVDCx5p33_ASAP7_75t_R g886 ( 
.A(n_834),
.Y(n_886)
);

INVx2_ASAP7_75t_L g887 ( 
.A(n_301),
.Y(n_887)
);

CKINVDCx5p33_ASAP7_75t_R g888 ( 
.A(n_277),
.Y(n_888)
);

CKINVDCx5p33_ASAP7_75t_R g889 ( 
.A(n_547),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_204),
.Y(n_890)
);

CKINVDCx5p33_ASAP7_75t_R g891 ( 
.A(n_625),
.Y(n_891)
);

INVx1_ASAP7_75t_L g892 ( 
.A(n_702),
.Y(n_892)
);

CKINVDCx5p33_ASAP7_75t_R g893 ( 
.A(n_64),
.Y(n_893)
);

CKINVDCx5p33_ASAP7_75t_R g894 ( 
.A(n_647),
.Y(n_894)
);

BUFx6f_ASAP7_75t_L g895 ( 
.A(n_105),
.Y(n_895)
);

CKINVDCx5p33_ASAP7_75t_R g896 ( 
.A(n_838),
.Y(n_896)
);

BUFx3_ASAP7_75t_L g897 ( 
.A(n_451),
.Y(n_897)
);

CKINVDCx5p33_ASAP7_75t_R g898 ( 
.A(n_782),
.Y(n_898)
);

CKINVDCx5p33_ASAP7_75t_R g899 ( 
.A(n_819),
.Y(n_899)
);

BUFx2_ASAP7_75t_SL g900 ( 
.A(n_834),
.Y(n_900)
);

CKINVDCx5p33_ASAP7_75t_R g901 ( 
.A(n_220),
.Y(n_901)
);

BUFx10_ASAP7_75t_L g902 ( 
.A(n_512),
.Y(n_902)
);

INVx2_ASAP7_75t_L g903 ( 
.A(n_292),
.Y(n_903)
);

BUFx6f_ASAP7_75t_L g904 ( 
.A(n_500),
.Y(n_904)
);

CKINVDCx5p33_ASAP7_75t_R g905 ( 
.A(n_806),
.Y(n_905)
);

CKINVDCx5p33_ASAP7_75t_R g906 ( 
.A(n_677),
.Y(n_906)
);

CKINVDCx5p33_ASAP7_75t_R g907 ( 
.A(n_816),
.Y(n_907)
);

CKINVDCx14_ASAP7_75t_R g908 ( 
.A(n_846),
.Y(n_908)
);

CKINVDCx5p33_ASAP7_75t_R g909 ( 
.A(n_288),
.Y(n_909)
);

CKINVDCx5p33_ASAP7_75t_R g910 ( 
.A(n_139),
.Y(n_910)
);

INVx2_ASAP7_75t_L g911 ( 
.A(n_19),
.Y(n_911)
);

INVx2_ASAP7_75t_SL g912 ( 
.A(n_746),
.Y(n_912)
);

CKINVDCx5p33_ASAP7_75t_R g913 ( 
.A(n_742),
.Y(n_913)
);

CKINVDCx5p33_ASAP7_75t_R g914 ( 
.A(n_368),
.Y(n_914)
);

BUFx10_ASAP7_75t_L g915 ( 
.A(n_148),
.Y(n_915)
);

CKINVDCx5p33_ASAP7_75t_R g916 ( 
.A(n_827),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_504),
.Y(n_917)
);

CKINVDCx20_ASAP7_75t_R g918 ( 
.A(n_580),
.Y(n_918)
);

CKINVDCx5p33_ASAP7_75t_R g919 ( 
.A(n_484),
.Y(n_919)
);

CKINVDCx5p33_ASAP7_75t_R g920 ( 
.A(n_452),
.Y(n_920)
);

CKINVDCx5p33_ASAP7_75t_R g921 ( 
.A(n_108),
.Y(n_921)
);

CKINVDCx20_ASAP7_75t_R g922 ( 
.A(n_91),
.Y(n_922)
);

INVx2_ASAP7_75t_SL g923 ( 
.A(n_648),
.Y(n_923)
);

CKINVDCx5p33_ASAP7_75t_R g924 ( 
.A(n_68),
.Y(n_924)
);

CKINVDCx5p33_ASAP7_75t_R g925 ( 
.A(n_813),
.Y(n_925)
);

CKINVDCx5p33_ASAP7_75t_R g926 ( 
.A(n_63),
.Y(n_926)
);

CKINVDCx5p33_ASAP7_75t_R g927 ( 
.A(n_414),
.Y(n_927)
);

CKINVDCx5p33_ASAP7_75t_R g928 ( 
.A(n_27),
.Y(n_928)
);

CKINVDCx5p33_ASAP7_75t_R g929 ( 
.A(n_749),
.Y(n_929)
);

BUFx6f_ASAP7_75t_L g930 ( 
.A(n_821),
.Y(n_930)
);

CKINVDCx5p33_ASAP7_75t_R g931 ( 
.A(n_836),
.Y(n_931)
);

CKINVDCx5p33_ASAP7_75t_R g932 ( 
.A(n_668),
.Y(n_932)
);

INVx1_ASAP7_75t_L g933 ( 
.A(n_593),
.Y(n_933)
);

CKINVDCx5p33_ASAP7_75t_R g934 ( 
.A(n_431),
.Y(n_934)
);

INVx1_ASAP7_75t_L g935 ( 
.A(n_561),
.Y(n_935)
);

INVx1_ASAP7_75t_L g936 ( 
.A(n_643),
.Y(n_936)
);

CKINVDCx5p33_ASAP7_75t_R g937 ( 
.A(n_534),
.Y(n_937)
);

CKINVDCx5p33_ASAP7_75t_R g938 ( 
.A(n_3),
.Y(n_938)
);

CKINVDCx5p33_ASAP7_75t_R g939 ( 
.A(n_529),
.Y(n_939)
);

CKINVDCx5p33_ASAP7_75t_R g940 ( 
.A(n_826),
.Y(n_940)
);

CKINVDCx20_ASAP7_75t_R g941 ( 
.A(n_479),
.Y(n_941)
);

CKINVDCx5p33_ASAP7_75t_R g942 ( 
.A(n_697),
.Y(n_942)
);

INVx1_ASAP7_75t_L g943 ( 
.A(n_796),
.Y(n_943)
);

INVx1_ASAP7_75t_L g944 ( 
.A(n_849),
.Y(n_944)
);

CKINVDCx5p33_ASAP7_75t_R g945 ( 
.A(n_339),
.Y(n_945)
);

BUFx3_ASAP7_75t_L g946 ( 
.A(n_270),
.Y(n_946)
);

CKINVDCx5p33_ASAP7_75t_R g947 ( 
.A(n_183),
.Y(n_947)
);

INVx1_ASAP7_75t_L g948 ( 
.A(n_706),
.Y(n_948)
);

INVx1_ASAP7_75t_L g949 ( 
.A(n_96),
.Y(n_949)
);

BUFx2_ASAP7_75t_L g950 ( 
.A(n_26),
.Y(n_950)
);

BUFx3_ASAP7_75t_L g951 ( 
.A(n_760),
.Y(n_951)
);

CKINVDCx5p33_ASAP7_75t_R g952 ( 
.A(n_807),
.Y(n_952)
);

INVx2_ASAP7_75t_L g953 ( 
.A(n_600),
.Y(n_953)
);

INVx1_ASAP7_75t_L g954 ( 
.A(n_840),
.Y(n_954)
);

CKINVDCx5p33_ASAP7_75t_R g955 ( 
.A(n_813),
.Y(n_955)
);

INVx1_ASAP7_75t_L g956 ( 
.A(n_699),
.Y(n_956)
);

INVx2_ASAP7_75t_L g957 ( 
.A(n_488),
.Y(n_957)
);

CKINVDCx5p33_ASAP7_75t_R g958 ( 
.A(n_99),
.Y(n_958)
);

INVx1_ASAP7_75t_L g959 ( 
.A(n_125),
.Y(n_959)
);

INVx1_ASAP7_75t_L g960 ( 
.A(n_381),
.Y(n_960)
);

CKINVDCx5p33_ASAP7_75t_R g961 ( 
.A(n_102),
.Y(n_961)
);

INVx1_ASAP7_75t_L g962 ( 
.A(n_372),
.Y(n_962)
);

CKINVDCx5p33_ASAP7_75t_R g963 ( 
.A(n_604),
.Y(n_963)
);

CKINVDCx5p33_ASAP7_75t_R g964 ( 
.A(n_491),
.Y(n_964)
);

CKINVDCx5p33_ASAP7_75t_R g965 ( 
.A(n_210),
.Y(n_965)
);

CKINVDCx5p33_ASAP7_75t_R g966 ( 
.A(n_383),
.Y(n_966)
);

CKINVDCx5p33_ASAP7_75t_R g967 ( 
.A(n_127),
.Y(n_967)
);

CKINVDCx5p33_ASAP7_75t_R g968 ( 
.A(n_648),
.Y(n_968)
);

INVx1_ASAP7_75t_L g969 ( 
.A(n_262),
.Y(n_969)
);

INVx1_ASAP7_75t_L g970 ( 
.A(n_159),
.Y(n_970)
);

INVx1_ASAP7_75t_L g971 ( 
.A(n_219),
.Y(n_971)
);

CKINVDCx5p33_ASAP7_75t_R g972 ( 
.A(n_845),
.Y(n_972)
);

HB1xp67_ASAP7_75t_L g973 ( 
.A(n_422),
.Y(n_973)
);

BUFx10_ASAP7_75t_L g974 ( 
.A(n_564),
.Y(n_974)
);

INVx1_ASAP7_75t_L g975 ( 
.A(n_227),
.Y(n_975)
);

CKINVDCx5p33_ASAP7_75t_R g976 ( 
.A(n_287),
.Y(n_976)
);

INVx1_ASAP7_75t_L g977 ( 
.A(n_210),
.Y(n_977)
);

INVx1_ASAP7_75t_L g978 ( 
.A(n_207),
.Y(n_978)
);

INVx1_ASAP7_75t_L g979 ( 
.A(n_433),
.Y(n_979)
);

CKINVDCx5p33_ASAP7_75t_R g980 ( 
.A(n_31),
.Y(n_980)
);

CKINVDCx5p33_ASAP7_75t_R g981 ( 
.A(n_205),
.Y(n_981)
);

CKINVDCx5p33_ASAP7_75t_R g982 ( 
.A(n_41),
.Y(n_982)
);

CKINVDCx5p33_ASAP7_75t_R g983 ( 
.A(n_830),
.Y(n_983)
);

CKINVDCx5p33_ASAP7_75t_R g984 ( 
.A(n_231),
.Y(n_984)
);

CKINVDCx5p33_ASAP7_75t_R g985 ( 
.A(n_407),
.Y(n_985)
);

INVx1_ASAP7_75t_L g986 ( 
.A(n_384),
.Y(n_986)
);

INVxp67_ASAP7_75t_L g987 ( 
.A(n_336),
.Y(n_987)
);

CKINVDCx5p33_ASAP7_75t_R g988 ( 
.A(n_810),
.Y(n_988)
);

CKINVDCx5p33_ASAP7_75t_R g989 ( 
.A(n_733),
.Y(n_989)
);

INVx1_ASAP7_75t_L g990 ( 
.A(n_792),
.Y(n_990)
);

CKINVDCx5p33_ASAP7_75t_R g991 ( 
.A(n_259),
.Y(n_991)
);

INVx1_ASAP7_75t_SL g992 ( 
.A(n_743),
.Y(n_992)
);

CKINVDCx5p33_ASAP7_75t_R g993 ( 
.A(n_331),
.Y(n_993)
);

BUFx10_ASAP7_75t_L g994 ( 
.A(n_608),
.Y(n_994)
);

BUFx3_ASAP7_75t_L g995 ( 
.A(n_83),
.Y(n_995)
);

CKINVDCx5p33_ASAP7_75t_R g996 ( 
.A(n_647),
.Y(n_996)
);

INVx1_ASAP7_75t_L g997 ( 
.A(n_357),
.Y(n_997)
);

CKINVDCx5p33_ASAP7_75t_R g998 ( 
.A(n_161),
.Y(n_998)
);

INVxp67_ASAP7_75t_SL g999 ( 
.A(n_358),
.Y(n_999)
);

CKINVDCx5p33_ASAP7_75t_R g1000 ( 
.A(n_9),
.Y(n_1000)
);

CKINVDCx5p33_ASAP7_75t_R g1001 ( 
.A(n_330),
.Y(n_1001)
);

CKINVDCx20_ASAP7_75t_R g1002 ( 
.A(n_417),
.Y(n_1002)
);

INVx1_ASAP7_75t_L g1003 ( 
.A(n_32),
.Y(n_1003)
);

CKINVDCx20_ASAP7_75t_R g1004 ( 
.A(n_13),
.Y(n_1004)
);

INVx1_ASAP7_75t_SL g1005 ( 
.A(n_386),
.Y(n_1005)
);

CKINVDCx5p33_ASAP7_75t_R g1006 ( 
.A(n_1),
.Y(n_1006)
);

INVx1_ASAP7_75t_L g1007 ( 
.A(n_61),
.Y(n_1007)
);

CKINVDCx5p33_ASAP7_75t_R g1008 ( 
.A(n_717),
.Y(n_1008)
);

CKINVDCx5p33_ASAP7_75t_R g1009 ( 
.A(n_131),
.Y(n_1009)
);

CKINVDCx5p33_ASAP7_75t_R g1010 ( 
.A(n_845),
.Y(n_1010)
);

INVx1_ASAP7_75t_L g1011 ( 
.A(n_178),
.Y(n_1011)
);

CKINVDCx5p33_ASAP7_75t_R g1012 ( 
.A(n_586),
.Y(n_1012)
);

CKINVDCx5p33_ASAP7_75t_R g1013 ( 
.A(n_629),
.Y(n_1013)
);

INVx1_ASAP7_75t_L g1014 ( 
.A(n_831),
.Y(n_1014)
);

INVx1_ASAP7_75t_L g1015 ( 
.A(n_80),
.Y(n_1015)
);

CKINVDCx5p33_ASAP7_75t_R g1016 ( 
.A(n_189),
.Y(n_1016)
);

BUFx2_ASAP7_75t_L g1017 ( 
.A(n_490),
.Y(n_1017)
);

INVx2_ASAP7_75t_L g1018 ( 
.A(n_478),
.Y(n_1018)
);

CKINVDCx5p33_ASAP7_75t_R g1019 ( 
.A(n_552),
.Y(n_1019)
);

CKINVDCx5p33_ASAP7_75t_R g1020 ( 
.A(n_757),
.Y(n_1020)
);

CKINVDCx5p33_ASAP7_75t_R g1021 ( 
.A(n_809),
.Y(n_1021)
);

INVx2_ASAP7_75t_L g1022 ( 
.A(n_429),
.Y(n_1022)
);

CKINVDCx5p33_ASAP7_75t_R g1023 ( 
.A(n_841),
.Y(n_1023)
);

BUFx10_ASAP7_75t_L g1024 ( 
.A(n_439),
.Y(n_1024)
);

CKINVDCx20_ASAP7_75t_R g1025 ( 
.A(n_291),
.Y(n_1025)
);

BUFx10_ASAP7_75t_L g1026 ( 
.A(n_192),
.Y(n_1026)
);

CKINVDCx5p33_ASAP7_75t_R g1027 ( 
.A(n_105),
.Y(n_1027)
);

CKINVDCx5p33_ASAP7_75t_R g1028 ( 
.A(n_119),
.Y(n_1028)
);

CKINVDCx5p33_ASAP7_75t_R g1029 ( 
.A(n_53),
.Y(n_1029)
);

INVx2_ASAP7_75t_L g1030 ( 
.A(n_808),
.Y(n_1030)
);

CKINVDCx5p33_ASAP7_75t_R g1031 ( 
.A(n_794),
.Y(n_1031)
);

CKINVDCx20_ASAP7_75t_R g1032 ( 
.A(n_801),
.Y(n_1032)
);

INVx1_ASAP7_75t_L g1033 ( 
.A(n_97),
.Y(n_1033)
);

CKINVDCx5p33_ASAP7_75t_R g1034 ( 
.A(n_26),
.Y(n_1034)
);

INVx1_ASAP7_75t_L g1035 ( 
.A(n_829),
.Y(n_1035)
);

CKINVDCx5p33_ASAP7_75t_R g1036 ( 
.A(n_584),
.Y(n_1036)
);

CKINVDCx5p33_ASAP7_75t_R g1037 ( 
.A(n_287),
.Y(n_1037)
);

CKINVDCx5p33_ASAP7_75t_R g1038 ( 
.A(n_839),
.Y(n_1038)
);

INVx1_ASAP7_75t_L g1039 ( 
.A(n_797),
.Y(n_1039)
);

CKINVDCx5p33_ASAP7_75t_R g1040 ( 
.A(n_155),
.Y(n_1040)
);

CKINVDCx5p33_ASAP7_75t_R g1041 ( 
.A(n_293),
.Y(n_1041)
);

BUFx6f_ASAP7_75t_L g1042 ( 
.A(n_60),
.Y(n_1042)
);

INVx2_ASAP7_75t_L g1043 ( 
.A(n_289),
.Y(n_1043)
);

CKINVDCx5p33_ASAP7_75t_R g1044 ( 
.A(n_733),
.Y(n_1044)
);

INVx2_ASAP7_75t_L g1045 ( 
.A(n_789),
.Y(n_1045)
);

CKINVDCx5p33_ASAP7_75t_R g1046 ( 
.A(n_602),
.Y(n_1046)
);

CKINVDCx5p33_ASAP7_75t_R g1047 ( 
.A(n_334),
.Y(n_1047)
);

CKINVDCx5p33_ASAP7_75t_R g1048 ( 
.A(n_404),
.Y(n_1048)
);

INVx2_ASAP7_75t_SL g1049 ( 
.A(n_22),
.Y(n_1049)
);

CKINVDCx5p33_ASAP7_75t_R g1050 ( 
.A(n_609),
.Y(n_1050)
);

CKINVDCx5p33_ASAP7_75t_R g1051 ( 
.A(n_37),
.Y(n_1051)
);

INVx1_ASAP7_75t_L g1052 ( 
.A(n_272),
.Y(n_1052)
);

CKINVDCx5p33_ASAP7_75t_R g1053 ( 
.A(n_123),
.Y(n_1053)
);

INVx1_ASAP7_75t_L g1054 ( 
.A(n_210),
.Y(n_1054)
);

CKINVDCx5p33_ASAP7_75t_R g1055 ( 
.A(n_482),
.Y(n_1055)
);

CKINVDCx5p33_ASAP7_75t_R g1056 ( 
.A(n_644),
.Y(n_1056)
);

INVx1_ASAP7_75t_L g1057 ( 
.A(n_456),
.Y(n_1057)
);

CKINVDCx5p33_ASAP7_75t_R g1058 ( 
.A(n_299),
.Y(n_1058)
);

BUFx10_ASAP7_75t_L g1059 ( 
.A(n_824),
.Y(n_1059)
);

INVx1_ASAP7_75t_SL g1060 ( 
.A(n_492),
.Y(n_1060)
);

INVx1_ASAP7_75t_L g1061 ( 
.A(n_97),
.Y(n_1061)
);

INVx1_ASAP7_75t_L g1062 ( 
.A(n_513),
.Y(n_1062)
);

CKINVDCx5p33_ASAP7_75t_R g1063 ( 
.A(n_823),
.Y(n_1063)
);

INVx1_ASAP7_75t_SL g1064 ( 
.A(n_59),
.Y(n_1064)
);

INVx2_ASAP7_75t_L g1065 ( 
.A(n_577),
.Y(n_1065)
);

CKINVDCx5p33_ASAP7_75t_R g1066 ( 
.A(n_383),
.Y(n_1066)
);

BUFx10_ASAP7_75t_L g1067 ( 
.A(n_793),
.Y(n_1067)
);

CKINVDCx5p33_ASAP7_75t_R g1068 ( 
.A(n_827),
.Y(n_1068)
);

CKINVDCx20_ASAP7_75t_R g1069 ( 
.A(n_832),
.Y(n_1069)
);

INVx1_ASAP7_75t_L g1070 ( 
.A(n_674),
.Y(n_1070)
);

CKINVDCx5p33_ASAP7_75t_R g1071 ( 
.A(n_126),
.Y(n_1071)
);

CKINVDCx5p33_ASAP7_75t_R g1072 ( 
.A(n_14),
.Y(n_1072)
);

CKINVDCx5p33_ASAP7_75t_R g1073 ( 
.A(n_819),
.Y(n_1073)
);

INVx2_ASAP7_75t_L g1074 ( 
.A(n_639),
.Y(n_1074)
);

INVx1_ASAP7_75t_SL g1075 ( 
.A(n_206),
.Y(n_1075)
);

INVx1_ASAP7_75t_L g1076 ( 
.A(n_401),
.Y(n_1076)
);

CKINVDCx5p33_ASAP7_75t_R g1077 ( 
.A(n_847),
.Y(n_1077)
);

CKINVDCx14_ASAP7_75t_R g1078 ( 
.A(n_786),
.Y(n_1078)
);

CKINVDCx5p33_ASAP7_75t_R g1079 ( 
.A(n_342),
.Y(n_1079)
);

CKINVDCx20_ASAP7_75t_R g1080 ( 
.A(n_738),
.Y(n_1080)
);

INVx1_ASAP7_75t_L g1081 ( 
.A(n_67),
.Y(n_1081)
);

CKINVDCx5p33_ASAP7_75t_R g1082 ( 
.A(n_640),
.Y(n_1082)
);

CKINVDCx5p33_ASAP7_75t_R g1083 ( 
.A(n_798),
.Y(n_1083)
);

INVx1_ASAP7_75t_L g1084 ( 
.A(n_43),
.Y(n_1084)
);

CKINVDCx5p33_ASAP7_75t_R g1085 ( 
.A(n_758),
.Y(n_1085)
);

CKINVDCx5p33_ASAP7_75t_R g1086 ( 
.A(n_213),
.Y(n_1086)
);

CKINVDCx5p33_ASAP7_75t_R g1087 ( 
.A(n_67),
.Y(n_1087)
);

INVx2_ASAP7_75t_L g1088 ( 
.A(n_520),
.Y(n_1088)
);

CKINVDCx5p33_ASAP7_75t_R g1089 ( 
.A(n_683),
.Y(n_1089)
);

INVx1_ASAP7_75t_SL g1090 ( 
.A(n_790),
.Y(n_1090)
);

INVx1_ASAP7_75t_L g1091 ( 
.A(n_402),
.Y(n_1091)
);

CKINVDCx5p33_ASAP7_75t_R g1092 ( 
.A(n_367),
.Y(n_1092)
);

CKINVDCx5p33_ASAP7_75t_R g1093 ( 
.A(n_419),
.Y(n_1093)
);

CKINVDCx5p33_ASAP7_75t_R g1094 ( 
.A(n_404),
.Y(n_1094)
);

CKINVDCx5p33_ASAP7_75t_R g1095 ( 
.A(n_522),
.Y(n_1095)
);

CKINVDCx5p33_ASAP7_75t_R g1096 ( 
.A(n_306),
.Y(n_1096)
);

INVx1_ASAP7_75t_L g1097 ( 
.A(n_1),
.Y(n_1097)
);

INVx1_ASAP7_75t_SL g1098 ( 
.A(n_271),
.Y(n_1098)
);

CKINVDCx5p33_ASAP7_75t_R g1099 ( 
.A(n_829),
.Y(n_1099)
);

INVx1_ASAP7_75t_L g1100 ( 
.A(n_131),
.Y(n_1100)
);

CKINVDCx5p33_ASAP7_75t_R g1101 ( 
.A(n_400),
.Y(n_1101)
);

BUFx6f_ASAP7_75t_L g1102 ( 
.A(n_546),
.Y(n_1102)
);

INVx1_ASAP7_75t_L g1103 ( 
.A(n_614),
.Y(n_1103)
);

CKINVDCx5p33_ASAP7_75t_R g1104 ( 
.A(n_5),
.Y(n_1104)
);

INVx1_ASAP7_75t_L g1105 ( 
.A(n_225),
.Y(n_1105)
);

BUFx6f_ASAP7_75t_L g1106 ( 
.A(n_196),
.Y(n_1106)
);

CKINVDCx14_ASAP7_75t_R g1107 ( 
.A(n_812),
.Y(n_1107)
);

CKINVDCx5p33_ASAP7_75t_R g1108 ( 
.A(n_606),
.Y(n_1108)
);

CKINVDCx5p33_ASAP7_75t_R g1109 ( 
.A(n_650),
.Y(n_1109)
);

INVx1_ASAP7_75t_L g1110 ( 
.A(n_741),
.Y(n_1110)
);

CKINVDCx5p33_ASAP7_75t_R g1111 ( 
.A(n_489),
.Y(n_1111)
);

CKINVDCx5p33_ASAP7_75t_R g1112 ( 
.A(n_344),
.Y(n_1112)
);

INVx1_ASAP7_75t_L g1113 ( 
.A(n_345),
.Y(n_1113)
);

INVx2_ASAP7_75t_L g1114 ( 
.A(n_490),
.Y(n_1114)
);

INVx1_ASAP7_75t_L g1115 ( 
.A(n_640),
.Y(n_1115)
);

INVx1_ASAP7_75t_L g1116 ( 
.A(n_796),
.Y(n_1116)
);

INVx2_ASAP7_75t_L g1117 ( 
.A(n_721),
.Y(n_1117)
);

CKINVDCx5p33_ASAP7_75t_R g1118 ( 
.A(n_720),
.Y(n_1118)
);

INVx1_ASAP7_75t_L g1119 ( 
.A(n_82),
.Y(n_1119)
);

CKINVDCx5p33_ASAP7_75t_R g1120 ( 
.A(n_623),
.Y(n_1120)
);

INVx1_ASAP7_75t_L g1121 ( 
.A(n_844),
.Y(n_1121)
);

INVx1_ASAP7_75t_L g1122 ( 
.A(n_377),
.Y(n_1122)
);

CKINVDCx5p33_ASAP7_75t_R g1123 ( 
.A(n_70),
.Y(n_1123)
);

INVx1_ASAP7_75t_SL g1124 ( 
.A(n_22),
.Y(n_1124)
);

INVx1_ASAP7_75t_SL g1125 ( 
.A(n_839),
.Y(n_1125)
);

CKINVDCx5p33_ASAP7_75t_R g1126 ( 
.A(n_34),
.Y(n_1126)
);

CKINVDCx5p33_ASAP7_75t_R g1127 ( 
.A(n_171),
.Y(n_1127)
);

CKINVDCx5p33_ASAP7_75t_R g1128 ( 
.A(n_119),
.Y(n_1128)
);

CKINVDCx5p33_ASAP7_75t_R g1129 ( 
.A(n_188),
.Y(n_1129)
);

HB1xp67_ASAP7_75t_L g1130 ( 
.A(n_802),
.Y(n_1130)
);

CKINVDCx5p33_ASAP7_75t_R g1131 ( 
.A(n_2),
.Y(n_1131)
);

INVx1_ASAP7_75t_L g1132 ( 
.A(n_343),
.Y(n_1132)
);

BUFx5_ASAP7_75t_L g1133 ( 
.A(n_783),
.Y(n_1133)
);

INVx1_ASAP7_75t_L g1134 ( 
.A(n_484),
.Y(n_1134)
);

CKINVDCx5p33_ASAP7_75t_R g1135 ( 
.A(n_617),
.Y(n_1135)
);

CKINVDCx5p33_ASAP7_75t_R g1136 ( 
.A(n_843),
.Y(n_1136)
);

INVx1_ASAP7_75t_L g1137 ( 
.A(n_787),
.Y(n_1137)
);

CKINVDCx20_ASAP7_75t_R g1138 ( 
.A(n_795),
.Y(n_1138)
);

CKINVDCx5p33_ASAP7_75t_R g1139 ( 
.A(n_784),
.Y(n_1139)
);

BUFx2_ASAP7_75t_L g1140 ( 
.A(n_93),
.Y(n_1140)
);

CKINVDCx20_ASAP7_75t_R g1141 ( 
.A(n_508),
.Y(n_1141)
);

CKINVDCx5p33_ASAP7_75t_R g1142 ( 
.A(n_235),
.Y(n_1142)
);

CKINVDCx5p33_ASAP7_75t_R g1143 ( 
.A(n_842),
.Y(n_1143)
);

CKINVDCx5p33_ASAP7_75t_R g1144 ( 
.A(n_381),
.Y(n_1144)
);

INVx2_ASAP7_75t_SL g1145 ( 
.A(n_632),
.Y(n_1145)
);

CKINVDCx5p33_ASAP7_75t_R g1146 ( 
.A(n_456),
.Y(n_1146)
);

CKINVDCx5p33_ASAP7_75t_R g1147 ( 
.A(n_481),
.Y(n_1147)
);

CKINVDCx5p33_ASAP7_75t_R g1148 ( 
.A(n_16),
.Y(n_1148)
);

CKINVDCx5p33_ASAP7_75t_R g1149 ( 
.A(n_764),
.Y(n_1149)
);

CKINVDCx5p33_ASAP7_75t_R g1150 ( 
.A(n_474),
.Y(n_1150)
);

CKINVDCx5p33_ASAP7_75t_R g1151 ( 
.A(n_281),
.Y(n_1151)
);

INVx1_ASAP7_75t_L g1152 ( 
.A(n_356),
.Y(n_1152)
);

BUFx10_ASAP7_75t_L g1153 ( 
.A(n_14),
.Y(n_1153)
);

CKINVDCx5p33_ASAP7_75t_R g1154 ( 
.A(n_43),
.Y(n_1154)
);

CKINVDCx5p33_ASAP7_75t_R g1155 ( 
.A(n_16),
.Y(n_1155)
);

CKINVDCx5p33_ASAP7_75t_R g1156 ( 
.A(n_204),
.Y(n_1156)
);

CKINVDCx5p33_ASAP7_75t_R g1157 ( 
.A(n_423),
.Y(n_1157)
);

CKINVDCx5p33_ASAP7_75t_R g1158 ( 
.A(n_303),
.Y(n_1158)
);

CKINVDCx5p33_ASAP7_75t_R g1159 ( 
.A(n_725),
.Y(n_1159)
);

CKINVDCx5p33_ASAP7_75t_R g1160 ( 
.A(n_201),
.Y(n_1160)
);

BUFx6f_ASAP7_75t_L g1161 ( 
.A(n_360),
.Y(n_1161)
);

CKINVDCx5p33_ASAP7_75t_R g1162 ( 
.A(n_521),
.Y(n_1162)
);

INVx1_ASAP7_75t_SL g1163 ( 
.A(n_8),
.Y(n_1163)
);

CKINVDCx5p33_ASAP7_75t_R g1164 ( 
.A(n_695),
.Y(n_1164)
);

CKINVDCx5p33_ASAP7_75t_R g1165 ( 
.A(n_658),
.Y(n_1165)
);

INVx1_ASAP7_75t_L g1166 ( 
.A(n_278),
.Y(n_1166)
);

INVx1_ASAP7_75t_L g1167 ( 
.A(n_711),
.Y(n_1167)
);

INVx1_ASAP7_75t_SL g1168 ( 
.A(n_187),
.Y(n_1168)
);

CKINVDCx5p33_ASAP7_75t_R g1169 ( 
.A(n_354),
.Y(n_1169)
);

INVx1_ASAP7_75t_SL g1170 ( 
.A(n_103),
.Y(n_1170)
);

CKINVDCx5p33_ASAP7_75t_R g1171 ( 
.A(n_596),
.Y(n_1171)
);

CKINVDCx5p33_ASAP7_75t_R g1172 ( 
.A(n_338),
.Y(n_1172)
);

CKINVDCx5p33_ASAP7_75t_R g1173 ( 
.A(n_557),
.Y(n_1173)
);

INVx1_ASAP7_75t_SL g1174 ( 
.A(n_433),
.Y(n_1174)
);

INVx1_ASAP7_75t_L g1175 ( 
.A(n_806),
.Y(n_1175)
);

BUFx6f_ASAP7_75t_L g1176 ( 
.A(n_586),
.Y(n_1176)
);

CKINVDCx5p33_ASAP7_75t_R g1177 ( 
.A(n_88),
.Y(n_1177)
);

CKINVDCx5p33_ASAP7_75t_R g1178 ( 
.A(n_160),
.Y(n_1178)
);

CKINVDCx5p33_ASAP7_75t_R g1179 ( 
.A(n_331),
.Y(n_1179)
);

INVx1_ASAP7_75t_L g1180 ( 
.A(n_775),
.Y(n_1180)
);

INVx1_ASAP7_75t_SL g1181 ( 
.A(n_814),
.Y(n_1181)
);

INVx1_ASAP7_75t_L g1182 ( 
.A(n_55),
.Y(n_1182)
);

INVx1_ASAP7_75t_L g1183 ( 
.A(n_687),
.Y(n_1183)
);

CKINVDCx5p33_ASAP7_75t_R g1184 ( 
.A(n_352),
.Y(n_1184)
);

INVx1_ASAP7_75t_L g1185 ( 
.A(n_130),
.Y(n_1185)
);

INVx2_ASAP7_75t_L g1186 ( 
.A(n_797),
.Y(n_1186)
);

CKINVDCx20_ASAP7_75t_R g1187 ( 
.A(n_162),
.Y(n_1187)
);

CKINVDCx5p33_ASAP7_75t_R g1188 ( 
.A(n_253),
.Y(n_1188)
);

CKINVDCx20_ASAP7_75t_R g1189 ( 
.A(n_814),
.Y(n_1189)
);

CKINVDCx5p33_ASAP7_75t_R g1190 ( 
.A(n_489),
.Y(n_1190)
);

CKINVDCx5p33_ASAP7_75t_R g1191 ( 
.A(n_736),
.Y(n_1191)
);

INVx1_ASAP7_75t_L g1192 ( 
.A(n_553),
.Y(n_1192)
);

INVx2_ASAP7_75t_L g1193 ( 
.A(n_498),
.Y(n_1193)
);

BUFx6f_ASAP7_75t_L g1194 ( 
.A(n_750),
.Y(n_1194)
);

BUFx6f_ASAP7_75t_L g1195 ( 
.A(n_367),
.Y(n_1195)
);

CKINVDCx5p33_ASAP7_75t_R g1196 ( 
.A(n_674),
.Y(n_1196)
);

BUFx6f_ASAP7_75t_L g1197 ( 
.A(n_281),
.Y(n_1197)
);

INVx1_ASAP7_75t_L g1198 ( 
.A(n_125),
.Y(n_1198)
);

CKINVDCx5p33_ASAP7_75t_R g1199 ( 
.A(n_521),
.Y(n_1199)
);

INVx1_ASAP7_75t_L g1200 ( 
.A(n_186),
.Y(n_1200)
);

CKINVDCx5p33_ASAP7_75t_R g1201 ( 
.A(n_407),
.Y(n_1201)
);

CKINVDCx5p33_ASAP7_75t_R g1202 ( 
.A(n_830),
.Y(n_1202)
);

INVx1_ASAP7_75t_L g1203 ( 
.A(n_508),
.Y(n_1203)
);

CKINVDCx5p33_ASAP7_75t_R g1204 ( 
.A(n_815),
.Y(n_1204)
);

CKINVDCx5p33_ASAP7_75t_R g1205 ( 
.A(n_660),
.Y(n_1205)
);

CKINVDCx5p33_ASAP7_75t_R g1206 ( 
.A(n_612),
.Y(n_1206)
);

CKINVDCx5p33_ASAP7_75t_R g1207 ( 
.A(n_787),
.Y(n_1207)
);

INVx1_ASAP7_75t_L g1208 ( 
.A(n_437),
.Y(n_1208)
);

CKINVDCx5p33_ASAP7_75t_R g1209 ( 
.A(n_800),
.Y(n_1209)
);

INVx1_ASAP7_75t_L g1210 ( 
.A(n_215),
.Y(n_1210)
);

CKINVDCx20_ASAP7_75t_R g1211 ( 
.A(n_76),
.Y(n_1211)
);

INVx1_ASAP7_75t_L g1212 ( 
.A(n_621),
.Y(n_1212)
);

CKINVDCx20_ASAP7_75t_R g1213 ( 
.A(n_831),
.Y(n_1213)
);

INVx1_ASAP7_75t_L g1214 ( 
.A(n_312),
.Y(n_1214)
);

INVx1_ASAP7_75t_L g1215 ( 
.A(n_53),
.Y(n_1215)
);

INVx1_ASAP7_75t_L g1216 ( 
.A(n_119),
.Y(n_1216)
);

CKINVDCx5p33_ASAP7_75t_R g1217 ( 
.A(n_272),
.Y(n_1217)
);

CKINVDCx5p33_ASAP7_75t_R g1218 ( 
.A(n_833),
.Y(n_1218)
);

BUFx10_ASAP7_75t_L g1219 ( 
.A(n_203),
.Y(n_1219)
);

CKINVDCx5p33_ASAP7_75t_R g1220 ( 
.A(n_192),
.Y(n_1220)
);

CKINVDCx16_ASAP7_75t_R g1221 ( 
.A(n_251),
.Y(n_1221)
);

INVx1_ASAP7_75t_L g1222 ( 
.A(n_131),
.Y(n_1222)
);

INVx1_ASAP7_75t_L g1223 ( 
.A(n_698),
.Y(n_1223)
);

CKINVDCx5p33_ASAP7_75t_R g1224 ( 
.A(n_353),
.Y(n_1224)
);

BUFx3_ASAP7_75t_L g1225 ( 
.A(n_857),
.Y(n_1225)
);

CKINVDCx20_ASAP7_75t_R g1226 ( 
.A(n_604),
.Y(n_1226)
);

INVx1_ASAP7_75t_L g1227 ( 
.A(n_374),
.Y(n_1227)
);

INVx1_ASAP7_75t_L g1228 ( 
.A(n_654),
.Y(n_1228)
);

CKINVDCx5p33_ASAP7_75t_R g1229 ( 
.A(n_86),
.Y(n_1229)
);

CKINVDCx5p33_ASAP7_75t_R g1230 ( 
.A(n_12),
.Y(n_1230)
);

INVx2_ASAP7_75t_L g1231 ( 
.A(n_410),
.Y(n_1231)
);

CKINVDCx5p33_ASAP7_75t_R g1232 ( 
.A(n_393),
.Y(n_1232)
);

CKINVDCx5p33_ASAP7_75t_R g1233 ( 
.A(n_616),
.Y(n_1233)
);

CKINVDCx5p33_ASAP7_75t_R g1234 ( 
.A(n_505),
.Y(n_1234)
);

CKINVDCx5p33_ASAP7_75t_R g1235 ( 
.A(n_481),
.Y(n_1235)
);

CKINVDCx5p33_ASAP7_75t_R g1236 ( 
.A(n_349),
.Y(n_1236)
);

INVx1_ASAP7_75t_L g1237 ( 
.A(n_64),
.Y(n_1237)
);

CKINVDCx20_ASAP7_75t_R g1238 ( 
.A(n_386),
.Y(n_1238)
);

CKINVDCx5p33_ASAP7_75t_R g1239 ( 
.A(n_805),
.Y(n_1239)
);

CKINVDCx5p33_ASAP7_75t_R g1240 ( 
.A(n_431),
.Y(n_1240)
);

CKINVDCx5p33_ASAP7_75t_R g1241 ( 
.A(n_825),
.Y(n_1241)
);

HB1xp67_ASAP7_75t_L g1242 ( 
.A(n_743),
.Y(n_1242)
);

INVxp67_ASAP7_75t_L g1243 ( 
.A(n_774),
.Y(n_1243)
);

INVxp67_ASAP7_75t_L g1244 ( 
.A(n_395),
.Y(n_1244)
);

INVx1_ASAP7_75t_L g1245 ( 
.A(n_799),
.Y(n_1245)
);

INVx1_ASAP7_75t_L g1246 ( 
.A(n_445),
.Y(n_1246)
);

CKINVDCx5p33_ASAP7_75t_R g1247 ( 
.A(n_492),
.Y(n_1247)
);

CKINVDCx5p33_ASAP7_75t_R g1248 ( 
.A(n_756),
.Y(n_1248)
);

INVx1_ASAP7_75t_L g1249 ( 
.A(n_847),
.Y(n_1249)
);

CKINVDCx20_ASAP7_75t_R g1250 ( 
.A(n_817),
.Y(n_1250)
);

INVx1_ASAP7_75t_L g1251 ( 
.A(n_486),
.Y(n_1251)
);

BUFx6f_ASAP7_75t_L g1252 ( 
.A(n_76),
.Y(n_1252)
);

CKINVDCx5p33_ASAP7_75t_R g1253 ( 
.A(n_836),
.Y(n_1253)
);

INVx2_ASAP7_75t_SL g1254 ( 
.A(n_574),
.Y(n_1254)
);

CKINVDCx5p33_ASAP7_75t_R g1255 ( 
.A(n_186),
.Y(n_1255)
);

BUFx6f_ASAP7_75t_L g1256 ( 
.A(n_90),
.Y(n_1256)
);

CKINVDCx20_ASAP7_75t_R g1257 ( 
.A(n_346),
.Y(n_1257)
);

CKINVDCx5p33_ASAP7_75t_R g1258 ( 
.A(n_618),
.Y(n_1258)
);

BUFx10_ASAP7_75t_L g1259 ( 
.A(n_55),
.Y(n_1259)
);

INVx2_ASAP7_75t_SL g1260 ( 
.A(n_509),
.Y(n_1260)
);

CKINVDCx5p33_ASAP7_75t_R g1261 ( 
.A(n_153),
.Y(n_1261)
);

INVx1_ASAP7_75t_L g1262 ( 
.A(n_137),
.Y(n_1262)
);

INVx1_ASAP7_75t_L g1263 ( 
.A(n_759),
.Y(n_1263)
);

BUFx3_ASAP7_75t_L g1264 ( 
.A(n_549),
.Y(n_1264)
);

INVx1_ASAP7_75t_L g1265 ( 
.A(n_593),
.Y(n_1265)
);

CKINVDCx5p33_ASAP7_75t_R g1266 ( 
.A(n_667),
.Y(n_1266)
);

CKINVDCx5p33_ASAP7_75t_R g1267 ( 
.A(n_533),
.Y(n_1267)
);

CKINVDCx5p33_ASAP7_75t_R g1268 ( 
.A(n_822),
.Y(n_1268)
);

INVx1_ASAP7_75t_L g1269 ( 
.A(n_693),
.Y(n_1269)
);

INVx1_ASAP7_75t_L g1270 ( 
.A(n_837),
.Y(n_1270)
);

CKINVDCx5p33_ASAP7_75t_R g1271 ( 
.A(n_86),
.Y(n_1271)
);

CKINVDCx5p33_ASAP7_75t_R g1272 ( 
.A(n_646),
.Y(n_1272)
);

INVx1_ASAP7_75t_L g1273 ( 
.A(n_77),
.Y(n_1273)
);

CKINVDCx5p33_ASAP7_75t_R g1274 ( 
.A(n_41),
.Y(n_1274)
);

CKINVDCx5p33_ASAP7_75t_R g1275 ( 
.A(n_487),
.Y(n_1275)
);

CKINVDCx5p33_ASAP7_75t_R g1276 ( 
.A(n_160),
.Y(n_1276)
);

CKINVDCx5p33_ASAP7_75t_R g1277 ( 
.A(n_559),
.Y(n_1277)
);

CKINVDCx5p33_ASAP7_75t_R g1278 ( 
.A(n_817),
.Y(n_1278)
);

BUFx5_ASAP7_75t_L g1279 ( 
.A(n_155),
.Y(n_1279)
);

CKINVDCx5p33_ASAP7_75t_R g1280 ( 
.A(n_52),
.Y(n_1280)
);

CKINVDCx5p33_ASAP7_75t_R g1281 ( 
.A(n_750),
.Y(n_1281)
);

CKINVDCx5p33_ASAP7_75t_R g1282 ( 
.A(n_515),
.Y(n_1282)
);

CKINVDCx5p33_ASAP7_75t_R g1283 ( 
.A(n_795),
.Y(n_1283)
);

CKINVDCx5p33_ASAP7_75t_R g1284 ( 
.A(n_153),
.Y(n_1284)
);

INVx2_ASAP7_75t_L g1285 ( 
.A(n_15),
.Y(n_1285)
);

CKINVDCx5p33_ASAP7_75t_R g1286 ( 
.A(n_713),
.Y(n_1286)
);

CKINVDCx5p33_ASAP7_75t_R g1287 ( 
.A(n_848),
.Y(n_1287)
);

CKINVDCx5p33_ASAP7_75t_R g1288 ( 
.A(n_756),
.Y(n_1288)
);

INVx2_ASAP7_75t_L g1289 ( 
.A(n_663),
.Y(n_1289)
);

CKINVDCx5p33_ASAP7_75t_R g1290 ( 
.A(n_605),
.Y(n_1290)
);

INVx1_ASAP7_75t_L g1291 ( 
.A(n_145),
.Y(n_1291)
);

INVx1_ASAP7_75t_L g1292 ( 
.A(n_7),
.Y(n_1292)
);

INVx2_ASAP7_75t_L g1293 ( 
.A(n_662),
.Y(n_1293)
);

BUFx3_ASAP7_75t_L g1294 ( 
.A(n_288),
.Y(n_1294)
);

INVx1_ASAP7_75t_L g1295 ( 
.A(n_835),
.Y(n_1295)
);

CKINVDCx5p33_ASAP7_75t_R g1296 ( 
.A(n_566),
.Y(n_1296)
);

CKINVDCx5p33_ASAP7_75t_R g1297 ( 
.A(n_568),
.Y(n_1297)
);

BUFx8_ASAP7_75t_SL g1298 ( 
.A(n_105),
.Y(n_1298)
);

INVx1_ASAP7_75t_L g1299 ( 
.A(n_740),
.Y(n_1299)
);

CKINVDCx5p33_ASAP7_75t_R g1300 ( 
.A(n_32),
.Y(n_1300)
);

INVx1_ASAP7_75t_L g1301 ( 
.A(n_387),
.Y(n_1301)
);

CKINVDCx16_ASAP7_75t_R g1302 ( 
.A(n_788),
.Y(n_1302)
);

INVx1_ASAP7_75t_L g1303 ( 
.A(n_581),
.Y(n_1303)
);

CKINVDCx5p33_ASAP7_75t_R g1304 ( 
.A(n_397),
.Y(n_1304)
);

INVx1_ASAP7_75t_L g1305 ( 
.A(n_581),
.Y(n_1305)
);

CKINVDCx5p33_ASAP7_75t_R g1306 ( 
.A(n_686),
.Y(n_1306)
);

CKINVDCx5p33_ASAP7_75t_R g1307 ( 
.A(n_794),
.Y(n_1307)
);

INVx1_ASAP7_75t_L g1308 ( 
.A(n_316),
.Y(n_1308)
);

CKINVDCx5p33_ASAP7_75t_R g1309 ( 
.A(n_282),
.Y(n_1309)
);

BUFx5_ASAP7_75t_L g1310 ( 
.A(n_111),
.Y(n_1310)
);

CKINVDCx5p33_ASAP7_75t_R g1311 ( 
.A(n_205),
.Y(n_1311)
);

CKINVDCx5p33_ASAP7_75t_R g1312 ( 
.A(n_816),
.Y(n_1312)
);

INVx1_ASAP7_75t_L g1313 ( 
.A(n_406),
.Y(n_1313)
);

CKINVDCx5p33_ASAP7_75t_R g1314 ( 
.A(n_186),
.Y(n_1314)
);

INVx1_ASAP7_75t_L g1315 ( 
.A(n_303),
.Y(n_1315)
);

INVx2_ASAP7_75t_L g1316 ( 
.A(n_164),
.Y(n_1316)
);

CKINVDCx5p33_ASAP7_75t_R g1317 ( 
.A(n_57),
.Y(n_1317)
);

CKINVDCx5p33_ASAP7_75t_R g1318 ( 
.A(n_162),
.Y(n_1318)
);

INVx2_ASAP7_75t_L g1319 ( 
.A(n_396),
.Y(n_1319)
);

INVx1_ASAP7_75t_SL g1320 ( 
.A(n_531),
.Y(n_1320)
);

BUFx6f_ASAP7_75t_L g1321 ( 
.A(n_825),
.Y(n_1321)
);

CKINVDCx5p33_ASAP7_75t_R g1322 ( 
.A(n_162),
.Y(n_1322)
);

INVx1_ASAP7_75t_L g1323 ( 
.A(n_408),
.Y(n_1323)
);

CKINVDCx5p33_ASAP7_75t_R g1324 ( 
.A(n_7),
.Y(n_1324)
);

INVx1_ASAP7_75t_L g1325 ( 
.A(n_667),
.Y(n_1325)
);

CKINVDCx20_ASAP7_75t_R g1326 ( 
.A(n_140),
.Y(n_1326)
);

BUFx2_ASAP7_75t_SL g1327 ( 
.A(n_244),
.Y(n_1327)
);

CKINVDCx5p33_ASAP7_75t_R g1328 ( 
.A(n_418),
.Y(n_1328)
);

CKINVDCx5p33_ASAP7_75t_R g1329 ( 
.A(n_579),
.Y(n_1329)
);

CKINVDCx5p33_ASAP7_75t_R g1330 ( 
.A(n_56),
.Y(n_1330)
);

CKINVDCx5p33_ASAP7_75t_R g1331 ( 
.A(n_51),
.Y(n_1331)
);

CKINVDCx5p33_ASAP7_75t_R g1332 ( 
.A(n_74),
.Y(n_1332)
);

CKINVDCx5p33_ASAP7_75t_R g1333 ( 
.A(n_149),
.Y(n_1333)
);

INVx2_ASAP7_75t_L g1334 ( 
.A(n_820),
.Y(n_1334)
);

CKINVDCx5p33_ASAP7_75t_R g1335 ( 
.A(n_552),
.Y(n_1335)
);

CKINVDCx5p33_ASAP7_75t_R g1336 ( 
.A(n_662),
.Y(n_1336)
);

INVx2_ASAP7_75t_SL g1337 ( 
.A(n_802),
.Y(n_1337)
);

INVx2_ASAP7_75t_SL g1338 ( 
.A(n_518),
.Y(n_1338)
);

HB1xp67_ASAP7_75t_L g1339 ( 
.A(n_368),
.Y(n_1339)
);

BUFx10_ASAP7_75t_L g1340 ( 
.A(n_679),
.Y(n_1340)
);

CKINVDCx5p33_ASAP7_75t_R g1341 ( 
.A(n_204),
.Y(n_1341)
);

INVx1_ASAP7_75t_L g1342 ( 
.A(n_785),
.Y(n_1342)
);

BUFx3_ASAP7_75t_L g1343 ( 
.A(n_687),
.Y(n_1343)
);

CKINVDCx5p33_ASAP7_75t_R g1344 ( 
.A(n_394),
.Y(n_1344)
);

CKINVDCx5p33_ASAP7_75t_R g1345 ( 
.A(n_78),
.Y(n_1345)
);

CKINVDCx5p33_ASAP7_75t_R g1346 ( 
.A(n_77),
.Y(n_1346)
);

INVx1_ASAP7_75t_L g1347 ( 
.A(n_171),
.Y(n_1347)
);

INVx1_ASAP7_75t_SL g1348 ( 
.A(n_185),
.Y(n_1348)
);

CKINVDCx5p33_ASAP7_75t_R g1349 ( 
.A(n_90),
.Y(n_1349)
);

CKINVDCx5p33_ASAP7_75t_R g1350 ( 
.A(n_161),
.Y(n_1350)
);

CKINVDCx5p33_ASAP7_75t_R g1351 ( 
.A(n_391),
.Y(n_1351)
);

CKINVDCx20_ASAP7_75t_R g1352 ( 
.A(n_818),
.Y(n_1352)
);

INVx1_ASAP7_75t_L g1353 ( 
.A(n_290),
.Y(n_1353)
);

CKINVDCx5p33_ASAP7_75t_R g1354 ( 
.A(n_624),
.Y(n_1354)
);

INVx1_ASAP7_75t_L g1355 ( 
.A(n_435),
.Y(n_1355)
);

BUFx3_ASAP7_75t_L g1356 ( 
.A(n_840),
.Y(n_1356)
);

CKINVDCx5p33_ASAP7_75t_R g1357 ( 
.A(n_747),
.Y(n_1357)
);

CKINVDCx5p33_ASAP7_75t_R g1358 ( 
.A(n_803),
.Y(n_1358)
);

BUFx6f_ASAP7_75t_L g1359 ( 
.A(n_243),
.Y(n_1359)
);

INVx1_ASAP7_75t_L g1360 ( 
.A(n_462),
.Y(n_1360)
);

CKINVDCx5p33_ASAP7_75t_R g1361 ( 
.A(n_154),
.Y(n_1361)
);

CKINVDCx5p33_ASAP7_75t_R g1362 ( 
.A(n_253),
.Y(n_1362)
);

CKINVDCx5p33_ASAP7_75t_R g1363 ( 
.A(n_804),
.Y(n_1363)
);

INVx1_ASAP7_75t_L g1364 ( 
.A(n_213),
.Y(n_1364)
);

CKINVDCx5p33_ASAP7_75t_R g1365 ( 
.A(n_445),
.Y(n_1365)
);

CKINVDCx5p33_ASAP7_75t_R g1366 ( 
.A(n_665),
.Y(n_1366)
);

INVx1_ASAP7_75t_L g1367 ( 
.A(n_313),
.Y(n_1367)
);

CKINVDCx20_ASAP7_75t_R g1368 ( 
.A(n_43),
.Y(n_1368)
);

CKINVDCx5p33_ASAP7_75t_R g1369 ( 
.A(n_161),
.Y(n_1369)
);

CKINVDCx5p33_ASAP7_75t_R g1370 ( 
.A(n_330),
.Y(n_1370)
);

CKINVDCx5p33_ASAP7_75t_R g1371 ( 
.A(n_563),
.Y(n_1371)
);

INVx1_ASAP7_75t_L g1372 ( 
.A(n_510),
.Y(n_1372)
);

INVx1_ASAP7_75t_L g1373 ( 
.A(n_62),
.Y(n_1373)
);

CKINVDCx5p33_ASAP7_75t_R g1374 ( 
.A(n_664),
.Y(n_1374)
);

INVx1_ASAP7_75t_L g1375 ( 
.A(n_372),
.Y(n_1375)
);

INVx1_ASAP7_75t_L g1376 ( 
.A(n_632),
.Y(n_1376)
);

CKINVDCx16_ASAP7_75t_R g1377 ( 
.A(n_60),
.Y(n_1377)
);

CKINVDCx5p33_ASAP7_75t_R g1378 ( 
.A(n_356),
.Y(n_1378)
);

BUFx10_ASAP7_75t_L g1379 ( 
.A(n_80),
.Y(n_1379)
);

CKINVDCx5p33_ASAP7_75t_R g1380 ( 
.A(n_791),
.Y(n_1380)
);

CKINVDCx20_ASAP7_75t_R g1381 ( 
.A(n_192),
.Y(n_1381)
);

CKINVDCx5p33_ASAP7_75t_R g1382 ( 
.A(n_231),
.Y(n_1382)
);

BUFx3_ASAP7_75t_L g1383 ( 
.A(n_94),
.Y(n_1383)
);

CKINVDCx5p33_ASAP7_75t_R g1384 ( 
.A(n_334),
.Y(n_1384)
);

CKINVDCx5p33_ASAP7_75t_R g1385 ( 
.A(n_17),
.Y(n_1385)
);

INVxp67_ASAP7_75t_SL g1386 ( 
.A(n_946),
.Y(n_1386)
);

INVxp67_ASAP7_75t_SL g1387 ( 
.A(n_946),
.Y(n_1387)
);

INVx2_ASAP7_75t_L g1388 ( 
.A(n_1133),
.Y(n_1388)
);

INVxp33_ASAP7_75t_SL g1389 ( 
.A(n_883),
.Y(n_1389)
);

INVx1_ASAP7_75t_L g1390 ( 
.A(n_950),
.Y(n_1390)
);

CKINVDCx20_ASAP7_75t_R g1391 ( 
.A(n_1298),
.Y(n_1391)
);

BUFx3_ASAP7_75t_L g1392 ( 
.A(n_897),
.Y(n_1392)
);

INVx1_ASAP7_75t_L g1393 ( 
.A(n_1140),
.Y(n_1393)
);

INVx1_ASAP7_75t_L g1394 ( 
.A(n_1049),
.Y(n_1394)
);

INVxp67_ASAP7_75t_SL g1395 ( 
.A(n_995),
.Y(n_1395)
);

INVx1_ASAP7_75t_L g1396 ( 
.A(n_1049),
.Y(n_1396)
);

CKINVDCx5p33_ASAP7_75t_R g1397 ( 
.A(n_1298),
.Y(n_1397)
);

INVxp67_ASAP7_75t_SL g1398 ( 
.A(n_995),
.Y(n_1398)
);

CKINVDCx5p33_ASAP7_75t_R g1399 ( 
.A(n_860),
.Y(n_1399)
);

INVx1_ASAP7_75t_L g1400 ( 
.A(n_873),
.Y(n_1400)
);

INVx1_ASAP7_75t_L g1401 ( 
.A(n_873),
.Y(n_1401)
);

CKINVDCx5p33_ASAP7_75t_R g1402 ( 
.A(n_860),
.Y(n_1402)
);

INVx2_ASAP7_75t_L g1403 ( 
.A(n_1133),
.Y(n_1403)
);

CKINVDCx5p33_ASAP7_75t_R g1404 ( 
.A(n_893),
.Y(n_1404)
);

INVx1_ASAP7_75t_L g1405 ( 
.A(n_912),
.Y(n_1405)
);

INVx2_ASAP7_75t_L g1406 ( 
.A(n_1133),
.Y(n_1406)
);

INVx1_ASAP7_75t_L g1407 ( 
.A(n_912),
.Y(n_1407)
);

CKINVDCx5p33_ASAP7_75t_R g1408 ( 
.A(n_893),
.Y(n_1408)
);

CKINVDCx5p33_ASAP7_75t_R g1409 ( 
.A(n_901),
.Y(n_1409)
);

INVx1_ASAP7_75t_L g1410 ( 
.A(n_923),
.Y(n_1410)
);

INVxp67_ASAP7_75t_L g1411 ( 
.A(n_1017),
.Y(n_1411)
);

INVxp67_ASAP7_75t_SL g1412 ( 
.A(n_1294),
.Y(n_1412)
);

CKINVDCx20_ASAP7_75t_R g1413 ( 
.A(n_922),
.Y(n_1413)
);

CKINVDCx16_ASAP7_75t_R g1414 ( 
.A(n_1221),
.Y(n_1414)
);

BUFx3_ASAP7_75t_L g1415 ( 
.A(n_897),
.Y(n_1415)
);

INVx1_ASAP7_75t_L g1416 ( 
.A(n_923),
.Y(n_1416)
);

INVx1_ASAP7_75t_L g1417 ( 
.A(n_1145),
.Y(n_1417)
);

CKINVDCx14_ASAP7_75t_R g1418 ( 
.A(n_908),
.Y(n_1418)
);

CKINVDCx20_ASAP7_75t_R g1419 ( 
.A(n_922),
.Y(n_1419)
);

INVx1_ASAP7_75t_L g1420 ( 
.A(n_1145),
.Y(n_1420)
);

CKINVDCx5p33_ASAP7_75t_R g1421 ( 
.A(n_901),
.Y(n_1421)
);

INVx1_ASAP7_75t_L g1422 ( 
.A(n_1254),
.Y(n_1422)
);

HB1xp67_ASAP7_75t_L g1423 ( 
.A(n_909),
.Y(n_1423)
);

INVx1_ASAP7_75t_L g1424 ( 
.A(n_1254),
.Y(n_1424)
);

INVxp33_ASAP7_75t_SL g1425 ( 
.A(n_973),
.Y(n_1425)
);

INVx1_ASAP7_75t_L g1426 ( 
.A(n_1260),
.Y(n_1426)
);

CKINVDCx5p33_ASAP7_75t_R g1427 ( 
.A(n_909),
.Y(n_1427)
);

CKINVDCx20_ASAP7_75t_R g1428 ( 
.A(n_1004),
.Y(n_1428)
);

CKINVDCx5p33_ASAP7_75t_R g1429 ( 
.A(n_910),
.Y(n_1429)
);

CKINVDCx5p33_ASAP7_75t_R g1430 ( 
.A(n_910),
.Y(n_1430)
);

CKINVDCx20_ASAP7_75t_R g1431 ( 
.A(n_1004),
.Y(n_1431)
);

BUFx6f_ASAP7_75t_L g1432 ( 
.A(n_895),
.Y(n_1432)
);

HB1xp67_ASAP7_75t_L g1433 ( 
.A(n_1370),
.Y(n_1433)
);

INVx1_ASAP7_75t_L g1434 ( 
.A(n_1260),
.Y(n_1434)
);

CKINVDCx20_ASAP7_75t_R g1435 ( 
.A(n_1025),
.Y(n_1435)
);

INVxp67_ASAP7_75t_SL g1436 ( 
.A(n_1294),
.Y(n_1436)
);

HB1xp67_ASAP7_75t_L g1437 ( 
.A(n_1370),
.Y(n_1437)
);

CKINVDCx5p33_ASAP7_75t_R g1438 ( 
.A(n_1382),
.Y(n_1438)
);

INVx2_ASAP7_75t_L g1439 ( 
.A(n_1133),
.Y(n_1439)
);

HB1xp67_ASAP7_75t_L g1440 ( 
.A(n_1382),
.Y(n_1440)
);

INVxp33_ASAP7_75t_L g1441 ( 
.A(n_1130),
.Y(n_1441)
);

INVx1_ASAP7_75t_L g1442 ( 
.A(n_1337),
.Y(n_1442)
);

INVx1_ASAP7_75t_L g1443 ( 
.A(n_1337),
.Y(n_1443)
);

INVx1_ASAP7_75t_L g1444 ( 
.A(n_1338),
.Y(n_1444)
);

BUFx6f_ASAP7_75t_L g1445 ( 
.A(n_895),
.Y(n_1445)
);

CKINVDCx20_ASAP7_75t_R g1446 ( 
.A(n_1025),
.Y(n_1446)
);

INVx1_ASAP7_75t_L g1447 ( 
.A(n_1338),
.Y(n_1447)
);

INVx1_ASAP7_75t_L g1448 ( 
.A(n_861),
.Y(n_1448)
);

CKINVDCx20_ASAP7_75t_R g1449 ( 
.A(n_1187),
.Y(n_1449)
);

INVx1_ASAP7_75t_L g1450 ( 
.A(n_862),
.Y(n_1450)
);

INVx1_ASAP7_75t_L g1451 ( 
.A(n_880),
.Y(n_1451)
);

CKINVDCx5p33_ASAP7_75t_R g1452 ( 
.A(n_1384),
.Y(n_1452)
);

INVx1_ASAP7_75t_L g1453 ( 
.A(n_890),
.Y(n_1453)
);

INVx1_ASAP7_75t_L g1454 ( 
.A(n_949),
.Y(n_1454)
);

INVxp67_ASAP7_75t_L g1455 ( 
.A(n_1242),
.Y(n_1455)
);

CKINVDCx5p33_ASAP7_75t_R g1456 ( 
.A(n_1384),
.Y(n_1456)
);

INVxp67_ASAP7_75t_SL g1457 ( 
.A(n_1383),
.Y(n_1457)
);

CKINVDCx20_ASAP7_75t_R g1458 ( 
.A(n_1187),
.Y(n_1458)
);

INVx1_ASAP7_75t_L g1459 ( 
.A(n_959),
.Y(n_1459)
);

CKINVDCx14_ASAP7_75t_R g1460 ( 
.A(n_1078),
.Y(n_1460)
);

INVx1_ASAP7_75t_L g1461 ( 
.A(n_969),
.Y(n_1461)
);

INVx1_ASAP7_75t_L g1462 ( 
.A(n_970),
.Y(n_1462)
);

INVx1_ASAP7_75t_L g1463 ( 
.A(n_971),
.Y(n_1463)
);

INVx1_ASAP7_75t_L g1464 ( 
.A(n_975),
.Y(n_1464)
);

HB1xp67_ASAP7_75t_L g1465 ( 
.A(n_1385),
.Y(n_1465)
);

INVx1_ASAP7_75t_L g1466 ( 
.A(n_977),
.Y(n_1466)
);

INVxp33_ASAP7_75t_SL g1467 ( 
.A(n_1339),
.Y(n_1467)
);

CKINVDCx5p33_ASAP7_75t_R g1468 ( 
.A(n_1385),
.Y(n_1468)
);

INVx1_ASAP7_75t_L g1469 ( 
.A(n_978),
.Y(n_1469)
);

INVxp67_ASAP7_75t_SL g1470 ( 
.A(n_1383),
.Y(n_1470)
);

HB1xp67_ASAP7_75t_L g1471 ( 
.A(n_1377),
.Y(n_1471)
);

INVx1_ASAP7_75t_L g1472 ( 
.A(n_1003),
.Y(n_1472)
);

CKINVDCx5p33_ASAP7_75t_R g1473 ( 
.A(n_1107),
.Y(n_1473)
);

BUFx6f_ASAP7_75t_SL g1474 ( 
.A(n_872),
.Y(n_1474)
);

CKINVDCx20_ASAP7_75t_R g1475 ( 
.A(n_1211),
.Y(n_1475)
);

CKINVDCx20_ASAP7_75t_R g1476 ( 
.A(n_1211),
.Y(n_1476)
);

BUFx6f_ASAP7_75t_L g1477 ( 
.A(n_895),
.Y(n_1477)
);

INVx1_ASAP7_75t_L g1478 ( 
.A(n_1007),
.Y(n_1478)
);

CKINVDCx5p33_ASAP7_75t_R g1479 ( 
.A(n_867),
.Y(n_1479)
);

INVx1_ASAP7_75t_L g1480 ( 
.A(n_1011),
.Y(n_1480)
);

CKINVDCx5p33_ASAP7_75t_R g1481 ( 
.A(n_869),
.Y(n_1481)
);

INVx1_ASAP7_75t_L g1482 ( 
.A(n_1015),
.Y(n_1482)
);

INVxp33_ASAP7_75t_SL g1483 ( 
.A(n_879),
.Y(n_1483)
);

CKINVDCx5p33_ASAP7_75t_R g1484 ( 
.A(n_884),
.Y(n_1484)
);

CKINVDCx5p33_ASAP7_75t_R g1485 ( 
.A(n_888),
.Y(n_1485)
);

INVx1_ASAP7_75t_L g1486 ( 
.A(n_1033),
.Y(n_1486)
);

CKINVDCx5p33_ASAP7_75t_R g1487 ( 
.A(n_921),
.Y(n_1487)
);

INVx1_ASAP7_75t_L g1488 ( 
.A(n_1052),
.Y(n_1488)
);

INVx1_ASAP7_75t_L g1489 ( 
.A(n_1054),
.Y(n_1489)
);

CKINVDCx5p33_ASAP7_75t_R g1490 ( 
.A(n_924),
.Y(n_1490)
);

INVx1_ASAP7_75t_L g1491 ( 
.A(n_1061),
.Y(n_1491)
);

INVx2_ASAP7_75t_L g1492 ( 
.A(n_1133),
.Y(n_1492)
);

INVx1_ASAP7_75t_L g1493 ( 
.A(n_1081),
.Y(n_1493)
);

INVx1_ASAP7_75t_L g1494 ( 
.A(n_1084),
.Y(n_1494)
);

INVxp67_ASAP7_75t_SL g1495 ( 
.A(n_987),
.Y(n_1495)
);

INVx1_ASAP7_75t_L g1496 ( 
.A(n_1097),
.Y(n_1496)
);

INVxp33_ASAP7_75t_SL g1497 ( 
.A(n_926),
.Y(n_1497)
);

CKINVDCx20_ASAP7_75t_R g1498 ( 
.A(n_1326),
.Y(n_1498)
);

CKINVDCx5p33_ASAP7_75t_R g1499 ( 
.A(n_928),
.Y(n_1499)
);

INVx1_ASAP7_75t_L g1500 ( 
.A(n_1100),
.Y(n_1500)
);

CKINVDCx20_ASAP7_75t_R g1501 ( 
.A(n_1326),
.Y(n_1501)
);

INVx1_ASAP7_75t_SL g1502 ( 
.A(n_872),
.Y(n_1502)
);

INVx1_ASAP7_75t_L g1503 ( 
.A(n_1105),
.Y(n_1503)
);

INVx1_ASAP7_75t_L g1504 ( 
.A(n_1119),
.Y(n_1504)
);

INVxp67_ASAP7_75t_L g1505 ( 
.A(n_872),
.Y(n_1505)
);

CKINVDCx5p33_ASAP7_75t_R g1506 ( 
.A(n_938),
.Y(n_1506)
);

HB1xp67_ASAP7_75t_L g1507 ( 
.A(n_945),
.Y(n_1507)
);

INVx1_ASAP7_75t_L g1508 ( 
.A(n_1166),
.Y(n_1508)
);

CKINVDCx20_ASAP7_75t_R g1509 ( 
.A(n_1381),
.Y(n_1509)
);

HB1xp67_ASAP7_75t_L g1510 ( 
.A(n_947),
.Y(n_1510)
);

INVxp67_ASAP7_75t_L g1511 ( 
.A(n_915),
.Y(n_1511)
);

CKINVDCx5p33_ASAP7_75t_R g1512 ( 
.A(n_958),
.Y(n_1512)
);

INVx1_ASAP7_75t_L g1513 ( 
.A(n_1182),
.Y(n_1513)
);

INVxp67_ASAP7_75t_L g1514 ( 
.A(n_915),
.Y(n_1514)
);

INVx1_ASAP7_75t_L g1515 ( 
.A(n_1185),
.Y(n_1515)
);

CKINVDCx20_ASAP7_75t_R g1516 ( 
.A(n_1381),
.Y(n_1516)
);

INVxp67_ASAP7_75t_SL g1517 ( 
.A(n_881),
.Y(n_1517)
);

INVx1_ASAP7_75t_L g1518 ( 
.A(n_1198),
.Y(n_1518)
);

INVx1_ASAP7_75t_L g1519 ( 
.A(n_1200),
.Y(n_1519)
);

INVx1_ASAP7_75t_L g1520 ( 
.A(n_1210),
.Y(n_1520)
);

CKINVDCx20_ASAP7_75t_R g1521 ( 
.A(n_1368),
.Y(n_1521)
);

INVx1_ASAP7_75t_L g1522 ( 
.A(n_1214),
.Y(n_1522)
);

INVx1_ASAP7_75t_L g1523 ( 
.A(n_1215),
.Y(n_1523)
);

CKINVDCx20_ASAP7_75t_R g1524 ( 
.A(n_1368),
.Y(n_1524)
);

INVx2_ASAP7_75t_L g1525 ( 
.A(n_1133),
.Y(n_1525)
);

CKINVDCx20_ASAP7_75t_R g1526 ( 
.A(n_1302),
.Y(n_1526)
);

BUFx6f_ASAP7_75t_L g1527 ( 
.A(n_895),
.Y(n_1527)
);

BUFx6f_ASAP7_75t_L g1528 ( 
.A(n_1432),
.Y(n_1528)
);

NAND2xp5_ASAP7_75t_L g1529 ( 
.A(n_1495),
.B(n_961),
.Y(n_1529)
);

INVx3_ASAP7_75t_L g1530 ( 
.A(n_1392),
.Y(n_1530)
);

INVx1_ASAP7_75t_L g1531 ( 
.A(n_1388),
.Y(n_1531)
);

AND2x4_ASAP7_75t_L g1532 ( 
.A(n_1390),
.B(n_951),
.Y(n_1532)
);

OAI22xp33_ASAP7_75t_L g1533 ( 
.A1(n_1414),
.A2(n_1441),
.B1(n_1471),
.B2(n_1397),
.Y(n_1533)
);

AND2x2_ASAP7_75t_L g1534 ( 
.A(n_1495),
.B(n_915),
.Y(n_1534)
);

AND2x2_ASAP7_75t_L g1535 ( 
.A(n_1502),
.B(n_1026),
.Y(n_1535)
);

INVx1_ASAP7_75t_L g1536 ( 
.A(n_1386),
.Y(n_1536)
);

BUFx6f_ASAP7_75t_L g1537 ( 
.A(n_1432),
.Y(n_1537)
);

AOI22xp5_ASAP7_75t_L g1538 ( 
.A1(n_1389),
.A2(n_967),
.B1(n_976),
.B2(n_965),
.Y(n_1538)
);

INVx1_ASAP7_75t_L g1539 ( 
.A(n_1386),
.Y(n_1539)
);

INVx3_ASAP7_75t_L g1540 ( 
.A(n_1415),
.Y(n_1540)
);

XOR2xp5_ASAP7_75t_L g1541 ( 
.A(n_1391),
.B(n_863),
.Y(n_1541)
);

AND2x2_ASAP7_75t_L g1542 ( 
.A(n_1455),
.B(n_1026),
.Y(n_1542)
);

INVx2_ASAP7_75t_L g1543 ( 
.A(n_1403),
.Y(n_1543)
);

INVx1_ASAP7_75t_L g1544 ( 
.A(n_1387),
.Y(n_1544)
);

INVx2_ASAP7_75t_L g1545 ( 
.A(n_1406),
.Y(n_1545)
);

INVx2_ASAP7_75t_L g1546 ( 
.A(n_1439),
.Y(n_1546)
);

INVx1_ASAP7_75t_L g1547 ( 
.A(n_1387),
.Y(n_1547)
);

AND2x4_ASAP7_75t_L g1548 ( 
.A(n_1393),
.B(n_1423),
.Y(n_1548)
);

INVx1_ASAP7_75t_L g1549 ( 
.A(n_1395),
.Y(n_1549)
);

INVx1_ASAP7_75t_L g1550 ( 
.A(n_1395),
.Y(n_1550)
);

INVx1_ASAP7_75t_L g1551 ( 
.A(n_1398),
.Y(n_1551)
);

CKINVDCx5p33_ASAP7_75t_R g1552 ( 
.A(n_1474),
.Y(n_1552)
);

INVx1_ASAP7_75t_L g1553 ( 
.A(n_1398),
.Y(n_1553)
);

BUFx3_ASAP7_75t_L g1554 ( 
.A(n_1394),
.Y(n_1554)
);

INVx2_ASAP7_75t_L g1555 ( 
.A(n_1492),
.Y(n_1555)
);

AND2x4_ASAP7_75t_L g1556 ( 
.A(n_1433),
.B(n_951),
.Y(n_1556)
);

INVx1_ASAP7_75t_L g1557 ( 
.A(n_1412),
.Y(n_1557)
);

INVx3_ASAP7_75t_L g1558 ( 
.A(n_1396),
.Y(n_1558)
);

INVx1_ASAP7_75t_L g1559 ( 
.A(n_1412),
.Y(n_1559)
);

BUFx6f_ASAP7_75t_L g1560 ( 
.A(n_1432),
.Y(n_1560)
);

INVx1_ASAP7_75t_L g1561 ( 
.A(n_1436),
.Y(n_1561)
);

BUFx6f_ASAP7_75t_L g1562 ( 
.A(n_1432),
.Y(n_1562)
);

CKINVDCx20_ASAP7_75t_R g1563 ( 
.A(n_1413),
.Y(n_1563)
);

HB1xp67_ASAP7_75t_L g1564 ( 
.A(n_1399),
.Y(n_1564)
);

INVx1_ASAP7_75t_L g1565 ( 
.A(n_1436),
.Y(n_1565)
);

CKINVDCx20_ASAP7_75t_R g1566 ( 
.A(n_1419),
.Y(n_1566)
);

BUFx6f_ASAP7_75t_L g1567 ( 
.A(n_1445),
.Y(n_1567)
);

BUFx8_ASAP7_75t_L g1568 ( 
.A(n_1474),
.Y(n_1568)
);

INVx1_ASAP7_75t_L g1569 ( 
.A(n_1457),
.Y(n_1569)
);

INVx2_ASAP7_75t_L g1570 ( 
.A(n_1525),
.Y(n_1570)
);

INVx1_ASAP7_75t_L g1571 ( 
.A(n_1457),
.Y(n_1571)
);

BUFx3_ASAP7_75t_L g1572 ( 
.A(n_1400),
.Y(n_1572)
);

NOR2xp33_ASAP7_75t_L g1573 ( 
.A(n_1505),
.B(n_1243),
.Y(n_1573)
);

INVx1_ASAP7_75t_L g1574 ( 
.A(n_1470),
.Y(n_1574)
);

NAND2xp5_ASAP7_75t_L g1575 ( 
.A(n_1511),
.B(n_980),
.Y(n_1575)
);

INVx1_ASAP7_75t_L g1576 ( 
.A(n_1470),
.Y(n_1576)
);

AND2x2_ASAP7_75t_L g1577 ( 
.A(n_1514),
.B(n_1026),
.Y(n_1577)
);

INVx1_ASAP7_75t_L g1578 ( 
.A(n_1517),
.Y(n_1578)
);

INVx3_ASAP7_75t_L g1579 ( 
.A(n_1401),
.Y(n_1579)
);

INVx1_ASAP7_75t_L g1580 ( 
.A(n_1517),
.Y(n_1580)
);

BUFx6f_ASAP7_75t_L g1581 ( 
.A(n_1445),
.Y(n_1581)
);

AND2x4_ASAP7_75t_L g1582 ( 
.A(n_1437),
.B(n_1225),
.Y(n_1582)
);

NAND2x1p5_ASAP7_75t_L g1583 ( 
.A(n_1405),
.B(n_1225),
.Y(n_1583)
);

INVx2_ASAP7_75t_L g1584 ( 
.A(n_1407),
.Y(n_1584)
);

INVx1_ASAP7_75t_L g1585 ( 
.A(n_1410),
.Y(n_1585)
);

BUFx6f_ASAP7_75t_L g1586 ( 
.A(n_1445),
.Y(n_1586)
);

INVx1_ASAP7_75t_L g1587 ( 
.A(n_1448),
.Y(n_1587)
);

INVx2_ASAP7_75t_L g1588 ( 
.A(n_1416),
.Y(n_1588)
);

INVx1_ASAP7_75t_L g1589 ( 
.A(n_1417),
.Y(n_1589)
);

INVx2_ASAP7_75t_L g1590 ( 
.A(n_1420),
.Y(n_1590)
);

OR2x2_ASAP7_75t_L g1591 ( 
.A(n_1411),
.B(n_1327),
.Y(n_1591)
);

INVx1_ASAP7_75t_L g1592 ( 
.A(n_1422),
.Y(n_1592)
);

BUFx6f_ASAP7_75t_L g1593 ( 
.A(n_1445),
.Y(n_1593)
);

CKINVDCx5p33_ASAP7_75t_R g1594 ( 
.A(n_1402),
.Y(n_1594)
);

AND2x2_ASAP7_75t_L g1595 ( 
.A(n_1440),
.B(n_1153),
.Y(n_1595)
);

AND2x2_ASAP7_75t_L g1596 ( 
.A(n_1465),
.B(n_1153),
.Y(n_1596)
);

CKINVDCx5p33_ASAP7_75t_R g1597 ( 
.A(n_1404),
.Y(n_1597)
);

BUFx3_ASAP7_75t_L g1598 ( 
.A(n_1424),
.Y(n_1598)
);

INVx2_ASAP7_75t_L g1599 ( 
.A(n_1426),
.Y(n_1599)
);

INVxp67_ASAP7_75t_L g1600 ( 
.A(n_1507),
.Y(n_1600)
);

INVx1_ASAP7_75t_L g1601 ( 
.A(n_1434),
.Y(n_1601)
);

INVx1_ASAP7_75t_L g1602 ( 
.A(n_1442),
.Y(n_1602)
);

OAI22xp5_ASAP7_75t_L g1603 ( 
.A1(n_1408),
.A2(n_1369),
.B1(n_982),
.B2(n_984),
.Y(n_1603)
);

BUFx8_ASAP7_75t_L g1604 ( 
.A(n_1483),
.Y(n_1604)
);

INVx1_ASAP7_75t_L g1605 ( 
.A(n_1443),
.Y(n_1605)
);

INVx1_ASAP7_75t_L g1606 ( 
.A(n_1444),
.Y(n_1606)
);

INVx1_ASAP7_75t_L g1607 ( 
.A(n_1447),
.Y(n_1607)
);

AND2x2_ASAP7_75t_L g1608 ( 
.A(n_1510),
.B(n_1153),
.Y(n_1608)
);

AND2x2_ASAP7_75t_L g1609 ( 
.A(n_1418),
.B(n_1219),
.Y(n_1609)
);

NAND2xp5_ASAP7_75t_L g1610 ( 
.A(n_1497),
.B(n_981),
.Y(n_1610)
);

CKINVDCx6p67_ASAP7_75t_R g1611 ( 
.A(n_1526),
.Y(n_1611)
);

CKINVDCx5p33_ASAP7_75t_R g1612 ( 
.A(n_1409),
.Y(n_1612)
);

INVx1_ASAP7_75t_L g1613 ( 
.A(n_1450),
.Y(n_1613)
);

AND2x4_ASAP7_75t_L g1614 ( 
.A(n_1421),
.B(n_1264),
.Y(n_1614)
);

CKINVDCx20_ASAP7_75t_R g1615 ( 
.A(n_1428),
.Y(n_1615)
);

CKINVDCx20_ASAP7_75t_R g1616 ( 
.A(n_1431),
.Y(n_1616)
);

INVx1_ASAP7_75t_L g1617 ( 
.A(n_1451),
.Y(n_1617)
);

AND2x4_ASAP7_75t_L g1618 ( 
.A(n_1427),
.B(n_1264),
.Y(n_1618)
);

INVx1_ASAP7_75t_L g1619 ( 
.A(n_1453),
.Y(n_1619)
);

INVx1_ASAP7_75t_L g1620 ( 
.A(n_1454),
.Y(n_1620)
);

BUFx6f_ASAP7_75t_L g1621 ( 
.A(n_1477),
.Y(n_1621)
);

AOI22xp5_ASAP7_75t_L g1622 ( 
.A1(n_1425),
.A2(n_993),
.B1(n_998),
.B2(n_991),
.Y(n_1622)
);

OAI22xp5_ASAP7_75t_SL g1623 ( 
.A1(n_1435),
.A2(n_918),
.B1(n_941),
.B2(n_863),
.Y(n_1623)
);

INVx2_ASAP7_75t_L g1624 ( 
.A(n_1459),
.Y(n_1624)
);

AND2x4_ASAP7_75t_L g1625 ( 
.A(n_1429),
.B(n_1343),
.Y(n_1625)
);

INVx1_ASAP7_75t_L g1626 ( 
.A(n_1461),
.Y(n_1626)
);

BUFx6f_ASAP7_75t_L g1627 ( 
.A(n_1477),
.Y(n_1627)
);

CKINVDCx5p33_ASAP7_75t_R g1628 ( 
.A(n_1430),
.Y(n_1628)
);

INVx3_ASAP7_75t_L g1629 ( 
.A(n_1462),
.Y(n_1629)
);

INVx2_ASAP7_75t_L g1630 ( 
.A(n_1463),
.Y(n_1630)
);

AND2x2_ASAP7_75t_L g1631 ( 
.A(n_1460),
.B(n_1219),
.Y(n_1631)
);

INVx1_ASAP7_75t_L g1632 ( 
.A(n_1464),
.Y(n_1632)
);

AND2x4_ASAP7_75t_L g1633 ( 
.A(n_1438),
.B(n_1343),
.Y(n_1633)
);

CKINVDCx20_ASAP7_75t_R g1634 ( 
.A(n_1446),
.Y(n_1634)
);

OA21x2_ASAP7_75t_L g1635 ( 
.A1(n_1466),
.A2(n_882),
.B(n_881),
.Y(n_1635)
);

NAND2xp33_ASAP7_75t_L g1636 ( 
.A(n_1469),
.B(n_1279),
.Y(n_1636)
);

CKINVDCx20_ASAP7_75t_R g1637 ( 
.A(n_1449),
.Y(n_1637)
);

CKINVDCx5p33_ASAP7_75t_R g1638 ( 
.A(n_1452),
.Y(n_1638)
);

INVx2_ASAP7_75t_L g1639 ( 
.A(n_1472),
.Y(n_1639)
);

AND2x4_ASAP7_75t_L g1640 ( 
.A(n_1456),
.B(n_1356),
.Y(n_1640)
);

HB1xp67_ASAP7_75t_L g1641 ( 
.A(n_1468),
.Y(n_1641)
);

INVx1_ASAP7_75t_L g1642 ( 
.A(n_1478),
.Y(n_1642)
);

INVx1_ASAP7_75t_L g1643 ( 
.A(n_1480),
.Y(n_1643)
);

INVx1_ASAP7_75t_L g1644 ( 
.A(n_1482),
.Y(n_1644)
);

INVx1_ASAP7_75t_L g1645 ( 
.A(n_1486),
.Y(n_1645)
);

AND2x2_ASAP7_75t_L g1646 ( 
.A(n_1479),
.B(n_1219),
.Y(n_1646)
);

INVx4_ASAP7_75t_L g1647 ( 
.A(n_1481),
.Y(n_1647)
);

INVx2_ASAP7_75t_L g1648 ( 
.A(n_1488),
.Y(n_1648)
);

AND2x2_ASAP7_75t_L g1649 ( 
.A(n_1484),
.B(n_1485),
.Y(n_1649)
);

INVx1_ASAP7_75t_L g1650 ( 
.A(n_1489),
.Y(n_1650)
);

INVx1_ASAP7_75t_L g1651 ( 
.A(n_1491),
.Y(n_1651)
);

AND2x2_ASAP7_75t_L g1652 ( 
.A(n_1487),
.B(n_1259),
.Y(n_1652)
);

INVx2_ASAP7_75t_L g1653 ( 
.A(n_1493),
.Y(n_1653)
);

INVx2_ASAP7_75t_L g1654 ( 
.A(n_1494),
.Y(n_1654)
);

CKINVDCx5p33_ASAP7_75t_R g1655 ( 
.A(n_1490),
.Y(n_1655)
);

INVx2_ASAP7_75t_L g1656 ( 
.A(n_1496),
.Y(n_1656)
);

HB1xp67_ASAP7_75t_L g1657 ( 
.A(n_1499),
.Y(n_1657)
);

CKINVDCx5p33_ASAP7_75t_R g1658 ( 
.A(n_1506),
.Y(n_1658)
);

INVx3_ASAP7_75t_L g1659 ( 
.A(n_1500),
.Y(n_1659)
);

NAND2x1_ASAP7_75t_L g1660 ( 
.A(n_1503),
.B(n_882),
.Y(n_1660)
);

INVx2_ASAP7_75t_L g1661 ( 
.A(n_1504),
.Y(n_1661)
);

NAND2xp5_ASAP7_75t_L g1662 ( 
.A(n_1508),
.B(n_1000),
.Y(n_1662)
);

NAND2xp5_ASAP7_75t_L g1663 ( 
.A(n_1513),
.B(n_1515),
.Y(n_1663)
);

INVx1_ASAP7_75t_L g1664 ( 
.A(n_1518),
.Y(n_1664)
);

BUFx6f_ASAP7_75t_L g1665 ( 
.A(n_1477),
.Y(n_1665)
);

INVx2_ASAP7_75t_L g1666 ( 
.A(n_1519),
.Y(n_1666)
);

INVx1_ASAP7_75t_L g1667 ( 
.A(n_1520),
.Y(n_1667)
);

INVx1_ASAP7_75t_L g1668 ( 
.A(n_1522),
.Y(n_1668)
);

BUFx6f_ASAP7_75t_L g1669 ( 
.A(n_1477),
.Y(n_1669)
);

INVx3_ASAP7_75t_L g1670 ( 
.A(n_1523),
.Y(n_1670)
);

INVx1_ASAP7_75t_L g1671 ( 
.A(n_1527),
.Y(n_1671)
);

HB1xp67_ASAP7_75t_L g1672 ( 
.A(n_1512),
.Y(n_1672)
);

CKINVDCx5p33_ASAP7_75t_R g1673 ( 
.A(n_1458),
.Y(n_1673)
);

CKINVDCx5p33_ASAP7_75t_R g1674 ( 
.A(n_1475),
.Y(n_1674)
);

INVx1_ASAP7_75t_L g1675 ( 
.A(n_1527),
.Y(n_1675)
);

NAND2xp5_ASAP7_75t_SL g1676 ( 
.A(n_1473),
.B(n_1467),
.Y(n_1676)
);

INVx1_ASAP7_75t_L g1677 ( 
.A(n_1527),
.Y(n_1677)
);

NAND2x1p5_ASAP7_75t_L g1678 ( 
.A(n_1527),
.B(n_1356),
.Y(n_1678)
);

AND2x2_ASAP7_75t_L g1679 ( 
.A(n_1476),
.B(n_1259),
.Y(n_1679)
);

NAND2xp5_ASAP7_75t_L g1680 ( 
.A(n_1498),
.B(n_1001),
.Y(n_1680)
);

INVx1_ASAP7_75t_L g1681 ( 
.A(n_1501),
.Y(n_1681)
);

AND2x4_ASAP7_75t_L g1682 ( 
.A(n_1509),
.B(n_877),
.Y(n_1682)
);

BUFx6f_ASAP7_75t_L g1683 ( 
.A(n_1516),
.Y(n_1683)
);

BUFx6f_ASAP7_75t_L g1684 ( 
.A(n_1521),
.Y(n_1684)
);

NAND2xp5_ASAP7_75t_L g1685 ( 
.A(n_1524),
.B(n_1006),
.Y(n_1685)
);

INVx1_ASAP7_75t_L g1686 ( 
.A(n_1386),
.Y(n_1686)
);

BUFx3_ASAP7_75t_L g1687 ( 
.A(n_1392),
.Y(n_1687)
);

OAI22xp5_ASAP7_75t_L g1688 ( 
.A1(n_1414),
.A2(n_1016),
.B1(n_1027),
.B2(n_1009),
.Y(n_1688)
);

INVx2_ASAP7_75t_L g1689 ( 
.A(n_1392),
.Y(n_1689)
);

BUFx6f_ASAP7_75t_L g1690 ( 
.A(n_1432),
.Y(n_1690)
);

AND2x4_ASAP7_75t_L g1691 ( 
.A(n_1390),
.B(n_877),
.Y(n_1691)
);

BUFx6f_ASAP7_75t_L g1692 ( 
.A(n_1432),
.Y(n_1692)
);

AND3x2_ASAP7_75t_L g1693 ( 
.A(n_1471),
.B(n_999),
.C(n_1244),
.Y(n_1693)
);

NOR2xp33_ASAP7_75t_L g1694 ( 
.A(n_1505),
.B(n_1028),
.Y(n_1694)
);

CKINVDCx5p33_ASAP7_75t_R g1695 ( 
.A(n_1474),
.Y(n_1695)
);

INVx2_ASAP7_75t_L g1696 ( 
.A(n_1392),
.Y(n_1696)
);

INVx1_ASAP7_75t_L g1697 ( 
.A(n_1386),
.Y(n_1697)
);

CKINVDCx5p33_ASAP7_75t_R g1698 ( 
.A(n_1474),
.Y(n_1698)
);

NAND2xp5_ASAP7_75t_L g1699 ( 
.A(n_1495),
.B(n_1029),
.Y(n_1699)
);

INVx2_ASAP7_75t_L g1700 ( 
.A(n_1392),
.Y(n_1700)
);

INVx1_ASAP7_75t_L g1701 ( 
.A(n_1386),
.Y(n_1701)
);

CKINVDCx5p33_ASAP7_75t_R g1702 ( 
.A(n_1474),
.Y(n_1702)
);

INVx2_ASAP7_75t_L g1703 ( 
.A(n_1392),
.Y(n_1703)
);

INVx1_ASAP7_75t_L g1704 ( 
.A(n_1386),
.Y(n_1704)
);

AND2x2_ASAP7_75t_L g1705 ( 
.A(n_1441),
.B(n_1259),
.Y(n_1705)
);

CKINVDCx5p33_ASAP7_75t_R g1706 ( 
.A(n_1474),
.Y(n_1706)
);

OAI22xp5_ASAP7_75t_L g1707 ( 
.A1(n_1414),
.A2(n_1037),
.B1(n_1040),
.B2(n_1034),
.Y(n_1707)
);

INVx3_ASAP7_75t_L g1708 ( 
.A(n_1392),
.Y(n_1708)
);

NAND2x1_ASAP7_75t_L g1709 ( 
.A(n_1448),
.B(n_887),
.Y(n_1709)
);

INVx1_ASAP7_75t_L g1710 ( 
.A(n_1386),
.Y(n_1710)
);

NOR2xp33_ASAP7_75t_L g1711 ( 
.A(n_1505),
.B(n_1041),
.Y(n_1711)
);

INVx1_ASAP7_75t_L g1712 ( 
.A(n_1386),
.Y(n_1712)
);

CKINVDCx5p33_ASAP7_75t_R g1713 ( 
.A(n_1474),
.Y(n_1713)
);

INVx3_ASAP7_75t_L g1714 ( 
.A(n_1392),
.Y(n_1714)
);

CKINVDCx5p33_ASAP7_75t_R g1715 ( 
.A(n_1474),
.Y(n_1715)
);

BUFx6f_ASAP7_75t_L g1716 ( 
.A(n_1432),
.Y(n_1716)
);

INVx1_ASAP7_75t_L g1717 ( 
.A(n_1386),
.Y(n_1717)
);

AND2x4_ASAP7_75t_L g1718 ( 
.A(n_1390),
.B(n_953),
.Y(n_1718)
);

INVx2_ASAP7_75t_L g1719 ( 
.A(n_1392),
.Y(n_1719)
);

OAI22xp5_ASAP7_75t_L g1720 ( 
.A1(n_1414),
.A2(n_1051),
.B1(n_1053),
.B2(n_1047),
.Y(n_1720)
);

NAND2xp5_ASAP7_75t_L g1721 ( 
.A(n_1495),
.B(n_1058),
.Y(n_1721)
);

INVx2_ASAP7_75t_L g1722 ( 
.A(n_1392),
.Y(n_1722)
);

INVx2_ASAP7_75t_L g1723 ( 
.A(n_1392),
.Y(n_1723)
);

NAND2xp5_ASAP7_75t_L g1724 ( 
.A(n_1495),
.B(n_1071),
.Y(n_1724)
);

INVx3_ASAP7_75t_L g1725 ( 
.A(n_1392),
.Y(n_1725)
);

BUFx6f_ASAP7_75t_L g1726 ( 
.A(n_1432),
.Y(n_1726)
);

INVxp67_ASAP7_75t_L g1727 ( 
.A(n_1471),
.Y(n_1727)
);

INVx2_ASAP7_75t_L g1728 ( 
.A(n_1392),
.Y(n_1728)
);

INVx2_ASAP7_75t_L g1729 ( 
.A(n_1392),
.Y(n_1729)
);

INVx3_ASAP7_75t_L g1730 ( 
.A(n_1392),
.Y(n_1730)
);

OAI22xp5_ASAP7_75t_SL g1731 ( 
.A1(n_1413),
.A2(n_941),
.B1(n_1002),
.B2(n_918),
.Y(n_1731)
);

OAI22xp5_ASAP7_75t_L g1732 ( 
.A1(n_1414),
.A2(n_1086),
.B1(n_1087),
.B2(n_1072),
.Y(n_1732)
);

AND2x2_ASAP7_75t_L g1733 ( 
.A(n_1441),
.B(n_1379),
.Y(n_1733)
);

INVx4_ASAP7_75t_L g1734 ( 
.A(n_1474),
.Y(n_1734)
);

INVx1_ASAP7_75t_L g1735 ( 
.A(n_1386),
.Y(n_1735)
);

AND2x4_ASAP7_75t_L g1736 ( 
.A(n_1390),
.B(n_953),
.Y(n_1736)
);

INVx3_ASAP7_75t_L g1737 ( 
.A(n_1392),
.Y(n_1737)
);

CKINVDCx8_ASAP7_75t_R g1738 ( 
.A(n_1397),
.Y(n_1738)
);

INVx2_ASAP7_75t_L g1739 ( 
.A(n_1392),
.Y(n_1739)
);

NOR2x1_ASAP7_75t_L g1740 ( 
.A(n_1390),
.B(n_1216),
.Y(n_1740)
);

NAND2x1_ASAP7_75t_L g1741 ( 
.A(n_1448),
.B(n_887),
.Y(n_1741)
);

NAND2xp33_ASAP7_75t_L g1742 ( 
.A(n_1502),
.B(n_1279),
.Y(n_1742)
);

AND2x4_ASAP7_75t_L g1743 ( 
.A(n_1390),
.B(n_957),
.Y(n_1743)
);

INVx1_ASAP7_75t_L g1744 ( 
.A(n_1386),
.Y(n_1744)
);

BUFx2_ASAP7_75t_L g1745 ( 
.A(n_1399),
.Y(n_1745)
);

OA21x2_ASAP7_75t_L g1746 ( 
.A1(n_1388),
.A2(n_911),
.B(n_903),
.Y(n_1746)
);

CKINVDCx20_ASAP7_75t_R g1747 ( 
.A(n_1413),
.Y(n_1747)
);

INVx2_ASAP7_75t_L g1748 ( 
.A(n_1392),
.Y(n_1748)
);

INVx2_ASAP7_75t_L g1749 ( 
.A(n_1635),
.Y(n_1749)
);

NAND2xp5_ASAP7_75t_L g1750 ( 
.A(n_1629),
.B(n_1279),
.Y(n_1750)
);

INVxp67_ASAP7_75t_SL g1751 ( 
.A(n_1635),
.Y(n_1751)
);

INVx1_ASAP7_75t_L g1752 ( 
.A(n_1558),
.Y(n_1752)
);

CKINVDCx5p33_ASAP7_75t_R g1753 ( 
.A(n_1568),
.Y(n_1753)
);

INVx1_ASAP7_75t_L g1754 ( 
.A(n_1558),
.Y(n_1754)
);

INVx2_ASAP7_75t_L g1755 ( 
.A(n_1746),
.Y(n_1755)
);

INVx2_ASAP7_75t_L g1756 ( 
.A(n_1746),
.Y(n_1756)
);

INVx2_ASAP7_75t_L g1757 ( 
.A(n_1579),
.Y(n_1757)
);

AND2x6_ASAP7_75t_L g1758 ( 
.A(n_1534),
.B(n_903),
.Y(n_1758)
);

BUFx10_ASAP7_75t_L g1759 ( 
.A(n_1552),
.Y(n_1759)
);

NAND2xp5_ASAP7_75t_L g1760 ( 
.A(n_1629),
.B(n_1659),
.Y(n_1760)
);

INVx2_ASAP7_75t_L g1761 ( 
.A(n_1579),
.Y(n_1761)
);

NAND2xp5_ASAP7_75t_L g1762 ( 
.A(n_1659),
.B(n_1670),
.Y(n_1762)
);

NAND2xp5_ASAP7_75t_L g1763 ( 
.A(n_1670),
.B(n_1279),
.Y(n_1763)
);

INVx1_ASAP7_75t_L g1764 ( 
.A(n_1578),
.Y(n_1764)
);

INVx1_ASAP7_75t_L g1765 ( 
.A(n_1580),
.Y(n_1765)
);

NAND2xp5_ASAP7_75t_SL g1766 ( 
.A(n_1577),
.B(n_1379),
.Y(n_1766)
);

INVx2_ASAP7_75t_L g1767 ( 
.A(n_1689),
.Y(n_1767)
);

NAND2xp5_ASAP7_75t_L g1768 ( 
.A(n_1587),
.B(n_1644),
.Y(n_1768)
);

INVx2_ASAP7_75t_L g1769 ( 
.A(n_1696),
.Y(n_1769)
);

INVx2_ASAP7_75t_L g1770 ( 
.A(n_1700),
.Y(n_1770)
);

INVx2_ASAP7_75t_L g1771 ( 
.A(n_1703),
.Y(n_1771)
);

NOR3xp33_ASAP7_75t_SL g1772 ( 
.A(n_1533),
.B(n_896),
.C(n_894),
.Y(n_1772)
);

INVx2_ASAP7_75t_L g1773 ( 
.A(n_1719),
.Y(n_1773)
);

NAND2xp5_ASAP7_75t_L g1774 ( 
.A(n_1587),
.B(n_1644),
.Y(n_1774)
);

INVx2_ASAP7_75t_L g1775 ( 
.A(n_1722),
.Y(n_1775)
);

INVx4_ASAP7_75t_L g1776 ( 
.A(n_1734),
.Y(n_1776)
);

INVx2_ASAP7_75t_L g1777 ( 
.A(n_1723),
.Y(n_1777)
);

INVx2_ASAP7_75t_SL g1778 ( 
.A(n_1705),
.Y(n_1778)
);

AOI22xp33_ASAP7_75t_L g1779 ( 
.A1(n_1536),
.A2(n_1310),
.B1(n_1279),
.B2(n_1237),
.Y(n_1779)
);

INVx2_ASAP7_75t_L g1780 ( 
.A(n_1728),
.Y(n_1780)
);

INVx1_ASAP7_75t_L g1781 ( 
.A(n_1584),
.Y(n_1781)
);

AOI21x1_ASAP7_75t_L g1782 ( 
.A1(n_1531),
.A2(n_1262),
.B(n_1222),
.Y(n_1782)
);

INVx2_ASAP7_75t_L g1783 ( 
.A(n_1729),
.Y(n_1783)
);

INVx2_ASAP7_75t_L g1784 ( 
.A(n_1739),
.Y(n_1784)
);

BUFx3_ASAP7_75t_L g1785 ( 
.A(n_1568),
.Y(n_1785)
);

NAND2xp5_ASAP7_75t_SL g1786 ( 
.A(n_1542),
.B(n_1379),
.Y(n_1786)
);

INVx1_ASAP7_75t_L g1787 ( 
.A(n_1588),
.Y(n_1787)
);

AND2x2_ASAP7_75t_L g1788 ( 
.A(n_1733),
.B(n_902),
.Y(n_1788)
);

INVx2_ASAP7_75t_L g1789 ( 
.A(n_1748),
.Y(n_1789)
);

INVx1_ASAP7_75t_L g1790 ( 
.A(n_1590),
.Y(n_1790)
);

INVx1_ASAP7_75t_L g1791 ( 
.A(n_1599),
.Y(n_1791)
);

AOI22xp33_ASAP7_75t_L g1792 ( 
.A1(n_1539),
.A2(n_1279),
.B1(n_1310),
.B2(n_1291),
.Y(n_1792)
);

CKINVDCx5p33_ASAP7_75t_R g1793 ( 
.A(n_1604),
.Y(n_1793)
);

INVx3_ASAP7_75t_L g1794 ( 
.A(n_1530),
.Y(n_1794)
);

NAND2xp5_ASAP7_75t_SL g1795 ( 
.A(n_1646),
.B(n_911),
.Y(n_1795)
);

BUFx10_ASAP7_75t_L g1796 ( 
.A(n_1695),
.Y(n_1796)
);

BUFx3_ASAP7_75t_L g1797 ( 
.A(n_1687),
.Y(n_1797)
);

INVx2_ASAP7_75t_L g1798 ( 
.A(n_1678),
.Y(n_1798)
);

NAND2xp33_ASAP7_75t_SL g1799 ( 
.A(n_1734),
.B(n_1698),
.Y(n_1799)
);

INVx2_ASAP7_75t_L g1800 ( 
.A(n_1660),
.Y(n_1800)
);

INVx2_ASAP7_75t_L g1801 ( 
.A(n_1709),
.Y(n_1801)
);

INVx2_ASAP7_75t_L g1802 ( 
.A(n_1741),
.Y(n_1802)
);

OR2x6_ASAP7_75t_L g1803 ( 
.A(n_1745),
.B(n_900),
.Y(n_1803)
);

NOR2xp33_ASAP7_75t_SL g1804 ( 
.A(n_1647),
.B(n_1096),
.Y(n_1804)
);

BUFx6f_ASAP7_75t_SL g1805 ( 
.A(n_1647),
.Y(n_1805)
);

AND2x4_ASAP7_75t_L g1806 ( 
.A(n_1535),
.B(n_864),
.Y(n_1806)
);

NAND2xp33_ASAP7_75t_L g1807 ( 
.A(n_1702),
.B(n_1706),
.Y(n_1807)
);

INVx2_ASAP7_75t_L g1808 ( 
.A(n_1624),
.Y(n_1808)
);

INVx2_ASAP7_75t_L g1809 ( 
.A(n_1630),
.Y(n_1809)
);

AOI22xp33_ASAP7_75t_L g1810 ( 
.A1(n_1544),
.A2(n_1279),
.B1(n_1310),
.B2(n_1292),
.Y(n_1810)
);

AND2x2_ASAP7_75t_L g1811 ( 
.A(n_1727),
.B(n_902),
.Y(n_1811)
);

INVx2_ASAP7_75t_L g1812 ( 
.A(n_1639),
.Y(n_1812)
);

INVx2_ASAP7_75t_L g1813 ( 
.A(n_1648),
.Y(n_1813)
);

BUFx3_ASAP7_75t_L g1814 ( 
.A(n_1604),
.Y(n_1814)
);

INVx2_ASAP7_75t_L g1815 ( 
.A(n_1653),
.Y(n_1815)
);

INVx2_ASAP7_75t_L g1816 ( 
.A(n_1654),
.Y(n_1816)
);

AND2x6_ASAP7_75t_L g1817 ( 
.A(n_1652),
.B(n_1043),
.Y(n_1817)
);

INVx1_ASAP7_75t_L g1818 ( 
.A(n_1585),
.Y(n_1818)
);

NAND2xp5_ASAP7_75t_SL g1819 ( 
.A(n_1608),
.B(n_1043),
.Y(n_1819)
);

INVxp67_ASAP7_75t_SL g1820 ( 
.A(n_1663),
.Y(n_1820)
);

NAND2xp5_ASAP7_75t_SL g1821 ( 
.A(n_1575),
.B(n_1285),
.Y(n_1821)
);

INVx2_ASAP7_75t_L g1822 ( 
.A(n_1656),
.Y(n_1822)
);

AO21x2_ASAP7_75t_L g1823 ( 
.A1(n_1636),
.A2(n_1645),
.B(n_1531),
.Y(n_1823)
);

NAND2xp5_ASAP7_75t_SL g1824 ( 
.A(n_1595),
.B(n_1596),
.Y(n_1824)
);

NAND3xp33_ASAP7_75t_L g1825 ( 
.A(n_1547),
.B(n_1123),
.C(n_1104),
.Y(n_1825)
);

INVx1_ASAP7_75t_L g1826 ( 
.A(n_1589),
.Y(n_1826)
);

INVx2_ASAP7_75t_L g1827 ( 
.A(n_1661),
.Y(n_1827)
);

INVx3_ASAP7_75t_L g1828 ( 
.A(n_1530),
.Y(n_1828)
);

OR2x6_ASAP7_75t_L g1829 ( 
.A(n_1679),
.B(n_957),
.Y(n_1829)
);

INVx1_ASAP7_75t_L g1830 ( 
.A(n_1592),
.Y(n_1830)
);

INVx1_ASAP7_75t_L g1831 ( 
.A(n_1601),
.Y(n_1831)
);

INVx3_ASAP7_75t_L g1832 ( 
.A(n_1540),
.Y(n_1832)
);

NAND2xp5_ASAP7_75t_L g1833 ( 
.A(n_1645),
.B(n_1310),
.Y(n_1833)
);

INVx1_ASAP7_75t_L g1834 ( 
.A(n_1602),
.Y(n_1834)
);

INVx2_ASAP7_75t_L g1835 ( 
.A(n_1666),
.Y(n_1835)
);

INVx4_ASAP7_75t_L g1836 ( 
.A(n_1713),
.Y(n_1836)
);

INVx2_ASAP7_75t_L g1837 ( 
.A(n_1554),
.Y(n_1837)
);

INVx2_ASAP7_75t_L g1838 ( 
.A(n_1540),
.Y(n_1838)
);

INVx2_ASAP7_75t_L g1839 ( 
.A(n_1708),
.Y(n_1839)
);

INVx2_ASAP7_75t_L g1840 ( 
.A(n_1708),
.Y(n_1840)
);

INVx1_ASAP7_75t_L g1841 ( 
.A(n_1605),
.Y(n_1841)
);

INVx2_ASAP7_75t_L g1842 ( 
.A(n_1714),
.Y(n_1842)
);

AOI22xp5_ASAP7_75t_L g1843 ( 
.A1(n_1549),
.A2(n_1127),
.B1(n_1128),
.B2(n_1126),
.Y(n_1843)
);

OAI22xp33_ASAP7_75t_SL g1844 ( 
.A1(n_1606),
.A2(n_1374),
.B1(n_1378),
.B2(n_1371),
.Y(n_1844)
);

INVx2_ASAP7_75t_L g1845 ( 
.A(n_1714),
.Y(n_1845)
);

INVx2_ASAP7_75t_L g1846 ( 
.A(n_1725),
.Y(n_1846)
);

INVx1_ASAP7_75t_L g1847 ( 
.A(n_1607),
.Y(n_1847)
);

INVx2_ASAP7_75t_L g1848 ( 
.A(n_1725),
.Y(n_1848)
);

INVx2_ASAP7_75t_L g1849 ( 
.A(n_1730),
.Y(n_1849)
);

AOI22xp33_ASAP7_75t_L g1850 ( 
.A1(n_1550),
.A2(n_1310),
.B1(n_1308),
.B2(n_1273),
.Y(n_1850)
);

NAND2xp5_ASAP7_75t_SL g1851 ( 
.A(n_1694),
.B(n_1285),
.Y(n_1851)
);

INVx2_ASAP7_75t_L g1852 ( 
.A(n_1730),
.Y(n_1852)
);

AND2x2_ASAP7_75t_L g1853 ( 
.A(n_1600),
.B(n_902),
.Y(n_1853)
);

INVx1_ASAP7_75t_SL g1854 ( 
.A(n_1649),
.Y(n_1854)
);

NAND2xp5_ASAP7_75t_L g1855 ( 
.A(n_1551),
.B(n_1310),
.Y(n_1855)
);

NAND2xp33_ASAP7_75t_L g1856 ( 
.A(n_1715),
.B(n_1310),
.Y(n_1856)
);

INVx2_ASAP7_75t_L g1857 ( 
.A(n_1737),
.Y(n_1857)
);

NAND2xp5_ASAP7_75t_L g1858 ( 
.A(n_1553),
.B(n_1133),
.Y(n_1858)
);

BUFx6f_ASAP7_75t_L g1859 ( 
.A(n_1572),
.Y(n_1859)
);

INVx2_ASAP7_75t_L g1860 ( 
.A(n_1737),
.Y(n_1860)
);

INVx2_ASAP7_75t_L g1861 ( 
.A(n_1598),
.Y(n_1861)
);

NAND2xp5_ASAP7_75t_SL g1862 ( 
.A(n_1711),
.B(n_1610),
.Y(n_1862)
);

BUFx6f_ASAP7_75t_L g1863 ( 
.A(n_1583),
.Y(n_1863)
);

BUFx8_ASAP7_75t_SL g1864 ( 
.A(n_1563),
.Y(n_1864)
);

NOR2xp33_ASAP7_75t_L g1865 ( 
.A(n_1557),
.B(n_1315),
.Y(n_1865)
);

INVx8_ASAP7_75t_L g1866 ( 
.A(n_1556),
.Y(n_1866)
);

INVx2_ASAP7_75t_L g1867 ( 
.A(n_1559),
.Y(n_1867)
);

INVx2_ASAP7_75t_L g1868 ( 
.A(n_1561),
.Y(n_1868)
);

INVx2_ASAP7_75t_L g1869 ( 
.A(n_1565),
.Y(n_1869)
);

INVx1_ASAP7_75t_L g1870 ( 
.A(n_1569),
.Y(n_1870)
);

NAND2xp5_ASAP7_75t_L g1871 ( 
.A(n_1571),
.B(n_1129),
.Y(n_1871)
);

INVx1_ASAP7_75t_L g1872 ( 
.A(n_1574),
.Y(n_1872)
);

INVx3_ASAP7_75t_L g1873 ( 
.A(n_1576),
.Y(n_1873)
);

INVx2_ASAP7_75t_L g1874 ( 
.A(n_1686),
.Y(n_1874)
);

INVx2_ASAP7_75t_L g1875 ( 
.A(n_1697),
.Y(n_1875)
);

INVx1_ASAP7_75t_L g1876 ( 
.A(n_1701),
.Y(n_1876)
);

INVx1_ASAP7_75t_L g1877 ( 
.A(n_1704),
.Y(n_1877)
);

NAND2xp5_ASAP7_75t_SL g1878 ( 
.A(n_1529),
.B(n_1316),
.Y(n_1878)
);

NOR3xp33_ASAP7_75t_L g1879 ( 
.A(n_1603),
.B(n_1064),
.C(n_885),
.Y(n_1879)
);

NAND2xp5_ASAP7_75t_SL g1880 ( 
.A(n_1699),
.B(n_1316),
.Y(n_1880)
);

INVx1_ASAP7_75t_L g1881 ( 
.A(n_1710),
.Y(n_1881)
);

BUFx3_ASAP7_75t_L g1882 ( 
.A(n_1655),
.Y(n_1882)
);

INVx2_ASAP7_75t_L g1883 ( 
.A(n_1712),
.Y(n_1883)
);

INVx2_ASAP7_75t_L g1884 ( 
.A(n_1717),
.Y(n_1884)
);

NOR2xp33_ASAP7_75t_L g1885 ( 
.A(n_1735),
.B(n_1347),
.Y(n_1885)
);

NOR2x1p5_ASAP7_75t_L g1886 ( 
.A(n_1611),
.B(n_1658),
.Y(n_1886)
);

NAND2xp5_ASAP7_75t_L g1887 ( 
.A(n_1744),
.B(n_1131),
.Y(n_1887)
);

AOI21x1_ASAP7_75t_L g1888 ( 
.A1(n_1543),
.A2(n_1364),
.B(n_1353),
.Y(n_1888)
);

INVx1_ASAP7_75t_L g1889 ( 
.A(n_1613),
.Y(n_1889)
);

AND2x6_ASAP7_75t_L g1890 ( 
.A(n_1609),
.B(n_1042),
.Y(n_1890)
);

NAND2xp33_ASAP7_75t_L g1891 ( 
.A(n_1617),
.B(n_1042),
.Y(n_1891)
);

INVx1_ASAP7_75t_L g1892 ( 
.A(n_1619),
.Y(n_1892)
);

NAND2xp5_ASAP7_75t_L g1893 ( 
.A(n_1721),
.B(n_1724),
.Y(n_1893)
);

NOR2xp33_ASAP7_75t_L g1894 ( 
.A(n_1662),
.B(n_1367),
.Y(n_1894)
);

INVx2_ASAP7_75t_SL g1895 ( 
.A(n_1631),
.Y(n_1895)
);

INVx4_ASAP7_75t_L g1896 ( 
.A(n_1556),
.Y(n_1896)
);

INVx1_ASAP7_75t_L g1897 ( 
.A(n_1620),
.Y(n_1897)
);

INVx1_ASAP7_75t_L g1898 ( 
.A(n_1626),
.Y(n_1898)
);

INVx2_ASAP7_75t_L g1899 ( 
.A(n_1632),
.Y(n_1899)
);

AND2x2_ASAP7_75t_L g1900 ( 
.A(n_1548),
.B(n_974),
.Y(n_1900)
);

INVx2_ASAP7_75t_L g1901 ( 
.A(n_1642),
.Y(n_1901)
);

INVx1_ASAP7_75t_L g1902 ( 
.A(n_1643),
.Y(n_1902)
);

INVx2_ASAP7_75t_L g1903 ( 
.A(n_1650),
.Y(n_1903)
);

AND2x2_ASAP7_75t_L g1904 ( 
.A(n_1548),
.B(n_974),
.Y(n_1904)
);

INVx1_ASAP7_75t_L g1905 ( 
.A(n_1651),
.Y(n_1905)
);

INVx4_ASAP7_75t_L g1906 ( 
.A(n_1582),
.Y(n_1906)
);

INVx1_ASAP7_75t_L g1907 ( 
.A(n_1664),
.Y(n_1907)
);

INVx1_ASAP7_75t_L g1908 ( 
.A(n_1667),
.Y(n_1908)
);

INVx2_ASAP7_75t_L g1909 ( 
.A(n_1668),
.Y(n_1909)
);

INVx3_ASAP7_75t_L g1910 ( 
.A(n_1532),
.Y(n_1910)
);

BUFx6f_ASAP7_75t_L g1911 ( 
.A(n_1528),
.Y(n_1911)
);

INVx2_ASAP7_75t_L g1912 ( 
.A(n_1545),
.Y(n_1912)
);

INVx3_ASAP7_75t_L g1913 ( 
.A(n_1532),
.Y(n_1913)
);

INVx2_ASAP7_75t_L g1914 ( 
.A(n_1546),
.Y(n_1914)
);

AOI22xp33_ASAP7_75t_SL g1915 ( 
.A1(n_1623),
.A2(n_1032),
.B1(n_1069),
.B2(n_1002),
.Y(n_1915)
);

INVx1_ASAP7_75t_L g1916 ( 
.A(n_1691),
.Y(n_1916)
);

INVx6_ASAP7_75t_L g1917 ( 
.A(n_1582),
.Y(n_1917)
);

INVx1_ASAP7_75t_L g1918 ( 
.A(n_1691),
.Y(n_1918)
);

NOR2xp33_ASAP7_75t_L g1919 ( 
.A(n_1573),
.B(n_1373),
.Y(n_1919)
);

BUFx6f_ASAP7_75t_L g1920 ( 
.A(n_1528),
.Y(n_1920)
);

AO21x2_ASAP7_75t_L g1921 ( 
.A1(n_1742),
.A2(n_874),
.B(n_868),
.Y(n_1921)
);

INVx1_ASAP7_75t_L g1922 ( 
.A(n_1718),
.Y(n_1922)
);

NAND2xp5_ASAP7_75t_L g1923 ( 
.A(n_1740),
.B(n_1148),
.Y(n_1923)
);

NOR2xp33_ASAP7_75t_L g1924 ( 
.A(n_1614),
.B(n_876),
.Y(n_1924)
);

INVx2_ASAP7_75t_L g1925 ( 
.A(n_1555),
.Y(n_1925)
);

AOI22xp5_ASAP7_75t_L g1926 ( 
.A1(n_1538),
.A2(n_1151),
.B1(n_1154),
.B2(n_1142),
.Y(n_1926)
);

INVx2_ASAP7_75t_L g1927 ( 
.A(n_1570),
.Y(n_1927)
);

INVx1_ASAP7_75t_L g1928 ( 
.A(n_1718),
.Y(n_1928)
);

INVx2_ASAP7_75t_SL g1929 ( 
.A(n_1591),
.Y(n_1929)
);

INVx1_ASAP7_75t_L g1930 ( 
.A(n_1736),
.Y(n_1930)
);

NAND2xp5_ASAP7_75t_L g1931 ( 
.A(n_1736),
.B(n_1155),
.Y(n_1931)
);

NAND2xp5_ASAP7_75t_L g1932 ( 
.A(n_1743),
.B(n_1156),
.Y(n_1932)
);

INVx1_ASAP7_75t_L g1933 ( 
.A(n_1743),
.Y(n_1933)
);

AOI22xp33_ASAP7_75t_L g1934 ( 
.A1(n_1682),
.A2(n_1106),
.B1(n_1197),
.B2(n_1042),
.Y(n_1934)
);

NAND2xp5_ASAP7_75t_SL g1935 ( 
.A(n_1614),
.B(n_1158),
.Y(n_1935)
);

NAND2xp33_ASAP7_75t_L g1936 ( 
.A(n_1594),
.B(n_1042),
.Y(n_1936)
);

INVx1_ASAP7_75t_L g1937 ( 
.A(n_1618),
.Y(n_1937)
);

INVx1_ASAP7_75t_L g1938 ( 
.A(n_1618),
.Y(n_1938)
);

AOI22xp5_ASAP7_75t_L g1939 ( 
.A1(n_1622),
.A2(n_1172),
.B1(n_1177),
.B2(n_1160),
.Y(n_1939)
);

INVx1_ASAP7_75t_L g1940 ( 
.A(n_1625),
.Y(n_1940)
);

INVx2_ASAP7_75t_L g1941 ( 
.A(n_1671),
.Y(n_1941)
);

INVx1_ASAP7_75t_L g1942 ( 
.A(n_1625),
.Y(n_1942)
);

CKINVDCx5p33_ASAP7_75t_R g1943 ( 
.A(n_1673),
.Y(n_1943)
);

INVx2_ASAP7_75t_L g1944 ( 
.A(n_1675),
.Y(n_1944)
);

INVx1_ASAP7_75t_L g1945 ( 
.A(n_1633),
.Y(n_1945)
);

INVx2_ASAP7_75t_L g1946 ( 
.A(n_1677),
.Y(n_1946)
);

INVx2_ASAP7_75t_L g1947 ( 
.A(n_1528),
.Y(n_1947)
);

BUFx3_ASAP7_75t_L g1948 ( 
.A(n_1738),
.Y(n_1948)
);

AOI22xp5_ASAP7_75t_L g1949 ( 
.A1(n_1688),
.A2(n_1179),
.B1(n_1188),
.B2(n_1178),
.Y(n_1949)
);

NAND2xp5_ASAP7_75t_SL g1950 ( 
.A(n_1633),
.B(n_1217),
.Y(n_1950)
);

NAND2xp5_ASAP7_75t_L g1951 ( 
.A(n_1640),
.B(n_1229),
.Y(n_1951)
);

OR2x6_ASAP7_75t_L g1952 ( 
.A(n_1657),
.B(n_1018),
.Y(n_1952)
);

AOI22xp33_ASAP7_75t_L g1953 ( 
.A1(n_1682),
.A2(n_1197),
.B1(n_1252),
.B2(n_1106),
.Y(n_1953)
);

BUFx3_ASAP7_75t_L g1954 ( 
.A(n_1597),
.Y(n_1954)
);

INVx1_ASAP7_75t_L g1955 ( 
.A(n_1640),
.Y(n_1955)
);

AND2x6_ASAP7_75t_L g1956 ( 
.A(n_1680),
.B(n_1106),
.Y(n_1956)
);

INVx2_ASAP7_75t_L g1957 ( 
.A(n_1537),
.Y(n_1957)
);

NOR2xp33_ASAP7_75t_L g1958 ( 
.A(n_1676),
.B(n_892),
.Y(n_1958)
);

NOR2xp33_ASAP7_75t_L g1959 ( 
.A(n_1707),
.B(n_917),
.Y(n_1959)
);

INVx2_ASAP7_75t_L g1960 ( 
.A(n_1537),
.Y(n_1960)
);

NAND2xp5_ASAP7_75t_SL g1961 ( 
.A(n_1720),
.B(n_1732),
.Y(n_1961)
);

INVx2_ASAP7_75t_L g1962 ( 
.A(n_1537),
.Y(n_1962)
);

INVx2_ASAP7_75t_L g1963 ( 
.A(n_1560),
.Y(n_1963)
);

INVx2_ASAP7_75t_L g1964 ( 
.A(n_1560),
.Y(n_1964)
);

INVx3_ASAP7_75t_L g1965 ( 
.A(n_1693),
.Y(n_1965)
);

INVx2_ASAP7_75t_L g1966 ( 
.A(n_1560),
.Y(n_1966)
);

INVx2_ASAP7_75t_SL g1967 ( 
.A(n_1564),
.Y(n_1967)
);

INVx2_ASAP7_75t_L g1968 ( 
.A(n_1562),
.Y(n_1968)
);

BUFx6f_ASAP7_75t_SL g1969 ( 
.A(n_1683),
.Y(n_1969)
);

INVx3_ASAP7_75t_L g1970 ( 
.A(n_1562),
.Y(n_1970)
);

HB1xp67_ASAP7_75t_L g1971 ( 
.A(n_1641),
.Y(n_1971)
);

BUFx3_ASAP7_75t_L g1972 ( 
.A(n_1612),
.Y(n_1972)
);

NOR2xp33_ASAP7_75t_L g1973 ( 
.A(n_1672),
.B(n_933),
.Y(n_1973)
);

OR2x2_ASAP7_75t_L g1974 ( 
.A(n_1685),
.B(n_894),
.Y(n_1974)
);

NAND2xp33_ASAP7_75t_L g1975 ( 
.A(n_1628),
.B(n_1106),
.Y(n_1975)
);

BUFx3_ASAP7_75t_L g1976 ( 
.A(n_1638),
.Y(n_1976)
);

INVx2_ASAP7_75t_L g1977 ( 
.A(n_1562),
.Y(n_1977)
);

INVx1_ASAP7_75t_L g1978 ( 
.A(n_1567),
.Y(n_1978)
);

NAND2xp5_ASAP7_75t_SL g1979 ( 
.A(n_1683),
.B(n_1220),
.Y(n_1979)
);

NOR2xp33_ASAP7_75t_SL g1980 ( 
.A(n_1567),
.B(n_1230),
.Y(n_1980)
);

INVx2_ASAP7_75t_L g1981 ( 
.A(n_1567),
.Y(n_1981)
);

BUFx3_ASAP7_75t_L g1982 ( 
.A(n_1683),
.Y(n_1982)
);

INVx2_ASAP7_75t_L g1983 ( 
.A(n_1581),
.Y(n_1983)
);

BUFx6f_ASAP7_75t_L g1984 ( 
.A(n_1581),
.Y(n_1984)
);

NAND2xp5_ASAP7_75t_SL g1985 ( 
.A(n_1684),
.B(n_1255),
.Y(n_1985)
);

INVx1_ASAP7_75t_L g1986 ( 
.A(n_1581),
.Y(n_1986)
);

INVx1_ASAP7_75t_L g1987 ( 
.A(n_1586),
.Y(n_1987)
);

INVx2_ASAP7_75t_L g1988 ( 
.A(n_1586),
.Y(n_1988)
);

NAND2xp5_ASAP7_75t_SL g1989 ( 
.A(n_1684),
.B(n_1361),
.Y(n_1989)
);

INVx2_ASAP7_75t_L g1990 ( 
.A(n_1586),
.Y(n_1990)
);

AND2x2_ASAP7_75t_L g1991 ( 
.A(n_1684),
.B(n_974),
.Y(n_1991)
);

INVx1_ASAP7_75t_L g1992 ( 
.A(n_1593),
.Y(n_1992)
);

NAND2xp5_ASAP7_75t_L g1993 ( 
.A(n_1593),
.B(n_1362),
.Y(n_1993)
);

NAND2xp5_ASAP7_75t_L g1994 ( 
.A(n_1593),
.B(n_1261),
.Y(n_1994)
);

INVx1_ASAP7_75t_L g1995 ( 
.A(n_1621),
.Y(n_1995)
);

NAND2xp33_ASAP7_75t_R g1996 ( 
.A(n_1674),
.B(n_896),
.Y(n_1996)
);

NAND2xp5_ASAP7_75t_SL g1997 ( 
.A(n_1681),
.B(n_1271),
.Y(n_1997)
);

INVx1_ASAP7_75t_L g1998 ( 
.A(n_1621),
.Y(n_1998)
);

INVx2_ASAP7_75t_SL g1999 ( 
.A(n_1566),
.Y(n_1999)
);

OAI22xp33_ASAP7_75t_L g2000 ( 
.A1(n_1615),
.A2(n_1276),
.B1(n_1280),
.B2(n_1274),
.Y(n_2000)
);

NOR2xp33_ASAP7_75t_L g2001 ( 
.A(n_1621),
.B(n_935),
.Y(n_2001)
);

BUFx6f_ASAP7_75t_L g2002 ( 
.A(n_1627),
.Y(n_2002)
);

NOR2x1p5_ASAP7_75t_L g2003 ( 
.A(n_1541),
.B(n_898),
.Y(n_2003)
);

NAND2xp5_ASAP7_75t_SL g2004 ( 
.A(n_1627),
.B(n_1284),
.Y(n_2004)
);

CKINVDCx5p33_ASAP7_75t_R g2005 ( 
.A(n_1616),
.Y(n_2005)
);

INVx2_ASAP7_75t_L g2006 ( 
.A(n_1627),
.Y(n_2006)
);

INVx2_ASAP7_75t_L g2007 ( 
.A(n_1665),
.Y(n_2007)
);

INVx1_ASAP7_75t_SL g2008 ( 
.A(n_1634),
.Y(n_2008)
);

INVx4_ASAP7_75t_L g2009 ( 
.A(n_1665),
.Y(n_2009)
);

NAND3xp33_ASAP7_75t_L g2010 ( 
.A(n_1665),
.B(n_1309),
.C(n_1300),
.Y(n_2010)
);

NOR2xp33_ASAP7_75t_L g2011 ( 
.A(n_1669),
.B(n_936),
.Y(n_2011)
);

NAND2xp5_ASAP7_75t_L g2012 ( 
.A(n_1669),
.B(n_1314),
.Y(n_2012)
);

INVx2_ASAP7_75t_SL g2013 ( 
.A(n_1637),
.Y(n_2013)
);

INVx2_ASAP7_75t_L g2014 ( 
.A(n_1669),
.Y(n_2014)
);

AND2x4_ASAP7_75t_L g2015 ( 
.A(n_1747),
.B(n_943),
.Y(n_2015)
);

INVx1_ASAP7_75t_L g2016 ( 
.A(n_1690),
.Y(n_2016)
);

INVx2_ASAP7_75t_L g2017 ( 
.A(n_1690),
.Y(n_2017)
);

NAND2xp5_ASAP7_75t_L g2018 ( 
.A(n_1690),
.B(n_1311),
.Y(n_2018)
);

CKINVDCx5p33_ASAP7_75t_R g2019 ( 
.A(n_1731),
.Y(n_2019)
);

NOR2xp33_ASAP7_75t_L g2020 ( 
.A(n_1692),
.B(n_944),
.Y(n_2020)
);

INVx1_ASAP7_75t_L g2021 ( 
.A(n_1692),
.Y(n_2021)
);

INVx3_ASAP7_75t_L g2022 ( 
.A(n_1692),
.Y(n_2022)
);

BUFx6f_ASAP7_75t_SL g2023 ( 
.A(n_1716),
.Y(n_2023)
);

INVx3_ASAP7_75t_L g2024 ( 
.A(n_1716),
.Y(n_2024)
);

INVx2_ASAP7_75t_L g2025 ( 
.A(n_1716),
.Y(n_2025)
);

AOI22xp33_ASAP7_75t_L g2026 ( 
.A1(n_1726),
.A2(n_1252),
.B1(n_1256),
.B2(n_1197),
.Y(n_2026)
);

BUFx6f_ASAP7_75t_L g2027 ( 
.A(n_1726),
.Y(n_2027)
);

NAND3xp33_ASAP7_75t_L g2028 ( 
.A(n_1726),
.B(n_1318),
.C(n_1317),
.Y(n_2028)
);

NAND2xp5_ASAP7_75t_L g2029 ( 
.A(n_1629),
.B(n_1322),
.Y(n_2029)
);

INVx2_ASAP7_75t_L g2030 ( 
.A(n_1635),
.Y(n_2030)
);

NOR2xp33_ASAP7_75t_L g2031 ( 
.A(n_1536),
.B(n_948),
.Y(n_2031)
);

INVx1_ASAP7_75t_L g2032 ( 
.A(n_1558),
.Y(n_2032)
);

AND2x6_ASAP7_75t_L g2033 ( 
.A(n_1534),
.B(n_1197),
.Y(n_2033)
);

INVx2_ASAP7_75t_SL g2034 ( 
.A(n_1705),
.Y(n_2034)
);

NAND2xp5_ASAP7_75t_L g2035 ( 
.A(n_1629),
.B(n_1324),
.Y(n_2035)
);

NAND2xp5_ASAP7_75t_L g2036 ( 
.A(n_1629),
.B(n_1330),
.Y(n_2036)
);

INVx1_ASAP7_75t_L g2037 ( 
.A(n_1558),
.Y(n_2037)
);

CKINVDCx11_ASAP7_75t_R g2038 ( 
.A(n_1738),
.Y(n_2038)
);

INVx3_ASAP7_75t_L g2039 ( 
.A(n_1558),
.Y(n_2039)
);

INVx2_ASAP7_75t_L g2040 ( 
.A(n_1635),
.Y(n_2040)
);

BUFx10_ASAP7_75t_L g2041 ( 
.A(n_1552),
.Y(n_2041)
);

BUFx3_ASAP7_75t_L g2042 ( 
.A(n_1568),
.Y(n_2042)
);

NAND2xp5_ASAP7_75t_L g2043 ( 
.A(n_1629),
.B(n_1331),
.Y(n_2043)
);

BUFx6f_ASAP7_75t_L g2044 ( 
.A(n_1635),
.Y(n_2044)
);

INVx1_ASAP7_75t_L g2045 ( 
.A(n_1558),
.Y(n_2045)
);

INVx2_ASAP7_75t_L g2046 ( 
.A(n_1635),
.Y(n_2046)
);

BUFx3_ASAP7_75t_L g2047 ( 
.A(n_1568),
.Y(n_2047)
);

NAND2xp5_ASAP7_75t_SL g2048 ( 
.A(n_1804),
.B(n_1820),
.Y(n_2048)
);

NAND2xp5_ASAP7_75t_SL g2049 ( 
.A(n_1804),
.B(n_1332),
.Y(n_2049)
);

NAND2xp5_ASAP7_75t_L g2050 ( 
.A(n_1820),
.B(n_1333),
.Y(n_2050)
);

INVx2_ASAP7_75t_L g2051 ( 
.A(n_1873),
.Y(n_2051)
);

NAND2xp5_ASAP7_75t_SL g2052 ( 
.A(n_1859),
.B(n_1350),
.Y(n_2052)
);

NAND2xp5_ASAP7_75t_L g2053 ( 
.A(n_1893),
.B(n_2029),
.Y(n_2053)
);

NAND2xp5_ASAP7_75t_SL g2054 ( 
.A(n_1859),
.B(n_1341),
.Y(n_2054)
);

AND3x4_ASAP7_75t_L g2055 ( 
.A(n_1814),
.B(n_1352),
.C(n_1069),
.Y(n_2055)
);

NOR2xp33_ASAP7_75t_L g2056 ( 
.A(n_1929),
.B(n_898),
.Y(n_2056)
);

NAND2xp5_ASAP7_75t_L g2057 ( 
.A(n_1893),
.B(n_1345),
.Y(n_2057)
);

NAND2xp5_ASAP7_75t_L g2058 ( 
.A(n_1768),
.B(n_1346),
.Y(n_2058)
);

NOR2xp33_ASAP7_75t_L g2059 ( 
.A(n_1896),
.B(n_899),
.Y(n_2059)
);

INVx1_ASAP7_75t_L g2060 ( 
.A(n_1768),
.Y(n_2060)
);

NAND2xp5_ASAP7_75t_SL g2061 ( 
.A(n_1859),
.B(n_1349),
.Y(n_2061)
);

AOI22xp5_ASAP7_75t_L g2062 ( 
.A1(n_1806),
.A2(n_905),
.B1(n_906),
.B2(n_899),
.Y(n_2062)
);

HB1xp67_ASAP7_75t_L g2063 ( 
.A(n_1971),
.Y(n_2063)
);

AOI22xp5_ASAP7_75t_L g2064 ( 
.A1(n_1806),
.A2(n_906),
.B1(n_907),
.B2(n_905),
.Y(n_2064)
);

NAND2xp5_ASAP7_75t_L g2065 ( 
.A(n_1774),
.B(n_1075),
.Y(n_2065)
);

NAND2xp5_ASAP7_75t_SL g2066 ( 
.A(n_1967),
.B(n_1854),
.Y(n_2066)
);

CKINVDCx5p33_ASAP7_75t_R g2067 ( 
.A(n_1864),
.Y(n_2067)
);

INVx1_ASAP7_75t_L g2068 ( 
.A(n_1774),
.Y(n_2068)
);

AND2x4_ASAP7_75t_L g2069 ( 
.A(n_1776),
.B(n_954),
.Y(n_2069)
);

INVx1_ASAP7_75t_L g2070 ( 
.A(n_1760),
.Y(n_2070)
);

INVx4_ASAP7_75t_L g2071 ( 
.A(n_1805),
.Y(n_2071)
);

INVxp33_ASAP7_75t_L g2072 ( 
.A(n_1971),
.Y(n_2072)
);

INVx2_ASAP7_75t_SL g2073 ( 
.A(n_1866),
.Y(n_2073)
);

INVx1_ASAP7_75t_L g2074 ( 
.A(n_1760),
.Y(n_2074)
);

INVx1_ASAP7_75t_L g2075 ( 
.A(n_1762),
.Y(n_2075)
);

NAND2xp33_ASAP7_75t_L g2076 ( 
.A(n_2044),
.B(n_1374),
.Y(n_2076)
);

BUFx3_ASAP7_75t_L g2077 ( 
.A(n_1785),
.Y(n_2077)
);

AND2x2_ASAP7_75t_L g2078 ( 
.A(n_1854),
.B(n_1032),
.Y(n_2078)
);

OAI22xp33_ASAP7_75t_L g2079 ( 
.A1(n_2000),
.A2(n_1138),
.B1(n_1141),
.B2(n_1080),
.Y(n_2079)
);

AND2x2_ASAP7_75t_L g2080 ( 
.A(n_1843),
.B(n_1080),
.Y(n_2080)
);

NAND3xp33_ASAP7_75t_L g2081 ( 
.A(n_1934),
.B(n_1256),
.C(n_1252),
.Y(n_2081)
);

BUFx6f_ASAP7_75t_SL g2082 ( 
.A(n_2042),
.Y(n_2082)
);

NOR2xp33_ASAP7_75t_SL g2083 ( 
.A(n_1751),
.B(n_1749),
.Y(n_2083)
);

NAND2xp5_ASAP7_75t_L g2084 ( 
.A(n_2029),
.B(n_1098),
.Y(n_2084)
);

NAND2xp5_ASAP7_75t_L g2085 ( 
.A(n_2035),
.B(n_2036),
.Y(n_2085)
);

NOR2xp33_ASAP7_75t_L g2086 ( 
.A(n_1896),
.B(n_907),
.Y(n_2086)
);

NOR2xp33_ASAP7_75t_L g2087 ( 
.A(n_1906),
.B(n_913),
.Y(n_2087)
);

NOR2xp33_ASAP7_75t_SL g2088 ( 
.A(n_1751),
.B(n_1138),
.Y(n_2088)
);

OR2x2_ASAP7_75t_L g2089 ( 
.A(n_2000),
.B(n_1380),
.Y(n_2089)
);

INVxp67_ASAP7_75t_L g2090 ( 
.A(n_1952),
.Y(n_2090)
);

NAND2xp5_ASAP7_75t_L g2091 ( 
.A(n_2035),
.B(n_1124),
.Y(n_2091)
);

NAND2xp5_ASAP7_75t_L g2092 ( 
.A(n_2036),
.B(n_1163),
.Y(n_2092)
);

NAND2xp5_ASAP7_75t_SL g2093 ( 
.A(n_2043),
.B(n_1168),
.Y(n_2093)
);

NOR2xp33_ASAP7_75t_L g2094 ( 
.A(n_1906),
.B(n_913),
.Y(n_2094)
);

INVx2_ASAP7_75t_L g2095 ( 
.A(n_1873),
.Y(n_2095)
);

NAND2xp5_ASAP7_75t_L g2096 ( 
.A(n_2043),
.B(n_1170),
.Y(n_2096)
);

NAND2xp5_ASAP7_75t_SL g2097 ( 
.A(n_1871),
.B(n_1348),
.Y(n_2097)
);

INVx1_ASAP7_75t_L g2098 ( 
.A(n_1762),
.Y(n_2098)
);

INVx1_ASAP7_75t_L g2099 ( 
.A(n_1764),
.Y(n_2099)
);

CKINVDCx5p33_ASAP7_75t_R g2100 ( 
.A(n_1793),
.Y(n_2100)
);

INVx1_ASAP7_75t_L g2101 ( 
.A(n_1765),
.Y(n_2101)
);

INVx2_ASAP7_75t_L g2102 ( 
.A(n_2039),
.Y(n_2102)
);

NAND2xp5_ASAP7_75t_SL g2103 ( 
.A(n_1871),
.B(n_914),
.Y(n_2103)
);

NAND2xp5_ASAP7_75t_SL g2104 ( 
.A(n_1887),
.B(n_914),
.Y(n_2104)
);

NAND2xp5_ASAP7_75t_L g2105 ( 
.A(n_1887),
.B(n_916),
.Y(n_2105)
);

NAND2xp5_ASAP7_75t_L g2106 ( 
.A(n_1894),
.B(n_916),
.Y(n_2106)
);

NAND2xp5_ASAP7_75t_L g2107 ( 
.A(n_1894),
.B(n_1919),
.Y(n_2107)
);

INVx1_ASAP7_75t_L g2108 ( 
.A(n_1870),
.Y(n_2108)
);

NAND2xp5_ASAP7_75t_SL g2109 ( 
.A(n_1980),
.B(n_1371),
.Y(n_2109)
);

OR2x2_ASAP7_75t_L g2110 ( 
.A(n_2008),
.B(n_1378),
.Y(n_2110)
);

NAND2xp5_ASAP7_75t_SL g2111 ( 
.A(n_1980),
.B(n_1380),
.Y(n_2111)
);

INVx2_ASAP7_75t_L g2112 ( 
.A(n_2039),
.Y(n_2112)
);

INVx2_ASAP7_75t_L g2113 ( 
.A(n_1757),
.Y(n_2113)
);

INVx2_ASAP7_75t_L g2114 ( 
.A(n_1761),
.Y(n_2114)
);

NOR2xp33_ASAP7_75t_L g2115 ( 
.A(n_1778),
.B(n_1141),
.Y(n_2115)
);

INVx1_ASAP7_75t_L g2116 ( 
.A(n_1872),
.Y(n_2116)
);

NOR2xp33_ASAP7_75t_L g2117 ( 
.A(n_2034),
.B(n_1189),
.Y(n_2117)
);

AOI22xp5_ASAP7_75t_L g2118 ( 
.A1(n_1961),
.A2(n_866),
.B1(n_870),
.B2(n_865),
.Y(n_2118)
);

NAND2xp5_ASAP7_75t_L g2119 ( 
.A(n_1919),
.B(n_871),
.Y(n_2119)
);

CKINVDCx5p33_ASAP7_75t_R g2120 ( 
.A(n_2038),
.Y(n_2120)
);

AOI22xp5_ASAP7_75t_L g2121 ( 
.A1(n_1824),
.A2(n_1788),
.B1(n_1758),
.B2(n_1959),
.Y(n_2121)
);

AND2x2_ASAP7_75t_L g2122 ( 
.A(n_1843),
.B(n_1949),
.Y(n_2122)
);

INVx2_ASAP7_75t_L g2123 ( 
.A(n_2044),
.Y(n_2123)
);

AOI22xp5_ASAP7_75t_L g2124 ( 
.A1(n_1758),
.A2(n_878),
.B1(n_886),
.B2(n_875),
.Y(n_2124)
);

O2A1O1Ixp33_ASAP7_75t_L g2125 ( 
.A1(n_1844),
.A2(n_960),
.B(n_962),
.C(n_956),
.Y(n_2125)
);

NAND2xp5_ASAP7_75t_L g2126 ( 
.A(n_1758),
.B(n_889),
.Y(n_2126)
);

AOI21xp5_ASAP7_75t_L g2127 ( 
.A1(n_1862),
.A2(n_986),
.B(n_979),
.Y(n_2127)
);

NAND2xp5_ASAP7_75t_L g2128 ( 
.A(n_1758),
.B(n_891),
.Y(n_2128)
);

AOI22xp33_ASAP7_75t_L g2129 ( 
.A1(n_1879),
.A2(n_1256),
.B1(n_1359),
.B2(n_1252),
.Y(n_2129)
);

NAND2xp5_ASAP7_75t_L g2130 ( 
.A(n_1889),
.B(n_919),
.Y(n_2130)
);

NAND2xp5_ASAP7_75t_SL g2131 ( 
.A(n_1825),
.B(n_920),
.Y(n_2131)
);

NAND2xp5_ASAP7_75t_L g2132 ( 
.A(n_1876),
.B(n_1877),
.Y(n_2132)
);

INVx1_ASAP7_75t_L g2133 ( 
.A(n_1881),
.Y(n_2133)
);

NAND2xp5_ASAP7_75t_L g2134 ( 
.A(n_1818),
.B(n_925),
.Y(n_2134)
);

NAND2xp5_ASAP7_75t_L g2135 ( 
.A(n_1826),
.B(n_927),
.Y(n_2135)
);

INVx8_ASAP7_75t_L g2136 ( 
.A(n_1805),
.Y(n_2136)
);

AND2x6_ASAP7_75t_L g2137 ( 
.A(n_2030),
.B(n_1256),
.Y(n_2137)
);

INVx1_ASAP7_75t_L g2138 ( 
.A(n_1867),
.Y(n_2138)
);

INVx2_ASAP7_75t_SL g2139 ( 
.A(n_1866),
.Y(n_2139)
);

NAND2xp5_ASAP7_75t_SL g2140 ( 
.A(n_1825),
.B(n_929),
.Y(n_2140)
);

AOI22xp33_ASAP7_75t_L g2141 ( 
.A1(n_1879),
.A2(n_1359),
.B1(n_1213),
.B2(n_1226),
.Y(n_2141)
);

INVx1_ASAP7_75t_L g2142 ( 
.A(n_1868),
.Y(n_2142)
);

AND2x2_ASAP7_75t_L g2143 ( 
.A(n_1949),
.B(n_1189),
.Y(n_2143)
);

NOR2xp33_ASAP7_75t_L g2144 ( 
.A(n_1895),
.B(n_1213),
.Y(n_2144)
);

INVxp67_ASAP7_75t_L g2145 ( 
.A(n_1952),
.Y(n_2145)
);

NAND2xp5_ASAP7_75t_L g2146 ( 
.A(n_1830),
.B(n_931),
.Y(n_2146)
);

NAND2xp5_ASAP7_75t_L g2147 ( 
.A(n_1831),
.B(n_932),
.Y(n_2147)
);

INVx2_ASAP7_75t_SL g2148 ( 
.A(n_1866),
.Y(n_2148)
);

NOR3xp33_ASAP7_75t_L g2149 ( 
.A(n_1915),
.B(n_1005),
.C(n_992),
.Y(n_2149)
);

NOR3xp33_ASAP7_75t_L g2150 ( 
.A(n_1915),
.B(n_1844),
.C(n_2008),
.Y(n_2150)
);

NAND2xp5_ASAP7_75t_SL g2151 ( 
.A(n_1863),
.B(n_934),
.Y(n_2151)
);

NOR2xp33_ASAP7_75t_L g2152 ( 
.A(n_1811),
.B(n_1226),
.Y(n_2152)
);

OR2x2_ASAP7_75t_L g2153 ( 
.A(n_1999),
.B(n_1060),
.Y(n_2153)
);

INVx2_ASAP7_75t_L g2154 ( 
.A(n_2044),
.Y(n_2154)
);

NAND2xp33_ASAP7_75t_L g2155 ( 
.A(n_1890),
.B(n_2033),
.Y(n_2155)
);

INVx2_ASAP7_75t_L g2156 ( 
.A(n_2040),
.Y(n_2156)
);

INVx1_ASAP7_75t_L g2157 ( 
.A(n_1869),
.Y(n_2157)
);

INVx1_ASAP7_75t_L g2158 ( 
.A(n_1874),
.Y(n_2158)
);

NOR3xp33_ASAP7_75t_L g2159 ( 
.A(n_2013),
.B(n_1125),
.C(n_1090),
.Y(n_2159)
);

NAND2xp5_ASAP7_75t_L g2160 ( 
.A(n_1834),
.B(n_937),
.Y(n_2160)
);

INVx1_ASAP7_75t_L g2161 ( 
.A(n_1875),
.Y(n_2161)
);

NAND2xp5_ASAP7_75t_L g2162 ( 
.A(n_1841),
.B(n_939),
.Y(n_2162)
);

INVx2_ASAP7_75t_L g2163 ( 
.A(n_2046),
.Y(n_2163)
);

AOI22xp5_ASAP7_75t_L g2164 ( 
.A1(n_1959),
.A2(n_942),
.B1(n_952),
.B2(n_940),
.Y(n_2164)
);

INVx2_ASAP7_75t_SL g2165 ( 
.A(n_1952),
.Y(n_2165)
);

INVx2_ASAP7_75t_SL g2166 ( 
.A(n_1803),
.Y(n_2166)
);

NAND2xp5_ASAP7_75t_L g2167 ( 
.A(n_1847),
.B(n_955),
.Y(n_2167)
);

INVx1_ASAP7_75t_L g2168 ( 
.A(n_1883),
.Y(n_2168)
);

AOI22xp5_ASAP7_75t_L g2169 ( 
.A1(n_1853),
.A2(n_964),
.B1(n_966),
.B2(n_963),
.Y(n_2169)
);

NAND2xp5_ASAP7_75t_SL g2170 ( 
.A(n_1863),
.B(n_968),
.Y(n_2170)
);

AOI22xp33_ASAP7_75t_L g2171 ( 
.A1(n_2033),
.A2(n_1359),
.B1(n_1250),
.B2(n_1257),
.Y(n_2171)
);

INVx2_ASAP7_75t_L g2172 ( 
.A(n_1884),
.Y(n_2172)
);

AOI22xp5_ASAP7_75t_L g2173 ( 
.A1(n_1926),
.A2(n_983),
.B1(n_985),
.B2(n_972),
.Y(n_2173)
);

AND2x2_ASAP7_75t_SL g2174 ( 
.A(n_1836),
.B(n_1238),
.Y(n_2174)
);

INVx2_ASAP7_75t_SL g2175 ( 
.A(n_1803),
.Y(n_2175)
);

OR2x2_ASAP7_75t_L g2176 ( 
.A(n_1882),
.B(n_1174),
.Y(n_2176)
);

NAND2xp5_ASAP7_75t_L g2177 ( 
.A(n_1892),
.B(n_988),
.Y(n_2177)
);

INVx1_ASAP7_75t_L g2178 ( 
.A(n_1897),
.Y(n_2178)
);

INVx1_ASAP7_75t_L g2179 ( 
.A(n_1898),
.Y(n_2179)
);

INVx1_ASAP7_75t_L g2180 ( 
.A(n_1902),
.Y(n_2180)
);

AND2x2_ASAP7_75t_L g2181 ( 
.A(n_1900),
.B(n_1238),
.Y(n_2181)
);

NOR2xp33_ASAP7_75t_L g2182 ( 
.A(n_1974),
.B(n_1250),
.Y(n_2182)
);

INVx1_ASAP7_75t_L g2183 ( 
.A(n_1905),
.Y(n_2183)
);

INVx1_ASAP7_75t_L g2184 ( 
.A(n_1907),
.Y(n_2184)
);

INVx1_ASAP7_75t_L g2185 ( 
.A(n_1908),
.Y(n_2185)
);

NAND2xp5_ASAP7_75t_SL g2186 ( 
.A(n_1863),
.B(n_989),
.Y(n_2186)
);

AND2x4_ASAP7_75t_L g2187 ( 
.A(n_1776),
.B(n_990),
.Y(n_2187)
);

INVx2_ASAP7_75t_L g2188 ( 
.A(n_1752),
.Y(n_2188)
);

NAND2xp5_ASAP7_75t_SL g2189 ( 
.A(n_1850),
.B(n_996),
.Y(n_2189)
);

NOR2xp33_ASAP7_75t_L g2190 ( 
.A(n_1786),
.B(n_1257),
.Y(n_2190)
);

NAND2xp33_ASAP7_75t_L g2191 ( 
.A(n_1890),
.B(n_1008),
.Y(n_2191)
);

NAND2xp5_ASAP7_75t_L g2192 ( 
.A(n_1899),
.B(n_1010),
.Y(n_2192)
);

NAND2xp5_ASAP7_75t_SL g2193 ( 
.A(n_1850),
.B(n_1012),
.Y(n_2193)
);

NAND2xp5_ASAP7_75t_SL g2194 ( 
.A(n_1934),
.B(n_1013),
.Y(n_2194)
);

NAND2xp5_ASAP7_75t_SL g2195 ( 
.A(n_1953),
.B(n_1019),
.Y(n_2195)
);

NOR3xp33_ASAP7_75t_L g2196 ( 
.A(n_2019),
.B(n_1320),
.C(n_1181),
.Y(n_2196)
);

INVx2_ASAP7_75t_L g2197 ( 
.A(n_1754),
.Y(n_2197)
);

NAND2xp33_ASAP7_75t_L g2198 ( 
.A(n_1890),
.B(n_1020),
.Y(n_2198)
);

NAND2xp5_ASAP7_75t_L g2199 ( 
.A(n_1901),
.B(n_1021),
.Y(n_2199)
);

AOI22xp5_ASAP7_75t_L g2200 ( 
.A1(n_1926),
.A2(n_1023),
.B1(n_1036),
.B2(n_1031),
.Y(n_2200)
);

INVx1_ASAP7_75t_L g2201 ( 
.A(n_1903),
.Y(n_2201)
);

NOR2xp33_ASAP7_75t_L g2202 ( 
.A(n_1917),
.B(n_1352),
.Y(n_2202)
);

INVx2_ASAP7_75t_SL g2203 ( 
.A(n_1803),
.Y(n_2203)
);

OR2x2_ASAP7_75t_L g2204 ( 
.A(n_1954),
.B(n_1038),
.Y(n_2204)
);

INVx2_ASAP7_75t_L g2205 ( 
.A(n_2032),
.Y(n_2205)
);

AOI22xp33_ASAP7_75t_L g2206 ( 
.A1(n_2033),
.A2(n_1359),
.B1(n_997),
.B2(n_1035),
.Y(n_2206)
);

NAND2xp5_ASAP7_75t_L g2207 ( 
.A(n_1909),
.B(n_1044),
.Y(n_2207)
);

NAND2xp5_ASAP7_75t_SL g2208 ( 
.A(n_1953),
.B(n_1046),
.Y(n_2208)
);

NAND2xp5_ASAP7_75t_L g2209 ( 
.A(n_1931),
.B(n_1048),
.Y(n_2209)
);

NAND2xp5_ASAP7_75t_L g2210 ( 
.A(n_1931),
.B(n_1050),
.Y(n_2210)
);

AOI22xp5_ASAP7_75t_L g2211 ( 
.A1(n_1939),
.A2(n_1056),
.B1(n_1063),
.B2(n_1055),
.Y(n_2211)
);

NAND2xp5_ASAP7_75t_L g2212 ( 
.A(n_1932),
.B(n_1066),
.Y(n_2212)
);

INVx1_ASAP7_75t_L g2213 ( 
.A(n_1916),
.Y(n_2213)
);

AOI22xp5_ASAP7_75t_L g2214 ( 
.A1(n_1939),
.A2(n_1073),
.B1(n_1077),
.B2(n_1068),
.Y(n_2214)
);

AND2x2_ASAP7_75t_L g2215 ( 
.A(n_1904),
.B(n_994),
.Y(n_2215)
);

INVxp67_ASAP7_75t_L g2216 ( 
.A(n_1996),
.Y(n_2216)
);

INVx1_ASAP7_75t_L g2217 ( 
.A(n_1918),
.Y(n_2217)
);

INVx2_ASAP7_75t_L g2218 ( 
.A(n_2037),
.Y(n_2218)
);

INVx1_ASAP7_75t_L g2219 ( 
.A(n_1922),
.Y(n_2219)
);

NOR2xp33_ASAP7_75t_L g2220 ( 
.A(n_1917),
.B(n_1079),
.Y(n_2220)
);

NAND2xp5_ASAP7_75t_L g2221 ( 
.A(n_1932),
.B(n_1082),
.Y(n_2221)
);

BUFx6f_ASAP7_75t_L g2222 ( 
.A(n_1755),
.Y(n_2222)
);

NOR2xp33_ASAP7_75t_L g2223 ( 
.A(n_1766),
.B(n_1083),
.Y(n_2223)
);

INVx1_ASAP7_75t_L g2224 ( 
.A(n_1928),
.Y(n_2224)
);

NAND2xp5_ASAP7_75t_L g2225 ( 
.A(n_1865),
.B(n_1085),
.Y(n_2225)
);

NAND2xp5_ASAP7_75t_L g2226 ( 
.A(n_1865),
.B(n_1089),
.Y(n_2226)
);

AND2x2_ASAP7_75t_L g2227 ( 
.A(n_1829),
.B(n_994),
.Y(n_2227)
);

INVx1_ASAP7_75t_L g2228 ( 
.A(n_1930),
.Y(n_2228)
);

INVx2_ASAP7_75t_L g2229 ( 
.A(n_2045),
.Y(n_2229)
);

BUFx5_ASAP7_75t_L g2230 ( 
.A(n_2033),
.Y(n_2230)
);

BUFx12f_ASAP7_75t_SL g2231 ( 
.A(n_1836),
.Y(n_2231)
);

NOR2x1p5_ASAP7_75t_L g2232 ( 
.A(n_2047),
.B(n_1099),
.Y(n_2232)
);

AOI22xp5_ASAP7_75t_L g2233 ( 
.A1(n_1973),
.A2(n_1093),
.B1(n_1094),
.B2(n_1092),
.Y(n_2233)
);

INVx2_ASAP7_75t_L g2234 ( 
.A(n_1756),
.Y(n_2234)
);

INVxp67_ASAP7_75t_L g2235 ( 
.A(n_1996),
.Y(n_2235)
);

NAND2xp5_ASAP7_75t_SL g2236 ( 
.A(n_1951),
.B(n_1095),
.Y(n_2236)
);

INVx2_ASAP7_75t_L g2237 ( 
.A(n_1808),
.Y(n_2237)
);

BUFx6f_ASAP7_75t_L g2238 ( 
.A(n_1911),
.Y(n_2238)
);

INVx2_ASAP7_75t_L g2239 ( 
.A(n_1809),
.Y(n_2239)
);

NAND2xp5_ASAP7_75t_L g2240 ( 
.A(n_1885),
.B(n_1101),
.Y(n_2240)
);

NAND2xp5_ASAP7_75t_L g2241 ( 
.A(n_1885),
.B(n_1108),
.Y(n_2241)
);

AND2x2_ASAP7_75t_SL g2242 ( 
.A(n_1807),
.B(n_1018),
.Y(n_2242)
);

NAND2xp5_ASAP7_75t_L g2243 ( 
.A(n_1781),
.B(n_1109),
.Y(n_2243)
);

AND2x2_ASAP7_75t_SL g2244 ( 
.A(n_1965),
.B(n_1022),
.Y(n_2244)
);

BUFx8_ASAP7_75t_L g2245 ( 
.A(n_1969),
.Y(n_2245)
);

NAND2xp5_ASAP7_75t_L g2246 ( 
.A(n_1787),
.B(n_1111),
.Y(n_2246)
);

INVxp67_ASAP7_75t_L g2247 ( 
.A(n_1972),
.Y(n_2247)
);

NAND2xp5_ASAP7_75t_SL g2248 ( 
.A(n_1951),
.B(n_1112),
.Y(n_2248)
);

NAND2xp5_ASAP7_75t_SL g2249 ( 
.A(n_1837),
.B(n_1118),
.Y(n_2249)
);

INVx2_ASAP7_75t_L g2250 ( 
.A(n_1812),
.Y(n_2250)
);

BUFx6f_ASAP7_75t_L g2251 ( 
.A(n_1911),
.Y(n_2251)
);

NAND2xp5_ASAP7_75t_L g2252 ( 
.A(n_1790),
.B(n_1120),
.Y(n_2252)
);

INVx2_ASAP7_75t_SL g2253 ( 
.A(n_1982),
.Y(n_2253)
);

NOR2xp33_ASAP7_75t_L g2254 ( 
.A(n_1935),
.B(n_1135),
.Y(n_2254)
);

INVx1_ASAP7_75t_L g2255 ( 
.A(n_1933),
.Y(n_2255)
);

INVx2_ASAP7_75t_L g2256 ( 
.A(n_1813),
.Y(n_2256)
);

INVx1_ASAP7_75t_L g2257 ( 
.A(n_1910),
.Y(n_2257)
);

NOR2xp33_ASAP7_75t_L g2258 ( 
.A(n_1950),
.B(n_1136),
.Y(n_2258)
);

HB1xp67_ASAP7_75t_L g2259 ( 
.A(n_1976),
.Y(n_2259)
);

BUFx2_ASAP7_75t_L g2260 ( 
.A(n_1829),
.Y(n_2260)
);

NOR3xp33_ASAP7_75t_L g2261 ( 
.A(n_1965),
.B(n_1795),
.C(n_1819),
.Y(n_2261)
);

NOR3xp33_ASAP7_75t_L g2262 ( 
.A(n_1979),
.B(n_1143),
.C(n_1139),
.Y(n_2262)
);

NOR2xp33_ASAP7_75t_L g2263 ( 
.A(n_1937),
.B(n_1938),
.Y(n_2263)
);

NAND2xp5_ASAP7_75t_L g2264 ( 
.A(n_1791),
.B(n_1144),
.Y(n_2264)
);

INVx2_ASAP7_75t_L g2265 ( 
.A(n_1815),
.Y(n_2265)
);

NAND2xp5_ASAP7_75t_L g2266 ( 
.A(n_1817),
.B(n_2031),
.Y(n_2266)
);

NAND2xp5_ASAP7_75t_L g2267 ( 
.A(n_1817),
.B(n_1146),
.Y(n_2267)
);

INVx2_ASAP7_75t_L g2268 ( 
.A(n_1816),
.Y(n_2268)
);

NAND2xp5_ASAP7_75t_L g2269 ( 
.A(n_1817),
.B(n_1147),
.Y(n_2269)
);

INVxp67_ASAP7_75t_L g2270 ( 
.A(n_1829),
.Y(n_2270)
);

NAND2xp5_ASAP7_75t_L g2271 ( 
.A(n_1817),
.B(n_1149),
.Y(n_2271)
);

NOR2xp33_ASAP7_75t_L g2272 ( 
.A(n_1940),
.B(n_1157),
.Y(n_2272)
);

NOR2xp33_ASAP7_75t_L g2273 ( 
.A(n_1942),
.B(n_1159),
.Y(n_2273)
);

BUFx3_ASAP7_75t_L g2274 ( 
.A(n_1797),
.Y(n_2274)
);

INVx1_ASAP7_75t_L g2275 ( 
.A(n_1910),
.Y(n_2275)
);

NAND2xp5_ASAP7_75t_L g2276 ( 
.A(n_1833),
.B(n_1150),
.Y(n_2276)
);

AOI22xp5_ASAP7_75t_L g2277 ( 
.A1(n_1973),
.A2(n_1958),
.B1(n_1955),
.B2(n_1945),
.Y(n_2277)
);

BUFx6f_ASAP7_75t_L g2278 ( 
.A(n_1911),
.Y(n_2278)
);

NAND2xp5_ASAP7_75t_L g2279 ( 
.A(n_1833),
.B(n_1162),
.Y(n_2279)
);

HB1xp67_ASAP7_75t_L g2280 ( 
.A(n_2005),
.Y(n_2280)
);

NAND2xp5_ASAP7_75t_L g2281 ( 
.A(n_2031),
.B(n_1164),
.Y(n_2281)
);

OAI22xp5_ASAP7_75t_L g2282 ( 
.A1(n_1779),
.A2(n_1039),
.B1(n_1057),
.B2(n_1014),
.Y(n_2282)
);

NOR2xp33_ASAP7_75t_L g2283 ( 
.A(n_1913),
.B(n_1165),
.Y(n_2283)
);

AOI22xp33_ASAP7_75t_L g2284 ( 
.A1(n_1913),
.A2(n_1958),
.B1(n_1890),
.B2(n_1923),
.Y(n_2284)
);

NAND2xp5_ASAP7_75t_L g2285 ( 
.A(n_1878),
.B(n_1880),
.Y(n_2285)
);

INVx1_ASAP7_75t_L g2286 ( 
.A(n_1858),
.Y(n_2286)
);

AOI22xp33_ASAP7_75t_L g2287 ( 
.A1(n_1923),
.A2(n_1956),
.B1(n_1924),
.B2(n_1792),
.Y(n_2287)
);

INVx2_ASAP7_75t_L g2288 ( 
.A(n_1822),
.Y(n_2288)
);

A2O1A1Ixp33_ASAP7_75t_L g2289 ( 
.A1(n_1855),
.A2(n_1070),
.B(n_1076),
.C(n_1062),
.Y(n_2289)
);

AND2x2_ASAP7_75t_L g2290 ( 
.A(n_1991),
.B(n_994),
.Y(n_2290)
);

AOI22xp33_ASAP7_75t_L g2291 ( 
.A1(n_1956),
.A2(n_1103),
.B1(n_1110),
.B2(n_1091),
.Y(n_2291)
);

NAND2xp5_ASAP7_75t_SL g2292 ( 
.A(n_1861),
.B(n_1169),
.Y(n_2292)
);

INVx1_ASAP7_75t_L g2293 ( 
.A(n_1858),
.Y(n_2293)
);

AND2x2_ASAP7_75t_L g2294 ( 
.A(n_1772),
.B(n_1024),
.Y(n_2294)
);

NAND2xp5_ASAP7_75t_SL g2295 ( 
.A(n_1779),
.B(n_1171),
.Y(n_2295)
);

NAND2xp5_ASAP7_75t_SL g2296 ( 
.A(n_1792),
.B(n_1173),
.Y(n_2296)
);

NAND2xp5_ASAP7_75t_L g2297 ( 
.A(n_1924),
.B(n_1184),
.Y(n_2297)
);

INVxp67_ASAP7_75t_L g2298 ( 
.A(n_1948),
.Y(n_2298)
);

INVx1_ASAP7_75t_L g2299 ( 
.A(n_1855),
.Y(n_2299)
);

INVx2_ASAP7_75t_L g2300 ( 
.A(n_1827),
.Y(n_2300)
);

INVx3_ASAP7_75t_L g2301 ( 
.A(n_1794),
.Y(n_2301)
);

NAND2xp5_ASAP7_75t_L g2302 ( 
.A(n_1835),
.B(n_1190),
.Y(n_2302)
);

INVx1_ASAP7_75t_L g2303 ( 
.A(n_1750),
.Y(n_2303)
);

NAND2xp5_ASAP7_75t_L g2304 ( 
.A(n_1821),
.B(n_1851),
.Y(n_2304)
);

INVx1_ASAP7_75t_L g2305 ( 
.A(n_1750),
.Y(n_2305)
);

NAND2xp5_ASAP7_75t_L g2306 ( 
.A(n_1794),
.B(n_1191),
.Y(n_2306)
);

NAND2xp5_ASAP7_75t_L g2307 ( 
.A(n_1828),
.B(n_1196),
.Y(n_2307)
);

INVx1_ASAP7_75t_L g2308 ( 
.A(n_1763),
.Y(n_2308)
);

NAND2xp5_ASAP7_75t_L g2309 ( 
.A(n_1828),
.B(n_1199),
.Y(n_2309)
);

NAND2xp5_ASAP7_75t_SL g2310 ( 
.A(n_1810),
.B(n_1201),
.Y(n_2310)
);

NAND2xp5_ASAP7_75t_SL g2311 ( 
.A(n_1810),
.B(n_1202),
.Y(n_2311)
);

INVx2_ASAP7_75t_L g2312 ( 
.A(n_1888),
.Y(n_2312)
);

NOR2xp33_ASAP7_75t_L g2313 ( 
.A(n_1997),
.B(n_1204),
.Y(n_2313)
);

NOR2xp33_ASAP7_75t_L g2314 ( 
.A(n_1985),
.B(n_1205),
.Y(n_2314)
);

AND2x6_ASAP7_75t_SL g2315 ( 
.A(n_2015),
.B(n_1342),
.Y(n_2315)
);

NAND2xp5_ASAP7_75t_L g2316 ( 
.A(n_1832),
.B(n_1206),
.Y(n_2316)
);

INVx1_ASAP7_75t_L g2317 ( 
.A(n_1763),
.Y(n_2317)
);

NAND2xp5_ASAP7_75t_SL g2318 ( 
.A(n_2010),
.B(n_1207),
.Y(n_2318)
);

INVx1_ASAP7_75t_L g2319 ( 
.A(n_1767),
.Y(n_2319)
);

INVx1_ASAP7_75t_L g2320 ( 
.A(n_1769),
.Y(n_2320)
);

NOR3xp33_ASAP7_75t_L g2321 ( 
.A(n_1989),
.B(n_1943),
.C(n_2015),
.Y(n_2321)
);

NAND2xp5_ASAP7_75t_SL g2322 ( 
.A(n_2010),
.B(n_1209),
.Y(n_2322)
);

NAND2xp5_ASAP7_75t_L g2323 ( 
.A(n_1832),
.B(n_1218),
.Y(n_2323)
);

BUFx3_ASAP7_75t_L g2324 ( 
.A(n_1753),
.Y(n_2324)
);

OAI221xp5_ASAP7_75t_L g2325 ( 
.A1(n_1772),
.A2(n_1233),
.B1(n_1234),
.B2(n_1232),
.C(n_1224),
.Y(n_2325)
);

INVx2_ASAP7_75t_SL g2326 ( 
.A(n_1759),
.Y(n_2326)
);

INVx1_ASAP7_75t_L g2327 ( 
.A(n_1770),
.Y(n_2327)
);

NAND2xp33_ASAP7_75t_L g2328 ( 
.A(n_1956),
.B(n_1235),
.Y(n_2328)
);

BUFx3_ASAP7_75t_L g2329 ( 
.A(n_1759),
.Y(n_2329)
);

OR2x6_ASAP7_75t_L g2330 ( 
.A(n_1886),
.B(n_1022),
.Y(n_2330)
);

AOI221xp5_ASAP7_75t_L g2331 ( 
.A1(n_1969),
.A2(n_1799),
.B1(n_1116),
.B2(n_1121),
.C(n_1115),
.Y(n_2331)
);

AND2x2_ASAP7_75t_L g2332 ( 
.A(n_1796),
.B(n_1024),
.Y(n_2332)
);

AND2x6_ASAP7_75t_L g2333 ( 
.A(n_1798),
.B(n_1030),
.Y(n_2333)
);

NAND3xp33_ASAP7_75t_L g2334 ( 
.A(n_2001),
.B(n_2020),
.C(n_2011),
.Y(n_2334)
);

NAND2xp5_ASAP7_75t_L g2335 ( 
.A(n_1838),
.B(n_1236),
.Y(n_2335)
);

CKINVDCx5p33_ASAP7_75t_R g2336 ( 
.A(n_1796),
.Y(n_2336)
);

NAND2xp5_ASAP7_75t_L g2337 ( 
.A(n_1839),
.B(n_1239),
.Y(n_2337)
);

INVx2_ASAP7_75t_L g2338 ( 
.A(n_1771),
.Y(n_2338)
);

INVx3_ASAP7_75t_L g2339 ( 
.A(n_2023),
.Y(n_2339)
);

OR2x2_ASAP7_75t_L g2340 ( 
.A(n_2003),
.B(n_1240),
.Y(n_2340)
);

NAND2xp5_ASAP7_75t_L g2341 ( 
.A(n_1782),
.B(n_1241),
.Y(n_2341)
);

NOR2xp33_ASAP7_75t_L g2342 ( 
.A(n_1840),
.B(n_1842),
.Y(n_2342)
);

NOR2xp33_ASAP7_75t_L g2343 ( 
.A(n_1845),
.B(n_1247),
.Y(n_2343)
);

AND2x2_ASAP7_75t_L g2344 ( 
.A(n_2041),
.B(n_1024),
.Y(n_2344)
);

INVx1_ASAP7_75t_L g2345 ( 
.A(n_1773),
.Y(n_2345)
);

BUFx6f_ASAP7_75t_L g2346 ( 
.A(n_1920),
.Y(n_2346)
);

NAND2xp5_ASAP7_75t_SL g2347 ( 
.A(n_2028),
.B(n_1248),
.Y(n_2347)
);

NAND2xp33_ASAP7_75t_L g2348 ( 
.A(n_1956),
.B(n_1253),
.Y(n_2348)
);

INVx1_ASAP7_75t_L g2349 ( 
.A(n_1775),
.Y(n_2349)
);

NAND2xp5_ASAP7_75t_SL g2350 ( 
.A(n_2028),
.B(n_1258),
.Y(n_2350)
);

NAND2xp5_ASAP7_75t_L g2351 ( 
.A(n_1846),
.B(n_1266),
.Y(n_2351)
);

NAND2xp5_ASAP7_75t_L g2352 ( 
.A(n_1848),
.B(n_1267),
.Y(n_2352)
);

AOI22xp5_ASAP7_75t_L g2353 ( 
.A1(n_1856),
.A2(n_1272),
.B1(n_1275),
.B2(n_1268),
.Y(n_2353)
);

AOI22xp33_ASAP7_75t_L g2354 ( 
.A1(n_1912),
.A2(n_1122),
.B1(n_1132),
.B2(n_1113),
.Y(n_2354)
);

INVx2_ASAP7_75t_L g2355 ( 
.A(n_1777),
.Y(n_2355)
);

INVx2_ASAP7_75t_L g2356 ( 
.A(n_1780),
.Y(n_2356)
);

NAND2xp5_ASAP7_75t_SL g2357 ( 
.A(n_1993),
.B(n_1277),
.Y(n_2357)
);

NAND3xp33_ASAP7_75t_L g2358 ( 
.A(n_2001),
.B(n_930),
.C(n_904),
.Y(n_2358)
);

NOR2xp33_ASAP7_75t_L g2359 ( 
.A(n_1849),
.B(n_1278),
.Y(n_2359)
);

A2O1A1Ixp33_ASAP7_75t_L g2360 ( 
.A1(n_2011),
.A2(n_1137),
.B(n_1152),
.C(n_1134),
.Y(n_2360)
);

OAI22xp5_ASAP7_75t_L g2361 ( 
.A1(n_1993),
.A2(n_1175),
.B1(n_1180),
.B2(n_1167),
.Y(n_2361)
);

NAND2xp5_ASAP7_75t_SL g2362 ( 
.A(n_1994),
.B(n_1281),
.Y(n_2362)
);

NAND2xp5_ASAP7_75t_L g2363 ( 
.A(n_1852),
.B(n_1282),
.Y(n_2363)
);

INVx2_ASAP7_75t_L g2364 ( 
.A(n_1783),
.Y(n_2364)
);

INVx2_ASAP7_75t_L g2365 ( 
.A(n_1784),
.Y(n_2365)
);

NAND2xp5_ASAP7_75t_SL g2366 ( 
.A(n_1994),
.B(n_1283),
.Y(n_2366)
);

NAND2xp5_ASAP7_75t_L g2367 ( 
.A(n_1857),
.B(n_1286),
.Y(n_2367)
);

NAND2xp5_ASAP7_75t_SL g2368 ( 
.A(n_2012),
.B(n_1287),
.Y(n_2368)
);

A2O1A1Ixp33_ASAP7_75t_L g2369 ( 
.A1(n_2020),
.A2(n_1192),
.B(n_1203),
.C(n_1183),
.Y(n_2369)
);

INVx2_ASAP7_75t_L g2370 ( 
.A(n_1789),
.Y(n_2370)
);

NAND2xp5_ASAP7_75t_L g2371 ( 
.A(n_1860),
.B(n_1288),
.Y(n_2371)
);

NAND3xp33_ASAP7_75t_L g2372 ( 
.A(n_1936),
.B(n_1975),
.C(n_2026),
.Y(n_2372)
);

NAND2xp5_ASAP7_75t_SL g2373 ( 
.A(n_2012),
.B(n_1290),
.Y(n_2373)
);

INVx2_ASAP7_75t_L g2374 ( 
.A(n_1914),
.Y(n_2374)
);

NAND2xp5_ASAP7_75t_SL g2375 ( 
.A(n_2018),
.B(n_1296),
.Y(n_2375)
);

NOR2xp67_ASAP7_75t_L g2376 ( 
.A(n_2018),
.B(n_0),
.Y(n_2376)
);

INVx2_ASAP7_75t_SL g2377 ( 
.A(n_2041),
.Y(n_2377)
);

AND2x2_ASAP7_75t_L g2378 ( 
.A(n_1800),
.B(n_1059),
.Y(n_2378)
);

INVx1_ASAP7_75t_L g2379 ( 
.A(n_1801),
.Y(n_2379)
);

AOI22xp5_ASAP7_75t_L g2380 ( 
.A1(n_1802),
.A2(n_1304),
.B1(n_1306),
.B2(n_1297),
.Y(n_2380)
);

NAND2xp5_ASAP7_75t_L g2381 ( 
.A(n_1925),
.B(n_1307),
.Y(n_2381)
);

NAND2xp5_ASAP7_75t_L g2382 ( 
.A(n_1927),
.B(n_1312),
.Y(n_2382)
);

NOR2xp33_ASAP7_75t_L g2383 ( 
.A(n_2004),
.B(n_1328),
.Y(n_2383)
);

NAND2xp5_ASAP7_75t_SL g2384 ( 
.A(n_2009),
.B(n_1329),
.Y(n_2384)
);

NAND2xp5_ASAP7_75t_SL g2385 ( 
.A(n_2009),
.B(n_1335),
.Y(n_2385)
);

NAND2xp5_ASAP7_75t_SL g2386 ( 
.A(n_1941),
.B(n_1336),
.Y(n_2386)
);

NAND2xp5_ASAP7_75t_L g2387 ( 
.A(n_1921),
.B(n_1344),
.Y(n_2387)
);

CKINVDCx5p33_ASAP7_75t_R g2388 ( 
.A(n_2023),
.Y(n_2388)
);

INVx1_ASAP7_75t_L g2389 ( 
.A(n_1823),
.Y(n_2389)
);

NAND2xp5_ASAP7_75t_SL g2390 ( 
.A(n_1944),
.B(n_1351),
.Y(n_2390)
);

NAND2xp5_ASAP7_75t_L g2391 ( 
.A(n_1823),
.B(n_1354),
.Y(n_2391)
);

AOI22xp33_ASAP7_75t_L g2392 ( 
.A1(n_1921),
.A2(n_1212),
.B1(n_1223),
.B2(n_1208),
.Y(n_2392)
);

NAND2xp5_ASAP7_75t_L g2393 ( 
.A(n_1946),
.B(n_1357),
.Y(n_2393)
);

INVx2_ASAP7_75t_L g2394 ( 
.A(n_1970),
.Y(n_2394)
);

INVx1_ASAP7_75t_L g2395 ( 
.A(n_1891),
.Y(n_2395)
);

INVx1_ASAP7_75t_L g2396 ( 
.A(n_1970),
.Y(n_2396)
);

INVx2_ASAP7_75t_SL g2397 ( 
.A(n_2136),
.Y(n_2397)
);

INVx1_ASAP7_75t_L g2398 ( 
.A(n_2178),
.Y(n_2398)
);

NAND2xp5_ASAP7_75t_L g2399 ( 
.A(n_2053),
.B(n_1358),
.Y(n_2399)
);

NAND2xp5_ASAP7_75t_SL g2400 ( 
.A(n_2088),
.B(n_1363),
.Y(n_2400)
);

INVx4_ASAP7_75t_L g2401 ( 
.A(n_2136),
.Y(n_2401)
);

AND2x4_ASAP7_75t_L g2402 ( 
.A(n_2060),
.B(n_2068),
.Y(n_2402)
);

AND2x4_ASAP7_75t_L g2403 ( 
.A(n_2329),
.B(n_1227),
.Y(n_2403)
);

INVx2_ASAP7_75t_L g2404 ( 
.A(n_2172),
.Y(n_2404)
);

NAND2xp5_ASAP7_75t_SL g2405 ( 
.A(n_2088),
.B(n_1365),
.Y(n_2405)
);

BUFx6f_ASAP7_75t_L g2406 ( 
.A(n_2238),
.Y(n_2406)
);

INVx1_ASAP7_75t_L g2407 ( 
.A(n_2179),
.Y(n_2407)
);

INVx2_ASAP7_75t_SL g2408 ( 
.A(n_2136),
.Y(n_2408)
);

AOI22xp33_ASAP7_75t_L g2409 ( 
.A1(n_2150),
.A2(n_1067),
.B1(n_1340),
.B2(n_1059),
.Y(n_2409)
);

NAND2xp5_ASAP7_75t_L g2410 ( 
.A(n_2057),
.B(n_1366),
.Y(n_2410)
);

AOI22xp33_ASAP7_75t_L g2411 ( 
.A1(n_2122),
.A2(n_1067),
.B1(n_1340),
.B2(n_1059),
.Y(n_2411)
);

BUFx2_ASAP7_75t_SL g2412 ( 
.A(n_2082),
.Y(n_2412)
);

BUFx2_ASAP7_75t_L g2413 ( 
.A(n_2063),
.Y(n_2413)
);

NAND2xp5_ASAP7_75t_L g2414 ( 
.A(n_2057),
.B(n_1228),
.Y(n_2414)
);

INVx1_ASAP7_75t_SL g2415 ( 
.A(n_2072),
.Y(n_2415)
);

NAND2xp5_ASAP7_75t_L g2416 ( 
.A(n_2065),
.B(n_1245),
.Y(n_2416)
);

INVx2_ASAP7_75t_L g2417 ( 
.A(n_2156),
.Y(n_2417)
);

INVx2_ASAP7_75t_SL g2418 ( 
.A(n_2245),
.Y(n_2418)
);

AND2x4_ASAP7_75t_L g2419 ( 
.A(n_2165),
.B(n_1246),
.Y(n_2419)
);

INVx2_ASAP7_75t_L g2420 ( 
.A(n_2163),
.Y(n_2420)
);

INVx1_ASAP7_75t_L g2421 ( 
.A(n_2180),
.Y(n_2421)
);

INVx1_ASAP7_75t_L g2422 ( 
.A(n_2183),
.Y(n_2422)
);

NAND2xp5_ASAP7_75t_SL g2423 ( 
.A(n_2174),
.B(n_1067),
.Y(n_2423)
);

NOR2xp33_ASAP7_75t_L g2424 ( 
.A(n_2182),
.B(n_1340),
.Y(n_2424)
);

AOI22xp5_ASAP7_75t_L g2425 ( 
.A1(n_2107),
.A2(n_1251),
.B1(n_1263),
.B2(n_1249),
.Y(n_2425)
);

AND2x6_ASAP7_75t_SL g2426 ( 
.A(n_2330),
.B(n_1265),
.Y(n_2426)
);

AND2x2_ASAP7_75t_SL g2427 ( 
.A(n_2244),
.B(n_904),
.Y(n_2427)
);

INVx2_ASAP7_75t_L g2428 ( 
.A(n_2099),
.Y(n_2428)
);

INVx1_ASAP7_75t_L g2429 ( 
.A(n_2184),
.Y(n_2429)
);

INVx2_ASAP7_75t_L g2430 ( 
.A(n_2101),
.Y(n_2430)
);

INVx1_ASAP7_75t_L g2431 ( 
.A(n_2185),
.Y(n_2431)
);

NAND2xp5_ASAP7_75t_L g2432 ( 
.A(n_2065),
.B(n_1269),
.Y(n_2432)
);

INVx2_ASAP7_75t_L g2433 ( 
.A(n_2108),
.Y(n_2433)
);

NAND2xp5_ASAP7_75t_L g2434 ( 
.A(n_2070),
.B(n_1270),
.Y(n_2434)
);

O2A1O1Ixp5_ASAP7_75t_L g2435 ( 
.A1(n_2048),
.A2(n_2021),
.B(n_2016),
.C(n_1986),
.Y(n_2435)
);

INVx5_ASAP7_75t_L g2436 ( 
.A(n_2339),
.Y(n_2436)
);

OR2x2_ASAP7_75t_L g2437 ( 
.A(n_2080),
.B(n_1295),
.Y(n_2437)
);

HB1xp67_ASAP7_75t_L g2438 ( 
.A(n_2259),
.Y(n_2438)
);

AOI22xp5_ASAP7_75t_L g2439 ( 
.A1(n_2085),
.A2(n_1301),
.B1(n_1303),
.B2(n_1299),
.Y(n_2439)
);

INVx2_ASAP7_75t_L g2440 ( 
.A(n_2116),
.Y(n_2440)
);

NAND2xp5_ASAP7_75t_L g2441 ( 
.A(n_2074),
.B(n_1305),
.Y(n_2441)
);

HB1xp67_ASAP7_75t_L g2442 ( 
.A(n_2078),
.Y(n_2442)
);

NAND2xp5_ASAP7_75t_L g2443 ( 
.A(n_2075),
.B(n_1313),
.Y(n_2443)
);

INVx2_ASAP7_75t_L g2444 ( 
.A(n_2133),
.Y(n_2444)
);

NAND2xp5_ASAP7_75t_SL g2445 ( 
.A(n_2050),
.B(n_1920),
.Y(n_2445)
);

BUFx3_ASAP7_75t_L g2446 ( 
.A(n_2245),
.Y(n_2446)
);

O2A1O1Ixp33_ASAP7_75t_L g2447 ( 
.A1(n_2125),
.A2(n_1325),
.B(n_1355),
.C(n_1323),
.Y(n_2447)
);

AOI22xp33_ASAP7_75t_SL g2448 ( 
.A1(n_2143),
.A2(n_1372),
.B1(n_1375),
.B2(n_1360),
.Y(n_2448)
);

NAND2xp5_ASAP7_75t_L g2449 ( 
.A(n_2098),
.B(n_1376),
.Y(n_2449)
);

NOR2x1p5_ASAP7_75t_L g2450 ( 
.A(n_2067),
.B(n_1030),
.Y(n_2450)
);

NAND2xp5_ASAP7_75t_L g2451 ( 
.A(n_2058),
.B(n_1045),
.Y(n_2451)
);

INVx2_ASAP7_75t_L g2452 ( 
.A(n_2234),
.Y(n_2452)
);

NAND2xp5_ASAP7_75t_L g2453 ( 
.A(n_2058),
.B(n_1045),
.Y(n_2453)
);

NAND2xp5_ASAP7_75t_L g2454 ( 
.A(n_2084),
.B(n_1065),
.Y(n_2454)
);

INVx5_ASAP7_75t_L g2455 ( 
.A(n_2339),
.Y(n_2455)
);

NAND2xp5_ASAP7_75t_SL g2456 ( 
.A(n_2171),
.B(n_1920),
.Y(n_2456)
);

BUFx2_ASAP7_75t_L g2457 ( 
.A(n_2260),
.Y(n_2457)
);

NAND2xp5_ASAP7_75t_L g2458 ( 
.A(n_2091),
.B(n_1065),
.Y(n_2458)
);

INVx1_ASAP7_75t_L g2459 ( 
.A(n_2201),
.Y(n_2459)
);

INVx1_ASAP7_75t_L g2460 ( 
.A(n_2132),
.Y(n_2460)
);

NOR2xp33_ASAP7_75t_L g2461 ( 
.A(n_2152),
.B(n_2190),
.Y(n_2461)
);

INVx2_ASAP7_75t_L g2462 ( 
.A(n_2138),
.Y(n_2462)
);

INVx2_ASAP7_75t_L g2463 ( 
.A(n_2142),
.Y(n_2463)
);

INVx1_ASAP7_75t_L g2464 ( 
.A(n_2157),
.Y(n_2464)
);

CKINVDCx9p33_ASAP7_75t_R g2465 ( 
.A(n_2055),
.Y(n_2465)
);

NAND2xp5_ASAP7_75t_L g2466 ( 
.A(n_2092),
.B(n_1074),
.Y(n_2466)
);

AOI22xp33_ASAP7_75t_L g2467 ( 
.A1(n_2149),
.A2(n_930),
.B1(n_1102),
.B2(n_904),
.Y(n_2467)
);

INVx1_ASAP7_75t_L g2468 ( 
.A(n_2158),
.Y(n_2468)
);

HB1xp67_ASAP7_75t_L g2469 ( 
.A(n_2247),
.Y(n_2469)
);

AOI22xp5_ASAP7_75t_L g2470 ( 
.A1(n_2121),
.A2(n_1088),
.B1(n_1114),
.B2(n_1074),
.Y(n_2470)
);

INVx2_ASAP7_75t_L g2471 ( 
.A(n_2161),
.Y(n_2471)
);

HB1xp67_ASAP7_75t_L g2472 ( 
.A(n_2231),
.Y(n_2472)
);

AOI22xp5_ASAP7_75t_L g2473 ( 
.A1(n_2282),
.A2(n_1114),
.B1(n_1117),
.B2(n_1088),
.Y(n_2473)
);

NOR3xp33_ASAP7_75t_L g2474 ( 
.A(n_2079),
.B(n_2321),
.C(n_2331),
.Y(n_2474)
);

INVx1_ASAP7_75t_L g2475 ( 
.A(n_2168),
.Y(n_2475)
);

NAND2xp5_ASAP7_75t_SL g2476 ( 
.A(n_2242),
.B(n_1984),
.Y(n_2476)
);

AND2x4_ASAP7_75t_L g2477 ( 
.A(n_2166),
.B(n_1117),
.Y(n_2477)
);

INVx5_ASAP7_75t_L g2478 ( 
.A(n_2071),
.Y(n_2478)
);

AOI22xp33_ASAP7_75t_L g2479 ( 
.A1(n_2089),
.A2(n_930),
.B1(n_1102),
.B2(n_904),
.Y(n_2479)
);

INVx2_ASAP7_75t_L g2480 ( 
.A(n_2188),
.Y(n_2480)
);

NAND2xp5_ASAP7_75t_SL g2481 ( 
.A(n_2090),
.B(n_1984),
.Y(n_2481)
);

INVx2_ASAP7_75t_L g2482 ( 
.A(n_2197),
.Y(n_2482)
);

NAND2x1p5_ASAP7_75t_L g2483 ( 
.A(n_2071),
.B(n_1984),
.Y(n_2483)
);

NAND2x1_ASAP7_75t_L g2484 ( 
.A(n_2137),
.B(n_2022),
.Y(n_2484)
);

INVx2_ASAP7_75t_SL g2485 ( 
.A(n_2388),
.Y(n_2485)
);

NAND2xp5_ASAP7_75t_L g2486 ( 
.A(n_2096),
.B(n_1186),
.Y(n_2486)
);

NAND2xp5_ASAP7_75t_L g2487 ( 
.A(n_2277),
.B(n_2106),
.Y(n_2487)
);

AND3x2_ASAP7_75t_SL g2488 ( 
.A(n_2120),
.B(n_1193),
.C(n_1186),
.Y(n_2488)
);

INVx3_ASAP7_75t_L g2489 ( 
.A(n_2051),
.Y(n_2489)
);

NAND2xp5_ASAP7_75t_SL g2490 ( 
.A(n_2145),
.B(n_2002),
.Y(n_2490)
);

INVx1_ASAP7_75t_L g2491 ( 
.A(n_2213),
.Y(n_2491)
);

BUFx12f_ASAP7_75t_L g2492 ( 
.A(n_2100),
.Y(n_2492)
);

AND2x4_ASAP7_75t_L g2493 ( 
.A(n_2175),
.B(n_1193),
.Y(n_2493)
);

INVx1_ASAP7_75t_L g2494 ( 
.A(n_2217),
.Y(n_2494)
);

NAND2xp5_ASAP7_75t_SL g2495 ( 
.A(n_2124),
.B(n_2002),
.Y(n_2495)
);

NAND2xp5_ASAP7_75t_SL g2496 ( 
.A(n_2073),
.B(n_2002),
.Y(n_2496)
);

BUFx4f_ASAP7_75t_L g2497 ( 
.A(n_2330),
.Y(n_2497)
);

INVx1_ASAP7_75t_L g2498 ( 
.A(n_2219),
.Y(n_2498)
);

INVx1_ASAP7_75t_L g2499 ( 
.A(n_2224),
.Y(n_2499)
);

INVx2_ASAP7_75t_L g2500 ( 
.A(n_2205),
.Y(n_2500)
);

NAND2xp5_ASAP7_75t_L g2501 ( 
.A(n_2105),
.B(n_1231),
.Y(n_2501)
);

AND2x4_ASAP7_75t_L g2502 ( 
.A(n_2203),
.B(n_1231),
.Y(n_2502)
);

INVx2_ASAP7_75t_SL g2503 ( 
.A(n_2077),
.Y(n_2503)
);

INVx1_ASAP7_75t_L g2504 ( 
.A(n_2228),
.Y(n_2504)
);

INVx2_ASAP7_75t_L g2505 ( 
.A(n_2218),
.Y(n_2505)
);

INVx2_ASAP7_75t_SL g2506 ( 
.A(n_2324),
.Y(n_2506)
);

AOI22xp33_ASAP7_75t_L g2507 ( 
.A1(n_2181),
.A2(n_1102),
.B1(n_1161),
.B2(n_930),
.Y(n_2507)
);

INVx1_ASAP7_75t_L g2508 ( 
.A(n_2255),
.Y(n_2508)
);

NAND2xp5_ASAP7_75t_SL g2509 ( 
.A(n_2139),
.B(n_2027),
.Y(n_2509)
);

INVx2_ASAP7_75t_L g2510 ( 
.A(n_2229),
.Y(n_2510)
);

INVx3_ASAP7_75t_L g2511 ( 
.A(n_2095),
.Y(n_2511)
);

AND2x4_ASAP7_75t_L g2512 ( 
.A(n_2326),
.B(n_1289),
.Y(n_2512)
);

CKINVDCx5p33_ASAP7_75t_R g2513 ( 
.A(n_2082),
.Y(n_2513)
);

NAND2xp5_ASAP7_75t_SL g2514 ( 
.A(n_2148),
.B(n_2027),
.Y(n_2514)
);

INVx3_ASAP7_75t_SL g2515 ( 
.A(n_2336),
.Y(n_2515)
);

NAND2xp5_ASAP7_75t_L g2516 ( 
.A(n_2299),
.B(n_1289),
.Y(n_2516)
);

AND2x2_ASAP7_75t_L g2517 ( 
.A(n_2141),
.B(n_1293),
.Y(n_2517)
);

INVx1_ASAP7_75t_L g2518 ( 
.A(n_2237),
.Y(n_2518)
);

CKINVDCx5p33_ASAP7_75t_R g2519 ( 
.A(n_2315),
.Y(n_2519)
);

INVx5_ASAP7_75t_L g2520 ( 
.A(n_2137),
.Y(n_2520)
);

BUFx2_ASAP7_75t_L g2521 ( 
.A(n_2315),
.Y(n_2521)
);

AND3x1_ASAP7_75t_L g2522 ( 
.A(n_2196),
.B(n_1319),
.C(n_1293),
.Y(n_2522)
);

INVx2_ASAP7_75t_L g2523 ( 
.A(n_2239),
.Y(n_2523)
);

AOI22xp5_ASAP7_75t_L g2524 ( 
.A1(n_2282),
.A2(n_1334),
.B1(n_1319),
.B2(n_1161),
.Y(n_2524)
);

NAND2x1p5_ASAP7_75t_L g2525 ( 
.A(n_2377),
.B(n_2027),
.Y(n_2525)
);

AND2x4_ASAP7_75t_L g2526 ( 
.A(n_2274),
.B(n_1334),
.Y(n_2526)
);

INVx5_ASAP7_75t_L g2527 ( 
.A(n_2137),
.Y(n_2527)
);

AOI22xp5_ASAP7_75t_L g2528 ( 
.A1(n_2097),
.A2(n_1161),
.B1(n_1176),
.B2(n_1102),
.Y(n_2528)
);

AOI22xp33_ASAP7_75t_L g2529 ( 
.A1(n_2215),
.A2(n_1176),
.B1(n_1194),
.B2(n_1161),
.Y(n_2529)
);

NAND2xp5_ASAP7_75t_SL g2530 ( 
.A(n_2176),
.B(n_2026),
.Y(n_2530)
);

INVxp67_ASAP7_75t_SL g2531 ( 
.A(n_2222),
.Y(n_2531)
);

NAND2xp5_ASAP7_75t_SL g2532 ( 
.A(n_2204),
.B(n_2022),
.Y(n_2532)
);

INVx1_ASAP7_75t_L g2533 ( 
.A(n_2250),
.Y(n_2533)
);

NAND2xp5_ASAP7_75t_L g2534 ( 
.A(n_2286),
.B(n_0),
.Y(n_2534)
);

INVx2_ASAP7_75t_L g2535 ( 
.A(n_2256),
.Y(n_2535)
);

NAND2xp5_ASAP7_75t_SL g2536 ( 
.A(n_2066),
.B(n_2024),
.Y(n_2536)
);

BUFx3_ASAP7_75t_L g2537 ( 
.A(n_2280),
.Y(n_2537)
);

NAND2xp5_ASAP7_75t_SL g2538 ( 
.A(n_2216),
.B(n_2024),
.Y(n_2538)
);

INVx2_ASAP7_75t_L g2539 ( 
.A(n_2265),
.Y(n_2539)
);

NAND2xp5_ASAP7_75t_L g2540 ( 
.A(n_2293),
.B(n_2303),
.Y(n_2540)
);

CKINVDCx5p33_ASAP7_75t_R g2541 ( 
.A(n_2330),
.Y(n_2541)
);

INVx1_ASAP7_75t_L g2542 ( 
.A(n_2268),
.Y(n_2542)
);

CKINVDCx5p33_ASAP7_75t_R g2543 ( 
.A(n_2232),
.Y(n_2543)
);

INVx2_ASAP7_75t_L g2544 ( 
.A(n_2288),
.Y(n_2544)
);

NAND2xp5_ASAP7_75t_SL g2545 ( 
.A(n_2235),
.B(n_1176),
.Y(n_2545)
);

HB1xp67_ASAP7_75t_L g2546 ( 
.A(n_2270),
.Y(n_2546)
);

INVx1_ASAP7_75t_L g2547 ( 
.A(n_2300),
.Y(n_2547)
);

AND2x2_ASAP7_75t_L g2548 ( 
.A(n_2062),
.B(n_0),
.Y(n_2548)
);

BUFx3_ASAP7_75t_L g2549 ( 
.A(n_2253),
.Y(n_2549)
);

NAND2xp5_ASAP7_75t_SL g2550 ( 
.A(n_2230),
.B(n_1176),
.Y(n_2550)
);

AND2x4_ASAP7_75t_L g2551 ( 
.A(n_2261),
.B(n_2257),
.Y(n_2551)
);

AND2x4_ASAP7_75t_L g2552 ( 
.A(n_2275),
.B(n_1),
.Y(n_2552)
);

NAND2xp5_ASAP7_75t_L g2553 ( 
.A(n_2130),
.B(n_2),
.Y(n_2553)
);

AOI21xp5_ASAP7_75t_L g2554 ( 
.A1(n_2083),
.A2(n_1987),
.B(n_1978),
.Y(n_2554)
);

BUFx2_ASAP7_75t_L g2555 ( 
.A(n_2333),
.Y(n_2555)
);

AND2x2_ASAP7_75t_SL g2556 ( 
.A(n_2155),
.B(n_1194),
.Y(n_2556)
);

INVx1_ASAP7_75t_L g2557 ( 
.A(n_2319),
.Y(n_2557)
);

BUFx3_ASAP7_75t_L g2558 ( 
.A(n_2333),
.Y(n_2558)
);

INVx1_ASAP7_75t_L g2559 ( 
.A(n_2320),
.Y(n_2559)
);

INVx3_ASAP7_75t_L g2560 ( 
.A(n_2301),
.Y(n_2560)
);

OR2x6_ASAP7_75t_L g2561 ( 
.A(n_2298),
.B(n_2227),
.Y(n_2561)
);

AND2x2_ASAP7_75t_L g2562 ( 
.A(n_2064),
.B(n_2),
.Y(n_2562)
);

NAND2xp5_ASAP7_75t_SL g2563 ( 
.A(n_2230),
.B(n_1194),
.Y(n_2563)
);

OR2x2_ASAP7_75t_L g2564 ( 
.A(n_2110),
.B(n_3),
.Y(n_2564)
);

INVx1_ASAP7_75t_L g2565 ( 
.A(n_2327),
.Y(n_2565)
);

NAND2xp5_ASAP7_75t_SL g2566 ( 
.A(n_2230),
.B(n_1194),
.Y(n_2566)
);

OR2x6_ASAP7_75t_L g2567 ( 
.A(n_2052),
.B(n_1195),
.Y(n_2567)
);

NAND2xp5_ASAP7_75t_L g2568 ( 
.A(n_2130),
.B(n_3),
.Y(n_2568)
);

INVx2_ASAP7_75t_L g2569 ( 
.A(n_2374),
.Y(n_2569)
);

AND2x6_ASAP7_75t_L g2570 ( 
.A(n_2305),
.B(n_1195),
.Y(n_2570)
);

INVx1_ASAP7_75t_L g2571 ( 
.A(n_2345),
.Y(n_2571)
);

INVx1_ASAP7_75t_L g2572 ( 
.A(n_2349),
.Y(n_2572)
);

AND2x4_ASAP7_75t_L g2573 ( 
.A(n_2290),
.B(n_4),
.Y(n_2573)
);

INVx2_ASAP7_75t_L g2574 ( 
.A(n_2338),
.Y(n_2574)
);

NAND2xp5_ASAP7_75t_SL g2575 ( 
.A(n_2230),
.B(n_1195),
.Y(n_2575)
);

INVx4_ASAP7_75t_L g2576 ( 
.A(n_2238),
.Y(n_2576)
);

AO22x1_ASAP7_75t_L g2577 ( 
.A1(n_2115),
.A2(n_1321),
.B1(n_1195),
.B2(n_6),
.Y(n_2577)
);

NAND2xp5_ASAP7_75t_L g2578 ( 
.A(n_2177),
.B(n_4),
.Y(n_2578)
);

INVx1_ASAP7_75t_L g2579 ( 
.A(n_2263),
.Y(n_2579)
);

INVx1_ASAP7_75t_L g2580 ( 
.A(n_2069),
.Y(n_2580)
);

O2A1O1Ixp5_ASAP7_75t_L g2581 ( 
.A1(n_2049),
.A2(n_1995),
.B(n_1998),
.C(n_1992),
.Y(n_2581)
);

AND2x2_ASAP7_75t_SL g2582 ( 
.A(n_2191),
.B(n_2198),
.Y(n_2582)
);

NAND2xp5_ASAP7_75t_L g2583 ( 
.A(n_2308),
.B(n_4),
.Y(n_2583)
);

INVx1_ASAP7_75t_L g2584 ( 
.A(n_2069),
.Y(n_2584)
);

INVx4_ASAP7_75t_L g2585 ( 
.A(n_2238),
.Y(n_2585)
);

INVx1_ASAP7_75t_L g2586 ( 
.A(n_2187),
.Y(n_2586)
);

NAND2xp5_ASAP7_75t_L g2587 ( 
.A(n_2177),
.B(n_5),
.Y(n_2587)
);

INVx2_ASAP7_75t_SL g2588 ( 
.A(n_2332),
.Y(n_2588)
);

AND2x6_ASAP7_75t_L g2589 ( 
.A(n_2317),
.B(n_2222),
.Y(n_2589)
);

BUFx3_ASAP7_75t_L g2590 ( 
.A(n_2333),
.Y(n_2590)
);

INVx1_ASAP7_75t_L g2591 ( 
.A(n_2187),
.Y(n_2591)
);

INVx1_ASAP7_75t_L g2592 ( 
.A(n_2285),
.Y(n_2592)
);

INVx3_ASAP7_75t_L g2593 ( 
.A(n_2301),
.Y(n_2593)
);

INVx3_ASAP7_75t_L g2594 ( 
.A(n_2251),
.Y(n_2594)
);

NAND2xp5_ASAP7_75t_SL g2595 ( 
.A(n_2230),
.B(n_1321),
.Y(n_2595)
);

NAND2xp5_ASAP7_75t_L g2596 ( 
.A(n_2289),
.B(n_5),
.Y(n_2596)
);

NAND2xp5_ASAP7_75t_L g2597 ( 
.A(n_2119),
.B(n_6),
.Y(n_2597)
);

INVx2_ASAP7_75t_SL g2598 ( 
.A(n_2344),
.Y(n_2598)
);

OR2x6_ASAP7_75t_L g2599 ( 
.A(n_2054),
.B(n_1321),
.Y(n_2599)
);

BUFx2_ASAP7_75t_L g2600 ( 
.A(n_2333),
.Y(n_2600)
);

NAND2xp5_ASAP7_75t_L g2601 ( 
.A(n_2192),
.B(n_6),
.Y(n_2601)
);

INVx1_ASAP7_75t_L g2602 ( 
.A(n_2192),
.Y(n_2602)
);

NAND2xp5_ASAP7_75t_L g2603 ( 
.A(n_2199),
.B(n_7),
.Y(n_2603)
);

NOR3xp33_ASAP7_75t_SL g2604 ( 
.A(n_2325),
.B(n_8),
.C(n_9),
.Y(n_2604)
);

NOR2xp33_ASAP7_75t_L g2605 ( 
.A(n_2202),
.B(n_8),
.Y(n_2605)
);

BUFx4f_ASAP7_75t_L g2606 ( 
.A(n_2137),
.Y(n_2606)
);

AND2x2_ASAP7_75t_L g2607 ( 
.A(n_2056),
.B(n_9),
.Y(n_2607)
);

INVx1_ASAP7_75t_L g2608 ( 
.A(n_2199),
.Y(n_2608)
);

INVxp33_ASAP7_75t_L g2609 ( 
.A(n_2144),
.Y(n_2609)
);

AOI22xp33_ASAP7_75t_L g2610 ( 
.A1(n_2159),
.A2(n_1321),
.B1(n_1957),
.B2(n_1947),
.Y(n_2610)
);

INVxp67_ASAP7_75t_SL g2611 ( 
.A(n_2222),
.Y(n_2611)
);

INVx1_ASAP7_75t_L g2612 ( 
.A(n_2355),
.Y(n_2612)
);

AOI22xp33_ASAP7_75t_L g2613 ( 
.A1(n_2117),
.A2(n_2294),
.B1(n_2266),
.B2(n_2093),
.Y(n_2613)
);

CKINVDCx20_ASAP7_75t_R g2614 ( 
.A(n_2153),
.Y(n_2614)
);

INVx5_ASAP7_75t_L g2615 ( 
.A(n_2251),
.Y(n_2615)
);

NAND2xp5_ASAP7_75t_L g2616 ( 
.A(n_2276),
.B(n_10),
.Y(n_2616)
);

NAND2xp5_ASAP7_75t_L g2617 ( 
.A(n_2361),
.B(n_10),
.Y(n_2617)
);

AND2x4_ASAP7_75t_L g2618 ( 
.A(n_2262),
.B(n_10),
.Y(n_2618)
);

NOR2xp33_ASAP7_75t_L g2619 ( 
.A(n_2340),
.B(n_11),
.Y(n_2619)
);

AOI22xp5_ASAP7_75t_L g2620 ( 
.A1(n_2361),
.A2(n_1962),
.B1(n_1963),
.B2(n_1960),
.Y(n_2620)
);

NAND2xp5_ASAP7_75t_L g2621 ( 
.A(n_2276),
.B(n_2279),
.Y(n_2621)
);

INVx2_ASAP7_75t_SL g2622 ( 
.A(n_2061),
.Y(n_2622)
);

NOR2x1_ASAP7_75t_R g2623 ( 
.A(n_2109),
.B(n_11),
.Y(n_2623)
);

A2O1A1Ixp33_ASAP7_75t_L g2624 ( 
.A1(n_2376),
.A2(n_1966),
.B(n_1968),
.C(n_1964),
.Y(n_2624)
);

INVx1_ASAP7_75t_L g2625 ( 
.A(n_2356),
.Y(n_2625)
);

AOI22xp33_ASAP7_75t_L g2626 ( 
.A1(n_2059),
.A2(n_2086),
.B1(n_2094),
.B2(n_2087),
.Y(n_2626)
);

INVx1_ASAP7_75t_L g2627 ( 
.A(n_2364),
.Y(n_2627)
);

BUFx6f_ASAP7_75t_L g2628 ( 
.A(n_2251),
.Y(n_2628)
);

OR2x6_ASAP7_75t_L g2629 ( 
.A(n_2151),
.B(n_1977),
.Y(n_2629)
);

INVx1_ASAP7_75t_L g2630 ( 
.A(n_2365),
.Y(n_2630)
);

BUFx12f_ASAP7_75t_L g2631 ( 
.A(n_2378),
.Y(n_2631)
);

INVx2_ASAP7_75t_L g2632 ( 
.A(n_2370),
.Y(n_2632)
);

AOI22xp33_ASAP7_75t_L g2633 ( 
.A1(n_2103),
.A2(n_1983),
.B1(n_1988),
.B2(n_1981),
.Y(n_2633)
);

INVx2_ASAP7_75t_L g2634 ( 
.A(n_2113),
.Y(n_2634)
);

INVx1_ASAP7_75t_L g2635 ( 
.A(n_2304),
.Y(n_2635)
);

NAND2x1_ASAP7_75t_L g2636 ( 
.A(n_2278),
.B(n_1990),
.Y(n_2636)
);

NAND2xp5_ASAP7_75t_L g2637 ( 
.A(n_2225),
.B(n_11),
.Y(n_2637)
);

OR2x6_ASAP7_75t_L g2638 ( 
.A(n_2170),
.B(n_2006),
.Y(n_2638)
);

NOR2xp33_ASAP7_75t_R g2639 ( 
.A(n_2328),
.B(n_12),
.Y(n_2639)
);

NAND2xp5_ASAP7_75t_L g2640 ( 
.A(n_2226),
.B(n_12),
.Y(n_2640)
);

NOR2xp33_ASAP7_75t_L g2641 ( 
.A(n_2169),
.B(n_13),
.Y(n_2641)
);

NAND2xp5_ASAP7_75t_L g2642 ( 
.A(n_2240),
.B(n_13),
.Y(n_2642)
);

INVx5_ASAP7_75t_L g2643 ( 
.A(n_2278),
.Y(n_2643)
);

INVxp67_ASAP7_75t_L g2644 ( 
.A(n_2104),
.Y(n_2644)
);

AND2x4_ASAP7_75t_L g2645 ( 
.A(n_2249),
.B(n_14),
.Y(n_2645)
);

NAND2xp5_ASAP7_75t_L g2646 ( 
.A(n_2241),
.B(n_15),
.Y(n_2646)
);

AND2x2_ASAP7_75t_L g2647 ( 
.A(n_2173),
.B(n_2200),
.Y(n_2647)
);

AND2x4_ASAP7_75t_L g2648 ( 
.A(n_2292),
.B(n_2186),
.Y(n_2648)
);

OAI21xp33_ASAP7_75t_SL g2649 ( 
.A1(n_2391),
.A2(n_23),
.B(n_15),
.Y(n_2649)
);

AOI22xp33_ASAP7_75t_L g2650 ( 
.A1(n_2272),
.A2(n_2014),
.B1(n_2017),
.B2(n_2007),
.Y(n_2650)
);

BUFx6f_ASAP7_75t_L g2651 ( 
.A(n_2278),
.Y(n_2651)
);

INVx2_ASAP7_75t_L g2652 ( 
.A(n_2114),
.Y(n_2652)
);

AOI22xp33_ASAP7_75t_L g2653 ( 
.A1(n_2273),
.A2(n_2025),
.B1(n_18),
.B2(n_16),
.Y(n_2653)
);

BUFx6f_ASAP7_75t_L g2654 ( 
.A(n_2346),
.Y(n_2654)
);

AND2x2_ASAP7_75t_L g2655 ( 
.A(n_2211),
.B(n_17),
.Y(n_2655)
);

AND2x4_ASAP7_75t_L g2656 ( 
.A(n_2379),
.B(n_17),
.Y(n_2656)
);

INVx1_ASAP7_75t_L g2657 ( 
.A(n_2393),
.Y(n_2657)
);

NAND2xp5_ASAP7_75t_L g2658 ( 
.A(n_2281),
.B(n_18),
.Y(n_2658)
);

INVxp67_ASAP7_75t_L g2659 ( 
.A(n_2220),
.Y(n_2659)
);

NAND2x1p5_ASAP7_75t_L g2660 ( 
.A(n_2346),
.B(n_18),
.Y(n_2660)
);

NAND2xp5_ASAP7_75t_SL g2661 ( 
.A(n_2346),
.B(n_20),
.Y(n_2661)
);

INVx2_ASAP7_75t_L g2662 ( 
.A(n_2312),
.Y(n_2662)
);

NOR2x2_ASAP7_75t_L g2663 ( 
.A(n_2102),
.B(n_19),
.Y(n_2663)
);

O2A1O1Ixp5_ASAP7_75t_L g2664 ( 
.A1(n_2318),
.A2(n_21),
.B(n_19),
.C(n_20),
.Y(n_2664)
);

INVx1_ASAP7_75t_L g2665 ( 
.A(n_2393),
.Y(n_2665)
);

NOR2xp33_ASAP7_75t_R g2666 ( 
.A(n_2348),
.B(n_21),
.Y(n_2666)
);

INVx2_ASAP7_75t_L g2667 ( 
.A(n_2112),
.Y(n_2667)
);

NOR2x2_ASAP7_75t_L g2668 ( 
.A(n_2214),
.B(n_21),
.Y(n_2668)
);

INVx2_ASAP7_75t_L g2669 ( 
.A(n_2389),
.Y(n_2669)
);

AOI22xp5_ASAP7_75t_L g2670 ( 
.A1(n_2129),
.A2(n_2083),
.B1(n_2287),
.B2(n_2210),
.Y(n_2670)
);

NAND2xp5_ASAP7_75t_SL g2671 ( 
.A(n_2126),
.B(n_23),
.Y(n_2671)
);

AND2x4_ASAP7_75t_L g2672 ( 
.A(n_2357),
.B(n_22),
.Y(n_2672)
);

NAND2xp5_ASAP7_75t_L g2673 ( 
.A(n_2279),
.B(n_23),
.Y(n_2673)
);

AND2x2_ASAP7_75t_L g2674 ( 
.A(n_2233),
.B(n_2164),
.Y(n_2674)
);

INVx2_ASAP7_75t_L g2675 ( 
.A(n_2341),
.Y(n_2675)
);

INVx2_ASAP7_75t_L g2676 ( 
.A(n_2341),
.Y(n_2676)
);

INVx1_ASAP7_75t_L g2677 ( 
.A(n_2207),
.Y(n_2677)
);

INVx2_ASAP7_75t_L g2678 ( 
.A(n_2395),
.Y(n_2678)
);

NAND2xp5_ASAP7_75t_L g2679 ( 
.A(n_2127),
.B(n_24),
.Y(n_2679)
);

AND3x2_ASAP7_75t_SL g2680 ( 
.A(n_2131),
.B(n_24),
.C(n_25),
.Y(n_2680)
);

NOR2x1p5_ASAP7_75t_L g2681 ( 
.A(n_2128),
.B(n_24),
.Y(n_2681)
);

NAND2xp5_ASAP7_75t_L g2682 ( 
.A(n_2209),
.B(n_25),
.Y(n_2682)
);

INVx1_ASAP7_75t_L g2683 ( 
.A(n_2134),
.Y(n_2683)
);

BUFx3_ASAP7_75t_L g2684 ( 
.A(n_2396),
.Y(n_2684)
);

INVx1_ASAP7_75t_L g2685 ( 
.A(n_2135),
.Y(n_2685)
);

NOR3xp33_ASAP7_75t_SL g2686 ( 
.A(n_2254),
.B(n_25),
.C(n_26),
.Y(n_2686)
);

NAND2xp33_ASAP7_75t_L g2687 ( 
.A(n_2391),
.B(n_28),
.Y(n_2687)
);

NAND2xp5_ASAP7_75t_L g2688 ( 
.A(n_2392),
.B(n_27),
.Y(n_2688)
);

NOR2xp67_ASAP7_75t_L g2689 ( 
.A(n_2334),
.B(n_27),
.Y(n_2689)
);

INVx1_ASAP7_75t_L g2690 ( 
.A(n_2146),
.Y(n_2690)
);

NAND2xp5_ASAP7_75t_SL g2691 ( 
.A(n_2267),
.B(n_29),
.Y(n_2691)
);

NAND2xp5_ASAP7_75t_SL g2692 ( 
.A(n_2269),
.B(n_2271),
.Y(n_2692)
);

NOR2xp33_ASAP7_75t_L g2693 ( 
.A(n_2236),
.B(n_28),
.Y(n_2693)
);

INVx1_ASAP7_75t_L g2694 ( 
.A(n_2147),
.Y(n_2694)
);

INVx1_ASAP7_75t_L g2695 ( 
.A(n_2160),
.Y(n_2695)
);

INVx2_ASAP7_75t_L g2696 ( 
.A(n_2394),
.Y(n_2696)
);

INVx1_ASAP7_75t_L g2697 ( 
.A(n_2162),
.Y(n_2697)
);

BUFx6f_ASAP7_75t_L g2698 ( 
.A(n_2123),
.Y(n_2698)
);

INVx1_ASAP7_75t_L g2699 ( 
.A(n_2167),
.Y(n_2699)
);

NAND2xp5_ASAP7_75t_L g2700 ( 
.A(n_2360),
.B(n_28),
.Y(n_2700)
);

OR2x6_ASAP7_75t_L g2701 ( 
.A(n_2384),
.B(n_29),
.Y(n_2701)
);

INVx2_ASAP7_75t_L g2702 ( 
.A(n_2154),
.Y(n_2702)
);

A2O1A1Ixp33_ASAP7_75t_L g2703 ( 
.A1(n_2334),
.A2(n_31),
.B(n_29),
.C(n_30),
.Y(n_2703)
);

AND2x2_ASAP7_75t_L g2704 ( 
.A(n_2212),
.B(n_30),
.Y(n_2704)
);

NAND2xp5_ASAP7_75t_L g2705 ( 
.A(n_2369),
.B(n_30),
.Y(n_2705)
);

NAND2xp5_ASAP7_75t_L g2706 ( 
.A(n_2118),
.B(n_2221),
.Y(n_2706)
);

AND2x6_ASAP7_75t_L g2707 ( 
.A(n_2342),
.B(n_31),
.Y(n_2707)
);

NAND2xp5_ASAP7_75t_L g2708 ( 
.A(n_2140),
.B(n_2387),
.Y(n_2708)
);

AOI22xp33_ASAP7_75t_L g2709 ( 
.A1(n_2283),
.A2(n_34),
.B1(n_32),
.B2(n_33),
.Y(n_2709)
);

INVx3_ASAP7_75t_L g2710 ( 
.A(n_2335),
.Y(n_2710)
);

INVx2_ASAP7_75t_SL g2711 ( 
.A(n_2385),
.Y(n_2711)
);

BUFx5_ASAP7_75t_L g2712 ( 
.A(n_2081),
.Y(n_2712)
);

NAND2xp33_ASAP7_75t_SL g2713 ( 
.A(n_2284),
.B(n_33),
.Y(n_2713)
);

AND2x4_ASAP7_75t_L g2714 ( 
.A(n_2362),
.B(n_33),
.Y(n_2714)
);

NAND2xp5_ASAP7_75t_L g2715 ( 
.A(n_2243),
.B(n_2246),
.Y(n_2715)
);

INVx4_ASAP7_75t_L g2716 ( 
.A(n_2111),
.Y(n_2716)
);

AOI22xp5_ASAP7_75t_L g2717 ( 
.A1(n_2297),
.A2(n_2248),
.B1(n_2189),
.B2(n_2193),
.Y(n_2717)
);

AND2x2_ASAP7_75t_L g2718 ( 
.A(n_2380),
.B(n_34),
.Y(n_2718)
);

INVxp67_ASAP7_75t_L g2719 ( 
.A(n_2306),
.Y(n_2719)
);

NAND2xp5_ASAP7_75t_SL g2720 ( 
.A(n_2353),
.B(n_36),
.Y(n_2720)
);

INVx2_ASAP7_75t_L g2721 ( 
.A(n_2252),
.Y(n_2721)
);

NAND2xp5_ASAP7_75t_SL g2722 ( 
.A(n_2258),
.B(n_36),
.Y(n_2722)
);

INVx1_ASAP7_75t_L g2723 ( 
.A(n_2264),
.Y(n_2723)
);

CKINVDCx6p67_ASAP7_75t_R g2724 ( 
.A(n_2386),
.Y(n_2724)
);

NAND2xp5_ASAP7_75t_SL g2725 ( 
.A(n_2314),
.B(n_36),
.Y(n_2725)
);

INVx5_ASAP7_75t_L g2726 ( 
.A(n_2076),
.Y(n_2726)
);

INVx2_ASAP7_75t_L g2727 ( 
.A(n_2302),
.Y(n_2727)
);

AOI22xp33_ASAP7_75t_L g2728 ( 
.A1(n_2223),
.A2(n_38),
.B1(n_35),
.B2(n_37),
.Y(n_2728)
);

NAND2xp5_ASAP7_75t_L g2729 ( 
.A(n_2354),
.B(n_35),
.Y(n_2729)
);

OR2x2_ASAP7_75t_L g2730 ( 
.A(n_2307),
.B(n_35),
.Y(n_2730)
);

OR2x2_ASAP7_75t_L g2731 ( 
.A(n_2309),
.B(n_37),
.Y(n_2731)
);

INVx1_ASAP7_75t_L g2732 ( 
.A(n_2381),
.Y(n_2732)
);

AND2x4_ASAP7_75t_L g2733 ( 
.A(n_2366),
.B(n_2368),
.Y(n_2733)
);

INVx2_ASAP7_75t_L g2734 ( 
.A(n_2382),
.Y(n_2734)
);

INVx1_ASAP7_75t_L g2735 ( 
.A(n_2316),
.Y(n_2735)
);

INVx1_ASAP7_75t_L g2736 ( 
.A(n_2323),
.Y(n_2736)
);

INVx1_ASAP7_75t_L g2737 ( 
.A(n_2337),
.Y(n_2737)
);

NOR2xp33_ASAP7_75t_L g2738 ( 
.A(n_2313),
.B(n_38),
.Y(n_2738)
);

AND2x2_ASAP7_75t_L g2739 ( 
.A(n_2343),
.B(n_38),
.Y(n_2739)
);

HB1xp67_ASAP7_75t_L g2740 ( 
.A(n_2194),
.Y(n_2740)
);

INVx1_ASAP7_75t_L g2741 ( 
.A(n_2351),
.Y(n_2741)
);

INVx1_ASAP7_75t_L g2742 ( 
.A(n_2352),
.Y(n_2742)
);

NOR2xp33_ASAP7_75t_L g2743 ( 
.A(n_2373),
.B(n_39),
.Y(n_2743)
);

AOI22xp33_ASAP7_75t_L g2744 ( 
.A1(n_2295),
.A2(n_41),
.B1(n_39),
.B2(n_40),
.Y(n_2744)
);

NAND2xp5_ASAP7_75t_SL g2745 ( 
.A(n_2291),
.B(n_42),
.Y(n_2745)
);

INVx4_ASAP7_75t_L g2746 ( 
.A(n_2206),
.Y(n_2746)
);

CKINVDCx5p33_ASAP7_75t_R g2747 ( 
.A(n_2383),
.Y(n_2747)
);

AND2x4_ASAP7_75t_L g2748 ( 
.A(n_2375),
.B(n_40),
.Y(n_2748)
);

NAND2xp5_ASAP7_75t_SL g2749 ( 
.A(n_2359),
.B(n_2363),
.Y(n_2749)
);

INVx2_ASAP7_75t_L g2750 ( 
.A(n_2358),
.Y(n_2750)
);

NAND2xp5_ASAP7_75t_L g2751 ( 
.A(n_2296),
.B(n_40),
.Y(n_2751)
);

NAND2xp5_ASAP7_75t_SL g2752 ( 
.A(n_2367),
.B(n_44),
.Y(n_2752)
);

INVx4_ASAP7_75t_L g2753 ( 
.A(n_2081),
.Y(n_2753)
);

BUFx2_ASAP7_75t_L g2754 ( 
.A(n_2371),
.Y(n_2754)
);

NOR2x1p5_ASAP7_75t_L g2755 ( 
.A(n_2372),
.B(n_42),
.Y(n_2755)
);

INVx3_ASAP7_75t_L g2756 ( 
.A(n_2322),
.Y(n_2756)
);

INVx2_ASAP7_75t_SL g2757 ( 
.A(n_2390),
.Y(n_2757)
);

NAND2xp5_ASAP7_75t_L g2758 ( 
.A(n_2310),
.B(n_44),
.Y(n_2758)
);

NAND2xp5_ASAP7_75t_L g2759 ( 
.A(n_2311),
.B(n_44),
.Y(n_2759)
);

HB1xp67_ASAP7_75t_L g2760 ( 
.A(n_2195),
.Y(n_2760)
);

INVx2_ASAP7_75t_L g2761 ( 
.A(n_2358),
.Y(n_2761)
);

INVx1_ASAP7_75t_L g2762 ( 
.A(n_2347),
.Y(n_2762)
);

NAND2xp5_ASAP7_75t_SL g2763 ( 
.A(n_2208),
.B(n_46),
.Y(n_2763)
);

AOI22xp5_ASAP7_75t_L g2764 ( 
.A1(n_2350),
.A2(n_47),
.B1(n_45),
.B2(n_46),
.Y(n_2764)
);

AOI22xp33_ASAP7_75t_L g2765 ( 
.A1(n_2372),
.A2(n_47),
.B1(n_45),
.B2(n_46),
.Y(n_2765)
);

BUFx6f_ASAP7_75t_L g2766 ( 
.A(n_2238),
.Y(n_2766)
);

CKINVDCx20_ASAP7_75t_R g2767 ( 
.A(n_2245),
.Y(n_2767)
);

NOR2xp33_ASAP7_75t_L g2768 ( 
.A(n_2072),
.B(n_45),
.Y(n_2768)
);

INVx2_ASAP7_75t_L g2769 ( 
.A(n_2172),
.Y(n_2769)
);

NAND2xp5_ASAP7_75t_L g2770 ( 
.A(n_2053),
.B(n_47),
.Y(n_2770)
);

INVx3_ASAP7_75t_L g2771 ( 
.A(n_2060),
.Y(n_2771)
);

BUFx6f_ASAP7_75t_L g2772 ( 
.A(n_2238),
.Y(n_2772)
);

AOI22xp5_ASAP7_75t_L g2773 ( 
.A1(n_2060),
.A2(n_50),
.B1(n_48),
.B2(n_49),
.Y(n_2773)
);

NAND2xp5_ASAP7_75t_L g2774 ( 
.A(n_2053),
.B(n_48),
.Y(n_2774)
);

BUFx3_ASAP7_75t_L g2775 ( 
.A(n_2245),
.Y(n_2775)
);

NAND2xp5_ASAP7_75t_SL g2776 ( 
.A(n_2088),
.B(n_49),
.Y(n_2776)
);

NAND3xp33_ASAP7_75t_L g2777 ( 
.A(n_2129),
.B(n_48),
.C(n_49),
.Y(n_2777)
);

AND2x2_ASAP7_75t_L g2778 ( 
.A(n_2122),
.B(n_50),
.Y(n_2778)
);

INVx2_ASAP7_75t_L g2779 ( 
.A(n_2172),
.Y(n_2779)
);

NAND2xp5_ASAP7_75t_L g2780 ( 
.A(n_2053),
.B(n_50),
.Y(n_2780)
);

AND2x4_ASAP7_75t_L g2781 ( 
.A(n_2060),
.B(n_51),
.Y(n_2781)
);

NAND2xp5_ASAP7_75t_L g2782 ( 
.A(n_2060),
.B(n_51),
.Y(n_2782)
);

INVx2_ASAP7_75t_L g2783 ( 
.A(n_2172),
.Y(n_2783)
);

AOI22xp5_ASAP7_75t_L g2784 ( 
.A1(n_2060),
.A2(n_54),
.B1(n_52),
.B2(n_53),
.Y(n_2784)
);

INVx1_ASAP7_75t_L g2785 ( 
.A(n_2178),
.Y(n_2785)
);

INVx1_ASAP7_75t_L g2786 ( 
.A(n_2178),
.Y(n_2786)
);

AND2x4_ASAP7_75t_L g2787 ( 
.A(n_2060),
.B(n_52),
.Y(n_2787)
);

INVx2_ASAP7_75t_L g2788 ( 
.A(n_2172),
.Y(n_2788)
);

NAND2xp5_ASAP7_75t_L g2789 ( 
.A(n_2060),
.B(n_54),
.Y(n_2789)
);

HB1xp67_ASAP7_75t_L g2790 ( 
.A(n_2063),
.Y(n_2790)
);

NAND2xp5_ASAP7_75t_L g2791 ( 
.A(n_2060),
.B(n_54),
.Y(n_2791)
);

OAI21xp33_ASAP7_75t_L g2792 ( 
.A1(n_2107),
.A2(n_55),
.B(n_56),
.Y(n_2792)
);

CKINVDCx5p33_ASAP7_75t_R g2793 ( 
.A(n_2067),
.Y(n_2793)
);

AO22x1_ASAP7_75t_L g2794 ( 
.A1(n_2055),
.A2(n_58),
.B1(n_59),
.B2(n_57),
.Y(n_2794)
);

NAND2xp5_ASAP7_75t_L g2795 ( 
.A(n_2053),
.B(n_56),
.Y(n_2795)
);

BUFx2_ASAP7_75t_L g2796 ( 
.A(n_2063),
.Y(n_2796)
);

INVx2_ASAP7_75t_L g2797 ( 
.A(n_2172),
.Y(n_2797)
);

BUFx6f_ASAP7_75t_L g2798 ( 
.A(n_2238),
.Y(n_2798)
);

INVx1_ASAP7_75t_L g2799 ( 
.A(n_2178),
.Y(n_2799)
);

INVx2_ASAP7_75t_L g2800 ( 
.A(n_2172),
.Y(n_2800)
);

NAND2xp5_ASAP7_75t_L g2801 ( 
.A(n_2053),
.B(n_57),
.Y(n_2801)
);

BUFx6f_ASAP7_75t_L g2802 ( 
.A(n_2238),
.Y(n_2802)
);

INVx1_ASAP7_75t_L g2803 ( 
.A(n_2178),
.Y(n_2803)
);

NOR2xp33_ASAP7_75t_L g2804 ( 
.A(n_2072),
.B(n_58),
.Y(n_2804)
);

NAND2xp5_ASAP7_75t_L g2805 ( 
.A(n_2053),
.B(n_58),
.Y(n_2805)
);

AND2x4_ASAP7_75t_L g2806 ( 
.A(n_2060),
.B(n_59),
.Y(n_2806)
);

NAND2xp5_ASAP7_75t_L g2807 ( 
.A(n_2053),
.B(n_60),
.Y(n_2807)
);

BUFx2_ASAP7_75t_L g2808 ( 
.A(n_2063),
.Y(n_2808)
);

INVx5_ASAP7_75t_L g2809 ( 
.A(n_2136),
.Y(n_2809)
);

INVx1_ASAP7_75t_L g2810 ( 
.A(n_2178),
.Y(n_2810)
);

NAND2xp5_ASAP7_75t_L g2811 ( 
.A(n_2060),
.B(n_61),
.Y(n_2811)
);

BUFx2_ASAP7_75t_L g2812 ( 
.A(n_2063),
.Y(n_2812)
);

NAND2xp5_ASAP7_75t_L g2813 ( 
.A(n_2060),
.B(n_61),
.Y(n_2813)
);

BUFx6f_ASAP7_75t_L g2814 ( 
.A(n_2238),
.Y(n_2814)
);

NAND2xp5_ASAP7_75t_L g2815 ( 
.A(n_2060),
.B(n_62),
.Y(n_2815)
);

NAND2xp5_ASAP7_75t_L g2816 ( 
.A(n_2053),
.B(n_62),
.Y(n_2816)
);

INVxp67_ASAP7_75t_L g2817 ( 
.A(n_2063),
.Y(n_2817)
);

BUFx6f_ASAP7_75t_L g2818 ( 
.A(n_2238),
.Y(n_2818)
);

INVx1_ASAP7_75t_L g2819 ( 
.A(n_2178),
.Y(n_2819)
);

NAND2xp5_ASAP7_75t_L g2820 ( 
.A(n_2053),
.B(n_63),
.Y(n_2820)
);

NAND2xp5_ASAP7_75t_L g2821 ( 
.A(n_2053),
.B(n_63),
.Y(n_2821)
);

INVx2_ASAP7_75t_L g2822 ( 
.A(n_2172),
.Y(n_2822)
);

NOR3xp33_ASAP7_75t_SL g2823 ( 
.A(n_2067),
.B(n_64),
.C(n_65),
.Y(n_2823)
);

NAND2xp5_ASAP7_75t_L g2824 ( 
.A(n_2053),
.B(n_65),
.Y(n_2824)
);

INVx1_ASAP7_75t_SL g2825 ( 
.A(n_2063),
.Y(n_2825)
);

NAND2xp5_ASAP7_75t_L g2826 ( 
.A(n_2053),
.B(n_65),
.Y(n_2826)
);

NAND2xp5_ASAP7_75t_L g2827 ( 
.A(n_2053),
.B(n_66),
.Y(n_2827)
);

NAND2xp5_ASAP7_75t_L g2828 ( 
.A(n_2053),
.B(n_66),
.Y(n_2828)
);

AOI22xp5_ASAP7_75t_L g2829 ( 
.A1(n_2060),
.A2(n_68),
.B1(n_66),
.B2(n_67),
.Y(n_2829)
);

NAND2xp5_ASAP7_75t_SL g2830 ( 
.A(n_2088),
.B(n_69),
.Y(n_2830)
);

NAND2xp5_ASAP7_75t_L g2831 ( 
.A(n_2053),
.B(n_68),
.Y(n_2831)
);

INVx1_ASAP7_75t_L g2832 ( 
.A(n_2178),
.Y(n_2832)
);

NAND2xp5_ASAP7_75t_SL g2833 ( 
.A(n_2088),
.B(n_70),
.Y(n_2833)
);

OAI22xp5_ASAP7_75t_SL g2834 ( 
.A1(n_2055),
.A2(n_71),
.B1(n_69),
.B2(n_70),
.Y(n_2834)
);

OAI22xp33_ASAP7_75t_L g2835 ( 
.A1(n_2088),
.A2(n_72),
.B1(n_69),
.B2(n_71),
.Y(n_2835)
);

NOR3xp33_ASAP7_75t_SL g2836 ( 
.A(n_2067),
.B(n_71),
.C(n_72),
.Y(n_2836)
);

CKINVDCx5p33_ASAP7_75t_R g2837 ( 
.A(n_2067),
.Y(n_2837)
);

CKINVDCx5p33_ASAP7_75t_R g2838 ( 
.A(n_2067),
.Y(n_2838)
);

AND2x4_ASAP7_75t_L g2839 ( 
.A(n_2060),
.B(n_72),
.Y(n_2839)
);

NAND2xp5_ASAP7_75t_L g2840 ( 
.A(n_2060),
.B(n_73),
.Y(n_2840)
);

NAND2xp5_ASAP7_75t_SL g2841 ( 
.A(n_2088),
.B(n_74),
.Y(n_2841)
);

AOI22xp33_ASAP7_75t_L g2842 ( 
.A1(n_2150),
.A2(n_75),
.B1(n_73),
.B2(n_74),
.Y(n_2842)
);

BUFx8_ASAP7_75t_L g2843 ( 
.A(n_2082),
.Y(n_2843)
);

NOR3xp33_ASAP7_75t_L g2844 ( 
.A(n_2107),
.B(n_76),
.C(n_75),
.Y(n_2844)
);

INVx3_ASAP7_75t_L g2845 ( 
.A(n_2060),
.Y(n_2845)
);

NOR2xp33_ASAP7_75t_L g2846 ( 
.A(n_2072),
.B(n_73),
.Y(n_2846)
);

NOR2x1p5_ASAP7_75t_L g2847 ( 
.A(n_2067),
.B(n_75),
.Y(n_2847)
);

NAND2xp5_ASAP7_75t_SL g2848 ( 
.A(n_2088),
.B(n_78),
.Y(n_2848)
);

AOI22xp33_ASAP7_75t_SL g2849 ( 
.A1(n_2088),
.A2(n_79),
.B1(n_77),
.B2(n_78),
.Y(n_2849)
);

INVx1_ASAP7_75t_L g2850 ( 
.A(n_2178),
.Y(n_2850)
);

BUFx2_ASAP7_75t_L g2851 ( 
.A(n_2063),
.Y(n_2851)
);

BUFx4f_ASAP7_75t_SL g2852 ( 
.A(n_2245),
.Y(n_2852)
);

OR2x2_ASAP7_75t_L g2853 ( 
.A(n_2080),
.B(n_79),
.Y(n_2853)
);

NOR2xp33_ASAP7_75t_SL g2854 ( 
.A(n_2088),
.B(n_79),
.Y(n_2854)
);

AOI22xp33_ASAP7_75t_L g2855 ( 
.A1(n_2150),
.A2(n_82),
.B1(n_80),
.B2(n_81),
.Y(n_2855)
);

NAND2xp5_ASAP7_75t_L g2856 ( 
.A(n_2053),
.B(n_81),
.Y(n_2856)
);

INVx2_ASAP7_75t_L g2857 ( 
.A(n_2172),
.Y(n_2857)
);

INVx3_ASAP7_75t_L g2858 ( 
.A(n_2060),
.Y(n_2858)
);

INVx2_ASAP7_75t_L g2859 ( 
.A(n_2172),
.Y(n_2859)
);

INVx2_ASAP7_75t_L g2860 ( 
.A(n_2172),
.Y(n_2860)
);

NAND2xp5_ASAP7_75t_SL g2861 ( 
.A(n_2088),
.B(n_82),
.Y(n_2861)
);

INVx1_ASAP7_75t_L g2862 ( 
.A(n_2178),
.Y(n_2862)
);

AND3x1_ASAP7_75t_L g2863 ( 
.A(n_2149),
.B(n_81),
.C(n_83),
.Y(n_2863)
);

INVx2_ASAP7_75t_L g2864 ( 
.A(n_2172),
.Y(n_2864)
);

BUFx6f_ASAP7_75t_L g2865 ( 
.A(n_2238),
.Y(n_2865)
);

NAND2xp5_ASAP7_75t_SL g2866 ( 
.A(n_2088),
.B(n_84),
.Y(n_2866)
);

AND2x6_ASAP7_75t_L g2867 ( 
.A(n_2060),
.B(n_83),
.Y(n_2867)
);

BUFx3_ASAP7_75t_L g2868 ( 
.A(n_2245),
.Y(n_2868)
);

NAND2xp5_ASAP7_75t_L g2869 ( 
.A(n_2053),
.B(n_84),
.Y(n_2869)
);

INVx2_ASAP7_75t_L g2870 ( 
.A(n_2172),
.Y(n_2870)
);

BUFx6f_ASAP7_75t_L g2871 ( 
.A(n_2238),
.Y(n_2871)
);

INVx2_ASAP7_75t_SL g2872 ( 
.A(n_2136),
.Y(n_2872)
);

INVx5_ASAP7_75t_L g2873 ( 
.A(n_2136),
.Y(n_2873)
);

INVx5_ASAP7_75t_L g2874 ( 
.A(n_2136),
.Y(n_2874)
);

INVx1_ASAP7_75t_L g2875 ( 
.A(n_2178),
.Y(n_2875)
);

HB1xp67_ASAP7_75t_L g2876 ( 
.A(n_2063),
.Y(n_2876)
);

OR2x2_ASAP7_75t_SL g2877 ( 
.A(n_2089),
.B(n_84),
.Y(n_2877)
);

INVxp67_ASAP7_75t_L g2878 ( 
.A(n_2063),
.Y(n_2878)
);

NOR2xp33_ASAP7_75t_L g2879 ( 
.A(n_2072),
.B(n_85),
.Y(n_2879)
);

AND2x4_ASAP7_75t_L g2880 ( 
.A(n_2060),
.B(n_85),
.Y(n_2880)
);

INVx1_ASAP7_75t_L g2881 ( 
.A(n_2178),
.Y(n_2881)
);

INVx2_ASAP7_75t_L g2882 ( 
.A(n_2172),
.Y(n_2882)
);

NAND2xp5_ASAP7_75t_L g2883 ( 
.A(n_2060),
.B(n_85),
.Y(n_2883)
);

AOI221xp5_ASAP7_75t_SL g2884 ( 
.A1(n_2125),
.A2(n_88),
.B1(n_86),
.B2(n_87),
.C(n_89),
.Y(n_2884)
);

INVx3_ASAP7_75t_L g2885 ( 
.A(n_2060),
.Y(n_2885)
);

INVx1_ASAP7_75t_L g2886 ( 
.A(n_2178),
.Y(n_2886)
);

NAND2xp5_ASAP7_75t_L g2887 ( 
.A(n_2060),
.B(n_87),
.Y(n_2887)
);

NAND2xp5_ASAP7_75t_L g2888 ( 
.A(n_2053),
.B(n_87),
.Y(n_2888)
);

BUFx3_ASAP7_75t_L g2889 ( 
.A(n_2245),
.Y(n_2889)
);

INVx1_ASAP7_75t_L g2890 ( 
.A(n_2178),
.Y(n_2890)
);

INVx2_ASAP7_75t_L g2891 ( 
.A(n_2172),
.Y(n_2891)
);

INVx1_ASAP7_75t_L g2892 ( 
.A(n_2178),
.Y(n_2892)
);

AND2x4_ASAP7_75t_L g2893 ( 
.A(n_2060),
.B(n_88),
.Y(n_2893)
);

AOI22xp33_ASAP7_75t_L g2894 ( 
.A1(n_2150),
.A2(n_91),
.B1(n_89),
.B2(n_90),
.Y(n_2894)
);

INVx3_ASAP7_75t_L g2895 ( 
.A(n_2060),
.Y(n_2895)
);

OR2x2_ASAP7_75t_L g2896 ( 
.A(n_2080),
.B(n_89),
.Y(n_2896)
);

AND2x6_ASAP7_75t_SL g2897 ( 
.A(n_2330),
.B(n_92),
.Y(n_2897)
);

NAND2xp5_ASAP7_75t_L g2898 ( 
.A(n_2060),
.B(n_91),
.Y(n_2898)
);

INVx1_ASAP7_75t_L g2899 ( 
.A(n_2178),
.Y(n_2899)
);

INVx2_ASAP7_75t_L g2900 ( 
.A(n_2172),
.Y(n_2900)
);

AND2x4_ASAP7_75t_L g2901 ( 
.A(n_2060),
.B(n_92),
.Y(n_2901)
);

A2O1A1Ixp33_ASAP7_75t_SL g2902 ( 
.A1(n_2159),
.A2(n_94),
.B(n_92),
.C(n_93),
.Y(n_2902)
);

INVx3_ASAP7_75t_L g2903 ( 
.A(n_2060),
.Y(n_2903)
);

NAND2xp33_ASAP7_75t_L g2904 ( 
.A(n_2060),
.B(n_94),
.Y(n_2904)
);

INVx1_ASAP7_75t_L g2905 ( 
.A(n_2178),
.Y(n_2905)
);

INVx1_ASAP7_75t_L g2906 ( 
.A(n_2428),
.Y(n_2906)
);

BUFx2_ASAP7_75t_L g2907 ( 
.A(n_2537),
.Y(n_2907)
);

NAND2xp5_ASAP7_75t_L g2908 ( 
.A(n_2402),
.B(n_2460),
.Y(n_2908)
);

AOI21xp5_ASAP7_75t_L g2909 ( 
.A1(n_2540),
.A2(n_93),
.B(n_95),
.Y(n_2909)
);

AOI22xp33_ASAP7_75t_L g2910 ( 
.A1(n_2474),
.A2(n_97),
.B1(n_95),
.B2(n_96),
.Y(n_2910)
);

OR2x2_ASAP7_75t_L g2911 ( 
.A(n_2825),
.B(n_2853),
.Y(n_2911)
);

NAND2xp5_ASAP7_75t_L g2912 ( 
.A(n_2402),
.B(n_95),
.Y(n_2912)
);

CKINVDCx5p33_ASAP7_75t_R g2913 ( 
.A(n_2852),
.Y(n_2913)
);

NAND2xp5_ASAP7_75t_SL g2914 ( 
.A(n_2427),
.B(n_341),
.Y(n_2914)
);

NAND2xp5_ASAP7_75t_L g2915 ( 
.A(n_2487),
.B(n_98),
.Y(n_2915)
);

AOI21xp5_ASAP7_75t_L g2916 ( 
.A1(n_2540),
.A2(n_98),
.B(n_99),
.Y(n_2916)
);

NAND2xp5_ASAP7_75t_SL g2917 ( 
.A(n_2854),
.B(n_341),
.Y(n_2917)
);

NAND2xp5_ASAP7_75t_L g2918 ( 
.A(n_2579),
.B(n_98),
.Y(n_2918)
);

INVx3_ASAP7_75t_L g2919 ( 
.A(n_2809),
.Y(n_2919)
);

OAI21xp33_ASAP7_75t_L g2920 ( 
.A1(n_2854),
.A2(n_99),
.B(n_100),
.Y(n_2920)
);

INVx1_ASAP7_75t_L g2921 ( 
.A(n_2430),
.Y(n_2921)
);

NOR2xp33_ASAP7_75t_L g2922 ( 
.A(n_2461),
.B(n_100),
.Y(n_2922)
);

AOI21xp5_ASAP7_75t_L g2923 ( 
.A1(n_2621),
.A2(n_100),
.B(n_101),
.Y(n_2923)
);

NOR2xp33_ASAP7_75t_L g2924 ( 
.A(n_2609),
.B(n_101),
.Y(n_2924)
);

NOR3xp33_ASAP7_75t_SL g2925 ( 
.A(n_2543),
.B(n_101),
.C(n_102),
.Y(n_2925)
);

AOI21xp5_ASAP7_75t_L g2926 ( 
.A1(n_2621),
.A2(n_102),
.B(n_103),
.Y(n_2926)
);

AOI21xp5_ASAP7_75t_L g2927 ( 
.A1(n_2445),
.A2(n_103),
.B(n_104),
.Y(n_2927)
);

NAND2xp5_ASAP7_75t_L g2928 ( 
.A(n_2778),
.B(n_104),
.Y(n_2928)
);

INVx1_ASAP7_75t_SL g2929 ( 
.A(n_2825),
.Y(n_2929)
);

AOI221x1_ASAP7_75t_L g2930 ( 
.A1(n_2792),
.A2(n_2844),
.B1(n_2713),
.B2(n_2703),
.C(n_2834),
.Y(n_2930)
);

NAND2xp5_ASAP7_75t_L g2931 ( 
.A(n_2602),
.B(n_104),
.Y(n_2931)
);

AO22x2_ASAP7_75t_L g2932 ( 
.A1(n_2781),
.A2(n_108),
.B1(n_106),
.B2(n_107),
.Y(n_2932)
);

OAI22xp5_ASAP7_75t_L g2933 ( 
.A1(n_2771),
.A2(n_108),
.B1(n_106),
.B2(n_107),
.Y(n_2933)
);

INVx3_ASAP7_75t_L g2934 ( 
.A(n_2809),
.Y(n_2934)
);

AO21x1_ASAP7_75t_L g2935 ( 
.A1(n_2904),
.A2(n_343),
.B(n_342),
.Y(n_2935)
);

BUFx2_ASAP7_75t_L g2936 ( 
.A(n_2413),
.Y(n_2936)
);

AOI21xp5_ASAP7_75t_L g2937 ( 
.A1(n_2749),
.A2(n_2554),
.B(n_2451),
.Y(n_2937)
);

NOR2xp33_ASAP7_75t_L g2938 ( 
.A(n_2614),
.B(n_106),
.Y(n_2938)
);

INVx1_ASAP7_75t_L g2939 ( 
.A(n_2433),
.Y(n_2939)
);

O2A1O1Ixp33_ASAP7_75t_L g2940 ( 
.A1(n_2902),
.A2(n_110),
.B(n_107),
.C(n_109),
.Y(n_2940)
);

NAND2xp33_ASAP7_75t_SL g2941 ( 
.A(n_2639),
.B(n_109),
.Y(n_2941)
);

NAND2xp5_ASAP7_75t_L g2942 ( 
.A(n_2608),
.B(n_109),
.Y(n_2942)
);

NAND2xp5_ASAP7_75t_SL g2943 ( 
.A(n_2497),
.B(n_344),
.Y(n_2943)
);

NOR2xp33_ASAP7_75t_L g2944 ( 
.A(n_2423),
.B(n_110),
.Y(n_2944)
);

AOI21xp5_ASAP7_75t_L g2945 ( 
.A1(n_2451),
.A2(n_110),
.B(n_111),
.Y(n_2945)
);

AOI21xp5_ASAP7_75t_L g2946 ( 
.A1(n_2715),
.A2(n_111),
.B(n_112),
.Y(n_2946)
);

AOI21xp5_ASAP7_75t_L g2947 ( 
.A1(n_2706),
.A2(n_112),
.B(n_113),
.Y(n_2947)
);

OAI22xp5_ASAP7_75t_L g2948 ( 
.A1(n_2771),
.A2(n_114),
.B1(n_112),
.B2(n_113),
.Y(n_2948)
);

INVx1_ASAP7_75t_L g2949 ( 
.A(n_2440),
.Y(n_2949)
);

INVx2_ASAP7_75t_L g2950 ( 
.A(n_2845),
.Y(n_2950)
);

BUFx3_ASAP7_75t_L g2951 ( 
.A(n_2809),
.Y(n_2951)
);

AOI22xp5_ASAP7_75t_L g2952 ( 
.A1(n_2647),
.A2(n_115),
.B1(n_113),
.B2(n_114),
.Y(n_2952)
);

AOI21xp5_ASAP7_75t_L g2953 ( 
.A1(n_2706),
.A2(n_114),
.B(n_115),
.Y(n_2953)
);

O2A1O1Ixp33_ASAP7_75t_L g2954 ( 
.A1(n_2722),
.A2(n_117),
.B(n_115),
.C(n_116),
.Y(n_2954)
);

OAI22xp5_ASAP7_75t_L g2955 ( 
.A1(n_2845),
.A2(n_118),
.B1(n_116),
.B2(n_117),
.Y(n_2955)
);

NAND3xp33_ASAP7_75t_L g2956 ( 
.A(n_2604),
.B(n_116),
.C(n_117),
.Y(n_2956)
);

AND2x2_ASAP7_75t_L g2957 ( 
.A(n_2796),
.B(n_118),
.Y(n_2957)
);

INVx3_ASAP7_75t_L g2958 ( 
.A(n_2873),
.Y(n_2958)
);

AOI21xp5_ASAP7_75t_L g2959 ( 
.A1(n_2453),
.A2(n_118),
.B(n_120),
.Y(n_2959)
);

NAND2xp5_ASAP7_75t_SL g2960 ( 
.A(n_2497),
.B(n_345),
.Y(n_2960)
);

BUFx2_ASAP7_75t_L g2961 ( 
.A(n_2808),
.Y(n_2961)
);

AOI33xp33_ASAP7_75t_L g2962 ( 
.A1(n_2448),
.A2(n_122),
.A3(n_124),
.B1(n_120),
.B2(n_121),
.B3(n_123),
.Y(n_2962)
);

INVx2_ASAP7_75t_L g2963 ( 
.A(n_2858),
.Y(n_2963)
);

INVx3_ASAP7_75t_L g2964 ( 
.A(n_2873),
.Y(n_2964)
);

NAND2xp5_ASAP7_75t_L g2965 ( 
.A(n_2657),
.B(n_120),
.Y(n_2965)
);

BUFx2_ASAP7_75t_L g2966 ( 
.A(n_2812),
.Y(n_2966)
);

AOI22xp5_ASAP7_75t_L g2967 ( 
.A1(n_2674),
.A2(n_123),
.B1(n_121),
.B2(n_122),
.Y(n_2967)
);

BUFx6f_ASAP7_75t_L g2968 ( 
.A(n_2406),
.Y(n_2968)
);

BUFx6f_ASAP7_75t_L g2969 ( 
.A(n_2406),
.Y(n_2969)
);

INVxp33_ASAP7_75t_SL g2970 ( 
.A(n_2623),
.Y(n_2970)
);

NAND2xp5_ASAP7_75t_L g2971 ( 
.A(n_2665),
.B(n_121),
.Y(n_2971)
);

NAND2xp5_ASAP7_75t_SL g2972 ( 
.A(n_2666),
.B(n_2556),
.Y(n_2972)
);

NAND2xp5_ASAP7_75t_L g2973 ( 
.A(n_2683),
.B(n_122),
.Y(n_2973)
);

NOR2xp33_ASAP7_75t_L g2974 ( 
.A(n_2659),
.B(n_124),
.Y(n_2974)
);

NAND2xp5_ASAP7_75t_L g2975 ( 
.A(n_2685),
.B(n_124),
.Y(n_2975)
);

AOI22xp33_ASAP7_75t_L g2976 ( 
.A1(n_2834),
.A2(n_127),
.B1(n_125),
.B2(n_126),
.Y(n_2976)
);

NAND2xp5_ASAP7_75t_SL g2977 ( 
.A(n_2858),
.B(n_346),
.Y(n_2977)
);

CKINVDCx5p33_ASAP7_75t_R g2978 ( 
.A(n_2767),
.Y(n_2978)
);

NOR2xp33_ASAP7_75t_L g2979 ( 
.A(n_2631),
.B(n_126),
.Y(n_2979)
);

NOR2xp33_ASAP7_75t_R g2980 ( 
.A(n_2873),
.B(n_127),
.Y(n_2980)
);

NAND3xp33_ASAP7_75t_SL g2981 ( 
.A(n_2519),
.B(n_128),
.C(n_129),
.Y(n_2981)
);

AOI21xp5_ASAP7_75t_L g2982 ( 
.A1(n_2708),
.A2(n_128),
.B(n_129),
.Y(n_2982)
);

NOR2xp33_ASAP7_75t_SL g2983 ( 
.A(n_2401),
.B(n_128),
.Y(n_2983)
);

AOI21xp5_ASAP7_75t_L g2984 ( 
.A1(n_2708),
.A2(n_129),
.B(n_130),
.Y(n_2984)
);

BUFx6f_ASAP7_75t_L g2985 ( 
.A(n_2406),
.Y(n_2985)
);

NAND2xp5_ASAP7_75t_SL g2986 ( 
.A(n_2885),
.B(n_347),
.Y(n_2986)
);

INVx1_ASAP7_75t_L g2987 ( 
.A(n_2444),
.Y(n_2987)
);

O2A1O1Ixp33_ASAP7_75t_L g2988 ( 
.A1(n_2725),
.A2(n_2447),
.B(n_2619),
.C(n_2617),
.Y(n_2988)
);

A2O1A1Ixp33_ASAP7_75t_L g2989 ( 
.A1(n_2649),
.A2(n_133),
.B(n_130),
.C(n_132),
.Y(n_2989)
);

AOI22xp33_ASAP7_75t_L g2990 ( 
.A1(n_2707),
.A2(n_134),
.B1(n_132),
.B2(n_133),
.Y(n_2990)
);

NOR2xp33_ASAP7_75t_L g2991 ( 
.A(n_2424),
.B(n_132),
.Y(n_2991)
);

OAI22xp5_ASAP7_75t_L g2992 ( 
.A1(n_2885),
.A2(n_2903),
.B1(n_2895),
.B2(n_2781),
.Y(n_2992)
);

BUFx2_ASAP7_75t_L g2993 ( 
.A(n_2851),
.Y(n_2993)
);

AOI21xp5_ASAP7_75t_L g2994 ( 
.A1(n_2662),
.A2(n_133),
.B(n_134),
.Y(n_2994)
);

O2A1O1Ixp33_ASAP7_75t_L g2995 ( 
.A1(n_2738),
.A2(n_136),
.B(n_134),
.C(n_135),
.Y(n_2995)
);

A2O1A1Ixp33_ASAP7_75t_L g2996 ( 
.A1(n_2649),
.A2(n_137),
.B(n_135),
.C(n_136),
.Y(n_2996)
);

INVx2_ASAP7_75t_L g2997 ( 
.A(n_2895),
.Y(n_2997)
);

INVx2_ASAP7_75t_L g2998 ( 
.A(n_2903),
.Y(n_2998)
);

NOR2xp33_ASAP7_75t_L g2999 ( 
.A(n_2415),
.B(n_135),
.Y(n_2999)
);

AOI21xp5_ASAP7_75t_L g3000 ( 
.A1(n_2692),
.A2(n_2495),
.B(n_2616),
.Y(n_3000)
);

OR2x6_ASAP7_75t_L g3001 ( 
.A(n_2401),
.B(n_2412),
.Y(n_3001)
);

INVx1_ASAP7_75t_L g3002 ( 
.A(n_2398),
.Y(n_3002)
);

OAI22xp5_ASAP7_75t_L g3003 ( 
.A1(n_2787),
.A2(n_138),
.B1(n_136),
.B2(n_137),
.Y(n_3003)
);

OAI22xp5_ASAP7_75t_L g3004 ( 
.A1(n_2787),
.A2(n_140),
.B1(n_138),
.B2(n_139),
.Y(n_3004)
);

BUFx6f_ASAP7_75t_L g3005 ( 
.A(n_2628),
.Y(n_3005)
);

O2A1O1Ixp33_ASAP7_75t_L g3006 ( 
.A1(n_2687),
.A2(n_140),
.B(n_138),
.C(n_139),
.Y(n_3006)
);

AOI22xp33_ASAP7_75t_L g3007 ( 
.A1(n_2707),
.A2(n_143),
.B1(n_141),
.B2(n_142),
.Y(n_3007)
);

CKINVDCx5p33_ASAP7_75t_R g3008 ( 
.A(n_2843),
.Y(n_3008)
);

CKINVDCx10_ASAP7_75t_R g3009 ( 
.A(n_2561),
.Y(n_3009)
);

NAND2xp5_ASAP7_75t_SL g3010 ( 
.A(n_2541),
.B(n_347),
.Y(n_3010)
);

INVx2_ASAP7_75t_L g3011 ( 
.A(n_2417),
.Y(n_3011)
);

BUFx6f_ASAP7_75t_L g3012 ( 
.A(n_2628),
.Y(n_3012)
);

NOR2xp33_ASAP7_75t_L g3013 ( 
.A(n_2415),
.B(n_141),
.Y(n_3013)
);

O2A1O1Ixp33_ASAP7_75t_L g3014 ( 
.A1(n_2605),
.A2(n_143),
.B(n_141),
.C(n_142),
.Y(n_3014)
);

BUFx6f_ASAP7_75t_SL g3015 ( 
.A(n_2446),
.Y(n_3015)
);

AND2x2_ASAP7_75t_L g3016 ( 
.A(n_2442),
.B(n_142),
.Y(n_3016)
);

HB1xp67_ASAP7_75t_L g3017 ( 
.A(n_2790),
.Y(n_3017)
);

NOR2xp33_ASAP7_75t_L g3018 ( 
.A(n_2437),
.B(n_143),
.Y(n_3018)
);

BUFx6f_ASAP7_75t_L g3019 ( 
.A(n_2628),
.Y(n_3019)
);

O2A1O1Ixp33_ASAP7_75t_L g3020 ( 
.A1(n_2682),
.A2(n_146),
.B(n_144),
.C(n_145),
.Y(n_3020)
);

INVx3_ASAP7_75t_L g3021 ( 
.A(n_2874),
.Y(n_3021)
);

INVx2_ASAP7_75t_L g3022 ( 
.A(n_2420),
.Y(n_3022)
);

AOI21xp5_ASAP7_75t_L g3023 ( 
.A1(n_2616),
.A2(n_144),
.B(n_145),
.Y(n_3023)
);

HB1xp67_ASAP7_75t_L g3024 ( 
.A(n_2876),
.Y(n_3024)
);

O2A1O1Ixp33_ASAP7_75t_L g3025 ( 
.A1(n_2752),
.A2(n_148),
.B(n_146),
.C(n_147),
.Y(n_3025)
);

NOR2xp33_ASAP7_75t_L g3026 ( 
.A(n_2719),
.B(n_2588),
.Y(n_3026)
);

AOI22xp33_ASAP7_75t_L g3027 ( 
.A1(n_2707),
.A2(n_148),
.B1(n_146),
.B2(n_147),
.Y(n_3027)
);

NAND2xp5_ASAP7_75t_L g3028 ( 
.A(n_2690),
.B(n_147),
.Y(n_3028)
);

AOI21xp5_ASAP7_75t_L g3029 ( 
.A1(n_2673),
.A2(n_2597),
.B(n_2770),
.Y(n_3029)
);

NAND2xp5_ASAP7_75t_SL g3030 ( 
.A(n_2521),
.B(n_348),
.Y(n_3030)
);

AND2x2_ASAP7_75t_L g3031 ( 
.A(n_2573),
.B(n_149),
.Y(n_3031)
);

AND2x2_ASAP7_75t_L g3032 ( 
.A(n_2573),
.B(n_149),
.Y(n_3032)
);

A2O1A1Ixp33_ASAP7_75t_L g3033 ( 
.A1(n_2689),
.A2(n_152),
.B(n_150),
.C(n_151),
.Y(n_3033)
);

NAND2xp33_ASAP7_75t_R g3034 ( 
.A(n_2513),
.B(n_150),
.Y(n_3034)
);

NAND2xp5_ASAP7_75t_SL g3035 ( 
.A(n_2806),
.B(n_348),
.Y(n_3035)
);

AOI21xp5_ASAP7_75t_L g3036 ( 
.A1(n_2774),
.A2(n_150),
.B(n_151),
.Y(n_3036)
);

NAND2xp5_ASAP7_75t_L g3037 ( 
.A(n_2694),
.B(n_151),
.Y(n_3037)
);

OAI22xp5_ASAP7_75t_L g3038 ( 
.A1(n_2806),
.A2(n_154),
.B1(n_152),
.B2(n_153),
.Y(n_3038)
);

NAND2xp5_ASAP7_75t_L g3039 ( 
.A(n_2695),
.B(n_152),
.Y(n_3039)
);

NAND2xp5_ASAP7_75t_L g3040 ( 
.A(n_2697),
.B(n_154),
.Y(n_3040)
);

INVx2_ASAP7_75t_L g3041 ( 
.A(n_2452),
.Y(n_3041)
);

OAI22xp5_ASAP7_75t_L g3042 ( 
.A1(n_2839),
.A2(n_157),
.B1(n_155),
.B2(n_156),
.Y(n_3042)
);

INVxp67_ASAP7_75t_L g3043 ( 
.A(n_2623),
.Y(n_3043)
);

NOR3xp33_ASAP7_75t_L g3044 ( 
.A(n_2794),
.B(n_156),
.C(n_157),
.Y(n_3044)
);

INVx4_ASAP7_75t_L g3045 ( 
.A(n_2874),
.Y(n_3045)
);

AOI21xp5_ASAP7_75t_L g3046 ( 
.A1(n_2780),
.A2(n_156),
.B(n_157),
.Y(n_3046)
);

INVx2_ASAP7_75t_L g3047 ( 
.A(n_2462),
.Y(n_3047)
);

INVxp67_ASAP7_75t_SL g3048 ( 
.A(n_2839),
.Y(n_3048)
);

NAND2xp5_ASAP7_75t_L g3049 ( 
.A(n_2699),
.B(n_158),
.Y(n_3049)
);

NOR2xp33_ASAP7_75t_L g3050 ( 
.A(n_2598),
.B(n_158),
.Y(n_3050)
);

INVx1_ASAP7_75t_L g3051 ( 
.A(n_2407),
.Y(n_3051)
);

AOI21xp5_ASAP7_75t_L g3052 ( 
.A1(n_2795),
.A2(n_158),
.B(n_159),
.Y(n_3052)
);

OAI22xp5_ASAP7_75t_SL g3053 ( 
.A1(n_2877),
.A2(n_163),
.B1(n_159),
.B2(n_160),
.Y(n_3053)
);

INVxp33_ASAP7_75t_SL g3054 ( 
.A(n_2775),
.Y(n_3054)
);

AND2x2_ASAP7_75t_L g3055 ( 
.A(n_2896),
.B(n_163),
.Y(n_3055)
);

INVxp67_ASAP7_75t_L g3056 ( 
.A(n_2438),
.Y(n_3056)
);

AOI21xp5_ASAP7_75t_L g3057 ( 
.A1(n_2801),
.A2(n_163),
.B(n_164),
.Y(n_3057)
);

OAI321xp33_ASAP7_75t_L g3058 ( 
.A1(n_2835),
.A2(n_2792),
.A3(n_2829),
.B1(n_2784),
.B2(n_2773),
.C(n_2409),
.Y(n_3058)
);

AND2x4_ASAP7_75t_L g3059 ( 
.A(n_2874),
.B(n_164),
.Y(n_3059)
);

INVx3_ASAP7_75t_L g3060 ( 
.A(n_2615),
.Y(n_3060)
);

NAND2xp33_ASAP7_75t_SL g3061 ( 
.A(n_2880),
.B(n_165),
.Y(n_3061)
);

NAND2xp5_ASAP7_75t_SL g3062 ( 
.A(n_2880),
.B(n_349),
.Y(n_3062)
);

INVx1_ASAP7_75t_L g3063 ( 
.A(n_2421),
.Y(n_3063)
);

OAI21xp5_ASAP7_75t_L g3064 ( 
.A1(n_2410),
.A2(n_165),
.B(n_166),
.Y(n_3064)
);

A2O1A1Ixp33_ASAP7_75t_L g3065 ( 
.A1(n_2689),
.A2(n_167),
.B(n_165),
.C(n_166),
.Y(n_3065)
);

NAND2xp5_ASAP7_75t_L g3066 ( 
.A(n_2439),
.B(n_166),
.Y(n_3066)
);

INVx2_ASAP7_75t_L g3067 ( 
.A(n_2463),
.Y(n_3067)
);

INVx1_ASAP7_75t_L g3068 ( 
.A(n_2422),
.Y(n_3068)
);

NAND2xp5_ASAP7_75t_SL g3069 ( 
.A(n_2893),
.B(n_350),
.Y(n_3069)
);

A2O1A1Ixp33_ASAP7_75t_L g3070 ( 
.A1(n_2723),
.A2(n_169),
.B(n_167),
.C(n_168),
.Y(n_3070)
);

A2O1A1Ixp33_ASAP7_75t_L g3071 ( 
.A1(n_2677),
.A2(n_2732),
.B(n_2736),
.C(n_2735),
.Y(n_3071)
);

AOI21xp5_ASAP7_75t_L g3072 ( 
.A1(n_2805),
.A2(n_167),
.B(n_168),
.Y(n_3072)
);

INVx1_ASAP7_75t_L g3073 ( 
.A(n_2429),
.Y(n_3073)
);

INVx4_ASAP7_75t_L g3074 ( 
.A(n_2868),
.Y(n_3074)
);

CKINVDCx14_ASAP7_75t_R g3075 ( 
.A(n_2793),
.Y(n_3075)
);

BUFx2_ASAP7_75t_L g3076 ( 
.A(n_2867),
.Y(n_3076)
);

CKINVDCx10_ASAP7_75t_R g3077 ( 
.A(n_2561),
.Y(n_3077)
);

AOI21xp5_ASAP7_75t_L g3078 ( 
.A1(n_2807),
.A2(n_168),
.B(n_169),
.Y(n_3078)
);

AOI22xp5_ASAP7_75t_L g3079 ( 
.A1(n_2893),
.A2(n_171),
.B1(n_169),
.B2(n_170),
.Y(n_3079)
);

NOR2xp33_ASAP7_75t_L g3080 ( 
.A(n_2817),
.B(n_170),
.Y(n_3080)
);

NAND2xp5_ASAP7_75t_SL g3081 ( 
.A(n_2901),
.B(n_350),
.Y(n_3081)
);

AOI21xp5_ASAP7_75t_L g3082 ( 
.A1(n_2816),
.A2(n_170),
.B(n_172),
.Y(n_3082)
);

NAND2xp5_ASAP7_75t_L g3083 ( 
.A(n_2439),
.B(n_172),
.Y(n_3083)
);

BUFx12f_ASAP7_75t_L g3084 ( 
.A(n_2843),
.Y(n_3084)
);

AOI22xp33_ASAP7_75t_SL g3085 ( 
.A1(n_2867),
.A2(n_174),
.B1(n_172),
.B2(n_173),
.Y(n_3085)
);

NAND2xp5_ASAP7_75t_L g3086 ( 
.A(n_2431),
.B(n_173),
.Y(n_3086)
);

AND2x6_ASAP7_75t_SL g3087 ( 
.A(n_2465),
.B(n_173),
.Y(n_3087)
);

NAND2xp5_ASAP7_75t_SL g3088 ( 
.A(n_2901),
.B(n_351),
.Y(n_3088)
);

A2O1A1Ixp33_ASAP7_75t_L g3089 ( 
.A1(n_2717),
.A2(n_176),
.B(n_174),
.C(n_175),
.Y(n_3089)
);

OAI22xp5_ASAP7_75t_L g3090 ( 
.A1(n_2524),
.A2(n_176),
.B1(n_174),
.B2(n_175),
.Y(n_3090)
);

A2O1A1Ixp33_ASAP7_75t_SL g3091 ( 
.A1(n_2743),
.A2(n_177),
.B(n_175),
.C(n_176),
.Y(n_3091)
);

CKINVDCx20_ASAP7_75t_R g3092 ( 
.A(n_2889),
.Y(n_3092)
);

NAND2xp5_ASAP7_75t_L g3093 ( 
.A(n_2785),
.B(n_177),
.Y(n_3093)
);

NAND2xp5_ASAP7_75t_L g3094 ( 
.A(n_2786),
.B(n_177),
.Y(n_3094)
);

NAND2xp5_ASAP7_75t_L g3095 ( 
.A(n_2799),
.B(n_178),
.Y(n_3095)
);

OAI21x1_ASAP7_75t_L g3096 ( 
.A1(n_2435),
.A2(n_178),
.B(n_179),
.Y(n_3096)
);

BUFx2_ASAP7_75t_L g3097 ( 
.A(n_2867),
.Y(n_3097)
);

INVx1_ASAP7_75t_L g3098 ( 
.A(n_2803),
.Y(n_3098)
);

NAND2xp5_ASAP7_75t_L g3099 ( 
.A(n_2810),
.B(n_179),
.Y(n_3099)
);

O2A1O1Ixp33_ASAP7_75t_L g3100 ( 
.A1(n_2553),
.A2(n_181),
.B(n_179),
.C(n_180),
.Y(n_3100)
);

A2O1A1Ixp33_ASAP7_75t_L g3101 ( 
.A1(n_2717),
.A2(n_182),
.B(n_180),
.C(n_181),
.Y(n_3101)
);

NAND2xp33_ASAP7_75t_R g3102 ( 
.A(n_2837),
.B(n_180),
.Y(n_3102)
);

INVx1_ASAP7_75t_L g3103 ( 
.A(n_2819),
.Y(n_3103)
);

NAND2xp5_ASAP7_75t_L g3104 ( 
.A(n_2832),
.B(n_181),
.Y(n_3104)
);

NAND2xp5_ASAP7_75t_L g3105 ( 
.A(n_2850),
.B(n_182),
.Y(n_3105)
);

INVx1_ASAP7_75t_SL g3106 ( 
.A(n_2469),
.Y(n_3106)
);

AOI21xp5_ASAP7_75t_L g3107 ( 
.A1(n_2820),
.A2(n_182),
.B(n_183),
.Y(n_3107)
);

AOI21xp5_ASAP7_75t_L g3108 ( 
.A1(n_2821),
.A2(n_183),
.B(n_184),
.Y(n_3108)
);

OAI22xp5_ASAP7_75t_L g3109 ( 
.A1(n_2524),
.A2(n_187),
.B1(n_184),
.B2(n_185),
.Y(n_3109)
);

OA21x2_ASAP7_75t_L g3110 ( 
.A1(n_2669),
.A2(n_2761),
.B(n_2750),
.Y(n_3110)
);

NAND2xp5_ASAP7_75t_L g3111 ( 
.A(n_2862),
.B(n_184),
.Y(n_3111)
);

INVx5_ASAP7_75t_L g3112 ( 
.A(n_2867),
.Y(n_3112)
);

INVx1_ASAP7_75t_L g3113 ( 
.A(n_2875),
.Y(n_3113)
);

NOR2xp33_ASAP7_75t_L g3114 ( 
.A(n_2878),
.B(n_185),
.Y(n_3114)
);

INVx1_ASAP7_75t_L g3115 ( 
.A(n_2881),
.Y(n_3115)
);

INVx2_ASAP7_75t_L g3116 ( 
.A(n_2471),
.Y(n_3116)
);

OAI22xp5_ASAP7_75t_L g3117 ( 
.A1(n_2534),
.A2(n_189),
.B1(n_187),
.B2(n_188),
.Y(n_3117)
);

OR2x2_ASAP7_75t_L g3118 ( 
.A(n_2564),
.B(n_188),
.Y(n_3118)
);

INVx2_ASAP7_75t_L g3119 ( 
.A(n_2886),
.Y(n_3119)
);

AOI22xp5_ASAP7_75t_L g3120 ( 
.A1(n_2641),
.A2(n_191),
.B1(n_189),
.B2(n_190),
.Y(n_3120)
);

INVx1_ASAP7_75t_L g3121 ( 
.A(n_2890),
.Y(n_3121)
);

AOI22xp33_ASAP7_75t_L g3122 ( 
.A1(n_2707),
.A2(n_193),
.B1(n_190),
.B2(n_191),
.Y(n_3122)
);

AOI21xp5_ASAP7_75t_L g3123 ( 
.A1(n_2824),
.A2(n_190),
.B(n_191),
.Y(n_3123)
);

INVx6_ASAP7_75t_L g3124 ( 
.A(n_2478),
.Y(n_3124)
);

AOI22xp5_ASAP7_75t_L g3125 ( 
.A1(n_2747),
.A2(n_195),
.B1(n_193),
.B2(n_194),
.Y(n_3125)
);

NOR3xp33_ASAP7_75t_SL g3126 ( 
.A(n_2838),
.B(n_193),
.C(n_194),
.Y(n_3126)
);

NAND2xp5_ASAP7_75t_L g3127 ( 
.A(n_2892),
.B(n_194),
.Y(n_3127)
);

O2A1O1Ixp33_ASAP7_75t_SL g3128 ( 
.A1(n_2484),
.A2(n_197),
.B(n_195),
.C(n_196),
.Y(n_3128)
);

INVx1_ASAP7_75t_L g3129 ( 
.A(n_2899),
.Y(n_3129)
);

INVx4_ASAP7_75t_L g3130 ( 
.A(n_2478),
.Y(n_3130)
);

BUFx6f_ASAP7_75t_L g3131 ( 
.A(n_2651),
.Y(n_3131)
);

INVx2_ASAP7_75t_L g3132 ( 
.A(n_2905),
.Y(n_3132)
);

INVx1_ASAP7_75t_L g3133 ( 
.A(n_2459),
.Y(n_3133)
);

AOI21xp5_ASAP7_75t_L g3134 ( 
.A1(n_2826),
.A2(n_195),
.B(n_196),
.Y(n_3134)
);

O2A1O1Ixp33_ASAP7_75t_L g3135 ( 
.A1(n_2568),
.A2(n_199),
.B(n_197),
.C(n_198),
.Y(n_3135)
);

NAND2xp5_ASAP7_75t_SL g3136 ( 
.A(n_2606),
.B(n_351),
.Y(n_3136)
);

O2A1O1Ixp33_ASAP7_75t_L g3137 ( 
.A1(n_2578),
.A2(n_199),
.B(n_197),
.C(n_198),
.Y(n_3137)
);

INVx2_ASAP7_75t_L g3138 ( 
.A(n_2480),
.Y(n_3138)
);

INVx3_ASAP7_75t_L g3139 ( 
.A(n_2615),
.Y(n_3139)
);

NAND2xp5_ASAP7_75t_L g3140 ( 
.A(n_2517),
.B(n_198),
.Y(n_3140)
);

INVx1_ASAP7_75t_L g3141 ( 
.A(n_2464),
.Y(n_3141)
);

NAND2xp5_ASAP7_75t_L g3142 ( 
.A(n_2548),
.B(n_199),
.Y(n_3142)
);

AOI21xp5_ASAP7_75t_L g3143 ( 
.A1(n_2827),
.A2(n_200),
.B(n_201),
.Y(n_3143)
);

BUFx4f_ASAP7_75t_L g3144 ( 
.A(n_2492),
.Y(n_3144)
);

INVx6_ASAP7_75t_L g3145 ( 
.A(n_2478),
.Y(n_3145)
);

NOR2xp33_ASAP7_75t_L g3146 ( 
.A(n_2754),
.B(n_200),
.Y(n_3146)
);

NOR2xp67_ASAP7_75t_L g3147 ( 
.A(n_2520),
.B(n_201),
.Y(n_3147)
);

AND2x4_ASAP7_75t_L g3148 ( 
.A(n_2721),
.B(n_200),
.Y(n_3148)
);

BUFx3_ASAP7_75t_L g3149 ( 
.A(n_2418),
.Y(n_3149)
);

BUFx6f_ASAP7_75t_L g3150 ( 
.A(n_2651),
.Y(n_3150)
);

AOI21xp5_ASAP7_75t_L g3151 ( 
.A1(n_2828),
.A2(n_202),
.B(n_203),
.Y(n_3151)
);

O2A1O1Ixp33_ASAP7_75t_L g3152 ( 
.A1(n_2587),
.A2(n_205),
.B(n_202),
.C(n_203),
.Y(n_3152)
);

OAI22xp5_ASAP7_75t_L g3153 ( 
.A1(n_2534),
.A2(n_207),
.B1(n_202),
.B2(n_206),
.Y(n_3153)
);

INVx2_ASAP7_75t_SL g3154 ( 
.A(n_2397),
.Y(n_3154)
);

NAND2xp5_ASAP7_75t_L g3155 ( 
.A(n_2562),
.B(n_206),
.Y(n_3155)
);

INVx2_ASAP7_75t_L g3156 ( 
.A(n_2482),
.Y(n_3156)
);

AOI21xp5_ASAP7_75t_L g3157 ( 
.A1(n_2831),
.A2(n_207),
.B(n_208),
.Y(n_3157)
);

INVx3_ASAP7_75t_L g3158 ( 
.A(n_2615),
.Y(n_3158)
);

INVxp67_ASAP7_75t_L g3159 ( 
.A(n_2768),
.Y(n_3159)
);

INVx1_ASAP7_75t_L g3160 ( 
.A(n_2468),
.Y(n_3160)
);

AOI21xp5_ASAP7_75t_L g3161 ( 
.A1(n_2856),
.A2(n_208),
.B(n_209),
.Y(n_3161)
);

NAND2xp5_ASAP7_75t_L g3162 ( 
.A(n_2491),
.B(n_208),
.Y(n_3162)
);

NOR2xp33_ASAP7_75t_R g3163 ( 
.A(n_2426),
.B(n_209),
.Y(n_3163)
);

INVx2_ASAP7_75t_L g3164 ( 
.A(n_2500),
.Y(n_3164)
);

A2O1A1Ixp33_ASAP7_75t_L g3165 ( 
.A1(n_2737),
.A2(n_212),
.B(n_209),
.C(n_211),
.Y(n_3165)
);

INVx1_ASAP7_75t_SL g3166 ( 
.A(n_2663),
.Y(n_3166)
);

OR2x2_ASAP7_75t_L g3167 ( 
.A(n_2399),
.B(n_211),
.Y(n_3167)
);

AOI21xp5_ASAP7_75t_L g3168 ( 
.A1(n_2869),
.A2(n_211),
.B(n_212),
.Y(n_3168)
);

A2O1A1Ixp33_ASAP7_75t_L g3169 ( 
.A1(n_2741),
.A2(n_214),
.B(n_212),
.C(n_213),
.Y(n_3169)
);

NOR2xp33_ASAP7_75t_L g3170 ( 
.A(n_2457),
.B(n_214),
.Y(n_3170)
);

NOR2xp33_ASAP7_75t_SL g3171 ( 
.A(n_2515),
.B(n_214),
.Y(n_3171)
);

OAI22xp5_ASAP7_75t_L g3172 ( 
.A1(n_2782),
.A2(n_2898),
.B1(n_2789),
.B2(n_2811),
.Y(n_3172)
);

INVx2_ASAP7_75t_L g3173 ( 
.A(n_2505),
.Y(n_3173)
);

HB1xp67_ASAP7_75t_L g3174 ( 
.A(n_2656),
.Y(n_3174)
);

AOI21xp5_ASAP7_75t_L g3175 ( 
.A1(n_2888),
.A2(n_215),
.B(n_216),
.Y(n_3175)
);

OAI21xp33_ASAP7_75t_L g3176 ( 
.A1(n_2626),
.A2(n_215),
.B(n_216),
.Y(n_3176)
);

AOI21xp5_ASAP7_75t_L g3177 ( 
.A1(n_2414),
.A2(n_216),
.B(n_217),
.Y(n_3177)
);

AND2x2_ASAP7_75t_L g3178 ( 
.A(n_2655),
.B(n_217),
.Y(n_3178)
);

AOI22xp33_ASAP7_75t_L g3179 ( 
.A1(n_2672),
.A2(n_219),
.B1(n_217),
.B2(n_218),
.Y(n_3179)
);

NAND2xp5_ASAP7_75t_L g3180 ( 
.A(n_2494),
.B(n_2498),
.Y(n_3180)
);

NOR2xp33_ASAP7_75t_L g3181 ( 
.A(n_2710),
.B(n_218),
.Y(n_3181)
);

A2O1A1Ixp33_ASAP7_75t_L g3182 ( 
.A1(n_2742),
.A2(n_220),
.B(n_218),
.C(n_219),
.Y(n_3182)
);

O2A1O1Ixp33_ASAP7_75t_SL g3183 ( 
.A1(n_2583),
.A2(n_222),
.B(n_220),
.C(n_221),
.Y(n_3183)
);

NOR3xp33_ASAP7_75t_SL g3184 ( 
.A(n_2693),
.B(n_221),
.C(n_222),
.Y(n_3184)
);

AOI22xp5_ASAP7_75t_L g3185 ( 
.A1(n_2522),
.A2(n_223),
.B1(n_221),
.B2(n_222),
.Y(n_3185)
);

AOI21xp5_ASAP7_75t_L g3186 ( 
.A1(n_2637),
.A2(n_223),
.B(n_224),
.Y(n_3186)
);

BUFx2_ASAP7_75t_L g3187 ( 
.A(n_2426),
.Y(n_3187)
);

OAI22x1_ASAP7_75t_L g3188 ( 
.A1(n_2847),
.A2(n_225),
.B1(n_223),
.B2(n_224),
.Y(n_3188)
);

INVx1_ASAP7_75t_L g3189 ( 
.A(n_2475),
.Y(n_3189)
);

NAND2xp5_ASAP7_75t_SL g3190 ( 
.A(n_2606),
.B(n_352),
.Y(n_3190)
);

NOR2xp33_ASAP7_75t_L g3191 ( 
.A(n_2710),
.B(n_224),
.Y(n_3191)
);

AO32x2_ASAP7_75t_L g3192 ( 
.A1(n_2753),
.A2(n_227),
.A3(n_225),
.B1(n_226),
.B2(n_228),
.Y(n_3192)
);

BUFx6f_ASAP7_75t_L g3193 ( 
.A(n_2651),
.Y(n_3193)
);

BUFx3_ASAP7_75t_L g3194 ( 
.A(n_2408),
.Y(n_3194)
);

NAND2xp5_ASAP7_75t_L g3195 ( 
.A(n_2499),
.B(n_226),
.Y(n_3195)
);

OAI22xp5_ASAP7_75t_L g3196 ( 
.A1(n_2782),
.A2(n_228),
.B1(n_226),
.B2(n_227),
.Y(n_3196)
);

NOR2xp33_ASAP7_75t_L g3197 ( 
.A(n_2644),
.B(n_228),
.Y(n_3197)
);

NAND2xp5_ASAP7_75t_L g3198 ( 
.A(n_2504),
.B(n_229),
.Y(n_3198)
);

AOI22xp33_ASAP7_75t_L g3199 ( 
.A1(n_2672),
.A2(n_231),
.B1(n_229),
.B2(n_230),
.Y(n_3199)
);

BUFx3_ASAP7_75t_L g3200 ( 
.A(n_2872),
.Y(n_3200)
);

AOI21xp33_ASAP7_75t_L g3201 ( 
.A1(n_2640),
.A2(n_229),
.B(n_230),
.Y(n_3201)
);

AOI21xp5_ASAP7_75t_L g3202 ( 
.A1(n_2642),
.A2(n_232),
.B(n_233),
.Y(n_3202)
);

NAND2x1p5_ASAP7_75t_L g3203 ( 
.A(n_2436),
.B(n_232),
.Y(n_3203)
);

OR2x2_ASAP7_75t_L g3204 ( 
.A(n_2432),
.B(n_232),
.Y(n_3204)
);

INVx1_ASAP7_75t_L g3205 ( 
.A(n_2557),
.Y(n_3205)
);

OAI21xp33_ASAP7_75t_SL g3206 ( 
.A1(n_2755),
.A2(n_235),
.B(n_234),
.Y(n_3206)
);

AOI21xp5_ASAP7_75t_L g3207 ( 
.A1(n_2646),
.A2(n_233),
.B(n_234),
.Y(n_3207)
);

NAND2xp5_ASAP7_75t_L g3208 ( 
.A(n_2508),
.B(n_233),
.Y(n_3208)
);

A2O1A1Ixp33_ASAP7_75t_L g3209 ( 
.A1(n_2670),
.A2(n_236),
.B(n_234),
.C(n_235),
.Y(n_3209)
);

INVx1_ASAP7_75t_L g3210 ( 
.A(n_2559),
.Y(n_3210)
);

OA21x2_ASAP7_75t_L g3211 ( 
.A1(n_2670),
.A2(n_236),
.B(n_237),
.Y(n_3211)
);

OR2x2_ASAP7_75t_L g3212 ( 
.A(n_2432),
.B(n_236),
.Y(n_3212)
);

INVx2_ASAP7_75t_SL g3213 ( 
.A(n_2436),
.Y(n_3213)
);

NOR2xp33_ASAP7_75t_L g3214 ( 
.A(n_2561),
.B(n_237),
.Y(n_3214)
);

AND2x4_ASAP7_75t_L g3215 ( 
.A(n_2727),
.B(n_237),
.Y(n_3215)
);

OAI21xp5_ASAP7_75t_L g3216 ( 
.A1(n_2601),
.A2(n_238),
.B(n_239),
.Y(n_3216)
);

OR2x6_ASAP7_75t_SL g3217 ( 
.A(n_2668),
.B(n_238),
.Y(n_3217)
);

NOR2xp33_ASAP7_75t_L g3218 ( 
.A(n_2734),
.B(n_238),
.Y(n_3218)
);

BUFx3_ASAP7_75t_L g3219 ( 
.A(n_2503),
.Y(n_3219)
);

NAND2xp5_ASAP7_75t_SL g3220 ( 
.A(n_2643),
.B(n_353),
.Y(n_3220)
);

AOI33xp33_ASAP7_75t_L g3221 ( 
.A1(n_2411),
.A2(n_241),
.A3(n_243),
.B1(n_239),
.B2(n_240),
.B3(n_242),
.Y(n_3221)
);

NAND2xp5_ASAP7_75t_L g3222 ( 
.A(n_2613),
.B(n_239),
.Y(n_3222)
);

AND3x4_ASAP7_75t_L g3223 ( 
.A(n_2823),
.B(n_2836),
.C(n_2686),
.Y(n_3223)
);

NOR2xp33_ASAP7_75t_L g3224 ( 
.A(n_2580),
.B(n_2584),
.Y(n_3224)
);

O2A1O1Ixp33_ASAP7_75t_L g3225 ( 
.A1(n_2658),
.A2(n_242),
.B(n_240),
.C(n_241),
.Y(n_3225)
);

CKINVDCx5p33_ASAP7_75t_R g3226 ( 
.A(n_2897),
.Y(n_3226)
);

NAND2xp5_ASAP7_75t_L g3227 ( 
.A(n_2425),
.B(n_240),
.Y(n_3227)
);

INVx1_ASAP7_75t_SL g3228 ( 
.A(n_2549),
.Y(n_3228)
);

OR2x2_ASAP7_75t_L g3229 ( 
.A(n_2416),
.B(n_241),
.Y(n_3229)
);

NAND2xp5_ASAP7_75t_L g3230 ( 
.A(n_2425),
.B(n_242),
.Y(n_3230)
);

NAND2xp5_ASAP7_75t_L g3231 ( 
.A(n_2704),
.B(n_244),
.Y(n_3231)
);

BUFx2_ASAP7_75t_L g3232 ( 
.A(n_2567),
.Y(n_3232)
);

AOI21xp5_ASAP7_75t_L g3233 ( 
.A1(n_2501),
.A2(n_244),
.B(n_245),
.Y(n_3233)
);

NAND2xp5_ASAP7_75t_L g3234 ( 
.A(n_2635),
.B(n_245),
.Y(n_3234)
);

CKINVDCx5p33_ASAP7_75t_R g3235 ( 
.A(n_2897),
.Y(n_3235)
);

BUFx3_ASAP7_75t_L g3236 ( 
.A(n_2506),
.Y(n_3236)
);

OAI22xp5_ASAP7_75t_L g3237 ( 
.A1(n_2789),
.A2(n_247),
.B1(n_245),
.B2(n_246),
.Y(n_3237)
);

INVx2_ASAP7_75t_L g3238 ( 
.A(n_2510),
.Y(n_3238)
);

INVx1_ASAP7_75t_L g3239 ( 
.A(n_2565),
.Y(n_3239)
);

NOR2xp67_ASAP7_75t_L g3240 ( 
.A(n_2520),
.B(n_247),
.Y(n_3240)
);

OAI22xp5_ASAP7_75t_L g3241 ( 
.A1(n_2791),
.A2(n_248),
.B1(n_246),
.B2(n_247),
.Y(n_3241)
);

NAND2xp5_ASAP7_75t_L g3242 ( 
.A(n_2592),
.B(n_2607),
.Y(n_3242)
);

A2O1A1Ixp33_ASAP7_75t_SL g3243 ( 
.A1(n_2804),
.A2(n_249),
.B(n_246),
.C(n_248),
.Y(n_3243)
);

INVx2_ASAP7_75t_SL g3244 ( 
.A(n_2436),
.Y(n_3244)
);

INVx1_ASAP7_75t_L g3245 ( 
.A(n_2571),
.Y(n_3245)
);

NOR2xp33_ASAP7_75t_L g3246 ( 
.A(n_2586),
.B(n_248),
.Y(n_3246)
);

OAI21xp5_ASAP7_75t_L g3247 ( 
.A1(n_2603),
.A2(n_249),
.B(n_250),
.Y(n_3247)
);

AOI21xp5_ASAP7_75t_L g3248 ( 
.A1(n_2624),
.A2(n_249),
.B(n_250),
.Y(n_3248)
);

BUFx3_ASAP7_75t_L g3249 ( 
.A(n_2472),
.Y(n_3249)
);

AOI22xp5_ASAP7_75t_L g3250 ( 
.A1(n_2522),
.A2(n_252),
.B1(n_250),
.B2(n_251),
.Y(n_3250)
);

A2O1A1Ixp33_ASAP7_75t_SL g3251 ( 
.A1(n_2846),
.A2(n_253),
.B(n_251),
.C(n_252),
.Y(n_3251)
);

OAI22xp5_ASAP7_75t_L g3252 ( 
.A1(n_2791),
.A2(n_255),
.B1(n_252),
.B2(n_254),
.Y(n_3252)
);

INVx2_ASAP7_75t_L g3253 ( 
.A(n_2404),
.Y(n_3253)
);

INVx1_ASAP7_75t_L g3254 ( 
.A(n_2572),
.Y(n_3254)
);

INVx1_ASAP7_75t_L g3255 ( 
.A(n_2811),
.Y(n_3255)
);

OR2x2_ASAP7_75t_L g3256 ( 
.A(n_2419),
.B(n_254),
.Y(n_3256)
);

INVx2_ASAP7_75t_L g3257 ( 
.A(n_2769),
.Y(n_3257)
);

NAND2xp5_ASAP7_75t_SL g3258 ( 
.A(n_2643),
.B(n_354),
.Y(n_3258)
);

INVx2_ASAP7_75t_L g3259 ( 
.A(n_2779),
.Y(n_3259)
);

CKINVDCx5p33_ASAP7_75t_R g3260 ( 
.A(n_2450),
.Y(n_3260)
);

BUFx6f_ASAP7_75t_L g3261 ( 
.A(n_2654),
.Y(n_3261)
);

NAND3xp33_ASAP7_75t_L g3262 ( 
.A(n_2467),
.B(n_254),
.C(n_255),
.Y(n_3262)
);

O2A1O1Ixp33_ASAP7_75t_L g3263 ( 
.A1(n_2776),
.A2(n_257),
.B(n_255),
.C(n_256),
.Y(n_3263)
);

NAND2xp5_ASAP7_75t_SL g3264 ( 
.A(n_2643),
.B(n_355),
.Y(n_3264)
);

AOI21xp5_ASAP7_75t_L g3265 ( 
.A1(n_2454),
.A2(n_256),
.B(n_257),
.Y(n_3265)
);

AO21x2_ASAP7_75t_L g3266 ( 
.A1(n_2470),
.A2(n_256),
.B(n_258),
.Y(n_3266)
);

O2A1O1Ixp33_ASAP7_75t_L g3267 ( 
.A1(n_2830),
.A2(n_260),
.B(n_258),
.C(n_259),
.Y(n_3267)
);

AOI21x1_ASAP7_75t_L g3268 ( 
.A1(n_2550),
.A2(n_258),
.B(n_260),
.Y(n_3268)
);

NAND2xp5_ASAP7_75t_L g3269 ( 
.A(n_2718),
.B(n_260),
.Y(n_3269)
);

NOR2xp33_ASAP7_75t_SL g3270 ( 
.A(n_2520),
.B(n_261),
.Y(n_3270)
);

BUFx2_ASAP7_75t_L g3271 ( 
.A(n_2567),
.Y(n_3271)
);

O2A1O1Ixp33_ASAP7_75t_L g3272 ( 
.A1(n_2833),
.A2(n_263),
.B(n_261),
.C(n_262),
.Y(n_3272)
);

AOI21xp5_ASAP7_75t_L g3273 ( 
.A1(n_2458),
.A2(n_261),
.B(n_262),
.Y(n_3273)
);

AND2x2_ASAP7_75t_L g3274 ( 
.A(n_2419),
.B(n_263),
.Y(n_3274)
);

NAND2xp5_ASAP7_75t_SL g3275 ( 
.A(n_2582),
.B(n_355),
.Y(n_3275)
);

NAND2xp5_ASAP7_75t_SL g3276 ( 
.A(n_2527),
.B(n_357),
.Y(n_3276)
);

BUFx2_ASAP7_75t_SL g3277 ( 
.A(n_2455),
.Y(n_3277)
);

INVx2_ASAP7_75t_L g3278 ( 
.A(n_2783),
.Y(n_3278)
);

AND2x2_ASAP7_75t_L g3279 ( 
.A(n_2656),
.B(n_263),
.Y(n_3279)
);

AND2x2_ASAP7_75t_L g3280 ( 
.A(n_2681),
.B(n_264),
.Y(n_3280)
);

AOI21xp5_ASAP7_75t_L g3281 ( 
.A1(n_2466),
.A2(n_264),
.B(n_265),
.Y(n_3281)
);

INVx1_ASAP7_75t_L g3282 ( 
.A(n_2813),
.Y(n_3282)
);

INVx3_ASAP7_75t_L g3283 ( 
.A(n_2589),
.Y(n_3283)
);

INVx1_ASAP7_75t_L g3284 ( 
.A(n_2813),
.Y(n_3284)
);

INVx1_ASAP7_75t_L g3285 ( 
.A(n_2815),
.Y(n_3285)
);

OR2x2_ASAP7_75t_L g3286 ( 
.A(n_2434),
.B(n_264),
.Y(n_3286)
);

INVx2_ASAP7_75t_L g3287 ( 
.A(n_2788),
.Y(n_3287)
);

AOI21xp5_ASAP7_75t_L g3288 ( 
.A1(n_2486),
.A2(n_265),
.B(n_266),
.Y(n_3288)
);

INVx2_ASAP7_75t_L g3289 ( 
.A(n_2797),
.Y(n_3289)
);

AOI21xp5_ASAP7_75t_L g3290 ( 
.A1(n_2675),
.A2(n_265),
.B(n_266),
.Y(n_3290)
);

A2O1A1Ixp33_ASAP7_75t_L g3291 ( 
.A1(n_2676),
.A2(n_268),
.B(n_266),
.C(n_267),
.Y(n_3291)
);

BUFx6f_ASAP7_75t_L g3292 ( 
.A(n_2654),
.Y(n_3292)
);

NAND2xp5_ASAP7_75t_L g3293 ( 
.A(n_2591),
.B(n_267),
.Y(n_3293)
);

NOR2xp67_ASAP7_75t_SL g3294 ( 
.A(n_2527),
.B(n_267),
.Y(n_3294)
);

NOR2xp33_ASAP7_75t_L g3295 ( 
.A(n_2546),
.B(n_268),
.Y(n_3295)
);

NAND2xp5_ASAP7_75t_L g3296 ( 
.A(n_2815),
.B(n_268),
.Y(n_3296)
);

NAND2xp5_ASAP7_75t_L g3297 ( 
.A(n_2840),
.B(n_269),
.Y(n_3297)
);

NAND2xp33_ASAP7_75t_R g3298 ( 
.A(n_2555),
.B(n_2600),
.Y(n_3298)
);

OAI22xp5_ASAP7_75t_L g3299 ( 
.A1(n_2840),
.A2(n_271),
.B1(n_269),
.B2(n_270),
.Y(n_3299)
);

AOI22xp33_ASAP7_75t_L g3300 ( 
.A1(n_2714),
.A2(n_271),
.B1(n_269),
.B2(n_270),
.Y(n_3300)
);

INVx2_ASAP7_75t_L g3301 ( 
.A(n_2800),
.Y(n_3301)
);

INVx1_ASAP7_75t_L g3302 ( 
.A(n_2883),
.Y(n_3302)
);

AOI21xp5_ASAP7_75t_L g3303 ( 
.A1(n_2516),
.A2(n_272),
.B(n_273),
.Y(n_3303)
);

A2O1A1Ixp33_ASAP7_75t_L g3304 ( 
.A1(n_2664),
.A2(n_275),
.B(n_273),
.C(n_274),
.Y(n_3304)
);

CKINVDCx5p33_ASAP7_75t_R g3305 ( 
.A(n_2485),
.Y(n_3305)
);

AOI221x1_ASAP7_75t_L g3306 ( 
.A1(n_2753),
.A2(n_275),
.B1(n_273),
.B2(n_274),
.C(n_276),
.Y(n_3306)
);

OAI22xp5_ASAP7_75t_L g3307 ( 
.A1(n_2883),
.A2(n_276),
.B1(n_274),
.B2(n_275),
.Y(n_3307)
);

NAND2xp5_ASAP7_75t_L g3308 ( 
.A(n_2887),
.B(n_2898),
.Y(n_3308)
);

AOI21x1_ASAP7_75t_L g3309 ( 
.A1(n_2563),
.A2(n_276),
.B(n_277),
.Y(n_3309)
);

AO21x1_ASAP7_75t_L g3310 ( 
.A1(n_2841),
.A2(n_359),
.B(n_358),
.Y(n_3310)
);

NOR2x1_ASAP7_75t_SL g3311 ( 
.A(n_2527),
.B(n_277),
.Y(n_3311)
);

AOI21xp5_ASAP7_75t_L g3312 ( 
.A1(n_2530),
.A2(n_278),
.B(n_279),
.Y(n_3312)
);

OAI22xp5_ASAP7_75t_L g3313 ( 
.A1(n_2887),
.A2(n_2583),
.B1(n_2473),
.B2(n_2773),
.Y(n_3313)
);

AOI21xp5_ASAP7_75t_L g3314 ( 
.A1(n_2434),
.A2(n_279),
.B(n_280),
.Y(n_3314)
);

INVx1_ASAP7_75t_L g3315 ( 
.A(n_2552),
.Y(n_3315)
);

NAND2xp5_ASAP7_75t_SL g3316 ( 
.A(n_2400),
.B(n_359),
.Y(n_3316)
);

CKINVDCx5p33_ASAP7_75t_R g3317 ( 
.A(n_2724),
.Y(n_3317)
);

OAI21x1_ASAP7_75t_L g3318 ( 
.A1(n_2636),
.A2(n_279),
.B(n_280),
.Y(n_3318)
);

AOI21xp5_ASAP7_75t_L g3319 ( 
.A1(n_2441),
.A2(n_280),
.B(n_281),
.Y(n_3319)
);

AOI22xp5_ASAP7_75t_L g3320 ( 
.A1(n_2714),
.A2(n_284),
.B1(n_282),
.B2(n_283),
.Y(n_3320)
);

BUFx6f_ASAP7_75t_SL g3321 ( 
.A(n_2618),
.Y(n_3321)
);

CKINVDCx5p33_ASAP7_75t_R g3322 ( 
.A(n_2701),
.Y(n_3322)
);

AND2x2_ASAP7_75t_L g3323 ( 
.A(n_2552),
.B(n_282),
.Y(n_3323)
);

NOR2xp33_ASAP7_75t_R g3324 ( 
.A(n_2558),
.B(n_283),
.Y(n_3324)
);

AND2x2_ASAP7_75t_L g3325 ( 
.A(n_2879),
.B(n_2618),
.Y(n_3325)
);

AOI221xp5_ASAP7_75t_L g3326 ( 
.A1(n_2863),
.A2(n_285),
.B1(n_283),
.B2(n_284),
.C(n_286),
.Y(n_3326)
);

NOR2xp33_ASAP7_75t_L g3327 ( 
.A(n_2733),
.B(n_284),
.Y(n_3327)
);

OAI21xp33_ASAP7_75t_SL g3328 ( 
.A1(n_2784),
.A2(n_287),
.B(n_286),
.Y(n_3328)
);

OAI22xp5_ASAP7_75t_L g3329 ( 
.A1(n_2473),
.A2(n_288),
.B1(n_285),
.B2(n_286),
.Y(n_3329)
);

OAI21xp33_ASAP7_75t_SL g3330 ( 
.A1(n_2829),
.A2(n_291),
.B(n_290),
.Y(n_3330)
);

NAND2xp5_ASAP7_75t_L g3331 ( 
.A(n_2441),
.B(n_289),
.Y(n_3331)
);

INVx1_ASAP7_75t_L g3332 ( 
.A(n_2518),
.Y(n_3332)
);

NAND2xp5_ASAP7_75t_SL g3333 ( 
.A(n_2405),
.B(n_360),
.Y(n_3333)
);

AOI21xp5_ASAP7_75t_L g3334 ( 
.A1(n_2443),
.A2(n_289),
.B(n_290),
.Y(n_3334)
);

NAND2xp5_ASAP7_75t_L g3335 ( 
.A(n_2443),
.B(n_291),
.Y(n_3335)
);

INVx1_ASAP7_75t_L g3336 ( 
.A(n_2533),
.Y(n_3336)
);

A2O1A1Ixp33_ASAP7_75t_L g3337 ( 
.A1(n_2470),
.A2(n_294),
.B(n_292),
.C(n_293),
.Y(n_3337)
);

BUFx3_ASAP7_75t_L g3338 ( 
.A(n_2455),
.Y(n_3338)
);

INVx4_ASAP7_75t_L g3339 ( 
.A(n_2455),
.Y(n_3339)
);

INVx1_ASAP7_75t_L g3340 ( 
.A(n_2542),
.Y(n_3340)
);

BUFx2_ASAP7_75t_L g3341 ( 
.A(n_2567),
.Y(n_3341)
);

AOI21xp5_ASAP7_75t_L g3342 ( 
.A1(n_2449),
.A2(n_292),
.B(n_293),
.Y(n_3342)
);

BUFx6f_ASAP7_75t_L g3343 ( 
.A(n_2654),
.Y(n_3343)
);

OAI22xp5_ASAP7_75t_L g3344 ( 
.A1(n_2849),
.A2(n_2449),
.B1(n_2731),
.B2(n_2730),
.Y(n_3344)
);

AOI21xp5_ASAP7_75t_L g3345 ( 
.A1(n_2545),
.A2(n_294),
.B(n_295),
.Y(n_3345)
);

INVx2_ASAP7_75t_L g3346 ( 
.A(n_2822),
.Y(n_3346)
);

AOI21xp5_ASAP7_75t_L g3347 ( 
.A1(n_2702),
.A2(n_294),
.B(n_295),
.Y(n_3347)
);

NOR2xp33_ASAP7_75t_L g3348 ( 
.A(n_2733),
.B(n_295),
.Y(n_3348)
);

AOI22xp5_ASAP7_75t_L g3349 ( 
.A1(n_2748),
.A2(n_298),
.B1(n_296),
.B2(n_297),
.Y(n_3349)
);

BUFx2_ASAP7_75t_R g3350 ( 
.A(n_2913),
.Y(n_3350)
);

NAND2xp5_ASAP7_75t_L g3351 ( 
.A(n_2908),
.B(n_2748),
.Y(n_3351)
);

NOR2x1_ASAP7_75t_L g3352 ( 
.A(n_3130),
.B(n_2701),
.Y(n_3352)
);

INVx2_ASAP7_75t_L g3353 ( 
.A(n_3047),
.Y(n_3353)
);

NAND2xp5_ASAP7_75t_L g3354 ( 
.A(n_3071),
.B(n_2922),
.Y(n_3354)
);

INVx2_ASAP7_75t_L g3355 ( 
.A(n_3067),
.Y(n_3355)
);

AND2x2_ASAP7_75t_L g3356 ( 
.A(n_3031),
.B(n_2701),
.Y(n_3356)
);

OAI21xp33_ASAP7_75t_SL g3357 ( 
.A1(n_2972),
.A2(n_2476),
.B(n_2866),
.Y(n_3357)
);

O2A1O1Ixp5_ASAP7_75t_L g3358 ( 
.A1(n_2914),
.A2(n_2577),
.B(n_2861),
.C(n_2848),
.Y(n_3358)
);

NAND2xp5_ASAP7_75t_L g3359 ( 
.A(n_3018),
.B(n_2645),
.Y(n_3359)
);

OAI21xp5_ASAP7_75t_L g3360 ( 
.A1(n_3313),
.A2(n_2777),
.B(n_2720),
.Y(n_3360)
);

AOI21xp5_ASAP7_75t_L g3361 ( 
.A1(n_3172),
.A2(n_2611),
.B(n_2531),
.Y(n_3361)
);

BUFx12f_ASAP7_75t_L g3362 ( 
.A(n_3084),
.Y(n_3362)
);

AND2x2_ASAP7_75t_L g3363 ( 
.A(n_3032),
.B(n_2645),
.Y(n_3363)
);

CKINVDCx20_ASAP7_75t_R g3364 ( 
.A(n_3092),
.Y(n_3364)
);

OAI21xp5_ASAP7_75t_L g3365 ( 
.A1(n_2988),
.A2(n_2777),
.B(n_2691),
.Y(n_3365)
);

OAI21x1_ASAP7_75t_L g3366 ( 
.A1(n_2937),
.A2(n_2594),
.B(n_2575),
.Y(n_3366)
);

INVx2_ASAP7_75t_L g3367 ( 
.A(n_3116),
.Y(n_3367)
);

INVx3_ASAP7_75t_L g3368 ( 
.A(n_3001),
.Y(n_3368)
);

NAND2xp5_ASAP7_75t_L g3369 ( 
.A(n_2911),
.B(n_2700),
.Y(n_3369)
);

CKINVDCx20_ASAP7_75t_R g3370 ( 
.A(n_2978),
.Y(n_3370)
);

O2A1O1Ixp33_ASAP7_75t_SL g3371 ( 
.A1(n_2989),
.A2(n_2661),
.B(n_2456),
.C(n_2700),
.Y(n_3371)
);

INVx3_ASAP7_75t_SL g3372 ( 
.A(n_3008),
.Y(n_3372)
);

BUFx2_ASAP7_75t_L g3373 ( 
.A(n_3001),
.Y(n_3373)
);

O2A1O1Ixp33_ASAP7_75t_SL g3374 ( 
.A1(n_2996),
.A2(n_2705),
.B(n_2688),
.C(n_2671),
.Y(n_3374)
);

NAND2xp5_ASAP7_75t_L g3375 ( 
.A(n_3255),
.B(n_2705),
.Y(n_3375)
);

INVx1_ASAP7_75t_L g3376 ( 
.A(n_3002),
.Y(n_3376)
);

INVx1_ASAP7_75t_L g3377 ( 
.A(n_3051),
.Y(n_3377)
);

NAND2xp5_ASAP7_75t_L g3378 ( 
.A(n_3282),
.B(n_2739),
.Y(n_3378)
);

NAND2xp33_ASAP7_75t_R g3379 ( 
.A(n_2980),
.B(n_2599),
.Y(n_3379)
);

OAI21x1_ASAP7_75t_L g3380 ( 
.A1(n_3000),
.A2(n_2594),
.B(n_2566),
.Y(n_3380)
);

AND2x2_ASAP7_75t_L g3381 ( 
.A(n_3178),
.B(n_3274),
.Y(n_3381)
);

NAND2xp5_ASAP7_75t_L g3382 ( 
.A(n_3284),
.B(n_2729),
.Y(n_3382)
);

INVx2_ASAP7_75t_L g3383 ( 
.A(n_3119),
.Y(n_3383)
);

AOI21xp5_ASAP7_75t_L g3384 ( 
.A1(n_3029),
.A2(n_2772),
.B(n_2766),
.Y(n_3384)
);

OA22x2_ASAP7_75t_L g3385 ( 
.A1(n_3166),
.A2(n_2599),
.B1(n_2764),
.B2(n_2488),
.Y(n_3385)
);

NAND2xp33_ASAP7_75t_R g3386 ( 
.A(n_3163),
.B(n_2599),
.Y(n_3386)
);

AOI21xp5_ASAP7_75t_L g3387 ( 
.A1(n_2992),
.A2(n_2772),
.B(n_2766),
.Y(n_3387)
);

NAND2xp5_ASAP7_75t_L g3388 ( 
.A(n_3285),
.B(n_2688),
.Y(n_3388)
);

BUFx6f_ASAP7_75t_L g3389 ( 
.A(n_2968),
.Y(n_3389)
);

O2A1O1Ixp5_ASAP7_75t_L g3390 ( 
.A1(n_3275),
.A2(n_2595),
.B(n_2763),
.C(n_2746),
.Y(n_3390)
);

INVx4_ASAP7_75t_L g3391 ( 
.A(n_3001),
.Y(n_3391)
);

INVx2_ASAP7_75t_L g3392 ( 
.A(n_3132),
.Y(n_3392)
);

AO31x2_ASAP7_75t_L g3393 ( 
.A1(n_2930),
.A2(n_2751),
.A3(n_2759),
.B(n_2758),
.Y(n_3393)
);

AOI21xp5_ASAP7_75t_L g3394 ( 
.A1(n_3308),
.A2(n_2871),
.B(n_2865),
.Y(n_3394)
);

OR2x2_ASAP7_75t_L g3395 ( 
.A(n_2929),
.B(n_2477),
.Y(n_3395)
);

OAI21x1_ASAP7_75t_L g3396 ( 
.A1(n_3096),
.A2(n_2581),
.B(n_2660),
.Y(n_3396)
);

O2A1O1Ixp33_ASAP7_75t_L g3397 ( 
.A1(n_3344),
.A2(n_3243),
.B(n_3251),
.C(n_3091),
.Y(n_3397)
);

INVx1_ASAP7_75t_L g3398 ( 
.A(n_3063),
.Y(n_3398)
);

INVx1_ASAP7_75t_L g3399 ( 
.A(n_3068),
.Y(n_3399)
);

AOI21xp5_ASAP7_75t_L g3400 ( 
.A1(n_3048),
.A2(n_2871),
.B(n_2865),
.Y(n_3400)
);

BUFx2_ASAP7_75t_L g3401 ( 
.A(n_2907),
.Y(n_3401)
);

OAI21x1_ASAP7_75t_L g3402 ( 
.A1(n_3283),
.A2(n_2483),
.B(n_2678),
.Y(n_3402)
);

AOI21xp5_ASAP7_75t_L g3403 ( 
.A1(n_3076),
.A2(n_2871),
.B(n_2865),
.Y(n_3403)
);

OAI21xp5_ASAP7_75t_L g3404 ( 
.A1(n_2991),
.A2(n_2479),
.B(n_2507),
.Y(n_3404)
);

NOR2xp67_ASAP7_75t_SL g3405 ( 
.A(n_3112),
.B(n_3277),
.Y(n_3405)
);

NAND2xp5_ASAP7_75t_L g3406 ( 
.A(n_3302),
.B(n_3073),
.Y(n_3406)
);

O2A1O1Ixp33_ASAP7_75t_L g3407 ( 
.A1(n_3159),
.A2(n_2596),
.B(n_2745),
.C(n_2532),
.Y(n_3407)
);

BUFx6f_ASAP7_75t_L g3408 ( 
.A(n_2968),
.Y(n_3408)
);

AOI21xp5_ASAP7_75t_L g3409 ( 
.A1(n_3097),
.A2(n_2772),
.B(n_2766),
.Y(n_3409)
);

INVx1_ASAP7_75t_L g3410 ( 
.A(n_3098),
.Y(n_3410)
);

NAND2xp5_ASAP7_75t_L g3411 ( 
.A(n_3103),
.B(n_2842),
.Y(n_3411)
);

INVx2_ASAP7_75t_L g3412 ( 
.A(n_2906),
.Y(n_3412)
);

A2O1A1Ixp33_ASAP7_75t_L g3413 ( 
.A1(n_3061),
.A2(n_2764),
.B(n_2894),
.C(n_2855),
.Y(n_3413)
);

NAND3xp33_ASAP7_75t_SL g3414 ( 
.A(n_3171),
.B(n_2728),
.C(n_2709),
.Y(n_3414)
);

AOI21xp5_ASAP7_75t_L g3415 ( 
.A1(n_3112),
.A2(n_2818),
.B(n_2802),
.Y(n_3415)
);

AOI21xp33_ASAP7_75t_L g3416 ( 
.A1(n_2940),
.A2(n_2758),
.B(n_2751),
.Y(n_3416)
);

OAI22xp5_ASAP7_75t_L g3417 ( 
.A1(n_3112),
.A2(n_2863),
.B1(n_2653),
.B2(n_2610),
.Y(n_3417)
);

NAND2x1p5_ASAP7_75t_L g3418 ( 
.A(n_3045),
.B(n_2590),
.Y(n_3418)
);

NAND2xp5_ASAP7_75t_L g3419 ( 
.A(n_3113),
.B(n_2526),
.Y(n_3419)
);

NAND2xp5_ASAP7_75t_SL g3420 ( 
.A(n_3322),
.B(n_2726),
.Y(n_3420)
);

A2O1A1Ixp33_ASAP7_75t_L g3421 ( 
.A1(n_2941),
.A2(n_2884),
.B(n_2679),
.C(n_2528),
.Y(n_3421)
);

INVx4_ASAP7_75t_L g3422 ( 
.A(n_3074),
.Y(n_3422)
);

AND2x2_ASAP7_75t_L g3423 ( 
.A(n_3279),
.B(n_2512),
.Y(n_3423)
);

OAI21x1_ASAP7_75t_L g3424 ( 
.A1(n_3283),
.A2(n_2525),
.B(n_2509),
.Y(n_3424)
);

INVx1_ASAP7_75t_L g3425 ( 
.A(n_3115),
.Y(n_3425)
);

A2O1A1Ixp33_ASAP7_75t_L g3426 ( 
.A1(n_3206),
.A2(n_2884),
.B(n_2528),
.C(n_2551),
.Y(n_3426)
);

BUFx3_ASAP7_75t_L g3427 ( 
.A(n_3054),
.Y(n_3427)
);

NAND2xp5_ASAP7_75t_SL g3428 ( 
.A(n_2970),
.B(n_2726),
.Y(n_3428)
);

AO21x2_ASAP7_75t_L g3429 ( 
.A1(n_3058),
.A2(n_2759),
.B(n_2490),
.Y(n_3429)
);

INVx3_ASAP7_75t_L g3430 ( 
.A(n_3045),
.Y(n_3430)
);

AOI21xp5_ASAP7_75t_L g3431 ( 
.A1(n_3110),
.A2(n_2802),
.B(n_2798),
.Y(n_3431)
);

HB1xp67_ASAP7_75t_L g3432 ( 
.A(n_2936),
.Y(n_3432)
);

OAI21xp5_ASAP7_75t_L g3433 ( 
.A1(n_3262),
.A2(n_2529),
.B(n_2744),
.Y(n_3433)
);

OAI21xp5_ASAP7_75t_L g3434 ( 
.A1(n_3304),
.A2(n_2512),
.B(n_2765),
.Y(n_3434)
);

BUFx6f_ASAP7_75t_L g3435 ( 
.A(n_2968),
.Y(n_3435)
);

BUFx2_ASAP7_75t_L g3436 ( 
.A(n_3130),
.Y(n_3436)
);

NAND2xp33_ASAP7_75t_L g3437 ( 
.A(n_3324),
.B(n_2570),
.Y(n_3437)
);

NAND2xp5_ASAP7_75t_L g3438 ( 
.A(n_3121),
.B(n_2526),
.Y(n_3438)
);

O2A1O1Ixp33_ASAP7_75t_L g3439 ( 
.A1(n_3030),
.A2(n_2622),
.B(n_2757),
.C(n_2711),
.Y(n_3439)
);

NAND2xp33_ASAP7_75t_R g3440 ( 
.A(n_3317),
.B(n_2403),
.Y(n_3440)
);

NAND2xp5_ASAP7_75t_L g3441 ( 
.A(n_3129),
.B(n_3204),
.Y(n_3441)
);

INVxp67_ASAP7_75t_SL g3442 ( 
.A(n_3174),
.Y(n_3442)
);

AO31x2_ASAP7_75t_L g3443 ( 
.A1(n_2935),
.A2(n_2585),
.A3(n_2576),
.B(n_2746),
.Y(n_3443)
);

NAND2xp5_ASAP7_75t_L g3444 ( 
.A(n_3212),
.B(n_2551),
.Y(n_3444)
);

AO31x2_ASAP7_75t_L g3445 ( 
.A1(n_3306),
.A2(n_2585),
.A3(n_2576),
.B(n_2857),
.Y(n_3445)
);

INVx2_ASAP7_75t_SL g3446 ( 
.A(n_3124),
.Y(n_3446)
);

NAND2xp5_ASAP7_75t_L g3447 ( 
.A(n_3066),
.B(n_2403),
.Y(n_3447)
);

NAND2xp5_ASAP7_75t_L g3448 ( 
.A(n_3083),
.B(n_2477),
.Y(n_3448)
);

NAND2xp5_ASAP7_75t_L g3449 ( 
.A(n_3286),
.B(n_2493),
.Y(n_3449)
);

AO21x2_ASAP7_75t_L g3450 ( 
.A1(n_3209),
.A2(n_2481),
.B(n_2620),
.Y(n_3450)
);

INVx1_ASAP7_75t_L g3451 ( 
.A(n_3133),
.Y(n_3451)
);

INVxp67_ASAP7_75t_SL g3452 ( 
.A(n_3148),
.Y(n_3452)
);

OAI21x1_ASAP7_75t_L g3453 ( 
.A1(n_3110),
.A2(n_2514),
.B(n_2496),
.Y(n_3453)
);

AOI21xp5_ASAP7_75t_L g3454 ( 
.A1(n_3296),
.A2(n_2802),
.B(n_2798),
.Y(n_3454)
);

NAND2xp5_ASAP7_75t_L g3455 ( 
.A(n_3227),
.B(n_2493),
.Y(n_3455)
);

NAND2xp5_ASAP7_75t_L g3456 ( 
.A(n_3230),
.B(n_2502),
.Y(n_3456)
);

AO31x2_ASAP7_75t_L g3457 ( 
.A1(n_3310),
.A2(n_2860),
.A3(n_2864),
.B(n_2859),
.Y(n_3457)
);

AOI21xp5_ASAP7_75t_L g3458 ( 
.A1(n_3297),
.A2(n_2814),
.B(n_2798),
.Y(n_3458)
);

NAND2xp5_ASAP7_75t_L g3459 ( 
.A(n_3180),
.B(n_2502),
.Y(n_3459)
);

OR2x2_ASAP7_75t_L g3460 ( 
.A(n_2961),
.B(n_2547),
.Y(n_3460)
);

INVx2_ASAP7_75t_L g3461 ( 
.A(n_2921),
.Y(n_3461)
);

AOI21x1_ASAP7_75t_L g3462 ( 
.A1(n_3232),
.A2(n_2538),
.B(n_2740),
.Y(n_3462)
);

INVx3_ASAP7_75t_L g3463 ( 
.A(n_2951),
.Y(n_3463)
);

AOI21xp5_ASAP7_75t_SL g3464 ( 
.A1(n_2920),
.A2(n_2818),
.B(n_2814),
.Y(n_3464)
);

OAI21x1_ASAP7_75t_L g3465 ( 
.A1(n_3268),
.A2(n_3309),
.B(n_3318),
.Y(n_3465)
);

INVx3_ASAP7_75t_L g3466 ( 
.A(n_3074),
.Y(n_3466)
);

OAI21xp5_ASAP7_75t_L g3467 ( 
.A1(n_3312),
.A2(n_2620),
.B(n_2762),
.Y(n_3467)
);

OAI21x1_ASAP7_75t_L g3468 ( 
.A1(n_3248),
.A2(n_2593),
.B(n_2560),
.Y(n_3468)
);

BUFx3_ASAP7_75t_L g3469 ( 
.A(n_3236),
.Y(n_3469)
);

AOI21xp5_ASAP7_75t_L g3470 ( 
.A1(n_2915),
.A2(n_2818),
.B(n_2814),
.Y(n_3470)
);

INVx1_ASAP7_75t_L g3471 ( 
.A(n_3141),
.Y(n_3471)
);

BUFx6f_ASAP7_75t_L g3472 ( 
.A(n_2969),
.Y(n_3472)
);

NOR2xp33_ASAP7_75t_L g3473 ( 
.A(n_3043),
.B(n_2648),
.Y(n_3473)
);

NAND2xp5_ASAP7_75t_SL g3474 ( 
.A(n_3271),
.B(n_2726),
.Y(n_3474)
);

OAI21x1_ASAP7_75t_L g3475 ( 
.A1(n_2950),
.A2(n_2997),
.B(n_2963),
.Y(n_3475)
);

AOI21xp5_ASAP7_75t_L g3476 ( 
.A1(n_2917),
.A2(n_2698),
.B(n_2536),
.Y(n_3476)
);

INVx1_ASAP7_75t_L g3477 ( 
.A(n_3160),
.Y(n_3477)
);

INVx6_ASAP7_75t_SL g3478 ( 
.A(n_3059),
.Y(n_3478)
);

AND2x2_ASAP7_75t_L g3479 ( 
.A(n_3323),
.B(n_2612),
.Y(n_3479)
);

BUFx3_ASAP7_75t_L g3480 ( 
.A(n_3144),
.Y(n_3480)
);

OAI21x1_ASAP7_75t_L g3481 ( 
.A1(n_2998),
.A2(n_2593),
.B(n_2560),
.Y(n_3481)
);

AOI21x1_ASAP7_75t_L g3482 ( 
.A1(n_3341),
.A2(n_2760),
.B(n_2638),
.Y(n_3482)
);

NAND3xp33_ASAP7_75t_L g3483 ( 
.A(n_3126),
.B(n_2925),
.C(n_3184),
.Y(n_3483)
);

AOI21xp5_ASAP7_75t_L g3484 ( 
.A1(n_3242),
.A2(n_2698),
.B(n_2870),
.Y(n_3484)
);

INVx2_ASAP7_75t_L g3485 ( 
.A(n_2939),
.Y(n_3485)
);

INVx5_ASAP7_75t_L g3486 ( 
.A(n_3124),
.Y(n_3486)
);

BUFx4f_ASAP7_75t_L g3487 ( 
.A(n_3059),
.Y(n_3487)
);

AOI21xp5_ASAP7_75t_L g3488 ( 
.A1(n_3331),
.A2(n_3335),
.B(n_3183),
.Y(n_3488)
);

NOR2xp33_ASAP7_75t_L g3489 ( 
.A(n_3321),
.B(n_2648),
.Y(n_3489)
);

INVx1_ASAP7_75t_L g3490 ( 
.A(n_3189),
.Y(n_3490)
);

OAI21x1_ASAP7_75t_L g3491 ( 
.A1(n_3060),
.A2(n_2511),
.B(n_2489),
.Y(n_3491)
);

OR2x2_ASAP7_75t_L g3492 ( 
.A(n_2966),
.B(n_2625),
.Y(n_3492)
);

AOI21xp5_ASAP7_75t_SL g3493 ( 
.A1(n_3033),
.A2(n_2570),
.B(n_2716),
.Y(n_3493)
);

AO31x2_ASAP7_75t_L g3494 ( 
.A1(n_3065),
.A2(n_2891),
.A3(n_2900),
.B(n_2882),
.Y(n_3494)
);

OA21x2_ASAP7_75t_L g3495 ( 
.A1(n_3176),
.A2(n_3247),
.B(n_3216),
.Y(n_3495)
);

NAND2xp5_ASAP7_75t_SL g3496 ( 
.A(n_3270),
.B(n_2716),
.Y(n_3496)
);

INVx2_ASAP7_75t_L g3497 ( 
.A(n_2949),
.Y(n_3497)
);

NAND3x1_ASAP7_75t_L g3498 ( 
.A(n_3217),
.B(n_2680),
.C(n_2756),
.Y(n_3498)
);

OAI21xp5_ASAP7_75t_L g3499 ( 
.A1(n_3303),
.A2(n_2570),
.B(n_2650),
.Y(n_3499)
);

CKINVDCx20_ASAP7_75t_R g3500 ( 
.A(n_3075),
.Y(n_3500)
);

INVx1_ASAP7_75t_L g3501 ( 
.A(n_3205),
.Y(n_3501)
);

INVx4_ASAP7_75t_L g3502 ( 
.A(n_3144),
.Y(n_3502)
);

NAND2xp5_ASAP7_75t_L g3503 ( 
.A(n_3055),
.B(n_2627),
.Y(n_3503)
);

BUFx2_ASAP7_75t_L g3504 ( 
.A(n_2919),
.Y(n_3504)
);

NAND2xp5_ASAP7_75t_L g3505 ( 
.A(n_3210),
.B(n_2630),
.Y(n_3505)
);

OAI21xp5_ASAP7_75t_L g3506 ( 
.A1(n_3064),
.A2(n_2570),
.B(n_2633),
.Y(n_3506)
);

INVx4_ASAP7_75t_L g3507 ( 
.A(n_3015),
.Y(n_3507)
);

OA21x2_ASAP7_75t_L g3508 ( 
.A1(n_2947),
.A2(n_2696),
.B(n_2667),
.Y(n_3508)
);

NAND2xp5_ASAP7_75t_L g3509 ( 
.A(n_3239),
.B(n_2634),
.Y(n_3509)
);

OAI21xp5_ASAP7_75t_L g3510 ( 
.A1(n_3233),
.A2(n_3273),
.B(n_3265),
.Y(n_3510)
);

OAI21x1_ASAP7_75t_L g3511 ( 
.A1(n_3060),
.A2(n_2511),
.B(n_2489),
.Y(n_3511)
);

OA21x2_ASAP7_75t_L g3512 ( 
.A1(n_2953),
.A2(n_2535),
.B(n_2523),
.Y(n_3512)
);

AOI221x1_ASAP7_75t_L g3513 ( 
.A1(n_3044),
.A2(n_2756),
.B1(n_2698),
.B2(n_2569),
.C(n_2574),
.Y(n_3513)
);

OAI21x1_ASAP7_75t_SL g3514 ( 
.A1(n_3311),
.A2(n_2544),
.B(n_2539),
.Y(n_3514)
);

OAI21x1_ASAP7_75t_L g3515 ( 
.A1(n_3139),
.A2(n_2632),
.B(n_2652),
.Y(n_3515)
);

AOI21xp5_ASAP7_75t_L g3516 ( 
.A1(n_2977),
.A2(n_2986),
.B(n_3006),
.Y(n_3516)
);

AOI21xp5_ASAP7_75t_L g3517 ( 
.A1(n_3128),
.A2(n_2638),
.B(n_2629),
.Y(n_3517)
);

O2A1O1Ixp5_ASAP7_75t_L g3518 ( 
.A1(n_3294),
.A2(n_2589),
.B(n_2712),
.C(n_2638),
.Y(n_3518)
);

NOR3xp33_ASAP7_75t_L g3519 ( 
.A(n_2981),
.B(n_2684),
.C(n_2629),
.Y(n_3519)
);

AOI21xp5_ASAP7_75t_L g3520 ( 
.A1(n_3035),
.A2(n_2629),
.B(n_2589),
.Y(n_3520)
);

AOI21xp5_ASAP7_75t_L g3521 ( 
.A1(n_3062),
.A2(n_2589),
.B(n_2712),
.Y(n_3521)
);

AND3x4_ASAP7_75t_L g3522 ( 
.A(n_3149),
.B(n_296),
.C(n_297),
.Y(n_3522)
);

INVx1_ASAP7_75t_L g3523 ( 
.A(n_3245),
.Y(n_3523)
);

OAI21x1_ASAP7_75t_SL g3524 ( 
.A1(n_2990),
.A2(n_2712),
.B(n_296),
.Y(n_3524)
);

INVxp67_ASAP7_75t_SL g3525 ( 
.A(n_3148),
.Y(n_3525)
);

AOI21xp5_ASAP7_75t_L g3526 ( 
.A1(n_3069),
.A2(n_2712),
.B(n_297),
.Y(n_3526)
);

NAND2xp5_ASAP7_75t_L g3527 ( 
.A(n_3254),
.B(n_298),
.Y(n_3527)
);

AND2x4_ASAP7_75t_L g3528 ( 
.A(n_3139),
.B(n_298),
.Y(n_3528)
);

NAND3xp33_ASAP7_75t_L g3529 ( 
.A(n_2983),
.B(n_2712),
.C(n_299),
.Y(n_3529)
);

NAND3x1_ASAP7_75t_L g3530 ( 
.A(n_2938),
.B(n_299),
.C(n_300),
.Y(n_3530)
);

INVx1_ASAP7_75t_L g3531 ( 
.A(n_2987),
.Y(n_3531)
);

AOI22xp5_ASAP7_75t_L g3532 ( 
.A1(n_3223),
.A2(n_302),
.B1(n_300),
.B2(n_301),
.Y(n_3532)
);

BUFx6f_ASAP7_75t_L g3533 ( 
.A(n_2969),
.Y(n_3533)
);

INVx1_ASAP7_75t_L g3534 ( 
.A(n_3332),
.Y(n_3534)
);

AOI21xp5_ASAP7_75t_L g3535 ( 
.A1(n_3081),
.A2(n_300),
.B(n_301),
.Y(n_3535)
);

AOI221x1_ASAP7_75t_L g3536 ( 
.A1(n_2932),
.A2(n_304),
.B1(n_302),
.B2(n_303),
.C(n_305),
.Y(n_3536)
);

INVx3_ASAP7_75t_L g3537 ( 
.A(n_3145),
.Y(n_3537)
);

NOR2xp67_ASAP7_75t_L g3538 ( 
.A(n_2919),
.B(n_302),
.Y(n_3538)
);

AO21x2_ASAP7_75t_L g3539 ( 
.A1(n_3147),
.A2(n_304),
.B(n_305),
.Y(n_3539)
);

AND2x2_ASAP7_75t_L g3540 ( 
.A(n_2957),
.B(n_304),
.Y(n_3540)
);

OAI21xp5_ASAP7_75t_L g3541 ( 
.A1(n_3281),
.A2(n_305),
.B(n_306),
.Y(n_3541)
);

AOI21x1_ASAP7_75t_L g3542 ( 
.A1(n_3211),
.A2(n_362),
.B(n_361),
.Y(n_3542)
);

NAND2xp5_ASAP7_75t_L g3543 ( 
.A(n_3325),
.B(n_306),
.Y(n_3543)
);

AND2x2_ASAP7_75t_L g3544 ( 
.A(n_2932),
.B(n_307),
.Y(n_3544)
);

OAI21x1_ASAP7_75t_L g3545 ( 
.A1(n_3158),
.A2(n_309),
.B(n_308),
.Y(n_3545)
);

NAND2xp5_ASAP7_75t_SL g3546 ( 
.A(n_3215),
.B(n_307),
.Y(n_3546)
);

CKINVDCx5p33_ASAP7_75t_R g3547 ( 
.A(n_3015),
.Y(n_3547)
);

NAND2xp5_ASAP7_75t_L g3548 ( 
.A(n_3016),
.B(n_307),
.Y(n_3548)
);

AOI21xp5_ASAP7_75t_L g3549 ( 
.A1(n_3088),
.A2(n_308),
.B(n_309),
.Y(n_3549)
);

A2O1A1Ixp33_ASAP7_75t_L g3550 ( 
.A1(n_3206),
.A2(n_310),
.B(n_308),
.C(n_309),
.Y(n_3550)
);

INVx1_ASAP7_75t_L g3551 ( 
.A(n_3336),
.Y(n_3551)
);

OAI21x1_ASAP7_75t_L g3552 ( 
.A1(n_3158),
.A2(n_312),
.B(n_311),
.Y(n_3552)
);

NAND2xp5_ASAP7_75t_L g3553 ( 
.A(n_3218),
.B(n_310),
.Y(n_3553)
);

INVx5_ASAP7_75t_L g3554 ( 
.A(n_3145),
.Y(n_3554)
);

AND2x2_ASAP7_75t_L g3555 ( 
.A(n_3256),
.B(n_310),
.Y(n_3555)
);

A2O1A1Ixp33_ASAP7_75t_L g3556 ( 
.A1(n_3328),
.A2(n_313),
.B(n_311),
.C(n_312),
.Y(n_3556)
);

INVx1_ASAP7_75t_L g3557 ( 
.A(n_3340),
.Y(n_3557)
);

OAI21x1_ASAP7_75t_L g3558 ( 
.A1(n_2927),
.A2(n_314),
.B(n_313),
.Y(n_3558)
);

AO31x2_ASAP7_75t_L g3559 ( 
.A1(n_3089),
.A2(n_315),
.A3(n_311),
.B(n_314),
.Y(n_3559)
);

INVx1_ASAP7_75t_L g3560 ( 
.A(n_3138),
.Y(n_3560)
);

AND2x2_ASAP7_75t_L g3561 ( 
.A(n_2993),
.B(n_3146),
.Y(n_3561)
);

AOI21xp5_ASAP7_75t_L g3562 ( 
.A1(n_2969),
.A2(n_314),
.B(n_315),
.Y(n_3562)
);

OAI21x1_ASAP7_75t_L g3563 ( 
.A1(n_3211),
.A2(n_317),
.B(n_316),
.Y(n_3563)
);

INVx1_ASAP7_75t_SL g3564 ( 
.A(n_3228),
.Y(n_3564)
);

AOI21x1_ASAP7_75t_L g3565 ( 
.A1(n_3147),
.A2(n_362),
.B(n_361),
.Y(n_3565)
);

NAND2xp5_ASAP7_75t_L g3566 ( 
.A(n_3229),
.B(n_315),
.Y(n_3566)
);

BUFx6f_ASAP7_75t_L g3567 ( 
.A(n_2985),
.Y(n_3567)
);

INVx1_ASAP7_75t_L g3568 ( 
.A(n_3156),
.Y(n_3568)
);

AOI21xp5_ASAP7_75t_L g3569 ( 
.A1(n_2985),
.A2(n_316),
.B(n_317),
.Y(n_3569)
);

AOI21x1_ASAP7_75t_SL g3570 ( 
.A1(n_3222),
.A2(n_317),
.B(n_318),
.Y(n_3570)
);

INVx2_ASAP7_75t_L g3571 ( 
.A(n_3164),
.Y(n_3571)
);

OAI21x1_ASAP7_75t_SL g3572 ( 
.A1(n_3007),
.A2(n_318),
.B(n_319),
.Y(n_3572)
);

NAND2xp5_ASAP7_75t_L g3573 ( 
.A(n_3026),
.B(n_318),
.Y(n_3573)
);

XOR2xp5_ASAP7_75t_L g3574 ( 
.A(n_3226),
.B(n_319),
.Y(n_3574)
);

AOI21xp5_ASAP7_75t_L g3575 ( 
.A1(n_2985),
.A2(n_319),
.B(n_320),
.Y(n_3575)
);

OAI21x1_ASAP7_75t_L g3576 ( 
.A1(n_3345),
.A2(n_322),
.B(n_321),
.Y(n_3576)
);

INVx1_ASAP7_75t_L g3577 ( 
.A(n_3173),
.Y(n_3577)
);

AO31x2_ASAP7_75t_L g3578 ( 
.A1(n_3101),
.A2(n_322),
.A3(n_320),
.B(n_321),
.Y(n_3578)
);

AOI21xp5_ASAP7_75t_L g3579 ( 
.A1(n_3005),
.A2(n_320),
.B(n_321),
.Y(n_3579)
);

NAND2xp5_ASAP7_75t_SL g3580 ( 
.A(n_3215),
.B(n_322),
.Y(n_3580)
);

BUFx6f_ASAP7_75t_L g3581 ( 
.A(n_3005),
.Y(n_3581)
);

NOR2xp67_ASAP7_75t_SL g3582 ( 
.A(n_2934),
.B(n_323),
.Y(n_3582)
);

INVx1_ASAP7_75t_SL g3583 ( 
.A(n_3106),
.Y(n_3583)
);

NAND2x1p5_ASAP7_75t_L g3584 ( 
.A(n_2934),
.B(n_323),
.Y(n_3584)
);

BUFx12f_ASAP7_75t_L g3585 ( 
.A(n_3087),
.Y(n_3585)
);

NAND2xp33_ASAP7_75t_R g3586 ( 
.A(n_3235),
.B(n_323),
.Y(n_3586)
);

INVxp67_ASAP7_75t_SL g3587 ( 
.A(n_3017),
.Y(n_3587)
);

INVx1_ASAP7_75t_L g3588 ( 
.A(n_3238),
.Y(n_3588)
);

AOI21x1_ASAP7_75t_L g3589 ( 
.A1(n_3240),
.A2(n_364),
.B(n_363),
.Y(n_3589)
);

AOI22xp5_ASAP7_75t_L g3590 ( 
.A1(n_3053),
.A2(n_326),
.B1(n_324),
.B2(n_325),
.Y(n_3590)
);

OAI22xp5_ASAP7_75t_L g3591 ( 
.A1(n_2976),
.A2(n_326),
.B1(n_324),
.B2(n_325),
.Y(n_3591)
);

AOI21xp5_ASAP7_75t_L g3592 ( 
.A1(n_3005),
.A2(n_324),
.B(n_325),
.Y(n_3592)
);

NAND2xp5_ASAP7_75t_L g3593 ( 
.A(n_2974),
.B(n_326),
.Y(n_3593)
);

INVx3_ASAP7_75t_L g3594 ( 
.A(n_2958),
.Y(n_3594)
);

INVx2_ASAP7_75t_L g3595 ( 
.A(n_3011),
.Y(n_3595)
);

INVx1_ASAP7_75t_L g3596 ( 
.A(n_2973),
.Y(n_3596)
);

A2O1A1Ixp33_ASAP7_75t_L g3597 ( 
.A1(n_3328),
.A2(n_3330),
.B(n_2995),
.C(n_3014),
.Y(n_3597)
);

INVx1_ASAP7_75t_L g3598 ( 
.A(n_2975),
.Y(n_3598)
);

INVx1_ASAP7_75t_L g3599 ( 
.A(n_3028),
.Y(n_3599)
);

HB1xp67_ASAP7_75t_L g3600 ( 
.A(n_3024),
.Y(n_3600)
);

AND2x2_ASAP7_75t_L g3601 ( 
.A(n_3280),
.B(n_327),
.Y(n_3601)
);

CKINVDCx5p33_ASAP7_75t_R g3602 ( 
.A(n_3009),
.Y(n_3602)
);

INVx8_ASAP7_75t_L g3603 ( 
.A(n_2958),
.Y(n_3603)
);

NAND2xp33_ASAP7_75t_L g3604 ( 
.A(n_2964),
.B(n_327),
.Y(n_3604)
);

OAI21xp5_ASAP7_75t_L g3605 ( 
.A1(n_3288),
.A2(n_327),
.B(n_328),
.Y(n_3605)
);

OAI21xp5_ASAP7_75t_L g3606 ( 
.A1(n_2959),
.A2(n_328),
.B(n_329),
.Y(n_3606)
);

OAI21x1_ASAP7_75t_L g3607 ( 
.A1(n_3022),
.A2(n_3253),
.B(n_3041),
.Y(n_3607)
);

NAND2x1p5_ASAP7_75t_L g3608 ( 
.A(n_2964),
.B(n_328),
.Y(n_3608)
);

BUFx2_ASAP7_75t_L g3609 ( 
.A(n_3021),
.Y(n_3609)
);

BUFx10_ASAP7_75t_L g3610 ( 
.A(n_3321),
.Y(n_3610)
);

INVx1_ASAP7_75t_SL g3611 ( 
.A(n_3009),
.Y(n_3611)
);

AND2x2_ASAP7_75t_L g3612 ( 
.A(n_3118),
.B(n_329),
.Y(n_3612)
);

AOI21xp5_ASAP7_75t_L g3613 ( 
.A1(n_3012),
.A2(n_330),
.B(n_331),
.Y(n_3613)
);

OAI21x1_ASAP7_75t_L g3614 ( 
.A1(n_3257),
.A2(n_334),
.B(n_333),
.Y(n_3614)
);

BUFx6f_ASAP7_75t_L g3615 ( 
.A(n_3012),
.Y(n_3615)
);

AO31x2_ASAP7_75t_L g3616 ( 
.A1(n_3291),
.A2(n_335),
.A3(n_332),
.B(n_333),
.Y(n_3616)
);

NAND2xp5_ASAP7_75t_L g3617 ( 
.A(n_3142),
.B(n_332),
.Y(n_3617)
);

AOI21x1_ASAP7_75t_SL g3618 ( 
.A1(n_3140),
.A2(n_332),
.B(n_333),
.Y(n_3618)
);

AOI21xp5_ASAP7_75t_L g3619 ( 
.A1(n_3012),
.A2(n_335),
.B(n_336),
.Y(n_3619)
);

NAND2xp5_ASAP7_75t_L g3620 ( 
.A(n_3155),
.B(n_335),
.Y(n_3620)
);

INVx1_ASAP7_75t_L g3621 ( 
.A(n_3037),
.Y(n_3621)
);

AOI21xp5_ASAP7_75t_L g3622 ( 
.A1(n_3019),
.A2(n_336),
.B(n_337),
.Y(n_3622)
);

OAI21xp5_ASAP7_75t_L g3623 ( 
.A1(n_2946),
.A2(n_337),
.B(n_338),
.Y(n_3623)
);

AND2x2_ASAP7_75t_L g3624 ( 
.A(n_3187),
.B(n_3080),
.Y(n_3624)
);

INVx1_ASAP7_75t_L g3625 ( 
.A(n_3039),
.Y(n_3625)
);

BUFx10_ASAP7_75t_L g3626 ( 
.A(n_3305),
.Y(n_3626)
);

NOR2xp33_ASAP7_75t_L g3627 ( 
.A(n_3214),
.B(n_337),
.Y(n_3627)
);

INVx2_ASAP7_75t_SL g3628 ( 
.A(n_3077),
.Y(n_3628)
);

OR2x2_ASAP7_75t_L g3629 ( 
.A(n_3056),
.B(n_338),
.Y(n_3629)
);

AOI21xp5_ASAP7_75t_L g3630 ( 
.A1(n_3019),
.A2(n_339),
.B(n_340),
.Y(n_3630)
);

AOI21xp5_ASAP7_75t_SL g3631 ( 
.A1(n_3337),
.A2(n_339),
.B(n_340),
.Y(n_3631)
);

NAND2xp5_ASAP7_75t_L g3632 ( 
.A(n_3269),
.B(n_340),
.Y(n_3632)
);

OR2x2_ASAP7_75t_L g3633 ( 
.A(n_2928),
.B(n_363),
.Y(n_3633)
);

CKINVDCx11_ASAP7_75t_R g3634 ( 
.A(n_3249),
.Y(n_3634)
);

OAI22xp5_ASAP7_75t_L g3635 ( 
.A1(n_3085),
.A2(n_366),
.B1(n_364),
.B2(n_365),
.Y(n_3635)
);

OAI21x1_ASAP7_75t_L g3636 ( 
.A1(n_3259),
.A2(n_365),
.B(n_366),
.Y(n_3636)
);

OAI21x1_ASAP7_75t_L g3637 ( 
.A1(n_3278),
.A2(n_369),
.B(n_370),
.Y(n_3637)
);

OA21x2_ASAP7_75t_L g3638 ( 
.A1(n_2982),
.A2(n_2984),
.B(n_3023),
.Y(n_3638)
);

OAI21xp5_ASAP7_75t_L g3639 ( 
.A1(n_2945),
.A2(n_369),
.B(n_370),
.Y(n_3639)
);

INVx1_ASAP7_75t_L g3640 ( 
.A(n_3040),
.Y(n_3640)
);

INVx1_ASAP7_75t_L g3641 ( 
.A(n_3049),
.Y(n_3641)
);

O2A1O1Ixp5_ASAP7_75t_L g3642 ( 
.A1(n_3136),
.A2(n_374),
.B(n_371),
.C(n_373),
.Y(n_3642)
);

BUFx10_ASAP7_75t_L g3643 ( 
.A(n_2979),
.Y(n_3643)
);

AOI21xp5_ASAP7_75t_L g3644 ( 
.A1(n_3019),
.A2(n_371),
.B(n_373),
.Y(n_3644)
);

OR2x2_ASAP7_75t_L g3645 ( 
.A(n_2912),
.B(n_375),
.Y(n_3645)
);

INVx6_ASAP7_75t_L g3646 ( 
.A(n_3339),
.Y(n_3646)
);

BUFx8_ASAP7_75t_L g3647 ( 
.A(n_3154),
.Y(n_3647)
);

INVx1_ASAP7_75t_L g3648 ( 
.A(n_2918),
.Y(n_3648)
);

NAND2xp5_ASAP7_75t_L g3649 ( 
.A(n_2962),
.B(n_375),
.Y(n_3649)
);

OAI21x1_ASAP7_75t_L g3650 ( 
.A1(n_3287),
.A2(n_376),
.B(n_377),
.Y(n_3650)
);

NAND2xp5_ASAP7_75t_L g3651 ( 
.A(n_3221),
.B(n_376),
.Y(n_3651)
);

INVx2_ASAP7_75t_L g3652 ( 
.A(n_3289),
.Y(n_3652)
);

AND2x2_ASAP7_75t_L g3653 ( 
.A(n_3114),
.B(n_378),
.Y(n_3653)
);

INVxp67_ASAP7_75t_SL g3654 ( 
.A(n_3315),
.Y(n_3654)
);

OAI21x1_ASAP7_75t_L g3655 ( 
.A1(n_3301),
.A2(n_378),
.B(n_379),
.Y(n_3655)
);

CKINVDCx11_ASAP7_75t_R g3656 ( 
.A(n_3219),
.Y(n_3656)
);

NAND2xp5_ASAP7_75t_L g3657 ( 
.A(n_3181),
.B(n_379),
.Y(n_3657)
);

OAI21x1_ASAP7_75t_SL g3658 ( 
.A1(n_3027),
.A2(n_851),
.B(n_850),
.Y(n_3658)
);

BUFx12f_ASAP7_75t_L g3659 ( 
.A(n_3260),
.Y(n_3659)
);

OA21x2_ASAP7_75t_L g3660 ( 
.A1(n_2994),
.A2(n_380),
.B(n_382),
.Y(n_3660)
);

AOI21xp5_ASAP7_75t_L g3661 ( 
.A1(n_3131),
.A2(n_380),
.B(n_382),
.Y(n_3661)
);

OAI22xp5_ASAP7_75t_L g3662 ( 
.A1(n_3122),
.A2(n_387),
.B1(n_384),
.B2(n_385),
.Y(n_3662)
);

INVxp67_ASAP7_75t_L g3663 ( 
.A(n_3170),
.Y(n_3663)
);

OR2x2_ASAP7_75t_L g3664 ( 
.A(n_3231),
.B(n_385),
.Y(n_3664)
);

OAI21x1_ASAP7_75t_L g3665 ( 
.A1(n_3346),
.A2(n_388),
.B(n_389),
.Y(n_3665)
);

AND2x2_ASAP7_75t_L g3666 ( 
.A(n_3327),
.B(n_388),
.Y(n_3666)
);

BUFx10_ASAP7_75t_L g3667 ( 
.A(n_3213),
.Y(n_3667)
);

NAND2xp5_ASAP7_75t_L g3668 ( 
.A(n_3191),
.B(n_389),
.Y(n_3668)
);

OAI22x1_ASAP7_75t_L g3669 ( 
.A1(n_3203),
.A2(n_392),
.B1(n_390),
.B2(n_391),
.Y(n_3669)
);

NAND2xp5_ASAP7_75t_SL g3670 ( 
.A(n_3240),
.B(n_390),
.Y(n_3670)
);

AO31x2_ASAP7_75t_L g3671 ( 
.A1(n_3117),
.A2(n_394),
.A3(n_392),
.B(n_393),
.Y(n_3671)
);

AO31x2_ASAP7_75t_L g3672 ( 
.A1(n_3153),
.A2(n_397),
.A3(n_395),
.B(n_396),
.Y(n_3672)
);

OAI21x1_ASAP7_75t_L g3673 ( 
.A1(n_3290),
.A2(n_398),
.B(n_399),
.Y(n_3673)
);

NAND2xp33_ASAP7_75t_L g3674 ( 
.A(n_3021),
.B(n_859),
.Y(n_3674)
);

AO32x2_ASAP7_75t_L g3675 ( 
.A1(n_3003),
.A2(n_400),
.A3(n_398),
.B1(n_399),
.B2(n_402),
.Y(n_3675)
);

INVxp67_ASAP7_75t_L g3676 ( 
.A(n_3050),
.Y(n_3676)
);

OAI21x1_ASAP7_75t_L g3677 ( 
.A1(n_3276),
.A2(n_403),
.B(n_405),
.Y(n_3677)
);

INVx1_ASAP7_75t_L g3678 ( 
.A(n_3086),
.Y(n_3678)
);

NAND2xp5_ASAP7_75t_L g3679 ( 
.A(n_2931),
.B(n_403),
.Y(n_3679)
);

CKINVDCx11_ASAP7_75t_R g3680 ( 
.A(n_3194),
.Y(n_3680)
);

INVx3_ASAP7_75t_L g3681 ( 
.A(n_3339),
.Y(n_3681)
);

CKINVDCx20_ASAP7_75t_R g3682 ( 
.A(n_3200),
.Y(n_3682)
);

AOI21xp5_ASAP7_75t_L g3683 ( 
.A1(n_3131),
.A2(n_405),
.B(n_406),
.Y(n_3683)
);

AO32x2_ASAP7_75t_L g3684 ( 
.A1(n_3004),
.A2(n_410),
.A3(n_408),
.B1(n_409),
.B2(n_411),
.Y(n_3684)
);

INVx1_ASAP7_75t_L g3685 ( 
.A(n_3093),
.Y(n_3685)
);

AND2x4_ASAP7_75t_L g3686 ( 
.A(n_3338),
.B(n_409),
.Y(n_3686)
);

A2O1A1Ixp33_ASAP7_75t_L g3687 ( 
.A1(n_3330),
.A2(n_413),
.B(n_411),
.C(n_412),
.Y(n_3687)
);

NAND2x1p5_ASAP7_75t_L g3688 ( 
.A(n_3244),
.B(n_858),
.Y(n_3688)
);

NOR2xp33_ASAP7_75t_L g3689 ( 
.A(n_3077),
.B(n_412),
.Y(n_3689)
);

AO21x1_ASAP7_75t_L g3690 ( 
.A1(n_3038),
.A2(n_413),
.B(n_414),
.Y(n_3690)
);

AOI21x1_ASAP7_75t_L g3691 ( 
.A1(n_3220),
.A2(n_415),
.B(n_416),
.Y(n_3691)
);

OR2x2_ASAP7_75t_L g3692 ( 
.A(n_3167),
.B(n_415),
.Y(n_3692)
);

NAND2xp5_ASAP7_75t_L g3693 ( 
.A(n_2942),
.B(n_858),
.Y(n_3693)
);

NAND2xp5_ASAP7_75t_L g3694 ( 
.A(n_2965),
.B(n_416),
.Y(n_3694)
);

INVx3_ASAP7_75t_SL g3695 ( 
.A(n_2943),
.Y(n_3695)
);

AOI22xp33_ASAP7_75t_L g3696 ( 
.A1(n_2924),
.A2(n_3326),
.B1(n_3348),
.B2(n_2944),
.Y(n_3696)
);

OAI21x1_ASAP7_75t_L g3697 ( 
.A1(n_3347),
.A2(n_417),
.B(n_418),
.Y(n_3697)
);

O2A1O1Ixp5_ASAP7_75t_SL g3698 ( 
.A1(n_3258),
.A2(n_421),
.B(n_419),
.C(n_420),
.Y(n_3698)
);

AND2x2_ASAP7_75t_L g3699 ( 
.A(n_2999),
.B(n_3013),
.Y(n_3699)
);

A2O1A1Ixp33_ASAP7_75t_L g3700 ( 
.A1(n_3100),
.A2(n_422),
.B(n_420),
.C(n_421),
.Y(n_3700)
);

AOI21x1_ASAP7_75t_L g3701 ( 
.A1(n_3264),
.A2(n_423),
.B(n_424),
.Y(n_3701)
);

AND2x2_ASAP7_75t_L g3702 ( 
.A(n_3295),
.B(n_424),
.Y(n_3702)
);

AND2x4_ASAP7_75t_L g3703 ( 
.A(n_3131),
.B(n_425),
.Y(n_3703)
);

NAND2xp5_ASAP7_75t_L g3704 ( 
.A(n_2971),
.B(n_3246),
.Y(n_3704)
);

A2O1A1Ixp33_ASAP7_75t_L g3705 ( 
.A1(n_3135),
.A2(n_427),
.B(n_425),
.C(n_426),
.Y(n_3705)
);

OAI21xp5_ASAP7_75t_L g3706 ( 
.A1(n_3314),
.A2(n_426),
.B(n_427),
.Y(n_3706)
);

A2O1A1Ixp33_ASAP7_75t_L g3707 ( 
.A1(n_3137),
.A2(n_430),
.B(n_428),
.C(n_429),
.Y(n_3707)
);

INVx3_ASAP7_75t_SL g3708 ( 
.A(n_2960),
.Y(n_3708)
);

NAND2xp5_ASAP7_75t_L g3709 ( 
.A(n_3234),
.B(n_857),
.Y(n_3709)
);

AOI21xp5_ASAP7_75t_L g3710 ( 
.A1(n_3150),
.A2(n_428),
.B(n_430),
.Y(n_3710)
);

OAI21xp5_ASAP7_75t_L g3711 ( 
.A1(n_3319),
.A2(n_432),
.B(n_434),
.Y(n_3711)
);

NOR2xp67_ASAP7_75t_L g3712 ( 
.A(n_3188),
.B(n_432),
.Y(n_3712)
);

OAI21x1_ASAP7_75t_L g3713 ( 
.A1(n_2923),
.A2(n_434),
.B(n_435),
.Y(n_3713)
);

INVx1_ASAP7_75t_L g3714 ( 
.A(n_3094),
.Y(n_3714)
);

OAI21x1_ASAP7_75t_L g3715 ( 
.A1(n_2926),
.A2(n_3046),
.B(n_3036),
.Y(n_3715)
);

OAI21x1_ASAP7_75t_L g3716 ( 
.A1(n_3052),
.A2(n_436),
.B(n_437),
.Y(n_3716)
);

AOI21x1_ASAP7_75t_L g3717 ( 
.A1(n_3190),
.A2(n_436),
.B(n_438),
.Y(n_3717)
);

OAI21x1_ASAP7_75t_L g3718 ( 
.A1(n_3431),
.A2(n_3072),
.B(n_3057),
.Y(n_3718)
);

AOI22xp5_ASAP7_75t_L g3719 ( 
.A1(n_3386),
.A2(n_3250),
.B1(n_3185),
.B2(n_3102),
.Y(n_3719)
);

INVx1_ASAP7_75t_L g3720 ( 
.A(n_3376),
.Y(n_3720)
);

HB1xp67_ASAP7_75t_L g3721 ( 
.A(n_3600),
.Y(n_3721)
);

OAI21x1_ASAP7_75t_L g3722 ( 
.A1(n_3453),
.A2(n_3082),
.B(n_3078),
.Y(n_3722)
);

OAI21xp5_ASAP7_75t_L g3723 ( 
.A1(n_3358),
.A2(n_3020),
.B(n_3225),
.Y(n_3723)
);

BUFx6f_ASAP7_75t_L g3724 ( 
.A(n_3603),
.Y(n_3724)
);

BUFx8_ASAP7_75t_L g3725 ( 
.A(n_3362),
.Y(n_3725)
);

NAND2xp5_ASAP7_75t_L g3726 ( 
.A(n_3441),
.B(n_2967),
.Y(n_3726)
);

NOR2x1_ASAP7_75t_R g3727 ( 
.A(n_3502),
.B(n_3602),
.Y(n_3727)
);

OAI21x1_ASAP7_75t_L g3728 ( 
.A1(n_3387),
.A2(n_3108),
.B(n_3107),
.Y(n_3728)
);

A2O1A1Ixp33_ASAP7_75t_L g3729 ( 
.A1(n_3604),
.A2(n_3487),
.B(n_3352),
.C(n_3437),
.Y(n_3729)
);

AO21x2_ASAP7_75t_L g3730 ( 
.A1(n_3384),
.A2(n_3266),
.B(n_3201),
.Y(n_3730)
);

OAI22xp33_ASAP7_75t_L g3731 ( 
.A1(n_3379),
.A2(n_3079),
.B1(n_3349),
.B2(n_3320),
.Y(n_3731)
);

INVxp33_ASAP7_75t_L g3732 ( 
.A(n_3634),
.Y(n_3732)
);

OAI21x1_ASAP7_75t_L g3733 ( 
.A1(n_3465),
.A2(n_3134),
.B(n_3123),
.Y(n_3733)
);

INVx2_ASAP7_75t_L g3734 ( 
.A(n_3353),
.Y(n_3734)
);

OAI21x1_ASAP7_75t_L g3735 ( 
.A1(n_3366),
.A2(n_3151),
.B(n_3143),
.Y(n_3735)
);

INVx1_ASAP7_75t_L g3736 ( 
.A(n_3377),
.Y(n_3736)
);

OAI21x1_ASAP7_75t_L g3737 ( 
.A1(n_3515),
.A2(n_3380),
.B(n_3481),
.Y(n_3737)
);

OAI21x1_ASAP7_75t_L g3738 ( 
.A1(n_3396),
.A2(n_3161),
.B(n_3157),
.Y(n_3738)
);

INVx1_ASAP7_75t_L g3739 ( 
.A(n_3398),
.Y(n_3739)
);

INVx8_ASAP7_75t_L g3740 ( 
.A(n_3603),
.Y(n_3740)
);

OAI21x1_ASAP7_75t_L g3741 ( 
.A1(n_3521),
.A2(n_3175),
.B(n_3168),
.Y(n_3741)
);

INVx3_ASAP7_75t_L g3742 ( 
.A(n_3391),
.Y(n_3742)
);

O2A1O1Ixp33_ASAP7_75t_SL g3743 ( 
.A1(n_3550),
.A2(n_3070),
.B(n_3169),
.C(n_3165),
.Y(n_3743)
);

OAI21xp5_ASAP7_75t_L g3744 ( 
.A1(n_3397),
.A2(n_3152),
.B(n_3342),
.Y(n_3744)
);

OAI21x1_ASAP7_75t_SL g3745 ( 
.A1(n_3391),
.A2(n_3042),
.B(n_2916),
.Y(n_3745)
);

INVx1_ASAP7_75t_SL g3746 ( 
.A(n_3680),
.Y(n_3746)
);

INVx2_ASAP7_75t_L g3747 ( 
.A(n_3355),
.Y(n_3747)
);

INVx4_ASAP7_75t_L g3748 ( 
.A(n_3422),
.Y(n_3748)
);

INVxp67_ASAP7_75t_L g3749 ( 
.A(n_3401),
.Y(n_3749)
);

AOI22xp33_ASAP7_75t_SL g3750 ( 
.A1(n_3385),
.A2(n_3266),
.B1(n_3329),
.B2(n_3090),
.Y(n_3750)
);

OA21x2_ASAP7_75t_L g3751 ( 
.A1(n_3513),
.A2(n_2909),
.B(n_3186),
.Y(n_3751)
);

INVx1_ASAP7_75t_L g3752 ( 
.A(n_3399),
.Y(n_3752)
);

HB1xp67_ASAP7_75t_L g3753 ( 
.A(n_3587),
.Y(n_3753)
);

OAI21x1_ASAP7_75t_SL g3754 ( 
.A1(n_3690),
.A2(n_3422),
.B(n_3482),
.Y(n_3754)
);

INVx1_ASAP7_75t_L g3755 ( 
.A(n_3410),
.Y(n_3755)
);

BUFx4f_ASAP7_75t_SL g3756 ( 
.A(n_3364),
.Y(n_3756)
);

INVx5_ASAP7_75t_L g3757 ( 
.A(n_3502),
.Y(n_3757)
);

NAND2xp5_ASAP7_75t_L g3758 ( 
.A(n_3369),
.B(n_2952),
.Y(n_3758)
);

INVx2_ASAP7_75t_L g3759 ( 
.A(n_3367),
.Y(n_3759)
);

INVx2_ASAP7_75t_SL g3760 ( 
.A(n_3647),
.Y(n_3760)
);

INVx4_ASAP7_75t_L g3761 ( 
.A(n_3466),
.Y(n_3761)
);

OAI21x1_ASAP7_75t_L g3762 ( 
.A1(n_3518),
.A2(n_3207),
.B(n_3202),
.Y(n_3762)
);

INVx1_ASAP7_75t_L g3763 ( 
.A(n_3425),
.Y(n_3763)
);

OAI21x1_ASAP7_75t_L g3764 ( 
.A1(n_3415),
.A2(n_3334),
.B(n_3177),
.Y(n_3764)
);

OA21x2_ASAP7_75t_L g3765 ( 
.A1(n_3563),
.A2(n_3182),
.B(n_2956),
.Y(n_3765)
);

OAI21x1_ASAP7_75t_L g3766 ( 
.A1(n_3470),
.A2(n_3025),
.B(n_3263),
.Y(n_3766)
);

INVx1_ASAP7_75t_L g3767 ( 
.A(n_3451),
.Y(n_3767)
);

OAI21x1_ASAP7_75t_SL g3768 ( 
.A1(n_3520),
.A2(n_3237),
.B(n_3196),
.Y(n_3768)
);

AND2x2_ASAP7_75t_L g3769 ( 
.A(n_3381),
.B(n_3197),
.Y(n_3769)
);

BUFx3_ASAP7_75t_L g3770 ( 
.A(n_3647),
.Y(n_3770)
);

OAI21x1_ASAP7_75t_L g3771 ( 
.A1(n_3491),
.A2(n_3272),
.B(n_3267),
.Y(n_3771)
);

BUFx3_ASAP7_75t_L g3772 ( 
.A(n_3682),
.Y(n_3772)
);

INVxp67_ASAP7_75t_SL g3773 ( 
.A(n_3452),
.Y(n_3773)
);

INVx1_ASAP7_75t_L g3774 ( 
.A(n_3471),
.Y(n_3774)
);

A2O1A1Ixp33_ASAP7_75t_L g3775 ( 
.A1(n_3674),
.A2(n_2954),
.B(n_3125),
.C(n_3120),
.Y(n_3775)
);

INVx3_ASAP7_75t_L g3776 ( 
.A(n_3646),
.Y(n_3776)
);

BUFx10_ASAP7_75t_L g3777 ( 
.A(n_3547),
.Y(n_3777)
);

INVxp67_ASAP7_75t_SL g3778 ( 
.A(n_3525),
.Y(n_3778)
);

BUFx6f_ASAP7_75t_L g3779 ( 
.A(n_3389),
.Y(n_3779)
);

OAI21x1_ASAP7_75t_L g3780 ( 
.A1(n_3511),
.A2(n_3099),
.B(n_3095),
.Y(n_3780)
);

OAI22xp5_ASAP7_75t_L g3781 ( 
.A1(n_3597),
.A2(n_3179),
.B1(n_3300),
.B2(n_3199),
.Y(n_3781)
);

NAND2xp5_ASAP7_75t_L g3782 ( 
.A(n_3648),
.B(n_3224),
.Y(n_3782)
);

OAI222xp33_ASAP7_75t_L g3783 ( 
.A1(n_3544),
.A2(n_3109),
.B1(n_3299),
.B2(n_3307),
.C1(n_3252),
.C2(n_3241),
.Y(n_3783)
);

AOI21xp5_ASAP7_75t_SL g3784 ( 
.A1(n_3687),
.A2(n_2948),
.B(n_2933),
.Y(n_3784)
);

BUFx3_ASAP7_75t_L g3785 ( 
.A(n_3427),
.Y(n_3785)
);

OR2x6_ASAP7_75t_L g3786 ( 
.A(n_3480),
.B(n_3010),
.Y(n_3786)
);

O2A1O1Ixp33_ASAP7_75t_L g3787 ( 
.A1(n_3704),
.A2(n_3333),
.B(n_3316),
.C(n_2955),
.Y(n_3787)
);

INVx2_ASAP7_75t_L g3788 ( 
.A(n_3571),
.Y(n_3788)
);

O2A1O1Ixp33_ASAP7_75t_L g3789 ( 
.A1(n_3359),
.A2(n_3556),
.B(n_3483),
.C(n_3447),
.Y(n_3789)
);

OA21x2_ASAP7_75t_L g3790 ( 
.A1(n_3517),
.A2(n_3105),
.B(n_3104),
.Y(n_3790)
);

OAI21xp5_ASAP7_75t_L g3791 ( 
.A1(n_3421),
.A2(n_2910),
.B(n_3111),
.Y(n_3791)
);

OAI21x1_ASAP7_75t_L g3792 ( 
.A1(n_3361),
.A2(n_3162),
.B(n_3127),
.Y(n_3792)
);

AOI221xp5_ASAP7_75t_L g3793 ( 
.A1(n_3696),
.A2(n_3198),
.B1(n_3208),
.B2(n_3195),
.C(n_3293),
.Y(n_3793)
);

BUFx2_ASAP7_75t_R g3794 ( 
.A(n_3372),
.Y(n_3794)
);

OAI21x1_ASAP7_75t_L g3795 ( 
.A1(n_3454),
.A2(n_3193),
.B(n_3150),
.Y(n_3795)
);

INVx6_ASAP7_75t_L g3796 ( 
.A(n_3626),
.Y(n_3796)
);

AOI21xp5_ASAP7_75t_L g3797 ( 
.A1(n_3464),
.A2(n_3193),
.B(n_3150),
.Y(n_3797)
);

INVx2_ASAP7_75t_SL g3798 ( 
.A(n_3626),
.Y(n_3798)
);

INVx2_ASAP7_75t_SL g3799 ( 
.A(n_3667),
.Y(n_3799)
);

AO31x2_ASAP7_75t_L g3800 ( 
.A1(n_3426),
.A2(n_3192),
.A3(n_3261),
.B(n_3193),
.Y(n_3800)
);

OAI21x1_ASAP7_75t_L g3801 ( 
.A1(n_3458),
.A2(n_3292),
.B(n_3261),
.Y(n_3801)
);

INVx5_ASAP7_75t_L g3802 ( 
.A(n_3667),
.Y(n_3802)
);

INVx5_ASAP7_75t_L g3803 ( 
.A(n_3646),
.Y(n_3803)
);

OA21x2_ASAP7_75t_L g3804 ( 
.A1(n_3488),
.A2(n_3192),
.B(n_3298),
.Y(n_3804)
);

HB1xp67_ASAP7_75t_L g3805 ( 
.A(n_3432),
.Y(n_3805)
);

INVx1_ASAP7_75t_L g3806 ( 
.A(n_3477),
.Y(n_3806)
);

NAND2x1p5_ASAP7_75t_L g3807 ( 
.A(n_3405),
.B(n_3261),
.Y(n_3807)
);

OAI21x1_ASAP7_75t_L g3808 ( 
.A1(n_3403),
.A2(n_3343),
.B(n_3292),
.Y(n_3808)
);

BUFx3_ASAP7_75t_L g3809 ( 
.A(n_3469),
.Y(n_3809)
);

INVx2_ASAP7_75t_L g3810 ( 
.A(n_3595),
.Y(n_3810)
);

INVx2_ASAP7_75t_L g3811 ( 
.A(n_3652),
.Y(n_3811)
);

A2O1A1Ixp33_ASAP7_75t_L g3812 ( 
.A1(n_3712),
.A2(n_3034),
.B(n_3343),
.C(n_3292),
.Y(n_3812)
);

INVx1_ASAP7_75t_L g3813 ( 
.A(n_3490),
.Y(n_3813)
);

INVx2_ASAP7_75t_SL g3814 ( 
.A(n_3610),
.Y(n_3814)
);

AOI221xp5_ASAP7_75t_L g3815 ( 
.A1(n_3593),
.A2(n_3354),
.B1(n_3591),
.B2(n_3627),
.C(n_3598),
.Y(n_3815)
);

NOR2xp33_ASAP7_75t_L g3816 ( 
.A(n_3611),
.B(n_3689),
.Y(n_3816)
);

AOI21xp5_ASAP7_75t_L g3817 ( 
.A1(n_3371),
.A2(n_3343),
.B(n_3192),
.Y(n_3817)
);

OA21x2_ASAP7_75t_L g3818 ( 
.A1(n_3467),
.A2(n_438),
.B(n_439),
.Y(n_3818)
);

AND2x2_ASAP7_75t_L g3819 ( 
.A(n_3540),
.B(n_856),
.Y(n_3819)
);

OAI21x1_ASAP7_75t_SL g3820 ( 
.A1(n_3542),
.A2(n_440),
.B(n_441),
.Y(n_3820)
);

AOI21x1_ASAP7_75t_L g3821 ( 
.A1(n_3496),
.A2(n_440),
.B(n_441),
.Y(n_3821)
);

AOI21xp5_ASAP7_75t_L g3822 ( 
.A1(n_3394),
.A2(n_442),
.B(n_443),
.Y(n_3822)
);

INVx1_ASAP7_75t_L g3823 ( 
.A(n_3501),
.Y(n_3823)
);

NAND2x1p5_ASAP7_75t_L g3824 ( 
.A(n_3486),
.B(n_3554),
.Y(n_3824)
);

BUFx6f_ASAP7_75t_L g3825 ( 
.A(n_3389),
.Y(n_3825)
);

OR2x6_ASAP7_75t_L g3826 ( 
.A(n_3628),
.B(n_442),
.Y(n_3826)
);

OAI21xp5_ASAP7_75t_L g3827 ( 
.A1(n_3642),
.A2(n_443),
.B(n_444),
.Y(n_3827)
);

AOI22xp33_ASAP7_75t_L g3828 ( 
.A1(n_3414),
.A2(n_447),
.B1(n_444),
.B2(n_446),
.Y(n_3828)
);

OAI21x1_ASAP7_75t_L g3829 ( 
.A1(n_3409),
.A2(n_3468),
.B(n_3570),
.Y(n_3829)
);

AND2x4_ASAP7_75t_L g3830 ( 
.A(n_3436),
.B(n_446),
.Y(n_3830)
);

INVx2_ASAP7_75t_L g3831 ( 
.A(n_3383),
.Y(n_3831)
);

BUFx10_ASAP7_75t_L g3832 ( 
.A(n_3686),
.Y(n_3832)
);

OAI21x1_ASAP7_75t_L g3833 ( 
.A1(n_3475),
.A2(n_3400),
.B(n_3618),
.Y(n_3833)
);

INVx1_ASAP7_75t_L g3834 ( 
.A(n_3523),
.Y(n_3834)
);

AND2x2_ASAP7_75t_L g3835 ( 
.A(n_3479),
.B(n_856),
.Y(n_3835)
);

OAI21xp5_ASAP7_75t_L g3836 ( 
.A1(n_3529),
.A2(n_447),
.B(n_448),
.Y(n_3836)
);

OAI21x1_ASAP7_75t_L g3837 ( 
.A1(n_3402),
.A2(n_448),
.B(n_449),
.Y(n_3837)
);

AOI22xp33_ASAP7_75t_L g3838 ( 
.A1(n_3699),
.A2(n_452),
.B1(n_450),
.B2(n_451),
.Y(n_3838)
);

AOI21x1_ASAP7_75t_L g3839 ( 
.A1(n_3462),
.A2(n_450),
.B(n_453),
.Y(n_3839)
);

AO21x2_ASAP7_75t_L g3840 ( 
.A1(n_3416),
.A2(n_453),
.B(n_454),
.Y(n_3840)
);

AO21x2_ASAP7_75t_L g3841 ( 
.A1(n_3670),
.A2(n_454),
.B(n_455),
.Y(n_3841)
);

OA21x2_ASAP7_75t_L g3842 ( 
.A1(n_3506),
.A2(n_455),
.B(n_457),
.Y(n_3842)
);

CKINVDCx16_ASAP7_75t_R g3843 ( 
.A(n_3370),
.Y(n_3843)
);

AOI21x1_ASAP7_75t_L g3844 ( 
.A1(n_3582),
.A2(n_457),
.B(n_458),
.Y(n_3844)
);

INVx2_ASAP7_75t_L g3845 ( 
.A(n_3392),
.Y(n_3845)
);

INVx1_ASAP7_75t_L g3846 ( 
.A(n_3534),
.Y(n_3846)
);

OAI21x1_ASAP7_75t_L g3847 ( 
.A1(n_3424),
.A2(n_458),
.B(n_459),
.Y(n_3847)
);

INVx1_ASAP7_75t_L g3848 ( 
.A(n_3551),
.Y(n_3848)
);

OAI22xp5_ASAP7_75t_L g3849 ( 
.A1(n_3522),
.A2(n_461),
.B1(n_459),
.B2(n_460),
.Y(n_3849)
);

OAI21x1_ASAP7_75t_L g3850 ( 
.A1(n_3715),
.A2(n_460),
.B(n_461),
.Y(n_3850)
);

BUFx2_ASAP7_75t_L g3851 ( 
.A(n_3478),
.Y(n_3851)
);

AOI21xp5_ASAP7_75t_L g3852 ( 
.A1(n_3493),
.A2(n_3374),
.B(n_3360),
.Y(n_3852)
);

OAI21x1_ASAP7_75t_L g3853 ( 
.A1(n_3476),
.A2(n_462),
.B(n_463),
.Y(n_3853)
);

OAI21xp5_ASAP7_75t_L g3854 ( 
.A1(n_3700),
.A2(n_855),
.B(n_463),
.Y(n_3854)
);

BUFx3_ASAP7_75t_L g3855 ( 
.A(n_3656),
.Y(n_3855)
);

INVxp67_ASAP7_75t_SL g3856 ( 
.A(n_3654),
.Y(n_3856)
);

AND2x4_ASAP7_75t_L g3857 ( 
.A(n_3373),
.B(n_464),
.Y(n_3857)
);

OAI21x1_ASAP7_75t_L g3858 ( 
.A1(n_3607),
.A2(n_464),
.B(n_465),
.Y(n_3858)
);

OAI21x1_ASAP7_75t_L g3859 ( 
.A1(n_3510),
.A2(n_3637),
.B(n_3636),
.Y(n_3859)
);

OAI21x1_ASAP7_75t_L g3860 ( 
.A1(n_3650),
.A2(n_465),
.B(n_466),
.Y(n_3860)
);

NOR2xp33_ASAP7_75t_L g3861 ( 
.A(n_3663),
.B(n_466),
.Y(n_3861)
);

AO21x2_ASAP7_75t_L g3862 ( 
.A1(n_3499),
.A2(n_467),
.B(n_468),
.Y(n_3862)
);

OAI21xp5_ASAP7_75t_L g3863 ( 
.A1(n_3705),
.A2(n_855),
.B(n_467),
.Y(n_3863)
);

O2A1O1Ixp5_ASAP7_75t_L g3864 ( 
.A1(n_3365),
.A2(n_470),
.B(n_468),
.C(n_469),
.Y(n_3864)
);

INVx1_ASAP7_75t_L g3865 ( 
.A(n_3557),
.Y(n_3865)
);

OAI21x1_ASAP7_75t_L g3866 ( 
.A1(n_3655),
.A2(n_469),
.B(n_470),
.Y(n_3866)
);

INVx2_ASAP7_75t_L g3867 ( 
.A(n_3412),
.Y(n_3867)
);

OAI21x1_ASAP7_75t_L g3868 ( 
.A1(n_3665),
.A2(n_471),
.B(n_472),
.Y(n_3868)
);

OAI21x1_ASAP7_75t_L g3869 ( 
.A1(n_3614),
.A2(n_471),
.B(n_472),
.Y(n_3869)
);

OAI21x1_ASAP7_75t_L g3870 ( 
.A1(n_3484),
.A2(n_473),
.B(n_474),
.Y(n_3870)
);

INVx1_ASAP7_75t_SL g3871 ( 
.A(n_3564),
.Y(n_3871)
);

OAI21xp5_ASAP7_75t_L g3872 ( 
.A1(n_3707),
.A2(n_854),
.B(n_473),
.Y(n_3872)
);

AO31x2_ASAP7_75t_L g3873 ( 
.A1(n_3417),
.A2(n_477),
.A3(n_475),
.B(n_476),
.Y(n_3873)
);

NOR2xp33_ASAP7_75t_L g3874 ( 
.A(n_3676),
.B(n_475),
.Y(n_3874)
);

OAI21xp33_ASAP7_75t_L g3875 ( 
.A1(n_3532),
.A2(n_476),
.B(n_477),
.Y(n_3875)
);

OAI21x1_ASAP7_75t_L g3876 ( 
.A1(n_3565),
.A2(n_478),
.B(n_479),
.Y(n_3876)
);

OAI21x1_ASAP7_75t_SL g3877 ( 
.A1(n_3706),
.A2(n_480),
.B(n_482),
.Y(n_3877)
);

OA21x2_ASAP7_75t_L g3878 ( 
.A1(n_3516),
.A2(n_480),
.B(n_483),
.Y(n_3878)
);

INVx1_ASAP7_75t_L g3879 ( 
.A(n_3531),
.Y(n_3879)
);

NAND3xp33_ASAP7_75t_L g3880 ( 
.A(n_3536),
.B(n_483),
.C(n_485),
.Y(n_3880)
);

INVxp67_ASAP7_75t_L g3881 ( 
.A(n_3583),
.Y(n_3881)
);

NOR2xp33_ASAP7_75t_L g3882 ( 
.A(n_3473),
.B(n_485),
.Y(n_3882)
);

NOR2xp67_ASAP7_75t_L g3883 ( 
.A(n_3507),
.B(n_486),
.Y(n_3883)
);

AOI22xp33_ASAP7_75t_L g3884 ( 
.A1(n_3624),
.A2(n_491),
.B1(n_487),
.B2(n_488),
.Y(n_3884)
);

AO31x2_ASAP7_75t_L g3885 ( 
.A1(n_3413),
.A2(n_3375),
.A3(n_3388),
.B(n_3526),
.Y(n_3885)
);

OAI21x1_ASAP7_75t_L g3886 ( 
.A1(n_3589),
.A2(n_493),
.B(n_494),
.Y(n_3886)
);

INVx2_ASAP7_75t_L g3887 ( 
.A(n_3461),
.Y(n_3887)
);

INVx2_ASAP7_75t_SL g3888 ( 
.A(n_3610),
.Y(n_3888)
);

HB1xp67_ASAP7_75t_L g3889 ( 
.A(n_3395),
.Y(n_3889)
);

OAI22xp5_ASAP7_75t_L g3890 ( 
.A1(n_3590),
.A2(n_3498),
.B1(n_3478),
.B2(n_3538),
.Y(n_3890)
);

INVx2_ASAP7_75t_L g3891 ( 
.A(n_3485),
.Y(n_3891)
);

AOI22xp33_ASAP7_75t_SL g3892 ( 
.A1(n_3368),
.A2(n_495),
.B1(n_493),
.B2(n_494),
.Y(n_3892)
);

INVx1_ASAP7_75t_L g3893 ( 
.A(n_3443),
.Y(n_3893)
);

INVx1_ASAP7_75t_L g3894 ( 
.A(n_3443),
.Y(n_3894)
);

INVx1_ASAP7_75t_L g3895 ( 
.A(n_3443),
.Y(n_3895)
);

INVx1_ASAP7_75t_L g3896 ( 
.A(n_3393),
.Y(n_3896)
);

INVx2_ASAP7_75t_L g3897 ( 
.A(n_3497),
.Y(n_3897)
);

INVx5_ASAP7_75t_L g3898 ( 
.A(n_3507),
.Y(n_3898)
);

INVx6_ASAP7_75t_L g3899 ( 
.A(n_3486),
.Y(n_3899)
);

OAI21x1_ASAP7_75t_L g3900 ( 
.A1(n_3514),
.A2(n_495),
.B(n_496),
.Y(n_3900)
);

INVx3_ASAP7_75t_L g3901 ( 
.A(n_3430),
.Y(n_3901)
);

OA21x2_ASAP7_75t_L g3902 ( 
.A1(n_3390),
.A2(n_496),
.B(n_497),
.Y(n_3902)
);

INVx2_ASAP7_75t_L g3903 ( 
.A(n_3560),
.Y(n_3903)
);

CKINVDCx20_ASAP7_75t_R g3904 ( 
.A(n_3500),
.Y(n_3904)
);

OA21x2_ASAP7_75t_L g3905 ( 
.A1(n_3677),
.A2(n_497),
.B(n_498),
.Y(n_3905)
);

AO21x2_ASAP7_75t_L g3906 ( 
.A1(n_3524),
.A2(n_499),
.B(n_500),
.Y(n_3906)
);

HB1xp67_ASAP7_75t_L g3907 ( 
.A(n_3460),
.Y(n_3907)
);

HB1xp67_ASAP7_75t_L g3908 ( 
.A(n_3492),
.Y(n_3908)
);

AO21x1_ASAP7_75t_L g3909 ( 
.A1(n_3528),
.A2(n_499),
.B(n_501),
.Y(n_3909)
);

OAI21x1_ASAP7_75t_L g3910 ( 
.A1(n_3508),
.A2(n_501),
.B(n_502),
.Y(n_3910)
);

BUFx3_ASAP7_75t_L g3911 ( 
.A(n_3463),
.Y(n_3911)
);

BUFx2_ASAP7_75t_L g3912 ( 
.A(n_3504),
.Y(n_3912)
);

BUFx4f_ASAP7_75t_L g3913 ( 
.A(n_3585),
.Y(n_3913)
);

NAND2xp5_ASAP7_75t_L g3914 ( 
.A(n_3406),
.B(n_502),
.Y(n_3914)
);

OAI21x1_ASAP7_75t_L g3915 ( 
.A1(n_3508),
.A2(n_503),
.B(n_505),
.Y(n_3915)
);

INVx1_ASAP7_75t_L g3916 ( 
.A(n_3393),
.Y(n_3916)
);

NOR2xp33_ASAP7_75t_L g3917 ( 
.A(n_3695),
.B(n_503),
.Y(n_3917)
);

BUFx2_ASAP7_75t_SL g3918 ( 
.A(n_3486),
.Y(n_3918)
);

BUFx2_ASAP7_75t_L g3919 ( 
.A(n_3609),
.Y(n_3919)
);

INVx2_ASAP7_75t_L g3920 ( 
.A(n_3568),
.Y(n_3920)
);

INVx4_ASAP7_75t_L g3921 ( 
.A(n_3554),
.Y(n_3921)
);

INVx4_ASAP7_75t_L g3922 ( 
.A(n_3554),
.Y(n_3922)
);

INVx2_ASAP7_75t_SL g3923 ( 
.A(n_3446),
.Y(n_3923)
);

AND2x4_ASAP7_75t_L g3924 ( 
.A(n_3681),
.B(n_506),
.Y(n_3924)
);

INVx1_ASAP7_75t_L g3925 ( 
.A(n_3505),
.Y(n_3925)
);

AOI22xp33_ASAP7_75t_L g3926 ( 
.A1(n_3519),
.A2(n_509),
.B1(n_506),
.B2(n_507),
.Y(n_3926)
);

OAI21x1_ASAP7_75t_L g3927 ( 
.A1(n_3512),
.A2(n_507),
.B(n_510),
.Y(n_3927)
);

AO21x2_ASAP7_75t_L g3928 ( 
.A1(n_3639),
.A2(n_511),
.B(n_512),
.Y(n_3928)
);

OAI22xp33_ASAP7_75t_L g3929 ( 
.A1(n_3584),
.A2(n_514),
.B1(n_511),
.B2(n_513),
.Y(n_3929)
);

OAI21x1_ASAP7_75t_L g3930 ( 
.A1(n_3512),
.A2(n_514),
.B(n_515),
.Y(n_3930)
);

INVx8_ASAP7_75t_L g3931 ( 
.A(n_3528),
.Y(n_3931)
);

O2A1O1Ixp33_ASAP7_75t_SL g3932 ( 
.A1(n_3546),
.A2(n_3580),
.B(n_3428),
.C(n_3420),
.Y(n_3932)
);

AOI22xp33_ASAP7_75t_L g3933 ( 
.A1(n_3356),
.A2(n_518),
.B1(n_516),
.B2(n_517),
.Y(n_3933)
);

NOR2xp33_ASAP7_75t_L g3934 ( 
.A(n_3708),
.B(n_516),
.Y(n_3934)
);

INVx1_ASAP7_75t_L g3935 ( 
.A(n_3393),
.Y(n_3935)
);

CKINVDCx20_ASAP7_75t_R g3936 ( 
.A(n_3659),
.Y(n_3936)
);

CKINVDCx20_ASAP7_75t_R g3937 ( 
.A(n_3574),
.Y(n_3937)
);

OAI21x1_ASAP7_75t_L g3938 ( 
.A1(n_3698),
.A2(n_517),
.B(n_519),
.Y(n_3938)
);

OAI21x1_ASAP7_75t_L g3939 ( 
.A1(n_3697),
.A2(n_519),
.B(n_520),
.Y(n_3939)
);

OA21x2_ASAP7_75t_L g3940 ( 
.A1(n_3545),
.A2(n_522),
.B(n_523),
.Y(n_3940)
);

BUFx12f_ASAP7_75t_L g3941 ( 
.A(n_3643),
.Y(n_3941)
);

AND2x2_ASAP7_75t_L g3942 ( 
.A(n_3363),
.B(n_3612),
.Y(n_3942)
);

AO31x2_ASAP7_75t_L g3943 ( 
.A1(n_3577),
.A2(n_525),
.A3(n_523),
.B(n_524),
.Y(n_3943)
);

OAI22xp33_ASAP7_75t_L g3944 ( 
.A1(n_3608),
.A2(n_526),
.B1(n_524),
.B2(n_525),
.Y(n_3944)
);

NAND2xp5_ASAP7_75t_SL g3945 ( 
.A(n_3357),
.B(n_526),
.Y(n_3945)
);

OAI21x1_ASAP7_75t_L g3946 ( 
.A1(n_3673),
.A2(n_527),
.B(n_528),
.Y(n_3946)
);

AO21x2_ASAP7_75t_L g3947 ( 
.A1(n_3711),
.A2(n_527),
.B(n_528),
.Y(n_3947)
);

OAI21x1_ASAP7_75t_L g3948 ( 
.A1(n_3552),
.A2(n_529),
.B(n_530),
.Y(n_3948)
);

OA21x2_ASAP7_75t_L g3949 ( 
.A1(n_3434),
.A2(n_530),
.B(n_531),
.Y(n_3949)
);

A2O1A1Ixp33_ASAP7_75t_L g3950 ( 
.A1(n_3623),
.A2(n_534),
.B(n_532),
.C(n_533),
.Y(n_3950)
);

BUFx3_ASAP7_75t_L g3951 ( 
.A(n_3537),
.Y(n_3951)
);

INVx1_ASAP7_75t_L g3952 ( 
.A(n_3588),
.Y(n_3952)
);

OAI21x1_ASAP7_75t_L g3953 ( 
.A1(n_3474),
.A2(n_532),
.B(n_535),
.Y(n_3953)
);

OAI21x1_ASAP7_75t_SL g3954 ( 
.A1(n_3606),
.A2(n_535),
.B(n_536),
.Y(n_3954)
);

AOI22xp33_ASAP7_75t_L g3955 ( 
.A1(n_3561),
.A2(n_538),
.B1(n_536),
.B2(n_537),
.Y(n_3955)
);

BUFx12f_ASAP7_75t_L g3956 ( 
.A(n_3643),
.Y(n_3956)
);

AO21x2_ASAP7_75t_L g3957 ( 
.A1(n_3658),
.A2(n_537),
.B(n_538),
.Y(n_3957)
);

INVx3_ASAP7_75t_L g3958 ( 
.A(n_3418),
.Y(n_3958)
);

OAI21x1_ASAP7_75t_L g3959 ( 
.A1(n_3558),
.A2(n_539),
.B(n_540),
.Y(n_3959)
);

INVx1_ASAP7_75t_L g3960 ( 
.A(n_3671),
.Y(n_3960)
);

OR2x6_ASAP7_75t_L g3961 ( 
.A(n_3688),
.B(n_539),
.Y(n_3961)
);

AND2x2_ASAP7_75t_L g3962 ( 
.A(n_3601),
.B(n_854),
.Y(n_3962)
);

INVx2_ASAP7_75t_L g3963 ( 
.A(n_3509),
.Y(n_3963)
);

AOI22xp5_ASAP7_75t_L g3964 ( 
.A1(n_3444),
.A2(n_542),
.B1(n_540),
.B2(n_541),
.Y(n_3964)
);

INVx2_ASAP7_75t_L g3965 ( 
.A(n_3703),
.Y(n_3965)
);

INVx1_ASAP7_75t_L g3966 ( 
.A(n_3671),
.Y(n_3966)
);

AOI21xp33_ASAP7_75t_L g3967 ( 
.A1(n_3407),
.A2(n_541),
.B(n_542),
.Y(n_3967)
);

AO21x2_ASAP7_75t_L g3968 ( 
.A1(n_3572),
.A2(n_543),
.B(n_544),
.Y(n_3968)
);

NOR2xp33_ASAP7_75t_SL g3969 ( 
.A(n_3350),
.B(n_543),
.Y(n_3969)
);

INVx1_ASAP7_75t_L g3970 ( 
.A(n_3419),
.Y(n_3970)
);

OAI21x1_ASAP7_75t_L g3971 ( 
.A1(n_3713),
.A2(n_544),
.B(n_545),
.Y(n_3971)
);

BUFx6f_ASAP7_75t_L g3972 ( 
.A(n_3389),
.Y(n_3972)
);

AOI21x1_ASAP7_75t_L g3973 ( 
.A1(n_3691),
.A2(n_545),
.B(n_546),
.Y(n_3973)
);

AO21x2_ASAP7_75t_L g3974 ( 
.A1(n_3701),
.A2(n_3539),
.B(n_3455),
.Y(n_3974)
);

AND2x4_ASAP7_75t_L g3975 ( 
.A(n_3703),
.B(n_547),
.Y(n_3975)
);

OAI21x1_ASAP7_75t_SL g3976 ( 
.A1(n_3541),
.A2(n_548),
.B(n_549),
.Y(n_3976)
);

AO21x2_ASAP7_75t_L g3977 ( 
.A1(n_3448),
.A2(n_548),
.B(n_550),
.Y(n_3977)
);

AOI21x1_ASAP7_75t_L g3978 ( 
.A1(n_3717),
.A2(n_550),
.B(n_551),
.Y(n_3978)
);

AOI22xp33_ASAP7_75t_L g3979 ( 
.A1(n_3423),
.A2(n_554),
.B1(n_551),
.B2(n_553),
.Y(n_3979)
);

INVx1_ASAP7_75t_SL g3980 ( 
.A(n_3686),
.Y(n_3980)
);

OAI21x1_ASAP7_75t_L g3981 ( 
.A1(n_3576),
.A2(n_554),
.B(n_555),
.Y(n_3981)
);

OAI222xp33_ASAP7_75t_L g3982 ( 
.A1(n_3635),
.A2(n_557),
.B1(n_559),
.B2(n_555),
.C1(n_556),
.C2(n_558),
.Y(n_3982)
);

O2A1O1Ixp33_ASAP7_75t_L g3983 ( 
.A1(n_3553),
.A2(n_560),
.B(n_556),
.C(n_558),
.Y(n_3983)
);

NAND2x1p5_ASAP7_75t_L g3984 ( 
.A(n_3594),
.B(n_560),
.Y(n_3984)
);

OAI21x1_ASAP7_75t_L g3985 ( 
.A1(n_3638),
.A2(n_561),
.B(n_562),
.Y(n_3985)
);

A2O1A1Ixp33_ASAP7_75t_L g3986 ( 
.A1(n_3605),
.A2(n_564),
.B(n_562),
.C(n_563),
.Y(n_3986)
);

INVx1_ASAP7_75t_L g3987 ( 
.A(n_3438),
.Y(n_3987)
);

NAND2x1p5_ASAP7_75t_L g3988 ( 
.A(n_3408),
.B(n_565),
.Y(n_3988)
);

INVx2_ASAP7_75t_L g3989 ( 
.A(n_3596),
.Y(n_3989)
);

NOR2xp33_ASAP7_75t_L g3990 ( 
.A(n_3543),
.B(n_565),
.Y(n_3990)
);

OA21x2_ASAP7_75t_L g3991 ( 
.A1(n_3716),
.A2(n_566),
.B(n_567),
.Y(n_3991)
);

INVx2_ASAP7_75t_L g3992 ( 
.A(n_3599),
.Y(n_3992)
);

BUFx2_ASAP7_75t_SL g3993 ( 
.A(n_3408),
.Y(n_3993)
);

OA21x2_ASAP7_75t_L g3994 ( 
.A1(n_3456),
.A2(n_567),
.B(n_568),
.Y(n_3994)
);

AND2x2_ASAP7_75t_L g3995 ( 
.A(n_3555),
.B(n_569),
.Y(n_3995)
);

OAI21x1_ASAP7_75t_L g3996 ( 
.A1(n_3638),
.A2(n_569),
.B(n_570),
.Y(n_3996)
);

OAI21x1_ASAP7_75t_L g3997 ( 
.A1(n_3660),
.A2(n_570),
.B(n_571),
.Y(n_3997)
);

CKINVDCx20_ASAP7_75t_R g3998 ( 
.A(n_3489),
.Y(n_3998)
);

BUFx2_ASAP7_75t_L g3999 ( 
.A(n_3442),
.Y(n_3999)
);

OR2x6_ASAP7_75t_L g4000 ( 
.A(n_3669),
.B(n_571),
.Y(n_4000)
);

A2O1A1Ixp33_ASAP7_75t_L g4001 ( 
.A1(n_3535),
.A2(n_574),
.B(n_572),
.C(n_573),
.Y(n_4001)
);

OAI21xp5_ASAP7_75t_L g4002 ( 
.A1(n_3549),
.A2(n_572),
.B(n_573),
.Y(n_4002)
);

HB1xp67_ASAP7_75t_L g4003 ( 
.A(n_3459),
.Y(n_4003)
);

AOI22xp5_ASAP7_75t_L g4004 ( 
.A1(n_3666),
.A2(n_577),
.B1(n_575),
.B2(n_576),
.Y(n_4004)
);

OAI21x1_ASAP7_75t_L g4005 ( 
.A1(n_3660),
.A2(n_575),
.B(n_576),
.Y(n_4005)
);

BUFx2_ASAP7_75t_R g4006 ( 
.A(n_3351),
.Y(n_4006)
);

INVx1_ASAP7_75t_L g4007 ( 
.A(n_3671),
.Y(n_4007)
);

OAI21x1_ASAP7_75t_SL g4008 ( 
.A1(n_3651),
.A2(n_578),
.B(n_579),
.Y(n_4008)
);

OAI21x1_ASAP7_75t_L g4009 ( 
.A1(n_3495),
.A2(n_578),
.B(n_580),
.Y(n_4009)
);

AOI21xp5_ASAP7_75t_L g4010 ( 
.A1(n_3495),
.A2(n_3429),
.B(n_3450),
.Y(n_4010)
);

OAI22xp33_ASAP7_75t_L g4011 ( 
.A1(n_3440),
.A2(n_584),
.B1(n_582),
.B2(n_583),
.Y(n_4011)
);

NOR2xp33_ASAP7_75t_L g4012 ( 
.A(n_3548),
.B(n_582),
.Y(n_4012)
);

OAI22xp5_ASAP7_75t_L g4013 ( 
.A1(n_3530),
.A2(n_587),
.B1(n_583),
.B2(n_585),
.Y(n_4013)
);

BUFx3_ASAP7_75t_L g4014 ( 
.A(n_3408),
.Y(n_4014)
);

INVx1_ASAP7_75t_L g4015 ( 
.A(n_3672),
.Y(n_4015)
);

NOR2xp33_ASAP7_75t_L g4016 ( 
.A(n_3573),
.B(n_585),
.Y(n_4016)
);

CKINVDCx5p33_ASAP7_75t_R g4017 ( 
.A(n_3586),
.Y(n_4017)
);

OAI21x1_ASAP7_75t_L g4018 ( 
.A1(n_3562),
.A2(n_587),
.B(n_588),
.Y(n_4018)
);

INVx2_ASAP7_75t_L g4019 ( 
.A(n_3621),
.Y(n_4019)
);

INVx2_ASAP7_75t_L g4020 ( 
.A(n_3625),
.Y(n_4020)
);

AOI21xp5_ASAP7_75t_SL g4021 ( 
.A1(n_3729),
.A2(n_3662),
.B(n_3649),
.Y(n_4021)
);

OR2x2_ASAP7_75t_L g4022 ( 
.A(n_3753),
.B(n_3503),
.Y(n_4022)
);

INVx1_ASAP7_75t_L g4023 ( 
.A(n_3736),
.Y(n_4023)
);

AOI21x1_ASAP7_75t_SL g4024 ( 
.A1(n_3830),
.A2(n_3702),
.B(n_3620),
.Y(n_4024)
);

O2A1O1Ixp33_ASAP7_75t_L g4025 ( 
.A1(n_3849),
.A2(n_3641),
.B(n_3640),
.C(n_3439),
.Y(n_4025)
);

AOI21x1_ASAP7_75t_SL g4026 ( 
.A1(n_3830),
.A2(n_3632),
.B(n_3617),
.Y(n_4026)
);

HB1xp67_ASAP7_75t_L g4027 ( 
.A(n_3999),
.Y(n_4027)
);

AOI21x1_ASAP7_75t_SL g4028 ( 
.A1(n_3924),
.A2(n_3566),
.B(n_3653),
.Y(n_4028)
);

CKINVDCx5p33_ASAP7_75t_R g4029 ( 
.A(n_3725),
.Y(n_4029)
);

OAI22xp5_ASAP7_75t_L g4030 ( 
.A1(n_3719),
.A2(n_3449),
.B1(n_3378),
.B2(n_3631),
.Y(n_4030)
);

OR2x2_ASAP7_75t_L g4031 ( 
.A(n_3907),
.B(n_3629),
.Y(n_4031)
);

NAND2xp5_ASAP7_75t_L g4032 ( 
.A(n_4003),
.B(n_3678),
.Y(n_4032)
);

O2A1O1Ixp33_ASAP7_75t_L g4033 ( 
.A1(n_4000),
.A2(n_3714),
.B(n_3685),
.C(n_3657),
.Y(n_4033)
);

BUFx2_ASAP7_75t_L g4034 ( 
.A(n_3748),
.Y(n_4034)
);

AND2x2_ASAP7_75t_L g4035 ( 
.A(n_3942),
.B(n_3675),
.Y(n_4035)
);

BUFx12f_ASAP7_75t_L g4036 ( 
.A(n_3725),
.Y(n_4036)
);

O2A1O1Ixp33_ASAP7_75t_L g4037 ( 
.A1(n_4000),
.A2(n_3668),
.B(n_3664),
.C(n_3709),
.Y(n_4037)
);

OA21x2_ASAP7_75t_L g4038 ( 
.A1(n_4010),
.A2(n_3661),
.B(n_3644),
.Y(n_4038)
);

O2A1O1Ixp33_ASAP7_75t_L g4039 ( 
.A1(n_4011),
.A2(n_3633),
.B(n_3692),
.C(n_3679),
.Y(n_4039)
);

OAI22xp5_ASAP7_75t_L g4040 ( 
.A1(n_3748),
.A2(n_3382),
.B1(n_3411),
.B2(n_3645),
.Y(n_4040)
);

AND2x2_ASAP7_75t_L g4041 ( 
.A(n_3908),
.B(n_3675),
.Y(n_4041)
);

OR2x2_ASAP7_75t_L g4042 ( 
.A(n_3721),
.B(n_3527),
.Y(n_4042)
);

INVx2_ASAP7_75t_SL g4043 ( 
.A(n_3740),
.Y(n_4043)
);

NAND2xp5_ASAP7_75t_L g4044 ( 
.A(n_3970),
.B(n_3672),
.Y(n_4044)
);

NAND2xp5_ASAP7_75t_L g4045 ( 
.A(n_3987),
.B(n_3672),
.Y(n_4045)
);

HB1xp67_ASAP7_75t_L g4046 ( 
.A(n_3856),
.Y(n_4046)
);

INVx1_ASAP7_75t_L g4047 ( 
.A(n_3736),
.Y(n_4047)
);

INVx2_ASAP7_75t_L g4048 ( 
.A(n_3867),
.Y(n_4048)
);

O2A1O1Ixp33_ASAP7_75t_L g4049 ( 
.A1(n_4013),
.A2(n_3694),
.B(n_3693),
.C(n_3569),
.Y(n_4049)
);

CKINVDCx5p33_ASAP7_75t_R g4050 ( 
.A(n_3913),
.Y(n_4050)
);

NAND2xp5_ASAP7_75t_L g4051 ( 
.A(n_3989),
.B(n_3559),
.Y(n_4051)
);

INVx1_ASAP7_75t_L g4052 ( 
.A(n_3739),
.Y(n_4052)
);

AOI21xp5_ASAP7_75t_L g4053 ( 
.A1(n_3852),
.A2(n_3404),
.B(n_3435),
.Y(n_4053)
);

NAND2x1_ASAP7_75t_L g4054 ( 
.A(n_3761),
.B(n_3435),
.Y(n_4054)
);

AND2x4_ASAP7_75t_L g4055 ( 
.A(n_3912),
.B(n_3435),
.Y(n_4055)
);

CKINVDCx20_ASAP7_75t_R g4056 ( 
.A(n_3904),
.Y(n_4056)
);

AND2x2_ASAP7_75t_L g4057 ( 
.A(n_3889),
.B(n_3675),
.Y(n_4057)
);

AND2x2_ASAP7_75t_L g4058 ( 
.A(n_3769),
.B(n_3684),
.Y(n_4058)
);

OA21x2_ASAP7_75t_L g4059 ( 
.A1(n_3817),
.A2(n_3710),
.B(n_3683),
.Y(n_4059)
);

AND2x2_ASAP7_75t_L g4060 ( 
.A(n_3992),
.B(n_3684),
.Y(n_4060)
);

OAI22xp5_ASAP7_75t_L g4061 ( 
.A1(n_3750),
.A2(n_3575),
.B1(n_3592),
.B2(n_3579),
.Y(n_4061)
);

OR2x2_ASAP7_75t_L g4062 ( 
.A(n_3805),
.B(n_3616),
.Y(n_4062)
);

AND2x2_ASAP7_75t_L g4063 ( 
.A(n_4019),
.B(n_3684),
.Y(n_4063)
);

OAI22xp5_ASAP7_75t_SL g4064 ( 
.A1(n_3770),
.A2(n_3826),
.B1(n_3843),
.B2(n_3760),
.Y(n_4064)
);

NAND2xp5_ASAP7_75t_L g4065 ( 
.A(n_4020),
.B(n_3559),
.Y(n_4065)
);

OA21x2_ASAP7_75t_L g4066 ( 
.A1(n_3829),
.A2(n_3630),
.B(n_3619),
.Y(n_4066)
);

AOI21x1_ASAP7_75t_SL g4067 ( 
.A1(n_3924),
.A2(n_3445),
.B(n_3559),
.Y(n_4067)
);

BUFx3_ASAP7_75t_L g4068 ( 
.A(n_3740),
.Y(n_4068)
);

OA21x2_ASAP7_75t_L g4069 ( 
.A1(n_3833),
.A2(n_3622),
.B(n_3613),
.Y(n_4069)
);

OA21x2_ASAP7_75t_L g4070 ( 
.A1(n_3859),
.A2(n_3433),
.B(n_3457),
.Y(n_4070)
);

OAI22xp5_ASAP7_75t_L g4071 ( 
.A1(n_3961),
.A2(n_3472),
.B1(n_3567),
.B2(n_3533),
.Y(n_4071)
);

BUFx12f_ASAP7_75t_L g4072 ( 
.A(n_3777),
.Y(n_4072)
);

OR2x2_ASAP7_75t_L g4073 ( 
.A(n_3919),
.B(n_3739),
.Y(n_4073)
);

NOR2xp33_ASAP7_75t_R g4074 ( 
.A(n_3913),
.B(n_588),
.Y(n_4074)
);

O2A1O1Ixp33_ASAP7_75t_L g4075 ( 
.A1(n_3890),
.A2(n_3578),
.B(n_3616),
.C(n_3457),
.Y(n_4075)
);

NAND2xp5_ASAP7_75t_L g4076 ( 
.A(n_3963),
.B(n_3578),
.Y(n_4076)
);

NAND2xp5_ASAP7_75t_L g4077 ( 
.A(n_3925),
.B(n_3578),
.Y(n_4077)
);

A2O1A1Ixp33_ASAP7_75t_L g4078 ( 
.A1(n_3812),
.A2(n_3883),
.B(n_3875),
.C(n_3917),
.Y(n_4078)
);

O2A1O1Ixp5_ASAP7_75t_L g4079 ( 
.A1(n_3761),
.A2(n_3616),
.B(n_3445),
.C(n_3457),
.Y(n_4079)
);

OAI22xp5_ASAP7_75t_L g4080 ( 
.A1(n_3961),
.A2(n_3472),
.B1(n_3567),
.B2(n_3533),
.Y(n_4080)
);

OR2x2_ASAP7_75t_L g4081 ( 
.A(n_3752),
.B(n_3494),
.Y(n_4081)
);

OA21x2_ASAP7_75t_L g4082 ( 
.A1(n_3896),
.A2(n_3445),
.B(n_3494),
.Y(n_4082)
);

AOI21x1_ASAP7_75t_SL g4083 ( 
.A1(n_3857),
.A2(n_589),
.B(n_590),
.Y(n_4083)
);

AND2x4_ASAP7_75t_L g4084 ( 
.A(n_3773),
.B(n_3472),
.Y(n_4084)
);

AND2x2_ASAP7_75t_L g4085 ( 
.A(n_3819),
.B(n_3494),
.Y(n_4085)
);

NAND2xp5_ASAP7_75t_L g4086 ( 
.A(n_3887),
.B(n_3891),
.Y(n_4086)
);

INVx4_ASAP7_75t_L g4087 ( 
.A(n_3802),
.Y(n_4087)
);

OAI22xp5_ASAP7_75t_L g4088 ( 
.A1(n_3931),
.A2(n_3567),
.B1(n_3581),
.B2(n_3533),
.Y(n_4088)
);

INVx1_ASAP7_75t_SL g4089 ( 
.A(n_3809),
.Y(n_4089)
);

O2A1O1Ixp33_ASAP7_75t_L g4090 ( 
.A1(n_3929),
.A2(n_591),
.B(n_589),
.C(n_590),
.Y(n_4090)
);

AND2x4_ASAP7_75t_L g4091 ( 
.A(n_3778),
.B(n_3581),
.Y(n_4091)
);

AND2x2_ASAP7_75t_L g4092 ( 
.A(n_3897),
.B(n_3581),
.Y(n_4092)
);

OAI31xp33_ASAP7_75t_SL g4093 ( 
.A1(n_3980),
.A2(n_594),
.A3(n_591),
.B(n_592),
.Y(n_4093)
);

NAND2xp5_ASAP7_75t_L g4094 ( 
.A(n_3903),
.B(n_3615),
.Y(n_4094)
);

AOI21x1_ASAP7_75t_SL g4095 ( 
.A1(n_3857),
.A2(n_3975),
.B(n_3914),
.Y(n_4095)
);

AND2x2_ASAP7_75t_L g4096 ( 
.A(n_3962),
.B(n_3615),
.Y(n_4096)
);

A2O1A1Ixp33_ASAP7_75t_L g4097 ( 
.A1(n_3934),
.A2(n_3615),
.B(n_595),
.C(n_592),
.Y(n_4097)
);

OA21x2_ASAP7_75t_L g4098 ( 
.A1(n_3896),
.A2(n_594),
.B(n_595),
.Y(n_4098)
);

AND2x4_ASAP7_75t_L g4099 ( 
.A(n_3802),
.B(n_596),
.Y(n_4099)
);

O2A1O1Ixp5_ASAP7_75t_L g4100 ( 
.A1(n_3909),
.A2(n_599),
.B(n_597),
.C(n_598),
.Y(n_4100)
);

AOI21xp5_ASAP7_75t_SL g4101 ( 
.A1(n_3975),
.A2(n_597),
.B(n_598),
.Y(n_4101)
);

INVxp67_ASAP7_75t_L g4102 ( 
.A(n_3799),
.Y(n_4102)
);

AND2x2_ASAP7_75t_L g4103 ( 
.A(n_3835),
.B(n_3720),
.Y(n_4103)
);

AOI21xp5_ASAP7_75t_SL g4104 ( 
.A1(n_3949),
.A2(n_599),
.B(n_600),
.Y(n_4104)
);

OAI22xp5_ASAP7_75t_L g4105 ( 
.A1(n_3931),
.A2(n_603),
.B1(n_601),
.B2(n_602),
.Y(n_4105)
);

INVx2_ASAP7_75t_L g4106 ( 
.A(n_3734),
.Y(n_4106)
);

OAI22xp5_ASAP7_75t_L g4107 ( 
.A1(n_3731),
.A2(n_605),
.B1(n_601),
.B2(n_603),
.Y(n_4107)
);

HB1xp67_ASAP7_75t_L g4108 ( 
.A(n_3749),
.Y(n_4108)
);

INVx1_ASAP7_75t_L g4109 ( 
.A(n_3752),
.Y(n_4109)
);

HB1xp67_ASAP7_75t_L g4110 ( 
.A(n_3881),
.Y(n_4110)
);

O2A1O1Ixp33_ASAP7_75t_L g4111 ( 
.A1(n_3944),
.A2(n_608),
.B(n_606),
.C(n_607),
.Y(n_4111)
);

OAI22xp5_ASAP7_75t_L g4112 ( 
.A1(n_4006),
.A2(n_610),
.B1(n_607),
.B2(n_609),
.Y(n_4112)
);

A2O1A1Ixp33_ASAP7_75t_SL g4113 ( 
.A1(n_4016),
.A2(n_612),
.B(n_610),
.C(n_611),
.Y(n_4113)
);

AOI21xp5_ASAP7_75t_L g4114 ( 
.A1(n_3797),
.A2(n_611),
.B(n_613),
.Y(n_4114)
);

HB1xp67_ASAP7_75t_L g4115 ( 
.A(n_3920),
.Y(n_4115)
);

NOR2xp33_ASAP7_75t_R g4116 ( 
.A(n_3756),
.B(n_614),
.Y(n_4116)
);

INVx1_ASAP7_75t_L g4117 ( 
.A(n_3763),
.Y(n_4117)
);

BUFx3_ASAP7_75t_L g4118 ( 
.A(n_3785),
.Y(n_4118)
);

O2A1O1Ixp5_ASAP7_75t_L g4119 ( 
.A1(n_3921),
.A2(n_618),
.B(n_615),
.C(n_617),
.Y(n_4119)
);

O2A1O1Ixp33_ASAP7_75t_L g4120 ( 
.A1(n_3982),
.A2(n_620),
.B(n_615),
.C(n_619),
.Y(n_4120)
);

INVx2_ASAP7_75t_SL g4121 ( 
.A(n_3802),
.Y(n_4121)
);

NOR2xp67_ASAP7_75t_L g4122 ( 
.A(n_3898),
.B(n_3757),
.Y(n_4122)
);

NAND2xp5_ASAP7_75t_L g4123 ( 
.A(n_3952),
.B(n_619),
.Y(n_4123)
);

OA21x2_ASAP7_75t_L g4124 ( 
.A1(n_3916),
.A2(n_3935),
.B(n_3894),
.Y(n_4124)
);

INVx1_ASAP7_75t_L g4125 ( 
.A(n_3763),
.Y(n_4125)
);

OAI22xp5_ASAP7_75t_L g4126 ( 
.A1(n_3826),
.A2(n_622),
.B1(n_620),
.B2(n_621),
.Y(n_4126)
);

O2A1O1Ixp33_ASAP7_75t_L g4127 ( 
.A1(n_3789),
.A2(n_624),
.B(n_622),
.C(n_623),
.Y(n_4127)
);

INVx2_ASAP7_75t_L g4128 ( 
.A(n_3747),
.Y(n_4128)
);

HB1xp67_ASAP7_75t_L g4129 ( 
.A(n_3831),
.Y(n_4129)
);

INVx1_ASAP7_75t_L g4130 ( 
.A(n_3767),
.Y(n_4130)
);

HB1xp67_ASAP7_75t_L g4131 ( 
.A(n_3845),
.Y(n_4131)
);

O2A1O1Ixp33_ASAP7_75t_L g4132 ( 
.A1(n_3882),
.A2(n_627),
.B(n_625),
.C(n_626),
.Y(n_4132)
);

OAI22xp5_ASAP7_75t_L g4133 ( 
.A1(n_3775),
.A2(n_628),
.B1(n_626),
.B2(n_627),
.Y(n_4133)
);

NAND2xp5_ASAP7_75t_L g4134 ( 
.A(n_3952),
.B(n_628),
.Y(n_4134)
);

HB1xp67_ASAP7_75t_L g4135 ( 
.A(n_3901),
.Y(n_4135)
);

AND2x4_ASAP7_75t_L g4136 ( 
.A(n_3803),
.B(n_629),
.Y(n_4136)
);

O2A1O1Ixp5_ASAP7_75t_L g4137 ( 
.A1(n_3921),
.A2(n_633),
.B(n_630),
.C(n_631),
.Y(n_4137)
);

AND2x4_ASAP7_75t_L g4138 ( 
.A(n_3803),
.B(n_630),
.Y(n_4138)
);

AOI21xp5_ASAP7_75t_SL g4139 ( 
.A1(n_3949),
.A2(n_3994),
.B(n_3878),
.Y(n_4139)
);

O2A1O1Ixp33_ASAP7_75t_L g4140 ( 
.A1(n_3983),
.A2(n_634),
.B(n_631),
.C(n_633),
.Y(n_4140)
);

HB1xp67_ASAP7_75t_L g4141 ( 
.A(n_3901),
.Y(n_4141)
);

OAI31xp33_ASAP7_75t_L g4142 ( 
.A1(n_3969),
.A2(n_636),
.A3(n_634),
.B(n_635),
.Y(n_4142)
);

AOI211xp5_ASAP7_75t_L g4143 ( 
.A1(n_3932),
.A2(n_637),
.B(n_635),
.C(n_636),
.Y(n_4143)
);

OA21x2_ASAP7_75t_L g4144 ( 
.A1(n_3916),
.A2(n_637),
.B(n_638),
.Y(n_4144)
);

CKINVDCx20_ASAP7_75t_R g4145 ( 
.A(n_3936),
.Y(n_4145)
);

HB1xp67_ASAP7_75t_L g4146 ( 
.A(n_3759),
.Y(n_4146)
);

AOI21xp5_ASAP7_75t_SL g4147 ( 
.A1(n_3994),
.A2(n_3878),
.B(n_3842),
.Y(n_4147)
);

AOI21x1_ASAP7_75t_SL g4148 ( 
.A1(n_3995),
.A2(n_638),
.B(n_639),
.Y(n_4148)
);

AND2x2_ASAP7_75t_L g4149 ( 
.A(n_3755),
.B(n_853),
.Y(n_4149)
);

O2A1O1Ixp33_ASAP7_75t_L g4150 ( 
.A1(n_3945),
.A2(n_643),
.B(n_641),
.C(n_642),
.Y(n_4150)
);

BUFx8_ASAP7_75t_L g4151 ( 
.A(n_3724),
.Y(n_4151)
);

AND2x2_ASAP7_75t_L g4152 ( 
.A(n_3834),
.B(n_641),
.Y(n_4152)
);

HB1xp67_ASAP7_75t_L g4153 ( 
.A(n_3788),
.Y(n_4153)
);

INVx1_ASAP7_75t_L g4154 ( 
.A(n_3767),
.Y(n_4154)
);

NOR2x1_ASAP7_75t_SL g4155 ( 
.A(n_3918),
.B(n_642),
.Y(n_4155)
);

A2O1A1Ixp33_ASAP7_75t_L g4156 ( 
.A1(n_3950),
.A2(n_646),
.B(n_644),
.C(n_645),
.Y(n_4156)
);

INVx1_ASAP7_75t_L g4157 ( 
.A(n_3774),
.Y(n_4157)
);

AND2x2_ASAP7_75t_L g4158 ( 
.A(n_3879),
.B(n_645),
.Y(n_4158)
);

OAI22xp5_ASAP7_75t_SL g4159 ( 
.A1(n_3732),
.A2(n_651),
.B1(n_649),
.B2(n_650),
.Y(n_4159)
);

AOI21x1_ASAP7_75t_SL g4160 ( 
.A1(n_3782),
.A2(n_649),
.B(n_651),
.Y(n_4160)
);

NAND2xp5_ASAP7_75t_L g4161 ( 
.A(n_3774),
.B(n_652),
.Y(n_4161)
);

AND2x2_ASAP7_75t_L g4162 ( 
.A(n_3806),
.B(n_652),
.Y(n_4162)
);

INVxp67_ASAP7_75t_L g4163 ( 
.A(n_3918),
.Y(n_4163)
);

NOR2xp67_ASAP7_75t_L g4164 ( 
.A(n_3898),
.B(n_653),
.Y(n_4164)
);

AOI21xp5_ASAP7_75t_L g4165 ( 
.A1(n_3790),
.A2(n_653),
.B(n_654),
.Y(n_4165)
);

AOI21x1_ASAP7_75t_SL g4166 ( 
.A1(n_3726),
.A2(n_3727),
.B(n_3758),
.Y(n_4166)
);

HB1xp67_ASAP7_75t_L g4167 ( 
.A(n_3810),
.Y(n_4167)
);

AOI21xp5_ASAP7_75t_L g4168 ( 
.A1(n_3790),
.A2(n_655),
.B(n_656),
.Y(n_4168)
);

NAND2xp5_ASAP7_75t_L g4169 ( 
.A(n_3806),
.B(n_655),
.Y(n_4169)
);

HB1xp67_ASAP7_75t_L g4170 ( 
.A(n_3811),
.Y(n_4170)
);

AOI21xp5_ASAP7_75t_L g4171 ( 
.A1(n_3784),
.A2(n_656),
.B(n_657),
.Y(n_4171)
);

NAND2xp5_ASAP7_75t_L g4172 ( 
.A(n_3813),
.B(n_657),
.Y(n_4172)
);

OAI22xp5_ASAP7_75t_L g4173 ( 
.A1(n_3926),
.A2(n_660),
.B1(n_658),
.B2(n_659),
.Y(n_4173)
);

AOI21x1_ASAP7_75t_SL g4174 ( 
.A1(n_3794),
.A2(n_659),
.B(n_661),
.Y(n_4174)
);

AND2x2_ASAP7_75t_L g4175 ( 
.A(n_3813),
.B(n_853),
.Y(n_4175)
);

OR2x2_ASAP7_75t_L g4176 ( 
.A(n_3823),
.B(n_661),
.Y(n_4176)
);

O2A1O1Ixp33_ASAP7_75t_L g4177 ( 
.A1(n_3986),
.A2(n_665),
.B(n_663),
.C(n_664),
.Y(n_4177)
);

AND2x2_ASAP7_75t_L g4178 ( 
.A(n_3823),
.B(n_666),
.Y(n_4178)
);

OAI22xp5_ASAP7_75t_L g4179 ( 
.A1(n_3892),
.A2(n_669),
.B1(n_666),
.B2(n_668),
.Y(n_4179)
);

A2O1A1Ixp33_ASAP7_75t_L g4180 ( 
.A1(n_3836),
.A2(n_671),
.B(n_669),
.C(n_670),
.Y(n_4180)
);

AND2x4_ASAP7_75t_L g4181 ( 
.A(n_3803),
.B(n_670),
.Y(n_4181)
);

O2A1O1Ixp5_ASAP7_75t_L g4182 ( 
.A1(n_3922),
.A2(n_673),
.B(n_671),
.C(n_672),
.Y(n_4182)
);

INVx2_ASAP7_75t_L g4183 ( 
.A(n_3846),
.Y(n_4183)
);

AOI221xp5_ASAP7_75t_L g4184 ( 
.A1(n_3815),
.A2(n_672),
.B1(n_673),
.B2(n_675),
.C(n_676),
.Y(n_4184)
);

HB1xp67_ASAP7_75t_L g4185 ( 
.A(n_3871),
.Y(n_4185)
);

AOI21xp5_ASAP7_75t_L g4186 ( 
.A1(n_3754),
.A2(n_675),
.B(n_676),
.Y(n_4186)
);

AOI21xp5_ASAP7_75t_L g4187 ( 
.A1(n_3768),
.A2(n_677),
.B(n_678),
.Y(n_4187)
);

NAND2xp5_ASAP7_75t_L g4188 ( 
.A(n_3846),
.B(n_678),
.Y(n_4188)
);

A2O1A1Ixp33_ASAP7_75t_L g4189 ( 
.A1(n_3880),
.A2(n_681),
.B(n_679),
.C(n_680),
.Y(n_4189)
);

INVx2_ASAP7_75t_L g4190 ( 
.A(n_3848),
.Y(n_4190)
);

AOI21x1_ASAP7_75t_SL g4191 ( 
.A1(n_3796),
.A2(n_681),
.B(n_682),
.Y(n_4191)
);

OR2x2_ASAP7_75t_L g4192 ( 
.A(n_3848),
.B(n_683),
.Y(n_4192)
);

OAI22xp5_ASAP7_75t_L g4193 ( 
.A1(n_3984),
.A2(n_4004),
.B1(n_3757),
.B2(n_3898),
.Y(n_4193)
);

OAI22xp5_ASAP7_75t_L g4194 ( 
.A1(n_3757),
.A2(n_686),
.B1(n_684),
.B2(n_685),
.Y(n_4194)
);

INVx2_ASAP7_75t_L g4195 ( 
.A(n_3865),
.Y(n_4195)
);

A2O1A1Ixp33_ASAP7_75t_L g4196 ( 
.A1(n_4002),
.A2(n_688),
.B(n_684),
.C(n_685),
.Y(n_4196)
);

NAND2xp5_ASAP7_75t_L g4197 ( 
.A(n_3865),
.B(n_688),
.Y(n_4197)
);

NAND2xp5_ASAP7_75t_L g4198 ( 
.A(n_3885),
.B(n_689),
.Y(n_4198)
);

AOI21xp5_ASAP7_75t_L g4199 ( 
.A1(n_3745),
.A2(n_3723),
.B(n_3791),
.Y(n_4199)
);

INVx1_ASAP7_75t_L g4200 ( 
.A(n_3943),
.Y(n_4200)
);

AND2x2_ASAP7_75t_L g4201 ( 
.A(n_3911),
.B(n_689),
.Y(n_4201)
);

BUFx3_ASAP7_75t_L g4202 ( 
.A(n_3724),
.Y(n_4202)
);

INVx1_ASAP7_75t_L g4203 ( 
.A(n_3943),
.Y(n_4203)
);

AND2x4_ASAP7_75t_L g4204 ( 
.A(n_3742),
.B(n_690),
.Y(n_4204)
);

INVx3_ASAP7_75t_L g4205 ( 
.A(n_3724),
.Y(n_4205)
);

INVxp67_ASAP7_75t_L g4206 ( 
.A(n_3923),
.Y(n_4206)
);

INVx1_ASAP7_75t_L g4207 ( 
.A(n_3943),
.Y(n_4207)
);

INVx1_ASAP7_75t_L g4208 ( 
.A(n_3960),
.Y(n_4208)
);

AND2x2_ASAP7_75t_L g4209 ( 
.A(n_3832),
.B(n_852),
.Y(n_4209)
);

AOI21xp5_ASAP7_75t_SL g4210 ( 
.A1(n_3842),
.A2(n_3922),
.B(n_3818),
.Y(n_4210)
);

AND2x2_ASAP7_75t_L g4211 ( 
.A(n_3832),
.B(n_852),
.Y(n_4211)
);

CKINVDCx20_ASAP7_75t_R g4212 ( 
.A(n_3855),
.Y(n_4212)
);

O2A1O1Ixp33_ASAP7_75t_L g4213 ( 
.A1(n_3787),
.A2(n_692),
.B(n_690),
.C(n_691),
.Y(n_4213)
);

AND2x4_ASAP7_75t_L g4214 ( 
.A(n_3742),
.B(n_691),
.Y(n_4214)
);

AND2x2_ASAP7_75t_L g4215 ( 
.A(n_3965),
.B(n_692),
.Y(n_4215)
);

AOI21xp5_ASAP7_75t_SL g4216 ( 
.A1(n_3818),
.A2(n_3940),
.B(n_3991),
.Y(n_4216)
);

BUFx10_ASAP7_75t_L g4217 ( 
.A(n_3796),
.Y(n_4217)
);

CKINVDCx20_ASAP7_75t_R g4218 ( 
.A(n_3772),
.Y(n_4218)
);

BUFx3_ASAP7_75t_L g4219 ( 
.A(n_3951),
.Y(n_4219)
);

AOI21xp5_ASAP7_75t_SL g4220 ( 
.A1(n_3940),
.A2(n_693),
.B(n_694),
.Y(n_4220)
);

AND2x2_ASAP7_75t_L g4221 ( 
.A(n_3885),
.B(n_694),
.Y(n_4221)
);

OA21x2_ASAP7_75t_L g4222 ( 
.A1(n_3935),
.A2(n_695),
.B(n_696),
.Y(n_4222)
);

INVx1_ASAP7_75t_SL g4223 ( 
.A(n_3899),
.Y(n_4223)
);

AOI21xp5_ASAP7_75t_SL g4224 ( 
.A1(n_3991),
.A2(n_3824),
.B(n_3902),
.Y(n_4224)
);

INVx5_ASAP7_75t_L g4225 ( 
.A(n_3899),
.Y(n_4225)
);

AOI21x1_ASAP7_75t_SL g4226 ( 
.A1(n_3941),
.A2(n_696),
.B(n_697),
.Y(n_4226)
);

NAND2xp5_ASAP7_75t_L g4227 ( 
.A(n_3885),
.B(n_698),
.Y(n_4227)
);

BUFx3_ASAP7_75t_L g4228 ( 
.A(n_4034),
.Y(n_4228)
);

OAI21x1_ASAP7_75t_L g4229 ( 
.A1(n_4079),
.A2(n_3996),
.B(n_3985),
.Y(n_4229)
);

INVx1_ASAP7_75t_L g4230 ( 
.A(n_4115),
.Y(n_4230)
);

INVx2_ASAP7_75t_L g4231 ( 
.A(n_4129),
.Y(n_4231)
);

INVx1_ASAP7_75t_L g4232 ( 
.A(n_4046),
.Y(n_4232)
);

OR2x6_ASAP7_75t_L g4233 ( 
.A(n_4210),
.B(n_3960),
.Y(n_4233)
);

INVx1_ASAP7_75t_L g4234 ( 
.A(n_4023),
.Y(n_4234)
);

AO21x2_ASAP7_75t_L g4235 ( 
.A1(n_4198),
.A2(n_3820),
.B(n_3966),
.Y(n_4235)
);

NAND2x1_ASAP7_75t_L g4236 ( 
.A(n_4087),
.B(n_3814),
.Y(n_4236)
);

INVx1_ASAP7_75t_L g4237 ( 
.A(n_4047),
.Y(n_4237)
);

OR2x2_ASAP7_75t_L g4238 ( 
.A(n_4027),
.B(n_3966),
.Y(n_4238)
);

INVx2_ASAP7_75t_L g4239 ( 
.A(n_4131),
.Y(n_4239)
);

AO21x2_ASAP7_75t_L g4240 ( 
.A1(n_4227),
.A2(n_4015),
.B(n_4007),
.Y(n_4240)
);

HB1xp67_ASAP7_75t_L g4241 ( 
.A(n_4146),
.Y(n_4241)
);

OAI21xp33_ASAP7_75t_L g4242 ( 
.A1(n_4093),
.A2(n_4015),
.B(n_4007),
.Y(n_4242)
);

INVx1_ASAP7_75t_L g4243 ( 
.A(n_4052),
.Y(n_4243)
);

CKINVDCx5p33_ASAP7_75t_R g4244 ( 
.A(n_4036),
.Y(n_4244)
);

OR2x6_ASAP7_75t_L g4245 ( 
.A(n_4224),
.B(n_3893),
.Y(n_4245)
);

AND2x2_ASAP7_75t_L g4246 ( 
.A(n_4103),
.B(n_3893),
.Y(n_4246)
);

AO21x2_ASAP7_75t_L g4247 ( 
.A1(n_4199),
.A2(n_3895),
.B(n_3894),
.Y(n_4247)
);

INVx2_ASAP7_75t_L g4248 ( 
.A(n_4124),
.Y(n_4248)
);

AO21x2_ASAP7_75t_L g4249 ( 
.A1(n_4221),
.A2(n_3895),
.B(n_4008),
.Y(n_4249)
);

INVx2_ASAP7_75t_SL g4250 ( 
.A(n_4151),
.Y(n_4250)
);

AND2x2_ASAP7_75t_L g4251 ( 
.A(n_4153),
.B(n_3851),
.Y(n_4251)
);

OR2x2_ASAP7_75t_L g4252 ( 
.A(n_4022),
.B(n_3746),
.Y(n_4252)
);

OAI21xp5_ASAP7_75t_L g4253 ( 
.A1(n_4119),
.A2(n_3864),
.B(n_3863),
.Y(n_4253)
);

INVx4_ASAP7_75t_SL g4254 ( 
.A(n_4064),
.Y(n_4254)
);

BUFx6f_ASAP7_75t_L g4255 ( 
.A(n_4054),
.Y(n_4255)
);

AND2x2_ASAP7_75t_L g4256 ( 
.A(n_4167),
.B(n_4014),
.Y(n_4256)
);

NAND2xp5_ASAP7_75t_L g4257 ( 
.A(n_4041),
.B(n_3800),
.Y(n_4257)
);

BUFx6f_ASAP7_75t_L g4258 ( 
.A(n_4087),
.Y(n_4258)
);

OA21x2_ASAP7_75t_L g4259 ( 
.A1(n_4053),
.A2(n_3737),
.B(n_3795),
.Y(n_4259)
);

INVx2_ASAP7_75t_L g4260 ( 
.A(n_4170),
.Y(n_4260)
);

AO21x2_ASAP7_75t_L g4261 ( 
.A1(n_4165),
.A2(n_3839),
.B(n_3877),
.Y(n_4261)
);

INVx1_ASAP7_75t_L g4262 ( 
.A(n_4109),
.Y(n_4262)
);

INVx1_ASAP7_75t_L g4263 ( 
.A(n_4117),
.Y(n_4263)
);

OA21x2_ASAP7_75t_L g4264 ( 
.A1(n_4200),
.A2(n_3801),
.B(n_3792),
.Y(n_4264)
);

INVx1_ASAP7_75t_L g4265 ( 
.A(n_4125),
.Y(n_4265)
);

HB1xp67_ASAP7_75t_L g4266 ( 
.A(n_4135),
.Y(n_4266)
);

HB1xp67_ASAP7_75t_L g4267 ( 
.A(n_4141),
.Y(n_4267)
);

AND2x2_ASAP7_75t_L g4268 ( 
.A(n_4096),
.B(n_3776),
.Y(n_4268)
);

HB1xp67_ASAP7_75t_L g4269 ( 
.A(n_4124),
.Y(n_4269)
);

INVx1_ASAP7_75t_L g4270 ( 
.A(n_4130),
.Y(n_4270)
);

INVx2_ASAP7_75t_L g4271 ( 
.A(n_4183),
.Y(n_4271)
);

OAI21x1_ASAP7_75t_L g4272 ( 
.A1(n_4067),
.A2(n_4216),
.B(n_4168),
.Y(n_4272)
);

AND2x2_ASAP7_75t_L g4273 ( 
.A(n_4185),
.B(n_3776),
.Y(n_4273)
);

NOR2xp33_ASAP7_75t_L g4274 ( 
.A(n_4033),
.B(n_3861),
.Y(n_4274)
);

OR2x6_ASAP7_75t_L g4275 ( 
.A(n_4122),
.B(n_3993),
.Y(n_4275)
);

BUFx3_ASAP7_75t_L g4276 ( 
.A(n_4118),
.Y(n_4276)
);

OR2x2_ASAP7_75t_L g4277 ( 
.A(n_4073),
.B(n_3873),
.Y(n_4277)
);

INVx2_ASAP7_75t_SL g4278 ( 
.A(n_4151),
.Y(n_4278)
);

INVx2_ASAP7_75t_L g4279 ( 
.A(n_4190),
.Y(n_4279)
);

AND2x2_ASAP7_75t_L g4280 ( 
.A(n_4108),
.B(n_3798),
.Y(n_4280)
);

INVx1_ASAP7_75t_L g4281 ( 
.A(n_4154),
.Y(n_4281)
);

AND2x2_ASAP7_75t_L g4282 ( 
.A(n_4110),
.B(n_4035),
.Y(n_4282)
);

OA21x2_ASAP7_75t_L g4283 ( 
.A1(n_4203),
.A2(n_3808),
.B(n_3910),
.Y(n_4283)
);

INVx1_ASAP7_75t_L g4284 ( 
.A(n_4157),
.Y(n_4284)
);

AND2x4_ASAP7_75t_L g4285 ( 
.A(n_4055),
.B(n_3800),
.Y(n_4285)
);

INVx2_ASAP7_75t_L g4286 ( 
.A(n_4195),
.Y(n_4286)
);

INVx2_ASAP7_75t_L g4287 ( 
.A(n_4208),
.Y(n_4287)
);

OR2x2_ASAP7_75t_L g4288 ( 
.A(n_4032),
.B(n_3873),
.Y(n_4288)
);

INVx1_ASAP7_75t_L g4289 ( 
.A(n_4086),
.Y(n_4289)
);

OA21x2_ASAP7_75t_L g4290 ( 
.A1(n_4207),
.A2(n_3927),
.B(n_3915),
.Y(n_4290)
);

INVx2_ASAP7_75t_L g4291 ( 
.A(n_4106),
.Y(n_4291)
);

OR2x2_ASAP7_75t_L g4292 ( 
.A(n_4031),
.B(n_3873),
.Y(n_4292)
);

OA21x2_ASAP7_75t_L g4293 ( 
.A1(n_4044),
.A2(n_3930),
.B(n_3997),
.Y(n_4293)
);

INVx2_ASAP7_75t_L g4294 ( 
.A(n_4128),
.Y(n_4294)
);

INVx1_ASAP7_75t_L g4295 ( 
.A(n_4048),
.Y(n_4295)
);

INVx1_ASAP7_75t_L g4296 ( 
.A(n_4042),
.Y(n_4296)
);

HB1xp67_ASAP7_75t_L g4297 ( 
.A(n_4084),
.Y(n_4297)
);

BUFx6f_ASAP7_75t_L g4298 ( 
.A(n_4225),
.Y(n_4298)
);

INVx2_ASAP7_75t_L g4299 ( 
.A(n_4081),
.Y(n_4299)
);

BUFx5_ASAP7_75t_L g4300 ( 
.A(n_4204),
.Y(n_4300)
);

INVx2_ASAP7_75t_L g4301 ( 
.A(n_4082),
.Y(n_4301)
);

INVx1_ASAP7_75t_L g4302 ( 
.A(n_4062),
.Y(n_4302)
);

BUFx3_ASAP7_75t_L g4303 ( 
.A(n_4202),
.Y(n_4303)
);

AND2x4_ASAP7_75t_L g4304 ( 
.A(n_4055),
.B(n_3800),
.Y(n_4304)
);

INVx2_ASAP7_75t_L g4305 ( 
.A(n_4082),
.Y(n_4305)
);

INVx3_ASAP7_75t_L g4306 ( 
.A(n_4084),
.Y(n_4306)
);

BUFx3_ASAP7_75t_L g4307 ( 
.A(n_4225),
.Y(n_4307)
);

NAND2xp5_ASAP7_75t_L g4308 ( 
.A(n_4057),
.B(n_4058),
.Y(n_4308)
);

INVx1_ASAP7_75t_L g4309 ( 
.A(n_4060),
.Y(n_4309)
);

INVxp67_ASAP7_75t_SL g4310 ( 
.A(n_4098),
.Y(n_4310)
);

BUFx2_ASAP7_75t_L g4311 ( 
.A(n_4163),
.Y(n_4311)
);

INVx1_ASAP7_75t_L g4312 ( 
.A(n_4063),
.Y(n_4312)
);

INVx1_ASAP7_75t_L g4313 ( 
.A(n_4051),
.Y(n_4313)
);

INVxp67_ASAP7_75t_L g4314 ( 
.A(n_4098),
.Y(n_4314)
);

INVx2_ASAP7_75t_SL g4315 ( 
.A(n_4217),
.Y(n_4315)
);

INVx1_ASAP7_75t_L g4316 ( 
.A(n_4065),
.Y(n_4316)
);

AND2x2_ASAP7_75t_L g4317 ( 
.A(n_4092),
.B(n_3888),
.Y(n_4317)
);

AO21x2_ASAP7_75t_L g4318 ( 
.A1(n_4139),
.A2(n_3976),
.B(n_3954),
.Y(n_4318)
);

INVx3_ASAP7_75t_L g4319 ( 
.A(n_4091),
.Y(n_4319)
);

AND2x2_ASAP7_75t_L g4320 ( 
.A(n_4085),
.B(n_3974),
.Y(n_4320)
);

AND2x2_ASAP7_75t_L g4321 ( 
.A(n_4206),
.B(n_3730),
.Y(n_4321)
);

INVx4_ASAP7_75t_L g4322 ( 
.A(n_4225),
.Y(n_4322)
);

INVx1_ASAP7_75t_L g4323 ( 
.A(n_4045),
.Y(n_4323)
);

AND2x2_ASAP7_75t_L g4324 ( 
.A(n_4091),
.B(n_3804),
.Y(n_4324)
);

INVx1_ASAP7_75t_L g4325 ( 
.A(n_4076),
.Y(n_4325)
);

INVx2_ASAP7_75t_L g4326 ( 
.A(n_4094),
.Y(n_4326)
);

INVx1_ASAP7_75t_L g4327 ( 
.A(n_4162),
.Y(n_4327)
);

INVx2_ASAP7_75t_L g4328 ( 
.A(n_4077),
.Y(n_4328)
);

INVx1_ASAP7_75t_L g4329 ( 
.A(n_4175),
.Y(n_4329)
);

AND2x2_ASAP7_75t_L g4330 ( 
.A(n_4282),
.B(n_4320),
.Y(n_4330)
);

OR2x2_ASAP7_75t_L g4331 ( 
.A(n_4308),
.B(n_4070),
.Y(n_4331)
);

NOR2x1_ASAP7_75t_L g4332 ( 
.A(n_4276),
.B(n_4219),
.Y(n_4332)
);

INVx2_ASAP7_75t_L g4333 ( 
.A(n_4248),
.Y(n_4333)
);

AND2x2_ASAP7_75t_L g4334 ( 
.A(n_4246),
.B(n_4070),
.Y(n_4334)
);

AND2x2_ASAP7_75t_L g4335 ( 
.A(n_4321),
.B(n_3804),
.Y(n_4335)
);

AND2x2_ASAP7_75t_L g4336 ( 
.A(n_4309),
.B(n_4038),
.Y(n_4336)
);

AND2x2_ASAP7_75t_L g4337 ( 
.A(n_4312),
.B(n_4038),
.Y(n_4337)
);

INVx2_ASAP7_75t_L g4338 ( 
.A(n_4248),
.Y(n_4338)
);

INVx2_ASAP7_75t_L g4339 ( 
.A(n_4287),
.Y(n_4339)
);

INVx2_ASAP7_75t_L g4340 ( 
.A(n_4287),
.Y(n_4340)
);

AND2x2_ASAP7_75t_L g4341 ( 
.A(n_4324),
.B(n_4059),
.Y(n_4341)
);

INVx2_ASAP7_75t_L g4342 ( 
.A(n_4271),
.Y(n_4342)
);

OR2x2_ASAP7_75t_L g4343 ( 
.A(n_4308),
.B(n_4089),
.Y(n_4343)
);

INVx1_ASAP7_75t_L g4344 ( 
.A(n_4269),
.Y(n_4344)
);

BUFx2_ASAP7_75t_L g4345 ( 
.A(n_4228),
.Y(n_4345)
);

INVx2_ASAP7_75t_L g4346 ( 
.A(n_4271),
.Y(n_4346)
);

INVx2_ASAP7_75t_L g4347 ( 
.A(n_4279),
.Y(n_4347)
);

INVx2_ASAP7_75t_L g4348 ( 
.A(n_4279),
.Y(n_4348)
);

AND2x2_ASAP7_75t_L g4349 ( 
.A(n_4328),
.B(n_4059),
.Y(n_4349)
);

INVx1_ASAP7_75t_L g4350 ( 
.A(n_4241),
.Y(n_4350)
);

AND2x2_ASAP7_75t_L g4351 ( 
.A(n_4328),
.B(n_4144),
.Y(n_4351)
);

INVx1_ASAP7_75t_L g4352 ( 
.A(n_4241),
.Y(n_4352)
);

INVx1_ASAP7_75t_L g4353 ( 
.A(n_4230),
.Y(n_4353)
);

INVxp67_ASAP7_75t_SL g4354 ( 
.A(n_4266),
.Y(n_4354)
);

AND2x2_ASAP7_75t_L g4355 ( 
.A(n_4323),
.B(n_4144),
.Y(n_4355)
);

AND2x2_ASAP7_75t_L g4356 ( 
.A(n_4299),
.B(n_4222),
.Y(n_4356)
);

INVxp67_ASAP7_75t_SL g4357 ( 
.A(n_4266),
.Y(n_4357)
);

INVx1_ASAP7_75t_L g4358 ( 
.A(n_4269),
.Y(n_4358)
);

OAI21xp5_ASAP7_75t_L g4359 ( 
.A1(n_4242),
.A2(n_4078),
.B(n_4101),
.Y(n_4359)
);

BUFx2_ASAP7_75t_L g4360 ( 
.A(n_4228),
.Y(n_4360)
);

INVx2_ASAP7_75t_SL g4361 ( 
.A(n_4276),
.Y(n_4361)
);

INVx2_ASAP7_75t_L g4362 ( 
.A(n_4286),
.Y(n_4362)
);

NOR2x1p5_ASAP7_75t_L g4363 ( 
.A(n_4236),
.B(n_4068),
.Y(n_4363)
);

INVx1_ASAP7_75t_L g4364 ( 
.A(n_4286),
.Y(n_4364)
);

AND2x2_ASAP7_75t_L g4365 ( 
.A(n_4299),
.B(n_4222),
.Y(n_4365)
);

AND2x2_ASAP7_75t_L g4366 ( 
.A(n_4313),
.B(n_4178),
.Y(n_4366)
);

AND2x2_ASAP7_75t_L g4367 ( 
.A(n_4316),
.B(n_4075),
.Y(n_4367)
);

AO31x2_ASAP7_75t_L g4368 ( 
.A1(n_4301),
.A2(n_4040),
.A3(n_4030),
.B(n_4071),
.Y(n_4368)
);

INVxp67_ASAP7_75t_L g4369 ( 
.A(n_4267),
.Y(n_4369)
);

OAI22xp5_ASAP7_75t_L g4370 ( 
.A1(n_4242),
.A2(n_4080),
.B1(n_4099),
.B2(n_4204),
.Y(n_4370)
);

INVx3_ASAP7_75t_L g4371 ( 
.A(n_4275),
.Y(n_4371)
);

INVx2_ASAP7_75t_L g4372 ( 
.A(n_4301),
.Y(n_4372)
);

NAND2xp5_ASAP7_75t_L g4373 ( 
.A(n_4302),
.B(n_4149),
.Y(n_4373)
);

AND2x4_ASAP7_75t_L g4374 ( 
.A(n_4285),
.B(n_4121),
.Y(n_4374)
);

INVx2_ASAP7_75t_L g4375 ( 
.A(n_4305),
.Y(n_4375)
);

INVx1_ASAP7_75t_L g4376 ( 
.A(n_4232),
.Y(n_4376)
);

INVx1_ASAP7_75t_L g4377 ( 
.A(n_4289),
.Y(n_4377)
);

INVx1_ASAP7_75t_L g4378 ( 
.A(n_4231),
.Y(n_4378)
);

INVx1_ASAP7_75t_L g4379 ( 
.A(n_4239),
.Y(n_4379)
);

AO31x2_ASAP7_75t_L g4380 ( 
.A1(n_4305),
.A2(n_4061),
.A3(n_4186),
.B(n_4187),
.Y(n_4380)
);

AND2x2_ASAP7_75t_L g4381 ( 
.A(n_4325),
.B(n_3862),
.Y(n_4381)
);

INVx2_ASAP7_75t_L g4382 ( 
.A(n_4291),
.Y(n_4382)
);

AND2x2_ASAP7_75t_L g4383 ( 
.A(n_4257),
.B(n_4069),
.Y(n_4383)
);

AND2x2_ASAP7_75t_L g4384 ( 
.A(n_4257),
.B(n_4069),
.Y(n_4384)
);

OR2x2_ASAP7_75t_L g4385 ( 
.A(n_4296),
.B(n_4102),
.Y(n_4385)
);

AND2x2_ASAP7_75t_L g4386 ( 
.A(n_4285),
.B(n_4147),
.Y(n_4386)
);

INVx1_ASAP7_75t_L g4387 ( 
.A(n_4234),
.Y(n_4387)
);

AND2x2_ASAP7_75t_L g4388 ( 
.A(n_4304),
.B(n_4066),
.Y(n_4388)
);

AND2x2_ASAP7_75t_L g4389 ( 
.A(n_4304),
.B(n_4066),
.Y(n_4389)
);

INVx2_ASAP7_75t_L g4390 ( 
.A(n_4294),
.Y(n_4390)
);

INVx2_ASAP7_75t_L g4391 ( 
.A(n_4295),
.Y(n_4391)
);

INVx1_ASAP7_75t_L g4392 ( 
.A(n_4260),
.Y(n_4392)
);

INVx1_ASAP7_75t_L g4393 ( 
.A(n_4237),
.Y(n_4393)
);

INVx1_ASAP7_75t_SL g4394 ( 
.A(n_4250),
.Y(n_4394)
);

HB1xp67_ASAP7_75t_L g4395 ( 
.A(n_4267),
.Y(n_4395)
);

CKINVDCx8_ASAP7_75t_R g4396 ( 
.A(n_4254),
.Y(n_4396)
);

BUFx2_ASAP7_75t_L g4397 ( 
.A(n_4275),
.Y(n_4397)
);

AND2x2_ASAP7_75t_L g4398 ( 
.A(n_4326),
.B(n_3902),
.Y(n_4398)
);

AOI22xp33_ASAP7_75t_SL g4399 ( 
.A1(n_4300),
.A2(n_4074),
.B1(n_4116),
.B2(n_4155),
.Y(n_4399)
);

AND2x2_ASAP7_75t_L g4400 ( 
.A(n_4297),
.B(n_4152),
.Y(n_4400)
);

INVx1_ASAP7_75t_L g4401 ( 
.A(n_4243),
.Y(n_4401)
);

AND2x2_ASAP7_75t_L g4402 ( 
.A(n_4297),
.B(n_4158),
.Y(n_4402)
);

INVx1_ASAP7_75t_L g4403 ( 
.A(n_4262),
.Y(n_4403)
);

NAND2xp5_ASAP7_75t_L g4404 ( 
.A(n_4292),
.B(n_4176),
.Y(n_4404)
);

NAND2xp5_ASAP7_75t_L g4405 ( 
.A(n_4288),
.B(n_4192),
.Y(n_4405)
);

HB1xp67_ASAP7_75t_L g4406 ( 
.A(n_4256),
.Y(n_4406)
);

AND2x2_ASAP7_75t_L g4407 ( 
.A(n_4247),
.B(n_3751),
.Y(n_4407)
);

OR2x2_ASAP7_75t_L g4408 ( 
.A(n_4343),
.B(n_4238),
.Y(n_4408)
);

AO21x2_ASAP7_75t_L g4409 ( 
.A1(n_4344),
.A2(n_4310),
.B(n_4314),
.Y(n_4409)
);

AOI221xp5_ASAP7_75t_L g4410 ( 
.A1(n_4359),
.A2(n_4274),
.B1(n_4107),
.B2(n_4126),
.C(n_4037),
.Y(n_4410)
);

HB1xp67_ASAP7_75t_L g4411 ( 
.A(n_4395),
.Y(n_4411)
);

INVx1_ASAP7_75t_L g4412 ( 
.A(n_4350),
.Y(n_4412)
);

INVxp67_ASAP7_75t_L g4413 ( 
.A(n_4345),
.Y(n_4413)
);

OR2x2_ASAP7_75t_L g4414 ( 
.A(n_4343),
.B(n_4277),
.Y(n_4414)
);

BUFx4f_ASAP7_75t_SL g4415 ( 
.A(n_4394),
.Y(n_4415)
);

INVx1_ASAP7_75t_L g4416 ( 
.A(n_4352),
.Y(n_4416)
);

HB1xp67_ASAP7_75t_L g4417 ( 
.A(n_4345),
.Y(n_4417)
);

INVx2_ASAP7_75t_L g4418 ( 
.A(n_4360),
.Y(n_4418)
);

OAI22xp5_ASAP7_75t_L g4419 ( 
.A1(n_4396),
.A2(n_4399),
.B1(n_4370),
.B2(n_4361),
.Y(n_4419)
);

INVx2_ASAP7_75t_L g4420 ( 
.A(n_4360),
.Y(n_4420)
);

INVx2_ASAP7_75t_L g4421 ( 
.A(n_4333),
.Y(n_4421)
);

INVx1_ASAP7_75t_L g4422 ( 
.A(n_4387),
.Y(n_4422)
);

INVx1_ASAP7_75t_L g4423 ( 
.A(n_4387),
.Y(n_4423)
);

INVx1_ASAP7_75t_L g4424 ( 
.A(n_4403),
.Y(n_4424)
);

OAI22xp33_ASAP7_75t_L g4425 ( 
.A1(n_4396),
.A2(n_4275),
.B1(n_4322),
.B2(n_4233),
.Y(n_4425)
);

AND2x2_ASAP7_75t_L g4426 ( 
.A(n_4330),
.B(n_4273),
.Y(n_4426)
);

INVx2_ASAP7_75t_L g4427 ( 
.A(n_4333),
.Y(n_4427)
);

HB1xp67_ASAP7_75t_L g4428 ( 
.A(n_4354),
.Y(n_4428)
);

AOI22xp33_ASAP7_75t_L g4429 ( 
.A1(n_4367),
.A2(n_4274),
.B1(n_4318),
.B2(n_4254),
.Y(n_4429)
);

INVx2_ASAP7_75t_L g4430 ( 
.A(n_4338),
.Y(n_4430)
);

INVx2_ASAP7_75t_L g4431 ( 
.A(n_4338),
.Y(n_4431)
);

OR2x6_ASAP7_75t_L g4432 ( 
.A(n_4363),
.B(n_4322),
.Y(n_4432)
);

NAND2xp5_ASAP7_75t_L g4433 ( 
.A(n_4367),
.B(n_4327),
.Y(n_4433)
);

AOI221xp5_ASAP7_75t_L g4434 ( 
.A1(n_4383),
.A2(n_4112),
.B1(n_4105),
.B2(n_4159),
.C(n_4133),
.Y(n_4434)
);

INVxp67_ASAP7_75t_SL g4435 ( 
.A(n_4357),
.Y(n_4435)
);

INVx2_ASAP7_75t_SL g4436 ( 
.A(n_4332),
.Y(n_4436)
);

OAI22xp33_ASAP7_75t_L g4437 ( 
.A1(n_4397),
.A2(n_4233),
.B1(n_4307),
.B2(n_4245),
.Y(n_4437)
);

AND2x2_ASAP7_75t_L g4438 ( 
.A(n_4330),
.B(n_4306),
.Y(n_4438)
);

AOI221xp5_ASAP7_75t_L g4439 ( 
.A1(n_4383),
.A2(n_4132),
.B1(n_4329),
.B2(n_3874),
.C(n_4311),
.Y(n_4439)
);

NOR4xp25_ASAP7_75t_SL g4440 ( 
.A(n_4397),
.B(n_4244),
.C(n_4029),
.D(n_4254),
.Y(n_4440)
);

OR2x2_ASAP7_75t_L g4441 ( 
.A(n_4331),
.B(n_4306),
.Y(n_4441)
);

NAND3xp33_ASAP7_75t_L g4442 ( 
.A(n_4344),
.B(n_4143),
.C(n_4142),
.Y(n_4442)
);

OR2x6_ASAP7_75t_L g4443 ( 
.A(n_4361),
.B(n_4371),
.Y(n_4443)
);

NAND3xp33_ASAP7_75t_L g4444 ( 
.A(n_4358),
.B(n_4171),
.C(n_4253),
.Y(n_4444)
);

BUFx3_ASAP7_75t_L g4445 ( 
.A(n_4406),
.Y(n_4445)
);

AO21x2_ASAP7_75t_L g4446 ( 
.A1(n_4358),
.A2(n_4310),
.B(n_4314),
.Y(n_4446)
);

AND2x2_ASAP7_75t_L g4447 ( 
.A(n_4374),
.B(n_4319),
.Y(n_4447)
);

NOR2xp33_ASAP7_75t_R g4448 ( 
.A(n_4371),
.B(n_4244),
.Y(n_4448)
);

OAI221xp5_ASAP7_75t_L g4449 ( 
.A1(n_4386),
.A2(n_4097),
.B1(n_4017),
.B2(n_4193),
.C(n_4315),
.Y(n_4449)
);

INVx1_ASAP7_75t_L g4450 ( 
.A(n_4403),
.Y(n_4450)
);

INVx1_ASAP7_75t_L g4451 ( 
.A(n_4377),
.Y(n_4451)
);

NAND2xp33_ASAP7_75t_R g4452 ( 
.A(n_4371),
.B(n_4050),
.Y(n_4452)
);

AND2x4_ASAP7_75t_L g4453 ( 
.A(n_4386),
.B(n_4245),
.Y(n_4453)
);

AND4x1_ASAP7_75t_L g4454 ( 
.A(n_4400),
.B(n_4201),
.C(n_4100),
.D(n_4209),
.Y(n_4454)
);

INVxp67_ASAP7_75t_SL g4455 ( 
.A(n_4369),
.Y(n_4455)
);

INVx2_ASAP7_75t_L g4456 ( 
.A(n_4372),
.Y(n_4456)
);

AND2x2_ASAP7_75t_L g4457 ( 
.A(n_4374),
.B(n_4319),
.Y(n_4457)
);

AND2x2_ASAP7_75t_L g4458 ( 
.A(n_4374),
.B(n_4251),
.Y(n_4458)
);

AOI222xp33_ASAP7_75t_SL g4459 ( 
.A1(n_4353),
.A2(n_4194),
.B1(n_4179),
.B2(n_3781),
.C1(n_4173),
.C2(n_4253),
.Y(n_4459)
);

OAI33xp33_ASAP7_75t_L g4460 ( 
.A1(n_4385),
.A2(n_4331),
.A3(n_4373),
.B1(n_4376),
.B2(n_4252),
.B3(n_4405),
.Y(n_4460)
);

AOI22xp33_ASAP7_75t_L g4461 ( 
.A1(n_4400),
.A2(n_4318),
.B1(n_4233),
.B2(n_4249),
.Y(n_4461)
);

INVx1_ASAP7_75t_L g4462 ( 
.A(n_4378),
.Y(n_4462)
);

NAND4xp25_ASAP7_75t_L g4463 ( 
.A(n_4385),
.B(n_3816),
.C(n_4039),
.D(n_4025),
.Y(n_4463)
);

AOI221xp5_ASAP7_75t_L g4464 ( 
.A1(n_4384),
.A2(n_4127),
.B1(n_4111),
.B2(n_4090),
.C(n_4213),
.Y(n_4464)
);

OA21x2_ASAP7_75t_L g4465 ( 
.A1(n_4341),
.A2(n_4272),
.B(n_4229),
.Y(n_4465)
);

INVx1_ASAP7_75t_L g4466 ( 
.A(n_4379),
.Y(n_4466)
);

NAND2xp5_ASAP7_75t_L g4467 ( 
.A(n_4384),
.B(n_4355),
.Y(n_4467)
);

AND2x2_ASAP7_75t_L g4468 ( 
.A(n_4402),
.B(n_4341),
.Y(n_4468)
);

CKINVDCx5p33_ASAP7_75t_R g4469 ( 
.A(n_4402),
.Y(n_4469)
);

INVxp67_ASAP7_75t_SL g4470 ( 
.A(n_4382),
.Y(n_4470)
);

AO21x2_ASAP7_75t_L g4471 ( 
.A1(n_4388),
.A2(n_4247),
.B(n_4169),
.Y(n_4471)
);

INVx1_ASAP7_75t_L g4472 ( 
.A(n_4392),
.Y(n_4472)
);

AO21x2_ASAP7_75t_L g4473 ( 
.A1(n_4388),
.A2(n_4172),
.B(n_4161),
.Y(n_4473)
);

INVx2_ASAP7_75t_L g4474 ( 
.A(n_4372),
.Y(n_4474)
);

INVx2_ASAP7_75t_L g4475 ( 
.A(n_4375),
.Y(n_4475)
);

INVx1_ASAP7_75t_L g4476 ( 
.A(n_4393),
.Y(n_4476)
);

INVx2_ASAP7_75t_L g4477 ( 
.A(n_4421),
.Y(n_4477)
);

NAND3xp33_ASAP7_75t_SL g4478 ( 
.A(n_4440),
.B(n_4212),
.C(n_4218),
.Y(n_4478)
);

HB1xp67_ASAP7_75t_L g4479 ( 
.A(n_4428),
.Y(n_4479)
);

NAND2xp5_ASAP7_75t_L g4480 ( 
.A(n_4473),
.B(n_4336),
.Y(n_4480)
);

INVx1_ASAP7_75t_L g4481 ( 
.A(n_4422),
.Y(n_4481)
);

INVx1_ASAP7_75t_L g4482 ( 
.A(n_4423),
.Y(n_4482)
);

INVx1_ASAP7_75t_L g4483 ( 
.A(n_4424),
.Y(n_4483)
);

NOR2xp33_ASAP7_75t_L g4484 ( 
.A(n_4415),
.B(n_4278),
.Y(n_4484)
);

INVx2_ASAP7_75t_L g4485 ( 
.A(n_4427),
.Y(n_4485)
);

INVxp67_ASAP7_75t_SL g4486 ( 
.A(n_4417),
.Y(n_4486)
);

INVx2_ASAP7_75t_L g4487 ( 
.A(n_4430),
.Y(n_4487)
);

INVx2_ASAP7_75t_L g4488 ( 
.A(n_4431),
.Y(n_4488)
);

NOR3xp33_ASAP7_75t_SL g4489 ( 
.A(n_4419),
.B(n_4196),
.C(n_3783),
.Y(n_4489)
);

INVx1_ASAP7_75t_L g4490 ( 
.A(n_4450),
.Y(n_4490)
);

INVx1_ASAP7_75t_L g4491 ( 
.A(n_4411),
.Y(n_4491)
);

INVx1_ASAP7_75t_L g4492 ( 
.A(n_4414),
.Y(n_4492)
);

BUFx3_ASAP7_75t_L g4493 ( 
.A(n_4432),
.Y(n_4493)
);

HB1xp67_ASAP7_75t_L g4494 ( 
.A(n_4435),
.Y(n_4494)
);

INVx2_ASAP7_75t_SL g4495 ( 
.A(n_4432),
.Y(n_4495)
);

INVx2_ASAP7_75t_L g4496 ( 
.A(n_4456),
.Y(n_4496)
);

INVx1_ASAP7_75t_L g4497 ( 
.A(n_4462),
.Y(n_4497)
);

INVx2_ASAP7_75t_L g4498 ( 
.A(n_4474),
.Y(n_4498)
);

OA21x2_ASAP7_75t_L g4499 ( 
.A1(n_4429),
.A2(n_4389),
.B(n_4349),
.Y(n_4499)
);

INVx2_ASAP7_75t_L g4500 ( 
.A(n_4475),
.Y(n_4500)
);

NAND2xp5_ASAP7_75t_SL g4501 ( 
.A(n_4419),
.B(n_4258),
.Y(n_4501)
);

AOI21xp5_ASAP7_75t_L g4502 ( 
.A1(n_4432),
.A2(n_4220),
.B(n_4104),
.Y(n_4502)
);

INVx1_ASAP7_75t_L g4503 ( 
.A(n_4409),
.Y(n_4503)
);

NAND2xp5_ASAP7_75t_L g4504 ( 
.A(n_4473),
.B(n_4336),
.Y(n_4504)
);

AND2x2_ASAP7_75t_L g4505 ( 
.A(n_4468),
.B(n_4438),
.Y(n_4505)
);

HB1xp67_ASAP7_75t_L g4506 ( 
.A(n_4445),
.Y(n_4506)
);

NOR3xp33_ASAP7_75t_L g4507 ( 
.A(n_4444),
.B(n_4182),
.C(n_4137),
.Y(n_4507)
);

BUFx8_ASAP7_75t_L g4508 ( 
.A(n_4436),
.Y(n_4508)
);

HB1xp67_ASAP7_75t_L g4509 ( 
.A(n_4413),
.Y(n_4509)
);

OA21x2_ASAP7_75t_L g4510 ( 
.A1(n_4461),
.A2(n_4389),
.B(n_4349),
.Y(n_4510)
);

OA21x2_ASAP7_75t_L g4511 ( 
.A1(n_4444),
.A2(n_4335),
.B(n_4375),
.Y(n_4511)
);

INVx1_ASAP7_75t_L g4512 ( 
.A(n_4466),
.Y(n_4512)
);

INVx1_ASAP7_75t_L g4513 ( 
.A(n_4472),
.Y(n_4513)
);

AOI21x1_ASAP7_75t_L g4514 ( 
.A1(n_4443),
.A2(n_4164),
.B(n_4043),
.Y(n_4514)
);

INVx2_ASAP7_75t_L g4515 ( 
.A(n_4409),
.Y(n_4515)
);

OA21x2_ASAP7_75t_L g4516 ( 
.A1(n_4418),
.A2(n_4335),
.B(n_4407),
.Y(n_4516)
);

AND2x4_ASAP7_75t_L g4517 ( 
.A(n_4453),
.B(n_4368),
.Y(n_4517)
);

INVx1_ASAP7_75t_L g4518 ( 
.A(n_4476),
.Y(n_4518)
);

INVx1_ASAP7_75t_L g4519 ( 
.A(n_4446),
.Y(n_4519)
);

INVx1_ASAP7_75t_L g4520 ( 
.A(n_4446),
.Y(n_4520)
);

INVx2_ASAP7_75t_L g4521 ( 
.A(n_4441),
.Y(n_4521)
);

OA21x2_ASAP7_75t_L g4522 ( 
.A1(n_4420),
.A2(n_4407),
.B(n_4337),
.Y(n_4522)
);

NAND2xp5_ASAP7_75t_SL g4523 ( 
.A(n_4501),
.B(n_4425),
.Y(n_4523)
);

NAND2xp5_ASAP7_75t_L g4524 ( 
.A(n_4494),
.B(n_4455),
.Y(n_4524)
);

AND2x2_ASAP7_75t_L g4525 ( 
.A(n_4495),
.B(n_4443),
.Y(n_4525)
);

INVx2_ASAP7_75t_L g4526 ( 
.A(n_4522),
.Y(n_4526)
);

INVx1_ASAP7_75t_L g4527 ( 
.A(n_4479),
.Y(n_4527)
);

OR2x2_ASAP7_75t_L g4528 ( 
.A(n_4480),
.B(n_4467),
.Y(n_4528)
);

NOR2xp67_ASAP7_75t_SL g4529 ( 
.A(n_4501),
.B(n_4072),
.Y(n_4529)
);

INVx1_ASAP7_75t_L g4530 ( 
.A(n_4509),
.Y(n_4530)
);

OR2x2_ASAP7_75t_L g4531 ( 
.A(n_4504),
.B(n_4433),
.Y(n_4531)
);

AND2x4_ASAP7_75t_L g4532 ( 
.A(n_4493),
.B(n_4495),
.Y(n_4532)
);

NAND2xp5_ASAP7_75t_L g4533 ( 
.A(n_4491),
.B(n_4337),
.Y(n_4533)
);

INVx1_ASAP7_75t_L g4534 ( 
.A(n_4486),
.Y(n_4534)
);

AND2x2_ASAP7_75t_L g4535 ( 
.A(n_4506),
.B(n_4443),
.Y(n_4535)
);

OR2x2_ASAP7_75t_L g4536 ( 
.A(n_4492),
.B(n_4408),
.Y(n_4536)
);

OAI221xp5_ASAP7_75t_L g4537 ( 
.A1(n_4489),
.A2(n_4410),
.B1(n_4463),
.B2(n_4439),
.C(n_4449),
.Y(n_4537)
);

AND2x2_ASAP7_75t_L g4538 ( 
.A(n_4493),
.B(n_4453),
.Y(n_4538)
);

INVx1_ASAP7_75t_L g4539 ( 
.A(n_4497),
.Y(n_4539)
);

INVx1_ASAP7_75t_L g4540 ( 
.A(n_4512),
.Y(n_4540)
);

AND2x2_ASAP7_75t_L g4541 ( 
.A(n_4505),
.B(n_4440),
.Y(n_4541)
);

AND2x2_ASAP7_75t_L g4542 ( 
.A(n_4505),
.B(n_4447),
.Y(n_4542)
);

AOI21xp5_ASAP7_75t_L g4543 ( 
.A1(n_4502),
.A2(n_4460),
.B(n_4437),
.Y(n_4543)
);

INVx1_ASAP7_75t_L g4544 ( 
.A(n_4513),
.Y(n_4544)
);

AND2x2_ASAP7_75t_L g4545 ( 
.A(n_4517),
.B(n_4426),
.Y(n_4545)
);

INVx2_ASAP7_75t_L g4546 ( 
.A(n_4522),
.Y(n_4546)
);

AND2x2_ASAP7_75t_L g4547 ( 
.A(n_4517),
.B(n_4457),
.Y(n_4547)
);

BUFx3_ASAP7_75t_L g4548 ( 
.A(n_4508),
.Y(n_4548)
);

AND2x2_ASAP7_75t_L g4549 ( 
.A(n_4517),
.B(n_4448),
.Y(n_4549)
);

NOR2xp33_ASAP7_75t_L g4550 ( 
.A(n_4478),
.B(n_4463),
.Y(n_4550)
);

INVx1_ASAP7_75t_L g4551 ( 
.A(n_4518),
.Y(n_4551)
);

AND2x2_ASAP7_75t_L g4552 ( 
.A(n_4521),
.B(n_4458),
.Y(n_4552)
);

INVx1_ASAP7_75t_L g4553 ( 
.A(n_4490),
.Y(n_4553)
);

BUFx3_ASAP7_75t_L g4554 ( 
.A(n_4508),
.Y(n_4554)
);

INVx2_ASAP7_75t_SL g4555 ( 
.A(n_4508),
.Y(n_4555)
);

NOR2xp33_ASAP7_75t_L g4556 ( 
.A(n_4484),
.B(n_4469),
.Y(n_4556)
);

INVx1_ASAP7_75t_L g4557 ( 
.A(n_4481),
.Y(n_4557)
);

INVx2_ASAP7_75t_L g4558 ( 
.A(n_4522),
.Y(n_4558)
);

NAND2xp5_ASAP7_75t_L g4559 ( 
.A(n_4481),
.B(n_4334),
.Y(n_4559)
);

AND2x2_ASAP7_75t_L g4560 ( 
.A(n_4521),
.B(n_4334),
.Y(n_4560)
);

BUFx2_ASAP7_75t_L g4561 ( 
.A(n_4516),
.Y(n_4561)
);

INVx1_ASAP7_75t_L g4562 ( 
.A(n_4482),
.Y(n_4562)
);

INVx1_ASAP7_75t_L g4563 ( 
.A(n_4482),
.Y(n_4563)
);

INVxp67_ASAP7_75t_SL g4564 ( 
.A(n_4503),
.Y(n_4564)
);

AND2x2_ASAP7_75t_L g4565 ( 
.A(n_4499),
.B(n_4280),
.Y(n_4565)
);

INVx1_ASAP7_75t_L g4566 ( 
.A(n_4483),
.Y(n_4566)
);

OR2x6_ASAP7_75t_L g4567 ( 
.A(n_4514),
.B(n_4307),
.Y(n_4567)
);

INVx2_ASAP7_75t_L g4568 ( 
.A(n_4526),
.Y(n_4568)
);

AOI21xp33_ASAP7_75t_SL g4569 ( 
.A1(n_4555),
.A2(n_4499),
.B(n_4511),
.Y(n_4569)
);

OR2x2_ASAP7_75t_L g4570 ( 
.A(n_4534),
.B(n_4499),
.Y(n_4570)
);

INVx1_ASAP7_75t_L g4571 ( 
.A(n_4524),
.Y(n_4571)
);

HB1xp67_ASAP7_75t_L g4572 ( 
.A(n_4527),
.Y(n_4572)
);

OR2x2_ASAP7_75t_L g4573 ( 
.A(n_4530),
.B(n_4559),
.Y(n_4573)
);

AND2x2_ASAP7_75t_L g4574 ( 
.A(n_4541),
.B(n_4511),
.Y(n_4574)
);

AOI22xp5_ASAP7_75t_L g4575 ( 
.A1(n_4537),
.A2(n_4459),
.B1(n_4434),
.B2(n_4507),
.Y(n_4575)
);

INVx1_ASAP7_75t_L g4576 ( 
.A(n_4564),
.Y(n_4576)
);

AOI33xp33_ASAP7_75t_L g4577 ( 
.A1(n_4532),
.A2(n_4503),
.A3(n_4520),
.B1(n_4519),
.B2(n_4515),
.B3(n_4211),
.Y(n_4577)
);

AND2x2_ASAP7_75t_L g4578 ( 
.A(n_4535),
.B(n_4511),
.Y(n_4578)
);

OR2x2_ASAP7_75t_L g4579 ( 
.A(n_4528),
.B(n_4483),
.Y(n_4579)
);

NAND2xp5_ASAP7_75t_L g4580 ( 
.A(n_4532),
.B(n_4471),
.Y(n_4580)
);

BUFx2_ASAP7_75t_L g4581 ( 
.A(n_4548),
.Y(n_4581)
);

INVx1_ASAP7_75t_L g4582 ( 
.A(n_4564),
.Y(n_4582)
);

INVx1_ASAP7_75t_L g4583 ( 
.A(n_4536),
.Y(n_4583)
);

INVx1_ASAP7_75t_L g4584 ( 
.A(n_4539),
.Y(n_4584)
);

INVx1_ASAP7_75t_L g4585 ( 
.A(n_4540),
.Y(n_4585)
);

INVx1_ASAP7_75t_L g4586 ( 
.A(n_4544),
.Y(n_4586)
);

NAND2xp33_ASAP7_75t_SL g4587 ( 
.A(n_4529),
.B(n_4523),
.Y(n_4587)
);

OR2x2_ASAP7_75t_L g4588 ( 
.A(n_4531),
.B(n_4510),
.Y(n_4588)
);

AND2x2_ASAP7_75t_L g4589 ( 
.A(n_4549),
.B(n_4510),
.Y(n_4589)
);

INVx2_ASAP7_75t_SL g4590 ( 
.A(n_4548),
.Y(n_4590)
);

OAI21xp33_ASAP7_75t_SL g4591 ( 
.A1(n_4523),
.A2(n_4520),
.B(n_4519),
.Y(n_4591)
);

OR2x2_ASAP7_75t_L g4592 ( 
.A(n_4533),
.B(n_4510),
.Y(n_4592)
);

NOR2x1_ASAP7_75t_L g4593 ( 
.A(n_4554),
.B(n_4145),
.Y(n_4593)
);

INVx1_ASAP7_75t_L g4594 ( 
.A(n_4551),
.Y(n_4594)
);

INVx1_ASAP7_75t_L g4595 ( 
.A(n_4553),
.Y(n_4595)
);

INVx1_ASAP7_75t_L g4596 ( 
.A(n_4557),
.Y(n_4596)
);

OAI22xp5_ASAP7_75t_L g4597 ( 
.A1(n_4550),
.A2(n_4514),
.B1(n_4516),
.B2(n_4442),
.Y(n_4597)
);

OR2x2_ASAP7_75t_L g4598 ( 
.A(n_4583),
.B(n_4532),
.Y(n_4598)
);

INVx1_ASAP7_75t_L g4599 ( 
.A(n_4581),
.Y(n_4599)
);

AOI22xp33_ASAP7_75t_L g4600 ( 
.A1(n_4587),
.A2(n_4550),
.B1(n_4537),
.B2(n_4554),
.Y(n_4600)
);

NAND2xp5_ASAP7_75t_SL g4601 ( 
.A(n_4591),
.B(n_4555),
.Y(n_4601)
);

INVx1_ASAP7_75t_L g4602 ( 
.A(n_4572),
.Y(n_4602)
);

INVx1_ASAP7_75t_L g4603 ( 
.A(n_4576),
.Y(n_4603)
);

INVxp67_ASAP7_75t_L g4604 ( 
.A(n_4590),
.Y(n_4604)
);

INVx1_ASAP7_75t_SL g4605 ( 
.A(n_4593),
.Y(n_4605)
);

INVx2_ASAP7_75t_L g4606 ( 
.A(n_4568),
.Y(n_4606)
);

NOR2x1_ASAP7_75t_L g4607 ( 
.A(n_4582),
.B(n_4567),
.Y(n_4607)
);

INVx2_ASAP7_75t_SL g4608 ( 
.A(n_4573),
.Y(n_4608)
);

INVx1_ASAP7_75t_L g4609 ( 
.A(n_4571),
.Y(n_4609)
);

NAND2xp5_ASAP7_75t_L g4610 ( 
.A(n_4575),
.B(n_4562),
.Y(n_4610)
);

INVx2_ASAP7_75t_SL g4611 ( 
.A(n_4578),
.Y(n_4611)
);

INVx1_ASAP7_75t_L g4612 ( 
.A(n_4579),
.Y(n_4612)
);

AND2x2_ASAP7_75t_L g4613 ( 
.A(n_4589),
.B(n_4525),
.Y(n_4613)
);

OR2x2_ASAP7_75t_L g4614 ( 
.A(n_4575),
.B(n_4543),
.Y(n_4614)
);

AND2x2_ASAP7_75t_L g4615 ( 
.A(n_4574),
.B(n_4538),
.Y(n_4615)
);

AND2x2_ASAP7_75t_L g4616 ( 
.A(n_4597),
.B(n_4547),
.Y(n_4616)
);

AND2x2_ASAP7_75t_L g4617 ( 
.A(n_4577),
.B(n_4545),
.Y(n_4617)
);

HB1xp67_ASAP7_75t_L g4618 ( 
.A(n_4584),
.Y(n_4618)
);

INVx1_ASAP7_75t_L g4619 ( 
.A(n_4585),
.Y(n_4619)
);

OR2x2_ASAP7_75t_L g4620 ( 
.A(n_4592),
.B(n_4543),
.Y(n_4620)
);

OR2x2_ASAP7_75t_L g4621 ( 
.A(n_4580),
.B(n_4565),
.Y(n_4621)
);

OR2x2_ASAP7_75t_L g4622 ( 
.A(n_4599),
.B(n_4588),
.Y(n_4622)
);

INVx1_ASAP7_75t_L g4623 ( 
.A(n_4604),
.Y(n_4623)
);

NAND2xp5_ASAP7_75t_L g4624 ( 
.A(n_4604),
.B(n_4591),
.Y(n_4624)
);

INVx3_ASAP7_75t_SL g4625 ( 
.A(n_4605),
.Y(n_4625)
);

INVxp67_ASAP7_75t_L g4626 ( 
.A(n_4601),
.Y(n_4626)
);

AOI221xp5_ASAP7_75t_L g4627 ( 
.A1(n_4600),
.A2(n_4569),
.B1(n_4594),
.B2(n_4595),
.C(n_4586),
.Y(n_4627)
);

AOI322xp5_ASAP7_75t_L g4628 ( 
.A1(n_4600),
.A2(n_4556),
.A3(n_4561),
.B1(n_4546),
.B2(n_4558),
.C1(n_4526),
.C2(n_4596),
.Y(n_4628)
);

AOI211xp5_ASAP7_75t_SL g4629 ( 
.A1(n_4614),
.A2(n_4570),
.B(n_4556),
.C(n_4099),
.Y(n_4629)
);

INVx1_ASAP7_75t_L g4630 ( 
.A(n_4598),
.Y(n_4630)
);

NOR3xp33_ASAP7_75t_L g4631 ( 
.A(n_4605),
.B(n_4610),
.C(n_4602),
.Y(n_4631)
);

NAND2xp5_ASAP7_75t_L g4632 ( 
.A(n_4620),
.B(n_4611),
.Y(n_4632)
);

INVx1_ASAP7_75t_L g4633 ( 
.A(n_4618),
.Y(n_4633)
);

INVx1_ASAP7_75t_L g4634 ( 
.A(n_4618),
.Y(n_4634)
);

A2O1A1Ixp33_ASAP7_75t_L g4635 ( 
.A1(n_4616),
.A2(n_4569),
.B(n_4546),
.C(n_4558),
.Y(n_4635)
);

INVx1_ASAP7_75t_L g4636 ( 
.A(n_4608),
.Y(n_4636)
);

INVx2_ASAP7_75t_L g4637 ( 
.A(n_4606),
.Y(n_4637)
);

NOR2x1_ASAP7_75t_L g4638 ( 
.A(n_4607),
.B(n_4603),
.Y(n_4638)
);

INVx1_ASAP7_75t_L g4639 ( 
.A(n_4612),
.Y(n_4639)
);

AOI21xp5_ASAP7_75t_L g4640 ( 
.A1(n_4610),
.A2(n_4567),
.B(n_4566),
.Y(n_4640)
);

BUFx2_ASAP7_75t_L g4641 ( 
.A(n_4615),
.Y(n_4641)
);

AOI21xp5_ASAP7_75t_L g4642 ( 
.A1(n_4609),
.A2(n_4567),
.B(n_4563),
.Y(n_4642)
);

INVx1_ASAP7_75t_L g4643 ( 
.A(n_4613),
.Y(n_4643)
);

INVx1_ASAP7_75t_SL g4644 ( 
.A(n_4619),
.Y(n_4644)
);

NAND2xp5_ASAP7_75t_L g4645 ( 
.A(n_4617),
.B(n_4545),
.Y(n_4645)
);

INVx2_ASAP7_75t_SL g4646 ( 
.A(n_4621),
.Y(n_4646)
);

INVx1_ASAP7_75t_L g4647 ( 
.A(n_4599),
.Y(n_4647)
);

INVx1_ASAP7_75t_L g4648 ( 
.A(n_4623),
.Y(n_4648)
);

AND2x2_ASAP7_75t_L g4649 ( 
.A(n_4641),
.B(n_4542),
.Y(n_4649)
);

NAND2xp5_ASAP7_75t_SL g4650 ( 
.A(n_4626),
.B(n_4515),
.Y(n_4650)
);

INVx1_ASAP7_75t_SL g4651 ( 
.A(n_4625),
.Y(n_4651)
);

INVx2_ASAP7_75t_L g4652 ( 
.A(n_4637),
.Y(n_4652)
);

AND2x2_ASAP7_75t_L g4653 ( 
.A(n_4643),
.B(n_4552),
.Y(n_4653)
);

NAND2xp5_ASAP7_75t_SL g4654 ( 
.A(n_4627),
.B(n_4056),
.Y(n_4654)
);

NOR2xp33_ASAP7_75t_L g4655 ( 
.A(n_4624),
.B(n_3937),
.Y(n_4655)
);

INVx1_ASAP7_75t_L g4656 ( 
.A(n_4622),
.Y(n_4656)
);

OR2x2_ASAP7_75t_L g4657 ( 
.A(n_4636),
.B(n_4632),
.Y(n_4657)
);

NOR2xp33_ASAP7_75t_L g4658 ( 
.A(n_4630),
.B(n_3956),
.Y(n_4658)
);

NOR2xp33_ASAP7_75t_L g4659 ( 
.A(n_4635),
.B(n_4217),
.Y(n_4659)
);

NOR2x1_ASAP7_75t_L g4660 ( 
.A(n_4638),
.B(n_4442),
.Y(n_4660)
);

INVx1_ASAP7_75t_SL g4661 ( 
.A(n_4647),
.Y(n_4661)
);

NOR2xp33_ASAP7_75t_L g4662 ( 
.A(n_4646),
.B(n_3777),
.Y(n_4662)
);

NAND3x1_ASAP7_75t_L g4663 ( 
.A(n_4631),
.B(n_4634),
.C(n_4633),
.Y(n_4663)
);

INVx1_ASAP7_75t_L g4664 ( 
.A(n_4639),
.Y(n_4664)
);

INVx1_ASAP7_75t_L g4665 ( 
.A(n_4644),
.Y(n_4665)
);

INVxp67_ASAP7_75t_SL g4666 ( 
.A(n_4640),
.Y(n_4666)
);

NAND2xp5_ASAP7_75t_L g4667 ( 
.A(n_4628),
.B(n_4451),
.Y(n_4667)
);

NAND2xp5_ASAP7_75t_L g4668 ( 
.A(n_4628),
.B(n_4471),
.Y(n_4668)
);

INVxp67_ASAP7_75t_L g4669 ( 
.A(n_4629),
.Y(n_4669)
);

INVx1_ASAP7_75t_L g4670 ( 
.A(n_4645),
.Y(n_4670)
);

INVx1_ASAP7_75t_L g4671 ( 
.A(n_4642),
.Y(n_4671)
);

INVx1_ASAP7_75t_L g4672 ( 
.A(n_4623),
.Y(n_4672)
);

NOR2xp67_ASAP7_75t_L g4673 ( 
.A(n_4623),
.B(n_4560),
.Y(n_4673)
);

NAND2xp5_ASAP7_75t_L g4674 ( 
.A(n_4628),
.B(n_4516),
.Y(n_4674)
);

NAND2xp33_ASAP7_75t_SL g4675 ( 
.A(n_4657),
.B(n_4452),
.Y(n_4675)
);

OR2x2_ASAP7_75t_L g4676 ( 
.A(n_4651),
.B(n_4412),
.Y(n_4676)
);

NOR3xp33_ASAP7_75t_L g4677 ( 
.A(n_4651),
.B(n_4184),
.C(n_4138),
.Y(n_4677)
);

AOI21xp5_ASAP7_75t_L g4678 ( 
.A1(n_4654),
.A2(n_4113),
.B(n_4140),
.Y(n_4678)
);

NAND4xp25_ASAP7_75t_SL g4679 ( 
.A(n_4660),
.B(n_4656),
.C(n_4670),
.D(n_4671),
.Y(n_4679)
);

NAND3xp33_ASAP7_75t_L g4680 ( 
.A(n_4665),
.B(n_4459),
.C(n_4138),
.Y(n_4680)
);

NAND2xp5_ASAP7_75t_L g4681 ( 
.A(n_4666),
.B(n_4649),
.Y(n_4681)
);

AOI322xp5_ASAP7_75t_L g4682 ( 
.A1(n_4669),
.A2(n_4464),
.A3(n_4012),
.B1(n_3998),
.B2(n_3990),
.C1(n_4470),
.C2(n_4416),
.Y(n_4682)
);

OAI221xp5_ASAP7_75t_L g4683 ( 
.A1(n_4674),
.A2(n_4454),
.B1(n_4223),
.B2(n_4180),
.C(n_3828),
.Y(n_4683)
);

NAND2xp5_ASAP7_75t_L g4684 ( 
.A(n_4655),
.B(n_4465),
.Y(n_4684)
);

INVxp67_ASAP7_75t_L g4685 ( 
.A(n_4658),
.Y(n_4685)
);

AOI22xp5_ASAP7_75t_L g4686 ( 
.A1(n_4662),
.A2(n_4465),
.B1(n_4136),
.B2(n_4181),
.Y(n_4686)
);

O2A1O1Ixp33_ASAP7_75t_L g4687 ( 
.A1(n_4648),
.A2(n_4672),
.B(n_4661),
.C(n_4652),
.Y(n_4687)
);

NAND3x1_ASAP7_75t_L g4688 ( 
.A(n_4664),
.B(n_4454),
.C(n_3964),
.Y(n_4688)
);

OAI21xp33_ASAP7_75t_L g4689 ( 
.A1(n_4659),
.A2(n_4303),
.B(n_4205),
.Y(n_4689)
);

NAND2xp5_ASAP7_75t_L g4690 ( 
.A(n_4673),
.B(n_4477),
.Y(n_4690)
);

AOI21xp5_ASAP7_75t_L g4691 ( 
.A1(n_4650),
.A2(n_4181),
.B(n_4136),
.Y(n_4691)
);

INVx1_ASAP7_75t_L g4692 ( 
.A(n_4653),
.Y(n_4692)
);

NAND3xp33_ASAP7_75t_SL g4693 ( 
.A(n_4661),
.B(n_3838),
.C(n_3884),
.Y(n_4693)
);

NOR2xp33_ASAP7_75t_SL g4694 ( 
.A(n_4667),
.B(n_4303),
.Y(n_4694)
);

OAI211xp5_ASAP7_75t_L g4695 ( 
.A1(n_4668),
.A2(n_3955),
.B(n_3933),
.C(n_3979),
.Y(n_4695)
);

INVx1_ASAP7_75t_L g4696 ( 
.A(n_4663),
.Y(n_4696)
);

OAI22xp5_ASAP7_75t_L g4697 ( 
.A1(n_4669),
.A2(n_4485),
.B1(n_4487),
.B2(n_4477),
.Y(n_4697)
);

AOI21xp5_ASAP7_75t_L g4698 ( 
.A1(n_4654),
.A2(n_4120),
.B(n_4189),
.Y(n_4698)
);

AOI221x1_ASAP7_75t_L g4699 ( 
.A1(n_4665),
.A2(n_4197),
.B1(n_4188),
.B2(n_4001),
.C(n_4123),
.Y(n_4699)
);

NOR3xp33_ASAP7_75t_SL g4700 ( 
.A(n_4666),
.B(n_4156),
.C(n_4150),
.Y(n_4700)
);

AOI221xp5_ASAP7_75t_L g4701 ( 
.A1(n_4651),
.A2(n_4214),
.B1(n_4049),
.B2(n_3967),
.C(n_4177),
.Y(n_4701)
);

AND4x1_ASAP7_75t_L g4702 ( 
.A(n_4655),
.B(n_4114),
.C(n_3793),
.D(n_3872),
.Y(n_4702)
);

AOI221xp5_ASAP7_75t_L g4703 ( 
.A1(n_4651),
.A2(n_4214),
.B1(n_4021),
.B2(n_4134),
.C(n_4485),
.Y(n_4703)
);

NAND5xp2_ASAP7_75t_L g4704 ( 
.A(n_4669),
.B(n_3988),
.C(n_3844),
.D(n_4174),
.E(n_3854),
.Y(n_4704)
);

NAND2xp5_ASAP7_75t_L g4705 ( 
.A(n_4651),
.B(n_4487),
.Y(n_4705)
);

O2A1O1Ixp5_ASAP7_75t_SL g4706 ( 
.A1(n_4665),
.A2(n_3958),
.B(n_4401),
.C(n_3827),
.Y(n_4706)
);

INVx1_ASAP7_75t_L g4707 ( 
.A(n_4651),
.Y(n_4707)
);

AOI22x1_ASAP7_75t_L g4708 ( 
.A1(n_4707),
.A2(n_4298),
.B1(n_3958),
.B2(n_4488),
.Y(n_4708)
);

NAND4xp75_ASAP7_75t_L g4709 ( 
.A(n_4681),
.B(n_3822),
.C(n_3744),
.D(n_4215),
.Y(n_4709)
);

NOR2xp67_ASAP7_75t_L g4710 ( 
.A(n_4679),
.B(n_699),
.Y(n_4710)
);

NAND2xp5_ASAP7_75t_L g4711 ( 
.A(n_4694),
.B(n_4368),
.Y(n_4711)
);

INVx1_ASAP7_75t_L g4712 ( 
.A(n_4705),
.Y(n_4712)
);

OAI322xp33_ASAP7_75t_L g4713 ( 
.A1(n_4696),
.A2(n_4500),
.A3(n_4498),
.B1(n_4496),
.B2(n_4488),
.C1(n_4226),
.C2(n_4404),
.Y(n_4713)
);

AOI22xp5_ASAP7_75t_L g4714 ( 
.A1(n_4675),
.A2(n_3786),
.B1(n_4498),
.B2(n_4496),
.Y(n_4714)
);

INVx1_ASAP7_75t_L g4715 ( 
.A(n_4676),
.Y(n_4715)
);

BUFx2_ASAP7_75t_L g4716 ( 
.A(n_4685),
.Y(n_4716)
);

OAI31xp33_ASAP7_75t_L g4717 ( 
.A1(n_4680),
.A2(n_3807),
.A3(n_4088),
.B(n_4500),
.Y(n_4717)
);

O2A1O1Ixp33_ASAP7_75t_SL g4718 ( 
.A1(n_4692),
.A2(n_4083),
.B(n_4166),
.C(n_4148),
.Y(n_4718)
);

BUFx2_ASAP7_75t_L g4719 ( 
.A(n_4690),
.Y(n_4719)
);

AOI222xp33_ASAP7_75t_L g4720 ( 
.A1(n_4697),
.A2(n_4317),
.B1(n_4355),
.B2(n_4365),
.C1(n_4356),
.C2(n_4366),
.Y(n_4720)
);

OAI21xp33_ASAP7_75t_SL g4721 ( 
.A1(n_4684),
.A2(n_3786),
.B(n_4268),
.Y(n_4721)
);

NAND2xp5_ASAP7_75t_L g4722 ( 
.A(n_4682),
.B(n_4368),
.Y(n_4722)
);

INVxp67_ASAP7_75t_L g4723 ( 
.A(n_4678),
.Y(n_4723)
);

O2A1O1Ixp33_ASAP7_75t_L g4724 ( 
.A1(n_4687),
.A2(n_3841),
.B(n_3977),
.C(n_3840),
.Y(n_4724)
);

AOI22xp33_ASAP7_75t_L g4725 ( 
.A1(n_4703),
.A2(n_4258),
.B1(n_4255),
.B2(n_4381),
.Y(n_4725)
);

OAI21xp5_ASAP7_75t_L g4726 ( 
.A1(n_4688),
.A2(n_3953),
.B(n_4018),
.Y(n_4726)
);

NAND2x1p5_ASAP7_75t_L g4727 ( 
.A(n_4702),
.B(n_4298),
.Y(n_4727)
);

NAND2xp5_ASAP7_75t_SL g4728 ( 
.A(n_4689),
.B(n_4255),
.Y(n_4728)
);

NAND2xp5_ASAP7_75t_SL g4729 ( 
.A(n_4700),
.B(n_4255),
.Y(n_4729)
);

INVx1_ASAP7_75t_L g4730 ( 
.A(n_4677),
.Y(n_4730)
);

AOI222xp33_ASAP7_75t_L g4731 ( 
.A1(n_4693),
.A2(n_4356),
.B1(n_4365),
.B2(n_4366),
.C1(n_4351),
.C2(n_4381),
.Y(n_4731)
);

INVx1_ASAP7_75t_L g4732 ( 
.A(n_4683),
.Y(n_4732)
);

AOI22xp5_ASAP7_75t_L g4733 ( 
.A1(n_4698),
.A2(n_4298),
.B1(n_4300),
.B2(n_4258),
.Y(n_4733)
);

A2O1A1Ixp33_ASAP7_75t_SL g4734 ( 
.A1(n_4686),
.A2(n_702),
.B(n_700),
.C(n_701),
.Y(n_4734)
);

OAI21xp5_ASAP7_75t_L g4735 ( 
.A1(n_4706),
.A2(n_3900),
.B(n_3948),
.Y(n_4735)
);

AOI21xp33_ASAP7_75t_SL g4736 ( 
.A1(n_4695),
.A2(n_700),
.B(n_701),
.Y(n_4736)
);

OAI221xp5_ASAP7_75t_L g4737 ( 
.A1(n_4727),
.A2(n_4701),
.B1(n_4691),
.B2(n_4699),
.C(n_4704),
.Y(n_4737)
);

NAND2xp5_ASAP7_75t_L g4738 ( 
.A(n_4710),
.B(n_4368),
.Y(n_4738)
);

INVx1_ASAP7_75t_L g4739 ( 
.A(n_4712),
.Y(n_4739)
);

INVxp67_ASAP7_75t_L g4740 ( 
.A(n_4716),
.Y(n_4740)
);

INVx2_ASAP7_75t_L g4741 ( 
.A(n_4727),
.Y(n_4741)
);

NOR2xp33_ASAP7_75t_L g4742 ( 
.A(n_4729),
.B(n_703),
.Y(n_4742)
);

NOR3x1_ASAP7_75t_L g4743 ( 
.A(n_4734),
.B(n_3981),
.C(n_3959),
.Y(n_4743)
);

INVx2_ASAP7_75t_SL g4744 ( 
.A(n_4728),
.Y(n_4744)
);

INVx1_ASAP7_75t_SL g4745 ( 
.A(n_4719),
.Y(n_4745)
);

NAND2xp5_ASAP7_75t_L g4746 ( 
.A(n_4732),
.B(n_4736),
.Y(n_4746)
);

AOI21xp5_ASAP7_75t_L g4747 ( 
.A1(n_4723),
.A2(n_4715),
.B(n_4730),
.Y(n_4747)
);

INVx1_ASAP7_75t_L g4748 ( 
.A(n_4713),
.Y(n_4748)
);

INVx1_ASAP7_75t_L g4749 ( 
.A(n_4718),
.Y(n_4749)
);

AOI21xp33_ASAP7_75t_SL g4750 ( 
.A1(n_4722),
.A2(n_703),
.B(n_704),
.Y(n_4750)
);

NAND2xp5_ASAP7_75t_L g4751 ( 
.A(n_4709),
.B(n_4368),
.Y(n_4751)
);

INVx1_ASAP7_75t_L g4752 ( 
.A(n_4711),
.Y(n_4752)
);

INVx1_ASAP7_75t_SL g4753 ( 
.A(n_4708),
.Y(n_4753)
);

NOR2x1_ASAP7_75t_L g4754 ( 
.A(n_4726),
.B(n_3928),
.Y(n_4754)
);

AND2x2_ASAP7_75t_L g4755 ( 
.A(n_4731),
.B(n_4380),
.Y(n_4755)
);

XNOR2x1_ASAP7_75t_L g4756 ( 
.A(n_4733),
.B(n_704),
.Y(n_4756)
);

AND2x2_ASAP7_75t_L g4757 ( 
.A(n_4725),
.B(n_4380),
.Y(n_4757)
);

AND2x2_ASAP7_75t_L g4758 ( 
.A(n_4721),
.B(n_4380),
.Y(n_4758)
);

NAND2xp5_ASAP7_75t_L g4759 ( 
.A(n_4717),
.B(n_4380),
.Y(n_4759)
);

INVx2_ASAP7_75t_SL g4760 ( 
.A(n_4714),
.Y(n_4760)
);

NAND2xp33_ASAP7_75t_R g4761 ( 
.A(n_4735),
.B(n_705),
.Y(n_4761)
);

INVx1_ASAP7_75t_L g4762 ( 
.A(n_4724),
.Y(n_4762)
);

AND2x2_ASAP7_75t_L g4763 ( 
.A(n_4720),
.B(n_4380),
.Y(n_4763)
);

OR2x2_ASAP7_75t_L g4764 ( 
.A(n_4712),
.B(n_4391),
.Y(n_4764)
);

NAND2xp5_ASAP7_75t_SL g4765 ( 
.A(n_4710),
.B(n_3821),
.Y(n_4765)
);

NOR2xp67_ASAP7_75t_L g4766 ( 
.A(n_4741),
.B(n_705),
.Y(n_4766)
);

NOR2xp33_ASAP7_75t_R g4767 ( 
.A(n_4749),
.B(n_706),
.Y(n_4767)
);

INVx1_ASAP7_75t_SL g4768 ( 
.A(n_4745),
.Y(n_4768)
);

AOI22xp5_ASAP7_75t_L g4769 ( 
.A1(n_4744),
.A2(n_3968),
.B1(n_3957),
.B2(n_3947),
.Y(n_4769)
);

O2A1O1Ixp33_ASAP7_75t_L g4770 ( 
.A1(n_4740),
.A2(n_3743),
.B(n_3906),
.C(n_709),
.Y(n_4770)
);

HB1xp67_ASAP7_75t_L g4771 ( 
.A(n_4756),
.Y(n_4771)
);

AOI21xp5_ASAP7_75t_L g4772 ( 
.A1(n_4746),
.A2(n_3886),
.B(n_3876),
.Y(n_4772)
);

AOI22xp33_ASAP7_75t_L g4773 ( 
.A1(n_4748),
.A2(n_4245),
.B1(n_4261),
.B2(n_4249),
.Y(n_4773)
);

AOI22xp33_ASAP7_75t_SL g4774 ( 
.A1(n_4745),
.A2(n_4300),
.B1(n_4261),
.B2(n_3905),
.Y(n_4774)
);

AOI322xp5_ASAP7_75t_L g4775 ( 
.A1(n_4760),
.A2(n_4351),
.A3(n_4095),
.B1(n_4024),
.B2(n_4398),
.C1(n_4028),
.C2(n_4026),
.Y(n_4775)
);

NAND2xp5_ASAP7_75t_L g4776 ( 
.A(n_4742),
.B(n_707),
.Y(n_4776)
);

AND2x4_ASAP7_75t_L g4777 ( 
.A(n_4739),
.B(n_4391),
.Y(n_4777)
);

BUFx6f_ASAP7_75t_L g4778 ( 
.A(n_4762),
.Y(n_4778)
);

INVx1_ASAP7_75t_SL g4779 ( 
.A(n_4753),
.Y(n_4779)
);

AOI221xp5_ASAP7_75t_L g4780 ( 
.A1(n_4750),
.A2(n_4364),
.B1(n_4263),
.B2(n_4281),
.C(n_4270),
.Y(n_4780)
);

INVx1_ASAP7_75t_L g4781 ( 
.A(n_4764),
.Y(n_4781)
);

AOI21xp5_ASAP7_75t_L g4782 ( 
.A1(n_4747),
.A2(n_3837),
.B(n_3971),
.Y(n_4782)
);

AOI22xp5_ASAP7_75t_L g4783 ( 
.A1(n_4737),
.A2(n_4300),
.B1(n_4235),
.B2(n_3905),
.Y(n_4783)
);

OAI221xp5_ASAP7_75t_L g4784 ( 
.A1(n_4765),
.A2(n_3978),
.B1(n_3973),
.B2(n_3993),
.C(n_4191),
.Y(n_4784)
);

AOI222xp33_ASAP7_75t_L g4785 ( 
.A1(n_4752),
.A2(n_3939),
.B1(n_3946),
.B2(n_4009),
.C1(n_4005),
.C2(n_4364),
.Y(n_4785)
);

AND2x2_ASAP7_75t_L g4786 ( 
.A(n_4755),
.B(n_4300),
.Y(n_4786)
);

XNOR2xp5_ASAP7_75t_SL g4787 ( 
.A(n_4761),
.B(n_707),
.Y(n_4787)
);

OAI22xp5_ASAP7_75t_L g4788 ( 
.A1(n_4751),
.A2(n_4390),
.B1(n_4382),
.B2(n_4346),
.Y(n_4788)
);

AOI22xp33_ASAP7_75t_SL g4789 ( 
.A1(n_4738),
.A2(n_4300),
.B1(n_3853),
.B2(n_3850),
.Y(n_4789)
);

AOI211xp5_ASAP7_75t_L g4790 ( 
.A1(n_4750),
.A2(n_710),
.B(n_708),
.C(n_709),
.Y(n_4790)
);

NAND2xp5_ASAP7_75t_L g4791 ( 
.A(n_4758),
.B(n_708),
.Y(n_4791)
);

AOI311xp33_ASAP7_75t_L g4792 ( 
.A1(n_4759),
.A2(n_4284),
.A3(n_4265),
.B(n_4160),
.C(n_712),
.Y(n_4792)
);

AOI22xp5_ASAP7_75t_L g4793 ( 
.A1(n_4754),
.A2(n_4235),
.B1(n_3765),
.B2(n_4398),
.Y(n_4793)
);

NAND5xp2_ASAP7_75t_L g4794 ( 
.A(n_4792),
.B(n_4757),
.C(n_4763),
.D(n_4743),
.E(n_712),
.Y(n_4794)
);

OAI222xp33_ASAP7_75t_L g4795 ( 
.A1(n_4768),
.A2(n_4390),
.B1(n_4362),
.B2(n_4348),
.C1(n_4347),
.C2(n_4346),
.Y(n_4795)
);

NAND3xp33_ASAP7_75t_SL g4796 ( 
.A(n_4779),
.B(n_710),
.C(n_711),
.Y(n_4796)
);

AOI211xp5_ASAP7_75t_L g4797 ( 
.A1(n_4766),
.A2(n_715),
.B(n_713),
.C(n_714),
.Y(n_4797)
);

AOI221xp5_ASAP7_75t_L g4798 ( 
.A1(n_4791),
.A2(n_4362),
.B1(n_4348),
.B2(n_4347),
.C(n_4342),
.Y(n_4798)
);

INVx2_ASAP7_75t_L g4799 ( 
.A(n_4777),
.Y(n_4799)
);

AND2x2_ASAP7_75t_L g4800 ( 
.A(n_4786),
.B(n_4339),
.Y(n_4800)
);

INVx1_ASAP7_75t_L g4801 ( 
.A(n_4787),
.Y(n_4801)
);

INVx1_ASAP7_75t_L g4802 ( 
.A(n_4776),
.Y(n_4802)
);

INVx2_ASAP7_75t_L g4803 ( 
.A(n_4781),
.Y(n_4803)
);

AND2x2_ASAP7_75t_SL g4804 ( 
.A(n_4771),
.B(n_3765),
.Y(n_4804)
);

NAND4xp25_ASAP7_75t_L g4805 ( 
.A(n_4790),
.B(n_4770),
.C(n_4772),
.D(n_4782),
.Y(n_4805)
);

NAND2xp5_ASAP7_75t_L g4806 ( 
.A(n_4778),
.B(n_714),
.Y(n_4806)
);

INVx2_ASAP7_75t_L g4807 ( 
.A(n_4778),
.Y(n_4807)
);

INVxp67_ASAP7_75t_L g4808 ( 
.A(n_4784),
.Y(n_4808)
);

NAND2xp5_ASAP7_75t_SL g4809 ( 
.A(n_4767),
.B(n_4773),
.Y(n_4809)
);

NAND4xp25_ASAP7_75t_SL g4810 ( 
.A(n_4783),
.B(n_4342),
.C(n_4340),
.D(n_4339),
.Y(n_4810)
);

NAND3xp33_ASAP7_75t_SL g4811 ( 
.A(n_4789),
.B(n_715),
.C(n_716),
.Y(n_4811)
);

NOR2x1_ASAP7_75t_L g4812 ( 
.A(n_4788),
.B(n_716),
.Y(n_4812)
);

NAND3xp33_ASAP7_75t_SL g4813 ( 
.A(n_4780),
.B(n_4775),
.C(n_4769),
.Y(n_4813)
);

AOI22xp33_ASAP7_75t_L g4814 ( 
.A1(n_4774),
.A2(n_4240),
.B1(n_4259),
.B2(n_4340),
.Y(n_4814)
);

NOR2x1_ASAP7_75t_L g4815 ( 
.A(n_4793),
.B(n_717),
.Y(n_4815)
);

NOR3xp33_ASAP7_75t_L g4816 ( 
.A(n_4785),
.B(n_718),
.C(n_719),
.Y(n_4816)
);

A2O1A1Ixp33_ASAP7_75t_L g4817 ( 
.A1(n_4768),
.A2(n_3870),
.B(n_3847),
.C(n_3858),
.Y(n_4817)
);

OAI22xp5_ASAP7_75t_L g4818 ( 
.A1(n_4808),
.A2(n_3779),
.B1(n_3972),
.B2(n_3825),
.Y(n_4818)
);

NOR2xp67_ASAP7_75t_L g4819 ( 
.A(n_4805),
.B(n_718),
.Y(n_4819)
);

NAND2x1p5_ASAP7_75t_L g4820 ( 
.A(n_4807),
.B(n_3779),
.Y(n_4820)
);

NAND4xp75_ASAP7_75t_L g4821 ( 
.A(n_4806),
.B(n_721),
.C(n_719),
.D(n_720),
.Y(n_4821)
);

NAND4xp75_ASAP7_75t_L g4822 ( 
.A(n_4801),
.B(n_4803),
.C(n_4809),
.D(n_4802),
.Y(n_4822)
);

AND2x4_ASAP7_75t_SL g4823 ( 
.A(n_4799),
.B(n_3779),
.Y(n_4823)
);

INVx1_ASAP7_75t_L g4824 ( 
.A(n_4796),
.Y(n_4824)
);

INVx1_ASAP7_75t_L g4825 ( 
.A(n_4797),
.Y(n_4825)
);

OAI22xp5_ASAP7_75t_SL g4826 ( 
.A1(n_4797),
.A2(n_3825),
.B1(n_3972),
.B2(n_3751),
.Y(n_4826)
);

OAI22xp5_ASAP7_75t_SL g4827 ( 
.A1(n_4804),
.A2(n_3972),
.B1(n_3825),
.B2(n_724),
.Y(n_4827)
);

NOR2x1_ASAP7_75t_L g4828 ( 
.A(n_4811),
.B(n_722),
.Y(n_4828)
);

NOR3xp33_ASAP7_75t_L g4829 ( 
.A(n_4816),
.B(n_4813),
.C(n_4794),
.Y(n_4829)
);

HB1xp67_ASAP7_75t_L g4830 ( 
.A(n_4812),
.Y(n_4830)
);

NOR3x1_ASAP7_75t_L g4831 ( 
.A(n_4815),
.B(n_3869),
.C(n_3866),
.Y(n_4831)
);

HB1xp67_ASAP7_75t_L g4832 ( 
.A(n_4810),
.Y(n_4832)
);

NOR2x1p5_ASAP7_75t_L g4833 ( 
.A(n_4800),
.B(n_722),
.Y(n_4833)
);

HB1xp67_ASAP7_75t_L g4834 ( 
.A(n_4795),
.Y(n_4834)
);

INVx1_ASAP7_75t_L g4835 ( 
.A(n_4814),
.Y(n_4835)
);

BUFx2_ASAP7_75t_L g4836 ( 
.A(n_4798),
.Y(n_4836)
);

AND3x1_ASAP7_75t_L g4837 ( 
.A(n_4817),
.B(n_723),
.C(n_724),
.Y(n_4837)
);

INVx1_ASAP7_75t_L g4838 ( 
.A(n_4819),
.Y(n_4838)
);

INVx1_ASAP7_75t_L g4839 ( 
.A(n_4820),
.Y(n_4839)
);

OAI221xp5_ASAP7_75t_SL g4840 ( 
.A1(n_4829),
.A2(n_723),
.B1(n_725),
.B2(n_726),
.C(n_727),
.Y(n_4840)
);

OAI322xp33_ASAP7_75t_L g4841 ( 
.A1(n_4824),
.A2(n_726),
.A3(n_727),
.B1(n_728),
.B2(n_729),
.C1(n_730),
.C2(n_731),
.Y(n_4841)
);

OAI221xp5_ASAP7_75t_L g4842 ( 
.A1(n_4828),
.A2(n_728),
.B1(n_729),
.B2(n_730),
.C(n_731),
.Y(n_4842)
);

OAI22xp33_ASAP7_75t_SL g4843 ( 
.A1(n_4835),
.A2(n_735),
.B1(n_732),
.B2(n_734),
.Y(n_4843)
);

A2O1A1Ixp33_ASAP7_75t_L g4844 ( 
.A1(n_4823),
.A2(n_3860),
.B(n_3868),
.C(n_3766),
.Y(n_4844)
);

OAI211xp5_ASAP7_75t_SL g4845 ( 
.A1(n_4825),
.A2(n_736),
.B(n_732),
.C(n_734),
.Y(n_4845)
);

AOI22xp5_ASAP7_75t_L g4846 ( 
.A1(n_4822),
.A2(n_4827),
.B1(n_4834),
.B2(n_4836),
.Y(n_4846)
);

OAI322xp33_ASAP7_75t_SL g4847 ( 
.A1(n_4837),
.A2(n_737),
.A3(n_738),
.B1(n_739),
.B2(n_740),
.C1(n_741),
.C2(n_742),
.Y(n_4847)
);

OAI211xp5_ASAP7_75t_L g4848 ( 
.A1(n_4830),
.A2(n_744),
.B(n_737),
.C(n_739),
.Y(n_4848)
);

OAI211xp5_ASAP7_75t_L g4849 ( 
.A1(n_4832),
.A2(n_748),
.B(n_745),
.C(n_746),
.Y(n_4849)
);

OAI22xp5_ASAP7_75t_L g4850 ( 
.A1(n_4833),
.A2(n_4259),
.B1(n_4293),
.B2(n_4290),
.Y(n_4850)
);

AOI322xp5_ASAP7_75t_L g4851 ( 
.A1(n_4821),
.A2(n_745),
.A3(n_748),
.B1(n_749),
.B2(n_751),
.C1(n_752),
.C2(n_753),
.Y(n_4851)
);

AOI322xp5_ASAP7_75t_L g4852 ( 
.A1(n_4818),
.A2(n_751),
.A3(n_752),
.B1(n_753),
.B2(n_754),
.C1(n_755),
.C2(n_757),
.Y(n_4852)
);

INVx2_ASAP7_75t_L g4853 ( 
.A(n_4831),
.Y(n_4853)
);

OAI322xp33_ASAP7_75t_SL g4854 ( 
.A1(n_4826),
.A2(n_754),
.A3(n_755),
.B1(n_758),
.B2(n_759),
.C1(n_760),
.C2(n_761),
.Y(n_4854)
);

AOI322xp5_ASAP7_75t_L g4855 ( 
.A1(n_4829),
.A2(n_761),
.A3(n_762),
.B1(n_763),
.B2(n_764),
.C1(n_765),
.C2(n_766),
.Y(n_4855)
);

INVx2_ASAP7_75t_L g4856 ( 
.A(n_4839),
.Y(n_4856)
);

INVx2_ASAP7_75t_L g4857 ( 
.A(n_4853),
.Y(n_4857)
);

BUFx2_ASAP7_75t_L g4858 ( 
.A(n_4846),
.Y(n_4858)
);

OAI22xp5_ASAP7_75t_L g4859 ( 
.A1(n_4838),
.A2(n_4293),
.B1(n_4290),
.B2(n_4264),
.Y(n_4859)
);

OA22x2_ASAP7_75t_L g4860 ( 
.A1(n_4849),
.A2(n_3938),
.B1(n_3771),
.B2(n_3764),
.Y(n_4860)
);

AOI22xp33_ASAP7_75t_L g4861 ( 
.A1(n_4845),
.A2(n_4842),
.B1(n_4841),
.B2(n_4843),
.Y(n_4861)
);

NAND2xp5_ASAP7_75t_L g4862 ( 
.A(n_4855),
.B(n_763),
.Y(n_4862)
);

INVx2_ASAP7_75t_L g4863 ( 
.A(n_4850),
.Y(n_4863)
);

CKINVDCx20_ASAP7_75t_R g4864 ( 
.A(n_4847),
.Y(n_4864)
);

XNOR2xp5_ASAP7_75t_L g4865 ( 
.A(n_4848),
.B(n_765),
.Y(n_4865)
);

OAI22xp33_ASAP7_75t_L g4866 ( 
.A1(n_4854),
.A2(n_4283),
.B1(n_4264),
.B2(n_768),
.Y(n_4866)
);

OAI21xp33_ASAP7_75t_L g4867 ( 
.A1(n_4840),
.A2(n_3728),
.B(n_3741),
.Y(n_4867)
);

HB1xp67_ASAP7_75t_L g4868 ( 
.A(n_4851),
.Y(n_4868)
);

AND2x4_ASAP7_75t_L g4869 ( 
.A(n_4852),
.B(n_766),
.Y(n_4869)
);

AOI21xp5_ASAP7_75t_L g4870 ( 
.A1(n_4862),
.A2(n_4844),
.B(n_767),
.Y(n_4870)
);

AOI21xp5_ASAP7_75t_L g4871 ( 
.A1(n_4856),
.A2(n_4865),
.B(n_4858),
.Y(n_4871)
);

NAND2xp5_ASAP7_75t_L g4872 ( 
.A(n_4857),
.B(n_767),
.Y(n_4872)
);

HB1xp67_ASAP7_75t_L g4873 ( 
.A(n_4868),
.Y(n_4873)
);

AOI21xp5_ASAP7_75t_L g4874 ( 
.A1(n_4866),
.A2(n_4869),
.B(n_4861),
.Y(n_4874)
);

NAND2xp5_ASAP7_75t_L g4875 ( 
.A(n_4867),
.B(n_768),
.Y(n_4875)
);

AOI22xp5_ASAP7_75t_L g4876 ( 
.A1(n_4864),
.A2(n_4240),
.B1(n_3762),
.B2(n_3733),
.Y(n_4876)
);

OAI21xp5_ASAP7_75t_L g4877 ( 
.A1(n_4863),
.A2(n_3780),
.B(n_3718),
.Y(n_4877)
);

AOI22x1_ASAP7_75t_L g4878 ( 
.A1(n_4859),
.A2(n_769),
.B1(n_770),
.B2(n_771),
.Y(n_4878)
);

INVx1_ASAP7_75t_L g4879 ( 
.A(n_4860),
.Y(n_4879)
);

INVx1_ASAP7_75t_L g4880 ( 
.A(n_4856),
.Y(n_4880)
);

OAI22xp5_ASAP7_75t_L g4881 ( 
.A1(n_4880),
.A2(n_4283),
.B1(n_770),
.B2(n_771),
.Y(n_4881)
);

AOI22xp5_ASAP7_75t_L g4882 ( 
.A1(n_4873),
.A2(n_3738),
.B1(n_3735),
.B2(n_3722),
.Y(n_4882)
);

OAI22x1_ASAP7_75t_L g4883 ( 
.A1(n_4878),
.A2(n_769),
.B1(n_772),
.B2(n_773),
.Y(n_4883)
);

OAI22xp5_ASAP7_75t_SL g4884 ( 
.A1(n_4872),
.A2(n_772),
.B1(n_773),
.B2(n_774),
.Y(n_4884)
);

INVx2_ASAP7_75t_L g4885 ( 
.A(n_4879),
.Y(n_4885)
);

AOI22xp5_ASAP7_75t_L g4886 ( 
.A1(n_4874),
.A2(n_775),
.B1(n_776),
.B2(n_777),
.Y(n_4886)
);

CKINVDCx20_ASAP7_75t_R g4887 ( 
.A(n_4871),
.Y(n_4887)
);

INVx1_ASAP7_75t_L g4888 ( 
.A(n_4885),
.Y(n_4888)
);

AOI22xp33_ASAP7_75t_L g4889 ( 
.A1(n_4887),
.A2(n_4875),
.B1(n_4870),
.B2(n_4877),
.Y(n_4889)
);

INVx1_ASAP7_75t_L g4890 ( 
.A(n_4884),
.Y(n_4890)
);

OR2x2_ASAP7_75t_L g4891 ( 
.A(n_4888),
.B(n_4886),
.Y(n_4891)
);

OAI221xp5_ASAP7_75t_L g4892 ( 
.A1(n_4889),
.A2(n_4881),
.B1(n_4876),
.B2(n_4883),
.C(n_4882),
.Y(n_4892)
);

AOI22xp33_ASAP7_75t_L g4893 ( 
.A1(n_4891),
.A2(n_4890),
.B1(n_777),
.B2(n_778),
.Y(n_4893)
);

AOI322xp5_ASAP7_75t_L g4894 ( 
.A1(n_4893),
.A2(n_4892),
.A3(n_778),
.B1(n_779),
.B2(n_780),
.C1(n_781),
.C2(n_782),
.Y(n_4894)
);

AOI22xp5_ASAP7_75t_L g4895 ( 
.A1(n_4894),
.A2(n_776),
.B1(n_779),
.B2(n_780),
.Y(n_4895)
);

AOI211xp5_ASAP7_75t_L g4896 ( 
.A1(n_4895),
.A2(n_781),
.B(n_783),
.C(n_784),
.Y(n_4896)
);


endmodule