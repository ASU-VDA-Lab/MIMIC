module fake_jpeg_2477_n_206 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_206);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_206;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_143;
wire n_202;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g48 ( 
.A(n_29),
.Y(n_48)
);

INVx11_ASAP7_75t_L g49 ( 
.A(n_21),
.Y(n_49)
);

INVx6_ASAP7_75t_SL g50 ( 
.A(n_39),
.Y(n_50)
);

BUFx10_ASAP7_75t_L g51 ( 
.A(n_32),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_30),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_19),
.B(n_7),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_0),
.Y(n_54)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_5),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_28),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_42),
.Y(n_57)
);

INVx1_ASAP7_75t_SL g58 ( 
.A(n_23),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_31),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_47),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_26),
.Y(n_61)
);

BUFx12_ASAP7_75t_L g62 ( 
.A(n_6),
.Y(n_62)
);

BUFx10_ASAP7_75t_L g63 ( 
.A(n_40),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_0),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_15),
.Y(n_65)
);

BUFx12f_ASAP7_75t_L g66 ( 
.A(n_9),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_27),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_16),
.Y(n_68)
);

CKINVDCx16_ASAP7_75t_R g69 ( 
.A(n_50),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_69),
.B(n_71),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_56),
.Y(n_70)
);

INVx6_ASAP7_75t_L g88 ( 
.A(n_70),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_58),
.B(n_1),
.Y(n_71)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_55),
.Y(n_72)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_72),
.Y(n_87)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_55),
.Y(n_73)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_73),
.Y(n_89)
);

INVx11_ASAP7_75t_L g74 ( 
.A(n_66),
.Y(n_74)
);

BUFx8_ASAP7_75t_L g84 ( 
.A(n_74),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_53),
.B(n_1),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_75),
.B(n_2),
.Y(n_90)
);

HB1xp67_ASAP7_75t_L g76 ( 
.A(n_66),
.Y(n_76)
);

CKINVDCx16_ASAP7_75t_R g85 ( 
.A(n_76),
.Y(n_85)
);

BUFx16f_ASAP7_75t_L g77 ( 
.A(n_69),
.Y(n_77)
);

BUFx3_ASAP7_75t_L g92 ( 
.A(n_77),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_74),
.A2(n_58),
.B1(n_49),
.B2(n_66),
.Y(n_78)
);

INVxp67_ASAP7_75t_L g91 ( 
.A(n_78),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_72),
.A2(n_56),
.B1(n_57),
.B2(n_66),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_79),
.A2(n_73),
.B1(n_70),
.B2(n_76),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_L g80 ( 
.A1(n_72),
.A2(n_49),
.B1(n_68),
.B2(n_64),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_80),
.A2(n_70),
.B1(n_54),
.B2(n_59),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_75),
.B(n_48),
.Y(n_81)
);

A2O1A1Ixp33_ASAP7_75t_L g97 ( 
.A1(n_81),
.A2(n_71),
.B(n_54),
.C(n_52),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_74),
.A2(n_68),
.B1(n_64),
.B2(n_65),
.Y(n_82)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_82),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_75),
.B(n_65),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_86),
.B(n_90),
.Y(n_101)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_89),
.Y(n_93)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_93),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_94),
.A2(n_100),
.B1(n_87),
.B2(n_52),
.Y(n_110)
);

BUFx2_ASAP7_75t_L g95 ( 
.A(n_84),
.Y(n_95)
);

CKINVDCx14_ASAP7_75t_R g123 ( 
.A(n_95),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_97),
.B(n_81),
.Y(n_112)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_89),
.Y(n_98)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_98),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_87),
.B(n_73),
.C(n_48),
.Y(n_99)
);

XNOR2xp5_ASAP7_75t_L g119 ( 
.A(n_99),
.B(n_63),
.Y(n_119)
);

HB1xp67_ASAP7_75t_L g102 ( 
.A(n_84),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_102),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_83),
.B(n_61),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_103),
.B(n_104),
.Y(n_111)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_85),
.Y(n_104)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_84),
.Y(n_105)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_105),
.Y(n_116)
);

O2A1O1Ixp33_ASAP7_75t_L g106 ( 
.A1(n_77),
.A2(n_50),
.B(n_67),
.C(n_61),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_106),
.B(n_88),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_79),
.A2(n_70),
.B1(n_67),
.B2(n_57),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_107),
.A2(n_88),
.B1(n_63),
.B2(n_51),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_83),
.B(n_59),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_108),
.B(n_60),
.Y(n_113)
);

O2A1O1Ixp33_ASAP7_75t_SL g109 ( 
.A1(n_96),
.A2(n_84),
.B(n_77),
.C(n_85),
.Y(n_109)
);

A2O1A1O1Ixp25_ASAP7_75t_L g144 ( 
.A1(n_109),
.A2(n_51),
.B(n_62),
.C(n_46),
.D(n_45),
.Y(n_144)
);

INVxp33_ASAP7_75t_L g139 ( 
.A(n_110),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_SL g145 ( 
.A(n_112),
.B(n_113),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_114),
.B(n_115),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_101),
.B(n_90),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_107),
.A2(n_88),
.B1(n_63),
.B2(n_51),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_117),
.A2(n_105),
.B1(n_95),
.B2(n_63),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_99),
.B(n_2),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_118),
.B(n_120),
.Y(n_140)
);

XOR2xp5_ASAP7_75t_L g135 ( 
.A(n_119),
.B(n_91),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_92),
.B(n_3),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_97),
.B(n_3),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_122),
.B(n_124),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_92),
.B(n_4),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_125),
.A2(n_117),
.B1(n_123),
.B2(n_116),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_100),
.B(n_4),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_126),
.B(n_5),
.Y(n_136)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_128),
.Y(n_129)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_129),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_119),
.B(n_96),
.C(n_94),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_131),
.B(n_135),
.C(n_141),
.Y(n_151)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_128),
.Y(n_132)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_132),
.Y(n_160)
);

AOI21xp5_ASAP7_75t_L g133 ( 
.A1(n_114),
.A2(n_91),
.B(n_106),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_L g162 ( 
.A1(n_133),
.A2(n_144),
.B(n_41),
.Y(n_162)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_127),
.Y(n_134)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_134),
.Y(n_163)
);

NOR3xp33_ASAP7_75t_L g158 ( 
.A(n_136),
.B(n_148),
.C(n_10),
.Y(n_158)
);

AOI22xp33_ASAP7_75t_SL g168 ( 
.A1(n_137),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_111),
.B(n_6),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_SL g161 ( 
.A(n_138),
.B(n_43),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_SL g141 ( 
.A(n_110),
.B(n_109),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_142),
.A2(n_147),
.B1(n_144),
.B2(n_137),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g146 ( 
.A(n_116),
.Y(n_146)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_146),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_125),
.A2(n_51),
.B1(n_62),
.B2(n_44),
.Y(n_147)
);

NOR2x1_ASAP7_75t_L g148 ( 
.A(n_109),
.B(n_62),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_127),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_149),
.B(n_8),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_130),
.B(n_121),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_150),
.B(n_153),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_139),
.A2(n_121),
.B1(n_8),
.B2(n_9),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_152),
.A2(n_154),
.B1(n_159),
.B2(n_168),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_146),
.Y(n_153)
);

AOI221xp5_ASAP7_75t_L g154 ( 
.A1(n_131),
.A2(n_135),
.B1(n_145),
.B2(n_148),
.C(n_141),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_140),
.B(n_7),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_155),
.B(n_158),
.Y(n_172)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_157),
.Y(n_171)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_161),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_SL g179 ( 
.A1(n_162),
.A2(n_166),
.B(n_25),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_139),
.B(n_38),
.C(n_37),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_164),
.B(n_35),
.C(n_34),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_143),
.B(n_10),
.Y(n_165)
);

CKINVDCx16_ASAP7_75t_R g177 ( 
.A(n_165),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_L g166 ( 
.A1(n_142),
.A2(n_11),
.B(n_12),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_147),
.B(n_36),
.Y(n_169)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_169),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g187 ( 
.A(n_170),
.B(n_180),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_L g175 ( 
.A(n_151),
.B(n_33),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_175),
.B(n_181),
.C(n_182),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_179),
.B(n_13),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_SL g180 ( 
.A1(n_150),
.A2(n_24),
.B(n_14),
.Y(n_180)
);

XOR2xp5_ASAP7_75t_L g181 ( 
.A(n_151),
.B(n_156),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g182 ( 
.A(n_160),
.B(n_163),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_173),
.A2(n_166),
.B1(n_152),
.B2(n_169),
.Y(n_183)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_183),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_L g184 ( 
.A1(n_178),
.A2(n_162),
.B1(n_164),
.B2(n_160),
.Y(n_184)
);

NOR4xp25_ASAP7_75t_L g196 ( 
.A(n_184),
.B(n_186),
.C(n_182),
.D(n_18),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_185),
.B(n_188),
.C(n_190),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_177),
.B(n_163),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_181),
.B(n_167),
.C(n_15),
.Y(n_188)
);

NAND3xp33_ASAP7_75t_L g189 ( 
.A(n_171),
.B(n_167),
.C(n_16),
.Y(n_189)
);

OAI31xp33_ASAP7_75t_L g194 ( 
.A1(n_189),
.A2(n_172),
.A3(n_176),
.B(n_19),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_175),
.B(n_14),
.C(n_17),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_191),
.B(n_174),
.C(n_170),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_193),
.B(n_194),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_196),
.B(n_197),
.Y(n_199)
);

A2O1A1Ixp33_ASAP7_75t_SL g197 ( 
.A1(n_191),
.A2(n_17),
.B(n_18),
.C(n_20),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_195),
.B(n_187),
.C(n_192),
.Y(n_200)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_200),
.B(n_197),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_SL g203 ( 
.A(n_201),
.B(n_202),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_SL g202 ( 
.A1(n_198),
.A2(n_189),
.B(n_21),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_203),
.B(n_199),
.C(n_22),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_L g205 ( 
.A1(n_204),
.A2(n_20),
.B(n_22),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_205),
.B(n_23),
.Y(n_206)
);


endmodule