module fake_netlist_6_4501_n_2157 (n_52, n_435, n_1, n_91, n_326, n_256, n_440, n_209, n_367, n_465, n_63, n_223, n_278, n_341, n_362, n_148, n_226, n_161, n_22, n_208, n_462, n_68, n_316, n_419, n_28, n_304, n_212, n_50, n_7, n_144, n_365, n_125, n_168, n_384, n_297, n_342, n_77, n_106, n_358, n_160, n_449, n_131, n_188, n_310, n_186, n_245, n_0, n_368, n_396, n_495, n_350, n_78, n_84, n_392, n_442, n_480, n_142, n_143, n_382, n_180, n_62, n_349, n_233, n_255, n_284, n_400, n_140, n_337, n_214, n_485, n_67, n_15, n_443, n_246, n_38, n_471, n_289, n_421, n_424, n_59, n_181, n_182, n_238, n_202, n_320, n_108, n_327, n_369, n_280, n_287, n_353, n_389, n_415, n_65, n_230, n_461, n_141, n_383, n_200, n_447, n_176, n_114, n_86, n_198, n_104, n_222, n_179, n_248, n_300, n_71, n_74, n_229, n_305, n_72, n_173, n_250, n_372, n_468, n_111, n_314, n_378, n_413, n_377, n_35, n_183, n_79, n_375, n_338, n_466, n_56, n_360, n_119, n_235, n_147, n_191, n_340, n_387, n_452, n_39, n_344, n_73, n_428, n_432, n_101, n_167, n_174, n_127, n_153, n_156, n_491, n_145, n_42, n_133, n_96, n_8, n_371, n_189, n_405, n_213, n_294, n_302, n_380, n_129, n_197, n_11, n_137, n_17, n_343, n_448, n_20, n_494, n_493, n_397, n_155, n_109, n_445, n_425, n_122, n_45, n_454, n_34, n_218, n_70, n_234, n_37, n_486, n_381, n_82, n_27, n_236, n_112, n_172, n_472, n_270, n_239, n_126, n_414, n_97, n_58, n_490, n_290, n_220, n_118, n_224, n_48, n_25, n_93, n_80, n_196, n_402, n_352, n_478, n_9, n_460, n_107, n_6, n_417, n_14, n_446, n_89, n_374, n_366, n_407, n_450, n_103, n_272, n_185, n_348, n_69, n_376, n_390, n_473, n_293, n_31, n_334, n_53, n_370, n_44, n_458, n_232, n_16, n_163, n_46, n_330, n_470, n_475, n_298, n_18, n_492, n_281, n_258, n_154, n_456, n_98, n_260, n_265, n_313, n_451, n_279, n_252, n_228, n_356, n_166, n_184, n_216, n_455, n_83, n_363, n_395, n_323, n_393, n_411, n_152, n_92, n_321, n_331, n_105, n_227, n_132, n_406, n_483, n_102, n_204, n_482, n_474, n_261, n_420, n_312, n_394, n_32, n_66, n_130, n_164, n_292, n_100, n_121, n_307, n_469, n_433, n_23, n_476, n_2, n_291, n_219, n_357, n_150, n_264, n_263, n_481, n_325, n_329, n_464, n_33, n_477, n_408, n_61, n_237, n_244, n_399, n_76, n_243, n_124, n_94, n_282, n_436, n_116, n_211, n_117, n_175, n_322, n_345, n_409, n_231, n_354, n_40, n_240, n_139, n_319, n_41, n_134, n_273, n_95, n_311, n_10, n_403, n_253, n_123, n_136, n_249, n_201, n_386, n_159, n_157, n_162, n_115, n_487, n_128, n_241, n_30, n_275, n_43, n_276, n_441, n_221, n_444, n_423, n_146, n_318, n_303, n_467, n_306, n_21, n_193, n_269, n_359, n_346, n_88, n_3, n_416, n_277, n_418, n_113, n_4, n_199, n_138, n_266, n_296, n_268, n_271, n_404, n_439, n_158, n_217, n_49, n_210, n_299, n_206, n_5, n_453, n_333, n_215, n_178, n_247, n_225, n_308, n_309, n_355, n_426, n_317, n_149, n_431, n_90, n_347, n_24, n_459, n_54, n_328, n_488, n_429, n_373, n_87, n_195, n_285, n_497, n_85, n_99, n_257, n_13, n_203, n_286, n_254, n_207, n_242, n_19, n_47, n_29, n_75, n_401, n_324, n_335, n_430, n_463, n_489, n_205, n_120, n_251, n_301, n_274, n_110, n_151, n_412, n_81, n_36, n_26, n_55, n_267, n_438, n_339, n_315, n_434, n_64, n_288, n_427, n_479, n_496, n_422, n_135, n_165, n_351, n_437, n_259, n_177, n_391, n_457, n_364, n_295, n_385, n_388, n_190, n_262, n_484, n_187, n_60, n_361, n_379, n_170, n_332, n_336, n_12, n_398, n_410, n_194, n_171, n_192, n_57, n_169, n_51, n_283, n_2157);

input n_52;
input n_435;
input n_1;
input n_91;
input n_326;
input n_256;
input n_440;
input n_209;
input n_367;
input n_465;
input n_63;
input n_223;
input n_278;
input n_341;
input n_362;
input n_148;
input n_226;
input n_161;
input n_22;
input n_208;
input n_462;
input n_68;
input n_316;
input n_419;
input n_28;
input n_304;
input n_212;
input n_50;
input n_7;
input n_144;
input n_365;
input n_125;
input n_168;
input n_384;
input n_297;
input n_342;
input n_77;
input n_106;
input n_358;
input n_160;
input n_449;
input n_131;
input n_188;
input n_310;
input n_186;
input n_245;
input n_0;
input n_368;
input n_396;
input n_495;
input n_350;
input n_78;
input n_84;
input n_392;
input n_442;
input n_480;
input n_142;
input n_143;
input n_382;
input n_180;
input n_62;
input n_349;
input n_233;
input n_255;
input n_284;
input n_400;
input n_140;
input n_337;
input n_214;
input n_485;
input n_67;
input n_15;
input n_443;
input n_246;
input n_38;
input n_471;
input n_289;
input n_421;
input n_424;
input n_59;
input n_181;
input n_182;
input n_238;
input n_202;
input n_320;
input n_108;
input n_327;
input n_369;
input n_280;
input n_287;
input n_353;
input n_389;
input n_415;
input n_65;
input n_230;
input n_461;
input n_141;
input n_383;
input n_200;
input n_447;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_222;
input n_179;
input n_248;
input n_300;
input n_71;
input n_74;
input n_229;
input n_305;
input n_72;
input n_173;
input n_250;
input n_372;
input n_468;
input n_111;
input n_314;
input n_378;
input n_413;
input n_377;
input n_35;
input n_183;
input n_79;
input n_375;
input n_338;
input n_466;
input n_56;
input n_360;
input n_119;
input n_235;
input n_147;
input n_191;
input n_340;
input n_387;
input n_452;
input n_39;
input n_344;
input n_73;
input n_428;
input n_432;
input n_101;
input n_167;
input n_174;
input n_127;
input n_153;
input n_156;
input n_491;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_371;
input n_189;
input n_405;
input n_213;
input n_294;
input n_302;
input n_380;
input n_129;
input n_197;
input n_11;
input n_137;
input n_17;
input n_343;
input n_448;
input n_20;
input n_494;
input n_493;
input n_397;
input n_155;
input n_109;
input n_445;
input n_425;
input n_122;
input n_45;
input n_454;
input n_34;
input n_218;
input n_70;
input n_234;
input n_37;
input n_486;
input n_381;
input n_82;
input n_27;
input n_236;
input n_112;
input n_172;
input n_472;
input n_270;
input n_239;
input n_126;
input n_414;
input n_97;
input n_58;
input n_490;
input n_290;
input n_220;
input n_118;
input n_224;
input n_48;
input n_25;
input n_93;
input n_80;
input n_196;
input n_402;
input n_352;
input n_478;
input n_9;
input n_460;
input n_107;
input n_6;
input n_417;
input n_14;
input n_446;
input n_89;
input n_374;
input n_366;
input n_407;
input n_450;
input n_103;
input n_272;
input n_185;
input n_348;
input n_69;
input n_376;
input n_390;
input n_473;
input n_293;
input n_31;
input n_334;
input n_53;
input n_370;
input n_44;
input n_458;
input n_232;
input n_16;
input n_163;
input n_46;
input n_330;
input n_470;
input n_475;
input n_298;
input n_18;
input n_492;
input n_281;
input n_258;
input n_154;
input n_456;
input n_98;
input n_260;
input n_265;
input n_313;
input n_451;
input n_279;
input n_252;
input n_228;
input n_356;
input n_166;
input n_184;
input n_216;
input n_455;
input n_83;
input n_363;
input n_395;
input n_323;
input n_393;
input n_411;
input n_152;
input n_92;
input n_321;
input n_331;
input n_105;
input n_227;
input n_132;
input n_406;
input n_483;
input n_102;
input n_204;
input n_482;
input n_474;
input n_261;
input n_420;
input n_312;
input n_394;
input n_32;
input n_66;
input n_130;
input n_164;
input n_292;
input n_100;
input n_121;
input n_307;
input n_469;
input n_433;
input n_23;
input n_476;
input n_2;
input n_291;
input n_219;
input n_357;
input n_150;
input n_264;
input n_263;
input n_481;
input n_325;
input n_329;
input n_464;
input n_33;
input n_477;
input n_408;
input n_61;
input n_237;
input n_244;
input n_399;
input n_76;
input n_243;
input n_124;
input n_94;
input n_282;
input n_436;
input n_116;
input n_211;
input n_117;
input n_175;
input n_322;
input n_345;
input n_409;
input n_231;
input n_354;
input n_40;
input n_240;
input n_139;
input n_319;
input n_41;
input n_134;
input n_273;
input n_95;
input n_311;
input n_10;
input n_403;
input n_253;
input n_123;
input n_136;
input n_249;
input n_201;
input n_386;
input n_159;
input n_157;
input n_162;
input n_115;
input n_487;
input n_128;
input n_241;
input n_30;
input n_275;
input n_43;
input n_276;
input n_441;
input n_221;
input n_444;
input n_423;
input n_146;
input n_318;
input n_303;
input n_467;
input n_306;
input n_21;
input n_193;
input n_269;
input n_359;
input n_346;
input n_88;
input n_3;
input n_416;
input n_277;
input n_418;
input n_113;
input n_4;
input n_199;
input n_138;
input n_266;
input n_296;
input n_268;
input n_271;
input n_404;
input n_439;
input n_158;
input n_217;
input n_49;
input n_210;
input n_299;
input n_206;
input n_5;
input n_453;
input n_333;
input n_215;
input n_178;
input n_247;
input n_225;
input n_308;
input n_309;
input n_355;
input n_426;
input n_317;
input n_149;
input n_431;
input n_90;
input n_347;
input n_24;
input n_459;
input n_54;
input n_328;
input n_488;
input n_429;
input n_373;
input n_87;
input n_195;
input n_285;
input n_497;
input n_85;
input n_99;
input n_257;
input n_13;
input n_203;
input n_286;
input n_254;
input n_207;
input n_242;
input n_19;
input n_47;
input n_29;
input n_75;
input n_401;
input n_324;
input n_335;
input n_430;
input n_463;
input n_489;
input n_205;
input n_120;
input n_251;
input n_301;
input n_274;
input n_110;
input n_151;
input n_412;
input n_81;
input n_36;
input n_26;
input n_55;
input n_267;
input n_438;
input n_339;
input n_315;
input n_434;
input n_64;
input n_288;
input n_427;
input n_479;
input n_496;
input n_422;
input n_135;
input n_165;
input n_351;
input n_437;
input n_259;
input n_177;
input n_391;
input n_457;
input n_364;
input n_295;
input n_385;
input n_388;
input n_190;
input n_262;
input n_484;
input n_187;
input n_60;
input n_361;
input n_379;
input n_170;
input n_332;
input n_336;
input n_12;
input n_398;
input n_410;
input n_194;
input n_171;
input n_192;
input n_57;
input n_169;
input n_51;
input n_283;

output n_2157;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_1212;
wire n_726;
wire n_700;
wire n_1307;
wire n_2003;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_1853;
wire n_783;
wire n_1738;
wire n_798;
wire n_1575;
wire n_1854;
wire n_1923;
wire n_509;
wire n_1342;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_1739;
wire n_2051;
wire n_1380;
wire n_1402;
wire n_1688;
wire n_1691;
wire n_1975;
wire n_1009;
wire n_1743;
wire n_1930;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1991;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_1844;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_1786;
wire n_830;
wire n_873;
wire n_1371;
wire n_1285;
wire n_1985;
wire n_1803;
wire n_1172;
wire n_852;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1867;
wire n_1704;
wire n_1078;
wire n_544;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_2019;
wire n_836;
wire n_2074;
wire n_522;
wire n_2129;
wire n_1261;
wire n_945;
wire n_1649;
wire n_2018;
wire n_2094;
wire n_1903;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_616;
wire n_658;
wire n_1874;
wire n_1119;
wire n_2013;
wire n_1433;
wire n_1902;
wire n_1842;
wire n_1620;
wire n_2044;
wire n_1954;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1798;
wire n_1550;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_1971;
wire n_2058;
wire n_2090;
wire n_538;
wire n_2004;
wire n_1106;
wire n_886;
wire n_1471;
wire n_953;
wire n_1094;
wire n_1345;
wire n_1820;
wire n_539;
wire n_2108;
wire n_1421;
wire n_1936;
wire n_638;
wire n_1404;
wire n_1211;
wire n_2124;
wire n_887;
wire n_1660;
wire n_1961;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_2155;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_1894;
wire n_1231;
wire n_1978;
wire n_2085;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_1815;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_1193;
wire n_1967;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1911;
wire n_1956;
wire n_1644;
wire n_2011;
wire n_1558;
wire n_1732;
wire n_551;
wire n_699;
wire n_1986;
wire n_564;
wire n_824;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_2113;
wire n_1918;
wire n_577;
wire n_1843;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_813;
wire n_1909;
wire n_2080;
wire n_1481;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_2104;
wire n_513;
wire n_645;
wire n_1381;
wire n_1699;
wire n_916;
wire n_2093;
wire n_1970;
wire n_608;
wire n_2101;
wire n_630;
wire n_2059;
wire n_541;
wire n_512;
wire n_2073;
wire n_792;
wire n_1328;
wire n_1957;
wire n_1907;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_982;
wire n_549;
wire n_1762;
wire n_1910;
wire n_1075;
wire n_932;
wire n_1876;
wire n_1895;
wire n_2123;
wire n_1697;
wire n_2143;
wire n_979;
wire n_1873;
wire n_905;
wire n_1866;
wire n_1680;
wire n_993;
wire n_689;
wire n_2031;
wire n_2130;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1988;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_2009;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_2068;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_2072;
wire n_1354;
wire n_586;
wire n_1875;
wire n_1865;
wire n_1701;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_1950;
wire n_530;
wire n_1563;
wire n_1912;
wire n_1982;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_1335;
wire n_1760;
wire n_1927;
wire n_2028;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_1165;
wire n_702;
wire n_2008;
wire n_1926;
wire n_1175;
wire n_1386;
wire n_1896;
wire n_1747;
wire n_1012;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1977;
wire n_1802;
wire n_1504;
wire n_1655;
wire n_835;
wire n_928;
wire n_1214;
wire n_850;
wire n_690;
wire n_1801;
wire n_1886;
wire n_2092;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_1813;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_1124;
wire n_1624;
wire n_515;
wire n_2096;
wire n_1965;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_697;
wire n_687;
wire n_890;
wire n_637;
wire n_701;
wire n_950;
wire n_2036;
wire n_2152;
wire n_1709;
wire n_1825;
wire n_1757;
wire n_1796;
wire n_1792;
wire n_891;
wire n_2067;
wire n_2136;
wire n_2082;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_2075;
wire n_1987;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_1990;
wire n_694;
wire n_2150;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_2078;
wire n_595;
wire n_627;
wire n_1767;
wire n_1779;
wire n_524;
wire n_1465;
wire n_1858;
wire n_1044;
wire n_2133;
wire n_1712;
wire n_1391;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_673;
wire n_1969;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_2145;
wire n_1968;
wire n_898;
wire n_1952;
wire n_865;
wire n_925;
wire n_1932;
wire n_1101;
wire n_1026;
wire n_1880;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_2151;
wire n_1451;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_1839;
wire n_685;
wire n_1765;
wire n_605;
wire n_1514;
wire n_1863;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_996;
wire n_532;
wire n_1308;
wire n_2089;
wire n_1376;
wire n_1513;
wire n_791;
wire n_1913;
wire n_510;
wire n_837;
wire n_2097;
wire n_1488;
wire n_1808;
wire n_948;
wire n_704;
wire n_2148;
wire n_977;
wire n_1005;
wire n_1947;
wire n_536;
wire n_1788;
wire n_1999;
wire n_622;
wire n_1469;
wire n_2060;
wire n_1838;
wire n_1835;
wire n_1776;
wire n_1766;
wire n_1959;
wire n_2002;
wire n_581;
wire n_2138;
wire n_765;
wire n_1492;
wire n_987;
wire n_1340;
wire n_1771;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_1878;
wire n_899;
wire n_738;
wire n_2012;
wire n_1304;
wire n_1035;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_2134;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_2069;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_1577;
wire n_1181;
wire n_2119;
wire n_1822;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_1992;
wire n_648;
wire n_657;
wire n_1049;
wire n_2057;
wire n_2103;
wire n_1666;
wire n_1505;
wire n_803;
wire n_1717;
wire n_926;
wire n_1817;
wire n_927;
wire n_1849;
wire n_919;
wire n_1698;
wire n_929;
wire n_1228;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_2127;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_1195;
wire n_2137;
wire n_1626;
wire n_1507;
wire n_552;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_912;
wire n_1857;
wire n_1519;
wire n_2144;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_1395;
wire n_2110;
wire n_731;
wire n_1502;
wire n_1659;
wire n_1955;
wire n_755;
wire n_931;
wire n_1021;
wire n_527;
wire n_683;
wire n_811;
wire n_1207;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_1250;
wire n_1137;
wire n_1897;
wire n_2064;
wire n_880;
wire n_2053;
wire n_2121;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_1942;
wire n_1966;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_1837;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_1440;
wire n_2132;
wire n_2063;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_1483;
wire n_1834;
wire n_1372;
wire n_1457;
wire n_505;
wire n_1719;
wire n_1339;
wire n_1787;
wire n_537;
wire n_1993;
wire n_1427;
wire n_1466;
wire n_1919;
wire n_1080;
wire n_723;
wire n_1877;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_1939;
wire n_2030;
wire n_1769;
wire n_1220;
wire n_1893;
wire n_556;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_2025;
wire n_1125;
wire n_970;
wire n_1980;
wire n_642;
wire n_995;
wire n_1159;
wire n_1092;
wire n_1060;
wire n_1951;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_511;
wire n_1286;
wire n_1773;
wire n_1775;
wire n_2115;
wire n_1053;
wire n_1681;
wire n_520;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_775;
wire n_651;
wire n_1153;
wire n_1618;
wire n_518;
wire n_1531;
wire n_1185;
wire n_1745;
wire n_914;
wire n_759;
wire n_1831;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_2146;
wire n_2131;
wire n_773;
wire n_1901;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1892;
wire n_1933;
wire n_1135;
wire n_1179;
wire n_1169;
wire n_1617;
wire n_1470;
wire n_1243;
wire n_848;
wire n_1096;
wire n_1091;
wire n_1917;
wire n_2000;
wire n_1580;
wire n_1425;
wire n_1881;
wire n_1267;
wire n_1281;
wire n_1806;
wire n_983;
wire n_2023;
wire n_1520;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_1731;
wire n_2087;
wire n_1855;
wire n_1636;
wire n_1437;
wire n_2135;
wire n_1645;
wire n_1832;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_2049;
wire n_1331;
wire n_736;
wire n_613;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_2100;
wire n_778;
wire n_1668;
wire n_1134;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1995;
wire n_1594;
wire n_664;
wire n_1869;
wire n_1764;
wire n_1429;
wire n_1610;
wire n_1889;
wire n_2016;
wire n_1905;
wire n_793;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_1937;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_1744;
wire n_828;
wire n_2139;
wire n_2142;
wire n_607;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_1254;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_724;
wire n_1934;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_1871;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_1549;
wire n_1510;
wire n_892;
wire n_768;
wire n_1468;
wire n_1859;
wire n_2102;
wire n_1095;
wire n_2024;
wire n_1595;
wire n_2156;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_1916;
wire n_597;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1852;
wire n_1024;
wire n_1768;
wire n_2153;
wire n_1847;
wire n_2052;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_750;
wire n_1115;
wire n_901;
wire n_1499;
wire n_923;
wire n_504;
wire n_1409;
wire n_1841;
wire n_1639;
wire n_1623;
wire n_1015;
wire n_1503;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_1126;
wire n_1997;
wire n_710;
wire n_1108;
wire n_1818;
wire n_1182;
wire n_1298;
wire n_2088;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1960;
wire n_2061;
wire n_1686;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1943;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_1694;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_1983;
wire n_1938;
wire n_1262;
wire n_1891;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_2037;
wire n_782;
wire n_1539;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_2120;
wire n_1472;
wire n_2050;
wire n_1081;
wire n_1870;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_1827;
wire n_1361;
wire n_1864;
wire n_2006;
wire n_1491;
wire n_662;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_2017;
wire n_1695;
wire n_1828;
wire n_2046;
wire n_650;
wire n_1046;
wire n_1940;
wire n_1979;
wire n_1145;
wire n_1121;
wire n_1102;
wire n_1963;
wire n_972;
wire n_1405;
wire n_1406;
wire n_1332;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_1569;
wire n_936;
wire n_1883;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_2084;
wire n_654;
wire n_1222;
wire n_599;
wire n_776;
wire n_1823;
wire n_1974;
wire n_1720;
wire n_934;
wire n_1637;
wire n_1407;
wire n_1795;
wire n_1341;
wire n_1456;
wire n_1845;
wire n_1489;
wire n_942;
wire n_1524;
wire n_543;
wire n_1964;
wire n_1920;
wire n_2099;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_2007;
wire n_2039;
wire n_1946;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_1640;
wire n_804;
wire n_1846;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_2141;
wire n_1343;
wire n_1522;
wire n_548;
wire n_1782;
wire n_1676;
wire n_833;
wire n_1830;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_1900;
wire n_799;
wire n_1548;
wire n_1155;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_2021;
wire n_2114;
wire n_1086;
wire n_1066;
wire n_1948;
wire n_2125;
wire n_2026;
wire n_1282;
wire n_550;
wire n_652;
wire n_2154;
wire n_560;
wire n_1906;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_1758;
wire n_1925;
wire n_737;
wire n_1318;
wire n_1914;
wire n_1235;
wire n_1229;
wire n_1292;
wire n_1373;
wire n_1029;
wire n_1447;
wire n_2056;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_1248;
wire n_1556;
wire n_902;
wire n_1047;
wire n_1984;
wire n_1385;
wire n_1269;
wire n_1931;
wire n_2083;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_1375;
wire n_1941;
wire n_2128;
wire n_655;
wire n_706;
wire n_1045;
wire n_1794;
wire n_786;
wire n_1650;
wire n_1236;
wire n_1962;
wire n_1559;
wire n_1725;
wire n_1928;
wire n_1872;
wire n_834;
wire n_743;
wire n_766;
wire n_1746;
wire n_1325;
wire n_1002;
wire n_1741;
wire n_1949;
wire n_545;
wire n_1804;
wire n_1727;
wire n_1019;
wire n_636;
wire n_2054;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_2062;
wire n_2041;
wire n_1477;
wire n_1360;
wire n_1860;
wire n_1904;
wire n_1200;
wire n_2070;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1908;
wire n_1454;
wire n_2126;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_1098;
wire n_1329;
wire n_2045;
wire n_817;
wire n_897;
wire n_846;
wire n_2066;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1800;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_1191;
wire n_1826;
wire n_566;
wire n_1023;
wire n_1882;
wire n_1076;
wire n_1118;
wire n_1007;
wire n_1807;
wire n_1929;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1814;
wire n_1631;
wire n_591;
wire n_1377;
wire n_1879;
wire n_853;
wire n_695;
wire n_1542;
wire n_875;
wire n_680;
wire n_1678;
wire n_661;
wire n_1716;
wire n_1256;
wire n_671;
wire n_1953;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_1976;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1824;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_2122;
wire n_2109;
wire n_1435;
wire n_969;
wire n_988;
wire n_2140;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_2029;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_955;
wire n_1379;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_1810;
wire n_573;
wire n_769;
wire n_676;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_814;
wire n_1643;
wire n_2020;
wire n_1729;
wire n_669;
wire n_2048;
wire n_2005;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_691;
wire n_535;
wire n_2076;
wire n_1408;
wire n_1196;
wire n_1598;
wire n_863;
wire n_601;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1848;
wire n_1147;
wire n_763;
wire n_1785;
wire n_1754;
wire n_2149;
wire n_1506;
wire n_1652;
wire n_1812;
wire n_957;
wire n_1994;
wire n_895;
wire n_866;
wire n_1227;
wire n_744;
wire n_971;
wire n_946;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_1173;
wire n_1924;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_1174;
wire n_1944;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_844;
wire n_1017;
wire n_2117;
wire n_1083;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_2081;
wire n_2022;
wire n_1945;
wire n_910;
wire n_1721;
wire n_1656;
wire n_1460;
wire n_911;
wire n_2112;
wire n_1464;
wire n_653;
wire n_1737;
wire n_1414;
wire n_908;
wire n_752;
wire n_944;
wire n_2034;
wire n_576;
wire n_1028;
wire n_2106;
wire n_1922;
wire n_563;
wire n_2032;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_1973;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1821;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_712;
wire n_1276;
wire n_2015;
wire n_2118;
wire n_2111;
wire n_1148;
wire n_1989;
wire n_1161;
wire n_1085;
wire n_2014;
wire n_2042;
wire n_1239;
wire n_771;
wire n_1584;
wire n_924;
wire n_1582;
wire n_1149;
wire n_1184;
wire n_719;
wire n_1972;
wire n_1525;
wire n_1585;
wire n_1851;
wire n_1799;
wire n_1090;
wire n_2147;
wire n_592;
wire n_1816;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_984;
wire n_1829;
wire n_503;
wire n_2035;
wire n_1450;
wire n_1638;
wire n_868;
wire n_859;
wire n_570;
wire n_2033;
wire n_735;
wire n_1789;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_1144;
wire n_2071;
wire n_985;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_2010;
wire n_1651;
wire n_1198;
wire n_2047;
wire n_2095;
wire n_1609;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1998;
wire n_1574;
wire n_756;
wire n_1619;
wire n_1981;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_1552;
wire n_583;
wire n_1996;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_2043;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_973;
wire n_1921;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_2065;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_2001;
wire n_2107;
wire n_1884;
wire n_2040;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_1260;
wire n_1819;
wire n_2055;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_2038;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_1861;
wire n_1632;
wire n_1890;
wire n_1805;
wire n_1557;
wire n_1888;
wire n_1833;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_1850;
wire n_1898;
wire n_1868;
wire n_2079;
wire n_1089;
wire n_1887;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_1242;
wire n_2086;
wire n_1836;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_640;
wire n_1322;
wire n_965;
wire n_1899;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_1856;
wire n_1862;
wire n_1958;
wire n_2077;
wire n_784;
wire n_1059;
wire n_1197;
wire n_722;
wire n_862;
wire n_2105;
wire n_2098;
wire n_540;
wire n_1423;
wire n_1935;
wire n_2027;
wire n_2091;
wire n_1915;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_827;
wire n_531;
wire n_1025;
wire n_2116;
wire n_1885;
wire n_1013;
wire n_1259;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g498 ( 
.A(n_84),
.Y(n_498)
);

CKINVDCx5p33_ASAP7_75t_R g499 ( 
.A(n_117),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_433),
.Y(n_500)
);

CKINVDCx5p33_ASAP7_75t_R g501 ( 
.A(n_26),
.Y(n_501)
);

CKINVDCx5p33_ASAP7_75t_R g502 ( 
.A(n_337),
.Y(n_502)
);

INVx2_ASAP7_75t_SL g503 ( 
.A(n_23),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_436),
.Y(n_504)
);

INVx1_ASAP7_75t_SL g505 ( 
.A(n_333),
.Y(n_505)
);

CKINVDCx5p33_ASAP7_75t_R g506 ( 
.A(n_243),
.Y(n_506)
);

CKINVDCx5p33_ASAP7_75t_R g507 ( 
.A(n_304),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_366),
.Y(n_508)
);

CKINVDCx5p33_ASAP7_75t_R g509 ( 
.A(n_292),
.Y(n_509)
);

CKINVDCx5p33_ASAP7_75t_R g510 ( 
.A(n_46),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_2),
.Y(n_511)
);

CKINVDCx5p33_ASAP7_75t_R g512 ( 
.A(n_462),
.Y(n_512)
);

CKINVDCx5p33_ASAP7_75t_R g513 ( 
.A(n_261),
.Y(n_513)
);

CKINVDCx5p33_ASAP7_75t_R g514 ( 
.A(n_489),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_452),
.Y(n_515)
);

CKINVDCx5p33_ASAP7_75t_R g516 ( 
.A(n_496),
.Y(n_516)
);

CKINVDCx20_ASAP7_75t_R g517 ( 
.A(n_313),
.Y(n_517)
);

BUFx6f_ASAP7_75t_L g518 ( 
.A(n_215),
.Y(n_518)
);

CKINVDCx5p33_ASAP7_75t_R g519 ( 
.A(n_228),
.Y(n_519)
);

CKINVDCx5p33_ASAP7_75t_R g520 ( 
.A(n_386),
.Y(n_520)
);

CKINVDCx5p33_ASAP7_75t_R g521 ( 
.A(n_71),
.Y(n_521)
);

CKINVDCx16_ASAP7_75t_R g522 ( 
.A(n_244),
.Y(n_522)
);

CKINVDCx5p33_ASAP7_75t_R g523 ( 
.A(n_497),
.Y(n_523)
);

CKINVDCx20_ASAP7_75t_R g524 ( 
.A(n_484),
.Y(n_524)
);

CKINVDCx5p33_ASAP7_75t_R g525 ( 
.A(n_415),
.Y(n_525)
);

CKINVDCx20_ASAP7_75t_R g526 ( 
.A(n_106),
.Y(n_526)
);

CKINVDCx20_ASAP7_75t_R g527 ( 
.A(n_157),
.Y(n_527)
);

BUFx6f_ASAP7_75t_L g528 ( 
.A(n_485),
.Y(n_528)
);

CKINVDCx5p33_ASAP7_75t_R g529 ( 
.A(n_320),
.Y(n_529)
);

CKINVDCx5p33_ASAP7_75t_R g530 ( 
.A(n_140),
.Y(n_530)
);

CKINVDCx5p33_ASAP7_75t_R g531 ( 
.A(n_447),
.Y(n_531)
);

CKINVDCx5p33_ASAP7_75t_R g532 ( 
.A(n_355),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_262),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_158),
.Y(n_534)
);

CKINVDCx5p33_ASAP7_75t_R g535 ( 
.A(n_327),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_234),
.Y(n_536)
);

CKINVDCx5p33_ASAP7_75t_R g537 ( 
.A(n_249),
.Y(n_537)
);

CKINVDCx5p33_ASAP7_75t_R g538 ( 
.A(n_345),
.Y(n_538)
);

CKINVDCx5p33_ASAP7_75t_R g539 ( 
.A(n_81),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_434),
.Y(n_540)
);

BUFx3_ASAP7_75t_L g541 ( 
.A(n_431),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_379),
.Y(n_542)
);

INVx2_ASAP7_75t_L g543 ( 
.A(n_162),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_295),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_487),
.Y(n_545)
);

CKINVDCx5p33_ASAP7_75t_R g546 ( 
.A(n_162),
.Y(n_546)
);

BUFx6f_ASAP7_75t_L g547 ( 
.A(n_268),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_358),
.Y(n_548)
);

CKINVDCx5p33_ASAP7_75t_R g549 ( 
.A(n_343),
.Y(n_549)
);

CKINVDCx5p33_ASAP7_75t_R g550 ( 
.A(n_387),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_450),
.Y(n_551)
);

INVx2_ASAP7_75t_L g552 ( 
.A(n_231),
.Y(n_552)
);

CKINVDCx5p33_ASAP7_75t_R g553 ( 
.A(n_285),
.Y(n_553)
);

INVx1_ASAP7_75t_SL g554 ( 
.A(n_53),
.Y(n_554)
);

CKINVDCx20_ASAP7_75t_R g555 ( 
.A(n_394),
.Y(n_555)
);

CKINVDCx5p33_ASAP7_75t_R g556 ( 
.A(n_478),
.Y(n_556)
);

CKINVDCx5p33_ASAP7_75t_R g557 ( 
.A(n_453),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_335),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_48),
.Y(n_559)
);

CKINVDCx20_ASAP7_75t_R g560 ( 
.A(n_99),
.Y(n_560)
);

CKINVDCx5p33_ASAP7_75t_R g561 ( 
.A(n_481),
.Y(n_561)
);

CKINVDCx5p33_ASAP7_75t_R g562 ( 
.A(n_200),
.Y(n_562)
);

BUFx5_ASAP7_75t_L g563 ( 
.A(n_491),
.Y(n_563)
);

CKINVDCx5p33_ASAP7_75t_R g564 ( 
.A(n_98),
.Y(n_564)
);

CKINVDCx20_ASAP7_75t_R g565 ( 
.A(n_430),
.Y(n_565)
);

CKINVDCx5p33_ASAP7_75t_R g566 ( 
.A(n_306),
.Y(n_566)
);

BUFx3_ASAP7_75t_L g567 ( 
.A(n_265),
.Y(n_567)
);

CKINVDCx5p33_ASAP7_75t_R g568 ( 
.A(n_44),
.Y(n_568)
);

CKINVDCx5p33_ASAP7_75t_R g569 ( 
.A(n_289),
.Y(n_569)
);

CKINVDCx5p33_ASAP7_75t_R g570 ( 
.A(n_477),
.Y(n_570)
);

CKINVDCx16_ASAP7_75t_R g571 ( 
.A(n_374),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_4),
.Y(n_572)
);

CKINVDCx5p33_ASAP7_75t_R g573 ( 
.A(n_417),
.Y(n_573)
);

CKINVDCx5p33_ASAP7_75t_R g574 ( 
.A(n_392),
.Y(n_574)
);

INVxp67_ASAP7_75t_L g575 ( 
.A(n_67),
.Y(n_575)
);

CKINVDCx14_ASAP7_75t_R g576 ( 
.A(n_143),
.Y(n_576)
);

BUFx5_ASAP7_75t_L g577 ( 
.A(n_133),
.Y(n_577)
);

INVx2_ASAP7_75t_L g578 ( 
.A(n_486),
.Y(n_578)
);

BUFx10_ASAP7_75t_L g579 ( 
.A(n_84),
.Y(n_579)
);

INVx2_ASAP7_75t_L g580 ( 
.A(n_45),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_2),
.Y(n_581)
);

CKINVDCx5p33_ASAP7_75t_R g582 ( 
.A(n_166),
.Y(n_582)
);

CKINVDCx5p33_ASAP7_75t_R g583 ( 
.A(n_300),
.Y(n_583)
);

CKINVDCx5p33_ASAP7_75t_R g584 ( 
.A(n_65),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_221),
.Y(n_585)
);

BUFx3_ASAP7_75t_L g586 ( 
.A(n_191),
.Y(n_586)
);

BUFx3_ASAP7_75t_L g587 ( 
.A(n_382),
.Y(n_587)
);

CKINVDCx5p33_ASAP7_75t_R g588 ( 
.A(n_381),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_323),
.Y(n_589)
);

BUFx3_ASAP7_75t_L g590 ( 
.A(n_239),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_413),
.Y(n_591)
);

CKINVDCx5p33_ASAP7_75t_R g592 ( 
.A(n_102),
.Y(n_592)
);

CKINVDCx5p33_ASAP7_75t_R g593 ( 
.A(n_27),
.Y(n_593)
);

CKINVDCx5p33_ASAP7_75t_R g594 ( 
.A(n_143),
.Y(n_594)
);

INVx4_ASAP7_75t_R g595 ( 
.A(n_321),
.Y(n_595)
);

CKINVDCx5p33_ASAP7_75t_R g596 ( 
.A(n_488),
.Y(n_596)
);

CKINVDCx5p33_ASAP7_75t_R g597 ( 
.A(n_92),
.Y(n_597)
);

CKINVDCx5p33_ASAP7_75t_R g598 ( 
.A(n_359),
.Y(n_598)
);

CKINVDCx5p33_ASAP7_75t_R g599 ( 
.A(n_137),
.Y(n_599)
);

CKINVDCx5p33_ASAP7_75t_R g600 ( 
.A(n_97),
.Y(n_600)
);

HB1xp67_ASAP7_75t_L g601 ( 
.A(n_204),
.Y(n_601)
);

CKINVDCx5p33_ASAP7_75t_R g602 ( 
.A(n_246),
.Y(n_602)
);

CKINVDCx5p33_ASAP7_75t_R g603 ( 
.A(n_35),
.Y(n_603)
);

CKINVDCx5p33_ASAP7_75t_R g604 ( 
.A(n_479),
.Y(n_604)
);

BUFx6f_ASAP7_75t_L g605 ( 
.A(n_90),
.Y(n_605)
);

CKINVDCx20_ASAP7_75t_R g606 ( 
.A(n_206),
.Y(n_606)
);

CKINVDCx5p33_ASAP7_75t_R g607 ( 
.A(n_224),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_466),
.Y(n_608)
);

CKINVDCx5p33_ASAP7_75t_R g609 ( 
.A(n_101),
.Y(n_609)
);

CKINVDCx5p33_ASAP7_75t_R g610 ( 
.A(n_102),
.Y(n_610)
);

CKINVDCx5p33_ASAP7_75t_R g611 ( 
.A(n_330),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_439),
.Y(n_612)
);

CKINVDCx5p33_ASAP7_75t_R g613 ( 
.A(n_181),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_172),
.Y(n_614)
);

CKINVDCx5p33_ASAP7_75t_R g615 ( 
.A(n_407),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_113),
.Y(n_616)
);

CKINVDCx20_ASAP7_75t_R g617 ( 
.A(n_401),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_112),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_269),
.Y(n_619)
);

CKINVDCx5p33_ASAP7_75t_R g620 ( 
.A(n_214),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_12),
.Y(n_621)
);

BUFx6f_ASAP7_75t_L g622 ( 
.A(n_119),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_410),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_294),
.Y(n_624)
);

CKINVDCx5p33_ASAP7_75t_R g625 ( 
.A(n_82),
.Y(n_625)
);

BUFx3_ASAP7_75t_L g626 ( 
.A(n_483),
.Y(n_626)
);

INVx1_ASAP7_75t_SL g627 ( 
.A(n_369),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_264),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_389),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_425),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_492),
.Y(n_631)
);

CKINVDCx5p33_ASAP7_75t_R g632 ( 
.A(n_225),
.Y(n_632)
);

CKINVDCx5p33_ASAP7_75t_R g633 ( 
.A(n_29),
.Y(n_633)
);

CKINVDCx5p33_ASAP7_75t_R g634 ( 
.A(n_42),
.Y(n_634)
);

INVx2_ASAP7_75t_L g635 ( 
.A(n_480),
.Y(n_635)
);

CKINVDCx20_ASAP7_75t_R g636 ( 
.A(n_119),
.Y(n_636)
);

CKINVDCx20_ASAP7_75t_R g637 ( 
.A(n_257),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_446),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_451),
.Y(n_639)
);

CKINVDCx5p33_ASAP7_75t_R g640 ( 
.A(n_108),
.Y(n_640)
);

CKINVDCx5p33_ASAP7_75t_R g641 ( 
.A(n_456),
.Y(n_641)
);

CKINVDCx5p33_ASAP7_75t_R g642 ( 
.A(n_164),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_1),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_42),
.Y(n_644)
);

CKINVDCx5p33_ASAP7_75t_R g645 ( 
.A(n_155),
.Y(n_645)
);

INVxp33_ASAP7_75t_R g646 ( 
.A(n_160),
.Y(n_646)
);

CKINVDCx5p33_ASAP7_75t_R g647 ( 
.A(n_175),
.Y(n_647)
);

INVx1_ASAP7_75t_SL g648 ( 
.A(n_86),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_35),
.Y(n_649)
);

CKINVDCx5p33_ASAP7_75t_R g650 ( 
.A(n_94),
.Y(n_650)
);

INVx2_ASAP7_75t_SL g651 ( 
.A(n_305),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_93),
.Y(n_652)
);

CKINVDCx20_ASAP7_75t_R g653 ( 
.A(n_472),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_474),
.Y(n_654)
);

CKINVDCx5p33_ASAP7_75t_R g655 ( 
.A(n_470),
.Y(n_655)
);

CKINVDCx5p33_ASAP7_75t_R g656 ( 
.A(n_288),
.Y(n_656)
);

INVx2_ASAP7_75t_L g657 ( 
.A(n_362),
.Y(n_657)
);

CKINVDCx20_ASAP7_75t_R g658 ( 
.A(n_399),
.Y(n_658)
);

CKINVDCx5p33_ASAP7_75t_R g659 ( 
.A(n_133),
.Y(n_659)
);

BUFx8_ASAP7_75t_SL g660 ( 
.A(n_191),
.Y(n_660)
);

CKINVDCx5p33_ASAP7_75t_R g661 ( 
.A(n_291),
.Y(n_661)
);

CKINVDCx16_ASAP7_75t_R g662 ( 
.A(n_216),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_82),
.Y(n_663)
);

CKINVDCx5p33_ASAP7_75t_R g664 ( 
.A(n_159),
.Y(n_664)
);

CKINVDCx5p33_ASAP7_75t_R g665 ( 
.A(n_147),
.Y(n_665)
);

CKINVDCx20_ASAP7_75t_R g666 ( 
.A(n_482),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_167),
.Y(n_667)
);

INVx2_ASAP7_75t_SL g668 ( 
.A(n_86),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_331),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_142),
.Y(n_670)
);

BUFx10_ASAP7_75t_L g671 ( 
.A(n_338),
.Y(n_671)
);

INVx2_ASAP7_75t_SL g672 ( 
.A(n_307),
.Y(n_672)
);

CKINVDCx14_ASAP7_75t_R g673 ( 
.A(n_124),
.Y(n_673)
);

CKINVDCx5p33_ASAP7_75t_R g674 ( 
.A(n_384),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_274),
.Y(n_675)
);

BUFx5_ASAP7_75t_L g676 ( 
.A(n_324),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_101),
.Y(n_677)
);

BUFx2_ASAP7_75t_SL g678 ( 
.A(n_303),
.Y(n_678)
);

CKINVDCx5p33_ASAP7_75t_R g679 ( 
.A(n_226),
.Y(n_679)
);

BUFx3_ASAP7_75t_L g680 ( 
.A(n_467),
.Y(n_680)
);

CKINVDCx5p33_ASAP7_75t_R g681 ( 
.A(n_280),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_93),
.Y(n_682)
);

BUFx10_ASAP7_75t_L g683 ( 
.A(n_252),
.Y(n_683)
);

BUFx10_ASAP7_75t_L g684 ( 
.A(n_88),
.Y(n_684)
);

CKINVDCx5p33_ASAP7_75t_R g685 ( 
.A(n_118),
.Y(n_685)
);

CKINVDCx5p33_ASAP7_75t_R g686 ( 
.A(n_229),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_361),
.Y(n_687)
);

CKINVDCx5p33_ASAP7_75t_R g688 ( 
.A(n_114),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_340),
.Y(n_689)
);

CKINVDCx5p33_ASAP7_75t_R g690 ( 
.A(n_293),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_577),
.Y(n_691)
);

INVx2_ASAP7_75t_SL g692 ( 
.A(n_579),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_577),
.Y(n_693)
);

CKINVDCx20_ASAP7_75t_R g694 ( 
.A(n_660),
.Y(n_694)
);

BUFx3_ASAP7_75t_L g695 ( 
.A(n_567),
.Y(n_695)
);

INVx2_ASAP7_75t_L g696 ( 
.A(n_577),
.Y(n_696)
);

INVx2_ASAP7_75t_L g697 ( 
.A(n_577),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_577),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_577),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_586),
.Y(n_700)
);

CKINVDCx20_ASAP7_75t_R g701 ( 
.A(n_526),
.Y(n_701)
);

INVx2_ASAP7_75t_L g702 ( 
.A(n_563),
.Y(n_702)
);

INVxp33_ASAP7_75t_SL g703 ( 
.A(n_601),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_586),
.Y(n_704)
);

INVxp33_ASAP7_75t_SL g705 ( 
.A(n_601),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_605),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_605),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_605),
.Y(n_708)
);

NOR2xp67_ASAP7_75t_L g709 ( 
.A(n_575),
.B(n_0),
.Y(n_709)
);

INVx2_ASAP7_75t_L g710 ( 
.A(n_563),
.Y(n_710)
);

INVxp67_ASAP7_75t_SL g711 ( 
.A(n_541),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_605),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_622),
.Y(n_713)
);

INVx2_ASAP7_75t_L g714 ( 
.A(n_563),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_622),
.Y(n_715)
);

INVxp67_ASAP7_75t_SL g716 ( 
.A(n_541),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_622),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_622),
.Y(n_718)
);

INVx2_ASAP7_75t_L g719 ( 
.A(n_563),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_511),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_534),
.Y(n_721)
);

CKINVDCx20_ASAP7_75t_R g722 ( 
.A(n_527),
.Y(n_722)
);

CKINVDCx16_ASAP7_75t_R g723 ( 
.A(n_522),
.Y(n_723)
);

INVxp67_ASAP7_75t_SL g724 ( 
.A(n_587),
.Y(n_724)
);

BUFx3_ASAP7_75t_L g725 ( 
.A(n_680),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_559),
.Y(n_726)
);

INVxp67_ASAP7_75t_SL g727 ( 
.A(n_587),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_572),
.Y(n_728)
);

INVxp33_ASAP7_75t_SL g729 ( 
.A(n_498),
.Y(n_729)
);

CKINVDCx20_ASAP7_75t_R g730 ( 
.A(n_560),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_581),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_614),
.Y(n_732)
);

CKINVDCx16_ASAP7_75t_R g733 ( 
.A(n_571),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_616),
.Y(n_734)
);

CKINVDCx5p33_ASAP7_75t_R g735 ( 
.A(n_502),
.Y(n_735)
);

CKINVDCx20_ASAP7_75t_R g736 ( 
.A(n_606),
.Y(n_736)
);

CKINVDCx5p33_ASAP7_75t_R g737 ( 
.A(n_506),
.Y(n_737)
);

INVxp67_ASAP7_75t_SL g738 ( 
.A(n_590),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_618),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_621),
.Y(n_740)
);

CKINVDCx20_ASAP7_75t_R g741 ( 
.A(n_636),
.Y(n_741)
);

CKINVDCx5p33_ASAP7_75t_R g742 ( 
.A(n_507),
.Y(n_742)
);

INVx3_ASAP7_75t_L g743 ( 
.A(n_543),
.Y(n_743)
);

INVxp33_ASAP7_75t_SL g744 ( 
.A(n_499),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_643),
.Y(n_745)
);

CKINVDCx20_ASAP7_75t_R g746 ( 
.A(n_576),
.Y(n_746)
);

CKINVDCx20_ASAP7_75t_R g747 ( 
.A(n_673),
.Y(n_747)
);

NAND2xp33_ASAP7_75t_R g748 ( 
.A(n_501),
.B(n_0),
.Y(n_748)
);

CKINVDCx5p33_ASAP7_75t_R g749 ( 
.A(n_509),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_644),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_649),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_652),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_663),
.Y(n_753)
);

INVxp67_ASAP7_75t_L g754 ( 
.A(n_579),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_667),
.Y(n_755)
);

INVxp67_ASAP7_75t_SL g756 ( 
.A(n_590),
.Y(n_756)
);

BUFx6f_ASAP7_75t_L g757 ( 
.A(n_518),
.Y(n_757)
);

CKINVDCx5p33_ASAP7_75t_R g758 ( 
.A(n_512),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_670),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_677),
.Y(n_760)
);

CKINVDCx5p33_ASAP7_75t_R g761 ( 
.A(n_513),
.Y(n_761)
);

INVxp33_ASAP7_75t_L g762 ( 
.A(n_682),
.Y(n_762)
);

INVx2_ASAP7_75t_L g763 ( 
.A(n_563),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_626),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_626),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_500),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_504),
.Y(n_767)
);

CKINVDCx5p33_ASAP7_75t_R g768 ( 
.A(n_514),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_508),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_515),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_533),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_536),
.Y(n_772)
);

CKINVDCx5p33_ASAP7_75t_R g773 ( 
.A(n_516),
.Y(n_773)
);

CKINVDCx5p33_ASAP7_75t_R g774 ( 
.A(n_519),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_540),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_542),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_544),
.Y(n_777)
);

CKINVDCx5p33_ASAP7_75t_R g778 ( 
.A(n_520),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_545),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_548),
.Y(n_780)
);

CKINVDCx5p33_ASAP7_75t_R g781 ( 
.A(n_523),
.Y(n_781)
);

INVxp67_ASAP7_75t_SL g782 ( 
.A(n_551),
.Y(n_782)
);

INVxp67_ASAP7_75t_SL g783 ( 
.A(n_558),
.Y(n_783)
);

NOR2xp67_ASAP7_75t_L g784 ( 
.A(n_503),
.B(n_1),
.Y(n_784)
);

AND2x2_ASAP7_75t_L g785 ( 
.A(n_711),
.B(n_580),
.Y(n_785)
);

HB1xp67_ASAP7_75t_L g786 ( 
.A(n_754),
.Y(n_786)
);

INVx2_ASAP7_75t_SL g787 ( 
.A(n_695),
.Y(n_787)
);

BUFx6f_ASAP7_75t_L g788 ( 
.A(n_757),
.Y(n_788)
);

INVx2_ASAP7_75t_SL g789 ( 
.A(n_695),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_706),
.Y(n_790)
);

AOI22xp5_ASAP7_75t_L g791 ( 
.A1(n_703),
.A2(n_662),
.B1(n_524),
.B2(n_555),
.Y(n_791)
);

NAND2x1p5_ASAP7_75t_L g792 ( 
.A(n_766),
.B(n_505),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_L g793 ( 
.A(n_735),
.B(n_651),
.Y(n_793)
);

BUFx6f_ASAP7_75t_L g794 ( 
.A(n_757),
.Y(n_794)
);

INVx2_ASAP7_75t_L g795 ( 
.A(n_757),
.Y(n_795)
);

INVx2_ASAP7_75t_L g796 ( 
.A(n_757),
.Y(n_796)
);

OAI21x1_ASAP7_75t_L g797 ( 
.A1(n_696),
.A2(n_578),
.B(n_552),
.Y(n_797)
);

AND2x2_ASAP7_75t_L g798 ( 
.A(n_716),
.B(n_668),
.Y(n_798)
);

BUFx6f_ASAP7_75t_L g799 ( 
.A(n_696),
.Y(n_799)
);

INVx2_ASAP7_75t_L g800 ( 
.A(n_697),
.Y(n_800)
);

CKINVDCx5p33_ASAP7_75t_R g801 ( 
.A(n_737),
.Y(n_801)
);

HB1xp67_ASAP7_75t_L g802 ( 
.A(n_742),
.Y(n_802)
);

CKINVDCx5p33_ASAP7_75t_R g803 ( 
.A(n_749),
.Y(n_803)
);

BUFx6f_ASAP7_75t_L g804 ( 
.A(n_697),
.Y(n_804)
);

AND2x2_ASAP7_75t_L g805 ( 
.A(n_724),
.B(n_671),
.Y(n_805)
);

BUFx3_ASAP7_75t_L g806 ( 
.A(n_725),
.Y(n_806)
);

INVx3_ASAP7_75t_L g807 ( 
.A(n_691),
.Y(n_807)
);

INVx2_ASAP7_75t_L g808 ( 
.A(n_693),
.Y(n_808)
);

OAI22x1_ASAP7_75t_R g809 ( 
.A1(n_694),
.A2(n_646),
.B1(n_521),
.B2(n_582),
.Y(n_809)
);

AND2x4_ASAP7_75t_L g810 ( 
.A(n_782),
.B(n_672),
.Y(n_810)
);

BUFx6f_ASAP7_75t_L g811 ( 
.A(n_707),
.Y(n_811)
);

OA21x2_ASAP7_75t_L g812 ( 
.A1(n_698),
.A2(n_589),
.B(n_585),
.Y(n_812)
);

BUFx6f_ASAP7_75t_L g813 ( 
.A(n_708),
.Y(n_813)
);

OAI22x1_ASAP7_75t_SL g814 ( 
.A1(n_701),
.A2(n_688),
.B1(n_685),
.B2(n_530),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_L g815 ( 
.A(n_758),
.B(n_635),
.Y(n_815)
);

HB1xp67_ASAP7_75t_L g816 ( 
.A(n_761),
.Y(n_816)
);

AND2x2_ASAP7_75t_L g817 ( 
.A(n_727),
.B(n_671),
.Y(n_817)
);

INVx4_ASAP7_75t_L g818 ( 
.A(n_768),
.Y(n_818)
);

BUFx6f_ASAP7_75t_L g819 ( 
.A(n_712),
.Y(n_819)
);

BUFx3_ASAP7_75t_L g820 ( 
.A(n_725),
.Y(n_820)
);

INVx1_ASAP7_75t_L g821 ( 
.A(n_713),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_715),
.Y(n_822)
);

INVx2_ASAP7_75t_L g823 ( 
.A(n_699),
.Y(n_823)
);

BUFx6f_ASAP7_75t_L g824 ( 
.A(n_717),
.Y(n_824)
);

OAI22xp5_ASAP7_75t_L g825 ( 
.A1(n_705),
.A2(n_539),
.B1(n_546),
.B2(n_510),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_718),
.Y(n_826)
);

AND2x2_ASAP7_75t_L g827 ( 
.A(n_738),
.B(n_683),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_767),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_L g829 ( 
.A(n_773),
.B(n_657),
.Y(n_829)
);

BUFx6f_ASAP7_75t_L g830 ( 
.A(n_720),
.Y(n_830)
);

INVx5_ASAP7_75t_L g831 ( 
.A(n_702),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_769),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_770),
.Y(n_833)
);

OAI22x1_ASAP7_75t_R g834 ( 
.A1(n_694),
.A2(n_722),
.B1(n_730),
.B2(n_701),
.Y(n_834)
);

INVxp67_ASAP7_75t_L g835 ( 
.A(n_692),
.Y(n_835)
);

INVx2_ASAP7_75t_L g836 ( 
.A(n_702),
.Y(n_836)
);

INVx5_ASAP7_75t_L g837 ( 
.A(n_710),
.Y(n_837)
);

INVx2_ASAP7_75t_SL g838 ( 
.A(n_764),
.Y(n_838)
);

INVx5_ASAP7_75t_L g839 ( 
.A(n_710),
.Y(n_839)
);

AND2x4_ASAP7_75t_L g840 ( 
.A(n_783),
.B(n_591),
.Y(n_840)
);

INVx2_ASAP7_75t_SL g841 ( 
.A(n_765),
.Y(n_841)
);

INVx4_ASAP7_75t_L g842 ( 
.A(n_774),
.Y(n_842)
);

INVx3_ASAP7_75t_L g843 ( 
.A(n_714),
.Y(n_843)
);

INVx3_ASAP7_75t_L g844 ( 
.A(n_714),
.Y(n_844)
);

BUFx12f_ASAP7_75t_L g845 ( 
.A(n_778),
.Y(n_845)
);

BUFx6f_ASAP7_75t_L g846 ( 
.A(n_719),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_771),
.Y(n_847)
);

AND2x2_ASAP7_75t_L g848 ( 
.A(n_785),
.B(n_756),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_836),
.Y(n_849)
);

INVx2_ASAP7_75t_L g850 ( 
.A(n_800),
.Y(n_850)
);

INVx3_ASAP7_75t_L g851 ( 
.A(n_846),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_L g852 ( 
.A(n_815),
.B(n_781),
.Y(n_852)
);

INVx3_ASAP7_75t_L g853 ( 
.A(n_846),
.Y(n_853)
);

BUFx3_ASAP7_75t_L g854 ( 
.A(n_806),
.Y(n_854)
);

INVx1_ASAP7_75t_SL g855 ( 
.A(n_806),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_836),
.Y(n_856)
);

OA21x2_ASAP7_75t_L g857 ( 
.A1(n_797),
.A2(n_763),
.B(n_719),
.Y(n_857)
);

INVx3_ASAP7_75t_L g858 ( 
.A(n_846),
.Y(n_858)
);

INVx2_ASAP7_75t_L g859 ( 
.A(n_800),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_L g860 ( 
.A(n_829),
.B(n_810),
.Y(n_860)
);

INVx1_ASAP7_75t_L g861 ( 
.A(n_808),
.Y(n_861)
);

INVx1_ASAP7_75t_L g862 ( 
.A(n_808),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_823),
.Y(n_863)
);

INVx2_ASAP7_75t_L g864 ( 
.A(n_843),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_L g865 ( 
.A(n_810),
.B(n_772),
.Y(n_865)
);

AND2x2_ASAP7_75t_L g866 ( 
.A(n_785),
.B(n_700),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_823),
.Y(n_867)
);

INVx2_ASAP7_75t_L g868 ( 
.A(n_843),
.Y(n_868)
);

INVx3_ASAP7_75t_L g869 ( 
.A(n_846),
.Y(n_869)
);

AND2x2_ASAP7_75t_L g870 ( 
.A(n_798),
.B(n_704),
.Y(n_870)
);

INVx2_ASAP7_75t_L g871 ( 
.A(n_843),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_807),
.Y(n_872)
);

INVx1_ASAP7_75t_L g873 ( 
.A(n_807),
.Y(n_873)
);

INVx2_ASAP7_75t_L g874 ( 
.A(n_844),
.Y(n_874)
);

BUFx6f_ASAP7_75t_L g875 ( 
.A(n_788),
.Y(n_875)
);

INVx1_ASAP7_75t_L g876 ( 
.A(n_807),
.Y(n_876)
);

HB1xp67_ASAP7_75t_L g877 ( 
.A(n_787),
.Y(n_877)
);

NOR2xp33_ASAP7_75t_L g878 ( 
.A(n_793),
.B(n_729),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_828),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_832),
.Y(n_880)
);

INVx1_ASAP7_75t_L g881 ( 
.A(n_833),
.Y(n_881)
);

INVx3_ASAP7_75t_L g882 ( 
.A(n_846),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_847),
.Y(n_883)
);

HB1xp67_ASAP7_75t_L g884 ( 
.A(n_787),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_830),
.Y(n_885)
);

INVx2_ASAP7_75t_L g886 ( 
.A(n_844),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_830),
.Y(n_887)
);

AND2x4_ASAP7_75t_L g888 ( 
.A(n_789),
.B(n_721),
.Y(n_888)
);

INVx2_ASAP7_75t_L g889 ( 
.A(n_844),
.Y(n_889)
);

BUFx6f_ASAP7_75t_L g890 ( 
.A(n_788),
.Y(n_890)
);

BUFx2_ASAP7_75t_L g891 ( 
.A(n_820),
.Y(n_891)
);

INVx1_ASAP7_75t_L g892 ( 
.A(n_790),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_821),
.Y(n_893)
);

INVx1_ASAP7_75t_L g894 ( 
.A(n_830),
.Y(n_894)
);

AND2x2_ASAP7_75t_L g895 ( 
.A(n_798),
.B(n_775),
.Y(n_895)
);

INVx2_ASAP7_75t_L g896 ( 
.A(n_799),
.Y(n_896)
);

OA21x2_ASAP7_75t_L g897 ( 
.A1(n_797),
.A2(n_763),
.B(n_776),
.Y(n_897)
);

HB1xp67_ASAP7_75t_L g898 ( 
.A(n_789),
.Y(n_898)
);

INVx1_ASAP7_75t_L g899 ( 
.A(n_830),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_L g900 ( 
.A(n_810),
.B(n_777),
.Y(n_900)
);

HB1xp67_ASAP7_75t_L g901 ( 
.A(n_820),
.Y(n_901)
);

INVx1_ASAP7_75t_L g902 ( 
.A(n_822),
.Y(n_902)
);

INVx2_ASAP7_75t_L g903 ( 
.A(n_799),
.Y(n_903)
);

INVx1_ASAP7_75t_L g904 ( 
.A(n_826),
.Y(n_904)
);

BUFx3_ASAP7_75t_L g905 ( 
.A(n_788),
.Y(n_905)
);

AND2x6_ASAP7_75t_L g906 ( 
.A(n_840),
.B(n_518),
.Y(n_906)
);

INVx1_ASAP7_75t_L g907 ( 
.A(n_811),
.Y(n_907)
);

AND2x4_ASAP7_75t_L g908 ( 
.A(n_838),
.B(n_726),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_SL g909 ( 
.A(n_792),
.B(n_723),
.Y(n_909)
);

INVx2_ASAP7_75t_L g910 ( 
.A(n_799),
.Y(n_910)
);

AND2x2_ASAP7_75t_L g911 ( 
.A(n_840),
.B(n_779),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_799),
.Y(n_912)
);

INVx2_ASAP7_75t_L g913 ( 
.A(n_799),
.Y(n_913)
);

OAI22xp5_ASAP7_75t_SL g914 ( 
.A1(n_791),
.A2(n_722),
.B1(n_736),
.B2(n_730),
.Y(n_914)
);

OAI21x1_ASAP7_75t_L g915 ( 
.A1(n_812),
.A2(n_780),
.B(n_612),
.Y(n_915)
);

AND2x2_ASAP7_75t_R g916 ( 
.A(n_809),
.B(n_834),
.Y(n_916)
);

OA21x2_ASAP7_75t_L g917 ( 
.A1(n_795),
.A2(n_619),
.B(n_608),
.Y(n_917)
);

INVx3_ASAP7_75t_L g918 ( 
.A(n_804),
.Y(n_918)
);

NAND2xp5_ASAP7_75t_L g919 ( 
.A(n_840),
.B(n_744),
.Y(n_919)
);

INVx1_ASAP7_75t_L g920 ( 
.A(n_804),
.Y(n_920)
);

INVx2_ASAP7_75t_L g921 ( 
.A(n_804),
.Y(n_921)
);

INVx1_ASAP7_75t_L g922 ( 
.A(n_804),
.Y(n_922)
);

NAND2xp5_ASAP7_75t_SL g923 ( 
.A(n_792),
.B(n_733),
.Y(n_923)
);

INVx1_ASAP7_75t_L g924 ( 
.A(n_804),
.Y(n_924)
);

INVx2_ASAP7_75t_L g925 ( 
.A(n_795),
.Y(n_925)
);

NAND2x1_ASAP7_75t_L g926 ( 
.A(n_812),
.B(n_595),
.Y(n_926)
);

INVxp67_ASAP7_75t_L g927 ( 
.A(n_786),
.Y(n_927)
);

INVx3_ASAP7_75t_L g928 ( 
.A(n_788),
.Y(n_928)
);

BUFx6f_ASAP7_75t_L g929 ( 
.A(n_794),
.Y(n_929)
);

INVx1_ASAP7_75t_L g930 ( 
.A(n_796),
.Y(n_930)
);

NOR2xp33_ASAP7_75t_L g931 ( 
.A(n_818),
.B(n_744),
.Y(n_931)
);

INVx1_ASAP7_75t_L g932 ( 
.A(n_796),
.Y(n_932)
);

OAI22xp5_ASAP7_75t_L g933 ( 
.A1(n_860),
.A2(n_792),
.B1(n_565),
.B2(n_617),
.Y(n_933)
);

INVx4_ASAP7_75t_L g934 ( 
.A(n_854),
.Y(n_934)
);

NOR2x1p5_ASAP7_75t_L g935 ( 
.A(n_919),
.B(n_845),
.Y(n_935)
);

INVx2_ASAP7_75t_L g936 ( 
.A(n_864),
.Y(n_936)
);

NAND2xp5_ASAP7_75t_L g937 ( 
.A(n_848),
.B(n_805),
.Y(n_937)
);

INVx2_ASAP7_75t_L g938 ( 
.A(n_864),
.Y(n_938)
);

INVx1_ASAP7_75t_L g939 ( 
.A(n_872),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_SL g940 ( 
.A(n_848),
.B(n_818),
.Y(n_940)
);

NOR2xp33_ASAP7_75t_SL g941 ( 
.A(n_931),
.B(n_845),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_L g942 ( 
.A(n_878),
.B(n_805),
.Y(n_942)
);

BUFx3_ASAP7_75t_L g943 ( 
.A(n_854),
.Y(n_943)
);

INVx2_ASAP7_75t_L g944 ( 
.A(n_868),
.Y(n_944)
);

AO22x2_ASAP7_75t_L g945 ( 
.A1(n_909),
.A2(n_825),
.B1(n_648),
.B2(n_554),
.Y(n_945)
);

AND2x2_ASAP7_75t_L g946 ( 
.A(n_895),
.B(n_817),
.Y(n_946)
);

INVx2_ASAP7_75t_L g947 ( 
.A(n_868),
.Y(n_947)
);

OR2x6_ASAP7_75t_L g948 ( 
.A(n_914),
.B(n_842),
.Y(n_948)
);

NAND2xp5_ASAP7_75t_SL g949 ( 
.A(n_888),
.B(n_842),
.Y(n_949)
);

INVx1_ASAP7_75t_L g950 ( 
.A(n_892),
.Y(n_950)
);

INVx1_ASAP7_75t_L g951 ( 
.A(n_892),
.Y(n_951)
);

AND3x2_ASAP7_75t_L g952 ( 
.A(n_927),
.B(n_835),
.C(n_816),
.Y(n_952)
);

BUFx3_ASAP7_75t_L g953 ( 
.A(n_891),
.Y(n_953)
);

AND2x2_ASAP7_75t_L g954 ( 
.A(n_895),
.B(n_817),
.Y(n_954)
);

INVx1_ASAP7_75t_SL g955 ( 
.A(n_855),
.Y(n_955)
);

OR2x6_ASAP7_75t_L g956 ( 
.A(n_891),
.B(n_802),
.Y(n_956)
);

INVx2_ASAP7_75t_L g957 ( 
.A(n_871),
.Y(n_957)
);

BUFx10_ASAP7_75t_L g958 ( 
.A(n_908),
.Y(n_958)
);

BUFx2_ASAP7_75t_L g959 ( 
.A(n_901),
.Y(n_959)
);

OAI22xp5_ASAP7_75t_L g960 ( 
.A1(n_852),
.A2(n_900),
.B1(n_865),
.B2(n_884),
.Y(n_960)
);

NAND2xp33_ASAP7_75t_R g961 ( 
.A(n_866),
.B(n_801),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_SL g962 ( 
.A(n_908),
.B(n_803),
.Y(n_962)
);

NAND2xp5_ASAP7_75t_SL g963 ( 
.A(n_908),
.B(n_803),
.Y(n_963)
);

INVx1_ASAP7_75t_L g964 ( 
.A(n_873),
.Y(n_964)
);

OR2x6_ASAP7_75t_L g965 ( 
.A(n_923),
.B(n_838),
.Y(n_965)
);

INVx3_ASAP7_75t_L g966 ( 
.A(n_925),
.Y(n_966)
);

HB1xp67_ASAP7_75t_L g967 ( 
.A(n_877),
.Y(n_967)
);

INVxp67_ASAP7_75t_SL g968 ( 
.A(n_851),
.Y(n_968)
);

OR2x6_ASAP7_75t_L g969 ( 
.A(n_866),
.B(n_841),
.Y(n_969)
);

INVxp33_ASAP7_75t_SL g970 ( 
.A(n_898),
.Y(n_970)
);

BUFx3_ASAP7_75t_L g971 ( 
.A(n_879),
.Y(n_971)
);

BUFx10_ASAP7_75t_L g972 ( 
.A(n_880),
.Y(n_972)
);

CKINVDCx5p33_ASAP7_75t_R g973 ( 
.A(n_881),
.Y(n_973)
);

INVx1_ASAP7_75t_L g974 ( 
.A(n_893),
.Y(n_974)
);

AOI22xp33_ASAP7_75t_L g975 ( 
.A1(n_911),
.A2(n_705),
.B1(n_812),
.B2(n_827),
.Y(n_975)
);

INVx2_ASAP7_75t_L g976 ( 
.A(n_871),
.Y(n_976)
);

XNOR2xp5_ASAP7_75t_L g977 ( 
.A(n_916),
.B(n_736),
.Y(n_977)
);

INVxp67_ASAP7_75t_SL g978 ( 
.A(n_851),
.Y(n_978)
);

NAND2xp5_ASAP7_75t_SL g979 ( 
.A(n_911),
.B(n_827),
.Y(n_979)
);

INVx2_ASAP7_75t_SL g980 ( 
.A(n_870),
.Y(n_980)
);

BUFx6f_ASAP7_75t_L g981 ( 
.A(n_905),
.Y(n_981)
);

INVx4_ASAP7_75t_L g982 ( 
.A(n_875),
.Y(n_982)
);

INVx2_ASAP7_75t_L g983 ( 
.A(n_874),
.Y(n_983)
);

BUFx6f_ASAP7_75t_L g984 ( 
.A(n_905),
.Y(n_984)
);

NAND2xp5_ASAP7_75t_L g985 ( 
.A(n_873),
.B(n_841),
.Y(n_985)
);

AND2x4_ASAP7_75t_L g986 ( 
.A(n_883),
.B(n_728),
.Y(n_986)
);

INVx4_ASAP7_75t_L g987 ( 
.A(n_875),
.Y(n_987)
);

INVx1_ASAP7_75t_SL g988 ( 
.A(n_870),
.Y(n_988)
);

AND2x2_ASAP7_75t_L g989 ( 
.A(n_893),
.B(n_762),
.Y(n_989)
);

AND2x4_ASAP7_75t_L g990 ( 
.A(n_902),
.B(n_731),
.Y(n_990)
);

NAND2xp5_ASAP7_75t_L g991 ( 
.A(n_876),
.B(n_811),
.Y(n_991)
);

BUFx4f_ASAP7_75t_L g992 ( 
.A(n_906),
.Y(n_992)
);

AO22x2_ASAP7_75t_L g993 ( 
.A1(n_904),
.A2(n_627),
.B1(n_678),
.B2(n_624),
.Y(n_993)
);

BUFx6f_ASAP7_75t_L g994 ( 
.A(n_875),
.Y(n_994)
);

NAND2xp5_ASAP7_75t_SL g995 ( 
.A(n_885),
.B(n_746),
.Y(n_995)
);

INVx1_ASAP7_75t_L g996 ( 
.A(n_876),
.Y(n_996)
);

NAND2xp5_ASAP7_75t_L g997 ( 
.A(n_887),
.B(n_811),
.Y(n_997)
);

NAND2xp5_ASAP7_75t_L g998 ( 
.A(n_894),
.B(n_811),
.Y(n_998)
);

INVx1_ASAP7_75t_L g999 ( 
.A(n_930),
.Y(n_999)
);

OAI22xp5_ASAP7_75t_L g1000 ( 
.A1(n_926),
.A2(n_637),
.B1(n_653),
.B2(n_517),
.Y(n_1000)
);

NAND2xp5_ASAP7_75t_L g1001 ( 
.A(n_899),
.B(n_813),
.Y(n_1001)
);

INVx2_ASAP7_75t_L g1002 ( 
.A(n_874),
.Y(n_1002)
);

INVx1_ASAP7_75t_L g1003 ( 
.A(n_930),
.Y(n_1003)
);

INVx1_ASAP7_75t_L g1004 ( 
.A(n_932),
.Y(n_1004)
);

BUFx4f_ASAP7_75t_L g1005 ( 
.A(n_906),
.Y(n_1005)
);

INVx1_ASAP7_75t_L g1006 ( 
.A(n_932),
.Y(n_1006)
);

NAND2xp5_ASAP7_75t_SL g1007 ( 
.A(n_861),
.B(n_747),
.Y(n_1007)
);

INVx1_ASAP7_75t_L g1008 ( 
.A(n_861),
.Y(n_1008)
);

INVx2_ASAP7_75t_SL g1009 ( 
.A(n_925),
.Y(n_1009)
);

INVx2_ASAP7_75t_SL g1010 ( 
.A(n_862),
.Y(n_1010)
);

INVx1_ASAP7_75t_L g1011 ( 
.A(n_862),
.Y(n_1011)
);

NAND2xp5_ASAP7_75t_SL g1012 ( 
.A(n_863),
.B(n_747),
.Y(n_1012)
);

INVx3_ASAP7_75t_L g1013 ( 
.A(n_928),
.Y(n_1013)
);

INVx1_ASAP7_75t_L g1014 ( 
.A(n_863),
.Y(n_1014)
);

INVx1_ASAP7_75t_L g1015 ( 
.A(n_849),
.Y(n_1015)
);

INVx3_ASAP7_75t_L g1016 ( 
.A(n_928),
.Y(n_1016)
);

INVx2_ASAP7_75t_L g1017 ( 
.A(n_886),
.Y(n_1017)
);

INVx2_ASAP7_75t_L g1018 ( 
.A(n_886),
.Y(n_1018)
);

INVx1_ASAP7_75t_L g1019 ( 
.A(n_849),
.Y(n_1019)
);

BUFx6f_ASAP7_75t_L g1020 ( 
.A(n_875),
.Y(n_1020)
);

NOR2xp33_ASAP7_75t_L g1021 ( 
.A(n_912),
.B(n_741),
.Y(n_1021)
);

INVx2_ASAP7_75t_SL g1022 ( 
.A(n_867),
.Y(n_1022)
);

INVx1_ASAP7_75t_L g1023 ( 
.A(n_856),
.Y(n_1023)
);

INVx1_ASAP7_75t_L g1024 ( 
.A(n_856),
.Y(n_1024)
);

AOI22xp33_ASAP7_75t_L g1025 ( 
.A1(n_906),
.A2(n_623),
.B1(n_629),
.B2(n_628),
.Y(n_1025)
);

INVx2_ASAP7_75t_L g1026 ( 
.A(n_889),
.Y(n_1026)
);

INVx1_ASAP7_75t_L g1027 ( 
.A(n_867),
.Y(n_1027)
);

NAND2xp5_ASAP7_75t_L g1028 ( 
.A(n_906),
.B(n_813),
.Y(n_1028)
);

INVx3_ASAP7_75t_L g1029 ( 
.A(n_928),
.Y(n_1029)
);

NAND2xp5_ASAP7_75t_SL g1030 ( 
.A(n_896),
.B(n_658),
.Y(n_1030)
);

OR2x2_ASAP7_75t_L g1031 ( 
.A(n_915),
.B(n_762),
.Y(n_1031)
);

OR2x6_ASAP7_75t_L g1032 ( 
.A(n_915),
.B(n_709),
.Y(n_1032)
);

AND2x2_ASAP7_75t_L g1033 ( 
.A(n_850),
.B(n_732),
.Y(n_1033)
);

BUFx2_ASAP7_75t_L g1034 ( 
.A(n_917),
.Y(n_1034)
);

NAND2xp5_ASAP7_75t_L g1035 ( 
.A(n_920),
.B(n_813),
.Y(n_1035)
);

BUFx8_ASAP7_75t_SL g1036 ( 
.A(n_889),
.Y(n_1036)
);

BUFx4f_ASAP7_75t_L g1037 ( 
.A(n_917),
.Y(n_1037)
);

NAND2xp5_ASAP7_75t_L g1038 ( 
.A(n_920),
.B(n_813),
.Y(n_1038)
);

AND2x4_ASAP7_75t_L g1039 ( 
.A(n_907),
.B(n_734),
.Y(n_1039)
);

INVx2_ASAP7_75t_L g1040 ( 
.A(n_850),
.Y(n_1040)
);

AND2x6_ASAP7_75t_L g1041 ( 
.A(n_896),
.B(n_518),
.Y(n_1041)
);

NAND2xp5_ASAP7_75t_L g1042 ( 
.A(n_922),
.B(n_819),
.Y(n_1042)
);

BUFx3_ASAP7_75t_L g1043 ( 
.A(n_917),
.Y(n_1043)
);

NAND2xp5_ASAP7_75t_L g1044 ( 
.A(n_922),
.B(n_819),
.Y(n_1044)
);

NAND2xp5_ASAP7_75t_SL g1045 ( 
.A(n_903),
.B(n_666),
.Y(n_1045)
);

NAND2xp5_ASAP7_75t_SL g1046 ( 
.A(n_903),
.B(n_525),
.Y(n_1046)
);

HB1xp67_ASAP7_75t_L g1047 ( 
.A(n_917),
.Y(n_1047)
);

INVx1_ASAP7_75t_L g1048 ( 
.A(n_859),
.Y(n_1048)
);

NAND2xp5_ASAP7_75t_L g1049 ( 
.A(n_924),
.B(n_819),
.Y(n_1049)
);

INVx1_ASAP7_75t_L g1050 ( 
.A(n_859),
.Y(n_1050)
);

INVx3_ASAP7_75t_L g1051 ( 
.A(n_897),
.Y(n_1051)
);

INVx2_ASAP7_75t_L g1052 ( 
.A(n_851),
.Y(n_1052)
);

AND2x2_ASAP7_75t_L g1053 ( 
.A(n_897),
.B(n_739),
.Y(n_1053)
);

AND2x2_ASAP7_75t_L g1054 ( 
.A(n_897),
.B(n_740),
.Y(n_1054)
);

INVx4_ASAP7_75t_L g1055 ( 
.A(n_875),
.Y(n_1055)
);

OR2x6_ASAP7_75t_L g1056 ( 
.A(n_926),
.B(n_784),
.Y(n_1056)
);

CKINVDCx20_ASAP7_75t_R g1057 ( 
.A(n_910),
.Y(n_1057)
);

NAND2xp33_ASAP7_75t_L g1058 ( 
.A(n_913),
.B(n_563),
.Y(n_1058)
);

INVx2_ASAP7_75t_L g1059 ( 
.A(n_853),
.Y(n_1059)
);

NAND2xp5_ASAP7_75t_L g1060 ( 
.A(n_942),
.B(n_921),
.Y(n_1060)
);

INVx1_ASAP7_75t_L g1061 ( 
.A(n_939),
.Y(n_1061)
);

NAND2xp5_ASAP7_75t_SL g1062 ( 
.A(n_937),
.B(n_890),
.Y(n_1062)
);

NAND2xp5_ASAP7_75t_L g1063 ( 
.A(n_946),
.B(n_921),
.Y(n_1063)
);

INVx2_ASAP7_75t_L g1064 ( 
.A(n_939),
.Y(n_1064)
);

NAND2xp5_ASAP7_75t_L g1065 ( 
.A(n_954),
.B(n_853),
.Y(n_1065)
);

NOR2x1p5_ASAP7_75t_L g1066 ( 
.A(n_953),
.B(n_814),
.Y(n_1066)
);

NAND2xp5_ASAP7_75t_L g1067 ( 
.A(n_950),
.B(n_858),
.Y(n_1067)
);

NAND2xp5_ASAP7_75t_L g1068 ( 
.A(n_951),
.B(n_858),
.Y(n_1068)
);

NAND2xp5_ASAP7_75t_L g1069 ( 
.A(n_974),
.B(n_858),
.Y(n_1069)
);

INVxp67_ASAP7_75t_L g1070 ( 
.A(n_967),
.Y(n_1070)
);

INVx2_ASAP7_75t_SL g1071 ( 
.A(n_955),
.Y(n_1071)
);

NAND2xp5_ASAP7_75t_L g1072 ( 
.A(n_1010),
.B(n_1022),
.Y(n_1072)
);

INVx1_ASAP7_75t_SL g1073 ( 
.A(n_988),
.Y(n_1073)
);

NAND2xp5_ASAP7_75t_L g1074 ( 
.A(n_960),
.B(n_869),
.Y(n_1074)
);

NAND2xp5_ASAP7_75t_L g1075 ( 
.A(n_989),
.B(n_869),
.Y(n_1075)
);

CKINVDCx5p33_ASAP7_75t_R g1076 ( 
.A(n_961),
.Y(n_1076)
);

INVx8_ASAP7_75t_L g1077 ( 
.A(n_956),
.Y(n_1077)
);

AOI22xp5_ASAP7_75t_L g1078 ( 
.A1(n_940),
.A2(n_882),
.B1(n_918),
.B2(n_869),
.Y(n_1078)
);

NOR2xp33_ASAP7_75t_L g1079 ( 
.A(n_970),
.B(n_882),
.Y(n_1079)
);

NAND2xp5_ASAP7_75t_L g1080 ( 
.A(n_975),
.B(n_882),
.Y(n_1080)
);

INVx1_ASAP7_75t_L g1081 ( 
.A(n_964),
.Y(n_1081)
);

INVx2_ASAP7_75t_SL g1082 ( 
.A(n_969),
.Y(n_1082)
);

NAND2xp5_ASAP7_75t_L g1083 ( 
.A(n_980),
.B(n_918),
.Y(n_1083)
);

INVxp67_ASAP7_75t_L g1084 ( 
.A(n_1021),
.Y(n_1084)
);

NAND2xp5_ASAP7_75t_SL g1085 ( 
.A(n_958),
.B(n_890),
.Y(n_1085)
);

NAND2xp5_ASAP7_75t_L g1086 ( 
.A(n_979),
.B(n_890),
.Y(n_1086)
);

NAND2xp5_ASAP7_75t_L g1087 ( 
.A(n_1008),
.B(n_890),
.Y(n_1087)
);

NAND2xp5_ASAP7_75t_L g1088 ( 
.A(n_1011),
.B(n_929),
.Y(n_1088)
);

AND2x2_ASAP7_75t_L g1089 ( 
.A(n_969),
.B(n_684),
.Y(n_1089)
);

OAI22xp5_ASAP7_75t_L g1090 ( 
.A1(n_945),
.A2(n_564),
.B1(n_568),
.B2(n_562),
.Y(n_1090)
);

NAND2xp5_ASAP7_75t_L g1091 ( 
.A(n_1014),
.B(n_929),
.Y(n_1091)
);

NAND2xp5_ASAP7_75t_L g1092 ( 
.A(n_1027),
.B(n_929),
.Y(n_1092)
);

NAND2xp5_ASAP7_75t_SL g1093 ( 
.A(n_973),
.B(n_929),
.Y(n_1093)
);

INVx1_ASAP7_75t_L g1094 ( 
.A(n_996),
.Y(n_1094)
);

NAND2xp5_ASAP7_75t_L g1095 ( 
.A(n_1027),
.B(n_929),
.Y(n_1095)
);

AND2x4_ASAP7_75t_L g1096 ( 
.A(n_934),
.B(n_745),
.Y(n_1096)
);

NAND2xp5_ASAP7_75t_SL g1097 ( 
.A(n_933),
.B(n_529),
.Y(n_1097)
);

INVx1_ASAP7_75t_L g1098 ( 
.A(n_996),
.Y(n_1098)
);

NAND2xp5_ASAP7_75t_L g1099 ( 
.A(n_1053),
.B(n_630),
.Y(n_1099)
);

INVx1_ASAP7_75t_L g1100 ( 
.A(n_1015),
.Y(n_1100)
);

BUFx6f_ASAP7_75t_L g1101 ( 
.A(n_981),
.Y(n_1101)
);

OR2x2_ASAP7_75t_L g1102 ( 
.A(n_959),
.B(n_750),
.Y(n_1102)
);

NAND2xp5_ASAP7_75t_L g1103 ( 
.A(n_1054),
.B(n_631),
.Y(n_1103)
);

NAND2xp5_ASAP7_75t_L g1104 ( 
.A(n_1051),
.B(n_1019),
.Y(n_1104)
);

AOI22xp33_ASAP7_75t_L g1105 ( 
.A1(n_1031),
.A2(n_639),
.B1(n_654),
.B2(n_638),
.Y(n_1105)
);

NAND2xp5_ASAP7_75t_L g1106 ( 
.A(n_1051),
.B(n_669),
.Y(n_1106)
);

INVx2_ASAP7_75t_L g1107 ( 
.A(n_1023),
.Y(n_1107)
);

INVx2_ASAP7_75t_L g1108 ( 
.A(n_1023),
.Y(n_1108)
);

INVx1_ASAP7_75t_L g1109 ( 
.A(n_1024),
.Y(n_1109)
);

NAND2x1_ASAP7_75t_L g1110 ( 
.A(n_982),
.B(n_857),
.Y(n_1110)
);

NOR2xp33_ASAP7_75t_L g1111 ( 
.A(n_1000),
.B(n_584),
.Y(n_1111)
);

NAND2xp5_ASAP7_75t_L g1112 ( 
.A(n_985),
.B(n_1009),
.Y(n_1112)
);

NAND2xp5_ASAP7_75t_L g1113 ( 
.A(n_1033),
.B(n_675),
.Y(n_1113)
);

INVx2_ASAP7_75t_L g1114 ( 
.A(n_1048),
.Y(n_1114)
);

INVx1_ASAP7_75t_L g1115 ( 
.A(n_999),
.Y(n_1115)
);

NAND2xp5_ASAP7_75t_L g1116 ( 
.A(n_1003),
.B(n_687),
.Y(n_1116)
);

INVx2_ASAP7_75t_L g1117 ( 
.A(n_1048),
.Y(n_1117)
);

NAND2xp5_ASAP7_75t_L g1118 ( 
.A(n_1004),
.B(n_689),
.Y(n_1118)
);

NAND2xp5_ASAP7_75t_SL g1119 ( 
.A(n_971),
.B(n_531),
.Y(n_1119)
);

INVx2_ASAP7_75t_L g1120 ( 
.A(n_1050),
.Y(n_1120)
);

NAND2xp5_ASAP7_75t_SL g1121 ( 
.A(n_972),
.B(n_532),
.Y(n_1121)
);

NAND2xp5_ASAP7_75t_L g1122 ( 
.A(n_1006),
.B(n_897),
.Y(n_1122)
);

NOR2xp33_ASAP7_75t_L g1123 ( 
.A(n_962),
.B(n_592),
.Y(n_1123)
);

NAND3xp33_ASAP7_75t_L g1124 ( 
.A(n_1030),
.B(n_857),
.C(n_748),
.Y(n_1124)
);

NAND2xp5_ASAP7_75t_L g1125 ( 
.A(n_1050),
.B(n_857),
.Y(n_1125)
);

NAND2xp5_ASAP7_75t_SL g1126 ( 
.A(n_972),
.B(n_535),
.Y(n_1126)
);

AND2x2_ASAP7_75t_L g1127 ( 
.A(n_956),
.B(n_684),
.Y(n_1127)
);

NOR2xp33_ASAP7_75t_L g1128 ( 
.A(n_963),
.B(n_593),
.Y(n_1128)
);

NAND2xp5_ASAP7_75t_SL g1129 ( 
.A(n_949),
.B(n_537),
.Y(n_1129)
);

INVx1_ASAP7_75t_L g1130 ( 
.A(n_1039),
.Y(n_1130)
);

INVxp67_ASAP7_75t_L g1131 ( 
.A(n_1007),
.Y(n_1131)
);

NOR2xp33_ASAP7_75t_L g1132 ( 
.A(n_1045),
.B(n_594),
.Y(n_1132)
);

NAND2xp5_ASAP7_75t_L g1133 ( 
.A(n_986),
.B(n_857),
.Y(n_1133)
);

A2O1A1Ixp33_ASAP7_75t_L g1134 ( 
.A1(n_1037),
.A2(n_549),
.B(n_550),
.C(n_538),
.Y(n_1134)
);

INVx1_ASAP7_75t_L g1135 ( 
.A(n_1039),
.Y(n_1135)
);

INVx1_ASAP7_75t_L g1136 ( 
.A(n_1040),
.Y(n_1136)
);

OA22x2_ASAP7_75t_L g1137 ( 
.A1(n_948),
.A2(n_599),
.B1(n_600),
.B2(n_597),
.Y(n_1137)
);

INVx2_ASAP7_75t_L g1138 ( 
.A(n_966),
.Y(n_1138)
);

NAND2xp5_ASAP7_75t_L g1139 ( 
.A(n_986),
.B(n_553),
.Y(n_1139)
);

INVx2_ASAP7_75t_SL g1140 ( 
.A(n_990),
.Y(n_1140)
);

O2A1O1Ixp5_ASAP7_75t_L g1141 ( 
.A1(n_1037),
.A2(n_752),
.B(n_753),
.C(n_751),
.Y(n_1141)
);

NAND2xp5_ASAP7_75t_SL g1142 ( 
.A(n_941),
.B(n_556),
.Y(n_1142)
);

INVx1_ASAP7_75t_L g1143 ( 
.A(n_936),
.Y(n_1143)
);

AOI22x1_ASAP7_75t_L g1144 ( 
.A1(n_1047),
.A2(n_1034),
.B1(n_968),
.B2(n_978),
.Y(n_1144)
);

NAND2xp5_ASAP7_75t_SL g1145 ( 
.A(n_981),
.B(n_557),
.Y(n_1145)
);

NOR2xp33_ASAP7_75t_L g1146 ( 
.A(n_1012),
.B(n_603),
.Y(n_1146)
);

NAND2xp5_ASAP7_75t_L g1147 ( 
.A(n_966),
.B(n_561),
.Y(n_1147)
);

NAND2xp5_ASAP7_75t_L g1148 ( 
.A(n_938),
.B(n_566),
.Y(n_1148)
);

OAI22xp33_ASAP7_75t_L g1149 ( 
.A1(n_965),
.A2(n_748),
.B1(n_528),
.B2(n_547),
.Y(n_1149)
);

NOR2xp33_ASAP7_75t_L g1150 ( 
.A(n_1057),
.B(n_609),
.Y(n_1150)
);

NAND2xp5_ASAP7_75t_L g1151 ( 
.A(n_944),
.B(n_569),
.Y(n_1151)
);

AOI22xp5_ASAP7_75t_L g1152 ( 
.A1(n_1056),
.A2(n_573),
.B1(n_574),
.B2(n_570),
.Y(n_1152)
);

NAND2xp5_ASAP7_75t_SL g1153 ( 
.A(n_981),
.B(n_984),
.Y(n_1153)
);

NAND2xp5_ASAP7_75t_L g1154 ( 
.A(n_947),
.B(n_583),
.Y(n_1154)
);

INVx1_ASAP7_75t_L g1155 ( 
.A(n_957),
.Y(n_1155)
);

INVx2_ASAP7_75t_L g1156 ( 
.A(n_976),
.Y(n_1156)
);

BUFx6f_ASAP7_75t_L g1157 ( 
.A(n_984),
.Y(n_1157)
);

INVx1_ASAP7_75t_L g1158 ( 
.A(n_983),
.Y(n_1158)
);

BUFx6f_ASAP7_75t_L g1159 ( 
.A(n_984),
.Y(n_1159)
);

NOR2xp33_ASAP7_75t_R g1160 ( 
.A(n_943),
.B(n_588),
.Y(n_1160)
);

NAND2xp5_ASAP7_75t_L g1161 ( 
.A(n_1002),
.B(n_596),
.Y(n_1161)
);

AND2x2_ASAP7_75t_L g1162 ( 
.A(n_965),
.B(n_755),
.Y(n_1162)
);

NOR2xp33_ASAP7_75t_L g1163 ( 
.A(n_995),
.B(n_610),
.Y(n_1163)
);

NOR2xp67_ASAP7_75t_L g1164 ( 
.A(n_1017),
.B(n_759),
.Y(n_1164)
);

NAND2xp5_ASAP7_75t_L g1165 ( 
.A(n_1018),
.B(n_598),
.Y(n_1165)
);

OR2x6_ASAP7_75t_L g1166 ( 
.A(n_948),
.B(n_760),
.Y(n_1166)
);

NAND2xp5_ASAP7_75t_L g1167 ( 
.A(n_1026),
.B(n_602),
.Y(n_1167)
);

NAND2xp5_ASAP7_75t_L g1168 ( 
.A(n_1013),
.B(n_1016),
.Y(n_1168)
);

AOI22xp33_ASAP7_75t_L g1169 ( 
.A1(n_945),
.A2(n_676),
.B1(n_528),
.B2(n_547),
.Y(n_1169)
);

NAND2xp5_ASAP7_75t_L g1170 ( 
.A(n_1013),
.B(n_604),
.Y(n_1170)
);

NAND2xp5_ASAP7_75t_SL g1171 ( 
.A(n_992),
.B(n_607),
.Y(n_1171)
);

INVx1_ASAP7_75t_L g1172 ( 
.A(n_1016),
.Y(n_1172)
);

INVx1_ASAP7_75t_L g1173 ( 
.A(n_1029),
.Y(n_1173)
);

NOR2xp33_ASAP7_75t_SL g1174 ( 
.A(n_1005),
.B(n_683),
.Y(n_1174)
);

AND2x2_ASAP7_75t_L g1175 ( 
.A(n_993),
.B(n_935),
.Y(n_1175)
);

AOI22xp5_ASAP7_75t_L g1176 ( 
.A1(n_1046),
.A2(n_615),
.B1(n_620),
.B2(n_611),
.Y(n_1176)
);

INVxp67_ASAP7_75t_SL g1177 ( 
.A(n_994),
.Y(n_1177)
);

NAND2xp5_ASAP7_75t_L g1178 ( 
.A(n_1029),
.B(n_632),
.Y(n_1178)
);

INVxp67_ASAP7_75t_L g1179 ( 
.A(n_1036),
.Y(n_1179)
);

AND2x2_ASAP7_75t_L g1180 ( 
.A(n_993),
.B(n_743),
.Y(n_1180)
);

NAND2xp5_ASAP7_75t_L g1181 ( 
.A(n_1043),
.B(n_641),
.Y(n_1181)
);

INVxp33_ASAP7_75t_SL g1182 ( 
.A(n_977),
.Y(n_1182)
);

INVx2_ASAP7_75t_SL g1183 ( 
.A(n_952),
.Y(n_1183)
);

NOR2xp33_ASAP7_75t_L g1184 ( 
.A(n_1052),
.B(n_613),
.Y(n_1184)
);

AOI22xp33_ASAP7_75t_L g1185 ( 
.A1(n_1032),
.A2(n_676),
.B1(n_547),
.B2(n_528),
.Y(n_1185)
);

CKINVDCx5p33_ASAP7_75t_R g1186 ( 
.A(n_1032),
.Y(n_1186)
);

OAI22xp33_ASAP7_75t_L g1187 ( 
.A1(n_1028),
.A2(n_633),
.B1(n_634),
.B2(n_625),
.Y(n_1187)
);

INVx2_ASAP7_75t_L g1188 ( 
.A(n_1059),
.Y(n_1188)
);

INVx2_ASAP7_75t_SL g1189 ( 
.A(n_997),
.Y(n_1189)
);

NOR2xp33_ASAP7_75t_L g1190 ( 
.A(n_991),
.B(n_640),
.Y(n_1190)
);

NAND2xp5_ASAP7_75t_SL g1191 ( 
.A(n_994),
.B(n_655),
.Y(n_1191)
);

NAND2xp5_ASAP7_75t_L g1192 ( 
.A(n_982),
.B(n_656),
.Y(n_1192)
);

AOI22xp33_ASAP7_75t_L g1193 ( 
.A1(n_1025),
.A2(n_1058),
.B1(n_998),
.B2(n_1001),
.Y(n_1193)
);

BUFx6f_ASAP7_75t_L g1194 ( 
.A(n_1020),
.Y(n_1194)
);

NAND2xp5_ASAP7_75t_L g1195 ( 
.A(n_987),
.B(n_661),
.Y(n_1195)
);

NAND2xp33_ASAP7_75t_L g1196 ( 
.A(n_1020),
.B(n_676),
.Y(n_1196)
);

AOI22xp33_ASAP7_75t_L g1197 ( 
.A1(n_1035),
.A2(n_676),
.B1(n_824),
.B2(n_819),
.Y(n_1197)
);

OR2x2_ASAP7_75t_L g1198 ( 
.A(n_1038),
.B(n_1042),
.Y(n_1198)
);

INVx2_ASAP7_75t_L g1199 ( 
.A(n_1044),
.Y(n_1199)
);

OR2x2_ASAP7_75t_L g1200 ( 
.A(n_1049),
.B(n_642),
.Y(n_1200)
);

BUFx6f_ASAP7_75t_L g1201 ( 
.A(n_1020),
.Y(n_1201)
);

NAND2xp33_ASAP7_75t_L g1202 ( 
.A(n_1041),
.B(n_676),
.Y(n_1202)
);

NAND2xp5_ASAP7_75t_L g1203 ( 
.A(n_1055),
.B(n_674),
.Y(n_1203)
);

NAND2xp5_ASAP7_75t_L g1204 ( 
.A(n_1041),
.B(n_679),
.Y(n_1204)
);

INVx1_ASAP7_75t_L g1205 ( 
.A(n_1041),
.Y(n_1205)
);

INVx2_ASAP7_75t_L g1206 ( 
.A(n_1041),
.Y(n_1206)
);

NAND2xp33_ASAP7_75t_L g1207 ( 
.A(n_937),
.B(n_681),
.Y(n_1207)
);

NOR2xp33_ASAP7_75t_L g1208 ( 
.A(n_942),
.B(n_645),
.Y(n_1208)
);

NAND2xp5_ASAP7_75t_L g1209 ( 
.A(n_942),
.B(n_686),
.Y(n_1209)
);

AOI22xp5_ASAP7_75t_L g1210 ( 
.A1(n_942),
.A2(n_690),
.B1(n_824),
.B2(n_647),
.Y(n_1210)
);

INVx3_ASAP7_75t_L g1211 ( 
.A(n_1013),
.Y(n_1211)
);

INVx2_ASAP7_75t_L g1212 ( 
.A(n_939),
.Y(n_1212)
);

INVx1_ASAP7_75t_L g1213 ( 
.A(n_939),
.Y(n_1213)
);

INVx2_ASAP7_75t_SL g1214 ( 
.A(n_955),
.Y(n_1214)
);

INVxp67_ASAP7_75t_L g1215 ( 
.A(n_967),
.Y(n_1215)
);

OAI22xp33_ASAP7_75t_L g1216 ( 
.A1(n_942),
.A2(n_659),
.B1(n_664),
.B2(n_650),
.Y(n_1216)
);

NAND2xp5_ASAP7_75t_L g1217 ( 
.A(n_942),
.B(n_665),
.Y(n_1217)
);

BUFx6f_ASAP7_75t_L g1218 ( 
.A(n_981),
.Y(n_1218)
);

NAND2xp5_ASAP7_75t_L g1219 ( 
.A(n_942),
.B(n_794),
.Y(n_1219)
);

NAND2xp5_ASAP7_75t_SL g1220 ( 
.A(n_937),
.B(n_794),
.Y(n_1220)
);

NAND2xp5_ASAP7_75t_L g1221 ( 
.A(n_942),
.B(n_794),
.Y(n_1221)
);

NOR2xp33_ASAP7_75t_L g1222 ( 
.A(n_942),
.B(n_3),
.Y(n_1222)
);

NAND2xp5_ASAP7_75t_L g1223 ( 
.A(n_942),
.B(n_831),
.Y(n_1223)
);

INVx1_ASAP7_75t_L g1224 ( 
.A(n_939),
.Y(n_1224)
);

NAND2xp5_ASAP7_75t_SL g1225 ( 
.A(n_937),
.B(n_839),
.Y(n_1225)
);

OAI22xp5_ASAP7_75t_L g1226 ( 
.A1(n_937),
.A2(n_743),
.B1(n_837),
.B2(n_831),
.Y(n_1226)
);

O2A1O1Ixp33_ASAP7_75t_L g1227 ( 
.A1(n_937),
.A2(n_5),
.B(n_3),
.C(n_4),
.Y(n_1227)
);

BUFx3_ASAP7_75t_L g1228 ( 
.A(n_1057),
.Y(n_1228)
);

AOI22xp33_ASAP7_75t_L g1229 ( 
.A1(n_1031),
.A2(n_837),
.B1(n_839),
.B2(n_831),
.Y(n_1229)
);

INVx1_ASAP7_75t_L g1230 ( 
.A(n_1061),
.Y(n_1230)
);

BUFx3_ASAP7_75t_L g1231 ( 
.A(n_1228),
.Y(n_1231)
);

INVx1_ASAP7_75t_L g1232 ( 
.A(n_1081),
.Y(n_1232)
);

NAND2xp5_ASAP7_75t_SL g1233 ( 
.A(n_1071),
.B(n_831),
.Y(n_1233)
);

AOI22xp33_ASAP7_75t_L g1234 ( 
.A1(n_1222),
.A2(n_839),
.B1(n_837),
.B2(n_7),
.Y(n_1234)
);

AND2x4_ASAP7_75t_L g1235 ( 
.A(n_1140),
.B(n_211),
.Y(n_1235)
);

INVx3_ASAP7_75t_L g1236 ( 
.A(n_1194),
.Y(n_1236)
);

NAND2xp5_ASAP7_75t_L g1237 ( 
.A(n_1208),
.B(n_5),
.Y(n_1237)
);

BUFx2_ASAP7_75t_L g1238 ( 
.A(n_1214),
.Y(n_1238)
);

INVx2_ASAP7_75t_L g1239 ( 
.A(n_1064),
.Y(n_1239)
);

INVx1_ASAP7_75t_L g1240 ( 
.A(n_1094),
.Y(n_1240)
);

NOR2xp33_ASAP7_75t_L g1241 ( 
.A(n_1084),
.B(n_6),
.Y(n_1241)
);

INVx2_ASAP7_75t_SL g1242 ( 
.A(n_1102),
.Y(n_1242)
);

INVx1_ASAP7_75t_L g1243 ( 
.A(n_1098),
.Y(n_1243)
);

NAND2xp5_ASAP7_75t_SL g1244 ( 
.A(n_1073),
.B(n_837),
.Y(n_1244)
);

BUFx6f_ASAP7_75t_L g1245 ( 
.A(n_1194),
.Y(n_1245)
);

AND2x2_ASAP7_75t_L g1246 ( 
.A(n_1073),
.B(n_6),
.Y(n_1246)
);

INVx1_ASAP7_75t_L g1247 ( 
.A(n_1213),
.Y(n_1247)
);

NOR3xp33_ASAP7_75t_SL g1248 ( 
.A(n_1076),
.B(n_7),
.C(n_8),
.Y(n_1248)
);

INVx3_ASAP7_75t_SL g1249 ( 
.A(n_1077),
.Y(n_1249)
);

INVxp67_ASAP7_75t_SL g1250 ( 
.A(n_1194),
.Y(n_1250)
);

INVx1_ASAP7_75t_L g1251 ( 
.A(n_1224),
.Y(n_1251)
);

NAND2xp5_ASAP7_75t_L g1252 ( 
.A(n_1112),
.B(n_8),
.Y(n_1252)
);

OAI22xp5_ASAP7_75t_L g1253 ( 
.A1(n_1100),
.A2(n_839),
.B1(n_213),
.B2(n_217),
.Y(n_1253)
);

BUFx2_ASAP7_75t_L g1254 ( 
.A(n_1070),
.Y(n_1254)
);

INVx1_ASAP7_75t_L g1255 ( 
.A(n_1212),
.Y(n_1255)
);

INVx1_ASAP7_75t_L g1256 ( 
.A(n_1109),
.Y(n_1256)
);

NAND2xp5_ASAP7_75t_L g1257 ( 
.A(n_1217),
.B(n_9),
.Y(n_1257)
);

NOR2xp33_ASAP7_75t_L g1258 ( 
.A(n_1131),
.B(n_10),
.Y(n_1258)
);

NAND2xp5_ASAP7_75t_L g1259 ( 
.A(n_1209),
.B(n_10),
.Y(n_1259)
);

BUFx3_ASAP7_75t_L g1260 ( 
.A(n_1077),
.Y(n_1260)
);

HB1xp67_ASAP7_75t_L g1261 ( 
.A(n_1215),
.Y(n_1261)
);

OAI22xp5_ASAP7_75t_SL g1262 ( 
.A1(n_1182),
.A2(n_13),
.B1(n_11),
.B2(n_12),
.Y(n_1262)
);

OR2x2_ASAP7_75t_L g1263 ( 
.A(n_1200),
.B(n_11),
.Y(n_1263)
);

NOR2xp33_ASAP7_75t_L g1264 ( 
.A(n_1150),
.B(n_14),
.Y(n_1264)
);

INVx5_ASAP7_75t_L g1265 ( 
.A(n_1201),
.Y(n_1265)
);

INVx2_ASAP7_75t_L g1266 ( 
.A(n_1107),
.Y(n_1266)
);

INVx2_ASAP7_75t_L g1267 ( 
.A(n_1108),
.Y(n_1267)
);

NAND2xp5_ASAP7_75t_L g1268 ( 
.A(n_1060),
.B(n_14),
.Y(n_1268)
);

INVx2_ASAP7_75t_L g1269 ( 
.A(n_1114),
.Y(n_1269)
);

INVx1_ASAP7_75t_L g1270 ( 
.A(n_1117),
.Y(n_1270)
);

NOR3xp33_ASAP7_75t_SL g1271 ( 
.A(n_1186),
.B(n_15),
.C(n_16),
.Y(n_1271)
);

CKINVDCx5p33_ASAP7_75t_R g1272 ( 
.A(n_1077),
.Y(n_1272)
);

INVxp67_ASAP7_75t_L g1273 ( 
.A(n_1162),
.Y(n_1273)
);

CKINVDCx5p33_ASAP7_75t_R g1274 ( 
.A(n_1160),
.Y(n_1274)
);

NAND2xp5_ASAP7_75t_SL g1275 ( 
.A(n_1101),
.B(n_839),
.Y(n_1275)
);

CKINVDCx5p33_ASAP7_75t_R g1276 ( 
.A(n_1179),
.Y(n_1276)
);

BUFx3_ASAP7_75t_L g1277 ( 
.A(n_1082),
.Y(n_1277)
);

O2A1O1Ixp33_ASAP7_75t_L g1278 ( 
.A1(n_1216),
.A2(n_17),
.B(n_15),
.C(n_16),
.Y(n_1278)
);

INVx1_ASAP7_75t_L g1279 ( 
.A(n_1120),
.Y(n_1279)
);

INVx1_ASAP7_75t_L g1280 ( 
.A(n_1115),
.Y(n_1280)
);

NAND2xp5_ASAP7_75t_L g1281 ( 
.A(n_1189),
.B(n_17),
.Y(n_1281)
);

INVx1_ASAP7_75t_L g1282 ( 
.A(n_1136),
.Y(n_1282)
);

AND2x4_ASAP7_75t_L g1283 ( 
.A(n_1130),
.B(n_212),
.Y(n_1283)
);

AOI22xp33_ASAP7_75t_L g1284 ( 
.A1(n_1111),
.A2(n_1124),
.B1(n_1132),
.B2(n_1169),
.Y(n_1284)
);

NAND2xp5_ASAP7_75t_L g1285 ( 
.A(n_1199),
.B(n_18),
.Y(n_1285)
);

AOI22xp33_ASAP7_75t_L g1286 ( 
.A1(n_1124),
.A2(n_20),
.B1(n_18),
.B2(n_19),
.Y(n_1286)
);

INVx1_ASAP7_75t_L g1287 ( 
.A(n_1063),
.Y(n_1287)
);

BUFx12f_ASAP7_75t_L g1288 ( 
.A(n_1183),
.Y(n_1288)
);

INVx3_ASAP7_75t_L g1289 ( 
.A(n_1201),
.Y(n_1289)
);

NOR2x2_ASAP7_75t_L g1290 ( 
.A(n_1166),
.B(n_19),
.Y(n_1290)
);

OAI22xp33_ASAP7_75t_L g1291 ( 
.A1(n_1174),
.A2(n_22),
.B1(n_20),
.B2(n_21),
.Y(n_1291)
);

BUFx8_ASAP7_75t_L g1292 ( 
.A(n_1089),
.Y(n_1292)
);

NOR2xp33_ASAP7_75t_L g1293 ( 
.A(n_1072),
.B(n_22),
.Y(n_1293)
);

NAND2xp5_ASAP7_75t_L g1294 ( 
.A(n_1075),
.B(n_24),
.Y(n_1294)
);

INVx2_ASAP7_75t_SL g1295 ( 
.A(n_1127),
.Y(n_1295)
);

OAI22xp5_ASAP7_75t_L g1296 ( 
.A1(n_1133),
.A2(n_219),
.B1(n_220),
.B2(n_218),
.Y(n_1296)
);

AOI22x1_ASAP7_75t_L g1297 ( 
.A1(n_1172),
.A2(n_223),
.B1(n_227),
.B2(n_222),
.Y(n_1297)
);

OR2x2_ASAP7_75t_L g1298 ( 
.A(n_1139),
.B(n_24),
.Y(n_1298)
);

AOI22xp5_ASAP7_75t_L g1299 ( 
.A1(n_1207),
.A2(n_232),
.B1(n_233),
.B2(n_230),
.Y(n_1299)
);

HB1xp67_ASAP7_75t_L g1300 ( 
.A(n_1101),
.Y(n_1300)
);

INVx1_ASAP7_75t_L g1301 ( 
.A(n_1143),
.Y(n_1301)
);

INVx1_ASAP7_75t_L g1302 ( 
.A(n_1155),
.Y(n_1302)
);

NAND2xp5_ASAP7_75t_SL g1303 ( 
.A(n_1157),
.B(n_235),
.Y(n_1303)
);

INVx3_ASAP7_75t_L g1304 ( 
.A(n_1201),
.Y(n_1304)
);

NAND2xp5_ASAP7_75t_L g1305 ( 
.A(n_1190),
.B(n_25),
.Y(n_1305)
);

NAND2xp5_ASAP7_75t_L g1306 ( 
.A(n_1065),
.B(n_25),
.Y(n_1306)
);

NAND2xp5_ASAP7_75t_SL g1307 ( 
.A(n_1157),
.B(n_236),
.Y(n_1307)
);

INVx2_ASAP7_75t_L g1308 ( 
.A(n_1138),
.Y(n_1308)
);

INVx2_ASAP7_75t_L g1309 ( 
.A(n_1156),
.Y(n_1309)
);

NAND2xp5_ASAP7_75t_SL g1310 ( 
.A(n_1157),
.B(n_237),
.Y(n_1310)
);

INVx1_ASAP7_75t_L g1311 ( 
.A(n_1158),
.Y(n_1311)
);

NOR2xp33_ASAP7_75t_L g1312 ( 
.A(n_1146),
.B(n_26),
.Y(n_1312)
);

INVx2_ASAP7_75t_L g1313 ( 
.A(n_1211),
.Y(n_1313)
);

AND2x2_ASAP7_75t_L g1314 ( 
.A(n_1180),
.B(n_27),
.Y(n_1314)
);

INVx1_ASAP7_75t_L g1315 ( 
.A(n_1067),
.Y(n_1315)
);

AOI22xp33_ASAP7_75t_L g1316 ( 
.A1(n_1097),
.A2(n_31),
.B1(n_28),
.B2(n_30),
.Y(n_1316)
);

NAND2xp5_ASAP7_75t_L g1317 ( 
.A(n_1198),
.B(n_31),
.Y(n_1317)
);

BUFx3_ASAP7_75t_L g1318 ( 
.A(n_1159),
.Y(n_1318)
);

INVx1_ASAP7_75t_L g1319 ( 
.A(n_1068),
.Y(n_1319)
);

NAND2xp5_ASAP7_75t_L g1320 ( 
.A(n_1113),
.B(n_32),
.Y(n_1320)
);

NAND2xp5_ASAP7_75t_L g1321 ( 
.A(n_1079),
.B(n_32),
.Y(n_1321)
);

INVx2_ASAP7_75t_L g1322 ( 
.A(n_1211),
.Y(n_1322)
);

NAND3xp33_ASAP7_75t_SL g1323 ( 
.A(n_1163),
.B(n_33),
.C(n_34),
.Y(n_1323)
);

NAND2xp5_ASAP7_75t_L g1324 ( 
.A(n_1219),
.B(n_33),
.Y(n_1324)
);

INVx1_ASAP7_75t_L g1325 ( 
.A(n_1069),
.Y(n_1325)
);

INVx1_ASAP7_75t_SL g1326 ( 
.A(n_1175),
.Y(n_1326)
);

AND2x4_ASAP7_75t_L g1327 ( 
.A(n_1135),
.B(n_238),
.Y(n_1327)
);

INVx1_ASAP7_75t_L g1328 ( 
.A(n_1173),
.Y(n_1328)
);

CKINVDCx5p33_ASAP7_75t_R g1329 ( 
.A(n_1166),
.Y(n_1329)
);

INVx4_ASAP7_75t_L g1330 ( 
.A(n_1159),
.Y(n_1330)
);

INVx1_ASAP7_75t_L g1331 ( 
.A(n_1083),
.Y(n_1331)
);

INVx1_ASAP7_75t_L g1332 ( 
.A(n_1188),
.Y(n_1332)
);

AOI22xp5_ASAP7_75t_L g1333 ( 
.A1(n_1123),
.A2(n_241),
.B1(n_242),
.B2(n_240),
.Y(n_1333)
);

INVx2_ASAP7_75t_L g1334 ( 
.A(n_1092),
.Y(n_1334)
);

AOI221xp5_ASAP7_75t_SL g1335 ( 
.A1(n_1090),
.A2(n_37),
.B1(n_34),
.B2(n_36),
.C(n_38),
.Y(n_1335)
);

INVx2_ASAP7_75t_L g1336 ( 
.A(n_1095),
.Y(n_1336)
);

NAND2xp5_ASAP7_75t_SL g1337 ( 
.A(n_1159),
.B(n_245),
.Y(n_1337)
);

INVx1_ASAP7_75t_L g1338 ( 
.A(n_1087),
.Y(n_1338)
);

BUFx6f_ASAP7_75t_L g1339 ( 
.A(n_1218),
.Y(n_1339)
);

INVx2_ASAP7_75t_L g1340 ( 
.A(n_1218),
.Y(n_1340)
);

OR2x6_ASAP7_75t_L g1341 ( 
.A(n_1166),
.B(n_36),
.Y(n_1341)
);

NAND2xp5_ASAP7_75t_L g1342 ( 
.A(n_1221),
.B(n_37),
.Y(n_1342)
);

INVx2_ASAP7_75t_L g1343 ( 
.A(n_1218),
.Y(n_1343)
);

BUFx4f_ASAP7_75t_L g1344 ( 
.A(n_1096),
.Y(n_1344)
);

INVx1_ASAP7_75t_L g1345 ( 
.A(n_1088),
.Y(n_1345)
);

INVx1_ASAP7_75t_L g1346 ( 
.A(n_1091),
.Y(n_1346)
);

INVx1_ASAP7_75t_L g1347 ( 
.A(n_1086),
.Y(n_1347)
);

INVx4_ASAP7_75t_L g1348 ( 
.A(n_1096),
.Y(n_1348)
);

INVx2_ASAP7_75t_L g1349 ( 
.A(n_1168),
.Y(n_1349)
);

NAND2xp5_ASAP7_75t_SL g1350 ( 
.A(n_1149),
.B(n_247),
.Y(n_1350)
);

INVx1_ASAP7_75t_L g1351 ( 
.A(n_1116),
.Y(n_1351)
);

BUFx4f_ASAP7_75t_L g1352 ( 
.A(n_1205),
.Y(n_1352)
);

INVx1_ASAP7_75t_L g1353 ( 
.A(n_1118),
.Y(n_1353)
);

HB1xp67_ASAP7_75t_L g1354 ( 
.A(n_1164),
.Y(n_1354)
);

INVx2_ASAP7_75t_SL g1355 ( 
.A(n_1137),
.Y(n_1355)
);

NAND2xp5_ASAP7_75t_L g1356 ( 
.A(n_1128),
.B(n_38),
.Y(n_1356)
);

BUFx3_ASAP7_75t_L g1357 ( 
.A(n_1184),
.Y(n_1357)
);

AOI22xp33_ASAP7_75t_L g1358 ( 
.A1(n_1105),
.A2(n_41),
.B1(n_39),
.B2(n_40),
.Y(n_1358)
);

BUFx2_ASAP7_75t_L g1359 ( 
.A(n_1066),
.Y(n_1359)
);

NAND2xp5_ASAP7_75t_L g1360 ( 
.A(n_1104),
.B(n_39),
.Y(n_1360)
);

INVx1_ASAP7_75t_L g1361 ( 
.A(n_1122),
.Y(n_1361)
);

INVx5_ASAP7_75t_L g1362 ( 
.A(n_1206),
.Y(n_1362)
);

INVx1_ASAP7_75t_L g1363 ( 
.A(n_1062),
.Y(n_1363)
);

INVx1_ASAP7_75t_L g1364 ( 
.A(n_1220),
.Y(n_1364)
);

NAND2xp5_ASAP7_75t_L g1365 ( 
.A(n_1181),
.B(n_1080),
.Y(n_1365)
);

NAND2xp5_ASAP7_75t_L g1366 ( 
.A(n_1099),
.B(n_1103),
.Y(n_1366)
);

NAND2xp33_ASAP7_75t_SL g1367 ( 
.A(n_1142),
.B(n_41),
.Y(n_1367)
);

NAND2xp5_ASAP7_75t_L g1368 ( 
.A(n_1223),
.B(n_43),
.Y(n_1368)
);

CKINVDCx5p33_ASAP7_75t_R g1369 ( 
.A(n_1152),
.Y(n_1369)
);

INVx2_ASAP7_75t_L g1370 ( 
.A(n_1125),
.Y(n_1370)
);

NAND2xp5_ASAP7_75t_SL g1371 ( 
.A(n_1174),
.B(n_1187),
.Y(n_1371)
);

INVx2_ASAP7_75t_L g1372 ( 
.A(n_1144),
.Y(n_1372)
);

INVx2_ASAP7_75t_L g1373 ( 
.A(n_1106),
.Y(n_1373)
);

BUFx5_ASAP7_75t_L g1374 ( 
.A(n_1110),
.Y(n_1374)
);

HB1xp67_ASAP7_75t_L g1375 ( 
.A(n_1153),
.Y(n_1375)
);

INVx1_ASAP7_75t_L g1376 ( 
.A(n_1074),
.Y(n_1376)
);

AND2x4_ASAP7_75t_L g1377 ( 
.A(n_1093),
.B(n_1145),
.Y(n_1377)
);

CKINVDCx5p33_ASAP7_75t_R g1378 ( 
.A(n_1210),
.Y(n_1378)
);

NOR2xp33_ASAP7_75t_L g1379 ( 
.A(n_1121),
.B(n_43),
.Y(n_1379)
);

CKINVDCx11_ASAP7_75t_R g1380 ( 
.A(n_1090),
.Y(n_1380)
);

INVx2_ASAP7_75t_L g1381 ( 
.A(n_1141),
.Y(n_1381)
);

INVx2_ASAP7_75t_SL g1382 ( 
.A(n_1119),
.Y(n_1382)
);

INVx1_ASAP7_75t_L g1383 ( 
.A(n_1148),
.Y(n_1383)
);

NAND2xp5_ASAP7_75t_SL g1384 ( 
.A(n_1192),
.B(n_248),
.Y(n_1384)
);

INVxp67_ASAP7_75t_L g1385 ( 
.A(n_1126),
.Y(n_1385)
);

INVx2_ASAP7_75t_L g1386 ( 
.A(n_1078),
.Y(n_1386)
);

INVx1_ASAP7_75t_L g1387 ( 
.A(n_1151),
.Y(n_1387)
);

BUFx3_ASAP7_75t_L g1388 ( 
.A(n_1154),
.Y(n_1388)
);

INVx3_ASAP7_75t_L g1389 ( 
.A(n_1170),
.Y(n_1389)
);

INVx3_ASAP7_75t_L g1390 ( 
.A(n_1178),
.Y(n_1390)
);

INVx1_ASAP7_75t_L g1391 ( 
.A(n_1161),
.Y(n_1391)
);

INVx1_ASAP7_75t_L g1392 ( 
.A(n_1177),
.Y(n_1392)
);

INVx1_ASAP7_75t_L g1393 ( 
.A(n_1225),
.Y(n_1393)
);

NAND2xp5_ASAP7_75t_L g1394 ( 
.A(n_1147),
.B(n_1195),
.Y(n_1394)
);

INVx1_ASAP7_75t_L g1395 ( 
.A(n_1165),
.Y(n_1395)
);

INVx1_ASAP7_75t_L g1396 ( 
.A(n_1167),
.Y(n_1396)
);

AOI22xp33_ASAP7_75t_L g1397 ( 
.A1(n_1185),
.A2(n_48),
.B1(n_46),
.B2(n_47),
.Y(n_1397)
);

INVx3_ASAP7_75t_L g1398 ( 
.A(n_1203),
.Y(n_1398)
);

INVx2_ASAP7_75t_L g1399 ( 
.A(n_1085),
.Y(n_1399)
);

BUFx8_ASAP7_75t_L g1400 ( 
.A(n_1227),
.Y(n_1400)
);

NAND2xp5_ASAP7_75t_L g1401 ( 
.A(n_1129),
.B(n_47),
.Y(n_1401)
);

INVx2_ASAP7_75t_L g1402 ( 
.A(n_1226),
.Y(n_1402)
);

INVx1_ASAP7_75t_L g1403 ( 
.A(n_1196),
.Y(n_1403)
);

INVx2_ASAP7_75t_SL g1404 ( 
.A(n_1191),
.Y(n_1404)
);

AOI22xp5_ASAP7_75t_L g1405 ( 
.A1(n_1176),
.A2(n_251),
.B1(n_253),
.B2(n_250),
.Y(n_1405)
);

NOR2x1p5_ASAP7_75t_L g1406 ( 
.A(n_1204),
.B(n_254),
.Y(n_1406)
);

INVx2_ASAP7_75t_L g1407 ( 
.A(n_1226),
.Y(n_1407)
);

BUFx12f_ASAP7_75t_L g1408 ( 
.A(n_1171),
.Y(n_1408)
);

OAI22xp5_ASAP7_75t_SL g1409 ( 
.A1(n_1193),
.A2(n_51),
.B1(n_49),
.B2(n_50),
.Y(n_1409)
);

BUFx6f_ASAP7_75t_L g1410 ( 
.A(n_1202),
.Y(n_1410)
);

OR2x6_ASAP7_75t_L g1411 ( 
.A(n_1238),
.B(n_1134),
.Y(n_1411)
);

INVx2_ASAP7_75t_L g1412 ( 
.A(n_1230),
.Y(n_1412)
);

AND2x2_ASAP7_75t_L g1413 ( 
.A(n_1273),
.B(n_1197),
.Y(n_1413)
);

AND2x2_ASAP7_75t_L g1414 ( 
.A(n_1242),
.B(n_50),
.Y(n_1414)
);

INVx1_ASAP7_75t_L g1415 ( 
.A(n_1232),
.Y(n_1415)
);

NAND2xp5_ASAP7_75t_L g1416 ( 
.A(n_1287),
.B(n_1229),
.Y(n_1416)
);

AND2x4_ASAP7_75t_L g1417 ( 
.A(n_1348),
.B(n_255),
.Y(n_1417)
);

INVx1_ASAP7_75t_L g1418 ( 
.A(n_1232),
.Y(n_1418)
);

INVxp67_ASAP7_75t_L g1419 ( 
.A(n_1261),
.Y(n_1419)
);

NAND2xp5_ASAP7_75t_L g1420 ( 
.A(n_1351),
.B(n_52),
.Y(n_1420)
);

INVx2_ASAP7_75t_L g1421 ( 
.A(n_1280),
.Y(n_1421)
);

BUFx6f_ASAP7_75t_L g1422 ( 
.A(n_1245),
.Y(n_1422)
);

NAND2xp5_ASAP7_75t_SL g1423 ( 
.A(n_1357),
.B(n_53),
.Y(n_1423)
);

NAND2xp5_ASAP7_75t_L g1424 ( 
.A(n_1353),
.B(n_54),
.Y(n_1424)
);

INVx2_ASAP7_75t_L g1425 ( 
.A(n_1239),
.Y(n_1425)
);

INVx4_ASAP7_75t_L g1426 ( 
.A(n_1265),
.Y(n_1426)
);

INVx1_ASAP7_75t_L g1427 ( 
.A(n_1240),
.Y(n_1427)
);

AOI22xp5_ASAP7_75t_L g1428 ( 
.A1(n_1312),
.A2(n_57),
.B1(n_55),
.B2(n_56),
.Y(n_1428)
);

INVx6_ASAP7_75t_L g1429 ( 
.A(n_1292),
.Y(n_1429)
);

AND2x4_ASAP7_75t_L g1430 ( 
.A(n_1348),
.B(n_495),
.Y(n_1430)
);

INVx1_ASAP7_75t_SL g1431 ( 
.A(n_1254),
.Y(n_1431)
);

INVx1_ASAP7_75t_SL g1432 ( 
.A(n_1326),
.Y(n_1432)
);

NAND2xp5_ASAP7_75t_SL g1433 ( 
.A(n_1378),
.B(n_55),
.Y(n_1433)
);

AOI22xp5_ASAP7_75t_L g1434 ( 
.A1(n_1264),
.A2(n_58),
.B1(n_56),
.B2(n_57),
.Y(n_1434)
);

INVxp67_ASAP7_75t_SL g1435 ( 
.A(n_1392),
.Y(n_1435)
);

OAI22xp5_ASAP7_75t_L g1436 ( 
.A1(n_1284),
.A2(n_60),
.B1(n_58),
.B2(n_59),
.Y(n_1436)
);

NAND2xp5_ASAP7_75t_L g1437 ( 
.A(n_1376),
.B(n_59),
.Y(n_1437)
);

INVx1_ASAP7_75t_L g1438 ( 
.A(n_1243),
.Y(n_1438)
);

OR2x6_ASAP7_75t_L g1439 ( 
.A(n_1288),
.B(n_256),
.Y(n_1439)
);

AND2x2_ASAP7_75t_L g1440 ( 
.A(n_1246),
.B(n_61),
.Y(n_1440)
);

INVx1_ASAP7_75t_L g1441 ( 
.A(n_1247),
.Y(n_1441)
);

HB1xp67_ASAP7_75t_L g1442 ( 
.A(n_1300),
.Y(n_1442)
);

INVx3_ASAP7_75t_L g1443 ( 
.A(n_1330),
.Y(n_1443)
);

CKINVDCx5p33_ASAP7_75t_R g1444 ( 
.A(n_1274),
.Y(n_1444)
);

OAI22xp5_ASAP7_75t_L g1445 ( 
.A1(n_1366),
.A2(n_64),
.B1(n_62),
.B2(n_63),
.Y(n_1445)
);

INVx1_ASAP7_75t_SL g1446 ( 
.A(n_1231),
.Y(n_1446)
);

NAND2xp5_ASAP7_75t_L g1447 ( 
.A(n_1383),
.B(n_64),
.Y(n_1447)
);

BUFx12f_ASAP7_75t_L g1448 ( 
.A(n_1272),
.Y(n_1448)
);

INVx3_ASAP7_75t_L g1449 ( 
.A(n_1330),
.Y(n_1449)
);

BUFx2_ASAP7_75t_L g1450 ( 
.A(n_1318),
.Y(n_1450)
);

OAI22xp5_ASAP7_75t_L g1451 ( 
.A1(n_1344),
.A2(n_67),
.B1(n_65),
.B2(n_66),
.Y(n_1451)
);

INVx2_ASAP7_75t_L g1452 ( 
.A(n_1266),
.Y(n_1452)
);

AND2x4_ASAP7_75t_L g1453 ( 
.A(n_1260),
.B(n_494),
.Y(n_1453)
);

AND2x2_ASAP7_75t_L g1454 ( 
.A(n_1314),
.B(n_66),
.Y(n_1454)
);

INVxp33_ASAP7_75t_L g1455 ( 
.A(n_1263),
.Y(n_1455)
);

BUFx6f_ASAP7_75t_L g1456 ( 
.A(n_1245),
.Y(n_1456)
);

INVx1_ASAP7_75t_L g1457 ( 
.A(n_1251),
.Y(n_1457)
);

BUFx2_ASAP7_75t_L g1458 ( 
.A(n_1340),
.Y(n_1458)
);

HB1xp67_ASAP7_75t_L g1459 ( 
.A(n_1375),
.Y(n_1459)
);

INVx1_ASAP7_75t_L g1460 ( 
.A(n_1256),
.Y(n_1460)
);

AOI22xp33_ASAP7_75t_L g1461 ( 
.A1(n_1356),
.A2(n_70),
.B1(n_68),
.B2(n_69),
.Y(n_1461)
);

AND2x4_ASAP7_75t_L g1462 ( 
.A(n_1283),
.B(n_258),
.Y(n_1462)
);

NAND2xp5_ASAP7_75t_L g1463 ( 
.A(n_1387),
.B(n_71),
.Y(n_1463)
);

NAND2xp5_ASAP7_75t_L g1464 ( 
.A(n_1391),
.B(n_72),
.Y(n_1464)
);

NOR2xp33_ASAP7_75t_L g1465 ( 
.A(n_1369),
.B(n_72),
.Y(n_1465)
);

NAND2xp5_ASAP7_75t_L g1466 ( 
.A(n_1395),
.B(n_73),
.Y(n_1466)
);

AO22x1_ASAP7_75t_L g1467 ( 
.A1(n_1379),
.A2(n_75),
.B1(n_73),
.B2(n_74),
.Y(n_1467)
);

CKINVDCx5p33_ASAP7_75t_R g1468 ( 
.A(n_1276),
.Y(n_1468)
);

INVx3_ASAP7_75t_L g1469 ( 
.A(n_1245),
.Y(n_1469)
);

AND2x2_ASAP7_75t_L g1470 ( 
.A(n_1258),
.B(n_74),
.Y(n_1470)
);

INVx2_ASAP7_75t_L g1471 ( 
.A(n_1267),
.Y(n_1471)
);

AND2x2_ASAP7_75t_L g1472 ( 
.A(n_1344),
.B(n_75),
.Y(n_1472)
);

NAND2xp5_ASAP7_75t_L g1473 ( 
.A(n_1395),
.B(n_76),
.Y(n_1473)
);

INVx2_ASAP7_75t_L g1474 ( 
.A(n_1269),
.Y(n_1474)
);

INVx2_ASAP7_75t_L g1475 ( 
.A(n_1255),
.Y(n_1475)
);

AND2x2_ASAP7_75t_L g1476 ( 
.A(n_1396),
.B(n_76),
.Y(n_1476)
);

NAND2xp5_ASAP7_75t_L g1477 ( 
.A(n_1396),
.B(n_1331),
.Y(n_1477)
);

BUFx5_ASAP7_75t_L g1478 ( 
.A(n_1361),
.Y(n_1478)
);

BUFx6f_ASAP7_75t_L g1479 ( 
.A(n_1339),
.Y(n_1479)
);

INVx5_ASAP7_75t_L g1480 ( 
.A(n_1339),
.Y(n_1480)
);

AND2x2_ASAP7_75t_L g1481 ( 
.A(n_1241),
.B(n_77),
.Y(n_1481)
);

NAND2xp5_ASAP7_75t_L g1482 ( 
.A(n_1373),
.B(n_77),
.Y(n_1482)
);

HB1xp67_ASAP7_75t_L g1483 ( 
.A(n_1265),
.Y(n_1483)
);

INVx1_ASAP7_75t_L g1484 ( 
.A(n_1270),
.Y(n_1484)
);

CKINVDCx5p33_ASAP7_75t_R g1485 ( 
.A(n_1249),
.Y(n_1485)
);

INVx1_ASAP7_75t_SL g1486 ( 
.A(n_1277),
.Y(n_1486)
);

INVx4_ASAP7_75t_L g1487 ( 
.A(n_1265),
.Y(n_1487)
);

NAND2xp5_ASAP7_75t_L g1488 ( 
.A(n_1347),
.B(n_78),
.Y(n_1488)
);

INVxp67_ASAP7_75t_SL g1489 ( 
.A(n_1392),
.Y(n_1489)
);

INVx1_ASAP7_75t_L g1490 ( 
.A(n_1279),
.Y(n_1490)
);

INVx2_ASAP7_75t_L g1491 ( 
.A(n_1282),
.Y(n_1491)
);

BUFx4f_ASAP7_75t_L g1492 ( 
.A(n_1339),
.Y(n_1492)
);

INVx1_ASAP7_75t_L g1493 ( 
.A(n_1301),
.Y(n_1493)
);

NOR2xp33_ASAP7_75t_L g1494 ( 
.A(n_1388),
.B(n_78),
.Y(n_1494)
);

A2O1A1Ixp33_ASAP7_75t_L g1495 ( 
.A1(n_1237),
.A2(n_81),
.B(n_79),
.C(n_80),
.Y(n_1495)
);

INVx1_ASAP7_75t_L g1496 ( 
.A(n_1302),
.Y(n_1496)
);

AND2x2_ASAP7_75t_L g1497 ( 
.A(n_1293),
.B(n_1295),
.Y(n_1497)
);

NAND2xp5_ASAP7_75t_SL g1498 ( 
.A(n_1385),
.B(n_80),
.Y(n_1498)
);

BUFx6f_ASAP7_75t_L g1499 ( 
.A(n_1236),
.Y(n_1499)
);

INVx4_ASAP7_75t_L g1500 ( 
.A(n_1236),
.Y(n_1500)
);

INVx2_ASAP7_75t_SL g1501 ( 
.A(n_1292),
.Y(n_1501)
);

INVx1_ASAP7_75t_L g1502 ( 
.A(n_1311),
.Y(n_1502)
);

INVx1_ASAP7_75t_L g1503 ( 
.A(n_1309),
.Y(n_1503)
);

INVx1_ASAP7_75t_L g1504 ( 
.A(n_1332),
.Y(n_1504)
);

NAND2xp5_ASAP7_75t_SL g1505 ( 
.A(n_1377),
.B(n_83),
.Y(n_1505)
);

INVx2_ASAP7_75t_L g1506 ( 
.A(n_1308),
.Y(n_1506)
);

INVx2_ASAP7_75t_L g1507 ( 
.A(n_1328),
.Y(n_1507)
);

CKINVDCx5p33_ASAP7_75t_R g1508 ( 
.A(n_1359),
.Y(n_1508)
);

A2O1A1Ixp33_ASAP7_75t_L g1509 ( 
.A1(n_1305),
.A2(n_87),
.B(n_83),
.C(n_85),
.Y(n_1509)
);

INVx2_ASAP7_75t_L g1510 ( 
.A(n_1334),
.Y(n_1510)
);

INVx4_ASAP7_75t_L g1511 ( 
.A(n_1289),
.Y(n_1511)
);

CKINVDCx5p33_ASAP7_75t_R g1512 ( 
.A(n_1329),
.Y(n_1512)
);

BUFx6f_ASAP7_75t_L g1513 ( 
.A(n_1289),
.Y(n_1513)
);

INVx1_ASAP7_75t_L g1514 ( 
.A(n_1349),
.Y(n_1514)
);

BUFx6f_ASAP7_75t_L g1515 ( 
.A(n_1304),
.Y(n_1515)
);

INVx1_ASAP7_75t_L g1516 ( 
.A(n_1285),
.Y(n_1516)
);

INVx1_ASAP7_75t_L g1517 ( 
.A(n_1336),
.Y(n_1517)
);

AOI22xp5_ASAP7_75t_L g1518 ( 
.A1(n_1377),
.A2(n_1382),
.B1(n_1367),
.B2(n_1404),
.Y(n_1518)
);

NAND2xp5_ASAP7_75t_L g1519 ( 
.A(n_1317),
.B(n_85),
.Y(n_1519)
);

NAND2xp5_ASAP7_75t_L g1520 ( 
.A(n_1315),
.B(n_87),
.Y(n_1520)
);

NAND2xp5_ASAP7_75t_L g1521 ( 
.A(n_1319),
.B(n_88),
.Y(n_1521)
);

BUFx2_ASAP7_75t_L g1522 ( 
.A(n_1343),
.Y(n_1522)
);

AND2x2_ASAP7_75t_L g1523 ( 
.A(n_1283),
.B(n_89),
.Y(n_1523)
);

NAND2x1p5_ASAP7_75t_L g1524 ( 
.A(n_1304),
.B(n_259),
.Y(n_1524)
);

BUFx3_ASAP7_75t_L g1525 ( 
.A(n_1355),
.Y(n_1525)
);

INVx2_ASAP7_75t_L g1526 ( 
.A(n_1313),
.Y(n_1526)
);

INVx2_ASAP7_75t_L g1527 ( 
.A(n_1322),
.Y(n_1527)
);

INVx1_ASAP7_75t_L g1528 ( 
.A(n_1360),
.Y(n_1528)
);

NOR2xp33_ASAP7_75t_L g1529 ( 
.A(n_1298),
.B(n_89),
.Y(n_1529)
);

INVx1_ASAP7_75t_L g1530 ( 
.A(n_1363),
.Y(n_1530)
);

INVx2_ASAP7_75t_L g1531 ( 
.A(n_1338),
.Y(n_1531)
);

INVx2_ASAP7_75t_L g1532 ( 
.A(n_1345),
.Y(n_1532)
);

NOR2x1_ASAP7_75t_L g1533 ( 
.A(n_1398),
.B(n_1323),
.Y(n_1533)
);

INVx2_ASAP7_75t_L g1534 ( 
.A(n_1346),
.Y(n_1534)
);

AOI22xp33_ASAP7_75t_L g1535 ( 
.A1(n_1409),
.A2(n_92),
.B1(n_90),
.B2(n_91),
.Y(n_1535)
);

NAND2xp5_ASAP7_75t_L g1536 ( 
.A(n_1325),
.B(n_91),
.Y(n_1536)
);

NOR2xp33_ASAP7_75t_L g1537 ( 
.A(n_1321),
.B(n_94),
.Y(n_1537)
);

INVx2_ASAP7_75t_L g1538 ( 
.A(n_1399),
.Y(n_1538)
);

INVx1_ASAP7_75t_L g1539 ( 
.A(n_1281),
.Y(n_1539)
);

NOR2xp67_ASAP7_75t_L g1540 ( 
.A(n_1408),
.B(n_260),
.Y(n_1540)
);

NAND2xp5_ASAP7_75t_L g1541 ( 
.A(n_1257),
.B(n_95),
.Y(n_1541)
);

NAND2xp5_ASAP7_75t_L g1542 ( 
.A(n_1252),
.B(n_95),
.Y(n_1542)
);

AND2x4_ASAP7_75t_L g1543 ( 
.A(n_1327),
.B(n_263),
.Y(n_1543)
);

AND2x2_ASAP7_75t_SL g1544 ( 
.A(n_1286),
.B(n_96),
.Y(n_1544)
);

BUFx8_ASAP7_75t_L g1545 ( 
.A(n_1327),
.Y(n_1545)
);

NAND2xp5_ASAP7_75t_L g1546 ( 
.A(n_1365),
.B(n_96),
.Y(n_1546)
);

NAND2xp5_ASAP7_75t_L g1547 ( 
.A(n_1370),
.B(n_97),
.Y(n_1547)
);

NOR2xp33_ASAP7_75t_L g1548 ( 
.A(n_1380),
.B(n_99),
.Y(n_1548)
);

HB1xp67_ASAP7_75t_L g1549 ( 
.A(n_1235),
.Y(n_1549)
);

NAND2xp5_ASAP7_75t_L g1550 ( 
.A(n_1389),
.B(n_100),
.Y(n_1550)
);

INVx2_ASAP7_75t_L g1551 ( 
.A(n_1364),
.Y(n_1551)
);

AND3x1_ASAP7_75t_SL g1552 ( 
.A(n_1262),
.B(n_1290),
.C(n_1406),
.Y(n_1552)
);

BUFx6f_ASAP7_75t_L g1553 ( 
.A(n_1352),
.Y(n_1553)
);

NOR3xp33_ASAP7_75t_L g1554 ( 
.A(n_1371),
.B(n_103),
.C(n_104),
.Y(n_1554)
);

INVx2_ASAP7_75t_L g1555 ( 
.A(n_1372),
.Y(n_1555)
);

AND2x2_ASAP7_75t_L g1556 ( 
.A(n_1235),
.B(n_103),
.Y(n_1556)
);

INVx2_ASAP7_75t_L g1557 ( 
.A(n_1362),
.Y(n_1557)
);

AND2x2_ASAP7_75t_L g1558 ( 
.A(n_1248),
.B(n_104),
.Y(n_1558)
);

INVx1_ASAP7_75t_L g1559 ( 
.A(n_1268),
.Y(n_1559)
);

INVx2_ASAP7_75t_L g1560 ( 
.A(n_1362),
.Y(n_1560)
);

BUFx6f_ASAP7_75t_L g1561 ( 
.A(n_1352),
.Y(n_1561)
);

INVx4_ASAP7_75t_L g1562 ( 
.A(n_1362),
.Y(n_1562)
);

INVx2_ASAP7_75t_L g1563 ( 
.A(n_1386),
.Y(n_1563)
);

BUFx6f_ASAP7_75t_L g1564 ( 
.A(n_1341),
.Y(n_1564)
);

INVx1_ASAP7_75t_L g1565 ( 
.A(n_1294),
.Y(n_1565)
);

AND2x4_ASAP7_75t_L g1566 ( 
.A(n_1250),
.B(n_493),
.Y(n_1566)
);

AO22x1_ASAP7_75t_L g1567 ( 
.A1(n_1400),
.A2(n_107),
.B1(n_105),
.B2(n_106),
.Y(n_1567)
);

INVx1_ASAP7_75t_L g1568 ( 
.A(n_1306),
.Y(n_1568)
);

INVxp67_ASAP7_75t_L g1569 ( 
.A(n_1341),
.Y(n_1569)
);

NAND2xp5_ASAP7_75t_L g1570 ( 
.A(n_1389),
.B(n_107),
.Y(n_1570)
);

NAND2xp5_ASAP7_75t_SL g1571 ( 
.A(n_1259),
.B(n_108),
.Y(n_1571)
);

NOR2x2_ASAP7_75t_L g1572 ( 
.A(n_1402),
.B(n_109),
.Y(n_1572)
);

HB1xp67_ASAP7_75t_L g1573 ( 
.A(n_1354),
.Y(n_1573)
);

INVx4_ASAP7_75t_L g1574 ( 
.A(n_1398),
.Y(n_1574)
);

INVx1_ASAP7_75t_L g1575 ( 
.A(n_1324),
.Y(n_1575)
);

INVx5_ASAP7_75t_L g1576 ( 
.A(n_1410),
.Y(n_1576)
);

NAND2xp5_ASAP7_75t_L g1577 ( 
.A(n_1390),
.B(n_110),
.Y(n_1577)
);

INVx1_ASAP7_75t_L g1578 ( 
.A(n_1342),
.Y(n_1578)
);

NAND2xp33_ASAP7_75t_SL g1579 ( 
.A(n_1271),
.B(n_111),
.Y(n_1579)
);

BUFx6f_ASAP7_75t_L g1580 ( 
.A(n_1410),
.Y(n_1580)
);

AND2x2_ASAP7_75t_L g1581 ( 
.A(n_1320),
.B(n_112),
.Y(n_1581)
);

NAND2xp5_ASAP7_75t_L g1582 ( 
.A(n_1394),
.B(n_113),
.Y(n_1582)
);

BUFx2_ASAP7_75t_L g1583 ( 
.A(n_1400),
.Y(n_1583)
);

BUFx2_ASAP7_75t_L g1584 ( 
.A(n_1431),
.Y(n_1584)
);

INVx1_ASAP7_75t_L g1585 ( 
.A(n_1415),
.Y(n_1585)
);

OAI21x1_ASAP7_75t_L g1586 ( 
.A1(n_1555),
.A2(n_1381),
.B(n_1297),
.Y(n_1586)
);

CKINVDCx20_ASAP7_75t_R g1587 ( 
.A(n_1468),
.Y(n_1587)
);

OAI21x1_ASAP7_75t_L g1588 ( 
.A1(n_1563),
.A2(n_1407),
.B(n_1384),
.Y(n_1588)
);

O2A1O1Ixp5_ASAP7_75t_L g1589 ( 
.A1(n_1537),
.A2(n_1350),
.B(n_1368),
.C(n_1291),
.Y(n_1589)
);

INVx1_ASAP7_75t_L g1590 ( 
.A(n_1418),
.Y(n_1590)
);

AO31x2_ASAP7_75t_L g1591 ( 
.A1(n_1436),
.A2(n_1296),
.A3(n_1253),
.B(n_1393),
.Y(n_1591)
);

OAI22xp5_ASAP7_75t_L g1592 ( 
.A1(n_1518),
.A2(n_1397),
.B1(n_1234),
.B2(n_1244),
.Y(n_1592)
);

AO221x2_ASAP7_75t_L g1593 ( 
.A1(n_1467),
.A2(n_1335),
.B1(n_1401),
.B2(n_1278),
.C(n_1316),
.Y(n_1593)
);

AOI21xp33_ASAP7_75t_L g1594 ( 
.A1(n_1455),
.A2(n_1358),
.B(n_1403),
.Y(n_1594)
);

NAND2xp5_ASAP7_75t_L g1595 ( 
.A(n_1559),
.B(n_1477),
.Y(n_1595)
);

OAI21x1_ASAP7_75t_L g1596 ( 
.A1(n_1412),
.A2(n_1403),
.B(n_1307),
.Y(n_1596)
);

OAI21xp5_ASAP7_75t_L g1597 ( 
.A1(n_1533),
.A2(n_1405),
.B(n_1333),
.Y(n_1597)
);

AO31x2_ASAP7_75t_L g1598 ( 
.A1(n_1528),
.A2(n_1374),
.A3(n_1299),
.B(n_1310),
.Y(n_1598)
);

OAI22xp5_ASAP7_75t_L g1599 ( 
.A1(n_1549),
.A2(n_1410),
.B1(n_1233),
.B2(n_1337),
.Y(n_1599)
);

NAND2xp5_ASAP7_75t_SL g1600 ( 
.A(n_1497),
.B(n_1303),
.Y(n_1600)
);

OAI21xp5_ASAP7_75t_L g1601 ( 
.A1(n_1582),
.A2(n_1275),
.B(n_1374),
.Y(n_1601)
);

INVx1_ASAP7_75t_L g1602 ( 
.A(n_1421),
.Y(n_1602)
);

NAND2xp5_ASAP7_75t_L g1603 ( 
.A(n_1565),
.B(n_1374),
.Y(n_1603)
);

BUFx6f_ASAP7_75t_L g1604 ( 
.A(n_1492),
.Y(n_1604)
);

BUFx6f_ASAP7_75t_L g1605 ( 
.A(n_1480),
.Y(n_1605)
);

OAI21xp5_ASAP7_75t_L g1606 ( 
.A1(n_1568),
.A2(n_1374),
.B(n_114),
.Y(n_1606)
);

INVx1_ASAP7_75t_L g1607 ( 
.A(n_1427),
.Y(n_1607)
);

INVx1_ASAP7_75t_L g1608 ( 
.A(n_1438),
.Y(n_1608)
);

NAND2xp5_ASAP7_75t_L g1609 ( 
.A(n_1575),
.B(n_115),
.Y(n_1609)
);

OAI21x1_ASAP7_75t_L g1610 ( 
.A1(n_1530),
.A2(n_267),
.B(n_266),
.Y(n_1610)
);

A2O1A1Ixp33_ASAP7_75t_L g1611 ( 
.A1(n_1578),
.A2(n_118),
.B(n_116),
.C(n_117),
.Y(n_1611)
);

NAND2xp5_ASAP7_75t_L g1612 ( 
.A(n_1516),
.B(n_120),
.Y(n_1612)
);

NAND2xp5_ASAP7_75t_L g1613 ( 
.A(n_1539),
.B(n_121),
.Y(n_1613)
);

NAND2xp5_ASAP7_75t_SL g1614 ( 
.A(n_1574),
.B(n_121),
.Y(n_1614)
);

AOI21xp5_ASAP7_75t_L g1615 ( 
.A1(n_1435),
.A2(n_271),
.B(n_270),
.Y(n_1615)
);

OAI21x1_ASAP7_75t_L g1616 ( 
.A1(n_1551),
.A2(n_273),
.B(n_272),
.Y(n_1616)
);

OAI21x1_ASAP7_75t_L g1617 ( 
.A1(n_1531),
.A2(n_276),
.B(n_275),
.Y(n_1617)
);

NAND2xp5_ASAP7_75t_SL g1618 ( 
.A(n_1574),
.B(n_122),
.Y(n_1618)
);

INVx4_ASAP7_75t_L g1619 ( 
.A(n_1480),
.Y(n_1619)
);

OAI21x1_ASAP7_75t_L g1620 ( 
.A1(n_1532),
.A2(n_278),
.B(n_277),
.Y(n_1620)
);

INVx5_ASAP7_75t_L g1621 ( 
.A(n_1426),
.Y(n_1621)
);

NAND2xp5_ASAP7_75t_L g1622 ( 
.A(n_1534),
.B(n_122),
.Y(n_1622)
);

AOI21xp33_ASAP7_75t_L g1623 ( 
.A1(n_1544),
.A2(n_123),
.B(n_124),
.Y(n_1623)
);

NAND2xp5_ASAP7_75t_SL g1624 ( 
.A(n_1447),
.B(n_123),
.Y(n_1624)
);

OAI21x1_ASAP7_75t_L g1625 ( 
.A1(n_1416),
.A2(n_1490),
.B(n_1484),
.Y(n_1625)
);

AO21x1_ASAP7_75t_L g1626 ( 
.A1(n_1541),
.A2(n_125),
.B(n_126),
.Y(n_1626)
);

INVx2_ASAP7_75t_L g1627 ( 
.A(n_1491),
.Y(n_1627)
);

OAI21x1_ASAP7_75t_L g1628 ( 
.A1(n_1475),
.A2(n_281),
.B(n_279),
.Y(n_1628)
);

NAND3x1_ASAP7_75t_L g1629 ( 
.A(n_1465),
.B(n_125),
.C(n_126),
.Y(n_1629)
);

CKINVDCx5p33_ASAP7_75t_R g1630 ( 
.A(n_1444),
.Y(n_1630)
);

OAI22xp5_ASAP7_75t_L g1631 ( 
.A1(n_1432),
.A2(n_129),
.B1(n_127),
.B2(n_128),
.Y(n_1631)
);

NAND2xp5_ASAP7_75t_L g1632 ( 
.A(n_1510),
.B(n_127),
.Y(n_1632)
);

CKINVDCx20_ASAP7_75t_R g1633 ( 
.A(n_1485),
.Y(n_1633)
);

AOI21x1_ASAP7_75t_L g1634 ( 
.A1(n_1546),
.A2(n_283),
.B(n_282),
.Y(n_1634)
);

OAI21x1_ASAP7_75t_L g1635 ( 
.A1(n_1550),
.A2(n_286),
.B(n_284),
.Y(n_1635)
);

NAND2xp5_ASAP7_75t_L g1636 ( 
.A(n_1517),
.B(n_128),
.Y(n_1636)
);

NAND2xp5_ASAP7_75t_L g1637 ( 
.A(n_1514),
.B(n_129),
.Y(n_1637)
);

OAI21xp5_ASAP7_75t_L g1638 ( 
.A1(n_1519),
.A2(n_130),
.B(n_131),
.Y(n_1638)
);

HB1xp67_ASAP7_75t_L g1639 ( 
.A(n_1419),
.Y(n_1639)
);

INVx2_ASAP7_75t_L g1640 ( 
.A(n_1507),
.Y(n_1640)
);

NAND2xp5_ASAP7_75t_L g1641 ( 
.A(n_1581),
.B(n_130),
.Y(n_1641)
);

HB1xp67_ASAP7_75t_L g1642 ( 
.A(n_1442),
.Y(n_1642)
);

OAI21x1_ASAP7_75t_L g1643 ( 
.A1(n_1570),
.A2(n_290),
.B(n_287),
.Y(n_1643)
);

INVx5_ASAP7_75t_L g1644 ( 
.A(n_1426),
.Y(n_1644)
);

AOI21xp5_ASAP7_75t_SL g1645 ( 
.A1(n_1462),
.A2(n_297),
.B(n_296),
.Y(n_1645)
);

NAND2xp5_ASAP7_75t_L g1646 ( 
.A(n_1529),
.B(n_131),
.Y(n_1646)
);

OAI21x1_ASAP7_75t_L g1647 ( 
.A1(n_1577),
.A2(n_299),
.B(n_298),
.Y(n_1647)
);

AOI21x1_ASAP7_75t_L g1648 ( 
.A1(n_1542),
.A2(n_302),
.B(n_301),
.Y(n_1648)
);

INVxp67_ASAP7_75t_SL g1649 ( 
.A(n_1489),
.Y(n_1649)
);

AOI22x1_ASAP7_75t_L g1650 ( 
.A1(n_1557),
.A2(n_135),
.B1(n_132),
.B2(n_134),
.Y(n_1650)
);

OAI21x1_ASAP7_75t_L g1651 ( 
.A1(n_1538),
.A2(n_309),
.B(n_308),
.Y(n_1651)
);

OAI21xp5_ASAP7_75t_L g1652 ( 
.A1(n_1554),
.A2(n_132),
.B(n_134),
.Y(n_1652)
);

AND2x2_ASAP7_75t_L g1653 ( 
.A(n_1476),
.B(n_136),
.Y(n_1653)
);

NAND2x1p5_ASAP7_75t_L g1654 ( 
.A(n_1576),
.B(n_310),
.Y(n_1654)
);

HB1xp67_ASAP7_75t_L g1655 ( 
.A(n_1459),
.Y(n_1655)
);

OAI21xp5_ASAP7_75t_L g1656 ( 
.A1(n_1547),
.A2(n_138),
.B(n_139),
.Y(n_1656)
);

AOI21x1_ASAP7_75t_L g1657 ( 
.A1(n_1437),
.A2(n_1411),
.B(n_1488),
.Y(n_1657)
);

INVx1_ASAP7_75t_L g1658 ( 
.A(n_1441),
.Y(n_1658)
);

OR2x2_ASAP7_75t_L g1659 ( 
.A(n_1463),
.B(n_141),
.Y(n_1659)
);

OAI21x1_ASAP7_75t_L g1660 ( 
.A1(n_1504),
.A2(n_312),
.B(n_311),
.Y(n_1660)
);

NAND2xp5_ASAP7_75t_L g1661 ( 
.A(n_1464),
.B(n_142),
.Y(n_1661)
);

AOI21xp5_ASAP7_75t_L g1662 ( 
.A1(n_1576),
.A2(n_315),
.B(n_314),
.Y(n_1662)
);

AOI21xp5_ASAP7_75t_L g1663 ( 
.A1(n_1462),
.A2(n_1543),
.B(n_1411),
.Y(n_1663)
);

OAI21x1_ASAP7_75t_L g1664 ( 
.A1(n_1524),
.A2(n_317),
.B(n_316),
.Y(n_1664)
);

AOI21xp5_ASAP7_75t_L g1665 ( 
.A1(n_1543),
.A2(n_319),
.B(n_318),
.Y(n_1665)
);

INVxp67_ASAP7_75t_L g1666 ( 
.A(n_1573),
.Y(n_1666)
);

NAND2xp5_ASAP7_75t_L g1667 ( 
.A(n_1466),
.B(n_144),
.Y(n_1667)
);

INVx1_ASAP7_75t_L g1668 ( 
.A(n_1457),
.Y(n_1668)
);

INVxp67_ASAP7_75t_L g1669 ( 
.A(n_1450),
.Y(n_1669)
);

AOI21xp33_ASAP7_75t_L g1670 ( 
.A1(n_1413),
.A2(n_144),
.B(n_145),
.Y(n_1670)
);

OAI21xp5_ASAP7_75t_L g1671 ( 
.A1(n_1495),
.A2(n_145),
.B(n_146),
.Y(n_1671)
);

AND2x2_ASAP7_75t_L g1672 ( 
.A(n_1440),
.B(n_146),
.Y(n_1672)
);

NAND2xp5_ASAP7_75t_L g1673 ( 
.A(n_1473),
.B(n_147),
.Y(n_1673)
);

AO31x2_ASAP7_75t_L g1674 ( 
.A1(n_1509),
.A2(n_150),
.A3(n_148),
.B(n_149),
.Y(n_1674)
);

AOI21xp5_ASAP7_75t_L g1675 ( 
.A1(n_1417),
.A2(n_325),
.B(n_322),
.Y(n_1675)
);

AOI21xp5_ASAP7_75t_L g1676 ( 
.A1(n_1417),
.A2(n_328),
.B(n_326),
.Y(n_1676)
);

OAI22xp5_ASAP7_75t_L g1677 ( 
.A1(n_1535),
.A2(n_150),
.B1(n_148),
.B2(n_149),
.Y(n_1677)
);

NAND2xp5_ASAP7_75t_L g1678 ( 
.A(n_1420),
.B(n_151),
.Y(n_1678)
);

OAI21x1_ASAP7_75t_SL g1679 ( 
.A1(n_1520),
.A2(n_151),
.B(n_152),
.Y(n_1679)
);

AND2x4_ASAP7_75t_L g1680 ( 
.A(n_1553),
.B(n_329),
.Y(n_1680)
);

OAI21x1_ASAP7_75t_L g1681 ( 
.A1(n_1460),
.A2(n_334),
.B(n_332),
.Y(n_1681)
);

AND2x4_ASAP7_75t_L g1682 ( 
.A(n_1553),
.B(n_336),
.Y(n_1682)
);

NAND3xp33_ASAP7_75t_L g1683 ( 
.A(n_1434),
.B(n_152),
.C(n_153),
.Y(n_1683)
);

INVx1_ASAP7_75t_L g1684 ( 
.A(n_1493),
.Y(n_1684)
);

NAND2xp5_ASAP7_75t_L g1685 ( 
.A(n_1424),
.B(n_153),
.Y(n_1685)
);

INVx1_ASAP7_75t_L g1686 ( 
.A(n_1496),
.Y(n_1686)
);

INVx5_ASAP7_75t_L g1687 ( 
.A(n_1487),
.Y(n_1687)
);

A2O1A1Ixp33_ASAP7_75t_L g1688 ( 
.A1(n_1428),
.A2(n_154),
.B(n_155),
.C(n_156),
.Y(n_1688)
);

INVx4_ASAP7_75t_L g1689 ( 
.A(n_1480),
.Y(n_1689)
);

AOI21xp5_ASAP7_75t_L g1690 ( 
.A1(n_1430),
.A2(n_1580),
.B(n_1562),
.Y(n_1690)
);

OAI21x1_ASAP7_75t_L g1691 ( 
.A1(n_1502),
.A2(n_341),
.B(n_339),
.Y(n_1691)
);

NAND2xp5_ASAP7_75t_L g1692 ( 
.A(n_1521),
.B(n_154),
.Y(n_1692)
);

NAND2xp5_ASAP7_75t_L g1693 ( 
.A(n_1536),
.B(n_156),
.Y(n_1693)
);

NAND2xp5_ASAP7_75t_L g1694 ( 
.A(n_1482),
.B(n_157),
.Y(n_1694)
);

AND2x2_ASAP7_75t_L g1695 ( 
.A(n_1481),
.B(n_158),
.Y(n_1695)
);

INVx1_ASAP7_75t_L g1696 ( 
.A(n_1503),
.Y(n_1696)
);

NAND2xp5_ASAP7_75t_L g1697 ( 
.A(n_1505),
.B(n_160),
.Y(n_1697)
);

AO31x2_ASAP7_75t_L g1698 ( 
.A1(n_1445),
.A2(n_161),
.A3(n_163),
.B(n_164),
.Y(n_1698)
);

OAI21xp5_ASAP7_75t_L g1699 ( 
.A1(n_1571),
.A2(n_161),
.B(n_163),
.Y(n_1699)
);

NAND2xp5_ASAP7_75t_SL g1700 ( 
.A(n_1553),
.B(n_165),
.Y(n_1700)
);

NOR2xp33_ASAP7_75t_L g1701 ( 
.A(n_1446),
.B(n_342),
.Y(n_1701)
);

NAND2xp5_ASAP7_75t_SL g1702 ( 
.A(n_1561),
.B(n_165),
.Y(n_1702)
);

OAI22xp5_ASAP7_75t_L g1703 ( 
.A1(n_1569),
.A2(n_166),
.B1(n_167),
.B2(n_168),
.Y(n_1703)
);

AND2x2_ASAP7_75t_L g1704 ( 
.A(n_1470),
.B(n_168),
.Y(n_1704)
);

NAND2xp5_ASAP7_75t_L g1705 ( 
.A(n_1545),
.B(n_169),
.Y(n_1705)
);

AO21x1_ASAP7_75t_L g1706 ( 
.A1(n_1451),
.A2(n_1579),
.B(n_1498),
.Y(n_1706)
);

NOR2xp67_ASAP7_75t_L g1707 ( 
.A(n_1425),
.B(n_344),
.Y(n_1707)
);

AO21x1_ASAP7_75t_L g1708 ( 
.A1(n_1562),
.A2(n_170),
.B(n_171),
.Y(n_1708)
);

AO31x2_ASAP7_75t_L g1709 ( 
.A1(n_1478),
.A2(n_170),
.A3(n_171),
.B(n_172),
.Y(n_1709)
);

AO31x2_ASAP7_75t_L g1710 ( 
.A1(n_1478),
.A2(n_173),
.A3(n_174),
.B(n_175),
.Y(n_1710)
);

NAND2xp5_ASAP7_75t_L g1711 ( 
.A(n_1545),
.B(n_173),
.Y(n_1711)
);

AOI21xp5_ASAP7_75t_SL g1712 ( 
.A1(n_1566),
.A2(n_347),
.B(n_346),
.Y(n_1712)
);

OAI21x1_ASAP7_75t_L g1713 ( 
.A1(n_1526),
.A2(n_349),
.B(n_348),
.Y(n_1713)
);

INVx3_ASAP7_75t_L g1714 ( 
.A(n_1561),
.Y(n_1714)
);

OAI22xp5_ASAP7_75t_L g1715 ( 
.A1(n_1525),
.A2(n_174),
.B1(n_176),
.B2(n_177),
.Y(n_1715)
);

AOI211x1_ASAP7_75t_L g1716 ( 
.A1(n_1567),
.A2(n_1558),
.B(n_1433),
.C(n_1423),
.Y(n_1716)
);

A2O1A1Ixp33_ASAP7_75t_L g1717 ( 
.A1(n_1494),
.A2(n_176),
.B(n_177),
.C(n_178),
.Y(n_1717)
);

OAI21xp5_ASAP7_75t_L g1718 ( 
.A1(n_1461),
.A2(n_178),
.B(n_179),
.Y(n_1718)
);

NAND2xp5_ASAP7_75t_L g1719 ( 
.A(n_1523),
.B(n_179),
.Y(n_1719)
);

NAND2xp33_ASAP7_75t_L g1720 ( 
.A(n_1561),
.B(n_180),
.Y(n_1720)
);

INVx1_ASAP7_75t_SL g1721 ( 
.A(n_1486),
.Y(n_1721)
);

OAI21x1_ASAP7_75t_L g1722 ( 
.A1(n_1527),
.A2(n_351),
.B(n_350),
.Y(n_1722)
);

AND2x4_ASAP7_75t_L g1723 ( 
.A(n_1458),
.B(n_352),
.Y(n_1723)
);

HB1xp67_ASAP7_75t_L g1724 ( 
.A(n_1522),
.Y(n_1724)
);

AOI22xp5_ASAP7_75t_L g1725 ( 
.A1(n_1472),
.A2(n_180),
.B1(n_181),
.B2(n_182),
.Y(n_1725)
);

AND2x4_ASAP7_75t_L g1726 ( 
.A(n_1453),
.B(n_353),
.Y(n_1726)
);

NAND2xp5_ASAP7_75t_L g1727 ( 
.A(n_1556),
.B(n_182),
.Y(n_1727)
);

AND2x2_ASAP7_75t_L g1728 ( 
.A(n_1454),
.B(n_183),
.Y(n_1728)
);

BUFx3_ASAP7_75t_L g1729 ( 
.A(n_1448),
.Y(n_1729)
);

NOR2xp67_ASAP7_75t_SL g1730 ( 
.A(n_1712),
.B(n_1429),
.Y(n_1730)
);

AOI21xp5_ASAP7_75t_L g1731 ( 
.A1(n_1597),
.A2(n_1580),
.B(n_1478),
.Y(n_1731)
);

AND2x4_ASAP7_75t_L g1732 ( 
.A(n_1663),
.B(n_1453),
.Y(n_1732)
);

O2A1O1Ixp5_ASAP7_75t_L g1733 ( 
.A1(n_1652),
.A2(n_1548),
.B(n_1560),
.C(n_1500),
.Y(n_1733)
);

AND2x4_ASAP7_75t_L g1734 ( 
.A(n_1724),
.B(n_1469),
.Y(n_1734)
);

INVx1_ASAP7_75t_SL g1735 ( 
.A(n_1721),
.Y(n_1735)
);

INVx2_ASAP7_75t_L g1736 ( 
.A(n_1627),
.Y(n_1736)
);

AOI22xp5_ASAP7_75t_L g1737 ( 
.A1(n_1706),
.A2(n_1552),
.B1(n_1583),
.B2(n_1564),
.Y(n_1737)
);

BUFx6f_ASAP7_75t_L g1738 ( 
.A(n_1604),
.Y(n_1738)
);

OR2x2_ASAP7_75t_L g1739 ( 
.A(n_1655),
.B(n_1452),
.Y(n_1739)
);

AOI22xp33_ASAP7_75t_L g1740 ( 
.A1(n_1623),
.A2(n_1564),
.B1(n_1439),
.B2(n_1429),
.Y(n_1740)
);

AND2x4_ASAP7_75t_L g1741 ( 
.A(n_1714),
.B(n_1723),
.Y(n_1741)
);

AOI22xp5_ASAP7_75t_L g1742 ( 
.A1(n_1683),
.A2(n_1564),
.B1(n_1508),
.B2(n_1540),
.Y(n_1742)
);

INVx1_ASAP7_75t_L g1743 ( 
.A(n_1585),
.Y(n_1743)
);

BUFx3_ASAP7_75t_L g1744 ( 
.A(n_1584),
.Y(n_1744)
);

INVx1_ASAP7_75t_SL g1745 ( 
.A(n_1639),
.Y(n_1745)
);

CKINVDCx5p33_ASAP7_75t_R g1746 ( 
.A(n_1630),
.Y(n_1746)
);

BUFx10_ASAP7_75t_L g1747 ( 
.A(n_1604),
.Y(n_1747)
);

AOI21xp5_ASAP7_75t_L g1748 ( 
.A1(n_1595),
.A2(n_1449),
.B(n_1443),
.Y(n_1748)
);

NAND2x1p5_ASAP7_75t_L g1749 ( 
.A(n_1621),
.B(n_1443),
.Y(n_1749)
);

NOR2xp33_ASAP7_75t_L g1750 ( 
.A(n_1669),
.B(n_1512),
.Y(n_1750)
);

AOI21xp5_ASAP7_75t_L g1751 ( 
.A1(n_1649),
.A2(n_1449),
.B(n_1471),
.Y(n_1751)
);

INVx2_ASAP7_75t_L g1752 ( 
.A(n_1640),
.Y(n_1752)
);

AOI22xp5_ASAP7_75t_L g1753 ( 
.A1(n_1593),
.A2(n_1439),
.B1(n_1501),
.B2(n_1414),
.Y(n_1753)
);

BUFx6f_ASAP7_75t_L g1754 ( 
.A(n_1604),
.Y(n_1754)
);

AOI21x1_ASAP7_75t_L g1755 ( 
.A1(n_1657),
.A2(n_1483),
.B(n_1474),
.Y(n_1755)
);

INVx1_ASAP7_75t_L g1756 ( 
.A(n_1590),
.Y(n_1756)
);

NAND2xp5_ASAP7_75t_L g1757 ( 
.A(n_1642),
.B(n_1506),
.Y(n_1757)
);

AND2x4_ASAP7_75t_L g1758 ( 
.A(n_1690),
.B(n_1469),
.Y(n_1758)
);

INVx1_ASAP7_75t_SL g1759 ( 
.A(n_1587),
.Y(n_1759)
);

INVx2_ASAP7_75t_SL g1760 ( 
.A(n_1729),
.Y(n_1760)
);

INVx1_ASAP7_75t_L g1761 ( 
.A(n_1607),
.Y(n_1761)
);

INVx3_ASAP7_75t_SL g1762 ( 
.A(n_1633),
.Y(n_1762)
);

AND2x2_ASAP7_75t_L g1763 ( 
.A(n_1653),
.B(n_1499),
.Y(n_1763)
);

OR2x6_ASAP7_75t_L g1764 ( 
.A(n_1645),
.B(n_1500),
.Y(n_1764)
);

AOI21xp5_ASAP7_75t_L g1765 ( 
.A1(n_1606),
.A2(n_1511),
.B(n_1456),
.Y(n_1765)
);

INVx2_ASAP7_75t_SL g1766 ( 
.A(n_1605),
.Y(n_1766)
);

AOI21xp5_ASAP7_75t_L g1767 ( 
.A1(n_1603),
.A2(n_1511),
.B(n_1456),
.Y(n_1767)
);

OA21x2_ASAP7_75t_L g1768 ( 
.A1(n_1586),
.A2(n_1625),
.B(n_1588),
.Y(n_1768)
);

INVx3_ASAP7_75t_SL g1769 ( 
.A(n_1723),
.Y(n_1769)
);

BUFx6f_ASAP7_75t_L g1770 ( 
.A(n_1605),
.Y(n_1770)
);

NAND2xp5_ASAP7_75t_L g1771 ( 
.A(n_1667),
.B(n_1499),
.Y(n_1771)
);

AO21x2_ASAP7_75t_L g1772 ( 
.A1(n_1601),
.A2(n_1572),
.B(n_1456),
.Y(n_1772)
);

NAND3xp33_ASAP7_75t_L g1773 ( 
.A(n_1638),
.B(n_1513),
.C(n_1499),
.Y(n_1773)
);

INVx1_ASAP7_75t_L g1774 ( 
.A(n_1608),
.Y(n_1774)
);

INVx3_ASAP7_75t_L g1775 ( 
.A(n_1605),
.Y(n_1775)
);

AOI21xp5_ASAP7_75t_L g1776 ( 
.A1(n_1589),
.A2(n_1479),
.B(n_1422),
.Y(n_1776)
);

INVx1_ASAP7_75t_L g1777 ( 
.A(n_1658),
.Y(n_1777)
);

AND2x2_ASAP7_75t_L g1778 ( 
.A(n_1695),
.B(n_1513),
.Y(n_1778)
);

NAND2xp5_ASAP7_75t_L g1779 ( 
.A(n_1673),
.B(n_1716),
.Y(n_1779)
);

OAI22xp33_ASAP7_75t_L g1780 ( 
.A1(n_1725),
.A2(n_1515),
.B1(n_1513),
.B2(n_1479),
.Y(n_1780)
);

AOI21xp5_ASAP7_75t_L g1781 ( 
.A1(n_1671),
.A2(n_1479),
.B(n_1422),
.Y(n_1781)
);

NAND2x1p5_ASAP7_75t_L g1782 ( 
.A(n_1621),
.B(n_1422),
.Y(n_1782)
);

A2O1A1Ixp33_ASAP7_75t_L g1783 ( 
.A1(n_1718),
.A2(n_1515),
.B(n_184),
.C(n_185),
.Y(n_1783)
);

OAI22xp5_ASAP7_75t_L g1784 ( 
.A1(n_1629),
.A2(n_183),
.B1(n_184),
.B2(n_185),
.Y(n_1784)
);

AND2x4_ASAP7_75t_L g1785 ( 
.A(n_1668),
.B(n_354),
.Y(n_1785)
);

NAND2xp5_ASAP7_75t_L g1786 ( 
.A(n_1602),
.B(n_186),
.Y(n_1786)
);

AOI21xp5_ASAP7_75t_L g1787 ( 
.A1(n_1615),
.A2(n_357),
.B(n_356),
.Y(n_1787)
);

INVx1_ASAP7_75t_SL g1788 ( 
.A(n_1672),
.Y(n_1788)
);

INVx1_ASAP7_75t_L g1789 ( 
.A(n_1684),
.Y(n_1789)
);

INVx1_ASAP7_75t_L g1790 ( 
.A(n_1686),
.Y(n_1790)
);

INVx2_ASAP7_75t_SL g1791 ( 
.A(n_1621),
.Y(n_1791)
);

AOI21xp5_ASAP7_75t_L g1792 ( 
.A1(n_1593),
.A2(n_363),
.B(n_360),
.Y(n_1792)
);

AND2x2_ASAP7_75t_L g1793 ( 
.A(n_1704),
.B(n_364),
.Y(n_1793)
);

INVx1_ASAP7_75t_L g1794 ( 
.A(n_1696),
.Y(n_1794)
);

BUFx4_ASAP7_75t_SL g1795 ( 
.A(n_1659),
.Y(n_1795)
);

NAND2xp5_ASAP7_75t_L g1796 ( 
.A(n_1666),
.B(n_186),
.Y(n_1796)
);

AO21x1_ASAP7_75t_L g1797 ( 
.A1(n_1656),
.A2(n_1670),
.B(n_1592),
.Y(n_1797)
);

OAI21xp5_ASAP7_75t_L g1798 ( 
.A1(n_1688),
.A2(n_187),
.B(n_188),
.Y(n_1798)
);

AOI22xp33_ASAP7_75t_L g1799 ( 
.A1(n_1677),
.A2(n_187),
.B1(n_188),
.B2(n_189),
.Y(n_1799)
);

AOI21xp5_ASAP7_75t_L g1800 ( 
.A1(n_1600),
.A2(n_367),
.B(n_365),
.Y(n_1800)
);

INVx1_ASAP7_75t_L g1801 ( 
.A(n_1709),
.Y(n_1801)
);

INVx2_ASAP7_75t_L g1802 ( 
.A(n_1632),
.Y(n_1802)
);

NAND2xp5_ASAP7_75t_SL g1803 ( 
.A(n_1707),
.B(n_368),
.Y(n_1803)
);

BUFx3_ASAP7_75t_L g1804 ( 
.A(n_1726),
.Y(n_1804)
);

AND2x4_ASAP7_75t_L g1805 ( 
.A(n_1726),
.B(n_370),
.Y(n_1805)
);

OAI22xp5_ASAP7_75t_L g1806 ( 
.A1(n_1646),
.A2(n_1697),
.B1(n_1661),
.B2(n_1685),
.Y(n_1806)
);

CKINVDCx16_ASAP7_75t_R g1807 ( 
.A(n_1728),
.Y(n_1807)
);

INVxp67_ASAP7_75t_SL g1808 ( 
.A(n_1596),
.Y(n_1808)
);

O2A1O1Ixp33_ASAP7_75t_L g1809 ( 
.A1(n_1717),
.A2(n_189),
.B(n_190),
.C(n_192),
.Y(n_1809)
);

BUFx8_ASAP7_75t_SL g1810 ( 
.A(n_1705),
.Y(n_1810)
);

OR2x6_ASAP7_75t_L g1811 ( 
.A(n_1654),
.B(n_1665),
.Y(n_1811)
);

NAND2xp5_ASAP7_75t_L g1812 ( 
.A(n_1678),
.B(n_192),
.Y(n_1812)
);

AOI21xp5_ASAP7_75t_L g1813 ( 
.A1(n_1675),
.A2(n_372),
.B(n_371),
.Y(n_1813)
);

INVx3_ASAP7_75t_L g1814 ( 
.A(n_1619),
.Y(n_1814)
);

AOI21xp5_ASAP7_75t_L g1815 ( 
.A1(n_1676),
.A2(n_443),
.B(n_490),
.Y(n_1815)
);

AND2x2_ASAP7_75t_L g1816 ( 
.A(n_1641),
.B(n_373),
.Y(n_1816)
);

OAI22xp5_ASAP7_75t_L g1817 ( 
.A1(n_1692),
.A2(n_193),
.B1(n_194),
.B2(n_195),
.Y(n_1817)
);

AND2x4_ASAP7_75t_L g1818 ( 
.A(n_1680),
.B(n_375),
.Y(n_1818)
);

INVx1_ASAP7_75t_L g1819 ( 
.A(n_1709),
.Y(n_1819)
);

BUFx6f_ASAP7_75t_L g1820 ( 
.A(n_1619),
.Y(n_1820)
);

NOR2xp33_ASAP7_75t_L g1821 ( 
.A(n_1719),
.B(n_376),
.Y(n_1821)
);

OAI22xp5_ASAP7_75t_L g1822 ( 
.A1(n_1693),
.A2(n_193),
.B1(n_194),
.B2(n_195),
.Y(n_1822)
);

HB1xp67_ASAP7_75t_L g1823 ( 
.A(n_1599),
.Y(n_1823)
);

INVx1_ASAP7_75t_L g1824 ( 
.A(n_1710),
.Y(n_1824)
);

NOR2xp33_ASAP7_75t_L g1825 ( 
.A(n_1727),
.B(n_377),
.Y(n_1825)
);

BUFx4_ASAP7_75t_SL g1826 ( 
.A(n_1720),
.Y(n_1826)
);

NAND2xp5_ASAP7_75t_SL g1827 ( 
.A(n_1699),
.B(n_378),
.Y(n_1827)
);

AND2x4_ASAP7_75t_L g1828 ( 
.A(n_1644),
.B(n_380),
.Y(n_1828)
);

INVx1_ASAP7_75t_L g1829 ( 
.A(n_1743),
.Y(n_1829)
);

INVx1_ASAP7_75t_L g1830 ( 
.A(n_1756),
.Y(n_1830)
);

AND2x2_ASAP7_75t_L g1831 ( 
.A(n_1763),
.B(n_1710),
.Y(n_1831)
);

NAND2xp5_ASAP7_75t_L g1832 ( 
.A(n_1761),
.B(n_1710),
.Y(n_1832)
);

NAND2xp5_ASAP7_75t_L g1833 ( 
.A(n_1774),
.B(n_1698),
.Y(n_1833)
);

A2O1A1Ixp33_ASAP7_75t_L g1834 ( 
.A1(n_1809),
.A2(n_1611),
.B(n_1624),
.C(n_1694),
.Y(n_1834)
);

NAND2xp5_ASAP7_75t_L g1835 ( 
.A(n_1777),
.B(n_1698),
.Y(n_1835)
);

INVx1_ASAP7_75t_L g1836 ( 
.A(n_1789),
.Y(n_1836)
);

CKINVDCx5p33_ASAP7_75t_R g1837 ( 
.A(n_1746),
.Y(n_1837)
);

A2O1A1Ixp33_ASAP7_75t_L g1838 ( 
.A1(n_1798),
.A2(n_1662),
.B(n_1701),
.C(n_1700),
.Y(n_1838)
);

AND2x2_ASAP7_75t_L g1839 ( 
.A(n_1778),
.B(n_1734),
.Y(n_1839)
);

NAND2xp5_ASAP7_75t_L g1840 ( 
.A(n_1790),
.B(n_1698),
.Y(n_1840)
);

NAND2xp5_ASAP7_75t_SL g1841 ( 
.A(n_1732),
.B(n_1626),
.Y(n_1841)
);

INVx1_ASAP7_75t_SL g1842 ( 
.A(n_1745),
.Y(n_1842)
);

BUFx3_ASAP7_75t_L g1843 ( 
.A(n_1738),
.Y(n_1843)
);

AND2x2_ASAP7_75t_L g1844 ( 
.A(n_1734),
.B(n_1674),
.Y(n_1844)
);

OA21x2_ASAP7_75t_L g1845 ( 
.A1(n_1801),
.A2(n_1643),
.B(n_1635),
.Y(n_1845)
);

NAND2xp5_ASAP7_75t_L g1846 ( 
.A(n_1794),
.B(n_1674),
.Y(n_1846)
);

INVx2_ASAP7_75t_L g1847 ( 
.A(n_1736),
.Y(n_1847)
);

O2A1O1Ixp33_ASAP7_75t_L g1848 ( 
.A1(n_1783),
.A2(n_1631),
.B(n_1703),
.C(n_1702),
.Y(n_1848)
);

OR2x2_ASAP7_75t_L g1849 ( 
.A(n_1739),
.B(n_1636),
.Y(n_1849)
);

INVx2_ASAP7_75t_L g1850 ( 
.A(n_1752),
.Y(n_1850)
);

NAND2xp5_ASAP7_75t_L g1851 ( 
.A(n_1823),
.B(n_1674),
.Y(n_1851)
);

OAI22xp5_ASAP7_75t_L g1852 ( 
.A1(n_1799),
.A2(n_1650),
.B1(n_1609),
.B2(n_1612),
.Y(n_1852)
);

BUFx2_ASAP7_75t_R g1853 ( 
.A(n_1762),
.Y(n_1853)
);

INVx2_ASAP7_75t_L g1854 ( 
.A(n_1757),
.Y(n_1854)
);

AND2x2_ASAP7_75t_L g1855 ( 
.A(n_1788),
.B(n_1613),
.Y(n_1855)
);

OR2x2_ASAP7_75t_L g1856 ( 
.A(n_1802),
.B(n_1637),
.Y(n_1856)
);

CKINVDCx5p33_ASAP7_75t_R g1857 ( 
.A(n_1810),
.Y(n_1857)
);

AOI21x1_ASAP7_75t_SL g1858 ( 
.A1(n_1779),
.A2(n_1711),
.B(n_1622),
.Y(n_1858)
);

A2O1A1Ixp33_ASAP7_75t_SL g1859 ( 
.A1(n_1730),
.A2(n_1715),
.B(n_1594),
.C(n_1708),
.Y(n_1859)
);

OAI211xp5_ASAP7_75t_L g1860 ( 
.A1(n_1784),
.A2(n_1614),
.B(n_1618),
.C(n_1648),
.Y(n_1860)
);

NAND2x1p5_ASAP7_75t_L g1861 ( 
.A(n_1755),
.B(n_1644),
.Y(n_1861)
);

BUFx3_ASAP7_75t_L g1862 ( 
.A(n_1738),
.Y(n_1862)
);

OA22x2_ASAP7_75t_L g1863 ( 
.A1(n_1742),
.A2(n_1679),
.B1(n_1680),
.B2(n_1682),
.Y(n_1863)
);

INVx1_ASAP7_75t_L g1864 ( 
.A(n_1819),
.Y(n_1864)
);

INVx1_ASAP7_75t_L g1865 ( 
.A(n_1824),
.Y(n_1865)
);

AOI21xp5_ASAP7_75t_SL g1866 ( 
.A1(n_1805),
.A2(n_1682),
.B(n_1689),
.Y(n_1866)
);

OR2x2_ASAP7_75t_L g1867 ( 
.A(n_1744),
.B(n_1598),
.Y(n_1867)
);

INVx2_ASAP7_75t_L g1868 ( 
.A(n_1786),
.Y(n_1868)
);

AND2x2_ASAP7_75t_L g1869 ( 
.A(n_1772),
.B(n_1598),
.Y(n_1869)
);

AND2x4_ASAP7_75t_L g1870 ( 
.A(n_1732),
.B(n_1644),
.Y(n_1870)
);

INVx1_ASAP7_75t_L g1871 ( 
.A(n_1808),
.Y(n_1871)
);

NAND2xp5_ASAP7_75t_L g1872 ( 
.A(n_1797),
.B(n_1591),
.Y(n_1872)
);

BUFx3_ASAP7_75t_L g1873 ( 
.A(n_1754),
.Y(n_1873)
);

CKINVDCx20_ASAP7_75t_R g1874 ( 
.A(n_1759),
.Y(n_1874)
);

AND2x4_ASAP7_75t_L g1875 ( 
.A(n_1758),
.B(n_1687),
.Y(n_1875)
);

A2O1A1Ixp33_ASAP7_75t_L g1876 ( 
.A1(n_1733),
.A2(n_1664),
.B(n_1681),
.C(n_1691),
.Y(n_1876)
);

A2O1A1Ixp33_ASAP7_75t_SL g1877 ( 
.A1(n_1821),
.A2(n_1634),
.B(n_1647),
.C(n_1610),
.Y(n_1877)
);

AND2x2_ASAP7_75t_L g1878 ( 
.A(n_1807),
.B(n_1660),
.Y(n_1878)
);

CKINVDCx5p33_ASAP7_75t_R g1879 ( 
.A(n_1754),
.Y(n_1879)
);

INVx2_ASAP7_75t_L g1880 ( 
.A(n_1864),
.Y(n_1880)
);

OAI221xp5_ASAP7_75t_L g1881 ( 
.A1(n_1838),
.A2(n_1740),
.B1(n_1806),
.B2(n_1792),
.C(n_1817),
.Y(n_1881)
);

HB1xp67_ASAP7_75t_L g1882 ( 
.A(n_1842),
.Y(n_1882)
);

INVx1_ASAP7_75t_L g1883 ( 
.A(n_1865),
.Y(n_1883)
);

INVx1_ASAP7_75t_L g1884 ( 
.A(n_1829),
.Y(n_1884)
);

NAND2xp5_ASAP7_75t_L g1885 ( 
.A(n_1854),
.B(n_1731),
.Y(n_1885)
);

INVx3_ASAP7_75t_L g1886 ( 
.A(n_1847),
.Y(n_1886)
);

CKINVDCx5p33_ASAP7_75t_R g1887 ( 
.A(n_1837),
.Y(n_1887)
);

INVx2_ASAP7_75t_L g1888 ( 
.A(n_1830),
.Y(n_1888)
);

AND2x4_ASAP7_75t_L g1889 ( 
.A(n_1844),
.B(n_1758),
.Y(n_1889)
);

AOI22xp33_ASAP7_75t_L g1890 ( 
.A1(n_1863),
.A2(n_1827),
.B1(n_1773),
.B2(n_1822),
.Y(n_1890)
);

INVx1_ASAP7_75t_L g1891 ( 
.A(n_1836),
.Y(n_1891)
);

NAND2x1p5_ASAP7_75t_L g1892 ( 
.A(n_1845),
.B(n_1768),
.Y(n_1892)
);

BUFx3_ASAP7_75t_L g1893 ( 
.A(n_1875),
.Y(n_1893)
);

BUFx2_ASAP7_75t_L g1894 ( 
.A(n_1867),
.Y(n_1894)
);

INVx1_ASAP7_75t_L g1895 ( 
.A(n_1846),
.Y(n_1895)
);

OR2x2_ASAP7_75t_L g1896 ( 
.A(n_1846),
.B(n_1735),
.Y(n_1896)
);

INVx1_ASAP7_75t_L g1897 ( 
.A(n_1832),
.Y(n_1897)
);

AO21x2_ASAP7_75t_L g1898 ( 
.A1(n_1872),
.A2(n_1776),
.B(n_1765),
.Y(n_1898)
);

INVx2_ASAP7_75t_L g1899 ( 
.A(n_1850),
.Y(n_1899)
);

AO21x2_ASAP7_75t_L g1900 ( 
.A1(n_1872),
.A2(n_1751),
.B(n_1781),
.Y(n_1900)
);

INVx2_ASAP7_75t_L g1901 ( 
.A(n_1832),
.Y(n_1901)
);

INVx2_ASAP7_75t_L g1902 ( 
.A(n_1871),
.Y(n_1902)
);

INVx8_ASAP7_75t_L g1903 ( 
.A(n_1870),
.Y(n_1903)
);

INVxp33_ASAP7_75t_L g1904 ( 
.A(n_1839),
.Y(n_1904)
);

HB1xp67_ASAP7_75t_L g1905 ( 
.A(n_1842),
.Y(n_1905)
);

INVx3_ASAP7_75t_L g1906 ( 
.A(n_1875),
.Y(n_1906)
);

BUFx2_ASAP7_75t_L g1907 ( 
.A(n_1869),
.Y(n_1907)
);

INVx2_ASAP7_75t_L g1908 ( 
.A(n_1833),
.Y(n_1908)
);

BUFx3_ASAP7_75t_L g1909 ( 
.A(n_1893),
.Y(n_1909)
);

INVx2_ASAP7_75t_L g1910 ( 
.A(n_1880),
.Y(n_1910)
);

INVx1_ASAP7_75t_SL g1911 ( 
.A(n_1894),
.Y(n_1911)
);

AND2x2_ASAP7_75t_L g1912 ( 
.A(n_1907),
.B(n_1831),
.Y(n_1912)
);

OAI222xp33_ASAP7_75t_L g1913 ( 
.A1(n_1881),
.A2(n_1841),
.B1(n_1863),
.B2(n_1878),
.C1(n_1753),
.C2(n_1852),
.Y(n_1913)
);

INVx1_ASAP7_75t_L g1914 ( 
.A(n_1880),
.Y(n_1914)
);

AND2x2_ASAP7_75t_L g1915 ( 
.A(n_1907),
.B(n_1851),
.Y(n_1915)
);

INVx2_ASAP7_75t_SL g1916 ( 
.A(n_1903),
.Y(n_1916)
);

AOI22xp33_ASAP7_75t_L g1917 ( 
.A1(n_1881),
.A2(n_1852),
.B1(n_1811),
.B2(n_1787),
.Y(n_1917)
);

BUFx3_ASAP7_75t_L g1918 ( 
.A(n_1893),
.Y(n_1918)
);

INVx2_ASAP7_75t_L g1919 ( 
.A(n_1880),
.Y(n_1919)
);

AND2x2_ASAP7_75t_L g1920 ( 
.A(n_1894),
.B(n_1851),
.Y(n_1920)
);

NAND2xp5_ASAP7_75t_L g1921 ( 
.A(n_1882),
.B(n_1868),
.Y(n_1921)
);

INVx2_ASAP7_75t_L g1922 ( 
.A(n_1908),
.Y(n_1922)
);

AND2x2_ASAP7_75t_L g1923 ( 
.A(n_1889),
.B(n_1833),
.Y(n_1923)
);

HB1xp67_ASAP7_75t_L g1924 ( 
.A(n_1905),
.Y(n_1924)
);

INVx1_ASAP7_75t_L g1925 ( 
.A(n_1883),
.Y(n_1925)
);

OR2x2_ASAP7_75t_L g1926 ( 
.A(n_1896),
.B(n_1835),
.Y(n_1926)
);

HB1xp67_ASAP7_75t_L g1927 ( 
.A(n_1908),
.Y(n_1927)
);

HB1xp67_ASAP7_75t_L g1928 ( 
.A(n_1908),
.Y(n_1928)
);

HB1xp67_ASAP7_75t_L g1929 ( 
.A(n_1901),
.Y(n_1929)
);

INVx2_ASAP7_75t_L g1930 ( 
.A(n_1910),
.Y(n_1930)
);

INVx2_ASAP7_75t_L g1931 ( 
.A(n_1910),
.Y(n_1931)
);

AND2x2_ASAP7_75t_L g1932 ( 
.A(n_1923),
.B(n_1906),
.Y(n_1932)
);

NAND2xp5_ASAP7_75t_L g1933 ( 
.A(n_1924),
.B(n_1896),
.Y(n_1933)
);

NAND2xp5_ASAP7_75t_L g1934 ( 
.A(n_1915),
.B(n_1897),
.Y(n_1934)
);

INVxp67_ASAP7_75t_SL g1935 ( 
.A(n_1927),
.Y(n_1935)
);

NAND2xp5_ASAP7_75t_L g1936 ( 
.A(n_1915),
.B(n_1897),
.Y(n_1936)
);

INVx3_ASAP7_75t_L g1937 ( 
.A(n_1909),
.Y(n_1937)
);

AND2x2_ASAP7_75t_L g1938 ( 
.A(n_1923),
.B(n_1906),
.Y(n_1938)
);

INVxp67_ASAP7_75t_R g1939 ( 
.A(n_1912),
.Y(n_1939)
);

INVx1_ASAP7_75t_L g1940 ( 
.A(n_1930),
.Y(n_1940)
);

AND2x2_ASAP7_75t_L g1941 ( 
.A(n_1939),
.B(n_1909),
.Y(n_1941)
);

INVx1_ASAP7_75t_L g1942 ( 
.A(n_1931),
.Y(n_1942)
);

INVx2_ASAP7_75t_L g1943 ( 
.A(n_1937),
.Y(n_1943)
);

OR2x6_ASAP7_75t_L g1944 ( 
.A(n_1937),
.B(n_1866),
.Y(n_1944)
);

NAND2xp5_ASAP7_75t_L g1945 ( 
.A(n_1933),
.B(n_1920),
.Y(n_1945)
);

AOI222xp33_ASAP7_75t_L g1946 ( 
.A1(n_1941),
.A2(n_1913),
.B1(n_1917),
.B2(n_1812),
.C1(n_1890),
.C2(n_1834),
.Y(n_1946)
);

INVxp67_ASAP7_75t_SL g1947 ( 
.A(n_1943),
.Y(n_1947)
);

HB1xp67_ASAP7_75t_L g1948 ( 
.A(n_1940),
.Y(n_1948)
);

INVx1_ASAP7_75t_L g1949 ( 
.A(n_1940),
.Y(n_1949)
);

INVx1_ASAP7_75t_L g1950 ( 
.A(n_1942),
.Y(n_1950)
);

OAI22xp5_ASAP7_75t_L g1951 ( 
.A1(n_1944),
.A2(n_1936),
.B1(n_1934),
.B2(n_1918),
.Y(n_1951)
);

INVxp67_ASAP7_75t_L g1952 ( 
.A(n_1944),
.Y(n_1952)
);

INVx1_ASAP7_75t_L g1953 ( 
.A(n_1945),
.Y(n_1953)
);

INVx2_ASAP7_75t_L g1954 ( 
.A(n_1940),
.Y(n_1954)
);

INVx1_ASAP7_75t_L g1955 ( 
.A(n_1940),
.Y(n_1955)
);

INVxp67_ASAP7_75t_SL g1956 ( 
.A(n_1948),
.Y(n_1956)
);

INVx2_ASAP7_75t_L g1957 ( 
.A(n_1954),
.Y(n_1957)
);

NAND2xp5_ASAP7_75t_L g1958 ( 
.A(n_1953),
.B(n_1934),
.Y(n_1958)
);

AOI21xp33_ASAP7_75t_L g1959 ( 
.A1(n_1946),
.A2(n_1859),
.B(n_1825),
.Y(n_1959)
);

INVx2_ASAP7_75t_SL g1960 ( 
.A(n_1948),
.Y(n_1960)
);

AND2x4_ASAP7_75t_L g1961 ( 
.A(n_1947),
.B(n_1909),
.Y(n_1961)
);

INVx2_ASAP7_75t_L g1962 ( 
.A(n_1954),
.Y(n_1962)
);

AND2x2_ASAP7_75t_L g1963 ( 
.A(n_1952),
.B(n_1932),
.Y(n_1963)
);

INVx1_ASAP7_75t_L g1964 ( 
.A(n_1949),
.Y(n_1964)
);

INVx1_ASAP7_75t_L g1965 ( 
.A(n_1955),
.Y(n_1965)
);

INVx1_ASAP7_75t_L g1966 ( 
.A(n_1950),
.Y(n_1966)
);

NOR2xp33_ASAP7_75t_L g1967 ( 
.A(n_1966),
.B(n_1857),
.Y(n_1967)
);

INVxp67_ASAP7_75t_SL g1968 ( 
.A(n_1956),
.Y(n_1968)
);

AND2x2_ASAP7_75t_L g1969 ( 
.A(n_1963),
.B(n_1951),
.Y(n_1969)
);

BUFx2_ASAP7_75t_SL g1970 ( 
.A(n_1960),
.Y(n_1970)
);

INVx1_ASAP7_75t_L g1971 ( 
.A(n_1956),
.Y(n_1971)
);

INVx1_ASAP7_75t_L g1972 ( 
.A(n_1957),
.Y(n_1972)
);

AND2x2_ASAP7_75t_L g1973 ( 
.A(n_1961),
.B(n_1938),
.Y(n_1973)
);

INVx1_ASAP7_75t_L g1974 ( 
.A(n_1962),
.Y(n_1974)
);

AND2x2_ASAP7_75t_L g1975 ( 
.A(n_1969),
.B(n_1961),
.Y(n_1975)
);

OR2x6_ASAP7_75t_L g1976 ( 
.A(n_1970),
.B(n_1760),
.Y(n_1976)
);

NAND2xp33_ASAP7_75t_SL g1977 ( 
.A(n_1971),
.B(n_1887),
.Y(n_1977)
);

OR2x2_ASAP7_75t_L g1978 ( 
.A(n_1968),
.B(n_1958),
.Y(n_1978)
);

NAND2xp5_ASAP7_75t_L g1979 ( 
.A(n_1975),
.B(n_1968),
.Y(n_1979)
);

INVx1_ASAP7_75t_L g1980 ( 
.A(n_1978),
.Y(n_1980)
);

AND2x2_ASAP7_75t_L g1981 ( 
.A(n_1976),
.B(n_1967),
.Y(n_1981)
);

INVx1_ASAP7_75t_L g1982 ( 
.A(n_1977),
.Y(n_1982)
);

NAND2x1p5_ASAP7_75t_L g1983 ( 
.A(n_1981),
.B(n_1967),
.Y(n_1983)
);

INVx2_ASAP7_75t_L g1984 ( 
.A(n_1979),
.Y(n_1984)
);

INVx1_ASAP7_75t_L g1985 ( 
.A(n_1980),
.Y(n_1985)
);

INVx1_ASAP7_75t_L g1986 ( 
.A(n_1982),
.Y(n_1986)
);

INVx1_ASAP7_75t_L g1987 ( 
.A(n_1979),
.Y(n_1987)
);

NOR2xp33_ASAP7_75t_L g1988 ( 
.A(n_1983),
.B(n_1972),
.Y(n_1988)
);

INVx1_ASAP7_75t_L g1989 ( 
.A(n_1985),
.Y(n_1989)
);

INVx1_ASAP7_75t_L g1990 ( 
.A(n_1985),
.Y(n_1990)
);

NOR2xp33_ASAP7_75t_L g1991 ( 
.A(n_1986),
.B(n_1974),
.Y(n_1991)
);

NAND2x1_ASAP7_75t_L g1992 ( 
.A(n_1984),
.B(n_1964),
.Y(n_1992)
);

AND2x2_ASAP7_75t_L g1993 ( 
.A(n_1987),
.B(n_1973),
.Y(n_1993)
);

NAND2xp5_ASAP7_75t_L g1994 ( 
.A(n_1986),
.B(n_1965),
.Y(n_1994)
);

INVx1_ASAP7_75t_L g1995 ( 
.A(n_1985),
.Y(n_1995)
);

NAND2xp5_ASAP7_75t_L g1996 ( 
.A(n_1986),
.B(n_1958),
.Y(n_1996)
);

INVx1_ASAP7_75t_L g1997 ( 
.A(n_1985),
.Y(n_1997)
);

XOR2x2_ASAP7_75t_L g1998 ( 
.A(n_1988),
.B(n_1750),
.Y(n_1998)
);

NAND2xp33_ASAP7_75t_SL g1999 ( 
.A(n_1992),
.B(n_1874),
.Y(n_1999)
);

INVx1_ASAP7_75t_L g2000 ( 
.A(n_1993),
.Y(n_2000)
);

AOI211xp5_ASAP7_75t_L g2001 ( 
.A1(n_1991),
.A2(n_1959),
.B(n_1796),
.C(n_1737),
.Y(n_2001)
);

INVx2_ASAP7_75t_L g2002 ( 
.A(n_1989),
.Y(n_2002)
);

INVxp33_ASAP7_75t_L g2003 ( 
.A(n_1996),
.Y(n_2003)
);

HB1xp67_ASAP7_75t_L g2004 ( 
.A(n_1990),
.Y(n_2004)
);

NAND2x1_ASAP7_75t_SL g2005 ( 
.A(n_1995),
.B(n_1689),
.Y(n_2005)
);

NAND2xp5_ASAP7_75t_L g2006 ( 
.A(n_1997),
.B(n_1959),
.Y(n_2006)
);

NAND2xp5_ASAP7_75t_L g2007 ( 
.A(n_1994),
.B(n_1935),
.Y(n_2007)
);

NAND2xp5_ASAP7_75t_L g2008 ( 
.A(n_1988),
.B(n_1936),
.Y(n_2008)
);

NAND2xp5_ASAP7_75t_L g2009 ( 
.A(n_1988),
.B(n_1911),
.Y(n_2009)
);

NAND2xp5_ASAP7_75t_L g2010 ( 
.A(n_1988),
.B(n_1911),
.Y(n_2010)
);

NAND3xp33_ASAP7_75t_L g2011 ( 
.A(n_2000),
.B(n_1879),
.C(n_1816),
.Y(n_2011)
);

AOI21xp5_ASAP7_75t_L g2012 ( 
.A1(n_1999),
.A2(n_1771),
.B(n_1848),
.Y(n_2012)
);

AOI211xp5_ASAP7_75t_L g2013 ( 
.A1(n_2003),
.A2(n_1828),
.B(n_1793),
.C(n_1805),
.Y(n_2013)
);

NOR3xp33_ASAP7_75t_L g2014 ( 
.A(n_2006),
.B(n_1853),
.C(n_1795),
.Y(n_2014)
);

NAND2xp5_ASAP7_75t_L g2015 ( 
.A(n_2004),
.B(n_1921),
.Y(n_2015)
);

AOI211xp5_ASAP7_75t_L g2016 ( 
.A1(n_2009),
.A2(n_1828),
.B(n_1818),
.C(n_1800),
.Y(n_2016)
);

AND2x2_ASAP7_75t_L g2017 ( 
.A(n_1998),
.B(n_1918),
.Y(n_2017)
);

OAI211xp5_ASAP7_75t_L g2018 ( 
.A1(n_2005),
.A2(n_1813),
.B(n_1815),
.C(n_1687),
.Y(n_2018)
);

AOI21xp5_ASAP7_75t_L g2019 ( 
.A1(n_2010),
.A2(n_1803),
.B(n_1877),
.Y(n_2019)
);

OAI211xp5_ASAP7_75t_SL g2020 ( 
.A1(n_2007),
.A2(n_1860),
.B(n_1849),
.C(n_1856),
.Y(n_2020)
);

NOR2xp33_ASAP7_75t_L g2021 ( 
.A(n_2008),
.B(n_1747),
.Y(n_2021)
);

NAND2xp5_ASAP7_75t_L g2022 ( 
.A(n_2002),
.B(n_1855),
.Y(n_2022)
);

NAND2xp5_ASAP7_75t_L g2023 ( 
.A(n_2001),
.B(n_1918),
.Y(n_2023)
);

NAND2xp5_ASAP7_75t_L g2024 ( 
.A(n_2017),
.B(n_1925),
.Y(n_2024)
);

NAND2xp5_ASAP7_75t_SL g2025 ( 
.A(n_2014),
.B(n_1820),
.Y(n_2025)
);

NAND3xp33_ASAP7_75t_L g2026 ( 
.A(n_2021),
.B(n_1687),
.C(n_1820),
.Y(n_2026)
);

NAND3xp33_ASAP7_75t_L g2027 ( 
.A(n_2011),
.B(n_1770),
.C(n_1843),
.Y(n_2027)
);

NAND3xp33_ASAP7_75t_SL g2028 ( 
.A(n_2018),
.B(n_1826),
.C(n_1782),
.Y(n_2028)
);

NAND2xp5_ASAP7_75t_SL g2029 ( 
.A(n_2015),
.B(n_1770),
.Y(n_2029)
);

NOR3xp33_ASAP7_75t_L g2030 ( 
.A(n_2023),
.B(n_1775),
.C(n_1766),
.Y(n_2030)
);

NOR5xp2_ASAP7_75t_L g2031 ( 
.A(n_2020),
.B(n_196),
.C(n_197),
.D(n_198),
.E(n_199),
.Y(n_2031)
);

AOI211xp5_ASAP7_75t_L g2032 ( 
.A1(n_2022),
.A2(n_1769),
.B(n_1780),
.C(n_198),
.Y(n_2032)
);

AOI211xp5_ASAP7_75t_L g2033 ( 
.A1(n_2019),
.A2(n_196),
.B(n_197),
.C(n_199),
.Y(n_2033)
);

NAND2xp5_ASAP7_75t_L g2034 ( 
.A(n_2013),
.B(n_1925),
.Y(n_2034)
);

NAND2xp5_ASAP7_75t_L g2035 ( 
.A(n_2012),
.B(n_1910),
.Y(n_2035)
);

INVxp67_ASAP7_75t_L g2036 ( 
.A(n_2025),
.Y(n_2036)
);

NAND3xp33_ASAP7_75t_L g2037 ( 
.A(n_2033),
.B(n_2016),
.C(n_201),
.Y(n_2037)
);

NAND2xp5_ASAP7_75t_L g2038 ( 
.A(n_2030),
.B(n_201),
.Y(n_2038)
);

INVx1_ASAP7_75t_L g2039 ( 
.A(n_2024),
.Y(n_2039)
);

NOR2x1_ASAP7_75t_L g2040 ( 
.A(n_2028),
.B(n_202),
.Y(n_2040)
);

OAI21xp33_ASAP7_75t_L g2041 ( 
.A1(n_2034),
.A2(n_1873),
.B(n_1862),
.Y(n_2041)
);

AOI321xp33_ASAP7_75t_L g2042 ( 
.A1(n_2029),
.A2(n_1785),
.A3(n_1741),
.B1(n_1885),
.B2(n_205),
.C(n_206),
.Y(n_2042)
);

AND2x4_ASAP7_75t_L g2043 ( 
.A(n_2027),
.B(n_2026),
.Y(n_2043)
);

AOI221xp5_ASAP7_75t_L g2044 ( 
.A1(n_2032),
.A2(n_1785),
.B1(n_203),
.B2(n_204),
.C(n_205),
.Y(n_2044)
);

OAI21xp33_ASAP7_75t_L g2045 ( 
.A1(n_2035),
.A2(n_2031),
.B(n_1920),
.Y(n_2045)
);

AOI22xp33_ASAP7_75t_L g2046 ( 
.A1(n_2028),
.A2(n_1916),
.B1(n_1814),
.B2(n_1898),
.Y(n_2046)
);

NAND3xp33_ASAP7_75t_L g2047 ( 
.A(n_2033),
.B(n_202),
.C(n_207),
.Y(n_2047)
);

AND2x2_ASAP7_75t_L g2048 ( 
.A(n_2030),
.B(n_1912),
.Y(n_2048)
);

AOI22xp5_ASAP7_75t_L g2049 ( 
.A1(n_2025),
.A2(n_1916),
.B1(n_1791),
.B2(n_1926),
.Y(n_2049)
);

NOR3xp33_ASAP7_75t_L g2050 ( 
.A(n_2025),
.B(n_207),
.C(n_208),
.Y(n_2050)
);

NOR2x1_ASAP7_75t_L g2051 ( 
.A(n_2047),
.B(n_208),
.Y(n_2051)
);

NOR2x1_ASAP7_75t_L g2052 ( 
.A(n_2040),
.B(n_209),
.Y(n_2052)
);

NOR3x2_ASAP7_75t_L g2053 ( 
.A(n_2050),
.B(n_209),
.C(n_210),
.Y(n_2053)
);

OAI222xp33_ASAP7_75t_L g2054 ( 
.A1(n_2036),
.A2(n_1764),
.B1(n_1811),
.B2(n_1926),
.C1(n_1749),
.C2(n_1861),
.Y(n_2054)
);

HB1xp67_ASAP7_75t_L g2055 ( 
.A(n_2038),
.Y(n_2055)
);

INVx1_ASAP7_75t_L g2056 ( 
.A(n_2045),
.Y(n_2056)
);

INVx1_ASAP7_75t_L g2057 ( 
.A(n_2037),
.Y(n_2057)
);

NOR3xp33_ASAP7_75t_L g2058 ( 
.A(n_2039),
.B(n_210),
.C(n_1628),
.Y(n_2058)
);

NAND3x2_ASAP7_75t_L g2059 ( 
.A(n_2043),
.B(n_1914),
.C(n_1858),
.Y(n_2059)
);

OR2x2_ASAP7_75t_L g2060 ( 
.A(n_2048),
.B(n_1900),
.Y(n_2060)
);

NAND2xp5_ASAP7_75t_SL g2061 ( 
.A(n_2042),
.B(n_1922),
.Y(n_2061)
);

NOR3xp33_ASAP7_75t_L g2062 ( 
.A(n_2044),
.B(n_1616),
.C(n_1617),
.Y(n_2062)
);

NOR3xp33_ASAP7_75t_L g2063 ( 
.A(n_2041),
.B(n_1620),
.C(n_1651),
.Y(n_2063)
);

NOR3xp33_ASAP7_75t_L g2064 ( 
.A(n_2049),
.B(n_1722),
.C(n_1713),
.Y(n_2064)
);

OAI21xp5_ASAP7_75t_SL g2065 ( 
.A1(n_2046),
.A2(n_1885),
.B(n_1861),
.Y(n_2065)
);

INVx2_ASAP7_75t_L g2066 ( 
.A(n_2048),
.Y(n_2066)
);

NAND4xp75_ASAP7_75t_L g2067 ( 
.A(n_2040),
.B(n_1748),
.C(n_1767),
.D(n_1895),
.Y(n_2067)
);

OAI21xp33_ASAP7_75t_L g2068 ( 
.A1(n_2045),
.A2(n_1893),
.B(n_1904),
.Y(n_2068)
);

INVx2_ASAP7_75t_L g2069 ( 
.A(n_2048),
.Y(n_2069)
);

AND2x4_ASAP7_75t_L g2070 ( 
.A(n_2040),
.B(n_1804),
.Y(n_2070)
);

NOR2x1_ASAP7_75t_L g2071 ( 
.A(n_2047),
.B(n_383),
.Y(n_2071)
);

NAND2xp5_ASAP7_75t_L g2072 ( 
.A(n_2070),
.B(n_1900),
.Y(n_2072)
);

NOR3xp33_ASAP7_75t_L g2073 ( 
.A(n_2056),
.B(n_1876),
.C(n_1906),
.Y(n_2073)
);

AND2x4_ASAP7_75t_L g2074 ( 
.A(n_2070),
.B(n_1906),
.Y(n_2074)
);

NOR3xp33_ASAP7_75t_L g2075 ( 
.A(n_2057),
.B(n_1840),
.C(n_1835),
.Y(n_2075)
);

NAND2xp5_ASAP7_75t_SL g2076 ( 
.A(n_2052),
.B(n_1919),
.Y(n_2076)
);

NOR3xp33_ASAP7_75t_L g2077 ( 
.A(n_2066),
.B(n_1840),
.C(n_385),
.Y(n_2077)
);

NAND3xp33_ASAP7_75t_SL g2078 ( 
.A(n_2069),
.B(n_2055),
.C(n_2068),
.Y(n_2078)
);

INVx1_ASAP7_75t_SL g2079 ( 
.A(n_2053),
.Y(n_2079)
);

HB1xp67_ASAP7_75t_L g2080 ( 
.A(n_2051),
.Y(n_2080)
);

NOR4xp25_ASAP7_75t_L g2081 ( 
.A(n_2061),
.B(n_1914),
.C(n_1919),
.D(n_1922),
.Y(n_2081)
);

NOR3xp33_ASAP7_75t_L g2082 ( 
.A(n_2071),
.B(n_388),
.C(n_390),
.Y(n_2082)
);

INVx1_ASAP7_75t_L g2083 ( 
.A(n_2067),
.Y(n_2083)
);

INVx1_ASAP7_75t_L g2084 ( 
.A(n_2060),
.Y(n_2084)
);

NAND2xp5_ASAP7_75t_L g2085 ( 
.A(n_2065),
.B(n_1900),
.Y(n_2085)
);

INVx1_ASAP7_75t_L g2086 ( 
.A(n_2080),
.Y(n_2086)
);

NOR2x1_ASAP7_75t_L g2087 ( 
.A(n_2078),
.B(n_2079),
.Y(n_2087)
);

AOI22xp5_ASAP7_75t_L g2088 ( 
.A1(n_2082),
.A2(n_2062),
.B1(n_2059),
.B2(n_2058),
.Y(n_2088)
);

INVx1_ASAP7_75t_L g2089 ( 
.A(n_2076),
.Y(n_2089)
);

OR2x2_ASAP7_75t_L g2090 ( 
.A(n_2074),
.B(n_2081),
.Y(n_2090)
);

XOR2x1_ASAP7_75t_L g2091 ( 
.A(n_2084),
.B(n_2054),
.Y(n_2091)
);

INVx1_ASAP7_75t_L g2092 ( 
.A(n_2083),
.Y(n_2092)
);

AND2x4_ASAP7_75t_L g2093 ( 
.A(n_2074),
.B(n_2073),
.Y(n_2093)
);

AOI22xp5_ASAP7_75t_L g2094 ( 
.A1(n_2077),
.A2(n_2075),
.B1(n_2072),
.B2(n_2085),
.Y(n_2094)
);

INVx2_ASAP7_75t_L g2095 ( 
.A(n_2074),
.Y(n_2095)
);

INVx1_ASAP7_75t_L g2096 ( 
.A(n_2080),
.Y(n_2096)
);

INVx2_ASAP7_75t_L g2097 ( 
.A(n_2074),
.Y(n_2097)
);

NAND2xp5_ASAP7_75t_L g2098 ( 
.A(n_2079),
.B(n_2064),
.Y(n_2098)
);

INVx2_ASAP7_75t_L g2099 ( 
.A(n_2074),
.Y(n_2099)
);

XNOR2xp5_ASAP7_75t_L g2100 ( 
.A(n_2078),
.B(n_2063),
.Y(n_2100)
);

NOR2x1_ASAP7_75t_L g2101 ( 
.A(n_2078),
.B(n_391),
.Y(n_2101)
);

INVx1_ASAP7_75t_L g2102 ( 
.A(n_2087),
.Y(n_2102)
);

NAND4xp25_ASAP7_75t_L g2103 ( 
.A(n_2086),
.B(n_1870),
.C(n_395),
.D(n_396),
.Y(n_2103)
);

AOI22xp33_ASAP7_75t_L g2104 ( 
.A1(n_2096),
.A2(n_1898),
.B1(n_1900),
.B2(n_1895),
.Y(n_2104)
);

AO22x2_ASAP7_75t_L g2105 ( 
.A1(n_2095),
.A2(n_1919),
.B1(n_1922),
.B2(n_1884),
.Y(n_2105)
);

INVx1_ASAP7_75t_L g2106 ( 
.A(n_2101),
.Y(n_2106)
);

CKINVDCx5p33_ASAP7_75t_R g2107 ( 
.A(n_2092),
.Y(n_2107)
);

NOR2xp67_ASAP7_75t_SL g2108 ( 
.A(n_2097),
.B(n_393),
.Y(n_2108)
);

CKINVDCx20_ASAP7_75t_R g2109 ( 
.A(n_2100),
.Y(n_2109)
);

NAND2xp5_ASAP7_75t_L g2110 ( 
.A(n_2099),
.B(n_397),
.Y(n_2110)
);

NAND2x1_ASAP7_75t_L g2111 ( 
.A(n_2090),
.B(n_1889),
.Y(n_2111)
);

HB1xp67_ASAP7_75t_L g2112 ( 
.A(n_2091),
.Y(n_2112)
);

AND2x4_ASAP7_75t_L g2113 ( 
.A(n_2093),
.B(n_1889),
.Y(n_2113)
);

NOR3xp33_ASAP7_75t_SL g2114 ( 
.A(n_2098),
.B(n_398),
.C(n_400),
.Y(n_2114)
);

AOI21xp5_ASAP7_75t_L g2115 ( 
.A1(n_2102),
.A2(n_2089),
.B(n_2094),
.Y(n_2115)
);

AOI322xp5_ASAP7_75t_L g2116 ( 
.A1(n_2112),
.A2(n_2088),
.A3(n_1929),
.B1(n_1928),
.B2(n_1901),
.C1(n_1891),
.C2(n_1884),
.Y(n_2116)
);

OAI221xp5_ASAP7_75t_SL g2117 ( 
.A1(n_2106),
.A2(n_1891),
.B1(n_1902),
.B2(n_1883),
.C(n_1901),
.Y(n_2117)
);

OAI22xp5_ASAP7_75t_L g2118 ( 
.A1(n_2109),
.A2(n_1902),
.B1(n_1886),
.B2(n_1888),
.Y(n_2118)
);

NAND2xp5_ASAP7_75t_L g2119 ( 
.A(n_2113),
.B(n_402),
.Y(n_2119)
);

AOI221xp5_ASAP7_75t_L g2120 ( 
.A1(n_2107),
.A2(n_1902),
.B1(n_1888),
.B2(n_1899),
.C(n_1886),
.Y(n_2120)
);

NAND3xp33_ASAP7_75t_SL g2121 ( 
.A(n_2110),
.B(n_403),
.C(n_404),
.Y(n_2121)
);

INVx2_ASAP7_75t_L g2122 ( 
.A(n_2111),
.Y(n_2122)
);

NOR4xp25_ASAP7_75t_L g2123 ( 
.A(n_2103),
.B(n_405),
.C(n_406),
.D(n_408),
.Y(n_2123)
);

NOR4xp25_ASAP7_75t_L g2124 ( 
.A(n_2114),
.B(n_409),
.C(n_411),
.D(n_412),
.Y(n_2124)
);

INVx1_ASAP7_75t_L g2125 ( 
.A(n_2108),
.Y(n_2125)
);

NOR3xp33_ASAP7_75t_L g2126 ( 
.A(n_2105),
.B(n_414),
.C(n_416),
.Y(n_2126)
);

OAI22xp5_ASAP7_75t_L g2127 ( 
.A1(n_2104),
.A2(n_1886),
.B1(n_1888),
.B2(n_1892),
.Y(n_2127)
);

O2A1O1Ixp33_ASAP7_75t_L g2128 ( 
.A1(n_2122),
.A2(n_418),
.B(n_419),
.C(n_420),
.Y(n_2128)
);

AOI22xp5_ASAP7_75t_L g2129 ( 
.A1(n_2125),
.A2(n_1898),
.B1(n_1889),
.B2(n_1903),
.Y(n_2129)
);

AOI221x1_ASAP7_75t_L g2130 ( 
.A1(n_2115),
.A2(n_421),
.B1(n_422),
.B2(n_423),
.C(n_424),
.Y(n_2130)
);

OAI22xp5_ASAP7_75t_SL g2131 ( 
.A1(n_2124),
.A2(n_426),
.B1(n_427),
.B2(n_428),
.Y(n_2131)
);

AOI22xp5_ASAP7_75t_L g2132 ( 
.A1(n_2121),
.A2(n_1898),
.B1(n_1903),
.B2(n_1886),
.Y(n_2132)
);

OAI221xp5_ASAP7_75t_L g2133 ( 
.A1(n_2123),
.A2(n_1892),
.B1(n_432),
.B2(n_435),
.C(n_437),
.Y(n_2133)
);

INVx2_ASAP7_75t_L g2134 ( 
.A(n_2119),
.Y(n_2134)
);

NAND4xp25_ASAP7_75t_L g2135 ( 
.A(n_2126),
.B(n_429),
.C(n_438),
.D(n_440),
.Y(n_2135)
);

INVx2_ASAP7_75t_L g2136 ( 
.A(n_2134),
.Y(n_2136)
);

OAI21xp5_ASAP7_75t_L g2137 ( 
.A1(n_2133),
.A2(n_2127),
.B(n_2116),
.Y(n_2137)
);

HB1xp67_ASAP7_75t_L g2138 ( 
.A(n_2131),
.Y(n_2138)
);

NAND2xp5_ASAP7_75t_L g2139 ( 
.A(n_2135),
.B(n_2118),
.Y(n_2139)
);

NAND2xp5_ASAP7_75t_L g2140 ( 
.A(n_2130),
.B(n_2120),
.Y(n_2140)
);

AO22x2_ASAP7_75t_L g2141 ( 
.A1(n_2128),
.A2(n_2117),
.B1(n_442),
.B2(n_444),
.Y(n_2141)
);

AOI21xp5_ASAP7_75t_L g2142 ( 
.A1(n_2132),
.A2(n_441),
.B(n_445),
.Y(n_2142)
);

NAND2xp5_ASAP7_75t_L g2143 ( 
.A(n_2129),
.B(n_448),
.Y(n_2143)
);

INVx1_ASAP7_75t_L g2144 ( 
.A(n_2131),
.Y(n_2144)
);

O2A1O1Ixp33_ASAP7_75t_L g2145 ( 
.A1(n_2138),
.A2(n_449),
.B(n_454),
.C(n_455),
.Y(n_2145)
);

NOR3x1_ASAP7_75t_L g2146 ( 
.A(n_2144),
.B(n_2137),
.C(n_2140),
.Y(n_2146)
);

INVxp67_ASAP7_75t_SL g2147 ( 
.A(n_2136),
.Y(n_2147)
);

XNOR2xp5_ASAP7_75t_L g2148 ( 
.A(n_2141),
.B(n_457),
.Y(n_2148)
);

NOR2x1_ASAP7_75t_L g2149 ( 
.A(n_2143),
.B(n_458),
.Y(n_2149)
);

OAI22xp5_ASAP7_75t_L g2150 ( 
.A1(n_2147),
.A2(n_2139),
.B1(n_2142),
.B2(n_1892),
.Y(n_2150)
);

AOI222xp33_ASAP7_75t_SL g2151 ( 
.A1(n_2146),
.A2(n_459),
.B1(n_460),
.B2(n_461),
.C1(n_463),
.C2(n_464),
.Y(n_2151)
);

AOI22xp33_ASAP7_75t_SL g2152 ( 
.A1(n_2150),
.A2(n_2148),
.B1(n_2149),
.B2(n_2145),
.Y(n_2152)
);

OAI21xp5_ASAP7_75t_L g2153 ( 
.A1(n_2152),
.A2(n_2151),
.B(n_468),
.Y(n_2153)
);

INVx1_ASAP7_75t_L g2154 ( 
.A(n_2153),
.Y(n_2154)
);

OR2x2_ASAP7_75t_L g2155 ( 
.A(n_2154),
.B(n_465),
.Y(n_2155)
);

AOI21xp33_ASAP7_75t_SL g2156 ( 
.A1(n_2155),
.A2(n_469),
.B(n_471),
.Y(n_2156)
);

AOI211xp5_ASAP7_75t_L g2157 ( 
.A1(n_2156),
.A2(n_473),
.B(n_475),
.C(n_476),
.Y(n_2157)
);


endmodule