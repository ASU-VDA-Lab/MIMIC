module fake_netlist_6_517_n_1119 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_193, n_147, n_154, n_191, n_88, n_3, n_209, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_199, n_138, n_22, n_161, n_208, n_68, n_166, n_28, n_184, n_212, n_50, n_158, n_49, n_7, n_210, n_216, n_83, n_206, n_217, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_215, n_178, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_188, n_102, n_186, n_204, n_0, n_87, n_195, n_189, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_213, n_164, n_100, n_129, n_13, n_121, n_197, n_11, n_137, n_17, n_23, n_203, n_142, n_20, n_143, n_207, n_2, n_180, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_205, n_34, n_140, n_218, n_70, n_120, n_214, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_181, n_76, n_36, n_182, n_26, n_124, n_55, n_126, n_202, n_94, n_97, n_108, n_58, n_116, n_211, n_64, n_117, n_118, n_175, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_196, n_200, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_198, n_104, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_6, n_190, n_14, n_123, n_136, n_72, n_187, n_89, n_173, n_201, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_185, n_35, n_183, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_194, n_171, n_31, n_192, n_57, n_169, n_53, n_51, n_44, n_56, n_1119);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_193;
input n_147;
input n_154;
input n_191;
input n_88;
input n_3;
input n_209;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_199;
input n_138;
input n_22;
input n_161;
input n_208;
input n_68;
input n_166;
input n_28;
input n_184;
input n_212;
input n_50;
input n_158;
input n_49;
input n_7;
input n_210;
input n_216;
input n_83;
input n_206;
input n_217;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_215;
input n_178;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_188;
input n_102;
input n_186;
input n_204;
input n_0;
input n_87;
input n_195;
input n_189;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_213;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_197;
input n_11;
input n_137;
input n_17;
input n_23;
input n_203;
input n_142;
input n_20;
input n_143;
input n_207;
input n_2;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_205;
input n_34;
input n_140;
input n_218;
input n_70;
input n_120;
input n_214;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_55;
input n_126;
input n_202;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_211;
input n_64;
input n_117;
input n_118;
input n_175;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_196;
input n_200;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_190;
input n_14;
input n_123;
input n_136;
input n_72;
input n_187;
input n_89;
input n_173;
input n_201;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_185;
input n_35;
input n_183;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_194;
input n_171;
input n_31;
input n_192;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1119;

wire n_992;
wire n_591;
wire n_435;
wire n_1115;
wire n_793;
wire n_326;
wire n_801;
wire n_256;
wire n_853;
wire n_440;
wire n_587;
wire n_695;
wire n_507;
wire n_968;
wire n_909;
wire n_580;
wire n_762;
wire n_1030;
wire n_881;
wire n_1008;
wire n_465;
wire n_367;
wire n_680;
wire n_741;
wire n_760;
wire n_875;
wire n_1027;
wire n_590;
wire n_625;
wire n_661;
wire n_223;
wire n_278;
wire n_1079;
wire n_341;
wire n_362;
wire n_226;
wire n_828;
wire n_462;
wire n_607;
wire n_671;
wire n_726;
wire n_1033;
wire n_316;
wire n_419;
wire n_304;
wire n_700;
wire n_694;
wire n_1103;
wire n_933;
wire n_740;
wire n_1038;
wire n_578;
wire n_703;
wire n_1003;
wire n_365;
wire n_978;
wire n_1061;
wire n_384;
wire n_297;
wire n_595;
wire n_627;
wire n_524;
wire n_342;
wire n_820;
wire n_1044;
wire n_951;
wire n_783;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_751;
wire n_449;
wire n_749;
wire n_798;
wire n_310;
wire n_509;
wire n_245;
wire n_368;
wire n_575;
wire n_994;
wire n_1072;
wire n_677;
wire n_988;
wire n_969;
wire n_805;
wire n_396;
wire n_495;
wire n_1065;
wire n_815;
wire n_350;
wire n_1100;
wire n_585;
wire n_732;
wire n_974;
wire n_568;
wire n_392;
wire n_840;
wire n_442;
wire n_480;
wire n_874;
wire n_724;
wire n_382;
wire n_673;
wire n_1020;
wire n_1009;
wire n_1042;
wire n_1071;
wire n_628;
wire n_1067;
wire n_883;
wire n_557;
wire n_823;
wire n_349;
wire n_643;
wire n_233;
wire n_617;
wire n_698;
wire n_898;
wire n_1074;
wire n_1032;
wire n_845;
wire n_255;
wire n_807;
wire n_1036;
wire n_739;
wire n_284;
wire n_400;
wire n_337;
wire n_955;
wire n_865;
wire n_893;
wire n_925;
wire n_485;
wire n_1099;
wire n_1026;
wire n_443;
wire n_1101;
wire n_246;
wire n_892;
wire n_768;
wire n_1097;
wire n_471;
wire n_289;
wire n_935;
wire n_421;
wire n_781;
wire n_424;
wire n_789;
wire n_615;
wire n_238;
wire n_1095;
wire n_573;
wire n_769;
wire n_320;
wire n_639;
wire n_676;
wire n_327;
wire n_794;
wire n_963;
wire n_727;
wire n_894;
wire n_369;
wire n_597;
wire n_685;
wire n_280;
wire n_287;
wire n_832;
wire n_353;
wire n_610;
wire n_555;
wire n_389;
wire n_814;
wire n_415;
wire n_830;
wire n_230;
wire n_605;
wire n_461;
wire n_873;
wire n_383;
wire n_826;
wire n_1024;
wire n_669;
wire n_447;
wire n_872;
wire n_300;
wire n_222;
wire n_718;
wire n_248;
wire n_517;
wire n_1018;
wire n_747;
wire n_852;
wire n_667;
wire n_229;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_1105;
wire n_621;
wire n_305;
wire n_1037;
wire n_721;
wire n_996;
wire n_750;
wire n_532;
wire n_742;
wire n_535;
wire n_691;
wire n_901;
wire n_250;
wire n_372;
wire n_468;
wire n_544;
wire n_1078;
wire n_504;
wire n_923;
wire n_314;
wire n_378;
wire n_413;
wire n_377;
wire n_791;
wire n_510;
wire n_837;
wire n_836;
wire n_1015;
wire n_863;
wire n_375;
wire n_601;
wire n_338;
wire n_522;
wire n_948;
wire n_466;
wire n_704;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_763;
wire n_1057;
wire n_360;
wire n_977;
wire n_945;
wire n_603;
wire n_1005;
wire n_991;
wire n_957;
wire n_235;
wire n_536;
wire n_895;
wire n_866;
wire n_622;
wire n_340;
wire n_710;
wire n_1108;
wire n_387;
wire n_452;
wire n_658;
wire n_616;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_581;
wire n_428;
wire n_785;
wire n_761;
wire n_746;
wire n_609;
wire n_765;
wire n_432;
wire n_987;
wire n_641;
wire n_822;
wire n_693;
wire n_1056;
wire n_631;
wire n_516;
wire n_720;
wire n_758;
wire n_525;
wire n_842;
wire n_1116;
wire n_611;
wire n_943;
wire n_491;
wire n_878;
wire n_772;
wire n_656;
wire n_843;
wire n_989;
wire n_797;
wire n_666;
wire n_1016;
wire n_371;
wire n_795;
wire n_770;
wire n_940;
wire n_567;
wire n_899;
wire n_738;
wire n_405;
wire n_538;
wire n_1035;
wire n_294;
wire n_302;
wire n_499;
wire n_380;
wire n_838;
wire n_705;
wire n_647;
wire n_343;
wire n_844;
wire n_448;
wire n_886;
wire n_953;
wire n_1004;
wire n_1017;
wire n_1094;
wire n_494;
wire n_539;
wire n_493;
wire n_397;
wire n_1022;
wire n_1083;
wire n_614;
wire n_529;
wire n_445;
wire n_425;
wire n_684;
wire n_930;
wire n_888;
wire n_1112;
wire n_454;
wire n_638;
wire n_234;
wire n_910;
wire n_486;
wire n_911;
wire n_381;
wire n_947;
wire n_236;
wire n_653;
wire n_887;
wire n_1117;
wire n_1087;
wire n_752;
wire n_908;
wire n_944;
wire n_713;
wire n_648;
wire n_657;
wire n_1049;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_239;
wire n_414;
wire n_563;
wire n_782;
wire n_976;
wire n_490;
wire n_803;
wire n_290;
wire n_220;
wire n_809;
wire n_1043;
wire n_1011;
wire n_224;
wire n_926;
wire n_927;
wire n_839;
wire n_986;
wire n_734;
wire n_1088;
wire n_708;
wire n_919;
wire n_1081;
wire n_402;
wire n_352;
wire n_917;
wire n_668;
wire n_478;
wire n_626;
wire n_990;
wire n_574;
wire n_800;
wire n_779;
wire n_929;
wire n_460;
wire n_1084;
wire n_1104;
wire n_907;
wire n_854;
wire n_1058;
wire n_417;
wire n_446;
wire n_498;
wire n_662;
wire n_374;
wire n_659;
wire n_709;
wire n_904;
wire n_366;
wire n_870;
wire n_777;
wire n_407;
wire n_913;
wire n_450;
wire n_808;
wire n_867;
wire n_272;
wire n_526;
wire n_1109;
wire n_921;
wire n_712;
wire n_348;
wire n_711;
wire n_579;
wire n_376;
wire n_937;
wire n_390;
wire n_473;
wire n_293;
wire n_1054;
wire n_334;
wire n_559;
wire n_370;
wire n_458;
wire n_1070;
wire n_1085;
wire n_232;
wire n_650;
wire n_998;
wire n_1046;
wire n_717;
wire n_330;
wire n_771;
wire n_470;
wire n_475;
wire n_924;
wire n_1102;
wire n_298;
wire n_492;
wire n_972;
wire n_281;
wire n_258;
wire n_551;
wire n_699;
wire n_456;
wire n_564;
wire n_260;
wire n_265;
wire n_313;
wire n_451;
wire n_624;
wire n_824;
wire n_962;
wire n_1073;
wire n_1000;
wire n_279;
wire n_686;
wire n_796;
wire n_1041;
wire n_252;
wire n_757;
wire n_228;
wire n_565;
wire n_594;
wire n_719;
wire n_356;
wire n_577;
wire n_936;
wire n_552;
wire n_1062;
wire n_619;
wire n_885;
wire n_455;
wire n_896;
wire n_521;
wire n_363;
wire n_572;
wire n_912;
wire n_395;
wire n_813;
wire n_592;
wire n_1090;
wire n_745;
wire n_654;
wire n_323;
wire n_829;
wire n_606;
wire n_393;
wire n_984;
wire n_818;
wire n_411;
wire n_503;
wire n_716;
wire n_623;
wire n_1048;
wire n_884;
wire n_599;
wire n_513;
wire n_855;
wire n_776;
wire n_321;
wire n_645;
wire n_331;
wire n_916;
wire n_227;
wire n_868;
wire n_570;
wire n_731;
wire n_859;
wire n_406;
wire n_483;
wire n_735;
wire n_482;
wire n_934;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_527;
wire n_261;
wire n_608;
wire n_620;
wire n_420;
wire n_683;
wire n_630;
wire n_312;
wire n_394;
wire n_519;
wire n_541;
wire n_512;
wire n_958;
wire n_292;
wire n_307;
wire n_469;
wire n_433;
wire n_500;
wire n_942;
wire n_792;
wire n_880;
wire n_476;
wire n_981;
wire n_714;
wire n_291;
wire n_219;
wire n_543;
wire n_889;
wire n_357;
wire n_264;
wire n_263;
wire n_985;
wire n_589;
wire n_860;
wire n_481;
wire n_788;
wire n_819;
wire n_939;
wire n_997;
wire n_821;
wire n_325;
wire n_938;
wire n_1068;
wire n_767;
wire n_804;
wire n_329;
wire n_464;
wire n_600;
wire n_831;
wire n_802;
wire n_964;
wire n_982;
wire n_561;
wire n_477;
wire n_549;
wire n_980;
wire n_533;
wire n_954;
wire n_1075;
wire n_408;
wire n_932;
wire n_806;
wire n_864;
wire n_879;
wire n_959;
wire n_237;
wire n_584;
wire n_1110;
wire n_244;
wire n_399;
wire n_243;
wire n_979;
wire n_548;
wire n_905;
wire n_282;
wire n_436;
wire n_833;
wire n_523;
wire n_322;
wire n_707;
wire n_993;
wire n_345;
wire n_409;
wire n_231;
wire n_354;
wire n_689;
wire n_799;
wire n_505;
wire n_240;
wire n_756;
wire n_319;
wire n_547;
wire n_537;
wire n_273;
wire n_558;
wire n_810;
wire n_635;
wire n_787;
wire n_311;
wire n_1064;
wire n_403;
wire n_1080;
wire n_723;
wire n_253;
wire n_634;
wire n_1051;
wire n_583;
wire n_596;
wire n_966;
wire n_546;
wire n_562;
wire n_249;
wire n_386;
wire n_764;
wire n_1039;
wire n_556;
wire n_1034;
wire n_1086;
wire n_1066;
wire n_692;
wire n_733;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_487;
wire n_550;
wire n_241;
wire n_275;
wire n_553;
wire n_652;
wire n_849;
wire n_970;
wire n_1107;
wire n_560;
wire n_1014;
wire n_753;
wire n_642;
wire n_995;
wire n_276;
wire n_569;
wire n_1092;
wire n_441;
wire n_221;
wire n_811;
wire n_1060;
wire n_882;
wire n_444;
wire n_586;
wire n_423;
wire n_737;
wire n_318;
wire n_1111;
wire n_303;
wire n_511;
wire n_715;
wire n_467;
wire n_306;
wire n_269;
wire n_359;
wire n_973;
wire n_346;
wire n_416;
wire n_1053;
wire n_530;
wire n_277;
wire n_520;
wire n_1029;
wire n_418;
wire n_1093;
wire n_618;
wire n_1055;
wire n_790;
wire n_1106;
wire n_582;
wire n_266;
wire n_296;
wire n_861;
wire n_674;
wire n_857;
wire n_871;
wire n_967;
wire n_775;
wire n_922;
wire n_571;
wire n_268;
wire n_271;
wire n_404;
wire n_651;
wire n_439;
wire n_299;
wire n_518;
wire n_679;
wire n_1069;
wire n_453;
wire n_612;
wire n_633;
wire n_665;
wire n_902;
wire n_333;
wire n_588;
wire n_247;
wire n_225;
wire n_308;
wire n_309;
wire n_914;
wire n_759;
wire n_1047;
wire n_1010;
wire n_355;
wire n_426;
wire n_317;
wire n_1040;
wire n_915;
wire n_632;
wire n_702;
wire n_431;
wire n_347;
wire n_812;
wire n_459;
wire n_1052;
wire n_502;
wire n_328;
wire n_672;
wire n_534;
wire n_488;
wire n_429;
wire n_1006;
wire n_373;
wire n_1012;
wire n_497;
wire n_285;
wire n_780;
wire n_773;
wire n_675;
wire n_920;
wire n_257;
wire n_903;
wire n_730;
wire n_655;
wire n_706;
wire n_1045;
wire n_786;
wire n_670;
wire n_286;
wire n_254;
wire n_834;
wire n_242;
wire n_835;
wire n_928;
wire n_690;
wire n_850;
wire n_1089;
wire n_401;
wire n_324;
wire n_766;
wire n_743;
wire n_816;
wire n_335;
wire n_430;
wire n_1002;
wire n_463;
wire n_545;
wire n_489;
wire n_877;
wire n_604;
wire n_848;
wire n_251;
wire n_1019;
wire n_301;
wire n_274;
wire n_636;
wire n_825;
wire n_728;
wire n_681;
wire n_1096;
wire n_1063;
wire n_729;
wire n_1091;
wire n_876;
wire n_774;
wire n_412;
wire n_640;
wire n_660;
wire n_965;
wire n_267;
wire n_438;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_515;
wire n_983;
wire n_288;
wire n_427;
wire n_1059;
wire n_479;
wire n_496;
wire n_598;
wire n_422;
wire n_696;
wire n_906;
wire n_722;
wire n_688;
wire n_1077;
wire n_961;
wire n_862;
wire n_351;
wire n_869;
wire n_437;
wire n_1082;
wire n_259;
wire n_1113;
wire n_540;
wire n_593;
wire n_514;
wire n_646;
wire n_528;
wire n_457;
wire n_391;
wire n_1098;
wire n_697;
wire n_687;
wire n_364;
wire n_890;
wire n_637;
wire n_295;
wire n_385;
wire n_701;
wire n_817;
wire n_950;
wire n_629;
wire n_388;
wire n_858;
wire n_262;
wire n_484;
wire n_613;
wire n_736;
wire n_897;
wire n_900;
wire n_846;
wire n_501;
wire n_841;
wire n_956;
wire n_960;
wire n_531;
wire n_1001;
wire n_827;
wire n_508;
wire n_361;
wire n_663;
wire n_856;
wire n_1050;
wire n_379;
wire n_778;
wire n_1025;
wire n_332;
wire n_891;
wire n_336;
wire n_398;
wire n_410;
wire n_566;
wire n_554;
wire n_602;
wire n_1013;
wire n_1023;
wire n_1076;
wire n_1118;
wire n_664;
wire n_949;
wire n_678;
wire n_1007;
wire n_649;
wire n_283;

BUFx2_ASAP7_75t_L g219 ( 
.A(n_33),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_139),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_143),
.Y(n_221)
);

BUFx6f_ASAP7_75t_L g222 ( 
.A(n_215),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_136),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_50),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_166),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_98),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_174),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_208),
.Y(n_228)
);

BUFx6f_ASAP7_75t_L g229 ( 
.A(n_76),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_111),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_13),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_54),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_116),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_190),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_185),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_52),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_218),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_106),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_184),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_124),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_201),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_129),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_99),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_78),
.Y(n_244)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_132),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_189),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_110),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_17),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_75),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_175),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_74),
.Y(n_251)
);

BUFx6f_ASAP7_75t_L g252 ( 
.A(n_23),
.Y(n_252)
);

INVxp67_ASAP7_75t_L g253 ( 
.A(n_117),
.Y(n_253)
);

BUFx3_ASAP7_75t_L g254 ( 
.A(n_144),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_5),
.Y(n_255)
);

BUFx2_ASAP7_75t_SL g256 ( 
.A(n_5),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_141),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_172),
.Y(n_258)
);

BUFx3_ASAP7_75t_L g259 ( 
.A(n_49),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_85),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_182),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_40),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_165),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_181),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_151),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_88),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_80),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_194),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_207),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_35),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_93),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_146),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_134),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_79),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_34),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_55),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_140),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_22),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_96),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_196),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_119),
.Y(n_281)
);

BUFx6f_ASAP7_75t_L g282 ( 
.A(n_63),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_84),
.Y(n_283)
);

INVx1_ASAP7_75t_SL g284 ( 
.A(n_210),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_43),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_66),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_41),
.Y(n_287)
);

INVx1_ASAP7_75t_SL g288 ( 
.A(n_125),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g289 ( 
.A(n_1),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_252),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_252),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_221),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_252),
.Y(n_293)
);

INVxp67_ASAP7_75t_SL g294 ( 
.A(n_219),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_223),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g296 ( 
.A(n_289),
.Y(n_296)
);

INVxp33_ASAP7_75t_L g297 ( 
.A(n_278),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_252),
.Y(n_298)
);

INVxp67_ASAP7_75t_SL g299 ( 
.A(n_254),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_254),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_259),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_259),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_220),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_226),
.Y(n_304)
);

CKINVDCx16_ASAP7_75t_R g305 ( 
.A(n_225),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_224),
.Y(n_306)
);

INVxp33_ASAP7_75t_SL g307 ( 
.A(n_256),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_232),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_231),
.Y(n_309)
);

INVxp67_ASAP7_75t_SL g310 ( 
.A(n_253),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_248),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_234),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_247),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_257),
.Y(n_314)
);

HB1xp67_ASAP7_75t_L g315 ( 
.A(n_255),
.Y(n_315)
);

INVxp67_ASAP7_75t_SL g316 ( 
.A(n_264),
.Y(n_316)
);

CKINVDCx16_ASAP7_75t_R g317 ( 
.A(n_239),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_242),
.Y(n_318)
);

BUFx6f_ASAP7_75t_L g319 ( 
.A(n_222),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_227),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_268),
.Y(n_321)
);

INVxp33_ASAP7_75t_SL g322 ( 
.A(n_228),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_230),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_272),
.Y(n_324)
);

CKINVDCx16_ASAP7_75t_R g325 ( 
.A(n_263),
.Y(n_325)
);

CKINVDCx16_ASAP7_75t_R g326 ( 
.A(n_270),
.Y(n_326)
);

CKINVDCx16_ASAP7_75t_R g327 ( 
.A(n_222),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g328 ( 
.A(n_233),
.Y(n_328)
);

BUFx3_ASAP7_75t_L g329 ( 
.A(n_275),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_277),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_283),
.Y(n_331)
);

INVxp67_ASAP7_75t_SL g332 ( 
.A(n_245),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_235),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_236),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_222),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_222),
.Y(n_336)
);

CKINVDCx20_ASAP7_75t_R g337 ( 
.A(n_237),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_335),
.Y(n_338)
);

BUFx6f_ASAP7_75t_L g339 ( 
.A(n_319),
.Y(n_339)
);

INVx2_ASAP7_75t_L g340 ( 
.A(n_319),
.Y(n_340)
);

INVx2_ASAP7_75t_L g341 ( 
.A(n_319),
.Y(n_341)
);

BUFx6f_ASAP7_75t_L g342 ( 
.A(n_319),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_L g343 ( 
.A(n_322),
.B(n_284),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_336),
.Y(n_344)
);

AND2x4_ASAP7_75t_L g345 ( 
.A(n_316),
.B(n_229),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_290),
.Y(n_346)
);

AND2x2_ASAP7_75t_L g347 ( 
.A(n_299),
.B(n_288),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_327),
.B(n_287),
.Y(n_348)
);

HB1xp67_ASAP7_75t_L g349 ( 
.A(n_315),
.Y(n_349)
);

BUFx3_ASAP7_75t_L g350 ( 
.A(n_291),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_293),
.Y(n_351)
);

OAI21x1_ASAP7_75t_L g352 ( 
.A1(n_303),
.A2(n_282),
.B(n_229),
.Y(n_352)
);

BUFx6f_ASAP7_75t_L g353 ( 
.A(n_298),
.Y(n_353)
);

OA21x2_ASAP7_75t_L g354 ( 
.A1(n_306),
.A2(n_312),
.B(n_308),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_313),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_292),
.Y(n_356)
);

INVx2_ASAP7_75t_L g357 ( 
.A(n_314),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_321),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_324),
.Y(n_359)
);

AND2x2_ASAP7_75t_L g360 ( 
.A(n_300),
.B(n_238),
.Y(n_360)
);

NOR2x1_ASAP7_75t_L g361 ( 
.A(n_329),
.B(n_229),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_330),
.Y(n_362)
);

AND2x2_ASAP7_75t_L g363 ( 
.A(n_301),
.B(n_240),
.Y(n_363)
);

OAI21x1_ASAP7_75t_L g364 ( 
.A1(n_331),
.A2(n_282),
.B(n_229),
.Y(n_364)
);

BUFx6f_ASAP7_75t_L g365 ( 
.A(n_329),
.Y(n_365)
);

INVx2_ASAP7_75t_L g366 ( 
.A(n_302),
.Y(n_366)
);

AOI22x1_ASAP7_75t_SL g367 ( 
.A1(n_296),
.A2(n_286),
.B1(n_285),
.B2(n_281),
.Y(n_367)
);

INVx2_ASAP7_75t_L g368 ( 
.A(n_332),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_310),
.Y(n_369)
);

AND2x4_ASAP7_75t_L g370 ( 
.A(n_294),
.B(n_282),
.Y(n_370)
);

INVx2_ASAP7_75t_L g371 ( 
.A(n_295),
.Y(n_371)
);

AND2x2_ASAP7_75t_SL g372 ( 
.A(n_305),
.B(n_282),
.Y(n_372)
);

AND2x2_ASAP7_75t_L g373 ( 
.A(n_297),
.B(n_241),
.Y(n_373)
);

OA21x2_ASAP7_75t_L g374 ( 
.A1(n_304),
.A2(n_244),
.B(n_243),
.Y(n_374)
);

AND2x4_ASAP7_75t_L g375 ( 
.A(n_320),
.B(n_246),
.Y(n_375)
);

OAI22xp5_ASAP7_75t_SL g376 ( 
.A1(n_296),
.A2(n_280),
.B1(n_279),
.B2(n_276),
.Y(n_376)
);

AND2x4_ASAP7_75t_L g377 ( 
.A(n_323),
.B(n_249),
.Y(n_377)
);

OA21x2_ASAP7_75t_L g378 ( 
.A1(n_334),
.A2(n_251),
.B(n_250),
.Y(n_378)
);

OAI21x1_ASAP7_75t_L g379 ( 
.A1(n_322),
.A2(n_260),
.B(n_258),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_297),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_307),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_307),
.B(n_274),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_328),
.Y(n_383)
);

AND2x2_ASAP7_75t_L g384 ( 
.A(n_328),
.B(n_261),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_333),
.Y(n_385)
);

OA21x2_ASAP7_75t_L g386 ( 
.A1(n_333),
.A2(n_265),
.B(n_262),
.Y(n_386)
);

NOR2xp33_ASAP7_75t_L g387 ( 
.A(n_337),
.B(n_266),
.Y(n_387)
);

AND2x2_ASAP7_75t_L g388 ( 
.A(n_337),
.B(n_267),
.Y(n_388)
);

BUFx2_ASAP7_75t_L g389 ( 
.A(n_309),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_309),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_311),
.Y(n_391)
);

BUFx3_ASAP7_75t_L g392 ( 
.A(n_365),
.Y(n_392)
);

INVx5_ASAP7_75t_L g393 ( 
.A(n_339),
.Y(n_393)
);

INVx3_ASAP7_75t_L g394 ( 
.A(n_339),
.Y(n_394)
);

INVx2_ASAP7_75t_L g395 ( 
.A(n_341),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_366),
.Y(n_396)
);

INVx2_ASAP7_75t_L g397 ( 
.A(n_341),
.Y(n_397)
);

NOR2xp33_ASAP7_75t_L g398 ( 
.A(n_343),
.B(n_311),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_366),
.Y(n_399)
);

AND2x2_ASAP7_75t_L g400 ( 
.A(n_380),
.B(n_317),
.Y(n_400)
);

INVx3_ASAP7_75t_L g401 ( 
.A(n_339),
.Y(n_401)
);

NOR2xp33_ASAP7_75t_L g402 ( 
.A(n_348),
.B(n_325),
.Y(n_402)
);

INVx2_ASAP7_75t_L g403 ( 
.A(n_341),
.Y(n_403)
);

INVx2_ASAP7_75t_L g404 ( 
.A(n_339),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_366),
.Y(n_405)
);

INVx2_ASAP7_75t_L g406 ( 
.A(n_353),
.Y(n_406)
);

AND2x2_ASAP7_75t_L g407 ( 
.A(n_380),
.B(n_326),
.Y(n_407)
);

INVxp67_ASAP7_75t_SL g408 ( 
.A(n_365),
.Y(n_408)
);

INVx2_ASAP7_75t_L g409 ( 
.A(n_353),
.Y(n_409)
);

INVx3_ASAP7_75t_L g410 ( 
.A(n_339),
.Y(n_410)
);

INVx2_ASAP7_75t_L g411 ( 
.A(n_339),
.Y(n_411)
);

INVx2_ASAP7_75t_L g412 ( 
.A(n_342),
.Y(n_412)
);

AOI22xp5_ASAP7_75t_L g413 ( 
.A1(n_376),
.A2(n_273),
.B1(n_271),
.B2(n_269),
.Y(n_413)
);

INVx2_ASAP7_75t_L g414 ( 
.A(n_353),
.Y(n_414)
);

INVxp33_ASAP7_75t_SL g415 ( 
.A(n_376),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_350),
.Y(n_416)
);

AOI22xp5_ASAP7_75t_L g417 ( 
.A1(n_381),
.A2(n_318),
.B1(n_1),
.B2(n_2),
.Y(n_417)
);

AND2x2_ASAP7_75t_L g418 ( 
.A(n_370),
.B(n_373),
.Y(n_418)
);

INVx2_ASAP7_75t_L g419 ( 
.A(n_342),
.Y(n_419)
);

INVx2_ASAP7_75t_L g420 ( 
.A(n_342),
.Y(n_420)
);

INVx2_ASAP7_75t_L g421 ( 
.A(n_342),
.Y(n_421)
);

AND3x2_ASAP7_75t_L g422 ( 
.A(n_387),
.B(n_0),
.C(n_2),
.Y(n_422)
);

INVx2_ASAP7_75t_L g423 ( 
.A(n_353),
.Y(n_423)
);

INVx2_ASAP7_75t_L g424 ( 
.A(n_353),
.Y(n_424)
);

AND3x2_ASAP7_75t_L g425 ( 
.A(n_349),
.B(n_0),
.C(n_3),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_350),
.Y(n_426)
);

INVx2_ASAP7_75t_L g427 ( 
.A(n_353),
.Y(n_427)
);

AND2x2_ASAP7_75t_L g428 ( 
.A(n_370),
.B(n_373),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_350),
.Y(n_429)
);

NOR2xp33_ASAP7_75t_L g430 ( 
.A(n_371),
.B(n_318),
.Y(n_430)
);

INVx2_ASAP7_75t_L g431 ( 
.A(n_340),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_338),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_SL g433 ( 
.A(n_372),
.B(n_3),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_338),
.Y(n_434)
);

AND2x2_ASAP7_75t_L g435 ( 
.A(n_370),
.B(n_32),
.Y(n_435)
);

INVx2_ASAP7_75t_L g436 ( 
.A(n_340),
.Y(n_436)
);

INVxp67_ASAP7_75t_R g437 ( 
.A(n_379),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_344),
.Y(n_438)
);

INVx3_ASAP7_75t_L g439 ( 
.A(n_342),
.Y(n_439)
);

BUFx6f_ASAP7_75t_L g440 ( 
.A(n_342),
.Y(n_440)
);

AND3x2_ASAP7_75t_L g441 ( 
.A(n_384),
.B(n_4),
.C(n_6),
.Y(n_441)
);

INVx2_ASAP7_75t_SL g442 ( 
.A(n_347),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_SL g443 ( 
.A(n_372),
.B(n_6),
.Y(n_443)
);

INVx2_ASAP7_75t_L g444 ( 
.A(n_346),
.Y(n_444)
);

INVx5_ASAP7_75t_L g445 ( 
.A(n_365),
.Y(n_445)
);

INVx2_ASAP7_75t_L g446 ( 
.A(n_346),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_SL g447 ( 
.A(n_347),
.B(n_7),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_368),
.B(n_36),
.Y(n_448)
);

INVx2_ASAP7_75t_L g449 ( 
.A(n_351),
.Y(n_449)
);

INVx2_ASAP7_75t_L g450 ( 
.A(n_351),
.Y(n_450)
);

INVx2_ASAP7_75t_L g451 ( 
.A(n_344),
.Y(n_451)
);

AND3x2_ASAP7_75t_L g452 ( 
.A(n_384),
.B(n_7),
.C(n_8),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_355),
.Y(n_453)
);

AND2x2_ASAP7_75t_L g454 ( 
.A(n_370),
.B(n_37),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_L g455 ( 
.A(n_368),
.B(n_38),
.Y(n_455)
);

BUFx2_ASAP7_75t_L g456 ( 
.A(n_381),
.Y(n_456)
);

NOR2xp33_ASAP7_75t_L g457 ( 
.A(n_371),
.B(n_8),
.Y(n_457)
);

INVx6_ASAP7_75t_L g458 ( 
.A(n_365),
.Y(n_458)
);

OR2x6_ASAP7_75t_L g459 ( 
.A(n_379),
.B(n_374),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_368),
.B(n_39),
.Y(n_460)
);

INVx2_ASAP7_75t_L g461 ( 
.A(n_357),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_SL g462 ( 
.A(n_382),
.B(n_9),
.Y(n_462)
);

INVx2_ASAP7_75t_L g463 ( 
.A(n_352),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_355),
.Y(n_464)
);

INVx2_ASAP7_75t_L g465 ( 
.A(n_461),
.Y(n_465)
);

INVxp33_ASAP7_75t_SL g466 ( 
.A(n_398),
.Y(n_466)
);

CKINVDCx20_ASAP7_75t_R g467 ( 
.A(n_430),
.Y(n_467)
);

CKINVDCx5p33_ASAP7_75t_R g468 ( 
.A(n_402),
.Y(n_468)
);

BUFx5_ASAP7_75t_L g469 ( 
.A(n_392),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_453),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_453),
.Y(n_471)
);

AND2x4_ASAP7_75t_L g472 ( 
.A(n_464),
.B(n_360),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_464),
.Y(n_473)
);

CKINVDCx5p33_ASAP7_75t_R g474 ( 
.A(n_415),
.Y(n_474)
);

INVx4_ASAP7_75t_SL g475 ( 
.A(n_459),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_432),
.Y(n_476)
);

AND2x2_ASAP7_75t_L g477 ( 
.A(n_442),
.B(n_369),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_432),
.Y(n_478)
);

INVx2_ASAP7_75t_L g479 ( 
.A(n_461),
.Y(n_479)
);

XOR2x2_ASAP7_75t_L g480 ( 
.A(n_413),
.B(n_386),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_L g481 ( 
.A(n_418),
.B(n_428),
.Y(n_481)
);

CKINVDCx20_ASAP7_75t_R g482 ( 
.A(n_400),
.Y(n_482)
);

XNOR2xp5_ASAP7_75t_L g483 ( 
.A(n_400),
.B(n_389),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_L g484 ( 
.A(n_418),
.B(n_345),
.Y(n_484)
);

OAI21xp5_ASAP7_75t_L g485 ( 
.A1(n_463),
.A2(n_369),
.B(n_364),
.Y(n_485)
);

NOR2xp33_ASAP7_75t_L g486 ( 
.A(n_456),
.B(n_356),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_434),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_434),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_438),
.Y(n_489)
);

INVxp33_ASAP7_75t_L g490 ( 
.A(n_407),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_438),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_416),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_416),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_426),
.Y(n_494)
);

BUFx2_ASAP7_75t_L g495 ( 
.A(n_407),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_426),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_429),
.Y(n_497)
);

NOR2xp33_ASAP7_75t_L g498 ( 
.A(n_456),
.B(n_375),
.Y(n_498)
);

NOR2xp33_ASAP7_75t_L g499 ( 
.A(n_428),
.B(n_375),
.Y(n_499)
);

INVxp67_ASAP7_75t_SL g500 ( 
.A(n_440),
.Y(n_500)
);

INVxp33_ASAP7_75t_SL g501 ( 
.A(n_413),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_429),
.Y(n_502)
);

AND2x2_ASAP7_75t_L g503 ( 
.A(n_457),
.B(n_388),
.Y(n_503)
);

XOR2xp5_ASAP7_75t_L g504 ( 
.A(n_433),
.B(n_389),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_444),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_444),
.Y(n_506)
);

OR2x6_ASAP7_75t_L g507 ( 
.A(n_443),
.B(n_383),
.Y(n_507)
);

AND2x2_ASAP7_75t_L g508 ( 
.A(n_447),
.B(n_360),
.Y(n_508)
);

CKINVDCx20_ASAP7_75t_R g509 ( 
.A(n_459),
.Y(n_509)
);

INVxp33_ASAP7_75t_SL g510 ( 
.A(n_437),
.Y(n_510)
);

CKINVDCx5p33_ASAP7_75t_R g511 ( 
.A(n_459),
.Y(n_511)
);

BUFx2_ASAP7_75t_L g512 ( 
.A(n_441),
.Y(n_512)
);

INVxp33_ASAP7_75t_L g513 ( 
.A(n_462),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_446),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_446),
.Y(n_515)
);

OAI21xp5_ASAP7_75t_L g516 ( 
.A1(n_463),
.A2(n_364),
.B(n_352),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_449),
.Y(n_517)
);

INVx2_ASAP7_75t_L g518 ( 
.A(n_449),
.Y(n_518)
);

CKINVDCx14_ASAP7_75t_R g519 ( 
.A(n_459),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_L g520 ( 
.A(n_435),
.B(n_345),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_L g521 ( 
.A(n_435),
.B(n_363),
.Y(n_521)
);

NOR2xp33_ASAP7_75t_L g522 ( 
.A(n_454),
.B(n_375),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_450),
.Y(n_523)
);

NOR2xp33_ASAP7_75t_L g524 ( 
.A(n_454),
.B(n_375),
.Y(n_524)
);

NOR2xp33_ASAP7_75t_L g525 ( 
.A(n_448),
.B(n_377),
.Y(n_525)
);

INVx2_ASAP7_75t_L g526 ( 
.A(n_450),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_451),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_451),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_396),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_396),
.Y(n_530)
);

CKINVDCx5p33_ASAP7_75t_R g531 ( 
.A(n_459),
.Y(n_531)
);

XOR2xp5_ASAP7_75t_L g532 ( 
.A(n_417),
.B(n_367),
.Y(n_532)
);

AND2x4_ASAP7_75t_L g533 ( 
.A(n_392),
.B(n_363),
.Y(n_533)
);

OR2x6_ASAP7_75t_L g534 ( 
.A(n_455),
.B(n_383),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_399),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_SL g536 ( 
.A(n_460),
.B(n_377),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_399),
.Y(n_537)
);

XNOR2xp5_ASAP7_75t_L g538 ( 
.A(n_417),
.B(n_367),
.Y(n_538)
);

AND2x2_ASAP7_75t_L g539 ( 
.A(n_405),
.B(n_377),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_431),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_431),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_436),
.Y(n_542)
);

NOR2xp33_ASAP7_75t_L g543 ( 
.A(n_392),
.B(n_377),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_436),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_395),
.Y(n_545)
);

NOR2xp33_ASAP7_75t_L g546 ( 
.A(n_408),
.B(n_386),
.Y(n_546)
);

NOR2xp33_ASAP7_75t_L g547 ( 
.A(n_466),
.B(n_386),
.Y(n_547)
);

OAI22xp5_ASAP7_75t_L g548 ( 
.A1(n_522),
.A2(n_437),
.B1(n_463),
.B2(n_386),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_L g549 ( 
.A(n_481),
.B(n_345),
.Y(n_549)
);

INVx2_ASAP7_75t_SL g550 ( 
.A(n_495),
.Y(n_550)
);

NOR2xp33_ASAP7_75t_L g551 ( 
.A(n_468),
.B(n_385),
.Y(n_551)
);

AOI22xp33_ASAP7_75t_L g552 ( 
.A1(n_501),
.A2(n_378),
.B1(n_374),
.B2(n_345),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_505),
.Y(n_553)
);

INVx2_ASAP7_75t_SL g554 ( 
.A(n_477),
.Y(n_554)
);

INVx2_ASAP7_75t_L g555 ( 
.A(n_465),
.Y(n_555)
);

AND2x4_ASAP7_75t_L g556 ( 
.A(n_533),
.B(n_452),
.Y(n_556)
);

AND2x2_ASAP7_75t_L g557 ( 
.A(n_486),
.B(n_385),
.Y(n_557)
);

INVx2_ASAP7_75t_L g558 ( 
.A(n_479),
.Y(n_558)
);

NOR2xp33_ASAP7_75t_L g559 ( 
.A(n_490),
.B(n_374),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_SL g560 ( 
.A(n_498),
.B(n_365),
.Y(n_560)
);

AND2x2_ASAP7_75t_L g561 ( 
.A(n_503),
.B(n_390),
.Y(n_561)
);

AOI22xp5_ASAP7_75t_L g562 ( 
.A1(n_499),
.A2(n_374),
.B1(n_378),
.B2(n_391),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_L g563 ( 
.A(n_481),
.B(n_378),
.Y(n_563)
);

AND2x4_ASAP7_75t_L g564 ( 
.A(n_533),
.B(n_422),
.Y(n_564)
);

INVx2_ASAP7_75t_SL g565 ( 
.A(n_482),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_SL g566 ( 
.A(n_472),
.B(n_365),
.Y(n_566)
);

OR2x2_ASAP7_75t_L g567 ( 
.A(n_483),
.B(n_358),
.Y(n_567)
);

AOI22xp33_ASAP7_75t_SL g568 ( 
.A1(n_467),
.A2(n_425),
.B1(n_358),
.B2(n_359),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_SL g569 ( 
.A(n_472),
.B(n_357),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_L g570 ( 
.A(n_484),
.B(n_394),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_L g571 ( 
.A(n_484),
.B(n_394),
.Y(n_571)
);

BUFx3_ASAP7_75t_L g572 ( 
.A(n_512),
.Y(n_572)
);

AOI22xp33_ASAP7_75t_L g573 ( 
.A1(n_480),
.A2(n_354),
.B1(n_403),
.B2(n_395),
.Y(n_573)
);

OR2x2_ASAP7_75t_L g574 ( 
.A(n_507),
.B(n_359),
.Y(n_574)
);

NOR2x1p5_ASAP7_75t_L g575 ( 
.A(n_474),
.B(n_362),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_L g576 ( 
.A(n_521),
.B(n_394),
.Y(n_576)
);

NOR2xp33_ASAP7_75t_L g577 ( 
.A(n_513),
.B(n_362),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_L g578 ( 
.A(n_539),
.B(n_394),
.Y(n_578)
);

AOI22xp33_ASAP7_75t_L g579 ( 
.A1(n_507),
.A2(n_354),
.B1(n_397),
.B2(n_403),
.Y(n_579)
);

BUFx3_ASAP7_75t_L g580 ( 
.A(n_534),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_506),
.Y(n_581)
);

AO22x1_ASAP7_75t_L g582 ( 
.A1(n_524),
.A2(n_361),
.B1(n_397),
.B2(n_412),
.Y(n_582)
);

O2A1O1Ixp33_ASAP7_75t_L g583 ( 
.A1(n_520),
.A2(n_354),
.B(n_412),
.C(n_411),
.Y(n_583)
);

INVx2_ASAP7_75t_L g584 ( 
.A(n_518),
.Y(n_584)
);

NAND2xp5_ASAP7_75t_L g585 ( 
.A(n_470),
.B(n_471),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_L g586 ( 
.A(n_473),
.B(n_476),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_SL g587 ( 
.A(n_508),
.B(n_361),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_SL g588 ( 
.A(n_510),
.B(n_440),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_L g589 ( 
.A(n_478),
.B(n_487),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_SL g590 ( 
.A(n_488),
.B(n_440),
.Y(n_590)
);

INVx3_ASAP7_75t_L g591 ( 
.A(n_526),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_L g592 ( 
.A(n_489),
.B(n_401),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_L g593 ( 
.A(n_491),
.B(n_401),
.Y(n_593)
);

AND2x6_ASAP7_75t_SL g594 ( 
.A(n_507),
.B(n_9),
.Y(n_594)
);

INVx5_ASAP7_75t_L g595 ( 
.A(n_534),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_SL g596 ( 
.A(n_525),
.B(n_440),
.Y(n_596)
);

AND2x2_ASAP7_75t_L g597 ( 
.A(n_534),
.B(n_354),
.Y(n_597)
);

AND2x2_ASAP7_75t_L g598 ( 
.A(n_504),
.B(n_406),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_514),
.Y(n_599)
);

AND2x2_ASAP7_75t_L g600 ( 
.A(n_543),
.B(n_406),
.Y(n_600)
);

NAND2x1p5_ASAP7_75t_L g601 ( 
.A(n_492),
.B(n_445),
.Y(n_601)
);

NOR2xp33_ASAP7_75t_L g602 ( 
.A(n_493),
.B(n_458),
.Y(n_602)
);

AOI22xp33_ASAP7_75t_L g603 ( 
.A1(n_520),
.A2(n_546),
.B1(n_494),
.B2(n_497),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_L g604 ( 
.A(n_496),
.B(n_401),
.Y(n_604)
);

INVx2_ASAP7_75t_L g605 ( 
.A(n_515),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_SL g606 ( 
.A(n_502),
.B(n_517),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_L g607 ( 
.A(n_523),
.B(n_401),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_527),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_528),
.Y(n_609)
);

AOI22xp5_ASAP7_75t_L g610 ( 
.A1(n_509),
.A2(n_458),
.B1(n_409),
.B2(n_427),
.Y(n_610)
);

INVx4_ASAP7_75t_L g611 ( 
.A(n_475),
.Y(n_611)
);

BUFx6f_ASAP7_75t_L g612 ( 
.A(n_529),
.Y(n_612)
);

NOR2xp33_ASAP7_75t_L g613 ( 
.A(n_530),
.B(n_458),
.Y(n_613)
);

INVx2_ASAP7_75t_SL g614 ( 
.A(n_565),
.Y(n_614)
);

BUFx6f_ASAP7_75t_L g615 ( 
.A(n_611),
.Y(n_615)
);

INVxp67_ASAP7_75t_SL g616 ( 
.A(n_612),
.Y(n_616)
);

BUFx6f_ASAP7_75t_L g617 ( 
.A(n_611),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_592),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_L g619 ( 
.A(n_554),
.B(n_535),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_553),
.Y(n_620)
);

HB1xp67_ASAP7_75t_L g621 ( 
.A(n_550),
.Y(n_621)
);

INVx4_ASAP7_75t_L g622 ( 
.A(n_612),
.Y(n_622)
);

BUFx6f_ASAP7_75t_L g623 ( 
.A(n_612),
.Y(n_623)
);

BUFx6f_ASAP7_75t_L g624 ( 
.A(n_580),
.Y(n_624)
);

NAND2xp33_ASAP7_75t_SL g625 ( 
.A(n_575),
.B(n_511),
.Y(n_625)
);

INVx4_ASAP7_75t_L g626 ( 
.A(n_595),
.Y(n_626)
);

AND2x4_ASAP7_75t_L g627 ( 
.A(n_556),
.B(n_475),
.Y(n_627)
);

AND2x4_ASAP7_75t_L g628 ( 
.A(n_556),
.B(n_475),
.Y(n_628)
);

NOR2xp33_ASAP7_75t_R g629 ( 
.A(n_547),
.B(n_519),
.Y(n_629)
);

BUFx4f_ASAP7_75t_L g630 ( 
.A(n_564),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_L g631 ( 
.A(n_549),
.B(n_537),
.Y(n_631)
);

INVx6_ASAP7_75t_L g632 ( 
.A(n_572),
.Y(n_632)
);

BUFx3_ASAP7_75t_L g633 ( 
.A(n_598),
.Y(n_633)
);

INVx4_ASAP7_75t_L g634 ( 
.A(n_595),
.Y(n_634)
);

AOI22xp5_ASAP7_75t_L g635 ( 
.A1(n_547),
.A2(n_536),
.B1(n_531),
.B2(n_538),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_581),
.Y(n_636)
);

OR2x2_ASAP7_75t_L g637 ( 
.A(n_567),
.B(n_485),
.Y(n_637)
);

AND2x4_ASAP7_75t_L g638 ( 
.A(n_595),
.B(n_500),
.Y(n_638)
);

INVx5_ASAP7_75t_L g639 ( 
.A(n_595),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_599),
.Y(n_640)
);

INVx3_ASAP7_75t_L g641 ( 
.A(n_601),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_608),
.Y(n_642)
);

NOR2xp33_ASAP7_75t_L g643 ( 
.A(n_551),
.B(n_532),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_609),
.Y(n_644)
);

INVx1_ASAP7_75t_SL g645 ( 
.A(n_557),
.Y(n_645)
);

NOR2xp33_ASAP7_75t_L g646 ( 
.A(n_551),
.B(n_561),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_L g647 ( 
.A(n_585),
.B(n_469),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_586),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_589),
.Y(n_649)
);

CKINVDCx16_ASAP7_75t_R g650 ( 
.A(n_564),
.Y(n_650)
);

BUFx6f_ASAP7_75t_L g651 ( 
.A(n_574),
.Y(n_651)
);

BUFx2_ASAP7_75t_SL g652 ( 
.A(n_584),
.Y(n_652)
);

INVx4_ASAP7_75t_L g653 ( 
.A(n_591),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_593),
.Y(n_654)
);

INVx2_ASAP7_75t_L g655 ( 
.A(n_605),
.Y(n_655)
);

OAI21xp33_ASAP7_75t_SL g656 ( 
.A1(n_579),
.A2(n_485),
.B(n_516),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_555),
.Y(n_657)
);

INVx3_ASAP7_75t_L g658 ( 
.A(n_601),
.Y(n_658)
);

CKINVDCx5p33_ASAP7_75t_R g659 ( 
.A(n_594),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_L g660 ( 
.A(n_577),
.B(n_469),
.Y(n_660)
);

NAND2x1p5_ASAP7_75t_L g661 ( 
.A(n_591),
.B(n_540),
.Y(n_661)
);

BUFx3_ASAP7_75t_L g662 ( 
.A(n_577),
.Y(n_662)
);

INVx3_ASAP7_75t_L g663 ( 
.A(n_558),
.Y(n_663)
);

HB1xp67_ASAP7_75t_L g664 ( 
.A(n_569),
.Y(n_664)
);

NOR2xp33_ASAP7_75t_L g665 ( 
.A(n_559),
.B(n_541),
.Y(n_665)
);

AND2x4_ASAP7_75t_L g666 ( 
.A(n_566),
.B(n_542),
.Y(n_666)
);

NAND2x1p5_ASAP7_75t_L g667 ( 
.A(n_588),
.B(n_606),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_604),
.Y(n_668)
);

NOR2xp33_ASAP7_75t_L g669 ( 
.A(n_559),
.B(n_544),
.Y(n_669)
);

INVx2_ASAP7_75t_L g670 ( 
.A(n_607),
.Y(n_670)
);

BUFx3_ASAP7_75t_L g671 ( 
.A(n_597),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_570),
.Y(n_672)
);

INVx2_ASAP7_75t_L g673 ( 
.A(n_576),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_571),
.Y(n_674)
);

BUFx4f_ASAP7_75t_L g675 ( 
.A(n_600),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_L g676 ( 
.A(n_603),
.B(n_573),
.Y(n_676)
);

INVx2_ASAP7_75t_SL g677 ( 
.A(n_632),
.Y(n_677)
);

OR2x6_ASAP7_75t_L g678 ( 
.A(n_632),
.B(n_587),
.Y(n_678)
);

INVx2_ASAP7_75t_L g679 ( 
.A(n_620),
.Y(n_679)
);

AOI21x1_ASAP7_75t_L g680 ( 
.A1(n_660),
.A2(n_582),
.B(n_596),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_L g681 ( 
.A(n_648),
.B(n_603),
.Y(n_681)
);

INVx2_ASAP7_75t_L g682 ( 
.A(n_636),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_L g683 ( 
.A(n_649),
.B(n_573),
.Y(n_683)
);

OAI21x1_ASAP7_75t_L g684 ( 
.A1(n_647),
.A2(n_583),
.B(n_516),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_640),
.Y(n_685)
);

BUFx6f_ASAP7_75t_L g686 ( 
.A(n_615),
.Y(n_686)
);

OAI21xp5_ASAP7_75t_L g687 ( 
.A1(n_665),
.A2(n_563),
.B(n_548),
.Y(n_687)
);

NAND2x1p5_ASAP7_75t_L g688 ( 
.A(n_639),
.B(n_590),
.Y(n_688)
);

BUFx6f_ASAP7_75t_L g689 ( 
.A(n_615),
.Y(n_689)
);

AND2x4_ASAP7_75t_L g690 ( 
.A(n_627),
.B(n_610),
.Y(n_690)
);

AOI21xp5_ASAP7_75t_L g691 ( 
.A1(n_631),
.A2(n_560),
.B(n_578),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_SL g692 ( 
.A(n_646),
.B(n_568),
.Y(n_692)
);

OAI21x1_ASAP7_75t_L g693 ( 
.A1(n_618),
.A2(n_583),
.B(n_579),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_L g694 ( 
.A(n_645),
.B(n_568),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_L g695 ( 
.A(n_662),
.B(n_552),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_SL g696 ( 
.A(n_675),
.B(n_562),
.Y(n_696)
);

AOI21xp5_ASAP7_75t_L g697 ( 
.A1(n_656),
.A2(n_613),
.B(n_552),
.Y(n_697)
);

OAI21x1_ASAP7_75t_L g698 ( 
.A1(n_618),
.A2(n_545),
.B(n_602),
.Y(n_698)
);

AOI21xp5_ASAP7_75t_L g699 ( 
.A1(n_669),
.A2(n_602),
.B(n_469),
.Y(n_699)
);

OAI21xp5_ASAP7_75t_L g700 ( 
.A1(n_672),
.A2(n_414),
.B(n_409),
.Y(n_700)
);

AOI21xp5_ASAP7_75t_L g701 ( 
.A1(n_672),
.A2(n_469),
.B(n_445),
.Y(n_701)
);

OAI21x1_ASAP7_75t_L g702 ( 
.A1(n_654),
.A2(n_411),
.B(n_404),
.Y(n_702)
);

AOI22xp5_ASAP7_75t_L g703 ( 
.A1(n_635),
.A2(n_458),
.B1(n_414),
.B2(n_423),
.Y(n_703)
);

OAI21x1_ASAP7_75t_L g704 ( 
.A1(n_654),
.A2(n_668),
.B(n_658),
.Y(n_704)
);

OAI21x1_ASAP7_75t_L g705 ( 
.A1(n_668),
.A2(n_411),
.B(n_404),
.Y(n_705)
);

INVx3_ASAP7_75t_L g706 ( 
.A(n_615),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_642),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_L g708 ( 
.A(n_674),
.B(n_469),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_L g709 ( 
.A(n_674),
.B(n_423),
.Y(n_709)
);

OR2x6_ASAP7_75t_L g710 ( 
.A(n_627),
.B(n_424),
.Y(n_710)
);

INVx2_ASAP7_75t_L g711 ( 
.A(n_644),
.Y(n_711)
);

OR2x2_ASAP7_75t_L g712 ( 
.A(n_637),
.B(n_424),
.Y(n_712)
);

AOI21xp5_ASAP7_75t_L g713 ( 
.A1(n_675),
.A2(n_445),
.B(n_440),
.Y(n_713)
);

AOI21xp5_ASAP7_75t_SL g714 ( 
.A1(n_676),
.A2(n_427),
.B(n_412),
.Y(n_714)
);

INVx2_ASAP7_75t_SL g715 ( 
.A(n_624),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_673),
.Y(n_716)
);

BUFx2_ASAP7_75t_L g717 ( 
.A(n_633),
.Y(n_717)
);

OAI21x1_ASAP7_75t_L g718 ( 
.A1(n_641),
.A2(n_419),
.B(n_404),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_L g719 ( 
.A(n_664),
.B(n_419),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_L g720 ( 
.A(n_671),
.B(n_419),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_670),
.Y(n_721)
);

INVx1_ASAP7_75t_SL g722 ( 
.A(n_621),
.Y(n_722)
);

AOI21xp5_ASAP7_75t_L g723 ( 
.A1(n_616),
.A2(n_445),
.B(n_393),
.Y(n_723)
);

AOI21xp5_ASAP7_75t_L g724 ( 
.A1(n_638),
.A2(n_445),
.B(n_393),
.Y(n_724)
);

OAI21x1_ASAP7_75t_L g725 ( 
.A1(n_641),
.A2(n_421),
.B(n_420),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_L g726 ( 
.A(n_651),
.B(n_420),
.Y(n_726)
);

BUFx6f_ASAP7_75t_L g727 ( 
.A(n_617),
.Y(n_727)
);

OAI21x1_ASAP7_75t_L g728 ( 
.A1(n_658),
.A2(n_421),
.B(n_420),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_L g729 ( 
.A(n_651),
.B(n_421),
.Y(n_729)
);

INVx2_ASAP7_75t_L g730 ( 
.A(n_655),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_L g731 ( 
.A(n_651),
.B(n_410),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_SL g732 ( 
.A(n_614),
.B(n_410),
.Y(n_732)
);

AOI21x1_ASAP7_75t_L g733 ( 
.A1(n_666),
.A2(n_445),
.B(n_439),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_L g734 ( 
.A(n_619),
.B(n_410),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_L g735 ( 
.A(n_663),
.B(n_410),
.Y(n_735)
);

AO31x2_ASAP7_75t_L g736 ( 
.A1(n_653),
.A2(n_439),
.A3(n_11),
.B(n_12),
.Y(n_736)
);

INVx2_ASAP7_75t_SL g737 ( 
.A(n_677),
.Y(n_737)
);

OAI21x1_ASAP7_75t_L g738 ( 
.A1(n_702),
.A2(n_667),
.B(n_661),
.Y(n_738)
);

A2O1A1Ixp33_ASAP7_75t_L g739 ( 
.A1(n_697),
.A2(n_643),
.B(n_625),
.C(n_657),
.Y(n_739)
);

CKINVDCx20_ASAP7_75t_R g740 ( 
.A(n_717),
.Y(n_740)
);

AOI21xp5_ASAP7_75t_L g741 ( 
.A1(n_687),
.A2(n_638),
.B(n_639),
.Y(n_741)
);

AOI221x1_ASAP7_75t_L g742 ( 
.A1(n_714),
.A2(n_666),
.B1(n_652),
.B2(n_634),
.C(n_626),
.Y(n_742)
);

NAND2x1_ASAP7_75t_L g743 ( 
.A(n_721),
.B(n_622),
.Y(n_743)
);

A2O1A1Ixp33_ASAP7_75t_L g744 ( 
.A1(n_692),
.A2(n_630),
.B(n_663),
.C(n_639),
.Y(n_744)
);

OA21x2_ASAP7_75t_L g745 ( 
.A1(n_684),
.A2(n_628),
.B(n_629),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_685),
.Y(n_746)
);

A2O1A1Ixp33_ASAP7_75t_L g747 ( 
.A1(n_696),
.A2(n_630),
.B(n_623),
.C(n_628),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_L g748 ( 
.A(n_716),
.B(n_650),
.Y(n_748)
);

OAI22xp5_ASAP7_75t_L g749 ( 
.A1(n_694),
.A2(n_623),
.B1(n_624),
.B2(n_659),
.Y(n_749)
);

NOR2xp67_ASAP7_75t_L g750 ( 
.A(n_730),
.B(n_624),
.Y(n_750)
);

OA21x2_ASAP7_75t_L g751 ( 
.A1(n_693),
.A2(n_623),
.B(n_439),
.Y(n_751)
);

BUFx10_ASAP7_75t_L g752 ( 
.A(n_715),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_L g753 ( 
.A(n_716),
.B(n_617),
.Y(n_753)
);

INVx3_ASAP7_75t_SL g754 ( 
.A(n_678),
.Y(n_754)
);

AOI21xp5_ASAP7_75t_L g755 ( 
.A1(n_699),
.A2(n_617),
.B(n_439),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_685),
.Y(n_756)
);

AO31x2_ASAP7_75t_L g757 ( 
.A1(n_701),
.A2(n_115),
.A3(n_217),
.B(n_216),
.Y(n_757)
);

AO31x2_ASAP7_75t_L g758 ( 
.A1(n_691),
.A2(n_681),
.A3(n_683),
.B(n_708),
.Y(n_758)
);

BUFx12f_ASAP7_75t_L g759 ( 
.A(n_686),
.Y(n_759)
);

AO31x2_ASAP7_75t_L g760 ( 
.A1(n_695),
.A2(n_114),
.A3(n_214),
.B(n_213),
.Y(n_760)
);

AO31x2_ASAP7_75t_L g761 ( 
.A1(n_709),
.A2(n_112),
.A3(n_212),
.B(n_211),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_707),
.Y(n_762)
);

O2A1O1Ixp33_ASAP7_75t_SL g763 ( 
.A1(n_732),
.A2(n_10),
.B(n_11),
.C(n_12),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_L g764 ( 
.A(n_721),
.B(n_722),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_L g765 ( 
.A(n_722),
.B(n_10),
.Y(n_765)
);

NOR2xp33_ASAP7_75t_L g766 ( 
.A(n_690),
.B(n_42),
.Y(n_766)
);

A2O1A1Ixp33_ASAP7_75t_L g767 ( 
.A1(n_690),
.A2(n_13),
.B(n_14),
.C(n_15),
.Y(n_767)
);

AOI21xp5_ASAP7_75t_L g768 ( 
.A1(n_700),
.A2(n_393),
.B(n_45),
.Y(n_768)
);

AOI21xp5_ASAP7_75t_L g769 ( 
.A1(n_704),
.A2(n_713),
.B(n_698),
.Y(n_769)
);

AO31x2_ASAP7_75t_L g770 ( 
.A1(n_724),
.A2(n_120),
.A3(n_209),
.B(n_206),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_679),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_682),
.Y(n_772)
);

A2O1A1Ixp33_ASAP7_75t_L g773 ( 
.A1(n_711),
.A2(n_14),
.B(n_15),
.C(n_16),
.Y(n_773)
);

OAI21x1_ASAP7_75t_L g774 ( 
.A1(n_705),
.A2(n_725),
.B(n_718),
.Y(n_774)
);

NOR2xp33_ASAP7_75t_L g775 ( 
.A(n_731),
.B(n_44),
.Y(n_775)
);

AOI221x1_ASAP7_75t_L g776 ( 
.A1(n_720),
.A2(n_16),
.B1(n_17),
.B2(n_18),
.C(n_19),
.Y(n_776)
);

AOI21xp5_ASAP7_75t_SL g777 ( 
.A1(n_712),
.A2(n_122),
.B(n_205),
.Y(n_777)
);

AO31x2_ASAP7_75t_L g778 ( 
.A1(n_723),
.A2(n_121),
.A3(n_204),
.B(n_203),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_L g779 ( 
.A(n_726),
.B(n_18),
.Y(n_779)
);

INVx5_ASAP7_75t_L g780 ( 
.A(n_686),
.Y(n_780)
);

AOI21xp5_ASAP7_75t_L g781 ( 
.A1(n_734),
.A2(n_393),
.B(n_118),
.Y(n_781)
);

AOI21xp5_ASAP7_75t_L g782 ( 
.A1(n_703),
.A2(n_393),
.B(n_113),
.Y(n_782)
);

AOI22xp5_ASAP7_75t_L g783 ( 
.A1(n_678),
.A2(n_393),
.B1(n_20),
.B2(n_21),
.Y(n_783)
);

O2A1O1Ixp33_ASAP7_75t_L g784 ( 
.A1(n_729),
.A2(n_19),
.B(n_20),
.C(n_21),
.Y(n_784)
);

AND2x2_ASAP7_75t_L g785 ( 
.A(n_710),
.B(n_22),
.Y(n_785)
);

BUFx12f_ASAP7_75t_L g786 ( 
.A(n_686),
.Y(n_786)
);

BUFx10_ASAP7_75t_L g787 ( 
.A(n_689),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_L g788 ( 
.A(n_719),
.B(n_23),
.Y(n_788)
);

OA21x2_ASAP7_75t_L g789 ( 
.A1(n_680),
.A2(n_127),
.B(n_200),
.Y(n_789)
);

OAI21xp5_ASAP7_75t_L g790 ( 
.A1(n_703),
.A2(n_735),
.B(n_733),
.Y(n_790)
);

INVx2_ASAP7_75t_L g791 ( 
.A(n_706),
.Y(n_791)
);

OA21x2_ASAP7_75t_L g792 ( 
.A1(n_728),
.A2(n_126),
.B(n_199),
.Y(n_792)
);

AOI21xp5_ASAP7_75t_L g793 ( 
.A1(n_688),
.A2(n_123),
.B(n_198),
.Y(n_793)
);

INVx2_ASAP7_75t_SL g794 ( 
.A(n_689),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_L g795 ( 
.A(n_706),
.B(n_24),
.Y(n_795)
);

AO31x2_ASAP7_75t_L g796 ( 
.A1(n_736),
.A2(n_109),
.A3(n_197),
.B(n_195),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_736),
.Y(n_797)
);

OAI22xp5_ASAP7_75t_L g798 ( 
.A1(n_710),
.A2(n_24),
.B1(n_25),
.B2(n_26),
.Y(n_798)
);

AOI21xp5_ASAP7_75t_L g799 ( 
.A1(n_689),
.A2(n_108),
.B(n_193),
.Y(n_799)
);

OAI21xp5_ASAP7_75t_L g800 ( 
.A1(n_736),
.A2(n_25),
.B(n_26),
.Y(n_800)
);

AOI21xp5_ASAP7_75t_L g801 ( 
.A1(n_727),
.A2(n_128),
.B(n_192),
.Y(n_801)
);

CKINVDCx16_ASAP7_75t_R g802 ( 
.A(n_727),
.Y(n_802)
);

AND2x2_ASAP7_75t_L g803 ( 
.A(n_748),
.B(n_727),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_746),
.Y(n_804)
);

INVx2_ASAP7_75t_L g805 ( 
.A(n_771),
.Y(n_805)
);

AOI22xp33_ASAP7_75t_L g806 ( 
.A1(n_766),
.A2(n_27),
.B1(n_28),
.B2(n_29),
.Y(n_806)
);

BUFx10_ASAP7_75t_L g807 ( 
.A(n_737),
.Y(n_807)
);

BUFx4f_ASAP7_75t_SL g808 ( 
.A(n_759),
.Y(n_808)
);

INVx6_ASAP7_75t_L g809 ( 
.A(n_780),
.Y(n_809)
);

OAI22xp5_ASAP7_75t_L g810 ( 
.A1(n_767),
.A2(n_27),
.B1(n_28),
.B2(n_29),
.Y(n_810)
);

CKINVDCx11_ASAP7_75t_R g811 ( 
.A(n_740),
.Y(n_811)
);

OAI21xp33_ASAP7_75t_L g812 ( 
.A1(n_739),
.A2(n_30),
.B(n_31),
.Y(n_812)
);

AOI22xp33_ASAP7_75t_SL g813 ( 
.A1(n_800),
.A2(n_798),
.B1(n_776),
.B2(n_765),
.Y(n_813)
);

AOI22xp33_ASAP7_75t_L g814 ( 
.A1(n_783),
.A2(n_30),
.B1(n_31),
.B2(n_46),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_756),
.Y(n_815)
);

AOI22xp5_ASAP7_75t_L g816 ( 
.A1(n_749),
.A2(n_47),
.B1(n_48),
.B2(n_51),
.Y(n_816)
);

BUFx12f_ASAP7_75t_L g817 ( 
.A(n_786),
.Y(n_817)
);

AOI22xp33_ASAP7_75t_L g818 ( 
.A1(n_754),
.A2(n_53),
.B1(n_56),
.B2(n_57),
.Y(n_818)
);

BUFx2_ASAP7_75t_SL g819 ( 
.A(n_750),
.Y(n_819)
);

BUFx3_ASAP7_75t_L g820 ( 
.A(n_752),
.Y(n_820)
);

CKINVDCx11_ASAP7_75t_R g821 ( 
.A(n_802),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_762),
.Y(n_822)
);

AOI22xp5_ASAP7_75t_L g823 ( 
.A1(n_775),
.A2(n_58),
.B1(n_59),
.B2(n_60),
.Y(n_823)
);

INVx2_ASAP7_75t_L g824 ( 
.A(n_772),
.Y(n_824)
);

AOI22xp33_ASAP7_75t_SL g825 ( 
.A1(n_785),
.A2(n_61),
.B1(n_62),
.B2(n_64),
.Y(n_825)
);

INVx2_ASAP7_75t_L g826 ( 
.A(n_791),
.Y(n_826)
);

AOI22xp33_ASAP7_75t_L g827 ( 
.A1(n_788),
.A2(n_65),
.B1(n_67),
.B2(n_68),
.Y(n_827)
);

INVx6_ASAP7_75t_L g828 ( 
.A(n_780),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_764),
.Y(n_829)
);

OAI22xp5_ASAP7_75t_L g830 ( 
.A1(n_773),
.A2(n_69),
.B1(n_70),
.B2(n_71),
.Y(n_830)
);

AOI22xp33_ASAP7_75t_L g831 ( 
.A1(n_779),
.A2(n_795),
.B1(n_782),
.B2(n_741),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_797),
.Y(n_832)
);

BUFx10_ASAP7_75t_L g833 ( 
.A(n_794),
.Y(n_833)
);

BUFx3_ASAP7_75t_L g834 ( 
.A(n_787),
.Y(n_834)
);

AO22x1_ASAP7_75t_L g835 ( 
.A1(n_780),
.A2(n_72),
.B1(n_73),
.B2(n_77),
.Y(n_835)
);

BUFx6f_ASAP7_75t_L g836 ( 
.A(n_753),
.Y(n_836)
);

AOI22xp33_ASAP7_75t_L g837 ( 
.A1(n_793),
.A2(n_81),
.B1(n_82),
.B2(n_83),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_758),
.Y(n_838)
);

BUFx2_ASAP7_75t_SL g839 ( 
.A(n_745),
.Y(n_839)
);

CKINVDCx6p67_ASAP7_75t_R g840 ( 
.A(n_777),
.Y(n_840)
);

INVx6_ASAP7_75t_L g841 ( 
.A(n_747),
.Y(n_841)
);

INVx2_ASAP7_75t_L g842 ( 
.A(n_743),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_796),
.Y(n_843)
);

OAI22xp33_ASAP7_75t_L g844 ( 
.A1(n_742),
.A2(n_86),
.B1(n_87),
.B2(n_89),
.Y(n_844)
);

AOI22xp33_ASAP7_75t_L g845 ( 
.A1(n_799),
.A2(n_90),
.B1(n_91),
.B2(n_92),
.Y(n_845)
);

AOI22xp33_ASAP7_75t_L g846 ( 
.A1(n_801),
.A2(n_94),
.B1(n_95),
.B2(n_97),
.Y(n_846)
);

AOI22xp33_ASAP7_75t_L g847 ( 
.A1(n_768),
.A2(n_100),
.B1(n_101),
.B2(n_102),
.Y(n_847)
);

INVx1_ASAP7_75t_L g848 ( 
.A(n_796),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_751),
.Y(n_849)
);

OAI21xp5_ASAP7_75t_SL g850 ( 
.A1(n_784),
.A2(n_103),
.B(n_104),
.Y(n_850)
);

CKINVDCx5p33_ASAP7_75t_R g851 ( 
.A(n_781),
.Y(n_851)
);

OAI21xp5_ASAP7_75t_SL g852 ( 
.A1(n_744),
.A2(n_105),
.B(n_107),
.Y(n_852)
);

INVx1_ASAP7_75t_L g853 ( 
.A(n_745),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_760),
.Y(n_854)
);

BUFx6f_ASAP7_75t_L g855 ( 
.A(n_738),
.Y(n_855)
);

CKINVDCx11_ASAP7_75t_R g856 ( 
.A(n_763),
.Y(n_856)
);

AOI22xp33_ASAP7_75t_SL g857 ( 
.A1(n_789),
.A2(n_130),
.B1(n_131),
.B2(n_133),
.Y(n_857)
);

AOI22xp33_ASAP7_75t_L g858 ( 
.A1(n_790),
.A2(n_135),
.B1(n_137),
.B2(n_138),
.Y(n_858)
);

INVx2_ASAP7_75t_L g859 ( 
.A(n_761),
.Y(n_859)
);

AOI22xp33_ASAP7_75t_L g860 ( 
.A1(n_755),
.A2(n_142),
.B1(n_145),
.B2(n_147),
.Y(n_860)
);

AOI22xp33_ASAP7_75t_L g861 ( 
.A1(n_792),
.A2(n_148),
.B1(n_149),
.B2(n_150),
.Y(n_861)
);

INVx1_ASAP7_75t_L g862 ( 
.A(n_832),
.Y(n_862)
);

INVx4_ASAP7_75t_L g863 ( 
.A(n_809),
.Y(n_863)
);

AOI21x1_ASAP7_75t_L g864 ( 
.A1(n_843),
.A2(n_769),
.B(n_792),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_L g865 ( 
.A(n_829),
.B(n_760),
.Y(n_865)
);

HB1xp67_ASAP7_75t_L g866 ( 
.A(n_836),
.Y(n_866)
);

INVx2_ASAP7_75t_L g867 ( 
.A(n_804),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_815),
.Y(n_868)
);

OA21x2_ASAP7_75t_L g869 ( 
.A1(n_848),
.A2(n_854),
.B(n_853),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_822),
.Y(n_870)
);

AND2x4_ASAP7_75t_L g871 ( 
.A(n_855),
.B(n_757),
.Y(n_871)
);

AND2x4_ASAP7_75t_L g872 ( 
.A(n_855),
.B(n_770),
.Y(n_872)
);

INVx3_ASAP7_75t_L g873 ( 
.A(n_855),
.Y(n_873)
);

AND2x2_ASAP7_75t_L g874 ( 
.A(n_838),
.B(n_770),
.Y(n_874)
);

CKINVDCx8_ASAP7_75t_R g875 ( 
.A(n_819),
.Y(n_875)
);

HB1xp67_ASAP7_75t_L g876 ( 
.A(n_836),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_849),
.Y(n_877)
);

INVx2_ASAP7_75t_L g878 ( 
.A(n_805),
.Y(n_878)
);

BUFx2_ASAP7_75t_L g879 ( 
.A(n_859),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_824),
.Y(n_880)
);

INVx4_ASAP7_75t_L g881 ( 
.A(n_809),
.Y(n_881)
);

OR2x2_ASAP7_75t_L g882 ( 
.A(n_839),
.B(n_778),
.Y(n_882)
);

INVxp67_ASAP7_75t_L g883 ( 
.A(n_803),
.Y(n_883)
);

AO21x1_ASAP7_75t_L g884 ( 
.A1(n_810),
.A2(n_774),
.B(n_778),
.Y(n_884)
);

BUFx12f_ASAP7_75t_L g885 ( 
.A(n_811),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_826),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_842),
.Y(n_887)
);

BUFx3_ASAP7_75t_L g888 ( 
.A(n_809),
.Y(n_888)
);

INVx2_ASAP7_75t_L g889 ( 
.A(n_841),
.Y(n_889)
);

INVx1_ASAP7_75t_SL g890 ( 
.A(n_821),
.Y(n_890)
);

HB1xp67_ASAP7_75t_L g891 ( 
.A(n_841),
.Y(n_891)
);

BUFx2_ASAP7_75t_L g892 ( 
.A(n_841),
.Y(n_892)
);

AOI22xp33_ASAP7_75t_L g893 ( 
.A1(n_812),
.A2(n_152),
.B1(n_153),
.B2(n_154),
.Y(n_893)
);

OR2x6_ASAP7_75t_L g894 ( 
.A(n_852),
.B(n_155),
.Y(n_894)
);

BUFx3_ASAP7_75t_L g895 ( 
.A(n_828),
.Y(n_895)
);

INVx1_ASAP7_75t_L g896 ( 
.A(n_857),
.Y(n_896)
);

INVx1_ASAP7_75t_L g897 ( 
.A(n_857),
.Y(n_897)
);

OA21x2_ASAP7_75t_L g898 ( 
.A1(n_831),
.A2(n_156),
.B(n_157),
.Y(n_898)
);

OAI21xp5_ASAP7_75t_L g899 ( 
.A1(n_850),
.A2(n_158),
.B(n_159),
.Y(n_899)
);

INVx1_ASAP7_75t_L g900 ( 
.A(n_851),
.Y(n_900)
);

OAI21x1_ASAP7_75t_L g901 ( 
.A1(n_861),
.A2(n_160),
.B(n_161),
.Y(n_901)
);

INVx2_ASAP7_75t_SL g902 ( 
.A(n_828),
.Y(n_902)
);

INVx2_ASAP7_75t_L g903 ( 
.A(n_828),
.Y(n_903)
);

INVx1_ASAP7_75t_L g904 ( 
.A(n_810),
.Y(n_904)
);

INVx2_ASAP7_75t_L g905 ( 
.A(n_833),
.Y(n_905)
);

INVx2_ASAP7_75t_L g906 ( 
.A(n_833),
.Y(n_906)
);

BUFx6f_ASAP7_75t_SL g907 ( 
.A(n_894),
.Y(n_907)
);

INVx2_ASAP7_75t_L g908 ( 
.A(n_867),
.Y(n_908)
);

INVx2_ASAP7_75t_L g909 ( 
.A(n_867),
.Y(n_909)
);

BUFx3_ASAP7_75t_L g910 ( 
.A(n_885),
.Y(n_910)
);

OR2x6_ASAP7_75t_L g911 ( 
.A(n_894),
.B(n_852),
.Y(n_911)
);

AO21x2_ASAP7_75t_L g912 ( 
.A1(n_864),
.A2(n_844),
.B(n_850),
.Y(n_912)
);

INVx1_ASAP7_75t_L g913 ( 
.A(n_862),
.Y(n_913)
);

INVx1_ASAP7_75t_L g914 ( 
.A(n_862),
.Y(n_914)
);

AND2x2_ASAP7_75t_L g915 ( 
.A(n_868),
.B(n_813),
.Y(n_915)
);

AND2x4_ASAP7_75t_L g916 ( 
.A(n_873),
.B(n_834),
.Y(n_916)
);

AOI221xp5_ASAP7_75t_L g917 ( 
.A1(n_904),
.A2(n_806),
.B1(n_813),
.B2(n_814),
.C(n_830),
.Y(n_917)
);

INVx2_ASAP7_75t_L g918 ( 
.A(n_878),
.Y(n_918)
);

NAND2xp5_ASAP7_75t_L g919 ( 
.A(n_880),
.B(n_825),
.Y(n_919)
);

NOR2xp33_ASAP7_75t_L g920 ( 
.A(n_900),
.B(n_820),
.Y(n_920)
);

INVxp67_ASAP7_75t_SL g921 ( 
.A(n_865),
.Y(n_921)
);

HB1xp67_ASAP7_75t_L g922 ( 
.A(n_866),
.Y(n_922)
);

AO21x2_ASAP7_75t_L g923 ( 
.A1(n_864),
.A2(n_830),
.B(n_816),
.Y(n_923)
);

INVx1_ASAP7_75t_SL g924 ( 
.A(n_876),
.Y(n_924)
);

INVx1_ASAP7_75t_L g925 ( 
.A(n_870),
.Y(n_925)
);

AO21x1_ASAP7_75t_L g926 ( 
.A1(n_896),
.A2(n_823),
.B(n_856),
.Y(n_926)
);

AND2x2_ASAP7_75t_L g927 ( 
.A(n_870),
.B(n_825),
.Y(n_927)
);

OR2x6_ASAP7_75t_L g928 ( 
.A(n_894),
.B(n_835),
.Y(n_928)
);

INVx2_ASAP7_75t_L g929 ( 
.A(n_880),
.Y(n_929)
);

INVx2_ASAP7_75t_L g930 ( 
.A(n_869),
.Y(n_930)
);

INVx2_ASAP7_75t_L g931 ( 
.A(n_869),
.Y(n_931)
);

INVx1_ASAP7_75t_L g932 ( 
.A(n_877),
.Y(n_932)
);

AO21x1_ASAP7_75t_SL g933 ( 
.A1(n_896),
.A2(n_858),
.B(n_847),
.Y(n_933)
);

HB1xp67_ASAP7_75t_L g934 ( 
.A(n_886),
.Y(n_934)
);

INVx2_ASAP7_75t_L g935 ( 
.A(n_930),
.Y(n_935)
);

INVx5_ASAP7_75t_L g936 ( 
.A(n_928),
.Y(n_936)
);

INVx1_ASAP7_75t_L g937 ( 
.A(n_932),
.Y(n_937)
);

AND2x2_ASAP7_75t_L g938 ( 
.A(n_922),
.B(n_883),
.Y(n_938)
);

INVx1_ASAP7_75t_L g939 ( 
.A(n_932),
.Y(n_939)
);

NAND3xp33_ASAP7_75t_L g940 ( 
.A(n_917),
.B(n_899),
.C(n_897),
.Y(n_940)
);

AND2x2_ASAP7_75t_L g941 ( 
.A(n_924),
.B(n_879),
.Y(n_941)
);

AND2x2_ASAP7_75t_L g942 ( 
.A(n_924),
.B(n_879),
.Y(n_942)
);

INVx2_ASAP7_75t_L g943 ( 
.A(n_930),
.Y(n_943)
);

NAND2xp5_ASAP7_75t_L g944 ( 
.A(n_915),
.B(n_887),
.Y(n_944)
);

INVx2_ASAP7_75t_L g945 ( 
.A(n_931),
.Y(n_945)
);

BUFx2_ASAP7_75t_L g946 ( 
.A(n_921),
.Y(n_946)
);

INVx2_ASAP7_75t_L g947 ( 
.A(n_931),
.Y(n_947)
);

INVx2_ASAP7_75t_L g948 ( 
.A(n_913),
.Y(n_948)
);

AND2x2_ASAP7_75t_L g949 ( 
.A(n_918),
.B(n_874),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_L g950 ( 
.A(n_915),
.B(n_887),
.Y(n_950)
);

OR2x2_ASAP7_75t_L g951 ( 
.A(n_934),
.B(n_869),
.Y(n_951)
);

OAI211xp5_ASAP7_75t_L g952 ( 
.A1(n_927),
.A2(n_897),
.B(n_904),
.C(n_893),
.Y(n_952)
);

BUFx3_ASAP7_75t_L g953 ( 
.A(n_910),
.Y(n_953)
);

AND2x2_ASAP7_75t_L g954 ( 
.A(n_918),
.B(n_874),
.Y(n_954)
);

INVxp67_ASAP7_75t_L g955 ( 
.A(n_920),
.Y(n_955)
);

INVx1_ASAP7_75t_L g956 ( 
.A(n_937),
.Y(n_956)
);

AND2x2_ASAP7_75t_L g957 ( 
.A(n_936),
.B(n_916),
.Y(n_957)
);

INVx2_ASAP7_75t_L g958 ( 
.A(n_935),
.Y(n_958)
);

AND2x2_ASAP7_75t_L g959 ( 
.A(n_936),
.B(n_916),
.Y(n_959)
);

OR2x2_ASAP7_75t_L g960 ( 
.A(n_946),
.B(n_908),
.Y(n_960)
);

NAND2xp5_ASAP7_75t_L g961 ( 
.A(n_944),
.B(n_927),
.Y(n_961)
);

AND2x2_ASAP7_75t_L g962 ( 
.A(n_936),
.B(n_916),
.Y(n_962)
);

BUFx2_ASAP7_75t_L g963 ( 
.A(n_936),
.Y(n_963)
);

NAND2xp5_ASAP7_75t_L g964 ( 
.A(n_950),
.B(n_929),
.Y(n_964)
);

AND2x2_ASAP7_75t_L g965 ( 
.A(n_936),
.B(n_916),
.Y(n_965)
);

INVx1_ASAP7_75t_L g966 ( 
.A(n_937),
.Y(n_966)
);

INVx1_ASAP7_75t_L g967 ( 
.A(n_939),
.Y(n_967)
);

AND2x2_ASAP7_75t_L g968 ( 
.A(n_936),
.B(n_908),
.Y(n_968)
);

AOI22xp33_ASAP7_75t_L g969 ( 
.A1(n_940),
.A2(n_907),
.B1(n_911),
.B2(n_926),
.Y(n_969)
);

NOR2xp33_ASAP7_75t_L g970 ( 
.A(n_953),
.B(n_910),
.Y(n_970)
);

AND2x2_ASAP7_75t_L g971 ( 
.A(n_946),
.B(n_909),
.Y(n_971)
);

INVx1_ASAP7_75t_L g972 ( 
.A(n_939),
.Y(n_972)
);

BUFx2_ASAP7_75t_L g973 ( 
.A(n_963),
.Y(n_973)
);

INVx1_ASAP7_75t_L g974 ( 
.A(n_956),
.Y(n_974)
);

HB1xp67_ASAP7_75t_L g975 ( 
.A(n_966),
.Y(n_975)
);

NAND2xp5_ASAP7_75t_L g976 ( 
.A(n_961),
.B(n_938),
.Y(n_976)
);

BUFx2_ASAP7_75t_L g977 ( 
.A(n_963),
.Y(n_977)
);

AND2x2_ASAP7_75t_L g978 ( 
.A(n_957),
.B(n_941),
.Y(n_978)
);

INVx1_ASAP7_75t_L g979 ( 
.A(n_967),
.Y(n_979)
);

AND2x2_ASAP7_75t_L g980 ( 
.A(n_957),
.B(n_938),
.Y(n_980)
);

AND2x4_ASAP7_75t_SL g981 ( 
.A(n_959),
.B(n_928),
.Y(n_981)
);

INVx1_ASAP7_75t_L g982 ( 
.A(n_972),
.Y(n_982)
);

INVx2_ASAP7_75t_L g983 ( 
.A(n_958),
.Y(n_983)
);

AND2x2_ASAP7_75t_L g984 ( 
.A(n_980),
.B(n_959),
.Y(n_984)
);

INVx2_ASAP7_75t_L g985 ( 
.A(n_973),
.Y(n_985)
);

INVx1_ASAP7_75t_L g986 ( 
.A(n_975),
.Y(n_986)
);

OR2x2_ASAP7_75t_L g987 ( 
.A(n_976),
.B(n_964),
.Y(n_987)
);

INVx1_ASAP7_75t_L g988 ( 
.A(n_975),
.Y(n_988)
);

AND3x2_ASAP7_75t_L g989 ( 
.A(n_977),
.B(n_970),
.C(n_891),
.Y(n_989)
);

AND2x2_ASAP7_75t_L g990 ( 
.A(n_981),
.B(n_962),
.Y(n_990)
);

INVx1_ASAP7_75t_L g991 ( 
.A(n_974),
.Y(n_991)
);

NAND2xp5_ASAP7_75t_L g992 ( 
.A(n_985),
.B(n_978),
.Y(n_992)
);

OR2x2_ASAP7_75t_L g993 ( 
.A(n_985),
.B(n_978),
.Y(n_993)
);

CKINVDCx20_ASAP7_75t_R g994 ( 
.A(n_990),
.Y(n_994)
);

INVxp67_ASAP7_75t_L g995 ( 
.A(n_986),
.Y(n_995)
);

NAND2xp5_ASAP7_75t_L g996 ( 
.A(n_991),
.B(n_979),
.Y(n_996)
);

CKINVDCx5p33_ASAP7_75t_R g997 ( 
.A(n_988),
.Y(n_997)
);

INVx2_ASAP7_75t_L g998 ( 
.A(n_994),
.Y(n_998)
);

INVx1_ASAP7_75t_SL g999 ( 
.A(n_993),
.Y(n_999)
);

NAND2x1p5_ASAP7_75t_L g1000 ( 
.A(n_992),
.B(n_890),
.Y(n_1000)
);

INVx2_ASAP7_75t_SL g1001 ( 
.A(n_997),
.Y(n_1001)
);

AND2x4_ASAP7_75t_L g1002 ( 
.A(n_995),
.B(n_984),
.Y(n_1002)
);

INVx1_ASAP7_75t_SL g1003 ( 
.A(n_996),
.Y(n_1003)
);

NOR2x1_ASAP7_75t_L g1004 ( 
.A(n_994),
.B(n_953),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_L g1005 ( 
.A(n_997),
.B(n_989),
.Y(n_1005)
);

NOR2xp33_ASAP7_75t_L g1006 ( 
.A(n_994),
.B(n_885),
.Y(n_1006)
);

NAND2xp5_ASAP7_75t_L g1007 ( 
.A(n_997),
.B(n_989),
.Y(n_1007)
);

INVxp67_ASAP7_75t_SL g1008 ( 
.A(n_1004),
.Y(n_1008)
);

NOR3xp33_ASAP7_75t_L g1009 ( 
.A(n_998),
.B(n_900),
.C(n_952),
.Y(n_1009)
);

INVx1_ASAP7_75t_L g1010 ( 
.A(n_999),
.Y(n_1010)
);

AOI22xp5_ASAP7_75t_L g1011 ( 
.A1(n_1001),
.A2(n_1002),
.B1(n_1007),
.B2(n_1005),
.Y(n_1011)
);

NOR4xp25_ASAP7_75t_L g1012 ( 
.A(n_1003),
.B(n_1006),
.C(n_969),
.D(n_1002),
.Y(n_1012)
);

INVx1_ASAP7_75t_L g1013 ( 
.A(n_1000),
.Y(n_1013)
);

AOI22xp5_ASAP7_75t_L g1014 ( 
.A1(n_998),
.A2(n_907),
.B1(n_926),
.B2(n_981),
.Y(n_1014)
);

INVx1_ASAP7_75t_L g1015 ( 
.A(n_999),
.Y(n_1015)
);

INVx2_ASAP7_75t_L g1016 ( 
.A(n_1013),
.Y(n_1016)
);

AOI22xp5_ASAP7_75t_L g1017 ( 
.A1(n_1009),
.A2(n_907),
.B1(n_962),
.B2(n_965),
.Y(n_1017)
);

NAND2xp5_ASAP7_75t_L g1018 ( 
.A(n_1008),
.B(n_987),
.Y(n_1018)
);

NAND2xp5_ASAP7_75t_L g1019 ( 
.A(n_1010),
.B(n_982),
.Y(n_1019)
);

OAI21xp5_ASAP7_75t_SL g1020 ( 
.A1(n_1011),
.A2(n_965),
.B(n_955),
.Y(n_1020)
);

AND2x2_ASAP7_75t_L g1021 ( 
.A(n_1015),
.B(n_983),
.Y(n_1021)
);

INVx1_ASAP7_75t_L g1022 ( 
.A(n_1014),
.Y(n_1022)
);

O2A1O1Ixp33_ASAP7_75t_L g1023 ( 
.A1(n_1012),
.A2(n_894),
.B(n_928),
.C(n_911),
.Y(n_1023)
);

INVx2_ASAP7_75t_L g1024 ( 
.A(n_1016),
.Y(n_1024)
);

AOI211xp5_ASAP7_75t_SL g1025 ( 
.A1(n_1022),
.A2(n_808),
.B(n_817),
.C(n_875),
.Y(n_1025)
);

OAI21xp5_ASAP7_75t_SL g1026 ( 
.A1(n_1023),
.A2(n_892),
.B(n_889),
.Y(n_1026)
);

OAI22xp5_ASAP7_75t_L g1027 ( 
.A1(n_1017),
.A2(n_875),
.B1(n_911),
.B2(n_928),
.Y(n_1027)
);

AOI322xp5_ASAP7_75t_L g1028 ( 
.A1(n_1018),
.A2(n_983),
.A3(n_942),
.B1(n_941),
.B2(n_919),
.C1(n_968),
.C2(n_892),
.Y(n_1028)
);

NAND3xp33_ASAP7_75t_L g1029 ( 
.A(n_1020),
.B(n_898),
.C(n_905),
.Y(n_1029)
);

OAI21xp33_ASAP7_75t_L g1030 ( 
.A1(n_1019),
.A2(n_928),
.B(n_889),
.Y(n_1030)
);

INVx1_ASAP7_75t_L g1031 ( 
.A(n_1024),
.Y(n_1031)
);

INVx1_ASAP7_75t_L g1032 ( 
.A(n_1026),
.Y(n_1032)
);

INVx1_ASAP7_75t_L g1033 ( 
.A(n_1030),
.Y(n_1033)
);

INVx1_ASAP7_75t_L g1034 ( 
.A(n_1029),
.Y(n_1034)
);

INVx1_ASAP7_75t_L g1035 ( 
.A(n_1027),
.Y(n_1035)
);

INVx2_ASAP7_75t_L g1036 ( 
.A(n_1025),
.Y(n_1036)
);

INVx1_ASAP7_75t_L g1037 ( 
.A(n_1028),
.Y(n_1037)
);

INVx1_ASAP7_75t_L g1038 ( 
.A(n_1024),
.Y(n_1038)
);

INVx1_ASAP7_75t_SL g1039 ( 
.A(n_1024),
.Y(n_1039)
);

INVx1_ASAP7_75t_L g1040 ( 
.A(n_1024),
.Y(n_1040)
);

INVxp67_ASAP7_75t_SL g1041 ( 
.A(n_1024),
.Y(n_1041)
);

NOR3x1_ASAP7_75t_L g1042 ( 
.A(n_1037),
.B(n_1021),
.C(n_902),
.Y(n_1042)
);

OAI211xp5_ASAP7_75t_SL g1043 ( 
.A1(n_1036),
.A2(n_846),
.B(n_845),
.C(n_827),
.Y(n_1043)
);

NAND5xp2_ASAP7_75t_L g1044 ( 
.A(n_1035),
.B(n_818),
.C(n_837),
.D(n_860),
.E(n_968),
.Y(n_1044)
);

INVx1_ASAP7_75t_L g1045 ( 
.A(n_1041),
.Y(n_1045)
);

AND2x4_ASAP7_75t_L g1046 ( 
.A(n_1039),
.B(n_971),
.Y(n_1046)
);

NAND3xp33_ASAP7_75t_L g1047 ( 
.A(n_1031),
.B(n_905),
.C(n_906),
.Y(n_1047)
);

NOR3xp33_ASAP7_75t_L g1048 ( 
.A(n_1038),
.B(n_906),
.C(n_863),
.Y(n_1048)
);

NOR2x1_ASAP7_75t_L g1049 ( 
.A(n_1039),
.B(n_960),
.Y(n_1049)
);

INVx1_ASAP7_75t_L g1050 ( 
.A(n_1040),
.Y(n_1050)
);

INVx1_ASAP7_75t_L g1051 ( 
.A(n_1033),
.Y(n_1051)
);

OA22x2_ASAP7_75t_SL g1052 ( 
.A1(n_1032),
.A2(n_958),
.B1(n_807),
.B2(n_903),
.Y(n_1052)
);

NAND2xp5_ASAP7_75t_L g1053 ( 
.A(n_1046),
.B(n_1034),
.Y(n_1053)
);

NOR3xp33_ASAP7_75t_L g1054 ( 
.A(n_1051),
.B(n_863),
.C(n_881),
.Y(n_1054)
);

AOI221xp5_ASAP7_75t_L g1055 ( 
.A1(n_1045),
.A2(n_1048),
.B1(n_1050),
.B2(n_1047),
.C(n_1052),
.Y(n_1055)
);

NOR2xp33_ASAP7_75t_L g1056 ( 
.A(n_1049),
.B(n_807),
.Y(n_1056)
);

OAI21xp5_ASAP7_75t_L g1057 ( 
.A1(n_1043),
.A2(n_894),
.B(n_960),
.Y(n_1057)
);

NAND2xp5_ASAP7_75t_L g1058 ( 
.A(n_1042),
.B(n_971),
.Y(n_1058)
);

INVx1_ASAP7_75t_L g1059 ( 
.A(n_1044),
.Y(n_1059)
);

AOI21xp33_ASAP7_75t_L g1060 ( 
.A1(n_1051),
.A2(n_898),
.B(n_911),
.Y(n_1060)
);

OAI221xp5_ASAP7_75t_SL g1061 ( 
.A1(n_1055),
.A2(n_1053),
.B1(n_1058),
.B2(n_1054),
.C(n_1059),
.Y(n_1061)
);

NAND2xp5_ASAP7_75t_L g1062 ( 
.A(n_1056),
.B(n_942),
.Y(n_1062)
);

NAND4xp25_ASAP7_75t_L g1063 ( 
.A(n_1057),
.B(n_895),
.C(n_888),
.D(n_863),
.Y(n_1063)
);

NOR2xp33_ASAP7_75t_L g1064 ( 
.A(n_1060),
.B(n_840),
.Y(n_1064)
);

OAI21xp5_ASAP7_75t_L g1065 ( 
.A1(n_1053),
.A2(n_911),
.B(n_898),
.Y(n_1065)
);

NOR3xp33_ASAP7_75t_L g1066 ( 
.A(n_1053),
.B(n_881),
.C(n_902),
.Y(n_1066)
);

INVx2_ASAP7_75t_L g1067 ( 
.A(n_1058),
.Y(n_1067)
);

OR3x1_ASAP7_75t_L g1068 ( 
.A(n_1056),
.B(n_913),
.C(n_925),
.Y(n_1068)
);

NAND2xp5_ASAP7_75t_SL g1069 ( 
.A(n_1056),
.B(n_895),
.Y(n_1069)
);

NAND2xp5_ASAP7_75t_L g1070 ( 
.A(n_1067),
.B(n_943),
.Y(n_1070)
);

NAND5xp2_ASAP7_75t_L g1071 ( 
.A(n_1061),
.B(n_933),
.C(n_886),
.D(n_898),
.E(n_167),
.Y(n_1071)
);

AND2x4_ASAP7_75t_L g1072 ( 
.A(n_1066),
.B(n_888),
.Y(n_1072)
);

NAND3xp33_ASAP7_75t_L g1073 ( 
.A(n_1064),
.B(n_951),
.C(n_881),
.Y(n_1073)
);

NAND2xp5_ASAP7_75t_L g1074 ( 
.A(n_1062),
.B(n_943),
.Y(n_1074)
);

AND2x4_ASAP7_75t_L g1075 ( 
.A(n_1069),
.B(n_903),
.Y(n_1075)
);

NOR2xp67_ASAP7_75t_SL g1076 ( 
.A(n_1063),
.B(n_162),
.Y(n_1076)
);

NOR2x1_ASAP7_75t_L g1077 ( 
.A(n_1068),
.B(n_912),
.Y(n_1077)
);

AND4x2_ASAP7_75t_L g1078 ( 
.A(n_1065),
.B(n_933),
.C(n_912),
.D(n_935),
.Y(n_1078)
);

AND2x2_ASAP7_75t_L g1079 ( 
.A(n_1067),
.B(n_954),
.Y(n_1079)
);

AND3x4_ASAP7_75t_L g1080 ( 
.A(n_1072),
.B(n_872),
.C(n_871),
.Y(n_1080)
);

XNOR2xp5_ASAP7_75t_L g1081 ( 
.A(n_1079),
.B(n_163),
.Y(n_1081)
);

NAND4xp75_ASAP7_75t_L g1082 ( 
.A(n_1070),
.B(n_1077),
.C(n_1074),
.D(n_1076),
.Y(n_1082)
);

NOR3xp33_ASAP7_75t_L g1083 ( 
.A(n_1073),
.B(n_901),
.C(n_873),
.Y(n_1083)
);

OAI21xp5_ASAP7_75t_L g1084 ( 
.A1(n_1075),
.A2(n_945),
.B(n_947),
.Y(n_1084)
);

INVx2_ASAP7_75t_SL g1085 ( 
.A(n_1078),
.Y(n_1085)
);

OAI22xp5_ASAP7_75t_L g1086 ( 
.A1(n_1073),
.A2(n_951),
.B1(n_945),
.B2(n_947),
.Y(n_1086)
);

AND3x1_ASAP7_75t_L g1087 ( 
.A(n_1071),
.B(n_948),
.C(n_949),
.Y(n_1087)
);

INVx1_ASAP7_75t_L g1088 ( 
.A(n_1079),
.Y(n_1088)
);

NAND2xp5_ASAP7_75t_SL g1089 ( 
.A(n_1072),
.B(n_948),
.Y(n_1089)
);

HB1xp67_ASAP7_75t_L g1090 ( 
.A(n_1070),
.Y(n_1090)
);

NOR2xp67_ASAP7_75t_L g1091 ( 
.A(n_1071),
.B(n_164),
.Y(n_1091)
);

BUFx2_ASAP7_75t_L g1092 ( 
.A(n_1088),
.Y(n_1092)
);

XNOR2x1_ASAP7_75t_L g1093 ( 
.A(n_1081),
.B(n_1082),
.Y(n_1093)
);

XNOR2x1_ASAP7_75t_L g1094 ( 
.A(n_1091),
.B(n_168),
.Y(n_1094)
);

OAI21xp5_ASAP7_75t_L g1095 ( 
.A1(n_1085),
.A2(n_882),
.B(n_872),
.Y(n_1095)
);

INVx1_ASAP7_75t_L g1096 ( 
.A(n_1087),
.Y(n_1096)
);

AOI21xp5_ASAP7_75t_L g1097 ( 
.A1(n_1090),
.A2(n_912),
.B(n_923),
.Y(n_1097)
);

INVx1_ASAP7_75t_L g1098 ( 
.A(n_1089),
.Y(n_1098)
);

XNOR2xp5_ASAP7_75t_L g1099 ( 
.A(n_1080),
.B(n_169),
.Y(n_1099)
);

INVx1_ASAP7_75t_L g1100 ( 
.A(n_1092),
.Y(n_1100)
);

INVx1_ASAP7_75t_SL g1101 ( 
.A(n_1094),
.Y(n_1101)
);

INVx3_ASAP7_75t_L g1102 ( 
.A(n_1098),
.Y(n_1102)
);

AOI22xp33_ASAP7_75t_L g1103 ( 
.A1(n_1096),
.A2(n_1083),
.B1(n_1086),
.B2(n_1084),
.Y(n_1103)
);

AND4x2_ASAP7_75t_L g1104 ( 
.A(n_1093),
.B(n_170),
.C(n_171),
.D(n_173),
.Y(n_1104)
);

INVx1_ASAP7_75t_L g1105 ( 
.A(n_1099),
.Y(n_1105)
);

NAND2xp5_ASAP7_75t_L g1106 ( 
.A(n_1100),
.B(n_1095),
.Y(n_1106)
);

INVxp33_ASAP7_75t_SL g1107 ( 
.A(n_1101),
.Y(n_1107)
);

INVx4_ASAP7_75t_L g1108 ( 
.A(n_1102),
.Y(n_1108)
);

INVx1_ASAP7_75t_L g1109 ( 
.A(n_1108),
.Y(n_1109)
);

INVx1_ASAP7_75t_L g1110 ( 
.A(n_1109),
.Y(n_1110)
);

NOR2xp67_ASAP7_75t_L g1111 ( 
.A(n_1110),
.B(n_1106),
.Y(n_1111)
);

OAI22xp5_ASAP7_75t_L g1112 ( 
.A1(n_1111),
.A2(n_1103),
.B1(n_1107),
.B2(n_1105),
.Y(n_1112)
);

OAI21x1_ASAP7_75t_L g1113 ( 
.A1(n_1111),
.A2(n_1104),
.B(n_1097),
.Y(n_1113)
);

OR2x6_ASAP7_75t_L g1114 ( 
.A(n_1112),
.B(n_1113),
.Y(n_1114)
);

AOI21x1_ASAP7_75t_L g1115 ( 
.A1(n_1112),
.A2(n_176),
.B(n_177),
.Y(n_1115)
);

AO221x2_ASAP7_75t_L g1116 ( 
.A1(n_1114),
.A2(n_178),
.B1(n_179),
.B2(n_180),
.C(n_183),
.Y(n_1116)
);

OAI21xp5_ASAP7_75t_L g1117 ( 
.A1(n_1115),
.A2(n_186),
.B(n_187),
.Y(n_1117)
);

AOI221xp5_ASAP7_75t_L g1118 ( 
.A1(n_1117),
.A2(n_188),
.B1(n_191),
.B2(n_202),
.C(n_914),
.Y(n_1118)
);

AOI211xp5_ASAP7_75t_L g1119 ( 
.A1(n_1118),
.A2(n_1116),
.B(n_884),
.C(n_871),
.Y(n_1119)
);


endmodule