module fake_jpeg_7922_n_269 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_269);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_269;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_140;
wire n_82;
wire n_128;
wire n_100;
wire n_258;
wire n_96;

INVx1_ASAP7_75t_L g15 ( 
.A(n_6),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_2),
.Y(n_16)
);

INVx4_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_7),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

HB1xp67_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

INVx1_ASAP7_75t_SL g24 ( 
.A(n_0),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_14),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_14),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_10),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_2),
.Y(n_30)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_21),
.Y(n_32)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_32),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_21),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_33),
.B(n_34),
.Y(n_56)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_21),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_18),
.Y(n_35)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_35),
.Y(n_55)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_22),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_36),
.B(n_37),
.Y(n_58)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_18),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_18),
.Y(n_38)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_38),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_18),
.Y(n_39)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_39),
.Y(n_66)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_15),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_40),
.B(n_42),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_20),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_41),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_30),
.B(n_0),
.Y(n_42)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_35),
.Y(n_43)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_43),
.Y(n_83)
);

OAI22xp33_ASAP7_75t_SL g44 ( 
.A1(n_36),
.A2(n_17),
.B1(n_31),
.B2(n_27),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_44),
.A2(n_28),
.B1(n_19),
.B2(n_25),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_37),
.A2(n_17),
.B1(n_24),
.B2(n_31),
.Y(n_45)
);

INVxp67_ASAP7_75t_L g68 ( 
.A(n_45),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g46 ( 
.A1(n_42),
.A2(n_31),
.B1(n_17),
.B2(n_30),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_46),
.A2(n_49),
.B1(n_50),
.B2(n_62),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_SL g47 ( 
.A(n_40),
.B(n_25),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_47),
.B(n_51),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_33),
.A2(n_24),
.B1(n_27),
.B2(n_15),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_34),
.A2(n_24),
.B1(n_27),
.B2(n_15),
.Y(n_50)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_35),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_SL g52 ( 
.A(n_32),
.B(n_29),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_52),
.B(n_54),
.Y(n_74)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_38),
.Y(n_59)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_59),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_39),
.B(n_23),
.Y(n_61)
);

AND2x2_ASAP7_75t_SL g69 ( 
.A(n_61),
.B(n_23),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_41),
.A2(n_29),
.B1(n_28),
.B2(n_19),
.Y(n_62)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_39),
.Y(n_63)
);

HB1xp67_ASAP7_75t_L g81 ( 
.A(n_63),
.Y(n_81)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_32),
.Y(n_64)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_64),
.B(n_65),
.Y(n_77)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_42),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_69),
.B(n_20),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_57),
.Y(n_70)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_70),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_L g72 ( 
.A1(n_65),
.A2(n_29),
.B1(n_28),
.B2(n_19),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_72),
.A2(n_78),
.B1(n_84),
.B2(n_16),
.Y(n_89)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_51),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_73),
.B(n_54),
.Y(n_104)
);

AND2x2_ASAP7_75t_SL g75 ( 
.A(n_60),
.B(n_23),
.Y(n_75)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_75),
.B(n_26),
.C(n_20),
.Y(n_105)
);

NAND2x1_ASAP7_75t_SL g76 ( 
.A(n_57),
.B(n_20),
.Y(n_76)
);

OAI21xp5_ASAP7_75t_L g103 ( 
.A1(n_76),
.A2(n_55),
.B(n_63),
.Y(n_103)
);

CKINVDCx14_ASAP7_75t_R g79 ( 
.A(n_47),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g91 ( 
.A(n_79),
.B(n_86),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_61),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_80),
.B(n_64),
.Y(n_95)
);

BUFx2_ASAP7_75t_L g82 ( 
.A(n_57),
.Y(n_82)
);

BUFx2_ASAP7_75t_L g101 ( 
.A(n_82),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_L g84 ( 
.A1(n_60),
.A2(n_25),
.B1(n_30),
.B2(n_16),
.Y(n_84)
);

OR2x2_ASAP7_75t_L g86 ( 
.A(n_52),
.B(n_56),
.Y(n_86)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_53),
.Y(n_87)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_87),
.Y(n_100)
);

AOI21xp5_ASAP7_75t_L g88 ( 
.A1(n_68),
.A2(n_46),
.B(n_58),
.Y(n_88)
);

OAI21xp5_ASAP7_75t_L g128 ( 
.A1(n_88),
.A2(n_98),
.B(n_103),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_89),
.B(n_92),
.Y(n_114)
);

AND2x6_ASAP7_75t_L g90 ( 
.A(n_77),
.B(n_11),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_90),
.Y(n_112)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_71),
.Y(n_92)
);

XNOR2xp5_ASAP7_75t_L g93 ( 
.A(n_85),
.B(n_56),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_93),
.B(n_75),
.C(n_69),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_85),
.A2(n_58),
.B1(n_55),
.B2(n_66),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_94),
.A2(n_55),
.B1(n_87),
.B2(n_76),
.Y(n_120)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_95),
.Y(n_113)
);

O2A1O1Ixp33_ASAP7_75t_L g96 ( 
.A1(n_74),
.A2(n_59),
.B(n_22),
.C(n_43),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_96),
.A2(n_67),
.B1(n_77),
.B2(n_26),
.Y(n_127)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_71),
.Y(n_99)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_99),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_86),
.B(n_53),
.Y(n_102)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_102),
.Y(n_119)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_104),
.Y(n_121)
);

AND2x2_ASAP7_75t_L g117 ( 
.A(n_105),
.B(n_76),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_86),
.B(n_53),
.Y(n_106)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_106),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_69),
.B(n_66),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_107),
.B(n_108),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_69),
.B(n_48),
.Y(n_108)
);

HB1xp67_ASAP7_75t_L g109 ( 
.A(n_82),
.Y(n_109)
);

INVx1_ASAP7_75t_SL g130 ( 
.A(n_109),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_110),
.B(n_111),
.C(n_122),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_93),
.B(n_80),
.C(n_75),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_88),
.A2(n_79),
.B1(n_74),
.B2(n_78),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_115),
.A2(n_120),
.B1(n_125),
.B2(n_96),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_SL g136 ( 
.A1(n_117),
.A2(n_103),
.B(n_106),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_91),
.B(n_99),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_SL g150 ( 
.A(n_118),
.B(n_12),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_107),
.B(n_75),
.C(n_77),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_101),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_123),
.B(n_124),
.Y(n_139)
);

CKINVDCx16_ASAP7_75t_R g124 ( 
.A(n_101),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_94),
.A2(n_48),
.B1(n_43),
.B2(n_87),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_108),
.B(n_77),
.C(n_67),
.Y(n_126)
);

XOR2xp5_ASAP7_75t_L g156 ( 
.A(n_126),
.B(n_129),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_L g151 ( 
.A1(n_127),
.A2(n_133),
.B(n_116),
.Y(n_151)
);

XOR2xp5_ASAP7_75t_L g129 ( 
.A(n_98),
.B(n_26),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_92),
.A2(n_11),
.B1(n_13),
.B2(n_3),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_114),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_134),
.B(n_137),
.Y(n_168)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_125),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_135),
.B(n_144),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_136),
.B(n_147),
.C(n_129),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_120),
.A2(n_119),
.B1(n_132),
.B2(n_112),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_138),
.A2(n_141),
.B1(n_113),
.B2(n_117),
.Y(n_160)
);

CKINVDCx16_ASAP7_75t_R g140 ( 
.A(n_130),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_140),
.B(n_157),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_119),
.A2(n_102),
.B1(n_89),
.B2(n_91),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_131),
.B(n_95),
.Y(n_142)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_142),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_131),
.B(n_105),
.Y(n_143)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_143),
.Y(n_163)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_130),
.Y(n_144)
);

AND2x2_ASAP7_75t_L g145 ( 
.A(n_132),
.B(n_90),
.Y(n_145)
);

AOI21xp5_ASAP7_75t_L g171 ( 
.A1(n_145),
.A2(n_152),
.B(n_117),
.Y(n_171)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_116),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_146),
.B(n_149),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_L g147 ( 
.A(n_110),
.B(n_81),
.Y(n_147)
);

AOI21xp5_ASAP7_75t_L g148 ( 
.A1(n_128),
.A2(n_100),
.B(n_83),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_SL g173 ( 
.A1(n_148),
.A2(n_151),
.B(n_82),
.Y(n_173)
);

OR2x2_ASAP7_75t_L g149 ( 
.A(n_127),
.B(n_83),
.Y(n_149)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_150),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_SL g152 ( 
.A1(n_128),
.A2(n_83),
.B(n_81),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_113),
.B(n_73),
.Y(n_153)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_153),
.Y(n_165)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_121),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_154),
.B(n_101),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_133),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_139),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_159),
.B(n_138),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_160),
.A2(n_178),
.B1(n_157),
.B2(n_149),
.Y(n_193)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_164),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g166 ( 
.A(n_156),
.B(n_111),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_166),
.B(n_167),
.C(n_155),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_142),
.B(n_126),
.Y(n_169)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_169),
.Y(n_188)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_153),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_170),
.B(n_174),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_L g201 ( 
.A1(n_171),
.A2(n_176),
.B(n_9),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_141),
.B(n_122),
.Y(n_172)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_172),
.Y(n_192)
);

AOI21xp5_ASAP7_75t_L g182 ( 
.A1(n_173),
.A2(n_152),
.B(n_136),
.Y(n_182)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_146),
.Y(n_174)
);

NOR2xp67_ASAP7_75t_SL g176 ( 
.A(n_145),
.B(n_9),
.Y(n_176)
);

INVx3_ASAP7_75t_L g177 ( 
.A(n_144),
.Y(n_177)
);

AOI22xp33_ASAP7_75t_L g184 ( 
.A1(n_177),
.A2(n_97),
.B1(n_154),
.B2(n_134),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_135),
.A2(n_97),
.B1(n_70),
.B2(n_0),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_150),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_180),
.Y(n_197)
);

AOI21xp5_ASAP7_75t_SL g181 ( 
.A1(n_162),
.A2(n_145),
.B(n_151),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_L g204 ( 
.A1(n_181),
.A2(n_182),
.B(n_201),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_183),
.B(n_190),
.C(n_172),
.Y(n_203)
);

OAI22xp33_ASAP7_75t_SL g212 ( 
.A1(n_184),
.A2(n_198),
.B1(n_165),
.B2(n_180),
.Y(n_212)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_187),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_161),
.B(n_143),
.Y(n_189)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_189),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_166),
.B(n_167),
.C(n_156),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_177),
.B(n_137),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_191),
.B(n_194),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_193),
.A2(n_196),
.B1(n_199),
.B2(n_192),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_164),
.B(n_149),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_161),
.B(n_148),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_195),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_168),
.A2(n_147),
.B1(n_155),
.B2(n_70),
.Y(n_196)
);

INVxp67_ASAP7_75t_L g198 ( 
.A(n_179),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_160),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_199)
);

CKINVDCx16_ASAP7_75t_R g200 ( 
.A(n_158),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_200),
.B(n_173),
.Y(n_216)
);

XOR2xp5_ASAP7_75t_L g202 ( 
.A(n_190),
.B(n_171),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_202),
.B(n_210),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_203),
.B(n_207),
.C(n_217),
.Y(n_220)
);

FAx1_ASAP7_75t_L g205 ( 
.A(n_195),
.B(n_162),
.CI(n_158),
.CON(n_205),
.SN(n_205)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_205),
.B(n_211),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_183),
.B(n_163),
.C(n_169),
.Y(n_207)
);

AO221x1_ASAP7_75t_L g208 ( 
.A1(n_198),
.A2(n_174),
.B1(n_178),
.B2(n_170),
.C(n_165),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_208),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g210 ( 
.A(n_196),
.B(n_182),
.Y(n_210)
);

HB1xp67_ASAP7_75t_L g211 ( 
.A(n_200),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_SL g221 ( 
.A(n_212),
.B(n_213),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_216),
.B(n_197),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_192),
.B(n_163),
.C(n_175),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_188),
.B(n_1),
.C(n_3),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_218),
.B(n_201),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_206),
.A2(n_193),
.B1(n_199),
.B2(n_197),
.Y(n_219)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_219),
.Y(n_235)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_222),
.Y(n_244)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_202),
.B(n_181),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_224),
.B(n_227),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_225),
.B(n_11),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_217),
.B(n_186),
.Y(n_226)
);

OAI21xp5_ASAP7_75t_SL g240 ( 
.A1(n_226),
.A2(n_231),
.B(n_4),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g227 ( 
.A(n_210),
.B(n_186),
.Y(n_227)
);

AND2x2_ASAP7_75t_L g229 ( 
.A(n_215),
.B(n_185),
.Y(n_229)
);

AOI21xp5_ASAP7_75t_L g237 ( 
.A1(n_229),
.A2(n_232),
.B(n_10),
.Y(n_237)
);

BUFx24_ASAP7_75t_SL g231 ( 
.A(n_205),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_SL g232 ( 
.A(n_218),
.B(n_185),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_220),
.B(n_207),
.C(n_203),
.Y(n_233)
);

OAI21xp5_ASAP7_75t_L g251 ( 
.A1(n_233),
.A2(n_236),
.B(n_238),
.Y(n_251)
);

FAx1_ASAP7_75t_SL g234 ( 
.A(n_230),
.B(n_205),
.CI(n_204),
.CON(n_234),
.SN(n_234)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_234),
.B(n_223),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_220),
.B(n_209),
.C(n_214),
.Y(n_236)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_237),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_227),
.B(n_10),
.C(n_4),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_239),
.B(n_224),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_240),
.B(n_242),
.Y(n_252)
);

AOI21xp5_ASAP7_75t_L g241 ( 
.A1(n_229),
.A2(n_4),
.B(n_5),
.Y(n_241)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_241),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_223),
.B(n_5),
.C(n_6),
.Y(n_242)
);

AOI21xp5_ASAP7_75t_SL g245 ( 
.A1(n_235),
.A2(n_221),
.B(n_228),
.Y(n_245)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_245),
.Y(n_254)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_247),
.Y(n_258)
);

MAJx2_ASAP7_75t_L g250 ( 
.A(n_243),
.B(n_5),
.C(n_6),
.Y(n_250)
);

OAI21xp5_ASAP7_75t_SL g256 ( 
.A1(n_250),
.A2(n_253),
.B(n_12),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_244),
.B(n_1),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_249),
.B(n_242),
.Y(n_255)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_255),
.Y(n_262)
);

AOI21xp5_ASAP7_75t_L g261 ( 
.A1(n_256),
.A2(n_259),
.B(n_253),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_251),
.B(n_233),
.C(n_236),
.Y(n_257)
);

OAI21xp5_ASAP7_75t_L g260 ( 
.A1(n_257),
.A2(n_238),
.B(n_234),
.Y(n_260)
);

OAI21xp5_ASAP7_75t_SL g259 ( 
.A1(n_246),
.A2(n_234),
.B(n_243),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_260),
.B(n_261),
.C(n_263),
.Y(n_264)
);

OAI21xp5_ASAP7_75t_L g263 ( 
.A1(n_257),
.A2(n_248),
.B(n_252),
.Y(n_263)
);

OAI21xp5_ASAP7_75t_L g265 ( 
.A1(n_262),
.A2(n_254),
.B(n_258),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_265),
.Y(n_266)
);

AOI21xp5_ASAP7_75t_L g267 ( 
.A1(n_264),
.A2(n_12),
.B(n_14),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_267),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_L g269 ( 
.A(n_268),
.B(n_266),
.Y(n_269)
);


endmodule