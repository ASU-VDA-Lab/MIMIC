module fake_aes_4986_n_45 (n_11, n_1, n_2, n_13, n_12, n_6, n_4, n_3, n_9, n_5, n_14, n_7, n_15, n_10, n_8, n_0, n_45);
input n_11;
input n_1;
input n_2;
input n_13;
input n_12;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_14;
input n_7;
input n_15;
input n_10;
input n_8;
input n_0;
output n_45;
wire n_20;
wire n_38;
wire n_44;
wire n_36;
wire n_37;
wire n_34;
wire n_23;
wire n_28;
wire n_31;
wire n_22;
wire n_25;
wire n_16;
wire n_26;
wire n_30;
wire n_33;
wire n_18;
wire n_32;
wire n_41;
wire n_35;
wire n_17;
wire n_42;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_43;
wire n_40;
wire n_27;
wire n_39;
OAI22xp5_ASAP7_75t_L g16 ( .A1(n_10), .A2(n_12), .B1(n_2), .B2(n_8), .Y(n_16) );
BUFx6f_ASAP7_75t_L g17 ( .A(n_5), .Y(n_17) );
NOR2xp33_ASAP7_75t_L g18 ( .A(n_11), .B(n_13), .Y(n_18) );
HB1xp67_ASAP7_75t_L g19 ( .A(n_0), .Y(n_19) );
AND2x4_ASAP7_75t_L g20 ( .A(n_15), .B(n_2), .Y(n_20) );
NAND2xp5_ASAP7_75t_L g21 ( .A(n_7), .B(n_9), .Y(n_21) );
NOR2xp33_ASAP7_75t_SL g22 ( .A(n_5), .B(n_3), .Y(n_22) );
AOI21xp5_ASAP7_75t_L g23 ( .A1(n_21), .A2(n_14), .B(n_1), .Y(n_23) );
INVx5_ASAP7_75t_L g24 ( .A(n_20), .Y(n_24) );
NAND2xp5_ASAP7_75t_L g25 ( .A(n_19), .B(n_0), .Y(n_25) );
AND2x2_ASAP7_75t_L g26 ( .A(n_20), .B(n_1), .Y(n_26) );
AO21x2_ASAP7_75t_L g27 ( .A1(n_23), .A2(n_16), .B(n_18), .Y(n_27) );
BUFx2_ASAP7_75t_L g28 ( .A(n_25), .Y(n_28) );
NAND2xp5_ASAP7_75t_L g29 ( .A(n_28), .B(n_26), .Y(n_29) );
BUFx3_ASAP7_75t_L g30 ( .A(n_27), .Y(n_30) );
AND2x2_ASAP7_75t_L g31 ( .A(n_29), .B(n_25), .Y(n_31) );
INVx1_ASAP7_75t_L g32 ( .A(n_30), .Y(n_32) );
NAND2xp5_ASAP7_75t_L g33 ( .A(n_31), .B(n_30), .Y(n_33) );
NAND2xp5_ASAP7_75t_L g34 ( .A(n_31), .B(n_27), .Y(n_34) );
AOI222xp33_ASAP7_75t_L g35 ( .A1(n_34), .A2(n_22), .B1(n_24), .B2(n_17), .C1(n_32), .C2(n_3), .Y(n_35) );
AOI31xp33_ASAP7_75t_L g36 ( .A1(n_33), .A2(n_32), .A3(n_22), .B(n_6), .Y(n_36) );
OAI211xp5_ASAP7_75t_L g37 ( .A1(n_34), .A2(n_24), .B(n_17), .C(n_6), .Y(n_37) );
INVx1_ASAP7_75t_L g38 ( .A(n_36), .Y(n_38) );
NAND2xp5_ASAP7_75t_L g39 ( .A(n_35), .B(n_36), .Y(n_39) );
INVx1_ASAP7_75t_L g40 ( .A(n_37), .Y(n_40) );
INVx1_ASAP7_75t_L g41 ( .A(n_38), .Y(n_41) );
AND2x2_ASAP7_75t_L g42 ( .A(n_40), .B(n_17), .Y(n_42) );
BUFx2_ASAP7_75t_L g43 ( .A(n_39), .Y(n_43) );
INVx2_ASAP7_75t_L g44 ( .A(n_41), .Y(n_44) );
AOI22x1_ASAP7_75t_L g45 ( .A1(n_44), .A2(n_43), .B1(n_42), .B2(n_4), .Y(n_45) );
endmodule