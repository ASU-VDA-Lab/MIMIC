module fake_jpeg_16751_n_267 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_267);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_267;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_127;
wire n_76;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_91;
wire n_54;
wire n_33;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_258;
wire n_96;

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_2),
.Y(n_15)
);

INVx11_ASAP7_75t_L g16 ( 
.A(n_14),
.Y(n_16)
);

BUFx16f_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

BUFx12_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

BUFx12_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_8),
.Y(n_22)
);

CKINVDCx16_ASAP7_75t_R g23 ( 
.A(n_3),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_12),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_12),
.Y(n_28)
);

INVx11_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_10),
.Y(n_33)
);

BUFx10_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_1),
.Y(n_35)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_14),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_6),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_13),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_37),
.Y(n_39)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_39),
.Y(n_64)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_31),
.Y(n_40)
);

INVx3_ASAP7_75t_SL g76 ( 
.A(n_40),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_24),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_41),
.Y(n_68)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_31),
.Y(n_42)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_42),
.Y(n_73)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_34),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_43),
.B(n_47),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_24),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_44),
.Y(n_80)
);

BUFx4f_ASAP7_75t_SL g45 ( 
.A(n_34),
.Y(n_45)
);

INVx5_ASAP7_75t_SL g93 ( 
.A(n_45),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_22),
.B(n_11),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_SL g67 ( 
.A(n_46),
.B(n_54),
.Y(n_67)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_31),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_34),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_21),
.Y(n_49)
);

INVx5_ASAP7_75t_L g74 ( 
.A(n_49),
.Y(n_74)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_50),
.Y(n_95)
);

CKINVDCx16_ASAP7_75t_R g51 ( 
.A(n_17),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_51),
.B(n_57),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_24),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_52),
.Y(n_98)
);

CKINVDCx9p33_ASAP7_75t_R g53 ( 
.A(n_17),
.Y(n_53)
);

BUFx2_ASAP7_75t_L g78 ( 
.A(n_53),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_22),
.B(n_11),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_19),
.B(n_0),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_55),
.B(n_27),
.Y(n_71)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_37),
.Y(n_56)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_56),
.Y(n_70)
);

CKINVDCx16_ASAP7_75t_R g57 ( 
.A(n_17),
.Y(n_57)
);

INVx5_ASAP7_75t_L g58 ( 
.A(n_31),
.Y(n_58)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_58),
.Y(n_81)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_31),
.Y(n_59)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_59),
.Y(n_83)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_21),
.Y(n_60)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_60),
.Y(n_82)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_31),
.Y(n_61)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_61),
.Y(n_88)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_34),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_62),
.B(n_30),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_50),
.A2(n_16),
.B1(n_29),
.B2(n_36),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_63),
.A2(n_75),
.B1(n_30),
.B2(n_20),
.Y(n_129)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_49),
.Y(n_65)
);

INVx5_ASAP7_75t_L g120 ( 
.A(n_65),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g66 ( 
.A(n_45),
.B(n_34),
.C(n_30),
.Y(n_66)
);

AND2x2_ASAP7_75t_L g124 ( 
.A(n_66),
.B(n_0),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_SL g112 ( 
.A(n_71),
.B(n_79),
.Y(n_112)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_49),
.Y(n_72)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_72),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_39),
.A2(n_16),
.B1(n_29),
.B2(n_36),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_L g77 ( 
.A1(n_56),
.A2(n_36),
.B1(n_16),
.B2(n_29),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_77),
.A2(n_100),
.B1(n_23),
.B2(n_35),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_45),
.B(n_19),
.Y(n_79)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_60),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_84),
.B(n_89),
.Y(n_113)
);

INVx6_ASAP7_75t_L g85 ( 
.A(n_60),
.Y(n_85)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_85),
.Y(n_136)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_59),
.Y(n_86)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_86),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_61),
.B(n_19),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_SL g123 ( 
.A(n_87),
.B(n_90),
.Y(n_123)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_53),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_41),
.B(n_27),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_44),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_91),
.B(n_96),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_52),
.B(n_27),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_SL g131 ( 
.A(n_94),
.B(n_99),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_40),
.Y(n_96)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_58),
.Y(n_97)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_97),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_62),
.B(n_38),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_L g100 ( 
.A1(n_43),
.A2(n_17),
.B1(n_21),
.B2(n_24),
.Y(n_100)
);

INVx6_ASAP7_75t_L g101 ( 
.A(n_48),
.Y(n_101)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_101),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_50),
.A2(n_38),
.B1(n_25),
.B2(n_33),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_102),
.A2(n_6),
.B1(n_9),
.B2(n_7),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_55),
.B(n_33),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_103),
.B(n_28),
.Y(n_110)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_104),
.Y(n_122)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_83),
.Y(n_105)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_105),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_L g156 ( 
.A1(n_106),
.A2(n_129),
.B1(n_72),
.B2(n_85),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_64),
.B(n_21),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_107),
.B(n_115),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_73),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_SL g166 ( 
.A(n_110),
.B(n_20),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_L g114 ( 
.A1(n_95),
.A2(n_23),
.B1(n_28),
.B2(n_35),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_114),
.A2(n_117),
.B1(n_100),
.B2(n_89),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_69),
.B(n_26),
.Y(n_115)
);

OAI22xp33_ASAP7_75t_L g117 ( 
.A1(n_70),
.A2(n_15),
.B1(n_26),
.B2(n_32),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_88),
.B(n_26),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_119),
.B(n_126),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_74),
.A2(n_15),
.B1(n_7),
.B2(n_9),
.Y(n_121)
);

AOI21xp5_ASAP7_75t_L g167 ( 
.A1(n_121),
.A2(n_124),
.B(n_130),
.Y(n_167)
);

INVxp67_ASAP7_75t_L g125 ( 
.A(n_92),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_86),
.B(n_0),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_127),
.A2(n_132),
.B1(n_141),
.B2(n_65),
.Y(n_168)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_81),
.Y(n_128)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_128),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_74),
.A2(n_9),
.B1(n_7),
.B2(n_32),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_75),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_132)
);

AOI32xp33_ASAP7_75t_L g133 ( 
.A1(n_101),
.A2(n_32),
.A3(n_20),
.B1(n_18),
.B2(n_5),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_133),
.B(n_134),
.Y(n_153)
);

HB1xp67_ASAP7_75t_L g134 ( 
.A(n_78),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_63),
.A2(n_20),
.B1(n_18),
.B2(n_4),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_135),
.A2(n_4),
.B1(n_5),
.B2(n_82),
.Y(n_169)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_81),
.Y(n_137)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_137),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_76),
.B(n_1),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_138),
.B(n_143),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_78),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_139),
.B(n_140),
.Y(n_154)
);

INVx1_ASAP7_75t_SL g140 ( 
.A(n_68),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_77),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_76),
.B(n_3),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_L g199 ( 
.A1(n_145),
.A2(n_156),
.B1(n_168),
.B2(n_120),
.Y(n_199)
);

INVx8_ASAP7_75t_L g146 ( 
.A(n_105),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_146),
.B(n_166),
.Y(n_193)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_142),
.Y(n_150)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_150),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_123),
.B(n_131),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_SL g182 ( 
.A(n_151),
.B(n_162),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_108),
.B(n_67),
.Y(n_157)
);

INVxp67_ASAP7_75t_L g186 ( 
.A(n_157),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_123),
.B(n_131),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_158),
.B(n_161),
.Y(n_178)
);

AO22x1_ASAP7_75t_L g159 ( 
.A1(n_132),
.A2(n_84),
.B1(n_82),
.B2(n_93),
.Y(n_159)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_159),
.Y(n_177)
);

INVx3_ASAP7_75t_L g160 ( 
.A(n_109),
.Y(n_160)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_160),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_112),
.B(n_98),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_112),
.B(n_97),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_126),
.B(n_68),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_163),
.B(n_149),
.Y(n_180)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_107),
.Y(n_164)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_164),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_119),
.B(n_93),
.C(n_98),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_165),
.B(n_118),
.C(n_137),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_169),
.A2(n_173),
.B1(n_167),
.B2(n_162),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_116),
.B(n_18),
.Y(n_170)
);

INVxp67_ASAP7_75t_L g201 ( 
.A(n_170),
.Y(n_201)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_142),
.Y(n_171)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_171),
.Y(n_185)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_111),
.Y(n_172)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_172),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_124),
.A2(n_80),
.B1(n_5),
.B2(n_18),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_111),
.Y(n_174)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_174),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_141),
.A2(n_80),
.B1(n_18),
.B2(n_5),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_175),
.A2(n_143),
.B1(n_138),
.B2(n_127),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_158),
.B(n_115),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_176),
.B(n_180),
.Y(n_210)
);

AOI221xp5_ASAP7_75t_L g205 ( 
.A1(n_181),
.A2(n_187),
.B1(n_168),
.B2(n_175),
.C(n_155),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_147),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_183),
.B(n_203),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_149),
.B(n_124),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_189),
.B(n_192),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_144),
.B(n_122),
.Y(n_192)
);

A2O1A1Ixp33_ASAP7_75t_L g194 ( 
.A1(n_153),
.A2(n_125),
.B(n_122),
.C(n_106),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_SL g220 ( 
.A(n_194),
.B(n_198),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_163),
.B(n_128),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_144),
.B(n_118),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_197),
.B(n_173),
.C(n_148),
.Y(n_212)
);

AOI21x1_ASAP7_75t_L g198 ( 
.A1(n_164),
.A2(n_117),
.B(n_140),
.Y(n_198)
);

INVxp67_ASAP7_75t_L g206 ( 
.A(n_199),
.Y(n_206)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_172),
.Y(n_200)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_200),
.Y(n_207)
);

INVx3_ASAP7_75t_L g202 ( 
.A(n_160),
.Y(n_202)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_202),
.Y(n_213)
);

INVxp67_ASAP7_75t_L g203 ( 
.A(n_150),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g204 ( 
.A(n_151),
.B(n_113),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_204),
.B(n_166),
.Y(n_216)
);

AOI322xp5_ASAP7_75t_L g234 ( 
.A1(n_205),
.A2(n_201),
.A3(n_200),
.B1(n_191),
.B2(n_186),
.C1(n_184),
.C2(n_183),
.Y(n_234)
);

AOI21xp33_ASAP7_75t_L g208 ( 
.A1(n_178),
.A2(n_161),
.B(n_155),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_L g209 ( 
.A1(n_177),
.A2(n_169),
.B1(n_165),
.B2(n_167),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_L g237 ( 
.A1(n_209),
.A2(n_214),
.B1(n_215),
.B2(n_220),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_212),
.B(n_217),
.C(n_219),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_L g214 ( 
.A1(n_177),
.A2(n_159),
.B1(n_120),
.B2(n_146),
.Y(n_214)
);

AOI21xp5_ASAP7_75t_L g215 ( 
.A1(n_198),
.A2(n_152),
.B(n_148),
.Y(n_215)
);

INVxp67_ASAP7_75t_L g227 ( 
.A(n_215),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_216),
.B(n_176),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_197),
.B(n_152),
.C(n_174),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_178),
.B(n_159),
.Y(n_218)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_218),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_180),
.B(n_145),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_189),
.B(n_154),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_221),
.B(n_193),
.C(n_204),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_SL g223 ( 
.A(n_182),
.B(n_147),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_SL g225 ( 
.A(n_223),
.B(n_182),
.Y(n_225)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_190),
.Y(n_224)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_224),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_225),
.B(n_226),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_206),
.A2(n_188),
.B1(n_196),
.B2(n_195),
.Y(n_228)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_228),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_230),
.B(n_232),
.C(n_212),
.Y(n_239)
);

XOR2xp5_ASAP7_75t_L g232 ( 
.A(n_217),
.B(n_187),
.Y(n_232)
);

MAJx2_ASAP7_75t_L g233 ( 
.A(n_220),
.B(n_194),
.C(n_181),
.Y(n_233)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_233),
.B(n_219),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_234),
.B(n_237),
.Y(n_247)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_222),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_207),
.A2(n_136),
.B1(n_179),
.B2(n_185),
.Y(n_238)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_239),
.B(n_241),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_229),
.B(n_221),
.C(n_210),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_229),
.B(n_210),
.C(n_211),
.Y(n_242)
);

OAI21xp5_ASAP7_75t_L g250 ( 
.A1(n_242),
.A2(n_244),
.B(n_246),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_SL g252 ( 
.A(n_243),
.B(n_233),
.Y(n_252)
);

AOI21xp5_ASAP7_75t_L g244 ( 
.A1(n_227),
.A2(n_218),
.B(n_214),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_232),
.B(n_230),
.C(n_231),
.Y(n_246)
);

AOI22xp33_ASAP7_75t_SL g248 ( 
.A1(n_244),
.A2(n_235),
.B1(n_236),
.B2(n_213),
.Y(n_248)
);

INVx11_ASAP7_75t_L g254 ( 
.A(n_248),
.Y(n_254)
);

AOI21xp5_ASAP7_75t_SL g249 ( 
.A1(n_245),
.A2(n_231),
.B(n_227),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_SL g251 ( 
.A(n_240),
.B(n_228),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_251),
.B(n_247),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_252),
.B(n_239),
.C(n_246),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_255),
.B(n_258),
.Y(n_260)
);

OAI21x1_ASAP7_75t_L g256 ( 
.A1(n_248),
.A2(n_250),
.B(n_249),
.Y(n_256)
);

AOI31xp67_ASAP7_75t_SL g259 ( 
.A1(n_256),
.A2(n_208),
.A3(n_252),
.B(n_243),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_257),
.B(n_253),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_253),
.B(n_238),
.Y(n_258)
);

INVxp67_ASAP7_75t_L g264 ( 
.A(n_259),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_261),
.B(n_262),
.C(n_257),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_258),
.B(n_241),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_263),
.B(n_261),
.C(n_260),
.Y(n_265)
);

OAI21x1_ASAP7_75t_SL g266 ( 
.A1(n_265),
.A2(n_264),
.B(n_254),
.Y(n_266)
);

XOR2xp5_ASAP7_75t_L g267 ( 
.A(n_266),
.B(n_254),
.Y(n_267)
);


endmodule