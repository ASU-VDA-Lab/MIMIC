module fake_jpeg_29348_n_63 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_7, n_63);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;
input n_7;

output n_63;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_23;
wire n_10;
wire n_27;
wire n_55;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_59;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_62;
wire n_25;
wire n_17;
wire n_31;
wire n_56;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_8;
wire n_15;

CKINVDCx20_ASAP7_75t_R g8 ( 
.A(n_6),
.Y(n_8)
);

INVx1_ASAP7_75t_L g9 ( 
.A(n_4),
.Y(n_9)
);

BUFx6f_ASAP7_75t_L g10 ( 
.A(n_6),
.Y(n_10)
);

INVx6_ASAP7_75t_L g11 ( 
.A(n_0),
.Y(n_11)
);

BUFx6f_ASAP7_75t_L g12 ( 
.A(n_0),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_0),
.Y(n_13)
);

BUFx12f_ASAP7_75t_L g14 ( 
.A(n_1),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_2),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_5),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_18),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_13),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_19),
.B(n_21),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_20),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_12),
.B(n_1),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_12),
.B(n_1),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_22),
.B(n_23),
.Y(n_27)
);

INVx8_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_L g24 ( 
.A1(n_21),
.A2(n_10),
.B1(n_15),
.B2(n_13),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_L g40 ( 
.A1(n_24),
.A2(n_8),
.B1(n_16),
.B2(n_9),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_19),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_SL g35 ( 
.A(n_25),
.B(n_30),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_SL g30 ( 
.A(n_22),
.B(n_17),
.Y(n_30)
);

OAI22xp33_ASAP7_75t_L g31 ( 
.A1(n_29),
.A2(n_20),
.B1(n_18),
.B2(n_23),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_L g43 ( 
.A1(n_31),
.A2(n_38),
.B1(n_40),
.B2(n_9),
.Y(n_43)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_28),
.Y(n_32)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_32),
.Y(n_41)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_29),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_33),
.B(n_36),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_26),
.B(n_15),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_34),
.B(n_5),
.Y(n_46)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_25),
.Y(n_36)
);

OA21x2_ASAP7_75t_L g37 ( 
.A1(n_27),
.A2(n_23),
.B(n_20),
.Y(n_37)
);

OA22x2_ASAP7_75t_L g45 ( 
.A1(n_37),
.A2(n_14),
.B1(n_8),
.B2(n_3),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_SL g38 ( 
.A1(n_28),
.A2(n_20),
.B1(n_14),
.B2(n_16),
.Y(n_38)
);

CKINVDCx16_ASAP7_75t_R g39 ( 
.A(n_28),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_39),
.B(n_14),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_43),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_SL g50 ( 
.A(n_44),
.B(n_46),
.Y(n_50)
);

MAJIxp5_ASAP7_75t_L g49 ( 
.A(n_45),
.B(n_47),
.C(n_40),
.Y(n_49)
);

AOI21xp5_ASAP7_75t_SL g47 ( 
.A1(n_34),
.A2(n_14),
.B(n_3),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_49),
.B(n_47),
.Y(n_53)
);

MAJIxp5_ASAP7_75t_L g51 ( 
.A(n_42),
.B(n_35),
.C(n_38),
.Y(n_51)
);

XNOR2xp5_ASAP7_75t_L g54 ( 
.A(n_51),
.B(n_46),
.Y(n_54)
);

INVxp33_ASAP7_75t_L g52 ( 
.A(n_50),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g55 ( 
.A1(n_52),
.A2(n_48),
.B1(n_45),
.B2(n_37),
.Y(n_55)
);

MAJIxp5_ASAP7_75t_L g56 ( 
.A(n_53),
.B(n_54),
.C(n_45),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_55),
.A2(n_52),
.B1(n_37),
.B2(n_41),
.Y(n_57)
);

MAJIxp5_ASAP7_75t_L g58 ( 
.A(n_56),
.B(n_41),
.C(n_32),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_57),
.B(n_58),
.Y(n_60)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_58),
.Y(n_59)
);

BUFx24_ASAP7_75t_SL g61 ( 
.A(n_59),
.Y(n_61)
);

AOI322xp5_ASAP7_75t_L g62 ( 
.A1(n_61),
.A2(n_2),
.A3(n_3),
.B1(n_7),
.B2(n_31),
.C1(n_60),
.C2(n_53),
.Y(n_62)
);

XNOR2xp5_ASAP7_75t_L g63 ( 
.A(n_62),
.B(n_7),
.Y(n_63)
);


endmodule