module fake_jpeg_23280_n_306 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_306);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_306;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_252;
wire n_273;
wire n_251;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_207;
wire n_155;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_301;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_298;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_303;
wire n_304;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_299;
wire n_294;
wire n_211;
wire n_300;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_302;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_305;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_297;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_256;
wire n_151;
wire n_221;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_181;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

BUFx4f_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_4),
.Y(n_20)
);

BUFx10_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_17),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_5),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_16),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_6),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_17),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

BUFx4f_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_8),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_6),
.Y(n_33)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_10),
.Y(n_34)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_9),
.Y(n_35)
);

BUFx16f_ASAP7_75t_L g36 ( 
.A(n_6),
.Y(n_36)
);

INVx6_ASAP7_75t_SL g37 ( 
.A(n_17),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_11),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_18),
.B(n_0),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_39),
.B(n_49),
.Y(n_53)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_19),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_40),
.B(n_41),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_26),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_19),
.Y(n_42)
);

INVx5_ASAP7_75t_L g63 ( 
.A(n_42),
.Y(n_63)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_31),
.Y(n_43)
);

BUFx4f_ASAP7_75t_L g66 ( 
.A(n_43),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_19),
.Y(n_44)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_44),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_26),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_45),
.B(n_48),
.Y(n_74)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_31),
.Y(n_46)
);

INVx5_ASAP7_75t_L g76 ( 
.A(n_46),
.Y(n_76)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_19),
.Y(n_47)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_47),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_SL g48 ( 
.A(n_20),
.B(n_24),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_31),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_39),
.A2(n_38),
.B1(n_22),
.B2(n_29),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_50),
.A2(n_71),
.B1(n_77),
.B2(n_36),
.Y(n_108)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_48),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_52),
.B(n_54),
.Y(n_81)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_48),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_L g55 ( 
.A1(n_41),
.A2(n_31),
.B1(n_23),
.B2(n_34),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_55),
.A2(n_68),
.B1(n_47),
.B2(n_45),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_39),
.B(n_30),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_56),
.B(n_57),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_39),
.B(n_30),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_42),
.Y(n_58)
);

INVx8_ASAP7_75t_L g83 ( 
.A(n_58),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_43),
.A2(n_38),
.B1(n_29),
.B2(n_22),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_59),
.A2(n_67),
.B1(n_44),
.B2(n_25),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_40),
.B(n_23),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_60),
.B(n_44),
.Y(n_90)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_42),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_61),
.B(n_72),
.Y(n_85)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_42),
.Y(n_62)
);

INVx6_ASAP7_75t_L g105 ( 
.A(n_62),
.Y(n_105)
);

A2O1A1Ixp33_ASAP7_75t_L g64 ( 
.A1(n_41),
.A2(n_21),
.B(n_37),
.C(n_25),
.Y(n_64)
);

A2O1A1Ixp33_ASAP7_75t_L g96 ( 
.A1(n_64),
.A2(n_69),
.B(n_21),
.C(n_33),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_43),
.A2(n_32),
.B1(n_35),
.B2(n_34),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g68 ( 
.A1(n_43),
.A2(n_46),
.B1(n_49),
.B2(n_40),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_46),
.A2(n_37),
.B1(n_35),
.B2(n_32),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_46),
.A2(n_28),
.B1(n_20),
.B2(n_24),
.Y(n_71)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_42),
.Y(n_72)
);

OAI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_49),
.A2(n_40),
.B1(n_47),
.B2(n_41),
.Y(n_73)
);

OAI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_73),
.A2(n_33),
.B1(n_27),
.B2(n_18),
.Y(n_102)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_47),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_75),
.B(n_78),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_49),
.A2(n_28),
.B1(n_27),
.B2(n_18),
.Y(n_77)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_47),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_60),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_79),
.B(n_87),
.Y(n_129)
);

OAI22xp33_ASAP7_75t_SL g145 ( 
.A1(n_80),
.A2(n_96),
.B1(n_102),
.B2(n_106),
.Y(n_145)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_66),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_82),
.B(n_91),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_L g84 ( 
.A1(n_53),
.A2(n_45),
.B(n_44),
.Y(n_84)
);

OAI21xp5_ASAP7_75t_L g123 ( 
.A1(n_84),
.A2(n_88),
.B(n_65),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_86),
.A2(n_9),
.B1(n_14),
.B2(n_13),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_70),
.Y(n_87)
);

NAND2xp33_ASAP7_75t_SL g88 ( 
.A(n_69),
.B(n_21),
.Y(n_88)
);

AND2x2_ASAP7_75t_L g133 ( 
.A(n_90),
.B(n_1),
.Y(n_133)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_66),
.Y(n_91)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_70),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_92),
.B(n_108),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_76),
.A2(n_25),
.B1(n_13),
.B2(n_16),
.Y(n_93)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_93),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_66),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_95),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_52),
.B(n_45),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g124 ( 
.A(n_97),
.B(n_112),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_66),
.Y(n_98)
);

CKINVDCx16_ASAP7_75t_R g119 ( 
.A(n_98),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_56),
.B(n_21),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_99),
.B(n_116),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_53),
.B(n_44),
.C(n_21),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_100),
.B(n_1),
.C(n_2),
.Y(n_138)
);

INVx8_ASAP7_75t_L g101 ( 
.A(n_58),
.Y(n_101)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_101),
.Y(n_127)
);

INVx13_ASAP7_75t_L g103 ( 
.A(n_58),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_103),
.B(n_104),
.Y(n_128)
);

CKINVDCx5p33_ASAP7_75t_R g104 ( 
.A(n_74),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_L g106 ( 
.A1(n_76),
.A2(n_50),
.B1(n_54),
.B2(n_65),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_64),
.A2(n_33),
.B1(n_27),
.B2(n_36),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_107),
.A2(n_77),
.B1(n_65),
.B2(n_63),
.Y(n_118)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_71),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_109),
.B(n_110),
.Y(n_136)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_68),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_74),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_111),
.B(n_115),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_57),
.B(n_36),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_61),
.B(n_0),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_SL g142 ( 
.A(n_113),
.B(n_114),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_51),
.B(n_0),
.Y(n_114)
);

INVx13_ASAP7_75t_L g115 ( 
.A(n_62),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_72),
.B(n_16),
.Y(n_116)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_105),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_117),
.B(n_137),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_118),
.A2(n_139),
.B1(n_92),
.B2(n_113),
.Y(n_158)
);

AND2x4_ASAP7_75t_L g122 ( 
.A(n_84),
.B(n_63),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_SL g168 ( 
.A1(n_122),
.A2(n_134),
.B(n_94),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_L g153 ( 
.A(n_123),
.B(n_80),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_89),
.B(n_51),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_126),
.B(n_131),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_89),
.B(n_0),
.Y(n_131)
);

INVx1_ASAP7_75t_SL g132 ( 
.A(n_116),
.Y(n_132)
);

INVx1_ASAP7_75t_SL g160 ( 
.A(n_132),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_133),
.B(n_141),
.Y(n_169)
);

AND2x2_ASAP7_75t_L g134 ( 
.A(n_90),
.B(n_1),
.Y(n_134)
);

A2O1A1Ixp33_ASAP7_75t_SL g135 ( 
.A1(n_107),
.A2(n_78),
.B(n_75),
.C(n_3),
.Y(n_135)
);

AOI21xp5_ASAP7_75t_L g161 ( 
.A1(n_135),
.A2(n_91),
.B(n_82),
.Y(n_161)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_85),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_138),
.B(n_144),
.C(n_148),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_110),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_139)
);

OR2x2_ASAP7_75t_L g141 ( 
.A(n_81),
.B(n_2),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_100),
.B(n_99),
.C(n_112),
.Y(n_144)
);

AND2x6_ASAP7_75t_L g146 ( 
.A(n_104),
.B(n_9),
.Y(n_146)
);

AOI221xp5_ASAP7_75t_L g178 ( 
.A1(n_146),
.A2(n_14),
.B1(n_15),
.B2(n_12),
.C(n_11),
.Y(n_178)
);

INVxp67_ASAP7_75t_L g163 ( 
.A(n_147),
.Y(n_163)
);

XOR2xp5_ASAP7_75t_L g148 ( 
.A(n_108),
.B(n_81),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_79),
.B(n_3),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_149),
.B(n_98),
.Y(n_175)
);

AND2x2_ASAP7_75t_SL g150 ( 
.A(n_122),
.B(n_87),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_150),
.B(n_138),
.C(n_120),
.Y(n_188)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_125),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_151),
.B(n_156),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_SL g152 ( 
.A(n_124),
.B(n_111),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_SL g186 ( 
.A(n_152),
.B(n_181),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g194 ( 
.A(n_153),
.B(n_168),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_122),
.A2(n_109),
.B1(n_96),
.B2(n_88),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_154),
.A2(n_173),
.B1(n_121),
.B2(n_120),
.Y(n_183)
);

CKINVDCx16_ASAP7_75t_R g156 ( 
.A(n_143),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_126),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_157),
.B(n_159),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_158),
.A2(n_172),
.B1(n_135),
.B2(n_132),
.Y(n_196)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_136),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_161),
.B(n_162),
.Y(n_190)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_129),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_149),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_164),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_128),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_165),
.B(n_166),
.Y(n_202)
);

BUFx2_ASAP7_75t_L g166 ( 
.A(n_140),
.Y(n_166)
);

OAI32xp33_ASAP7_75t_L g167 ( 
.A1(n_122),
.A2(n_114),
.A3(n_94),
.B1(n_85),
.B2(n_97),
.Y(n_167)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_167),
.B(n_177),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_137),
.B(n_115),
.Y(n_171)
);

CKINVDCx14_ASAP7_75t_R g189 ( 
.A(n_171),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_122),
.A2(n_118),
.B1(n_130),
.B2(n_145),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_148),
.A2(n_105),
.B1(n_115),
.B2(n_101),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_139),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_174),
.B(n_176),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_175),
.B(n_134),
.Y(n_192)
);

CKINVDCx16_ASAP7_75t_R g176 ( 
.A(n_140),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_SL g177 ( 
.A1(n_123),
.A2(n_98),
.B(n_95),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_178),
.A2(n_121),
.B1(n_131),
.B2(n_146),
.Y(n_187)
);

INVx3_ASAP7_75t_L g180 ( 
.A(n_117),
.Y(n_180)
);

BUFx6f_ASAP7_75t_L g204 ( 
.A(n_180),
.Y(n_204)
);

CKINVDCx14_ASAP7_75t_R g181 ( 
.A(n_142),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_183),
.A2(n_163),
.B1(n_168),
.B2(n_157),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_SL g184 ( 
.A(n_154),
.B(n_144),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_184),
.B(n_203),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_187),
.B(n_193),
.Y(n_218)
);

OAI21xp5_ASAP7_75t_SL g232 ( 
.A1(n_188),
.A2(n_119),
.B(n_176),
.Y(n_232)
);

NOR2x1_ASAP7_75t_L g191 ( 
.A(n_150),
.B(n_141),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_191),
.B(n_192),
.Y(n_213)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_170),
.Y(n_193)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_170),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_195),
.B(n_207),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_L g228 ( 
.A1(n_196),
.A2(n_197),
.B1(n_198),
.B2(n_205),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_172),
.A2(n_135),
.B1(n_124),
.B2(n_142),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_174),
.A2(n_135),
.B1(n_105),
.B2(n_134),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_L g201 ( 
.A(n_179),
.B(n_153),
.Y(n_201)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_201),
.B(n_160),
.Y(n_229)
);

AOI322xp5_ASAP7_75t_L g203 ( 
.A1(n_179),
.A2(n_133),
.A3(n_135),
.B1(n_147),
.B2(n_141),
.C1(n_101),
.C2(n_83),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_158),
.A2(n_133),
.B1(n_83),
.B2(n_127),
.Y(n_205)
);

INVxp33_ASAP7_75t_L g207 ( 
.A(n_171),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_175),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_208),
.B(n_155),
.Y(n_223)
);

BUFx6f_ASAP7_75t_L g209 ( 
.A(n_166),
.Y(n_209)
);

INVx4_ASAP7_75t_L g216 ( 
.A(n_209),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_L g249 ( 
.A1(n_210),
.A2(n_214),
.B1(n_226),
.B2(n_227),
.Y(n_249)
);

AOI21xp5_ASAP7_75t_SL g211 ( 
.A1(n_191),
.A2(n_177),
.B(n_150),
.Y(n_211)
);

OAI21xp5_ASAP7_75t_L g234 ( 
.A1(n_211),
.A2(n_223),
.B(n_225),
.Y(n_234)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_206),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_212),
.B(n_215),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_183),
.A2(n_161),
.B1(n_150),
.B2(n_152),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_202),
.Y(n_215)
);

AND2x2_ASAP7_75t_L g217 ( 
.A(n_199),
.B(n_169),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_217),
.A2(n_219),
.B1(n_224),
.B2(n_192),
.Y(n_235)
);

AND2x2_ASAP7_75t_L g219 ( 
.A(n_199),
.B(n_169),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_184),
.B(n_155),
.C(n_173),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_220),
.B(n_229),
.C(n_230),
.Y(n_242)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_185),
.Y(n_224)
);

OAI21xp5_ASAP7_75t_L g225 ( 
.A1(n_190),
.A2(n_160),
.B(n_167),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_182),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_208),
.A2(n_165),
.B1(n_162),
.B2(n_159),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_201),
.B(n_164),
.C(n_151),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_196),
.A2(n_156),
.B1(n_127),
.B2(n_180),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_231),
.A2(n_193),
.B1(n_195),
.B2(n_189),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_232),
.B(n_188),
.C(n_198),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_233),
.B(n_238),
.Y(n_259)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_235),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_220),
.B(n_194),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_L g258 ( 
.A(n_236),
.B(n_240),
.Y(n_258)
);

NOR3xp33_ASAP7_75t_SL g238 ( 
.A(n_225),
.B(n_200),
.C(n_187),
.Y(n_238)
);

XOR2xp5_ASAP7_75t_L g239 ( 
.A(n_229),
.B(n_194),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_239),
.B(n_244),
.C(n_245),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_SL g240 ( 
.A(n_217),
.B(n_197),
.Y(n_240)
);

HB1xp67_ASAP7_75t_L g241 ( 
.A(n_216),
.Y(n_241)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_241),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_231),
.A2(n_186),
.B1(n_200),
.B2(n_205),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_243),
.A2(n_246),
.B1(n_222),
.B2(n_213),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_230),
.B(n_207),
.C(n_119),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_228),
.A2(n_83),
.B1(n_103),
.B2(n_204),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_SL g247 ( 
.A(n_217),
.B(n_219),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_247),
.B(n_248),
.C(n_210),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_232),
.B(n_204),
.C(n_209),
.Y(n_248)
);

XOR2x2_ASAP7_75t_SL g250 ( 
.A(n_218),
.B(n_12),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_250),
.B(n_219),
.Y(n_261)
);

AO22x1_ASAP7_75t_L g252 ( 
.A1(n_234),
.A2(n_211),
.B1(n_214),
.B2(n_213),
.Y(n_252)
);

OAI21xp5_ASAP7_75t_SL g269 ( 
.A1(n_252),
.A2(n_266),
.B(n_242),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_254),
.A2(n_262),
.B1(n_244),
.B2(n_240),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_L g272 ( 
.A(n_255),
.B(n_3),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_SL g256 ( 
.A(n_237),
.B(n_224),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_256),
.B(n_257),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_238),
.B(n_223),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_SL g260 ( 
.A(n_245),
.B(n_227),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_260),
.B(n_261),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_235),
.A2(n_215),
.B1(n_212),
.B2(n_216),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_242),
.B(n_221),
.C(n_166),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_264),
.B(n_4),
.C(n_5),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_SL g265 ( 
.A(n_249),
.B(n_248),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_265),
.B(n_11),
.Y(n_274)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_247),
.Y(n_266)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_268),
.Y(n_286)
);

OAI21xp5_ASAP7_75t_SL g280 ( 
.A1(n_269),
.A2(n_274),
.B(n_277),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_L g270 ( 
.A1(n_253),
.A2(n_250),
.B1(n_239),
.B2(n_103),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_270),
.B(n_271),
.C(n_272),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_L g271 ( 
.A1(n_259),
.A2(n_221),
.B1(n_140),
.B2(n_95),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_273),
.B(n_255),
.C(n_251),
.Y(n_284)
);

INVxp67_ASAP7_75t_L g275 ( 
.A(n_262),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_275),
.B(n_252),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_254),
.A2(n_5),
.B1(n_7),
.B2(n_8),
.Y(n_277)
);

OAI21xp5_ASAP7_75t_SL g278 ( 
.A1(n_252),
.A2(n_5),
.B(n_7),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_278),
.B(n_263),
.C(n_266),
.Y(n_285)
);

OR2x2_ASAP7_75t_L g292 ( 
.A(n_279),
.B(n_281),
.Y(n_292)
);

OR2x2_ASAP7_75t_L g281 ( 
.A(n_278),
.B(n_275),
.Y(n_281)
);

NOR3xp33_ASAP7_75t_SL g282 ( 
.A(n_267),
.B(n_257),
.C(n_258),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_282),
.B(n_268),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_SL g287 ( 
.A(n_284),
.B(n_272),
.Y(n_287)
);

OAI21xp5_ASAP7_75t_L g291 ( 
.A1(n_285),
.A2(n_276),
.B(n_273),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_287),
.B(n_288),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_279),
.B(n_277),
.Y(n_288)
);

XOR2xp5_ASAP7_75t_L g289 ( 
.A(n_283),
.B(n_269),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_289),
.B(n_286),
.Y(n_295)
);

AOI21xp5_ASAP7_75t_L g296 ( 
.A1(n_290),
.A2(n_291),
.B(n_293),
.Y(n_296)
);

AOI21x1_ASAP7_75t_L g293 ( 
.A1(n_280),
.A2(n_258),
.B(n_251),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_295),
.B(n_298),
.C(n_7),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_SL g297 ( 
.A1(n_292),
.A2(n_281),
.B1(n_263),
.B2(n_264),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_297),
.B(n_289),
.Y(n_299)
);

AOI21xp5_ASAP7_75t_L g298 ( 
.A1(n_292),
.A2(n_14),
.B(n_15),
.Y(n_298)
);

INVxp67_ASAP7_75t_L g303 ( 
.A(n_299),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_294),
.B(n_15),
.Y(n_300)
);

OAI21xp5_ASAP7_75t_L g302 ( 
.A1(n_300),
.A2(n_301),
.B(n_296),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_302),
.B(n_7),
.C(n_8),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_SL g305 ( 
.A(n_304),
.B(n_8),
.Y(n_305)
);

OR2x2_ASAP7_75t_L g306 ( 
.A(n_305),
.B(n_303),
.Y(n_306)
);


endmodule