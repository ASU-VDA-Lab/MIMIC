module real_jpeg_14848_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_146;
wire n_247;
wire n_78;
wire n_83;
wire n_249;
wire n_215;
wire n_166;
wire n_221;
wire n_176;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_243;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_200;
wire n_48;
wire n_164;
wire n_184;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_113;
wire n_155;
wire n_120;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_44;
wire n_28;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_211;
wire n_172;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_203;
wire n_192;
wire n_100;
wire n_198;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_205;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_241;
wire n_103;
wire n_225;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_185;
wire n_125;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_97;
wire n_75;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_216;
wire n_202;
wire n_128;
wire n_179;
wire n_167;
wire n_244;
wire n_133;
wire n_213;
wire n_138;
wire n_25;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;

BUFx2_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

BUFx4f_ASAP7_75t_L g41 ( 
.A(n_1),
.Y(n_41)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_2),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g30 ( 
.A1(n_3),
.A2(n_25),
.B1(n_31),
.B2(n_32),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_3),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_3),
.A2(n_31),
.B1(n_43),
.B2(n_44),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g67 ( 
.A1(n_4),
.A2(n_61),
.B1(n_62),
.B2(n_68),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_4),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_4),
.A2(n_56),
.B1(n_57),
.B2(n_68),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_4),
.A2(n_43),
.B1(n_44),
.B2(n_68),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_4),
.A2(n_25),
.B1(n_32),
.B2(n_68),
.Y(n_217)
);

O2A1O1Ixp33_ASAP7_75t_L g99 ( 
.A1(n_5),
.A2(n_55),
.B(n_61),
.C(n_100),
.Y(n_99)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_5),
.Y(n_101)
);

OAI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_5),
.A2(n_61),
.B1(n_62),
.B2(n_101),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_5),
.B(n_130),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_5),
.B(n_56),
.Y(n_186)
);

AOI21xp33_ASAP7_75t_SL g200 ( 
.A1(n_5),
.A2(n_56),
.B(n_186),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_5),
.B(n_25),
.C(n_39),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_L g211 ( 
.A1(n_5),
.A2(n_43),
.B1(n_44),
.B2(n_101),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_L g222 ( 
.A1(n_5),
.A2(n_24),
.B1(n_27),
.B2(n_223),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_5),
.B(n_79),
.Y(n_235)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_6),
.Y(n_44)
);

INVx11_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_8),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g42 ( 
.A1(n_9),
.A2(n_43),
.B1(n_44),
.B2(n_45),
.Y(n_42)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_9),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_9),
.A2(n_25),
.B1(n_32),
.B2(n_45),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_9),
.A2(n_45),
.B1(n_56),
.B2(n_57),
.Y(n_125)
);

BUFx12_ASAP7_75t_L g75 ( 
.A(n_10),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_11),
.A2(n_61),
.B1(n_62),
.B2(n_108),
.Y(n_107)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_11),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_L g162 ( 
.A1(n_11),
.A2(n_56),
.B1(n_57),
.B2(n_108),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g212 ( 
.A1(n_11),
.A2(n_43),
.B1(n_44),
.B2(n_108),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_11),
.A2(n_25),
.B1(n_32),
.B2(n_108),
.Y(n_223)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_12),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_13),
.A2(n_61),
.B1(n_62),
.B2(n_66),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_13),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_13),
.A2(n_56),
.B1(n_57),
.B2(n_66),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g202 ( 
.A1(n_13),
.A2(n_43),
.B1(n_44),
.B2(n_66),
.Y(n_202)
);

AOI22xp33_ASAP7_75t_L g215 ( 
.A1(n_13),
.A2(n_25),
.B1(n_32),
.B2(n_66),
.Y(n_215)
);

AOI22xp33_ASAP7_75t_L g70 ( 
.A1(n_14),
.A2(n_56),
.B1(n_57),
.B2(n_71),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_14),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_14),
.A2(n_25),
.B1(n_32),
.B2(n_71),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_14),
.A2(n_61),
.B1(n_62),
.B2(n_71),
.Y(n_131)
);

OAI22xp33_ASAP7_75t_SL g151 ( 
.A1(n_14),
.A2(n_43),
.B1(n_44),
.B2(n_71),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g35 ( 
.A1(n_15),
.A2(n_25),
.B1(n_32),
.B2(n_36),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_15),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_L g47 ( 
.A1(n_15),
.A2(n_36),
.B1(n_43),
.B2(n_44),
.Y(n_47)
);

OAI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_15),
.A2(n_36),
.B1(n_56),
.B2(n_57),
.Y(n_78)
);

XNOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_136),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_135),
.Y(n_17)
);

INVxp67_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_109),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_20),
.B(n_109),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_81),
.C(n_93),
.Y(n_20)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_21),
.B(n_81),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_50),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_22),
.B(n_51),
.C(n_80),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_37),
.Y(n_22)
);

XOR2xp5_ASAP7_75t_L g167 ( 
.A(n_23),
.B(n_37),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_29),
.B(n_33),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_24),
.B(n_35),
.Y(n_87)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_24),
.Y(n_96)
);

AOI21xp5_ASAP7_75t_L g113 ( 
.A1(n_24),
.A2(n_27),
.B(n_114),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g225 ( 
.A1(n_24),
.A2(n_27),
.B1(n_215),
.B2(n_223),
.Y(n_225)
);

OAI21xp5_ASAP7_75t_L g232 ( 
.A1(n_24),
.A2(n_85),
.B(n_217),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_27),
.Y(n_24)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_25),
.Y(n_32)
);

AOI22xp5_ASAP7_75t_L g38 ( 
.A1(n_25),
.A2(n_32),
.B1(n_39),
.B2(n_40),
.Y(n_38)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_27),
.B(n_35),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_SL g221 ( 
.A(n_27),
.B(n_101),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_28),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_28),
.B(n_86),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_28),
.A2(n_30),
.B1(n_96),
.B2(n_97),
.Y(n_95)
);

AOI21xp5_ASAP7_75t_L g158 ( 
.A1(n_28),
.A2(n_87),
.B(n_97),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_28),
.A2(n_96),
.B1(n_214),
.B2(n_216),
.Y(n_213)
);

CKINVDCx16_ASAP7_75t_R g29 ( 
.A(n_30),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_32),
.B(n_221),
.Y(n_220)
);

INVxp67_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

AOI21xp5_ASAP7_75t_L g189 ( 
.A1(n_34),
.A2(n_86),
.B(n_96),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_L g37 ( 
.A1(n_38),
.A2(n_42),
.B(n_46),
.Y(n_37)
);

AND2x2_ASAP7_75t_L g48 ( 
.A(n_38),
.B(n_49),
.Y(n_48)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_38),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_38),
.B(n_101),
.Y(n_226)
);

OAI22xp33_ASAP7_75t_L g49 ( 
.A1(n_39),
.A2(n_40),
.B1(n_43),
.B2(n_44),
.Y(n_49)
);

CKINVDCx14_ASAP7_75t_SL g39 ( 
.A(n_40),
.Y(n_39)
);

INVx13_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_42),
.Y(n_89)
);

OA22x2_ASAP7_75t_L g73 ( 
.A1(n_43),
.A2(n_44),
.B1(n_74),
.B2(n_75),
.Y(n_73)
);

NAND3xp33_ASAP7_75t_SL g187 ( 
.A(n_43),
.B(n_57),
.C(n_74),
.Y(n_187)
);

INVx4_ASAP7_75t_SL g43 ( 
.A(n_44),
.Y(n_43)
);

A2O1A1Ixp33_ASAP7_75t_L g184 ( 
.A1(n_44),
.A2(n_75),
.B(n_185),
.C(n_187),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_44),
.B(n_209),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_47),
.B(n_48),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_47),
.B(n_90),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_48),
.A2(n_89),
.B1(n_90),
.B2(n_91),
.Y(n_88)
);

AOI21xp5_ASAP7_75t_L g116 ( 
.A1(n_48),
.A2(n_91),
.B(n_117),
.Y(n_116)
);

CKINVDCx16_ASAP7_75t_R g149 ( 
.A(n_48),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_48),
.A2(n_90),
.B1(n_180),
.B2(n_202),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_48),
.A2(n_90),
.B1(n_211),
.B2(n_212),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_48),
.A2(n_90),
.B1(n_202),
.B2(n_212),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_51),
.A2(n_52),
.B1(n_69),
.B2(n_80),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g52 ( 
.A1(n_53),
.A2(n_54),
.B1(n_65),
.B2(n_67),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_53),
.A2(n_54),
.B1(n_65),
.B2(n_107),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_SL g128 ( 
.A1(n_53),
.A2(n_67),
.B(n_129),
.Y(n_128)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_53),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_54),
.B(n_60),
.Y(n_53)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_54),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g54 ( 
.A1(n_55),
.A2(n_56),
.B1(n_57),
.B2(n_59),
.Y(n_54)
);

INVx1_ASAP7_75t_SL g59 ( 
.A(n_55),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_55),
.A2(n_59),
.B1(n_61),
.B2(n_62),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_56),
.A2(n_57),
.B1(n_74),
.B2(n_75),
.Y(n_76)
);

OAI21xp33_ASAP7_75t_L g100 ( 
.A1(n_56),
.A2(n_59),
.B(n_101),
.Y(n_100)
);

INVx5_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

BUFx12f_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_69),
.Y(n_80)
);

OAI21xp5_ASAP7_75t_L g69 ( 
.A1(n_70),
.A2(n_72),
.B(n_77),
.Y(n_69)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_70),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_L g102 ( 
.A1(n_72),
.A2(n_103),
.B(n_104),
.Y(n_102)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_72),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_72),
.A2(n_73),
.B1(n_103),
.B2(n_146),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_72),
.A2(n_73),
.B1(n_146),
.B2(n_162),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g199 ( 
.A1(n_72),
.A2(n_73),
.B1(n_162),
.B2(n_200),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_73),
.B(n_76),
.Y(n_72)
);

CKINVDCx14_ASAP7_75t_R g79 ( 
.A(n_73),
.Y(n_79)
);

OAI21xp5_ASAP7_75t_L g124 ( 
.A1(n_73),
.A2(n_125),
.B(n_126),
.Y(n_124)
);

INVx8_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_78),
.B(n_79),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_78),
.B(n_127),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_79),
.B(n_105),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_82),
.A2(n_83),
.B1(n_88),
.B2(n_92),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_82),
.B(n_92),
.Y(n_121)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_SL g83 ( 
.A(n_84),
.B(n_87),
.Y(n_83)
);

CKINVDCx16_ASAP7_75t_R g84 ( 
.A(n_85),
.Y(n_84)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_86),
.Y(n_114)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_88),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_90),
.B(n_151),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_93),
.B(n_250),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_102),
.C(n_106),
.Y(n_93)
);

XNOR2xp5_ASAP7_75t_SL g164 ( 
.A(n_94),
.B(n_165),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_98),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_95),
.A2(n_98),
.B1(n_99),
.B2(n_155),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_95),
.Y(n_155)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

XNOR2xp5_ASAP7_75t_L g165 ( 
.A(n_102),
.B(n_106),
.Y(n_165)
);

CKINVDCx14_ASAP7_75t_R g143 ( 
.A(n_107),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_L g109 ( 
.A(n_110),
.B(n_134),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_111),
.A2(n_119),
.B1(n_132),
.B2(n_133),
.Y(n_110)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_111),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_112),
.A2(n_113),
.B1(n_115),
.B2(n_116),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_113),
.Y(n_112)
);

CKINVDCx14_ASAP7_75t_R g115 ( 
.A(n_116),
.Y(n_115)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_SL g148 ( 
.A1(n_118),
.A2(n_149),
.B(n_150),
.Y(n_148)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_119),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_120),
.A2(n_121),
.B1(n_122),
.B2(n_123),
.Y(n_119)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

XOR2xp5_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_128),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_131),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_130),
.A2(n_141),
.B1(n_142),
.B2(n_143),
.Y(n_140)
);

O2A1O1Ixp33_ASAP7_75t_L g136 ( 
.A1(n_137),
.A2(n_169),
.B(n_248),
.C(n_252),
.Y(n_136)
);

AND2x2_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_163),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_SL g247 ( 
.A(n_138),
.B(n_163),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_153),
.C(n_156),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_L g172 ( 
.A(n_139),
.B(n_173),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_SL g139 ( 
.A(n_140),
.B(n_144),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_140),
.B(n_147),
.C(n_152),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_145),
.A2(n_147),
.B1(n_148),
.B2(n_152),
.Y(n_144)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_145),
.Y(n_152)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_SL g178 ( 
.A1(n_149),
.A2(n_179),
.B(n_181),
.Y(n_178)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_153),
.A2(n_154),
.B1(n_156),
.B2(n_174),
.Y(n_173)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_156),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_159),
.C(n_161),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_157),
.A2(n_158),
.B1(n_159),
.B2(n_160),
.Y(n_177)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_SL g176 ( 
.A(n_161),
.B(n_177),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_L g163 ( 
.A(n_164),
.B(n_166),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_164),
.B(n_167),
.C(n_168),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g166 ( 
.A(n_167),
.B(n_168),
.Y(n_166)
);

AOI21xp5_ASAP7_75t_L g169 ( 
.A1(n_170),
.A2(n_246),
.B(n_247),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_190),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_172),
.B(n_175),
.Y(n_171)
);

OR2x2_ASAP7_75t_L g246 ( 
.A(n_172),
.B(n_175),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_176),
.B(n_178),
.C(n_182),
.Y(n_175)
);

XOR2xp5_ASAP7_75t_L g192 ( 
.A(n_176),
.B(n_193),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_178),
.A2(n_182),
.B1(n_183),
.B2(n_194),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_178),
.Y(n_194)
);

CKINVDCx16_ASAP7_75t_R g179 ( 
.A(n_180),
.Y(n_179)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_188),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_184),
.A2(n_188),
.B1(n_189),
.B2(n_197),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_184),
.Y(n_197)
);

INVxp67_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_L g190 ( 
.A1(n_191),
.A2(n_203),
.B(n_245),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_SL g191 ( 
.A(n_192),
.B(n_195),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_192),
.B(n_195),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_198),
.C(n_201),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_196),
.B(n_241),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_198),
.A2(n_199),
.B1(n_201),
.B2(n_242),
.Y(n_241)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_201),
.Y(n_242)
);

AOI21xp5_ASAP7_75t_SL g203 ( 
.A1(n_204),
.A2(n_239),
.B(n_244),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_L g204 ( 
.A1(n_205),
.A2(n_229),
.B(n_238),
.Y(n_204)
);

AOI21xp5_ASAP7_75t_L g205 ( 
.A1(n_206),
.A2(n_218),
.B(n_228),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_207),
.B(n_213),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_207),
.B(n_213),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_210),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_208),
.B(n_210),
.Y(n_230)
);

INVxp67_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_L g218 ( 
.A1(n_219),
.A2(n_224),
.B(n_227),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_220),
.B(n_222),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_SL g224 ( 
.A(n_225),
.B(n_226),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_225),
.B(n_226),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_230),
.B(n_231),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_230),
.B(n_231),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_232),
.B(n_233),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_232),
.B(n_234),
.C(n_237),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_234),
.A2(n_235),
.B1(n_236),
.B2(n_237),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_236),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_240),
.B(n_243),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_240),
.B(n_243),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_249),
.B(n_251),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_249),
.B(n_251),
.Y(n_252)
);


endmodule