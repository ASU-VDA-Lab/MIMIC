module fake_jpeg_19692_n_175 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_175);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_175;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_14;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx6_ASAP7_75t_L g13 ( 
.A(n_5),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_1),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_3),
.Y(n_15)
);

INVx11_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_12),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_12),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_3),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

INVx8_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_4),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

INVx6_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

INVx3_ASAP7_75t_SL g28 ( 
.A(n_20),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_28),
.B(n_30),
.Y(n_41)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_20),
.Y(n_29)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_29),
.Y(n_52)
);

INVx5_ASAP7_75t_L g30 ( 
.A(n_20),
.Y(n_30)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_20),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_31),
.B(n_32),
.Y(n_42)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_20),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_20),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_33),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_17),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_34),
.Y(n_49)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_21),
.Y(n_35)
);

INVx5_ASAP7_75t_L g50 ( 
.A(n_35),
.Y(n_50)
);

CKINVDCx16_ASAP7_75t_R g36 ( 
.A(n_15),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_36),
.B(n_38),
.Y(n_48)
);

BUFx24_ASAP7_75t_L g37 ( 
.A(n_24),
.Y(n_37)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_37),
.Y(n_46)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_21),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_34),
.B(n_13),
.Y(n_39)
);

MAJIxp5_ASAP7_75t_L g79 ( 
.A(n_39),
.B(n_44),
.C(n_47),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g40 ( 
.A1(n_28),
.A2(n_13),
.B1(n_25),
.B2(n_21),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_40),
.A2(n_45),
.B1(n_37),
.B2(n_35),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_34),
.B(n_13),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_28),
.A2(n_13),
.B1(n_25),
.B2(n_21),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_36),
.B(n_25),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_L g51 ( 
.A1(n_29),
.A2(n_16),
.B1(n_26),
.B2(n_22),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g53 ( 
.A1(n_51),
.A2(n_26),
.B1(n_15),
.B2(n_22),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_53),
.A2(n_58),
.B1(n_68),
.B2(n_74),
.Y(n_97)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_49),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_54),
.B(n_65),
.Y(n_85)
);

NOR2x1_ASAP7_75t_L g55 ( 
.A(n_51),
.B(n_37),
.Y(n_55)
);

OR2x2_ASAP7_75t_L g98 ( 
.A(n_55),
.B(n_56),
.Y(n_98)
);

OAI21xp33_ASAP7_75t_L g56 ( 
.A1(n_47),
.A2(n_37),
.B(n_18),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_48),
.B(n_18),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_SL g94 ( 
.A(n_57),
.B(n_69),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g58 ( 
.A1(n_39),
.A2(n_32),
.B1(n_31),
.B2(n_30),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_42),
.Y(n_59)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_59),
.Y(n_86)
);

BUFx2_ASAP7_75t_L g60 ( 
.A(n_46),
.Y(n_60)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_60),
.Y(n_99)
);

BUFx2_ASAP7_75t_L g61 ( 
.A(n_46),
.Y(n_61)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_61),
.Y(n_102)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_46),
.Y(n_62)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_62),
.Y(n_84)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_42),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_63),
.Y(n_87)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_41),
.Y(n_64)
);

AND2x2_ASAP7_75t_L g92 ( 
.A(n_64),
.B(n_72),
.Y(n_92)
);

CKINVDCx14_ASAP7_75t_R g65 ( 
.A(n_48),
.Y(n_65)
);

BUFx4f_ASAP7_75t_SL g66 ( 
.A(n_43),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_66),
.B(n_70),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_40),
.A2(n_15),
.B1(n_22),
.B2(n_26),
.Y(n_67)
);

INVxp67_ASAP7_75t_L g91 ( 
.A(n_67),
.Y(n_91)
);

OR2x2_ASAP7_75t_L g69 ( 
.A(n_41),
.B(n_23),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_52),
.B(n_23),
.Y(n_70)
);

INVxp67_ASAP7_75t_L g71 ( 
.A(n_45),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_71),
.A2(n_75),
.B1(n_17),
.B2(n_2),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_52),
.B(n_19),
.Y(n_72)
);

XOR2xp5_ASAP7_75t_L g73 ( 
.A(n_39),
.B(n_24),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_73),
.B(n_17),
.C(n_2),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_44),
.A2(n_35),
.B1(n_38),
.B2(n_16),
.Y(n_74)
);

INVx6_ASAP7_75t_L g75 ( 
.A(n_50),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_52),
.B(n_14),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_76),
.B(n_78),
.Y(n_100)
);

CKINVDCx16_ASAP7_75t_R g77 ( 
.A(n_43),
.Y(n_77)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_77),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_44),
.B(n_19),
.Y(n_78)
);

OAI22xp33_ASAP7_75t_L g80 ( 
.A1(n_50),
.A2(n_16),
.B1(n_33),
.B2(n_27),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_80),
.A2(n_50),
.B1(n_49),
.B2(n_27),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_L g113 ( 
.A1(n_81),
.A2(n_89),
.B1(n_86),
.B2(n_54),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_71),
.A2(n_49),
.B1(n_33),
.B2(n_27),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_82),
.A2(n_67),
.B1(n_64),
.B2(n_55),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_59),
.A2(n_14),
.B1(n_17),
.B2(n_24),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_83),
.A2(n_101),
.B1(n_4),
.B2(n_5),
.Y(n_117)
);

AOI21xp5_ASAP7_75t_L g89 ( 
.A1(n_68),
.A2(n_43),
.B(n_1),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_SL g106 ( 
.A1(n_89),
.A2(n_74),
.B(n_53),
.Y(n_106)
);

CKINVDCx16_ASAP7_75t_R g111 ( 
.A(n_90),
.Y(n_111)
);

XOR2xp5_ASAP7_75t_L g116 ( 
.A(n_95),
.B(n_96),
.Y(n_116)
);

XNOR2xp5_ASAP7_75t_L g96 ( 
.A(n_73),
.B(n_0),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_63),
.A2(n_0),
.B1(n_4),
.B2(n_5),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_103),
.A2(n_113),
.B1(n_117),
.B2(n_119),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_96),
.B(n_79),
.C(n_58),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_104),
.B(n_88),
.C(n_81),
.Y(n_134)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_99),
.Y(n_105)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_105),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_SL g128 ( 
.A1(n_106),
.A2(n_92),
.B(n_98),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_87),
.B(n_69),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_107),
.B(n_109),
.Y(n_124)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_99),
.Y(n_108)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_108),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_87),
.B(n_79),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_86),
.B(n_61),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_110),
.B(n_118),
.Y(n_122)
);

AO21x1_ASAP7_75t_L g112 ( 
.A1(n_91),
.A2(n_80),
.B(n_75),
.Y(n_112)
);

AOI21xp5_ASAP7_75t_L g121 ( 
.A1(n_112),
.A2(n_91),
.B(n_82),
.Y(n_121)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_102),
.Y(n_114)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_114),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_95),
.B(n_60),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_115),
.B(n_120),
.Y(n_133)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_84),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_97),
.A2(n_66),
.B1(n_62),
.B2(n_8),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_97),
.A2(n_66),
.B1(n_7),
.B2(n_8),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_L g145 ( 
.A1(n_121),
.A2(n_126),
.B(n_128),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_105),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_123),
.B(n_118),
.Y(n_137)
);

NOR2xp67_ASAP7_75t_R g126 ( 
.A(n_103),
.B(n_98),
.Y(n_126)
);

AOI21x1_ASAP7_75t_L g130 ( 
.A1(n_115),
.A2(n_92),
.B(n_100),
.Y(n_130)
);

XNOR2xp5_ASAP7_75t_L g141 ( 
.A(n_130),
.B(n_116),
.Y(n_141)
);

OAI32xp33_ASAP7_75t_L g132 ( 
.A1(n_106),
.A2(n_100),
.A3(n_94),
.B1(n_85),
.B2(n_92),
.Y(n_132)
);

XOR2xp5_ASAP7_75t_L g142 ( 
.A(n_132),
.B(n_116),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_134),
.B(n_128),
.C(n_126),
.Y(n_146)
);

AOI21xp5_ASAP7_75t_L g135 ( 
.A1(n_112),
.A2(n_111),
.B(n_119),
.Y(n_135)
);

CKINVDCx14_ASAP7_75t_R g140 ( 
.A(n_135),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g136 ( 
.A1(n_131),
.A2(n_111),
.B1(n_120),
.B2(n_104),
.Y(n_136)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_136),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_137),
.B(n_138),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_124),
.B(n_93),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_133),
.A2(n_117),
.B1(n_112),
.B2(n_114),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_139),
.B(n_143),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_141),
.B(n_142),
.C(n_146),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_131),
.A2(n_108),
.B1(n_93),
.B2(n_102),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_122),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_SL g151 ( 
.A1(n_144),
.A2(n_127),
.B(n_129),
.Y(n_151)
);

HB1xp67_ASAP7_75t_L g149 ( 
.A(n_145),
.Y(n_149)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_149),
.Y(n_159)
);

AOI21xp5_ASAP7_75t_L g150 ( 
.A1(n_145),
.A2(n_132),
.B(n_133),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_150),
.B(n_151),
.Y(n_158)
);

AOI21xp5_ASAP7_75t_L g153 ( 
.A1(n_144),
.A2(n_130),
.B(n_129),
.Y(n_153)
);

XOR2xp5_ASAP7_75t_L g155 ( 
.A(n_153),
.B(n_134),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_155),
.B(n_6),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_152),
.A2(n_140),
.B1(n_139),
.B2(n_135),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_156),
.A2(n_157),
.B1(n_160),
.B2(n_147),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_152),
.A2(n_143),
.B1(n_141),
.B2(n_121),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_148),
.A2(n_146),
.B1(n_142),
.B2(n_125),
.Y(n_160)
);

AOI21xp5_ASAP7_75t_L g161 ( 
.A1(n_154),
.A2(n_125),
.B(n_84),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_SL g164 ( 
.A1(n_161),
.A2(n_7),
.B(n_9),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_162),
.B(n_157),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_163),
.B(n_155),
.C(n_159),
.Y(n_167)
);

AOI21xp5_ASAP7_75t_L g169 ( 
.A1(n_164),
.A2(n_165),
.B(n_166),
.Y(n_169)
);

INVxp67_ASAP7_75t_L g165 ( 
.A(n_158),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_L g166 ( 
.A1(n_160),
.A2(n_9),
.B(n_10),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_SL g170 ( 
.A1(n_167),
.A2(n_168),
.B(n_165),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_170),
.B(n_171),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_SL g171 ( 
.A1(n_169),
.A2(n_156),
.B(n_10),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_170),
.B(n_9),
.C(n_10),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_172),
.B(n_11),
.C(n_173),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_174),
.B(n_11),
.Y(n_175)
);


endmodule