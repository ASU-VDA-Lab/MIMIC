module real_aes_14941_n_77 (n_17, n_28, n_76, n_56, n_34, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_43, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_44, n_7, n_4, n_6, n_12, n_68, n_69, n_46, n_59, n_25, n_73, n_48, n_37, n_70, n_50, n_26, n_13, n_24, n_2, n_55, n_62, n_67, n_33, n_14, n_11, n_16, n_39, n_5, n_45, n_60, n_38, n_0, n_63, n_1, n_53, n_36, n_77);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_43;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_44;
input n_7;
input n_4;
input n_6;
input n_12;
input n_68;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_48;
input n_37;
input n_70;
input n_50;
input n_26;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_67;
input n_33;
input n_14;
input n_11;
input n_16;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_0;
input n_63;
input n_1;
input n_53;
input n_36;
output n_77;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_90;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_83;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_364;
wire n_319;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_97;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_548;
wire n_678;
wire n_427;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_92;
wire n_564;
wire n_519;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_94;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_98;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_82;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_178;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_80;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_339;
wire n_398;
wire n_89;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_93;
wire n_182;
wire n_449;
wire n_417;
wire n_363;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_505;
wire n_434;
wire n_502;
wire n_527;
wire n_600;
wire n_250;
wire n_85;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_87;
wire n_171;
wire n_658;
wire n_676;
wire n_78;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_96;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_95;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_81;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_88;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_653;
wire n_365;
wire n_290;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_420;
wire n_336;
wire n_349;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_249;
wire n_623;
wire n_446;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_99;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_79;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_566;
wire n_474;
wire n_170;
wire n_86;
wire n_375;
wire n_597;
wire n_640;
wire n_340;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_84;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
wire n_91;
INVx1_ASAP7_75t_L g90 ( .A(n_0), .Y(n_90) );
OA21x2_ASAP7_75t_L g164 ( .A1(n_0), .A2(n_40), .B(n_92), .Y(n_164) );
NAND2xp5_ASAP7_75t_L g157 ( .A(n_1), .B(n_158), .Y(n_157) );
NAND2xp33_ASAP7_75t_L g182 ( .A(n_2), .B(n_183), .Y(n_182) );
INVx1_ASAP7_75t_L g511 ( .A(n_3), .Y(n_511) );
AOI22xp33_ASAP7_75t_L g610 ( .A1(n_3), .A2(n_64), .B1(n_611), .B2(n_614), .Y(n_610) );
BUFx3_ASAP7_75t_L g581 ( .A(n_4), .Y(n_581) );
INVx3_ASAP7_75t_L g572 ( .A(n_5), .Y(n_572) );
NAND2xp5_ASAP7_75t_L g212 ( .A(n_6), .B(n_106), .Y(n_212) );
INVx2_ASAP7_75t_L g588 ( .A(n_7), .Y(n_588) );
INVx1_ASAP7_75t_L g604 ( .A(n_7), .Y(n_604) );
CKINVDCx5p33_ASAP7_75t_R g87 ( .A(n_8), .Y(n_87) );
BUFx3_ASAP7_75t_L g108 ( .A(n_9), .Y(n_108) );
INVx1_ASAP7_75t_L g125 ( .A(n_9), .Y(n_125) );
A2O1A1Ixp33_ASAP7_75t_L g138 ( .A1(n_10), .A2(n_139), .B(n_140), .C(n_142), .Y(n_138) );
BUFx10_ASAP7_75t_L g689 ( .A(n_11), .Y(n_689) );
CKINVDCx5p33_ASAP7_75t_R g198 ( .A(n_12), .Y(n_198) );
NAND2xp5_ASAP7_75t_L g216 ( .A(n_13), .B(n_217), .Y(n_216) );
NAND2xp5_ASAP7_75t_L g174 ( .A(n_14), .B(n_175), .Y(n_174) );
NAND2xp5_ASAP7_75t_L g262 ( .A(n_15), .B(n_205), .Y(n_262) );
A2O1A1Ixp33_ASAP7_75t_L g121 ( .A1(n_16), .A2(n_122), .B(n_126), .C(n_129), .Y(n_121) );
AND2x2_ASAP7_75t_L g195 ( .A(n_17), .B(n_194), .Y(n_195) );
AND2x2_ASAP7_75t_L g500 ( .A(n_18), .B(n_501), .Y(n_500) );
AND2x2_ASAP7_75t_L g508 ( .A(n_18), .B(n_29), .Y(n_508) );
INVx1_ASAP7_75t_L g538 ( .A(n_18), .Y(n_538) );
NAND2xp5_ASAP7_75t_L g220 ( .A(n_19), .B(n_185), .Y(n_220) );
AOI22xp33_ASAP7_75t_L g113 ( .A1(n_20), .A2(n_55), .B1(n_109), .B2(n_114), .Y(n_113) );
INVx1_ASAP7_75t_L g98 ( .A(n_21), .Y(n_98) );
INVx2_ASAP7_75t_L g505 ( .A(n_22), .Y(n_505) );
INVx1_ASAP7_75t_L g540 ( .A(n_23), .Y(n_540) );
INVx1_ASAP7_75t_L g162 ( .A(n_24), .Y(n_162) );
NAND2xp5_ASAP7_75t_SL g211 ( .A(n_25), .B(n_109), .Y(n_211) );
NAND2xp5_ASAP7_75t_L g184 ( .A(n_26), .B(n_185), .Y(n_184) );
AOI22xp33_ASAP7_75t_L g543 ( .A1(n_27), .A2(n_68), .B1(n_544), .B2(n_545), .Y(n_543) );
OAI22xp5_ASAP7_75t_L g639 ( .A1(n_27), .A2(n_640), .B1(n_643), .B2(n_653), .Y(n_639) );
NAND2xp5_ASAP7_75t_SL g261 ( .A(n_28), .B(n_123), .Y(n_261) );
INVx2_ASAP7_75t_L g501 ( .A(n_29), .Y(n_501) );
NAND2xp5_ASAP7_75t_L g551 ( .A(n_29), .B(n_538), .Y(n_551) );
OAI22xp33_ASAP7_75t_L g497 ( .A1(n_30), .A2(n_42), .B1(n_498), .B2(n_506), .Y(n_497) );
AOI22xp33_ASAP7_75t_L g617 ( .A1(n_30), .A2(n_43), .B1(n_618), .B2(n_621), .Y(n_617) );
OAI22xp5_ASAP7_75t_L g676 ( .A1(n_31), .A2(n_55), .B1(n_677), .B2(n_678), .Y(n_676) );
INVx1_ASAP7_75t_L g678 ( .A(n_31), .Y(n_678) );
NAND2xp5_ASAP7_75t_L g234 ( .A(n_32), .B(n_185), .Y(n_234) );
NAND2xp5_ASAP7_75t_SL g202 ( .A(n_33), .B(n_203), .Y(n_202) );
INVx1_ASAP7_75t_L g522 ( .A(n_34), .Y(n_522) );
CKINVDCx5p33_ASAP7_75t_R g141 ( .A(n_35), .Y(n_141) );
AND2x4_ASAP7_75t_L g97 ( .A(n_36), .B(n_98), .Y(n_97) );
HB1xp67_ASAP7_75t_L g664 ( .A(n_36), .Y(n_664) );
AOI21xp33_ASAP7_75t_L g547 ( .A1(n_37), .A2(n_548), .B(n_550), .Y(n_547) );
INVxp67_ASAP7_75t_SL g638 ( .A(n_37), .Y(n_638) );
INVx1_ASAP7_75t_L g586 ( .A(n_38), .Y(n_586) );
INVx1_ASAP7_75t_L g594 ( .A(n_38), .Y(n_594) );
AOI22xp33_ASAP7_75t_L g105 ( .A1(n_39), .A2(n_63), .B1(n_106), .B2(n_109), .Y(n_105) );
INVx1_ASAP7_75t_L g89 ( .A(n_40), .Y(n_89) );
INVx1_ASAP7_75t_L g92 ( .A(n_41), .Y(n_92) );
INVx1_ASAP7_75t_L g575 ( .A(n_42), .Y(n_575) );
AOI22xp33_ASAP7_75t_L g528 ( .A1(n_43), .A2(n_70), .B1(n_518), .B2(n_529), .Y(n_528) );
AND2x2_ASAP7_75t_L g269 ( .A(n_44), .B(n_186), .Y(n_269) );
INVx1_ASAP7_75t_L g671 ( .A(n_45), .Y(n_671) );
NAND2xp5_ASAP7_75t_L g204 ( .A(n_46), .B(n_205), .Y(n_204) );
NAND2x1_ASAP7_75t_L g232 ( .A(n_47), .B(n_139), .Y(n_232) );
NAND2xp5_ASAP7_75t_L g180 ( .A(n_48), .B(n_181), .Y(n_180) );
HB1xp67_ASAP7_75t_L g674 ( .A(n_49), .Y(n_674) );
INVx1_ASAP7_75t_L g516 ( .A(n_50), .Y(n_516) );
NAND2xp5_ASAP7_75t_L g149 ( .A(n_51), .B(n_150), .Y(n_149) );
NAND2xp5_ASAP7_75t_SL g214 ( .A(n_52), .B(n_215), .Y(n_214) );
NAND2xp5_ASAP7_75t_SL g226 ( .A(n_53), .B(n_227), .Y(n_226) );
NAND2xp5_ASAP7_75t_L g135 ( .A(n_54), .B(n_136), .Y(n_135) );
INVx1_ASAP7_75t_L g677 ( .A(n_55), .Y(n_677) );
HB1xp67_ASAP7_75t_L g669 ( .A(n_56), .Y(n_669) );
NAND2xp5_ASAP7_75t_SL g268 ( .A(n_57), .B(n_123), .Y(n_268) );
CKINVDCx5p33_ASAP7_75t_R g230 ( .A(n_58), .Y(n_230) );
NAND2xp5_ASAP7_75t_L g228 ( .A(n_59), .B(n_217), .Y(n_228) );
NAND2xp33_ASAP7_75t_SL g155 ( .A(n_60), .B(n_156), .Y(n_155) );
NAND2xp5_ASAP7_75t_SL g146 ( .A(n_61), .B(n_147), .Y(n_146) );
OAI211xp5_ASAP7_75t_L g552 ( .A1(n_62), .A2(n_553), .B(n_557), .C(n_562), .Y(n_552) );
AOI22xp33_ASAP7_75t_L g649 ( .A1(n_62), .A2(n_70), .B1(n_650), .B2(n_651), .Y(n_649) );
AOI21xp33_ASAP7_75t_L g531 ( .A1(n_64), .A2(n_532), .B(n_536), .Y(n_531) );
INVx1_ASAP7_75t_L g102 ( .A(n_65), .Y(n_102) );
BUFx3_ASAP7_75t_L g131 ( .A(n_65), .Y(n_131) );
INVx1_ASAP7_75t_L g153 ( .A(n_65), .Y(n_153) );
CKINVDCx5p33_ASAP7_75t_R g127 ( .A(n_66), .Y(n_127) );
NAND2xp5_ASAP7_75t_L g266 ( .A(n_67), .B(n_267), .Y(n_266) );
INVxp67_ASAP7_75t_SL g633 ( .A(n_68), .Y(n_633) );
INVx2_ASAP7_75t_L g504 ( .A(n_69), .Y(n_504) );
AND2x2_ASAP7_75t_L g515 ( .A(n_69), .B(n_505), .Y(n_515) );
INVxp67_ASAP7_75t_SL g534 ( .A(n_69), .Y(n_534) );
XNOR2xp5_ASAP7_75t_L g494 ( .A(n_71), .B(n_495), .Y(n_494) );
NAND2xp33_ASAP7_75t_L g176 ( .A(n_72), .B(n_177), .Y(n_176) );
INVx1_ASAP7_75t_L g569 ( .A(n_73), .Y(n_569) );
INVx2_ASAP7_75t_L g580 ( .A(n_74), .Y(n_580) );
INVx1_ASAP7_75t_L g565 ( .A(n_75), .Y(n_565) );
NAND2xp5_ASAP7_75t_SL g200 ( .A(n_76), .B(n_147), .Y(n_200) );
AOI21xp33_ASAP7_75t_L g77 ( .A1(n_78), .A2(n_483), .B(n_493), .Y(n_77) );
INVx2_ASAP7_75t_L g78 ( .A(n_79), .Y(n_78) );
AND2x2_ASAP7_75t_L g79 ( .A(n_80), .B(n_387), .Y(n_79) );
NOR3xp33_ASAP7_75t_L g80 ( .A(n_81), .B(n_296), .C(n_360), .Y(n_80) );
OAI221xp5_ASAP7_75t_L g81 ( .A1(n_82), .A2(n_188), .B1(n_235), .B2(n_246), .C(n_251), .Y(n_81) );
NAND2xp5_ASAP7_75t_L g82 ( .A(n_83), .B(n_116), .Y(n_82) );
INVx2_ASAP7_75t_L g83 ( .A(n_84), .Y(n_83) );
AND2x2_ASAP7_75t_L g308 ( .A(n_84), .B(n_309), .Y(n_308) );
AND2x2_ASAP7_75t_L g323 ( .A(n_84), .B(n_324), .Y(n_323) );
AND2x2_ASAP7_75t_L g396 ( .A(n_84), .B(n_143), .Y(n_396) );
INVx1_ASAP7_75t_L g84 ( .A(n_85), .Y(n_84) );
INVx1_ASAP7_75t_L g243 ( .A(n_85), .Y(n_243) );
INVx1_ASAP7_75t_L g275 ( .A(n_85), .Y(n_275) );
AND2x2_ASAP7_75t_L g294 ( .A(n_85), .B(n_295), .Y(n_294) );
AND2x2_ASAP7_75t_L g321 ( .A(n_85), .B(n_311), .Y(n_321) );
INVxp67_ASAP7_75t_L g336 ( .A(n_85), .Y(n_336) );
AND2x2_ASAP7_75t_L g359 ( .A(n_85), .B(n_170), .Y(n_359) );
HB1xp67_ASAP7_75t_L g386 ( .A(n_85), .Y(n_386) );
OR2x2_ASAP7_75t_L g85 ( .A(n_86), .B(n_93), .Y(n_85) );
NOR2xp33_ASAP7_75t_L g86 ( .A(n_87), .B(n_88), .Y(n_86) );
NAND2xp5_ASAP7_75t_L g132 ( .A(n_88), .B(n_133), .Y(n_132) );
INVx2_ASAP7_75t_L g136 ( .A(n_88), .Y(n_136) );
AO21x2_ASAP7_75t_L g88 ( .A1(n_89), .A2(n_90), .B(n_91), .Y(n_88) );
AOI21x1_ASAP7_75t_L g104 ( .A1(n_89), .A2(n_90), .B(n_91), .Y(n_104) );
INVx1_ASAP7_75t_L g91 ( .A(n_92), .Y(n_91) );
OAI22xp5_ASAP7_75t_L g93 ( .A1(n_94), .A2(n_105), .B1(n_111), .B2(n_113), .Y(n_93) );
NAND3xp33_ASAP7_75t_L g94 ( .A(n_95), .B(n_99), .C(n_103), .Y(n_94) );
NAND3xp33_ASAP7_75t_L g111 ( .A(n_95), .B(n_103), .C(n_112), .Y(n_111) );
BUFx2_ASAP7_75t_L g486 ( .A(n_95), .Y(n_486) );
INVx1_ASAP7_75t_L g95 ( .A(n_96), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_97), .Y(n_96) );
INVx2_ASAP7_75t_L g134 ( .A(n_97), .Y(n_134) );
BUFx6f_ASAP7_75t_SL g168 ( .A(n_97), .Y(n_168) );
INVx1_ASAP7_75t_L g259 ( .A(n_97), .Y(n_259) );
HB1xp67_ASAP7_75t_L g662 ( .A(n_98), .Y(n_662) );
INVx1_ASAP7_75t_L g99 ( .A(n_100), .Y(n_99) );
INVx2_ASAP7_75t_L g100 ( .A(n_101), .Y(n_100) );
INVx2_ASAP7_75t_L g142 ( .A(n_101), .Y(n_142) );
INVx2_ASAP7_75t_L g101 ( .A(n_102), .Y(n_101) );
BUFx3_ASAP7_75t_L g112 ( .A(n_102), .Y(n_112) );
INVx2_ASAP7_75t_L g103 ( .A(n_104), .Y(n_103) );
INVx2_ASAP7_75t_L g106 ( .A(n_107), .Y(n_106) );
INVx2_ASAP7_75t_L g158 ( .A(n_107), .Y(n_158) );
INVx2_ASAP7_75t_L g181 ( .A(n_107), .Y(n_181) );
INVx2_ASAP7_75t_L g205 ( .A(n_107), .Y(n_205) );
BUFx6f_ASAP7_75t_L g107 ( .A(n_108), .Y(n_107) );
INVx2_ASAP7_75t_L g110 ( .A(n_108), .Y(n_110) );
BUFx6f_ASAP7_75t_L g115 ( .A(n_108), .Y(n_115) );
INVx2_ASAP7_75t_L g109 ( .A(n_110), .Y(n_109) );
INVx2_ASAP7_75t_L g183 ( .A(n_110), .Y(n_183) );
INVx1_ASAP7_75t_L g227 ( .A(n_110), .Y(n_227) );
O2A1O1Ixp5_ASAP7_75t_L g229 ( .A1(n_112), .A2(n_230), .B(n_231), .C(n_232), .Y(n_229) );
INVx2_ASAP7_75t_L g263 ( .A(n_112), .Y(n_263) );
INVx2_ASAP7_75t_L g114 ( .A(n_115), .Y(n_114) );
INVx1_ASAP7_75t_L g150 ( .A(n_115), .Y(n_150) );
INVx2_ASAP7_75t_L g175 ( .A(n_115), .Y(n_175) );
INVx2_ASAP7_75t_L g267 ( .A(n_115), .Y(n_267) );
OAI21xp33_ASAP7_75t_L g364 ( .A1(n_116), .A2(n_365), .B(n_369), .Y(n_364) );
AND2x2_ASAP7_75t_L g116 ( .A(n_117), .B(n_143), .Y(n_116) );
AND2x2_ASAP7_75t_L g466 ( .A(n_117), .B(n_359), .Y(n_466) );
INVx1_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
BUFx2_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
INVx1_ASAP7_75t_L g239 ( .A(n_119), .Y(n_239) );
INVx1_ASAP7_75t_L g277 ( .A(n_119), .Y(n_277) );
AND2x2_ASAP7_75t_L g305 ( .A(n_119), .B(n_242), .Y(n_305) );
HB1xp67_ASAP7_75t_L g334 ( .A(n_119), .Y(n_334) );
NAND2x1p5_ASAP7_75t_L g119 ( .A(n_120), .B(n_137), .Y(n_119) );
NAND2x1p5_ASAP7_75t_L g295 ( .A(n_120), .B(n_137), .Y(n_295) );
OA21x2_ASAP7_75t_L g120 ( .A1(n_121), .A2(n_132), .B(n_135), .Y(n_120) );
INVx1_ASAP7_75t_L g122 ( .A(n_123), .Y(n_122) );
NOR2xp33_ASAP7_75t_L g140 ( .A(n_123), .B(n_141), .Y(n_140) );
BUFx6f_ASAP7_75t_L g123 ( .A(n_124), .Y(n_123) );
INVx3_ASAP7_75t_L g128 ( .A(n_124), .Y(n_128) );
INVx2_ASAP7_75t_L g124 ( .A(n_125), .Y(n_124) );
BUFx6f_ASAP7_75t_L g148 ( .A(n_125), .Y(n_148) );
NOR2xp33_ASAP7_75t_L g126 ( .A(n_127), .B(n_128), .Y(n_126) );
INVx2_ASAP7_75t_L g139 ( .A(n_128), .Y(n_139) );
INVx2_ASAP7_75t_L g199 ( .A(n_128), .Y(n_199) );
INVx2_ASAP7_75t_L g215 ( .A(n_128), .Y(n_215) );
AOI21xp5_ASAP7_75t_L g179 ( .A1(n_129), .A2(n_180), .B(n_182), .Y(n_179) );
INVx1_ASAP7_75t_L g129 ( .A(n_130), .Y(n_129) );
INVx2_ASAP7_75t_L g130 ( .A(n_131), .Y(n_130) );
INVx2_ASAP7_75t_L g159 ( .A(n_131), .Y(n_159) );
INVx1_ASAP7_75t_L g178 ( .A(n_131), .Y(n_178) );
AOI211x1_ASAP7_75t_L g196 ( .A1(n_131), .A2(n_195), .B(n_197), .C(n_201), .Y(n_196) );
OR2x2_ASAP7_75t_L g137 ( .A(n_132), .B(n_138), .Y(n_137) );
INVx2_ASAP7_75t_SL g133 ( .A(n_134), .Y(n_133) );
INVx1_ASAP7_75t_L g233 ( .A(n_134), .Y(n_233) );
INVx1_ASAP7_75t_L g701 ( .A(n_141), .Y(n_701) );
AND2x2_ASAP7_75t_L g293 ( .A(n_143), .B(n_294), .Y(n_293) );
INVx3_ASAP7_75t_L g482 ( .A(n_143), .Y(n_482) );
AND2x2_ASAP7_75t_L g143 ( .A(n_144), .B(n_169), .Y(n_143) );
INVx2_ASAP7_75t_L g242 ( .A(n_144), .Y(n_242) );
AND2x2_ASAP7_75t_L g276 ( .A(n_144), .B(n_277), .Y(n_276) );
INVx1_ASAP7_75t_L g287 ( .A(n_144), .Y(n_287) );
OR2x2_ASAP7_75t_L g325 ( .A(n_144), .B(n_295), .Y(n_325) );
AND2x2_ASAP7_75t_L g337 ( .A(n_144), .B(n_295), .Y(n_337) );
AND2x2_ASAP7_75t_L g407 ( .A(n_144), .B(n_170), .Y(n_407) );
AO31x2_ASAP7_75t_L g144 ( .A1(n_145), .A2(n_154), .A3(n_160), .B(n_165), .Y(n_144) );
AO21x1_ASAP7_75t_L g145 ( .A1(n_146), .A2(n_149), .B(n_151), .Y(n_145) );
INVx2_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
INVx2_ASAP7_75t_L g156 ( .A(n_148), .Y(n_156) );
INVx1_ASAP7_75t_L g177 ( .A(n_148), .Y(n_177) );
INVx2_ASAP7_75t_L g203 ( .A(n_148), .Y(n_203) );
INVx2_ASAP7_75t_L g231 ( .A(n_150), .Y(n_231) );
AOI21xp5_ASAP7_75t_L g201 ( .A1(n_151), .A2(n_202), .B(n_204), .Y(n_201) );
AOI21xp5_ASAP7_75t_L g213 ( .A1(n_151), .A2(n_214), .B(n_216), .Y(n_213) );
AOI21xp5_ASAP7_75t_L g225 ( .A1(n_151), .A2(n_226), .B(n_228), .Y(n_225) );
BUFx10_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
INVx1_ASAP7_75t_L g152 ( .A(n_153), .Y(n_152) );
BUFx3_ASAP7_75t_L g489 ( .A(n_153), .Y(n_489) );
AO21x1_ASAP7_75t_L g154 ( .A1(n_155), .A2(n_157), .B(n_159), .Y(n_154) );
INVx2_ASAP7_75t_L g217 ( .A(n_156), .Y(n_217) );
AOI21xp5_ASAP7_75t_L g210 ( .A1(n_159), .A2(n_211), .B(n_212), .Y(n_210) );
INVx1_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
AOI21xp5_ASAP7_75t_L g165 ( .A1(n_161), .A2(n_166), .B(n_168), .Y(n_165) );
NOR2xp33_ASAP7_75t_L g161 ( .A(n_162), .B(n_163), .Y(n_161) );
INVxp33_ASAP7_75t_L g163 ( .A(n_164), .Y(n_163) );
BUFx2_ASAP7_75t_L g167 ( .A(n_164), .Y(n_167) );
INVx1_ASAP7_75t_L g187 ( .A(n_164), .Y(n_187) );
BUFx6f_ASAP7_75t_L g194 ( .A(n_164), .Y(n_194) );
INVx1_ASAP7_75t_L g166 ( .A(n_167), .Y(n_166) );
BUFx3_ASAP7_75t_L g171 ( .A(n_167), .Y(n_171) );
OAI21x1_ASAP7_75t_L g172 ( .A1(n_168), .A2(n_173), .B(n_179), .Y(n_172) );
AOI21xp5_ASAP7_75t_L g192 ( .A1(n_168), .A2(n_193), .B(n_195), .Y(n_192) );
OAI21x1_ASAP7_75t_L g209 ( .A1(n_168), .A2(n_210), .B(n_213), .Y(n_209) );
INVx1_ASAP7_75t_L g169 ( .A(n_170), .Y(n_169) );
INVx1_ASAP7_75t_L g245 ( .A(n_170), .Y(n_245) );
INVx1_ASAP7_75t_L g311 ( .A(n_170), .Y(n_311) );
AND2x2_ASAP7_75t_L g333 ( .A(n_170), .B(n_243), .Y(n_333) );
AND2x2_ASAP7_75t_L g416 ( .A(n_170), .B(n_310), .Y(n_416) );
OAI21x1_ASAP7_75t_L g170 ( .A1(n_171), .A2(n_172), .B(n_184), .Y(n_170) );
AOI21xp5_ASAP7_75t_L g173 ( .A1(n_174), .A2(n_176), .B(n_178), .Y(n_173) );
AOI21xp5_ASAP7_75t_L g265 ( .A1(n_178), .A2(n_266), .B(n_268), .Y(n_265) );
BUFx6f_ASAP7_75t_L g185 ( .A(n_186), .Y(n_185) );
INVx2_ASAP7_75t_L g186 ( .A(n_187), .Y(n_186) );
NAND2xp5_ASAP7_75t_L g188 ( .A(n_189), .B(n_206), .Y(n_188) );
AND2x2_ASAP7_75t_L g339 ( .A(n_189), .B(n_330), .Y(n_339) );
OR2x2_ASAP7_75t_L g355 ( .A(n_189), .B(n_290), .Y(n_355) );
INVx2_ASAP7_75t_L g367 ( .A(n_189), .Y(n_367) );
NAND2xp5_ASAP7_75t_L g370 ( .A(n_189), .B(n_303), .Y(n_370) );
AND2x2_ASAP7_75t_L g467 ( .A(n_189), .B(n_382), .Y(n_467) );
BUFx3_ASAP7_75t_L g189 ( .A(n_190), .Y(n_189) );
AND2x2_ASAP7_75t_L g247 ( .A(n_190), .B(n_248), .Y(n_247) );
OR2x2_ASAP7_75t_L g377 ( .A(n_190), .B(n_282), .Y(n_377) );
INVx2_ASAP7_75t_L g190 ( .A(n_191), .Y(n_190) );
AND2x2_ASAP7_75t_L g270 ( .A(n_191), .B(n_208), .Y(n_270) );
INVx2_ASAP7_75t_L g301 ( .A(n_191), .Y(n_301) );
BUFx2_ASAP7_75t_L g328 ( .A(n_191), .Y(n_328) );
HB1xp67_ASAP7_75t_L g345 ( .A(n_191), .Y(n_345) );
INVx1_ASAP7_75t_L g352 ( .A(n_191), .Y(n_352) );
AND2x2_ASAP7_75t_L g411 ( .A(n_191), .B(n_354), .Y(n_411) );
INVx1_ASAP7_75t_L g472 ( .A(n_191), .Y(n_472) );
OR2x6_ASAP7_75t_L g191 ( .A(n_192), .B(n_196), .Y(n_191) );
INVxp67_ASAP7_75t_SL g193 ( .A(n_194), .Y(n_193) );
BUFx6f_ASAP7_75t_L g219 ( .A(n_194), .Y(n_219) );
NOR2xp67_ASAP7_75t_SL g258 ( .A(n_194), .B(n_259), .Y(n_258) );
OAI21xp5_ASAP7_75t_L g197 ( .A1(n_198), .A2(n_199), .B(n_200), .Y(n_197) );
INVx2_ASAP7_75t_L g492 ( .A(n_203), .Y(n_492) );
AND2x2_ASAP7_75t_L g206 ( .A(n_207), .B(n_221), .Y(n_206) );
NAND2xp5_ASAP7_75t_L g427 ( .A(n_207), .B(n_428), .Y(n_427) );
INVx1_ASAP7_75t_L g207 ( .A(n_208), .Y(n_207) );
AND2x2_ASAP7_75t_L g281 ( .A(n_208), .B(n_282), .Y(n_281) );
OAI21xp5_ASAP7_75t_L g208 ( .A1(n_209), .A2(n_218), .B(n_220), .Y(n_208) );
OAI21x1_ASAP7_75t_L g250 ( .A1(n_209), .A2(n_218), .B(n_220), .Y(n_250) );
OAI21x1_ASAP7_75t_L g223 ( .A1(n_218), .A2(n_224), .B(n_234), .Y(n_223) );
BUFx6f_ASAP7_75t_L g218 ( .A(n_219), .Y(n_218) );
INVx2_ASAP7_75t_L g437 ( .A(n_221), .Y(n_437) );
INVx1_ASAP7_75t_L g221 ( .A(n_222), .Y(n_221) );
INVx2_ASAP7_75t_L g354 ( .A(n_222), .Y(n_354) );
INVx1_ASAP7_75t_L g222 ( .A(n_223), .Y(n_222) );
INVx1_ASAP7_75t_L g280 ( .A(n_223), .Y(n_280) );
INVx1_ASAP7_75t_L g317 ( .A(n_223), .Y(n_317) );
OAI21xp5_ASAP7_75t_L g224 ( .A1(n_225), .A2(n_229), .B(n_233), .Y(n_224) );
OAI211xp5_ASAP7_75t_L g360 ( .A1(n_235), .A2(n_361), .B(n_364), .C(n_371), .Y(n_360) );
INVx1_ASAP7_75t_L g235 ( .A(n_236), .Y(n_235) );
INVx2_ASAP7_75t_L g236 ( .A(n_237), .Y(n_236) );
NAND2x1p5_ASAP7_75t_L g237 ( .A(n_238), .B(n_240), .Y(n_237) );
INVx2_ASAP7_75t_L g238 ( .A(n_239), .Y(n_238) );
HB1xp67_ASAP7_75t_L g284 ( .A(n_239), .Y(n_284) );
AND2x2_ASAP7_75t_L g403 ( .A(n_239), .B(n_333), .Y(n_403) );
AND2x2_ASAP7_75t_L g240 ( .A(n_241), .B(n_244), .Y(n_240) );
AND2x2_ASAP7_75t_L g313 ( .A(n_241), .B(n_309), .Y(n_313) );
AND2x2_ASAP7_75t_L g241 ( .A(n_242), .B(n_243), .Y(n_241) );
INVx1_ASAP7_75t_L g374 ( .A(n_242), .Y(n_374) );
INVx2_ASAP7_75t_L g347 ( .A(n_244), .Y(n_347) );
BUFx3_ASAP7_75t_L g244 ( .A(n_245), .Y(n_244) );
NAND2xp5_ASAP7_75t_L g286 ( .A(n_245), .B(n_287), .Y(n_286) );
INVxp67_ASAP7_75t_SL g449 ( .A(n_245), .Y(n_449) );
INVx1_ASAP7_75t_L g246 ( .A(n_247), .Y(n_246) );
AND2x2_ASAP7_75t_L g303 ( .A(n_248), .B(n_280), .Y(n_303) );
INVx1_ASAP7_75t_L g248 ( .A(n_249), .Y(n_248) );
OR2x2_ASAP7_75t_L g316 ( .A(n_249), .B(n_317), .Y(n_316) );
AND2x2_ASAP7_75t_L g330 ( .A(n_249), .B(n_256), .Y(n_330) );
AND2x2_ASAP7_75t_L g453 ( .A(n_249), .B(n_280), .Y(n_453) );
INVx2_ASAP7_75t_L g249 ( .A(n_250), .Y(n_249) );
OR2x2_ASAP7_75t_L g291 ( .A(n_250), .B(n_256), .Y(n_291) );
AOI221xp5_ASAP7_75t_L g251 ( .A1(n_252), .A2(n_271), .B1(n_278), .B2(n_283), .C(n_288), .Y(n_251) );
AOI222xp33_ASAP7_75t_L g445 ( .A1(n_252), .A2(n_383), .B1(n_446), .B2(n_451), .C1(n_454), .C2(n_455), .Y(n_445) );
INVx1_ASAP7_75t_L g252 ( .A(n_253), .Y(n_252) );
NAND2x1_ASAP7_75t_L g253 ( .A(n_254), .B(n_270), .Y(n_253) );
INVx4_ASAP7_75t_R g254 ( .A(n_255), .Y(n_254) );
NAND2xp5_ASAP7_75t_L g363 ( .A(n_255), .B(n_346), .Y(n_363) );
INVx1_ASAP7_75t_L g255 ( .A(n_256), .Y(n_255) );
INVx2_ASAP7_75t_L g282 ( .A(n_256), .Y(n_282) );
NAND2xp5_ASAP7_75t_L g290 ( .A(n_256), .B(n_280), .Y(n_290) );
AND2x4_ASAP7_75t_L g351 ( .A(n_256), .B(n_352), .Y(n_351) );
AND2x4_ASAP7_75t_L g256 ( .A(n_257), .B(n_264), .Y(n_256) );
NAND2xp5_ASAP7_75t_L g257 ( .A(n_258), .B(n_260), .Y(n_257) );
AOI21xp5_ASAP7_75t_L g264 ( .A1(n_258), .A2(n_265), .B(n_269), .Y(n_264) );
AOI21xp5_ASAP7_75t_L g260 ( .A1(n_261), .A2(n_262), .B(n_263), .Y(n_260) );
INVx1_ASAP7_75t_L g306 ( .A(n_270), .Y(n_306) );
INVx1_ASAP7_75t_L g271 ( .A(n_272), .Y(n_271) );
NAND2xp5_ASAP7_75t_L g272 ( .A(n_273), .B(n_276), .Y(n_272) );
NAND3xp33_ASAP7_75t_L g458 ( .A(n_273), .B(n_459), .C(n_462), .Y(n_458) );
OR2x2_ASAP7_75t_L g474 ( .A(n_273), .B(n_462), .Y(n_474) );
INVx2_ASAP7_75t_L g273 ( .A(n_274), .Y(n_273) );
OAI21xp33_ASAP7_75t_L g419 ( .A1(n_274), .A2(n_344), .B(n_420), .Y(n_419) );
INVx1_ASAP7_75t_L g274 ( .A(n_275), .Y(n_274) );
AND2x2_ASAP7_75t_L g408 ( .A(n_275), .B(n_295), .Y(n_408) );
NAND2xp5_ASAP7_75t_L g379 ( .A(n_276), .B(n_359), .Y(n_379) );
AND2x2_ASAP7_75t_L g278 ( .A(n_279), .B(n_281), .Y(n_278) );
OR2x2_ASAP7_75t_L g422 ( .A(n_279), .B(n_291), .Y(n_422) );
INVx1_ASAP7_75t_L g279 ( .A(n_280), .Y(n_279) );
INVx1_ASAP7_75t_L g400 ( .A(n_281), .Y(n_400) );
NAND2xp5_ASAP7_75t_L g405 ( .A(n_281), .B(n_327), .Y(n_405) );
NAND2xp5_ASAP7_75t_L g410 ( .A(n_281), .B(n_411), .Y(n_410) );
HB1xp67_ASAP7_75t_L g431 ( .A(n_281), .Y(n_431) );
NAND2xp5_ASAP7_75t_L g465 ( .A(n_281), .B(n_437), .Y(n_465) );
AND2x4_ASAP7_75t_SL g300 ( .A(n_282), .B(n_301), .Y(n_300) );
NOR2x1p5_ASAP7_75t_L g283 ( .A(n_284), .B(n_285), .Y(n_283) );
BUFx3_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
INVx1_ASAP7_75t_L g358 ( .A(n_287), .Y(n_358) );
NAND2xp5_ASAP7_75t_L g448 ( .A(n_287), .B(n_449), .Y(n_448) );
AOI21xp33_ASAP7_75t_L g288 ( .A1(n_289), .A2(n_291), .B(n_292), .Y(n_288) );
HB1xp67_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
INVx4_ASAP7_75t_L g382 ( .A(n_291), .Y(n_382) );
NOR2x1_ASAP7_75t_L g479 ( .A(n_291), .B(n_471), .Y(n_479) );
INVx1_ASAP7_75t_L g292 ( .A(n_293), .Y(n_292) );
AND2x2_ASAP7_75t_L g414 ( .A(n_294), .B(n_407), .Y(n_414) );
INVx2_ASAP7_75t_L g310 ( .A(n_295), .Y(n_310) );
NAND2xp5_ASAP7_75t_SL g296 ( .A(n_297), .B(n_340), .Y(n_296) );
NOR3xp33_ASAP7_75t_L g297 ( .A(n_298), .B(n_318), .C(n_331), .Y(n_297) );
OAI322xp33_ASAP7_75t_L g298 ( .A1(n_299), .A2(n_302), .A3(n_304), .B1(n_306), .B2(n_307), .C1(n_312), .C2(n_314), .Y(n_298) );
INVx1_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
INVx1_ASAP7_75t_L g438 ( .A(n_300), .Y(n_438) );
OAI22xp5_ASAP7_75t_L g412 ( .A1(n_302), .A2(n_413), .B1(n_415), .B2(n_417), .Y(n_412) );
INVx1_ASAP7_75t_L g302 ( .A(n_303), .Y(n_302) );
NAND2xp5_ASAP7_75t_L g456 ( .A(n_303), .B(n_351), .Y(n_456) );
INVx1_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
AND2x4_ASAP7_75t_SL g320 ( .A(n_305), .B(n_321), .Y(n_320) );
AND2x2_ASAP7_75t_L g401 ( .A(n_305), .B(n_359), .Y(n_401) );
NAND2xp5_ASAP7_75t_L g477 ( .A(n_305), .B(n_336), .Y(n_477) );
INVx2_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
AND2x2_ASAP7_75t_L g433 ( .A(n_308), .B(n_374), .Y(n_433) );
AND2x2_ASAP7_75t_L g309 ( .A(n_310), .B(n_311), .Y(n_309) );
INVx1_ASAP7_75t_L g312 ( .A(n_313), .Y(n_312) );
AOI322xp5_ASAP7_75t_L g371 ( .A1(n_314), .A2(n_351), .A3(n_372), .B1(n_375), .B2(n_378), .C1(n_380), .C2(n_383), .Y(n_371) );
INVx1_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
NAND2xp33_ASAP7_75t_L g376 ( .A(n_315), .B(n_377), .Y(n_376) );
INVx2_ASAP7_75t_SL g315 ( .A(n_316), .Y(n_315) );
INVx2_ASAP7_75t_L g368 ( .A(n_316), .Y(n_368) );
OR2x2_ASAP7_75t_L g391 ( .A(n_316), .B(n_377), .Y(n_391) );
BUFx2_ASAP7_75t_L g346 ( .A(n_317), .Y(n_346) );
AOI21xp33_ASAP7_75t_L g318 ( .A1(n_319), .A2(n_322), .B(n_326), .Y(n_318) );
OAI22xp5_ASAP7_75t_L g348 ( .A1(n_319), .A2(n_349), .B1(n_355), .B2(n_356), .Y(n_348) );
INVx1_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
INVx1_ASAP7_75t_L g441 ( .A(n_321), .Y(n_441) );
INVx1_ASAP7_75t_L g322 ( .A(n_323), .Y(n_322) );
INVx2_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
OR2x2_ASAP7_75t_L g344 ( .A(n_325), .B(n_345), .Y(n_344) );
OR2x2_ASAP7_75t_L g384 ( .A(n_325), .B(n_385), .Y(n_384) );
OR2x2_ASAP7_75t_L g424 ( .A(n_325), .B(n_425), .Y(n_424) );
OR2x2_ASAP7_75t_L g440 ( .A(n_325), .B(n_441), .Y(n_440) );
OR2x2_ASAP7_75t_L g326 ( .A(n_327), .B(n_329), .Y(n_326) );
INVx1_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
NAND2xp5_ASAP7_75t_L g381 ( .A(n_328), .B(n_382), .Y(n_381) );
INVx1_ASAP7_75t_L g399 ( .A(n_328), .Y(n_399) );
OR2x2_ASAP7_75t_L g417 ( .A(n_329), .B(n_353), .Y(n_417) );
OR2x2_ASAP7_75t_L g443 ( .A(n_329), .B(n_437), .Y(n_443) );
INVx2_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
AOI21xp33_ASAP7_75t_L g331 ( .A1(n_332), .A2(n_335), .B(n_338), .Y(n_331) );
NAND2xp5_ASAP7_75t_L g332 ( .A(n_333), .B(n_334), .Y(n_332) );
NAND2xp5_ASAP7_75t_L g373 ( .A(n_333), .B(n_374), .Y(n_373) );
NAND2xp5_ASAP7_75t_L g335 ( .A(n_336), .B(n_337), .Y(n_335) );
INVx2_ASAP7_75t_L g462 ( .A(n_337), .Y(n_462) );
INVx1_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
AOI21xp5_ASAP7_75t_L g340 ( .A1(n_341), .A2(n_347), .B(n_348), .Y(n_340) );
INVx1_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
NAND2xp5_ASAP7_75t_L g342 ( .A(n_343), .B(n_346), .Y(n_342) );
INVx2_ASAP7_75t_SL g343 ( .A(n_344), .Y(n_343) );
INVx2_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
AND2x2_ASAP7_75t_L g350 ( .A(n_351), .B(n_353), .Y(n_350) );
NAND2xp5_ASAP7_75t_L g452 ( .A(n_351), .B(n_453), .Y(n_452) );
HB1xp67_ASAP7_75t_L g428 ( .A(n_352), .Y(n_428) );
HB1xp67_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
OR2x2_ASAP7_75t_L g471 ( .A(n_354), .B(n_472), .Y(n_471) );
NAND2xp5_ASAP7_75t_L g439 ( .A(n_356), .B(n_440), .Y(n_439) );
INVx2_ASAP7_75t_SL g356 ( .A(n_357), .Y(n_356) );
AND2x2_ASAP7_75t_L g357 ( .A(n_358), .B(n_359), .Y(n_357) );
INVx1_ASAP7_75t_L g394 ( .A(n_358), .Y(n_394) );
NAND2xp5_ASAP7_75t_L g393 ( .A(n_359), .B(n_394), .Y(n_393) );
INVx2_ASAP7_75t_L g425 ( .A(n_359), .Y(n_425) );
NAND2xp5_ASAP7_75t_L g426 ( .A(n_361), .B(n_427), .Y(n_426) );
INVx1_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
INVx1_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
INVx1_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
NAND2xp5_ASAP7_75t_L g366 ( .A(n_367), .B(n_368), .Y(n_366) );
INVx1_ASAP7_75t_L g444 ( .A(n_367), .Y(n_444) );
NAND3xp33_ASAP7_75t_L g460 ( .A(n_367), .B(n_382), .C(n_461), .Y(n_460) );
INVx1_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
INVx1_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
INVxp67_ASAP7_75t_SL g375 ( .A(n_376), .Y(n_375) );
INVx1_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
INVx1_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
INVx1_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
OR2x2_ASAP7_75t_L g481 ( .A(n_385), .B(n_482), .Y(n_481) );
INVx1_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
NOR3xp33_ASAP7_75t_SL g387 ( .A(n_388), .B(n_429), .C(n_457), .Y(n_387) );
NAND3xp33_ASAP7_75t_SL g388 ( .A(n_389), .B(n_402), .C(n_418), .Y(n_388) );
AOI22xp5_ASAP7_75t_L g389 ( .A1(n_390), .A2(n_392), .B1(n_397), .B2(n_401), .Y(n_389) );
INVx1_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
NAND2xp5_ASAP7_75t_L g392 ( .A(n_393), .B(n_395), .Y(n_392) );
INVx1_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
AOI22xp33_ASAP7_75t_SL g463 ( .A1(n_396), .A2(n_464), .B1(n_466), .B2(n_467), .Y(n_463) );
INVx1_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
OR2x2_ASAP7_75t_L g398 ( .A(n_399), .B(n_400), .Y(n_398) );
AOI221xp5_ASAP7_75t_L g402 ( .A1(n_403), .A2(n_404), .B1(n_406), .B2(n_409), .C(n_412), .Y(n_402) );
INVx1_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
INVx1_ASAP7_75t_L g420 ( .A(n_406), .Y(n_420) );
AND2x2_ASAP7_75t_L g406 ( .A(n_407), .B(n_408), .Y(n_406) );
INVx2_ASAP7_75t_L g450 ( .A(n_408), .Y(n_450) );
INVxp67_ASAP7_75t_SL g409 ( .A(n_410), .Y(n_409) );
INVx2_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
INVxp33_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
INVx1_ASAP7_75t_L g478 ( .A(n_417), .Y(n_478) );
AOI22xp33_ASAP7_75t_L g418 ( .A1(n_419), .A2(n_421), .B1(n_423), .B2(n_426), .Y(n_418) );
INVx1_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
INVx2_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
OAI211xp5_ASAP7_75t_SL g429 ( .A1(n_430), .A2(n_432), .B(n_434), .C(n_445), .Y(n_429) );
INVx1_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
INVx1_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
AOI22xp5_ASAP7_75t_L g434 ( .A1(n_433), .A2(n_435), .B1(n_439), .B2(n_442), .Y(n_434) );
INVx2_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
OR2x2_ASAP7_75t_L g436 ( .A(n_437), .B(n_438), .Y(n_436) );
INVx1_ASAP7_75t_L g461 ( .A(n_437), .Y(n_461) );
NAND2xp5_ASAP7_75t_SL g442 ( .A(n_443), .B(n_444), .Y(n_442) );
INVx2_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
OR2x2_ASAP7_75t_L g447 ( .A(n_448), .B(n_450), .Y(n_447) );
INVxp67_ASAP7_75t_SL g454 ( .A(n_448), .Y(n_454) );
INVx1_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
INVxp67_ASAP7_75t_SL g455 ( .A(n_456), .Y(n_455) );
NAND4xp25_ASAP7_75t_L g457 ( .A(n_458), .B(n_463), .C(n_468), .D(n_475), .Y(n_457) );
INVx1_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
INVx1_ASAP7_75t_L g464 ( .A(n_465), .Y(n_464) );
NAND2xp5_ASAP7_75t_L g468 ( .A(n_469), .B(n_473), .Y(n_468) );
HB1xp67_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
INVx1_ASAP7_75t_L g470 ( .A(n_471), .Y(n_470) );
INVxp67_ASAP7_75t_SL g473 ( .A(n_474), .Y(n_473) );
AOI22xp33_ASAP7_75t_L g475 ( .A1(n_476), .A2(n_478), .B1(n_479), .B2(n_480), .Y(n_475) );
INVx1_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
INVx2_ASAP7_75t_L g480 ( .A(n_481), .Y(n_480) );
CKINVDCx6p67_ASAP7_75t_R g483 ( .A(n_484), .Y(n_483) );
CKINVDCx20_ASAP7_75t_R g484 ( .A(n_485), .Y(n_484) );
AND2x2_ASAP7_75t_L g485 ( .A(n_486), .B(n_487), .Y(n_485) );
INVxp67_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
AO21x2_ASAP7_75t_L g714 ( .A1(n_488), .A2(n_661), .B(n_715), .Y(n_714) );
NAND2xp5_ASAP7_75t_L g488 ( .A(n_489), .B(n_490), .Y(n_488) );
INVx1_ASAP7_75t_L g490 ( .A(n_491), .Y(n_490) );
INVx1_ASAP7_75t_L g491 ( .A(n_492), .Y(n_491) );
OAI221xp5_ASAP7_75t_L g493 ( .A1(n_494), .A2(n_495), .B1(n_655), .B2(n_665), .C(n_708), .Y(n_493) );
AOI22xp5_ASAP7_75t_L g708 ( .A1(n_495), .A2(n_701), .B1(n_709), .B2(n_712), .Y(n_708) );
AND3x2_ASAP7_75t_L g495 ( .A(n_496), .B(n_573), .C(n_631), .Y(n_495) );
OAI31xp33_ASAP7_75t_SL g496 ( .A1(n_497), .A2(n_509), .A3(n_552), .B(n_570), .Y(n_496) );
OR2x2_ASAP7_75t_L g498 ( .A(n_499), .B(n_502), .Y(n_498) );
INVx1_ASAP7_75t_L g513 ( .A(n_499), .Y(n_513) );
INVx1_ASAP7_75t_L g554 ( .A(n_499), .Y(n_554) );
INVx1_ASAP7_75t_L g499 ( .A(n_500), .Y(n_499) );
AND2x2_ASAP7_75t_L g537 ( .A(n_501), .B(n_538), .Y(n_537) );
OR2x6_ASAP7_75t_L g506 ( .A(n_502), .B(n_507), .Y(n_506) );
BUFx6f_ASAP7_75t_L g502 ( .A(n_503), .Y(n_502) );
NAND2xp5_ASAP7_75t_L g503 ( .A(n_504), .B(n_505), .Y(n_503) );
AND2x4_ASAP7_75t_L g519 ( .A(n_504), .B(n_520), .Y(n_519) );
INVx2_ASAP7_75t_L g526 ( .A(n_504), .Y(n_526) );
INVx2_ASAP7_75t_L g520 ( .A(n_505), .Y(n_520) );
INVx2_ASAP7_75t_L g527 ( .A(n_505), .Y(n_527) );
INVx1_ASAP7_75t_L g561 ( .A(n_507), .Y(n_561) );
INVx1_ASAP7_75t_L g507 ( .A(n_508), .Y(n_507) );
AND2x2_ASAP7_75t_L g563 ( .A(n_508), .B(n_564), .Y(n_563) );
AND2x2_ASAP7_75t_L g566 ( .A(n_508), .B(n_567), .Y(n_566) );
NAND3xp33_ASAP7_75t_L g509 ( .A(n_510), .B(n_521), .C(n_539), .Y(n_509) );
AOI22xp33_ASAP7_75t_L g510 ( .A1(n_511), .A2(n_512), .B1(n_516), .B2(n_517), .Y(n_510) );
AND2x4_ASAP7_75t_L g512 ( .A(n_513), .B(n_514), .Y(n_512) );
AND2x2_ASAP7_75t_L g517 ( .A(n_513), .B(n_518), .Y(n_517) );
BUFx4f_ASAP7_75t_L g514 ( .A(n_515), .Y(n_514) );
BUFx6f_ASAP7_75t_L g530 ( .A(n_515), .Y(n_530) );
OAI221xp5_ASAP7_75t_L g643 ( .A1(n_516), .A2(n_522), .B1(n_644), .B2(n_647), .C(n_649), .Y(n_643) );
BUFx6f_ASAP7_75t_L g518 ( .A(n_519), .Y(n_518) );
INVx5_ASAP7_75t_L g546 ( .A(n_519), .Y(n_546) );
INVx1_ASAP7_75t_L g535 ( .A(n_520), .Y(n_535) );
OAI211xp5_ASAP7_75t_L g521 ( .A1(n_522), .A2(n_523), .B(n_528), .C(n_531), .Y(n_521) );
BUFx6f_ASAP7_75t_L g523 ( .A(n_524), .Y(n_523) );
BUFx12f_ASAP7_75t_L g524 ( .A(n_525), .Y(n_524) );
BUFx6f_ASAP7_75t_L g542 ( .A(n_525), .Y(n_542) );
NAND2x1p5_ASAP7_75t_L g525 ( .A(n_526), .B(n_527), .Y(n_525) );
AND2x4_ASAP7_75t_L g556 ( .A(n_526), .B(n_527), .Y(n_556) );
INVx1_ASAP7_75t_L g568 ( .A(n_526), .Y(n_568) );
BUFx3_ASAP7_75t_L g564 ( .A(n_527), .Y(n_564) );
BUFx12f_ASAP7_75t_SL g529 ( .A(n_530), .Y(n_529) );
BUFx3_ASAP7_75t_L g544 ( .A(n_530), .Y(n_544) );
BUFx2_ASAP7_75t_L g532 ( .A(n_533), .Y(n_532) );
INVx5_ASAP7_75t_L g549 ( .A(n_533), .Y(n_549) );
AND2x4_ASAP7_75t_L g533 ( .A(n_534), .B(n_535), .Y(n_533) );
INVx2_ASAP7_75t_L g536 ( .A(n_537), .Y(n_536) );
OAI211xp5_ASAP7_75t_L g539 ( .A1(n_540), .A2(n_541), .B(n_543), .C(n_547), .Y(n_539) );
AOI22xp5_ASAP7_75t_L g596 ( .A1(n_540), .A2(n_565), .B1(n_597), .B2(n_605), .Y(n_596) );
HB1xp67_ASAP7_75t_L g541 ( .A(n_542), .Y(n_541) );
INVx3_ASAP7_75t_L g545 ( .A(n_546), .Y(n_545) );
INVx2_ASAP7_75t_L g548 ( .A(n_549), .Y(n_548) );
BUFx4_ASAP7_75t_L g550 ( .A(n_551), .Y(n_550) );
NAND2x1p5_ASAP7_75t_L g553 ( .A(n_554), .B(n_555), .Y(n_553) );
BUFx4f_ASAP7_75t_L g555 ( .A(n_556), .Y(n_555) );
INVx2_ASAP7_75t_L g560 ( .A(n_556), .Y(n_560) );
BUFx2_ASAP7_75t_L g557 ( .A(n_558), .Y(n_557) );
NAND2xp5_ASAP7_75t_L g558 ( .A(n_559), .B(n_561), .Y(n_558) );
INVx1_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
AOI22xp33_ASAP7_75t_L g562 ( .A1(n_563), .A2(n_565), .B1(n_566), .B2(n_569), .Y(n_562) );
INVx1_ASAP7_75t_L g567 ( .A(n_568), .Y(n_567) );
AO22x1_ASAP7_75t_L g574 ( .A1(n_569), .A2(n_575), .B1(n_576), .B2(n_589), .Y(n_574) );
INVx1_ASAP7_75t_L g570 ( .A(n_571), .Y(n_570) );
INVx2_ASAP7_75t_L g571 ( .A(n_572), .Y(n_571) );
OR2x2_ASAP7_75t_L g578 ( .A(n_572), .B(n_579), .Y(n_578) );
INVx1_ASAP7_75t_L g599 ( .A(n_572), .Y(n_599) );
INVx2_ASAP7_75t_L g625 ( .A(n_572), .Y(n_625) );
NOR2xp33_ASAP7_75t_L g573 ( .A(n_574), .B(n_595), .Y(n_573) );
AND2x4_ASAP7_75t_L g576 ( .A(n_577), .B(n_582), .Y(n_576) );
AND2x2_ASAP7_75t_L g589 ( .A(n_577), .B(n_590), .Y(n_589) );
AND2x2_ASAP7_75t_L g632 ( .A(n_577), .B(n_618), .Y(n_632) );
INVx2_ASAP7_75t_L g577 ( .A(n_578), .Y(n_577) );
OR2x6_ASAP7_75t_L g635 ( .A(n_578), .B(n_636), .Y(n_635) );
OR2x6_ASAP7_75t_L g579 ( .A(n_580), .B(n_581), .Y(n_579) );
INVx1_ASAP7_75t_L g601 ( .A(n_580), .Y(n_601) );
BUFx2_ASAP7_75t_L g627 ( .A(n_580), .Y(n_627) );
AND2x2_ASAP7_75t_L g600 ( .A(n_581), .B(n_601), .Y(n_600) );
INVx1_ASAP7_75t_L g628 ( .A(n_581), .Y(n_628) );
AND2x4_ASAP7_75t_L g642 ( .A(n_581), .B(n_627), .Y(n_642) );
OR2x2_ASAP7_75t_L g692 ( .A(n_581), .B(n_601), .Y(n_692) );
INVx1_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
INVx1_ASAP7_75t_L g583 ( .A(n_584), .Y(n_583) );
BUFx3_ASAP7_75t_L g584 ( .A(n_585), .Y(n_584) );
INVx4_ASAP7_75t_L g623 ( .A(n_585), .Y(n_623) );
BUFx6f_ASAP7_75t_L g648 ( .A(n_585), .Y(n_648) );
AND2x4_ASAP7_75t_L g585 ( .A(n_586), .B(n_587), .Y(n_585) );
INVx1_ASAP7_75t_L g608 ( .A(n_586), .Y(n_608) );
AND2x4_ASAP7_75t_L g637 ( .A(n_586), .B(n_604), .Y(n_637) );
AND2x4_ASAP7_75t_L g592 ( .A(n_587), .B(n_593), .Y(n_592) );
INVx2_ASAP7_75t_L g587 ( .A(n_588), .Y(n_587) );
AND2x2_ASAP7_75t_L g613 ( .A(n_588), .B(n_594), .Y(n_613) );
AND2x2_ASAP7_75t_L g620 ( .A(n_588), .B(n_593), .Y(n_620) );
BUFx6f_ASAP7_75t_L g590 ( .A(n_591), .Y(n_590) );
BUFx6f_ASAP7_75t_L g591 ( .A(n_592), .Y(n_591) );
INVx2_ASAP7_75t_L g616 ( .A(n_592), .Y(n_616) );
BUFx6f_ASAP7_75t_L g630 ( .A(n_592), .Y(n_630) );
INVx2_ASAP7_75t_L g593 ( .A(n_594), .Y(n_593) );
NAND2xp5_ASAP7_75t_L g595 ( .A(n_596), .B(n_609), .Y(n_595) );
AND2x2_ASAP7_75t_L g597 ( .A(n_598), .B(n_602), .Y(n_597) );
AND2x4_ASAP7_75t_L g605 ( .A(n_598), .B(n_606), .Y(n_605) );
AND2x4_ASAP7_75t_L g629 ( .A(n_598), .B(n_630), .Y(n_629) );
INVx2_ASAP7_75t_L g654 ( .A(n_598), .Y(n_654) );
AND2x4_ASAP7_75t_L g598 ( .A(n_599), .B(n_600), .Y(n_598) );
AND2x6_ASAP7_75t_L g641 ( .A(n_599), .B(n_642), .Y(n_641) );
INVx1_ASAP7_75t_L g700 ( .A(n_600), .Y(n_700) );
INVx2_ASAP7_75t_L g602 ( .A(n_603), .Y(n_602) );
HB1xp67_ASAP7_75t_L g603 ( .A(n_604), .Y(n_603) );
AND2x2_ASAP7_75t_L g646 ( .A(n_604), .B(n_608), .Y(n_646) );
INVx1_ASAP7_75t_L g690 ( .A(n_604), .Y(n_690) );
INVx1_ASAP7_75t_L g606 ( .A(n_607), .Y(n_606) );
INVx1_ASAP7_75t_L g607 ( .A(n_608), .Y(n_607) );
AOI31xp33_ASAP7_75t_L g609 ( .A1(n_610), .A2(n_617), .A3(n_624), .B(n_629), .Y(n_609) );
INVx3_ASAP7_75t_L g611 ( .A(n_612), .Y(n_611) );
INVx2_ASAP7_75t_L g612 ( .A(n_613), .Y(n_612) );
BUFx6f_ASAP7_75t_L g650 ( .A(n_613), .Y(n_650) );
INVx2_ASAP7_75t_SL g614 ( .A(n_615), .Y(n_614) );
BUFx3_ASAP7_75t_L g615 ( .A(n_616), .Y(n_615) );
INVx5_ASAP7_75t_L g618 ( .A(n_619), .Y(n_618) );
INVx3_ASAP7_75t_L g619 ( .A(n_620), .Y(n_619) );
INVx2_ASAP7_75t_L g621 ( .A(n_622), .Y(n_621) );
BUFx2_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
AND2x6_ASAP7_75t_L g624 ( .A(n_625), .B(n_626), .Y(n_624) );
AND2x2_ASAP7_75t_L g626 ( .A(n_627), .B(n_628), .Y(n_626) );
INVx3_ASAP7_75t_L g652 ( .A(n_630), .Y(n_652) );
AOI221xp5_ASAP7_75t_L g631 ( .A1(n_632), .A2(n_633), .B1(n_634), .B2(n_638), .C(n_639), .Y(n_631) );
CKINVDCx5p33_ASAP7_75t_R g634 ( .A(n_635), .Y(n_634) );
OR2x2_ASAP7_75t_L g653 ( .A(n_636), .B(n_654), .Y(n_653) );
INVx8_ASAP7_75t_L g636 ( .A(n_637), .Y(n_636) );
CKINVDCx8_ASAP7_75t_R g640 ( .A(n_641), .Y(n_640) );
INVx2_ASAP7_75t_L g644 ( .A(n_645), .Y(n_644) );
BUFx6f_ASAP7_75t_L g645 ( .A(n_646), .Y(n_645) );
INVx2_ASAP7_75t_SL g647 ( .A(n_648), .Y(n_647) );
INVx2_ASAP7_75t_L g651 ( .A(n_652), .Y(n_651) );
CKINVDCx16_ASAP7_75t_R g655 ( .A(n_656), .Y(n_655) );
CKINVDCx16_ASAP7_75t_R g656 ( .A(n_657), .Y(n_656) );
HB1xp67_ASAP7_75t_SL g657 ( .A(n_658), .Y(n_657) );
BUFx6f_ASAP7_75t_L g658 ( .A(n_659), .Y(n_658) );
NAND2xp5_ASAP7_75t_L g659 ( .A(n_660), .B(n_663), .Y(n_659) );
INVx1_ASAP7_75t_L g660 ( .A(n_661), .Y(n_660) );
BUFx2_ASAP7_75t_L g661 ( .A(n_662), .Y(n_661) );
INVx1_ASAP7_75t_L g685 ( .A(n_662), .Y(n_685) );
AND2x2_ASAP7_75t_L g715 ( .A(n_663), .B(n_716), .Y(n_715) );
INVx1_ASAP7_75t_L g663 ( .A(n_664), .Y(n_663) );
NAND2xp5_ASAP7_75t_L g684 ( .A(n_664), .B(n_685), .Y(n_684) );
AOI22xp33_ASAP7_75t_L g665 ( .A1(n_666), .A2(n_679), .B1(n_701), .B2(n_702), .Y(n_665) );
OAI22xp5_ASAP7_75t_L g709 ( .A1(n_666), .A2(n_701), .B1(n_710), .B2(n_711), .Y(n_709) );
XOR2xp5_ASAP7_75t_L g666 ( .A(n_667), .B(n_672), .Y(n_666) );
XNOR2xp5_ASAP7_75t_L g667 ( .A(n_668), .B(n_670), .Y(n_667) );
INVx1_ASAP7_75t_L g668 ( .A(n_669), .Y(n_668) );
INVx1_ASAP7_75t_L g670 ( .A(n_671), .Y(n_670) );
AOI22xp5_ASAP7_75t_L g672 ( .A1(n_673), .A2(n_674), .B1(n_675), .B2(n_676), .Y(n_672) );
INVx1_ASAP7_75t_L g673 ( .A(n_674), .Y(n_673) );
INVx1_ASAP7_75t_L g675 ( .A(n_676), .Y(n_675) );
INVx3_ASAP7_75t_L g679 ( .A(n_680), .Y(n_679) );
BUFx3_ASAP7_75t_L g680 ( .A(n_681), .Y(n_680) );
INVx5_ASAP7_75t_L g681 ( .A(n_682), .Y(n_681) );
CKINVDCx16_ASAP7_75t_R g710 ( .A(n_682), .Y(n_710) );
AND2x6_ASAP7_75t_L g682 ( .A(n_683), .B(n_693), .Y(n_682) );
NOR2xp33_ASAP7_75t_L g683 ( .A(n_684), .B(n_686), .Y(n_683) );
INVxp67_ASAP7_75t_L g706 ( .A(n_684), .Y(n_706) );
INVx1_ASAP7_75t_L g716 ( .A(n_685), .Y(n_716) );
INVxp67_ASAP7_75t_SL g686 ( .A(n_687), .Y(n_686) );
NAND2xp5_ASAP7_75t_L g707 ( .A(n_687), .B(n_697), .Y(n_707) );
NAND3xp33_ASAP7_75t_L g687 ( .A(n_688), .B(n_690), .C(n_691), .Y(n_687) );
INVx2_ASAP7_75t_L g688 ( .A(n_689), .Y(n_688) );
CKINVDCx11_ASAP7_75t_R g695 ( .A(n_689), .Y(n_695) );
AND2x4_ASAP7_75t_L g698 ( .A(n_690), .B(n_699), .Y(n_698) );
BUFx6f_ASAP7_75t_L g691 ( .A(n_692), .Y(n_691) );
NAND2xp5_ASAP7_75t_L g693 ( .A(n_694), .B(n_696), .Y(n_693) );
CKINVDCx5p33_ASAP7_75t_R g694 ( .A(n_695), .Y(n_694) );
INVx2_ASAP7_75t_SL g696 ( .A(n_697), .Y(n_696) );
INVx2_ASAP7_75t_SL g697 ( .A(n_698), .Y(n_697) );
INVx1_ASAP7_75t_L g699 ( .A(n_700), .Y(n_699) );
INVx2_ASAP7_75t_L g702 ( .A(n_703), .Y(n_702) );
BUFx4f_ASAP7_75t_SL g703 ( .A(n_704), .Y(n_703) );
BUFx6f_ASAP7_75t_L g711 ( .A(n_704), .Y(n_711) );
INVx4_ASAP7_75t_L g704 ( .A(n_705), .Y(n_704) );
AND2x2_ASAP7_75t_L g705 ( .A(n_706), .B(n_707), .Y(n_705) );
CKINVDCx20_ASAP7_75t_R g712 ( .A(n_713), .Y(n_712) );
CKINVDCx20_ASAP7_75t_R g713 ( .A(n_714), .Y(n_713) );
endmodule