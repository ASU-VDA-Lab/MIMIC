module fake_jpeg_24860_n_131 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_131);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_131;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_11),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_11),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_10),
.Y(n_16)
);

BUFx4f_ASAP7_75t_SL g17 ( 
.A(n_8),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_5),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

INVx11_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_2),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_5),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_1),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_7),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_4),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_20),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_29),
.B(n_33),
.Y(n_43)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_17),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_30),
.B(n_31),
.Y(n_54)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_17),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_19),
.B(n_0),
.Y(n_32)
);

AND2x2_ASAP7_75t_L g52 ( 
.A(n_32),
.B(n_37),
.Y(n_52)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_20),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_L g34 ( 
.A1(n_21),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_34)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_34),
.A2(n_42),
.B1(n_24),
.B2(n_22),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_17),
.Y(n_35)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_35),
.Y(n_56)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_27),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_36),
.B(n_38),
.Y(n_44)
);

NAND2xp33_ASAP7_75t_SL g37 ( 
.A(n_21),
.B(n_1),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_14),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_27),
.Y(n_39)
);

INVx5_ASAP7_75t_L g51 ( 
.A(n_39),
.Y(n_51)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_19),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_40),
.B(n_41),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_22),
.Y(n_41)
);

OAI22xp33_ASAP7_75t_SL g42 ( 
.A1(n_14),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_42)
);

AOI21xp5_ASAP7_75t_L g80 ( 
.A1(n_45),
.A2(n_55),
.B(n_44),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_41),
.B(n_16),
.Y(n_47)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_47),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_39),
.Y(n_48)
);

CKINVDCx16_ASAP7_75t_R g66 ( 
.A(n_48),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_32),
.B(n_16),
.Y(n_49)
);

CKINVDCx16_ASAP7_75t_R g70 ( 
.A(n_49),
.Y(n_70)
);

OR2x2_ASAP7_75t_L g50 ( 
.A(n_37),
.B(n_15),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_SL g81 ( 
.A(n_50),
.B(n_61),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_34),
.B(n_28),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_53),
.B(n_25),
.Y(n_67)
);

MAJIxp5_ASAP7_75t_L g55 ( 
.A(n_30),
.B(n_24),
.C(n_28),
.Y(n_55)
);

MAJIxp5_ASAP7_75t_L g68 ( 
.A(n_55),
.B(n_23),
.C(n_18),
.Y(n_68)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_35),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_57),
.B(n_62),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_38),
.B(n_26),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_58),
.B(n_60),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_36),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_59),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_31),
.B(n_26),
.Y(n_60)
);

AND2x2_ASAP7_75t_L g61 ( 
.A(n_35),
.B(n_40),
.Y(n_61)
);

OAI21xp5_ASAP7_75t_SL g74 ( 
.A1(n_61),
.A2(n_3),
.B(n_6),
.Y(n_74)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_29),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_33),
.B(n_25),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_63),
.B(n_15),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_67),
.A2(n_79),
.B1(n_80),
.B2(n_54),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_68),
.B(n_73),
.Y(n_85)
);

XNOR2xp5_ASAP7_75t_L g69 ( 
.A(n_52),
.B(n_23),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_69),
.B(n_71),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_52),
.B(n_18),
.Y(n_71)
);

OAI21xp5_ASAP7_75t_SL g91 ( 
.A1(n_74),
.A2(n_78),
.B(n_43),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_52),
.B(n_7),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_75),
.B(n_61),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_46),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_76),
.B(n_65),
.Y(n_87)
);

MAJx2_ASAP7_75t_L g78 ( 
.A(n_50),
.B(n_9),
.C(n_12),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_53),
.A2(n_9),
.B1(n_12),
.B2(n_13),
.Y(n_79)
);

CKINVDCx14_ASAP7_75t_R g83 ( 
.A(n_81),
.Y(n_83)
);

INVx2_ASAP7_75t_SL g82 ( 
.A(n_66),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_82),
.B(n_89),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_67),
.A2(n_51),
.B1(n_62),
.B2(n_56),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_86),
.A2(n_51),
.B1(n_56),
.B2(n_72),
.Y(n_99)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_87),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_88),
.B(n_93),
.Y(n_98)
);

CKINVDCx16_ASAP7_75t_R g89 ( 
.A(n_77),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_65),
.B(n_54),
.Y(n_90)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_90),
.Y(n_103)
);

AND2x2_ASAP7_75t_L g96 ( 
.A(n_91),
.B(n_95),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_64),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_92),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_79),
.B(n_68),
.Y(n_93)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_71),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_94),
.B(n_75),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_97),
.B(n_104),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_L g111 ( 
.A1(n_99),
.A2(n_72),
.B1(n_57),
.B2(n_105),
.Y(n_111)
);

XOR2xp5_ASAP7_75t_L g100 ( 
.A(n_95),
.B(n_69),
.Y(n_100)
);

XOR2xp5_ASAP7_75t_L g108 ( 
.A(n_100),
.B(n_101),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_84),
.B(n_80),
.C(n_78),
.Y(n_101)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_86),
.Y(n_104)
);

XOR2xp5_ASAP7_75t_L g109 ( 
.A(n_100),
.B(n_101),
.Y(n_109)
);

XNOR2xp5_ASAP7_75t_L g115 ( 
.A(n_109),
.B(n_113),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_104),
.A2(n_83),
.B1(n_94),
.B2(n_91),
.Y(n_110)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_110),
.Y(n_118)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_111),
.Y(n_119)
);

AND2x2_ASAP7_75t_L g112 ( 
.A(n_97),
.B(n_84),
.Y(n_112)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_112),
.Y(n_120)
);

XNOR2xp5_ASAP7_75t_L g113 ( 
.A(n_96),
.B(n_98),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_103),
.B(n_82),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_114),
.Y(n_117)
);

XNOR2xp5_ASAP7_75t_L g116 ( 
.A(n_108),
.B(n_96),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_116),
.B(n_109),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_SL g121 ( 
.A1(n_118),
.A2(n_107),
.B(n_106),
.Y(n_121)
);

XOR2xp5_ASAP7_75t_L g127 ( 
.A(n_121),
.B(n_122),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_119),
.A2(n_92),
.B1(n_102),
.B2(n_113),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_123),
.A2(n_124),
.B1(n_120),
.B2(n_85),
.Y(n_125)
);

A2O1A1Ixp33_ASAP7_75t_SL g124 ( 
.A1(n_117),
.A2(n_112),
.B(n_108),
.C(n_74),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_125),
.B(n_82),
.C(n_59),
.Y(n_129)
);

AOI31xp67_ASAP7_75t_L g126 ( 
.A1(n_124),
.A2(n_116),
.A3(n_115),
.B(n_70),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_126),
.B(n_115),
.Y(n_128)
);

NOR3xp33_ASAP7_75t_L g130 ( 
.A(n_128),
.B(n_129),
.C(n_127),
.Y(n_130)
);

XNOR2xp5_ASAP7_75t_L g131 ( 
.A(n_130),
.B(n_48),
.Y(n_131)
);


endmodule