module fake_jpeg_10984_n_61 (n_13, n_21, n_1, n_10, n_6, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_61);

input n_13;
input n_21;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_61;

wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_45;
wire n_23;
wire n_27;
wire n_55;
wire n_47;
wire n_22;
wire n_51;
wire n_40;
wire n_59;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_24;
wire n_28;
wire n_44;
wire n_26;
wire n_38;
wire n_36;
wire n_31;
wire n_25;
wire n_56;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_32;

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_21),
.Y(n_22)
);

AND2x2_ASAP7_75t_L g23 ( 
.A(n_2),
.B(n_8),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_18),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_16),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

BUFx2_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_27),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_29),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_SL g30 ( 
.A1(n_27),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_30)
);

AOI22xp5_ASAP7_75t_L g41 ( 
.A1(n_30),
.A2(n_33),
.B1(n_23),
.B2(n_28),
.Y(n_41)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_26),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_31),
.B(n_24),
.Y(n_37)
);

INVx2_ASAP7_75t_SL g32 ( 
.A(n_23),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_SL g36 ( 
.A(n_32),
.B(n_34),
.Y(n_36)
);

AOI22xp33_ASAP7_75t_SL g33 ( 
.A1(n_28),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_33)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_25),
.Y(n_34)
);

AND2x4_ASAP7_75t_SL g35 ( 
.A(n_32),
.B(n_25),
.Y(n_35)
);

AND2x2_ASAP7_75t_L g47 ( 
.A(n_35),
.B(n_41),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_37),
.B(n_22),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_31),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_SL g46 ( 
.A(n_39),
.B(n_40),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_34),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_L g42 ( 
.A1(n_36),
.A2(n_30),
.B1(n_29),
.B2(n_32),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_L g50 ( 
.A1(n_42),
.A2(n_48),
.B1(n_47),
.B2(n_46),
.Y(n_50)
);

MAJIxp5_ASAP7_75t_L g51 ( 
.A(n_43),
.B(n_44),
.C(n_4),
.Y(n_51)
);

AOI22x1_ASAP7_75t_L g44 ( 
.A1(n_35),
.A2(n_38),
.B1(n_23),
.B2(n_14),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_38),
.Y(n_45)
);

INVxp67_ASAP7_75t_L g49 ( 
.A(n_45),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_SL g48 ( 
.A(n_35),
.B(n_3),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_L g54 ( 
.A1(n_50),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_54)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_51),
.Y(n_56)
);

XOR2x2_ASAP7_75t_L g52 ( 
.A(n_47),
.B(n_43),
.Y(n_52)
);

XOR2xp5_ASAP7_75t_L g55 ( 
.A(n_52),
.B(n_53),
.Y(n_55)
);

XOR2xp5_ASAP7_75t_L g53 ( 
.A(n_47),
.B(n_13),
.Y(n_53)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_54),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_57),
.B(n_49),
.Y(n_58)
);

AOI322xp5_ASAP7_75t_L g59 ( 
.A1(n_58),
.A2(n_56),
.A3(n_52),
.B1(n_55),
.B2(n_5),
.C1(n_6),
.C2(n_7),
.Y(n_59)
);

AOI322xp5_ASAP7_75t_L g60 ( 
.A1(n_59),
.A2(n_55),
.A3(n_11),
.B1(n_15),
.B2(n_17),
.C1(n_10),
.C2(n_20),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_60),
.B(n_19),
.Y(n_61)
);


endmodule