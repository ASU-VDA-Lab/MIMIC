module fake_jpeg_20113_n_211 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_211);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_211;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx5_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_1),
.B(n_3),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

BUFx16f_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_6),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_12),
.Y(n_22)
);

INVx5_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_16),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_1),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

INVx1_ASAP7_75t_SL g27 ( 
.A(n_0),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_14),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_2),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_15),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_11),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_5),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_28),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_36),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_28),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_37),
.Y(n_64)
);

HB1xp67_ASAP7_75t_L g38 ( 
.A(n_20),
.Y(n_38)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_38),
.Y(n_51)
);

INVx2_ASAP7_75t_SL g39 ( 
.A(n_19),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_39),
.B(n_40),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_18),
.B(n_0),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_35),
.Y(n_41)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_41),
.Y(n_71)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_20),
.Y(n_42)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_42),
.Y(n_52)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_35),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_43),
.B(n_32),
.Y(n_74)
);

INVx11_ASAP7_75t_SL g44 ( 
.A(n_17),
.Y(n_44)
);

INVx11_ASAP7_75t_L g61 ( 
.A(n_44),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_28),
.Y(n_45)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_45),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_29),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_46),
.A2(n_27),
.B1(n_21),
.B2(n_25),
.Y(n_53)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_17),
.Y(n_47)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_47),
.Y(n_56)
);

INVx11_ASAP7_75t_L g48 ( 
.A(n_20),
.Y(n_48)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_48),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_26),
.Y(n_49)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_49),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_SL g50 ( 
.A(n_40),
.B(n_18),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_SL g80 ( 
.A(n_50),
.B(n_54),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_53),
.A2(n_39),
.B1(n_25),
.B2(n_46),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_SL g54 ( 
.A(n_41),
.B(n_33),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_43),
.B(n_33),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_57),
.B(n_59),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_L g58 ( 
.A1(n_47),
.A2(n_27),
.B1(n_23),
.B2(n_29),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_58),
.A2(n_62),
.B1(n_24),
.B2(n_49),
.Y(n_84)
);

INVx5_ASAP7_75t_L g59 ( 
.A(n_48),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_L g62 ( 
.A1(n_47),
.A2(n_23),
.B1(n_32),
.B2(n_21),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_36),
.B(n_19),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_65),
.B(n_66),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_36),
.B(n_19),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_42),
.B(n_30),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_67),
.B(n_70),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_SL g69 ( 
.A(n_39),
.B(n_30),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g98 ( 
.A(n_69),
.B(n_74),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_42),
.B(n_22),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_48),
.B(n_22),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_73),
.B(n_20),
.Y(n_85)
);

CKINVDCx14_ASAP7_75t_R g75 ( 
.A(n_74),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_75),
.B(n_81),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_L g108 ( 
.A1(n_77),
.A2(n_88),
.B(n_51),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_65),
.A2(n_39),
.B1(n_45),
.B2(n_37),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_78),
.A2(n_92),
.B1(n_93),
.B2(n_97),
.Y(n_105)
);

INVx1_ASAP7_75t_SL g81 ( 
.A(n_52),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_54),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_82),
.B(n_84),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_85),
.B(n_91),
.Y(n_106)
);

AND2x2_ASAP7_75t_SL g86 ( 
.A(n_71),
.B(n_45),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_86),
.B(n_95),
.Y(n_114)
);

OR2x2_ASAP7_75t_SL g87 ( 
.A(n_68),
.B(n_19),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_SL g107 ( 
.A(n_87),
.B(n_55),
.Y(n_107)
);

AOI21xp5_ASAP7_75t_L g88 ( 
.A1(n_66),
.A2(n_38),
.B(n_49),
.Y(n_88)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_72),
.Y(n_89)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_89),
.Y(n_113)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_68),
.B(n_37),
.Y(n_90)
);

INVx1_ASAP7_75t_SL g100 ( 
.A(n_90),
.Y(n_100)
);

INVx5_ASAP7_75t_L g91 ( 
.A(n_56),
.Y(n_91)
);

OAI22xp33_ASAP7_75t_L g92 ( 
.A1(n_63),
.A2(n_45),
.B1(n_37),
.B2(n_36),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_71),
.A2(n_24),
.B1(n_34),
.B2(n_26),
.Y(n_93)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_56),
.Y(n_94)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_94),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_50),
.B(n_34),
.Y(n_95)
);

XOR2xp5_ASAP7_75t_L g96 ( 
.A(n_69),
.B(n_31),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_96),
.B(n_31),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_55),
.A2(n_26),
.B1(n_34),
.B2(n_4),
.Y(n_97)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_60),
.Y(n_99)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_99),
.Y(n_112)
);

AND2x2_ASAP7_75t_L g132 ( 
.A(n_101),
.B(n_96),
.Y(n_132)
);

INVx1_ASAP7_75t_SL g102 ( 
.A(n_86),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_102),
.B(n_103),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_99),
.Y(n_103)
);

BUFx24_ASAP7_75t_L g104 ( 
.A(n_81),
.Y(n_104)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_104),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_L g128 ( 
.A1(n_107),
.A2(n_77),
.B(n_90),
.Y(n_128)
);

AOI21xp5_ASAP7_75t_L g139 ( 
.A1(n_108),
.A2(n_94),
.B(n_3),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_87),
.A2(n_52),
.B1(n_72),
.B2(n_59),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_109),
.A2(n_64),
.B1(n_60),
.B2(n_5),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_79),
.B(n_51),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_111),
.B(n_83),
.Y(n_124)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_86),
.Y(n_115)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_115),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_76),
.B(n_64),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_116),
.B(n_118),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_80),
.B(n_61),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_80),
.B(n_82),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_119),
.B(n_120),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_95),
.B(n_61),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_112),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_122),
.B(n_124),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_108),
.B(n_76),
.C(n_88),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_126),
.B(n_105),
.C(n_121),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_104),
.Y(n_127)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_127),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_L g156 ( 
.A1(n_128),
.A2(n_103),
.B(n_104),
.Y(n_156)
);

NAND2x1_ASAP7_75t_L g129 ( 
.A(n_100),
.B(n_90),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_SL g148 ( 
.A1(n_129),
.A2(n_132),
.B(n_139),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_117),
.A2(n_78),
.B1(n_92),
.B2(n_84),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_131),
.A2(n_136),
.B1(n_140),
.B2(n_141),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_118),
.B(n_98),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_133),
.B(n_137),
.Y(n_160)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_112),
.Y(n_134)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_134),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_117),
.A2(n_63),
.B1(n_93),
.B2(n_97),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_106),
.B(n_98),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_115),
.A2(n_100),
.B1(n_102),
.B2(n_114),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_114),
.A2(n_89),
.B1(n_91),
.B2(n_64),
.Y(n_141)
);

AND2x2_ASAP7_75t_L g161 ( 
.A(n_142),
.B(n_60),
.Y(n_161)
);

BUFx24_ASAP7_75t_SL g143 ( 
.A(n_135),
.Y(n_143)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_143),
.Y(n_172)
);

NAND3xp33_ASAP7_75t_L g145 ( 
.A(n_135),
.B(n_119),
.C(n_116),
.Y(n_145)
);

AOI322xp5_ASAP7_75t_L g166 ( 
.A1(n_145),
.A2(n_129),
.A3(n_130),
.B1(n_132),
.B2(n_123),
.C1(n_104),
.C2(n_127),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_SL g146 ( 
.A(n_125),
.B(n_110),
.Y(n_146)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_146),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g147 ( 
.A(n_126),
.B(n_101),
.Y(n_147)
);

XOR2xp5_ASAP7_75t_L g175 ( 
.A(n_147),
.B(n_156),
.Y(n_175)
);

AOI21xp5_ASAP7_75t_L g149 ( 
.A1(n_128),
.A2(n_107),
.B(n_110),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_SL g165 ( 
.A1(n_149),
.A2(n_161),
.B(n_129),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_125),
.B(n_120),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_151),
.B(n_153),
.Y(n_164)
);

INVxp67_ASAP7_75t_L g153 ( 
.A(n_138),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_134),
.Y(n_154)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_154),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_157),
.B(n_159),
.C(n_139),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_141),
.B(n_121),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_158),
.A2(n_136),
.B1(n_131),
.B2(n_123),
.Y(n_163)
);

XOR2xp5_ASAP7_75t_L g159 ( 
.A(n_140),
.B(n_105),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_162),
.B(n_165),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_163),
.B(n_155),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_SL g180 ( 
.A(n_166),
.B(n_156),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_161),
.A2(n_132),
.B1(n_130),
.B2(n_113),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_168),
.B(n_170),
.Y(n_182)
);

HB1xp67_ASAP7_75t_L g169 ( 
.A(n_157),
.Y(n_169)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_169),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_161),
.A2(n_113),
.B1(n_10),
.B2(n_11),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_147),
.B(n_9),
.C(n_14),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_171),
.B(n_160),
.C(n_150),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_155),
.A2(n_8),
.B1(n_13),
.B2(n_10),
.Y(n_173)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_173),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_176),
.B(n_177),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_180),
.B(n_185),
.Y(n_192)
);

NAND2xp33_ASAP7_75t_SL g181 ( 
.A(n_165),
.B(n_148),
.Y(n_181)
);

NAND2xp33_ASAP7_75t_SL g194 ( 
.A(n_181),
.B(n_167),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_175),
.B(n_148),
.C(n_159),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_184),
.B(n_175),
.C(n_171),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_164),
.B(n_153),
.Y(n_185)
);

AOI21xp5_ASAP7_75t_L g186 ( 
.A1(n_168),
.A2(n_152),
.B(n_149),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_186),
.B(n_173),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_186),
.A2(n_162),
.B1(n_164),
.B2(n_170),
.Y(n_187)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_187),
.Y(n_196)
);

XOR2xp5_ASAP7_75t_L g195 ( 
.A(n_188),
.B(n_193),
.Y(n_195)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_189),
.Y(n_198)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_182),
.Y(n_191)
);

OAI31xp33_ASAP7_75t_L g200 ( 
.A1(n_191),
.A2(n_144),
.A3(n_177),
.B(n_172),
.Y(n_200)
);

XOR2xp5_ASAP7_75t_L g193 ( 
.A(n_179),
.B(n_174),
.Y(n_193)
);

A2O1A1Ixp33_ASAP7_75t_SL g199 ( 
.A1(n_194),
.A2(n_181),
.B(n_167),
.C(n_179),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_188),
.A2(n_184),
.B1(n_178),
.B2(n_183),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_197),
.B(n_200),
.Y(n_202)
);

NAND3xp33_ASAP7_75t_L g204 ( 
.A(n_199),
.B(n_4),
.C(n_5),
.Y(n_204)
);

AOI322xp5_ASAP7_75t_L g201 ( 
.A1(n_198),
.A2(n_192),
.A3(n_190),
.B1(n_191),
.B2(n_187),
.C1(n_193),
.C2(n_15),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_201),
.B(n_203),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_196),
.B(n_2),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_204),
.B(n_205),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_196),
.A2(n_7),
.B1(n_9),
.B2(n_199),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_202),
.B(n_195),
.C(n_7),
.Y(n_206)
);

XOR2xp5_ASAP7_75t_L g209 ( 
.A(n_206),
.B(n_204),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_209),
.B(n_210),
.Y(n_211)
);

AOI21xp5_ASAP7_75t_L g210 ( 
.A1(n_207),
.A2(n_7),
.B(n_208),
.Y(n_210)
);


endmodule