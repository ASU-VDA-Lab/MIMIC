module fake_jpeg_14691_n_62 (n_3, n_2, n_1, n_0, n_4, n_8, n_6, n_5, n_7, n_62);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_6;
input n_5;
input n_7;

output n_62;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_23;
wire n_10;
wire n_27;
wire n_55;
wire n_22;
wire n_51;
wire n_47;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_59;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_56;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_15;

INVx2_ASAP7_75t_L g9 ( 
.A(n_4),
.Y(n_9)
);

INVx2_ASAP7_75t_L g10 ( 
.A(n_1),
.Y(n_10)
);

INVx2_ASAP7_75t_L g11 ( 
.A(n_1),
.Y(n_11)
);

BUFx6f_ASAP7_75t_L g12 ( 
.A(n_6),
.Y(n_12)
);

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_7),
.Y(n_13)
);

BUFx2_ASAP7_75t_L g14 ( 
.A(n_1),
.Y(n_14)
);

INVx11_ASAP7_75t_L g15 ( 
.A(n_7),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_9),
.B(n_0),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_SL g32 ( 
.A(n_19),
.B(n_23),
.Y(n_32)
);

AOI22xp5_ASAP7_75t_SL g20 ( 
.A1(n_9),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_20)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_17),
.B(n_0),
.C(n_2),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g29 ( 
.A(n_21),
.B(n_17),
.C(n_12),
.Y(n_29)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_22),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_10),
.B(n_3),
.Y(n_23)
);

AOI22xp5_ASAP7_75t_L g24 ( 
.A1(n_11),
.A2(n_3),
.B1(n_5),
.B2(n_6),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_SL g25 ( 
.A(n_18),
.B(n_8),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_SL g35 ( 
.A(n_25),
.B(n_15),
.Y(n_35)
);

INVxp67_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_26),
.B(n_14),
.Y(n_33)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_18),
.Y(n_27)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_27),
.Y(n_37)
);

AOI22xp33_ASAP7_75t_L g28 ( 
.A1(n_22),
.A2(n_15),
.B1(n_14),
.B2(n_13),
.Y(n_28)
);

OAI21xp5_ASAP7_75t_SL g42 ( 
.A1(n_28),
.A2(n_34),
.B(n_30),
.Y(n_42)
);

MAJIxp5_ASAP7_75t_L g40 ( 
.A(n_29),
.B(n_36),
.C(n_38),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_L g31 ( 
.A1(n_24),
.A2(n_8),
.B1(n_12),
.B2(n_13),
.Y(n_31)
);

XNOR2xp5_ASAP7_75t_L g41 ( 
.A(n_31),
.B(n_38),
.Y(n_41)
);

CKINVDCx14_ASAP7_75t_R g45 ( 
.A(n_33),
.Y(n_45)
);

AND2x4_ASAP7_75t_L g34 ( 
.A(n_20),
.B(n_17),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_SL g43 ( 
.A(n_35),
.B(n_32),
.Y(n_43)
);

MAJIxp5_ASAP7_75t_L g36 ( 
.A(n_21),
.B(n_16),
.C(n_27),
.Y(n_36)
);

XNOR2xp5_ASAP7_75t_L g38 ( 
.A(n_23),
.B(n_21),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_37),
.Y(n_39)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_39),
.Y(n_47)
);

XNOR2xp5_ASAP7_75t_L g46 ( 
.A(n_40),
.B(n_29),
.Y(n_46)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_43),
.Y(n_49)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_36),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_46),
.B(n_48),
.Y(n_52)
);

XNOR2xp5_ASAP7_75t_L g48 ( 
.A(n_40),
.B(n_34),
.Y(n_48)
);

MAJIxp5_ASAP7_75t_L g50 ( 
.A(n_44),
.B(n_34),
.C(n_41),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_50),
.B(n_51),
.Y(n_55)
);

XOR2xp5_ASAP7_75t_L g51 ( 
.A(n_41),
.B(n_42),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_51),
.B(n_50),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_53),
.B(n_55),
.Y(n_58)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_47),
.Y(n_54)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_49),
.Y(n_56)
);

NOR2x1_ASAP7_75t_L g57 ( 
.A(n_56),
.B(n_45),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_57),
.B(n_54),
.Y(n_59)
);

OAI21xp5_ASAP7_75t_L g61 ( 
.A1(n_59),
.A2(n_60),
.B(n_57),
.Y(n_61)
);

XNOR2xp5_ASAP7_75t_L g60 ( 
.A(n_58),
.B(n_52),
.Y(n_60)
);

MAJIxp5_ASAP7_75t_L g62 ( 
.A(n_61),
.B(n_60),
.C(n_58),
.Y(n_62)
);


endmodule