module real_jpeg_16990_n_11 (n_5, n_4, n_8, n_0, n_1, n_2, n_6, n_7, n_3, n_10, n_9, n_11);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_11;

wire n_17;
wire n_21;
wire n_33;
wire n_29;
wire n_31;
wire n_12;
wire n_24;
wire n_34;
wire n_28;
wire n_23;
wire n_14;
wire n_25;
wire n_22;
wire n_18;
wire n_26;
wire n_27;
wire n_20;
wire n_19;
wire n_32;
wire n_30;
wire n_16;
wire n_15;
wire n_13;

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_0),
.Y(n_14)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_1),
.B(n_6),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_1),
.B(n_6),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_2),
.B(n_14),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_2),
.B(n_14),
.Y(n_16)
);

CKINVDCx16_ASAP7_75t_R g22 ( 
.A(n_3),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_3),
.B(n_7),
.Y(n_30)
);

MAJIxp5_ASAP7_75t_L g18 ( 
.A(n_4),
.B(n_19),
.C(n_25),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_4),
.B(n_5),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_4),
.B(n_5),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_5),
.Y(n_25)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_6),
.B(n_21),
.C(n_23),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_SL g21 ( 
.A(n_7),
.B(n_22),
.Y(n_21)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

MAJIxp5_ASAP7_75t_L g27 ( 
.A(n_8),
.B(n_9),
.C(n_28),
.Y(n_27)
);

MAJIxp5_ASAP7_75t_L g19 ( 
.A(n_9),
.B(n_20),
.C(n_24),
.Y(n_19)
);

OAI22xp5_ASAP7_75t_SL g17 ( 
.A1(n_10),
.A2(n_18),
.B1(n_26),
.B2(n_34),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_10),
.Y(n_34)
);

XOR2xp5_ASAP7_75t_L g11 ( 
.A(n_12),
.B(n_17),
.Y(n_11)
);

NAND2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_15),
.Y(n_12)
);

INVxp67_ASAP7_75t_L g15 ( 
.A(n_16),
.Y(n_15)
);

AOI21xp5_ASAP7_75t_L g26 ( 
.A1(n_27),
.A2(n_32),
.B(n_33),
.Y(n_26)
);

AOI21xp5_ASAP7_75t_L g28 ( 
.A1(n_29),
.A2(n_30),
.B(n_31),
.Y(n_28)
);


endmodule