module real_jpeg_16955_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_195;
wire n_110;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_18;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

AND2x2_ASAP7_75t_L g36 ( 
.A(n_0),
.B(n_37),
.Y(n_36)
);

AND2x2_ASAP7_75t_L g58 ( 
.A(n_0),
.B(n_59),
.Y(n_58)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_0),
.B(n_85),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_0),
.B(n_107),
.Y(n_106)
);

AND2x2_ASAP7_75t_L g165 ( 
.A(n_0),
.B(n_166),
.Y(n_165)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_1),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g89 ( 
.A(n_1),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g167 ( 
.A(n_1),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_2),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_2),
.Y(n_60)
);

BUFx5_ASAP7_75t_L g95 ( 
.A(n_2),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g247 ( 
.A(n_2),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_3),
.B(n_42),
.Y(n_41)
);

AND2x2_ASAP7_75t_SL g63 ( 
.A(n_3),
.B(n_64),
.Y(n_63)
);

AND2x2_ASAP7_75t_SL g90 ( 
.A(n_3),
.B(n_91),
.Y(n_90)
);

AND2x2_ASAP7_75t_L g163 ( 
.A(n_3),
.B(n_164),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_3),
.B(n_245),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_SL g249 ( 
.A(n_3),
.B(n_250),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_3),
.B(n_82),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_4),
.B(n_27),
.Y(n_26)
);

AND2x2_ASAP7_75t_SL g88 ( 
.A(n_4),
.B(n_89),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_4),
.A2(n_9),
.B1(n_113),
.B2(n_116),
.Y(n_112)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_4),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_4),
.B(n_264),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_4),
.B(n_275),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_SL g305 ( 
.A(n_4),
.B(n_306),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_5),
.B(n_55),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_5),
.B(n_148),
.Y(n_147)
);

AND2x2_ASAP7_75t_L g223 ( 
.A(n_5),
.B(n_224),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_5),
.B(n_259),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_5),
.B(n_268),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_SL g314 ( 
.A(n_5),
.B(n_315),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_SL g319 ( 
.A(n_5),
.B(n_320),
.Y(n_319)
);

AND2x2_ASAP7_75t_L g29 ( 
.A(n_6),
.B(n_30),
.Y(n_29)
);

AND2x2_ASAP7_75t_L g51 ( 
.A(n_6),
.B(n_52),
.Y(n_51)
);

AND2x2_ASAP7_75t_L g94 ( 
.A(n_6),
.B(n_95),
.Y(n_94)
);

AND2x2_ASAP7_75t_L g140 ( 
.A(n_6),
.B(n_141),
.Y(n_140)
);

AND2x2_ASAP7_75t_L g174 ( 
.A(n_6),
.B(n_115),
.Y(n_174)
);

NAND2x1p5_ASAP7_75t_L g186 ( 
.A(n_6),
.B(n_187),
.Y(n_186)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_7),
.Y(n_83)
);

BUFx5_ASAP7_75t_L g107 ( 
.A(n_7),
.Y(n_107)
);

BUFx5_ASAP7_75t_L g115 ( 
.A(n_7),
.Y(n_115)
);

BUFx3_ASAP7_75t_L g137 ( 
.A(n_7),
.Y(n_137)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_8),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_8),
.Y(n_53)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_8),
.Y(n_93)
);

BUFx3_ASAP7_75t_L g161 ( 
.A(n_8),
.Y(n_161)
);

BUFx3_ASAP7_75t_L g222 ( 
.A(n_8),
.Y(n_222)
);

AND2x2_ASAP7_75t_L g102 ( 
.A(n_9),
.B(n_103),
.Y(n_102)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_9),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_9),
.B(n_95),
.Y(n_190)
);

INVx6_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_10),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_11),
.B(n_46),
.Y(n_45)
);

AND2x2_ASAP7_75t_L g69 ( 
.A(n_11),
.B(n_70),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_11),
.B(n_81),
.Y(n_80)
);

AND2x2_ASAP7_75t_L g158 ( 
.A(n_11),
.B(n_159),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_12),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g188 ( 
.A(n_12),
.Y(n_188)
);

AND2x2_ASAP7_75t_L g73 ( 
.A(n_13),
.B(n_74),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_13),
.B(n_99),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_13),
.B(n_145),
.Y(n_144)
);

AND2x2_ASAP7_75t_L g216 ( 
.A(n_13),
.B(n_217),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_13),
.B(n_267),
.Y(n_266)
);

AND2x2_ASAP7_75t_L g293 ( 
.A(n_13),
.B(n_59),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_13),
.B(n_302),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_SL g324 ( 
.A(n_13),
.B(n_306),
.Y(n_324)
);

BUFx12f_ASAP7_75t_L g72 ( 
.A(n_14),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_14),
.Y(n_105)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_15),
.Y(n_57)
);

BUFx8_ASAP7_75t_L g99 ( 
.A(n_15),
.Y(n_99)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_199),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_198),
.Y(n_17)
);

INVxp67_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

AND2x2_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_150),
.Y(n_19)
);

OR2x2_ASAP7_75t_L g198 ( 
.A(n_20),
.B(n_150),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_96),
.C(n_121),
.Y(n_20)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_21),
.B(n_228),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_61),
.Y(n_21)
);

XNOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_39),
.Y(n_22)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_23),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g23 ( 
.A1(n_24),
.A2(n_25),
.B1(n_35),
.B2(n_36),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

AOI22xp33_ASAP7_75t_SL g25 ( 
.A1(n_26),
.A2(n_29),
.B1(n_33),
.B2(n_34),
.Y(n_25)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_26),
.Y(n_33)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_26),
.B(n_34),
.C(n_35),
.Y(n_176)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_28),
.Y(n_164)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_29),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g262 ( 
.A(n_32),
.Y(n_262)
);

INVx1_ASAP7_75t_SL g35 ( 
.A(n_36),
.Y(n_35)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_39),
.Y(n_153)
);

XOR2xp5_ASAP7_75t_L g39 ( 
.A(n_40),
.B(n_50),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_L g40 ( 
.A1(n_41),
.A2(n_44),
.B1(n_45),
.B2(n_49),
.Y(n_40)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_41),
.Y(n_49)
);

A2O1A1Ixp33_ASAP7_75t_L g194 ( 
.A1(n_41),
.A2(n_45),
.B(n_50),
.C(n_195),
.Y(n_194)
);

BUFx5_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_43),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_43),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g226 ( 
.A(n_43),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_44),
.B(n_49),
.Y(n_195)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

MAJIxp5_ASAP7_75t_L g50 ( 
.A(n_51),
.B(n_54),
.C(n_58),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_51),
.A2(n_58),
.B1(n_124),
.B2(n_125),
.Y(n_123)
);

INVx1_ASAP7_75t_SL g124 ( 
.A(n_51),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

XOR2xp5_ASAP7_75t_L g122 ( 
.A(n_54),
.B(n_123),
.Y(n_122)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_58),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_61),
.B(n_152),
.C(n_153),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g61 ( 
.A(n_62),
.B(n_77),
.C(n_87),
.Y(n_61)
);

XNOR2xp5_ASAP7_75t_SL g206 ( 
.A(n_62),
.B(n_207),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g62 ( 
.A(n_63),
.B(n_68),
.Y(n_62)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_63),
.B(n_69),
.C(n_73),
.Y(n_110)
);

HB1xp67_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

XNOR2xp5_ASAP7_75t_L g68 ( 
.A(n_69),
.B(n_73),
.Y(n_68)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx3_ASAP7_75t_L g304 ( 
.A(n_71),
.Y(n_304)
);

INVx5_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx2_ASAP7_75t_SL g86 ( 
.A(n_72),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g250 ( 
.A(n_72),
.Y(n_250)
);

INVx3_ASAP7_75t_L g276 ( 
.A(n_72),
.Y(n_276)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx4_ASAP7_75t_L g149 ( 
.A(n_76),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_77),
.A2(n_78),
.B1(n_87),
.B2(n_208),
.Y(n_207)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_79),
.B(n_84),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_79),
.A2(n_80),
.B1(n_84),
.B2(n_173),
.Y(n_214)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

BUFx3_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx2_ASAP7_75t_L g308 ( 
.A(n_83),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_84),
.A2(n_173),
.B1(n_174),
.B2(n_175),
.Y(n_172)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_84),
.Y(n_173)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_87),
.Y(n_208)
);

MAJx2_ASAP7_75t_L g87 ( 
.A(n_88),
.B(n_90),
.C(n_94),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_88),
.A2(n_94),
.B1(n_212),
.B2(n_213),
.Y(n_211)
);

CKINVDCx14_ASAP7_75t_R g212 ( 
.A(n_88),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_L g210 ( 
.A(n_90),
.B(n_211),
.Y(n_210)
);

BUFx3_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

BUFx3_ASAP7_75t_L g269 ( 
.A(n_93),
.Y(n_269)
);

INVx1_ASAP7_75t_SL g213 ( 
.A(n_94),
.Y(n_213)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_95),
.Y(n_265)
);

INVx2_ASAP7_75t_SL g316 ( 
.A(n_95),
.Y(n_316)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_96),
.B(n_121),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_109),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_97),
.B(n_111),
.C(n_120),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g97 ( 
.A(n_98),
.B(n_100),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_98),
.B(n_102),
.C(n_106),
.Y(n_192)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_99),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_101),
.A2(n_102),
.B1(n_106),
.B2(n_108),
.Y(n_100)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx2_ASAP7_75t_L g323 ( 
.A(n_104),
.Y(n_323)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_105),
.Y(n_142)
);

INVx1_ASAP7_75t_SL g108 ( 
.A(n_106),
.Y(n_108)
);

AND2x2_ASAP7_75t_L g139 ( 
.A(n_106),
.B(n_140),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_108),
.B(n_140),
.Y(n_242)
);

AOI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_110),
.A2(n_111),
.B1(n_112),
.B2(n_120),
.Y(n_109)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_110),
.Y(n_120)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

AOI21xp5_ASAP7_75t_L g126 ( 
.A1(n_112),
.A2(n_127),
.B(n_133),
.Y(n_126)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_118),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_122),
.B(n_126),
.C(n_138),
.Y(n_121)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_122),
.B(n_126),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_128),
.B(n_129),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_SL g170 ( 
.A(n_128),
.B(n_171),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_128),
.B(n_221),
.Y(n_220)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

BUFx3_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_134),
.B(n_135),
.Y(n_133)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

BUFx3_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_SL g203 ( 
.A(n_138),
.B(n_204),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_143),
.C(n_146),
.Y(n_138)
);

XOR2xp5_ASAP7_75t_L g239 ( 
.A(n_139),
.B(n_240),
.Y(n_239)
);

INVx5_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_143),
.A2(n_144),
.B1(n_146),
.B2(n_147),
.Y(n_240)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

INVx4_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

XNOR2xp5_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_154),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_155),
.A2(n_156),
.B1(n_179),
.B2(n_180),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_168),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_162),
.Y(n_157)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_SL g162 ( 
.A(n_163),
.B(n_165),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g219 ( 
.A(n_167),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_169),
.A2(n_176),
.B1(n_177),
.B2(n_178),
.Y(n_168)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_169),
.Y(n_177)
);

XNOR2x1_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_172),
.Y(n_169)
);

INVx1_ASAP7_75t_SL g175 ( 
.A(n_174),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_174),
.B(n_249),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_175),
.B(n_249),
.Y(n_248)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_176),
.Y(n_178)
);

INVx1_ASAP7_75t_SL g179 ( 
.A(n_180),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_182),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_183),
.A2(n_194),
.B1(n_196),
.B2(n_197),
.Y(n_182)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_183),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_184),
.A2(n_185),
.B1(n_192),
.B2(n_193),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_186),
.A2(n_189),
.B1(n_190),
.B2(n_191),
.Y(n_185)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_186),
.Y(n_191)
);

BUFx6f_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

INVx1_ASAP7_75t_SL g189 ( 
.A(n_190),
.Y(n_189)
);

INVx1_ASAP7_75t_SL g193 ( 
.A(n_192),
.Y(n_193)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_194),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_L g199 ( 
.A1(n_200),
.A2(n_229),
.B(n_336),
.Y(n_199)
);

HB1xp67_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_202),
.B(n_227),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_202),
.B(n_227),
.Y(n_336)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_203),
.B(n_205),
.C(n_209),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g232 ( 
.A(n_203),
.B(n_233),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_205),
.A2(n_206),
.B1(n_209),
.B2(n_234),
.Y(n_233)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_209),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_210),
.B(n_214),
.C(n_215),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_L g237 ( 
.A(n_210),
.B(n_238),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_214),
.B(n_215),
.Y(n_238)
);

MAJx2_ASAP7_75t_L g215 ( 
.A(n_216),
.B(n_220),
.C(n_223),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_216),
.B(n_223),
.Y(n_283)
);

INVx3_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_220),
.B(n_283),
.Y(n_282)
);

INVx5_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

OAI21x1_ASAP7_75t_SL g230 ( 
.A1(n_231),
.A2(n_251),
.B(n_335),
.Y(n_230)
);

NOR2xp67_ASAP7_75t_SL g231 ( 
.A(n_232),
.B(n_235),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_SL g335 ( 
.A(n_232),
.B(n_235),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_236),
.B(n_239),
.C(n_241),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_SL g331 ( 
.A1(n_236),
.A2(n_237),
.B1(n_332),
.B2(n_333),
.Y(n_331)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_SL g333 ( 
.A(n_239),
.B(n_241),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_243),
.C(n_248),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_242),
.A2(n_243),
.B1(n_244),
.B2(n_286),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_242),
.Y(n_286)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

INVx4_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

INVx6_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_SL g284 ( 
.A(n_248),
.B(n_285),
.Y(n_284)
);

AOI21x1_ASAP7_75t_SL g251 ( 
.A1(n_252),
.A2(n_329),
.B(n_334),
.Y(n_251)
);

OAI21xp5_ASAP7_75t_L g252 ( 
.A1(n_253),
.A2(n_287),
.B(n_328),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_254),
.B(n_279),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_SL g328 ( 
.A(n_254),
.B(n_279),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_255),
.B(n_270),
.C(n_277),
.Y(n_254)
);

AOI22xp33_ASAP7_75t_SL g294 ( 
.A1(n_255),
.A2(n_256),
.B1(n_295),
.B2(n_297),
.Y(n_294)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_257),
.B(n_266),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_258),
.B(n_263),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_258),
.B(n_263),
.C(n_266),
.Y(n_281)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

BUFx3_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_270),
.A2(n_277),
.B1(n_278),
.B2(n_296),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_270),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_271),
.B(n_273),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_271),
.A2(n_272),
.B1(n_273),
.B2(n_274),
.Y(n_290)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

INVx4_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_280),
.B(n_284),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_281),
.B(n_282),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_281),
.B(n_282),
.C(n_284),
.Y(n_330)
);

AOI21xp5_ASAP7_75t_L g287 ( 
.A1(n_288),
.A2(n_298),
.B(n_327),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_289),
.B(n_294),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_SL g327 ( 
.A(n_289),
.B(n_294),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_290),
.B(n_291),
.C(n_293),
.Y(n_289)
);

XOR2xp5_ASAP7_75t_L g309 ( 
.A(n_290),
.B(n_310),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_SL g310 ( 
.A1(n_291),
.A2(n_292),
.B1(n_293),
.B2(n_311),
.Y(n_310)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

CKINVDCx16_ASAP7_75t_R g311 ( 
.A(n_293),
.Y(n_311)
);

INVxp67_ASAP7_75t_SL g297 ( 
.A(n_295),
.Y(n_297)
);

OAI21xp5_ASAP7_75t_SL g298 ( 
.A1(n_299),
.A2(n_312),
.B(n_326),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_300),
.B(n_309),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_SL g326 ( 
.A(n_300),
.B(n_309),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_301),
.B(n_305),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_L g317 ( 
.A(n_301),
.B(n_305),
.Y(n_317)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_303),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_304),
.Y(n_303)
);

INVx2_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_308),
.Y(n_307)
);

AOI21xp5_ASAP7_75t_L g312 ( 
.A1(n_313),
.A2(n_318),
.B(n_325),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_314),
.B(n_317),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_SL g325 ( 
.A(n_314),
.B(n_317),
.Y(n_325)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_316),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_319),
.B(n_324),
.Y(n_318)
);

INVx2_ASAP7_75t_L g320 ( 
.A(n_321),
.Y(n_320)
);

BUFx2_ASAP7_75t_L g321 ( 
.A(n_322),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_323),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_330),
.B(n_331),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_SL g334 ( 
.A(n_330),
.B(n_331),
.Y(n_334)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_333),
.Y(n_332)
);


endmodule