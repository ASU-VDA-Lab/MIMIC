module fake_jpeg_14022_n_158 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_158);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_158;

wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_51;
wire n_147;
wire n_73;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_35),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_23),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_46),
.Y(n_50)
);

BUFx5_ASAP7_75t_L g51 ( 
.A(n_19),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_47),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_17),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_34),
.B(n_18),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_7),
.Y(n_55)
);

BUFx12f_ASAP7_75t_L g56 ( 
.A(n_9),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_38),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_31),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_6),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_13),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_40),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_41),
.Y(n_62)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_43),
.Y(n_63)
);

OR2x2_ASAP7_75t_L g64 ( 
.A(n_29),
.B(n_6),
.Y(n_64)
);

BUFx10_ASAP7_75t_L g65 ( 
.A(n_12),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_45),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_9),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_36),
.Y(n_68)
);

BUFx10_ASAP7_75t_L g69 ( 
.A(n_12),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_26),
.Y(n_70)
);

CKINVDCx12_ASAP7_75t_R g71 ( 
.A(n_65),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_71),
.B(n_72),
.Y(n_82)
);

AND2x2_ASAP7_75t_L g72 ( 
.A(n_54),
.B(n_0),
.Y(n_72)
);

INVx2_ASAP7_75t_R g73 ( 
.A(n_65),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_73),
.B(n_55),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_59),
.B(n_0),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_74),
.B(n_80),
.Y(n_84)
);

HB1xp67_ASAP7_75t_L g75 ( 
.A(n_65),
.Y(n_75)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_75),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_63),
.A2(n_21),
.B1(n_42),
.B2(n_39),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_76),
.A2(n_66),
.B1(n_69),
.B2(n_57),
.Y(n_96)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_58),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_77),
.B(n_78),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_64),
.B(n_1),
.Y(n_78)
);

BUFx12f_ASAP7_75t_L g79 ( 
.A(n_51),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_79),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_60),
.B(n_1),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_83),
.B(n_95),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_79),
.Y(n_86)
);

INVx1_ASAP7_75t_SL g110 ( 
.A(n_86),
.Y(n_110)
);

AOI21xp5_ASAP7_75t_SL g88 ( 
.A1(n_73),
.A2(n_64),
.B(n_69),
.Y(n_88)
);

OAI21xp5_ASAP7_75t_L g114 ( 
.A1(n_88),
.A2(n_2),
.B(n_3),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_72),
.A2(n_69),
.B1(n_63),
.B2(n_66),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_89),
.A2(n_96),
.B1(n_61),
.B2(n_57),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_77),
.B(n_67),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_90),
.B(n_93),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_76),
.B(n_52),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_91),
.B(n_55),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_79),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_78),
.B(n_48),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_78),
.B(n_49),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_94),
.B(n_2),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_SL g95 ( 
.A(n_78),
.B(n_62),
.Y(n_95)
);

AND2x2_ASAP7_75t_L g117 ( 
.A(n_97),
.B(n_113),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_98),
.B(n_114),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_96),
.A2(n_61),
.B1(n_70),
.B2(n_68),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_99),
.A2(n_109),
.B1(n_5),
.B2(n_7),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_87),
.B(n_50),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_100),
.B(n_105),
.Y(n_118)
);

INVx13_ASAP7_75t_L g102 ( 
.A(n_81),
.Y(n_102)
);

CKINVDCx16_ASAP7_75t_R g120 ( 
.A(n_102),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_84),
.B(n_53),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_SL g126 ( 
.A(n_104),
.B(n_107),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_82),
.Y(n_105)
);

AOI21xp5_ASAP7_75t_L g106 ( 
.A1(n_88),
.A2(n_55),
.B(n_56),
.Y(n_106)
);

AOI21xp5_ASAP7_75t_L g132 ( 
.A1(n_106),
.A2(n_44),
.B(n_24),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_92),
.B(n_56),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_85),
.B(n_56),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_108),
.B(n_112),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_85),
.A2(n_86),
.B1(n_51),
.B2(n_4),
.Y(n_109)
);

BUFx24_ASAP7_75t_SL g111 ( 
.A(n_95),
.Y(n_111)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_111),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_91),
.B(n_20),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_95),
.B(n_3),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_115),
.B(n_8),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_SL g116 ( 
.A(n_112),
.B(n_4),
.C(n_5),
.Y(n_116)
);

XNOR2xp5_ASAP7_75t_L g141 ( 
.A(n_116),
.B(n_125),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_119),
.A2(n_117),
.B1(n_118),
.B2(n_127),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_106),
.B(n_100),
.C(n_99),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_123),
.B(n_127),
.C(n_130),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_124),
.B(n_128),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_114),
.B(n_8),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_97),
.B(n_25),
.C(n_37),
.Y(n_127)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_110),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_103),
.B(n_10),
.Y(n_130)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_102),
.Y(n_131)
);

AND2x2_ASAP7_75t_L g139 ( 
.A(n_131),
.B(n_133),
.Y(n_139)
);

AOI21xp5_ASAP7_75t_L g137 ( 
.A1(n_132),
.A2(n_27),
.B(n_14),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_109),
.B(n_10),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_134),
.B(n_137),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_117),
.A2(n_101),
.B1(n_13),
.B2(n_11),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_L g146 ( 
.A(n_136),
.B(n_140),
.Y(n_146)
);

XOR2xp5_ASAP7_75t_L g138 ( 
.A(n_123),
.B(n_28),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_138),
.B(n_129),
.C(n_32),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_121),
.A2(n_11),
.B1(n_15),
.B2(n_16),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_122),
.A2(n_126),
.B1(n_120),
.B2(n_131),
.Y(n_143)
);

BUFx2_ASAP7_75t_L g149 ( 
.A(n_143),
.Y(n_149)
);

A2O1A1O1Ixp25_ASAP7_75t_L g144 ( 
.A1(n_142),
.A2(n_132),
.B(n_116),
.C(n_129),
.D(n_33),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_144),
.B(n_147),
.Y(n_151)
);

AOI21xp33_ASAP7_75t_L g147 ( 
.A1(n_139),
.A2(n_22),
.B(n_30),
.Y(n_147)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_148),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_145),
.Y(n_150)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_150),
.Y(n_154)
);

AOI21xp5_ASAP7_75t_L g153 ( 
.A1(n_151),
.A2(n_149),
.B(n_141),
.Y(n_153)
);

AOI31xp67_ASAP7_75t_L g155 ( 
.A1(n_153),
.A2(n_149),
.A3(n_138),
.B(n_146),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_L g156 ( 
.A1(n_155),
.A2(n_154),
.B(n_152),
.Y(n_156)
);

INVxp67_ASAP7_75t_L g157 ( 
.A(n_156),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_157),
.B(n_135),
.Y(n_158)
);


endmodule