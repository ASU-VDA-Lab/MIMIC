module fake_jpeg_2048_n_211 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_211);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_211;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_207;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_143;
wire n_202;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_91;
wire n_93;
wire n_54;
wire n_161;
wire n_209;
wire n_208;
wire n_138;
wire n_101;
wire n_210;
wire n_149;
wire n_157;
wire n_87;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_0),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_49),
.Y(n_51)
);

BUFx4f_ASAP7_75t_L g52 ( 
.A(n_21),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_27),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_45),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_0),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_22),
.B(n_47),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_24),
.Y(n_57)
);

INVx1_ASAP7_75t_SL g58 ( 
.A(n_12),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_16),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_34),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_4),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_12),
.Y(n_62)
);

BUFx5_ASAP7_75t_L g63 ( 
.A(n_28),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_3),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_10),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_48),
.Y(n_66)
);

BUFx4f_ASAP7_75t_L g67 ( 
.A(n_25),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_37),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_5),
.Y(n_69)
);

BUFx24_ASAP7_75t_L g70 ( 
.A(n_32),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_20),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_26),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_2),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_62),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_74),
.Y(n_84)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_52),
.Y(n_75)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_75),
.Y(n_91)
);

BUFx3_ASAP7_75t_L g76 ( 
.A(n_70),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_76),
.Y(n_94)
);

INVx11_ASAP7_75t_L g77 ( 
.A(n_70),
.Y(n_77)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_77),
.Y(n_88)
);

BUFx12_ASAP7_75t_L g78 ( 
.A(n_70),
.Y(n_78)
);

INVx3_ASAP7_75t_SL g86 ( 
.A(n_78),
.Y(n_86)
);

INVx11_ASAP7_75t_L g79 ( 
.A(n_55),
.Y(n_79)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_79),
.Y(n_90)
);

OR2x2_ASAP7_75t_L g80 ( 
.A(n_58),
.B(n_1),
.Y(n_80)
);

AND2x2_ASAP7_75t_L g82 ( 
.A(n_80),
.B(n_81),
.Y(n_82)
);

BUFx12f_ASAP7_75t_L g81 ( 
.A(n_62),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_80),
.B(n_56),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_83),
.B(n_85),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_80),
.B(n_73),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_SL g87 ( 
.A(n_76),
.B(n_56),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g102 ( 
.A(n_87),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_76),
.A2(n_58),
.B1(n_71),
.B2(n_61),
.Y(n_89)
);

XNOR2xp5_ASAP7_75t_L g104 ( 
.A(n_89),
.B(n_82),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_L g92 ( 
.A1(n_74),
.A2(n_71),
.B1(n_67),
.B2(n_52),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_92),
.A2(n_93),
.B1(n_67),
.B2(n_55),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_74),
.A2(n_52),
.B1(n_67),
.B2(n_57),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_77),
.A2(n_55),
.B1(n_69),
.B2(n_50),
.Y(n_95)
);

OAI21xp33_ASAP7_75t_SL g101 ( 
.A1(n_95),
.A2(n_78),
.B(n_79),
.Y(n_101)
);

INVx1_ASAP7_75t_SL g97 ( 
.A(n_90),
.Y(n_97)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_97),
.Y(n_134)
);

O2A1O1Ixp33_ASAP7_75t_L g98 ( 
.A1(n_88),
.A2(n_77),
.B(n_78),
.C(n_75),
.Y(n_98)
);

AOI21xp5_ASAP7_75t_L g128 ( 
.A1(n_98),
.A2(n_81),
.B(n_63),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_99),
.A2(n_101),
.B1(n_104),
.B2(n_94),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_93),
.A2(n_57),
.B1(n_81),
.B2(n_72),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_100),
.A2(n_104),
.B1(n_108),
.B2(n_94),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_82),
.A2(n_79),
.B1(n_64),
.B2(n_59),
.Y(n_103)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_103),
.Y(n_123)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_91),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_105),
.B(n_106),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_83),
.B(n_82),
.C(n_91),
.Y(n_106)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_90),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_107),
.B(n_109),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_89),
.A2(n_81),
.B1(n_51),
.B2(n_53),
.Y(n_108)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_86),
.Y(n_109)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_84),
.Y(n_110)
);

INVx4_ASAP7_75t_L g132 ( 
.A(n_110),
.Y(n_132)
);

INVxp33_ASAP7_75t_SL g111 ( 
.A(n_88),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_111),
.B(n_97),
.Y(n_116)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_86),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_112),
.B(n_113),
.Y(n_129)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_84),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_98),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_114),
.B(n_115),
.Y(n_138)
);

NOR3xp33_ASAP7_75t_SL g115 ( 
.A(n_102),
.B(n_78),
.C(n_65),
.Y(n_115)
);

CKINVDCx16_ASAP7_75t_R g136 ( 
.A(n_116),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_111),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_118),
.B(n_120),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_119),
.A2(n_133),
.B1(n_5),
.B2(n_6),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_106),
.B(n_54),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_SL g121 ( 
.A(n_96),
.B(n_60),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_121),
.B(n_124),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_110),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_102),
.B(n_66),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_125),
.B(n_126),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_106),
.B(n_68),
.Y(n_126)
);

AND2x2_ASAP7_75t_L g140 ( 
.A(n_127),
.B(n_131),
.Y(n_140)
);

CKINVDCx16_ASAP7_75t_R g150 ( 
.A(n_128),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_96),
.B(n_1),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_130),
.B(n_9),
.Y(n_155)
);

NAND3xp33_ASAP7_75t_SL g131 ( 
.A(n_96),
.B(n_81),
.C(n_63),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_104),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_133)
);

A2O1A1O1Ixp25_ASAP7_75t_L g135 ( 
.A1(n_117),
.A2(n_38),
.B(n_44),
.C(n_43),
.D(n_42),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_135),
.B(n_141),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_119),
.A2(n_46),
.B1(n_41),
.B2(n_40),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_137),
.A2(n_11),
.B1(n_13),
.B2(n_14),
.Y(n_170)
);

INVxp67_ASAP7_75t_L g141 ( 
.A(n_129),
.Y(n_141)
);

INVxp67_ASAP7_75t_L g142 ( 
.A(n_122),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_142),
.B(n_144),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_143),
.B(n_152),
.Y(n_166)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_132),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_132),
.Y(n_145)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_145),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_120),
.B(n_39),
.C(n_36),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_146),
.B(n_147),
.C(n_128),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_L g147 ( 
.A(n_126),
.B(n_35),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_114),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_148),
.A2(n_124),
.B1(n_134),
.B2(n_115),
.Y(n_168)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_134),
.Y(n_149)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_149),
.Y(n_172)
);

AOI21xp5_ASAP7_75t_SL g152 ( 
.A1(n_123),
.A2(n_7),
.B(n_8),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_125),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_153),
.B(n_156),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_155),
.B(n_23),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_133),
.B(n_9),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_123),
.B(n_10),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_157),
.B(n_13),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_151),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_159),
.B(n_161),
.Y(n_178)
);

CKINVDCx16_ASAP7_75t_R g161 ( 
.A(n_139),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_162),
.B(n_164),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g163 ( 
.A(n_154),
.B(n_116),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_163),
.B(n_169),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_168),
.A2(n_138),
.B1(n_140),
.B2(n_150),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_141),
.Y(n_169)
);

AND2x2_ASAP7_75t_L g181 ( 
.A(n_170),
.B(n_171),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_142),
.B(n_11),
.Y(n_171)
);

BUFx6f_ASAP7_75t_L g173 ( 
.A(n_140),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_173),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_L g174 ( 
.A(n_147),
.B(n_33),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_L g177 ( 
.A1(n_174),
.A2(n_135),
.B(n_152),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_SL g182 ( 
.A1(n_175),
.A2(n_176),
.B(n_137),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_136),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_SL g188 ( 
.A(n_177),
.B(n_164),
.Y(n_188)
);

CKINVDCx14_ASAP7_75t_R g193 ( 
.A(n_179),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_182),
.B(n_168),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_173),
.A2(n_146),
.B1(n_15),
.B2(n_16),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_183),
.B(n_184),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_166),
.A2(n_14),
.B1(n_15),
.B2(n_17),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_L g187 ( 
.A1(n_167),
.A2(n_17),
.B(n_18),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_L g194 ( 
.A1(n_187),
.A2(n_166),
.B(n_160),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_188),
.B(n_192),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_189),
.A2(n_191),
.B1(n_194),
.B2(n_187),
.Y(n_197)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_178),
.Y(n_190)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_190),
.Y(n_198)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_185),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_180),
.B(n_163),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_194),
.B(n_186),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_196),
.B(n_197),
.Y(n_201)
);

AO21x1_ASAP7_75t_L g200 ( 
.A1(n_193),
.A2(n_181),
.B(n_177),
.Y(n_200)
);

AOI21xp5_ASAP7_75t_L g202 ( 
.A1(n_200),
.A2(n_181),
.B(n_184),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_202),
.B(n_203),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_L g203 ( 
.A1(n_198),
.A2(n_195),
.B1(n_165),
.B2(n_172),
.Y(n_203)
);

NOR2xp67_ASAP7_75t_SL g204 ( 
.A(n_201),
.B(n_196),
.Y(n_204)
);

AOI31xp33_ASAP7_75t_L g206 ( 
.A1(n_204),
.A2(n_200),
.A3(n_199),
.B(n_195),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_206),
.B(n_205),
.Y(n_207)
);

O2A1O1Ixp33_ASAP7_75t_SL g208 ( 
.A1(n_207),
.A2(n_158),
.B(n_30),
.C(n_31),
.Y(n_208)
);

NOR3xp33_ASAP7_75t_L g209 ( 
.A(n_208),
.B(n_29),
.C(n_19),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_L g210 ( 
.A1(n_209),
.A2(n_174),
.B1(n_170),
.B2(n_183),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_210),
.B(n_18),
.Y(n_211)
);


endmodule