module fake_netlist_5_1918_n_12 (n_4, n_0, n_2, n_3, n_1, n_12);

input n_4;
input n_0;
input n_2;
input n_3;
input n_1;

output n_12;

wire n_8;
wire n_10;
wire n_5;
wire n_9;
wire n_6;
wire n_11;
wire n_7;

INVx2_ASAP7_75t_L g5 ( 
.A(n_4),
.Y(n_5)
);

INVx2_ASAP7_75t_L g6 ( 
.A(n_2),
.Y(n_6)
);

OAI21x1_ASAP7_75t_L g7 ( 
.A1(n_5),
.A2(n_1),
.B(n_3),
.Y(n_7)
);

INVx2_ASAP7_75t_L g8 ( 
.A(n_7),
.Y(n_8)
);

NAND2xp5_ASAP7_75t_L g9 ( 
.A(n_8),
.B(n_6),
.Y(n_9)
);

BUFx6f_ASAP7_75t_L g10 ( 
.A(n_9),
.Y(n_10)
);

INVx1_ASAP7_75t_L g11 ( 
.A(n_10),
.Y(n_11)
);

NAND2xp33_ASAP7_75t_R g12 ( 
.A(n_11),
.B(n_0),
.Y(n_12)
);


endmodule