module fake_jpeg_32103_n_503 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_503);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_503;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_490;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx2_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

INVx4_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

INVx8_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

BUFx10_ASAP7_75t_L g22 ( 
.A(n_16),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

INVx6_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_16),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_2),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

INVx6_ASAP7_75t_SL g30 ( 
.A(n_14),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_4),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_12),
.Y(n_33)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_5),
.Y(n_34)
);

BUFx12_ASAP7_75t_L g35 ( 
.A(n_4),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_5),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_12),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_3),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_1),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_8),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_8),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_3),
.Y(n_42)
);

CKINVDCx16_ASAP7_75t_R g43 ( 
.A(n_7),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_9),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_6),
.Y(n_45)
);

CKINVDCx16_ASAP7_75t_R g46 ( 
.A(n_1),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_4),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_2),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_16),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_0),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_15),
.Y(n_51)
);

BUFx5_ASAP7_75t_L g52 ( 
.A(n_28),
.Y(n_52)
);

INVx5_ASAP7_75t_L g111 ( 
.A(n_52),
.Y(n_111)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_19),
.Y(n_53)
);

INVx5_ASAP7_75t_L g128 ( 
.A(n_53),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_25),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_54),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_25),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_55),
.Y(n_110)
);

INVx2_ASAP7_75t_SL g56 ( 
.A(n_40),
.Y(n_56)
);

INVx1_ASAP7_75t_SL g113 ( 
.A(n_56),
.Y(n_113)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_19),
.Y(n_57)
);

INVx5_ASAP7_75t_L g147 ( 
.A(n_57),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g58 ( 
.A(n_23),
.B(n_9),
.C(n_15),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_58),
.B(n_67),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_25),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_59),
.Y(n_127)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_23),
.Y(n_60)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_60),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_25),
.Y(n_61)
);

INVx6_ASAP7_75t_L g118 ( 
.A(n_61),
.Y(n_118)
);

BUFx5_ASAP7_75t_L g62 ( 
.A(n_28),
.Y(n_62)
);

INVx5_ASAP7_75t_L g152 ( 
.A(n_62),
.Y(n_152)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_17),
.Y(n_63)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_63),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_33),
.B(n_37),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_64),
.B(n_93),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_45),
.Y(n_65)
);

INVx6_ASAP7_75t_L g131 ( 
.A(n_65),
.Y(n_131)
);

BUFx5_ASAP7_75t_L g66 ( 
.A(n_28),
.Y(n_66)
);

BUFx3_ASAP7_75t_L g148 ( 
.A(n_66),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_43),
.B(n_7),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_45),
.Y(n_68)
);

INVx6_ASAP7_75t_L g156 ( 
.A(n_68),
.Y(n_156)
);

INVx8_ASAP7_75t_L g69 ( 
.A(n_19),
.Y(n_69)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_69),
.Y(n_103)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_17),
.Y(n_70)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_70),
.Y(n_116)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_32),
.Y(n_71)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_71),
.Y(n_126)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_18),
.Y(n_72)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_72),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_45),
.Y(n_73)
);

INVx3_ASAP7_75t_L g133 ( 
.A(n_73),
.Y(n_133)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_40),
.Y(n_74)
);

INVx3_ASAP7_75t_L g153 ( 
.A(n_74),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_45),
.Y(n_75)
);

INVx4_ASAP7_75t_L g117 ( 
.A(n_75),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_43),
.B(n_7),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_76),
.B(n_81),
.Y(n_114)
);

BUFx3_ASAP7_75t_L g77 ( 
.A(n_40),
.Y(n_77)
);

INVx4_ASAP7_75t_L g139 ( 
.A(n_77),
.Y(n_139)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_32),
.Y(n_78)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_78),
.Y(n_129)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_44),
.Y(n_79)
);

INVx4_ASAP7_75t_L g143 ( 
.A(n_79),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_51),
.Y(n_80)
);

INVx4_ASAP7_75t_L g145 ( 
.A(n_80),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_22),
.Y(n_81)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_44),
.Y(n_82)
);

INVx4_ASAP7_75t_L g149 ( 
.A(n_82),
.Y(n_149)
);

INVx11_ASAP7_75t_L g83 ( 
.A(n_39),
.Y(n_83)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_83),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_51),
.Y(n_84)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_84),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_51),
.Y(n_85)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_85),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_24),
.Y(n_86)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_86),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_33),
.B(n_10),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_87),
.B(n_90),
.Y(n_124)
);

INVx8_ASAP7_75t_L g88 ( 
.A(n_18),
.Y(n_88)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_88),
.Y(n_142)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_18),
.Y(n_89)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_89),
.Y(n_150)
);

BUFx12f_ASAP7_75t_L g90 ( 
.A(n_39),
.Y(n_90)
);

INVx2_ASAP7_75t_SL g91 ( 
.A(n_44),
.Y(n_91)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_91),
.Y(n_121)
);

BUFx5_ASAP7_75t_L g92 ( 
.A(n_28),
.Y(n_92)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_92),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_37),
.B(n_10),
.Y(n_93)
);

INVx6_ASAP7_75t_L g94 ( 
.A(n_39),
.Y(n_94)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_94),
.Y(n_155)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_28),
.Y(n_95)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_95),
.Y(n_132)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_26),
.Y(n_96)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_96),
.Y(n_140)
);

BUFx12f_ASAP7_75t_L g97 ( 
.A(n_39),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_97),
.B(n_98),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_27),
.B(n_38),
.Y(n_98)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_36),
.Y(n_99)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_99),
.Y(n_146)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_36),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_100),
.B(n_22),
.Y(n_134)
);

OAI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_86),
.A2(n_24),
.B1(n_34),
.B2(n_48),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_101),
.A2(n_108),
.B1(n_137),
.B2(n_22),
.Y(n_195)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_77),
.A2(n_30),
.B1(n_24),
.B2(n_21),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g165 ( 
.A1(n_102),
.A2(n_144),
.B1(n_154),
.B2(n_53),
.Y(n_165)
);

AOI22xp33_ASAP7_75t_L g104 ( 
.A1(n_80),
.A2(n_34),
.B1(n_48),
.B2(n_47),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_104),
.A2(n_106),
.B1(n_120),
.B2(n_46),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_84),
.A2(n_34),
.B1(n_49),
.B2(n_26),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_85),
.A2(n_48),
.B1(n_47),
.B2(n_27),
.Y(n_108)
);

OA22x2_ASAP7_75t_L g119 ( 
.A1(n_100),
.A2(n_49),
.B1(n_41),
.B2(n_29),
.Y(n_119)
);

OA22x2_ASAP7_75t_L g161 ( 
.A1(n_119),
.A2(n_113),
.B1(n_137),
.B2(n_125),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_94),
.A2(n_41),
.B1(n_29),
.B2(n_42),
.Y(n_120)
);

OR2x2_ASAP7_75t_SL g123 ( 
.A(n_74),
.B(n_46),
.Y(n_123)
);

CKINVDCx16_ASAP7_75t_R g171 ( 
.A(n_123),
.Y(n_171)
);

AND2x2_ASAP7_75t_L g166 ( 
.A(n_134),
.B(n_52),
.Y(n_166)
);

OAI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_54),
.A2(n_47),
.B1(n_30),
.B2(n_21),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_72),
.B(n_31),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_141),
.B(n_31),
.Y(n_164)
);

AOI22xp33_ASAP7_75t_SL g144 ( 
.A1(n_79),
.A2(n_30),
.B1(n_21),
.B2(n_47),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_SL g154 ( 
.A1(n_82),
.A2(n_50),
.B1(n_20),
.B2(n_38),
.Y(n_154)
);

BUFx4f_ASAP7_75t_SL g157 ( 
.A(n_111),
.Y(n_157)
);

BUFx3_ASAP7_75t_L g226 ( 
.A(n_157),
.Y(n_226)
);

INVx4_ASAP7_75t_L g158 ( 
.A(n_103),
.Y(n_158)
);

INVx4_ASAP7_75t_L g225 ( 
.A(n_158),
.Y(n_225)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_132),
.Y(n_159)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_159),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_114),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g221 ( 
.A(n_160),
.B(n_180),
.Y(n_221)
);

AND2x2_ASAP7_75t_L g254 ( 
.A(n_161),
.B(n_166),
.Y(n_254)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_140),
.Y(n_162)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_162),
.Y(n_237)
);

INVx3_ASAP7_75t_L g163 ( 
.A(n_142),
.Y(n_163)
);

INVx4_ASAP7_75t_L g231 ( 
.A(n_163),
.Y(n_231)
);

AO21x1_ASAP7_75t_L g241 ( 
.A1(n_164),
.A2(n_165),
.B(n_169),
.Y(n_241)
);

AOI22xp33_ASAP7_75t_L g167 ( 
.A1(n_119),
.A2(n_55),
.B1(n_59),
.B2(n_61),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_167),
.A2(n_191),
.B1(n_198),
.B2(n_208),
.Y(n_239)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_109),
.Y(n_168)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_168),
.Y(n_244)
);

AOI22xp33_ASAP7_75t_SL g169 ( 
.A1(n_145),
.A2(n_89),
.B1(n_88),
.B2(n_91),
.Y(n_169)
);

INVx6_ASAP7_75t_L g170 ( 
.A(n_107),
.Y(n_170)
);

INVx6_ASAP7_75t_L g240 ( 
.A(n_170),
.Y(n_240)
);

INVx4_ASAP7_75t_L g172 ( 
.A(n_149),
.Y(n_172)
);

INVx4_ASAP7_75t_L g238 ( 
.A(n_172),
.Y(n_238)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_146),
.Y(n_173)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_173),
.Y(n_219)
);

AND2x2_ASAP7_75t_L g174 ( 
.A(n_122),
.B(n_66),
.Y(n_174)
);

OR2x2_ASAP7_75t_L g215 ( 
.A(n_174),
.B(n_189),
.Y(n_215)
);

AOI22xp33_ASAP7_75t_SL g175 ( 
.A1(n_145),
.A2(n_56),
.B1(n_57),
.B2(n_69),
.Y(n_175)
);

INVxp67_ASAP7_75t_L g228 ( 
.A(n_175),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_124),
.B(n_95),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_SL g216 ( 
.A(n_176),
.B(n_178),
.Y(n_216)
);

BUFx3_ASAP7_75t_L g177 ( 
.A(n_148),
.Y(n_177)
);

INVx3_ASAP7_75t_L g210 ( 
.A(n_177),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_115),
.B(n_20),
.Y(n_178)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_116),
.Y(n_179)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_179),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_154),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_112),
.B(n_42),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_181),
.B(n_207),
.Y(n_211)
);

CKINVDCx16_ASAP7_75t_R g182 ( 
.A(n_119),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_182),
.B(n_206),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_183),
.A2(n_188),
.B1(n_202),
.B2(n_131),
.Y(n_217)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_126),
.Y(n_184)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_184),
.Y(n_250)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_129),
.Y(n_185)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_185),
.Y(n_253)
);

INVx5_ASAP7_75t_L g186 ( 
.A(n_152),
.Y(n_186)
);

INVx3_ASAP7_75t_L g223 ( 
.A(n_186),
.Y(n_223)
);

AOI21xp5_ASAP7_75t_L g187 ( 
.A1(n_101),
.A2(n_50),
.B(n_14),
.Y(n_187)
);

AOI21xp5_ASAP7_75t_L g220 ( 
.A1(n_187),
.A2(n_144),
.B(n_131),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_104),
.A2(n_73),
.B1(n_65),
.B2(n_68),
.Y(n_188)
);

A2O1A1Ixp33_ASAP7_75t_L g189 ( 
.A1(n_121),
.A2(n_92),
.B(n_62),
.C(n_22),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_150),
.B(n_75),
.C(n_90),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_190),
.B(n_205),
.C(n_143),
.Y(n_218)
);

AOI22xp33_ASAP7_75t_L g191 ( 
.A1(n_138),
.A2(n_83),
.B1(n_90),
.B2(n_97),
.Y(n_191)
);

BUFx6f_ASAP7_75t_L g192 ( 
.A(n_107),
.Y(n_192)
);

INVx6_ASAP7_75t_L g242 ( 
.A(n_192),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_SL g193 ( 
.A(n_113),
.B(n_11),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_SL g235 ( 
.A(n_193),
.B(n_197),
.Y(n_235)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_155),
.Y(n_194)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_194),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_L g222 ( 
.A1(n_195),
.A2(n_187),
.B1(n_198),
.B2(n_171),
.Y(n_222)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_130),
.Y(n_196)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_196),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_SL g197 ( 
.A(n_121),
.B(n_11),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_135),
.A2(n_97),
.B1(n_11),
.B2(n_12),
.Y(n_198)
);

BUFx4f_ASAP7_75t_SL g199 ( 
.A(n_128),
.Y(n_199)
);

INVxp67_ASAP7_75t_L g230 ( 
.A(n_199),
.Y(n_230)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_149),
.Y(n_200)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_200),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_153),
.B(n_35),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_SL g236 ( 
.A(n_201),
.B(n_143),
.Y(n_236)
);

OAI22xp33_ASAP7_75t_SL g202 ( 
.A1(n_136),
.A2(n_22),
.B1(n_35),
.B2(n_10),
.Y(n_202)
);

BUFx3_ASAP7_75t_L g203 ( 
.A(n_148),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_203),
.Y(n_232)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_105),
.Y(n_204)
);

HB1xp67_ASAP7_75t_L g245 ( 
.A(n_204),
.Y(n_245)
);

AND2x2_ASAP7_75t_L g205 ( 
.A(n_139),
.B(n_22),
.Y(n_205)
);

INVx3_ASAP7_75t_L g206 ( 
.A(n_139),
.Y(n_206)
);

INVx5_ASAP7_75t_L g207 ( 
.A(n_147),
.Y(n_207)
);

AO22x1_ASAP7_75t_SL g208 ( 
.A1(n_117),
.A2(n_35),
.B1(n_1),
.B2(n_2),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_117),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_209),
.B(n_156),
.Y(n_212)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_212),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_174),
.B(n_156),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_213),
.B(n_227),
.Y(n_260)
);

XOR2xp5_ASAP7_75t_L g214 ( 
.A(n_174),
.B(n_102),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_214),
.B(n_247),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_L g289 ( 
.A1(n_217),
.A2(n_13),
.B1(n_15),
.B2(n_14),
.Y(n_289)
);

INVxp67_ASAP7_75t_L g256 ( 
.A(n_218),
.Y(n_256)
);

OAI21x1_ASAP7_75t_L g278 ( 
.A1(n_220),
.A2(n_199),
.B(n_157),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_222),
.A2(n_248),
.B1(n_252),
.B2(n_10),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_166),
.B(n_118),
.Y(n_227)
);

INVxp67_ASAP7_75t_L g275 ( 
.A(n_236),
.Y(n_275)
);

AOI22xp33_ASAP7_75t_L g243 ( 
.A1(n_161),
.A2(n_133),
.B1(n_118),
.B2(n_127),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_243),
.A2(n_249),
.B1(n_192),
.B2(n_170),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_166),
.B(n_181),
.C(n_190),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_195),
.A2(n_127),
.B1(n_110),
.B2(n_151),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_183),
.A2(n_110),
.B1(n_11),
.B2(n_13),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_161),
.A2(n_35),
.B1(n_2),
.B2(n_3),
.Y(n_252)
);

BUFx8_ASAP7_75t_L g255 ( 
.A(n_226),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_255),
.Y(n_308)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_244),
.Y(n_257)
);

CKINVDCx14_ASAP7_75t_R g326 ( 
.A(n_257),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_SL g258 ( 
.A(n_211),
.B(n_173),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_SL g311 ( 
.A(n_258),
.B(n_276),
.Y(n_311)
);

INVx1_ASAP7_75t_SL g261 ( 
.A(n_226),
.Y(n_261)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_261),
.Y(n_302)
);

AOI21xp5_ASAP7_75t_L g262 ( 
.A1(n_254),
.A2(n_161),
.B(n_205),
.Y(n_262)
);

AOI21xp5_ASAP7_75t_L g297 ( 
.A1(n_262),
.A2(n_288),
.B(n_252),
.Y(n_297)
);

INVx11_ASAP7_75t_L g263 ( 
.A(n_230),
.Y(n_263)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_263),
.Y(n_306)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_219),
.Y(n_264)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_264),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_265),
.A2(n_268),
.B1(n_280),
.B2(n_286),
.Y(n_307)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_219),
.Y(n_266)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_266),
.Y(n_316)
);

HB1xp67_ASAP7_75t_L g267 ( 
.A(n_225),
.Y(n_267)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_267),
.Y(n_320)
);

OAI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_217),
.A2(n_188),
.B1(n_208),
.B2(n_184),
.Y(n_268)
);

A2O1A1Ixp33_ASAP7_75t_L g269 ( 
.A1(n_211),
.A2(n_189),
.B(n_208),
.C(n_194),
.Y(n_269)
);

OAI21xp5_ASAP7_75t_SL g317 ( 
.A1(n_269),
.A2(n_270),
.B(n_278),
.Y(n_317)
);

A2O1A1Ixp33_ASAP7_75t_L g270 ( 
.A1(n_215),
.A2(n_205),
.B(n_209),
.C(n_196),
.Y(n_270)
);

INVx3_ASAP7_75t_L g271 ( 
.A(n_242),
.Y(n_271)
);

INVx3_ASAP7_75t_L g322 ( 
.A(n_271),
.Y(n_322)
);

OAI32xp33_ASAP7_75t_L g272 ( 
.A1(n_234),
.A2(n_179),
.A3(n_168),
.B1(n_185),
.B2(n_159),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_272),
.B(n_274),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_221),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_273),
.Y(n_309)
);

INVxp33_ASAP7_75t_L g274 ( 
.A(n_212),
.Y(n_274)
);

FAx1_ASAP7_75t_SL g276 ( 
.A(n_254),
.B(n_163),
.CI(n_199),
.CON(n_276),
.SN(n_276)
);

AOI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_228),
.A2(n_158),
.B1(n_206),
.B2(n_172),
.Y(n_277)
);

INVxp67_ASAP7_75t_L g327 ( 
.A(n_277),
.Y(n_327)
);

OAI22xp33_ASAP7_75t_SL g280 ( 
.A1(n_228),
.A2(n_200),
.B1(n_204),
.B2(n_207),
.Y(n_280)
);

OAI32xp33_ASAP7_75t_L g281 ( 
.A1(n_213),
.A2(n_157),
.A3(n_186),
.B1(n_177),
.B2(n_203),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_281),
.B(n_291),
.Y(n_312)
);

BUFx4f_ASAP7_75t_SL g282 ( 
.A(n_230),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g332 ( 
.A(n_282),
.Y(n_332)
);

OAI22xp5_ASAP7_75t_SL g313 ( 
.A1(n_283),
.A2(n_285),
.B1(n_290),
.B2(n_249),
.Y(n_313)
);

INVx3_ASAP7_75t_L g284 ( 
.A(n_242),
.Y(n_284)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_284),
.Y(n_330)
);

AOI22xp33_ASAP7_75t_L g285 ( 
.A1(n_239),
.A2(n_35),
.B1(n_13),
.B2(n_14),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_SL g286 ( 
.A1(n_215),
.A2(n_0),
.B1(n_3),
.B2(n_4),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_254),
.B(n_0),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_287),
.B(n_292),
.Y(n_296)
);

OAI21xp5_ASAP7_75t_SL g288 ( 
.A1(n_220),
.A2(n_13),
.B(n_15),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_289),
.A2(n_248),
.B1(n_237),
.B2(n_240),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_239),
.A2(n_6),
.B1(n_16),
.B2(n_5),
.Y(n_290)
);

INVxp67_ASAP7_75t_L g291 ( 
.A(n_210),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_SL g292 ( 
.A(n_216),
.B(n_6),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_247),
.B(n_0),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_293),
.B(n_233),
.Y(n_304)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_233),
.Y(n_294)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_294),
.Y(n_331)
);

OR2x2_ASAP7_75t_L g295 ( 
.A(n_214),
.B(n_0),
.Y(n_295)
);

CKINVDCx16_ASAP7_75t_R g310 ( 
.A(n_295),
.Y(n_310)
);

OAI21xp5_ASAP7_75t_L g339 ( 
.A1(n_297),
.A2(n_269),
.B(n_275),
.Y(n_339)
);

XOR2xp5_ASAP7_75t_L g299 ( 
.A(n_279),
.B(n_218),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g344 ( 
.A(n_299),
.B(n_300),
.C(n_301),
.Y(n_344)
);

XOR2xp5_ASAP7_75t_L g300 ( 
.A(n_279),
.B(n_227),
.Y(n_300)
);

XOR2xp5_ASAP7_75t_L g301 ( 
.A(n_293),
.B(n_241),
.Y(n_301)
);

XOR2xp5_ASAP7_75t_L g303 ( 
.A(n_256),
.B(n_241),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g351 ( 
.A(n_303),
.B(n_319),
.C(n_321),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_SL g343 ( 
.A(n_304),
.B(n_286),
.Y(n_343)
);

HAxp5_ASAP7_75t_SL g305 ( 
.A(n_287),
.B(n_235),
.CON(n_305),
.SN(n_305)
);

AOI22xp5_ASAP7_75t_SL g353 ( 
.A1(n_305),
.A2(n_261),
.B1(n_282),
.B2(n_210),
.Y(n_353)
);

AOI22xp5_ASAP7_75t_L g345 ( 
.A1(n_313),
.A2(n_265),
.B1(n_272),
.B2(n_266),
.Y(n_345)
);

OAI22xp5_ASAP7_75t_L g360 ( 
.A1(n_314),
.A2(n_284),
.B1(n_271),
.B2(n_223),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_258),
.B(n_224),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_318),
.B(n_323),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_256),
.B(n_224),
.C(n_251),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_295),
.B(n_251),
.C(n_232),
.Y(n_321)
);

AO22x2_ASAP7_75t_L g323 ( 
.A1(n_259),
.A2(n_240),
.B1(n_225),
.B2(n_231),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_295),
.B(n_253),
.C(n_245),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g358 ( 
.A(n_324),
.B(n_329),
.C(n_246),
.Y(n_358)
);

AOI22xp5_ASAP7_75t_L g325 ( 
.A1(n_268),
.A2(n_223),
.B1(n_231),
.B2(n_244),
.Y(n_325)
);

OAI22xp5_ASAP7_75t_SL g336 ( 
.A1(n_325),
.A2(n_314),
.B1(n_307),
.B2(n_277),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_259),
.B(n_250),
.Y(n_328)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_328),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_260),
.B(n_262),
.C(n_270),
.Y(n_329)
);

OAI22xp5_ASAP7_75t_L g333 ( 
.A1(n_297),
.A2(n_283),
.B1(n_290),
.B2(n_260),
.Y(n_333)
);

AOI22xp5_ASAP7_75t_L g371 ( 
.A1(n_333),
.A2(n_336),
.B1(n_346),
.B2(n_349),
.Y(n_371)
);

CKINVDCx20_ASAP7_75t_R g335 ( 
.A(n_328),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g375 ( 
.A(n_335),
.Y(n_375)
);

AO21x2_ASAP7_75t_L g338 ( 
.A1(n_317),
.A2(n_288),
.B(n_278),
.Y(n_338)
);

OAI22xp5_ASAP7_75t_SL g367 ( 
.A1(n_338),
.A2(n_362),
.B1(n_364),
.B2(n_332),
.Y(n_367)
);

OAI21xp5_ASAP7_75t_L g388 ( 
.A1(n_339),
.A2(n_342),
.B(n_348),
.Y(n_388)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_315),
.Y(n_340)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_340),
.Y(n_370)
);

CKINVDCx20_ASAP7_75t_R g341 ( 
.A(n_309),
.Y(n_341)
);

CKINVDCx20_ASAP7_75t_R g380 ( 
.A(n_341),
.Y(n_380)
);

OAI21xp5_ASAP7_75t_L g342 ( 
.A1(n_312),
.A2(n_275),
.B(n_273),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_SL g369 ( 
.A(n_343),
.B(n_354),
.Y(n_369)
);

OAI22xp5_ASAP7_75t_L g366 ( 
.A1(n_345),
.A2(n_353),
.B1(n_363),
.B2(n_332),
.Y(n_366)
);

OAI22xp5_ASAP7_75t_L g346 ( 
.A1(n_307),
.A2(n_281),
.B1(n_264),
.B2(n_276),
.Y(n_346)
);

XOR2xp5_ASAP7_75t_L g347 ( 
.A(n_299),
.B(n_276),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_L g378 ( 
.A(n_347),
.B(n_303),
.C(n_321),
.Y(n_378)
);

AND2x2_ASAP7_75t_L g348 ( 
.A(n_298),
.B(n_294),
.Y(n_348)
);

OAI22xp5_ASAP7_75t_SL g349 ( 
.A1(n_329),
.A2(n_325),
.B1(n_327),
.B2(n_309),
.Y(n_349)
);

CKINVDCx20_ASAP7_75t_R g350 ( 
.A(n_318),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_L g373 ( 
.A(n_350),
.B(n_352),
.Y(n_373)
);

AOI21xp5_ASAP7_75t_L g352 ( 
.A1(n_317),
.A2(n_291),
.B(n_282),
.Y(n_352)
);

CKINVDCx20_ASAP7_75t_R g354 ( 
.A(n_326),
.Y(n_354)
);

CKINVDCx20_ASAP7_75t_R g355 ( 
.A(n_315),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_SL g392 ( 
.A(n_355),
.B(n_357),
.Y(n_392)
);

XNOR2xp5_ASAP7_75t_L g356 ( 
.A(n_300),
.B(n_282),
.Y(n_356)
);

XNOR2xp5_ASAP7_75t_L g374 ( 
.A(n_356),
.B(n_324),
.Y(n_374)
);

OAI21xp5_ASAP7_75t_L g357 ( 
.A1(n_311),
.A2(n_263),
.B(n_255),
.Y(n_357)
);

XNOR2xp5_ASAP7_75t_SL g368 ( 
.A(n_358),
.B(n_319),
.Y(n_368)
);

NOR2xp33_ASAP7_75t_L g359 ( 
.A(n_304),
.B(n_255),
.Y(n_359)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_359),
.Y(n_394)
);

AOI22xp5_ASAP7_75t_L g389 ( 
.A1(n_360),
.A2(n_308),
.B1(n_302),
.B2(n_330),
.Y(n_389)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_316),
.Y(n_361)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_361),
.Y(n_372)
);

AOI22xp5_ASAP7_75t_L g362 ( 
.A1(n_313),
.A2(n_257),
.B1(n_238),
.B2(n_246),
.Y(n_362)
);

NOR2xp33_ASAP7_75t_SL g363 ( 
.A(n_311),
.B(n_255),
.Y(n_363)
);

AOI22xp5_ASAP7_75t_L g364 ( 
.A1(n_327),
.A2(n_238),
.B1(n_250),
.B2(n_229),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_316),
.Y(n_365)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_365),
.Y(n_384)
);

AOI22xp5_ASAP7_75t_SL g415 ( 
.A1(n_366),
.A2(n_336),
.B1(n_333),
.B2(n_338),
.Y(n_415)
);

AOI22xp5_ASAP7_75t_L g403 ( 
.A1(n_367),
.A2(n_376),
.B1(n_381),
.B2(n_346),
.Y(n_403)
);

MAJIxp5_ASAP7_75t_L g400 ( 
.A(n_368),
.B(n_379),
.C(n_385),
.Y(n_400)
);

XOR2xp5_ASAP7_75t_L g401 ( 
.A(n_374),
.B(n_377),
.Y(n_401)
);

OAI22xp5_ASAP7_75t_SL g376 ( 
.A1(n_334),
.A2(n_345),
.B1(n_339),
.B2(n_342),
.Y(n_376)
);

XOR2xp5_ASAP7_75t_L g377 ( 
.A(n_344),
.B(n_301),
.Y(n_377)
);

XNOR2xp5_ASAP7_75t_L g399 ( 
.A(n_378),
.B(n_383),
.Y(n_399)
);

MAJIxp5_ASAP7_75t_L g379 ( 
.A(n_344),
.B(n_310),
.C(n_306),
.Y(n_379)
);

OAI22xp5_ASAP7_75t_SL g381 ( 
.A1(n_334),
.A2(n_335),
.B1(n_337),
.B2(n_350),
.Y(n_381)
);

OAI22xp5_ASAP7_75t_L g382 ( 
.A1(n_348),
.A2(n_331),
.B1(n_296),
.B2(n_310),
.Y(n_382)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_382),
.Y(n_417)
);

XNOR2xp5_ASAP7_75t_L g383 ( 
.A(n_351),
.B(n_296),
.Y(n_383)
);

XOR2xp5_ASAP7_75t_L g385 ( 
.A(n_351),
.B(n_306),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_340),
.Y(n_386)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_386),
.Y(n_395)
);

MAJIxp5_ASAP7_75t_L g387 ( 
.A(n_347),
.B(n_320),
.C(n_331),
.Y(n_387)
);

MAJIxp5_ASAP7_75t_L g404 ( 
.A(n_387),
.B(n_391),
.C(n_356),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_389),
.B(n_323),
.Y(n_396)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_361),
.Y(n_390)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_390),
.Y(n_398)
);

MAJIxp5_ASAP7_75t_L g391 ( 
.A(n_358),
.B(n_320),
.C(n_323),
.Y(n_391)
);

OAI22xp5_ASAP7_75t_L g393 ( 
.A1(n_348),
.A2(n_323),
.B1(n_308),
.B2(n_330),
.Y(n_393)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_393),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_396),
.B(n_403),
.Y(n_425)
);

HB1xp67_ASAP7_75t_L g397 ( 
.A(n_394),
.Y(n_397)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_397),
.Y(n_424)
);

MAJIxp5_ASAP7_75t_L g427 ( 
.A(n_404),
.B(n_414),
.C(n_378),
.Y(n_427)
);

CKINVDCx20_ASAP7_75t_R g405 ( 
.A(n_380),
.Y(n_405)
);

NOR2xp33_ASAP7_75t_L g426 ( 
.A(n_405),
.B(n_408),
.Y(n_426)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_370),
.Y(n_406)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_406),
.Y(n_431)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_370),
.Y(n_407)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_407),
.Y(n_435)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_372),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_372),
.Y(n_409)
);

NOR2xp33_ASAP7_75t_L g436 ( 
.A(n_409),
.B(n_411),
.Y(n_436)
);

INVx2_ASAP7_75t_L g410 ( 
.A(n_394),
.Y(n_410)
);

HB1xp67_ASAP7_75t_L g422 ( 
.A(n_410),
.Y(n_422)
);

NOR2xp33_ASAP7_75t_L g411 ( 
.A(n_380),
.B(n_363),
.Y(n_411)
);

NOR2xp33_ASAP7_75t_SL g412 ( 
.A(n_383),
.B(n_341),
.Y(n_412)
);

NOR2xp33_ASAP7_75t_L g438 ( 
.A(n_412),
.B(n_413),
.Y(n_438)
);

CKINVDCx20_ASAP7_75t_R g413 ( 
.A(n_381),
.Y(n_413)
);

MAJIxp5_ASAP7_75t_L g414 ( 
.A(n_385),
.B(n_349),
.C(n_357),
.Y(n_414)
);

XNOR2xp5_ASAP7_75t_L g437 ( 
.A(n_415),
.B(n_338),
.Y(n_437)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_384),
.Y(n_416)
);

AO21x1_ASAP7_75t_L g439 ( 
.A1(n_416),
.A2(n_406),
.B(n_395),
.Y(n_439)
);

CKINVDCx20_ASAP7_75t_R g418 ( 
.A(n_373),
.Y(n_418)
);

AOI22xp5_ASAP7_75t_L g423 ( 
.A1(n_418),
.A2(n_369),
.B1(n_376),
.B2(n_392),
.Y(n_423)
);

AOI21xp5_ASAP7_75t_SL g419 ( 
.A1(n_388),
.A2(n_352),
.B(n_338),
.Y(n_419)
);

OAI21xp5_ASAP7_75t_SL g434 ( 
.A1(n_419),
.A2(n_396),
.B(n_402),
.Y(n_434)
);

XNOR2xp5_ASAP7_75t_SL g420 ( 
.A(n_414),
.B(n_377),
.Y(n_420)
);

XOR2xp5_ASAP7_75t_L g442 ( 
.A(n_420),
.B(n_421),
.Y(n_442)
);

XOR2xp5_ASAP7_75t_L g421 ( 
.A(n_401),
.B(n_374),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_423),
.B(n_415),
.Y(n_451)
);

XNOR2xp5_ASAP7_75t_L g450 ( 
.A(n_427),
.B(n_429),
.Y(n_450)
);

MAJIxp5_ASAP7_75t_L g428 ( 
.A(n_400),
.B(n_368),
.C(n_387),
.Y(n_428)
);

MAJIxp5_ASAP7_75t_L g440 ( 
.A(n_428),
.B(n_432),
.C(n_433),
.Y(n_440)
);

XOR2xp5_ASAP7_75t_L g429 ( 
.A(n_401),
.B(n_379),
.Y(n_429)
);

AOI22xp5_ASAP7_75t_L g430 ( 
.A1(n_402),
.A2(n_367),
.B1(n_375),
.B2(n_371),
.Y(n_430)
);

INVxp67_ASAP7_75t_L g454 ( 
.A(n_430),
.Y(n_454)
);

MAJx2_ASAP7_75t_L g432 ( 
.A(n_404),
.B(n_391),
.C(n_388),
.Y(n_432)
);

MAJIxp5_ASAP7_75t_L g433 ( 
.A(n_400),
.B(n_371),
.C(n_337),
.Y(n_433)
);

XOR2x1_ASAP7_75t_L g455 ( 
.A(n_434),
.B(n_338),
.Y(n_455)
);

AOI22xp5_ASAP7_75t_L g445 ( 
.A1(n_437),
.A2(n_417),
.B1(n_375),
.B2(n_419),
.Y(n_445)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_439),
.Y(n_443)
);

NOR2xp33_ASAP7_75t_L g441 ( 
.A(n_436),
.B(n_426),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_441),
.B(n_448),
.Y(n_456)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_431),
.Y(n_444)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_444),
.Y(n_468)
);

OAI22xp5_ASAP7_75t_SL g465 ( 
.A1(n_445),
.A2(n_453),
.B1(n_454),
.B2(n_455),
.Y(n_465)
);

MAJIxp5_ASAP7_75t_L g446 ( 
.A(n_433),
.B(n_399),
.C(n_403),
.Y(n_446)
);

MAJIxp5_ASAP7_75t_L g457 ( 
.A(n_446),
.B(n_447),
.C(n_432),
.Y(n_457)
);

MAJIxp5_ASAP7_75t_L g447 ( 
.A(n_427),
.B(n_399),
.C(n_410),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_435),
.Y(n_448)
);

HB1xp67_ASAP7_75t_L g449 ( 
.A(n_434),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_449),
.B(n_451),
.Y(n_459)
);

NOR2xp33_ASAP7_75t_L g452 ( 
.A(n_438),
.B(n_354),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_L g461 ( 
.A(n_452),
.B(n_423),
.Y(n_461)
);

OR2x2_ASAP7_75t_L g453 ( 
.A(n_439),
.B(n_355),
.Y(n_453)
);

AOI21xp5_ASAP7_75t_L g458 ( 
.A1(n_453),
.A2(n_395),
.B(n_398),
.Y(n_458)
);

AOI22xp5_ASAP7_75t_SL g462 ( 
.A1(n_455),
.A2(n_437),
.B1(n_430),
.B2(n_422),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_457),
.B(n_460),
.Y(n_475)
);

OAI21xp5_ASAP7_75t_L g476 ( 
.A1(n_458),
.A2(n_386),
.B(n_384),
.Y(n_476)
);

MAJIxp5_ASAP7_75t_L g460 ( 
.A(n_447),
.B(n_428),
.C(n_429),
.Y(n_460)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_461),
.Y(n_470)
);

OR2x2_ASAP7_75t_L g471 ( 
.A(n_462),
.B(n_469),
.Y(n_471)
);

MAJIxp5_ASAP7_75t_L g463 ( 
.A(n_440),
.B(n_421),
.C(n_420),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_463),
.B(n_465),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_L g464 ( 
.A(n_443),
.B(n_424),
.Y(n_464)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_464),
.Y(n_477)
);

XNOR2xp5_ASAP7_75t_L g466 ( 
.A(n_446),
.B(n_425),
.Y(n_466)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_466),
.Y(n_478)
);

OAI22xp5_ASAP7_75t_SL g467 ( 
.A1(n_454),
.A2(n_425),
.B1(n_440),
.B2(n_389),
.Y(n_467)
);

AOI22xp5_ASAP7_75t_L g480 ( 
.A1(n_467),
.A2(n_442),
.B1(n_323),
.B2(n_322),
.Y(n_480)
);

MAJIxp5_ASAP7_75t_L g469 ( 
.A(n_450),
.B(n_409),
.C(n_408),
.Y(n_469)
);

OAI21xp5_ASAP7_75t_SL g472 ( 
.A1(n_458),
.A2(n_416),
.B(n_407),
.Y(n_472)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_472),
.Y(n_482)
);

OAI22xp5_ASAP7_75t_SL g473 ( 
.A1(n_462),
.A2(n_398),
.B1(n_353),
.B2(n_390),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g485 ( 
.A(n_473),
.B(n_479),
.Y(n_485)
);

A2O1A1Ixp33_ASAP7_75t_SL g483 ( 
.A1(n_476),
.A2(n_467),
.B(n_468),
.C(n_469),
.Y(n_483)
);

OAI22xp5_ASAP7_75t_SL g479 ( 
.A1(n_459),
.A2(n_362),
.B1(n_365),
.B2(n_364),
.Y(n_479)
);

INVxp67_ASAP7_75t_L g488 ( 
.A(n_480),
.Y(n_488)
);

OAI22xp5_ASAP7_75t_SL g481 ( 
.A1(n_465),
.A2(n_442),
.B1(n_322),
.B2(n_302),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_L g486 ( 
.A(n_481),
.B(n_466),
.Y(n_486)
);

OAI21x1_ASAP7_75t_L g491 ( 
.A1(n_483),
.A2(n_474),
.B(n_471),
.Y(n_491)
);

AND2x2_ASAP7_75t_L g484 ( 
.A(n_475),
.B(n_457),
.Y(n_484)
);

AOI21xp5_ASAP7_75t_L g493 ( 
.A1(n_484),
.A2(n_489),
.B(n_471),
.Y(n_493)
);

NOR2xp33_ASAP7_75t_L g490 ( 
.A(n_486),
.B(n_487),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_L g487 ( 
.A(n_470),
.B(n_456),
.Y(n_487)
);

OAI21xp5_ASAP7_75t_SL g489 ( 
.A1(n_474),
.A2(n_463),
.B(n_460),
.Y(n_489)
);

A2O1A1Ixp33_ASAP7_75t_L g497 ( 
.A1(n_491),
.A2(n_483),
.B(n_476),
.C(n_473),
.Y(n_497)
);

NOR2xp33_ASAP7_75t_SL g492 ( 
.A(n_482),
.B(n_477),
.Y(n_492)
);

AOI21xp5_ASAP7_75t_L g496 ( 
.A1(n_492),
.A2(n_494),
.B(n_472),
.Y(n_496)
);

OAI21xp5_ASAP7_75t_L g495 ( 
.A1(n_493),
.A2(n_488),
.B(n_480),
.Y(n_495)
);

MAJIxp5_ASAP7_75t_L g494 ( 
.A(n_485),
.B(n_478),
.C(n_481),
.Y(n_494)
);

INVxp67_ASAP7_75t_L g498 ( 
.A(n_495),
.Y(n_498)
);

INVxp67_ASAP7_75t_L g499 ( 
.A(n_496),
.Y(n_499)
);

NAND3xp33_ASAP7_75t_SL g500 ( 
.A(n_498),
.B(n_490),
.C(n_497),
.Y(n_500)
);

OAI31xp33_ASAP7_75t_L g501 ( 
.A1(n_500),
.A2(n_499),
.A3(n_479),
.B(n_229),
.Y(n_501)
);

AOI21xp5_ASAP7_75t_SL g502 ( 
.A1(n_501),
.A2(n_6),
.B(n_3),
.Y(n_502)
);

XOR2xp5_ASAP7_75t_L g503 ( 
.A(n_502),
.B(n_5),
.Y(n_503)
);


endmodule