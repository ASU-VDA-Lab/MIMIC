module fake_jpeg_11976_n_526 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_526);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_526;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_349;
wire n_21;
wire n_288;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_442;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx11_ASAP7_75t_SL g18 ( 
.A(n_13),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_17),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

INVx8_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

CKINVDCx16_ASAP7_75t_R g24 ( 
.A(n_7),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_17),
.Y(n_26)
);

INVx6_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_13),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_17),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_3),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_13),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_3),
.Y(n_36)
);

INVx2_ASAP7_75t_SL g37 ( 
.A(n_1),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_14),
.Y(n_38)
);

BUFx10_ASAP7_75t_L g39 ( 
.A(n_0),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_14),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_2),
.Y(n_41)
);

INVx13_ASAP7_75t_L g42 ( 
.A(n_6),
.Y(n_42)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_2),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_2),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_1),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_6),
.Y(n_46)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_5),
.Y(n_47)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_15),
.Y(n_48)
);

BUFx4f_ASAP7_75t_L g49 ( 
.A(n_4),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_3),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_0),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_10),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_12),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_11),
.Y(n_54)
);

BUFx5_ASAP7_75t_L g55 ( 
.A(n_16),
.Y(n_55)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_15),
.Y(n_56)
);

INVx11_ASAP7_75t_L g57 ( 
.A(n_39),
.Y(n_57)
);

INVx11_ASAP7_75t_L g190 ( 
.A(n_57),
.Y(n_190)
);

INVx4_ASAP7_75t_SL g58 ( 
.A(n_39),
.Y(n_58)
);

CKINVDCx6p67_ASAP7_75t_R g129 ( 
.A(n_58),
.Y(n_129)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_32),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g150 ( 
.A(n_59),
.Y(n_150)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_43),
.Y(n_60)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_60),
.Y(n_156)
);

BUFx12_ASAP7_75t_L g61 ( 
.A(n_39),
.Y(n_61)
);

INVx13_ASAP7_75t_L g183 ( 
.A(n_61),
.Y(n_183)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_55),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g142 ( 
.A(n_62),
.Y(n_142)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_32),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g176 ( 
.A(n_63),
.Y(n_176)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_55),
.Y(n_64)
);

INVx3_ASAP7_75t_L g144 ( 
.A(n_64),
.Y(n_144)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_55),
.Y(n_65)
);

INVx3_ASAP7_75t_L g159 ( 
.A(n_65),
.Y(n_159)
);

INVx11_ASAP7_75t_L g66 ( 
.A(n_39),
.Y(n_66)
);

BUFx5_ASAP7_75t_L g177 ( 
.A(n_66),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_43),
.B(n_1),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_67),
.B(n_90),
.Y(n_130)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_33),
.Y(n_68)
);

INVx2_ASAP7_75t_SL g185 ( 
.A(n_68),
.Y(n_185)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_28),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g196 ( 
.A(n_69),
.Y(n_196)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_33),
.Y(n_70)
);

INVx1_ASAP7_75t_SL g201 ( 
.A(n_70),
.Y(n_201)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_28),
.Y(n_71)
);

INVx6_ASAP7_75t_L g141 ( 
.A(n_71),
.Y(n_141)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_47),
.Y(n_72)
);

INVx3_ASAP7_75t_L g160 ( 
.A(n_72),
.Y(n_160)
);

INVx11_ASAP7_75t_L g73 ( 
.A(n_39),
.Y(n_73)
);

BUFx24_ASAP7_75t_L g153 ( 
.A(n_73),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_28),
.Y(n_74)
);

INVx6_ASAP7_75t_L g179 ( 
.A(n_74),
.Y(n_179)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_29),
.Y(n_75)
);

INVx6_ASAP7_75t_L g195 ( 
.A(n_75),
.Y(n_195)
);

INVx6_ASAP7_75t_L g76 ( 
.A(n_32),
.Y(n_76)
);

INVx5_ASAP7_75t_L g124 ( 
.A(n_76),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_29),
.Y(n_77)
);

BUFx3_ASAP7_75t_L g145 ( 
.A(n_77),
.Y(n_145)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_47),
.Y(n_78)
);

INVx3_ASAP7_75t_L g184 ( 
.A(n_78),
.Y(n_184)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_49),
.Y(n_79)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_79),
.Y(n_165)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_29),
.Y(n_80)
);

BUFx3_ASAP7_75t_L g147 ( 
.A(n_80),
.Y(n_147)
);

INVx2_ASAP7_75t_SL g81 ( 
.A(n_22),
.Y(n_81)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_81),
.Y(n_139)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_49),
.Y(n_82)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_82),
.Y(n_175)
);

INVx13_ASAP7_75t_L g83 ( 
.A(n_42),
.Y(n_83)
);

BUFx16f_ASAP7_75t_L g149 ( 
.A(n_83),
.Y(n_149)
);

INVx8_ASAP7_75t_L g84 ( 
.A(n_46),
.Y(n_84)
);

INVx4_ASAP7_75t_L g137 ( 
.A(n_84),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_21),
.B(n_16),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_SL g151 ( 
.A(n_85),
.B(n_111),
.Y(n_151)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_47),
.Y(n_86)
);

INVx4_ASAP7_75t_L g154 ( 
.A(n_86),
.Y(n_154)
);

BUFx3_ASAP7_75t_L g87 ( 
.A(n_22),
.Y(n_87)
);

BUFx12f_ASAP7_75t_L g131 ( 
.A(n_87),
.Y(n_131)
);

CKINVDCx6p67_ASAP7_75t_R g88 ( 
.A(n_18),
.Y(n_88)
);

BUFx12f_ASAP7_75t_L g158 ( 
.A(n_88),
.Y(n_158)
);

AOI21xp33_ASAP7_75t_SL g89 ( 
.A1(n_42),
.A2(n_16),
.B(n_15),
.Y(n_89)
);

NAND2x1_ASAP7_75t_L g126 ( 
.A(n_89),
.B(n_108),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_21),
.B(n_12),
.Y(n_90)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_33),
.Y(n_91)
);

INVx4_ASAP7_75t_L g180 ( 
.A(n_91),
.Y(n_180)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_46),
.Y(n_92)
);

BUFx12f_ASAP7_75t_L g182 ( 
.A(n_92),
.Y(n_182)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_49),
.Y(n_93)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_93),
.Y(n_194)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_35),
.Y(n_94)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_94),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_SL g95 ( 
.A(n_30),
.B(n_12),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_95),
.B(n_101),
.Y(n_125)
);

INVx6_ASAP7_75t_L g96 ( 
.A(n_46),
.Y(n_96)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_96),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_49),
.Y(n_97)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_97),
.Y(n_171)
);

BUFx12f_ASAP7_75t_L g98 ( 
.A(n_35),
.Y(n_98)
);

BUFx12_ASAP7_75t_L g140 ( 
.A(n_98),
.Y(n_140)
);

BUFx3_ASAP7_75t_L g99 ( 
.A(n_22),
.Y(n_99)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_99),
.Y(n_186)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_26),
.Y(n_100)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_100),
.Y(n_128)
);

CKINVDCx16_ASAP7_75t_R g101 ( 
.A(n_42),
.Y(n_101)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_22),
.Y(n_102)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_102),
.Y(n_157)
);

INVx11_ASAP7_75t_L g103 ( 
.A(n_24),
.Y(n_103)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_103),
.Y(n_197)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_22),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_104),
.B(n_106),
.Y(n_135)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_26),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_105),
.B(n_107),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_23),
.Y(n_106)
);

BUFx3_ASAP7_75t_L g107 ( 
.A(n_35),
.Y(n_107)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_19),
.Y(n_108)
);

INVx6_ASAP7_75t_SL g109 ( 
.A(n_48),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_109),
.B(n_110),
.Y(n_133)
);

INVx8_ASAP7_75t_L g110 ( 
.A(n_27),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_30),
.B(n_1),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_23),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_112),
.B(n_114),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_38),
.B(n_4),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_SL g170 ( 
.A(n_113),
.B(n_121),
.Y(n_170)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_23),
.Y(n_114)
);

INVx8_ASAP7_75t_L g115 ( 
.A(n_27),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_115),
.B(n_116),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_27),
.Y(n_116)
);

INVx6_ASAP7_75t_L g117 ( 
.A(n_40),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_117),
.B(n_118),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_40),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_SL g119 ( 
.A(n_38),
.B(n_4),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_119),
.B(n_120),
.Y(n_163)
);

INVx6_ASAP7_75t_L g120 ( 
.A(n_40),
.Y(n_120)
);

OR2x4_ASAP7_75t_L g121 ( 
.A(n_24),
.B(n_4),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_56),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_122),
.B(n_37),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_85),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_SL g230 ( 
.A(n_123),
.B(n_166),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_67),
.B(n_53),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_127),
.B(n_152),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_117),
.A2(n_56),
.B1(n_48),
.B2(n_52),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g235 ( 
.A1(n_134),
.A2(n_136),
.B1(n_161),
.B2(n_8),
.Y(n_235)
);

AOI22xp33_ASAP7_75t_L g136 ( 
.A1(n_80),
.A2(n_56),
.B1(n_36),
.B2(n_45),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_SL g138 ( 
.A1(n_84),
.A2(n_48),
.B1(n_37),
.B2(n_53),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_SL g216 ( 
.A1(n_138),
.A2(n_77),
.B1(n_75),
.B2(n_34),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_L g146 ( 
.A1(n_111),
.A2(n_37),
.B(n_52),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_146),
.B(n_174),
.C(n_152),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_113),
.B(n_31),
.Y(n_152)
);

OAI22xp33_ASAP7_75t_L g161 ( 
.A1(n_96),
.A2(n_37),
.B1(n_50),
.B2(n_41),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_110),
.B(n_31),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_164),
.B(n_168),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_61),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_83),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_SL g241 ( 
.A(n_167),
.B(n_173),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_115),
.B(n_25),
.Y(n_168)
);

AND2x2_ASAP7_75t_L g206 ( 
.A(n_169),
.B(n_92),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_116),
.B(n_25),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_172),
.B(n_124),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_88),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_120),
.A2(n_20),
.B1(n_50),
.B2(n_41),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_88),
.B(n_54),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g221 ( 
.A(n_178),
.B(n_187),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_81),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_181),
.B(n_188),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_98),
.B(n_54),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_122),
.B(n_51),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_97),
.B(n_51),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_189),
.B(n_191),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_SL g191 ( 
.A(n_58),
.B(n_45),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_106),
.B(n_44),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_192),
.B(n_193),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_112),
.B(n_44),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_114),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_198),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_118),
.B(n_36),
.Y(n_199)
);

INVxp67_ASAP7_75t_L g236 ( 
.A(n_199),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_69),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_202),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_71),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_203),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_SL g204 ( 
.A(n_74),
.B(n_34),
.Y(n_204)
);

CKINVDCx14_ASAP7_75t_R g223 ( 
.A(n_204),
.Y(n_223)
);

OAI21xp33_ASAP7_75t_L g282 ( 
.A1(n_206),
.A2(n_211),
.B(n_217),
.Y(n_282)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_171),
.Y(n_207)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_207),
.Y(n_276)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_171),
.Y(n_208)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_208),
.Y(n_278)
);

INVx3_ASAP7_75t_L g210 ( 
.A(n_149),
.Y(n_210)
);

BUFx2_ASAP7_75t_L g281 ( 
.A(n_210),
.Y(n_281)
);

AND2x2_ASAP7_75t_L g211 ( 
.A(n_127),
.B(n_164),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_139),
.Y(n_212)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_212),
.Y(n_280)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_139),
.Y(n_213)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_213),
.Y(n_284)
);

INVx4_ASAP7_75t_L g214 ( 
.A(n_182),
.Y(n_214)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_214),
.Y(n_302)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_165),
.Y(n_215)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_215),
.Y(n_289)
);

INVxp67_ASAP7_75t_L g274 ( 
.A(n_216),
.Y(n_274)
);

AND2x2_ASAP7_75t_L g217 ( 
.A(n_168),
.B(n_5),
.Y(n_217)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_165),
.Y(n_219)
);

INVx2_ASAP7_75t_L g308 ( 
.A(n_219),
.Y(n_308)
);

CKINVDCx16_ASAP7_75t_R g220 ( 
.A(n_153),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_SL g322 ( 
.A(n_220),
.B(n_246),
.Y(n_322)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_175),
.Y(n_222)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_222),
.Y(n_299)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_128),
.Y(n_224)
);

INVxp67_ASAP7_75t_SL g287 ( 
.A(n_224),
.Y(n_287)
);

INVx6_ASAP7_75t_L g226 ( 
.A(n_196),
.Y(n_226)
);

INVx2_ASAP7_75t_L g310 ( 
.A(n_226),
.Y(n_310)
);

INVx8_ASAP7_75t_L g227 ( 
.A(n_196),
.Y(n_227)
);

INVxp67_ASAP7_75t_L g295 ( 
.A(n_227),
.Y(n_295)
);

AND2x2_ASAP7_75t_L g228 ( 
.A(n_172),
.B(n_5),
.Y(n_228)
);

AND2x2_ASAP7_75t_L g275 ( 
.A(n_228),
.B(n_239),
.Y(n_275)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_175),
.Y(n_229)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_229),
.Y(n_301)
);

AOI22xp33_ASAP7_75t_L g232 ( 
.A1(n_143),
.A2(n_20),
.B1(n_19),
.B2(n_7),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_L g279 ( 
.A1(n_232),
.A2(n_244),
.B1(n_270),
.B2(n_272),
.Y(n_279)
);

AOI22xp33_ASAP7_75t_SL g233 ( 
.A1(n_170),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_233)
);

INVxp67_ASAP7_75t_L g304 ( 
.A(n_233),
.Y(n_304)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_132),
.Y(n_234)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_234),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_235),
.A2(n_247),
.B1(n_256),
.B2(n_259),
.Y(n_305)
);

A2O1A1Ixp33_ASAP7_75t_L g237 ( 
.A1(n_126),
.A2(n_8),
.B(n_9),
.C(n_10),
.Y(n_237)
);

AOI21xp33_ASAP7_75t_L g307 ( 
.A1(n_237),
.A2(n_255),
.B(n_262),
.Y(n_307)
);

BUFx6f_ASAP7_75t_L g238 ( 
.A(n_141),
.Y(n_238)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_238),
.Y(n_318)
);

INVx3_ASAP7_75t_L g239 ( 
.A(n_149),
.Y(n_239)
);

AND2x2_ASAP7_75t_L g240 ( 
.A(n_156),
.B(n_8),
.Y(n_240)
);

OAI21xp5_ASAP7_75t_SL g314 ( 
.A1(n_240),
.A2(n_242),
.B(n_251),
.Y(n_314)
);

AND2x2_ASAP7_75t_L g242 ( 
.A(n_156),
.B(n_9),
.Y(n_242)
);

AOI22xp33_ASAP7_75t_SL g243 ( 
.A1(n_201),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_243)
);

CKINVDCx16_ASAP7_75t_R g285 ( 
.A(n_243),
.Y(n_285)
);

AOI22xp33_ASAP7_75t_L g244 ( 
.A1(n_143),
.A2(n_10),
.B1(n_11),
.B2(n_148),
.Y(n_244)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_194),
.Y(n_246)
);

OAI22xp33_ASAP7_75t_SL g247 ( 
.A1(n_134),
.A2(n_174),
.B1(n_146),
.B2(n_126),
.Y(n_247)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_194),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_248),
.B(n_249),
.Y(n_288)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_200),
.Y(n_249)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_155),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_252),
.B(n_257),
.Y(n_277)
);

BUFx2_ASAP7_75t_L g253 ( 
.A(n_137),
.Y(n_253)
);

CKINVDCx16_ASAP7_75t_R g313 ( 
.A(n_253),
.Y(n_313)
);

NAND3xp33_ASAP7_75t_SL g254 ( 
.A(n_163),
.B(n_125),
.C(n_130),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_254),
.B(n_258),
.Y(n_293)
);

AOI22xp33_ASAP7_75t_SL g255 ( 
.A1(n_201),
.A2(n_158),
.B1(n_142),
.B2(n_151),
.Y(n_255)
);

OAI22xp33_ASAP7_75t_SL g256 ( 
.A1(n_150),
.A2(n_176),
.B1(n_161),
.B2(n_147),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_135),
.Y(n_257)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_200),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_L g259 ( 
.A1(n_162),
.A2(n_133),
.B1(n_150),
.B2(n_176),
.Y(n_259)
);

INVx4_ASAP7_75t_L g261 ( 
.A(n_182),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_261),
.B(n_263),
.Y(n_297)
);

AOI22xp33_ASAP7_75t_SL g262 ( 
.A1(n_158),
.A2(n_142),
.B1(n_144),
.B2(n_159),
.Y(n_262)
);

BUFx3_ASAP7_75t_L g263 ( 
.A(n_131),
.Y(n_263)
);

AOI32xp33_ASAP7_75t_L g264 ( 
.A1(n_197),
.A2(n_185),
.A3(n_153),
.B1(n_190),
.B2(n_186),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_264),
.B(n_267),
.Y(n_315)
);

AOI22xp33_ASAP7_75t_SL g265 ( 
.A1(n_158),
.A2(n_159),
.B1(n_144),
.B2(n_180),
.Y(n_265)
);

OAI21xp5_ASAP7_75t_L g317 ( 
.A1(n_265),
.A2(n_129),
.B(n_183),
.Y(n_317)
);

INVx3_ASAP7_75t_L g266 ( 
.A(n_149),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_266),
.Y(n_283)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_157),
.Y(n_267)
);

BUFx6f_ASAP7_75t_L g268 ( 
.A(n_141),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_268),
.B(n_226),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_269),
.B(n_271),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_L g270 ( 
.A1(n_179),
.A2(n_195),
.B1(n_124),
.B2(n_145),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_186),
.B(n_180),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_L g272 ( 
.A1(n_179),
.A2(n_195),
.B1(n_145),
.B2(n_147),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_245),
.A2(n_137),
.B1(n_185),
.B2(n_160),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g341 ( 
.A1(n_273),
.A2(n_294),
.B1(n_319),
.B2(n_242),
.Y(n_341)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_271),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_286),
.B(n_291),
.Y(n_332)
);

XNOR2xp5_ASAP7_75t_L g290 ( 
.A(n_211),
.B(n_160),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g349 ( 
.A(n_290),
.B(n_312),
.C(n_229),
.Y(n_349)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_205),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_L g294 ( 
.A1(n_245),
.A2(n_184),
.B1(n_154),
.B2(n_153),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_211),
.B(n_154),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_296),
.B(n_298),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_217),
.B(n_184),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_217),
.B(n_182),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_300),
.B(n_321),
.Y(n_329)
);

AOI22xp33_ASAP7_75t_L g303 ( 
.A1(n_257),
.A2(n_252),
.B1(n_228),
.B2(n_206),
.Y(n_303)
);

OAI21xp33_ASAP7_75t_SL g355 ( 
.A1(n_303),
.A2(n_219),
.B(n_248),
.Y(n_355)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_225),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g337 ( 
.A(n_309),
.B(n_311),
.Y(n_337)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_250),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_L g312 ( 
.A(n_209),
.B(n_251),
.Y(n_312)
);

O2A1O1Ixp33_ASAP7_75t_SL g316 ( 
.A1(n_269),
.A2(n_129),
.B(n_190),
.C(n_183),
.Y(n_316)
);

OA22x2_ASAP7_75t_L g347 ( 
.A1(n_316),
.A2(n_239),
.B1(n_210),
.B2(n_214),
.Y(n_347)
);

INVxp67_ASAP7_75t_L g330 ( 
.A(n_317),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_L g319 ( 
.A1(n_223),
.A2(n_209),
.B1(n_236),
.B2(n_231),
.Y(n_319)
);

OAI21xp5_ASAP7_75t_L g320 ( 
.A1(n_236),
.A2(n_129),
.B(n_140),
.Y(n_320)
);

OAI21xp5_ASAP7_75t_L g335 ( 
.A1(n_320),
.A2(n_129),
.B(n_266),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_228),
.B(n_131),
.Y(n_321)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_323),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_R g324 ( 
.A(n_290),
.B(n_218),
.Y(n_324)
);

OAI21xp5_ASAP7_75t_SL g367 ( 
.A1(n_324),
.A2(n_332),
.B(n_343),
.Y(n_367)
);

INVx2_ASAP7_75t_L g325 ( 
.A(n_308),
.Y(n_325)
);

INVx2_ASAP7_75t_L g364 ( 
.A(n_325),
.Y(n_364)
);

FAx1_ASAP7_75t_SL g327 ( 
.A(n_292),
.B(n_237),
.CI(n_221),
.CON(n_327),
.SN(n_327)
);

NOR2xp33_ASAP7_75t_SL g381 ( 
.A(n_327),
.B(n_331),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_SL g331 ( 
.A(n_291),
.B(n_230),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_292),
.B(n_240),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_333),
.B(n_342),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_SL g334 ( 
.A(n_277),
.B(n_241),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_SL g386 ( 
.A(n_334),
.B(n_336),
.Y(n_386)
);

INVxp67_ASAP7_75t_L g391 ( 
.A(n_335),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_SL g336 ( 
.A(n_277),
.B(n_260),
.Y(n_336)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_276),
.Y(n_338)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_338),
.Y(n_368)
);

AND2x2_ASAP7_75t_L g339 ( 
.A(n_316),
.B(n_206),
.Y(n_339)
);

CKINVDCx14_ASAP7_75t_R g385 ( 
.A(n_339),
.Y(n_385)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_276),
.Y(n_340)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_340),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_SL g365 ( 
.A(n_341),
.B(n_343),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_286),
.B(n_240),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_SL g343 ( 
.A(n_312),
.B(n_242),
.Y(n_343)
);

OAI22xp33_ASAP7_75t_SL g344 ( 
.A1(n_305),
.A2(n_213),
.B1(n_212),
.B2(n_208),
.Y(n_344)
);

AOI22xp5_ASAP7_75t_L g369 ( 
.A1(n_344),
.A2(n_345),
.B1(n_355),
.B2(n_294),
.Y(n_369)
);

OAI22xp33_ASAP7_75t_SL g345 ( 
.A1(n_305),
.A2(n_207),
.B1(n_253),
.B2(n_258),
.Y(n_345)
);

INVx2_ASAP7_75t_L g346 ( 
.A(n_308),
.Y(n_346)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_346),
.Y(n_377)
);

AND2x2_ASAP7_75t_L g379 ( 
.A(n_347),
.B(n_360),
.Y(n_379)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_278),
.Y(n_348)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_348),
.Y(n_390)
);

XNOR2xp5_ASAP7_75t_L g389 ( 
.A(n_349),
.B(n_321),
.Y(n_389)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_278),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_L g363 ( 
.A(n_350),
.B(n_352),
.Y(n_363)
);

AOI21xp33_ASAP7_75t_L g351 ( 
.A1(n_304),
.A2(n_246),
.B(n_215),
.Y(n_351)
);

INVxp67_ASAP7_75t_L g393 ( 
.A(n_351),
.Y(n_393)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_280),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_280),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_L g384 ( 
.A(n_353),
.B(n_354),
.Y(n_384)
);

NOR2xp33_ASAP7_75t_L g354 ( 
.A(n_309),
.B(n_222),
.Y(n_354)
);

INVx4_ASAP7_75t_L g356 ( 
.A(n_310),
.Y(n_356)
);

INVx13_ASAP7_75t_L g382 ( 
.A(n_356),
.Y(n_382)
);

CKINVDCx20_ASAP7_75t_R g357 ( 
.A(n_288),
.Y(n_357)
);

NOR2xp33_ASAP7_75t_L g387 ( 
.A(n_357),
.B(n_358),
.Y(n_387)
);

NOR2xp33_ASAP7_75t_L g358 ( 
.A(n_311),
.B(n_306),
.Y(n_358)
);

OAI21xp5_ASAP7_75t_SL g359 ( 
.A1(n_315),
.A2(n_140),
.B(n_131),
.Y(n_359)
);

AOI21xp5_ASAP7_75t_L g375 ( 
.A1(n_359),
.A2(n_320),
.B(n_317),
.Y(n_375)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_284),
.Y(n_360)
);

AOI22xp5_ASAP7_75t_L g361 ( 
.A1(n_274),
.A2(n_238),
.B1(n_268),
.B2(n_227),
.Y(n_361)
);

OAI22xp5_ASAP7_75t_L g388 ( 
.A1(n_361),
.A2(n_362),
.B1(n_318),
.B2(n_295),
.Y(n_388)
);

INVx1_ASAP7_75t_SL g362 ( 
.A(n_281),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_SL g373 ( 
.A(n_362),
.B(n_283),
.Y(n_373)
);

MAJIxp5_ASAP7_75t_L g366 ( 
.A(n_349),
.B(n_314),
.C(n_296),
.Y(n_366)
);

MAJIxp5_ASAP7_75t_L g402 ( 
.A(n_366),
.B(n_378),
.C(n_380),
.Y(n_402)
);

NOR2xp33_ASAP7_75t_SL g400 ( 
.A(n_367),
.B(n_328),
.Y(n_400)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_369),
.Y(n_406)
);

OR2x2_ASAP7_75t_L g372 ( 
.A(n_327),
.B(n_316),
.Y(n_372)
);

OR2x2_ASAP7_75t_L g403 ( 
.A(n_372),
.B(n_327),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_373),
.B(n_284),
.Y(n_405)
);

AOI22xp5_ASAP7_75t_SL g374 ( 
.A1(n_330),
.A2(n_274),
.B1(n_285),
.B2(n_307),
.Y(n_374)
);

OAI21xp5_ASAP7_75t_SL g414 ( 
.A1(n_374),
.A2(n_375),
.B(n_376),
.Y(n_414)
);

AOI21xp5_ASAP7_75t_L g376 ( 
.A1(n_330),
.A2(n_304),
.B(n_297),
.Y(n_376)
);

XOR2xp5_ASAP7_75t_L g378 ( 
.A(n_324),
.B(n_314),
.Y(n_378)
);

MAJIxp5_ASAP7_75t_L g380 ( 
.A(n_333),
.B(n_319),
.C(n_275),
.Y(n_380)
);

AOI22xp5_ASAP7_75t_L g383 ( 
.A1(n_339),
.A2(n_279),
.B1(n_282),
.B2(n_273),
.Y(n_383)
);

OAI22xp5_ASAP7_75t_SL g399 ( 
.A1(n_383),
.A2(n_341),
.B1(n_328),
.B2(n_329),
.Y(n_399)
);

AOI22xp5_ASAP7_75t_SL g396 ( 
.A1(n_388),
.A2(n_326),
.B1(n_360),
.B2(n_353),
.Y(n_396)
);

MAJIxp5_ASAP7_75t_L g421 ( 
.A(n_389),
.B(n_300),
.C(n_298),
.Y(n_421)
);

OAI21xp5_ASAP7_75t_SL g392 ( 
.A1(n_339),
.A2(n_293),
.B(n_322),
.Y(n_392)
);

OAI21xp5_ASAP7_75t_L g404 ( 
.A1(n_392),
.A2(n_394),
.B(n_359),
.Y(n_404)
);

AOI21xp5_ASAP7_75t_L g394 ( 
.A1(n_335),
.A2(n_275),
.B(n_283),
.Y(n_394)
);

NOR2xp33_ASAP7_75t_L g395 ( 
.A(n_387),
.B(n_337),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_395),
.B(n_398),
.Y(n_424)
);

OAI22xp5_ASAP7_75t_SL g430 ( 
.A1(n_396),
.A2(n_400),
.B1(n_391),
.B2(n_394),
.Y(n_430)
);

XNOR2xp5_ASAP7_75t_L g397 ( 
.A(n_378),
.B(n_342),
.Y(n_397)
);

MAJIxp5_ASAP7_75t_L g427 ( 
.A(n_397),
.B(n_401),
.C(n_411),
.Y(n_427)
);

CKINVDCx20_ASAP7_75t_R g398 ( 
.A(n_363),
.Y(n_398)
);

AOI22xp5_ASAP7_75t_L g437 ( 
.A1(n_399),
.A2(n_409),
.B1(n_379),
.B2(n_380),
.Y(n_437)
);

XOR2xp5_ASAP7_75t_L g401 ( 
.A(n_378),
.B(n_329),
.Y(n_401)
);

OAI21xp5_ASAP7_75t_L g431 ( 
.A1(n_403),
.A2(n_385),
.B(n_381),
.Y(n_431)
);

AND2x2_ASAP7_75t_L g425 ( 
.A(n_404),
.B(n_418),
.Y(n_425)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_405),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_384),
.B(n_357),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g439 ( 
.A(n_407),
.B(n_408),
.Y(n_439)
);

CKINVDCx20_ASAP7_75t_R g408 ( 
.A(n_363),
.Y(n_408)
);

OAI22xp5_ASAP7_75t_SL g409 ( 
.A1(n_372),
.A2(n_326),
.B1(n_361),
.B2(n_347),
.Y(n_409)
);

NOR2xp33_ASAP7_75t_L g410 ( 
.A(n_387),
.B(n_386),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_410),
.B(n_413),
.Y(n_440)
);

XNOR2xp5_ASAP7_75t_L g411 ( 
.A(n_366),
.B(n_275),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_368),
.Y(n_412)
);

INVx1_ASAP7_75t_SL g428 ( 
.A(n_412),
.Y(n_428)
);

CKINVDCx20_ASAP7_75t_R g413 ( 
.A(n_384),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_371),
.B(n_338),
.Y(n_415)
);

HB1xp67_ASAP7_75t_L g441 ( 
.A(n_415),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_371),
.B(n_352),
.Y(n_416)
);

NOR2xp33_ASAP7_75t_L g429 ( 
.A(n_416),
.B(n_419),
.Y(n_429)
);

NOR2xp33_ASAP7_75t_L g417 ( 
.A(n_386),
.B(n_340),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_SL g426 ( 
.A(n_417),
.B(n_420),
.Y(n_426)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_368),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_370),
.B(n_350),
.Y(n_419)
);

AOI221xp5_ASAP7_75t_L g420 ( 
.A1(n_381),
.A2(n_393),
.B1(n_385),
.B2(n_367),
.C(n_365),
.Y(n_420)
);

XNOR2xp5_ASAP7_75t_L g432 ( 
.A(n_421),
.B(n_389),
.Y(n_432)
);

OAI22xp5_ASAP7_75t_SL g422 ( 
.A1(n_406),
.A2(n_365),
.B1(n_372),
.B2(n_383),
.Y(n_422)
);

AOI22xp5_ASAP7_75t_L g458 ( 
.A1(n_422),
.A2(n_409),
.B1(n_415),
.B2(n_379),
.Y(n_458)
);

XOR2xp5_ASAP7_75t_L g423 ( 
.A(n_402),
.B(n_411),
.Y(n_423)
);

XOR2xp5_ASAP7_75t_L g463 ( 
.A(n_423),
.B(n_432),
.Y(n_463)
);

NOR2xp33_ASAP7_75t_L g450 ( 
.A(n_430),
.B(n_408),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_431),
.B(n_444),
.Y(n_456)
);

XOR2xp5_ASAP7_75t_L g433 ( 
.A(n_402),
.B(n_366),
.Y(n_433)
);

MAJIxp5_ASAP7_75t_L g461 ( 
.A(n_433),
.B(n_435),
.C(n_407),
.Y(n_461)
);

NOR2xp33_ASAP7_75t_L g434 ( 
.A(n_400),
.B(n_306),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_SL g452 ( 
.A(n_434),
.B(n_436),
.Y(n_452)
);

XOR2xp5_ASAP7_75t_L g435 ( 
.A(n_401),
.B(n_380),
.Y(n_435)
);

NOR2xp33_ASAP7_75t_L g436 ( 
.A(n_413),
.B(n_287),
.Y(n_436)
);

OAI22xp5_ASAP7_75t_SL g454 ( 
.A1(n_437),
.A2(n_445),
.B1(n_396),
.B2(n_405),
.Y(n_454)
);

XNOR2xp5_ASAP7_75t_SL g442 ( 
.A(n_397),
.B(n_392),
.Y(n_442)
);

XNOR2xp5_ASAP7_75t_SL g448 ( 
.A(n_442),
.B(n_399),
.Y(n_448)
);

OAI21xp5_ASAP7_75t_L g443 ( 
.A1(n_414),
.A2(n_375),
.B(n_374),
.Y(n_443)
);

AOI21xp5_ASAP7_75t_L g449 ( 
.A1(n_443),
.A2(n_414),
.B(n_374),
.Y(n_449)
);

BUFx6f_ASAP7_75t_L g444 ( 
.A(n_398),
.Y(n_444)
);

AOI22xp5_ASAP7_75t_L g445 ( 
.A1(n_406),
.A2(n_379),
.B1(n_388),
.B2(n_390),
.Y(n_445)
);

INVx5_ASAP7_75t_L g446 ( 
.A(n_395),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_446),
.B(n_373),
.Y(n_462)
);

XNOR2xp5_ASAP7_75t_L g447 ( 
.A(n_432),
.B(n_404),
.Y(n_447)
);

XNOR2xp5_ASAP7_75t_L g481 ( 
.A(n_447),
.B(n_453),
.Y(n_481)
);

XOR2xp5_ASAP7_75t_L g469 ( 
.A(n_448),
.B(n_449),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_L g472 ( 
.A(n_450),
.B(n_451),
.Y(n_472)
);

CKINVDCx20_ASAP7_75t_R g451 ( 
.A(n_439),
.Y(n_451)
);

XNOR2xp5_ASAP7_75t_L g453 ( 
.A(n_423),
.B(n_421),
.Y(n_453)
);

AOI22xp5_ASAP7_75t_L g478 ( 
.A1(n_454),
.A2(n_460),
.B1(n_465),
.B2(n_446),
.Y(n_478)
);

XNOR2xp5_ASAP7_75t_SL g455 ( 
.A(n_442),
.B(n_403),
.Y(n_455)
);

XOR2xp5_ASAP7_75t_L g476 ( 
.A(n_455),
.B(n_457),
.Y(n_476)
);

XNOR2xp5_ASAP7_75t_L g457 ( 
.A(n_427),
.B(n_416),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g473 ( 
.A(n_458),
.B(n_464),
.Y(n_473)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_440),
.Y(n_459)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_459),
.Y(n_468)
);

OAI22xp5_ASAP7_75t_SL g460 ( 
.A1(n_437),
.A2(n_403),
.B1(n_410),
.B2(n_369),
.Y(n_460)
);

MAJIxp5_ASAP7_75t_L g467 ( 
.A(n_461),
.B(n_427),
.C(n_435),
.Y(n_467)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_462),
.Y(n_477)
);

AOI22xp5_ASAP7_75t_L g464 ( 
.A1(n_422),
.A2(n_379),
.B1(n_418),
.B2(n_412),
.Y(n_464)
);

OAI22xp5_ASAP7_75t_SL g465 ( 
.A1(n_445),
.A2(n_438),
.B1(n_426),
.B2(n_441),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_L g466 ( 
.A(n_424),
.B(n_417),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_L g479 ( 
.A(n_466),
.B(n_428),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_L g483 ( 
.A(n_467),
.B(n_470),
.Y(n_483)
);

MAJIxp5_ASAP7_75t_L g470 ( 
.A(n_463),
.B(n_433),
.C(n_425),
.Y(n_470)
);

MAJIxp5_ASAP7_75t_L g471 ( 
.A(n_463),
.B(n_425),
.C(n_443),
.Y(n_471)
);

MAJIxp5_ASAP7_75t_L g482 ( 
.A(n_471),
.B(n_474),
.C(n_475),
.Y(n_482)
);

MAJIxp5_ASAP7_75t_L g474 ( 
.A(n_461),
.B(n_425),
.C(n_444),
.Y(n_474)
);

MAJIxp5_ASAP7_75t_L g475 ( 
.A(n_453),
.B(n_431),
.C(n_429),
.Y(n_475)
);

OAI22xp5_ASAP7_75t_SL g493 ( 
.A1(n_478),
.A2(n_376),
.B1(n_390),
.B2(n_370),
.Y(n_493)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_479),
.Y(n_489)
);

NOR2xp33_ASAP7_75t_SL g480 ( 
.A(n_452),
.B(n_419),
.Y(n_480)
);

NOR2xp33_ASAP7_75t_L g490 ( 
.A(n_480),
.B(n_428),
.Y(n_490)
);

AOI21xp5_ASAP7_75t_L g484 ( 
.A1(n_474),
.A2(n_456),
.B(n_447),
.Y(n_484)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_484),
.Y(n_502)
);

INVxp33_ASAP7_75t_L g485 ( 
.A(n_472),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_L g501 ( 
.A(n_485),
.B(n_490),
.Y(n_501)
);

AOI22xp33_ASAP7_75t_SL g486 ( 
.A1(n_477),
.A2(n_460),
.B1(n_465),
.B2(n_454),
.Y(n_486)
);

OAI22xp5_ASAP7_75t_L g499 ( 
.A1(n_486),
.A2(n_347),
.B1(n_348),
.B2(n_377),
.Y(n_499)
);

XNOR2xp5_ASAP7_75t_SL g487 ( 
.A(n_469),
.B(n_448),
.Y(n_487)
);

XOR2xp5_ASAP7_75t_L g500 ( 
.A(n_487),
.B(n_493),
.Y(n_500)
);

AOI22xp5_ASAP7_75t_SL g488 ( 
.A1(n_471),
.A2(n_455),
.B1(n_458),
.B2(n_464),
.Y(n_488)
);

OAI22xp5_ASAP7_75t_SL g496 ( 
.A1(n_488),
.A2(n_473),
.B1(n_469),
.B2(n_476),
.Y(n_496)
);

XOR2xp5_ASAP7_75t_L g491 ( 
.A(n_481),
.B(n_457),
.Y(n_491)
);

XNOR2xp5_ASAP7_75t_L g497 ( 
.A(n_491),
.B(n_492),
.Y(n_497)
);

XOR2xp5_ASAP7_75t_L g492 ( 
.A(n_470),
.B(n_476),
.Y(n_492)
);

MAJIxp5_ASAP7_75t_L g494 ( 
.A(n_482),
.B(n_467),
.C(n_475),
.Y(n_494)
);

MAJIxp5_ASAP7_75t_L g506 ( 
.A(n_494),
.B(n_503),
.C(n_497),
.Y(n_506)
);

NOR2xp33_ASAP7_75t_SL g495 ( 
.A(n_485),
.B(n_468),
.Y(n_495)
);

NOR2xp33_ASAP7_75t_L g507 ( 
.A(n_495),
.B(n_498),
.Y(n_507)
);

AOI22xp5_ASAP7_75t_L g504 ( 
.A1(n_496),
.A2(n_499),
.B1(n_493),
.B2(n_488),
.Y(n_504)
);

NOR2xp33_ASAP7_75t_L g498 ( 
.A(n_489),
.B(n_356),
.Y(n_498)
);

MAJIxp5_ASAP7_75t_L g503 ( 
.A(n_482),
.B(n_377),
.C(n_364),
.Y(n_503)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_504),
.Y(n_512)
);

AOI322xp5_ASAP7_75t_L g505 ( 
.A1(n_502),
.A2(n_382),
.A3(n_483),
.B1(n_487),
.B2(n_491),
.C1(n_364),
.C2(n_492),
.Y(n_505)
);

AO21x1_ASAP7_75t_L g514 ( 
.A1(n_505),
.A2(n_510),
.B(n_511),
.Y(n_514)
);

NOR2xp33_ASAP7_75t_SL g513 ( 
.A(n_506),
.B(n_508),
.Y(n_513)
);

NOR2xp33_ASAP7_75t_L g508 ( 
.A(n_494),
.B(n_318),
.Y(n_508)
);

OAI21xp5_ASAP7_75t_SL g509 ( 
.A1(n_503),
.A2(n_382),
.B(n_347),
.Y(n_509)
);

AOI31xp67_ASAP7_75t_L g517 ( 
.A1(n_509),
.A2(n_281),
.A3(n_313),
.B(n_263),
.Y(n_517)
);

AOI322xp5_ASAP7_75t_L g510 ( 
.A1(n_501),
.A2(n_382),
.A3(n_310),
.B1(n_325),
.B2(n_346),
.C1(n_295),
.C2(n_302),
.Y(n_510)
);

NOR2xp33_ASAP7_75t_L g511 ( 
.A(n_497),
.B(n_301),
.Y(n_511)
);

OAI22xp33_ASAP7_75t_L g515 ( 
.A1(n_504),
.A2(n_500),
.B1(n_496),
.B2(n_279),
.Y(n_515)
);

OR2x2_ASAP7_75t_L g520 ( 
.A(n_515),
.B(n_516),
.Y(n_520)
);

OAI21xp5_ASAP7_75t_SL g516 ( 
.A1(n_506),
.A2(n_500),
.B(n_302),
.Y(n_516)
);

MAJIxp5_ASAP7_75t_L g518 ( 
.A(n_517),
.B(n_507),
.C(n_281),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_SL g523 ( 
.A(n_518),
.B(n_519),
.Y(n_523)
);

BUFx2_ASAP7_75t_L g519 ( 
.A(n_512),
.Y(n_519)
);

OAI21xp5_ASAP7_75t_SL g521 ( 
.A1(n_513),
.A2(n_289),
.B(n_299),
.Y(n_521)
);

AO21x1_ASAP7_75t_L g522 ( 
.A1(n_521),
.A2(n_289),
.B(n_299),
.Y(n_522)
);

MAJIxp5_ASAP7_75t_L g524 ( 
.A(n_522),
.B(n_514),
.C(n_301),
.Y(n_524)
);

OAI321xp33_ASAP7_75t_L g525 ( 
.A1(n_524),
.A2(n_523),
.A3(n_520),
.B1(n_261),
.B2(n_140),
.C(n_177),
.Y(n_525)
);

XNOR2x2_ASAP7_75t_SL g526 ( 
.A(n_525),
.B(n_177),
.Y(n_526)
);


endmodule