module real_jpeg_17371_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_356;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_288;
wire n_83;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_360;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;
wire n_364;

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_0),
.A2(n_161),
.B1(n_162),
.B2(n_163),
.Y(n_160)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_0),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g216 ( 
.A1(n_0),
.A2(n_162),
.B1(n_217),
.B2(n_219),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_0),
.A2(n_162),
.B1(n_280),
.B2(n_282),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_1),
.A2(n_111),
.B1(n_115),
.B2(n_116),
.Y(n_110)
);

CKINVDCx16_ASAP7_75t_R g115 ( 
.A(n_1),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_1),
.A2(n_115),
.B1(n_294),
.B2(n_297),
.Y(n_293)
);

AOI22xp33_ASAP7_75t_SL g304 ( 
.A1(n_1),
.A2(n_115),
.B1(n_305),
.B2(n_307),
.Y(n_304)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_2),
.Y(n_80)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_2),
.Y(n_90)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_3),
.Y(n_182)
);

BUFx5_ASAP7_75t_L g188 ( 
.A(n_3),
.Y(n_188)
);

BUFx6f_ASAP7_75t_L g196 ( 
.A(n_3),
.Y(n_196)
);

BUFx6f_ASAP7_75t_L g198 ( 
.A(n_3),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_SL g40 ( 
.A1(n_4),
.A2(n_41),
.B1(n_45),
.B2(n_47),
.Y(n_40)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_4),
.Y(n_47)
);

OAI22x1_ASAP7_75t_SL g120 ( 
.A1(n_5),
.A2(n_121),
.B1(n_123),
.B2(n_124),
.Y(n_120)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_5),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_5),
.A2(n_123),
.B1(n_202),
.B2(n_204),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_6),
.A2(n_169),
.B1(n_170),
.B2(n_173),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_6),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_6),
.A2(n_169),
.B1(n_235),
.B2(n_240),
.Y(n_234)
);

AOI22xp33_ASAP7_75t_L g102 ( 
.A1(n_7),
.A2(n_103),
.B1(n_107),
.B2(n_108),
.Y(n_102)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_7),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_7),
.A2(n_108),
.B1(n_147),
.B2(n_155),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_7),
.A2(n_108),
.B1(n_270),
.B2(n_275),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_SL g327 ( 
.A1(n_7),
.A2(n_46),
.B1(n_108),
.B2(n_328),
.Y(n_327)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_8),
.Y(n_130)
);

BUFx5_ASAP7_75t_L g333 ( 
.A(n_8),
.Y(n_333)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_9),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_9),
.B(n_132),
.Y(n_131)
);

OAI32xp33_ASAP7_75t_L g226 ( 
.A1(n_9),
.A2(n_77),
.A3(n_170),
.B1(n_227),
.B2(n_230),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_9),
.B(n_109),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_SL g326 ( 
.A1(n_9),
.A2(n_23),
.B1(n_311),
.B2(n_327),
.Y(n_326)
);

AOI22xp33_ASAP7_75t_SL g346 ( 
.A1(n_9),
.A2(n_50),
.B1(n_347),
.B2(n_349),
.Y(n_346)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_10),
.Y(n_95)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_10),
.Y(n_100)
);

INVx3_ASAP7_75t_L g177 ( 
.A(n_10),
.Y(n_177)
);

BUFx6f_ASAP7_75t_L g193 ( 
.A(n_10),
.Y(n_193)
);

BUFx3_ASAP7_75t_L g206 ( 
.A(n_10),
.Y(n_206)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_10),
.Y(n_274)
);

OAI22xp33_ASAP7_75t_L g30 ( 
.A1(n_11),
.A2(n_31),
.B1(n_32),
.B2(n_33),
.Y(n_30)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

BUFx5_ASAP7_75t_L g58 ( 
.A(n_12),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_12),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g143 ( 
.A(n_12),
.Y(n_143)
);

INVx6_ASAP7_75t_L g153 ( 
.A(n_12),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_13),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_13),
.Y(n_85)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_14),
.Y(n_37)
);

BUFx4f_ASAP7_75t_L g44 ( 
.A(n_14),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g186 ( 
.A(n_14),
.Y(n_186)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_15),
.Y(n_54)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_15),
.Y(n_72)
);

BUFx8_ASAP7_75t_L g148 ( 
.A(n_15),
.Y(n_148)
);

BUFx5_ASAP7_75t_L g157 ( 
.A(n_15),
.Y(n_157)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_244),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_242),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_SL g18 ( 
.A(n_19),
.B(n_209),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_19),
.B(n_209),
.Y(n_243)
);

XOR2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_144),
.Y(n_19)
);

XNOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_73),
.Y(n_20)
);

XOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_48),
.Y(n_21)
);

OAI22xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_29),
.B1(n_38),
.B2(n_40),
.Y(n_22)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_23),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g278 ( 
.A1(n_23),
.A2(n_279),
.B1(n_287),
.B2(n_288),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_SL g330 ( 
.A1(n_23),
.A2(n_304),
.B1(n_327),
.B2(n_331),
.Y(n_330)
);

OR2x2_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_27),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_26),
.Y(n_39)
);

INVx2_ASAP7_75t_L g287 ( 
.A(n_26),
.Y(n_287)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_27),
.Y(n_31)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_27),
.Y(n_252)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_28),
.Y(n_46)
);

INVx4_ASAP7_75t_L g122 ( 
.A(n_28),
.Y(n_122)
);

INVx3_ASAP7_75t_L g183 ( 
.A(n_28),
.Y(n_183)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_28),
.Y(n_239)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

AOI22x1_ASAP7_75t_SL g118 ( 
.A1(n_30),
.A2(n_119),
.B1(n_120),
.B2(n_127),
.Y(n_118)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_35),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx3_ASAP7_75t_L g309 ( 
.A(n_36),
.Y(n_309)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g240 ( 
.A(n_43),
.Y(n_240)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx3_ASAP7_75t_L g262 ( 
.A(n_44),
.Y(n_262)
);

BUFx6f_ASAP7_75t_L g281 ( 
.A(n_44),
.Y(n_281)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g48 ( 
.A1(n_49),
.A2(n_55),
.B1(n_66),
.B2(n_68),
.Y(n_48)
);

OAI21xp33_ASAP7_75t_SL g146 ( 
.A1(n_49),
.A2(n_50),
.B(n_147),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_50),
.B(n_51),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_50),
.B(n_231),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_50),
.B(n_255),
.Y(n_254)
);

OAI21xp33_ASAP7_75t_SL g265 ( 
.A1(n_50),
.A2(n_254),
.B(n_266),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_SL g325 ( 
.A(n_50),
.B(n_128),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_50),
.B(n_208),
.Y(n_334)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_56),
.B(n_59),
.Y(n_55)
);

BUFx2_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

AND2x2_ASAP7_75t_L g69 ( 
.A(n_57),
.B(n_70),
.Y(n_69)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

BUFx2_ASAP7_75t_L g107 ( 
.A(n_62),
.Y(n_107)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx8_ASAP7_75t_L g67 ( 
.A(n_63),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g166 ( 
.A(n_64),
.Y(n_166)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_65),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_65),
.Y(n_114)
);

BUFx5_ASAP7_75t_L g138 ( 
.A(n_65),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g141 ( 
.A(n_65),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVxp67_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

OA21x2_ASAP7_75t_L g149 ( 
.A1(n_69),
.A2(n_133),
.B(n_150),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_70),
.B(n_151),
.Y(n_150)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

MAJIxp5_ASAP7_75t_L g73 ( 
.A(n_74),
.B(n_118),
.C(n_131),
.Y(n_73)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_74),
.B(n_212),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_75),
.A2(n_101),
.B1(n_109),
.B2(n_110),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_75),
.A2(n_109),
.B1(n_110),
.B2(n_160),
.Y(n_159)
);

INVx1_ASAP7_75t_SL g75 ( 
.A(n_76),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g345 ( 
.A1(n_76),
.A2(n_102),
.B1(n_346),
.B2(n_354),
.Y(n_345)
);

AO21x2_ASAP7_75t_SL g76 ( 
.A1(n_77),
.A2(n_86),
.B(n_94),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_78),
.B(n_81),
.Y(n_77)
);

INVx6_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_80),
.Y(n_97)
);

BUFx5_ASAP7_75t_L g98 ( 
.A(n_80),
.Y(n_98)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

BUFx3_ASAP7_75t_L g161 ( 
.A(n_83),
.Y(n_161)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_85),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_91),
.Y(n_86)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVx6_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

BUFx2_ASAP7_75t_L g109 ( 
.A(n_94),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_95),
.A2(n_96),
.B1(n_98),
.B2(n_99),
.Y(n_94)
);

BUFx3_ASAP7_75t_L g203 ( 
.A(n_95),
.Y(n_203)
);

INVx4_ASAP7_75t_L g218 ( 
.A(n_95),
.Y(n_218)
);

INVx5_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx6_ASAP7_75t_L g251 ( 
.A(n_99),
.Y(n_251)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVxp67_ASAP7_75t_SL g172 ( 
.A(n_100),
.Y(n_172)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

HB1xp67_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

BUFx2_ASAP7_75t_SL g104 ( 
.A(n_105),
.Y(n_104)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

BUFx3_ASAP7_75t_L g229 ( 
.A(n_106),
.Y(n_229)
);

INVx2_ASAP7_75t_L g354 ( 
.A(n_109),
.Y(n_354)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_114),
.Y(n_117)
);

INVx2_ASAP7_75t_L g353 ( 
.A(n_114),
.Y(n_353)
);

BUFx2_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

XOR2xp5_ASAP7_75t_L g212 ( 
.A(n_118),
.B(n_131),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_119),
.A2(n_120),
.B1(n_234),
.B2(n_241),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g302 ( 
.A1(n_119),
.A2(n_303),
.B1(n_310),
.B2(n_312),
.Y(n_302)
);

BUFx2_ASAP7_75t_L g328 ( 
.A(n_121),
.Y(n_328)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

HB1xp67_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVx6_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVx6_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g241 ( 
.A(n_129),
.Y(n_241)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_132),
.A2(n_146),
.B1(n_149),
.B2(n_154),
.Y(n_145)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

AOI22x1_ASAP7_75t_L g133 ( 
.A1(n_134),
.A2(n_137),
.B1(n_139),
.B2(n_142),
.Y(n_133)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx3_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

INVx3_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVx3_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

XOR2xp5_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_158),
.Y(n_144)
);

BUFx12f_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

INVx3_ASAP7_75t_SL g152 ( 
.A(n_153),
.Y(n_152)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

BUFx2_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_167),
.Y(n_158)
);

INVx8_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g348 ( 
.A(n_166),
.Y(n_348)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_168),
.A2(n_178),
.B1(n_200),
.B2(n_207),
.Y(n_167)
);

INVxp67_ASAP7_75t_L g223 ( 
.A(n_168),
.Y(n_223)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

HB1xp67_ASAP7_75t_L g231 ( 
.A(n_175),
.Y(n_231)
);

INVx5_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_178),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_178),
.A2(n_207),
.B1(n_265),
.B2(n_269),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_178),
.A2(n_207),
.B1(n_269),
.B2(n_293),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_L g356 ( 
.A1(n_178),
.A2(n_207),
.B1(n_216),
.B2(n_293),
.Y(n_356)
);

AND2x2_ASAP7_75t_SL g178 ( 
.A(n_179),
.B(n_189),
.Y(n_178)
);

BUFx3_ASAP7_75t_L g208 ( 
.A(n_179),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_180),
.A2(n_183),
.B1(n_184),
.B2(n_187),
.Y(n_179)
);

INVx8_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

BUFx6f_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

INVx5_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_186),
.Y(n_286)
);

BUFx3_ASAP7_75t_L g306 ( 
.A(n_186),
.Y(n_306)
);

INVx3_ASAP7_75t_L g324 ( 
.A(n_186),
.Y(n_324)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_188),
.Y(n_259)
);

OAI22xp33_ASAP7_75t_L g189 ( 
.A1(n_190),
.A2(n_194),
.B1(n_197),
.B2(n_199),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_192),
.Y(n_199)
);

INVx6_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_193),
.Y(n_222)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

INVx6_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

INVx4_ASAP7_75t_L g253 ( 
.A(n_197),
.Y(n_253)
);

INVx6_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

INVxp67_ASAP7_75t_SL g200 ( 
.A(n_201),
.Y(n_200)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

INVx2_ASAP7_75t_L g298 ( 
.A(n_205),
.Y(n_298)
);

INVx3_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_208),
.A2(n_214),
.B1(n_215),
.B2(n_223),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_210),
.B(n_213),
.C(n_224),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g359 ( 
.A1(n_210),
.A2(n_211),
.B1(n_360),
.B2(n_361),
.Y(n_359)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g361 ( 
.A1(n_213),
.A2(n_224),
.B1(n_225),
.B2(n_362),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_213),
.Y(n_362)
);

INVxp67_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_218),
.Y(n_268)
);

INVx4_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

BUFx6f_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

INVx5_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_232),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g341 ( 
.A1(n_226),
.A2(n_232),
.B1(n_233),
.B2(n_342),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_226),
.Y(n_342)
);

INVx3_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

BUFx6f_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_231),
.Y(n_255)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

INVxp67_ASAP7_75t_L g288 ( 
.A(n_234),
.Y(n_288)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

HB1xp67_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

INVx2_ASAP7_75t_L g311 ( 
.A(n_241),
.Y(n_311)
);

INVxp67_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

OAI21x1_ASAP7_75t_L g244 ( 
.A1(n_245),
.A2(n_358),
.B(n_364),
.Y(n_244)
);

AOI21x1_ASAP7_75t_SL g245 ( 
.A1(n_246),
.A2(n_338),
.B(n_357),
.Y(n_245)
);

OAI21x1_ASAP7_75t_L g246 ( 
.A1(n_247),
.A2(n_300),
.B(n_337),
.Y(n_246)
);

AND2x2_ASAP7_75t_L g247 ( 
.A(n_248),
.B(n_277),
.Y(n_247)
);

OR2x2_ASAP7_75t_L g337 ( 
.A(n_248),
.B(n_277),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_249),
.B(n_263),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g313 ( 
.A1(n_249),
.A2(n_263),
.B1(n_264),
.B2(n_314),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_249),
.Y(n_314)
);

OAI32xp33_ASAP7_75t_L g249 ( 
.A1(n_250),
.A2(n_252),
.A3(n_253),
.B1(n_254),
.B2(n_256),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_257),
.B(n_260),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

BUFx3_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

INVx3_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_274),
.Y(n_276)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_274),
.Y(n_296)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_278),
.B(n_289),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g339 ( 
.A(n_278),
.B(n_291),
.C(n_299),
.Y(n_339)
);

INVxp67_ASAP7_75t_L g312 ( 
.A(n_279),
.Y(n_312)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

BUFx2_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_L g289 ( 
.A1(n_290),
.A2(n_291),
.B1(n_292),
.B2(n_299),
.Y(n_289)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_290),
.Y(n_299)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

INVx3_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

AOI21xp5_ASAP7_75t_L g300 ( 
.A1(n_301),
.A2(n_315),
.B(n_336),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_302),
.B(n_313),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_302),
.B(n_313),
.Y(n_336)
);

INVxp67_ASAP7_75t_L g303 ( 
.A(n_304),
.Y(n_303)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_306),
.Y(n_305)
);

INVx2_ASAP7_75t_L g307 ( 
.A(n_308),
.Y(n_307)
);

INVx2_ASAP7_75t_SL g308 ( 
.A(n_309),
.Y(n_308)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_311),
.Y(n_310)
);

OAI21xp5_ASAP7_75t_L g315 ( 
.A1(n_316),
.A2(n_329),
.B(n_335),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_317),
.B(n_326),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_318),
.B(n_325),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_319),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

HB1xp67_ASAP7_75t_L g320 ( 
.A(n_321),
.Y(n_320)
);

INVx2_ASAP7_75t_L g321 ( 
.A(n_322),
.Y(n_321)
);

BUFx6f_ASAP7_75t_L g322 ( 
.A(n_323),
.Y(n_322)
);

INVx2_ASAP7_75t_L g323 ( 
.A(n_324),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_330),
.B(n_334),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_330),
.B(n_334),
.Y(n_335)
);

INVx6_ASAP7_75t_L g331 ( 
.A(n_332),
.Y(n_331)
);

BUFx12f_ASAP7_75t_L g332 ( 
.A(n_333),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_339),
.B(n_340),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g357 ( 
.A(n_339),
.B(n_340),
.Y(n_357)
);

XOR2xp5_ASAP7_75t_L g340 ( 
.A(n_341),
.B(n_343),
.Y(n_340)
);

MAJIxp5_ASAP7_75t_L g363 ( 
.A(n_341),
.B(n_344),
.C(n_356),
.Y(n_363)
);

OAI22xp5_ASAP7_75t_SL g343 ( 
.A1(n_344),
.A2(n_345),
.B1(n_355),
.B2(n_356),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_345),
.Y(n_344)
);

BUFx2_ASAP7_75t_L g347 ( 
.A(n_348),
.Y(n_347)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_350),
.Y(n_349)
);

BUFx2_ASAP7_75t_L g350 ( 
.A(n_351),
.Y(n_350)
);

INVx2_ASAP7_75t_L g351 ( 
.A(n_352),
.Y(n_351)
);

INVx2_ASAP7_75t_L g352 ( 
.A(n_353),
.Y(n_352)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_356),
.Y(n_355)
);

NOR2xp67_ASAP7_75t_SL g358 ( 
.A(n_359),
.B(n_363),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_359),
.B(n_363),
.Y(n_364)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_361),
.Y(n_360)
);


endmodule