module fake_jpeg_27822_n_313 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_313);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_313;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx11_ASAP7_75t_L g16 ( 
.A(n_13),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_2),
.Y(n_18)
);

CKINVDCx16_ASAP7_75t_R g19 ( 
.A(n_8),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_9),
.Y(n_20)
);

INVx11_ASAP7_75t_SL g21 ( 
.A(n_7),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

INVx6_ASAP7_75t_SL g24 ( 
.A(n_1),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

INVx11_ASAP7_75t_SL g27 ( 
.A(n_9),
.Y(n_27)
);

INVx13_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_8),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_17),
.Y(n_33)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_33),
.Y(n_55)
);

INVx4_ASAP7_75t_SL g34 ( 
.A(n_21),
.Y(n_34)
);

INVxp67_ASAP7_75t_L g62 ( 
.A(n_34),
.Y(n_62)
);

INVx5_ASAP7_75t_L g35 ( 
.A(n_28),
.Y(n_35)
);

INVx11_ASAP7_75t_L g43 ( 
.A(n_35),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_16),
.Y(n_37)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_37),
.Y(n_44)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_16),
.Y(n_38)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_38),
.Y(n_47)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_21),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_39),
.B(n_19),
.Y(n_60)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_17),
.Y(n_40)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_40),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_16),
.Y(n_41)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_41),
.Y(n_45)
);

BUFx2_ASAP7_75t_L g42 ( 
.A(n_27),
.Y(n_42)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_42),
.Y(n_59)
);

INVx5_ASAP7_75t_L g46 ( 
.A(n_38),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_46),
.Y(n_87)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_37),
.Y(n_48)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_48),
.Y(n_85)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_37),
.Y(n_49)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_49),
.Y(n_88)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_50),
.Y(n_80)
);

INVx6_ASAP7_75t_SL g52 ( 
.A(n_34),
.Y(n_52)
);

CKINVDCx14_ASAP7_75t_R g78 ( 
.A(n_52),
.Y(n_78)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_41),
.Y(n_53)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_53),
.Y(n_70)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_54),
.B(n_56),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_42),
.Y(n_56)
);

HB1xp67_ASAP7_75t_L g57 ( 
.A(n_34),
.Y(n_57)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_57),
.Y(n_64)
);

AND2x2_ASAP7_75t_L g66 ( 
.A(n_60),
.B(n_28),
.Y(n_66)
);

BUFx5_ASAP7_75t_L g61 ( 
.A(n_42),
.Y(n_61)
);

CKINVDCx14_ASAP7_75t_R g82 ( 
.A(n_61),
.Y(n_82)
);

NOR2xp67_ASAP7_75t_L g63 ( 
.A(n_41),
.B(n_26),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_SL g77 ( 
.A(n_63),
.B(n_26),
.Y(n_77)
);

A2O1A1Ixp33_ASAP7_75t_L g65 ( 
.A1(n_60),
.A2(n_20),
.B(n_29),
.C(n_19),
.Y(n_65)
);

XOR2xp5_ASAP7_75t_L g107 ( 
.A(n_65),
.B(n_25),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_66),
.B(n_69),
.Y(n_115)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_48),
.Y(n_67)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_67),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_59),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_68),
.B(n_73),
.Y(n_101)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_58),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_58),
.B(n_22),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_71),
.B(n_81),
.Y(n_91)
);

INVx8_ASAP7_75t_L g72 ( 
.A(n_47),
.Y(n_72)
);

INVx5_ASAP7_75t_L g108 ( 
.A(n_72),
.Y(n_108)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_43),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_55),
.A2(n_40),
.B1(n_33),
.B2(n_22),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_74),
.A2(n_75),
.B1(n_83),
.B2(n_34),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_55),
.A2(n_40),
.B1(n_33),
.B2(n_22),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_77),
.B(n_79),
.Y(n_104)
);

INVx1_ASAP7_75t_SL g79 ( 
.A(n_52),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_59),
.B(n_25),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_L g83 ( 
.A1(n_51),
.A2(n_28),
.B1(n_27),
.B2(n_26),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_61),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_84),
.B(n_90),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_44),
.B(n_18),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_86),
.B(n_18),
.Y(n_98)
);

INVx5_ASAP7_75t_L g89 ( 
.A(n_43),
.Y(n_89)
);

INVx2_ASAP7_75t_SL g99 ( 
.A(n_89),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_62),
.B(n_20),
.Y(n_90)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_86),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_92),
.B(n_93),
.Y(n_121)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_71),
.Y(n_93)
);

AOI21xp5_ASAP7_75t_L g95 ( 
.A1(n_66),
.A2(n_0),
.B(n_1),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_95),
.B(n_98),
.Y(n_124)
);

NAND2xp33_ASAP7_75t_SL g96 ( 
.A(n_66),
.B(n_42),
.Y(n_96)
);

OR2x2_ASAP7_75t_L g136 ( 
.A(n_96),
.B(n_103),
.Y(n_136)
);

INVx13_ASAP7_75t_L g97 ( 
.A(n_79),
.Y(n_97)
);

INVx5_ASAP7_75t_L g142 ( 
.A(n_97),
.Y(n_142)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_85),
.Y(n_100)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_100),
.Y(n_119)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_70),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_102),
.B(n_106),
.Y(n_125)
);

NAND2xp33_ASAP7_75t_SL g103 ( 
.A(n_77),
.B(n_35),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_72),
.A2(n_29),
.B1(n_20),
.B2(n_46),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_105),
.A2(n_110),
.B1(n_51),
.B2(n_49),
.Y(n_120)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_70),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_107),
.B(n_112),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_89),
.A2(n_29),
.B1(n_54),
.B2(n_35),
.Y(n_110)
);

INVx4_ASAP7_75t_L g111 ( 
.A(n_87),
.Y(n_111)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_111),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_81),
.B(n_50),
.Y(n_112)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_76),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_113),
.B(n_114),
.Y(n_133)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_78),
.Y(n_114)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_85),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_116),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_117),
.A2(n_74),
.B1(n_69),
.B2(n_67),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_68),
.B(n_28),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_118),
.B(n_98),
.Y(n_138)
);

OAI21xp33_ASAP7_75t_SL g147 ( 
.A1(n_120),
.A2(n_111),
.B(n_94),
.Y(n_147)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_101),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_122),
.B(n_123),
.Y(n_160)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_118),
.Y(n_123)
);

AND2x6_ASAP7_75t_L g126 ( 
.A(n_103),
.B(n_65),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_126),
.B(n_135),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_109),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_129),
.Y(n_152)
);

CKINVDCx5p33_ASAP7_75t_R g131 ( 
.A(n_97),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_131),
.B(n_139),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_132),
.A2(n_137),
.B1(n_141),
.B2(n_127),
.Y(n_162)
);

INVx3_ASAP7_75t_L g134 ( 
.A(n_99),
.Y(n_134)
);

INVx6_ASAP7_75t_L g150 ( 
.A(n_134),
.Y(n_150)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_112),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_93),
.B(n_64),
.C(n_75),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_L g166 ( 
.A(n_137),
.B(n_141),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_138),
.B(n_140),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_113),
.B(n_104),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_91),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_115),
.B(n_64),
.C(n_87),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_92),
.A2(n_53),
.B1(n_45),
.B2(n_44),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_143),
.A2(n_117),
.B1(n_106),
.B2(n_102),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_132),
.A2(n_91),
.B1(n_108),
.B2(n_115),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_144),
.A2(n_149),
.B1(n_155),
.B2(n_168),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_L g177 ( 
.A1(n_145),
.A2(n_156),
.B1(n_162),
.B2(n_164),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_SL g179 ( 
.A1(n_147),
.A2(n_161),
.B(n_19),
.Y(n_179)
);

CKINVDCx16_ASAP7_75t_R g148 ( 
.A(n_125),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_148),
.B(n_157),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_135),
.A2(n_107),
.B1(n_108),
.B2(n_94),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_140),
.B(n_95),
.Y(n_153)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_153),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_L g154 ( 
.A1(n_136),
.A2(n_96),
.B(n_25),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_L g171 ( 
.A1(n_154),
.A2(n_124),
.B(n_122),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_123),
.A2(n_88),
.B1(n_45),
.B2(n_99),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_SL g156 ( 
.A1(n_134),
.A2(n_99),
.B1(n_97),
.B2(n_84),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_128),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_143),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_158),
.B(n_163),
.Y(n_193)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_119),
.Y(n_159)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_159),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_SL g161 ( 
.A1(n_136),
.A2(n_82),
.B(n_62),
.Y(n_161)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_119),
.Y(n_163)
);

AOI22xp33_ASAP7_75t_SL g164 ( 
.A1(n_142),
.A2(n_73),
.B1(n_47),
.B2(n_88),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_129),
.B(n_116),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_SL g184 ( 
.A(n_167),
.B(n_128),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_121),
.A2(n_100),
.B1(n_87),
.B2(n_80),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_126),
.A2(n_80),
.B1(n_39),
.B2(n_32),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_169),
.A2(n_24),
.B1(n_30),
.B2(n_17),
.Y(n_196)
);

AND2x4_ASAP7_75t_SL g170 ( 
.A(n_161),
.B(n_127),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_170),
.B(n_181),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_171),
.B(n_190),
.Y(n_205)
);

AOI21xp5_ASAP7_75t_L g173 ( 
.A1(n_165),
.A2(n_124),
.B(n_133),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_173),
.B(n_176),
.Y(n_209)
);

AOI22xp33_ASAP7_75t_SL g175 ( 
.A1(n_150),
.A2(n_142),
.B1(n_130),
.B2(n_131),
.Y(n_175)
);

CKINVDCx16_ASAP7_75t_R g201 ( 
.A(n_175),
.Y(n_201)
);

AND2x6_ASAP7_75t_L g176 ( 
.A(n_162),
.B(n_14),
.Y(n_176)
);

CKINVDCx12_ASAP7_75t_R g178 ( 
.A(n_152),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_178),
.B(n_179),
.Y(n_199)
);

AND2x2_ASAP7_75t_L g180 ( 
.A(n_149),
.B(n_130),
.Y(n_180)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_180),
.Y(n_202)
);

INVxp67_ASAP7_75t_L g181 ( 
.A(n_146),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_168),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_182),
.B(n_186),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_184),
.B(n_185),
.Y(n_212)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_155),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_160),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_158),
.A2(n_32),
.B1(n_23),
.B2(n_18),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_187),
.A2(n_196),
.B1(n_24),
.B2(n_30),
.Y(n_208)
);

INVx5_ASAP7_75t_SL g188 ( 
.A(n_150),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_188),
.B(n_31),
.Y(n_217)
);

OAI21xp5_ASAP7_75t_L g190 ( 
.A1(n_154),
.A2(n_32),
.B(n_23),
.Y(n_190)
);

OAI21xp33_ASAP7_75t_L g191 ( 
.A1(n_152),
.A2(n_23),
.B(n_12),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_191),
.Y(n_211)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_169),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_192),
.B(n_30),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_SL g194 ( 
.A(n_151),
.B(n_26),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_SL g200 ( 
.A(n_194),
.B(n_151),
.Y(n_200)
);

XOR2xp5_ASAP7_75t_L g195 ( 
.A(n_166),
.B(n_30),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_195),
.B(n_166),
.C(n_145),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_200),
.B(n_203),
.Y(n_233)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_193),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_L g237 ( 
.A(n_204),
.B(n_206),
.Y(n_237)
);

A2O1A1O1Ixp25_ASAP7_75t_L g206 ( 
.A1(n_171),
.A2(n_153),
.B(n_144),
.C(n_24),
.D(n_157),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_195),
.B(n_163),
.C(n_159),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_207),
.B(n_219),
.C(n_31),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_L g224 ( 
.A1(n_208),
.A2(n_213),
.B1(n_182),
.B2(n_190),
.Y(n_224)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_189),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_210),
.B(n_215),
.Y(n_228)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_172),
.Y(n_214)
);

AOI22xp33_ASAP7_75t_L g223 ( 
.A1(n_214),
.A2(n_217),
.B1(n_188),
.B2(n_172),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_SL g215 ( 
.A(n_186),
.B(n_10),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_180),
.Y(n_216)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_216),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_181),
.B(n_174),
.Y(n_218)
);

HB1xp67_ASAP7_75t_L g238 ( 
.A(n_218),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_174),
.B(n_36),
.C(n_31),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_204),
.B(n_173),
.Y(n_220)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_220),
.B(n_229),
.Y(n_242)
);

AOI21xp5_ASAP7_75t_SL g221 ( 
.A1(n_197),
.A2(n_179),
.B(n_176),
.Y(n_221)
);

CKINVDCx14_ASAP7_75t_R g245 ( 
.A(n_221),
.Y(n_245)
);

XOR2x2_ASAP7_75t_L g222 ( 
.A(n_197),
.B(n_170),
.Y(n_222)
);

INVxp67_ASAP7_75t_L g240 ( 
.A(n_222),
.Y(n_240)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_223),
.Y(n_255)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_224),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_201),
.A2(n_177),
.B1(n_183),
.B2(n_180),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_L g241 ( 
.A1(n_226),
.A2(n_227),
.B1(n_234),
.B2(n_208),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_212),
.A2(n_183),
.B1(n_170),
.B2(n_187),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_SL g229 ( 
.A(n_205),
.B(n_30),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_207),
.B(n_31),
.Y(n_230)
);

XOR2xp5_ASAP7_75t_L g252 ( 
.A(n_230),
.B(n_235),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_231),
.B(n_239),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_L g232 ( 
.A1(n_209),
.A2(n_9),
.B1(n_15),
.B2(n_3),
.Y(n_232)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_232),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_202),
.A2(n_17),
.B1(n_31),
.B2(n_3),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g235 ( 
.A(n_205),
.B(n_17),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_L g236 ( 
.A1(n_211),
.A2(n_8),
.B1(n_15),
.B2(n_4),
.Y(n_236)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_236),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_199),
.B(n_7),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_241),
.A2(n_203),
.B1(n_211),
.B2(n_206),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_225),
.A2(n_202),
.B1(n_216),
.B2(n_222),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_244),
.A2(n_198),
.B1(n_218),
.B2(n_219),
.Y(n_264)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_238),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_247),
.B(n_249),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_233),
.B(n_210),
.Y(n_248)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_248),
.Y(n_257)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_223),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_228),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_250),
.B(n_253),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_221),
.Y(n_253)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_256),
.Y(n_282)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_244),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_259),
.B(n_260),
.Y(n_280)
);

INVx13_ASAP7_75t_L g260 ( 
.A(n_245),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_255),
.A2(n_198),
.B1(n_237),
.B2(n_231),
.Y(n_261)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_261),
.Y(n_274)
);

AOI21xp5_ASAP7_75t_L g262 ( 
.A1(n_240),
.A2(n_254),
.B(n_255),
.Y(n_262)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_262),
.Y(n_278)
);

XNOR2x1_ASAP7_75t_L g263 ( 
.A(n_242),
.B(n_240),
.Y(n_263)
);

MAJx2_ASAP7_75t_L g271 ( 
.A(n_263),
.B(n_266),
.C(n_269),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_264),
.A2(n_252),
.B1(n_2),
.B2(n_0),
.Y(n_272)
);

XOR2x1_ASAP7_75t_SL g266 ( 
.A(n_242),
.B(n_229),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_251),
.B(n_230),
.Y(n_267)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_267),
.Y(n_281)
);

OAI21xp5_ASAP7_75t_L g268 ( 
.A1(n_246),
.A2(n_217),
.B(n_214),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_268),
.B(n_252),
.C(n_36),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_243),
.A2(n_220),
.B1(n_235),
.B2(n_4),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_257),
.B(n_251),
.Y(n_270)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_270),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_SL g291 ( 
.A1(n_272),
.A2(n_279),
.B1(n_276),
.B2(n_271),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_264),
.B(n_260),
.Y(n_273)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_273),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_275),
.B(n_256),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_261),
.B(n_11),
.C(n_5),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_276),
.B(n_277),
.C(n_279),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_263),
.B(n_11),
.C(n_5),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_269),
.B(n_11),
.C(n_5),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_SL g298 ( 
.A(n_284),
.B(n_291),
.Y(n_298)
);

XOR2xp5_ASAP7_75t_L g285 ( 
.A(n_277),
.B(n_266),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_285),
.B(n_288),
.C(n_289),
.Y(n_295)
);

AOI21xp5_ASAP7_75t_L g286 ( 
.A1(n_278),
.A2(n_265),
.B(n_258),
.Y(n_286)
);

OAI21xp5_ASAP7_75t_SL g293 ( 
.A1(n_286),
.A2(n_271),
.B(n_6),
.Y(n_293)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_280),
.B(n_268),
.Y(n_288)
);

XOR2xp5_ASAP7_75t_L g289 ( 
.A(n_274),
.B(n_282),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_281),
.A2(n_6),
.B1(n_7),
.B2(n_12),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_292),
.B(n_6),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_293),
.B(n_294),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_L g294 ( 
.A(n_285),
.B(n_14),
.Y(n_294)
);

BUFx24_ASAP7_75t_SL g296 ( 
.A(n_283),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_296),
.B(n_297),
.Y(n_305)
);

INVx1_ASAP7_75t_SL g297 ( 
.A(n_288),
.Y(n_297)
);

INVxp33_ASAP7_75t_SL g303 ( 
.A(n_299),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_287),
.B(n_12),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_300),
.B(n_287),
.C(n_290),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_301),
.B(n_302),
.Y(n_306)
);

NOR2xp67_ASAP7_75t_L g302 ( 
.A(n_298),
.B(n_289),
.Y(n_302)
);

INVxp67_ASAP7_75t_L g307 ( 
.A(n_305),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_307),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_308),
.B(n_303),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_SL g310 ( 
.A1(n_309),
.A2(n_306),
.B1(n_295),
.B2(n_304),
.Y(n_310)
);

BUFx24_ASAP7_75t_SL g311 ( 
.A(n_310),
.Y(n_311)
);

A2O1A1O1Ixp25_ASAP7_75t_L g312 ( 
.A1(n_311),
.A2(n_0),
.B(n_13),
.C(n_14),
.D(n_306),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_312),
.B(n_13),
.Y(n_313)
);


endmodule