module fake_aes_985_n_1320 (n_117, n_219, n_44, n_133, n_149, n_289, n_220, n_81, n_69, n_214, n_267, n_204, n_221, n_249, n_185, n_22, n_203, n_57, n_88, n_52, n_244, n_26, n_50, n_33, n_102, n_73, n_49, n_119, n_141, n_115, n_97, n_80, n_167, n_284, n_107, n_158, n_278, n_60, n_114, n_121, n_41, n_35, n_94, n_65, n_171, n_196, n_125, n_192, n_240, n_254, n_9, n_161, n_262, n_10, n_177, n_130, n_189, n_103, n_239, n_19, n_87, n_137, n_180, n_104, n_277, n_160, n_98, n_74, n_206, n_276, n_154, n_272, n_7, n_29, n_285, n_195, n_165, n_146, n_45, n_85, n_250, n_237, n_181, n_101, n_62, n_255, n_36, n_47, n_215, n_37, n_34, n_5, n_23, n_8, n_91, n_108, n_116, n_155, n_209, n_217, n_139, n_229, n_230, n_274, n_16, n_13, n_198, n_169, n_193, n_273, n_282, n_252, n_152, n_113, n_241, n_95, n_124, n_156, n_238, n_128, n_120, n_129, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_135, n_42, n_188, n_24, n_78, n_247, n_197, n_201, n_242, n_260, n_6, n_4, n_127, n_170, n_40, n_111, n_157, n_79, n_202, n_210, n_38, n_64, n_142, n_184, n_245, n_265, n_191, n_264, n_281, n_232, n_200, n_46, n_31, n_208, n_211, n_58, n_122, n_187, n_138, n_126, n_275, n_178, n_118, n_258, n_253, n_32, n_0, n_179, n_84, n_131, n_112, n_266, n_55, n_205, n_12, n_86, n_143, n_213, n_235, n_243, n_182, n_263, n_166, n_162, n_186, n_75, n_163, n_226, n_105, n_159, n_174, n_227, n_248, n_268, n_231, n_72, n_136, n_283, n_43, n_76, n_89, n_176, n_68, n_144, n_27, n_53, n_183, n_256, n_67, n_77, n_216, n_20, n_2, n_147, n_199, n_54, n_148, n_123, n_83, n_172, n_28, n_48, n_100, n_212, n_228, n_92, n_11, n_223, n_251, n_25, n_30, n_59, n_236, n_150, n_218, n_168, n_194, n_3, n_287, n_18, n_110, n_261, n_66, n_134, n_222, n_234, n_1, n_164, n_233, n_271, n_82, n_106, n_175, n_15, n_173, n_190, n_286, n_145, n_270, n_246, n_153, n_61, n_259, n_280, n_21, n_99, n_109, n_93, n_132, n_288, n_151, n_51, n_140, n_207, n_257, n_224, n_96, n_269, n_225, n_39, n_279, n_1320);
input n_117;
input n_219;
input n_44;
input n_133;
input n_149;
input n_289;
input n_220;
input n_81;
input n_69;
input n_214;
input n_267;
input n_204;
input n_221;
input n_249;
input n_185;
input n_22;
input n_203;
input n_57;
input n_88;
input n_52;
input n_244;
input n_26;
input n_50;
input n_33;
input n_102;
input n_73;
input n_49;
input n_119;
input n_141;
input n_115;
input n_97;
input n_80;
input n_167;
input n_284;
input n_107;
input n_158;
input n_278;
input n_60;
input n_114;
input n_121;
input n_41;
input n_35;
input n_94;
input n_65;
input n_171;
input n_196;
input n_125;
input n_192;
input n_240;
input n_254;
input n_9;
input n_161;
input n_262;
input n_10;
input n_177;
input n_130;
input n_189;
input n_103;
input n_239;
input n_19;
input n_87;
input n_137;
input n_180;
input n_104;
input n_277;
input n_160;
input n_98;
input n_74;
input n_206;
input n_276;
input n_154;
input n_272;
input n_7;
input n_29;
input n_285;
input n_195;
input n_165;
input n_146;
input n_45;
input n_85;
input n_250;
input n_237;
input n_181;
input n_101;
input n_62;
input n_255;
input n_36;
input n_47;
input n_215;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_108;
input n_116;
input n_155;
input n_209;
input n_217;
input n_139;
input n_229;
input n_230;
input n_274;
input n_16;
input n_13;
input n_198;
input n_169;
input n_193;
input n_273;
input n_282;
input n_252;
input n_152;
input n_113;
input n_241;
input n_95;
input n_124;
input n_156;
input n_238;
input n_128;
input n_120;
input n_129;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_135;
input n_42;
input n_188;
input n_24;
input n_78;
input n_247;
input n_197;
input n_201;
input n_242;
input n_260;
input n_6;
input n_4;
input n_127;
input n_170;
input n_40;
input n_111;
input n_157;
input n_79;
input n_202;
input n_210;
input n_38;
input n_64;
input n_142;
input n_184;
input n_245;
input n_265;
input n_191;
input n_264;
input n_281;
input n_232;
input n_200;
input n_46;
input n_31;
input n_208;
input n_211;
input n_58;
input n_122;
input n_187;
input n_138;
input n_126;
input n_275;
input n_178;
input n_118;
input n_258;
input n_253;
input n_32;
input n_0;
input n_179;
input n_84;
input n_131;
input n_112;
input n_266;
input n_55;
input n_205;
input n_12;
input n_86;
input n_143;
input n_213;
input n_235;
input n_243;
input n_182;
input n_263;
input n_166;
input n_162;
input n_186;
input n_75;
input n_163;
input n_226;
input n_105;
input n_159;
input n_174;
input n_227;
input n_248;
input n_268;
input n_231;
input n_72;
input n_136;
input n_283;
input n_43;
input n_76;
input n_89;
input n_176;
input n_68;
input n_144;
input n_27;
input n_53;
input n_183;
input n_256;
input n_67;
input n_77;
input n_216;
input n_20;
input n_2;
input n_147;
input n_199;
input n_54;
input n_148;
input n_123;
input n_83;
input n_172;
input n_28;
input n_48;
input n_100;
input n_212;
input n_228;
input n_92;
input n_11;
input n_223;
input n_251;
input n_25;
input n_30;
input n_59;
input n_236;
input n_150;
input n_218;
input n_168;
input n_194;
input n_3;
input n_287;
input n_18;
input n_110;
input n_261;
input n_66;
input n_134;
input n_222;
input n_234;
input n_1;
input n_164;
input n_233;
input n_271;
input n_82;
input n_106;
input n_175;
input n_15;
input n_173;
input n_190;
input n_286;
input n_145;
input n_270;
input n_246;
input n_153;
input n_61;
input n_259;
input n_280;
input n_21;
input n_99;
input n_109;
input n_93;
input n_132;
input n_288;
input n_151;
input n_51;
input n_140;
input n_207;
input n_257;
input n_224;
input n_96;
input n_269;
input n_225;
input n_39;
input n_279;
output n_1320;
wire n_1309;
wire n_963;
wire n_1034;
wire n_949;
wire n_1277;
wire n_1312;
wire n_858;
wire n_646;
wire n_829;
wire n_1198;
wire n_667;
wire n_988;
wire n_311;
wire n_655;
wire n_1298;
wire n_903;
wire n_965;
wire n_918;
wire n_770;
wire n_1211;
wire n_878;
wire n_637;
wire n_564;
wire n_779;
wire n_528;
wire n_1128;
wire n_850;
wire n_672;
wire n_627;
wire n_1118;
wire n_1161;
wire n_1030;
wire n_807;
wire n_877;
wire n_545;
wire n_896;
wire n_334;
wire n_588;
wire n_1019;
wire n_940;
wire n_789;
wire n_1197;
wire n_1163;
wire n_387;
wire n_452;
wire n_518;
wire n_298;
wire n_411;
wire n_860;
wire n_1208;
wire n_305;
wire n_1201;
wire n_340;
wire n_373;
wire n_1194;
wire n_922;
wire n_465;
wire n_636;
wire n_914;
wire n_1005;
wire n_1097;
wire n_1125;
wire n_1017;
wire n_324;
wire n_773;
wire n_847;
wire n_668;
wire n_437;
wire n_680;
wire n_642;
wire n_1267;
wire n_830;
wire n_1112;
wire n_517;
wire n_1295;
wire n_1297;
wire n_502;
wire n_543;
wire n_312;
wire n_1159;
wire n_1250;
wire n_1002;
wire n_915;
wire n_367;
wire n_314;
wire n_999;
wire n_769;
wire n_624;
wire n_725;
wire n_1018;
wire n_979;
wire n_319;
wire n_499;
wire n_1033;
wire n_1063;
wire n_1010;
wire n_533;
wire n_490;
wire n_613;
wire n_648;
wire n_304;
wire n_892;
wire n_571;
wire n_610;
wire n_771;
wire n_474;
wire n_402;
wire n_413;
wire n_676;
wire n_950;
wire n_995;
wire n_938;
wire n_331;
wire n_746;
wire n_1307;
wire n_619;
wire n_501;
wire n_299;
wire n_699;
wire n_338;
wire n_551;
wire n_404;
wire n_1061;
wire n_509;
wire n_849;
wire n_864;
wire n_961;
wire n_1140;
wire n_611;
wire n_990;
wire n_800;
wire n_626;
wire n_1209;
wire n_926;
wire n_1274;
wire n_537;
wire n_660;
wire n_839;
wire n_1210;
wire n_1001;
wire n_1129;
wire n_450;
wire n_1099;
wire n_556;
wire n_1214;
wire n_379;
wire n_641;
wire n_966;
wire n_527;
wire n_797;
wire n_666;
wire n_1313;
wire n_954;
wire n_574;
wire n_823;
wire n_706;
wire n_822;
wire n_1181;
wire n_390;
wire n_514;
wire n_486;
wire n_568;
wire n_716;
wire n_899;
wire n_1066;
wire n_1251;
wire n_1199;
wire n_883;
wire n_573;
wire n_1308;
wire n_673;
wire n_1071;
wire n_1079;
wire n_409;
wire n_315;
wire n_295;
wire n_677;
wire n_1242;
wire n_756;
wire n_1240;
wire n_1139;
wire n_577;
wire n_870;
wire n_790;
wire n_761;
wire n_1287;
wire n_472;
wire n_1100;
wire n_419;
wire n_1193;
wire n_1119;
wire n_825;
wire n_477;
wire n_815;
wire n_908;
wire n_429;
wire n_488;
wire n_821;
wire n_745;
wire n_684;
wire n_1281;
wire n_327;
wire n_1102;
wire n_723;
wire n_972;
wire n_997;
wire n_1244;
wire n_1184;
wire n_947;
wire n_620;
wire n_1141;
wire n_1213;
wire n_359;
wire n_1189;
wire n_1316;
wire n_923;
wire n_1205;
wire n_1172;
wire n_741;
wire n_1142;
wire n_1228;
wire n_831;
wire n_859;
wire n_1165;
wire n_1300;
wire n_994;
wire n_930;
wire n_410;
wire n_774;
wire n_1207;
wire n_377;
wire n_510;
wire n_1075;
wire n_1282;
wire n_493;
wire n_855;
wire n_722;
wire n_1083;
wire n_690;
wire n_1164;
wire n_451;
wire n_487;
wire n_748;
wire n_824;
wire n_793;
wire n_753;
wire n_355;
wire n_382;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_1226;
wire n_1233;
wire n_1067;
wire n_866;
wire n_1108;
wire n_350;
wire n_433;
wire n_1311;
wire n_483;
wire n_395;
wire n_992;
wire n_361;
wire n_1077;
wire n_838;
wire n_705;
wire n_964;
wire n_590;
wire n_407;
wire n_1229;
wire n_792;
wire n_925;
wire n_1289;
wire n_957;
wire n_808;
wire n_431;
wire n_484;
wire n_862;
wire n_852;
wire n_1306;
wire n_958;
wire n_468;
wire n_917;
wire n_523;
wire n_920;
wire n_1202;
wire n_911;
wire n_980;
wire n_817;
wire n_1056;
wire n_856;
wire n_661;
wire n_890;
wire n_787;
wire n_1015;
wire n_548;
wire n_1048;
wire n_973;
wire n_587;
wire n_476;
wire n_434;
wire n_489;
wire n_752;
wire n_1098;
wire n_1012;
wire n_461;
wire n_857;
wire n_1090;
wire n_786;
wire n_1121;
wire n_576;
wire n_1179;
wire n_796;
wire n_1216;
wire n_927;
wire n_840;
wire n_846;
wire n_968;
wire n_512;
wire n_586;
wire n_1246;
wire n_1276;
wire n_560;
wire n_697;
wire n_780;
wire n_447;
wire n_897;
wire n_1188;
wire n_580;
wire n_1009;
wire n_921;
wire n_854;
wire n_1011;
wire n_1155;
wire n_511;
wire n_467;
wire n_692;
wire n_644;
wire n_1116;
wire n_818;
wire n_738;
wire n_1225;
wire n_575;
wire n_711;
wire n_977;
wire n_884;
wire n_767;
wire n_293;
wire n_393;
wire n_550;
wire n_826;
wire n_399;
wire n_1235;
wire n_1171;
wire n_294;
wire n_459;
wire n_907;
wire n_310;
wire n_1062;
wire n_708;
wire n_1271;
wire n_307;
wire n_634;
wire n_696;
wire n_1203;
wire n_1013;
wire n_1000;
wire n_939;
wire n_953;
wire n_391;
wire n_478;
wire n_482;
wire n_394;
wire n_442;
wire n_485;
wire n_1248;
wire n_519;
wire n_329;
wire n_1020;
wire n_1106;
wire n_635;
wire n_731;
wire n_986;
wire n_507;
wire n_605;
wire n_704;
wire n_633;
wire n_873;
wire n_751;
wire n_1147;
wire n_466;
wire n_900;
wire n_952;
wire n_685;
wire n_308;
wire n_565;
wire n_1035;
wire n_475;
wire n_578;
wire n_542;
wire n_430;
wire n_943;
wire n_557;
wire n_842;
wire n_1269;
wire n_439;
wire n_614;
wire n_1107;
wire n_446;
wire n_423;
wire n_342;
wire n_799;
wire n_1050;
wire n_643;
wire n_874;
wire n_1049;
wire n_454;
wire n_687;
wire n_970;
wire n_984;
wire n_720;
wire n_806;
wire n_1157;
wire n_539;
wire n_1153;
wire n_317;
wire n_816;
wire n_522;
wire n_898;
wire n_1135;
wire n_669;
wire n_541;
wire n_363;
wire n_733;
wire n_894;
wire n_376;
wire n_744;
wire n_520;
wire n_681;
wire n_942;
wire n_1029;
wire n_508;
wire n_721;
wire n_1060;
wire n_438;
wire n_640;
wire n_1037;
wire n_686;
wire n_944;
wire n_1110;
wire n_498;
wire n_1069;
wire n_1123;
wire n_811;
wire n_530;
wire n_737;
wire n_1266;
wire n_795;
wire n_1232;
wire n_449;
wire n_734;
wire n_919;
wire n_763;
wire n_1174;
wire n_657;
wire n_583;
wire n_841;
wire n_582;
wire n_836;
wire n_561;
wire n_1096;
wire n_594;
wire n_531;
wire n_1136;
wire n_306;
wire n_1007;
wire n_1117;
wire n_424;
wire n_714;
wire n_932;
wire n_837;
wire n_1315;
wire n_867;
wire n_1070;
wire n_1270;
wire n_675;
wire n_504;
wire n_581;
wire n_698;
wire n_555;
wire n_834;
wire n_901;
wire n_727;
wire n_1038;
wire n_1162;
wire n_1103;
wire n_785;
wire n_375;
wire n_688;
wire n_323;
wire n_347;
wire n_515;
wire n_1290;
wire n_1234;
wire n_592;
wire n_1045;
wire n_1115;
wire n_521;
wire n_625;
wire n_585;
wire n_1190;
wire n_1237;
wire n_713;
wire n_457;
wire n_736;
wire n_606;
wire n_332;
wire n_1292;
wire n_421;
wire n_1148;
wire n_739;
wire n_1166;
wire n_987;
wire n_1086;
wire n_406;
wire n_1236;
wire n_791;
wire n_707;
wire n_603;
wire n_1261;
wire n_885;
wire n_500;
wire n_607;
wire n_496;
wire n_801;
wire n_1059;
wire n_309;
wire n_701;
wire n_612;
wire n_1032;
wire n_1284;
wire n_336;
wire n_464;
wire n_1243;
wire n_1196;
wire n_814;
wire n_985;
wire n_1191;
wire n_971;
wire n_904;
wire n_1301;
wire n_532;
wire n_400;
wire n_386;
wire n_432;
wire n_659;
wire n_316;
wire n_1185;
wire n_389;
wire n_436;
wire n_1217;
wire n_715;
wire n_330;
wire n_1087;
wire n_662;
wire n_617;
wire n_598;
wire n_732;
wire n_724;
wire n_599;
wire n_301;
wire n_609;
wire n_909;
wire n_1273;
wire n_366;
wire n_1319;
wire n_596;
wire n_1215;
wire n_951;
wire n_321;
wire n_1024;
wire n_1016;
wire n_652;
wire n_333;
wire n_638;
wire n_563;
wire n_479;
wire n_623;
wire n_1222;
wire n_593;
wire n_872;
wire n_809;
wire n_1101;
wire n_1072;
wire n_865;
wire n_1064;
wire n_1254;
wire n_764;
wire n_426;
wire n_969;
wire n_417;
wire n_1253;
wire n_632;
wire n_1182;
wire n_828;
wire n_1138;
wire n_506;
wire n_381;
wire n_1255;
wire n_313;
wire n_322;
wire n_1299;
wire n_427;
wire n_703;
wire n_415;
wire n_1272;
wire n_928;
wire n_352;
wire n_882;
wire n_871;
wire n_803;
wire n_729;
wire n_805;
wire n_693;
wire n_1036;
wire n_1145;
wire n_651;
wire n_1303;
wire n_747;
wire n_905;
wire n_525;
wire n_876;
wire n_886;
wire n_959;
wire n_719;
wire n_1206;
wire n_1257;
wire n_710;
wire n_1178;
wire n_546;
wire n_412;
wire n_664;
wire n_1249;
wire n_788;
wire n_403;
wire n_516;
wire n_549;
wire n_832;
wire n_996;
wire n_420;
wire n_1089;
wire n_1058;
wire n_388;
wire n_1082;
wire n_1052;
wire n_1055;
wire n_974;
wire n_591;
wire n_933;
wire n_1252;
wire n_416;
wire n_536;
wire n_1256;
wire n_1259;
wire n_1318;
wire n_956;
wire n_989;
wire n_754;
wire n_775;
wire n_616;
wire n_1227;
wire n_365;
wire n_495;
wire n_364;
wire n_566;
wire n_1144;
wire n_344;
wire n_503;
wire n_1279;
wire n_1152;
wire n_1068;
wire n_1149;
wire n_615;
wire n_1170;
wire n_804;
wire n_570;
wire n_1133;
wire n_1317;
wire n_440;
wire n_422;
wire n_679;
wire n_1131;
wire n_597;
wire n_1039;
wire n_835;
wire n_778;
wire n_1156;
wire n_1288;
wire n_300;
wire n_1042;
wire n_584;
wire n_1130;
wire n_912;
wire n_1043;
wire n_1283;
wire n_346;
wire n_397;
wire n_1008;
wire n_1109;
wire n_1026;
wire n_1027;
wire n_1040;
wire n_569;
wire n_946;
wire n_960;
wire n_1168;
wire n_343;
wire n_458;
wire n_1084;
wire n_618;
wire n_341;
wire n_470;
wire n_1085;
wire n_1073;
wire n_868;
wire n_473;
wire n_991;
wire n_843;
wire n_1263;
wire n_538;
wire n_492;
wire n_1150;
wire n_368;
wire n_650;
wire n_469;
wire n_1187;
wire n_742;
wire n_913;
wire n_845;
wire n_891;
wire n_1134;
wire n_494;
wire n_372;
wire n_631;
wire n_934;
wire n_425;
wire n_562;
wire n_1192;
wire n_983;
wire n_781;
wire n_709;
wire n_1105;
wire n_408;
wire n_290;
wire n_385;
wire n_1127;
wire n_1173;
wire n_663;
wire n_513;
wire n_1092;
wire n_1124;
wire n_1278;
wire n_998;
wire n_604;
wire n_1260;
wire n_755;
wire n_848;
wire n_1031;
wire n_1293;
wire n_1280;
wire n_292;
wire n_1158;
wire n_328;
wire n_743;
wire n_757;
wire n_750;
wire n_448;
wire n_645;
wire n_348;
wire n_1022;
wire n_802;
wire n_353;
wire n_993;
wire n_1122;
wire n_1224;
wire n_383;
wire n_762;
wire n_981;
wire n_1095;
wire n_758;
wire n_544;
wire n_1175;
wire n_853;
wire n_296;
wire n_765;
wire n_1177;
wire n_1310;
wire n_462;
wire n_783;
wire n_1074;
wire n_463;
wire n_1003;
wire n_678;
wire n_1200;
wire n_384;
wire n_978;
wire n_547;
wire n_1247;
wire n_628;
wire n_812;
wire n_777;
wire n_351;
wire n_401;
wire n_345;
wire n_360;
wire n_481;
wire n_443;
wire n_694;
wire n_1262;
wire n_1078;
wire n_702;
wire n_572;
wire n_1094;
wire n_1204;
wire n_392;
wire n_1169;
wire n_975;
wire n_303;
wire n_326;
wire n_1081;
wire n_671;
wire n_540;
wire n_937;
wire n_1093;
wire n_955;
wire n_1275;
wire n_945;
wire n_554;
wire n_726;
wire n_712;
wire n_608;
wire n_567;
wire n_888;
wire n_455;
wire n_529;
wire n_1025;
wire n_1132;
wire n_630;
wire n_1180;
wire n_647;
wire n_844;
wire n_1160;
wire n_1245;
wire n_1195;
wire n_1241;
wire n_1302;
wire n_895;
wire n_798;
wire n_318;
wire n_887;
wire n_471;
wire n_1014;
wire n_665;
wire n_1154;
wire n_863;
wire n_1265;
wire n_730;
wire n_1212;
wire n_735;
wire n_1091;
wire n_784;
wire n_354;
wire n_1220;
wire n_893;
wire n_1028;
wire n_910;
wire n_935;
wire n_1046;
wire n_1183;
wire n_460;
wire n_813;
wire n_1076;
wire n_369;
wire n_1186;
wire n_1167;
wire n_674;
wire n_810;
wire n_982;
wire n_889;
wire n_689;
wire n_902;
wire n_1113;
wire n_1264;
wire n_760;
wire n_941;
wire n_302;
wire n_362;
wire n_931;
wire n_827;
wire n_1218;
wire n_1041;
wire n_1080;
wire n_1126;
wire n_1151;
wire n_936;
wire n_579;
wire n_776;
wire n_879;
wire n_1065;
wire n_622;
wire n_601;
wire n_1176;
wire n_649;
wire n_526;
wire n_1047;
wire n_320;
wire n_768;
wire n_869;
wire n_880;
wire n_621;
wire n_370;
wire n_589;
wire n_505;
wire n_682;
wire n_906;
wire n_357;
wire n_653;
wire n_881;
wire n_374;
wire n_718;
wire n_1238;
wire n_1114;
wire n_1286;
wire n_948;
wire n_1304;
wire n_1314;
wire n_717;
wire n_861;
wire n_654;
wire n_1221;
wire n_428;
wire n_794;
wire n_1268;
wire n_639;
wire n_1305;
wire n_552;
wire n_1023;
wire n_1057;
wire n_435;
wire n_1294;
wire n_1051;
wire n_1088;
wire n_851;
wire n_396;
wire n_398;
wire n_445;
wire n_656;
wire n_1230;
wire n_553;
wire n_325;
wire n_349;
wire n_1021;
wire n_749;
wire n_535;
wire n_1006;
wire n_1054;
wire n_1231;
wire n_358;
wire n_456;
wire n_962;
wire n_782;
wire n_524;
wire n_1044;
wire n_875;
wire n_497;
wire n_728;
wire n_339;
wire n_1239;
wire n_924;
wire n_378;
wire n_441;
wire n_1285;
wire n_335;
wire n_700;
wire n_534;
wire n_1296;
wire n_766;
wire n_602;
wire n_1143;
wire n_629;
wire n_297;
wire n_1053;
wire n_1223;
wire n_967;
wire n_1258;
wire n_291;
wire n_418;
wire n_380;
wire n_356;
wire n_600;
wire n_371;
wire n_820;
wire n_558;
wire n_670;
wire n_1004;
wire n_683;
wire n_929;
wire n_1111;
wire n_976;
wire n_695;
wire n_1104;
wire n_1120;
wire n_1219;
wire n_595;
wire n_759;
wire n_559;
wire n_480;
wire n_453;
wire n_833;
wire n_1146;
wire n_414;
wire n_1137;
wire n_916;
wire n_740;
wire n_772;
wire n_819;
wire n_405;
wire n_491;
wire n_1291;
INVx1_ASAP7_75t_L g290 ( .A(n_180), .Y(n_290) );
INVx1_ASAP7_75t_L g291 ( .A(n_35), .Y(n_291) );
CKINVDCx16_ASAP7_75t_R g292 ( .A(n_259), .Y(n_292) );
INVx1_ASAP7_75t_SL g293 ( .A(n_146), .Y(n_293) );
INVx1_ASAP7_75t_L g294 ( .A(n_64), .Y(n_294) );
INVx2_ASAP7_75t_L g295 ( .A(n_2), .Y(n_295) );
INVx2_ASAP7_75t_L g296 ( .A(n_34), .Y(n_296) );
INVx1_ASAP7_75t_L g297 ( .A(n_123), .Y(n_297) );
INVx1_ASAP7_75t_L g298 ( .A(n_215), .Y(n_298) );
CKINVDCx16_ASAP7_75t_R g299 ( .A(n_245), .Y(n_299) );
CKINVDCx5p33_ASAP7_75t_R g300 ( .A(n_257), .Y(n_300) );
BUFx3_ASAP7_75t_L g301 ( .A(n_116), .Y(n_301) );
CKINVDCx5p33_ASAP7_75t_R g302 ( .A(n_254), .Y(n_302) );
INVx1_ASAP7_75t_SL g303 ( .A(n_225), .Y(n_303) );
BUFx6f_ASAP7_75t_L g304 ( .A(n_273), .Y(n_304) );
INVxp67_ASAP7_75t_SL g305 ( .A(n_287), .Y(n_305) );
INVx2_ASAP7_75t_SL g306 ( .A(n_227), .Y(n_306) );
INVx1_ASAP7_75t_L g307 ( .A(n_241), .Y(n_307) );
INVx1_ASAP7_75t_L g308 ( .A(n_30), .Y(n_308) );
INVx1_ASAP7_75t_L g309 ( .A(n_87), .Y(n_309) );
BUFx3_ASAP7_75t_L g310 ( .A(n_31), .Y(n_310) );
BUFx6f_ASAP7_75t_L g311 ( .A(n_150), .Y(n_311) );
INVx1_ASAP7_75t_L g312 ( .A(n_94), .Y(n_312) );
CKINVDCx16_ASAP7_75t_R g313 ( .A(n_189), .Y(n_313) );
INVxp67_ASAP7_75t_L g314 ( .A(n_49), .Y(n_314) );
INVx1_ASAP7_75t_L g315 ( .A(n_253), .Y(n_315) );
INVx1_ASAP7_75t_L g316 ( .A(n_275), .Y(n_316) );
INVx1_ASAP7_75t_L g317 ( .A(n_156), .Y(n_317) );
CKINVDCx20_ASAP7_75t_R g318 ( .A(n_73), .Y(n_318) );
INVx1_ASAP7_75t_L g319 ( .A(n_31), .Y(n_319) );
INVx1_ASAP7_75t_L g320 ( .A(n_139), .Y(n_320) );
INVx1_ASAP7_75t_L g321 ( .A(n_53), .Y(n_321) );
INVx1_ASAP7_75t_L g322 ( .A(n_127), .Y(n_322) );
INVx1_ASAP7_75t_L g323 ( .A(n_278), .Y(n_323) );
INVx1_ASAP7_75t_SL g324 ( .A(n_272), .Y(n_324) );
INVx1_ASAP7_75t_L g325 ( .A(n_104), .Y(n_325) );
CKINVDCx20_ASAP7_75t_R g326 ( .A(n_221), .Y(n_326) );
INVx1_ASAP7_75t_L g327 ( .A(n_12), .Y(n_327) );
INVx1_ASAP7_75t_L g328 ( .A(n_208), .Y(n_328) );
INVx1_ASAP7_75t_L g329 ( .A(n_171), .Y(n_329) );
CKINVDCx16_ASAP7_75t_R g330 ( .A(n_35), .Y(n_330) );
INVx2_ASAP7_75t_L g331 ( .A(n_22), .Y(n_331) );
BUFx6f_ASAP7_75t_L g332 ( .A(n_205), .Y(n_332) );
INVx1_ASAP7_75t_L g333 ( .A(n_223), .Y(n_333) );
INVx1_ASAP7_75t_L g334 ( .A(n_95), .Y(n_334) );
INVxp67_ASAP7_75t_SL g335 ( .A(n_233), .Y(n_335) );
INVx1_ASAP7_75t_SL g336 ( .A(n_16), .Y(n_336) );
BUFx3_ASAP7_75t_L g337 ( .A(n_144), .Y(n_337) );
INVx1_ASAP7_75t_L g338 ( .A(n_269), .Y(n_338) );
INVx1_ASAP7_75t_L g339 ( .A(n_136), .Y(n_339) );
INVx1_ASAP7_75t_L g340 ( .A(n_44), .Y(n_340) );
INVxp67_ASAP7_75t_L g341 ( .A(n_102), .Y(n_341) );
INVx1_ASAP7_75t_L g342 ( .A(n_41), .Y(n_342) );
INVx1_ASAP7_75t_L g343 ( .A(n_264), .Y(n_343) );
INVx1_ASAP7_75t_L g344 ( .A(n_2), .Y(n_344) );
INVx1_ASAP7_75t_L g345 ( .A(n_220), .Y(n_345) );
INVx1_ASAP7_75t_L g346 ( .A(n_159), .Y(n_346) );
CKINVDCx5p33_ASAP7_75t_R g347 ( .A(n_113), .Y(n_347) );
INVx1_ASAP7_75t_L g348 ( .A(n_61), .Y(n_348) );
INVx1_ASAP7_75t_L g349 ( .A(n_281), .Y(n_349) );
INVx1_ASAP7_75t_L g350 ( .A(n_77), .Y(n_350) );
HB1xp67_ASAP7_75t_L g351 ( .A(n_243), .Y(n_351) );
INVx1_ASAP7_75t_L g352 ( .A(n_54), .Y(n_352) );
INVx1_ASAP7_75t_L g353 ( .A(n_234), .Y(n_353) );
INVx2_ASAP7_75t_L g354 ( .A(n_110), .Y(n_354) );
INVx1_ASAP7_75t_L g355 ( .A(n_232), .Y(n_355) );
INVx1_ASAP7_75t_L g356 ( .A(n_174), .Y(n_356) );
INVx1_ASAP7_75t_L g357 ( .A(n_247), .Y(n_357) );
INVx1_ASAP7_75t_L g358 ( .A(n_172), .Y(n_358) );
CKINVDCx16_ASAP7_75t_R g359 ( .A(n_41), .Y(n_359) );
INVx1_ASAP7_75t_L g360 ( .A(n_165), .Y(n_360) );
INVx1_ASAP7_75t_L g361 ( .A(n_140), .Y(n_361) );
CKINVDCx20_ASAP7_75t_R g362 ( .A(n_149), .Y(n_362) );
BUFx6f_ASAP7_75t_L g363 ( .A(n_251), .Y(n_363) );
INVx1_ASAP7_75t_L g364 ( .A(n_203), .Y(n_364) );
INVx1_ASAP7_75t_L g365 ( .A(n_106), .Y(n_365) );
BUFx3_ASAP7_75t_L g366 ( .A(n_280), .Y(n_366) );
INVx1_ASAP7_75t_L g367 ( .A(n_24), .Y(n_367) );
INVx1_ASAP7_75t_L g368 ( .A(n_228), .Y(n_368) );
INVx1_ASAP7_75t_L g369 ( .A(n_256), .Y(n_369) );
CKINVDCx5p33_ASAP7_75t_R g370 ( .A(n_38), .Y(n_370) );
CKINVDCx5p33_ASAP7_75t_R g371 ( .A(n_242), .Y(n_371) );
CKINVDCx16_ASAP7_75t_R g372 ( .A(n_126), .Y(n_372) );
INVx1_ASAP7_75t_L g373 ( .A(n_219), .Y(n_373) );
INVxp33_ASAP7_75t_SL g374 ( .A(n_145), .Y(n_374) );
BUFx2_ASAP7_75t_L g375 ( .A(n_10), .Y(n_375) );
INVx1_ASAP7_75t_L g376 ( .A(n_96), .Y(n_376) );
CKINVDCx20_ASAP7_75t_R g377 ( .A(n_270), .Y(n_377) );
INVx2_ASAP7_75t_L g378 ( .A(n_276), .Y(n_378) );
CKINVDCx16_ASAP7_75t_R g379 ( .A(n_206), .Y(n_379) );
INVx1_ASAP7_75t_L g380 ( .A(n_83), .Y(n_380) );
INVx2_ASAP7_75t_L g381 ( .A(n_130), .Y(n_381) );
CKINVDCx5p33_ASAP7_75t_R g382 ( .A(n_138), .Y(n_382) );
NOR2xp67_ASAP7_75t_L g383 ( .A(n_10), .B(n_119), .Y(n_383) );
INVx1_ASAP7_75t_L g384 ( .A(n_177), .Y(n_384) );
INVx2_ASAP7_75t_SL g385 ( .A(n_282), .Y(n_385) );
NOR2xp33_ASAP7_75t_L g386 ( .A(n_34), .B(n_4), .Y(n_386) );
INVxp33_ASAP7_75t_L g387 ( .A(n_279), .Y(n_387) );
INVxp67_ASAP7_75t_SL g388 ( .A(n_5), .Y(n_388) );
INVx2_ASAP7_75t_L g389 ( .A(n_133), .Y(n_389) );
INVxp67_ASAP7_75t_L g390 ( .A(n_137), .Y(n_390) );
CKINVDCx5p33_ASAP7_75t_R g391 ( .A(n_54), .Y(n_391) );
CKINVDCx20_ASAP7_75t_R g392 ( .A(n_128), .Y(n_392) );
CKINVDCx16_ASAP7_75t_R g393 ( .A(n_129), .Y(n_393) );
INVx1_ASAP7_75t_L g394 ( .A(n_46), .Y(n_394) );
INVxp67_ASAP7_75t_SL g395 ( .A(n_131), .Y(n_395) );
INVxp33_ASAP7_75t_SL g396 ( .A(n_29), .Y(n_396) );
BUFx6f_ASAP7_75t_L g397 ( .A(n_100), .Y(n_397) );
CKINVDCx5p33_ASAP7_75t_R g398 ( .A(n_196), .Y(n_398) );
INVx1_ASAP7_75t_L g399 ( .A(n_236), .Y(n_399) );
INVx2_ASAP7_75t_L g400 ( .A(n_202), .Y(n_400) );
CKINVDCx5p33_ASAP7_75t_R g401 ( .A(n_86), .Y(n_401) );
INVx2_ASAP7_75t_L g402 ( .A(n_188), .Y(n_402) );
INVx1_ASAP7_75t_L g403 ( .A(n_224), .Y(n_403) );
BUFx3_ASAP7_75t_L g404 ( .A(n_118), .Y(n_404) );
NOR2xp67_ASAP7_75t_L g405 ( .A(n_151), .B(n_190), .Y(n_405) );
CKINVDCx16_ASAP7_75t_R g406 ( .A(n_99), .Y(n_406) );
CKINVDCx5p33_ASAP7_75t_R g407 ( .A(n_182), .Y(n_407) );
INVxp67_ASAP7_75t_SL g408 ( .A(n_155), .Y(n_408) );
CKINVDCx20_ASAP7_75t_R g409 ( .A(n_218), .Y(n_409) );
INVx1_ASAP7_75t_L g410 ( .A(n_111), .Y(n_410) );
INVxp33_ASAP7_75t_L g411 ( .A(n_36), .Y(n_411) );
INVx1_ASAP7_75t_L g412 ( .A(n_213), .Y(n_412) );
INVxp33_ASAP7_75t_L g413 ( .A(n_11), .Y(n_413) );
INVxp67_ASAP7_75t_SL g414 ( .A(n_18), .Y(n_414) );
CKINVDCx16_ASAP7_75t_R g415 ( .A(n_101), .Y(n_415) );
INVx1_ASAP7_75t_L g416 ( .A(n_162), .Y(n_416) );
CKINVDCx20_ASAP7_75t_R g417 ( .A(n_65), .Y(n_417) );
INVx1_ASAP7_75t_L g418 ( .A(n_37), .Y(n_418) );
CKINVDCx16_ASAP7_75t_R g419 ( .A(n_0), .Y(n_419) );
INVx2_ASAP7_75t_L g420 ( .A(n_50), .Y(n_420) );
INVx1_ASAP7_75t_L g421 ( .A(n_199), .Y(n_421) );
CKINVDCx5p33_ASAP7_75t_R g422 ( .A(n_37), .Y(n_422) );
INVxp33_ASAP7_75t_SL g423 ( .A(n_214), .Y(n_423) );
INVxp67_ASAP7_75t_L g424 ( .A(n_57), .Y(n_424) );
INVx2_ASAP7_75t_L g425 ( .A(n_147), .Y(n_425) );
INVx1_ASAP7_75t_L g426 ( .A(n_56), .Y(n_426) );
CKINVDCx5p33_ASAP7_75t_R g427 ( .A(n_18), .Y(n_427) );
INVx1_ASAP7_75t_L g428 ( .A(n_173), .Y(n_428) );
INVx1_ASAP7_75t_L g429 ( .A(n_181), .Y(n_429) );
INVx1_ASAP7_75t_L g430 ( .A(n_120), .Y(n_430) );
INVx1_ASAP7_75t_L g431 ( .A(n_261), .Y(n_431) );
BUFx3_ASAP7_75t_L g432 ( .A(n_56), .Y(n_432) );
INVxp67_ASAP7_75t_SL g433 ( .A(n_92), .Y(n_433) );
INVxp67_ASAP7_75t_SL g434 ( .A(n_24), .Y(n_434) );
INVxp33_ASAP7_75t_L g435 ( .A(n_135), .Y(n_435) );
INVxp67_ASAP7_75t_SL g436 ( .A(n_112), .Y(n_436) );
INVx2_ASAP7_75t_L g437 ( .A(n_132), .Y(n_437) );
INVxp67_ASAP7_75t_SL g438 ( .A(n_271), .Y(n_438) );
INVx1_ASAP7_75t_L g439 ( .A(n_32), .Y(n_439) );
INVx1_ASAP7_75t_L g440 ( .A(n_240), .Y(n_440) );
CKINVDCx5p33_ASAP7_75t_R g441 ( .A(n_14), .Y(n_441) );
INVx1_ASAP7_75t_L g442 ( .A(n_134), .Y(n_442) );
INVx1_ASAP7_75t_L g443 ( .A(n_117), .Y(n_443) );
CKINVDCx5p33_ASAP7_75t_R g444 ( .A(n_197), .Y(n_444) );
CKINVDCx5p33_ASAP7_75t_R g445 ( .A(n_216), .Y(n_445) );
NOR2xp33_ASAP7_75t_L g446 ( .A(n_93), .B(n_109), .Y(n_446) );
INVx1_ASAP7_75t_L g447 ( .A(n_66), .Y(n_447) );
INVx2_ASAP7_75t_L g448 ( .A(n_82), .Y(n_448) );
INVx2_ASAP7_75t_L g449 ( .A(n_304), .Y(n_449) );
INVx1_ASAP7_75t_L g450 ( .A(n_295), .Y(n_450) );
AND2x2_ASAP7_75t_L g451 ( .A(n_411), .B(n_0), .Y(n_451) );
HB1xp67_ASAP7_75t_L g452 ( .A(n_411), .Y(n_452) );
INVx2_ASAP7_75t_L g453 ( .A(n_304), .Y(n_453) );
INVx1_ASAP7_75t_L g454 ( .A(n_295), .Y(n_454) );
CKINVDCx5p33_ASAP7_75t_R g455 ( .A(n_292), .Y(n_455) );
INVx6_ASAP7_75t_L g456 ( .A(n_301), .Y(n_456) );
HB1xp67_ASAP7_75t_L g457 ( .A(n_413), .Y(n_457) );
INVx1_ASAP7_75t_L g458 ( .A(n_296), .Y(n_458) );
INVx3_ASAP7_75t_L g459 ( .A(n_310), .Y(n_459) );
AND2x2_ASAP7_75t_L g460 ( .A(n_413), .B(n_1), .Y(n_460) );
INVx1_ASAP7_75t_L g461 ( .A(n_296), .Y(n_461) );
BUFx3_ASAP7_75t_L g462 ( .A(n_301), .Y(n_462) );
OAI22xp5_ASAP7_75t_L g463 ( .A1(n_330), .A2(n_4), .B1(n_1), .B2(n_3), .Y(n_463) );
NAND2xp5_ASAP7_75t_L g464 ( .A(n_306), .B(n_3), .Y(n_464) );
BUFx6f_ASAP7_75t_L g465 ( .A(n_304), .Y(n_465) );
AND2x4_ASAP7_75t_L g466 ( .A(n_310), .B(n_5), .Y(n_466) );
NAND2xp5_ASAP7_75t_L g467 ( .A(n_385), .B(n_6), .Y(n_467) );
AND2x2_ASAP7_75t_L g468 ( .A(n_387), .B(n_6), .Y(n_468) );
INVx1_ASAP7_75t_L g469 ( .A(n_331), .Y(n_469) );
CKINVDCx5p33_ASAP7_75t_R g470 ( .A(n_299), .Y(n_470) );
AND3x2_ASAP7_75t_L g471 ( .A(n_375), .B(n_7), .C(n_8), .Y(n_471) );
BUFx6f_ASAP7_75t_L g472 ( .A(n_304), .Y(n_472) );
CKINVDCx5p33_ASAP7_75t_R g473 ( .A(n_313), .Y(n_473) );
INVx1_ASAP7_75t_L g474 ( .A(n_331), .Y(n_474) );
CKINVDCx16_ASAP7_75t_R g475 ( .A(n_372), .Y(n_475) );
NAND2xp5_ASAP7_75t_L g476 ( .A(n_351), .B(n_7), .Y(n_476) );
NAND2xp5_ASAP7_75t_L g477 ( .A(n_291), .B(n_8), .Y(n_477) );
NAND2xp5_ASAP7_75t_L g478 ( .A(n_294), .B(n_9), .Y(n_478) );
INVxp67_ASAP7_75t_L g479 ( .A(n_432), .Y(n_479) );
INVx2_ASAP7_75t_L g480 ( .A(n_311), .Y(n_480) );
INVx1_ASAP7_75t_L g481 ( .A(n_420), .Y(n_481) );
AOI22xp5_ASAP7_75t_L g482 ( .A1(n_396), .A2(n_9), .B1(n_11), .B2(n_12), .Y(n_482) );
AND2x2_ASAP7_75t_L g483 ( .A(n_387), .B(n_435), .Y(n_483) );
INVx2_ASAP7_75t_L g484 ( .A(n_311), .Y(n_484) );
NAND2xp5_ASAP7_75t_SL g485 ( .A(n_311), .B(n_13), .Y(n_485) );
INVx2_ASAP7_75t_L g486 ( .A(n_465), .Y(n_486) );
AND2x6_ASAP7_75t_L g487 ( .A(n_466), .B(n_337), .Y(n_487) );
INVx1_ASAP7_75t_L g488 ( .A(n_459), .Y(n_488) );
CKINVDCx5p33_ASAP7_75t_R g489 ( .A(n_475), .Y(n_489) );
OR2x2_ASAP7_75t_L g490 ( .A(n_452), .B(n_359), .Y(n_490) );
INVx4_ASAP7_75t_L g491 ( .A(n_466), .Y(n_491) );
INVx2_ASAP7_75t_SL g492 ( .A(n_483), .Y(n_492) );
BUFx3_ASAP7_75t_L g493 ( .A(n_456), .Y(n_493) );
NAND2xp5_ASAP7_75t_L g494 ( .A(n_483), .B(n_435), .Y(n_494) );
INVx1_ASAP7_75t_L g495 ( .A(n_459), .Y(n_495) );
BUFx3_ASAP7_75t_L g496 ( .A(n_456), .Y(n_496) );
INVx1_ASAP7_75t_L g497 ( .A(n_459), .Y(n_497) );
NAND2xp5_ASAP7_75t_L g498 ( .A(n_452), .B(n_379), .Y(n_498) );
NOR2xp33_ASAP7_75t_L g499 ( .A(n_457), .B(n_341), .Y(n_499) );
INVx1_ASAP7_75t_L g500 ( .A(n_459), .Y(n_500) );
INVx3_ASAP7_75t_L g501 ( .A(n_466), .Y(n_501) );
INVx1_ASAP7_75t_L g502 ( .A(n_466), .Y(n_502) );
INVx1_ASAP7_75t_L g503 ( .A(n_449), .Y(n_503) );
NOR2xp33_ASAP7_75t_L g504 ( .A(n_457), .B(n_390), .Y(n_504) );
AND2x2_ASAP7_75t_L g505 ( .A(n_468), .B(n_393), .Y(n_505) );
BUFx3_ASAP7_75t_L g506 ( .A(n_456), .Y(n_506) );
INVx1_ASAP7_75t_L g507 ( .A(n_449), .Y(n_507) );
AND2x4_ASAP7_75t_L g508 ( .A(n_479), .B(n_432), .Y(n_508) );
INVx1_ASAP7_75t_L g509 ( .A(n_449), .Y(n_509) );
INVx1_ASAP7_75t_L g510 ( .A(n_453), .Y(n_510) );
INVx1_ASAP7_75t_L g511 ( .A(n_453), .Y(n_511) );
OAI22xp33_ASAP7_75t_L g512 ( .A1(n_475), .A2(n_419), .B1(n_370), .B2(n_391), .Y(n_512) );
NAND2xp5_ASAP7_75t_L g513 ( .A(n_479), .B(n_406), .Y(n_513) );
NAND2xp5_ASAP7_75t_SL g514 ( .A(n_455), .B(n_415), .Y(n_514) );
AND2x2_ASAP7_75t_L g515 ( .A(n_468), .B(n_420), .Y(n_515) );
OR2x2_ASAP7_75t_L g516 ( .A(n_451), .B(n_370), .Y(n_516) );
AND2x4_ASAP7_75t_L g517 ( .A(n_451), .B(n_308), .Y(n_517) );
BUFx3_ASAP7_75t_L g518 ( .A(n_456), .Y(n_518) );
NOR2xp33_ASAP7_75t_L g519 ( .A(n_470), .B(n_374), .Y(n_519) );
INVx4_ASAP7_75t_L g520 ( .A(n_456), .Y(n_520) );
NAND2xp5_ASAP7_75t_L g521 ( .A(n_462), .B(n_391), .Y(n_521) );
CKINVDCx5p33_ASAP7_75t_R g522 ( .A(n_473), .Y(n_522) );
BUFx2_ASAP7_75t_L g523 ( .A(n_460), .Y(n_523) );
AOI22xp5_ASAP7_75t_L g524 ( .A1(n_460), .A2(n_396), .B1(n_326), .B2(n_377), .Y(n_524) );
INVx2_ASAP7_75t_L g525 ( .A(n_465), .Y(n_525) );
NOR3xp33_ASAP7_75t_L g526 ( .A(n_463), .B(n_424), .C(n_314), .Y(n_526) );
NAND2xp5_ASAP7_75t_L g527 ( .A(n_462), .B(n_422), .Y(n_527) );
NAND2xp5_ASAP7_75t_L g528 ( .A(n_462), .B(n_422), .Y(n_528) );
INVx2_ASAP7_75t_L g529 ( .A(n_465), .Y(n_529) );
BUFx3_ASAP7_75t_L g530 ( .A(n_450), .Y(n_530) );
INVx3_ASAP7_75t_L g531 ( .A(n_472), .Y(n_531) );
NAND2xp5_ASAP7_75t_L g532 ( .A(n_450), .B(n_441), .Y(n_532) );
INVx2_ASAP7_75t_L g533 ( .A(n_465), .Y(n_533) );
INVx6_ASAP7_75t_L g534 ( .A(n_472), .Y(n_534) );
BUFx3_ASAP7_75t_L g535 ( .A(n_454), .Y(n_535) );
NAND2xp5_ASAP7_75t_SL g536 ( .A(n_491), .B(n_476), .Y(n_536) );
INVx2_ASAP7_75t_L g537 ( .A(n_530), .Y(n_537) );
INVx3_ASAP7_75t_L g538 ( .A(n_491), .Y(n_538) );
INVx1_ASAP7_75t_L g539 ( .A(n_530), .Y(n_539) );
OR2x2_ASAP7_75t_L g540 ( .A(n_490), .B(n_476), .Y(n_540) );
AOI22xp5_ASAP7_75t_L g541 ( .A1(n_492), .A2(n_362), .B1(n_377), .B2(n_326), .Y(n_541) );
INVx2_ASAP7_75t_L g542 ( .A(n_530), .Y(n_542) );
OR2x6_ASAP7_75t_L g543 ( .A(n_490), .B(n_463), .Y(n_543) );
INVx3_ASAP7_75t_L g544 ( .A(n_491), .Y(n_544) );
INVx1_ASAP7_75t_L g545 ( .A(n_535), .Y(n_545) );
NAND2xp5_ASAP7_75t_L g546 ( .A(n_494), .B(n_464), .Y(n_546) );
AOI22xp5_ASAP7_75t_L g547 ( .A1(n_492), .A2(n_362), .B1(n_409), .B2(n_392), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g548 ( .A(n_513), .B(n_464), .Y(n_548) );
AND2x4_ASAP7_75t_L g549 ( .A(n_523), .B(n_471), .Y(n_549) );
INVxp67_ASAP7_75t_L g550 ( .A(n_516), .Y(n_550) );
NAND3xp33_ASAP7_75t_L g551 ( .A(n_499), .B(n_467), .C(n_482), .Y(n_551) );
INVx1_ASAP7_75t_L g552 ( .A(n_535), .Y(n_552) );
NAND2xp5_ASAP7_75t_SL g553 ( .A(n_517), .B(n_302), .Y(n_553) );
INVx1_ASAP7_75t_L g554 ( .A(n_488), .Y(n_554) );
AOI22xp5_ASAP7_75t_L g555 ( .A1(n_505), .A2(n_409), .B1(n_392), .B2(n_467), .Y(n_555) );
INVx1_ASAP7_75t_L g556 ( .A(n_523), .Y(n_556) );
BUFx5_ASAP7_75t_L g557 ( .A(n_487), .Y(n_557) );
NOR2xp33_ASAP7_75t_L g558 ( .A(n_498), .B(n_374), .Y(n_558) );
AND2x6_ASAP7_75t_L g559 ( .A(n_501), .B(n_482), .Y(n_559) );
NAND2xp5_ASAP7_75t_L g560 ( .A(n_508), .B(n_371), .Y(n_560) );
NOR2xp33_ASAP7_75t_L g561 ( .A(n_504), .B(n_423), .Y(n_561) );
AOI21xp5_ASAP7_75t_L g562 ( .A1(n_502), .A2(n_485), .B(n_378), .Y(n_562) );
AOI22xp5_ASAP7_75t_L g563 ( .A1(n_505), .A2(n_441), .B1(n_427), .B2(n_423), .Y(n_563) );
INVx3_ASAP7_75t_L g564 ( .A(n_501), .Y(n_564) );
NAND2xp5_ASAP7_75t_SL g565 ( .A(n_517), .B(n_508), .Y(n_565) );
INVxp67_ASAP7_75t_L g566 ( .A(n_516), .Y(n_566) );
INVx2_ASAP7_75t_SL g567 ( .A(n_508), .Y(n_567) );
INVx3_ASAP7_75t_L g568 ( .A(n_501), .Y(n_568) );
AND2x6_ASAP7_75t_SL g569 ( .A(n_519), .B(n_477), .Y(n_569) );
AOI22xp33_ASAP7_75t_L g570 ( .A1(n_487), .A2(n_478), .B1(n_477), .B2(n_321), .Y(n_570) );
NAND2x1_ASAP7_75t_L g571 ( .A(n_487), .B(n_290), .Y(n_571) );
INVx1_ASAP7_75t_L g572 ( .A(n_508), .Y(n_572) );
INVx1_ASAP7_75t_SL g573 ( .A(n_521), .Y(n_573) );
INVx1_ASAP7_75t_L g574 ( .A(n_488), .Y(n_574) );
NAND2xp5_ASAP7_75t_L g575 ( .A(n_515), .B(n_371), .Y(n_575) );
INVx1_ASAP7_75t_L g576 ( .A(n_495), .Y(n_576) );
NAND2xp5_ASAP7_75t_L g577 ( .A(n_515), .B(n_382), .Y(n_577) );
INVx1_ASAP7_75t_SL g578 ( .A(n_527), .Y(n_578) );
INVx5_ASAP7_75t_L g579 ( .A(n_487), .Y(n_579) );
NAND2xp5_ASAP7_75t_SL g580 ( .A(n_517), .B(n_382), .Y(n_580) );
NAND2x1p5_ASAP7_75t_L g581 ( .A(n_514), .B(n_336), .Y(n_581) );
AND2x4_ASAP7_75t_L g582 ( .A(n_517), .B(n_471), .Y(n_582) );
AND2x6_ASAP7_75t_L g583 ( .A(n_501), .B(n_337), .Y(n_583) );
AOI21x1_ASAP7_75t_L g584 ( .A1(n_502), .A2(n_298), .B(n_297), .Y(n_584) );
BUFx2_ASAP7_75t_L g585 ( .A(n_489), .Y(n_585) );
AND2x2_ASAP7_75t_L g586 ( .A(n_524), .B(n_478), .Y(n_586) );
NAND2xp5_ASAP7_75t_SL g587 ( .A(n_528), .B(n_398), .Y(n_587) );
NAND2xp5_ASAP7_75t_L g588 ( .A(n_532), .B(n_398), .Y(n_588) );
AOI22xp5_ASAP7_75t_L g589 ( .A1(n_487), .A2(n_388), .B1(n_434), .B2(n_414), .Y(n_589) );
INVx1_ASAP7_75t_L g590 ( .A(n_495), .Y(n_590) );
BUFx6f_ASAP7_75t_L g591 ( .A(n_487), .Y(n_591) );
AND2x2_ASAP7_75t_SL g592 ( .A(n_524), .B(n_386), .Y(n_592) );
CKINVDCx5p33_ASAP7_75t_R g593 ( .A(n_522), .Y(n_593) );
AOI22xp5_ASAP7_75t_L g594 ( .A1(n_526), .A2(n_386), .B1(n_327), .B2(n_340), .Y(n_594) );
OR2x6_ASAP7_75t_L g595 ( .A(n_512), .B(n_318), .Y(n_595) );
INVx1_ASAP7_75t_L g596 ( .A(n_497), .Y(n_596) );
INVx1_ASAP7_75t_L g597 ( .A(n_497), .Y(n_597) );
NAND2xp5_ASAP7_75t_L g598 ( .A(n_500), .B(n_401), .Y(n_598) );
BUFx3_ASAP7_75t_L g599 ( .A(n_500), .Y(n_599) );
NAND3xp33_ASAP7_75t_SL g600 ( .A(n_520), .B(n_417), .C(n_318), .Y(n_600) );
INVx1_ASAP7_75t_L g601 ( .A(n_503), .Y(n_601) );
CKINVDCx16_ASAP7_75t_R g602 ( .A(n_493), .Y(n_602) );
NAND2xp5_ASAP7_75t_L g603 ( .A(n_520), .B(n_407), .Y(n_603) );
NAND2xp5_ASAP7_75t_L g604 ( .A(n_520), .B(n_407), .Y(n_604) );
INVx1_ASAP7_75t_L g605 ( .A(n_503), .Y(n_605) );
INVx1_ASAP7_75t_L g606 ( .A(n_507), .Y(n_606) );
AOI22xp5_ASAP7_75t_L g607 ( .A1(n_520), .A2(n_319), .B1(n_344), .B2(n_342), .Y(n_607) );
AOI22xp33_ASAP7_75t_L g608 ( .A1(n_496), .A2(n_352), .B1(n_367), .B2(n_348), .Y(n_608) );
AOI22xp5_ASAP7_75t_L g609 ( .A1(n_496), .A2(n_418), .B1(n_426), .B2(n_394), .Y(n_609) );
AND2x4_ASAP7_75t_L g610 ( .A(n_496), .B(n_454), .Y(n_610) );
INVx1_ASAP7_75t_L g611 ( .A(n_507), .Y(n_611) );
NAND2xp5_ASAP7_75t_SL g612 ( .A(n_506), .B(n_444), .Y(n_612) );
OR2x6_ASAP7_75t_L g613 ( .A(n_506), .B(n_417), .Y(n_613) );
INVx2_ASAP7_75t_L g614 ( .A(n_518), .Y(n_614) );
BUFx2_ASAP7_75t_L g615 ( .A(n_518), .Y(n_615) );
NOR3xp33_ASAP7_75t_SL g616 ( .A(n_509), .B(n_445), .C(n_439), .Y(n_616) );
NAND2xp5_ASAP7_75t_L g617 ( .A(n_518), .B(n_445), .Y(n_617) );
AND2x4_ASAP7_75t_L g618 ( .A(n_509), .B(n_458), .Y(n_618) );
INVx1_ASAP7_75t_L g619 ( .A(n_510), .Y(n_619) );
AOI21xp5_ASAP7_75t_L g620 ( .A1(n_510), .A2(n_378), .B(n_354), .Y(n_620) );
INVx1_ASAP7_75t_L g621 ( .A(n_511), .Y(n_621) );
INVx5_ASAP7_75t_L g622 ( .A(n_534), .Y(n_622) );
INVx1_ASAP7_75t_L g623 ( .A(n_511), .Y(n_623) );
NAND2xp5_ASAP7_75t_L g624 ( .A(n_531), .B(n_458), .Y(n_624) );
BUFx4f_ASAP7_75t_L g625 ( .A(n_534), .Y(n_625) );
INVx1_ASAP7_75t_L g626 ( .A(n_534), .Y(n_626) );
INVx2_ASAP7_75t_L g627 ( .A(n_531), .Y(n_627) );
NOR2xp67_ASAP7_75t_L g628 ( .A(n_531), .B(n_461), .Y(n_628) );
INVx2_ASAP7_75t_L g629 ( .A(n_564), .Y(n_629) );
OAI21xp33_ASAP7_75t_L g630 ( .A1(n_548), .A2(n_447), .B(n_347), .Y(n_630) );
AOI22xp33_ASAP7_75t_L g631 ( .A1(n_559), .A2(n_469), .B1(n_474), .B2(n_461), .Y(n_631) );
BUFx12f_ASAP7_75t_L g632 ( .A(n_593), .Y(n_632) );
BUFx8_ASAP7_75t_SL g633 ( .A(n_585), .Y(n_633) );
INVx3_ASAP7_75t_L g634 ( .A(n_538), .Y(n_634) );
BUFx12f_ASAP7_75t_L g635 ( .A(n_613), .Y(n_635) );
AOI21xp5_ASAP7_75t_L g636 ( .A1(n_536), .A2(n_335), .B(n_305), .Y(n_636) );
INVx1_ASAP7_75t_L g637 ( .A(n_572), .Y(n_637) );
AND2x2_ASAP7_75t_L g638 ( .A(n_550), .B(n_469), .Y(n_638) );
AOI21x1_ASAP7_75t_L g639 ( .A1(n_584), .A2(n_525), .B(n_486), .Y(n_639) );
BUFx2_ASAP7_75t_L g640 ( .A(n_613), .Y(n_640) );
CKINVDCx5p33_ASAP7_75t_R g641 ( .A(n_595), .Y(n_641) );
INVx2_ASAP7_75t_L g642 ( .A(n_564), .Y(n_642) );
INVx4_ASAP7_75t_L g643 ( .A(n_579), .Y(n_643) );
INVx1_ASAP7_75t_L g644 ( .A(n_567), .Y(n_644) );
NAND2xp5_ASAP7_75t_SL g645 ( .A(n_591), .B(n_300), .Y(n_645) );
AND2x4_ASAP7_75t_SL g646 ( .A(n_582), .B(n_474), .Y(n_646) );
INVx3_ASAP7_75t_L g647 ( .A(n_538), .Y(n_647) );
AND2x4_ASAP7_75t_SL g648 ( .A(n_582), .B(n_481), .Y(n_648) );
INVx1_ASAP7_75t_L g649 ( .A(n_565), .Y(n_649) );
INVx5_ASAP7_75t_L g650 ( .A(n_591), .Y(n_650) );
AND2x4_ASAP7_75t_L g651 ( .A(n_549), .B(n_481), .Y(n_651) );
A2O1A1Ixp33_ASAP7_75t_SL g652 ( .A1(n_558), .A2(n_446), .B(n_531), .C(n_480), .Y(n_652) );
NOR2xp33_ASAP7_75t_L g653 ( .A(n_566), .B(n_293), .Y(n_653) );
INVx2_ASAP7_75t_L g654 ( .A(n_568), .Y(n_654) );
INVx3_ASAP7_75t_L g655 ( .A(n_544), .Y(n_655) );
BUFx6f_ASAP7_75t_L g656 ( .A(n_591), .Y(n_656) );
HB1xp67_ASAP7_75t_L g657 ( .A(n_602), .Y(n_657) );
INVx5_ASAP7_75t_L g658 ( .A(n_579), .Y(n_658) );
INVxp67_ASAP7_75t_L g659 ( .A(n_540), .Y(n_659) );
BUFx2_ASAP7_75t_SL g660 ( .A(n_579), .Y(n_660) );
A2O1A1Ixp33_ASAP7_75t_L g661 ( .A1(n_546), .A2(n_383), .B(n_307), .C(n_312), .Y(n_661) );
INVx4_ASAP7_75t_L g662 ( .A(n_544), .Y(n_662) );
INVx4_ASAP7_75t_L g663 ( .A(n_557), .Y(n_663) );
INVx2_ASAP7_75t_L g664 ( .A(n_568), .Y(n_664) );
INVx2_ASAP7_75t_L g665 ( .A(n_537), .Y(n_665) );
BUFx3_ASAP7_75t_L g666 ( .A(n_549), .Y(n_666) );
NOR2xp33_ASAP7_75t_L g667 ( .A(n_563), .B(n_303), .Y(n_667) );
OAI22xp5_ASAP7_75t_L g668 ( .A1(n_570), .A2(n_408), .B1(n_433), .B2(n_395), .Y(n_668) );
BUFx2_ASAP7_75t_L g669 ( .A(n_595), .Y(n_669) );
INVx3_ASAP7_75t_L g670 ( .A(n_599), .Y(n_670) );
AOI22xp33_ASAP7_75t_L g671 ( .A1(n_559), .A2(n_315), .B1(n_316), .B2(n_309), .Y(n_671) );
INVx2_ASAP7_75t_L g672 ( .A(n_542), .Y(n_672) );
INVx1_ASAP7_75t_L g673 ( .A(n_610), .Y(n_673) );
AOI21xp5_ASAP7_75t_L g674 ( .A1(n_554), .A2(n_438), .B(n_436), .Y(n_674) );
O2A1O1Ixp5_ASAP7_75t_L g675 ( .A1(n_571), .A2(n_446), .B(n_381), .C(n_389), .Y(n_675) );
BUFx6f_ASAP7_75t_L g676 ( .A(n_625), .Y(n_676) );
NAND2xp5_ASAP7_75t_L g677 ( .A(n_573), .B(n_578), .Y(n_677) );
CKINVDCx6p67_ASAP7_75t_R g678 ( .A(n_543), .Y(n_678) );
INVx2_ASAP7_75t_L g679 ( .A(n_539), .Y(n_679) );
INVx2_ASAP7_75t_L g680 ( .A(n_545), .Y(n_680) );
OAI22xp33_ASAP7_75t_L g681 ( .A1(n_541), .A2(n_317), .B1(n_322), .B2(n_320), .Y(n_681) );
BUFx3_ASAP7_75t_L g682 ( .A(n_610), .Y(n_682) );
A2O1A1Ixp33_ASAP7_75t_L g683 ( .A1(n_551), .A2(n_323), .B(n_328), .C(n_325), .Y(n_683) );
NAND2xp5_ASAP7_75t_L g684 ( .A(n_559), .B(n_329), .Y(n_684) );
INVx2_ASAP7_75t_L g685 ( .A(n_552), .Y(n_685) );
BUFx2_ASAP7_75t_L g686 ( .A(n_547), .Y(n_686) );
INVx1_ASAP7_75t_L g687 ( .A(n_618), .Y(n_687) );
INVx2_ASAP7_75t_L g688 ( .A(n_554), .Y(n_688) );
INVx2_ASAP7_75t_L g689 ( .A(n_574), .Y(n_689) );
AND2x4_ASAP7_75t_L g690 ( .A(n_556), .B(n_333), .Y(n_690) );
A2O1A1Ixp33_ASAP7_75t_L g691 ( .A1(n_561), .A2(n_338), .B(n_339), .C(n_334), .Y(n_691) );
INVx1_ASAP7_75t_L g692 ( .A(n_618), .Y(n_692) );
INVx5_ASAP7_75t_L g693 ( .A(n_583), .Y(n_693) );
INVx1_ASAP7_75t_L g694 ( .A(n_576), .Y(n_694) );
NOR2xp33_ASAP7_75t_L g695 ( .A(n_569), .B(n_324), .Y(n_695) );
INVx3_ASAP7_75t_L g696 ( .A(n_625), .Y(n_696) );
AOI222xp33_ASAP7_75t_L g697 ( .A1(n_592), .A2(n_376), .B1(n_431), .B2(n_343), .C1(n_345), .C2(n_346), .Y(n_697) );
HB1xp67_ASAP7_75t_L g698 ( .A(n_575), .Y(n_698) );
INVx2_ASAP7_75t_L g699 ( .A(n_590), .Y(n_699) );
NAND2xp5_ASAP7_75t_SL g700 ( .A(n_557), .B(n_349), .Y(n_700) );
OAI22xp5_ASAP7_75t_L g701 ( .A1(n_543), .A2(n_353), .B1(n_355), .B2(n_350), .Y(n_701) );
NOR2xp33_ASAP7_75t_R g702 ( .A(n_600), .B(n_13), .Y(n_702) );
AOI22xp5_ASAP7_75t_L g703 ( .A1(n_559), .A2(n_356), .B1(n_358), .B2(n_357), .Y(n_703) );
BUFx6f_ASAP7_75t_L g704 ( .A(n_583), .Y(n_704) );
AOI22xp33_ASAP7_75t_L g705 ( .A1(n_586), .A2(n_360), .B1(n_364), .B2(n_361), .Y(n_705) );
AND2x2_ASAP7_75t_L g706 ( .A(n_555), .B(n_14), .Y(n_706) );
INVx2_ASAP7_75t_L g707 ( .A(n_596), .Y(n_707) );
O2A1O1Ixp33_ASAP7_75t_L g708 ( .A1(n_577), .A2(n_365), .B(n_369), .C(n_368), .Y(n_708) );
INVxp67_ASAP7_75t_SL g709 ( .A(n_557), .Y(n_709) );
INVx1_ASAP7_75t_L g710 ( .A(n_597), .Y(n_710) );
AOI21xp5_ASAP7_75t_L g711 ( .A1(n_562), .A2(n_380), .B(n_373), .Y(n_711) );
INVx2_ASAP7_75t_L g712 ( .A(n_601), .Y(n_712) );
O2A1O1Ixp33_ASAP7_75t_L g713 ( .A1(n_560), .A2(n_399), .B(n_403), .C(n_384), .Y(n_713) );
INVx2_ASAP7_75t_L g714 ( .A(n_605), .Y(n_714) );
CKINVDCx8_ASAP7_75t_R g715 ( .A(n_583), .Y(n_715) );
AND2x4_ASAP7_75t_L g716 ( .A(n_553), .B(n_410), .Y(n_716) );
INVx2_ASAP7_75t_SL g717 ( .A(n_581), .Y(n_717) );
BUFx2_ASAP7_75t_L g718 ( .A(n_583), .Y(n_718) );
INVx1_ASAP7_75t_L g719 ( .A(n_624), .Y(n_719) );
INVx2_ASAP7_75t_L g720 ( .A(n_606), .Y(n_720) );
INVx1_ASAP7_75t_L g721 ( .A(n_611), .Y(n_721) );
INVx2_ASAP7_75t_L g722 ( .A(n_619), .Y(n_722) );
INVx1_ASAP7_75t_L g723 ( .A(n_621), .Y(n_723) );
INVx2_ASAP7_75t_L g724 ( .A(n_623), .Y(n_724) );
NAND2xp5_ASAP7_75t_L g725 ( .A(n_589), .B(n_412), .Y(n_725) );
BUFx6f_ASAP7_75t_L g726 ( .A(n_615), .Y(n_726) );
HB1xp67_ASAP7_75t_SL g727 ( .A(n_616), .Y(n_727) );
AND2x2_ASAP7_75t_L g728 ( .A(n_594), .B(n_15), .Y(n_728) );
AOI21xp5_ASAP7_75t_L g729 ( .A1(n_598), .A2(n_421), .B(n_416), .Y(n_729) );
OAI21xp33_ASAP7_75t_L g730 ( .A1(n_588), .A2(n_429), .B(n_428), .Y(n_730) );
INVx8_ASAP7_75t_L g731 ( .A(n_622), .Y(n_731) );
INVx5_ASAP7_75t_L g732 ( .A(n_622), .Y(n_732) );
INVx1_ASAP7_75t_L g733 ( .A(n_607), .Y(n_733) );
INVxp67_ASAP7_75t_L g734 ( .A(n_580), .Y(n_734) );
INVx1_ASAP7_75t_L g735 ( .A(n_609), .Y(n_735) );
A2O1A1Ixp33_ASAP7_75t_L g736 ( .A1(n_620), .A2(n_440), .B(n_442), .C(n_430), .Y(n_736) );
NAND3xp33_ASAP7_75t_L g737 ( .A(n_608), .B(n_443), .C(n_381), .Y(n_737) );
BUFx2_ASAP7_75t_L g738 ( .A(n_603), .Y(n_738) );
CKINVDCx20_ASAP7_75t_R g739 ( .A(n_557), .Y(n_739) );
INVx3_ASAP7_75t_L g740 ( .A(n_614), .Y(n_740) );
NAND2xp5_ASAP7_75t_SL g741 ( .A(n_557), .B(n_354), .Y(n_741) );
O2A1O1Ixp33_ASAP7_75t_L g742 ( .A1(n_587), .A2(n_389), .B(n_402), .C(n_400), .Y(n_742) );
INVx6_ASAP7_75t_L g743 ( .A(n_622), .Y(n_743) );
AOI21xp5_ASAP7_75t_L g744 ( .A1(n_604), .A2(n_437), .B(n_425), .Y(n_744) );
NAND2xp5_ASAP7_75t_L g745 ( .A(n_617), .B(n_448), .Y(n_745) );
CKINVDCx5p33_ASAP7_75t_R g746 ( .A(n_612), .Y(n_746) );
AOI21xp5_ASAP7_75t_L g747 ( .A1(n_627), .A2(n_448), .B(n_486), .Y(n_747) );
BUFx12f_ASAP7_75t_L g748 ( .A(n_628), .Y(n_748) );
INVxp67_ASAP7_75t_L g749 ( .A(n_626), .Y(n_749) );
AND2x4_ASAP7_75t_L g750 ( .A(n_582), .B(n_405), .Y(n_750) );
INVx3_ASAP7_75t_L g751 ( .A(n_538), .Y(n_751) );
BUFx12f_ASAP7_75t_L g752 ( .A(n_593), .Y(n_752) );
AOI21x1_ASAP7_75t_L g753 ( .A1(n_584), .A2(n_525), .B(n_486), .Y(n_753) );
NAND2xp5_ASAP7_75t_L g754 ( .A(n_546), .B(n_366), .Y(n_754) );
INVx1_ASAP7_75t_L g755 ( .A(n_572), .Y(n_755) );
HB1xp67_ASAP7_75t_L g756 ( .A(n_550), .Y(n_756) );
NOR2xp33_ASAP7_75t_L g757 ( .A(n_550), .B(n_15), .Y(n_757) );
NAND2xp5_ASAP7_75t_SL g758 ( .A(n_591), .B(n_366), .Y(n_758) );
AOI21xp33_ASAP7_75t_L g759 ( .A1(n_571), .A2(n_404), .B(n_332), .Y(n_759) );
OAI22xp33_ASAP7_75t_L g760 ( .A1(n_541), .A2(n_404), .B1(n_332), .B2(n_363), .Y(n_760) );
O2A1O1Ixp33_ASAP7_75t_L g761 ( .A1(n_550), .A2(n_480), .B(n_484), .C(n_453), .Y(n_761) );
NAND2xp5_ASAP7_75t_SL g762 ( .A(n_591), .B(n_311), .Y(n_762) );
NAND2xp5_ASAP7_75t_L g763 ( .A(n_546), .B(n_480), .Y(n_763) );
AOI21xp5_ASAP7_75t_L g764 ( .A1(n_548), .A2(n_529), .B(n_525), .Y(n_764) );
AOI21xp5_ASAP7_75t_L g765 ( .A1(n_548), .A2(n_533), .B(n_529), .Y(n_765) );
INVx3_ASAP7_75t_L g766 ( .A(n_538), .Y(n_766) );
INVxp67_ASAP7_75t_SL g767 ( .A(n_591), .Y(n_767) );
A2O1A1Ixp33_ASAP7_75t_L g768 ( .A1(n_548), .A2(n_484), .B(n_363), .C(n_332), .Y(n_768) );
NAND2xp5_ASAP7_75t_L g769 ( .A(n_546), .B(n_484), .Y(n_769) );
NAND2xp5_ASAP7_75t_SL g770 ( .A(n_591), .B(n_332), .Y(n_770) );
INVx1_ASAP7_75t_L g771 ( .A(n_572), .Y(n_771) );
AOI21xp5_ASAP7_75t_L g772 ( .A1(n_548), .A2(n_533), .B(n_529), .Y(n_772) );
OAI21x1_ASAP7_75t_L g773 ( .A1(n_639), .A2(n_533), .B(n_397), .Y(n_773) );
AOI22xp33_ASAP7_75t_SL g774 ( .A1(n_669), .A2(n_363), .B1(n_397), .B2(n_19), .Y(n_774) );
INVx1_ASAP7_75t_L g775 ( .A(n_677), .Y(n_775) );
INVx1_ASAP7_75t_L g776 ( .A(n_677), .Y(n_776) );
OA21x2_ASAP7_75t_L g777 ( .A1(n_753), .A2(n_397), .B(n_363), .Y(n_777) );
INVx2_ASAP7_75t_L g778 ( .A(n_688), .Y(n_778) );
NOR2xp33_ASAP7_75t_L g779 ( .A(n_659), .B(n_686), .Y(n_779) );
HB1xp67_ASAP7_75t_L g780 ( .A(n_756), .Y(n_780) );
INVx4_ASAP7_75t_L g781 ( .A(n_731), .Y(n_781) );
OAI21x1_ASAP7_75t_L g782 ( .A1(n_747), .A2(n_397), .B(n_465), .Y(n_782) );
AOI22xp33_ASAP7_75t_L g783 ( .A1(n_706), .A2(n_472), .B1(n_465), .B2(n_19), .Y(n_783) );
HB1xp67_ASAP7_75t_L g784 ( .A(n_651), .Y(n_784) );
BUFx3_ASAP7_75t_L g785 ( .A(n_633), .Y(n_785) );
NOR2xp67_ASAP7_75t_L g786 ( .A(n_632), .B(n_16), .Y(n_786) );
BUFx6f_ASAP7_75t_L g787 ( .A(n_656), .Y(n_787) );
INVx1_ASAP7_75t_L g788 ( .A(n_721), .Y(n_788) );
INVx3_ASAP7_75t_SL g789 ( .A(n_731), .Y(n_789) );
NAND2xp5_ASAP7_75t_L g790 ( .A(n_733), .B(n_17), .Y(n_790) );
OAI21xp5_ASAP7_75t_L g791 ( .A1(n_744), .A2(n_472), .B(n_17), .Y(n_791) );
BUFx10_ASAP7_75t_L g792 ( .A(n_646), .Y(n_792) );
AOI21xp5_ASAP7_75t_L g793 ( .A1(n_711), .A2(n_79), .B(n_78), .Y(n_793) );
NAND2x1p5_ASAP7_75t_L g794 ( .A(n_693), .B(n_20), .Y(n_794) );
OAI22xp5_ASAP7_75t_L g795 ( .A1(n_631), .A2(n_20), .B1(n_21), .B2(n_22), .Y(n_795) );
OAI22xp5_ASAP7_75t_L g796 ( .A1(n_703), .A2(n_21), .B1(n_23), .B2(n_25), .Y(n_796) );
INVx1_ASAP7_75t_L g797 ( .A(n_723), .Y(n_797) );
INVx2_ASAP7_75t_L g798 ( .A(n_689), .Y(n_798) );
NAND2xp5_ASAP7_75t_L g799 ( .A(n_735), .B(n_23), .Y(n_799) );
OA21x2_ASAP7_75t_L g800 ( .A1(n_768), .A2(n_81), .B(n_80), .Y(n_800) );
OAI222xp33_ASAP7_75t_L g801 ( .A1(n_641), .A2(n_25), .B1(n_26), .B2(n_27), .C1(n_28), .C2(n_29), .Y(n_801) );
NOR2xp33_ASAP7_75t_L g802 ( .A(n_678), .B(n_26), .Y(n_802) );
INVx1_ASAP7_75t_L g803 ( .A(n_763), .Y(n_803) );
AOI21xp5_ASAP7_75t_L g804 ( .A1(n_711), .A2(n_85), .B(n_84), .Y(n_804) );
NOR2xp33_ASAP7_75t_L g805 ( .A(n_640), .B(n_27), .Y(n_805) );
INVx4_ASAP7_75t_L g806 ( .A(n_731), .Y(n_806) );
OAI21x1_ASAP7_75t_L g807 ( .A1(n_772), .A2(n_89), .B(n_88), .Y(n_807) );
AO31x2_ASAP7_75t_L g808 ( .A1(n_683), .A2(n_28), .A3(n_30), .B(n_32), .Y(n_808) );
OAI21x1_ASAP7_75t_L g809 ( .A1(n_764), .A2(n_91), .B(n_90), .Y(n_809) );
INVx1_ASAP7_75t_L g810 ( .A(n_763), .Y(n_810) );
BUFx2_ASAP7_75t_L g811 ( .A(n_657), .Y(n_811) );
NAND2x1p5_ASAP7_75t_L g812 ( .A(n_693), .B(n_33), .Y(n_812) );
BUFx4f_ASAP7_75t_L g813 ( .A(n_752), .Y(n_813) );
INVx1_ASAP7_75t_L g814 ( .A(n_769), .Y(n_814) );
AOI22xp33_ASAP7_75t_L g815 ( .A1(n_728), .A2(n_33), .B1(n_36), .B2(n_38), .Y(n_815) );
NOR2xp33_ASAP7_75t_L g816 ( .A(n_666), .B(n_39), .Y(n_816) );
INVx1_ASAP7_75t_L g817 ( .A(n_769), .Y(n_817) );
NAND2xp5_ASAP7_75t_L g818 ( .A(n_694), .B(n_39), .Y(n_818) );
O2A1O1Ixp33_ASAP7_75t_SL g819 ( .A1(n_736), .A2(n_169), .B(n_288), .C(n_286), .Y(n_819) );
AO31x2_ASAP7_75t_L g820 ( .A1(n_661), .A2(n_40), .A3(n_42), .B(n_43), .Y(n_820) );
INVx1_ASAP7_75t_L g821 ( .A(n_712), .Y(n_821) );
BUFx6f_ASAP7_75t_L g822 ( .A(n_656), .Y(n_822) );
AOI22xp33_ASAP7_75t_L g823 ( .A1(n_697), .A2(n_40), .B1(n_42), .B2(n_43), .Y(n_823) );
NOR2x1_ASAP7_75t_R g824 ( .A(n_635), .B(n_44), .Y(n_824) );
AO22x2_ASAP7_75t_L g825 ( .A1(n_701), .A2(n_45), .B1(n_46), .B2(n_47), .Y(n_825) );
A2O1A1Ixp33_ASAP7_75t_L g826 ( .A1(n_713), .A2(n_708), .B(n_729), .C(n_742), .Y(n_826) );
INVx2_ASAP7_75t_L g827 ( .A(n_699), .Y(n_827) );
INVx1_ASAP7_75t_L g828 ( .A(n_714), .Y(n_828) );
INVx1_ASAP7_75t_L g829 ( .A(n_720), .Y(n_829) );
OAI21x1_ASAP7_75t_L g830 ( .A1(n_764), .A2(n_98), .B(n_97), .Y(n_830) );
OAI21x1_ASAP7_75t_L g831 ( .A1(n_765), .A2(n_105), .B(n_103), .Y(n_831) );
AOI22xp33_ASAP7_75t_L g832 ( .A1(n_697), .A2(n_45), .B1(n_47), .B2(n_48), .Y(n_832) );
OAI21x1_ASAP7_75t_L g833 ( .A1(n_765), .A2(n_108), .B(n_107), .Y(n_833) );
AND2x4_ASAP7_75t_L g834 ( .A(n_648), .B(n_48), .Y(n_834) );
INVx2_ASAP7_75t_L g835 ( .A(n_707), .Y(n_835) );
AOI22xp33_ASAP7_75t_L g836 ( .A1(n_667), .A2(n_49), .B1(n_50), .B2(n_51), .Y(n_836) );
OAI22xp5_ASAP7_75t_L g837 ( .A1(n_671), .A2(n_51), .B1(n_52), .B2(n_53), .Y(n_837) );
CKINVDCx5p33_ASAP7_75t_R g838 ( .A(n_727), .Y(n_838) );
OAI21x1_ASAP7_75t_SL g839 ( .A1(n_722), .A2(n_52), .B(n_55), .Y(n_839) );
NAND2xp5_ASAP7_75t_L g840 ( .A(n_710), .B(n_724), .Y(n_840) );
AOI22xp33_ASAP7_75t_L g841 ( .A1(n_698), .A2(n_55), .B1(n_57), .B2(n_58), .Y(n_841) );
INVx1_ASAP7_75t_L g842 ( .A(n_649), .Y(n_842) );
OA21x2_ASAP7_75t_L g843 ( .A1(n_675), .A2(n_185), .B(n_285), .Y(n_843) );
INVx2_ASAP7_75t_L g844 ( .A(n_679), .Y(n_844) );
NAND2xp5_ASAP7_75t_L g845 ( .A(n_637), .B(n_58), .Y(n_845) );
INVxp67_ASAP7_75t_L g846 ( .A(n_651), .Y(n_846) );
INVx1_ASAP7_75t_L g847 ( .A(n_638), .Y(n_847) );
INVx2_ASAP7_75t_L g848 ( .A(n_680), .Y(n_848) );
NAND2xp5_ASAP7_75t_L g849 ( .A(n_755), .B(n_59), .Y(n_849) );
OAI211xp5_ASAP7_75t_SL g850 ( .A1(n_705), .A2(n_59), .B(n_60), .C(n_61), .Y(n_850) );
AOI32xp33_ASAP7_75t_L g851 ( .A1(n_701), .A2(n_60), .A3(n_62), .B1(n_63), .B2(n_64), .Y(n_851) );
OAI21xp5_ASAP7_75t_L g852 ( .A1(n_674), .A2(n_62), .B(n_63), .Y(n_852) );
AND2x2_ASAP7_75t_L g853 ( .A(n_653), .B(n_65), .Y(n_853) );
INVx1_ASAP7_75t_L g854 ( .A(n_687), .Y(n_854) );
OAI21x1_ASAP7_75t_L g855 ( .A1(n_741), .A2(n_191), .B(n_284), .Y(n_855) );
OAI21x1_ASAP7_75t_L g856 ( .A1(n_758), .A2(n_187), .B(n_283), .Y(n_856) );
NAND2xp5_ASAP7_75t_L g857 ( .A(n_771), .B(n_66), .Y(n_857) );
INVx1_ASAP7_75t_L g858 ( .A(n_692), .Y(n_858) );
AOI22xp33_ASAP7_75t_L g859 ( .A1(n_695), .A2(n_67), .B1(n_68), .B2(n_69), .Y(n_859) );
AOI22xp33_ASAP7_75t_L g860 ( .A1(n_757), .A2(n_67), .B1(n_68), .B2(n_69), .Y(n_860) );
AND2x2_ASAP7_75t_L g861 ( .A(n_690), .B(n_70), .Y(n_861) );
OAI21xp5_ASAP7_75t_L g862 ( .A1(n_674), .A2(n_70), .B(n_71), .Y(n_862) );
OAI21x1_ASAP7_75t_L g863 ( .A1(n_762), .A2(n_186), .B(n_277), .Y(n_863) );
INVx2_ASAP7_75t_L g864 ( .A(n_685), .Y(n_864) );
INVx1_ASAP7_75t_L g865 ( .A(n_754), .Y(n_865) );
INVx5_ASAP7_75t_L g866 ( .A(n_704), .Y(n_866) );
A2O1A1Ixp33_ASAP7_75t_L g867 ( .A1(n_713), .A2(n_71), .B(n_72), .C(n_73), .Y(n_867) );
AND2x2_ASAP7_75t_L g868 ( .A(n_690), .B(n_72), .Y(n_868) );
CKINVDCx5p33_ASAP7_75t_R g869 ( .A(n_702), .Y(n_869) );
NAND2xp5_ASAP7_75t_L g870 ( .A(n_719), .B(n_74), .Y(n_870) );
AOI22xp33_ASAP7_75t_L g871 ( .A1(n_684), .A2(n_74), .B1(n_75), .B2(n_76), .Y(n_871) );
INVx2_ASAP7_75t_L g872 ( .A(n_665), .Y(n_872) );
OAI21x1_ASAP7_75t_L g873 ( .A1(n_770), .A2(n_192), .B(n_274), .Y(n_873) );
INVx3_ASAP7_75t_L g874 ( .A(n_670), .Y(n_874) );
BUFx3_ASAP7_75t_L g875 ( .A(n_748), .Y(n_875) );
OR2x2_ASAP7_75t_L g876 ( .A(n_684), .B(n_75), .Y(n_876) );
OAI22x1_ASAP7_75t_L g877 ( .A1(n_717), .A2(n_76), .B1(n_114), .B2(n_115), .Y(n_877) );
BUFx6f_ASAP7_75t_L g878 ( .A(n_656), .Y(n_878) );
AND2x2_ASAP7_75t_L g879 ( .A(n_682), .B(n_121), .Y(n_879) );
AOI21xp5_ASAP7_75t_L g880 ( .A1(n_745), .A2(n_122), .B(n_124), .Y(n_880) );
NOR2xp67_ASAP7_75t_SL g881 ( .A(n_715), .B(n_125), .Y(n_881) );
INVx1_ASAP7_75t_SL g882 ( .A(n_726), .Y(n_882) );
BUFx6f_ASAP7_75t_L g883 ( .A(n_650), .Y(n_883) );
INVx2_ASAP7_75t_L g884 ( .A(n_672), .Y(n_884) );
A2O1A1Ixp33_ASAP7_75t_L g885 ( .A1(n_729), .A2(n_141), .B(n_142), .C(n_143), .Y(n_885) );
INVxp67_ASAP7_75t_SL g886 ( .A(n_704), .Y(n_886) );
NAND2xp5_ASAP7_75t_L g887 ( .A(n_754), .B(n_725), .Y(n_887) );
CKINVDCx16_ASAP7_75t_R g888 ( .A(n_750), .Y(n_888) );
OAI21xp5_ASAP7_75t_L g889 ( .A1(n_691), .A2(n_148), .B(n_152), .Y(n_889) );
OAI21x1_ASAP7_75t_L g890 ( .A1(n_740), .A2(n_153), .B(n_154), .Y(n_890) );
OA21x2_ASAP7_75t_L g891 ( .A1(n_759), .A2(n_157), .B(n_158), .Y(n_891) );
AOI22xp33_ASAP7_75t_L g892 ( .A1(n_716), .A2(n_160), .B1(n_161), .B2(n_163), .Y(n_892) );
INVxp67_ASAP7_75t_L g893 ( .A(n_738), .Y(n_893) );
AO31x2_ASAP7_75t_L g894 ( .A1(n_668), .A2(n_164), .A3(n_166), .B(n_167), .Y(n_894) );
OAI21x1_ASAP7_75t_L g895 ( .A1(n_700), .A2(n_168), .B(n_170), .Y(n_895) );
AOI221xp5_ASAP7_75t_L g896 ( .A1(n_681), .A2(n_668), .B1(n_725), .B2(n_760), .C(n_750), .Y(n_896) );
NOR2x1_ASAP7_75t_R g897 ( .A(n_693), .B(n_175), .Y(n_897) );
INVxp67_ASAP7_75t_SL g898 ( .A(n_704), .Y(n_898) );
OAI22xp33_ASAP7_75t_L g899 ( .A1(n_693), .A2(n_176), .B1(n_178), .B2(n_179), .Y(n_899) );
NAND2xp5_ASAP7_75t_L g900 ( .A(n_716), .B(n_183), .Y(n_900) );
NOR2xp67_ASAP7_75t_L g901 ( .A(n_734), .B(n_184), .Y(n_901) );
OAI21x1_ASAP7_75t_L g902 ( .A1(n_742), .A2(n_193), .B(n_194), .Y(n_902) );
INVx1_ASAP7_75t_L g903 ( .A(n_673), .Y(n_903) );
OAI21xp5_ASAP7_75t_L g904 ( .A1(n_737), .A2(n_195), .B(n_198), .Y(n_904) );
OAI21xp5_ASAP7_75t_L g905 ( .A1(n_737), .A2(n_200), .B(n_201), .Y(n_905) );
A2O1A1Ixp33_ASAP7_75t_L g906 ( .A1(n_730), .A2(n_204), .B(n_207), .C(n_209), .Y(n_906) );
AOI22xp33_ASAP7_75t_L g907 ( .A1(n_726), .A2(n_210), .B1(n_211), .B2(n_212), .Y(n_907) );
AOI22xp5_ASAP7_75t_L g908 ( .A1(n_630), .A2(n_217), .B1(n_222), .B2(n_226), .Y(n_908) );
CKINVDCx6p67_ASAP7_75t_R g909 ( .A(n_732), .Y(n_909) );
INVx1_ASAP7_75t_L g910 ( .A(n_644), .Y(n_910) );
BUFx6f_ASAP7_75t_L g911 ( .A(n_650), .Y(n_911) );
OR2x6_ASAP7_75t_L g912 ( .A(n_660), .B(n_229), .Y(n_912) );
AO21x2_ASAP7_75t_L g913 ( .A1(n_636), .A2(n_230), .B(n_231), .Y(n_913) );
AOI22xp33_ASAP7_75t_L g914 ( .A1(n_726), .A2(n_235), .B1(n_237), .B2(n_238), .Y(n_914) );
AO21x2_ASAP7_75t_L g915 ( .A1(n_636), .A2(n_239), .B(n_244), .Y(n_915) );
NAND2xp5_ASAP7_75t_L g916 ( .A(n_670), .B(n_246), .Y(n_916) );
INVx1_ASAP7_75t_L g917 ( .A(n_761), .Y(n_917) );
INVx1_ASAP7_75t_L g918 ( .A(n_629), .Y(n_918) );
INVx1_ASAP7_75t_L g919 ( .A(n_642), .Y(n_919) );
INVx1_ASAP7_75t_SL g920 ( .A(n_650), .Y(n_920) );
AOI22xp33_ASAP7_75t_L g921 ( .A1(n_634), .A2(n_248), .B1(n_249), .B2(n_250), .Y(n_921) );
AND2x2_ASAP7_75t_L g922 ( .A(n_746), .B(n_252), .Y(n_922) );
INVx1_ASAP7_75t_L g923 ( .A(n_775), .Y(n_923) );
AOI221xp5_ASAP7_75t_L g924 ( .A1(n_779), .A2(n_655), .B1(n_766), .B2(n_751), .C(n_647), .Y(n_924) );
AND2x4_ASAP7_75t_SL g925 ( .A(n_781), .B(n_676), .Y(n_925) );
INVx2_ASAP7_75t_L g926 ( .A(n_798), .Y(n_926) );
OA21x2_ASAP7_75t_L g927 ( .A1(n_773), .A2(n_749), .B(n_709), .Y(n_927) );
AND2x4_ASAP7_75t_L g928 ( .A(n_781), .B(n_806), .Y(n_928) );
AOI22xp33_ASAP7_75t_L g929 ( .A1(n_896), .A2(n_634), .B1(n_766), .B2(n_751), .Y(n_929) );
OAI22xp33_ASAP7_75t_L g930 ( .A1(n_893), .A2(n_718), .B1(n_739), .B2(n_663), .Y(n_930) );
AOI21xp5_ASAP7_75t_L g931 ( .A1(n_887), .A2(n_645), .B(n_767), .Y(n_931) );
CKINVDCx20_ASAP7_75t_R g932 ( .A(n_785), .Y(n_932) );
HB1xp67_ASAP7_75t_L g933 ( .A(n_780), .Y(n_933) );
INVx1_ASAP7_75t_L g934 ( .A(n_776), .Y(n_934) );
NAND2xp5_ASAP7_75t_L g935 ( .A(n_810), .B(n_654), .Y(n_935) );
AND2x2_ASAP7_75t_L g936 ( .A(n_893), .B(n_732), .Y(n_936) );
OAI21xp5_ASAP7_75t_L g937 ( .A1(n_865), .A2(n_664), .B(n_663), .Y(n_937) );
INVx3_ASAP7_75t_L g938 ( .A(n_806), .Y(n_938) );
AOI22xp33_ASAP7_75t_L g939 ( .A1(n_896), .A2(n_655), .B1(n_647), .B2(n_662), .Y(n_939) );
OAI221xp5_ASAP7_75t_L g940 ( .A1(n_823), .A2(n_662), .B1(n_696), .B2(n_743), .C(n_643), .Y(n_940) );
AOI22xp33_ASAP7_75t_SL g941 ( .A1(n_834), .A2(n_658), .B1(n_676), .B2(n_643), .Y(n_941) );
INVx2_ASAP7_75t_L g942 ( .A(n_827), .Y(n_942) );
INVx1_ASAP7_75t_L g943 ( .A(n_788), .Y(n_943) );
NAND3xp33_ASAP7_75t_L g944 ( .A(n_774), .B(n_791), .C(n_867), .Y(n_944) );
INVx2_ASAP7_75t_L g945 ( .A(n_835), .Y(n_945) );
OAI22xp33_ASAP7_75t_L g946 ( .A1(n_780), .A2(n_658), .B1(n_676), .B2(n_732), .Y(n_946) );
NAND2xp5_ASAP7_75t_L g947 ( .A(n_814), .B(n_658), .Y(n_947) );
AOI221xp5_ASAP7_75t_L g948 ( .A1(n_847), .A2(n_732), .B1(n_658), .B2(n_743), .C(n_262), .Y(n_948) );
AND2x2_ASAP7_75t_L g949 ( .A(n_789), .B(n_255), .Y(n_949) );
OAI22xp5_ASAP7_75t_L g950 ( .A1(n_817), .A2(n_258), .B1(n_260), .B2(n_263), .Y(n_950) );
INVx1_ASAP7_75t_L g951 ( .A(n_797), .Y(n_951) );
NAND2xp5_ASAP7_75t_L g952 ( .A(n_887), .B(n_265), .Y(n_952) );
A2O1A1Ixp33_ASAP7_75t_L g953 ( .A1(n_826), .A2(n_266), .B(n_267), .C(n_268), .Y(n_953) );
BUFx6f_ASAP7_75t_L g954 ( .A(n_789), .Y(n_954) );
INVx1_ASAP7_75t_L g955 ( .A(n_821), .Y(n_955) );
AOI22xp33_ASAP7_75t_L g956 ( .A1(n_861), .A2(n_289), .B1(n_868), .B2(n_853), .Y(n_956) );
OAI33xp33_ASAP7_75t_L g957 ( .A1(n_796), .A2(n_837), .A3(n_795), .B1(n_799), .B2(n_790), .B3(n_850), .Y(n_957) );
AND2x2_ASAP7_75t_L g958 ( .A(n_834), .B(n_784), .Y(n_958) );
INVx2_ASAP7_75t_L g959 ( .A(n_778), .Y(n_959) );
INVx4_ASAP7_75t_L g960 ( .A(n_909), .Y(n_960) );
AOI221xp5_ASAP7_75t_L g961 ( .A1(n_832), .A2(n_796), .B1(n_851), .B2(n_837), .C(n_795), .Y(n_961) );
INVxp67_ASAP7_75t_L g962 ( .A(n_824), .Y(n_962) );
AOI221xp5_ASAP7_75t_L g963 ( .A1(n_825), .A2(n_801), .B1(n_799), .B2(n_790), .C(n_850), .Y(n_963) );
AND2x4_ASAP7_75t_L g964 ( .A(n_912), .B(n_840), .Y(n_964) );
AOI221x1_ASAP7_75t_SL g965 ( .A1(n_786), .A2(n_802), .B1(n_805), .B2(n_858), .C(n_854), .Y(n_965) );
AO22x1_ASAP7_75t_L g966 ( .A1(n_869), .A2(n_862), .B1(n_852), .B2(n_838), .Y(n_966) );
AND2x2_ASAP7_75t_L g967 ( .A(n_784), .B(n_846), .Y(n_967) );
OAI22xp33_ASAP7_75t_L g968 ( .A1(n_912), .A2(n_888), .B1(n_840), .B2(n_870), .Y(n_968) );
OAI211xp5_ASAP7_75t_L g969 ( .A1(n_774), .A2(n_859), .B(n_815), .C(n_836), .Y(n_969) );
OAI21xp5_ASAP7_75t_L g970 ( .A1(n_791), .A2(n_870), .B(n_818), .Y(n_970) );
AOI211xp5_ASAP7_75t_L g971 ( .A1(n_801), .A2(n_816), .B(n_852), .C(n_862), .Y(n_971) );
INVx2_ASAP7_75t_L g972 ( .A(n_828), .Y(n_972) );
AOI22xp33_ASAP7_75t_L g973 ( .A1(n_811), .A2(n_876), .B1(n_846), .B2(n_917), .Y(n_973) );
AND2x2_ASAP7_75t_L g974 ( .A(n_829), .B(n_792), .Y(n_974) );
AOI22xp33_ASAP7_75t_L g975 ( .A1(n_912), .A2(n_825), .B1(n_818), .B2(n_857), .Y(n_975) );
AND2x2_ASAP7_75t_L g976 ( .A(n_792), .B(n_825), .Y(n_976) );
NAND2xp5_ASAP7_75t_L g977 ( .A(n_842), .B(n_844), .Y(n_977) );
NAND2xp5_ASAP7_75t_L g978 ( .A(n_848), .B(n_864), .Y(n_978) );
BUFx4f_ASAP7_75t_L g979 ( .A(n_794), .Y(n_979) );
HB1xp67_ASAP7_75t_L g980 ( .A(n_882), .Y(n_980) );
INVx1_ASAP7_75t_L g981 ( .A(n_845), .Y(n_981) );
INVx1_ASAP7_75t_L g982 ( .A(n_845), .Y(n_982) );
HB1xp67_ASAP7_75t_L g983 ( .A(n_882), .Y(n_983) );
AOI21xp5_ASAP7_75t_L g984 ( .A1(n_880), .A2(n_777), .B(n_916), .Y(n_984) );
INVx1_ASAP7_75t_L g985 ( .A(n_849), .Y(n_985) );
OR2x6_ASAP7_75t_L g986 ( .A(n_794), .B(n_812), .Y(n_986) );
AOI22xp33_ASAP7_75t_L g987 ( .A1(n_849), .A2(n_857), .B1(n_910), .B2(n_783), .Y(n_987) );
INVx1_ASAP7_75t_L g988 ( .A(n_903), .Y(n_988) );
INVx2_ASAP7_75t_L g989 ( .A(n_872), .Y(n_989) );
INVx1_ASAP7_75t_L g990 ( .A(n_808), .Y(n_990) );
OAI221xp5_ASAP7_75t_L g991 ( .A1(n_841), .A2(n_860), .B1(n_871), .B2(n_889), .C(n_900), .Y(n_991) );
CKINVDCx8_ASAP7_75t_R g992 ( .A(n_813), .Y(n_992) );
AND2x2_ASAP7_75t_L g993 ( .A(n_922), .B(n_874), .Y(n_993) );
AOI22xp33_ASAP7_75t_L g994 ( .A1(n_900), .A2(n_879), .B1(n_874), .B2(n_919), .Y(n_994) );
AND2x2_ASAP7_75t_L g995 ( .A(n_918), .B(n_884), .Y(n_995) );
INVx1_ASAP7_75t_L g996 ( .A(n_808), .Y(n_996) );
AOI22xp33_ASAP7_75t_L g997 ( .A1(n_901), .A2(n_889), .B1(n_812), .B2(n_839), .Y(n_997) );
INVx2_ASAP7_75t_SL g998 ( .A(n_813), .Y(n_998) );
OAI33xp33_ASAP7_75t_L g999 ( .A1(n_899), .A2(n_820), .A3(n_916), .B1(n_808), .B2(n_877), .B3(n_894), .Y(n_999) );
INVx1_ASAP7_75t_L g1000 ( .A(n_820), .Y(n_1000) );
AND2x4_ASAP7_75t_L g1001 ( .A(n_866), .B(n_883), .Y(n_1001) );
CKINVDCx5p33_ASAP7_75t_R g1002 ( .A(n_875), .Y(n_1002) );
AOI22xp33_ASAP7_75t_L g1003 ( .A1(n_920), .A2(n_883), .B1(n_911), .B2(n_904), .Y(n_1003) );
INVx1_ASAP7_75t_L g1004 ( .A(n_820), .Y(n_1004) );
CKINVDCx20_ASAP7_75t_R g1005 ( .A(n_920), .Y(n_1005) );
A2O1A1Ixp33_ASAP7_75t_L g1006 ( .A1(n_904), .A2(n_905), .B(n_804), .C(n_793), .Y(n_1006) );
INVx2_ASAP7_75t_L g1007 ( .A(n_913), .Y(n_1007) );
OAI22xp33_ASAP7_75t_L g1008 ( .A1(n_899), .A2(n_905), .B1(n_866), .B2(n_883), .Y(n_1008) );
OAI21xp33_ASAP7_75t_L g1009 ( .A1(n_892), .A2(n_885), .B(n_908), .Y(n_1009) );
HB1xp67_ASAP7_75t_L g1010 ( .A(n_911), .Y(n_1010) );
INVx2_ASAP7_75t_L g1011 ( .A(n_913), .Y(n_1011) );
HB1xp67_ASAP7_75t_L g1012 ( .A(n_911), .Y(n_1012) );
INVx1_ASAP7_75t_L g1013 ( .A(n_894), .Y(n_1013) );
AO22x1_ASAP7_75t_L g1014 ( .A1(n_866), .A2(n_898), .B1(n_886), .B2(n_897), .Y(n_1014) );
OAI211xp5_ASAP7_75t_L g1015 ( .A1(n_804), .A2(n_906), .B(n_921), .C(n_914), .Y(n_1015) );
AOI221xp5_ASAP7_75t_L g1016 ( .A1(n_819), .A2(n_881), .B1(n_907), .B2(n_886), .C(n_898), .Y(n_1016) );
INVx1_ASAP7_75t_L g1017 ( .A(n_894), .Y(n_1017) );
AND2x2_ASAP7_75t_L g1018 ( .A(n_866), .B(n_915), .Y(n_1018) );
OAI22x1_ASAP7_75t_L g1019 ( .A1(n_891), .A2(n_800), .B1(n_843), .B2(n_915), .Y(n_1019) );
AOI222xp33_ASAP7_75t_L g1020 ( .A1(n_902), .A2(n_830), .B1(n_833), .B2(n_831), .C1(n_807), .C2(n_809), .Y(n_1020) );
NAND2xp5_ASAP7_75t_L g1021 ( .A(n_787), .B(n_878), .Y(n_1021) );
A2O1A1Ixp33_ASAP7_75t_L g1022 ( .A1(n_895), .A2(n_855), .B(n_890), .C(n_856), .Y(n_1022) );
AOI22xp33_ASAP7_75t_L g1023 ( .A1(n_878), .A2(n_822), .B1(n_800), .B2(n_863), .Y(n_1023) );
OAI221xp5_ASAP7_75t_L g1024 ( .A1(n_822), .A2(n_631), .B1(n_671), .B2(n_779), .C(n_896), .Y(n_1024) );
OAI22xp33_ASAP7_75t_L g1025 ( .A1(n_873), .A2(n_595), .B1(n_547), .B2(n_541), .Y(n_1025) );
AOI221xp5_ASAP7_75t_L g1026 ( .A1(n_779), .A2(n_659), .B1(n_550), .B2(n_566), .C(n_551), .Y(n_1026) );
NAND2xp5_ASAP7_75t_L g1027 ( .A(n_803), .B(n_810), .Y(n_1027) );
AOI22xp33_ASAP7_75t_L g1028 ( .A1(n_779), .A2(n_595), .B1(n_543), .B2(n_559), .Y(n_1028) );
OAI21xp33_ASAP7_75t_L g1029 ( .A1(n_779), .A2(n_677), .B(n_558), .Y(n_1029) );
OAI22xp5_ASAP7_75t_L g1030 ( .A1(n_803), .A2(n_814), .B1(n_817), .B2(n_810), .Y(n_1030) );
OAI21x1_ASAP7_75t_L g1031 ( .A1(n_773), .A2(n_782), .B(n_777), .Y(n_1031) );
HB1xp67_ASAP7_75t_L g1032 ( .A(n_780), .Y(n_1032) );
AOI22xp5_ASAP7_75t_L g1033 ( .A1(n_779), .A2(n_677), .B1(n_595), .B2(n_659), .Y(n_1033) );
BUFx2_ASAP7_75t_L g1034 ( .A(n_789), .Y(n_1034) );
AOI21xp5_ASAP7_75t_L g1035 ( .A1(n_887), .A2(n_744), .B(n_652), .Y(n_1035) );
INVx2_ASAP7_75t_L g1036 ( .A(n_798), .Y(n_1036) );
AND2x4_ASAP7_75t_L g1037 ( .A(n_781), .B(n_806), .Y(n_1037) );
BUFx12f_ASAP7_75t_L g1038 ( .A(n_785), .Y(n_1038) );
OAI211xp5_ASAP7_75t_L g1039 ( .A1(n_774), .A2(n_823), .B(n_832), .C(n_697), .Y(n_1039) );
INVx1_ASAP7_75t_L g1040 ( .A(n_775), .Y(n_1040) );
AND2x4_ASAP7_75t_L g1041 ( .A(n_781), .B(n_806), .Y(n_1041) );
AOI22xp33_ASAP7_75t_L g1042 ( .A1(n_779), .A2(n_595), .B1(n_543), .B2(n_559), .Y(n_1042) );
AND2x4_ASAP7_75t_L g1043 ( .A(n_781), .B(n_806), .Y(n_1043) );
INVx1_ASAP7_75t_L g1044 ( .A(n_775), .Y(n_1044) );
AOI22xp33_ASAP7_75t_L g1045 ( .A1(n_779), .A2(n_595), .B1(n_543), .B2(n_559), .Y(n_1045) );
NAND2xp5_ASAP7_75t_L g1046 ( .A(n_803), .B(n_810), .Y(n_1046) );
INVx1_ASAP7_75t_L g1047 ( .A(n_775), .Y(n_1047) );
INVx1_ASAP7_75t_L g1048 ( .A(n_775), .Y(n_1048) );
INVx3_ASAP7_75t_L g1049 ( .A(n_781), .Y(n_1049) );
NAND2xp5_ASAP7_75t_L g1050 ( .A(n_803), .B(n_810), .Y(n_1050) );
NOR2xp33_ASAP7_75t_L g1051 ( .A(n_779), .B(n_686), .Y(n_1051) );
BUFx3_ASAP7_75t_L g1052 ( .A(n_954), .Y(n_1052) );
BUFx6f_ASAP7_75t_L g1053 ( .A(n_986), .Y(n_1053) );
NAND2xp5_ASAP7_75t_L g1054 ( .A(n_1026), .B(n_1051), .Y(n_1054) );
OR2x2_ASAP7_75t_L g1055 ( .A(n_1030), .B(n_1027), .Y(n_1055) );
INVx1_ASAP7_75t_L g1056 ( .A(n_990), .Y(n_1056) );
INVx3_ASAP7_75t_L g1057 ( .A(n_979), .Y(n_1057) );
INVx1_ASAP7_75t_L g1058 ( .A(n_996), .Y(n_1058) );
INVx4_ASAP7_75t_L g1059 ( .A(n_979), .Y(n_1059) );
INVx1_ASAP7_75t_L g1060 ( .A(n_943), .Y(n_1060) );
INVx1_ASAP7_75t_SL g1061 ( .A(n_1034), .Y(n_1061) );
INVx2_ASAP7_75t_L g1062 ( .A(n_1027), .Y(n_1062) );
OR2x2_ASAP7_75t_L g1063 ( .A(n_1030), .B(n_1050), .Y(n_1063) );
INVxp67_ASAP7_75t_SL g1064 ( .A(n_1046), .Y(n_1064) );
AND2x2_ASAP7_75t_L g1065 ( .A(n_1046), .B(n_1050), .Y(n_1065) );
AND2x2_ASAP7_75t_L g1066 ( .A(n_959), .B(n_926), .Y(n_1066) );
INVxp67_ASAP7_75t_L g1067 ( .A(n_933), .Y(n_1067) );
OR2x2_ASAP7_75t_L g1068 ( .A(n_964), .B(n_978), .Y(n_1068) );
NAND2xp5_ASAP7_75t_L g1069 ( .A(n_923), .B(n_934), .Y(n_1069) );
INVx3_ASAP7_75t_L g1070 ( .A(n_986), .Y(n_1070) );
INVx1_ASAP7_75t_L g1071 ( .A(n_1000), .Y(n_1071) );
NAND2xp5_ASAP7_75t_L g1072 ( .A(n_1040), .B(n_1044), .Y(n_1072) );
INVx2_ASAP7_75t_L g1073 ( .A(n_978), .Y(n_1073) );
INVx1_ASAP7_75t_L g1074 ( .A(n_951), .Y(n_1074) );
INVx2_ASAP7_75t_L g1075 ( .A(n_955), .Y(n_1075) );
INVx1_ASAP7_75t_L g1076 ( .A(n_1047), .Y(n_1076) );
AND2x2_ASAP7_75t_L g1077 ( .A(n_942), .B(n_945), .Y(n_1077) );
NOR2x1_ASAP7_75t_L g1078 ( .A(n_960), .B(n_1005), .Y(n_1078) );
AND2x2_ASAP7_75t_L g1079 ( .A(n_1036), .B(n_972), .Y(n_1079) );
HB1xp67_ASAP7_75t_L g1080 ( .A(n_1032), .Y(n_1080) );
INVx1_ASAP7_75t_L g1081 ( .A(n_1004), .Y(n_1081) );
INVx1_ASAP7_75t_L g1082 ( .A(n_977), .Y(n_1082) );
BUFx3_ASAP7_75t_L g1083 ( .A(n_954), .Y(n_1083) );
INVx1_ASAP7_75t_L g1084 ( .A(n_977), .Y(n_1084) );
BUFx3_ASAP7_75t_L g1085 ( .A(n_954), .Y(n_1085) );
INVx1_ASAP7_75t_L g1086 ( .A(n_1048), .Y(n_1086) );
INVx1_ASAP7_75t_L g1087 ( .A(n_1013), .Y(n_1087) );
INVx3_ASAP7_75t_L g1088 ( .A(n_986), .Y(n_1088) );
INVx2_ASAP7_75t_L g1089 ( .A(n_989), .Y(n_1089) );
HB1xp67_ASAP7_75t_L g1090 ( .A(n_974), .Y(n_1090) );
AOI322xp5_ASAP7_75t_L g1091 ( .A1(n_1028), .A2(n_1042), .A3(n_1045), .B1(n_1025), .B2(n_1033), .C1(n_976), .C2(n_961), .Y(n_1091) );
AND2x2_ASAP7_75t_L g1092 ( .A(n_995), .B(n_964), .Y(n_1092) );
INVx1_ASAP7_75t_L g1093 ( .A(n_1017), .Y(n_1093) );
INVx1_ASAP7_75t_L g1094 ( .A(n_981), .Y(n_1094) );
HB1xp67_ASAP7_75t_L g1095 ( .A(n_936), .Y(n_1095) );
AND2x2_ASAP7_75t_L g1096 ( .A(n_982), .B(n_985), .Y(n_1096) );
AND2x2_ASAP7_75t_L g1097 ( .A(n_988), .B(n_929), .Y(n_1097) );
INVx2_ASAP7_75t_SL g1098 ( .A(n_928), .Y(n_1098) );
INVx2_ASAP7_75t_L g1099 ( .A(n_927), .Y(n_1099) );
INVx4_ASAP7_75t_R g1100 ( .A(n_998), .Y(n_1100) );
NOR2x1_ASAP7_75t_SL g1101 ( .A(n_950), .B(n_947), .Y(n_1101) );
INVx2_ASAP7_75t_SL g1102 ( .A(n_928), .Y(n_1102) );
NAND2xp5_ASAP7_75t_L g1103 ( .A(n_1029), .B(n_958), .Y(n_1103) );
BUFx2_ASAP7_75t_L g1104 ( .A(n_980), .Y(n_1104) );
NAND2xp5_ASAP7_75t_L g1105 ( .A(n_1039), .B(n_973), .Y(n_1105) );
INVx1_ASAP7_75t_L g1106 ( .A(n_935), .Y(n_1106) );
AOI22xp5_ASAP7_75t_L g1107 ( .A1(n_961), .A2(n_968), .B1(n_1024), .B2(n_969), .Y(n_1107) );
CKINVDCx6p67_ASAP7_75t_R g1108 ( .A(n_960), .Y(n_1108) );
AND2x4_ASAP7_75t_L g1109 ( .A(n_1001), .B(n_937), .Y(n_1109) );
AND2x4_ASAP7_75t_SL g1110 ( .A(n_1037), .B(n_1041), .Y(n_1110) );
OR2x2_ASAP7_75t_L g1111 ( .A(n_975), .B(n_983), .Y(n_1111) );
AND2x4_ASAP7_75t_L g1112 ( .A(n_937), .B(n_1018), .Y(n_1112) );
INVxp67_ASAP7_75t_SL g1113 ( .A(n_1010), .Y(n_1113) );
BUFx3_ASAP7_75t_L g1114 ( .A(n_1037), .Y(n_1114) );
INVx3_ASAP7_75t_L g1115 ( .A(n_1041), .Y(n_1115) );
INVx1_ASAP7_75t_L g1116 ( .A(n_970), .Y(n_1116) );
INVx1_ASAP7_75t_L g1117 ( .A(n_952), .Y(n_1117) );
AND2x2_ASAP7_75t_L g1118 ( .A(n_939), .B(n_967), .Y(n_1118) );
INVx2_ASAP7_75t_SL g1119 ( .A(n_1043), .Y(n_1119) );
INVx2_ASAP7_75t_L g1120 ( .A(n_1007), .Y(n_1120) );
INVx2_ASAP7_75t_L g1121 ( .A(n_1011), .Y(n_1121) );
AO21x2_ASAP7_75t_L g1122 ( .A1(n_984), .A2(n_1006), .B(n_1008), .Y(n_1122) );
AND2x2_ASAP7_75t_L g1123 ( .A(n_1012), .B(n_987), .Y(n_1123) );
AOI22xp33_ASAP7_75t_L g1124 ( .A1(n_957), .A2(n_1024), .B1(n_963), .B2(n_944), .Y(n_1124) );
INVx1_ASAP7_75t_L g1125 ( .A(n_1049), .Y(n_1125) );
BUFx2_ASAP7_75t_L g1126 ( .A(n_1021), .Y(n_1126) );
NAND2xp5_ASAP7_75t_L g1127 ( .A(n_1043), .B(n_965), .Y(n_1127) );
INVx1_ASAP7_75t_L g1128 ( .A(n_938), .Y(n_1128) );
AND2x2_ASAP7_75t_L g1129 ( .A(n_971), .B(n_993), .Y(n_1129) );
INVx1_ASAP7_75t_L g1130 ( .A(n_938), .Y(n_1130) );
HB1xp67_ASAP7_75t_L g1131 ( .A(n_1049), .Y(n_1131) );
NAND2xp5_ASAP7_75t_L g1132 ( .A(n_965), .B(n_963), .Y(n_1132) );
INVx1_ASAP7_75t_L g1133 ( .A(n_1021), .Y(n_1133) );
INVx1_ASAP7_75t_L g1134 ( .A(n_966), .Y(n_1134) );
AND2x2_ASAP7_75t_L g1135 ( .A(n_994), .B(n_949), .Y(n_1135) );
OR2x2_ASAP7_75t_L g1136 ( .A(n_956), .B(n_930), .Y(n_1136) );
AND2x2_ASAP7_75t_L g1137 ( .A(n_924), .B(n_1035), .Y(n_1137) );
AND2x2_ASAP7_75t_L g1138 ( .A(n_924), .B(n_941), .Y(n_1138) );
BUFx2_ASAP7_75t_L g1139 ( .A(n_1014), .Y(n_1139) );
AND2x4_ASAP7_75t_L g1140 ( .A(n_925), .B(n_931), .Y(n_1140) );
AND2x4_ASAP7_75t_L g1141 ( .A(n_997), .B(n_953), .Y(n_1141) );
INVx1_ASAP7_75t_L g1142 ( .A(n_950), .Y(n_1142) );
CKINVDCx5p33_ASAP7_75t_R g1143 ( .A(n_992), .Y(n_1143) );
OAI33xp33_ASAP7_75t_L g1144 ( .A1(n_1132), .A2(n_962), .A3(n_946), .B1(n_1002), .B2(n_1009), .B3(n_999), .Y(n_1144) );
AND2x2_ASAP7_75t_L g1145 ( .A(n_1065), .B(n_1003), .Y(n_1145) );
OR2x2_ASAP7_75t_L g1146 ( .A(n_1055), .B(n_940), .Y(n_1146) );
NAND2xp5_ASAP7_75t_L g1147 ( .A(n_1065), .B(n_991), .Y(n_1147) );
INVx1_ASAP7_75t_L g1148 ( .A(n_1056), .Y(n_1148) );
NAND2xp5_ASAP7_75t_L g1149 ( .A(n_1096), .B(n_991), .Y(n_1149) );
INVx1_ASAP7_75t_L g1150 ( .A(n_1056), .Y(n_1150) );
AOI22xp33_ASAP7_75t_L g1151 ( .A1(n_1136), .A2(n_940), .B1(n_948), .B2(n_1016), .Y(n_1151) );
INVx1_ASAP7_75t_L g1152 ( .A(n_1058), .Y(n_1152) );
AND2x4_ASAP7_75t_L g1153 ( .A(n_1112), .B(n_1022), .Y(n_1153) );
INVx1_ASAP7_75t_L g1154 ( .A(n_1058), .Y(n_1154) );
INVx1_ASAP7_75t_L g1155 ( .A(n_1071), .Y(n_1155) );
NAND2xp5_ASAP7_75t_L g1156 ( .A(n_1096), .B(n_932), .Y(n_1156) );
OR2x6_ASAP7_75t_L g1157 ( .A(n_1139), .B(n_1019), .Y(n_1157) );
INVx1_ASAP7_75t_L g1158 ( .A(n_1081), .Y(n_1158) );
AND2x2_ASAP7_75t_L g1159 ( .A(n_1062), .B(n_1023), .Y(n_1159) );
AND2x2_ASAP7_75t_SL g1160 ( .A(n_1055), .B(n_1020), .Y(n_1160) );
INVx1_ASAP7_75t_SL g1161 ( .A(n_1108), .Y(n_1161) );
INVx1_ASAP7_75t_L g1162 ( .A(n_1087), .Y(n_1162) );
AOI22xp33_ASAP7_75t_L g1163 ( .A1(n_1136), .A2(n_1038), .B1(n_1020), .B2(n_1031), .Y(n_1163) );
NAND2xp5_ASAP7_75t_L g1164 ( .A(n_1105), .B(n_1015), .Y(n_1164) );
NOR2x1_ASAP7_75t_L g1165 ( .A(n_1139), .B(n_1070), .Y(n_1165) );
AND2x2_ASAP7_75t_L g1166 ( .A(n_1073), .B(n_1129), .Y(n_1166) );
INVx1_ASAP7_75t_L g1167 ( .A(n_1087), .Y(n_1167) );
AND2x2_ASAP7_75t_L g1168 ( .A(n_1073), .B(n_1129), .Y(n_1168) );
INVx1_ASAP7_75t_L g1169 ( .A(n_1093), .Y(n_1169) );
OAI33xp33_ASAP7_75t_L g1170 ( .A1(n_1127), .A2(n_1067), .A3(n_1054), .B1(n_1103), .B2(n_1074), .B3(n_1060), .Y(n_1170) );
AOI22xp33_ASAP7_75t_L g1171 ( .A1(n_1107), .A2(n_1138), .B1(n_1135), .B2(n_1118), .Y(n_1171) );
BUFx6f_ASAP7_75t_L g1172 ( .A(n_1140), .Y(n_1172) );
BUFx2_ASAP7_75t_L g1173 ( .A(n_1126), .Y(n_1173) );
INVxp67_ASAP7_75t_SL g1174 ( .A(n_1064), .Y(n_1174) );
HB1xp67_ASAP7_75t_L g1175 ( .A(n_1080), .Y(n_1175) );
AND2x2_ASAP7_75t_L g1176 ( .A(n_1092), .B(n_1133), .Y(n_1176) );
INVx1_ASAP7_75t_L g1177 ( .A(n_1116), .Y(n_1177) );
AOI221xp5_ASAP7_75t_L g1178 ( .A1(n_1124), .A2(n_1094), .B1(n_1076), .B2(n_1097), .C(n_1086), .Y(n_1178) );
INVx2_ASAP7_75t_L g1179 ( .A(n_1099), .Y(n_1179) );
OAI21xp5_ASAP7_75t_SL g1180 ( .A1(n_1110), .A2(n_1078), .B(n_1057), .Y(n_1180) );
BUFx3_ASAP7_75t_L g1181 ( .A(n_1114), .Y(n_1181) );
BUFx10_ASAP7_75t_L g1182 ( .A(n_1143), .Y(n_1182) );
AOI221xp5_ASAP7_75t_L g1183 ( .A1(n_1094), .A2(n_1097), .B1(n_1086), .B2(n_1072), .C(n_1069), .Y(n_1183) );
OR2x2_ASAP7_75t_L g1184 ( .A(n_1063), .B(n_1111), .Y(n_1184) );
INVxp67_ASAP7_75t_L g1185 ( .A(n_1090), .Y(n_1185) );
NAND3xp33_ASAP7_75t_L g1186 ( .A(n_1091), .B(n_1134), .C(n_1131), .Y(n_1186) );
INVx1_ASAP7_75t_L g1187 ( .A(n_1120), .Y(n_1187) );
AND2x2_ASAP7_75t_L g1188 ( .A(n_1075), .B(n_1079), .Y(n_1188) );
INVx5_ASAP7_75t_L g1189 ( .A(n_1053), .Y(n_1189) );
INVx1_ASAP7_75t_L g1190 ( .A(n_1121), .Y(n_1190) );
OAI211xp5_ASAP7_75t_L g1191 ( .A1(n_1134), .A2(n_1059), .B(n_1061), .C(n_1095), .Y(n_1191) );
AND2x2_ASAP7_75t_L g1192 ( .A(n_1066), .B(n_1077), .Y(n_1192) );
AND2x2_ASAP7_75t_L g1193 ( .A(n_1066), .B(n_1077), .Y(n_1193) );
INVx1_ASAP7_75t_L g1194 ( .A(n_1148), .Y(n_1194) );
AND2x2_ASAP7_75t_L g1195 ( .A(n_1166), .B(n_1137), .Y(n_1195) );
INVx2_ASAP7_75t_L g1196 ( .A(n_1179), .Y(n_1196) );
INVx1_ASAP7_75t_L g1197 ( .A(n_1175), .Y(n_1197) );
BUFx3_ASAP7_75t_L g1198 ( .A(n_1181), .Y(n_1198) );
NAND2xp5_ASAP7_75t_L g1199 ( .A(n_1192), .B(n_1082), .Y(n_1199) );
INVx1_ASAP7_75t_L g1200 ( .A(n_1150), .Y(n_1200) );
AND2x2_ASAP7_75t_L g1201 ( .A(n_1166), .B(n_1137), .Y(n_1201) );
BUFx2_ASAP7_75t_L g1202 ( .A(n_1174), .Y(n_1202) );
BUFx3_ASAP7_75t_L g1203 ( .A(n_1181), .Y(n_1203) );
AND2x2_ASAP7_75t_L g1204 ( .A(n_1168), .B(n_1122), .Y(n_1204) );
AOI221xp5_ASAP7_75t_L g1205 ( .A1(n_1170), .A2(n_1123), .B1(n_1084), .B2(n_1104), .C(n_1106), .Y(n_1205) );
AND2x2_ASAP7_75t_L g1206 ( .A(n_1168), .B(n_1122), .Y(n_1206) );
INVx1_ASAP7_75t_L g1207 ( .A(n_1152), .Y(n_1207) );
CKINVDCx20_ASAP7_75t_R g1208 ( .A(n_1161), .Y(n_1208) );
OR2x2_ASAP7_75t_L g1209 ( .A(n_1184), .B(n_1068), .Y(n_1209) );
INVx1_ASAP7_75t_L g1210 ( .A(n_1154), .Y(n_1210) );
NAND2xp5_ASAP7_75t_L g1211 ( .A(n_1193), .B(n_1106), .Y(n_1211) );
AOI22xp33_ASAP7_75t_L g1212 ( .A1(n_1160), .A2(n_1135), .B1(n_1142), .B2(n_1118), .Y(n_1212) );
AND2x4_ASAP7_75t_L g1213 ( .A(n_1153), .B(n_1109), .Y(n_1213) );
AND2x2_ASAP7_75t_L g1214 ( .A(n_1155), .B(n_1123), .Y(n_1214) );
NOR2xp33_ASAP7_75t_L g1215 ( .A(n_1156), .B(n_1108), .Y(n_1215) );
INVx3_ASAP7_75t_SL g1216 ( .A(n_1189), .Y(n_1216) );
INVx1_ASAP7_75t_L g1217 ( .A(n_1155), .Y(n_1217) );
HB1xp67_ASAP7_75t_L g1218 ( .A(n_1173), .Y(n_1218) );
NAND2xp67_ASAP7_75t_L g1219 ( .A(n_1188), .B(n_1089), .Y(n_1219) );
INVx1_ASAP7_75t_L g1220 ( .A(n_1158), .Y(n_1220) );
INVx1_ASAP7_75t_L g1221 ( .A(n_1158), .Y(n_1221) );
OR2x2_ASAP7_75t_L g1222 ( .A(n_1173), .B(n_1126), .Y(n_1222) );
AND2x4_ASAP7_75t_L g1223 ( .A(n_1153), .B(n_1172), .Y(n_1223) );
INVx1_ASAP7_75t_L g1224 ( .A(n_1162), .Y(n_1224) );
OR2x2_ASAP7_75t_L g1225 ( .A(n_1146), .B(n_1113), .Y(n_1225) );
OR2x2_ASAP7_75t_L g1226 ( .A(n_1146), .B(n_1089), .Y(n_1226) );
INVx1_ASAP7_75t_L g1227 ( .A(n_1162), .Y(n_1227) );
OR2x2_ASAP7_75t_L g1228 ( .A(n_1167), .B(n_1117), .Y(n_1228) );
INVxp67_ASAP7_75t_SL g1229 ( .A(n_1185), .Y(n_1229) );
INVx2_ASAP7_75t_L g1230 ( .A(n_1196), .Y(n_1230) );
AND2x2_ASAP7_75t_SL g1231 ( .A(n_1202), .B(n_1160), .Y(n_1231) );
INVx1_ASAP7_75t_L g1232 ( .A(n_1194), .Y(n_1232) );
NAND4xp25_ASAP7_75t_L g1233 ( .A(n_1212), .B(n_1171), .C(n_1163), .D(n_1186), .Y(n_1233) );
INVx1_ASAP7_75t_L g1234 ( .A(n_1194), .Y(n_1234) );
AOI22xp33_ASAP7_75t_L g1235 ( .A1(n_1197), .A2(n_1144), .B1(n_1147), .B2(n_1149), .Y(n_1235) );
NAND2xp5_ASAP7_75t_L g1236 ( .A(n_1195), .B(n_1183), .Y(n_1236) );
NAND2xp5_ASAP7_75t_L g1237 ( .A(n_1195), .B(n_1176), .Y(n_1237) );
INVx4_ASAP7_75t_L g1238 ( .A(n_1216), .Y(n_1238) );
NAND2x1_ASAP7_75t_L g1239 ( .A(n_1202), .B(n_1165), .Y(n_1239) );
NAND2xp5_ASAP7_75t_L g1240 ( .A(n_1201), .B(n_1176), .Y(n_1240) );
NOR2xp33_ASAP7_75t_L g1241 ( .A(n_1229), .B(n_1164), .Y(n_1241) );
OR2x2_ASAP7_75t_L g1242 ( .A(n_1209), .B(n_1187), .Y(n_1242) );
OR2x2_ASAP7_75t_L g1243 ( .A(n_1209), .B(n_1187), .Y(n_1243) );
NAND2xp5_ASAP7_75t_L g1244 ( .A(n_1201), .B(n_1178), .Y(n_1244) );
INVx1_ASAP7_75t_L g1245 ( .A(n_1200), .Y(n_1245) );
AND2x2_ASAP7_75t_L g1246 ( .A(n_1204), .B(n_1159), .Y(n_1246) );
NOR2xp33_ASAP7_75t_L g1247 ( .A(n_1199), .B(n_1191), .Y(n_1247) );
OR2x2_ASAP7_75t_L g1248 ( .A(n_1211), .B(n_1190), .Y(n_1248) );
AND2x2_ASAP7_75t_L g1249 ( .A(n_1204), .B(n_1169), .Y(n_1249) );
INVxp33_ASAP7_75t_L g1250 ( .A(n_1218), .Y(n_1250) );
NAND2xp5_ASAP7_75t_L g1251 ( .A(n_1214), .B(n_1145), .Y(n_1251) );
AND2x2_ASAP7_75t_L g1252 ( .A(n_1206), .B(n_1177), .Y(n_1252) );
INVx1_ASAP7_75t_L g1253 ( .A(n_1207), .Y(n_1253) );
INVx1_ASAP7_75t_L g1254 ( .A(n_1207), .Y(n_1254) );
INVx3_ASAP7_75t_SL g1255 ( .A(n_1208), .Y(n_1255) );
INVx1_ASAP7_75t_L g1256 ( .A(n_1210), .Y(n_1256) );
INVx1_ASAP7_75t_L g1257 ( .A(n_1210), .Y(n_1257) );
AND2x2_ASAP7_75t_L g1258 ( .A(n_1246), .B(n_1206), .Y(n_1258) );
OAI22xp33_ASAP7_75t_L g1259 ( .A1(n_1238), .A2(n_1216), .B1(n_1180), .B2(n_1208), .Y(n_1259) );
AOI22xp5_ASAP7_75t_L g1260 ( .A1(n_1233), .A2(n_1247), .B1(n_1231), .B2(n_1241), .Y(n_1260) );
NAND2xp5_ASAP7_75t_L g1261 ( .A(n_1249), .B(n_1236), .Y(n_1261) );
NAND2xp5_ASAP7_75t_L g1262 ( .A(n_1249), .B(n_1205), .Y(n_1262) );
NAND2xp5_ASAP7_75t_L g1263 ( .A(n_1244), .B(n_1252), .Y(n_1263) );
NAND2xp5_ASAP7_75t_SL g1264 ( .A(n_1238), .B(n_1198), .Y(n_1264) );
AOI22xp33_ASAP7_75t_L g1265 ( .A1(n_1241), .A2(n_1225), .B1(n_1215), .B2(n_1213), .Y(n_1265) );
INVx1_ASAP7_75t_L g1266 ( .A(n_1232), .Y(n_1266) );
INVx2_ASAP7_75t_SL g1267 ( .A(n_1238), .Y(n_1267) );
INVx2_ASAP7_75t_L g1268 ( .A(n_1230), .Y(n_1268) );
INVx1_ASAP7_75t_SL g1269 ( .A(n_1255), .Y(n_1269) );
OAI22x1_ASAP7_75t_L g1270 ( .A1(n_1255), .A2(n_1165), .B1(n_1213), .B2(n_1222), .Y(n_1270) );
INVx1_ASAP7_75t_L g1271 ( .A(n_1234), .Y(n_1271) );
INVx2_ASAP7_75t_L g1272 ( .A(n_1230), .Y(n_1272) );
AOI322xp5_ASAP7_75t_L g1273 ( .A1(n_1235), .A2(n_1151), .A3(n_1220), .B1(n_1221), .B2(n_1227), .C1(n_1217), .C2(n_1224), .Y(n_1273) );
INVx1_ASAP7_75t_L g1274 ( .A(n_1266), .Y(n_1274) );
NAND2x1_ASAP7_75t_SL g1275 ( .A(n_1260), .B(n_1059), .Y(n_1275) );
O2A1O1Ixp33_ASAP7_75t_SL g1276 ( .A1(n_1264), .A2(n_1239), .B(n_1219), .C(n_1250), .Y(n_1276) );
OAI322xp33_ASAP7_75t_L g1277 ( .A1(n_1262), .A2(n_1240), .A3(n_1237), .B1(n_1251), .B2(n_1248), .C1(n_1242), .C2(n_1243), .Y(n_1277) );
XNOR2x1_ASAP7_75t_L g1278 ( .A(n_1269), .B(n_1143), .Y(n_1278) );
INVx1_ASAP7_75t_L g1279 ( .A(n_1271), .Y(n_1279) );
AND2x2_ASAP7_75t_L g1280 ( .A(n_1258), .B(n_1223), .Y(n_1280) );
AOI221xp5_ASAP7_75t_L g1281 ( .A1(n_1265), .A2(n_1257), .B1(n_1256), .B2(n_1254), .C(n_1253), .Y(n_1281) );
INVx2_ASAP7_75t_L g1282 ( .A(n_1268), .Y(n_1282) );
NAND2xp5_ASAP7_75t_L g1283 ( .A(n_1263), .B(n_1245), .Y(n_1283) );
INVxp67_ASAP7_75t_SL g1284 ( .A(n_1268), .Y(n_1284) );
INVx1_ASAP7_75t_SL g1285 ( .A(n_1267), .Y(n_1285) );
NOR2xp33_ASAP7_75t_L g1286 ( .A(n_1261), .B(n_1198), .Y(n_1286) );
OAI211xp5_ASAP7_75t_L g1287 ( .A1(n_1273), .A2(n_1059), .B(n_1203), .C(n_1114), .Y(n_1287) );
NAND2x1p5_ASAP7_75t_L g1288 ( .A(n_1285), .B(n_1267), .Y(n_1288) );
INVx1_ASAP7_75t_L g1289 ( .A(n_1274), .Y(n_1289) );
INVx1_ASAP7_75t_L g1290 ( .A(n_1279), .Y(n_1290) );
NOR2x1_ASAP7_75t_L g1291 ( .A(n_1287), .B(n_1259), .Y(n_1291) );
NOR3xp33_ASAP7_75t_L g1292 ( .A(n_1281), .B(n_1115), .C(n_1088), .Y(n_1292) );
OAI21xp5_ASAP7_75t_SL g1293 ( .A1(n_1278), .A2(n_1057), .B(n_1115), .Y(n_1293) );
A2O1A1Ixp33_ASAP7_75t_L g1294 ( .A1(n_1275), .A2(n_1203), .B(n_1057), .C(n_1088), .Y(n_1294) );
INVx1_ASAP7_75t_L g1295 ( .A(n_1283), .Y(n_1295) );
AOI211xp5_ASAP7_75t_SL g1296 ( .A1(n_1293), .A2(n_1276), .B(n_1277), .C(n_1286), .Y(n_1296) );
CKINVDCx6p67_ASAP7_75t_R g1297 ( .A(n_1288), .Y(n_1297) );
OAI221xp5_ASAP7_75t_SL g1298 ( .A1(n_1294), .A2(n_1284), .B1(n_1280), .B2(n_1157), .C(n_1226), .Y(n_1298) );
AOI222xp33_ASAP7_75t_L g1299 ( .A1(n_1291), .A2(n_1270), .B1(n_1282), .B2(n_1182), .C1(n_1272), .C2(n_1227), .Y(n_1299) );
OAI221xp5_ASAP7_75t_SL g1300 ( .A1(n_1292), .A2(n_1157), .B1(n_1102), .B2(n_1098), .C(n_1119), .Y(n_1300) );
OAI221xp5_ASAP7_75t_SL g1301 ( .A1(n_1295), .A2(n_1157), .B1(n_1119), .B2(n_1098), .C(n_1228), .Y(n_1301) );
AND2x2_ASAP7_75t_L g1302 ( .A(n_1297), .B(n_1290), .Y(n_1302) );
HB1xp67_ASAP7_75t_L g1303 ( .A(n_1296), .Y(n_1303) );
AND2x2_ASAP7_75t_L g1304 ( .A(n_1299), .B(n_1289), .Y(n_1304) );
NOR3xp33_ASAP7_75t_L g1305 ( .A(n_1298), .B(n_1052), .C(n_1083), .Y(n_1305) );
OR4x2_ASAP7_75t_L g1306 ( .A(n_1303), .B(n_1300), .C(n_1301), .D(n_1100), .Y(n_1306) );
BUFx6f_ASAP7_75t_L g1307 ( .A(n_1302), .Y(n_1307) );
NOR3xp33_ASAP7_75t_L g1308 ( .A(n_1304), .B(n_1301), .C(n_1085), .Y(n_1308) );
CKINVDCx20_ASAP7_75t_R g1309 ( .A(n_1307), .Y(n_1309) );
HB1xp67_ASAP7_75t_L g1310 ( .A(n_1307), .Y(n_1310) );
INVx1_ASAP7_75t_L g1311 ( .A(n_1310), .Y(n_1311) );
XNOR2xp5_ASAP7_75t_L g1312 ( .A(n_1309), .B(n_1308), .Y(n_1312) );
OAI22xp5_ASAP7_75t_SL g1313 ( .A1(n_1309), .A2(n_1306), .B1(n_1305), .B2(n_1157), .Y(n_1313) );
INVx1_ASAP7_75t_SL g1314 ( .A(n_1311), .Y(n_1314) );
HB1xp67_ASAP7_75t_L g1315 ( .A(n_1312), .Y(n_1315) );
INVx1_ASAP7_75t_L g1316 ( .A(n_1313), .Y(n_1316) );
AOI222xp33_ASAP7_75t_L g1317 ( .A1(n_1314), .A2(n_1128), .B1(n_1125), .B2(n_1130), .C1(n_1141), .C2(n_1101), .Y(n_1317) );
INVx2_ASAP7_75t_SL g1318 ( .A(n_1315), .Y(n_1318) );
OAI22xp5_ASAP7_75t_L g1319 ( .A1(n_1318), .A2(n_1316), .B1(n_1189), .B2(n_1141), .Y(n_1319) );
AOI22xp5_ASAP7_75t_L g1320 ( .A1(n_1319), .A2(n_1317), .B1(n_1223), .B2(n_1140), .Y(n_1320) );
endmodule