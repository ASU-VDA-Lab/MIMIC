module real_jpeg_15378_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_366;
wire n_456;
wire n_259;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_483;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_464;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_233;
wire n_73;
wire n_516;
wire n_348;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_288;
wire n_83;
wire n_393;
wire n_221;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_21;
wire n_476;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_195;
wire n_110;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_25;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_515;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_487;
wire n_242;
wire n_493;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_196;
wire n_375;
wire n_330;
wire n_298;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_512;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_444;
wire n_178;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_509;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

AOI21xp5_ASAP7_75t_L g18 ( 
.A1(n_0),
.A2(n_19),
.B(n_515),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g515 ( 
.A(n_0),
.B(n_516),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_1),
.B(n_61),
.Y(n_60)
);

AND2x2_ASAP7_75t_L g64 ( 
.A(n_1),
.B(n_65),
.Y(n_64)
);

AND2x2_ASAP7_75t_L g69 ( 
.A(n_1),
.B(n_70),
.Y(n_69)
);

AND2x2_ASAP7_75t_L g89 ( 
.A(n_1),
.B(n_90),
.Y(n_89)
);

AND2x2_ASAP7_75t_L g92 ( 
.A(n_1),
.B(n_93),
.Y(n_92)
);

AND2x2_ASAP7_75t_L g118 ( 
.A(n_1),
.B(n_119),
.Y(n_118)
);

AND2x2_ASAP7_75t_L g183 ( 
.A(n_1),
.B(n_184),
.Y(n_183)
);

AND2x2_ASAP7_75t_L g236 ( 
.A(n_1),
.B(n_237),
.Y(n_236)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_2),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_2),
.Y(n_66)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_2),
.Y(n_270)
);

BUFx3_ASAP7_75t_L g288 ( 
.A(n_2),
.Y(n_288)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_3),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g259 ( 
.A(n_3),
.Y(n_259)
);

BUFx6f_ASAP7_75t_L g423 ( 
.A(n_3),
.Y(n_423)
);

AND2x2_ASAP7_75t_L g195 ( 
.A(n_4),
.B(n_196),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_4),
.B(n_198),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_4),
.B(n_254),
.Y(n_253)
);

AND2x2_ASAP7_75t_SL g266 ( 
.A(n_4),
.B(n_267),
.Y(n_266)
);

AND2x2_ASAP7_75t_SL g289 ( 
.A(n_4),
.B(n_290),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_4),
.B(n_421),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_SL g425 ( 
.A(n_4),
.B(n_426),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_4),
.B(n_284),
.Y(n_448)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_5),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_5),
.B(n_220),
.Y(n_219)
);

AND2x2_ASAP7_75t_SL g287 ( 
.A(n_5),
.B(n_288),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_5),
.A2(n_11),
.B1(n_302),
.B2(n_304),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g439 ( 
.A(n_5),
.B(n_440),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_5),
.B(n_451),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_SL g481 ( 
.A(n_5),
.B(n_482),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_SL g262 ( 
.A(n_6),
.B(n_263),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_6),
.B(n_330),
.Y(n_329)
);

AND2x2_ASAP7_75t_L g373 ( 
.A(n_6),
.B(n_374),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_6),
.B(n_435),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g468 ( 
.A(n_6),
.B(n_444),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_SL g490 ( 
.A(n_6),
.B(n_491),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_SL g495 ( 
.A(n_6),
.B(n_496),
.Y(n_495)
);

AND2x2_ASAP7_75t_L g29 ( 
.A(n_7),
.B(n_30),
.Y(n_29)
);

AND2x2_ASAP7_75t_L g36 ( 
.A(n_7),
.B(n_37),
.Y(n_36)
);

AND2x2_ASAP7_75t_L g45 ( 
.A(n_7),
.B(n_46),
.Y(n_45)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_7),
.B(n_98),
.Y(n_97)
);

AND2x2_ASAP7_75t_L g133 ( 
.A(n_7),
.B(n_134),
.Y(n_133)
);

AND2x2_ASAP7_75t_L g135 ( 
.A(n_7),
.B(n_136),
.Y(n_135)
);

AND2x2_ASAP7_75t_L g139 ( 
.A(n_7),
.B(n_43),
.Y(n_139)
);

NAND2x1p5_ASAP7_75t_L g148 ( 
.A(n_7),
.B(n_149),
.Y(n_148)
);

BUFx5_ASAP7_75t_L g134 ( 
.A(n_8),
.Y(n_134)
);

BUFx5_ASAP7_75t_L g237 ( 
.A(n_8),
.Y(n_237)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_8),
.Y(n_285)
);

BUFx3_ASAP7_75t_L g322 ( 
.A(n_8),
.Y(n_322)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_9),
.Y(n_38)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_9),
.Y(n_91)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_9),
.Y(n_114)
);

BUFx3_ASAP7_75t_L g194 ( 
.A(n_9),
.Y(n_194)
);

INVx3_ASAP7_75t_L g292 ( 
.A(n_9),
.Y(n_292)
);

BUFx3_ASAP7_75t_L g372 ( 
.A(n_9),
.Y(n_372)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_10),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_11),
.B(n_56),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_11),
.B(n_75),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_11),
.B(n_86),
.Y(n_85)
);

AND2x2_ASAP7_75t_L g111 ( 
.A(n_11),
.B(n_112),
.Y(n_111)
);

NAND2x1_ASAP7_75t_SL g151 ( 
.A(n_11),
.B(n_152),
.Y(n_151)
);

AND2x2_ASAP7_75t_L g232 ( 
.A(n_11),
.B(n_233),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_11),
.B(n_30),
.Y(n_239)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_11),
.Y(n_319)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

AND2x2_ASAP7_75t_L g116 ( 
.A(n_12),
.B(n_88),
.Y(n_116)
);

AND2x2_ASAP7_75t_L g191 ( 
.A(n_12),
.B(n_192),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_12),
.B(n_257),
.Y(n_256)
);

AND2x2_ASAP7_75t_L g272 ( 
.A(n_12),
.B(n_273),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_12),
.B(n_283),
.Y(n_282)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_13),
.Y(n_35)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_13),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_13),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g278 ( 
.A(n_13),
.Y(n_278)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_14),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_14),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_15),
.B(n_43),
.Y(n_235)
);

AND2x2_ASAP7_75t_L g275 ( 
.A(n_15),
.B(n_276),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_15),
.B(n_327),
.Y(n_326)
);

AND2x2_ASAP7_75t_L g366 ( 
.A(n_15),
.B(n_367),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_15),
.B(n_443),
.Y(n_442)
);

AND2x2_ASAP7_75t_L g469 ( 
.A(n_15),
.B(n_119),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_L g477 ( 
.A(n_15),
.B(n_478),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_SL g500 ( 
.A(n_15),
.B(n_482),
.Y(n_500)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_16),
.Y(n_100)
);

BUFx12f_ASAP7_75t_L g186 ( 
.A(n_16),
.Y(n_186)
);

BUFx8_ASAP7_75t_L g43 ( 
.A(n_17),
.Y(n_43)
);

BUFx5_ASAP7_75t_L g63 ( 
.A(n_17),
.Y(n_63)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_17),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_160),
.Y(n_19)
);

NAND2xp33_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_159),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_140),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_23),
.B(n_140),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_80),
.C(n_105),
.Y(n_23)
);

XNOR2xp5_ASAP7_75t_L g167 ( 
.A(n_24),
.B(n_80),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g24 ( 
.A1(n_25),
.A2(n_26),
.B1(n_51),
.B2(n_52),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

XNOR2xp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_39),
.Y(n_26)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_27),
.B(n_39),
.C(n_51),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_31),
.C(n_36),
.Y(n_27)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_28),
.A2(n_29),
.B1(n_36),
.B2(n_49),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_28),
.A2(n_29),
.B1(n_96),
.B2(n_97),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g362 ( 
.A1(n_28),
.A2(n_29),
.B1(n_287),
.B2(n_363),
.Y(n_362)
);

INVx1_ASAP7_75t_SL g28 ( 
.A(n_29),
.Y(n_28)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_29),
.B(n_96),
.C(n_101),
.Y(n_95)
);

MAJx2_ASAP7_75t_L g286 ( 
.A(n_29),
.B(n_287),
.C(n_289),
.Y(n_286)
);

INVx2_ASAP7_75t_L g441 ( 
.A(n_30),
.Y(n_441)
);

INVx2_ASAP7_75t_SL g492 ( 
.A(n_30),
.Y(n_492)
);

XOR2xp5_ASAP7_75t_L g81 ( 
.A(n_31),
.B(n_82),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_32),
.B(n_33),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_32),
.B(n_41),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_32),
.B(n_102),
.Y(n_101)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_35),
.Y(n_196)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_35),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g44 ( 
.A1(n_36),
.A2(n_45),
.B1(n_49),
.B2(n_50),
.Y(n_44)
);

INVx1_ASAP7_75t_SL g49 ( 
.A(n_36),
.Y(n_49)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_36),
.B(n_118),
.C(n_262),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g311 ( 
.A1(n_36),
.A2(n_49),
.B1(n_117),
.B2(n_118),
.Y(n_311)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

XNOR2xp5_ASAP7_75t_L g39 ( 
.A(n_40),
.B(n_44),
.Y(n_39)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_40),
.Y(n_154)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_43),
.Y(n_181)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_45),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_45),
.A2(n_50),
.B1(n_147),
.B2(n_148),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_45),
.B(n_49),
.C(n_154),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_SL g249 ( 
.A1(n_45),
.A2(n_50),
.B1(n_219),
.B2(n_250),
.Y(n_249)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g438 ( 
.A(n_48),
.Y(n_438)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_50),
.B(n_123),
.C(n_219),
.Y(n_218)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

XNOR2xp5_ASAP7_75t_SL g52 ( 
.A(n_53),
.B(n_67),
.Y(n_52)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_53),
.B(n_68),
.C(n_74),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g53 ( 
.A(n_54),
.B(n_60),
.C(n_64),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_54),
.A2(n_55),
.B1(n_64),
.B2(n_127),
.Y(n_126)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

BUFx5_ASAP7_75t_L g254 ( 
.A(n_59),
.Y(n_254)
);

INVx2_ASAP7_75t_L g307 ( 
.A(n_59),
.Y(n_307)
);

BUFx6f_ASAP7_75t_L g317 ( 
.A(n_59),
.Y(n_317)
);

BUFx6f_ASAP7_75t_L g376 ( 
.A(n_59),
.Y(n_376)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_60),
.A2(n_125),
.B1(n_126),
.B2(n_128),
.Y(n_124)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_60),
.Y(n_128)
);

INVx1_ASAP7_75t_SL g61 ( 
.A(n_62),
.Y(n_61)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_62),
.Y(n_152)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_64),
.Y(n_127)
);

MAJx2_ASAP7_75t_L g190 ( 
.A(n_64),
.B(n_191),
.C(n_195),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_SL g217 ( 
.A(n_64),
.B(n_195),
.Y(n_217)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_66),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g369 ( 
.A(n_66),
.Y(n_369)
);

OAI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_68),
.A2(n_69),
.B1(n_73),
.B2(n_74),
.Y(n_67)
);

MAJx2_ASAP7_75t_L g189 ( 
.A(n_68),
.B(n_190),
.C(n_197),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_L g226 ( 
.A1(n_68),
.A2(n_69),
.B1(n_197),
.B2(n_227),
.Y(n_226)
);

INVx2_ASAP7_75t_SL g68 ( 
.A(n_69),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_69),
.B(n_130),
.C(n_138),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_69),
.B(n_139),
.Y(n_202)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_72),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g149 ( 
.A(n_72),
.Y(n_149)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

HB1xp67_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_81),
.B(n_83),
.C(n_95),
.Y(n_80)
);

XNOR2xp5_ASAP7_75t_L g171 ( 
.A(n_81),
.B(n_172),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_L g172 ( 
.A(n_83),
.B(n_95),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_84),
.B(n_89),
.C(n_92),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_84),
.A2(n_85),
.B1(n_89),
.B2(n_123),
.Y(n_122)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx5_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx5_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx1_ASAP7_75t_SL g123 ( 
.A(n_89),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_89),
.A2(n_123),
.B1(n_248),
.B2(n_249),
.Y(n_247)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

XNOR2xp5_ASAP7_75t_L g121 ( 
.A(n_92),
.B(n_122),
.Y(n_121)
);

XOR2xp5_ASAP7_75t_SL g145 ( 
.A(n_92),
.B(n_146),
.Y(n_145)
);

HB1xp67_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx6_ASAP7_75t_L g137 ( 
.A(n_94),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_96),
.A2(n_97),
.B1(n_132),
.B2(n_133),
.Y(n_177)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_97),
.B(n_132),
.C(n_135),
.Y(n_131)
);

AND2x2_ASAP7_75t_L g324 ( 
.A(n_97),
.B(n_236),
.Y(n_324)
);

XNOR2xp5_ASAP7_75t_L g418 ( 
.A(n_97),
.B(n_297),
.Y(n_418)
);

INVx5_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_100),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_SL g107 ( 
.A(n_101),
.B(n_108),
.Y(n_107)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx2_ASAP7_75t_SL g103 ( 
.A(n_104),
.Y(n_103)
);

XNOR2xp5_ASAP7_75t_L g166 ( 
.A(n_105),
.B(n_167),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_106),
.B(n_124),
.C(n_129),
.Y(n_105)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_106),
.B(n_170),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_107),
.B(n_109),
.C(n_121),
.Y(n_106)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_107),
.B(n_212),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g212 ( 
.A(n_109),
.B(n_121),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_110),
.B(n_115),
.C(n_117),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_110),
.A2(n_111),
.B1(n_115),
.B2(n_116),
.Y(n_188)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVx6_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

CKINVDCx16_ASAP7_75t_R g115 ( 
.A(n_116),
.Y(n_115)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

XNOR2xp5_ASAP7_75t_L g187 ( 
.A(n_118),
.B(n_188),
.Y(n_187)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

XNOR2xp5_ASAP7_75t_L g170 ( 
.A(n_124),
.B(n_129),
.Y(n_170)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

AO22x1_ASAP7_75t_SL g201 ( 
.A1(n_130),
.A2(n_131),
.B1(n_202),
.B2(n_203),
.Y(n_201)
);

INVx1_ASAP7_75t_SL g130 ( 
.A(n_131),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_132),
.B(n_179),
.C(n_182),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_132),
.A2(n_133),
.B1(n_182),
.B2(n_183),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g424 ( 
.A(n_132),
.B(n_425),
.Y(n_424)
);

INVx1_ASAP7_75t_SL g132 ( 
.A(n_133),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_L g454 ( 
.A(n_133),
.B(n_425),
.Y(n_454)
);

INVx3_ASAP7_75t_L g303 ( 
.A(n_134),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_135),
.B(n_177),
.Y(n_176)
);

INVx4_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

CKINVDCx14_ASAP7_75t_R g138 ( 
.A(n_139),
.Y(n_138)
);

XOR2xp5_ASAP7_75t_L g140 ( 
.A(n_141),
.B(n_142),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_143),
.A2(n_144),
.B1(n_157),
.B2(n_158),
.Y(n_142)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_143),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_144),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_SL g144 ( 
.A(n_145),
.B(n_150),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_147),
.B(n_230),
.C(n_238),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g347 ( 
.A1(n_147),
.A2(n_148),
.B1(n_238),
.B2(n_239),
.Y(n_347)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_151),
.A2(n_153),
.B1(n_155),
.B2(n_156),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_151),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_153),
.Y(n_156)
);

INVxp67_ASAP7_75t_SL g160 ( 
.A(n_161),
.Y(n_160)
);

AOI21xp5_ASAP7_75t_L g161 ( 
.A1(n_162),
.A2(n_240),
.B(n_512),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_164),
.B(n_204),
.Y(n_163)
);

INVxp67_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_L g512 ( 
.A1(n_165),
.A2(n_513),
.B(n_514),
.Y(n_512)
);

NOR2xp67_ASAP7_75t_SL g165 ( 
.A(n_166),
.B(n_168),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g514 ( 
.A(n_166),
.B(n_168),
.Y(n_514)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_171),
.C(n_173),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_L g206 ( 
.A(n_169),
.B(n_171),
.Y(n_206)
);

XOR2xp5_ASAP7_75t_L g205 ( 
.A(n_173),
.B(n_206),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_189),
.C(n_201),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_174),
.A2(n_175),
.B1(n_209),
.B2(n_210),
.Y(n_208)
);

INVx1_ASAP7_75t_SL g174 ( 
.A(n_175),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_176),
.B(n_178),
.C(n_187),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_L g392 ( 
.A(n_176),
.B(n_393),
.Y(n_392)
);

XNOR2xp5_ASAP7_75t_L g393 ( 
.A(n_178),
.B(n_187),
.Y(n_393)
);

XNOR2x1_ASAP7_75t_L g222 ( 
.A(n_179),
.B(n_223),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_SL g179 ( 
.A(n_180),
.B(n_181),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_180),
.B(n_314),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g370 ( 
.A(n_180),
.B(n_371),
.Y(n_370)
);

OAI22xp5_ASAP7_75t_SL g364 ( 
.A1(n_182),
.A2(n_183),
.B1(n_281),
.B2(n_282),
.Y(n_364)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_183),
.B(n_281),
.Y(n_280)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

INVx2_ASAP7_75t_SL g185 ( 
.A(n_186),
.Y(n_185)
);

INVx5_ASAP7_75t_L g274 ( 
.A(n_186),
.Y(n_274)
);

BUFx6f_ASAP7_75t_L g426 ( 
.A(n_186),
.Y(n_426)
);

INVx3_ASAP7_75t_L g452 ( 
.A(n_186),
.Y(n_452)
);

XNOR2xp5_ASAP7_75t_SL g209 ( 
.A(n_189),
.B(n_201),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_190),
.B(n_226),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_L g216 ( 
.A(n_191),
.B(n_217),
.Y(n_216)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_197),
.Y(n_227)
);

INVx8_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

INVx4_ASAP7_75t_L g263 ( 
.A(n_199),
.Y(n_263)
);

BUFx6f_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_202),
.Y(n_203)
);

OR2x6_ASAP7_75t_L g204 ( 
.A(n_205),
.B(n_207),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g513 ( 
.A(n_205),
.B(n_207),
.Y(n_513)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_211),
.C(n_213),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_L g401 ( 
.A(n_208),
.B(n_211),
.Y(n_401)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_209),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_L g400 ( 
.A(n_213),
.B(n_401),
.Y(n_400)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_214),
.B(n_224),
.C(n_228),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g389 ( 
.A1(n_214),
.A2(n_215),
.B1(n_390),
.B2(n_391),
.Y(n_389)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_216),
.B(n_218),
.C(n_221),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_L g338 ( 
.A(n_216),
.B(n_339),
.Y(n_338)
);

AOI22xp5_ASAP7_75t_SL g339 ( 
.A1(n_218),
.A2(n_221),
.B1(n_222),
.B2(n_340),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_218),
.Y(n_340)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_219),
.Y(n_250)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g390 ( 
.A1(n_224),
.A2(n_225),
.B1(n_228),
.B2(n_229),
.Y(n_390)
);

INVx1_ASAP7_75t_SL g224 ( 
.A(n_225),
.Y(n_224)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_SL g345 ( 
.A1(n_230),
.A2(n_231),
.B1(n_346),
.B2(n_347),
.Y(n_345)
);

INVx1_ASAP7_75t_SL g230 ( 
.A(n_231),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_232),
.B(n_235),
.C(n_236),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_232),
.A2(n_236),
.B1(n_296),
.B2(n_297),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_232),
.Y(n_296)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

INVx2_ASAP7_75t_L g499 ( 
.A(n_234),
.Y(n_499)
);

XNOR2xp5_ASAP7_75t_L g294 ( 
.A(n_235),
.B(n_295),
.Y(n_294)
);

INVx1_ASAP7_75t_SL g297 ( 
.A(n_236),
.Y(n_297)
);

INVx1_ASAP7_75t_SL g238 ( 
.A(n_239),
.Y(n_238)
);

NAND2x1_ASAP7_75t_L g240 ( 
.A(n_241),
.B(n_403),
.Y(n_240)
);

A2O1A1O1Ixp25_ASAP7_75t_L g241 ( 
.A1(n_242),
.A2(n_380),
.B(n_396),
.C(n_397),
.D(n_402),
.Y(n_241)
);

OAI21x1_ASAP7_75t_L g242 ( 
.A1(n_243),
.A2(n_352),
.B(n_379),
.Y(n_242)
);

NOR2x1_ASAP7_75t_L g404 ( 
.A(n_243),
.B(n_405),
.Y(n_404)
);

AND2x2_ASAP7_75t_L g243 ( 
.A(n_244),
.B(n_332),
.Y(n_243)
);

OR2x2_ASAP7_75t_L g379 ( 
.A(n_244),
.B(n_332),
.Y(n_379)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_245),
.B(n_293),
.C(n_309),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g377 ( 
.A(n_245),
.B(n_378),
.Y(n_377)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_246),
.B(n_264),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_247),
.B(n_251),
.Y(n_246)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_247),
.Y(n_334)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_251),
.Y(n_335)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_252),
.B(n_261),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_253),
.A2(n_255),
.B1(n_256),
.B2(n_260),
.Y(n_252)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_253),
.Y(n_260)
);

A2O1A1Ixp33_ASAP7_75t_L g348 ( 
.A1(n_253),
.A2(n_256),
.B(n_261),
.C(n_349),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_255),
.B(n_260),
.Y(n_349)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

INVx4_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

INVx8_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g310 ( 
.A(n_262),
.B(n_311),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_264),
.B(n_334),
.C(n_335),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_265),
.B(n_279),
.C(n_286),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_SL g357 ( 
.A(n_265),
.B(n_358),
.Y(n_357)
);

XNOR2xp5_ASAP7_75t_L g265 ( 
.A(n_266),
.B(n_271),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_266),
.B(n_272),
.C(n_275),
.Y(n_299)
);

HB1xp67_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

BUFx6f_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_272),
.B(n_275),
.Y(n_271)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

INVx3_ASAP7_75t_L g480 ( 
.A(n_274),
.Y(n_480)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

INVx3_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

INVx4_ASAP7_75t_L g331 ( 
.A(n_278),
.Y(n_331)
);

AOI22xp5_ASAP7_75t_L g358 ( 
.A1(n_279),
.A2(n_280),
.B1(n_286),
.B2(n_359),
.Y(n_358)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

BUFx3_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

INVx3_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

INVx2_ASAP7_75t_L g484 ( 
.A(n_285),
.Y(n_484)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_286),
.Y(n_359)
);

CKINVDCx14_ASAP7_75t_R g363 ( 
.A(n_287),
.Y(n_363)
);

XNOR2xp5_ASAP7_75t_L g361 ( 
.A(n_289),
.B(n_362),
.Y(n_361)
);

BUFx3_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

INVx2_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

BUFx3_ASAP7_75t_L g445 ( 
.A(n_292),
.Y(n_445)
);

XNOR2xp5_ASAP7_75t_L g378 ( 
.A(n_293),
.B(n_309),
.Y(n_378)
);

XNOR2xp5_ASAP7_75t_L g293 ( 
.A(n_294),
.B(n_298),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g343 ( 
.A(n_294),
.B(n_300),
.C(n_308),
.Y(n_343)
);

AOI22xp33_ASAP7_75t_SL g298 ( 
.A1(n_299),
.A2(n_300),
.B1(n_301),
.B2(n_308),
.Y(n_298)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_299),
.Y(n_308)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

AOI21xp5_ASAP7_75t_L g312 ( 
.A1(n_301),
.A2(n_313),
.B(n_318),
.Y(n_312)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_303),
.Y(n_302)
);

INVx3_ASAP7_75t_L g304 ( 
.A(n_305),
.Y(n_304)
);

BUFx6f_ASAP7_75t_L g305 ( 
.A(n_306),
.Y(n_305)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_306),
.Y(n_327)
);

BUFx6f_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_310),
.B(n_312),
.C(n_323),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_L g355 ( 
.A(n_310),
.B(n_312),
.Y(n_355)
);

INVx2_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

BUFx3_ASAP7_75t_L g315 ( 
.A(n_316),
.Y(n_315)
);

BUFx6f_ASAP7_75t_L g316 ( 
.A(n_317),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_319),
.B(n_320),
.Y(n_318)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_321),
.Y(n_320)
);

BUFx3_ASAP7_75t_L g321 ( 
.A(n_322),
.Y(n_321)
);

XNOR2xp5_ASAP7_75t_SL g354 ( 
.A(n_323),
.B(n_355),
.Y(n_354)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_324),
.B(n_325),
.C(n_328),
.Y(n_323)
);

XOR2xp5_ASAP7_75t_L g415 ( 
.A(n_324),
.B(n_416),
.Y(n_415)
);

AOI22xp5_ASAP7_75t_L g416 ( 
.A1(n_325),
.A2(n_326),
.B1(n_328),
.B2(n_329),
.Y(n_416)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_326),
.Y(n_325)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_329),
.Y(n_328)
);

INVx4_ASAP7_75t_L g330 ( 
.A(n_331),
.Y(n_330)
);

XNOR2xp5_ASAP7_75t_L g332 ( 
.A(n_333),
.B(n_336),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_L g381 ( 
.A(n_333),
.B(n_341),
.C(n_382),
.Y(n_381)
);

OAI22xp5_ASAP7_75t_SL g336 ( 
.A1(n_337),
.A2(n_338),
.B1(n_341),
.B2(n_342),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_338),
.Y(n_337)
);

HB1xp67_ASAP7_75t_L g382 ( 
.A(n_338),
.Y(n_382)
);

INVx1_ASAP7_75t_SL g341 ( 
.A(n_342),
.Y(n_341)
);

XNOR2xp5_ASAP7_75t_L g342 ( 
.A(n_343),
.B(n_344),
.Y(n_342)
);

INVxp67_ASAP7_75t_L g385 ( 
.A(n_343),
.Y(n_385)
);

AOI22xp5_ASAP7_75t_SL g344 ( 
.A1(n_345),
.A2(n_348),
.B1(n_350),
.B2(n_351),
.Y(n_344)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_345),
.Y(n_350)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_347),
.Y(n_346)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_348),
.Y(n_351)
);

HB1xp67_ASAP7_75t_L g386 ( 
.A(n_348),
.Y(n_386)
);

HB1xp67_ASAP7_75t_L g387 ( 
.A(n_350),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_353),
.B(n_377),
.Y(n_352)
);

NOR2xp33_ASAP7_75t_L g405 ( 
.A(n_353),
.B(n_377),
.Y(n_405)
);

MAJIxp5_ASAP7_75t_L g353 ( 
.A(n_354),
.B(n_356),
.C(n_360),
.Y(n_353)
);

XOR2xp5_ASAP7_75t_L g408 ( 
.A(n_354),
.B(n_409),
.Y(n_408)
);

AOI22xp5_ASAP7_75t_L g409 ( 
.A1(n_356),
.A2(n_357),
.B1(n_360),
.B2(n_410),
.Y(n_409)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_357),
.Y(n_356)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_360),
.Y(n_410)
);

MAJIxp5_ASAP7_75t_L g360 ( 
.A(n_361),
.B(n_364),
.C(n_365),
.Y(n_360)
);

XNOR2xp5_ASAP7_75t_L g413 ( 
.A(n_361),
.B(n_414),
.Y(n_413)
);

XNOR2xp5_ASAP7_75t_L g414 ( 
.A(n_364),
.B(n_365),
.Y(n_414)
);

MAJx2_ASAP7_75t_L g365 ( 
.A(n_366),
.B(n_370),
.C(n_373),
.Y(n_365)
);

XNOR2xp5_ASAP7_75t_L g459 ( 
.A(n_366),
.B(n_373),
.Y(n_459)
);

INVx3_ASAP7_75t_L g367 ( 
.A(n_368),
.Y(n_367)
);

INVx2_ASAP7_75t_L g368 ( 
.A(n_369),
.Y(n_368)
);

XNOR2xp5_ASAP7_75t_L g458 ( 
.A(n_370),
.B(n_459),
.Y(n_458)
);

INVx5_ASAP7_75t_L g371 ( 
.A(n_372),
.Y(n_371)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_375),
.Y(n_374)
);

INVx2_ASAP7_75t_L g375 ( 
.A(n_376),
.Y(n_375)
);

NAND4xp25_ASAP7_75t_SL g403 ( 
.A(n_380),
.B(n_397),
.C(n_404),
.D(n_406),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_381),
.B(n_383),
.Y(n_380)
);

NOR2xp33_ASAP7_75t_L g396 ( 
.A(n_381),
.B(n_383),
.Y(n_396)
);

XNOR2xp5_ASAP7_75t_L g383 ( 
.A(n_384),
.B(n_388),
.Y(n_383)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_384),
.Y(n_399)
);

MAJIxp5_ASAP7_75t_L g384 ( 
.A(n_385),
.B(n_386),
.C(n_387),
.Y(n_384)
);

AOI22xp5_ASAP7_75t_SL g388 ( 
.A1(n_389),
.A2(n_392),
.B1(n_394),
.B2(n_395),
.Y(n_388)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_389),
.Y(n_394)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_390),
.Y(n_391)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_392),
.Y(n_395)
);

MAJIxp5_ASAP7_75t_L g398 ( 
.A(n_392),
.B(n_394),
.C(n_399),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_398),
.B(n_400),
.Y(n_397)
);

NOR2xp33_ASAP7_75t_L g402 ( 
.A(n_398),
.B(n_400),
.Y(n_402)
);

OAI21x1_ASAP7_75t_SL g406 ( 
.A1(n_407),
.A2(n_427),
.B(n_511),
.Y(n_406)
);

NOR2xp67_ASAP7_75t_SL g407 ( 
.A(n_408),
.B(n_411),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_SL g511 ( 
.A(n_408),
.B(n_411),
.Y(n_511)
);

MAJIxp5_ASAP7_75t_L g411 ( 
.A(n_412),
.B(n_415),
.C(n_417),
.Y(n_411)
);

AOI22xp5_ASAP7_75t_SL g507 ( 
.A1(n_412),
.A2(n_413),
.B1(n_508),
.B2(n_509),
.Y(n_507)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_413),
.Y(n_412)
);

XNOR2xp5_ASAP7_75t_SL g509 ( 
.A(n_415),
.B(n_417),
.Y(n_509)
);

MAJIxp5_ASAP7_75t_L g417 ( 
.A(n_418),
.B(n_419),
.C(n_424),
.Y(n_417)
);

AOI22xp5_ASAP7_75t_L g461 ( 
.A1(n_418),
.A2(n_419),
.B1(n_420),
.B2(n_462),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_418),
.Y(n_462)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_420),
.Y(n_419)
);

INVx4_ASAP7_75t_L g421 ( 
.A(n_422),
.Y(n_421)
);

INVx6_ASAP7_75t_L g422 ( 
.A(n_423),
.Y(n_422)
);

XNOR2xp5_ASAP7_75t_SL g460 ( 
.A(n_424),
.B(n_461),
.Y(n_460)
);

AOI21x1_ASAP7_75t_SL g427 ( 
.A1(n_428),
.A2(n_505),
.B(n_510),
.Y(n_427)
);

OAI21xp5_ASAP7_75t_L g428 ( 
.A1(n_429),
.A2(n_463),
.B(n_504),
.Y(n_428)
);

NOR2xp33_ASAP7_75t_L g429 ( 
.A(n_430),
.B(n_455),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_SL g504 ( 
.A(n_430),
.B(n_455),
.Y(n_504)
);

MAJIxp5_ASAP7_75t_L g430 ( 
.A(n_431),
.B(n_446),
.C(n_453),
.Y(n_430)
);

AOI22xp33_ASAP7_75t_SL g470 ( 
.A1(n_431),
.A2(n_432),
.B1(n_471),
.B2(n_473),
.Y(n_470)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_432),
.Y(n_431)
);

XOR2xp5_ASAP7_75t_L g432 ( 
.A(n_433),
.B(n_442),
.Y(n_432)
);

XNOR2xp5_ASAP7_75t_L g433 ( 
.A(n_434),
.B(n_439),
.Y(n_433)
);

MAJIxp5_ASAP7_75t_L g457 ( 
.A(n_434),
.B(n_439),
.C(n_442),
.Y(n_457)
);

INVx2_ASAP7_75t_L g435 ( 
.A(n_436),
.Y(n_435)
);

INVx2_ASAP7_75t_L g436 ( 
.A(n_437),
.Y(n_436)
);

INVx2_ASAP7_75t_L g437 ( 
.A(n_438),
.Y(n_437)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_441),
.Y(n_440)
);

BUFx3_ASAP7_75t_L g443 ( 
.A(n_444),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_445),
.Y(n_444)
);

AOI22xp5_ASAP7_75t_L g471 ( 
.A1(n_446),
.A2(n_453),
.B1(n_454),
.B2(n_472),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_446),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_L g446 ( 
.A(n_447),
.B(n_449),
.Y(n_446)
);

OAI22xp5_ASAP7_75t_SL g466 ( 
.A1(n_447),
.A2(n_448),
.B1(n_449),
.B2(n_450),
.Y(n_466)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_448),
.Y(n_447)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_450),
.Y(n_449)
);

INVx4_ASAP7_75t_L g451 ( 
.A(n_452),
.Y(n_451)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_454),
.Y(n_453)
);

XNOR2xp5_ASAP7_75t_L g455 ( 
.A(n_456),
.B(n_460),
.Y(n_455)
);

XNOR2xp5_ASAP7_75t_L g456 ( 
.A(n_457),
.B(n_458),
.Y(n_456)
);

MAJIxp5_ASAP7_75t_L g506 ( 
.A(n_457),
.B(n_458),
.C(n_460),
.Y(n_506)
);

AOI21xp5_ASAP7_75t_L g463 ( 
.A1(n_464),
.A2(n_474),
.B(n_503),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_L g464 ( 
.A(n_465),
.B(n_470),
.Y(n_464)
);

NOR2xp33_ASAP7_75t_SL g503 ( 
.A(n_465),
.B(n_470),
.Y(n_503)
);

MAJIxp5_ASAP7_75t_L g465 ( 
.A(n_466),
.B(n_467),
.C(n_469),
.Y(n_465)
);

XOR2xp5_ASAP7_75t_L g485 ( 
.A(n_466),
.B(n_486),
.Y(n_485)
);

OAI22xp5_ASAP7_75t_SL g486 ( 
.A1(n_467),
.A2(n_468),
.B1(n_469),
.B2(n_487),
.Y(n_486)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_468),
.Y(n_467)
);

CKINVDCx16_ASAP7_75t_R g487 ( 
.A(n_469),
.Y(n_487)
);

INVxp67_ASAP7_75t_SL g473 ( 
.A(n_471),
.Y(n_473)
);

OAI21xp5_ASAP7_75t_SL g474 ( 
.A1(n_475),
.A2(n_488),
.B(n_502),
.Y(n_474)
);

NOR2xp33_ASAP7_75t_L g475 ( 
.A(n_476),
.B(n_485),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_SL g502 ( 
.A(n_476),
.B(n_485),
.Y(n_502)
);

NOR2xp33_ASAP7_75t_L g476 ( 
.A(n_477),
.B(n_481),
.Y(n_476)
);

XNOR2xp5_ASAP7_75t_L g493 ( 
.A(n_477),
.B(n_481),
.Y(n_493)
);

INVx2_ASAP7_75t_L g478 ( 
.A(n_479),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_480),
.Y(n_479)
);

INVx2_ASAP7_75t_L g482 ( 
.A(n_483),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_484),
.Y(n_483)
);

AOI21xp5_ASAP7_75t_L g488 ( 
.A1(n_489),
.A2(n_494),
.B(n_501),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_L g489 ( 
.A(n_490),
.B(n_493),
.Y(n_489)
);

NOR2xp33_ASAP7_75t_SL g501 ( 
.A(n_490),
.B(n_493),
.Y(n_501)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_492),
.Y(n_491)
);

NOR2xp33_ASAP7_75t_L g494 ( 
.A(n_495),
.B(n_500),
.Y(n_494)
);

INVx2_ASAP7_75t_L g496 ( 
.A(n_497),
.Y(n_496)
);

BUFx2_ASAP7_75t_L g497 ( 
.A(n_498),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_499),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_L g505 ( 
.A(n_506),
.B(n_507),
.Y(n_505)
);

NOR2xp33_ASAP7_75t_SL g510 ( 
.A(n_506),
.B(n_507),
.Y(n_510)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_509),
.Y(n_508)
);


endmodule