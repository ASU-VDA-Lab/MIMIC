module fake_jpeg_11286_n_115 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_115);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_115;

wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_93;
wire n_91;
wire n_101;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_100;
wire n_82;
wire n_96;

INVx3_ASAP7_75t_L g34 ( 
.A(n_7),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_5),
.B(n_21),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_31),
.Y(n_36)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_4),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_24),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_15),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_33),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_20),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_2),
.Y(n_42)
);

BUFx5_ASAP7_75t_L g43 ( 
.A(n_6),
.Y(n_43)
);

BUFx16f_ASAP7_75t_L g44 ( 
.A(n_23),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_16),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_5),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_9),
.B(n_4),
.Y(n_47)
);

BUFx16f_ASAP7_75t_L g48 ( 
.A(n_46),
.Y(n_48)
);

INVx5_ASAP7_75t_SL g70 ( 
.A(n_48),
.Y(n_70)
);

BUFx10_ASAP7_75t_L g49 ( 
.A(n_44),
.Y(n_49)
);

CKINVDCx16_ASAP7_75t_R g58 ( 
.A(n_49),
.Y(n_58)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_44),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_50),
.B(n_51),
.Y(n_59)
);

INVx11_ASAP7_75t_L g51 ( 
.A(n_44),
.Y(n_51)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_34),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_52),
.B(n_53),
.Y(n_69)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_43),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_35),
.B(n_0),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_54),
.B(n_34),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_35),
.B(n_0),
.Y(n_55)
);

AND2x2_ASAP7_75t_L g62 ( 
.A(n_55),
.B(n_37),
.Y(n_62)
);

BUFx12f_ASAP7_75t_L g56 ( 
.A(n_43),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_56),
.B(n_57),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_SL g57 ( 
.A(n_47),
.B(n_42),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_61),
.B(n_64),
.Y(n_74)
);

AND2x2_ASAP7_75t_L g79 ( 
.A(n_62),
.B(n_1),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_48),
.B(n_39),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_SL g80 ( 
.A(n_63),
.B(n_66),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_50),
.B(n_36),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_49),
.B(n_38),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_65),
.B(n_67),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_48),
.B(n_41),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_49),
.B(n_40),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_51),
.B(n_45),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_68),
.B(n_22),
.Y(n_85)
);

AOI21xp5_ASAP7_75t_L g71 ( 
.A1(n_69),
.A2(n_37),
.B(n_56),
.Y(n_71)
);

OAI21xp5_ASAP7_75t_SL g98 ( 
.A1(n_71),
.A2(n_12),
.B(n_13),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_69),
.A2(n_46),
.B1(n_53),
.B2(n_56),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_72),
.A2(n_78),
.B1(n_82),
.B2(n_76),
.Y(n_96)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_59),
.Y(n_73)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_73),
.Y(n_95)
);

CKINVDCx16_ASAP7_75t_R g75 ( 
.A(n_70),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_75),
.B(n_79),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_59),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_77),
.B(n_85),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_58),
.A2(n_46),
.B1(n_2),
.B2(n_3),
.Y(n_78)
);

INVx5_ASAP7_75t_L g81 ( 
.A(n_60),
.Y(n_81)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_81),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_61),
.A2(n_1),
.B1(n_3),
.B2(n_6),
.Y(n_82)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_64),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_83),
.B(n_84),
.Y(n_87)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_64),
.Y(n_84)
);

XNOR2xp5_ASAP7_75t_SL g86 ( 
.A(n_61),
.B(n_25),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_86),
.B(n_17),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_SL g88 ( 
.A(n_79),
.B(n_7),
.C(n_8),
.Y(n_88)
);

AOI21xp5_ASAP7_75t_L g105 ( 
.A1(n_88),
.A2(n_90),
.B(n_97),
.Y(n_105)
);

INVxp33_ASAP7_75t_SL g90 ( 
.A(n_72),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_74),
.B(n_8),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_92),
.B(n_93),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_81),
.B(n_9),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_96),
.B(n_99),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_SL g97 ( 
.A(n_80),
.B(n_10),
.C(n_11),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_L g102 ( 
.A1(n_98),
.A2(n_100),
.B(n_82),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_86),
.B(n_14),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_87),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_101),
.B(n_102),
.C(n_91),
.Y(n_109)
);

O2A1O1Ixp33_ASAP7_75t_L g106 ( 
.A1(n_90),
.A2(n_78),
.B(n_19),
.C(n_26),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_106),
.A2(n_89),
.B1(n_94),
.B2(n_98),
.Y(n_108)
);

XOR2xp5_ASAP7_75t_L g107 ( 
.A(n_104),
.B(n_95),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_107),
.A2(n_108),
.B1(n_109),
.B2(n_89),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_110),
.A2(n_107),
.B1(n_105),
.B2(n_103),
.Y(n_111)
);

AOI21xp5_ASAP7_75t_L g112 ( 
.A1(n_111),
.A2(n_18),
.B(n_27),
.Y(n_112)
);

AOI21xp5_ASAP7_75t_L g113 ( 
.A1(n_112),
.A2(n_28),
.B(n_29),
.Y(n_113)
);

XOR2xp5_ASAP7_75t_L g114 ( 
.A(n_113),
.B(n_30),
.Y(n_114)
);

XOR2xp5_ASAP7_75t_L g115 ( 
.A(n_114),
.B(n_32),
.Y(n_115)
);


endmodule