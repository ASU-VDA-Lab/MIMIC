module real_jpeg_33869_n_8 (n_5, n_4, n_0, n_1, n_2, n_6, n_7, n_3, n_8);

input n_5;
input n_4;
input n_0;
input n_1;
input n_2;
input n_6;
input n_7;
input n_3;

output n_8;

wire n_17;
wire n_43;
wire n_54;
wire n_37;
wire n_21;
wire n_33;
wire n_35;
wire n_38;
wire n_50;
wire n_29;
wire n_55;
wire n_49;
wire n_52;
wire n_31;
wire n_9;
wire n_10;
wire n_12;
wire n_24;
wire n_34;
wire n_28;
wire n_44;
wire n_46;
wire n_23;
wire n_11;
wire n_14;
wire n_51;
wire n_47;
wire n_45;
wire n_25;
wire n_42;
wire n_22;
wire n_18;
wire n_53;
wire n_39;
wire n_40;
wire n_36;
wire n_41;
wire n_27;
wire n_32;
wire n_20;
wire n_48;
wire n_19;
wire n_26;
wire n_30;
wire n_16;
wire n_15;
wire n_13;

AND2x2_ASAP7_75t_L g21 ( 
.A(n_0),
.B(n_1),
.Y(n_21)
);

CKINVDCx11_ASAP7_75t_R g36 ( 
.A(n_0),
.Y(n_36)
);

AND2x2_ASAP7_75t_L g40 ( 
.A(n_0),
.B(n_41),
.Y(n_40)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_1),
.Y(n_41)
);

BUFx2_ASAP7_75t_R g19 ( 
.A(n_2),
.Y(n_19)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

NAND2x1p5_ASAP7_75t_L g29 ( 
.A(n_2),
.B(n_17),
.Y(n_29)
);

AND2x4_ASAP7_75t_SL g11 ( 
.A(n_3),
.B(n_12),
.Y(n_11)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_3),
.B(n_23),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_3),
.B(n_52),
.Y(n_54)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

OA22x2_ASAP7_75t_L g15 ( 
.A1(n_5),
.A2(n_6),
.B1(n_16),
.B2(n_17),
.Y(n_15)
);

INVx2_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

AO21x1_ASAP7_75t_L g52 ( 
.A1(n_5),
.A2(n_27),
.B(n_29),
.Y(n_52)
);

INVx3_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

AND2x2_ASAP7_75t_L g27 ( 
.A(n_6),
.B(n_28),
.Y(n_27)
);

AOI221xp5_ASAP7_75t_L g31 ( 
.A1(n_7),
.A2(n_32),
.B1(n_33),
.B2(n_34),
.C(n_37),
.Y(n_31)
);

OAI211xp5_ASAP7_75t_L g8 ( 
.A1(n_9),
.A2(n_24),
.B(n_31),
.C(n_55),
.Y(n_8)
);

NAND2xp5_ASAP7_75t_SL g9 ( 
.A(n_10),
.B(n_20),
.Y(n_9)
);

INVx2_ASAP7_75t_SL g10 ( 
.A(n_11),
.Y(n_10)
);

NAND2xp5_ASAP7_75t_SL g55 ( 
.A(n_11),
.B(n_48),
.Y(n_55)
);

AOI21xp5_ASAP7_75t_L g38 ( 
.A1(n_12),
.A2(n_39),
.B(n_42),
.Y(n_38)
);

INVx2_ASAP7_75t_L g12 ( 
.A(n_13),
.Y(n_12)
);

AND2x2_ASAP7_75t_L g32 ( 
.A(n_13),
.B(n_30),
.Y(n_32)
);

OA22x2_ASAP7_75t_L g13 ( 
.A1(n_14),
.A2(n_15),
.B1(n_18),
.B2(n_19),
.Y(n_13)
);

INVx2_ASAP7_75t_L g14 ( 
.A(n_15),
.Y(n_14)
);

OA21x2_ASAP7_75t_L g26 ( 
.A1(n_16),
.A2(n_27),
.B(n_29),
.Y(n_26)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

AND2x4_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_22),
.Y(n_20)
);

AND2x2_ASAP7_75t_L g33 ( 
.A(n_21),
.B(n_23),
.Y(n_33)
);

AND2x4_ASAP7_75t_L g48 ( 
.A(n_22),
.B(n_40),
.Y(n_48)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

AND2x2_ASAP7_75t_SL g39 ( 
.A(n_23),
.B(n_40),
.Y(n_39)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_SL g25 ( 
.A(n_26),
.B(n_30),
.Y(n_25)
);

OR2x2_ASAP7_75t_L g46 ( 
.A(n_26),
.B(n_30),
.Y(n_46)
);

NAND2xp67_ASAP7_75t_SL g50 ( 
.A(n_30),
.B(n_51),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g47 ( 
.A1(n_33),
.A2(n_48),
.B1(n_49),
.B2(n_53),
.Y(n_47)
);

BUFx12f_ASAP7_75t_SL g34 ( 
.A(n_35),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

OAI21xp33_ASAP7_75t_L g37 ( 
.A1(n_38),
.A2(n_45),
.B(n_47),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_40),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_43),
.B(n_44),
.Y(n_42)
);

CKINVDCx16_ASAP7_75t_R g45 ( 
.A(n_46),
.Y(n_45)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);


endmodule