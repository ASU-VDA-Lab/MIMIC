module real_aes_2574_n_104 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_822, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_103, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_104);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_822;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_103;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_104;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_571;
wire n_376;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_537;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_578;
wire n_528;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_559;
wire n_466;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_535;
wire n_732;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_755;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_746;
wire n_178;
wire n_409;
wire n_748;
wire n_781;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_504;
wire n_310;
wire n_455;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_812;
wire n_817;
wire n_443;
wire n_565;
wire n_782;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_808;
wire n_770;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_502;
wire n_505;
wire n_434;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_552;
wire n_402;
wire n_617;
wire n_733;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_807;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_790;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_288;
wire n_147;
wire n_150;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_810;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_749;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_765;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_809;
wire n_482;
wire n_520;
wire n_679;
wire n_633;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_623;
wire n_249;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_771;
wire n_524;
wire n_219;
wire n_705;
wire n_180;
wire n_212;
wire n_575;
wire n_210;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_393;
wire n_294;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_804;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_802;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_554;
wire n_475;
wire n_264;
wire n_798;
wire n_237;
wire n_668;
wire n_797;
NAND2xp5_ASAP7_75t_L g574 ( .A(n_0), .B(n_268), .Y(n_574) );
NAND2xp5_ASAP7_75t_L g817 ( .A(n_1), .B(n_818), .Y(n_817) );
INVx1_ASAP7_75t_L g157 ( .A(n_2), .Y(n_157) );
NAND2xp5_ASAP7_75t_L g531 ( .A(n_3), .B(n_524), .Y(n_531) );
NAND2xp33_ASAP7_75t_SL g567 ( .A(n_4), .B(n_169), .Y(n_567) );
NAND2xp5_ASAP7_75t_SL g260 ( .A(n_5), .B(n_176), .Y(n_260) );
INVx1_ASAP7_75t_L g560 ( .A(n_6), .Y(n_560) );
INVx1_ASAP7_75t_L g240 ( .A(n_7), .Y(n_240) );
OAI22xp5_ASAP7_75t_SL g501 ( .A1(n_8), .A2(n_502), .B1(n_503), .B2(n_505), .Y(n_501) );
CKINVDCx20_ASAP7_75t_R g502 ( .A(n_8), .Y(n_502) );
CKINVDCx16_ASAP7_75t_R g818 ( .A(n_9), .Y(n_818) );
NAND2xp5_ASAP7_75t_L g489 ( .A(n_10), .B(n_490), .Y(n_489) );
CKINVDCx5p33_ASAP7_75t_R g205 ( .A(n_11), .Y(n_205) );
AND2x2_ASAP7_75t_L g529 ( .A(n_12), .B(n_181), .Y(n_529) );
INVx2_ASAP7_75t_L g146 ( .A(n_13), .Y(n_146) );
CKINVDCx20_ASAP7_75t_R g504 ( .A(n_14), .Y(n_504) );
CKINVDCx16_ASAP7_75t_R g117 ( .A(n_15), .Y(n_117) );
NOR2xp33_ASAP7_75t_L g801 ( .A(n_15), .B(n_25), .Y(n_801) );
NOR3xp33_ASAP7_75t_L g816 ( .A(n_15), .B(n_817), .C(n_819), .Y(n_816) );
OAI22xp5_ASAP7_75t_SL g127 ( .A1(n_16), .A2(n_25), .B1(n_128), .B2(n_129), .Y(n_127) );
CKINVDCx20_ASAP7_75t_R g128 ( .A(n_16), .Y(n_128) );
INVx1_ASAP7_75t_L g269 ( .A(n_17), .Y(n_269) );
AOI221x1_ASAP7_75t_L g563 ( .A1(n_18), .A2(n_143), .B1(n_519), .B2(n_564), .C(n_566), .Y(n_563) );
NAND2xp5_ASAP7_75t_SL g550 ( .A(n_19), .B(n_524), .Y(n_550) );
INVx1_ASAP7_75t_L g121 ( .A(n_20), .Y(n_121) );
INVx1_ASAP7_75t_L g266 ( .A(n_21), .Y(n_266) );
INVx1_ASAP7_75t_SL g186 ( .A(n_22), .Y(n_186) );
NAND2xp5_ASAP7_75t_SL g256 ( .A(n_23), .B(n_163), .Y(n_256) );
AOI33xp33_ASAP7_75t_L g226 ( .A1(n_24), .A2(n_55), .A3(n_152), .B1(n_161), .B2(n_227), .B3(n_228), .Y(n_226) );
INVx1_ASAP7_75t_L g129 ( .A(n_25), .Y(n_129) );
AOI21xp5_ASAP7_75t_L g532 ( .A1(n_26), .A2(n_519), .B(n_533), .Y(n_532) );
NAND2xp5_ASAP7_75t_L g534 ( .A(n_27), .B(n_268), .Y(n_534) );
AOI221xp5_ASAP7_75t_SL g542 ( .A1(n_28), .A2(n_44), .B1(n_519), .B2(n_524), .C(n_543), .Y(n_542) );
INVx1_ASAP7_75t_L g197 ( .A(n_29), .Y(n_197) );
OA21x2_ASAP7_75t_L g145 ( .A1(n_30), .A2(n_93), .B(n_146), .Y(n_145) );
OR2x2_ASAP7_75t_L g177 ( .A(n_30), .B(n_93), .Y(n_177) );
NAND2xp5_ASAP7_75t_L g554 ( .A(n_31), .B(n_271), .Y(n_554) );
INVxp67_ASAP7_75t_L g562 ( .A(n_32), .Y(n_562) );
AND2x2_ASAP7_75t_L g590 ( .A(n_33), .B(n_180), .Y(n_590) );
NAND2xp5_ASAP7_75t_L g183 ( .A(n_34), .B(n_171), .Y(n_183) );
AOI21xp5_ASAP7_75t_L g572 ( .A1(n_35), .A2(n_519), .B(n_573), .Y(n_572) );
AOI22xp5_ASAP7_75t_L g104 ( .A1(n_36), .A2(n_105), .B1(n_812), .B2(n_813), .Y(n_104) );
NAND2xp5_ASAP7_75t_L g544 ( .A(n_37), .B(n_271), .Y(n_544) );
INVx1_ASAP7_75t_L g151 ( .A(n_38), .Y(n_151) );
AND2x2_ASAP7_75t_L g169 ( .A(n_38), .B(n_157), .Y(n_169) );
AND2x2_ASAP7_75t_L g175 ( .A(n_38), .B(n_154), .Y(n_175) );
OR2x6_ASAP7_75t_L g119 ( .A(n_39), .B(n_120), .Y(n_119) );
INVxp67_ASAP7_75t_L g819 ( .A(n_39), .Y(n_819) );
CKINVDCx20_ASAP7_75t_R g200 ( .A(n_40), .Y(n_200) );
NAND2xp5_ASAP7_75t_L g212 ( .A(n_41), .B(n_171), .Y(n_212) );
AOI22xp5_ASAP7_75t_L g249 ( .A1(n_42), .A2(n_144), .B1(n_176), .B2(n_250), .Y(n_249) );
NAND2xp5_ASAP7_75t_L g257 ( .A(n_43), .B(n_258), .Y(n_257) );
AOI22xp5_ASAP7_75t_L g625 ( .A1(n_45), .A2(n_84), .B1(n_149), .B2(n_519), .Y(n_625) );
NAND2xp5_ASAP7_75t_L g187 ( .A(n_46), .B(n_163), .Y(n_187) );
NAND2xp5_ASAP7_75t_L g588 ( .A(n_47), .B(n_268), .Y(n_588) );
XNOR2xp5_ASAP7_75t_L g131 ( .A(n_48), .B(n_88), .Y(n_131) );
NAND2xp5_ASAP7_75t_SL g242 ( .A(n_49), .B(n_221), .Y(n_242) );
NAND2xp5_ASAP7_75t_L g241 ( .A(n_50), .B(n_163), .Y(n_241) );
CKINVDCx5p33_ASAP7_75t_R g253 ( .A(n_51), .Y(n_253) );
AND2x2_ASAP7_75t_L g577 ( .A(n_52), .B(n_180), .Y(n_577) );
CKINVDCx20_ASAP7_75t_R g809 ( .A(n_53), .Y(n_809) );
NAND2xp5_ASAP7_75t_L g546 ( .A(n_54), .B(n_180), .Y(n_546) );
NAND2xp5_ASAP7_75t_L g216 ( .A(n_56), .B(n_163), .Y(n_216) );
INVx1_ASAP7_75t_L g156 ( .A(n_57), .Y(n_156) );
INVx1_ASAP7_75t_L g165 ( .A(n_57), .Y(n_165) );
AND2x2_ASAP7_75t_L g217 ( .A(n_58), .B(n_180), .Y(n_217) );
AOI221xp5_ASAP7_75t_L g238 ( .A1(n_59), .A2(n_77), .B1(n_149), .B2(n_171), .C(n_239), .Y(n_238) );
NAND2xp5_ASAP7_75t_L g170 ( .A(n_60), .B(n_171), .Y(n_170) );
NAND2xp5_ASAP7_75t_SL g589 ( .A(n_61), .B(n_524), .Y(n_589) );
NAND2xp5_ASAP7_75t_L g207 ( .A(n_62), .B(n_144), .Y(n_207) );
AOI21xp5_ASAP7_75t_SL g148 ( .A1(n_63), .A2(n_149), .B(n_158), .Y(n_148) );
AND2x2_ASAP7_75t_L g525 ( .A(n_64), .B(n_180), .Y(n_525) );
NAND2xp5_ASAP7_75t_L g575 ( .A(n_65), .B(n_271), .Y(n_575) );
INVx1_ASAP7_75t_L g263 ( .A(n_66), .Y(n_263) );
NAND2xp5_ASAP7_75t_L g522 ( .A(n_67), .B(n_268), .Y(n_522) );
AND2x2_ASAP7_75t_SL g555 ( .A(n_68), .B(n_181), .Y(n_555) );
XNOR2xp5_ASAP7_75t_L g503 ( .A(n_69), .B(n_504), .Y(n_503) );
AOI21xp5_ASAP7_75t_L g585 ( .A1(n_70), .A2(n_519), .B(n_586), .Y(n_585) );
INVx1_ASAP7_75t_L g215 ( .A(n_71), .Y(n_215) );
NAND2xp5_ASAP7_75t_L g535 ( .A(n_72), .B(n_271), .Y(n_535) );
AND2x2_ASAP7_75t_SL g626 ( .A(n_73), .B(n_221), .Y(n_626) );
AOI21xp5_ASAP7_75t_L g213 ( .A1(n_74), .A2(n_149), .B(n_214), .Y(n_213) );
INVx1_ASAP7_75t_L g154 ( .A(n_75), .Y(n_154) );
INVx1_ASAP7_75t_L g167 ( .A(n_75), .Y(n_167) );
NAND2xp5_ASAP7_75t_L g229 ( .A(n_76), .B(n_171), .Y(n_229) );
AND2x2_ASAP7_75t_L g188 ( .A(n_78), .B(n_143), .Y(n_188) );
INVx1_ASAP7_75t_L g264 ( .A(n_79), .Y(n_264) );
AOI21xp5_ASAP7_75t_L g184 ( .A1(n_80), .A2(n_149), .B(n_185), .Y(n_184) );
A2O1A1Ixp33_ASAP7_75t_L g254 ( .A1(n_81), .A2(n_149), .B(n_220), .C(n_255), .Y(n_254) );
NAND2xp5_ASAP7_75t_SL g523 ( .A(n_82), .B(n_524), .Y(n_523) );
AOI22xp5_ASAP7_75t_L g624 ( .A1(n_83), .A2(n_87), .B1(n_171), .B2(n_524), .Y(n_624) );
INVx1_ASAP7_75t_L g122 ( .A(n_85), .Y(n_122) );
AND2x2_ASAP7_75t_SL g142 ( .A(n_86), .B(n_143), .Y(n_142) );
AOI22xp5_ASAP7_75t_L g223 ( .A1(n_89), .A2(n_149), .B1(n_224), .B2(n_225), .Y(n_223) );
NAND2xp5_ASAP7_75t_L g553 ( .A(n_90), .B(n_268), .Y(n_553) );
NAND2xp5_ASAP7_75t_L g545 ( .A(n_91), .B(n_268), .Y(n_545) );
AOI21xp5_ASAP7_75t_L g518 ( .A1(n_92), .A2(n_519), .B(n_520), .Y(n_518) );
INVx1_ASAP7_75t_L g159 ( .A(n_94), .Y(n_159) );
NAND2xp5_ASAP7_75t_L g521 ( .A(n_95), .B(n_271), .Y(n_521) );
AND2x2_ASAP7_75t_L g230 ( .A(n_96), .B(n_143), .Y(n_230) );
A2O1A1Ixp33_ASAP7_75t_L g194 ( .A1(n_97), .A2(n_195), .B(n_196), .C(n_199), .Y(n_194) );
INVxp67_ASAP7_75t_L g565 ( .A(n_98), .Y(n_565) );
NAND2xp5_ASAP7_75t_L g576 ( .A(n_99), .B(n_524), .Y(n_576) );
NAND2xp5_ASAP7_75t_L g587 ( .A(n_100), .B(n_271), .Y(n_587) );
AOI21xp5_ASAP7_75t_L g551 ( .A1(n_101), .A2(n_519), .B(n_552), .Y(n_551) );
BUFx2_ASAP7_75t_SL g110 ( .A(n_102), .Y(n_110) );
BUFx2_ASAP7_75t_L g497 ( .A(n_102), .Y(n_497) );
NAND2xp5_ASAP7_75t_L g162 ( .A(n_103), .B(n_163), .Y(n_162) );
OA21x2_ASAP7_75t_L g105 ( .A1(n_106), .A2(n_111), .B(n_493), .Y(n_105) );
INVx1_ASAP7_75t_SL g106 ( .A(n_107), .Y(n_106) );
CKINVDCx5p33_ASAP7_75t_R g107 ( .A(n_108), .Y(n_107) );
CKINVDCx11_ASAP7_75t_R g108 ( .A(n_109), .Y(n_108) );
CKINVDCx8_ASAP7_75t_R g109 ( .A(n_110), .Y(n_109) );
OAI21xp5_ASAP7_75t_L g111 ( .A1(n_112), .A2(n_123), .B(n_489), .Y(n_111) );
CKINVDCx11_ASAP7_75t_R g112 ( .A(n_113), .Y(n_112) );
INVx1_ASAP7_75t_SL g113 ( .A(n_114), .Y(n_113) );
INVx1_ASAP7_75t_SL g114 ( .A(n_115), .Y(n_114) );
BUFx2_ASAP7_75t_L g115 ( .A(n_116), .Y(n_115) );
BUFx3_ASAP7_75t_L g492 ( .A(n_116), .Y(n_492) );
NAND2xp5_ASAP7_75t_L g116 ( .A(n_117), .B(n_118), .Y(n_116) );
HB1xp67_ASAP7_75t_L g507 ( .A(n_117), .Y(n_507) );
CKINVDCx16_ASAP7_75t_R g806 ( .A(n_117), .Y(n_806) );
OR2x2_ASAP7_75t_L g811 ( .A(n_117), .B(n_119), .Y(n_811) );
CKINVDCx5p33_ASAP7_75t_R g118 ( .A(n_119), .Y(n_118) );
AOI21xp5_ASAP7_75t_L g498 ( .A1(n_119), .A2(n_499), .B(n_808), .Y(n_498) );
NAND2xp5_ASAP7_75t_L g120 ( .A(n_121), .B(n_122), .Y(n_120) );
NOR2xp33_ASAP7_75t_L g820 ( .A(n_121), .B(n_122), .Y(n_820) );
AOI22xp33_ASAP7_75t_SL g123 ( .A1(n_124), .A2(n_125), .B1(n_132), .B2(n_133), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_125), .Y(n_124) );
OAI22xp5_ASAP7_75t_L g125 ( .A1(n_126), .A2(n_127), .B1(n_130), .B2(n_131), .Y(n_125) );
INVx1_ASAP7_75t_L g126 ( .A(n_127), .Y(n_126) );
NOR2xp33_ASAP7_75t_L g805 ( .A(n_129), .B(n_806), .Y(n_805) );
CKINVDCx5p33_ASAP7_75t_R g130 ( .A(n_131), .Y(n_130) );
INVx1_ASAP7_75t_L g132 ( .A(n_133), .Y(n_132) );
AND3x2_ASAP7_75t_L g133 ( .A(n_134), .B(n_379), .C(n_442), .Y(n_133) );
INVx1_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
OAI21xp5_ASAP7_75t_L g800 ( .A1(n_135), .A2(n_443), .B(n_801), .Y(n_800) );
NOR3xp33_ASAP7_75t_L g803 ( .A(n_135), .B(n_380), .C(n_804), .Y(n_803) );
NAND2xp5_ASAP7_75t_L g135 ( .A(n_136), .B(n_343), .Y(n_135) );
NOR3xp33_ASAP7_75t_L g136 ( .A(n_137), .B(n_284), .C(n_313), .Y(n_136) );
NAND2xp5_ASAP7_75t_SL g137 ( .A(n_138), .B(n_273), .Y(n_137) );
AOI22xp5_ASAP7_75t_L g138 ( .A1(n_139), .A2(n_189), .B1(n_231), .B2(n_243), .Y(n_138) );
NAND2x1_ASAP7_75t_L g428 ( .A(n_139), .B(n_274), .Y(n_428) );
INVx2_ASAP7_75t_SL g139 ( .A(n_140), .Y(n_139) );
OR2x2_ASAP7_75t_L g140 ( .A(n_141), .B(n_178), .Y(n_140) );
INVx2_ASAP7_75t_L g245 ( .A(n_141), .Y(n_245) );
INVx4_ASAP7_75t_L g289 ( .A(n_141), .Y(n_289) );
BUFx6f_ASAP7_75t_L g309 ( .A(n_141), .Y(n_309) );
AND2x4_ASAP7_75t_L g320 ( .A(n_141), .B(n_288), .Y(n_320) );
AND2x2_ASAP7_75t_L g326 ( .A(n_141), .B(n_248), .Y(n_326) );
NOR2x1_ASAP7_75t_SL g456 ( .A(n_141), .B(n_259), .Y(n_456) );
OR2x6_ASAP7_75t_L g141 ( .A(n_142), .B(n_147), .Y(n_141) );
OAI22xp5_ASAP7_75t_L g193 ( .A1(n_143), .A2(n_194), .B1(n_200), .B2(n_201), .Y(n_193) );
INVx3_ASAP7_75t_L g201 ( .A(n_143), .Y(n_201) );
INVx4_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
NAND2xp5_ASAP7_75t_L g203 ( .A(n_144), .B(n_204), .Y(n_203) );
AOI21x1_ASAP7_75t_L g570 ( .A1(n_144), .A2(n_571), .B(n_577), .Y(n_570) );
INVx3_ASAP7_75t_L g144 ( .A(n_145), .Y(n_144) );
BUFx4f_ASAP7_75t_L g221 ( .A(n_145), .Y(n_221) );
AND2x4_ASAP7_75t_L g176 ( .A(n_146), .B(n_177), .Y(n_176) );
AND2x2_ASAP7_75t_SL g181 ( .A(n_146), .B(n_177), .Y(n_181) );
AOI21xp5_ASAP7_75t_L g147 ( .A1(n_148), .A2(n_170), .B(n_176), .Y(n_147) );
INVxp67_ASAP7_75t_L g206 ( .A(n_149), .Y(n_206) );
AOI22xp5_ASAP7_75t_L g558 ( .A1(n_149), .A2(n_171), .B1(n_559), .B2(n_561), .Y(n_558) );
AND2x4_ASAP7_75t_L g149 ( .A(n_150), .B(n_155), .Y(n_149) );
NOR2x1p5_ASAP7_75t_L g150 ( .A(n_151), .B(n_152), .Y(n_150) );
INVx1_ASAP7_75t_L g228 ( .A(n_152), .Y(n_228) );
INVx3_ASAP7_75t_L g152 ( .A(n_153), .Y(n_152) );
OR2x6_ASAP7_75t_L g160 ( .A(n_153), .B(n_161), .Y(n_160) );
INVx2_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
AND2x6_ASAP7_75t_L g268 ( .A(n_154), .B(n_164), .Y(n_268) );
AND2x6_ASAP7_75t_L g519 ( .A(n_155), .B(n_175), .Y(n_519) );
AND2x2_ASAP7_75t_L g155 ( .A(n_156), .B(n_157), .Y(n_155) );
INVx2_ASAP7_75t_L g161 ( .A(n_156), .Y(n_161) );
AND2x4_ASAP7_75t_L g271 ( .A(n_156), .B(n_166), .Y(n_271) );
HB1xp67_ASAP7_75t_L g173 ( .A(n_157), .Y(n_173) );
O2A1O1Ixp33_ASAP7_75t_L g158 ( .A1(n_159), .A2(n_160), .B(n_162), .C(n_168), .Y(n_158) );
O2A1O1Ixp33_ASAP7_75t_SL g185 ( .A1(n_160), .A2(n_168), .B(n_186), .C(n_187), .Y(n_185) );
INVxp67_ASAP7_75t_L g195 ( .A(n_160), .Y(n_195) );
O2A1O1Ixp33_ASAP7_75t_L g214 ( .A1(n_160), .A2(n_168), .B(n_215), .C(n_216), .Y(n_214) );
O2A1O1Ixp33_ASAP7_75t_SL g239 ( .A1(n_160), .A2(n_168), .B(n_240), .C(n_241), .Y(n_239) );
INVx2_ASAP7_75t_L g258 ( .A(n_160), .Y(n_258) );
OAI22xp5_ASAP7_75t_L g262 ( .A1(n_160), .A2(n_198), .B1(n_263), .B2(n_264), .Y(n_262) );
AND2x2_ASAP7_75t_L g172 ( .A(n_161), .B(n_173), .Y(n_172) );
INVxp33_ASAP7_75t_L g227 ( .A(n_161), .Y(n_227) );
INVx1_ASAP7_75t_L g198 ( .A(n_163), .Y(n_198) );
AND2x4_ASAP7_75t_L g524 ( .A(n_163), .B(n_169), .Y(n_524) );
AND2x4_ASAP7_75t_L g163 ( .A(n_164), .B(n_166), .Y(n_163) );
INVx2_ASAP7_75t_L g164 ( .A(n_165), .Y(n_164) );
INVx2_ASAP7_75t_L g166 ( .A(n_167), .Y(n_166) );
INVx1_ASAP7_75t_L g224 ( .A(n_168), .Y(n_224) );
AOI21xp5_ASAP7_75t_L g255 ( .A1(n_168), .A2(n_256), .B(n_257), .Y(n_255) );
NOR2xp33_ASAP7_75t_L g272 ( .A(n_168), .B(n_176), .Y(n_272) );
AOI21xp5_ASAP7_75t_L g520 ( .A1(n_168), .A2(n_521), .B(n_522), .Y(n_520) );
AOI21xp5_ASAP7_75t_L g533 ( .A1(n_168), .A2(n_534), .B(n_535), .Y(n_533) );
AOI21xp5_ASAP7_75t_L g543 ( .A1(n_168), .A2(n_544), .B(n_545), .Y(n_543) );
AOI21xp5_ASAP7_75t_L g552 ( .A1(n_168), .A2(n_553), .B(n_554), .Y(n_552) );
AOI21xp5_ASAP7_75t_L g573 ( .A1(n_168), .A2(n_574), .B(n_575), .Y(n_573) );
AOI21xp5_ASAP7_75t_L g586 ( .A1(n_168), .A2(n_587), .B(n_588), .Y(n_586) );
INVx5_ASAP7_75t_L g168 ( .A(n_169), .Y(n_168) );
HB1xp67_ASAP7_75t_L g199 ( .A(n_169), .Y(n_199) );
INVx1_ASAP7_75t_L g208 ( .A(n_171), .Y(n_208) );
AND2x4_ASAP7_75t_L g171 ( .A(n_172), .B(n_174), .Y(n_171) );
INVx1_ASAP7_75t_L g251 ( .A(n_172), .Y(n_251) );
INVx1_ASAP7_75t_L g252 ( .A(n_174), .Y(n_252) );
BUFx3_ASAP7_75t_L g174 ( .A(n_175), .Y(n_174) );
AOI21xp5_ASAP7_75t_L g530 ( .A1(n_176), .A2(n_531), .B(n_532), .Y(n_530) );
NOR2xp33_ASAP7_75t_L g559 ( .A(n_176), .B(n_560), .Y(n_559) );
NOR2xp33_ASAP7_75t_L g561 ( .A(n_176), .B(n_562), .Y(n_561) );
NOR2xp33_ASAP7_75t_L g564 ( .A(n_176), .B(n_565), .Y(n_564) );
NOR3xp33_ASAP7_75t_L g566 ( .A(n_176), .B(n_198), .C(n_567), .Y(n_566) );
INVx2_ASAP7_75t_L g292 ( .A(n_178), .Y(n_292) );
HB1xp67_ASAP7_75t_L g306 ( .A(n_178), .Y(n_306) );
INVx1_ASAP7_75t_L g317 ( .A(n_178), .Y(n_317) );
HB1xp67_ASAP7_75t_L g329 ( .A(n_178), .Y(n_329) );
AND2x2_ASAP7_75t_L g361 ( .A(n_178), .B(n_259), .Y(n_361) );
AND2x2_ASAP7_75t_L g393 ( .A(n_178), .B(n_277), .Y(n_393) );
INVx1_ASAP7_75t_L g400 ( .A(n_178), .Y(n_400) );
AO21x2_ASAP7_75t_L g178 ( .A1(n_179), .A2(n_182), .B(n_188), .Y(n_178) );
AO21x2_ASAP7_75t_L g516 ( .A1(n_179), .A2(n_517), .B(n_525), .Y(n_516) );
AO21x2_ASAP7_75t_L g583 ( .A1(n_179), .A2(n_584), .B(n_590), .Y(n_583) );
AO21x2_ASAP7_75t_L g598 ( .A1(n_179), .A2(n_584), .B(n_590), .Y(n_598) );
CKINVDCx5p33_ASAP7_75t_R g179 ( .A(n_180), .Y(n_179) );
OA21x2_ASAP7_75t_L g541 ( .A1(n_180), .A2(n_542), .B(n_546), .Y(n_541) );
BUFx6f_ASAP7_75t_L g180 ( .A(n_181), .Y(n_180) );
NAND2xp5_ASAP7_75t_L g182 ( .A(n_183), .B(n_184), .Y(n_182) );
AND2x2_ASAP7_75t_L g189 ( .A(n_190), .B(n_209), .Y(n_189) );
INVx1_ASAP7_75t_L g190 ( .A(n_191), .Y(n_190) );
AND2x2_ASAP7_75t_L g342 ( .A(n_191), .B(n_281), .Y(n_342) );
INVx2_ASAP7_75t_L g416 ( .A(n_191), .Y(n_416) );
AND2x2_ASAP7_75t_L g439 ( .A(n_191), .B(n_209), .Y(n_439) );
INVx1_ASAP7_75t_L g191 ( .A(n_192), .Y(n_191) );
NAND2xp5_ASAP7_75t_L g280 ( .A(n_192), .B(n_234), .Y(n_280) );
INVx2_ASAP7_75t_L g301 ( .A(n_192), .Y(n_301) );
AND2x4_ASAP7_75t_L g323 ( .A(n_192), .B(n_324), .Y(n_323) );
INVx1_ASAP7_75t_L g358 ( .A(n_192), .Y(n_358) );
AND2x2_ASAP7_75t_L g435 ( .A(n_192), .B(n_237), .Y(n_435) );
OR2x2_ASAP7_75t_L g192 ( .A(n_193), .B(n_202), .Y(n_192) );
NOR2xp33_ASAP7_75t_L g196 ( .A(n_197), .B(n_198), .Y(n_196) );
AO21x2_ASAP7_75t_L g210 ( .A1(n_201), .A2(n_211), .B(n_217), .Y(n_210) );
AO21x2_ASAP7_75t_L g234 ( .A1(n_201), .A2(n_211), .B(n_217), .Y(n_234) );
OAI22xp5_ASAP7_75t_L g202 ( .A1(n_203), .A2(n_206), .B1(n_207), .B2(n_208), .Y(n_202) );
INVx1_ASAP7_75t_L g204 ( .A(n_205), .Y(n_204) );
INVx1_ASAP7_75t_L g406 ( .A(n_209), .Y(n_406) );
AND2x2_ASAP7_75t_L g209 ( .A(n_210), .B(n_218), .Y(n_209) );
NOR2xp67_ASAP7_75t_L g331 ( .A(n_210), .B(n_301), .Y(n_331) );
AND2x2_ASAP7_75t_L g336 ( .A(n_210), .B(n_301), .Y(n_336) );
INVx2_ASAP7_75t_L g349 ( .A(n_210), .Y(n_349) );
NOR2x1_ASAP7_75t_L g397 ( .A(n_210), .B(n_398), .Y(n_397) );
NAND2xp5_ASAP7_75t_L g211 ( .A(n_212), .B(n_213), .Y(n_211) );
AND2x4_ASAP7_75t_L g322 ( .A(n_218), .B(n_233), .Y(n_322) );
AND2x2_ASAP7_75t_L g337 ( .A(n_218), .B(n_338), .Y(n_337) );
INVx1_ASAP7_75t_L g390 ( .A(n_218), .Y(n_390) );
INVx2_ASAP7_75t_L g218 ( .A(n_219), .Y(n_218) );
NAND2xp5_ASAP7_75t_L g312 ( .A(n_219), .B(n_237), .Y(n_312) );
NAND2xp5_ASAP7_75t_L g394 ( .A(n_219), .B(n_234), .Y(n_394) );
AO21x2_ASAP7_75t_L g219 ( .A1(n_220), .A2(n_222), .B(n_230), .Y(n_219) );
AO21x2_ASAP7_75t_L g283 ( .A1(n_220), .A2(n_222), .B(n_230), .Y(n_283) );
AOI21x1_ASAP7_75t_L g622 ( .A1(n_220), .A2(n_623), .B(n_626), .Y(n_622) );
INVx2_ASAP7_75t_SL g220 ( .A(n_221), .Y(n_220) );
OA21x2_ASAP7_75t_L g237 ( .A1(n_221), .A2(n_238), .B(n_242), .Y(n_237) );
AOI21xp5_ASAP7_75t_L g549 ( .A1(n_221), .A2(n_550), .B(n_551), .Y(n_549) );
NAND2xp5_ASAP7_75t_SL g222 ( .A(n_223), .B(n_229), .Y(n_222) );
INVx1_ASAP7_75t_L g225 ( .A(n_226), .Y(n_225) );
INVxp33_ASAP7_75t_L g231 ( .A(n_232), .Y(n_231) );
NAND2x1p5_ASAP7_75t_L g232 ( .A(n_233), .B(n_235), .Y(n_232) );
INVx3_ASAP7_75t_L g298 ( .A(n_233), .Y(n_298) );
INVx3_ASAP7_75t_L g233 ( .A(n_234), .Y(n_233) );
HB1xp67_ASAP7_75t_L g296 ( .A(n_234), .Y(n_296) );
AND2x2_ASAP7_75t_L g465 ( .A(n_234), .B(n_466), .Y(n_465) );
INVx3_ASAP7_75t_L g353 ( .A(n_235), .Y(n_353) );
NAND2xp5_ASAP7_75t_L g485 ( .A(n_235), .B(n_390), .Y(n_485) );
BUFx3_ASAP7_75t_L g235 ( .A(n_236), .Y(n_235) );
AND2x2_ASAP7_75t_L g300 ( .A(n_236), .B(n_301), .Y(n_300) );
INVx1_ASAP7_75t_L g236 ( .A(n_237), .Y(n_236) );
AND2x4_ASAP7_75t_L g281 ( .A(n_237), .B(n_282), .Y(n_281) );
INVx2_ASAP7_75t_L g324 ( .A(n_237), .Y(n_324) );
INVxp67_ASAP7_75t_L g338 ( .A(n_237), .Y(n_338) );
INVx1_ASAP7_75t_L g398 ( .A(n_237), .Y(n_398) );
HB1xp67_ASAP7_75t_L g466 ( .A(n_237), .Y(n_466) );
INVx1_ASAP7_75t_L g450 ( .A(n_243), .Y(n_450) );
NOR2x1_ASAP7_75t_L g243 ( .A(n_244), .B(n_246), .Y(n_243) );
NOR2x1_ASAP7_75t_L g370 ( .A(n_244), .B(n_371), .Y(n_370) );
INVx1_ASAP7_75t_L g244 ( .A(n_245), .Y(n_244) );
AND2x2_ASAP7_75t_L g404 ( .A(n_245), .B(n_276), .Y(n_404) );
OR2x2_ASAP7_75t_L g440 ( .A(n_246), .B(n_441), .Y(n_440) );
INVx2_ASAP7_75t_L g246 ( .A(n_247), .Y(n_246) );
AND2x2_ASAP7_75t_L g422 ( .A(n_247), .B(n_400), .Y(n_422) );
AND2x2_ASAP7_75t_L g474 ( .A(n_247), .B(n_309), .Y(n_474) );
AND2x2_ASAP7_75t_L g247 ( .A(n_248), .B(n_259), .Y(n_247) );
AND2x4_ASAP7_75t_L g276 ( .A(n_248), .B(n_277), .Y(n_276) );
INVx1_ASAP7_75t_L g288 ( .A(n_248), .Y(n_288) );
INVx2_ASAP7_75t_L g305 ( .A(n_248), .Y(n_305) );
HB1xp67_ASAP7_75t_L g483 ( .A(n_248), .Y(n_483) );
AND2x2_ASAP7_75t_L g248 ( .A(n_249), .B(n_254), .Y(n_248) );
NOR3xp33_ASAP7_75t_L g250 ( .A(n_251), .B(n_252), .C(n_253), .Y(n_250) );
INVx3_ASAP7_75t_L g277 ( .A(n_259), .Y(n_277) );
INVx2_ASAP7_75t_L g371 ( .A(n_259), .Y(n_371) );
AND2x4_ASAP7_75t_L g259 ( .A(n_260), .B(n_261), .Y(n_259) );
OAI21xp5_ASAP7_75t_L g261 ( .A1(n_262), .A2(n_265), .B(n_272), .Y(n_261) );
OAI22xp5_ASAP7_75t_L g265 ( .A1(n_266), .A2(n_267), .B1(n_269), .B2(n_270), .Y(n_265) );
INVxp67_ASAP7_75t_L g267 ( .A(n_268), .Y(n_267) );
INVxp67_ASAP7_75t_L g270 ( .A(n_271), .Y(n_270) );
NAND2xp5_ASAP7_75t_L g273 ( .A(n_274), .B(n_278), .Y(n_273) );
INVx2_ASAP7_75t_L g274 ( .A(n_275), .Y(n_274) );
NOR2xp33_ASAP7_75t_L g368 ( .A(n_275), .B(n_351), .Y(n_368) );
NOR2x1_ASAP7_75t_L g410 ( .A(n_275), .B(n_289), .Y(n_410) );
INVx4_ASAP7_75t_L g275 ( .A(n_276), .Y(n_275) );
NAND2xp5_ASAP7_75t_L g488 ( .A(n_276), .B(n_351), .Y(n_488) );
AND2x2_ASAP7_75t_L g304 ( .A(n_277), .B(n_305), .Y(n_304) );
INVx1_ASAP7_75t_L g318 ( .A(n_277), .Y(n_318) );
AOI22xp5_ASAP7_75t_SL g366 ( .A1(n_278), .A2(n_367), .B1(n_368), .B2(n_369), .Y(n_366) );
AND2x2_ASAP7_75t_L g278 ( .A(n_279), .B(n_281), .Y(n_278) );
NAND2x1p5_ASAP7_75t_L g363 ( .A(n_279), .B(n_337), .Y(n_363) );
INVx2_ASAP7_75t_SL g279 ( .A(n_280), .Y(n_279) );
OR2x2_ASAP7_75t_L g424 ( .A(n_280), .B(n_312), .Y(n_424) );
AND2x2_ASAP7_75t_L g294 ( .A(n_281), .B(n_295), .Y(n_294) );
AND2x4_ASAP7_75t_L g330 ( .A(n_281), .B(n_331), .Y(n_330) );
AND2x2_ASAP7_75t_L g426 ( .A(n_281), .B(n_416), .Y(n_426) );
INVx2_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
AND2x4_ASAP7_75t_L g348 ( .A(n_283), .B(n_349), .Y(n_348) );
INVx1_ASAP7_75t_L g374 ( .A(n_283), .Y(n_374) );
AND2x2_ASAP7_75t_L g464 ( .A(n_283), .B(n_301), .Y(n_464) );
OAI221xp5_ASAP7_75t_L g284 ( .A1(n_285), .A2(n_293), .B1(n_297), .B2(n_302), .C(n_307), .Y(n_284) );
INVx1_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
AND2x2_ASAP7_75t_L g286 ( .A(n_287), .B(n_290), .Y(n_286) );
INVx1_ASAP7_75t_L g365 ( .A(n_287), .Y(n_365) );
NAND2xp5_ASAP7_75t_L g392 ( .A(n_287), .B(n_393), .Y(n_392) );
NAND2xp5_ASAP7_75t_L g480 ( .A(n_287), .B(n_361), .Y(n_480) );
AND2x4_ASAP7_75t_L g287 ( .A(n_288), .B(n_289), .Y(n_287) );
NOR2xp67_ASAP7_75t_SL g333 ( .A(n_289), .B(n_334), .Y(n_333) );
HB1xp67_ASAP7_75t_L g346 ( .A(n_289), .Y(n_346) );
OR2x2_ASAP7_75t_L g430 ( .A(n_289), .B(n_431), .Y(n_430) );
AND2x4_ASAP7_75t_SL g482 ( .A(n_289), .B(n_483), .Y(n_482) );
HB1xp67_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
INVx3_ASAP7_75t_L g351 ( .A(n_291), .Y(n_351) );
INVx2_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
HB1xp67_ASAP7_75t_L g441 ( .A(n_292), .Y(n_441) );
INVx1_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
AOI221x1_ASAP7_75t_L g381 ( .A1(n_294), .A2(n_382), .B1(n_384), .B2(n_387), .C(n_391), .Y(n_381) );
AND2x2_ASAP7_75t_L g367 ( .A(n_295), .B(n_323), .Y(n_367) );
INVx1_ASAP7_75t_L g295 ( .A(n_296), .Y(n_295) );
OR2x2_ASAP7_75t_L g297 ( .A(n_298), .B(n_299), .Y(n_297) );
AND2x2_ASAP7_75t_L g310 ( .A(n_298), .B(n_311), .Y(n_310) );
NAND2xp5_ASAP7_75t_L g437 ( .A(n_298), .B(n_300), .Y(n_437) );
INVx2_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
INVx2_ASAP7_75t_L g302 ( .A(n_303), .Y(n_302) );
AND2x2_ASAP7_75t_L g303 ( .A(n_304), .B(n_306), .Y(n_303) );
AND2x2_ASAP7_75t_SL g308 ( .A(n_304), .B(n_309), .Y(n_308) );
NAND2xp5_ASAP7_75t_L g334 ( .A(n_304), .B(n_317), .Y(n_334) );
INVx2_ASAP7_75t_L g341 ( .A(n_304), .Y(n_341) );
INVx1_ASAP7_75t_L g386 ( .A(n_305), .Y(n_386) );
BUFx2_ASAP7_75t_L g475 ( .A(n_306), .Y(n_475) );
NAND2xp33_ASAP7_75t_SL g307 ( .A(n_308), .B(n_310), .Y(n_307) );
OR2x6_ASAP7_75t_L g340 ( .A(n_309), .B(n_341), .Y(n_340) );
AND2x2_ASAP7_75t_L g421 ( .A(n_309), .B(n_361), .Y(n_421) );
INVx2_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
NAND2xp5_ASAP7_75t_L g313 ( .A(n_314), .B(n_332), .Y(n_313) );
AOI22xp5_ASAP7_75t_L g314 ( .A1(n_315), .A2(n_321), .B1(n_325), .B2(n_330), .Y(n_314) );
NOR2xp33_ASAP7_75t_L g315 ( .A(n_316), .B(n_319), .Y(n_315) );
AND2x2_ASAP7_75t_SL g378 ( .A(n_316), .B(n_320), .Y(n_378) );
AND2x4_ASAP7_75t_L g384 ( .A(n_316), .B(n_385), .Y(n_384) );
AND2x4_ASAP7_75t_SL g316 ( .A(n_317), .B(n_318), .Y(n_316) );
HB1xp67_ASAP7_75t_L g409 ( .A(n_317), .Y(n_409) );
INVx2_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
NOR2xp33_ASAP7_75t_L g359 ( .A(n_320), .B(n_360), .Y(n_359) );
NAND2xp5_ASAP7_75t_L g383 ( .A(n_320), .B(n_351), .Y(n_383) );
HB1xp67_ASAP7_75t_L g467 ( .A(n_320), .Y(n_467) );
AND2x2_ASAP7_75t_L g321 ( .A(n_322), .B(n_323), .Y(n_321) );
AND2x2_ASAP7_75t_L g414 ( .A(n_322), .B(n_415), .Y(n_414) );
INVx3_ASAP7_75t_L g375 ( .A(n_323), .Y(n_375) );
NAND2x1_ASAP7_75t_SL g419 ( .A(n_323), .B(n_374), .Y(n_419) );
AND2x2_ASAP7_75t_L g453 ( .A(n_323), .B(n_348), .Y(n_453) );
AND2x2_ASAP7_75t_L g325 ( .A(n_326), .B(n_327), .Y(n_325) );
INVx1_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
INVx1_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
AOI22xp5_ASAP7_75t_L g332 ( .A1(n_333), .A2(n_335), .B1(n_339), .B2(n_342), .Y(n_332) );
BUFx2_ASAP7_75t_L g448 ( .A(n_334), .Y(n_448) );
AOI22xp33_ASAP7_75t_L g486 ( .A1(n_335), .A2(n_404), .B1(n_478), .B2(n_487), .Y(n_486) );
AND2x2_ASAP7_75t_L g335 ( .A(n_336), .B(n_337), .Y(n_335) );
NAND2x1p5_ASAP7_75t_L g389 ( .A(n_336), .B(n_390), .Y(n_389) );
AND2x2_ASAP7_75t_L g356 ( .A(n_337), .B(n_357), .Y(n_356) );
INVx2_ASAP7_75t_L g339 ( .A(n_340), .Y(n_339) );
NAND3xp33_ASAP7_75t_L g472 ( .A(n_341), .B(n_473), .C(n_475), .Y(n_472) );
INVx1_ASAP7_75t_L g376 ( .A(n_342), .Y(n_376) );
AOI211x1_ASAP7_75t_L g343 ( .A1(n_344), .A2(n_352), .B(n_354), .C(n_372), .Y(n_343) );
INVx1_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
NAND2xp5_ASAP7_75t_L g345 ( .A(n_346), .B(n_347), .Y(n_345) );
NAND2xp5_ASAP7_75t_SL g403 ( .A(n_347), .B(n_404), .Y(n_403) );
AND2x2_ASAP7_75t_L g347 ( .A(n_348), .B(n_350), .Y(n_347) );
AND2x2_ASAP7_75t_L g434 ( .A(n_348), .B(n_435), .Y(n_434) );
NAND2xp5_ASAP7_75t_L g446 ( .A(n_348), .B(n_415), .Y(n_446) );
AND2x2_ASAP7_75t_L g478 ( .A(n_348), .B(n_416), .Y(n_478) );
INVx1_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
INVx1_ASAP7_75t_L g459 ( .A(n_351), .Y(n_459) );
INVx1_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
OR2x2_ASAP7_75t_L g388 ( .A(n_353), .B(n_389), .Y(n_388) );
NAND2xp5_ASAP7_75t_L g354 ( .A(n_355), .B(n_366), .Y(n_354) );
AOI22xp5_ASAP7_75t_SL g355 ( .A1(n_356), .A2(n_359), .B1(n_362), .B2(n_364), .Y(n_355) );
BUFx2_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
AND2x2_ASAP7_75t_L g396 ( .A(n_358), .B(n_397), .Y(n_396) );
INVx1_ASAP7_75t_SL g411 ( .A(n_358), .Y(n_411) );
INVx1_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
AND2x2_ASAP7_75t_SL g481 ( .A(n_361), .B(n_482), .Y(n_481) );
INVx3_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
INVxp67_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
HB1xp67_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
AND2x2_ASAP7_75t_L g417 ( .A(n_370), .B(n_400), .Y(n_417) );
AOI21xp5_ASAP7_75t_L g372 ( .A1(n_373), .A2(n_376), .B(n_377), .Y(n_372) );
OR2x2_ASAP7_75t_L g373 ( .A(n_374), .B(n_375), .Y(n_373) );
NAND2xp5_ASAP7_75t_L g471 ( .A(n_374), .B(n_396), .Y(n_471) );
OR2x2_ASAP7_75t_L g449 ( .A(n_375), .B(n_394), .Y(n_449) );
INVx1_ASAP7_75t_SL g377 ( .A(n_378), .Y(n_377) );
INVx1_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
NAND2xp33_ASAP7_75t_L g802 ( .A(n_380), .B(n_801), .Y(n_802) );
NAND3x1_ASAP7_75t_L g380 ( .A(n_381), .B(n_401), .C(n_425), .Y(n_380) );
INVx1_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
AOI22xp5_ASAP7_75t_L g413 ( .A1(n_384), .A2(n_414), .B1(n_417), .B2(n_418), .Y(n_413) );
NAND2xp5_ASAP7_75t_SL g399 ( .A(n_385), .B(n_400), .Y(n_399) );
INVx2_ASAP7_75t_SL g458 ( .A(n_385), .Y(n_458) );
NAND2xp5_ASAP7_75t_L g462 ( .A(n_385), .B(n_459), .Y(n_462) );
INVx2_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
INVx1_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
OAI222xp33_ASAP7_75t_L g445 ( .A1(n_389), .A2(n_446), .B1(n_447), .B2(n_448), .C1(n_449), .C2(n_450), .Y(n_445) );
OAI22xp5_ASAP7_75t_L g391 ( .A1(n_392), .A2(n_394), .B1(n_395), .B2(n_399), .Y(n_391) );
INVx1_ASAP7_75t_SL g431 ( .A(n_393), .Y(n_431) );
INVx1_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
AND2x2_ASAP7_75t_L g468 ( .A(n_397), .B(n_464), .Y(n_468) );
NOR2x1_ASAP7_75t_L g401 ( .A(n_402), .B(n_412), .Y(n_401) );
AOI21xp5_ASAP7_75t_SL g402 ( .A1(n_403), .A2(n_405), .B(n_411), .Y(n_402) );
NAND2xp5_ASAP7_75t_L g405 ( .A(n_406), .B(n_407), .Y(n_405) );
INVx1_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
NAND2xp5_ASAP7_75t_L g408 ( .A(n_409), .B(n_410), .Y(n_408) );
NAND2xp5_ASAP7_75t_L g412 ( .A(n_413), .B(n_420), .Y(n_412) );
INVx1_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
INVx2_ASAP7_75t_SL g418 ( .A(n_419), .Y(n_418) );
NAND2xp5_ASAP7_75t_L g432 ( .A(n_419), .B(n_433), .Y(n_432) );
OAI21xp5_ASAP7_75t_SL g420 ( .A1(n_421), .A2(n_422), .B(n_423), .Y(n_420) );
INVx1_ASAP7_75t_L g447 ( .A(n_422), .Y(n_447) );
INVx1_ASAP7_75t_SL g423 ( .A(n_424), .Y(n_423) );
AOI221xp5_ASAP7_75t_L g425 ( .A1(n_426), .A2(n_427), .B1(n_429), .B2(n_432), .C(n_436), .Y(n_425) );
INVx1_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
INVxp67_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
INVx2_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
AOI21xp5_ASAP7_75t_L g436 ( .A1(n_437), .A2(n_438), .B(n_440), .Y(n_436) );
INVx1_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
INVxp67_ASAP7_75t_SL g442 ( .A(n_443), .Y(n_442) );
NAND3x1_ASAP7_75t_L g443 ( .A(n_444), .B(n_469), .C(n_476), .Y(n_443) );
NAND4xp25_ASAP7_75t_L g804 ( .A(n_444), .B(n_469), .C(n_476), .D(n_805), .Y(n_804) );
NOR2x1_ASAP7_75t_L g444 ( .A(n_445), .B(n_451), .Y(n_444) );
NAND2xp5_ASAP7_75t_L g451 ( .A(n_452), .B(n_460), .Y(n_451) );
NAND2xp5_ASAP7_75t_SL g452 ( .A(n_453), .B(n_454), .Y(n_452) );
NAND2xp5_ASAP7_75t_L g454 ( .A(n_455), .B(n_457), .Y(n_454) );
NAND2xp5_ASAP7_75t_L g461 ( .A(n_455), .B(n_462), .Y(n_461) );
INVx1_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
NAND2xp5_ASAP7_75t_L g457 ( .A(n_458), .B(n_459), .Y(n_457) );
AOI22xp5_ASAP7_75t_L g460 ( .A1(n_461), .A2(n_463), .B1(n_467), .B2(n_468), .Y(n_460) );
AND2x4_ASAP7_75t_L g463 ( .A(n_464), .B(n_465), .Y(n_463) );
NAND2xp5_ASAP7_75t_SL g469 ( .A(n_470), .B(n_472), .Y(n_469) );
INVx1_ASAP7_75t_L g470 ( .A(n_471), .Y(n_470) );
INVx1_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
AND2x2_ASAP7_75t_L g476 ( .A(n_477), .B(n_486), .Y(n_476) );
AOI22xp5_ASAP7_75t_SL g477 ( .A1(n_478), .A2(n_479), .B1(n_481), .B2(n_484), .Y(n_477) );
INVx1_ASAP7_75t_L g479 ( .A(n_480), .Y(n_479) );
INVxp67_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
INVx1_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
AND2x2_ASAP7_75t_L g494 ( .A(n_489), .B(n_495), .Y(n_494) );
INVx1_ASAP7_75t_L g490 ( .A(n_491), .Y(n_490) );
HB1xp67_ASAP7_75t_L g491 ( .A(n_492), .Y(n_491) );
NAND2xp5_ASAP7_75t_L g493 ( .A(n_494), .B(n_498), .Y(n_493) );
CKINVDCx5p33_ASAP7_75t_R g495 ( .A(n_496), .Y(n_495) );
CKINVDCx20_ASAP7_75t_R g496 ( .A(n_497), .Y(n_496) );
OAI22xp5_ASAP7_75t_L g499 ( .A1(n_500), .A2(n_501), .B1(n_506), .B2(n_807), .Y(n_499) );
INVxp33_ASAP7_75t_L g500 ( .A(n_501), .Y(n_500) );
INVx1_ASAP7_75t_L g505 ( .A(n_503), .Y(n_505) );
INVx2_ASAP7_75t_L g807 ( .A(n_506), .Y(n_807) );
OAI21x1_ASAP7_75t_L g506 ( .A1(n_507), .A2(n_508), .B(n_798), .Y(n_506) );
AND2x4_ASAP7_75t_L g508 ( .A(n_509), .B(n_737), .Y(n_508) );
NOR3xp33_ASAP7_75t_L g509 ( .A(n_510), .B(n_630), .C(n_681), .Y(n_509) );
OAI211xp5_ASAP7_75t_SL g510 ( .A1(n_511), .A2(n_536), .B(n_578), .C(n_609), .Y(n_510) );
INVxp67_ASAP7_75t_L g511 ( .A(n_512), .Y(n_511) );
NOR2xp33_ASAP7_75t_L g512 ( .A(n_513), .B(n_526), .Y(n_512) );
INVx1_ASAP7_75t_L g513 ( .A(n_514), .Y(n_513) );
HB1xp67_ASAP7_75t_L g514 ( .A(n_515), .Y(n_514) );
NAND2xp5_ASAP7_75t_L g745 ( .A(n_515), .B(n_583), .Y(n_745) );
INVx1_ASAP7_75t_L g515 ( .A(n_516), .Y(n_515) );
AND2x2_ASAP7_75t_L g591 ( .A(n_516), .B(n_528), .Y(n_591) );
NAND2xp5_ASAP7_75t_L g597 ( .A(n_516), .B(n_598), .Y(n_597) );
OR2x2_ASAP7_75t_L g608 ( .A(n_516), .B(n_598), .Y(n_608) );
NAND2xp5_ASAP7_75t_L g628 ( .A(n_516), .B(n_629), .Y(n_628) );
AND2x2_ASAP7_75t_L g644 ( .A(n_516), .B(n_621), .Y(n_644) );
INVx2_ASAP7_75t_L g670 ( .A(n_516), .Y(n_670) );
AND2x4_ASAP7_75t_L g679 ( .A(n_516), .B(n_680), .Y(n_679) );
AND2x2_ASAP7_75t_L g784 ( .A(n_516), .B(n_651), .Y(n_784) );
NAND2xp5_ASAP7_75t_L g517 ( .A(n_518), .B(n_523), .Y(n_517) );
AND2x2_ASAP7_75t_L g668 ( .A(n_526), .B(n_669), .Y(n_668) );
OAI32xp33_ASAP7_75t_L g751 ( .A1(n_526), .A2(n_673), .A3(n_677), .B1(n_684), .B2(n_752), .Y(n_751) );
NAND2xp5_ASAP7_75t_L g783 ( .A(n_526), .B(n_784), .Y(n_783) );
INVx2_ASAP7_75t_L g526 ( .A(n_527), .Y(n_526) );
AND2x2_ASAP7_75t_L g606 ( .A(n_527), .B(n_607), .Y(n_606) );
NAND3xp33_ASAP7_75t_L g678 ( .A(n_527), .B(n_601), .C(n_679), .Y(n_678) );
OR2x2_ASAP7_75t_L g704 ( .A(n_527), .B(n_608), .Y(n_704) );
INVx2_ASAP7_75t_L g527 ( .A(n_528), .Y(n_527) );
HB1xp67_ASAP7_75t_L g595 ( .A(n_528), .Y(n_595) );
INVx5_ASAP7_75t_L g629 ( .A(n_528), .Y(n_629) );
AND2x4_ASAP7_75t_L g685 ( .A(n_528), .B(n_598), .Y(n_685) );
OR2x2_ASAP7_75t_L g700 ( .A(n_528), .B(n_621), .Y(n_700) );
OR2x2_ASAP7_75t_L g726 ( .A(n_528), .B(n_583), .Y(n_726) );
AND2x2_ASAP7_75t_L g734 ( .A(n_528), .B(n_680), .Y(n_734) );
AND2x4_ASAP7_75t_SL g759 ( .A(n_528), .B(n_679), .Y(n_759) );
OR2x6_ASAP7_75t_L g528 ( .A(n_529), .B(n_530), .Y(n_528) );
INVx1_ASAP7_75t_L g536 ( .A(n_537), .Y(n_536) );
NAND2xp5_ASAP7_75t_L g755 ( .A(n_537), .B(n_679), .Y(n_755) );
AND2x2_ASAP7_75t_L g537 ( .A(n_538), .B(n_547), .Y(n_537) );
NAND2xp5_ASAP7_75t_L g653 ( .A(n_538), .B(n_654), .Y(n_653) );
INVx1_ASAP7_75t_L g538 ( .A(n_539), .Y(n_538) );
OR2x6_ASAP7_75t_SL g580 ( .A(n_539), .B(n_581), .Y(n_580) );
INVxp67_ASAP7_75t_SL g539 ( .A(n_540), .Y(n_539) );
INVx1_ASAP7_75t_L g605 ( .A(n_540), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g657 ( .A(n_540), .B(n_639), .Y(n_657) );
HB1xp67_ASAP7_75t_L g795 ( .A(n_540), .Y(n_795) );
INVx1_ASAP7_75t_L g540 ( .A(n_541), .Y(n_540) );
INVx2_ASAP7_75t_L g613 ( .A(n_541), .Y(n_613) );
AND2x2_ASAP7_75t_L g637 ( .A(n_541), .B(n_569), .Y(n_637) );
INVx2_ASAP7_75t_L g665 ( .A(n_541), .Y(n_665) );
NAND2xp5_ASAP7_75t_L g706 ( .A(n_541), .B(n_548), .Y(n_706) );
BUFx3_ASAP7_75t_L g730 ( .A(n_541), .Y(n_730) );
OR2x2_ASAP7_75t_L g742 ( .A(n_541), .B(n_548), .Y(n_742) );
HB1xp67_ASAP7_75t_L g750 ( .A(n_541), .Y(n_750) );
AOI22xp5_ASAP7_75t_L g772 ( .A1(n_547), .A2(n_773), .B1(n_776), .B2(n_777), .Y(n_772) );
AND2x2_ASAP7_75t_L g547 ( .A(n_548), .B(n_556), .Y(n_547) );
INVx1_ASAP7_75t_L g601 ( .A(n_548), .Y(n_601) );
OR2x2_ASAP7_75t_L g612 ( .A(n_548), .B(n_613), .Y(n_612) );
INVx2_ASAP7_75t_L g619 ( .A(n_548), .Y(n_619) );
AND2x4_ASAP7_75t_SL g635 ( .A(n_548), .B(n_557), .Y(n_635) );
AND2x4_ASAP7_75t_L g640 ( .A(n_548), .B(n_641), .Y(n_640) );
INVx2_ASAP7_75t_L g649 ( .A(n_548), .Y(n_649) );
OR2x2_ASAP7_75t_L g655 ( .A(n_548), .B(n_557), .Y(n_655) );
OR2x2_ASAP7_75t_L g656 ( .A(n_548), .B(n_657), .Y(n_656) );
HB1xp67_ASAP7_75t_L g767 ( .A(n_548), .Y(n_767) );
NAND2xp5_ASAP7_75t_L g771 ( .A(n_548), .B(n_637), .Y(n_771) );
OR2x2_ASAP7_75t_L g787 ( .A(n_548), .B(n_690), .Y(n_787) );
OR2x6_ASAP7_75t_L g548 ( .A(n_549), .B(n_555), .Y(n_548) );
NAND2xp5_ASAP7_75t_L g600 ( .A(n_556), .B(n_601), .Y(n_600) );
INVx1_ASAP7_75t_L g614 ( .A(n_556), .Y(n_614) );
AND2x2_ASAP7_75t_SL g720 ( .A(n_556), .B(n_605), .Y(n_720) );
AND2x4_ASAP7_75t_L g556 ( .A(n_557), .B(n_568), .Y(n_556) );
NAND2xp5_ASAP7_75t_L g581 ( .A(n_557), .B(n_569), .Y(n_581) );
NOR2xp33_ASAP7_75t_L g602 ( .A(n_557), .B(n_603), .Y(n_602) );
NAND2xp5_ASAP7_75t_L g617 ( .A(n_557), .B(n_613), .Y(n_617) );
INVx3_ASAP7_75t_L g641 ( .A(n_557), .Y(n_641) );
INVx1_ASAP7_75t_L g674 ( .A(n_557), .Y(n_674) );
AND2x2_ASAP7_75t_L g754 ( .A(n_557), .B(n_619), .Y(n_754) );
AND2x4_ASAP7_75t_L g557 ( .A(n_558), .B(n_563), .Y(n_557) );
INVx2_ASAP7_75t_L g568 ( .A(n_569), .Y(n_568) );
NAND2xp5_ASAP7_75t_L g618 ( .A(n_569), .B(n_619), .Y(n_618) );
INVx1_ASAP7_75t_L g639 ( .A(n_569), .Y(n_639) );
AND2x2_ASAP7_75t_L g664 ( .A(n_569), .B(n_665), .Y(n_664) );
OR2x2_ASAP7_75t_L g690 ( .A(n_569), .B(n_613), .Y(n_690) );
NAND2xp5_ASAP7_75t_L g707 ( .A(n_569), .B(n_641), .Y(n_707) );
INVx1_ASAP7_75t_L g713 ( .A(n_569), .Y(n_713) );
INVx3_ASAP7_75t_L g569 ( .A(n_570), .Y(n_569) );
NAND2xp5_ASAP7_75t_L g571 ( .A(n_572), .B(n_576), .Y(n_571) );
AOI222xp33_ASAP7_75t_SL g578 ( .A1(n_579), .A2(n_582), .B1(n_592), .B2(n_599), .C1(n_602), .C2(n_606), .Y(n_578) );
CKINVDCx16_ASAP7_75t_R g579 ( .A(n_580), .Y(n_579) );
AND2x2_ASAP7_75t_L g582 ( .A(n_583), .B(n_591), .Y(n_582) );
NOR2xp33_ASAP7_75t_L g702 ( .A(n_583), .B(n_651), .Y(n_702) );
AND2x4_ASAP7_75t_L g718 ( .A(n_583), .B(n_629), .Y(n_718) );
NAND2xp5_ASAP7_75t_L g584 ( .A(n_585), .B(n_589), .Y(n_584) );
INVx2_ASAP7_75t_L g592 ( .A(n_593), .Y(n_592) );
NAND2xp5_ASAP7_75t_SL g593 ( .A(n_594), .B(n_596), .Y(n_593) );
INVx1_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
AND2x2_ASAP7_75t_L g643 ( .A(n_595), .B(n_644), .Y(n_643) );
AOI222xp33_ASAP7_75t_L g609 ( .A1(n_596), .A2(n_610), .B1(n_615), .B2(n_620), .C1(n_627), .C2(n_822), .Y(n_609) );
INVx1_ASAP7_75t_L g596 ( .A(n_597), .Y(n_596) );
OR2x2_ASAP7_75t_L g747 ( .A(n_597), .B(n_651), .Y(n_747) );
OR2x2_ASAP7_75t_L g790 ( .A(n_597), .B(n_696), .Y(n_790) );
AND2x2_ASAP7_75t_L g620 ( .A(n_598), .B(n_621), .Y(n_620) );
INVx2_ASAP7_75t_L g680 ( .A(n_598), .Y(n_680) );
HB1xp67_ASAP7_75t_L g695 ( .A(n_598), .Y(n_695) );
O2A1O1Ixp33_ASAP7_75t_L g708 ( .A1(n_599), .A2(n_709), .B(n_714), .C(n_715), .Y(n_708) );
INVx1_ASAP7_75t_SL g599 ( .A(n_600), .Y(n_599) );
INVx1_ASAP7_75t_L g736 ( .A(n_601), .Y(n_736) );
INVx1_ASAP7_75t_L g603 ( .A(n_604), .Y(n_603) );
HB1xp67_ASAP7_75t_L g604 ( .A(n_605), .Y(n_604) );
INVx2_ASAP7_75t_L g666 ( .A(n_606), .Y(n_666) );
AND2x2_ASAP7_75t_L g650 ( .A(n_607), .B(n_651), .Y(n_650) );
AND2x2_ASAP7_75t_L g659 ( .A(n_607), .B(n_660), .Y(n_659) );
INVx2_ASAP7_75t_L g607 ( .A(n_608), .Y(n_607) );
OAI31xp33_ASAP7_75t_L g701 ( .A1(n_610), .A2(n_627), .A3(n_702), .B(n_703), .Y(n_701) );
INVx1_ASAP7_75t_L g610 ( .A(n_611), .Y(n_610) );
A2O1A1Ixp33_ASAP7_75t_L g703 ( .A1(n_611), .A2(n_660), .B(n_704), .C(n_705), .Y(n_703) );
OR2x2_ASAP7_75t_L g611 ( .A(n_612), .B(n_614), .Y(n_611) );
OR2x2_ASAP7_75t_L g692 ( .A(n_612), .B(n_641), .Y(n_692) );
INVx2_ASAP7_75t_SL g615 ( .A(n_616), .Y(n_615) );
OR2x2_ASAP7_75t_L g616 ( .A(n_617), .B(n_618), .Y(n_616) );
BUFx2_ASAP7_75t_L g660 ( .A(n_621), .Y(n_660) );
AND2x2_ASAP7_75t_L g669 ( .A(n_621), .B(n_670), .Y(n_669) );
INVx2_ASAP7_75t_L g621 ( .A(n_622), .Y(n_621) );
BUFx6f_ASAP7_75t_L g651 ( .A(n_622), .Y(n_651) );
NAND2xp5_ASAP7_75t_L g623 ( .A(n_624), .B(n_625), .Y(n_623) );
INVx1_ASAP7_75t_L g627 ( .A(n_628), .Y(n_627) );
NAND2xp5_ASAP7_75t_L g778 ( .A(n_629), .B(n_686), .Y(n_778) );
OAI211xp5_ASAP7_75t_L g630 ( .A1(n_631), .A2(n_642), .B(n_645), .C(n_667), .Y(n_630) );
INVxp33_ASAP7_75t_L g631 ( .A(n_632), .Y(n_631) );
NAND2xp5_ASAP7_75t_SL g632 ( .A(n_633), .B(n_638), .Y(n_632) );
OR2x2_ASAP7_75t_L g633 ( .A(n_634), .B(n_636), .Y(n_633) );
INVx1_ASAP7_75t_SL g634 ( .A(n_635), .Y(n_634) );
AND2x2_ASAP7_75t_L g671 ( .A(n_635), .B(n_664), .Y(n_671) );
OR2x2_ASAP7_75t_L g647 ( .A(n_636), .B(n_648), .Y(n_647) );
OR2x2_ASAP7_75t_L g677 ( .A(n_636), .B(n_651), .Y(n_677) );
INVx2_ASAP7_75t_L g636 ( .A(n_637), .Y(n_636) );
AND2x2_ASAP7_75t_L g753 ( .A(n_637), .B(n_754), .Y(n_753) );
INVx1_ASAP7_75t_L g776 ( .A(n_638), .Y(n_776) );
NAND2xp5_ASAP7_75t_L g638 ( .A(n_639), .B(n_640), .Y(n_638) );
NAND2xp5_ASAP7_75t_L g688 ( .A(n_640), .B(n_689), .Y(n_688) );
NAND2xp5_ASAP7_75t_L g710 ( .A(n_640), .B(n_711), .Y(n_710) );
AND2x2_ASAP7_75t_L g788 ( .A(n_640), .B(n_664), .Y(n_788) );
NAND2xp5_ASAP7_75t_L g793 ( .A(n_640), .B(n_794), .Y(n_793) );
AND2x2_ASAP7_75t_L g731 ( .A(n_641), .B(n_713), .Y(n_731) );
INVx1_ASAP7_75t_SL g642 ( .A(n_643), .Y(n_642) );
AOI322xp5_ASAP7_75t_L g785 ( .A1(n_644), .A2(n_664), .A3(n_718), .B1(n_743), .B2(n_786), .C1(n_788), .C2(n_789), .Y(n_785) );
AOI211xp5_ASAP7_75t_SL g645 ( .A1(n_646), .A2(n_650), .B(n_652), .C(n_661), .Y(n_645) );
INVx1_ASAP7_75t_L g646 ( .A(n_647), .Y(n_646) );
NAND2xp5_ASAP7_75t_L g698 ( .A(n_648), .B(n_676), .Y(n_698) );
INVx1_ASAP7_75t_L g648 ( .A(n_649), .Y(n_648) );
AND2x2_ASAP7_75t_L g663 ( .A(n_649), .B(n_664), .Y(n_663) );
NOR2x1p5_ASAP7_75t_L g729 ( .A(n_649), .B(n_730), .Y(n_729) );
HB1xp67_ASAP7_75t_L g762 ( .A(n_649), .Y(n_762) );
O2A1O1Ixp33_ASAP7_75t_L g667 ( .A1(n_650), .A2(n_668), .B(n_671), .C(n_672), .Y(n_667) );
AND2x4_ASAP7_75t_L g686 ( .A(n_651), .B(n_670), .Y(n_686) );
INVx2_ASAP7_75t_L g696 ( .A(n_651), .Y(n_696) );
NAND2xp5_ASAP7_75t_SL g716 ( .A(n_651), .B(n_685), .Y(n_716) );
AND2x2_ASAP7_75t_L g758 ( .A(n_651), .B(n_759), .Y(n_758) );
NOR2xp33_ASAP7_75t_L g796 ( .A(n_651), .B(n_775), .Y(n_796) );
AND2x2_ASAP7_75t_L g797 ( .A(n_651), .B(n_679), .Y(n_797) );
AOI21xp33_ASAP7_75t_L g652 ( .A1(n_653), .A2(n_656), .B(n_658), .Y(n_652) );
AND2x2_ASAP7_75t_L g748 ( .A(n_654), .B(n_749), .Y(n_748) );
INVx1_ASAP7_75t_SL g654 ( .A(n_655), .Y(n_654) );
INVx1_ASAP7_75t_L g676 ( .A(n_657), .Y(n_676) );
INVx2_ASAP7_75t_L g658 ( .A(n_659), .Y(n_658) );
NOR2xp33_ASAP7_75t_L g661 ( .A(n_662), .B(n_666), .Y(n_661) );
INVx1_ASAP7_75t_L g662 ( .A(n_663), .Y(n_662) );
NAND2xp5_ASAP7_75t_L g724 ( .A(n_669), .B(n_725), .Y(n_724) );
INVx1_ASAP7_75t_L g763 ( .A(n_669), .Y(n_763) );
O2A1O1Ixp33_ASAP7_75t_SL g672 ( .A1(n_673), .A2(n_675), .B(n_677), .C(n_678), .Y(n_672) );
INVx1_ASAP7_75t_L g673 ( .A(n_674), .Y(n_673) );
INVx1_ASAP7_75t_L g675 ( .A(n_676), .Y(n_675) );
HB1xp67_ASAP7_75t_L g760 ( .A(n_676), .Y(n_760) );
INVx3_ASAP7_75t_SL g775 ( .A(n_679), .Y(n_775) );
NAND5xp2_ASAP7_75t_L g681 ( .A(n_682), .B(n_701), .C(n_708), .D(n_721), .E(n_732), .Y(n_681) );
AOI222xp33_ASAP7_75t_L g682 ( .A1(n_683), .A2(n_687), .B1(n_691), .B2(n_693), .C1(n_697), .C2(n_699), .Y(n_682) );
NOR2xp33_ASAP7_75t_L g683 ( .A(n_684), .B(n_686), .Y(n_683) );
AOI22xp5_ASAP7_75t_L g764 ( .A1(n_684), .A2(n_765), .B1(n_769), .B2(n_770), .Y(n_764) );
INVx2_ASAP7_75t_SL g684 ( .A(n_685), .Y(n_684) );
AND2x2_ASAP7_75t_L g714 ( .A(n_685), .B(n_686), .Y(n_714) );
INVx1_ASAP7_75t_L g687 ( .A(n_688), .Y(n_687) );
INVx1_ASAP7_75t_L g689 ( .A(n_690), .Y(n_689) );
INVx1_ASAP7_75t_SL g691 ( .A(n_692), .Y(n_691) );
NOR2xp33_ASAP7_75t_L g693 ( .A(n_694), .B(n_696), .Y(n_693) );
INVx1_ASAP7_75t_L g694 ( .A(n_695), .Y(n_694) );
NAND2xp5_ASAP7_75t_SL g781 ( .A(n_695), .B(n_782), .Y(n_781) );
NAND2xp5_ASAP7_75t_L g717 ( .A(n_696), .B(n_718), .Y(n_717) );
AND2x2_ASAP7_75t_L g733 ( .A(n_696), .B(n_734), .Y(n_733) );
OR2x2_ASAP7_75t_L g744 ( .A(n_696), .B(n_745), .Y(n_744) );
INVx1_ASAP7_75t_L g697 ( .A(n_698), .Y(n_697) );
INVx1_ASAP7_75t_SL g699 ( .A(n_700), .Y(n_699) );
OR2x2_ASAP7_75t_L g774 ( .A(n_700), .B(n_775), .Y(n_774) );
OR2x2_ASAP7_75t_L g705 ( .A(n_706), .B(n_707), .Y(n_705) );
INVx1_ASAP7_75t_L g722 ( .A(n_707), .Y(n_722) );
INVxp67_ASAP7_75t_L g709 ( .A(n_710), .Y(n_709) );
INVxp67_ASAP7_75t_L g711 ( .A(n_712), .Y(n_711) );
HB1xp67_ASAP7_75t_L g712 ( .A(n_713), .Y(n_712) );
AOI21xp33_ASAP7_75t_L g715 ( .A1(n_716), .A2(n_717), .B(n_719), .Y(n_715) );
AOI22xp33_ASAP7_75t_L g721 ( .A1(n_718), .A2(n_722), .B1(n_723), .B2(n_727), .Y(n_721) );
HB1xp67_ASAP7_75t_L g769 ( .A(n_718), .Y(n_769) );
INVx2_ASAP7_75t_SL g719 ( .A(n_720), .Y(n_719) );
AND2x2_ASAP7_75t_L g735 ( .A(n_720), .B(n_736), .Y(n_735) );
AND2x2_ASAP7_75t_L g740 ( .A(n_722), .B(n_741), .Y(n_740) );
INVx1_ASAP7_75t_L g723 ( .A(n_724), .Y(n_723) );
INVx1_ASAP7_75t_SL g725 ( .A(n_726), .Y(n_725) );
INVx1_ASAP7_75t_L g727 ( .A(n_728), .Y(n_727) );
NAND2xp5_ASAP7_75t_L g728 ( .A(n_729), .B(n_731), .Y(n_728) );
INVx1_ASAP7_75t_SL g768 ( .A(n_731), .Y(n_768) );
NAND2xp5_ASAP7_75t_L g732 ( .A(n_733), .B(n_735), .Y(n_732) );
NOR3xp33_ASAP7_75t_L g737 ( .A(n_738), .B(n_756), .C(n_779), .Y(n_737) );
NAND2xp5_ASAP7_75t_SL g738 ( .A(n_739), .B(n_755), .Y(n_738) );
AOI221xp5_ASAP7_75t_L g739 ( .A1(n_740), .A2(n_743), .B1(n_746), .B2(n_748), .C(n_751), .Y(n_739) );
INVx1_ASAP7_75t_SL g741 ( .A(n_742), .Y(n_741) );
OR2x2_ASAP7_75t_L g780 ( .A(n_742), .B(n_768), .Y(n_780) );
INVx1_ASAP7_75t_SL g743 ( .A(n_744), .Y(n_743) );
INVx1_ASAP7_75t_SL g746 ( .A(n_747), .Y(n_746) );
HB1xp67_ASAP7_75t_L g749 ( .A(n_750), .Y(n_749) );
INVx1_ASAP7_75t_SL g752 ( .A(n_753), .Y(n_752) );
OAI321xp33_ASAP7_75t_L g756 ( .A1(n_757), .A2(n_760), .A3(n_761), .B1(n_763), .B2(n_764), .C(n_772), .Y(n_756) );
INVx1_ASAP7_75t_SL g757 ( .A(n_758), .Y(n_757) );
INVx1_ASAP7_75t_L g761 ( .A(n_762), .Y(n_761) );
INVx1_ASAP7_75t_SL g765 ( .A(n_766), .Y(n_765) );
OR2x2_ASAP7_75t_L g766 ( .A(n_767), .B(n_768), .Y(n_766) );
AOI22xp33_ASAP7_75t_L g791 ( .A1(n_770), .A2(n_792), .B1(n_796), .B2(n_797), .Y(n_791) );
INVx1_ASAP7_75t_SL g770 ( .A(n_771), .Y(n_770) );
INVx1_ASAP7_75t_L g773 ( .A(n_774), .Y(n_773) );
INVx1_ASAP7_75t_L g777 ( .A(n_778), .Y(n_777) );
OAI211xp5_ASAP7_75t_SL g779 ( .A1(n_780), .A2(n_781), .B(n_785), .C(n_791), .Y(n_779) );
INVx1_ASAP7_75t_L g782 ( .A(n_783), .Y(n_782) );
INVx1_ASAP7_75t_L g786 ( .A(n_787), .Y(n_786) );
INVx1_ASAP7_75t_SL g789 ( .A(n_790), .Y(n_789) );
INVx1_ASAP7_75t_L g792 ( .A(n_793), .Y(n_792) );
INVxp67_ASAP7_75t_L g794 ( .A(n_795), .Y(n_794) );
NOR2x1_ASAP7_75t_L g798 ( .A(n_799), .B(n_803), .Y(n_798) );
NAND2xp5_ASAP7_75t_L g799 ( .A(n_800), .B(n_802), .Y(n_799) );
NOR2xp33_ASAP7_75t_L g808 ( .A(n_809), .B(n_810), .Y(n_808) );
BUFx2_ASAP7_75t_L g810 ( .A(n_811), .Y(n_810) );
CKINVDCx5p33_ASAP7_75t_R g812 ( .A(n_813), .Y(n_812) );
CKINVDCx20_ASAP7_75t_R g813 ( .A(n_814), .Y(n_813) );
INVx3_ASAP7_75t_SL g814 ( .A(n_815), .Y(n_814) );
NAND2xp5_ASAP7_75t_SL g815 ( .A(n_816), .B(n_820), .Y(n_815) );
endmodule