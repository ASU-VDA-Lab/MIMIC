module fake_jpeg_14897_n_361 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_361);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_361;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx6_ASAP7_75t_L g14 ( 
.A(n_9),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_0),
.Y(n_15)
);

INVx4_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

INVx5_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_12),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_11),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_13),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_5),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_3),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_5),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

BUFx10_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_12),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_1),
.Y(n_35)
);

INVx11_ASAP7_75t_SL g36 ( 
.A(n_4),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_12),
.Y(n_37)
);

INVx11_ASAP7_75t_L g38 ( 
.A(n_36),
.Y(n_38)
);

INVx8_ASAP7_75t_L g77 ( 
.A(n_38),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_15),
.B(n_0),
.Y(n_39)
);

AND2x2_ASAP7_75t_L g88 ( 
.A(n_39),
.B(n_42),
.Y(n_88)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_16),
.Y(n_40)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_40),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_34),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_41),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_15),
.B(n_1),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_16),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_43),
.B(n_51),
.Y(n_79)
);

OR2x2_ASAP7_75t_L g44 ( 
.A(n_19),
.B(n_1),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_SL g91 ( 
.A(n_44),
.B(n_48),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_34),
.Y(n_45)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_45),
.Y(n_70)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_18),
.Y(n_46)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_46),
.Y(n_84)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_18),
.Y(n_47)
);

INVx8_ASAP7_75t_L g109 ( 
.A(n_47),
.Y(n_109)
);

OR2x2_ASAP7_75t_L g48 ( 
.A(n_19),
.B(n_1),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_17),
.Y(n_49)
);

AND2x2_ASAP7_75t_L g102 ( 
.A(n_49),
.B(n_55),
.Y(n_102)
);

INVx11_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

INVx8_ASAP7_75t_L g113 ( 
.A(n_50),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_17),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g52 ( 
.A1(n_14),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_52),
.A2(n_4),
.B1(n_6),
.B2(n_7),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_20),
.B(n_2),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_53),
.B(n_59),
.Y(n_83)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_14),
.Y(n_54)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_54),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_26),
.B(n_2),
.Y(n_55)
);

INVx2_ASAP7_75t_SL g56 ( 
.A(n_33),
.Y(n_56)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_56),
.Y(n_89)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_14),
.Y(n_57)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_57),
.Y(n_100)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_26),
.Y(n_58)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_58),
.Y(n_101)
);

HB1xp67_ASAP7_75t_L g59 ( 
.A(n_33),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_34),
.Y(n_60)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_60),
.Y(n_92)
);

AND2x2_ASAP7_75t_L g61 ( 
.A(n_29),
.B(n_2),
.Y(n_61)
);

OR2x2_ASAP7_75t_L g106 ( 
.A(n_61),
.B(n_21),
.Y(n_106)
);

INVx5_ASAP7_75t_L g62 ( 
.A(n_18),
.Y(n_62)
);

INVx5_ASAP7_75t_L g95 ( 
.A(n_62),
.Y(n_95)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_34),
.Y(n_63)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_63),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_35),
.Y(n_64)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_64),
.Y(n_108)
);

INVx8_ASAP7_75t_L g65 ( 
.A(n_22),
.Y(n_65)
);

INVx8_ASAP7_75t_L g117 ( 
.A(n_65),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_35),
.Y(n_66)
);

INVx4_ASAP7_75t_L g111 ( 
.A(n_66),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_20),
.B(n_3),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_67),
.B(n_28),
.Y(n_85)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_33),
.Y(n_68)
);

INVx8_ASAP7_75t_L g118 ( 
.A(n_68),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_35),
.Y(n_69)
);

INVx4_ASAP7_75t_L g115 ( 
.A(n_69),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_62),
.A2(n_16),
.B1(n_29),
.B2(n_31),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_71),
.A2(n_74),
.B1(n_87),
.B2(n_96),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_54),
.A2(n_31),
.B1(n_35),
.B2(n_27),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_72),
.A2(n_78),
.B1(n_80),
.B2(n_99),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_39),
.B(n_42),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_73),
.B(n_103),
.Y(n_154)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_46),
.A2(n_25),
.B1(n_23),
.B2(n_28),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_75),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_125)
);

INVx4_ASAP7_75t_SL g76 ( 
.A(n_38),
.Y(n_76)
);

INVx13_ASAP7_75t_L g139 ( 
.A(n_76),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_52),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_57),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_44),
.B(n_23),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_82),
.B(n_86),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_85),
.B(n_93),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_48),
.B(n_25),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_47),
.A2(n_24),
.B1(n_27),
.B2(n_30),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_63),
.A2(n_24),
.B1(n_27),
.B2(n_37),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_90),
.A2(n_66),
.B1(n_64),
.B2(n_60),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_51),
.B(n_37),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_55),
.B(n_37),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_94),
.B(n_110),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_50),
.A2(n_30),
.B1(n_21),
.B2(n_9),
.Y(n_96)
);

INVx6_ASAP7_75t_L g97 ( 
.A(n_41),
.Y(n_97)
);

INVx8_ASAP7_75t_L g159 ( 
.A(n_97),
.Y(n_159)
);

BUFx3_ASAP7_75t_L g98 ( 
.A(n_41),
.Y(n_98)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_98),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_L g99 ( 
.A1(n_68),
.A2(n_33),
.B1(n_30),
.B2(n_21),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_61),
.B(n_32),
.Y(n_103)
);

INVx5_ASAP7_75t_L g105 ( 
.A(n_65),
.Y(n_105)
);

INVx5_ASAP7_75t_L g138 ( 
.A(n_105),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_L g165 ( 
.A1(n_106),
.A2(n_76),
.B(n_116),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_49),
.B(n_33),
.Y(n_110)
);

BUFx3_ASAP7_75t_L g112 ( 
.A(n_69),
.Y(n_112)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_112),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_56),
.A2(n_6),
.B1(n_8),
.B2(n_9),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g136 ( 
.A1(n_114),
.A2(n_10),
.B1(n_11),
.B2(n_13),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_102),
.A2(n_61),
.B1(n_58),
.B2(n_56),
.Y(n_122)
);

OR2x2_ASAP7_75t_L g188 ( 
.A(n_122),
.B(n_140),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_73),
.B(n_40),
.C(n_43),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_124),
.B(n_141),
.C(n_113),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_125),
.A2(n_149),
.B1(n_151),
.B2(n_158),
.Y(n_186)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_89),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_126),
.B(n_130),
.Y(n_177)
);

INVx4_ASAP7_75t_L g128 ( 
.A(n_77),
.Y(n_128)
);

BUFx3_ASAP7_75t_L g202 ( 
.A(n_128),
.Y(n_202)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_89),
.Y(n_129)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_129),
.Y(n_169)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_101),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_131),
.A2(n_132),
.B1(n_136),
.B2(n_142),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_88),
.A2(n_102),
.B1(n_90),
.B2(n_103),
.Y(n_132)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_101),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_134),
.B(n_150),
.Y(n_203)
);

OR2x2_ASAP7_75t_L g135 ( 
.A(n_91),
.B(n_33),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_135),
.B(n_156),
.Y(n_170)
);

INVx3_ASAP7_75t_L g137 ( 
.A(n_84),
.Y(n_137)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_137),
.Y(n_172)
);

CKINVDCx16_ASAP7_75t_R g140 ( 
.A(n_104),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_L g141 ( 
.A(n_88),
.B(n_22),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_88),
.A2(n_69),
.B1(n_45),
.B2(n_13),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_102),
.A2(n_32),
.B1(n_22),
.B2(n_10),
.Y(n_144)
);

INVxp67_ASAP7_75t_L g167 ( 
.A(n_144),
.Y(n_167)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_81),
.Y(n_145)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_145),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_79),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_146),
.B(n_152),
.Y(n_206)
);

AOI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_95),
.A2(n_22),
.B1(n_32),
.B2(n_109),
.Y(n_147)
);

INVxp67_ASAP7_75t_L g168 ( 
.A(n_147),
.Y(n_168)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_81),
.Y(n_148)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_148),
.Y(n_178)
);

O2A1O1Ixp33_ASAP7_75t_SL g149 ( 
.A1(n_91),
.A2(n_22),
.B(n_32),
.C(n_78),
.Y(n_149)
);

INVxp67_ASAP7_75t_L g150 ( 
.A(n_100),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_75),
.A2(n_32),
.B1(n_80),
.B2(n_97),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_104),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_83),
.B(n_106),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_SL g184 ( 
.A(n_153),
.B(n_155),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_84),
.B(n_109),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_100),
.B(n_107),
.Y(n_156)
);

AOI21xp5_ASAP7_75t_L g157 ( 
.A1(n_95),
.A2(n_105),
.B(n_70),
.Y(n_157)
);

NOR3xp33_ASAP7_75t_L g171 ( 
.A(n_157),
.B(n_163),
.C(n_113),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_L g158 ( 
.A1(n_70),
.A2(n_111),
.B1(n_108),
.B2(n_92),
.Y(n_158)
);

AOI22xp33_ASAP7_75t_SL g160 ( 
.A1(n_92),
.A2(n_111),
.B1(n_108),
.B2(n_115),
.Y(n_160)
);

INVxp67_ASAP7_75t_L g197 ( 
.A(n_160),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_72),
.B(n_117),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_SL g194 ( 
.A(n_161),
.B(n_142),
.Y(n_194)
);

INVxp67_ASAP7_75t_L g162 ( 
.A(n_107),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_162),
.B(n_164),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_115),
.A2(n_118),
.B1(n_117),
.B2(n_116),
.Y(n_163)
);

INVx4_ASAP7_75t_L g164 ( 
.A(n_77),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_L g209 ( 
.A(n_165),
.B(n_149),
.Y(n_209)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_98),
.Y(n_166)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_166),
.Y(n_183)
);

AOI22xp33_ASAP7_75t_L g246 ( 
.A1(n_171),
.A2(n_208),
.B1(n_186),
.B2(n_203),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_154),
.B(n_118),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_SL g222 ( 
.A(n_173),
.B(n_179),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_156),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_174),
.B(n_175),
.Y(n_214)
);

CKINVDCx16_ASAP7_75t_R g175 ( 
.A(n_119),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_154),
.B(n_112),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g235 ( 
.A(n_180),
.B(n_209),
.Y(n_235)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_129),
.Y(n_181)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_181),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_141),
.B(n_124),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_SL g236 ( 
.A(n_182),
.B(n_194),
.Y(n_236)
);

NAND2x1_ASAP7_75t_L g185 ( 
.A(n_165),
.B(n_144),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_SL g218 ( 
.A1(n_185),
.A2(n_135),
.B(n_130),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_132),
.B(n_122),
.C(n_143),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_189),
.B(n_123),
.C(n_157),
.Y(n_212)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_145),
.Y(n_190)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_190),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_148),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_191),
.B(n_192),
.Y(n_215)
);

CKINVDCx16_ASAP7_75t_R g192 ( 
.A(n_119),
.Y(n_192)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_133),
.Y(n_193)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_193),
.Y(n_223)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_133),
.Y(n_195)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_195),
.Y(n_224)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_137),
.Y(n_196)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_196),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_SL g198 ( 
.A(n_127),
.B(n_146),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_SL g241 ( 
.A(n_198),
.B(n_204),
.Y(n_241)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_158),
.Y(n_199)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_199),
.Y(n_231)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_163),
.Y(n_200)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_200),
.Y(n_232)
);

BUFx6f_ASAP7_75t_L g201 ( 
.A(n_159),
.Y(n_201)
);

INVx4_ASAP7_75t_L g211 ( 
.A(n_201),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_135),
.B(n_152),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_166),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_207),
.B(n_208),
.Y(n_219)
);

INVx3_ASAP7_75t_L g208 ( 
.A(n_138),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_187),
.A2(n_151),
.B1(n_123),
.B2(n_125),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_210),
.A2(n_216),
.B1(n_225),
.B2(n_231),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_212),
.B(n_213),
.C(n_238),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_182),
.B(n_140),
.C(n_121),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_200),
.A2(n_149),
.B1(n_120),
.B2(n_131),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_SL g254 ( 
.A1(n_218),
.A2(n_229),
.B(n_244),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_206),
.B(n_134),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_SL g260 ( 
.A(n_221),
.B(n_227),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_186),
.A2(n_159),
.B1(n_138),
.B2(n_150),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_184),
.B(n_126),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_174),
.B(n_139),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_228),
.B(n_245),
.Y(n_248)
);

AOI21xp5_ASAP7_75t_L g229 ( 
.A1(n_168),
.A2(n_162),
.B(n_128),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_169),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_SL g269 ( 
.A(n_230),
.B(n_233),
.Y(n_269)
);

INVxp67_ASAP7_75t_L g233 ( 
.A(n_205),
.Y(n_233)
);

INVx2_ASAP7_75t_SL g234 ( 
.A(n_181),
.Y(n_234)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_234),
.Y(n_255)
);

INVx4_ASAP7_75t_L g237 ( 
.A(n_172),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_237),
.B(n_240),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_180),
.B(n_164),
.C(n_139),
.Y(n_238)
);

NOR2x1_ASAP7_75t_L g239 ( 
.A(n_185),
.B(n_139),
.Y(n_239)
);

OAI21xp5_ASAP7_75t_L g256 ( 
.A1(n_239),
.A2(n_191),
.B(n_207),
.Y(n_256)
);

NOR3xp33_ASAP7_75t_SL g240 ( 
.A(n_185),
.B(n_167),
.C(n_188),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_167),
.A2(n_168),
.B1(n_197),
.B2(n_199),
.Y(n_242)
);

INVxp67_ASAP7_75t_L g267 ( 
.A(n_242),
.Y(n_267)
);

NOR3xp33_ASAP7_75t_L g243 ( 
.A(n_189),
.B(n_204),
.C(n_188),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_243),
.B(n_246),
.Y(n_249)
);

AOI21xp5_ASAP7_75t_L g244 ( 
.A1(n_209),
.A2(n_197),
.B(n_170),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_179),
.B(n_170),
.Y(n_245)
);

AND2x2_ASAP7_75t_L g250 ( 
.A(n_239),
.B(n_242),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_250),
.A2(n_266),
.B1(n_271),
.B2(n_232),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_222),
.B(n_173),
.Y(n_251)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_251),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_221),
.B(n_202),
.Y(n_252)
);

CKINVDCx14_ASAP7_75t_R g286 ( 
.A(n_252),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_235),
.B(n_177),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_253),
.B(n_261),
.C(n_264),
.Y(n_283)
);

AOI22xp33_ASAP7_75t_L g282 ( 
.A1(n_256),
.A2(n_265),
.B1(n_229),
.B2(n_232),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_237),
.B(n_202),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_SL g292 ( 
.A(n_258),
.B(n_262),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_231),
.A2(n_183),
.B1(n_176),
.B2(n_178),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_SL g299 ( 
.A1(n_259),
.A2(n_220),
.B1(n_230),
.B2(n_224),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_235),
.B(n_183),
.C(n_176),
.Y(n_261)
);

CKINVDCx16_ASAP7_75t_R g262 ( 
.A(n_215),
.Y(n_262)
);

OAI21xp5_ASAP7_75t_SL g263 ( 
.A1(n_244),
.A2(n_172),
.B(n_196),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_263),
.B(n_268),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g264 ( 
.A(n_238),
.B(n_178),
.Y(n_264)
);

OAI21xp5_ASAP7_75t_L g265 ( 
.A1(n_239),
.A2(n_190),
.B(n_169),
.Y(n_265)
);

AND2x2_ASAP7_75t_L g266 ( 
.A(n_212),
.B(n_193),
.Y(n_266)
);

OAI21xp5_ASAP7_75t_SL g268 ( 
.A1(n_218),
.A2(n_195),
.B(n_201),
.Y(n_268)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_220),
.Y(n_270)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_270),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_213),
.B(n_245),
.C(n_236),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_272),
.B(n_275),
.C(n_276),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_215),
.B(n_227),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_273),
.B(n_219),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_222),
.B(n_241),
.Y(n_274)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_274),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_236),
.B(n_214),
.C(n_210),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_240),
.B(n_214),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_241),
.B(n_228),
.Y(n_277)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_277),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_255),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_278),
.B(n_289),
.Y(n_303)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_280),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_282),
.B(n_293),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_260),
.B(n_219),
.Y(n_285)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_285),
.Y(n_316)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_270),
.Y(n_289)
);

INVx1_ASAP7_75t_SL g290 ( 
.A(n_250),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_290),
.B(n_291),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_260),
.B(n_226),
.Y(n_291)
);

BUFx24_ASAP7_75t_SL g293 ( 
.A(n_274),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_262),
.B(n_226),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_SL g320 ( 
.A(n_294),
.B(n_298),
.Y(n_320)
);

AND2x2_ASAP7_75t_L g318 ( 
.A(n_295),
.B(n_300),
.Y(n_318)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_264),
.B(n_216),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_297),
.B(n_257),
.C(n_261),
.Y(n_309)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_255),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_L g313 ( 
.A1(n_299),
.A2(n_301),
.B1(n_302),
.B2(n_248),
.Y(n_313)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_259),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_269),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_248),
.B(n_223),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_SL g304 ( 
.A1(n_290),
.A2(n_267),
.B1(n_250),
.B2(n_266),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_SL g328 ( 
.A1(n_304),
.A2(n_306),
.B1(n_310),
.B2(n_292),
.Y(n_328)
);

XNOR2xp5_ASAP7_75t_L g305 ( 
.A(n_297),
.B(n_257),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_305),
.B(n_311),
.C(n_317),
.Y(n_322)
);

AOI22xp5_ASAP7_75t_SL g306 ( 
.A1(n_300),
.A2(n_267),
.B1(n_266),
.B2(n_254),
.Y(n_306)
);

OR2x2_ASAP7_75t_L g308 ( 
.A(n_288),
.B(n_277),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_308),
.B(n_284),
.Y(n_333)
);

XOR2xp5_ASAP7_75t_L g327 ( 
.A(n_309),
.B(n_319),
.Y(n_327)
);

AOI22xp5_ASAP7_75t_L g310 ( 
.A1(n_287),
.A2(n_271),
.B1(n_275),
.B2(n_249),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_283),
.B(n_253),
.C(n_272),
.Y(n_311)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_313),
.Y(n_329)
);

AOI321xp33_ASAP7_75t_L g315 ( 
.A1(n_287),
.A2(n_276),
.A3(n_265),
.B1(n_256),
.B2(n_247),
.C(n_254),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_L g332 ( 
.A1(n_315),
.A2(n_284),
.B1(n_225),
.B2(n_223),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_283),
.B(n_263),
.C(n_251),
.Y(n_317)
);

XOR2xp5_ASAP7_75t_L g319 ( 
.A(n_296),
.B(n_268),
.Y(n_319)
);

AOI21xp5_ASAP7_75t_L g321 ( 
.A1(n_318),
.A2(n_279),
.B(n_295),
.Y(n_321)
);

XNOR2xp5_ASAP7_75t_L g344 ( 
.A(n_321),
.B(n_326),
.Y(n_344)
);

XNOR2xp5_ASAP7_75t_SL g323 ( 
.A(n_305),
.B(n_279),
.Y(n_323)
);

XOR2xp5_ASAP7_75t_L g339 ( 
.A(n_323),
.B(n_328),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_309),
.B(n_296),
.C(n_288),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_324),
.B(n_330),
.Y(n_336)
);

AOI22xp5_ASAP7_75t_L g325 ( 
.A1(n_318),
.A2(n_281),
.B1(n_278),
.B2(n_286),
.Y(n_325)
);

AOI22xp5_ASAP7_75t_L g335 ( 
.A1(n_325),
.A2(n_314),
.B1(n_316),
.B2(n_306),
.Y(n_335)
);

AOI21xp5_ASAP7_75t_L g326 ( 
.A1(n_303),
.A2(n_281),
.B(n_298),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_319),
.B(n_301),
.C(n_289),
.Y(n_330)
);

XNOR2xp5_ASAP7_75t_L g331 ( 
.A(n_317),
.B(n_299),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_331),
.B(n_333),
.Y(n_337)
);

AOI321xp33_ASAP7_75t_L g343 ( 
.A1(n_332),
.A2(n_304),
.A3(n_311),
.B1(n_217),
.B2(n_234),
.C(n_211),
.Y(n_343)
);

OAI22xp5_ASAP7_75t_L g334 ( 
.A1(n_310),
.A2(n_211),
.B1(n_224),
.B2(n_234),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_SL g340 ( 
.A(n_334),
.B(n_312),
.Y(n_340)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_335),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_333),
.B(n_320),
.Y(n_338)
);

HB1xp67_ASAP7_75t_L g349 ( 
.A(n_338),
.Y(n_349)
);

AOI22xp5_ASAP7_75t_L g348 ( 
.A1(n_340),
.A2(n_343),
.B1(n_330),
.B2(n_325),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_326),
.B(n_308),
.Y(n_341)
);

AOI31xp67_ASAP7_75t_SL g350 ( 
.A1(n_341),
.A2(n_342),
.A3(n_335),
.B(n_344),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_SL g342 ( 
.A(n_329),
.B(n_307),
.Y(n_342)
);

AOI21x1_ASAP7_75t_L g345 ( 
.A1(n_344),
.A2(n_321),
.B(n_328),
.Y(n_345)
);

AOI22xp5_ASAP7_75t_SL g351 ( 
.A1(n_345),
.A2(n_339),
.B1(n_331),
.B2(n_323),
.Y(n_351)
);

AOI21xp5_ASAP7_75t_SL g346 ( 
.A1(n_337),
.A2(n_336),
.B(n_343),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_346),
.B(n_339),
.Y(n_352)
);

MAJIxp5_ASAP7_75t_L g353 ( 
.A(n_348),
.B(n_324),
.C(n_322),
.Y(n_353)
);

OR2x2_ASAP7_75t_L g354 ( 
.A(n_350),
.B(n_322),
.Y(n_354)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_351),
.Y(n_356)
);

MAJIxp5_ASAP7_75t_L g355 ( 
.A(n_352),
.B(n_353),
.C(n_354),
.Y(n_355)
);

MAJIxp5_ASAP7_75t_L g357 ( 
.A(n_355),
.B(n_356),
.C(n_327),
.Y(n_357)
);

AOI21xp5_ASAP7_75t_L g359 ( 
.A1(n_357),
.A2(n_358),
.B(n_327),
.Y(n_359)
);

OR2x2_ASAP7_75t_L g358 ( 
.A(n_355),
.B(n_349),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_359),
.B(n_354),
.Y(n_360)
);

XOR2xp5_ASAP7_75t_L g361 ( 
.A(n_360),
.B(n_347),
.Y(n_361)
);


endmodule