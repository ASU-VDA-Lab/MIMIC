module fake_netlist_6_1057_n_1902 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_161, n_68, n_166, n_28, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_178, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_180, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_181, n_76, n_36, n_182, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_175, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_104, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_173, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_171, n_31, n_57, n_169, n_53, n_51, n_44, n_56, n_1902);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_161;
input n_68;
input n_166;
input n_28;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_178;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_175;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_104;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_173;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_171;
input n_31;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1902;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_1853;
wire n_783;
wire n_1738;
wire n_798;
wire n_188;
wire n_1575;
wire n_1854;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1688;
wire n_1691;
wire n_1009;
wire n_1743;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_1844;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_1786;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_200;
wire n_447;
wire n_1803;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1867;
wire n_1704;
wire n_1078;
wire n_250;
wire n_544;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_658;
wire n_616;
wire n_1874;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1842;
wire n_1620;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1798;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_1820;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_1894;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_1815;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1644;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_577;
wire n_1843;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1762;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1876;
wire n_1895;
wire n_1697;
wire n_243;
wire n_979;
wire n_1873;
wire n_905;
wire n_1866;
wire n_1680;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1865;
wire n_1875;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_530;
wire n_1563;
wire n_277;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_1760;
wire n_210;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_1896;
wire n_429;
wire n_1747;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1802;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_835;
wire n_1214;
wire n_928;
wire n_690;
wire n_850;
wire n_1801;
wire n_1886;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_1813;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_1709;
wire n_1825;
wire n_1757;
wire n_1796;
wire n_1792;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_462;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_297;
wire n_595;
wire n_627;
wire n_1767;
wire n_1779;
wire n_524;
wire n_1465;
wire n_342;
wire n_1858;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_1880;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_1839;
wire n_685;
wire n_1765;
wire n_353;
wire n_605;
wire n_1514;
wire n_1863;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_1808;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_1788;
wire n_622;
wire n_1469;
wire n_1838;
wire n_1835;
wire n_1766;
wire n_1776;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_1771;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_1878;
wire n_899;
wire n_189;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_1577;
wire n_1181;
wire n_1822;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_1817;
wire n_927;
wire n_1849;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_184;
wire n_552;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_216;
wire n_912;
wire n_1857;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_755;
wire n_931;
wire n_1021;
wire n_527;
wire n_474;
wire n_811;
wire n_683;
wire n_1207;
wire n_312;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_1897;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_1837;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1736;
wire n_1564;
wire n_211;
wire n_1483;
wire n_1834;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_1787;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_1877;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1769;
wire n_1220;
wire n_1893;
wire n_556;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1775;
wire n_1773;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_1745;
wire n_914;
wire n_759;
wire n_1831;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_1901;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1892;
wire n_1135;
wire n_1179;
wire n_1169;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1580;
wire n_1425;
wire n_1881;
wire n_1267;
wire n_1281;
wire n_1806;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_1855;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_1832;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1594;
wire n_664;
wire n_1869;
wire n_1764;
wire n_1429;
wire n_1610;
wire n_1889;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_186;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_1871;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_1859;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1852;
wire n_1024;
wire n_1768;
wire n_198;
wire n_1847;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1841;
wire n_1639;
wire n_1623;
wire n_183;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1818;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1686;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1262;
wire n_218;
wire n_1891;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_1870;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1827;
wire n_1361;
wire n_1864;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_370;
wire n_1695;
wire n_1828;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1883;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_1823;
wire n_227;
wire n_1720;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_1795;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1845;
wire n_1489;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_1846;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_1782;
wire n_282;
wire n_1676;
wire n_833;
wire n_1830;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_1900;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_1086;
wire n_1066;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_1758;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1794;
wire n_1236;
wire n_1559;
wire n_1725;
wire n_1872;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1746;
wire n_1325;
wire n_1002;
wire n_1741;
wire n_545;
wire n_489;
wire n_1804;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1860;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_187;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1800;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_1826;
wire n_566;
wire n_1023;
wire n_1882;
wire n_1118;
wire n_1076;
wire n_194;
wire n_1007;
wire n_1807;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1814;
wire n_1631;
wire n_591;
wire n_1377;
wire n_1879;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1824;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_1810;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_1729;
wire n_669;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1848;
wire n_763;
wire n_1147;
wire n_1785;
wire n_360;
wire n_1754;
wire n_1506;
wire n_1652;
wire n_1812;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_1173;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1821;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_185;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1525;
wire n_455;
wire n_1585;
wire n_1851;
wire n_363;
wire n_1799;
wire n_1090;
wire n_592;
wire n_1816;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_1829;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_1789;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_404;
wire n_271;
wire n_1884;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1819;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_1861;
wire n_373;
wire n_1632;
wire n_1890;
wire n_1805;
wire n_257;
wire n_1557;
wire n_1888;
wire n_1833;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_1850;
wire n_1898;
wire n_1868;
wire n_207;
wire n_1089;
wire n_1887;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_1836;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1899;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_1856;
wire n_1862;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1885;
wire n_1013;
wire n_1259;
wire n_192;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

INVx1_ASAP7_75t_L g183 ( 
.A(n_93),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_170),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_34),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_21),
.Y(n_186)
);

INVx2_ASAP7_75t_SL g187 ( 
.A(n_172),
.Y(n_187)
);

INVx1_ASAP7_75t_SL g188 ( 
.A(n_140),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_124),
.Y(n_189)
);

BUFx3_ASAP7_75t_L g190 ( 
.A(n_148),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_65),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_54),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_111),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_63),
.Y(n_194)
);

INVx2_ASAP7_75t_SL g195 ( 
.A(n_29),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_138),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_29),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_4),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_110),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_35),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_127),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_94),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_149),
.Y(n_203)
);

INVx1_ASAP7_75t_SL g204 ( 
.A(n_5),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_117),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_160),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_126),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_116),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_120),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_112),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_28),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_146),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_168),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_113),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_121),
.Y(n_215)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_68),
.Y(n_216)
);

BUFx2_ASAP7_75t_L g217 ( 
.A(n_132),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_67),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_100),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_34),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_91),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_163),
.Y(n_222)
);

BUFx6f_ASAP7_75t_L g223 ( 
.A(n_159),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_44),
.Y(n_224)
);

INVx1_ASAP7_75t_SL g225 ( 
.A(n_47),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_167),
.Y(n_226)
);

BUFx3_ASAP7_75t_L g227 ( 
.A(n_102),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_83),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_105),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_144),
.Y(n_230)
);

HB1xp67_ASAP7_75t_L g231 ( 
.A(n_125),
.Y(n_231)
);

BUFx3_ASAP7_75t_L g232 ( 
.A(n_176),
.Y(n_232)
);

BUFx6f_ASAP7_75t_L g233 ( 
.A(n_1),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_58),
.Y(n_234)
);

INVx1_ASAP7_75t_SL g235 ( 
.A(n_7),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_25),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_182),
.Y(n_237)
);

CKINVDCx14_ASAP7_75t_R g238 ( 
.A(n_7),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_48),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_51),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_118),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_40),
.Y(n_242)
);

HB1xp67_ASAP7_75t_L g243 ( 
.A(n_12),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_47),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_139),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_71),
.Y(n_246)
);

BUFx3_ASAP7_75t_L g247 ( 
.A(n_56),
.Y(n_247)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_31),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_55),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_6),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_39),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_74),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_54),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_95),
.Y(n_254)
);

INVxp67_ASAP7_75t_L g255 ( 
.A(n_52),
.Y(n_255)
);

BUFx3_ASAP7_75t_L g256 ( 
.A(n_75),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_64),
.Y(n_257)
);

BUFx10_ASAP7_75t_L g258 ( 
.A(n_19),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_130),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_98),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_4),
.Y(n_261)
);

BUFx6f_ASAP7_75t_L g262 ( 
.A(n_92),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_90),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_96),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_28),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_64),
.Y(n_266)
);

INVx1_ASAP7_75t_SL g267 ( 
.A(n_51),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_178),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_151),
.Y(n_269)
);

BUFx3_ASAP7_75t_L g270 ( 
.A(n_114),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_158),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_123),
.Y(n_272)
);

INVx2_ASAP7_75t_SL g273 ( 
.A(n_11),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_42),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_38),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_21),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_77),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_57),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_142),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_10),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_104),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_122),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_80),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_103),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_41),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_169),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_152),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_37),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_12),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_107),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_46),
.Y(n_291)
);

BUFx3_ASAP7_75t_L g292 ( 
.A(n_155),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_44),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_137),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_48),
.Y(n_295)
);

BUFx3_ASAP7_75t_L g296 ( 
.A(n_22),
.Y(n_296)
);

INVx2_ASAP7_75t_L g297 ( 
.A(n_97),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_0),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g299 ( 
.A(n_65),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g300 ( 
.A(n_57),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_38),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_10),
.Y(n_302)
);

BUFx8_ASAP7_75t_SL g303 ( 
.A(n_175),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_115),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_41),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_82),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_87),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_128),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_157),
.Y(n_309)
);

BUFx3_ASAP7_75t_L g310 ( 
.A(n_89),
.Y(n_310)
);

INVx2_ASAP7_75t_L g311 ( 
.A(n_17),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_43),
.Y(n_312)
);

BUFx6f_ASAP7_75t_L g313 ( 
.A(n_141),
.Y(n_313)
);

BUFx10_ASAP7_75t_L g314 ( 
.A(n_43),
.Y(n_314)
);

BUFx6f_ASAP7_75t_L g315 ( 
.A(n_108),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_66),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_32),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_153),
.Y(n_318)
);

INVx1_ASAP7_75t_SL g319 ( 
.A(n_2),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_25),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_99),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_119),
.Y(n_322)
);

INVx2_ASAP7_75t_L g323 ( 
.A(n_166),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_150),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_69),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_164),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_156),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_15),
.Y(n_328)
);

BUFx6f_ASAP7_75t_L g329 ( 
.A(n_79),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_81),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_2),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_45),
.Y(n_332)
);

BUFx6f_ASAP7_75t_L g333 ( 
.A(n_165),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_58),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_59),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_32),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_52),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_173),
.Y(n_338)
);

CKINVDCx20_ASAP7_75t_R g339 ( 
.A(n_179),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_70),
.Y(n_340)
);

INVx2_ASAP7_75t_L g341 ( 
.A(n_106),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_9),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_62),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_9),
.Y(n_344)
);

INVxp67_ASAP7_75t_L g345 ( 
.A(n_45),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_60),
.Y(n_346)
);

BUFx10_ASAP7_75t_L g347 ( 
.A(n_86),
.Y(n_347)
);

INVx1_ASAP7_75t_SL g348 ( 
.A(n_180),
.Y(n_348)
);

CKINVDCx20_ASAP7_75t_R g349 ( 
.A(n_174),
.Y(n_349)
);

INVx1_ASAP7_75t_SL g350 ( 
.A(n_14),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_72),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_177),
.Y(n_352)
);

BUFx10_ASAP7_75t_L g353 ( 
.A(n_134),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_30),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_101),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_73),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_37),
.Y(n_357)
);

INVx2_ASAP7_75t_SL g358 ( 
.A(n_84),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_23),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_136),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_50),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_36),
.Y(n_362)
);

CKINVDCx20_ASAP7_75t_R g363 ( 
.A(n_50),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_162),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_135),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_53),
.Y(n_366)
);

BUFx6f_ASAP7_75t_L g367 ( 
.A(n_223),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_247),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_238),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_236),
.Y(n_370)
);

CKINVDCx20_ASAP7_75t_R g371 ( 
.A(n_207),
.Y(n_371)
);

CKINVDCx20_ASAP7_75t_R g372 ( 
.A(n_208),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_247),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_296),
.Y(n_374)
);

NOR2xp67_ASAP7_75t_L g375 ( 
.A(n_255),
.B(n_0),
.Y(n_375)
);

BUFx2_ASAP7_75t_L g376 ( 
.A(n_296),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_233),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_233),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_233),
.Y(n_379)
);

NOR2xp33_ASAP7_75t_L g380 ( 
.A(n_217),
.B(n_1),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_239),
.Y(n_381)
);

NOR2xp33_ASAP7_75t_L g382 ( 
.A(n_231),
.B(n_3),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_240),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_233),
.Y(n_384)
);

NOR2xp33_ASAP7_75t_L g385 ( 
.A(n_187),
.B(n_358),
.Y(n_385)
);

INVxp67_ASAP7_75t_L g386 ( 
.A(n_243),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_233),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_185),
.Y(n_388)
);

HB1xp67_ASAP7_75t_L g389 ( 
.A(n_194),
.Y(n_389)
);

CKINVDCx20_ASAP7_75t_R g390 ( 
.A(n_212),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_242),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_244),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_248),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_248),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_311),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_249),
.Y(n_396)
);

BUFx6f_ASAP7_75t_SL g397 ( 
.A(n_347),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_191),
.Y(n_398)
);

XOR2xp5_ASAP7_75t_L g399 ( 
.A(n_186),
.B(n_3),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_192),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_234),
.Y(n_401)
);

OR2x2_ASAP7_75t_L g402 ( 
.A(n_250),
.B(n_5),
.Y(n_402)
);

INVxp67_ASAP7_75t_L g403 ( 
.A(n_258),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_276),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_280),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_251),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_257),
.Y(n_407)
);

CKINVDCx16_ASAP7_75t_R g408 ( 
.A(n_258),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_261),
.Y(n_409)
);

INVxp67_ASAP7_75t_SL g410 ( 
.A(n_190),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_291),
.Y(n_411)
);

CKINVDCx20_ASAP7_75t_R g412 ( 
.A(n_264),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_311),
.Y(n_413)
);

INVxp67_ASAP7_75t_SL g414 ( 
.A(n_190),
.Y(n_414)
);

NOR2xp67_ASAP7_75t_L g415 ( 
.A(n_345),
.B(n_6),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_265),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_293),
.Y(n_417)
);

NOR2xp67_ASAP7_75t_L g418 ( 
.A(n_195),
.B(n_8),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_266),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_274),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_278),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_301),
.Y(n_422)
);

INVx3_ASAP7_75t_L g423 ( 
.A(n_227),
.Y(n_423)
);

CKINVDCx20_ASAP7_75t_R g424 ( 
.A(n_279),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_317),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_328),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_285),
.Y(n_427)
);

NOR2xp33_ASAP7_75t_L g428 ( 
.A(n_187),
.B(n_8),
.Y(n_428)
);

CKINVDCx20_ASAP7_75t_R g429 ( 
.A(n_284),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_288),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_289),
.Y(n_431)
);

CKINVDCx5p33_ASAP7_75t_R g432 ( 
.A(n_295),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_332),
.Y(n_433)
);

CKINVDCx16_ASAP7_75t_R g434 ( 
.A(n_258),
.Y(n_434)
);

CKINVDCx20_ASAP7_75t_R g435 ( 
.A(n_326),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_335),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_336),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_337),
.Y(n_438)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_298),
.Y(n_439)
);

BUFx2_ASAP7_75t_L g440 ( 
.A(n_194),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_302),
.Y(n_441)
);

CKINVDCx16_ASAP7_75t_R g442 ( 
.A(n_314),
.Y(n_442)
);

INVx2_ASAP7_75t_L g443 ( 
.A(n_342),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_354),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_227),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_232),
.Y(n_446)
);

CKINVDCx5p33_ASAP7_75t_R g447 ( 
.A(n_366),
.Y(n_447)
);

CKINVDCx20_ASAP7_75t_R g448 ( 
.A(n_339),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_232),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_256),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_256),
.Y(n_451)
);

CKINVDCx20_ASAP7_75t_R g452 ( 
.A(n_349),
.Y(n_452)
);

CKINVDCx5p33_ASAP7_75t_R g453 ( 
.A(n_197),
.Y(n_453)
);

CKINVDCx20_ASAP7_75t_R g454 ( 
.A(n_303),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_270),
.Y(n_455)
);

BUFx2_ASAP7_75t_SL g456 ( 
.A(n_358),
.Y(n_456)
);

INVxp67_ASAP7_75t_SL g457 ( 
.A(n_270),
.Y(n_457)
);

CKINVDCx16_ASAP7_75t_R g458 ( 
.A(n_314),
.Y(n_458)
);

INVx2_ASAP7_75t_L g459 ( 
.A(n_367),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_377),
.Y(n_460)
);

AND2x4_ASAP7_75t_L g461 ( 
.A(n_378),
.B(n_292),
.Y(n_461)
);

BUFx6f_ASAP7_75t_L g462 ( 
.A(n_367),
.Y(n_462)
);

BUFx6f_ASAP7_75t_L g463 ( 
.A(n_367),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_L g464 ( 
.A(n_385),
.B(n_184),
.Y(n_464)
);

INVx2_ASAP7_75t_L g465 ( 
.A(n_367),
.Y(n_465)
);

BUFx2_ASAP7_75t_L g466 ( 
.A(n_453),
.Y(n_466)
);

INVx3_ASAP7_75t_L g467 ( 
.A(n_367),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_379),
.Y(n_468)
);

INVxp33_ASAP7_75t_SL g469 ( 
.A(n_369),
.Y(n_469)
);

NOR2xp33_ASAP7_75t_L g470 ( 
.A(n_456),
.B(n_188),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_384),
.Y(n_471)
);

AND2x2_ASAP7_75t_L g472 ( 
.A(n_445),
.B(n_446),
.Y(n_472)
);

INVx2_ASAP7_75t_L g473 ( 
.A(n_387),
.Y(n_473)
);

INVx3_ASAP7_75t_L g474 ( 
.A(n_393),
.Y(n_474)
);

INVx2_ASAP7_75t_L g475 ( 
.A(n_393),
.Y(n_475)
);

OA21x2_ASAP7_75t_L g476 ( 
.A1(n_394),
.A2(n_297),
.B(n_216),
.Y(n_476)
);

INVx6_ASAP7_75t_L g477 ( 
.A(n_402),
.Y(n_477)
);

INVx3_ASAP7_75t_L g478 ( 
.A(n_394),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_395),
.Y(n_479)
);

AND2x2_ASAP7_75t_L g480 ( 
.A(n_449),
.B(n_292),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_395),
.Y(n_481)
);

NOR2xp33_ASAP7_75t_L g482 ( 
.A(n_456),
.B(n_348),
.Y(n_482)
);

INVx3_ASAP7_75t_L g483 ( 
.A(n_413),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_413),
.Y(n_484)
);

INVxp67_ASAP7_75t_L g485 ( 
.A(n_389),
.Y(n_485)
);

OA21x2_ASAP7_75t_L g486 ( 
.A1(n_443),
.A2(n_297),
.B(n_216),
.Y(n_486)
);

INVx2_ASAP7_75t_L g487 ( 
.A(n_443),
.Y(n_487)
);

AND2x2_ASAP7_75t_L g488 ( 
.A(n_450),
.B(n_310),
.Y(n_488)
);

CKINVDCx14_ASAP7_75t_R g489 ( 
.A(n_369),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_388),
.Y(n_490)
);

INVx2_ASAP7_75t_L g491 ( 
.A(n_398),
.Y(n_491)
);

AOI22xp5_ASAP7_75t_SL g492 ( 
.A1(n_399),
.A2(n_363),
.B1(n_200),
.B2(n_253),
.Y(n_492)
);

NAND2xp33_ASAP7_75t_R g493 ( 
.A(n_453),
.B(n_197),
.Y(n_493)
);

AND2x4_ASAP7_75t_L g494 ( 
.A(n_423),
.B(n_310),
.Y(n_494)
);

NOR2xp33_ASAP7_75t_L g495 ( 
.A(n_380),
.B(n_195),
.Y(n_495)
);

INVxp67_ASAP7_75t_L g496 ( 
.A(n_440),
.Y(n_496)
);

NAND2xp33_ASAP7_75t_L g497 ( 
.A(n_402),
.B(n_273),
.Y(n_497)
);

INVx3_ASAP7_75t_L g498 ( 
.A(n_423),
.Y(n_498)
);

INVxp67_ASAP7_75t_L g499 ( 
.A(n_440),
.Y(n_499)
);

INVx2_ASAP7_75t_L g500 ( 
.A(n_400),
.Y(n_500)
);

INVx3_ASAP7_75t_L g501 ( 
.A(n_423),
.Y(n_501)
);

INVx2_ASAP7_75t_L g502 ( 
.A(n_401),
.Y(n_502)
);

INVx2_ASAP7_75t_L g503 ( 
.A(n_404),
.Y(n_503)
);

BUFx12f_ASAP7_75t_L g504 ( 
.A(n_370),
.Y(n_504)
);

INVx2_ASAP7_75t_L g505 ( 
.A(n_405),
.Y(n_505)
);

INVx2_ASAP7_75t_L g506 ( 
.A(n_411),
.Y(n_506)
);

AND3x2_ASAP7_75t_L g507 ( 
.A(n_428),
.B(n_341),
.C(n_323),
.Y(n_507)
);

INVx2_ASAP7_75t_L g508 ( 
.A(n_417),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_422),
.Y(n_509)
);

HB1xp67_ASAP7_75t_L g510 ( 
.A(n_376),
.Y(n_510)
);

AND2x4_ASAP7_75t_L g511 ( 
.A(n_451),
.B(n_323),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_425),
.Y(n_512)
);

AND2x2_ASAP7_75t_L g513 ( 
.A(n_455),
.B(n_341),
.Y(n_513)
);

INVx4_ASAP7_75t_L g514 ( 
.A(n_370),
.Y(n_514)
);

BUFx6f_ASAP7_75t_L g515 ( 
.A(n_426),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_433),
.Y(n_516)
);

CKINVDCx11_ASAP7_75t_R g517 ( 
.A(n_454),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_436),
.Y(n_518)
);

INVx2_ASAP7_75t_L g519 ( 
.A(n_437),
.Y(n_519)
);

INVx3_ASAP7_75t_L g520 ( 
.A(n_438),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_444),
.Y(n_521)
);

INVx2_ASAP7_75t_L g522 ( 
.A(n_368),
.Y(n_522)
);

INVx2_ASAP7_75t_L g523 ( 
.A(n_373),
.Y(n_523)
);

INVxp67_ASAP7_75t_L g524 ( 
.A(n_376),
.Y(n_524)
);

HB1xp67_ASAP7_75t_L g525 ( 
.A(n_418),
.Y(n_525)
);

CKINVDCx5p33_ASAP7_75t_R g526 ( 
.A(n_381),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_410),
.Y(n_527)
);

INVxp67_ASAP7_75t_L g528 ( 
.A(n_414),
.Y(n_528)
);

INVx2_ASAP7_75t_L g529 ( 
.A(n_374),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_457),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_375),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_415),
.Y(n_532)
);

NOR2xp33_ASAP7_75t_L g533 ( 
.A(n_382),
.B(n_273),
.Y(n_533)
);

INVx2_ASAP7_75t_L g534 ( 
.A(n_386),
.Y(n_534)
);

AND2x4_ASAP7_75t_L g535 ( 
.A(n_403),
.B(n_223),
.Y(n_535)
);

AND2x4_ASAP7_75t_L g536 ( 
.A(n_381),
.B(n_223),
.Y(n_536)
);

BUFx8_ASAP7_75t_L g537 ( 
.A(n_397),
.Y(n_537)
);

INVx2_ASAP7_75t_SL g538 ( 
.A(n_477),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_L g539 ( 
.A(n_536),
.B(n_383),
.Y(n_539)
);

AOI22xp33_ASAP7_75t_L g540 ( 
.A1(n_495),
.A2(n_315),
.B1(n_329),
.B2(n_333),
.Y(n_540)
);

INVxp67_ASAP7_75t_SL g541 ( 
.A(n_498),
.Y(n_541)
);

OR2x2_ASAP7_75t_L g542 ( 
.A(n_510),
.B(n_408),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_520),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_SL g544 ( 
.A(n_470),
.B(n_434),
.Y(n_544)
);

INVx2_ASAP7_75t_L g545 ( 
.A(n_473),
.Y(n_545)
);

OAI22x1_ASAP7_75t_L g546 ( 
.A1(n_496),
.A2(n_399),
.B1(n_224),
.B2(n_362),
.Y(n_546)
);

INVx3_ASAP7_75t_L g547 ( 
.A(n_462),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_L g548 ( 
.A(n_536),
.B(n_383),
.Y(n_548)
);

BUFx3_ASAP7_75t_L g549 ( 
.A(n_461),
.Y(n_549)
);

INVx2_ASAP7_75t_L g550 ( 
.A(n_473),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_520),
.Y(n_551)
);

AOI22xp33_ASAP7_75t_L g552 ( 
.A1(n_495),
.A2(n_533),
.B1(n_477),
.B2(n_530),
.Y(n_552)
);

HB1xp67_ASAP7_75t_L g553 ( 
.A(n_510),
.Y(n_553)
);

NOR2xp33_ASAP7_75t_L g554 ( 
.A(n_528),
.B(n_391),
.Y(n_554)
);

BUFx3_ASAP7_75t_L g555 ( 
.A(n_461),
.Y(n_555)
);

NAND3xp33_ASAP7_75t_L g556 ( 
.A(n_533),
.B(n_189),
.C(n_183),
.Y(n_556)
);

INVxp67_ASAP7_75t_SL g557 ( 
.A(n_498),
.Y(n_557)
);

INVx3_ASAP7_75t_L g558 ( 
.A(n_462),
.Y(n_558)
);

INVx3_ASAP7_75t_L g559 ( 
.A(n_462),
.Y(n_559)
);

AND2x2_ASAP7_75t_SL g560 ( 
.A(n_497),
.B(n_223),
.Y(n_560)
);

INVx2_ASAP7_75t_L g561 ( 
.A(n_473),
.Y(n_561)
);

INVx2_ASAP7_75t_L g562 ( 
.A(n_473),
.Y(n_562)
);

AOI22xp5_ASAP7_75t_L g563 ( 
.A1(n_497),
.A2(n_300),
.B1(n_299),
.B2(n_267),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_520),
.Y(n_564)
);

OR2x6_ASAP7_75t_L g565 ( 
.A(n_477),
.B(n_196),
.Y(n_565)
);

AND2x2_ASAP7_75t_L g566 ( 
.A(n_513),
.B(n_392),
.Y(n_566)
);

INVx1_ASAP7_75t_SL g567 ( 
.A(n_466),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_520),
.Y(n_568)
);

INVx1_ASAP7_75t_SL g569 ( 
.A(n_525),
.Y(n_569)
);

AOI22xp33_ASAP7_75t_L g570 ( 
.A1(n_477),
.A2(n_262),
.B1(n_329),
.B2(n_333),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_520),
.Y(n_571)
);

INVx2_ASAP7_75t_L g572 ( 
.A(n_468),
.Y(n_572)
);

INVx4_ASAP7_75t_SL g573 ( 
.A(n_477),
.Y(n_573)
);

INVx2_ASAP7_75t_L g574 ( 
.A(n_468),
.Y(n_574)
);

INVx2_ASAP7_75t_L g575 ( 
.A(n_468),
.Y(n_575)
);

AOI22xp33_ASAP7_75t_L g576 ( 
.A1(n_477),
.A2(n_262),
.B1(n_329),
.B2(n_333),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_460),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_460),
.Y(n_578)
);

CKINVDCx5p33_ASAP7_75t_R g579 ( 
.A(n_504),
.Y(n_579)
);

NOR2xp33_ASAP7_75t_L g580 ( 
.A(n_528),
.B(n_527),
.Y(n_580)
);

BUFx3_ASAP7_75t_L g581 ( 
.A(n_461),
.Y(n_581)
);

AOI22xp33_ASAP7_75t_L g582 ( 
.A1(n_477),
.A2(n_262),
.B1(n_329),
.B2(n_333),
.Y(n_582)
);

INVx2_ASAP7_75t_L g583 ( 
.A(n_471),
.Y(n_583)
);

BUFx6f_ASAP7_75t_L g584 ( 
.A(n_462),
.Y(n_584)
);

NAND2xp5_ASAP7_75t_SL g585 ( 
.A(n_470),
.B(n_442),
.Y(n_585)
);

INVx3_ASAP7_75t_L g586 ( 
.A(n_462),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_L g587 ( 
.A(n_536),
.B(n_392),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_L g588 ( 
.A(n_536),
.B(n_396),
.Y(n_588)
);

OR2x6_ASAP7_75t_L g589 ( 
.A(n_504),
.B(n_199),
.Y(n_589)
);

INVx2_ASAP7_75t_L g590 ( 
.A(n_471),
.Y(n_590)
);

AND2x6_ASAP7_75t_L g591 ( 
.A(n_536),
.B(n_223),
.Y(n_591)
);

AND2x4_ASAP7_75t_L g592 ( 
.A(n_494),
.B(n_201),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_L g593 ( 
.A(n_482),
.B(n_396),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_SL g594 ( 
.A(n_482),
.B(n_458),
.Y(n_594)
);

INVx2_ASAP7_75t_SL g595 ( 
.A(n_525),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_L g596 ( 
.A(n_527),
.B(n_530),
.Y(n_596)
);

BUFx3_ASAP7_75t_L g597 ( 
.A(n_461),
.Y(n_597)
);

OAI22xp33_ASAP7_75t_L g598 ( 
.A1(n_534),
.A2(n_350),
.B1(n_204),
.B2(n_225),
.Y(n_598)
);

AOI22xp33_ASAP7_75t_L g599 ( 
.A1(n_527),
.A2(n_262),
.B1(n_313),
.B2(n_315),
.Y(n_599)
);

OR2x6_ASAP7_75t_L g600 ( 
.A(n_504),
.B(n_213),
.Y(n_600)
);

INVx4_ASAP7_75t_L g601 ( 
.A(n_486),
.Y(n_601)
);

INVx2_ASAP7_75t_L g602 ( 
.A(n_471),
.Y(n_602)
);

INVx3_ASAP7_75t_L g603 ( 
.A(n_462),
.Y(n_603)
);

BUFx3_ASAP7_75t_L g604 ( 
.A(n_461),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_SL g605 ( 
.A(n_534),
.B(n_406),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_522),
.Y(n_606)
);

OAI21xp33_ASAP7_75t_SL g607 ( 
.A1(n_530),
.A2(n_319),
.B(n_235),
.Y(n_607)
);

OR2x6_ASAP7_75t_L g608 ( 
.A(n_504),
.B(n_218),
.Y(n_608)
);

INVx2_ASAP7_75t_L g609 ( 
.A(n_475),
.Y(n_609)
);

AOI22xp33_ASAP7_75t_L g610 ( 
.A1(n_511),
.A2(n_315),
.B1(n_329),
.B2(n_333),
.Y(n_610)
);

INVx2_ASAP7_75t_L g611 ( 
.A(n_475),
.Y(n_611)
);

INVx2_ASAP7_75t_SL g612 ( 
.A(n_507),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_522),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_SL g614 ( 
.A(n_534),
.B(n_406),
.Y(n_614)
);

AO21x2_ASAP7_75t_L g615 ( 
.A1(n_464),
.A2(n_222),
.B(n_219),
.Y(n_615)
);

INVx3_ASAP7_75t_L g616 ( 
.A(n_462),
.Y(n_616)
);

INVx2_ASAP7_75t_L g617 ( 
.A(n_475),
.Y(n_617)
);

BUFx10_ASAP7_75t_L g618 ( 
.A(n_526),
.Y(n_618)
);

INVx3_ASAP7_75t_L g619 ( 
.A(n_462),
.Y(n_619)
);

NOR2xp33_ASAP7_75t_L g620 ( 
.A(n_464),
.B(n_407),
.Y(n_620)
);

BUFx3_ASAP7_75t_L g621 ( 
.A(n_461),
.Y(n_621)
);

INVx2_ASAP7_75t_L g622 ( 
.A(n_475),
.Y(n_622)
);

INVx2_ASAP7_75t_L g623 ( 
.A(n_487),
.Y(n_623)
);

BUFx6f_ASAP7_75t_L g624 ( 
.A(n_462),
.Y(n_624)
);

INVx3_ASAP7_75t_L g625 ( 
.A(n_463),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_SL g626 ( 
.A(n_534),
.B(n_514),
.Y(n_626)
);

OR2x6_ASAP7_75t_L g627 ( 
.A(n_514),
.B(n_228),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_L g628 ( 
.A(n_494),
.B(n_409),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_522),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_SL g630 ( 
.A(n_514),
.B(n_409),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_522),
.Y(n_631)
);

NOR2xp33_ASAP7_75t_SL g632 ( 
.A(n_514),
.B(n_347),
.Y(n_632)
);

AO22x2_ASAP7_75t_L g633 ( 
.A1(n_496),
.A2(n_246),
.B1(n_252),
.B2(n_230),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_L g634 ( 
.A(n_494),
.B(n_416),
.Y(n_634)
);

INVx2_ASAP7_75t_L g635 ( 
.A(n_487),
.Y(n_635)
);

INVx3_ASAP7_75t_L g636 ( 
.A(n_463),
.Y(n_636)
);

INVx2_ASAP7_75t_L g637 ( 
.A(n_487),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_523),
.Y(n_638)
);

AND2x2_ASAP7_75t_SL g639 ( 
.A(n_486),
.B(n_262),
.Y(n_639)
);

INVxp33_ASAP7_75t_SL g640 ( 
.A(n_492),
.Y(n_640)
);

INVx2_ASAP7_75t_L g641 ( 
.A(n_487),
.Y(n_641)
);

BUFx3_ASAP7_75t_L g642 ( 
.A(n_494),
.Y(n_642)
);

OR2x6_ASAP7_75t_L g643 ( 
.A(n_514),
.B(n_254),
.Y(n_643)
);

INVx5_ASAP7_75t_L g644 ( 
.A(n_463),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_L g645 ( 
.A(n_494),
.B(n_416),
.Y(n_645)
);

INVx2_ASAP7_75t_L g646 ( 
.A(n_474),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_SL g647 ( 
.A(n_514),
.B(n_419),
.Y(n_647)
);

AOI22xp33_ASAP7_75t_L g648 ( 
.A1(n_511),
.A2(n_313),
.B1(n_315),
.B2(n_397),
.Y(n_648)
);

AND2x6_ASAP7_75t_L g649 ( 
.A(n_535),
.B(n_313),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_523),
.Y(n_650)
);

AND2x2_ASAP7_75t_SL g651 ( 
.A(n_486),
.B(n_313),
.Y(n_651)
);

AND2x2_ASAP7_75t_SL g652 ( 
.A(n_486),
.B(n_313),
.Y(n_652)
);

INVx2_ASAP7_75t_L g653 ( 
.A(n_474),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_523),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_523),
.Y(n_655)
);

INVx2_ASAP7_75t_L g656 ( 
.A(n_474),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_529),
.Y(n_657)
);

INVx2_ASAP7_75t_L g658 ( 
.A(n_474),
.Y(n_658)
);

INVx2_ASAP7_75t_L g659 ( 
.A(n_474),
.Y(n_659)
);

INVx2_ASAP7_75t_L g660 ( 
.A(n_478),
.Y(n_660)
);

INVxp67_ASAP7_75t_SL g661 ( 
.A(n_498),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_529),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_529),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_L g664 ( 
.A(n_498),
.B(n_419),
.Y(n_664)
);

AND3x2_ASAP7_75t_L g665 ( 
.A(n_466),
.B(n_268),
.C(n_263),
.Y(n_665)
);

INVx4_ASAP7_75t_L g666 ( 
.A(n_486),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_SL g667 ( 
.A(n_537),
.B(n_420),
.Y(n_667)
);

NAND2xp33_ASAP7_75t_L g668 ( 
.A(n_531),
.B(n_420),
.Y(n_668)
);

BUFx2_ASAP7_75t_L g669 ( 
.A(n_524),
.Y(n_669)
);

NAND2xp33_ASAP7_75t_L g670 ( 
.A(n_531),
.B(n_421),
.Y(n_670)
);

NOR2xp33_ASAP7_75t_L g671 ( 
.A(n_524),
.B(n_421),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_529),
.Y(n_672)
);

NAND2xp33_ASAP7_75t_SL g673 ( 
.A(n_493),
.B(n_427),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_498),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_L g675 ( 
.A(n_501),
.B(n_427),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_L g676 ( 
.A(n_501),
.B(n_507),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_SL g677 ( 
.A(n_537),
.B(n_430),
.Y(n_677)
);

INVx2_ASAP7_75t_L g678 ( 
.A(n_478),
.Y(n_678)
);

BUFx6f_ASAP7_75t_L g679 ( 
.A(n_463),
.Y(n_679)
);

OAI22xp33_ASAP7_75t_L g680 ( 
.A1(n_499),
.A2(n_485),
.B1(n_493),
.B2(n_532),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_SL g681 ( 
.A(n_537),
.B(n_430),
.Y(n_681)
);

INVx4_ASAP7_75t_L g682 ( 
.A(n_486),
.Y(n_682)
);

BUFx6f_ASAP7_75t_L g683 ( 
.A(n_463),
.Y(n_683)
);

AND2x6_ASAP7_75t_L g684 ( 
.A(n_535),
.B(n_315),
.Y(n_684)
);

INVx2_ASAP7_75t_L g685 ( 
.A(n_478),
.Y(n_685)
);

AND2x2_ASAP7_75t_L g686 ( 
.A(n_513),
.B(n_431),
.Y(n_686)
);

AND2x2_ASAP7_75t_SL g687 ( 
.A(n_476),
.B(n_269),
.Y(n_687)
);

OR2x2_ASAP7_75t_L g688 ( 
.A(n_499),
.B(n_431),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_SL g689 ( 
.A(n_560),
.B(n_501),
.Y(n_689)
);

AOI22xp5_ASAP7_75t_L g690 ( 
.A1(n_620),
.A2(n_466),
.B1(n_485),
.B2(n_412),
.Y(n_690)
);

AOI22xp5_ASAP7_75t_L g691 ( 
.A1(n_632),
.A2(n_424),
.B1(n_372),
.B2(n_371),
.Y(n_691)
);

NAND2xp33_ASAP7_75t_L g692 ( 
.A(n_570),
.B(n_282),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_SL g693 ( 
.A(n_560),
.B(n_501),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_L g694 ( 
.A(n_552),
.B(n_501),
.Y(n_694)
);

INVx2_ASAP7_75t_L g695 ( 
.A(n_572),
.Y(n_695)
);

NOR2xp33_ASAP7_75t_L g696 ( 
.A(n_593),
.B(n_469),
.Y(n_696)
);

INVx2_ASAP7_75t_L g697 ( 
.A(n_572),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_674),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_L g699 ( 
.A(n_580),
.B(n_535),
.Y(n_699)
);

AND2x4_ASAP7_75t_L g700 ( 
.A(n_642),
.B(n_472),
.Y(n_700)
);

AND2x6_ASAP7_75t_L g701 ( 
.A(n_642),
.B(n_535),
.Y(n_701)
);

NOR3xp33_ASAP7_75t_L g702 ( 
.A(n_673),
.B(n_489),
.C(n_439),
.Y(n_702)
);

NOR2xp33_ASAP7_75t_L g703 ( 
.A(n_554),
.B(n_469),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_L g704 ( 
.A(n_560),
.B(n_541),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_SL g705 ( 
.A(n_687),
.B(n_535),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_SL g706 ( 
.A(n_687),
.B(n_535),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_642),
.Y(n_707)
);

OAI221xp5_ASAP7_75t_L g708 ( 
.A1(n_556),
.A2(n_532),
.B1(n_531),
.B2(n_509),
.C(n_521),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_577),
.Y(n_709)
);

INVx2_ASAP7_75t_L g710 ( 
.A(n_574),
.Y(n_710)
);

INVx3_ASAP7_75t_L g711 ( 
.A(n_549),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_577),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_L g713 ( 
.A(n_557),
.B(n_532),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_L g714 ( 
.A(n_661),
.B(n_513),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_SL g715 ( 
.A(n_687),
.B(n_537),
.Y(n_715)
);

AOI22xp33_ASAP7_75t_L g716 ( 
.A1(n_615),
.A2(n_511),
.B1(n_476),
.B2(n_472),
.Y(n_716)
);

AOI22xp33_ASAP7_75t_L g717 ( 
.A1(n_615),
.A2(n_511),
.B1(n_476),
.B2(n_472),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_L g718 ( 
.A(n_538),
.B(n_511),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_SL g719 ( 
.A(n_632),
.B(n_537),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_L g720 ( 
.A(n_538),
.B(n_511),
.Y(n_720)
);

NAND3xp33_ASAP7_75t_L g721 ( 
.A(n_668),
.B(n_439),
.C(n_432),
.Y(n_721)
);

NOR3xp33_ASAP7_75t_L g722 ( 
.A(n_544),
.B(n_489),
.C(n_441),
.Y(n_722)
);

INVxp67_ASAP7_75t_L g723 ( 
.A(n_671),
.Y(n_723)
);

AND2x4_ASAP7_75t_L g724 ( 
.A(n_549),
.B(n_480),
.Y(n_724)
);

INVx2_ASAP7_75t_L g725 ( 
.A(n_574),
.Y(n_725)
);

NOR2xp33_ASAP7_75t_L g726 ( 
.A(n_569),
.B(n_432),
.Y(n_726)
);

INVx2_ASAP7_75t_L g727 ( 
.A(n_575),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_L g728 ( 
.A(n_596),
.B(n_515),
.Y(n_728)
);

INVx3_ASAP7_75t_L g729 ( 
.A(n_549),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_L g730 ( 
.A(n_626),
.B(n_515),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_L g731 ( 
.A(n_664),
.B(n_515),
.Y(n_731)
);

INVx2_ASAP7_75t_L g732 ( 
.A(n_575),
.Y(n_732)
);

INVx2_ASAP7_75t_L g733 ( 
.A(n_583),
.Y(n_733)
);

NOR2xp33_ASAP7_75t_L g734 ( 
.A(n_569),
.B(n_441),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_L g735 ( 
.A(n_675),
.B(n_515),
.Y(n_735)
);

OR2x2_ASAP7_75t_L g736 ( 
.A(n_553),
.B(n_447),
.Y(n_736)
);

INVxp67_ASAP7_75t_L g737 ( 
.A(n_669),
.Y(n_737)
);

INVx2_ASAP7_75t_L g738 ( 
.A(n_583),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_L g739 ( 
.A(n_639),
.B(n_515),
.Y(n_739)
);

NAND3xp33_ASAP7_75t_L g740 ( 
.A(n_670),
.B(n_447),
.C(n_480),
.Y(n_740)
);

INVx3_ASAP7_75t_L g741 ( 
.A(n_555),
.Y(n_741)
);

AOI22xp5_ASAP7_75t_L g742 ( 
.A1(n_539),
.A2(n_390),
.B1(n_429),
.B2(n_435),
.Y(n_742)
);

INVx2_ASAP7_75t_SL g743 ( 
.A(n_595),
.Y(n_743)
);

OR2x6_ASAP7_75t_L g744 ( 
.A(n_589),
.B(n_480),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_SL g745 ( 
.A(n_548),
.B(n_537),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_L g746 ( 
.A(n_639),
.B(n_651),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_L g747 ( 
.A(n_639),
.B(n_515),
.Y(n_747)
);

NAND2xp33_ASAP7_75t_L g748 ( 
.A(n_576),
.B(n_287),
.Y(n_748)
);

NOR3xp33_ASAP7_75t_L g749 ( 
.A(n_585),
.B(n_517),
.C(n_488),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_578),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_L g751 ( 
.A(n_651),
.B(n_515),
.Y(n_751)
);

AOI22xp33_ASAP7_75t_L g752 ( 
.A1(n_615),
.A2(n_476),
.B1(n_515),
.B2(n_488),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_578),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_555),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_L g755 ( 
.A(n_651),
.B(n_488),
.Y(n_755)
);

AOI22xp5_ASAP7_75t_L g756 ( 
.A1(n_587),
.A2(n_452),
.B1(n_448),
.B2(n_271),
.Y(n_756)
);

NAND2xp33_ASAP7_75t_L g757 ( 
.A(n_582),
.B(n_306),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_555),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_L g759 ( 
.A(n_652),
.B(n_478),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_L g760 ( 
.A(n_652),
.B(n_483),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_L g761 ( 
.A(n_592),
.B(n_588),
.Y(n_761)
);

INVx2_ASAP7_75t_L g762 ( 
.A(n_590),
.Y(n_762)
);

AND2x2_ASAP7_75t_L g763 ( 
.A(n_595),
.B(n_512),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_L g764 ( 
.A(n_592),
.B(n_483),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_L g765 ( 
.A(n_592),
.B(n_483),
.Y(n_765)
);

INVxp67_ASAP7_75t_SL g766 ( 
.A(n_584),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_SL g767 ( 
.A(n_581),
.B(n_308),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_581),
.Y(n_768)
);

INVxp33_ASAP7_75t_L g769 ( 
.A(n_566),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_L g770 ( 
.A(n_628),
.B(n_483),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_L g771 ( 
.A(n_634),
.B(n_483),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_581),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_L g773 ( 
.A(n_645),
.B(n_491),
.Y(n_773)
);

NOR2xp33_ASAP7_75t_L g774 ( 
.A(n_688),
.B(n_397),
.Y(n_774)
);

INVx2_ASAP7_75t_L g775 ( 
.A(n_590),
.Y(n_775)
);

OAI22xp5_ASAP7_75t_SL g776 ( 
.A1(n_640),
.A2(n_492),
.B1(n_211),
.B2(n_220),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_597),
.Y(n_777)
);

INVx2_ASAP7_75t_L g778 ( 
.A(n_602),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_L g779 ( 
.A(n_601),
.B(n_491),
.Y(n_779)
);

INVx3_ASAP7_75t_L g780 ( 
.A(n_597),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_SL g781 ( 
.A(n_597),
.B(n_309),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_L g782 ( 
.A(n_601),
.B(n_491),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_L g783 ( 
.A(n_601),
.B(n_491),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_L g784 ( 
.A(n_601),
.B(n_500),
.Y(n_784)
);

INVxp67_ASAP7_75t_L g785 ( 
.A(n_669),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_604),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_604),
.Y(n_787)
);

AND2x2_ASAP7_75t_L g788 ( 
.A(n_566),
.B(n_512),
.Y(n_788)
);

BUFx12f_ASAP7_75t_L g789 ( 
.A(n_618),
.Y(n_789)
);

BUFx8_ASAP7_75t_L g790 ( 
.A(n_542),
.Y(n_790)
);

BUFx2_ASAP7_75t_L g791 ( 
.A(n_542),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_SL g792 ( 
.A(n_604),
.B(n_324),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_L g793 ( 
.A(n_666),
.B(n_500),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_L g794 ( 
.A(n_666),
.B(n_500),
.Y(n_794)
);

NOR2xp33_ASAP7_75t_L g795 ( 
.A(n_688),
.B(n_184),
.Y(n_795)
);

NAND2x1_ASAP7_75t_L g796 ( 
.A(n_547),
.B(n_476),
.Y(n_796)
);

AOI22xp33_ASAP7_75t_L g797 ( 
.A1(n_556),
.A2(n_476),
.B1(n_355),
.B2(n_327),
.Y(n_797)
);

INVx2_ASAP7_75t_L g798 ( 
.A(n_602),
.Y(n_798)
);

OR2x6_ASAP7_75t_L g799 ( 
.A(n_589),
.B(n_516),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_L g800 ( 
.A(n_666),
.B(n_500),
.Y(n_800)
);

NOR2xp33_ASAP7_75t_L g801 ( 
.A(n_594),
.B(n_193),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_L g802 ( 
.A(n_666),
.B(n_502),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_L g803 ( 
.A(n_682),
.B(n_502),
.Y(n_803)
);

NOR2xp33_ASAP7_75t_L g804 ( 
.A(n_605),
.B(n_193),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_SL g805 ( 
.A(n_621),
.B(n_364),
.Y(n_805)
);

INVx2_ASAP7_75t_SL g806 ( 
.A(n_686),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_621),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_L g808 ( 
.A(n_682),
.B(n_502),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_L g809 ( 
.A(n_682),
.B(n_502),
.Y(n_809)
);

AND2x4_ASAP7_75t_L g810 ( 
.A(n_621),
.B(n_516),
.Y(n_810)
);

NOR2xp33_ASAP7_75t_L g811 ( 
.A(n_614),
.B(n_680),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_L g812 ( 
.A(n_682),
.B(n_503),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_SL g813 ( 
.A(n_676),
.B(n_237),
.Y(n_813)
);

AOI22xp33_ASAP7_75t_L g814 ( 
.A1(n_591),
.A2(n_503),
.B1(n_519),
.B2(n_505),
.Y(n_814)
);

INVx4_ASAP7_75t_L g815 ( 
.A(n_573),
.Y(n_815)
);

NOR2xp33_ASAP7_75t_L g816 ( 
.A(n_612),
.B(n_202),
.Y(n_816)
);

NOR2xp67_ASAP7_75t_L g817 ( 
.A(n_579),
.B(n_490),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_SL g818 ( 
.A(n_543),
.B(n_241),
.Y(n_818)
);

AND2x2_ASAP7_75t_L g819 ( 
.A(n_686),
.B(n_490),
.Y(n_819)
);

AOI221xp5_ASAP7_75t_L g820 ( 
.A1(n_598),
.A2(n_224),
.B1(n_362),
.B2(n_361),
.C(n_359),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_L g821 ( 
.A(n_551),
.B(n_503),
.Y(n_821)
);

AND2x2_ASAP7_75t_L g822 ( 
.A(n_567),
.B(n_490),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_L g823 ( 
.A(n_551),
.B(n_505),
.Y(n_823)
);

CKINVDCx5p33_ASAP7_75t_R g824 ( 
.A(n_618),
.Y(n_824)
);

OAI21xp5_ASAP7_75t_L g825 ( 
.A1(n_564),
.A2(n_465),
.B(n_459),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_SL g826 ( 
.A(n_564),
.B(n_245),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_SL g827 ( 
.A(n_568),
.B(n_259),
.Y(n_827)
);

O2A1O1Ixp33_ASAP7_75t_L g828 ( 
.A1(n_607),
.A2(n_521),
.B(n_509),
.C(n_518),
.Y(n_828)
);

O2A1O1Ixp5_ASAP7_75t_L g829 ( 
.A1(n_568),
.A2(n_465),
.B(n_459),
.C(n_519),
.Y(n_829)
);

NOR2xp33_ASAP7_75t_L g830 ( 
.A(n_612),
.B(n_202),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_571),
.Y(n_831)
);

INVx2_ASAP7_75t_L g832 ( 
.A(n_623),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_SL g833 ( 
.A(n_571),
.B(n_573),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_L g834 ( 
.A(n_540),
.B(n_505),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_646),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_L g836 ( 
.A(n_646),
.B(n_505),
.Y(n_836)
);

OR2x2_ASAP7_75t_L g837 ( 
.A(n_563),
.B(n_546),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_653),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_L g839 ( 
.A(n_656),
.B(n_506),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_L g840 ( 
.A(n_656),
.B(n_506),
.Y(n_840)
);

INVx2_ASAP7_75t_L g841 ( 
.A(n_623),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_L g842 ( 
.A(n_658),
.B(n_506),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_SL g843 ( 
.A(n_573),
.B(n_260),
.Y(n_843)
);

NOR2x1p5_ASAP7_75t_L g844 ( 
.A(n_579),
.B(n_198),
.Y(n_844)
);

CKINVDCx5p33_ASAP7_75t_R g845 ( 
.A(n_618),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_L g846 ( 
.A(n_658),
.B(n_506),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_SL g847 ( 
.A(n_573),
.B(n_272),
.Y(n_847)
);

AND2x2_ASAP7_75t_L g848 ( 
.A(n_563),
.B(n_509),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_L g849 ( 
.A(n_659),
.B(n_508),
.Y(n_849)
);

NAND2xp33_ASAP7_75t_SL g850 ( 
.A(n_648),
.B(n_198),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_SL g851 ( 
.A(n_659),
.B(n_277),
.Y(n_851)
);

INVxp67_ASAP7_75t_L g852 ( 
.A(n_546),
.Y(n_852)
);

AOI22xp33_ASAP7_75t_SL g853 ( 
.A1(n_640),
.A2(n_347),
.B1(n_353),
.B2(n_314),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_660),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_SL g855 ( 
.A(n_660),
.B(n_281),
.Y(n_855)
);

AOI21xp5_ASAP7_75t_L g856 ( 
.A1(n_746),
.A2(n_565),
.B(n_678),
.Y(n_856)
);

AOI21x1_ASAP7_75t_L g857 ( 
.A1(n_796),
.A2(n_565),
.B(n_606),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_SL g858 ( 
.A(n_723),
.B(n_726),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_L g859 ( 
.A(n_699),
.B(n_630),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_L g860 ( 
.A(n_709),
.B(n_647),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_L g861 ( 
.A(n_712),
.B(n_591),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_L g862 ( 
.A(n_750),
.B(n_591),
.Y(n_862)
);

AOI21xp5_ASAP7_75t_L g863 ( 
.A1(n_739),
.A2(n_565),
.B(n_678),
.Y(n_863)
);

NOR2xp33_ASAP7_75t_L g864 ( 
.A(n_703),
.B(n_696),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_L g865 ( 
.A(n_753),
.B(n_591),
.Y(n_865)
);

AOI21xp5_ASAP7_75t_L g866 ( 
.A1(n_747),
.A2(n_565),
.B(n_685),
.Y(n_866)
);

AOI21xp5_ASAP7_75t_L g867 ( 
.A1(n_751),
.A2(n_565),
.B(n_685),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_L g868 ( 
.A(n_714),
.B(n_591),
.Y(n_868)
);

AOI21xp5_ASAP7_75t_L g869 ( 
.A1(n_705),
.A2(n_610),
.B(n_606),
.Y(n_869)
);

AOI21xp5_ASAP7_75t_L g870 ( 
.A1(n_705),
.A2(n_629),
.B(n_613),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_L g871 ( 
.A(n_713),
.B(n_755),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_831),
.Y(n_872)
);

AOI21xp5_ASAP7_75t_L g873 ( 
.A1(n_706),
.A2(n_629),
.B(n_613),
.Y(n_873)
);

AOI21xp5_ASAP7_75t_L g874 ( 
.A1(n_706),
.A2(n_638),
.B(n_631),
.Y(n_874)
);

INVx3_ASAP7_75t_L g875 ( 
.A(n_729),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_L g876 ( 
.A(n_819),
.B(n_591),
.Y(n_876)
);

AND2x2_ASAP7_75t_L g877 ( 
.A(n_822),
.B(n_618),
.Y(n_877)
);

INVx2_ASAP7_75t_L g878 ( 
.A(n_695),
.Y(n_878)
);

AOI21xp5_ASAP7_75t_L g879 ( 
.A1(n_761),
.A2(n_624),
.B(n_584),
.Y(n_879)
);

A2O1A1Ixp33_ASAP7_75t_L g880 ( 
.A1(n_811),
.A2(n_804),
.B(n_795),
.C(n_801),
.Y(n_880)
);

OAI21xp5_ASAP7_75t_L g881 ( 
.A1(n_759),
.A2(n_643),
.B(n_627),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_698),
.Y(n_882)
);

NAND2xp5_ASAP7_75t_L g883 ( 
.A(n_763),
.B(n_591),
.Y(n_883)
);

OAI21xp33_ASAP7_75t_L g884 ( 
.A1(n_734),
.A2(n_607),
.B(n_633),
.Y(n_884)
);

INVx3_ASAP7_75t_L g885 ( 
.A(n_729),
.Y(n_885)
);

AOI21xp5_ASAP7_75t_L g886 ( 
.A1(n_731),
.A2(n_624),
.B(n_584),
.Y(n_886)
);

NOR2xp33_ASAP7_75t_L g887 ( 
.A(n_769),
.B(n_667),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_L g888 ( 
.A(n_724),
.B(n_627),
.Y(n_888)
);

INVx2_ASAP7_75t_SL g889 ( 
.A(n_743),
.Y(n_889)
);

AOI21xp5_ASAP7_75t_L g890 ( 
.A1(n_735),
.A2(n_624),
.B(n_584),
.Y(n_890)
);

NOR2xp33_ASAP7_75t_L g891 ( 
.A(n_769),
.B(n_677),
.Y(n_891)
);

O2A1O1Ixp33_ASAP7_75t_L g892 ( 
.A1(n_694),
.A2(n_643),
.B(n_627),
.C(n_681),
.Y(n_892)
);

AND2x4_ASAP7_75t_SL g893 ( 
.A(n_724),
.B(n_589),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_L g894 ( 
.A(n_724),
.B(n_810),
.Y(n_894)
);

AOI21xp5_ASAP7_75t_L g895 ( 
.A1(n_773),
.A2(n_679),
.B(n_624),
.Y(n_895)
);

AND2x2_ASAP7_75t_L g896 ( 
.A(n_788),
.B(n_589),
.Y(n_896)
);

INVx2_ASAP7_75t_L g897 ( 
.A(n_695),
.Y(n_897)
);

CKINVDCx5p33_ASAP7_75t_R g898 ( 
.A(n_789),
.Y(n_898)
);

NAND2xp5_ASAP7_75t_SL g899 ( 
.A(n_806),
.B(n_203),
.Y(n_899)
);

OAI22xp5_ASAP7_75t_L g900 ( 
.A1(n_704),
.A2(n_627),
.B1(n_643),
.B2(n_599),
.Y(n_900)
);

BUFx6f_ASAP7_75t_L g901 ( 
.A(n_700),
.Y(n_901)
);

NAND2xp33_ASAP7_75t_R g902 ( 
.A(n_791),
.B(n_736),
.Y(n_902)
);

INVx2_ASAP7_75t_L g903 ( 
.A(n_697),
.Y(n_903)
);

AOI21xp5_ASAP7_75t_L g904 ( 
.A1(n_779),
.A2(n_683),
.B(n_679),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_L g905 ( 
.A(n_810),
.B(n_627),
.Y(n_905)
);

AOI22xp5_ASAP7_75t_L g906 ( 
.A1(n_700),
.A2(n_643),
.B1(n_600),
.B2(n_589),
.Y(n_906)
);

NOR3xp33_ASAP7_75t_L g907 ( 
.A(n_721),
.B(n_517),
.C(n_518),
.Y(n_907)
);

AOI21xp5_ASAP7_75t_L g908 ( 
.A1(n_782),
.A2(n_683),
.B(n_679),
.Y(n_908)
);

AOI33xp33_ASAP7_75t_L g909 ( 
.A1(n_853),
.A2(n_665),
.A3(n_521),
.B1(n_518),
.B2(n_479),
.B3(n_484),
.Y(n_909)
);

AOI21xp5_ASAP7_75t_L g910 ( 
.A1(n_783),
.A2(n_683),
.B(n_679),
.Y(n_910)
);

NAND2xp5_ASAP7_75t_L g911 ( 
.A(n_810),
.B(n_643),
.Y(n_911)
);

NOR2xp67_ASAP7_75t_L g912 ( 
.A(n_824),
.B(n_650),
.Y(n_912)
);

INVx2_ASAP7_75t_L g913 ( 
.A(n_697),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_SL g914 ( 
.A(n_700),
.B(n_203),
.Y(n_914)
);

NOR2xp33_ASAP7_75t_L g915 ( 
.A(n_737),
.B(n_600),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_L g916 ( 
.A(n_711),
.B(n_633),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_L g917 ( 
.A(n_711),
.B(n_633),
.Y(n_917)
);

A2O1A1Ixp33_ASAP7_75t_L g918 ( 
.A1(n_816),
.A2(n_655),
.B(n_654),
.C(n_657),
.Y(n_918)
);

INVx3_ASAP7_75t_L g919 ( 
.A(n_729),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_L g920 ( 
.A(n_741),
.B(n_633),
.Y(n_920)
);

INVx3_ASAP7_75t_L g921 ( 
.A(n_780),
.Y(n_921)
);

AOI21xp5_ASAP7_75t_L g922 ( 
.A1(n_784),
.A2(n_683),
.B(n_679),
.Y(n_922)
);

BUFx12f_ASAP7_75t_L g923 ( 
.A(n_790),
.Y(n_923)
);

INVx11_ASAP7_75t_L g924 ( 
.A(n_789),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_SL g925 ( 
.A(n_817),
.B(n_205),
.Y(n_925)
);

AND2x2_ASAP7_75t_SL g926 ( 
.A(n_691),
.B(n_600),
.Y(n_926)
);

NAND2xp5_ASAP7_75t_L g927 ( 
.A(n_741),
.B(n_547),
.Y(n_927)
);

AOI21xp5_ASAP7_75t_L g928 ( 
.A1(n_793),
.A2(n_683),
.B(n_644),
.Y(n_928)
);

OAI21xp5_ASAP7_75t_L g929 ( 
.A1(n_760),
.A2(n_663),
.B(n_662),
.Y(n_929)
);

BUFx6f_ASAP7_75t_L g930 ( 
.A(n_780),
.Y(n_930)
);

NAND2xp5_ASAP7_75t_SL g931 ( 
.A(n_690),
.B(n_205),
.Y(n_931)
);

AOI21xp5_ASAP7_75t_L g932 ( 
.A1(n_794),
.A2(n_644),
.B(n_547),
.Y(n_932)
);

AOI22xp5_ASAP7_75t_L g933 ( 
.A1(n_754),
.A2(n_600),
.B1(n_608),
.B2(n_649),
.Y(n_933)
);

O2A1O1Ixp33_ASAP7_75t_L g934 ( 
.A1(n_708),
.A2(n_672),
.B(n_663),
.C(n_609),
.Y(n_934)
);

NAND2xp5_ASAP7_75t_L g935 ( 
.A(n_780),
.B(n_558),
.Y(n_935)
);

NAND2xp5_ASAP7_75t_SL g936 ( 
.A(n_848),
.B(n_206),
.Y(n_936)
);

INVx2_ASAP7_75t_L g937 ( 
.A(n_710),
.Y(n_937)
);

NOR2xp33_ASAP7_75t_L g938 ( 
.A(n_785),
.B(n_600),
.Y(n_938)
);

AOI22xp33_ASAP7_75t_L g939 ( 
.A1(n_701),
.A2(n_684),
.B1(n_649),
.B2(n_672),
.Y(n_939)
);

AOI21xp5_ASAP7_75t_L g940 ( 
.A1(n_800),
.A2(n_644),
.B(n_619),
.Y(n_940)
);

NOR2xp33_ASAP7_75t_L g941 ( 
.A(n_830),
.B(n_608),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_L g942 ( 
.A(n_770),
.B(n_558),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_SL g943 ( 
.A(n_740),
.B(n_206),
.Y(n_943)
);

INVxp67_ASAP7_75t_L g944 ( 
.A(n_774),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_L g945 ( 
.A(n_771),
.B(n_558),
.Y(n_945)
);

INVxp67_ASAP7_75t_L g946 ( 
.A(n_742),
.Y(n_946)
);

NAND2xp5_ASAP7_75t_L g947 ( 
.A(n_802),
.B(n_559),
.Y(n_947)
);

AND2x4_ASAP7_75t_L g948 ( 
.A(n_707),
.B(n_758),
.Y(n_948)
);

INVx5_ASAP7_75t_L g949 ( 
.A(n_815),
.Y(n_949)
);

CKINVDCx10_ASAP7_75t_R g950 ( 
.A(n_790),
.Y(n_950)
);

AOI21xp5_ASAP7_75t_L g951 ( 
.A1(n_803),
.A2(n_603),
.B(n_586),
.Y(n_951)
);

INVx3_ASAP7_75t_L g952 ( 
.A(n_701),
.Y(n_952)
);

AOI21xp5_ASAP7_75t_L g953 ( 
.A1(n_808),
.A2(n_603),
.B(n_586),
.Y(n_953)
);

AND2x2_ASAP7_75t_L g954 ( 
.A(n_756),
.B(n_608),
.Y(n_954)
);

INVx1_ASAP7_75t_L g955 ( 
.A(n_835),
.Y(n_955)
);

AOI21xp5_ASAP7_75t_L g956 ( 
.A1(n_809),
.A2(n_603),
.B(n_586),
.Y(n_956)
);

O2A1O1Ixp33_ASAP7_75t_L g957 ( 
.A1(n_828),
.A2(n_611),
.B(n_609),
.C(n_617),
.Y(n_957)
);

AOI22xp5_ASAP7_75t_L g958 ( 
.A1(n_768),
.A2(n_772),
.B1(n_786),
.B2(n_777),
.Y(n_958)
);

O2A1O1Ixp33_ASAP7_75t_L g959 ( 
.A1(n_813),
.A2(n_617),
.B(n_622),
.C(n_611),
.Y(n_959)
);

AOI22xp5_ASAP7_75t_L g960 ( 
.A1(n_787),
.A2(n_608),
.B1(n_684),
.B2(n_649),
.Y(n_960)
);

AOI21xp5_ASAP7_75t_L g961 ( 
.A1(n_812),
.A2(n_559),
.B(n_616),
.Y(n_961)
);

OAI21xp5_ASAP7_75t_L g962 ( 
.A1(n_689),
.A2(n_559),
.B(n_616),
.Y(n_962)
);

NOR2xp33_ASAP7_75t_L g963 ( 
.A(n_852),
.B(n_608),
.Y(n_963)
);

NAND2xp5_ASAP7_75t_SL g964 ( 
.A(n_845),
.B(n_209),
.Y(n_964)
);

NOR2xp33_ASAP7_75t_L g965 ( 
.A(n_837),
.B(n_209),
.Y(n_965)
);

NAND2xp5_ASAP7_75t_L g966 ( 
.A(n_807),
.B(n_710),
.Y(n_966)
);

AOI21xp5_ASAP7_75t_L g967 ( 
.A1(n_689),
.A2(n_616),
.B(n_619),
.Y(n_967)
);

AND2x4_ASAP7_75t_L g968 ( 
.A(n_799),
.B(n_508),
.Y(n_968)
);

BUFx4f_ASAP7_75t_L g969 ( 
.A(n_744),
.Y(n_969)
);

NOR2xp33_ASAP7_75t_L g970 ( 
.A(n_813),
.B(n_210),
.Y(n_970)
);

O2A1O1Ixp33_ASAP7_75t_L g971 ( 
.A1(n_693),
.A2(n_622),
.B(n_508),
.C(n_519),
.Y(n_971)
);

O2A1O1Ixp5_ASAP7_75t_L g972 ( 
.A1(n_745),
.A2(n_619),
.B(n_636),
.C(n_625),
.Y(n_972)
);

BUFx6f_ASAP7_75t_L g973 ( 
.A(n_701),
.Y(n_973)
);

NAND2xp5_ASAP7_75t_SL g974 ( 
.A(n_722),
.B(n_210),
.Y(n_974)
);

BUFx6f_ASAP7_75t_L g975 ( 
.A(n_701),
.Y(n_975)
);

INVx3_ASAP7_75t_L g976 ( 
.A(n_725),
.Y(n_976)
);

NAND2xp5_ASAP7_75t_SL g977 ( 
.A(n_815),
.B(n_214),
.Y(n_977)
);

NOR2xp33_ASAP7_75t_L g978 ( 
.A(n_776),
.B(n_214),
.Y(n_978)
);

OAI21xp33_ASAP7_75t_L g979 ( 
.A1(n_820),
.A2(n_346),
.B(n_220),
.Y(n_979)
);

NAND2xp5_ASAP7_75t_L g980 ( 
.A(n_725),
.B(n_625),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_L g981 ( 
.A(n_727),
.B(n_625),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_L g982 ( 
.A(n_727),
.B(n_636),
.Y(n_982)
);

NAND2xp5_ASAP7_75t_SL g983 ( 
.A(n_815),
.B(n_215),
.Y(n_983)
);

INVx1_ASAP7_75t_L g984 ( 
.A(n_838),
.Y(n_984)
);

BUFx6f_ASAP7_75t_L g985 ( 
.A(n_799),
.Y(n_985)
);

OAI22xp33_ASAP7_75t_L g986 ( 
.A1(n_799),
.A2(n_229),
.B1(n_226),
.B2(n_221),
.Y(n_986)
);

NAND2xp5_ASAP7_75t_SL g987 ( 
.A(n_719),
.B(n_702),
.Y(n_987)
);

INVx2_ASAP7_75t_L g988 ( 
.A(n_732),
.Y(n_988)
);

NOR2xp33_ASAP7_75t_L g989 ( 
.A(n_818),
.B(n_215),
.Y(n_989)
);

CKINVDCx5p33_ASAP7_75t_R g990 ( 
.A(n_790),
.Y(n_990)
);

INVx2_ASAP7_75t_L g991 ( 
.A(n_732),
.Y(n_991)
);

AOI21xp5_ASAP7_75t_L g992 ( 
.A1(n_693),
.A2(n_728),
.B(n_720),
.Y(n_992)
);

NAND2xp5_ASAP7_75t_L g993 ( 
.A(n_733),
.B(n_636),
.Y(n_993)
);

INVx2_ASAP7_75t_L g994 ( 
.A(n_733),
.Y(n_994)
);

NAND2x1p5_ASAP7_75t_L g995 ( 
.A(n_833),
.B(n_644),
.Y(n_995)
);

AOI22xp5_ASAP7_75t_L g996 ( 
.A1(n_818),
.A2(n_684),
.B1(n_649),
.B2(n_294),
.Y(n_996)
);

OAI22xp5_ASAP7_75t_L g997 ( 
.A1(n_715),
.A2(n_226),
.B1(n_221),
.B2(n_229),
.Y(n_997)
);

AOI21xp5_ASAP7_75t_L g998 ( 
.A1(n_718),
.A2(n_765),
.B(n_764),
.Y(n_998)
);

NAND2xp5_ASAP7_75t_L g999 ( 
.A(n_738),
.B(n_649),
.Y(n_999)
);

O2A1O1Ixp33_ASAP7_75t_L g1000 ( 
.A1(n_719),
.A2(n_508),
.B(n_519),
.C(n_641),
.Y(n_1000)
);

NAND2xp5_ASAP7_75t_SL g1001 ( 
.A(n_826),
.B(n_304),
.Y(n_1001)
);

AOI21xp5_ASAP7_75t_L g1002 ( 
.A1(n_730),
.A2(n_635),
.B(n_637),
.Y(n_1002)
);

NAND2xp5_ASAP7_75t_SL g1003 ( 
.A(n_826),
.B(n_304),
.Y(n_1003)
);

NAND2xp5_ASAP7_75t_L g1004 ( 
.A(n_738),
.B(n_649),
.Y(n_1004)
);

OR2x6_ASAP7_75t_L g1005 ( 
.A(n_744),
.B(n_479),
.Y(n_1005)
);

AOI21xp5_ASAP7_75t_L g1006 ( 
.A1(n_834),
.A2(n_637),
.B(n_635),
.Y(n_1006)
);

AND2x4_ASAP7_75t_L g1007 ( 
.A(n_744),
.B(n_479),
.Y(n_1007)
);

NAND2xp5_ASAP7_75t_L g1008 ( 
.A(n_762),
.B(n_649),
.Y(n_1008)
);

INVx2_ASAP7_75t_SL g1009 ( 
.A(n_844),
.Y(n_1009)
);

OR2x2_ASAP7_75t_L g1010 ( 
.A(n_749),
.B(n_211),
.Y(n_1010)
);

NAND2xp5_ASAP7_75t_SL g1011 ( 
.A(n_827),
.B(n_307),
.Y(n_1011)
);

OAI21xp5_ASAP7_75t_L g1012 ( 
.A1(n_829),
.A2(n_641),
.B(n_545),
.Y(n_1012)
);

INVx2_ASAP7_75t_SL g1013 ( 
.A(n_851),
.Y(n_1013)
);

NAND2xp5_ASAP7_75t_L g1014 ( 
.A(n_762),
.B(n_684),
.Y(n_1014)
);

HB1xp67_ASAP7_75t_L g1015 ( 
.A(n_827),
.Y(n_1015)
);

BUFx12f_ASAP7_75t_L g1016 ( 
.A(n_850),
.Y(n_1016)
);

OAI21xp5_ASAP7_75t_L g1017 ( 
.A1(n_825),
.A2(n_550),
.B(n_545),
.Y(n_1017)
);

OAI22xp5_ASAP7_75t_L g1018 ( 
.A1(n_715),
.A2(n_745),
.B1(n_797),
.B2(n_752),
.Y(n_1018)
);

AOI21xp5_ASAP7_75t_L g1019 ( 
.A1(n_766),
.A2(n_550),
.B(n_562),
.Y(n_1019)
);

AOI21xp5_ASAP7_75t_L g1020 ( 
.A1(n_821),
.A2(n_561),
.B(n_644),
.Y(n_1020)
);

OAI22xp5_ASAP7_75t_L g1021 ( 
.A1(n_716),
.A2(n_365),
.B1(n_352),
.B2(n_340),
.Y(n_1021)
);

NOR2xp33_ASAP7_75t_L g1022 ( 
.A(n_855),
.B(n_307),
.Y(n_1022)
);

A2O1A1Ixp33_ASAP7_75t_L g1023 ( 
.A1(n_850),
.A2(n_322),
.B(n_351),
.C(n_352),
.Y(n_1023)
);

AOI21xp33_ASAP7_75t_L g1024 ( 
.A1(n_767),
.A2(n_334),
.B(n_361),
.Y(n_1024)
);

OAI21xp5_ASAP7_75t_L g1025 ( 
.A1(n_717),
.A2(n_684),
.B(n_465),
.Y(n_1025)
);

OAI21xp5_ASAP7_75t_L g1026 ( 
.A1(n_823),
.A2(n_684),
.B(n_465),
.Y(n_1026)
);

AOI21xp5_ASAP7_75t_L g1027 ( 
.A1(n_767),
.A2(n_644),
.B(n_463),
.Y(n_1027)
);

O2A1O1Ixp33_ASAP7_75t_L g1028 ( 
.A1(n_781),
.A2(n_484),
.B(n_481),
.C(n_459),
.Y(n_1028)
);

NOR2xp33_ASAP7_75t_L g1029 ( 
.A(n_851),
.B(n_316),
.Y(n_1029)
);

INVxp67_ASAP7_75t_L g1030 ( 
.A(n_855),
.Y(n_1030)
);

NAND2xp5_ASAP7_75t_L g1031 ( 
.A(n_775),
.B(n_684),
.Y(n_1031)
);

OAI21xp5_ASAP7_75t_L g1032 ( 
.A1(n_775),
.A2(n_459),
.B(n_467),
.Y(n_1032)
);

NAND2xp5_ASAP7_75t_L g1033 ( 
.A(n_778),
.B(n_283),
.Y(n_1033)
);

AOI21xp5_ASAP7_75t_L g1034 ( 
.A1(n_781),
.A2(n_463),
.B(n_467),
.Y(n_1034)
);

INVx2_ASAP7_75t_L g1035 ( 
.A(n_778),
.Y(n_1035)
);

AO21x2_ASAP7_75t_L g1036 ( 
.A1(n_792),
.A2(n_484),
.B(n_481),
.Y(n_1036)
);

NAND2xp5_ASAP7_75t_L g1037 ( 
.A(n_798),
.B(n_854),
.Y(n_1037)
);

O2A1O1Ixp5_ASAP7_75t_L g1038 ( 
.A1(n_792),
.A2(n_481),
.B(n_467),
.C(n_353),
.Y(n_1038)
);

O2A1O1Ixp5_ASAP7_75t_L g1039 ( 
.A1(n_805),
.A2(n_847),
.B(n_843),
.C(n_833),
.Y(n_1039)
);

AOI21xp5_ASAP7_75t_L g1040 ( 
.A1(n_805),
.A2(n_463),
.B(n_467),
.Y(n_1040)
);

INVx3_ASAP7_75t_L g1041 ( 
.A(n_930),
.Y(n_1041)
);

NOR3xp33_ASAP7_75t_SL g1042 ( 
.A(n_902),
.B(n_343),
.C(n_305),
.Y(n_1042)
);

A2O1A1Ixp33_ASAP7_75t_L g1043 ( 
.A1(n_880),
.A2(n_692),
.B(n_748),
.C(n_757),
.Y(n_1043)
);

INVx1_ASAP7_75t_L g1044 ( 
.A(n_872),
.Y(n_1044)
);

A2O1A1Ixp33_ASAP7_75t_L g1045 ( 
.A1(n_864),
.A2(n_692),
.B(n_748),
.C(n_757),
.Y(n_1045)
);

NAND2xp5_ASAP7_75t_SL g1046 ( 
.A(n_877),
.B(n_814),
.Y(n_1046)
);

NAND2xp5_ASAP7_75t_L g1047 ( 
.A(n_871),
.B(n_832),
.Y(n_1047)
);

NOR2xp33_ASAP7_75t_L g1048 ( 
.A(n_858),
.B(n_836),
.Y(n_1048)
);

O2A1O1Ixp33_ASAP7_75t_L g1049 ( 
.A1(n_936),
.A2(n_849),
.B(n_846),
.C(n_842),
.Y(n_1049)
);

AND2x4_ASAP7_75t_L g1050 ( 
.A(n_985),
.B(n_832),
.Y(n_1050)
);

NAND2xp5_ASAP7_75t_L g1051 ( 
.A(n_859),
.B(n_841),
.Y(n_1051)
);

O2A1O1Ixp33_ASAP7_75t_L g1052 ( 
.A1(n_884),
.A2(n_840),
.B(n_839),
.C(n_847),
.Y(n_1052)
);

OAI22xp5_ASAP7_75t_L g1053 ( 
.A1(n_1018),
.A2(n_841),
.B1(n_843),
.B2(n_275),
.Y(n_1053)
);

NAND2xp5_ASAP7_75t_L g1054 ( 
.A(n_1030),
.B(n_316),
.Y(n_1054)
);

BUFx3_ASAP7_75t_L g1055 ( 
.A(n_923),
.Y(n_1055)
);

NOR3xp33_ASAP7_75t_L g1056 ( 
.A(n_978),
.B(n_334),
.C(n_305),
.Y(n_1056)
);

OAI22xp5_ASAP7_75t_L g1057 ( 
.A1(n_969),
.A2(n_275),
.B1(n_312),
.B2(n_320),
.Y(n_1057)
);

OAI21xp5_ASAP7_75t_L g1058 ( 
.A1(n_992),
.A2(n_467),
.B(n_286),
.Y(n_1058)
);

HB1xp67_ASAP7_75t_L g1059 ( 
.A(n_889),
.Y(n_1059)
);

AOI21xp5_ASAP7_75t_L g1060 ( 
.A1(n_949),
.A2(n_463),
.B(n_290),
.Y(n_1060)
);

NAND2xp5_ASAP7_75t_L g1061 ( 
.A(n_1015),
.B(n_365),
.Y(n_1061)
);

INVx1_ASAP7_75t_SL g1062 ( 
.A(n_896),
.Y(n_1062)
);

A2O1A1Ixp33_ASAP7_75t_L g1063 ( 
.A1(n_941),
.A2(n_989),
.B(n_970),
.C(n_892),
.Y(n_1063)
);

OAI22xp5_ASAP7_75t_L g1064 ( 
.A1(n_969),
.A2(n_312),
.B1(n_359),
.B2(n_357),
.Y(n_1064)
);

A2O1A1Ixp33_ASAP7_75t_L g1065 ( 
.A1(n_887),
.A2(n_360),
.B(n_318),
.C(n_356),
.Y(n_1065)
);

AND2x2_ASAP7_75t_L g1066 ( 
.A(n_946),
.B(n_353),
.Y(n_1066)
);

NOR2xp33_ASAP7_75t_L g1067 ( 
.A(n_944),
.B(n_965),
.Y(n_1067)
);

CKINVDCx8_ASAP7_75t_R g1068 ( 
.A(n_950),
.Y(n_1068)
);

AOI21xp5_ASAP7_75t_L g1069 ( 
.A1(n_949),
.A2(n_360),
.B(n_356),
.Y(n_1069)
);

OAI22xp5_ASAP7_75t_L g1070 ( 
.A1(n_906),
.A2(n_357),
.B1(n_331),
.B2(n_346),
.Y(n_1070)
);

OR2x2_ASAP7_75t_L g1071 ( 
.A(n_931),
.B(n_320),
.Y(n_1071)
);

AOI21xp5_ASAP7_75t_L g1072 ( 
.A1(n_949),
.A2(n_351),
.B(n_318),
.Y(n_1072)
);

CKINVDCx8_ASAP7_75t_R g1073 ( 
.A(n_898),
.Y(n_1073)
);

AOI21xp5_ASAP7_75t_L g1074 ( 
.A1(n_949),
.A2(n_321),
.B(n_322),
.Y(n_1074)
);

AND2x2_ASAP7_75t_L g1075 ( 
.A(n_891),
.B(n_344),
.Y(n_1075)
);

CKINVDCx5p33_ASAP7_75t_R g1076 ( 
.A(n_924),
.Y(n_1076)
);

NAND2xp5_ASAP7_75t_L g1077 ( 
.A(n_882),
.B(n_321),
.Y(n_1077)
);

NAND2xp5_ASAP7_75t_SL g1078 ( 
.A(n_901),
.B(n_926),
.Y(n_1078)
);

AOI21xp5_ASAP7_75t_L g1079 ( 
.A1(n_879),
.A2(n_325),
.B(n_330),
.Y(n_1079)
);

NOR2xp33_ASAP7_75t_L g1080 ( 
.A(n_915),
.B(n_344),
.Y(n_1080)
);

NOR2xp67_ASAP7_75t_SL g1081 ( 
.A(n_973),
.B(n_340),
.Y(n_1081)
);

NAND2xp5_ASAP7_75t_L g1082 ( 
.A(n_875),
.B(n_338),
.Y(n_1082)
);

OR2x2_ASAP7_75t_L g1083 ( 
.A(n_1010),
.B(n_343),
.Y(n_1083)
);

BUFx6f_ASAP7_75t_L g1084 ( 
.A(n_985),
.Y(n_1084)
);

NAND2xp5_ASAP7_75t_SL g1085 ( 
.A(n_901),
.B(n_338),
.Y(n_1085)
);

INVx2_ASAP7_75t_L g1086 ( 
.A(n_976),
.Y(n_1086)
);

INVx2_ASAP7_75t_SL g1087 ( 
.A(n_1009),
.Y(n_1087)
);

NAND3xp33_ASAP7_75t_SL g1088 ( 
.A(n_954),
.B(n_331),
.C(n_330),
.Y(n_1088)
);

NOR2xp33_ASAP7_75t_L g1089 ( 
.A(n_938),
.B(n_325),
.Y(n_1089)
);

BUFx3_ASAP7_75t_L g1090 ( 
.A(n_990),
.Y(n_1090)
);

NOR2xp67_ASAP7_75t_L g1091 ( 
.A(n_1013),
.B(n_181),
.Y(n_1091)
);

AND2x2_ASAP7_75t_L g1092 ( 
.A(n_1007),
.B(n_11),
.Y(n_1092)
);

NAND2xp5_ASAP7_75t_L g1093 ( 
.A(n_875),
.B(n_171),
.Y(n_1093)
);

INVx1_ASAP7_75t_L g1094 ( 
.A(n_878),
.Y(n_1094)
);

INVx3_ASAP7_75t_L g1095 ( 
.A(n_930),
.Y(n_1095)
);

NAND2x1p5_ASAP7_75t_L g1096 ( 
.A(n_973),
.B(n_161),
.Y(n_1096)
);

NAND2xp5_ASAP7_75t_SL g1097 ( 
.A(n_901),
.B(n_154),
.Y(n_1097)
);

INVx2_ASAP7_75t_SL g1098 ( 
.A(n_968),
.Y(n_1098)
);

AOI21xp5_ASAP7_75t_L g1099 ( 
.A1(n_992),
.A2(n_147),
.B(n_145),
.Y(n_1099)
);

NAND2xp5_ASAP7_75t_SL g1100 ( 
.A(n_912),
.B(n_143),
.Y(n_1100)
);

NAND2xp5_ASAP7_75t_SL g1101 ( 
.A(n_894),
.B(n_133),
.Y(n_1101)
);

CKINVDCx5p33_ASAP7_75t_R g1102 ( 
.A(n_1016),
.Y(n_1102)
);

O2A1O1Ixp33_ASAP7_75t_L g1103 ( 
.A1(n_1023),
.A2(n_13),
.B(n_14),
.C(n_15),
.Y(n_1103)
);

OAI22xp5_ASAP7_75t_L g1104 ( 
.A1(n_916),
.A2(n_13),
.B1(n_16),
.B2(n_17),
.Y(n_1104)
);

NOR2xp33_ASAP7_75t_L g1105 ( 
.A(n_964),
.B(n_16),
.Y(n_1105)
);

BUFx2_ASAP7_75t_SL g1106 ( 
.A(n_985),
.Y(n_1106)
);

INVx1_ASAP7_75t_L g1107 ( 
.A(n_897),
.Y(n_1107)
);

NAND2xp5_ASAP7_75t_L g1108 ( 
.A(n_885),
.B(n_919),
.Y(n_1108)
);

A2O1A1Ixp33_ASAP7_75t_L g1109 ( 
.A1(n_1022),
.A2(n_18),
.B(n_19),
.C(n_20),
.Y(n_1109)
);

NAND2xp5_ASAP7_75t_L g1110 ( 
.A(n_860),
.B(n_18),
.Y(n_1110)
);

NOR2xp33_ASAP7_75t_L g1111 ( 
.A(n_899),
.B(n_20),
.Y(n_1111)
);

NAND2xp5_ASAP7_75t_SL g1112 ( 
.A(n_973),
.B(n_131),
.Y(n_1112)
);

OAI22xp5_ASAP7_75t_L g1113 ( 
.A1(n_917),
.A2(n_22),
.B1(n_23),
.B2(n_24),
.Y(n_1113)
);

AOI21xp5_ASAP7_75t_L g1114 ( 
.A1(n_998),
.A2(n_129),
.B(n_109),
.Y(n_1114)
);

INVx3_ASAP7_75t_SL g1115 ( 
.A(n_1005),
.Y(n_1115)
);

BUFx6f_ASAP7_75t_L g1116 ( 
.A(n_1005),
.Y(n_1116)
);

AOI21xp5_ASAP7_75t_L g1117 ( 
.A1(n_998),
.A2(n_88),
.B(n_85),
.Y(n_1117)
);

INVx2_ASAP7_75t_SL g1118 ( 
.A(n_968),
.Y(n_1118)
);

BUFx6f_ASAP7_75t_L g1119 ( 
.A(n_975),
.Y(n_1119)
);

AOI21xp5_ASAP7_75t_L g1120 ( 
.A1(n_869),
.A2(n_78),
.B(n_76),
.Y(n_1120)
);

O2A1O1Ixp33_ASAP7_75t_L g1121 ( 
.A1(n_1024),
.A2(n_24),
.B(n_26),
.C(n_27),
.Y(n_1121)
);

AND2x4_ASAP7_75t_L g1122 ( 
.A(n_1007),
.B(n_26),
.Y(n_1122)
);

O2A1O1Ixp33_ASAP7_75t_L g1123 ( 
.A1(n_943),
.A2(n_27),
.B(n_30),
.C(n_31),
.Y(n_1123)
);

OAI22xp5_ASAP7_75t_L g1124 ( 
.A1(n_920),
.A2(n_33),
.B1(n_35),
.B2(n_36),
.Y(n_1124)
);

INVxp67_ASAP7_75t_L g1125 ( 
.A(n_963),
.Y(n_1125)
);

NOR2xp33_ASAP7_75t_L g1126 ( 
.A(n_979),
.B(n_33),
.Y(n_1126)
);

AOI21xp5_ASAP7_75t_L g1127 ( 
.A1(n_869),
.A2(n_63),
.B(n_40),
.Y(n_1127)
);

NAND2xp5_ASAP7_75t_L g1128 ( 
.A(n_885),
.B(n_39),
.Y(n_1128)
);

AOI21xp5_ASAP7_75t_L g1129 ( 
.A1(n_886),
.A2(n_890),
.B(n_947),
.Y(n_1129)
);

NOR2xp33_ASAP7_75t_L g1130 ( 
.A(n_1029),
.B(n_42),
.Y(n_1130)
);

INVx1_ASAP7_75t_L g1131 ( 
.A(n_903),
.Y(n_1131)
);

BUFx3_ASAP7_75t_L g1132 ( 
.A(n_948),
.Y(n_1132)
);

O2A1O1Ixp33_ASAP7_75t_L g1133 ( 
.A1(n_997),
.A2(n_46),
.B(n_49),
.C(n_53),
.Y(n_1133)
);

INVx1_ASAP7_75t_L g1134 ( 
.A(n_913),
.Y(n_1134)
);

AOI21xp5_ASAP7_75t_L g1135 ( 
.A1(n_1025),
.A2(n_62),
.B(n_55),
.Y(n_1135)
);

INVx1_ASAP7_75t_L g1136 ( 
.A(n_937),
.Y(n_1136)
);

AND2x4_ASAP7_75t_L g1137 ( 
.A(n_893),
.B(n_49),
.Y(n_1137)
);

AND2x2_ASAP7_75t_L g1138 ( 
.A(n_909),
.B(n_56),
.Y(n_1138)
);

INVx1_ASAP7_75t_L g1139 ( 
.A(n_988),
.Y(n_1139)
);

AOI21xp5_ASAP7_75t_L g1140 ( 
.A1(n_863),
.A2(n_59),
.B(n_60),
.Y(n_1140)
);

INVx1_ASAP7_75t_L g1141 ( 
.A(n_991),
.Y(n_1141)
);

AOI21xp5_ASAP7_75t_L g1142 ( 
.A1(n_863),
.A2(n_61),
.B(n_866),
.Y(n_1142)
);

INVx3_ASAP7_75t_L g1143 ( 
.A(n_930),
.Y(n_1143)
);

BUFx6f_ASAP7_75t_L g1144 ( 
.A(n_975),
.Y(n_1144)
);

AOI22xp5_ASAP7_75t_L g1145 ( 
.A1(n_987),
.A2(n_61),
.B1(n_1001),
.B2(n_1003),
.Y(n_1145)
);

INVx1_ASAP7_75t_L g1146 ( 
.A(n_994),
.Y(n_1146)
);

HAxp5_ASAP7_75t_L g1147 ( 
.A(n_907),
.B(n_974),
.CON(n_1147),
.SN(n_1147)
);

AOI21xp5_ASAP7_75t_L g1148 ( 
.A1(n_866),
.A2(n_867),
.B(n_904),
.Y(n_1148)
);

INVx1_ASAP7_75t_L g1149 ( 
.A(n_1035),
.Y(n_1149)
);

OR2x2_ASAP7_75t_L g1150 ( 
.A(n_914),
.B(n_1021),
.Y(n_1150)
);

NOR2xp33_ASAP7_75t_R g1151 ( 
.A(n_975),
.B(n_952),
.Y(n_1151)
);

AOI21xp5_ASAP7_75t_L g1152 ( 
.A1(n_867),
.A2(n_922),
.B(n_910),
.Y(n_1152)
);

NAND2xp5_ASAP7_75t_L g1153 ( 
.A(n_919),
.B(n_921),
.Y(n_1153)
);

O2A1O1Ixp33_ASAP7_75t_L g1154 ( 
.A1(n_1011),
.A2(n_925),
.B(n_986),
.C(n_918),
.Y(n_1154)
);

AOI21xp5_ASAP7_75t_L g1155 ( 
.A1(n_908),
.A2(n_945),
.B(n_942),
.Y(n_1155)
);

INVx2_ASAP7_75t_L g1156 ( 
.A(n_976),
.Y(n_1156)
);

OAI22xp5_ASAP7_75t_L g1157 ( 
.A1(n_881),
.A2(n_900),
.B1(n_939),
.B2(n_911),
.Y(n_1157)
);

INVx1_ASAP7_75t_L g1158 ( 
.A(n_966),
.Y(n_1158)
);

NOR2xp67_ASAP7_75t_L g1159 ( 
.A(n_955),
.B(n_984),
.Y(n_1159)
);

NOR2xp33_ASAP7_75t_L g1160 ( 
.A(n_948),
.B(n_883),
.Y(n_1160)
);

AOI21xp5_ASAP7_75t_L g1161 ( 
.A1(n_935),
.A2(n_895),
.B(n_929),
.Y(n_1161)
);

NOR2xp33_ASAP7_75t_L g1162 ( 
.A(n_876),
.B(n_958),
.Y(n_1162)
);

INVx1_ASAP7_75t_L g1163 ( 
.A(n_1037),
.Y(n_1163)
);

NAND2xp5_ASAP7_75t_L g1164 ( 
.A(n_1033),
.B(n_868),
.Y(n_1164)
);

AOI22xp5_ASAP7_75t_L g1165 ( 
.A1(n_905),
.A2(n_888),
.B1(n_977),
.B2(n_983),
.Y(n_1165)
);

AOI21xp5_ASAP7_75t_L g1166 ( 
.A1(n_927),
.A2(n_856),
.B(n_928),
.Y(n_1166)
);

INVx3_ASAP7_75t_L g1167 ( 
.A(n_995),
.Y(n_1167)
);

AOI21xp5_ASAP7_75t_L g1168 ( 
.A1(n_856),
.A2(n_962),
.B(n_951),
.Y(n_1168)
);

INVx4_ASAP7_75t_L g1169 ( 
.A(n_995),
.Y(n_1169)
);

AOI22xp33_ASAP7_75t_L g1170 ( 
.A1(n_1036),
.A2(n_861),
.B1(n_862),
.B2(n_865),
.Y(n_1170)
);

AOI21xp5_ASAP7_75t_L g1171 ( 
.A1(n_951),
.A2(n_961),
.B(n_953),
.Y(n_1171)
);

INVx1_ASAP7_75t_L g1172 ( 
.A(n_957),
.Y(n_1172)
);

AOI21xp5_ASAP7_75t_L g1173 ( 
.A1(n_953),
.A2(n_956),
.B(n_961),
.Y(n_1173)
);

INVx1_ASAP7_75t_SL g1174 ( 
.A(n_1036),
.Y(n_1174)
);

INVx2_ASAP7_75t_L g1175 ( 
.A(n_980),
.Y(n_1175)
);

NOR2xp67_ASAP7_75t_L g1176 ( 
.A(n_933),
.B(n_960),
.Y(n_1176)
);

INVx1_ASAP7_75t_L g1177 ( 
.A(n_971),
.Y(n_1177)
);

NOR2xp33_ASAP7_75t_L g1178 ( 
.A(n_981),
.B(n_982),
.Y(n_1178)
);

AOI22xp5_ASAP7_75t_L g1179 ( 
.A1(n_996),
.A2(n_1004),
.B1(n_1014),
.B2(n_1031),
.Y(n_1179)
);

INVx3_ASAP7_75t_SL g1180 ( 
.A(n_1038),
.Y(n_1180)
);

A2O1A1Ixp33_ASAP7_75t_L g1181 ( 
.A1(n_1039),
.A2(n_870),
.B(n_873),
.C(n_874),
.Y(n_1181)
);

NOR2xp33_ASAP7_75t_L g1182 ( 
.A(n_993),
.B(n_999),
.Y(n_1182)
);

INVx4_ASAP7_75t_L g1183 ( 
.A(n_870),
.Y(n_1183)
);

AND2x2_ASAP7_75t_L g1184 ( 
.A(n_873),
.B(n_874),
.Y(n_1184)
);

AOI21xp5_ASAP7_75t_L g1185 ( 
.A1(n_956),
.A2(n_967),
.B(n_940),
.Y(n_1185)
);

AOI21xp5_ASAP7_75t_L g1186 ( 
.A1(n_967),
.A2(n_932),
.B(n_1017),
.Y(n_1186)
);

BUFx6f_ASAP7_75t_L g1187 ( 
.A(n_857),
.Y(n_1187)
);

A2O1A1Ixp33_ASAP7_75t_L g1188 ( 
.A1(n_972),
.A2(n_959),
.B(n_1000),
.C(n_934),
.Y(n_1188)
);

NOR2xp33_ASAP7_75t_L g1189 ( 
.A(n_1008),
.B(n_1020),
.Y(n_1189)
);

O2A1O1Ixp5_ASAP7_75t_L g1190 ( 
.A1(n_1020),
.A2(n_1006),
.B(n_1012),
.C(n_1026),
.Y(n_1190)
);

INVx2_ASAP7_75t_L g1191 ( 
.A(n_1032),
.Y(n_1191)
);

AND2x2_ASAP7_75t_L g1192 ( 
.A(n_1006),
.B(n_1002),
.Y(n_1192)
);

NOR2xp67_ASAP7_75t_SL g1193 ( 
.A(n_1027),
.B(n_1019),
.Y(n_1193)
);

NOR2xp33_ASAP7_75t_L g1194 ( 
.A(n_1028),
.B(n_1027),
.Y(n_1194)
);

OAI21xp5_ASAP7_75t_L g1195 ( 
.A1(n_1063),
.A2(n_1034),
.B(n_1040),
.Y(n_1195)
);

AND2x4_ASAP7_75t_L g1196 ( 
.A(n_1132),
.B(n_1034),
.Y(n_1196)
);

AO31x2_ASAP7_75t_L g1197 ( 
.A1(n_1148),
.A2(n_1040),
.A3(n_1168),
.B(n_1181),
.Y(n_1197)
);

AOI21xp5_ASAP7_75t_L g1198 ( 
.A1(n_1161),
.A2(n_1155),
.B(n_1164),
.Y(n_1198)
);

BUFx6f_ASAP7_75t_L g1199 ( 
.A(n_1084),
.Y(n_1199)
);

O2A1O1Ixp33_ASAP7_75t_L g1200 ( 
.A1(n_1130),
.A2(n_1067),
.B(n_1109),
.C(n_1147),
.Y(n_1200)
);

OA21x2_ASAP7_75t_L g1201 ( 
.A1(n_1142),
.A2(n_1190),
.B(n_1173),
.Y(n_1201)
);

NOR2xp67_ASAP7_75t_L g1202 ( 
.A(n_1082),
.B(n_1165),
.Y(n_1202)
);

OAI22xp5_ASAP7_75t_L g1203 ( 
.A1(n_1150),
.A2(n_1062),
.B1(n_1176),
.B2(n_1125),
.Y(n_1203)
);

NAND2xp5_ASAP7_75t_L g1204 ( 
.A(n_1158),
.B(n_1163),
.Y(n_1204)
);

NAND2xp5_ASAP7_75t_L g1205 ( 
.A(n_1048),
.B(n_1075),
.Y(n_1205)
);

OA21x2_ASAP7_75t_L g1206 ( 
.A1(n_1171),
.A2(n_1186),
.B(n_1185),
.Y(n_1206)
);

INVx1_ASAP7_75t_SL g1207 ( 
.A(n_1062),
.Y(n_1207)
);

AO31x2_ASAP7_75t_L g1208 ( 
.A1(n_1157),
.A2(n_1188),
.A3(n_1152),
.B(n_1194),
.Y(n_1208)
);

OR2x6_ASAP7_75t_L g1209 ( 
.A(n_1106),
.B(n_1116),
.Y(n_1209)
);

O2A1O1Ixp5_ASAP7_75t_L g1210 ( 
.A1(n_1135),
.A2(n_1089),
.B(n_1127),
.C(n_1078),
.Y(n_1210)
);

OAI21x1_ASAP7_75t_L g1211 ( 
.A1(n_1129),
.A2(n_1093),
.B(n_1192),
.Y(n_1211)
);

NAND2xp5_ASAP7_75t_L g1212 ( 
.A(n_1080),
.B(n_1047),
.Y(n_1212)
);

OAI21x1_ASAP7_75t_L g1213 ( 
.A1(n_1093),
.A2(n_1120),
.B(n_1099),
.Y(n_1213)
);

NAND2xp5_ASAP7_75t_L g1214 ( 
.A(n_1047),
.B(n_1160),
.Y(n_1214)
);

NAND2xp5_ASAP7_75t_L g1215 ( 
.A(n_1162),
.B(n_1138),
.Y(n_1215)
);

A2O1A1Ixp33_ASAP7_75t_L g1216 ( 
.A1(n_1154),
.A2(n_1145),
.B(n_1045),
.C(n_1126),
.Y(n_1216)
);

AOI21xp5_ASAP7_75t_L g1217 ( 
.A1(n_1051),
.A2(n_1157),
.B(n_1178),
.Y(n_1217)
);

AOI21xp5_ASAP7_75t_L g1218 ( 
.A1(n_1051),
.A2(n_1052),
.B(n_1189),
.Y(n_1218)
);

AOI21xp5_ASAP7_75t_L g1219 ( 
.A1(n_1182),
.A2(n_1046),
.B(n_1184),
.Y(n_1219)
);

BUFx10_ASAP7_75t_L g1220 ( 
.A(n_1105),
.Y(n_1220)
);

OAI21x1_ASAP7_75t_L g1221 ( 
.A1(n_1114),
.A2(n_1117),
.B(n_1170),
.Y(n_1221)
);

OA21x2_ASAP7_75t_L g1222 ( 
.A1(n_1058),
.A2(n_1174),
.B(n_1177),
.Y(n_1222)
);

OAI21xp5_ASAP7_75t_L g1223 ( 
.A1(n_1043),
.A2(n_1053),
.B(n_1179),
.Y(n_1223)
);

AND2x4_ASAP7_75t_L g1224 ( 
.A(n_1098),
.B(n_1118),
.Y(n_1224)
);

O2A1O1Ixp5_ASAP7_75t_L g1225 ( 
.A1(n_1100),
.A2(n_1053),
.B(n_1081),
.C(n_1110),
.Y(n_1225)
);

OAI22xp5_ASAP7_75t_L g1226 ( 
.A1(n_1159),
.A2(n_1082),
.B1(n_1183),
.B2(n_1054),
.Y(n_1226)
);

NOR2xp33_ASAP7_75t_L g1227 ( 
.A(n_1066),
.B(n_1088),
.Y(n_1227)
);

NAND2xp5_ASAP7_75t_L g1228 ( 
.A(n_1175),
.B(n_1061),
.Y(n_1228)
);

A2O1A1Ixp33_ASAP7_75t_L g1229 ( 
.A1(n_1111),
.A2(n_1065),
.B(n_1140),
.C(n_1133),
.Y(n_1229)
);

NAND2xp5_ASAP7_75t_SL g1230 ( 
.A(n_1056),
.B(n_1042),
.Y(n_1230)
);

OAI21xp5_ASAP7_75t_L g1231 ( 
.A1(n_1049),
.A2(n_1058),
.B(n_1128),
.Y(n_1231)
);

AOI21xp5_ASAP7_75t_L g1232 ( 
.A1(n_1183),
.A2(n_1187),
.B(n_1191),
.Y(n_1232)
);

INVx1_ASAP7_75t_L g1233 ( 
.A(n_1094),
.Y(n_1233)
);

INVx1_ASAP7_75t_L g1234 ( 
.A(n_1107),
.Y(n_1234)
);

NAND2xp5_ASAP7_75t_L g1235 ( 
.A(n_1077),
.B(n_1092),
.Y(n_1235)
);

INVx3_ASAP7_75t_L g1236 ( 
.A(n_1119),
.Y(n_1236)
);

NOR2xp33_ASAP7_75t_L g1237 ( 
.A(n_1083),
.B(n_1071),
.Y(n_1237)
);

AOI21xp5_ASAP7_75t_L g1238 ( 
.A1(n_1187),
.A2(n_1172),
.B(n_1108),
.Y(n_1238)
);

AOI21x1_ASAP7_75t_L g1239 ( 
.A1(n_1128),
.A2(n_1101),
.B(n_1060),
.Y(n_1239)
);

BUFx12f_ASAP7_75t_L g1240 ( 
.A(n_1076),
.Y(n_1240)
);

BUFx6f_ASAP7_75t_L g1241 ( 
.A(n_1084),
.Y(n_1241)
);

NAND2xp5_ASAP7_75t_L g1242 ( 
.A(n_1122),
.B(n_1050),
.Y(n_1242)
);

INVx1_ASAP7_75t_L g1243 ( 
.A(n_1131),
.Y(n_1243)
);

INVxp67_ASAP7_75t_L g1244 ( 
.A(n_1059),
.Y(n_1244)
);

O2A1O1Ixp33_ASAP7_75t_SL g1245 ( 
.A1(n_1112),
.A2(n_1097),
.B(n_1153),
.C(n_1174),
.Y(n_1245)
);

O2A1O1Ixp33_ASAP7_75t_L g1246 ( 
.A1(n_1121),
.A2(n_1070),
.B(n_1124),
.C(n_1113),
.Y(n_1246)
);

AOI21xp5_ASAP7_75t_SL g1247 ( 
.A1(n_1096),
.A2(n_1187),
.B(n_1119),
.Y(n_1247)
);

A2O1A1Ixp33_ASAP7_75t_L g1248 ( 
.A1(n_1123),
.A2(n_1103),
.B(n_1091),
.C(n_1079),
.Y(n_1248)
);

INVx1_ASAP7_75t_L g1249 ( 
.A(n_1134),
.Y(n_1249)
);

INVx4_ASAP7_75t_L g1250 ( 
.A(n_1119),
.Y(n_1250)
);

INVx1_ASAP7_75t_L g1251 ( 
.A(n_1136),
.Y(n_1251)
);

AO31x2_ASAP7_75t_L g1252 ( 
.A1(n_1104),
.A2(n_1124),
.A3(n_1113),
.B(n_1070),
.Y(n_1252)
);

INVx3_ASAP7_75t_L g1253 ( 
.A(n_1144),
.Y(n_1253)
);

CKINVDCx12_ASAP7_75t_R g1254 ( 
.A(n_1073),
.Y(n_1254)
);

AO31x2_ASAP7_75t_L g1255 ( 
.A1(n_1104),
.A2(n_1169),
.A3(n_1141),
.B(n_1139),
.Y(n_1255)
);

A2O1A1Ixp33_ASAP7_75t_L g1256 ( 
.A1(n_1085),
.A2(n_1146),
.B(n_1149),
.C(n_1050),
.Y(n_1256)
);

AOI21xp5_ASAP7_75t_L g1257 ( 
.A1(n_1169),
.A2(n_1167),
.B(n_1156),
.Y(n_1257)
);

INVx1_ASAP7_75t_L g1258 ( 
.A(n_1086),
.Y(n_1258)
);

AOI21xp5_ASAP7_75t_L g1259 ( 
.A1(n_1167),
.A2(n_1041),
.B(n_1143),
.Y(n_1259)
);

INVxp67_ASAP7_75t_L g1260 ( 
.A(n_1087),
.Y(n_1260)
);

NAND2xp5_ASAP7_75t_L g1261 ( 
.A(n_1137),
.B(n_1116),
.Y(n_1261)
);

NAND2xp5_ASAP7_75t_SL g1262 ( 
.A(n_1137),
.B(n_1116),
.Y(n_1262)
);

OAI21xp5_ASAP7_75t_L g1263 ( 
.A1(n_1096),
.A2(n_1074),
.B(n_1072),
.Y(n_1263)
);

OAI22xp33_ASAP7_75t_L g1264 ( 
.A1(n_1115),
.A2(n_1102),
.B1(n_1057),
.B2(n_1064),
.Y(n_1264)
);

OAI21xp5_ASAP7_75t_L g1265 ( 
.A1(n_1069),
.A2(n_1041),
.B(n_1143),
.Y(n_1265)
);

AOI21xp5_ASAP7_75t_L g1266 ( 
.A1(n_1095),
.A2(n_1144),
.B(n_1180),
.Y(n_1266)
);

CKINVDCx16_ASAP7_75t_R g1267 ( 
.A(n_1055),
.Y(n_1267)
);

AND2x4_ASAP7_75t_L g1268 ( 
.A(n_1144),
.B(n_1095),
.Y(n_1268)
);

OAI21x1_ASAP7_75t_L g1269 ( 
.A1(n_1151),
.A2(n_1057),
.B(n_1064),
.Y(n_1269)
);

A2O1A1Ixp33_ASAP7_75t_L g1270 ( 
.A1(n_1090),
.A2(n_864),
.B(n_880),
.C(n_1063),
.Y(n_1270)
);

AOI21xp5_ASAP7_75t_L g1271 ( 
.A1(n_1068),
.A2(n_949),
.B(n_1063),
.Y(n_1271)
);

OAI21x1_ASAP7_75t_L g1272 ( 
.A1(n_1166),
.A2(n_1152),
.B(n_1171),
.Y(n_1272)
);

INVx4_ASAP7_75t_L g1273 ( 
.A(n_1084),
.Y(n_1273)
);

AND2x6_ASAP7_75t_L g1274 ( 
.A(n_1119),
.B(n_973),
.Y(n_1274)
);

NAND2xp5_ASAP7_75t_L g1275 ( 
.A(n_1067),
.B(n_864),
.Y(n_1275)
);

OAI21xp5_ASAP7_75t_L g1276 ( 
.A1(n_1063),
.A2(n_880),
.B(n_864),
.Y(n_1276)
);

OAI22xp5_ASAP7_75t_L g1277 ( 
.A1(n_1063),
.A2(n_864),
.B1(n_880),
.B2(n_1067),
.Y(n_1277)
);

AOI21xp5_ASAP7_75t_L g1278 ( 
.A1(n_1063),
.A2(n_949),
.B(n_1168),
.Y(n_1278)
);

BUFx6f_ASAP7_75t_L g1279 ( 
.A(n_1084),
.Y(n_1279)
);

AO31x2_ASAP7_75t_L g1280 ( 
.A1(n_1148),
.A2(n_1168),
.A3(n_1063),
.B(n_1181),
.Y(n_1280)
);

OAI21x1_ASAP7_75t_L g1281 ( 
.A1(n_1166),
.A2(n_1152),
.B(n_1171),
.Y(n_1281)
);

O2A1O1Ixp33_ASAP7_75t_SL g1282 ( 
.A1(n_1063),
.A2(n_880),
.B(n_719),
.C(n_1043),
.Y(n_1282)
);

AND2x2_ASAP7_75t_L g1283 ( 
.A(n_1075),
.B(n_877),
.Y(n_1283)
);

NAND2xp5_ASAP7_75t_L g1284 ( 
.A(n_1067),
.B(n_864),
.Y(n_1284)
);

CKINVDCx20_ASAP7_75t_R g1285 ( 
.A(n_1073),
.Y(n_1285)
);

O2A1O1Ixp33_ASAP7_75t_SL g1286 ( 
.A1(n_1063),
.A2(n_880),
.B(n_719),
.C(n_1043),
.Y(n_1286)
);

O2A1O1Ixp5_ASAP7_75t_L g1287 ( 
.A1(n_1130),
.A2(n_864),
.B(n_880),
.C(n_719),
.Y(n_1287)
);

AOI21x1_ASAP7_75t_L g1288 ( 
.A1(n_1193),
.A2(n_987),
.B(n_1168),
.Y(n_1288)
);

OA21x2_ASAP7_75t_L g1289 ( 
.A1(n_1148),
.A2(n_1168),
.B(n_1142),
.Y(n_1289)
);

NAND2xp5_ASAP7_75t_L g1290 ( 
.A(n_1067),
.B(n_864),
.Y(n_1290)
);

NOR2xp33_ASAP7_75t_L g1291 ( 
.A(n_1067),
.B(n_864),
.Y(n_1291)
);

A2O1A1Ixp33_ASAP7_75t_L g1292 ( 
.A1(n_1063),
.A2(n_864),
.B(n_880),
.C(n_1130),
.Y(n_1292)
);

OAI21x1_ASAP7_75t_L g1293 ( 
.A1(n_1166),
.A2(n_1152),
.B(n_1171),
.Y(n_1293)
);

AOI21xp5_ASAP7_75t_L g1294 ( 
.A1(n_1063),
.A2(n_949),
.B(n_1168),
.Y(n_1294)
);

NAND2x1p5_ASAP7_75t_L g1295 ( 
.A(n_1084),
.B(n_901),
.Y(n_1295)
);

A2O1A1Ixp33_ASAP7_75t_L g1296 ( 
.A1(n_1063),
.A2(n_864),
.B(n_880),
.C(n_1130),
.Y(n_1296)
);

AND2x2_ASAP7_75t_L g1297 ( 
.A(n_1075),
.B(n_877),
.Y(n_1297)
);

INVx2_ASAP7_75t_SL g1298 ( 
.A(n_1084),
.Y(n_1298)
);

AND2x2_ASAP7_75t_L g1299 ( 
.A(n_1075),
.B(n_877),
.Y(n_1299)
);

AOI221x1_ASAP7_75t_L g1300 ( 
.A1(n_1063),
.A2(n_880),
.B1(n_864),
.B2(n_1130),
.C(n_1135),
.Y(n_1300)
);

AOI21xp5_ASAP7_75t_L g1301 ( 
.A1(n_1063),
.A2(n_949),
.B(n_1168),
.Y(n_1301)
);

A2O1A1Ixp33_ASAP7_75t_L g1302 ( 
.A1(n_1063),
.A2(n_864),
.B(n_880),
.C(n_1130),
.Y(n_1302)
);

AO31x2_ASAP7_75t_L g1303 ( 
.A1(n_1148),
.A2(n_1168),
.A3(n_1063),
.B(n_1181),
.Y(n_1303)
);

INVx2_ASAP7_75t_L g1304 ( 
.A(n_1044),
.Y(n_1304)
);

NAND2xp5_ASAP7_75t_L g1305 ( 
.A(n_1067),
.B(n_864),
.Y(n_1305)
);

AOI22xp33_ASAP7_75t_L g1306 ( 
.A1(n_1130),
.A2(n_864),
.B1(n_1056),
.B2(n_811),
.Y(n_1306)
);

AO31x2_ASAP7_75t_L g1307 ( 
.A1(n_1148),
.A2(n_1168),
.A3(n_1063),
.B(n_1181),
.Y(n_1307)
);

INVx2_ASAP7_75t_L g1308 ( 
.A(n_1044),
.Y(n_1308)
);

BUFx6f_ASAP7_75t_L g1309 ( 
.A(n_1084),
.Y(n_1309)
);

AO31x2_ASAP7_75t_L g1310 ( 
.A1(n_1148),
.A2(n_1168),
.A3(n_1063),
.B(n_1181),
.Y(n_1310)
);

INVxp67_ASAP7_75t_L g1311 ( 
.A(n_1059),
.Y(n_1311)
);

NAND3xp33_ASAP7_75t_L g1312 ( 
.A(n_1130),
.B(n_864),
.C(n_880),
.Y(n_1312)
);

INVx3_ASAP7_75t_L g1313 ( 
.A(n_1119),
.Y(n_1313)
);

NAND3x1_ASAP7_75t_L g1314 ( 
.A(n_1130),
.B(n_864),
.C(n_691),
.Y(n_1314)
);

NOR2xp33_ASAP7_75t_L g1315 ( 
.A(n_1067),
.B(n_864),
.Y(n_1315)
);

AOI21xp5_ASAP7_75t_L g1316 ( 
.A1(n_1063),
.A2(n_949),
.B(n_1168),
.Y(n_1316)
);

OAI21x1_ASAP7_75t_L g1317 ( 
.A1(n_1166),
.A2(n_1152),
.B(n_1171),
.Y(n_1317)
);

OAI21xp5_ASAP7_75t_L g1318 ( 
.A1(n_1063),
.A2(n_880),
.B(n_1135),
.Y(n_1318)
);

OAI21x1_ASAP7_75t_L g1319 ( 
.A1(n_1166),
.A2(n_1152),
.B(n_1171),
.Y(n_1319)
);

BUFx3_ASAP7_75t_L g1320 ( 
.A(n_1084),
.Y(n_1320)
);

AO31x2_ASAP7_75t_L g1321 ( 
.A1(n_1148),
.A2(n_1168),
.A3(n_1063),
.B(n_1181),
.Y(n_1321)
);

AO21x2_ASAP7_75t_L g1322 ( 
.A1(n_1148),
.A2(n_1168),
.B(n_1063),
.Y(n_1322)
);

NAND2xp5_ASAP7_75t_L g1323 ( 
.A(n_1067),
.B(n_864),
.Y(n_1323)
);

OAI21xp5_ASAP7_75t_L g1324 ( 
.A1(n_1063),
.A2(n_880),
.B(n_864),
.Y(n_1324)
);

NAND2xp5_ASAP7_75t_L g1325 ( 
.A(n_1067),
.B(n_864),
.Y(n_1325)
);

AOI21xp5_ASAP7_75t_L g1326 ( 
.A1(n_1063),
.A2(n_949),
.B(n_1168),
.Y(n_1326)
);

AO31x2_ASAP7_75t_L g1327 ( 
.A1(n_1148),
.A2(n_1168),
.A3(n_1063),
.B(n_1181),
.Y(n_1327)
);

INVx1_ASAP7_75t_SL g1328 ( 
.A(n_1062),
.Y(n_1328)
);

OAI21xp5_ASAP7_75t_L g1329 ( 
.A1(n_1063),
.A2(n_880),
.B(n_1135),
.Y(n_1329)
);

NOR2xp67_ASAP7_75t_L g1330 ( 
.A(n_1082),
.B(n_1030),
.Y(n_1330)
);

OAI21x1_ASAP7_75t_SL g1331 ( 
.A1(n_1135),
.A2(n_1127),
.B(n_1140),
.Y(n_1331)
);

AND2x4_ASAP7_75t_L g1332 ( 
.A(n_1132),
.B(n_1098),
.Y(n_1332)
);

A2O1A1Ixp33_ASAP7_75t_L g1333 ( 
.A1(n_1063),
.A2(n_864),
.B(n_880),
.C(n_1130),
.Y(n_1333)
);

OAI22xp5_ASAP7_75t_L g1334 ( 
.A1(n_1063),
.A2(n_864),
.B1(n_880),
.B2(n_1067),
.Y(n_1334)
);

AOI21xp5_ASAP7_75t_L g1335 ( 
.A1(n_1063),
.A2(n_949),
.B(n_1168),
.Y(n_1335)
);

AOI22xp33_ASAP7_75t_L g1336 ( 
.A1(n_1130),
.A2(n_864),
.B1(n_1056),
.B2(n_811),
.Y(n_1336)
);

AND2x4_ASAP7_75t_L g1337 ( 
.A(n_1132),
.B(n_1098),
.Y(n_1337)
);

AO31x2_ASAP7_75t_L g1338 ( 
.A1(n_1148),
.A2(n_1168),
.A3(n_1063),
.B(n_1181),
.Y(n_1338)
);

NAND2xp5_ASAP7_75t_L g1339 ( 
.A(n_1067),
.B(n_864),
.Y(n_1339)
);

AOI21xp5_ASAP7_75t_L g1340 ( 
.A1(n_1063),
.A2(n_949),
.B(n_1168),
.Y(n_1340)
);

AOI21xp5_ASAP7_75t_L g1341 ( 
.A1(n_1063),
.A2(n_949),
.B(n_1168),
.Y(n_1341)
);

AND2x4_ASAP7_75t_L g1342 ( 
.A(n_1132),
.B(n_1098),
.Y(n_1342)
);

NAND2xp5_ASAP7_75t_SL g1343 ( 
.A(n_1067),
.B(n_877),
.Y(n_1343)
);

NOR2xp33_ASAP7_75t_L g1344 ( 
.A(n_1067),
.B(n_864),
.Y(n_1344)
);

OAI21x1_ASAP7_75t_L g1345 ( 
.A1(n_1166),
.A2(n_1152),
.B(n_1171),
.Y(n_1345)
);

AOI21xp5_ASAP7_75t_L g1346 ( 
.A1(n_1063),
.A2(n_949),
.B(n_1168),
.Y(n_1346)
);

AOI22xp33_ASAP7_75t_SL g1347 ( 
.A1(n_1291),
.A2(n_1315),
.B1(n_1344),
.B2(n_1220),
.Y(n_1347)
);

CKINVDCx5p33_ASAP7_75t_R g1348 ( 
.A(n_1285),
.Y(n_1348)
);

BUFx3_ASAP7_75t_L g1349 ( 
.A(n_1240),
.Y(n_1349)
);

OAI21xp5_ASAP7_75t_SL g1350 ( 
.A1(n_1306),
.A2(n_1336),
.B(n_1200),
.Y(n_1350)
);

INVx4_ASAP7_75t_L g1351 ( 
.A(n_1209),
.Y(n_1351)
);

BUFx12f_ASAP7_75t_L g1352 ( 
.A(n_1199),
.Y(n_1352)
);

NAND2xp5_ASAP7_75t_L g1353 ( 
.A(n_1214),
.B(n_1212),
.Y(n_1353)
);

OR2x2_ASAP7_75t_L g1354 ( 
.A(n_1205),
.B(n_1215),
.Y(n_1354)
);

INVx2_ASAP7_75t_L g1355 ( 
.A(n_1308),
.Y(n_1355)
);

BUFx12f_ASAP7_75t_L g1356 ( 
.A(n_1199),
.Y(n_1356)
);

CKINVDCx5p33_ASAP7_75t_R g1357 ( 
.A(n_1254),
.Y(n_1357)
);

BUFx3_ASAP7_75t_L g1358 ( 
.A(n_1320),
.Y(n_1358)
);

OAI22xp33_ASAP7_75t_L g1359 ( 
.A1(n_1275),
.A2(n_1323),
.B1(n_1284),
.B2(n_1305),
.Y(n_1359)
);

CKINVDCx20_ASAP7_75t_R g1360 ( 
.A(n_1267),
.Y(n_1360)
);

OAI22xp33_ASAP7_75t_L g1361 ( 
.A1(n_1290),
.A2(n_1325),
.B1(n_1339),
.B2(n_1312),
.Y(n_1361)
);

OAI22xp33_ASAP7_75t_L g1362 ( 
.A1(n_1312),
.A2(n_1277),
.B1(n_1334),
.B2(n_1300),
.Y(n_1362)
);

INVx8_ASAP7_75t_L g1363 ( 
.A(n_1274),
.Y(n_1363)
);

CKINVDCx6p67_ASAP7_75t_R g1364 ( 
.A(n_1209),
.Y(n_1364)
);

CKINVDCx11_ASAP7_75t_R g1365 ( 
.A(n_1220),
.Y(n_1365)
);

BUFx4f_ASAP7_75t_SL g1366 ( 
.A(n_1199),
.Y(n_1366)
);

AOI22xp33_ASAP7_75t_SL g1367 ( 
.A1(n_1227),
.A2(n_1324),
.B1(n_1276),
.B2(n_1329),
.Y(n_1367)
);

BUFx10_ASAP7_75t_L g1368 ( 
.A(n_1332),
.Y(n_1368)
);

HB1xp67_ASAP7_75t_L g1369 ( 
.A(n_1207),
.Y(n_1369)
);

BUFx8_ASAP7_75t_L g1370 ( 
.A(n_1241),
.Y(n_1370)
);

AOI22xp33_ASAP7_75t_SL g1371 ( 
.A1(n_1318),
.A2(n_1329),
.B1(n_1237),
.B2(n_1223),
.Y(n_1371)
);

OAI22xp33_ASAP7_75t_L g1372 ( 
.A1(n_1235),
.A2(n_1203),
.B1(n_1330),
.B2(n_1228),
.Y(n_1372)
);

AOI22xp5_ASAP7_75t_L g1373 ( 
.A1(n_1314),
.A2(n_1292),
.B1(n_1333),
.B2(n_1302),
.Y(n_1373)
);

AOI22xp33_ASAP7_75t_SL g1374 ( 
.A1(n_1318),
.A2(n_1299),
.B1(n_1297),
.B2(n_1283),
.Y(n_1374)
);

AOI22xp33_ASAP7_75t_L g1375 ( 
.A1(n_1230),
.A2(n_1343),
.B1(n_1330),
.B2(n_1202),
.Y(n_1375)
);

BUFx12f_ASAP7_75t_L g1376 ( 
.A(n_1241),
.Y(n_1376)
);

INVx3_ASAP7_75t_L g1377 ( 
.A(n_1268),
.Y(n_1377)
);

INVx6_ASAP7_75t_L g1378 ( 
.A(n_1209),
.Y(n_1378)
);

NAND2xp5_ASAP7_75t_L g1379 ( 
.A(n_1296),
.B(n_1270),
.Y(n_1379)
);

INVx4_ASAP7_75t_L g1380 ( 
.A(n_1274),
.Y(n_1380)
);

OAI22xp33_ASAP7_75t_L g1381 ( 
.A1(n_1204),
.A2(n_1264),
.B1(n_1328),
.B2(n_1207),
.Y(n_1381)
);

AOI22xp33_ASAP7_75t_L g1382 ( 
.A1(n_1202),
.A2(n_1271),
.B1(n_1196),
.B2(n_1269),
.Y(n_1382)
);

BUFx4f_ASAP7_75t_L g1383 ( 
.A(n_1274),
.Y(n_1383)
);

AOI22xp33_ASAP7_75t_L g1384 ( 
.A1(n_1196),
.A2(n_1226),
.B1(n_1231),
.B2(n_1331),
.Y(n_1384)
);

AOI22xp33_ASAP7_75t_L g1385 ( 
.A1(n_1328),
.A2(n_1322),
.B1(n_1262),
.B2(n_1242),
.Y(n_1385)
);

NAND2x1p5_ASAP7_75t_L g1386 ( 
.A(n_1273),
.B(n_1250),
.Y(n_1386)
);

INVx3_ASAP7_75t_SL g1387 ( 
.A(n_1332),
.Y(n_1387)
);

AOI22xp33_ASAP7_75t_SL g1388 ( 
.A1(n_1322),
.A2(n_1263),
.B1(n_1261),
.B2(n_1340),
.Y(n_1388)
);

CKINVDCx20_ASAP7_75t_R g1389 ( 
.A(n_1260),
.Y(n_1389)
);

OAI22xp5_ASAP7_75t_L g1390 ( 
.A1(n_1216),
.A2(n_1229),
.B1(n_1246),
.B2(n_1219),
.Y(n_1390)
);

BUFx2_ASAP7_75t_R g1391 ( 
.A(n_1236),
.Y(n_1391)
);

CKINVDCx11_ASAP7_75t_R g1392 ( 
.A(n_1279),
.Y(n_1392)
);

OAI22xp5_ASAP7_75t_L g1393 ( 
.A1(n_1217),
.A2(n_1218),
.B1(n_1248),
.B2(n_1249),
.Y(n_1393)
);

INVxp67_ASAP7_75t_L g1394 ( 
.A(n_1244),
.Y(n_1394)
);

INVx8_ASAP7_75t_L g1395 ( 
.A(n_1274),
.Y(n_1395)
);

OAI22xp5_ASAP7_75t_L g1396 ( 
.A1(n_1233),
.A2(n_1243),
.B1(n_1234),
.B2(n_1251),
.Y(n_1396)
);

INVx2_ASAP7_75t_L g1397 ( 
.A(n_1258),
.Y(n_1397)
);

OAI22xp5_ASAP7_75t_L g1398 ( 
.A1(n_1222),
.A2(n_1256),
.B1(n_1341),
.B2(n_1335),
.Y(n_1398)
);

BUFx4f_ASAP7_75t_SL g1399 ( 
.A(n_1279),
.Y(n_1399)
);

INVx2_ASAP7_75t_L g1400 ( 
.A(n_1268),
.Y(n_1400)
);

OAI22x1_ASAP7_75t_SL g1401 ( 
.A1(n_1273),
.A2(n_1298),
.B1(n_1250),
.B2(n_1236),
.Y(n_1401)
);

BUFx10_ASAP7_75t_L g1402 ( 
.A(n_1337),
.Y(n_1402)
);

BUFx12f_ASAP7_75t_L g1403 ( 
.A(n_1309),
.Y(n_1403)
);

CKINVDCx20_ASAP7_75t_R g1404 ( 
.A(n_1311),
.Y(n_1404)
);

AOI22xp33_ASAP7_75t_L g1405 ( 
.A1(n_1224),
.A2(n_1342),
.B1(n_1346),
.B2(n_1326),
.Y(n_1405)
);

INVx1_ASAP7_75t_L g1406 ( 
.A(n_1255),
.Y(n_1406)
);

INVx6_ASAP7_75t_L g1407 ( 
.A(n_1309),
.Y(n_1407)
);

INVx2_ASAP7_75t_L g1408 ( 
.A(n_1253),
.Y(n_1408)
);

OAI22xp33_ASAP7_75t_L g1409 ( 
.A1(n_1278),
.A2(n_1316),
.B1(n_1301),
.B2(n_1294),
.Y(n_1409)
);

INVx3_ASAP7_75t_L g1410 ( 
.A(n_1253),
.Y(n_1410)
);

AOI22xp33_ASAP7_75t_L g1411 ( 
.A1(n_1224),
.A2(n_1263),
.B1(n_1195),
.B2(n_1238),
.Y(n_1411)
);

BUFx2_ASAP7_75t_SL g1412 ( 
.A(n_1309),
.Y(n_1412)
);

AOI22xp33_ASAP7_75t_SL g1413 ( 
.A1(n_1221),
.A2(n_1222),
.B1(n_1287),
.B2(n_1252),
.Y(n_1413)
);

CKINVDCx6p67_ASAP7_75t_R g1414 ( 
.A(n_1295),
.Y(n_1414)
);

AOI22xp33_ASAP7_75t_SL g1415 ( 
.A1(n_1252),
.A2(n_1289),
.B1(n_1195),
.B2(n_1286),
.Y(n_1415)
);

AOI22xp33_ASAP7_75t_SL g1416 ( 
.A1(n_1252),
.A2(n_1289),
.B1(n_1282),
.B2(n_1213),
.Y(n_1416)
);

CKINVDCx5p33_ASAP7_75t_R g1417 ( 
.A(n_1313),
.Y(n_1417)
);

INVx2_ASAP7_75t_L g1418 ( 
.A(n_1313),
.Y(n_1418)
);

INVx1_ASAP7_75t_L g1419 ( 
.A(n_1255),
.Y(n_1419)
);

AOI22xp5_ASAP7_75t_L g1420 ( 
.A1(n_1245),
.A2(n_1265),
.B1(n_1232),
.B2(n_1266),
.Y(n_1420)
);

AOI22xp33_ASAP7_75t_L g1421 ( 
.A1(n_1265),
.A2(n_1201),
.B1(n_1257),
.B2(n_1211),
.Y(n_1421)
);

NAND2xp5_ASAP7_75t_L g1422 ( 
.A(n_1208),
.B(n_1280),
.Y(n_1422)
);

INVx6_ASAP7_75t_L g1423 ( 
.A(n_1247),
.Y(n_1423)
);

NAND2xp5_ASAP7_75t_L g1424 ( 
.A(n_1208),
.B(n_1303),
.Y(n_1424)
);

INVx1_ASAP7_75t_L g1425 ( 
.A(n_1208),
.Y(n_1425)
);

AOI22xp33_ASAP7_75t_L g1426 ( 
.A1(n_1201),
.A2(n_1206),
.B1(n_1198),
.B2(n_1259),
.Y(n_1426)
);

INVx6_ASAP7_75t_L g1427 ( 
.A(n_1225),
.Y(n_1427)
);

AOI22xp33_ASAP7_75t_SL g1428 ( 
.A1(n_1210),
.A2(n_1206),
.B1(n_1319),
.B2(n_1345),
.Y(n_1428)
);

NAND2xp5_ASAP7_75t_L g1429 ( 
.A(n_1338),
.B(n_1327),
.Y(n_1429)
);

INVx1_ASAP7_75t_L g1430 ( 
.A(n_1197),
.Y(n_1430)
);

INVx4_ASAP7_75t_L g1431 ( 
.A(n_1288),
.Y(n_1431)
);

BUFx12f_ASAP7_75t_L g1432 ( 
.A(n_1239),
.Y(n_1432)
);

INVx3_ASAP7_75t_SL g1433 ( 
.A(n_1197),
.Y(n_1433)
);

NAND2xp5_ASAP7_75t_L g1434 ( 
.A(n_1280),
.B(n_1338),
.Y(n_1434)
);

INVx1_ASAP7_75t_L g1435 ( 
.A(n_1280),
.Y(n_1435)
);

CKINVDCx5p33_ASAP7_75t_R g1436 ( 
.A(n_1303),
.Y(n_1436)
);

OAI21xp33_ASAP7_75t_SL g1437 ( 
.A1(n_1272),
.A2(n_1281),
.B(n_1293),
.Y(n_1437)
);

NAND2xp5_ASAP7_75t_L g1438 ( 
.A(n_1307),
.B(n_1310),
.Y(n_1438)
);

OAI22xp33_ASAP7_75t_L g1439 ( 
.A1(n_1307),
.A2(n_1310),
.B1(n_1321),
.B2(n_1327),
.Y(n_1439)
);

BUFx2_ASAP7_75t_L g1440 ( 
.A(n_1307),
.Y(n_1440)
);

INVx3_ASAP7_75t_L g1441 ( 
.A(n_1310),
.Y(n_1441)
);

AOI22xp33_ASAP7_75t_SL g1442 ( 
.A1(n_1317),
.A2(n_1321),
.B1(n_1327),
.B2(n_1338),
.Y(n_1442)
);

CKINVDCx20_ASAP7_75t_R g1443 ( 
.A(n_1321),
.Y(n_1443)
);

INVx2_ASAP7_75t_SL g1444 ( 
.A(n_1320),
.Y(n_1444)
);

INVx3_ASAP7_75t_L g1445 ( 
.A(n_1268),
.Y(n_1445)
);

CKINVDCx11_ASAP7_75t_R g1446 ( 
.A(n_1285),
.Y(n_1446)
);

AOI22xp33_ASAP7_75t_L g1447 ( 
.A1(n_1312),
.A2(n_864),
.B1(n_1130),
.B2(n_1306),
.Y(n_1447)
);

AOI22xp5_ASAP7_75t_L g1448 ( 
.A1(n_1291),
.A2(n_864),
.B1(n_1344),
.B2(n_1315),
.Y(n_1448)
);

BUFx10_ASAP7_75t_L g1449 ( 
.A(n_1332),
.Y(n_1449)
);

INVx1_ASAP7_75t_L g1450 ( 
.A(n_1304),
.Y(n_1450)
);

CKINVDCx5p33_ASAP7_75t_R g1451 ( 
.A(n_1285),
.Y(n_1451)
);

CKINVDCx10_ASAP7_75t_R g1452 ( 
.A(n_1267),
.Y(n_1452)
);

AND2x2_ASAP7_75t_L g1453 ( 
.A(n_1283),
.B(n_1297),
.Y(n_1453)
);

CKINVDCx20_ASAP7_75t_R g1454 ( 
.A(n_1285),
.Y(n_1454)
);

NAND2xp5_ASAP7_75t_L g1455 ( 
.A(n_1214),
.B(n_1212),
.Y(n_1455)
);

BUFx2_ASAP7_75t_SL g1456 ( 
.A(n_1285),
.Y(n_1456)
);

AOI22xp5_ASAP7_75t_L g1457 ( 
.A1(n_1291),
.A2(n_864),
.B1(n_1344),
.B2(n_1315),
.Y(n_1457)
);

INVx6_ASAP7_75t_L g1458 ( 
.A(n_1240),
.Y(n_1458)
);

CKINVDCx20_ASAP7_75t_R g1459 ( 
.A(n_1285),
.Y(n_1459)
);

AOI22xp33_ASAP7_75t_SL g1460 ( 
.A1(n_1291),
.A2(n_864),
.B1(n_1130),
.B2(n_926),
.Y(n_1460)
);

AOI22xp33_ASAP7_75t_SL g1461 ( 
.A1(n_1291),
.A2(n_864),
.B1(n_1130),
.B2(n_926),
.Y(n_1461)
);

AO22x1_ASAP7_75t_L g1462 ( 
.A1(n_1291),
.A2(n_864),
.B1(n_1130),
.B2(n_1315),
.Y(n_1462)
);

INVx6_ASAP7_75t_L g1463 ( 
.A(n_1240),
.Y(n_1463)
);

INVx1_ASAP7_75t_SL g1464 ( 
.A(n_1207),
.Y(n_1464)
);

AOI22xp33_ASAP7_75t_L g1465 ( 
.A1(n_1312),
.A2(n_864),
.B1(n_1130),
.B2(n_1306),
.Y(n_1465)
);

INVx1_ASAP7_75t_L g1466 ( 
.A(n_1304),
.Y(n_1466)
);

BUFx3_ASAP7_75t_L g1467 ( 
.A(n_1240),
.Y(n_1467)
);

BUFx8_ASAP7_75t_L g1468 ( 
.A(n_1240),
.Y(n_1468)
);

INVx2_ASAP7_75t_SL g1469 ( 
.A(n_1320),
.Y(n_1469)
);

AOI21xp5_ASAP7_75t_SL g1470 ( 
.A1(n_1292),
.A2(n_1063),
.B(n_1296),
.Y(n_1470)
);

AOI21xp5_ASAP7_75t_SL g1471 ( 
.A1(n_1292),
.A2(n_1063),
.B(n_1296),
.Y(n_1471)
);

AOI22xp33_ASAP7_75t_L g1472 ( 
.A1(n_1312),
.A2(n_864),
.B1(n_1130),
.B2(n_1306),
.Y(n_1472)
);

AOI22xp5_ASAP7_75t_L g1473 ( 
.A1(n_1291),
.A2(n_864),
.B1(n_1344),
.B2(n_1315),
.Y(n_1473)
);

INVx4_ASAP7_75t_L g1474 ( 
.A(n_1209),
.Y(n_1474)
);

AOI22xp33_ASAP7_75t_L g1475 ( 
.A1(n_1312),
.A2(n_864),
.B1(n_1130),
.B2(n_1306),
.Y(n_1475)
);

NOR2xp33_ASAP7_75t_L g1476 ( 
.A(n_1448),
.B(n_1457),
.Y(n_1476)
);

HB1xp67_ASAP7_75t_L g1477 ( 
.A(n_1369),
.Y(n_1477)
);

INVx1_ASAP7_75t_L g1478 ( 
.A(n_1406),
.Y(n_1478)
);

OAI21x1_ASAP7_75t_L g1479 ( 
.A1(n_1426),
.A2(n_1421),
.B(n_1398),
.Y(n_1479)
);

AO21x2_ASAP7_75t_L g1480 ( 
.A1(n_1409),
.A2(n_1362),
.B(n_1398),
.Y(n_1480)
);

INVx2_ASAP7_75t_L g1481 ( 
.A(n_1430),
.Y(n_1481)
);

INVx2_ASAP7_75t_L g1482 ( 
.A(n_1435),
.Y(n_1482)
);

BUFx3_ASAP7_75t_L g1483 ( 
.A(n_1423),
.Y(n_1483)
);

NAND2xp5_ASAP7_75t_L g1484 ( 
.A(n_1361),
.B(n_1353),
.Y(n_1484)
);

INVx1_ASAP7_75t_L g1485 ( 
.A(n_1419),
.Y(n_1485)
);

INVx1_ASAP7_75t_L g1486 ( 
.A(n_1425),
.Y(n_1486)
);

HB1xp67_ASAP7_75t_L g1487 ( 
.A(n_1464),
.Y(n_1487)
);

INVx1_ASAP7_75t_L g1488 ( 
.A(n_1440),
.Y(n_1488)
);

INVx1_ASAP7_75t_L g1489 ( 
.A(n_1436),
.Y(n_1489)
);

NAND4xp25_ASAP7_75t_L g1490 ( 
.A(n_1448),
.B(n_1473),
.C(n_1457),
.D(n_1447),
.Y(n_1490)
);

INVx1_ASAP7_75t_L g1491 ( 
.A(n_1429),
.Y(n_1491)
);

BUFx3_ASAP7_75t_L g1492 ( 
.A(n_1423),
.Y(n_1492)
);

NAND2xp5_ASAP7_75t_L g1493 ( 
.A(n_1353),
.B(n_1455),
.Y(n_1493)
);

OA21x2_ASAP7_75t_L g1494 ( 
.A1(n_1429),
.A2(n_1434),
.B(n_1424),
.Y(n_1494)
);

AND2x2_ASAP7_75t_L g1495 ( 
.A(n_1367),
.B(n_1371),
.Y(n_1495)
);

BUFx3_ASAP7_75t_L g1496 ( 
.A(n_1378),
.Y(n_1496)
);

NOR2xp33_ASAP7_75t_L g1497 ( 
.A(n_1473),
.B(n_1462),
.Y(n_1497)
);

INVx1_ASAP7_75t_L g1498 ( 
.A(n_1434),
.Y(n_1498)
);

INVx1_ASAP7_75t_L g1499 ( 
.A(n_1422),
.Y(n_1499)
);

CKINVDCx5p33_ASAP7_75t_R g1500 ( 
.A(n_1446),
.Y(n_1500)
);

INVx1_ASAP7_75t_L g1501 ( 
.A(n_1422),
.Y(n_1501)
);

BUFx12f_ASAP7_75t_L g1502 ( 
.A(n_1348),
.Y(n_1502)
);

INVx2_ASAP7_75t_L g1503 ( 
.A(n_1441),
.Y(n_1503)
);

BUFx3_ASAP7_75t_L g1504 ( 
.A(n_1378),
.Y(n_1504)
);

BUFx2_ASAP7_75t_L g1505 ( 
.A(n_1443),
.Y(n_1505)
);

OR2x2_ASAP7_75t_L g1506 ( 
.A(n_1424),
.B(n_1438),
.Y(n_1506)
);

OAI21xp33_ASAP7_75t_SL g1507 ( 
.A1(n_1373),
.A2(n_1470),
.B(n_1471),
.Y(n_1507)
);

INVx1_ASAP7_75t_L g1508 ( 
.A(n_1439),
.Y(n_1508)
);

AOI22xp33_ASAP7_75t_L g1509 ( 
.A1(n_1465),
.A2(n_1475),
.B1(n_1472),
.B2(n_1461),
.Y(n_1509)
);

BUFx2_ASAP7_75t_L g1510 ( 
.A(n_1432),
.Y(n_1510)
);

CKINVDCx5p33_ASAP7_75t_R g1511 ( 
.A(n_1452),
.Y(n_1511)
);

INVx2_ASAP7_75t_L g1512 ( 
.A(n_1433),
.Y(n_1512)
);

INVx1_ASAP7_75t_L g1513 ( 
.A(n_1393),
.Y(n_1513)
);

INVx1_ASAP7_75t_L g1514 ( 
.A(n_1393),
.Y(n_1514)
);

AND2x6_ASAP7_75t_L g1515 ( 
.A(n_1373),
.B(n_1379),
.Y(n_1515)
);

HB1xp67_ASAP7_75t_L g1516 ( 
.A(n_1396),
.Y(n_1516)
);

NOR2xp33_ASAP7_75t_L g1517 ( 
.A(n_1359),
.B(n_1354),
.Y(n_1517)
);

AOI21x1_ASAP7_75t_L g1518 ( 
.A1(n_1390),
.A2(n_1379),
.B(n_1396),
.Y(n_1518)
);

AND2x2_ASAP7_75t_L g1519 ( 
.A(n_1415),
.B(n_1413),
.Y(n_1519)
);

INVx3_ASAP7_75t_L g1520 ( 
.A(n_1431),
.Y(n_1520)
);

AOI22xp33_ASAP7_75t_L g1521 ( 
.A1(n_1460),
.A2(n_1390),
.B1(n_1374),
.B2(n_1372),
.Y(n_1521)
);

INVx2_ASAP7_75t_L g1522 ( 
.A(n_1431),
.Y(n_1522)
);

AOI21xp5_ASAP7_75t_L g1523 ( 
.A1(n_1437),
.A2(n_1411),
.B(n_1428),
.Y(n_1523)
);

INVx2_ASAP7_75t_SL g1524 ( 
.A(n_1368),
.Y(n_1524)
);

AND2x4_ASAP7_75t_L g1525 ( 
.A(n_1420),
.B(n_1384),
.Y(n_1525)
);

INVx1_ASAP7_75t_L g1526 ( 
.A(n_1442),
.Y(n_1526)
);

INVx1_ASAP7_75t_L g1527 ( 
.A(n_1416),
.Y(n_1527)
);

INVx1_ASAP7_75t_L g1528 ( 
.A(n_1388),
.Y(n_1528)
);

AND2x2_ASAP7_75t_L g1529 ( 
.A(n_1453),
.B(n_1450),
.Y(n_1529)
);

OAI21x1_ASAP7_75t_L g1530 ( 
.A1(n_1382),
.A2(n_1405),
.B(n_1385),
.Y(n_1530)
);

BUFx2_ASAP7_75t_L g1531 ( 
.A(n_1427),
.Y(n_1531)
);

AOI22xp33_ASAP7_75t_SL g1532 ( 
.A1(n_1427),
.A2(n_1350),
.B1(n_1455),
.B2(n_1474),
.Y(n_1532)
);

INVx2_ASAP7_75t_L g1533 ( 
.A(n_1466),
.Y(n_1533)
);

INVx1_ASAP7_75t_SL g1534 ( 
.A(n_1404),
.Y(n_1534)
);

BUFx2_ASAP7_75t_L g1535 ( 
.A(n_1437),
.Y(n_1535)
);

OAI21x1_ASAP7_75t_L g1536 ( 
.A1(n_1397),
.A2(n_1375),
.B(n_1355),
.Y(n_1536)
);

NAND2xp5_ASAP7_75t_SL g1537 ( 
.A(n_1347),
.B(n_1381),
.Y(n_1537)
);

OAI21x1_ASAP7_75t_L g1538 ( 
.A1(n_1410),
.A2(n_1408),
.B(n_1418),
.Y(n_1538)
);

INVx1_ASAP7_75t_L g1539 ( 
.A(n_1350),
.Y(n_1539)
);

OR2x6_ASAP7_75t_L g1540 ( 
.A(n_1363),
.B(n_1395),
.Y(n_1540)
);

INVx1_ASAP7_75t_L g1541 ( 
.A(n_1400),
.Y(n_1541)
);

INVx1_ASAP7_75t_L g1542 ( 
.A(n_1380),
.Y(n_1542)
);

INVx4_ASAP7_75t_L g1543 ( 
.A(n_1363),
.Y(n_1543)
);

BUFx2_ASAP7_75t_L g1544 ( 
.A(n_1351),
.Y(n_1544)
);

INVx1_ASAP7_75t_L g1545 ( 
.A(n_1380),
.Y(n_1545)
);

OAI21x1_ASAP7_75t_L g1546 ( 
.A1(n_1377),
.A2(n_1445),
.B(n_1386),
.Y(n_1546)
);

OR2x2_ASAP7_75t_L g1547 ( 
.A(n_1351),
.B(n_1474),
.Y(n_1547)
);

AND2x2_ASAP7_75t_L g1548 ( 
.A(n_1445),
.B(n_1364),
.Y(n_1548)
);

INVx1_ASAP7_75t_L g1549 ( 
.A(n_1363),
.Y(n_1549)
);

OAI22xp5_ASAP7_75t_L g1550 ( 
.A1(n_1383),
.A2(n_1391),
.B1(n_1394),
.B2(n_1387),
.Y(n_1550)
);

INVx2_ASAP7_75t_L g1551 ( 
.A(n_1368),
.Y(n_1551)
);

INVx2_ASAP7_75t_L g1552 ( 
.A(n_1402),
.Y(n_1552)
);

A2O1A1Ixp33_ASAP7_75t_L g1553 ( 
.A1(n_1383),
.A2(n_1395),
.B(n_1417),
.C(n_1444),
.Y(n_1553)
);

INVx1_ASAP7_75t_L g1554 ( 
.A(n_1395),
.Y(n_1554)
);

CKINVDCx20_ASAP7_75t_R g1555 ( 
.A(n_1454),
.Y(n_1555)
);

INVx1_ASAP7_75t_L g1556 ( 
.A(n_1401),
.Y(n_1556)
);

OAI21xp5_ASAP7_75t_L g1557 ( 
.A1(n_1386),
.A2(n_1389),
.B(n_1469),
.Y(n_1557)
);

OA21x2_ASAP7_75t_L g1558 ( 
.A1(n_1357),
.A2(n_1414),
.B(n_1412),
.Y(n_1558)
);

OAI21x1_ASAP7_75t_L g1559 ( 
.A1(n_1370),
.A2(n_1402),
.B(n_1449),
.Y(n_1559)
);

CKINVDCx5p33_ASAP7_75t_R g1560 ( 
.A(n_1452),
.Y(n_1560)
);

OAI21xp5_ASAP7_75t_L g1561 ( 
.A1(n_1459),
.A2(n_1360),
.B(n_1451),
.Y(n_1561)
);

INVx2_ASAP7_75t_L g1562 ( 
.A(n_1449),
.Y(n_1562)
);

OR2x2_ASAP7_75t_L g1563 ( 
.A(n_1456),
.B(n_1358),
.Y(n_1563)
);

INVx3_ASAP7_75t_L g1564 ( 
.A(n_1352),
.Y(n_1564)
);

AND2x2_ASAP7_75t_L g1565 ( 
.A(n_1505),
.B(n_1365),
.Y(n_1565)
);

AND2x4_ASAP7_75t_L g1566 ( 
.A(n_1512),
.B(n_1349),
.Y(n_1566)
);

AOI22xp5_ASAP7_75t_L g1567 ( 
.A1(n_1507),
.A2(n_1463),
.B1(n_1458),
.B2(n_1467),
.Y(n_1567)
);

AND2x2_ASAP7_75t_L g1568 ( 
.A(n_1505),
.B(n_1392),
.Y(n_1568)
);

NAND2xp5_ASAP7_75t_L g1569 ( 
.A(n_1517),
.B(n_1370),
.Y(n_1569)
);

OA21x2_ASAP7_75t_L g1570 ( 
.A1(n_1479),
.A2(n_1407),
.B(n_1403),
.Y(n_1570)
);

INVx4_ASAP7_75t_L g1571 ( 
.A(n_1558),
.Y(n_1571)
);

HB1xp67_ASAP7_75t_L g1572 ( 
.A(n_1487),
.Y(n_1572)
);

OAI22xp5_ASAP7_75t_L g1573 ( 
.A1(n_1509),
.A2(n_1458),
.B1(n_1463),
.B2(n_1399),
.Y(n_1573)
);

OR2x2_ASAP7_75t_L g1574 ( 
.A(n_1489),
.B(n_1468),
.Y(n_1574)
);

A2O1A1Ixp33_ASAP7_75t_L g1575 ( 
.A1(n_1507),
.A2(n_1366),
.B(n_1356),
.C(n_1376),
.Y(n_1575)
);

AND2x2_ASAP7_75t_L g1576 ( 
.A(n_1489),
.B(n_1468),
.Y(n_1576)
);

NAND2xp5_ASAP7_75t_L g1577 ( 
.A(n_1493),
.B(n_1476),
.Y(n_1577)
);

AND2x2_ASAP7_75t_L g1578 ( 
.A(n_1526),
.B(n_1508),
.Y(n_1578)
);

AO32x2_ASAP7_75t_L g1579 ( 
.A1(n_1524),
.A2(n_1550),
.A3(n_1506),
.B1(n_1516),
.B2(n_1494),
.Y(n_1579)
);

NOR2x1_ASAP7_75t_R g1580 ( 
.A(n_1511),
.B(n_1560),
.Y(n_1580)
);

OAI21xp5_ASAP7_75t_L g1581 ( 
.A1(n_1537),
.A2(n_1497),
.B(n_1490),
.Y(n_1581)
);

AND2x2_ASAP7_75t_L g1582 ( 
.A(n_1529),
.B(n_1477),
.Y(n_1582)
);

OAI21x1_ASAP7_75t_L g1583 ( 
.A1(n_1479),
.A2(n_1523),
.B(n_1538),
.Y(n_1583)
);

OAI21xp5_ASAP7_75t_L g1584 ( 
.A1(n_1521),
.A2(n_1495),
.B(n_1532),
.Y(n_1584)
);

AND2x2_ASAP7_75t_L g1585 ( 
.A(n_1526),
.B(n_1508),
.Y(n_1585)
);

A2O1A1Ixp33_ASAP7_75t_L g1586 ( 
.A1(n_1495),
.A2(n_1525),
.B(n_1539),
.C(n_1484),
.Y(n_1586)
);

AOI221xp5_ASAP7_75t_L g1587 ( 
.A1(n_1539),
.A2(n_1528),
.B1(n_1513),
.B2(n_1514),
.C(n_1525),
.Y(n_1587)
);

HB1xp67_ASAP7_75t_L g1588 ( 
.A(n_1488),
.Y(n_1588)
);

OAI22xp5_ASAP7_75t_L g1589 ( 
.A1(n_1556),
.A2(n_1531),
.B1(n_1553),
.B2(n_1510),
.Y(n_1589)
);

HB1xp67_ASAP7_75t_L g1590 ( 
.A(n_1488),
.Y(n_1590)
);

AO32x2_ASAP7_75t_L g1591 ( 
.A1(n_1524),
.A2(n_1506),
.A3(n_1494),
.B1(n_1499),
.B2(n_1501),
.Y(n_1591)
);

AND2x2_ASAP7_75t_L g1592 ( 
.A(n_1528),
.B(n_1531),
.Y(n_1592)
);

BUFx10_ASAP7_75t_L g1593 ( 
.A(n_1500),
.Y(n_1593)
);

A2O1A1Ixp33_ASAP7_75t_L g1594 ( 
.A1(n_1525),
.A2(n_1514),
.B(n_1513),
.C(n_1530),
.Y(n_1594)
);

A2O1A1Ixp33_ASAP7_75t_L g1595 ( 
.A1(n_1525),
.A2(n_1530),
.B(n_1519),
.C(n_1527),
.Y(n_1595)
);

INVx4_ASAP7_75t_L g1596 ( 
.A(n_1558),
.Y(n_1596)
);

AOI22xp5_ASAP7_75t_SL g1597 ( 
.A1(n_1515),
.A2(n_1556),
.B1(n_1510),
.B2(n_1555),
.Y(n_1597)
);

AOI21x1_ASAP7_75t_L g1598 ( 
.A1(n_1522),
.A2(n_1518),
.B(n_1545),
.Y(n_1598)
);

INVx5_ASAP7_75t_L g1599 ( 
.A(n_1540),
.Y(n_1599)
);

A2O1A1Ixp33_ASAP7_75t_L g1600 ( 
.A1(n_1527),
.A2(n_1515),
.B(n_1480),
.C(n_1492),
.Y(n_1600)
);

NOR2xp33_ASAP7_75t_L g1601 ( 
.A(n_1518),
.B(n_1515),
.Y(n_1601)
);

OA21x2_ASAP7_75t_L g1602 ( 
.A1(n_1535),
.A2(n_1478),
.B(n_1485),
.Y(n_1602)
);

OR2x6_ASAP7_75t_L g1603 ( 
.A(n_1540),
.B(n_1522),
.Y(n_1603)
);

INVx1_ASAP7_75t_SL g1604 ( 
.A(n_1563),
.Y(n_1604)
);

AOI21xp5_ASAP7_75t_L g1605 ( 
.A1(n_1494),
.A2(n_1492),
.B(n_1483),
.Y(n_1605)
);

CKINVDCx20_ASAP7_75t_R g1606 ( 
.A(n_1502),
.Y(n_1606)
);

OAI22xp5_ASAP7_75t_L g1607 ( 
.A1(n_1483),
.A2(n_1492),
.B1(n_1557),
.B2(n_1504),
.Y(n_1607)
);

INVx4_ASAP7_75t_L g1608 ( 
.A(n_1558),
.Y(n_1608)
);

NOR2x1_ASAP7_75t_R g1609 ( 
.A(n_1502),
.B(n_1483),
.Y(n_1609)
);

AOI211xp5_ASAP7_75t_SL g1610 ( 
.A1(n_1542),
.A2(n_1545),
.B(n_1520),
.C(n_1547),
.Y(n_1610)
);

OAI21xp5_ASAP7_75t_L g1611 ( 
.A1(n_1536),
.A2(n_1515),
.B(n_1542),
.Y(n_1611)
);

NOR2xp33_ASAP7_75t_L g1612 ( 
.A(n_1515),
.B(n_1496),
.Y(n_1612)
);

AND2x2_ASAP7_75t_SL g1613 ( 
.A(n_1558),
.B(n_1494),
.Y(n_1613)
);

AO32x2_ASAP7_75t_L g1614 ( 
.A1(n_1491),
.A2(n_1498),
.A3(n_1543),
.B1(n_1482),
.B2(n_1486),
.Y(n_1614)
);

AND2x2_ASAP7_75t_L g1615 ( 
.A(n_1491),
.B(n_1498),
.Y(n_1615)
);

INVx2_ASAP7_75t_L g1616 ( 
.A(n_1481),
.Y(n_1616)
);

NAND2xp33_ASAP7_75t_R g1617 ( 
.A(n_1540),
.B(n_1544),
.Y(n_1617)
);

OAI21xp5_ASAP7_75t_L g1618 ( 
.A1(n_1536),
.A2(n_1559),
.B(n_1546),
.Y(n_1618)
);

AND2x2_ASAP7_75t_L g1619 ( 
.A(n_1481),
.B(n_1482),
.Y(n_1619)
);

AOI22xp33_ASAP7_75t_L g1620 ( 
.A1(n_1581),
.A2(n_1584),
.B1(n_1577),
.B2(n_1587),
.Y(n_1620)
);

HB1xp67_ASAP7_75t_L g1621 ( 
.A(n_1602),
.Y(n_1621)
);

AOI22xp33_ASAP7_75t_L g1622 ( 
.A1(n_1573),
.A2(n_1534),
.B1(n_1563),
.B2(n_1504),
.Y(n_1622)
);

AND2x2_ASAP7_75t_L g1623 ( 
.A(n_1614),
.B(n_1535),
.Y(n_1623)
);

HB1xp67_ASAP7_75t_L g1624 ( 
.A(n_1602),
.Y(n_1624)
);

INVx2_ASAP7_75t_L g1625 ( 
.A(n_1616),
.Y(n_1625)
);

AND2x2_ASAP7_75t_L g1626 ( 
.A(n_1614),
.B(n_1481),
.Y(n_1626)
);

AND2x2_ASAP7_75t_L g1627 ( 
.A(n_1614),
.B(n_1482),
.Y(n_1627)
);

BUFx4f_ASAP7_75t_SL g1628 ( 
.A(n_1606),
.Y(n_1628)
);

HB1xp67_ASAP7_75t_L g1629 ( 
.A(n_1602),
.Y(n_1629)
);

INVx3_ASAP7_75t_SL g1630 ( 
.A(n_1613),
.Y(n_1630)
);

OAI21xp5_ASAP7_75t_SL g1631 ( 
.A1(n_1586),
.A2(n_1561),
.B(n_1548),
.Y(n_1631)
);

AND2x2_ASAP7_75t_L g1632 ( 
.A(n_1614),
.B(n_1486),
.Y(n_1632)
);

AND2x2_ASAP7_75t_L g1633 ( 
.A(n_1613),
.B(n_1591),
.Y(n_1633)
);

AND2x2_ASAP7_75t_L g1634 ( 
.A(n_1591),
.B(n_1619),
.Y(n_1634)
);

BUFx3_ASAP7_75t_L g1635 ( 
.A(n_1599),
.Y(n_1635)
);

AOI22xp33_ASAP7_75t_L g1636 ( 
.A1(n_1601),
.A2(n_1504),
.B1(n_1541),
.B2(n_1533),
.Y(n_1636)
);

NOR2x1_ASAP7_75t_SL g1637 ( 
.A(n_1603),
.B(n_1540),
.Y(n_1637)
);

INVx2_ASAP7_75t_L g1638 ( 
.A(n_1616),
.Y(n_1638)
);

HB1xp67_ASAP7_75t_L g1639 ( 
.A(n_1588),
.Y(n_1639)
);

AOI22xp33_ASAP7_75t_L g1640 ( 
.A1(n_1568),
.A2(n_1551),
.B1(n_1552),
.B2(n_1562),
.Y(n_1640)
);

AND2x2_ASAP7_75t_L g1641 ( 
.A(n_1579),
.B(n_1503),
.Y(n_1641)
);

AND2x2_ASAP7_75t_L g1642 ( 
.A(n_1579),
.B(n_1503),
.Y(n_1642)
);

HB1xp67_ASAP7_75t_L g1643 ( 
.A(n_1590),
.Y(n_1643)
);

AND2x2_ASAP7_75t_L g1644 ( 
.A(n_1579),
.B(n_1615),
.Y(n_1644)
);

AOI22xp33_ASAP7_75t_SL g1645 ( 
.A1(n_1628),
.A2(n_1597),
.B1(n_1586),
.B2(n_1565),
.Y(n_1645)
);

AND2x2_ASAP7_75t_L g1646 ( 
.A(n_1634),
.B(n_1579),
.Y(n_1646)
);

INVx3_ASAP7_75t_L g1647 ( 
.A(n_1625),
.Y(n_1647)
);

NAND3xp33_ASAP7_75t_L g1648 ( 
.A(n_1620),
.B(n_1595),
.C(n_1600),
.Y(n_1648)
);

NAND2xp5_ASAP7_75t_L g1649 ( 
.A(n_1644),
.B(n_1572),
.Y(n_1649)
);

AOI33xp33_ASAP7_75t_L g1650 ( 
.A1(n_1620),
.A2(n_1568),
.A3(n_1585),
.B1(n_1578),
.B2(n_1565),
.B3(n_1604),
.Y(n_1650)
);

NOR2xp33_ASAP7_75t_L g1651 ( 
.A(n_1631),
.B(n_1569),
.Y(n_1651)
);

INVx2_ASAP7_75t_L g1652 ( 
.A(n_1626),
.Y(n_1652)
);

INVx2_ASAP7_75t_L g1653 ( 
.A(n_1626),
.Y(n_1653)
);

OAI21x1_ASAP7_75t_SL g1654 ( 
.A1(n_1637),
.A2(n_1605),
.B(n_1611),
.Y(n_1654)
);

INVx2_ASAP7_75t_L g1655 ( 
.A(n_1626),
.Y(n_1655)
);

OAI221xp5_ASAP7_75t_L g1656 ( 
.A1(n_1631),
.A2(n_1595),
.B1(n_1600),
.B2(n_1567),
.C(n_1594),
.Y(n_1656)
);

INVx1_ASAP7_75t_L g1657 ( 
.A(n_1625),
.Y(n_1657)
);

INVx2_ASAP7_75t_L g1658 ( 
.A(n_1627),
.Y(n_1658)
);

AND2x2_ASAP7_75t_L g1659 ( 
.A(n_1634),
.B(n_1583),
.Y(n_1659)
);

OR2x2_ASAP7_75t_L g1660 ( 
.A(n_1634),
.B(n_1571),
.Y(n_1660)
);

NAND2xp5_ASAP7_75t_L g1661 ( 
.A(n_1644),
.B(n_1594),
.Y(n_1661)
);

AND2x2_ASAP7_75t_L g1662 ( 
.A(n_1633),
.B(n_1583),
.Y(n_1662)
);

AOI22xp33_ASAP7_75t_L g1663 ( 
.A1(n_1622),
.A2(n_1612),
.B1(n_1592),
.B2(n_1578),
.Y(n_1663)
);

AOI221xp5_ASAP7_75t_L g1664 ( 
.A1(n_1633),
.A2(n_1589),
.B1(n_1585),
.B2(n_1582),
.C(n_1607),
.Y(n_1664)
);

INVx1_ASAP7_75t_L g1665 ( 
.A(n_1625),
.Y(n_1665)
);

INVx1_ASAP7_75t_L g1666 ( 
.A(n_1638),
.Y(n_1666)
);

AO21x2_ASAP7_75t_L g1667 ( 
.A1(n_1621),
.A2(n_1618),
.B(n_1598),
.Y(n_1667)
);

HB1xp67_ASAP7_75t_L g1668 ( 
.A(n_1621),
.Y(n_1668)
);

HB1xp67_ASAP7_75t_L g1669 ( 
.A(n_1624),
.Y(n_1669)
);

AND2x2_ASAP7_75t_L g1670 ( 
.A(n_1633),
.B(n_1570),
.Y(n_1670)
);

INVxp67_ASAP7_75t_SL g1671 ( 
.A(n_1624),
.Y(n_1671)
);

INVx1_ASAP7_75t_L g1672 ( 
.A(n_1632),
.Y(n_1672)
);

OAI221xp5_ASAP7_75t_L g1673 ( 
.A1(n_1622),
.A2(n_1640),
.B1(n_1575),
.B2(n_1636),
.C(n_1630),
.Y(n_1673)
);

OAI211xp5_ASAP7_75t_SL g1674 ( 
.A1(n_1640),
.A2(n_1574),
.B(n_1575),
.C(n_1610),
.Y(n_1674)
);

OR2x2_ASAP7_75t_L g1675 ( 
.A(n_1623),
.B(n_1571),
.Y(n_1675)
);

INVx1_ASAP7_75t_SL g1676 ( 
.A(n_1639),
.Y(n_1676)
);

INVx1_ASAP7_75t_L g1677 ( 
.A(n_1632),
.Y(n_1677)
);

INVx1_ASAP7_75t_L g1678 ( 
.A(n_1632),
.Y(n_1678)
);

AOI22xp33_ASAP7_75t_L g1679 ( 
.A1(n_1628),
.A2(n_1612),
.B1(n_1576),
.B2(n_1566),
.Y(n_1679)
);

AND2x2_ASAP7_75t_L g1680 ( 
.A(n_1644),
.B(n_1570),
.Y(n_1680)
);

BUFx3_ASAP7_75t_L g1681 ( 
.A(n_1635),
.Y(n_1681)
);

INVx1_ASAP7_75t_L g1682 ( 
.A(n_1657),
.Y(n_1682)
);

INVx3_ASAP7_75t_L g1683 ( 
.A(n_1647),
.Y(n_1683)
);

HB1xp67_ASAP7_75t_L g1684 ( 
.A(n_1668),
.Y(n_1684)
);

NAND2xp5_ASAP7_75t_L g1685 ( 
.A(n_1661),
.B(n_1643),
.Y(n_1685)
);

AND2x2_ASAP7_75t_L g1686 ( 
.A(n_1652),
.B(n_1623),
.Y(n_1686)
);

BUFx2_ASAP7_75t_L g1687 ( 
.A(n_1681),
.Y(n_1687)
);

NAND2xp5_ASAP7_75t_L g1688 ( 
.A(n_1661),
.B(n_1641),
.Y(n_1688)
);

AND2x2_ASAP7_75t_L g1689 ( 
.A(n_1652),
.B(n_1623),
.Y(n_1689)
);

HB1xp67_ASAP7_75t_L g1690 ( 
.A(n_1668),
.Y(n_1690)
);

NAND2xp5_ASAP7_75t_L g1691 ( 
.A(n_1676),
.B(n_1641),
.Y(n_1691)
);

AND2x2_ASAP7_75t_L g1692 ( 
.A(n_1652),
.B(n_1630),
.Y(n_1692)
);

INVx1_ASAP7_75t_L g1693 ( 
.A(n_1669),
.Y(n_1693)
);

AND2x2_ASAP7_75t_L g1694 ( 
.A(n_1652),
.B(n_1630),
.Y(n_1694)
);

AND2x2_ASAP7_75t_L g1695 ( 
.A(n_1653),
.B(n_1630),
.Y(n_1695)
);

INVx2_ASAP7_75t_SL g1696 ( 
.A(n_1681),
.Y(n_1696)
);

NOR2x1_ASAP7_75t_L g1697 ( 
.A(n_1648),
.B(n_1571),
.Y(n_1697)
);

OR2x2_ASAP7_75t_L g1698 ( 
.A(n_1653),
.B(n_1629),
.Y(n_1698)
);

INVx1_ASAP7_75t_L g1699 ( 
.A(n_1669),
.Y(n_1699)
);

INVxp67_ASAP7_75t_L g1700 ( 
.A(n_1676),
.Y(n_1700)
);

OR2x2_ASAP7_75t_L g1701 ( 
.A(n_1653),
.B(n_1655),
.Y(n_1701)
);

AND2x4_ASAP7_75t_L g1702 ( 
.A(n_1653),
.B(n_1637),
.Y(n_1702)
);

AND2x2_ASAP7_75t_L g1703 ( 
.A(n_1655),
.B(n_1641),
.Y(n_1703)
);

AND2x4_ASAP7_75t_L g1704 ( 
.A(n_1655),
.B(n_1635),
.Y(n_1704)
);

BUFx3_ASAP7_75t_L g1705 ( 
.A(n_1681),
.Y(n_1705)
);

AND2x2_ASAP7_75t_L g1706 ( 
.A(n_1655),
.B(n_1642),
.Y(n_1706)
);

NAND2xp5_ASAP7_75t_SL g1707 ( 
.A(n_1648),
.B(n_1596),
.Y(n_1707)
);

INVx1_ASAP7_75t_L g1708 ( 
.A(n_1657),
.Y(n_1708)
);

INVx1_ASAP7_75t_L g1709 ( 
.A(n_1657),
.Y(n_1709)
);

AND2x2_ASAP7_75t_L g1710 ( 
.A(n_1658),
.B(n_1642),
.Y(n_1710)
);

INVx1_ASAP7_75t_L g1711 ( 
.A(n_1665),
.Y(n_1711)
);

INVx2_ASAP7_75t_L g1712 ( 
.A(n_1647),
.Y(n_1712)
);

HB1xp67_ASAP7_75t_L g1713 ( 
.A(n_1671),
.Y(n_1713)
);

INVx1_ASAP7_75t_L g1714 ( 
.A(n_1666),
.Y(n_1714)
);

INVx2_ASAP7_75t_L g1715 ( 
.A(n_1647),
.Y(n_1715)
);

INVx1_ASAP7_75t_L g1716 ( 
.A(n_1684),
.Y(n_1716)
);

AND2x2_ASAP7_75t_L g1717 ( 
.A(n_1697),
.B(n_1680),
.Y(n_1717)
);

AND2x4_ASAP7_75t_L g1718 ( 
.A(n_1705),
.B(n_1681),
.Y(n_1718)
);

OR2x2_ASAP7_75t_L g1719 ( 
.A(n_1685),
.B(n_1675),
.Y(n_1719)
);

NAND2x1_ASAP7_75t_L g1720 ( 
.A(n_1697),
.B(n_1654),
.Y(n_1720)
);

INVx1_ASAP7_75t_L g1721 ( 
.A(n_1684),
.Y(n_1721)
);

INVx1_ASAP7_75t_L g1722 ( 
.A(n_1690),
.Y(n_1722)
);

INVx2_ASAP7_75t_SL g1723 ( 
.A(n_1705),
.Y(n_1723)
);

NAND2xp5_ASAP7_75t_SL g1724 ( 
.A(n_1707),
.B(n_1645),
.Y(n_1724)
);

INVxp67_ASAP7_75t_L g1725 ( 
.A(n_1707),
.Y(n_1725)
);

OR2x2_ASAP7_75t_L g1726 ( 
.A(n_1685),
.B(n_1688),
.Y(n_1726)
);

INVx1_ASAP7_75t_L g1727 ( 
.A(n_1690),
.Y(n_1727)
);

AND2x2_ASAP7_75t_L g1728 ( 
.A(n_1705),
.B(n_1680),
.Y(n_1728)
);

AOI21xp5_ASAP7_75t_L g1729 ( 
.A1(n_1700),
.A2(n_1656),
.B(n_1645),
.Y(n_1729)
);

AND2x2_ASAP7_75t_L g1730 ( 
.A(n_1705),
.B(n_1680),
.Y(n_1730)
);

INVx1_ASAP7_75t_L g1731 ( 
.A(n_1713),
.Y(n_1731)
);

INVx1_ASAP7_75t_L g1732 ( 
.A(n_1713),
.Y(n_1732)
);

OR2x2_ASAP7_75t_L g1733 ( 
.A(n_1688),
.B(n_1675),
.Y(n_1733)
);

INVx2_ASAP7_75t_L g1734 ( 
.A(n_1698),
.Y(n_1734)
);

INVx2_ASAP7_75t_L g1735 ( 
.A(n_1698),
.Y(n_1735)
);

INVx1_ASAP7_75t_L g1736 ( 
.A(n_1693),
.Y(n_1736)
);

NOR2xp33_ASAP7_75t_L g1737 ( 
.A(n_1700),
.B(n_1651),
.Y(n_1737)
);

INVx1_ASAP7_75t_L g1738 ( 
.A(n_1693),
.Y(n_1738)
);

AND2x2_ASAP7_75t_L g1739 ( 
.A(n_1687),
.B(n_1670),
.Y(n_1739)
);

AND2x2_ASAP7_75t_L g1740 ( 
.A(n_1687),
.B(n_1692),
.Y(n_1740)
);

INVx1_ASAP7_75t_L g1741 ( 
.A(n_1699),
.Y(n_1741)
);

NOR2xp33_ASAP7_75t_L g1742 ( 
.A(n_1687),
.B(n_1651),
.Y(n_1742)
);

AND2x4_ASAP7_75t_L g1743 ( 
.A(n_1696),
.B(n_1658),
.Y(n_1743)
);

NAND2x1p5_ASAP7_75t_L g1744 ( 
.A(n_1696),
.B(n_1596),
.Y(n_1744)
);

AOI22xp33_ASAP7_75t_L g1745 ( 
.A1(n_1692),
.A2(n_1656),
.B1(n_1664),
.B2(n_1673),
.Y(n_1745)
);

AOI32xp33_ASAP7_75t_L g1746 ( 
.A1(n_1692),
.A2(n_1664),
.A3(n_1674),
.B1(n_1646),
.B2(n_1662),
.Y(n_1746)
);

INVx2_ASAP7_75t_L g1747 ( 
.A(n_1698),
.Y(n_1747)
);

INVx1_ASAP7_75t_L g1748 ( 
.A(n_1699),
.Y(n_1748)
);

NAND2xp5_ASAP7_75t_L g1749 ( 
.A(n_1696),
.B(n_1650),
.Y(n_1749)
);

OR2x2_ASAP7_75t_L g1750 ( 
.A(n_1691),
.B(n_1675),
.Y(n_1750)
);

INVx1_ASAP7_75t_L g1751 ( 
.A(n_1708),
.Y(n_1751)
);

NAND2x1p5_ASAP7_75t_L g1752 ( 
.A(n_1694),
.B(n_1596),
.Y(n_1752)
);

INVx1_ASAP7_75t_L g1753 ( 
.A(n_1708),
.Y(n_1753)
);

NAND2xp5_ASAP7_75t_L g1754 ( 
.A(n_1694),
.B(n_1650),
.Y(n_1754)
);

NAND2xp5_ASAP7_75t_L g1755 ( 
.A(n_1694),
.B(n_1649),
.Y(n_1755)
);

INVx2_ASAP7_75t_L g1756 ( 
.A(n_1695),
.Y(n_1756)
);

HB1xp67_ASAP7_75t_L g1757 ( 
.A(n_1695),
.Y(n_1757)
);

NAND2xp5_ASAP7_75t_L g1758 ( 
.A(n_1695),
.B(n_1649),
.Y(n_1758)
);

NAND2xp5_ASAP7_75t_L g1759 ( 
.A(n_1737),
.B(n_1670),
.Y(n_1759)
);

AND2x2_ASAP7_75t_L g1760 ( 
.A(n_1740),
.B(n_1702),
.Y(n_1760)
);

OA21x2_ASAP7_75t_L g1761 ( 
.A1(n_1724),
.A2(n_1709),
.B(n_1682),
.Y(n_1761)
);

AND2x4_ASAP7_75t_L g1762 ( 
.A(n_1740),
.B(n_1702),
.Y(n_1762)
);

INVx1_ASAP7_75t_L g1763 ( 
.A(n_1751),
.Y(n_1763)
);

AND2x2_ASAP7_75t_L g1764 ( 
.A(n_1718),
.B(n_1702),
.Y(n_1764)
);

NOR2xp33_ASAP7_75t_L g1765 ( 
.A(n_1724),
.B(n_1580),
.Y(n_1765)
);

AND2x2_ASAP7_75t_L g1766 ( 
.A(n_1718),
.B(n_1702),
.Y(n_1766)
);

NOR3xp33_ASAP7_75t_SL g1767 ( 
.A(n_1729),
.B(n_1674),
.C(n_1673),
.Y(n_1767)
);

OR2x2_ASAP7_75t_L g1768 ( 
.A(n_1726),
.B(n_1701),
.Y(n_1768)
);

INVx1_ASAP7_75t_SL g1769 ( 
.A(n_1718),
.Y(n_1769)
);

NAND2xp5_ASAP7_75t_L g1770 ( 
.A(n_1742),
.B(n_1670),
.Y(n_1770)
);

INVx1_ASAP7_75t_L g1771 ( 
.A(n_1753),
.Y(n_1771)
);

NOR3xp33_ASAP7_75t_L g1772 ( 
.A(n_1746),
.B(n_1609),
.C(n_1576),
.Y(n_1772)
);

AND2x2_ASAP7_75t_L g1773 ( 
.A(n_1717),
.B(n_1702),
.Y(n_1773)
);

AND2x2_ASAP7_75t_L g1774 ( 
.A(n_1717),
.B(n_1702),
.Y(n_1774)
);

AND2x2_ASAP7_75t_L g1775 ( 
.A(n_1756),
.B(n_1757),
.Y(n_1775)
);

OR2x2_ASAP7_75t_L g1776 ( 
.A(n_1726),
.B(n_1701),
.Y(n_1776)
);

AND2x2_ASAP7_75t_L g1777 ( 
.A(n_1756),
.B(n_1686),
.Y(n_1777)
);

INVx1_ASAP7_75t_SL g1778 ( 
.A(n_1749),
.Y(n_1778)
);

NAND2xp5_ASAP7_75t_L g1779 ( 
.A(n_1745),
.B(n_1725),
.Y(n_1779)
);

NAND2xp5_ASAP7_75t_L g1780 ( 
.A(n_1754),
.B(n_1662),
.Y(n_1780)
);

OAI21x1_ASAP7_75t_L g1781 ( 
.A1(n_1720),
.A2(n_1671),
.B(n_1683),
.Y(n_1781)
);

INVx2_ASAP7_75t_SL g1782 ( 
.A(n_1723),
.Y(n_1782)
);

INVx1_ASAP7_75t_L g1783 ( 
.A(n_1736),
.Y(n_1783)
);

CKINVDCx20_ASAP7_75t_R g1784 ( 
.A(n_1755),
.Y(n_1784)
);

OR2x2_ASAP7_75t_L g1785 ( 
.A(n_1719),
.B(n_1701),
.Y(n_1785)
);

OR2x2_ASAP7_75t_L g1786 ( 
.A(n_1719),
.B(n_1691),
.Y(n_1786)
);

INVx2_ASAP7_75t_SL g1787 ( 
.A(n_1723),
.Y(n_1787)
);

BUFx3_ASAP7_75t_L g1788 ( 
.A(n_1716),
.Y(n_1788)
);

AND2x2_ASAP7_75t_L g1789 ( 
.A(n_1728),
.B(n_1686),
.Y(n_1789)
);

NAND2xp5_ASAP7_75t_L g1790 ( 
.A(n_1731),
.B(n_1662),
.Y(n_1790)
);

HB1xp67_ASAP7_75t_L g1791 ( 
.A(n_1721),
.Y(n_1791)
);

OR2x2_ASAP7_75t_L g1792 ( 
.A(n_1722),
.B(n_1660),
.Y(n_1792)
);

OR2x2_ASAP7_75t_L g1793 ( 
.A(n_1727),
.B(n_1660),
.Y(n_1793)
);

OR2x2_ASAP7_75t_L g1794 ( 
.A(n_1732),
.B(n_1660),
.Y(n_1794)
);

OAI22xp33_ASAP7_75t_L g1795 ( 
.A1(n_1779),
.A2(n_1720),
.B1(n_1608),
.B2(n_1733),
.Y(n_1795)
);

INVx1_ASAP7_75t_L g1796 ( 
.A(n_1763),
.Y(n_1796)
);

BUFx3_ASAP7_75t_L g1797 ( 
.A(n_1788),
.Y(n_1797)
);

NAND2xp5_ASAP7_75t_L g1798 ( 
.A(n_1767),
.B(n_1738),
.Y(n_1798)
);

OAI22xp33_ASAP7_75t_L g1799 ( 
.A1(n_1778),
.A2(n_1608),
.B1(n_1733),
.B2(n_1617),
.Y(n_1799)
);

AOI22xp5_ASAP7_75t_L g1800 ( 
.A1(n_1772),
.A2(n_1784),
.B1(n_1765),
.B2(n_1761),
.Y(n_1800)
);

O2A1O1Ixp33_ASAP7_75t_L g1801 ( 
.A1(n_1791),
.A2(n_1741),
.B(n_1748),
.C(n_1654),
.Y(n_1801)
);

INVx1_ASAP7_75t_L g1802 ( 
.A(n_1763),
.Y(n_1802)
);

OAI321xp33_ASAP7_75t_L g1803 ( 
.A1(n_1775),
.A2(n_1752),
.A3(n_1744),
.B1(n_1734),
.B2(n_1747),
.C(n_1735),
.Y(n_1803)
);

INVx1_ASAP7_75t_L g1804 ( 
.A(n_1771),
.Y(n_1804)
);

O2A1O1Ixp33_ASAP7_75t_L g1805 ( 
.A1(n_1761),
.A2(n_1654),
.B(n_1752),
.C(n_1758),
.Y(n_1805)
);

INVx1_ASAP7_75t_L g1806 ( 
.A(n_1771),
.Y(n_1806)
);

INVxp67_ASAP7_75t_SL g1807 ( 
.A(n_1761),
.Y(n_1807)
);

AOI22xp33_ASAP7_75t_SL g1808 ( 
.A1(n_1761),
.A2(n_1728),
.B1(n_1730),
.B2(n_1739),
.Y(n_1808)
);

AND2x2_ASAP7_75t_L g1809 ( 
.A(n_1764),
.B(n_1730),
.Y(n_1809)
);

NOR2xp33_ASAP7_75t_L g1810 ( 
.A(n_1769),
.B(n_1606),
.Y(n_1810)
);

OAI22xp5_ASAP7_75t_L g1811 ( 
.A1(n_1769),
.A2(n_1679),
.B1(n_1663),
.B2(n_1646),
.Y(n_1811)
);

NAND3xp33_ASAP7_75t_L g1812 ( 
.A(n_1788),
.B(n_1735),
.C(n_1734),
.Y(n_1812)
);

AOI211x1_ASAP7_75t_SL g1813 ( 
.A1(n_1780),
.A2(n_1747),
.B(n_1715),
.C(n_1712),
.Y(n_1813)
);

AND2x2_ASAP7_75t_L g1814 ( 
.A(n_1764),
.B(n_1739),
.Y(n_1814)
);

INVx1_ASAP7_75t_SL g1815 ( 
.A(n_1775),
.Y(n_1815)
);

NAND2xp5_ASAP7_75t_L g1816 ( 
.A(n_1788),
.B(n_1743),
.Y(n_1816)
);

NAND2xp5_ASAP7_75t_L g1817 ( 
.A(n_1782),
.B(n_1743),
.Y(n_1817)
);

INVx1_ASAP7_75t_L g1818 ( 
.A(n_1783),
.Y(n_1818)
);

OAI22xp5_ASAP7_75t_L g1819 ( 
.A1(n_1759),
.A2(n_1679),
.B1(n_1663),
.B2(n_1646),
.Y(n_1819)
);

NAND4xp25_ASAP7_75t_L g1820 ( 
.A(n_1783),
.B(n_1750),
.C(n_1636),
.D(n_1608),
.Y(n_1820)
);

AOI311xp33_ASAP7_75t_L g1821 ( 
.A1(n_1790),
.A2(n_1677),
.A3(n_1678),
.B(n_1672),
.C(n_1709),
.Y(n_1821)
);

INVx1_ASAP7_75t_L g1822 ( 
.A(n_1807),
.Y(n_1822)
);

OAI221xp5_ASAP7_75t_SL g1823 ( 
.A1(n_1800),
.A2(n_1770),
.B1(n_1786),
.B2(n_1773),
.C(n_1774),
.Y(n_1823)
);

INVxp67_ASAP7_75t_L g1824 ( 
.A(n_1810),
.Y(n_1824)
);

AND2x2_ASAP7_75t_L g1825 ( 
.A(n_1809),
.B(n_1782),
.Y(n_1825)
);

NAND4xp25_ASAP7_75t_L g1826 ( 
.A(n_1798),
.B(n_1760),
.C(n_1762),
.D(n_1766),
.Y(n_1826)
);

INVxp67_ASAP7_75t_SL g1827 ( 
.A(n_1797),
.Y(n_1827)
);

INVx1_ASAP7_75t_L g1828 ( 
.A(n_1807),
.Y(n_1828)
);

INVx1_ASAP7_75t_L g1829 ( 
.A(n_1796),
.Y(n_1829)
);

AOI21xp33_ASAP7_75t_L g1830 ( 
.A1(n_1810),
.A2(n_1787),
.B(n_1792),
.Y(n_1830)
);

INVx1_ASAP7_75t_L g1831 ( 
.A(n_1802),
.Y(n_1831)
);

INVx1_ASAP7_75t_L g1832 ( 
.A(n_1804),
.Y(n_1832)
);

HB1xp67_ASAP7_75t_L g1833 ( 
.A(n_1815),
.Y(n_1833)
);

INVx1_ASAP7_75t_SL g1834 ( 
.A(n_1816),
.Y(n_1834)
);

INVx1_ASAP7_75t_L g1835 ( 
.A(n_1806),
.Y(n_1835)
);

AOI321xp33_ASAP7_75t_L g1836 ( 
.A1(n_1803),
.A2(n_1762),
.A3(n_1760),
.B1(n_1774),
.B2(n_1773),
.C(n_1766),
.Y(n_1836)
);

AOI22xp33_ASAP7_75t_L g1837 ( 
.A1(n_1819),
.A2(n_1762),
.B1(n_1777),
.B2(n_1787),
.Y(n_1837)
);

HB1xp67_ASAP7_75t_L g1838 ( 
.A(n_1812),
.Y(n_1838)
);

INVxp67_ASAP7_75t_L g1839 ( 
.A(n_1817),
.Y(n_1839)
);

AOI21xp5_ASAP7_75t_L g1840 ( 
.A1(n_1801),
.A2(n_1781),
.B(n_1762),
.Y(n_1840)
);

AND2x2_ASAP7_75t_L g1841 ( 
.A(n_1814),
.B(n_1808),
.Y(n_1841)
);

OR2x2_ASAP7_75t_L g1842 ( 
.A(n_1811),
.B(n_1792),
.Y(n_1842)
);

INVx1_ASAP7_75t_L g1843 ( 
.A(n_1833),
.Y(n_1843)
);

AND2x2_ASAP7_75t_L g1844 ( 
.A(n_1825),
.B(n_1789),
.Y(n_1844)
);

A2O1A1Ixp33_ASAP7_75t_L g1845 ( 
.A1(n_1836),
.A2(n_1805),
.B(n_1820),
.C(n_1781),
.Y(n_1845)
);

NAND2xp5_ASAP7_75t_L g1846 ( 
.A(n_1827),
.B(n_1818),
.Y(n_1846)
);

NAND3xp33_ASAP7_75t_SL g1847 ( 
.A(n_1838),
.B(n_1813),
.C(n_1752),
.Y(n_1847)
);

OAI221xp5_ASAP7_75t_L g1848 ( 
.A1(n_1823),
.A2(n_1821),
.B1(n_1786),
.B2(n_1793),
.C(n_1794),
.Y(n_1848)
);

INVxp67_ASAP7_75t_L g1849 ( 
.A(n_1825),
.Y(n_1849)
);

INVx2_ASAP7_75t_L g1850 ( 
.A(n_1822),
.Y(n_1850)
);

AOI32xp33_ASAP7_75t_L g1851 ( 
.A1(n_1841),
.A2(n_1795),
.A3(n_1799),
.B1(n_1777),
.B2(n_1789),
.Y(n_1851)
);

OAI21xp33_ASAP7_75t_L g1852 ( 
.A1(n_1830),
.A2(n_1795),
.B(n_1799),
.Y(n_1852)
);

XNOR2x1_ASAP7_75t_L g1853 ( 
.A(n_1834),
.B(n_1841),
.Y(n_1853)
);

INVx1_ASAP7_75t_L g1854 ( 
.A(n_1822),
.Y(n_1854)
);

INVx1_ASAP7_75t_SL g1855 ( 
.A(n_1842),
.Y(n_1855)
);

NAND2xp5_ASAP7_75t_L g1856 ( 
.A(n_1824),
.B(n_1839),
.Y(n_1856)
);

INVxp67_ASAP7_75t_L g1857 ( 
.A(n_1853),
.Y(n_1857)
);

INVx2_ASAP7_75t_L g1858 ( 
.A(n_1844),
.Y(n_1858)
);

INVx1_ASAP7_75t_L g1859 ( 
.A(n_1850),
.Y(n_1859)
);

AO22x2_ASAP7_75t_L g1860 ( 
.A1(n_1855),
.A2(n_1828),
.B1(n_1832),
.B2(n_1829),
.Y(n_1860)
);

AND2x2_ASAP7_75t_L g1861 ( 
.A(n_1849),
.B(n_1837),
.Y(n_1861)
);

AND2x2_ASAP7_75t_L g1862 ( 
.A(n_1843),
.B(n_1842),
.Y(n_1862)
);

NAND2xp5_ASAP7_75t_L g1863 ( 
.A(n_1846),
.B(n_1828),
.Y(n_1863)
);

NAND2xp5_ASAP7_75t_L g1864 ( 
.A(n_1856),
.B(n_1826),
.Y(n_1864)
);

OR2x2_ASAP7_75t_L g1865 ( 
.A(n_1848),
.B(n_1831),
.Y(n_1865)
);

NOR2xp33_ASAP7_75t_L g1866 ( 
.A(n_1852),
.B(n_1829),
.Y(n_1866)
);

AOI22xp33_ASAP7_75t_L g1867 ( 
.A1(n_1852),
.A2(n_1840),
.B1(n_1835),
.B2(n_1832),
.Y(n_1867)
);

NAND4xp25_ASAP7_75t_L g1868 ( 
.A(n_1857),
.B(n_1845),
.C(n_1851),
.D(n_1854),
.Y(n_1868)
);

AOI211x1_ASAP7_75t_SL g1869 ( 
.A1(n_1864),
.A2(n_1847),
.B(n_1835),
.C(n_1715),
.Y(n_1869)
);

AOI222xp33_ASAP7_75t_L g1870 ( 
.A1(n_1866),
.A2(n_1743),
.B1(n_1659),
.B2(n_1704),
.C1(n_1629),
.C2(n_1672),
.Y(n_1870)
);

INVx1_ASAP7_75t_L g1871 ( 
.A(n_1860),
.Y(n_1871)
);

NOR4xp25_ASAP7_75t_L g1872 ( 
.A(n_1867),
.B(n_1776),
.C(n_1768),
.D(n_1785),
.Y(n_1872)
);

NOR2x1p5_ASAP7_75t_L g1873 ( 
.A(n_1858),
.B(n_1863),
.Y(n_1873)
);

NOR4xp25_ASAP7_75t_SL g1874 ( 
.A(n_1871),
.B(n_1859),
.C(n_1860),
.D(n_1862),
.Y(n_1874)
);

A2O1A1Ixp33_ASAP7_75t_L g1875 ( 
.A1(n_1868),
.A2(n_1865),
.B(n_1861),
.C(n_1859),
.Y(n_1875)
);

NAND4xp25_ASAP7_75t_L g1876 ( 
.A(n_1869),
.B(n_1564),
.C(n_1785),
.D(n_1776),
.Y(n_1876)
);

AOI322xp5_ASAP7_75t_L g1877 ( 
.A1(n_1872),
.A2(n_1659),
.A3(n_1689),
.B1(n_1686),
.B2(n_1710),
.C1(n_1706),
.C2(n_1703),
.Y(n_1877)
);

OAI22xp5_ASAP7_75t_L g1878 ( 
.A1(n_1873),
.A2(n_1793),
.B1(n_1794),
.B2(n_1744),
.Y(n_1878)
);

AOI221xp5_ASAP7_75t_L g1879 ( 
.A1(n_1870),
.A2(n_1768),
.B1(n_1704),
.B2(n_1744),
.C(n_1750),
.Y(n_1879)
);

O2A1O1Ixp33_ASAP7_75t_L g1880 ( 
.A1(n_1871),
.A2(n_1564),
.B(n_1704),
.C(n_1667),
.Y(n_1880)
);

INVx1_ASAP7_75t_L g1881 ( 
.A(n_1875),
.Y(n_1881)
);

INVx2_ASAP7_75t_L g1882 ( 
.A(n_1878),
.Y(n_1882)
);

NOR2x1_ASAP7_75t_L g1883 ( 
.A(n_1874),
.B(n_1564),
.Y(n_1883)
);

NAND2xp33_ASAP7_75t_L g1884 ( 
.A(n_1879),
.B(n_1564),
.Y(n_1884)
);

INVx1_ASAP7_75t_L g1885 ( 
.A(n_1876),
.Y(n_1885)
);

NOR2xp67_ASAP7_75t_L g1886 ( 
.A(n_1880),
.B(n_1593),
.Y(n_1886)
);

NAND2xp5_ASAP7_75t_L g1887 ( 
.A(n_1883),
.B(n_1877),
.Y(n_1887)
);

NAND2xp5_ASAP7_75t_L g1888 ( 
.A(n_1881),
.B(n_1704),
.Y(n_1888)
);

NOR2x1p5_ASAP7_75t_L g1889 ( 
.A(n_1882),
.B(n_1593),
.Y(n_1889)
);

INVxp67_ASAP7_75t_SL g1890 ( 
.A(n_1889),
.Y(n_1890)
);

INVx2_ASAP7_75t_L g1891 ( 
.A(n_1890),
.Y(n_1891)
);

INVx2_ASAP7_75t_L g1892 ( 
.A(n_1891),
.Y(n_1892)
);

XNOR2xp5_ASAP7_75t_L g1893 ( 
.A(n_1891),
.B(n_1885),
.Y(n_1893)
);

AOI21xp33_ASAP7_75t_SL g1894 ( 
.A1(n_1893),
.A2(n_1887),
.B(n_1888),
.Y(n_1894)
);

OAI22x1_ASAP7_75t_L g1895 ( 
.A1(n_1892),
.A2(n_1884),
.B1(n_1886),
.B2(n_1593),
.Y(n_1895)
);

AO21x2_ASAP7_75t_L g1896 ( 
.A1(n_1894),
.A2(n_1715),
.B(n_1712),
.Y(n_1896)
);

OAI21xp33_ASAP7_75t_L g1897 ( 
.A1(n_1895),
.A2(n_1704),
.B(n_1566),
.Y(n_1897)
);

AOI22xp33_ASAP7_75t_SL g1898 ( 
.A1(n_1896),
.A2(n_1704),
.B1(n_1683),
.B2(n_1566),
.Y(n_1898)
);

O2A1O1Ixp5_ASAP7_75t_SL g1899 ( 
.A1(n_1898),
.A2(n_1897),
.B(n_1683),
.C(n_1711),
.Y(n_1899)
);

HB1xp67_ASAP7_75t_L g1900 ( 
.A(n_1899),
.Y(n_1900)
);

AOI221xp5_ASAP7_75t_L g1901 ( 
.A1(n_1900),
.A2(n_1709),
.B1(n_1711),
.B2(n_1682),
.C(n_1714),
.Y(n_1901)
);

AOI211xp5_ASAP7_75t_L g1902 ( 
.A1(n_1901),
.A2(n_1559),
.B(n_1554),
.C(n_1549),
.Y(n_1902)
);


endmodule