module fake_jpeg_24161_n_41 (n_3, n_2, n_1, n_0, n_4, n_5, n_41);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_41;

wire n_13;
wire n_21;
wire n_33;
wire n_10;
wire n_23;
wire n_27;
wire n_6;
wire n_22;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_34;
wire n_30;
wire n_39;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_31;
wire n_25;
wire n_29;
wire n_37;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

CKINVDCx20_ASAP7_75t_R g6 ( 
.A(n_1),
.Y(n_6)
);

BUFx6f_ASAP7_75t_L g7 ( 
.A(n_1),
.Y(n_7)
);

INVx8_ASAP7_75t_L g8 ( 
.A(n_5),
.Y(n_8)
);

BUFx3_ASAP7_75t_L g9 ( 
.A(n_2),
.Y(n_9)
);

INVx2_ASAP7_75t_SL g10 ( 
.A(n_3),
.Y(n_10)
);

BUFx6f_ASAP7_75t_L g11 ( 
.A(n_0),
.Y(n_11)
);

NOR2xp33_ASAP7_75t_L g12 ( 
.A(n_4),
.B(n_5),
.Y(n_12)
);

AND2x2_ASAP7_75t_L g13 ( 
.A(n_3),
.B(n_0),
.Y(n_13)
);

O2A1O1Ixp33_ASAP7_75t_L g14 ( 
.A1(n_9),
.A2(n_0),
.B(n_1),
.C(n_2),
.Y(n_14)
);

AOI21xp5_ASAP7_75t_L g24 ( 
.A1(n_14),
.A2(n_17),
.B(n_10),
.Y(n_24)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_9),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_15),
.B(n_19),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g16 ( 
.A(n_13),
.B(n_4),
.Y(n_16)
);

AND2x2_ASAP7_75t_L g26 ( 
.A(n_16),
.B(n_8),
.Y(n_26)
);

A2O1A1Ixp33_ASAP7_75t_L g17 ( 
.A1(n_13),
.A2(n_12),
.B(n_6),
.C(n_11),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_6),
.B(n_10),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_SL g25 ( 
.A(n_18),
.B(n_21),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_20),
.Y(n_22)
);

INVxp67_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_19),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_23),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_24),
.Y(n_29)
);

XNOR2xp5_ASAP7_75t_SL g30 ( 
.A(n_26),
.B(n_17),
.Y(n_30)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_30),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_28),
.B(n_22),
.Y(n_31)
);

MAJIxp5_ASAP7_75t_L g34 ( 
.A(n_31),
.B(n_30),
.C(n_25),
.Y(n_34)
);

INVxp67_ASAP7_75t_L g33 ( 
.A(n_29),
.Y(n_33)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_33),
.Y(n_36)
);

MAJIxp5_ASAP7_75t_L g37 ( 
.A(n_34),
.B(n_35),
.C(n_32),
.Y(n_37)
);

AOI21xp5_ASAP7_75t_L g35 ( 
.A1(n_33),
.A2(n_25),
.B(n_27),
.Y(n_35)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_37),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_L g38 ( 
.A1(n_36),
.A2(n_14),
.B1(n_8),
.B2(n_19),
.Y(n_38)
);

AOI21xp5_ASAP7_75t_L g40 ( 
.A1(n_39),
.A2(n_38),
.B(n_7),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_40),
.B(n_11),
.Y(n_41)
);


endmodule