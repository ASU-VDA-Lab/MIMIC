module real_jpeg_29557_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_313, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_313;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_163;
wire n_22;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_13;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_80;
wire n_30;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_16;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_100;
wire n_51;
wire n_14;
wire n_205;
wire n_261;
wire n_86;
wire n_70;
wire n_32;
wire n_228;
wire n_15;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_0),
.B(n_47),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_0),
.B(n_110),
.Y(n_109)
);

INVx11_ASAP7_75t_L g142 ( 
.A(n_0),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_0),
.B(n_206),
.Y(n_211)
);

BUFx12_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_2),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_L g29 ( 
.A1(n_3),
.A2(n_4),
.B1(n_20),
.B2(n_30),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_3),
.Y(n_30)
);

OAI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_3),
.A2(n_24),
.B1(n_25),
.B2(n_30),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_3),
.A2(n_30),
.B1(n_45),
.B2(n_47),
.Y(n_110)
);

OAI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_3),
.A2(n_30),
.B1(n_39),
.B2(n_43),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g19 ( 
.A1(n_4),
.A2(n_6),
.B1(n_20),
.B2(n_21),
.Y(n_19)
);

INVx13_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_4),
.A2(n_5),
.B1(n_20),
.B2(n_119),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_5),
.Y(n_119)
);

OAI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_5),
.A2(n_24),
.B1(n_25),
.B2(n_119),
.Y(n_123)
);

OAI22xp33_ASAP7_75t_SL g176 ( 
.A1(n_5),
.A2(n_39),
.B1(n_43),
.B2(n_119),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_5),
.A2(n_45),
.B1(n_47),
.B2(n_119),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_6),
.Y(n_21)
);

AOI22xp33_ASAP7_75t_L g79 ( 
.A1(n_6),
.A2(n_21),
.B1(n_24),
.B2(n_25),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_6),
.A2(n_21),
.B1(n_45),
.B2(n_47),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g248 ( 
.A1(n_6),
.A2(n_21),
.B1(n_39),
.B2(n_43),
.Y(n_248)
);

INVx11_ASAP7_75t_L g41 ( 
.A(n_7),
.Y(n_41)
);

AOI21xp33_ASAP7_75t_L g196 ( 
.A1(n_7),
.A2(n_10),
.B(n_45),
.Y(n_196)
);

BUFx24_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_9),
.Y(n_56)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_9),
.Y(n_63)
);

AOI21xp33_ASAP7_75t_SL g166 ( 
.A1(n_9),
.A2(n_10),
.B(n_39),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_10),
.A2(n_39),
.B1(n_43),
.B2(n_51),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_10),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_10),
.A2(n_24),
.B1(n_25),
.B2(n_51),
.Y(n_59)
);

AOI21xp5_ASAP7_75t_L g73 ( 
.A1(n_10),
.A2(n_20),
.B(n_74),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_10),
.B(n_20),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_10),
.B(n_69),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_10),
.A2(n_45),
.B1(n_47),
.B2(n_51),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_10),
.B(n_55),
.Y(n_200)
);

INVx11_ASAP7_75t_SL g46 ( 
.A(n_11),
.Y(n_46)
);

XOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_97),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_SL g13 ( 
.A(n_14),
.B(n_95),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_SL g14 ( 
.A(n_15),
.B(n_82),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_15),
.B(n_82),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_67),
.C(n_75),
.Y(n_15)
);

OAI22xp5_ASAP7_75t_SL g305 ( 
.A1(n_16),
.A2(n_17),
.B1(n_67),
.B2(n_300),
.Y(n_305)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_17),
.Y(n_16)
);

AOI22xp5_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_33),
.B1(n_34),
.B2(n_66),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_18),
.Y(n_66)
);

OAI21xp5_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_22),
.B(n_27),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_19),
.Y(n_87)
);

A2O1A1Ixp33_ASAP7_75t_L g31 ( 
.A1(n_20),
.A2(n_22),
.B(n_23),
.C(n_32),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_20),
.B(n_23),
.Y(n_32)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_22),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_22),
.B(n_118),
.Y(n_117)
);

AOI21xp5_ASAP7_75t_L g293 ( 
.A1(n_22),
.A2(n_31),
.B(n_73),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_24),
.B1(n_25),
.B2(n_26),
.Y(n_22)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_23),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_24),
.B(n_26),
.Y(n_136)
);

INVx8_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

O2A1O1Ixp33_ASAP7_75t_L g62 ( 
.A1(n_25),
.A2(n_55),
.B(n_63),
.C(n_64),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_25),
.B(n_63),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_25),
.A2(n_136),
.B1(n_137),
.B2(n_138),
.Y(n_135)
);

A2O1A1Ixp33_ASAP7_75t_L g165 ( 
.A1(n_25),
.A2(n_51),
.B(n_56),
.C(n_166),
.Y(n_165)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_28),
.B(n_117),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_31),
.Y(n_28)
);

CKINVDCx16_ASAP7_75t_R g70 ( 
.A(n_29),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_SL g72 ( 
.A(n_31),
.B(n_73),
.Y(n_72)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_31),
.Y(n_86)
);

CKINVDCx16_ASAP7_75t_R g138 ( 
.A(n_32),
.Y(n_138)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

XOR2xp5_ASAP7_75t_L g34 ( 
.A(n_35),
.B(n_52),
.Y(n_34)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_35),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_35),
.B(n_52),
.C(n_66),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_35),
.A2(n_76),
.B1(n_120),
.B2(n_121),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_SL g302 ( 
.A(n_35),
.B(n_77),
.Y(n_302)
);

AOI21xp5_ASAP7_75t_SL g35 ( 
.A1(n_36),
.A2(n_48),
.B(n_49),
.Y(n_35)
);

OAI21xp5_ASAP7_75t_SL g274 ( 
.A1(n_36),
.A2(n_112),
.B(n_248),
.Y(n_274)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_37),
.B(n_50),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_37),
.B(n_113),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_37),
.B(n_176),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_38),
.B(n_44),
.Y(n_37)
);

AOI22xp33_ASAP7_75t_L g38 ( 
.A1(n_39),
.A2(n_41),
.B1(n_42),
.B2(n_43),
.Y(n_38)
);

INVx4_ASAP7_75t_SL g43 ( 
.A(n_39),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_L g55 ( 
.A1(n_39),
.A2(n_43),
.B1(n_56),
.B2(n_57),
.Y(n_55)
);

A2O1A1Ixp33_ASAP7_75t_L g195 ( 
.A1(n_39),
.A2(n_41),
.B(n_51),
.C(n_196),
.Y(n_195)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx11_ASAP7_75t_L g42 ( 
.A(n_41),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_SL g44 ( 
.A1(n_41),
.A2(n_42),
.B1(n_45),
.B2(n_47),
.Y(n_44)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_44),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_44),
.B(n_113),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_44),
.B(n_176),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_44),
.B(n_50),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_45),
.Y(n_47)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_47),
.B(n_221),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_SL g216 ( 
.A(n_48),
.B(n_51),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_L g247 ( 
.A1(n_48),
.A2(n_177),
.B(n_248),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_50),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_51),
.B(n_222),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_53),
.B(n_60),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_53),
.B(n_132),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_54),
.B(n_58),
.Y(n_53)
);

AOI21xp5_ASAP7_75t_L g89 ( 
.A1(n_54),
.A2(n_58),
.B(n_90),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_SL g285 ( 
.A1(n_54),
.A2(n_61),
.B(n_79),
.Y(n_285)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_55),
.B(n_65),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_55),
.B(n_123),
.Y(n_122)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_56),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_59),
.B(n_62),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_61),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_61),
.B(n_122),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_62),
.B(n_65),
.Y(n_61)
);

AOI21xp5_ASAP7_75t_L g77 ( 
.A1(n_62),
.A2(n_78),
.B(n_80),
.Y(n_77)
);

INVxp67_ASAP7_75t_L g90 ( 
.A(n_62),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_62),
.B(n_123),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g75 ( 
.A(n_67),
.B(n_76),
.C(n_77),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g299 ( 
.A1(n_67),
.A2(n_300),
.B1(n_301),
.B2(n_302),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g300 ( 
.A(n_67),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_68),
.B(n_71),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_68),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_68),
.B(n_128),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_69),
.B(n_70),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g267 ( 
.A(n_69),
.B(n_268),
.Y(n_267)
);

INVxp67_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_72),
.B(n_117),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_73),
.Y(n_268)
);

INVxp67_ASAP7_75t_L g137 ( 
.A(n_74),
.Y(n_137)
);

XOR2xp5_ASAP7_75t_L g304 ( 
.A(n_75),
.B(n_305),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_76),
.B(n_116),
.C(n_120),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_79),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_80),
.B(n_271),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_81),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_81),
.B(n_133),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_83),
.A2(n_92),
.B1(n_93),
.B2(n_94),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_83),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_84),
.A2(n_85),
.B1(n_89),
.B2(n_91),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_85),
.Y(n_84)
);

AOI21xp5_ASAP7_75t_L g85 ( 
.A1(n_86),
.A2(n_87),
.B(n_88),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_86),
.B(n_129),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_89),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_89),
.A2(n_91),
.B1(n_252),
.B2(n_253),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_91),
.B(n_250),
.C(n_253),
.Y(n_276)
);

CKINVDCx16_ASAP7_75t_R g92 ( 
.A(n_93),
.Y(n_92)
);

INVxp67_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

OAI321xp33_ASAP7_75t_L g97 ( 
.A1(n_98),
.A2(n_297),
.A3(n_306),
.B1(n_309),
.B2(n_310),
.C(n_313),
.Y(n_97)
);

AOI21xp5_ASAP7_75t_L g98 ( 
.A1(n_99),
.A2(n_278),
.B(n_296),
.Y(n_98)
);

OAI21xp5_ASAP7_75t_SL g99 ( 
.A1(n_100),
.A2(n_257),
.B(n_277),
.Y(n_99)
);

O2A1O1Ixp33_ASAP7_75t_SL g100 ( 
.A1(n_101),
.A2(n_159),
.B(n_240),
.C(n_256),
.Y(n_100)
);

AND2x2_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_146),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_102),
.B(n_146),
.Y(n_239)
);

XOR2xp5_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_124),
.Y(n_102)
);

XOR2xp5_ASAP7_75t_L g103 ( 
.A(n_104),
.B(n_115),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_104),
.B(n_115),
.C(n_124),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g104 ( 
.A(n_105),
.B(n_111),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_105),
.B(n_111),
.Y(n_250)
);

OAI21xp5_ASAP7_75t_L g105 ( 
.A1(n_106),
.A2(n_108),
.B(n_109),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_SL g144 ( 
.A(n_106),
.B(n_145),
.Y(n_144)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_107),
.B(n_158),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_SL g168 ( 
.A1(n_107),
.A2(n_141),
.B(n_158),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g205 ( 
.A(n_107),
.B(n_206),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_L g139 ( 
.A1(n_108),
.A2(n_140),
.B(n_143),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_109),
.B(n_157),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_109),
.B(n_205),
.Y(n_217)
);

INVxp33_ASAP7_75t_L g145 ( 
.A(n_110),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_112),
.B(n_114),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_112),
.B(n_187),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_114),
.B(n_175),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g148 ( 
.A(n_116),
.B(n_149),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_118),
.Y(n_129)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_122),
.B(n_172),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_SL g124 ( 
.A(n_125),
.B(n_134),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_126),
.A2(n_127),
.B1(n_130),
.B2(n_131),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_126),
.B(n_131),
.C(n_134),
.Y(n_254)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_128),
.B(n_267),
.Y(n_266)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_133),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_135),
.B(n_139),
.Y(n_134)
);

XOR2xp5_ASAP7_75t_L g151 ( 
.A(n_135),
.B(n_139),
.Y(n_151)
);

INVx11_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g204 ( 
.A(n_141),
.B(n_158),
.Y(n_204)
);

INVx5_ASAP7_75t_SL g222 ( 
.A(n_141),
.Y(n_222)
);

INVx11_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_143),
.B(n_204),
.Y(n_246)
);

CKINVDCx16_ASAP7_75t_R g143 ( 
.A(n_144),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_144),
.B(n_210),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_150),
.C(n_152),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_147),
.A2(n_148),
.B1(n_235),
.B2(n_236),
.Y(n_234)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g236 ( 
.A1(n_150),
.A2(n_151),
.B1(n_152),
.B2(n_237),
.Y(n_236)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_152),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_154),
.C(n_156),
.Y(n_152)
);

XOR2xp5_ASAP7_75t_L g180 ( 
.A(n_153),
.B(n_181),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_154),
.A2(n_155),
.B1(n_156),
.B2(n_182),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_155),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_156),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_157),
.B(n_211),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_SL g159 ( 
.A(n_160),
.B(n_239),
.Y(n_159)
);

AOI21xp5_ASAP7_75t_L g160 ( 
.A1(n_161),
.A2(n_232),
.B(n_238),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_L g161 ( 
.A1(n_162),
.A2(n_189),
.B(n_231),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_178),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_163),
.B(n_178),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_164),
.B(n_170),
.C(n_173),
.Y(n_163)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_164),
.B(n_229),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_165),
.A2(n_167),
.B1(n_168),
.B2(n_169),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_165),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_165),
.B(n_168),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g273 ( 
.A1(n_167),
.A2(n_168),
.B1(n_274),
.B2(n_275),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_167),
.B(n_274),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_L g291 ( 
.A1(n_167),
.A2(n_168),
.B1(n_292),
.B2(n_293),
.Y(n_291)
);

CKINVDCx16_ASAP7_75t_R g167 ( 
.A(n_168),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_L g303 ( 
.A1(n_168),
.A2(n_288),
.B(n_293),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_170),
.A2(n_171),
.B1(n_173),
.B2(n_174),
.Y(n_229)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_172),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_174),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_175),
.B(n_177),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_177),
.B(n_186),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_179),
.A2(n_180),
.B1(n_183),
.B2(n_184),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_179),
.B(n_185),
.C(n_188),
.Y(n_233)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

XOR2xp5_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_188),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_187),
.Y(n_185)
);

AOI21xp5_ASAP7_75t_L g189 ( 
.A1(n_190),
.A2(n_226),
.B(n_230),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_L g190 ( 
.A1(n_191),
.A2(n_207),
.B(n_225),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_192),
.B(n_197),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g225 ( 
.A(n_192),
.B(n_197),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_SL g192 ( 
.A(n_193),
.B(n_195),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_193),
.A2(n_194),
.B1(n_195),
.B2(n_213),
.Y(n_212)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_195),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_203),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_199),
.A2(n_200),
.B1(n_201),
.B2(n_202),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_199),
.B(n_202),
.C(n_203),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_200),
.Y(n_199)
);

CKINVDCx16_ASAP7_75t_R g201 ( 
.A(n_202),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_204),
.B(n_205),
.Y(n_203)
);

AOI21xp5_ASAP7_75t_L g207 ( 
.A1(n_208),
.A2(n_214),
.B(n_224),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_209),
.B(n_212),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_SL g224 ( 
.A(n_209),
.B(n_212),
.Y(n_224)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

OAI21xp5_ASAP7_75t_SL g214 ( 
.A1(n_215),
.A2(n_218),
.B(n_223),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_216),
.B(n_217),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_SL g223 ( 
.A(n_216),
.B(n_217),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_219),
.B(n_220),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_227),
.B(n_228),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_SL g230 ( 
.A(n_227),
.B(n_228),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_233),
.B(n_234),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_SL g238 ( 
.A(n_233),
.B(n_234),
.Y(n_238)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_241),
.B(n_242),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_SL g256 ( 
.A(n_241),
.B(n_242),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_243),
.A2(n_244),
.B1(n_254),
.B2(n_255),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_245),
.B(n_249),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_245),
.B(n_249),
.C(n_255),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_246),
.B(n_247),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_246),
.B(n_247),
.Y(n_263)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_250),
.B(n_251),
.Y(n_249)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_254),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_258),
.B(n_259),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_SL g277 ( 
.A(n_258),
.B(n_259),
.Y(n_277)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_260),
.B(n_276),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_261),
.A2(n_262),
.B1(n_272),
.B2(n_273),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_261),
.B(n_273),
.C(n_276),
.Y(n_279)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

XOR2xp5_ASAP7_75t_L g262 ( 
.A(n_263),
.B(n_264),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_263),
.B(n_265),
.C(n_270),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_265),
.A2(n_266),
.B1(n_269),
.B2(n_270),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_266),
.Y(n_265)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_273),
.Y(n_272)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_274),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_279),
.B(n_280),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_SL g296 ( 
.A(n_279),
.B(n_280),
.Y(n_296)
);

AOI22xp33_ASAP7_75t_SL g280 ( 
.A1(n_281),
.A2(n_282),
.B1(n_294),
.B2(n_295),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

XOR2xp5_ASAP7_75t_L g282 ( 
.A(n_283),
.B(n_287),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_283),
.B(n_287),
.C(n_295),
.Y(n_307)
);

AOI21xp5_ASAP7_75t_L g283 ( 
.A1(n_284),
.A2(n_285),
.B(n_286),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_284),
.B(n_285),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_286),
.B(n_299),
.C(n_303),
.Y(n_298)
);

FAx1_ASAP7_75t_SL g308 ( 
.A(n_286),
.B(n_299),
.CI(n_303),
.CON(n_308),
.SN(n_308)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_288),
.A2(n_289),
.B1(n_290),
.B2(n_291),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_289),
.Y(n_288)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g292 ( 
.A(n_293),
.Y(n_292)
);

CKINVDCx16_ASAP7_75t_R g295 ( 
.A(n_294),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_298),
.B(n_304),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_298),
.B(n_304),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g301 ( 
.A(n_302),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_307),
.B(n_308),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_SL g309 ( 
.A(n_307),
.B(n_308),
.Y(n_309)
);

BUFx24_ASAP7_75t_SL g312 ( 
.A(n_308),
.Y(n_312)
);


endmodule