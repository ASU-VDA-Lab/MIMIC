module fake_jpeg_12729_n_362 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_362);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_362;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx2_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

CKINVDCx16_ASAP7_75t_R g19 ( 
.A(n_9),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_6),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_14),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_3),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

INVx13_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_11),
.Y(n_33)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_16),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_11),
.Y(n_35)
);

BUFx5_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_5),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_15),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_2),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_10),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_15),
.Y(n_41)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_13),
.Y(n_42)
);

INVx11_ASAP7_75t_SL g43 ( 
.A(n_9),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_39),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_44),
.Y(n_80)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_29),
.Y(n_45)
);

HB1xp67_ASAP7_75t_L g122 ( 
.A(n_45),
.Y(n_122)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_29),
.Y(n_46)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_46),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_39),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_47),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_39),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_48),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_26),
.B(n_9),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_49),
.B(n_72),
.Y(n_119)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_29),
.Y(n_50)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_50),
.Y(n_111)
);

AND2x2_ASAP7_75t_L g51 ( 
.A(n_17),
.B(n_8),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_51),
.B(n_71),
.Y(n_94)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_36),
.Y(n_52)
);

INVx5_ASAP7_75t_L g77 ( 
.A(n_52),
.Y(n_77)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_36),
.Y(n_53)
);

INVx5_ASAP7_75t_L g112 ( 
.A(n_53),
.Y(n_112)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_34),
.Y(n_54)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_54),
.Y(n_113)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_23),
.Y(n_55)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_55),
.Y(n_96)
);

BUFx5_ASAP7_75t_L g56 ( 
.A(n_18),
.Y(n_56)
);

BUFx12f_ASAP7_75t_L g110 ( 
.A(n_56),
.Y(n_110)
);

INVx2_ASAP7_75t_SL g57 ( 
.A(n_34),
.Y(n_57)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_57),
.Y(n_95)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_34),
.Y(n_58)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_58),
.Y(n_82)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_22),
.Y(n_59)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_59),
.Y(n_104)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_18),
.Y(n_60)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_60),
.Y(n_115)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_22),
.Y(n_61)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_61),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_18),
.Y(n_62)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_62),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_20),
.Y(n_63)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_63),
.Y(n_87)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_23),
.Y(n_64)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_64),
.Y(n_108)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_20),
.Y(n_65)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_65),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_20),
.Y(n_66)
);

BUFx10_ASAP7_75t_L g86 ( 
.A(n_66),
.Y(n_86)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_22),
.Y(n_67)
);

BUFx4f_ASAP7_75t_SL g83 ( 
.A(n_67),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_25),
.Y(n_68)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_68),
.B(n_69),
.Y(n_97)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_17),
.Y(n_69)
);

INVx13_ASAP7_75t_L g70 ( 
.A(n_32),
.Y(n_70)
);

INVx6_ASAP7_75t_SL g98 ( 
.A(n_70),
.Y(n_98)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_25),
.Y(n_71)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_42),
.Y(n_72)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_42),
.Y(n_73)
);

OR2x2_ASAP7_75t_L g100 ( 
.A(n_73),
.B(n_41),
.Y(n_100)
);

BUFx3_ASAP7_75t_L g74 ( 
.A(n_25),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_74),
.B(n_75),
.Y(n_102)
);

BUFx12f_ASAP7_75t_L g75 ( 
.A(n_30),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_24),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_76),
.B(n_38),
.Y(n_103)
);

INVx11_ASAP7_75t_L g78 ( 
.A(n_70),
.Y(n_78)
);

INVxp67_ASAP7_75t_L g138 ( 
.A(n_78),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_51),
.B(n_31),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_79),
.B(n_88),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_57),
.A2(n_43),
.B1(n_24),
.B2(n_35),
.Y(n_81)
);

OAI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_81),
.A2(n_21),
.B1(n_19),
.B2(n_40),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_SL g84 ( 
.A(n_52),
.B(n_37),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_SL g145 ( 
.A(n_84),
.B(n_85),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_60),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_65),
.B(n_35),
.Y(n_88)
);

OR2x2_ASAP7_75t_SL g89 ( 
.A(n_52),
.B(n_32),
.Y(n_89)
);

AND2x2_ASAP7_75t_L g152 ( 
.A(n_89),
.B(n_100),
.Y(n_152)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_53),
.A2(n_41),
.B1(n_33),
.B2(n_30),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g132 ( 
.A1(n_92),
.A2(n_105),
.B1(n_0),
.B2(n_1),
.Y(n_132)
);

INVx11_ASAP7_75t_L g93 ( 
.A(n_75),
.Y(n_93)
);

CKINVDCx16_ASAP7_75t_R g143 ( 
.A(n_93),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_75),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_101),
.B(n_103),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_44),
.A2(n_41),
.B1(n_33),
.B2(n_30),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_SL g107 ( 
.A(n_62),
.B(n_38),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_107),
.B(n_114),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_47),
.B(n_31),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_109),
.B(n_0),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_63),
.B(n_37),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_66),
.B(n_27),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_117),
.B(n_118),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_68),
.B(n_28),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_48),
.B(n_28),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_121),
.B(n_112),
.Y(n_163)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_108),
.Y(n_123)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_123),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_125),
.A2(n_127),
.B1(n_129),
.B2(n_135),
.Y(n_167)
);

INVx2_ASAP7_75t_SL g126 ( 
.A(n_98),
.Y(n_126)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_126),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_100),
.A2(n_33),
.B1(n_40),
.B2(n_27),
.Y(n_127)
);

INVx6_ASAP7_75t_L g128 ( 
.A(n_80),
.Y(n_128)
);

INVx6_ASAP7_75t_L g182 ( 
.A(n_128),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_119),
.A2(n_26),
.B1(n_19),
.B2(n_21),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_L g130 ( 
.A1(n_97),
.A2(n_32),
.B1(n_1),
.B2(n_2),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_130),
.A2(n_132),
.B1(n_140),
.B2(n_149),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_98),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_131),
.B(n_157),
.Y(n_195)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_120),
.Y(n_133)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_133),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_88),
.A2(n_8),
.B1(n_15),
.B2(n_14),
.Y(n_135)
);

INVx6_ASAP7_75t_L g136 ( 
.A(n_80),
.Y(n_136)
);

INVx3_ASAP7_75t_L g170 ( 
.A(n_136),
.Y(n_170)
);

INVx4_ASAP7_75t_L g137 ( 
.A(n_93),
.Y(n_137)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_137),
.Y(n_187)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_96),
.Y(n_139)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_139),
.Y(n_175)
);

AOI22xp33_ASAP7_75t_L g140 ( 
.A1(n_97),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_140)
);

AND2x2_ASAP7_75t_SL g174 ( 
.A(n_141),
.B(n_104),
.Y(n_174)
);

HB1xp67_ASAP7_75t_L g142 ( 
.A(n_95),
.Y(n_142)
);

CKINVDCx16_ASAP7_75t_R g197 ( 
.A(n_142),
.Y(n_197)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_96),
.Y(n_144)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_144),
.Y(n_190)
);

HB1xp67_ASAP7_75t_L g146 ( 
.A(n_95),
.Y(n_146)
);

CKINVDCx16_ASAP7_75t_R g199 ( 
.A(n_146),
.Y(n_199)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_116),
.Y(n_148)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_148),
.Y(n_196)
);

OAI22xp33_ASAP7_75t_SL g149 ( 
.A1(n_81),
.A2(n_12),
.B1(n_4),
.B2(n_7),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_109),
.B(n_1),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_150),
.B(n_151),
.Y(n_165)
);

AO22x2_ASAP7_75t_L g151 ( 
.A1(n_89),
.A2(n_4),
.B1(n_7),
.B2(n_8),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_SL g153 ( 
.A1(n_122),
.A2(n_4),
.B1(n_7),
.B2(n_12),
.Y(n_153)
);

INVxp67_ASAP7_75t_L g181 ( 
.A(n_153),
.Y(n_181)
);

BUFx12_ASAP7_75t_L g154 ( 
.A(n_78),
.Y(n_154)
);

CKINVDCx14_ASAP7_75t_R g171 ( 
.A(n_154),
.Y(n_171)
);

AOI22xp33_ASAP7_75t_SL g155 ( 
.A1(n_99),
.A2(n_13),
.B1(n_14),
.B2(n_16),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_SL g189 ( 
.A1(n_155),
.A2(n_158),
.B1(n_110),
.B2(n_86),
.Y(n_189)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_116),
.Y(n_156)
);

BUFx3_ASAP7_75t_L g186 ( 
.A(n_156),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_86),
.Y(n_157)
);

AOI22xp33_ASAP7_75t_SL g158 ( 
.A1(n_99),
.A2(n_13),
.B1(n_111),
.B2(n_112),
.Y(n_158)
);

INVx4_ASAP7_75t_L g159 ( 
.A(n_77),
.Y(n_159)
);

CKINVDCx16_ASAP7_75t_R g200 ( 
.A(n_159),
.Y(n_200)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_87),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_161),
.Y(n_173)
);

AND2x2_ASAP7_75t_L g162 ( 
.A(n_94),
.B(n_79),
.Y(n_162)
);

XOR2xp5_ASAP7_75t_SL g176 ( 
.A(n_162),
.B(n_152),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_163),
.B(n_102),
.Y(n_179)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_104),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_164),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_174),
.B(n_180),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_176),
.B(n_177),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_124),
.B(n_162),
.C(n_152),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_124),
.A2(n_90),
.B1(n_91),
.B2(n_115),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_178),
.A2(n_194),
.B1(n_139),
.B2(n_143),
.Y(n_216)
);

NAND3xp33_ASAP7_75t_L g218 ( 
.A(n_179),
.B(n_198),
.C(n_154),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_162),
.B(n_97),
.C(n_106),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_SL g183 ( 
.A(n_147),
.B(n_145),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_SL g203 ( 
.A(n_183),
.B(n_138),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_152),
.B(n_141),
.C(n_150),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_184),
.B(n_144),
.Y(n_215)
);

AOI21xp5_ASAP7_75t_L g185 ( 
.A1(n_131),
.A2(n_77),
.B(n_111),
.Y(n_185)
);

AOI21xp5_ASAP7_75t_L g205 ( 
.A1(n_185),
.A2(n_126),
.B(n_138),
.Y(n_205)
);

INVxp67_ASAP7_75t_L g210 ( 
.A(n_189),
.Y(n_210)
);

XOR2xp5_ASAP7_75t_L g191 ( 
.A(n_160),
.B(n_115),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_191),
.B(n_151),
.Y(n_209)
);

AOI22xp33_ASAP7_75t_L g192 ( 
.A1(n_127),
.A2(n_91),
.B1(n_90),
.B2(n_86),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_L g227 ( 
.A1(n_192),
.A2(n_201),
.B1(n_185),
.B2(n_171),
.Y(n_227)
);

AOI22xp33_ASAP7_75t_SL g193 ( 
.A1(n_129),
.A2(n_113),
.B1(n_106),
.B2(n_82),
.Y(n_193)
);

CKINVDCx16_ASAP7_75t_R g221 ( 
.A(n_193),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_123),
.A2(n_86),
.B1(n_82),
.B2(n_113),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_SL g198 ( 
.A(n_134),
.B(n_83),
.Y(n_198)
);

AOI22xp33_ASAP7_75t_SL g201 ( 
.A1(n_164),
.A2(n_83),
.B1(n_110),
.B2(n_161),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_172),
.Y(n_202)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_202),
.Y(n_236)
);

OR2x2_ASAP7_75t_L g239 ( 
.A(n_203),
.B(n_207),
.Y(n_239)
);

INVx4_ASAP7_75t_L g204 ( 
.A(n_170),
.Y(n_204)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_204),
.Y(n_249)
);

A2O1A1Ixp33_ASAP7_75t_SL g260 ( 
.A1(n_205),
.A2(n_227),
.B(n_224),
.C(n_212),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_183),
.B(n_133),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_206),
.B(n_213),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_SL g207 ( 
.A(n_177),
.B(n_151),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_172),
.Y(n_208)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_208),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_SL g241 ( 
.A(n_209),
.B(n_194),
.Y(n_241)
);

INVx3_ASAP7_75t_L g211 ( 
.A(n_170),
.Y(n_211)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_211),
.Y(n_246)
);

OAI21xp5_ASAP7_75t_SL g212 ( 
.A1(n_165),
.A2(n_151),
.B(n_126),
.Y(n_212)
);

INVxp67_ASAP7_75t_L g235 ( 
.A(n_212),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_165),
.B(n_151),
.Y(n_213)
);

INVx5_ASAP7_75t_L g214 ( 
.A(n_182),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_214),
.B(n_215),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_L g237 ( 
.A1(n_216),
.A2(n_223),
.B1(n_224),
.B2(n_234),
.Y(n_237)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_175),
.Y(n_217)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_217),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_218),
.B(n_228),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_169),
.B(n_156),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_219),
.B(n_226),
.Y(n_252)
);

OAI21xp33_ASAP7_75t_L g220 ( 
.A1(n_176),
.A2(n_154),
.B(n_148),
.Y(n_220)
);

AND2x2_ASAP7_75t_L g257 ( 
.A(n_220),
.B(n_227),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_178),
.A2(n_128),
.B1(n_136),
.B2(n_159),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_174),
.A2(n_137),
.B1(n_83),
.B2(n_110),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_167),
.A2(n_184),
.B1(n_180),
.B2(n_181),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_225),
.A2(n_190),
.B1(n_196),
.B2(n_173),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_169),
.B(n_191),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_195),
.B(n_198),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_174),
.B(n_166),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_229),
.B(n_230),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_166),
.B(n_197),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_188),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_232),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_188),
.Y(n_233)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_233),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_SL g234 ( 
.A(n_167),
.B(n_168),
.Y(n_234)
);

AND2x6_ASAP7_75t_L g240 ( 
.A(n_225),
.B(n_181),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_240),
.B(n_251),
.Y(n_276)
);

XOR2xp5_ASAP7_75t_L g281 ( 
.A(n_241),
.B(n_243),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_231),
.B(n_199),
.C(n_175),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_242),
.B(n_244),
.C(n_259),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_231),
.B(n_190),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_L g245 ( 
.A1(n_234),
.A2(n_210),
.B1(n_221),
.B2(n_216),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_L g266 ( 
.A1(n_245),
.A2(n_256),
.B1(n_205),
.B2(n_230),
.Y(n_266)
);

A2O1A1O1Ixp25_ASAP7_75t_L g250 ( 
.A1(n_209),
.A2(n_196),
.B(n_173),
.C(n_200),
.D(n_187),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_SL g268 ( 
.A(n_250),
.B(n_219),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_213),
.A2(n_182),
.B1(n_186),
.B2(n_187),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_253),
.A2(n_255),
.B1(n_237),
.B2(n_257),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_222),
.A2(n_186),
.B1(n_207),
.B2(n_229),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_L g256 ( 
.A1(n_221),
.A2(n_206),
.B1(n_223),
.B2(n_203),
.Y(n_256)
);

XOR2x2_ASAP7_75t_L g259 ( 
.A(n_222),
.B(n_226),
.Y(n_259)
);

AOI21xp5_ASAP7_75t_SL g280 ( 
.A1(n_260),
.A2(n_243),
.B(n_239),
.Y(n_280)
);

OAI21xp5_ASAP7_75t_L g263 ( 
.A1(n_235),
.A2(n_257),
.B(n_239),
.Y(n_263)
);

INVxp67_ASAP7_75t_L g289 ( 
.A(n_263),
.Y(n_289)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_262),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_265),
.B(n_267),
.Y(n_286)
);

CKINVDCx14_ASAP7_75t_R g294 ( 
.A(n_266),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_235),
.A2(n_233),
.B1(n_232),
.B2(n_208),
.Y(n_267)
);

CKINVDCx14_ASAP7_75t_R g301 ( 
.A(n_268),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_244),
.B(n_202),
.C(n_217),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_269),
.B(n_273),
.C(n_249),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_254),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_270),
.B(n_271),
.Y(n_295)
);

INVxp67_ASAP7_75t_L g271 ( 
.A(n_257),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_236),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_272),
.B(n_274),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_259),
.B(n_211),
.C(n_204),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_261),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_261),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_275),
.B(n_282),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_276),
.B(n_277),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_SL g277 ( 
.A(n_247),
.B(n_214),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_SL g278 ( 
.A(n_248),
.B(n_252),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_278),
.B(n_283),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_SL g298 ( 
.A(n_279),
.B(n_284),
.Y(n_298)
);

OAI21xp5_ASAP7_75t_L g292 ( 
.A1(n_280),
.A2(n_260),
.B(n_250),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_L g282 ( 
.A1(n_260),
.A2(n_248),
.B1(n_241),
.B2(n_240),
.Y(n_282)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_238),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_258),
.Y(n_284)
);

XOR2xp5_ASAP7_75t_L g285 ( 
.A(n_264),
.B(n_255),
.Y(n_285)
);

XOR2xp5_ASAP7_75t_L g308 ( 
.A(n_285),
.B(n_290),
.Y(n_308)
);

CKINVDCx16_ASAP7_75t_R g287 ( 
.A(n_263),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_SL g312 ( 
.A(n_287),
.B(n_291),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_279),
.A2(n_260),
.B1(n_252),
.B2(n_242),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_L g306 ( 
.A1(n_288),
.A2(n_281),
.B1(n_271),
.B2(n_273),
.Y(n_306)
);

XOR2xp5_ASAP7_75t_L g290 ( 
.A(n_264),
.B(n_253),
.Y(n_290)
);

CKINVDCx16_ASAP7_75t_R g291 ( 
.A(n_270),
.Y(n_291)
);

AOI21xp5_ASAP7_75t_L g314 ( 
.A1(n_292),
.A2(n_265),
.B(n_272),
.Y(n_314)
);

XOR2xp5_ASAP7_75t_L g293 ( 
.A(n_269),
.B(n_246),
.Y(n_293)
);

XOR2xp5_ASAP7_75t_L g316 ( 
.A(n_293),
.B(n_283),
.Y(n_316)
);

XOR2xp5_ASAP7_75t_SL g296 ( 
.A(n_282),
.B(n_249),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_L g311 ( 
.A(n_296),
.B(n_267),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_303),
.B(n_290),
.C(n_293),
.Y(n_317)
);

OAI22xp5_ASAP7_75t_L g304 ( 
.A1(n_301),
.A2(n_294),
.B1(n_300),
.B2(n_275),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_L g320 ( 
.A1(n_304),
.A2(n_309),
.B1(n_310),
.B2(n_287),
.Y(n_320)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_295),
.Y(n_305)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_305),
.Y(n_321)
);

INVxp67_ASAP7_75t_L g325 ( 
.A(n_306),
.Y(n_325)
);

BUFx2_ASAP7_75t_L g307 ( 
.A(n_295),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_307),
.B(n_313),
.Y(n_327)
);

OAI22xp5_ASAP7_75t_L g309 ( 
.A1(n_299),
.A2(n_274),
.B1(n_298),
.B2(n_276),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_SL g310 ( 
.A1(n_298),
.A2(n_280),
.B1(n_278),
.B2(n_281),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_L g328 ( 
.A(n_311),
.B(n_314),
.Y(n_328)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_302),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_L g315 ( 
.A(n_285),
.B(n_284),
.Y(n_315)
);

XOR2xp5_ASAP7_75t_L g323 ( 
.A(n_315),
.B(n_316),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_317),
.B(n_319),
.C(n_296),
.Y(n_326)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_297),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_318),
.B(n_297),
.Y(n_322)
);

XOR2xp5_ASAP7_75t_L g319 ( 
.A(n_303),
.B(n_288),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_320),
.B(n_324),
.Y(n_333)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_322),
.Y(n_341)
);

AOI22xp5_ASAP7_75t_L g324 ( 
.A1(n_310),
.A2(n_299),
.B1(n_292),
.B2(n_289),
.Y(n_324)
);

XNOR2xp5_ASAP7_75t_L g336 ( 
.A(n_326),
.B(n_312),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_316),
.B(n_291),
.Y(n_329)
);

OAI21xp5_ASAP7_75t_L g337 ( 
.A1(n_329),
.A2(n_330),
.B(n_331),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_SL g330 ( 
.A(n_317),
.B(n_289),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_315),
.B(n_286),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_326),
.B(n_319),
.C(n_308),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_332),
.B(n_334),
.Y(n_342)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_325),
.B(n_308),
.C(n_306),
.Y(n_334)
);

XOR2xp5_ASAP7_75t_L g335 ( 
.A(n_323),
.B(n_311),
.Y(n_335)
);

XOR2xp5_ASAP7_75t_L g347 ( 
.A(n_335),
.B(n_336),
.Y(n_347)
);

XNOR2x1_ASAP7_75t_L g338 ( 
.A(n_328),
.B(n_314),
.Y(n_338)
);

AND2x2_ASAP7_75t_L g343 ( 
.A(n_338),
.B(n_339),
.Y(n_343)
);

XOR2xp5_ASAP7_75t_L g339 ( 
.A(n_323),
.B(n_286),
.Y(n_339)
);

FAx1_ASAP7_75t_SL g340 ( 
.A(n_324),
.B(n_328),
.CI(n_327),
.CON(n_340),
.SN(n_340)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_340),
.B(n_325),
.Y(n_345)
);

INVx11_ASAP7_75t_L g344 ( 
.A(n_341),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_SL g350 ( 
.A(n_344),
.B(n_348),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_SL g352 ( 
.A(n_345),
.B(n_346),
.Y(n_352)
);

INVx3_ASAP7_75t_L g346 ( 
.A(n_337),
.Y(n_346)
);

NOR2xp33_ASAP7_75t_L g348 ( 
.A(n_340),
.B(n_321),
.Y(n_348)
);

AOI21xp5_ASAP7_75t_L g349 ( 
.A1(n_336),
.A2(n_307),
.B(n_333),
.Y(n_349)
);

OAI22xp5_ASAP7_75t_L g353 ( 
.A1(n_349),
.A2(n_334),
.B1(n_338),
.B2(n_332),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_L g351 ( 
.A(n_342),
.B(n_339),
.Y(n_351)
);

NOR2xp33_ASAP7_75t_L g355 ( 
.A(n_351),
.B(n_354),
.Y(n_355)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_353),
.Y(n_357)
);

NOR2xp33_ASAP7_75t_L g354 ( 
.A(n_346),
.B(n_335),
.Y(n_354)
);

NOR2xp33_ASAP7_75t_L g356 ( 
.A(n_350),
.B(n_344),
.Y(n_356)
);

MAJIxp5_ASAP7_75t_L g358 ( 
.A(n_356),
.B(n_352),
.C(n_347),
.Y(n_358)
);

MAJIxp5_ASAP7_75t_L g359 ( 
.A(n_358),
.B(n_357),
.C(n_355),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_SL g360 ( 
.A(n_359),
.B(n_357),
.Y(n_360)
);

AOI21xp5_ASAP7_75t_L g361 ( 
.A1(n_360),
.A2(n_350),
.B(n_343),
.Y(n_361)
);

NOR2xp33_ASAP7_75t_L g362 ( 
.A(n_361),
.B(n_343),
.Y(n_362)
);


endmodule