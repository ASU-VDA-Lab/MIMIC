module fake_netlist_5_1070_n_1686 (n_137, n_91, n_82, n_122, n_142, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_60, n_152, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_125, n_35, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_29, n_79, n_131, n_151, n_47, n_25, n_53, n_8, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_85, n_95, n_119, n_59, n_26, n_133, n_55, n_99, n_2, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_12, n_67, n_121, n_36, n_76, n_87, n_150, n_27, n_64, n_77, n_102, n_106, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_134, n_32, n_41, n_104, n_103, n_56, n_51, n_63, n_97, n_141, n_11, n_153, n_7, n_15, n_145, n_48, n_50, n_52, n_88, n_110, n_1686);

input n_137;
input n_91;
input n_82;
input n_122;
input n_142;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_60;
input n_152;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_125;
input n_35;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_29;
input n_79;
input n_131;
input n_151;
input n_47;
input n_25;
input n_53;
input n_8;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_85;
input n_95;
input n_119;
input n_59;
input n_26;
input n_133;
input n_55;
input n_99;
input n_2;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_150;
input n_27;
input n_64;
input n_77;
input n_102;
input n_106;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_134;
input n_32;
input n_41;
input n_104;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_11;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_1686;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1166;
wire n_469;
wire n_1508;
wire n_785;
wire n_549;
wire n_532;
wire n_1161;
wire n_1677;
wire n_1150;
wire n_226;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_1501;
wire n_880;
wire n_544;
wire n_1007;
wire n_155;
wire n_552;
wire n_1528;
wire n_1370;
wire n_1292;
wire n_1198;
wire n_1360;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1021;
wire n_551;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1353;
wire n_800;
wire n_1347;
wire n_1535;
wire n_1666;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_915;
wire n_1545;
wire n_864;
wire n_173;
wire n_859;
wire n_951;
wire n_1264;
wire n_447;
wire n_247;
wire n_1494;
wire n_292;
wire n_625;
wire n_854;
wire n_1462;
wire n_1580;
wire n_674;
wire n_417;
wire n_516;
wire n_933;
wire n_1152;
wire n_497;
wire n_1607;
wire n_1563;
wire n_606;
wire n_275;
wire n_877;
wire n_755;
wire n_1118;
wire n_947;
wire n_1285;
wire n_373;
wire n_307;
wire n_1359;
wire n_530;
wire n_1107;
wire n_556;
wire n_1230;
wire n_668;
wire n_375;
wire n_301;
wire n_929;
wire n_1124;
wire n_902;
wire n_1576;
wire n_191;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1257;
wire n_171;
wire n_1182;
wire n_579;
wire n_1261;
wire n_938;
wire n_1098;
wire n_320;
wire n_1154;
wire n_1242;
wire n_1135;
wire n_406;
wire n_519;
wire n_1016;
wire n_1243;
wire n_546;
wire n_1280;
wire n_281;
wire n_240;
wire n_291;
wire n_231;
wire n_257;
wire n_731;
wire n_371;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_317;
wire n_1236;
wire n_1633;
wire n_569;
wire n_227;
wire n_920;
wire n_1289;
wire n_1517;
wire n_335;
wire n_1669;
wire n_370;
wire n_976;
wire n_343;
wire n_1449;
wire n_308;
wire n_1566;
wire n_297;
wire n_156;
wire n_1078;
wire n_1670;
wire n_775;
wire n_219;
wire n_157;
wire n_600;
wire n_1484;
wire n_1374;
wire n_1328;
wire n_223;
wire n_264;
wire n_1598;
wire n_955;
wire n_163;
wire n_339;
wire n_1146;
wire n_882;
wire n_183;
wire n_243;
wire n_1036;
wire n_1097;
wire n_347;
wire n_550;
wire n_696;
wire n_897;
wire n_215;
wire n_350;
wire n_196;
wire n_798;
wire n_646;
wire n_1428;
wire n_436;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_290;
wire n_580;
wire n_1040;
wire n_578;
wire n_926;
wire n_344;
wire n_1218;
wire n_422;
wire n_475;
wire n_777;
wire n_1070;
wire n_1547;
wire n_1030;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_1561;
wire n_496;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_1600;
wire n_521;
wire n_663;
wire n_845;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_680;
wire n_1473;
wire n_1587;
wire n_395;
wire n_164;
wire n_553;
wire n_901;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_214;
wire n_1672;
wire n_675;
wire n_888;
wire n_1167;
wire n_1626;
wire n_637;
wire n_1384;
wire n_1556;
wire n_184;
wire n_446;
wire n_1064;
wire n_858;
wire n_923;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_468;
wire n_213;
wire n_342;
wire n_464;
wire n_363;
wire n_1582;
wire n_197;
wire n_1069;
wire n_1075;
wire n_1450;
wire n_1322;
wire n_1471;
wire n_1459;
wire n_460;
wire n_889;
wire n_973;
wire n_477;
wire n_571;
wire n_1585;
wire n_461;
wire n_1599;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_907;
wire n_1447;
wire n_1377;
wire n_190;
wire n_989;
wire n_1039;
wire n_228;
wire n_283;
wire n_1403;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_1002;
wire n_1463;
wire n_1581;
wire n_310;
wire n_593;
wire n_748;
wire n_586;
wire n_1058;
wire n_1667;
wire n_838;
wire n_332;
wire n_1053;
wire n_1224;
wire n_349;
wire n_1248;
wire n_230;
wire n_1331;
wire n_953;
wire n_279;
wire n_1014;
wire n_1241;
wire n_289;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_440;
wire n_793;
wire n_478;
wire n_476;
wire n_1527;
wire n_534;
wire n_884;
wire n_345;
wire n_944;
wire n_1623;
wire n_1565;
wire n_182;
wire n_647;
wire n_237;
wire n_407;
wire n_1072;
wire n_832;
wire n_857;
wire n_207;
wire n_561;
wire n_1319;
wire n_1387;
wire n_1532;
wire n_1027;
wire n_971;
wire n_1156;
wire n_326;
wire n_794;
wire n_404;
wire n_686;
wire n_847;
wire n_1393;
wire n_596;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_728;
wire n_266;
wire n_1162;
wire n_272;
wire n_1538;
wire n_1199;
wire n_352;
wire n_1038;
wire n_520;
wire n_1369;
wire n_409;
wire n_1660;
wire n_887;
wire n_300;
wire n_809;
wire n_870;
wire n_931;
wire n_599;
wire n_1662;
wire n_1481;
wire n_434;
wire n_1544;
wire n_868;
wire n_639;
wire n_914;
wire n_411;
wire n_414;
wire n_1629;
wire n_1293;
wire n_965;
wire n_935;
wire n_1175;
wire n_817;
wire n_360;
wire n_1479;
wire n_759;
wire n_806;
wire n_1477;
wire n_324;
wire n_1635;
wire n_1571;
wire n_187;
wire n_1189;
wire n_1259;
wire n_706;
wire n_746;
wire n_1649;
wire n_747;
wire n_784;
wire n_1244;
wire n_431;
wire n_1194;
wire n_615;
wire n_851;
wire n_843;
wire n_523;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_1679;
wire n_776;
wire n_1415;
wire n_367;
wire n_452;
wire n_525;
wire n_1260;
wire n_1647;
wire n_1464;
wire n_649;
wire n_547;
wire n_1444;
wire n_1191;
wire n_1674;
wire n_284;
wire n_1128;
wire n_744;
wire n_590;
wire n_629;
wire n_1308;
wire n_254;
wire n_1680;
wire n_1233;
wire n_1615;
wire n_1529;
wire n_526;
wire n_372;
wire n_293;
wire n_677;
wire n_244;
wire n_1333;
wire n_1121;
wire n_314;
wire n_368;
wire n_433;
wire n_604;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_1001;
wire n_1503;
wire n_498;
wire n_1468;
wire n_1559;
wire n_689;
wire n_738;
wire n_1624;
wire n_640;
wire n_1510;
wire n_252;
wire n_624;
wire n_1380;
wire n_1617;
wire n_295;
wire n_1010;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_1195;
wire n_610;
wire n_936;
wire n_568;
wire n_1500;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_448;
wire n_259;
wire n_758;
wire n_999;
wire n_1656;
wire n_1158;
wire n_1509;
wire n_563;
wire n_1145;
wire n_878;
wire n_524;
wire n_394;
wire n_204;
wire n_1678;
wire n_1049;
wire n_1153;
wire n_741;
wire n_1639;
wire n_1306;
wire n_1068;
wire n_331;
wire n_906;
wire n_1163;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_658;
wire n_1362;
wire n_1586;
wire n_456;
wire n_959;
wire n_535;
wire n_940;
wire n_1445;
wire n_1492;
wire n_592;
wire n_1169;
wire n_1596;
wire n_1017;
wire n_978;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_1095;
wire n_1614;
wire n_267;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_603;
wire n_1431;
wire n_484;
wire n_1593;
wire n_1033;
wire n_442;
wire n_636;
wire n_660;
wire n_1640;
wire n_1009;
wire n_1148;
wire n_742;
wire n_750;
wire n_995;
wire n_454;
wire n_1609;
wire n_374;
wire n_185;
wire n_396;
wire n_1383;
wire n_1073;
wire n_255;
wire n_662;
wire n_459;
wire n_218;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1065;
wire n_1592;
wire n_1336;
wire n_1574;
wire n_473;
wire n_1309;
wire n_1426;
wire n_1043;
wire n_355;
wire n_486;
wire n_1548;
wire n_614;
wire n_337;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_168;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_208;
wire n_743;
wire n_299;
wire n_303;
wire n_296;
wire n_613;
wire n_1119;
wire n_1240;
wire n_829;
wire n_1612;
wire n_1416;
wire n_361;
wire n_700;
wire n_1237;
wire n_573;
wire n_1420;
wire n_1132;
wire n_388;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_761;
wire n_1568;
wire n_1006;
wire n_329;
wire n_274;
wire n_1270;
wire n_1664;
wire n_1486;
wire n_582;
wire n_1332;
wire n_1390;
wire n_309;
wire n_512;
wire n_1591;
wire n_322;
wire n_1682;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1349;
wire n_1093;
wire n_288;
wire n_1031;
wire n_263;
wire n_609;
wire n_1041;
wire n_1265;
wire n_224;
wire n_1562;
wire n_383;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_239;
wire n_630;
wire n_504;
wire n_511;
wire n_874;
wire n_358;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_1304;
wire n_1324;
wire n_987;
wire n_261;
wire n_174;
wire n_1455;
wire n_767;
wire n_993;
wire n_1407;
wire n_1551;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_429;
wire n_948;
wire n_1217;
wire n_628;
wire n_365;
wire n_729;
wire n_1131;
wire n_1084;
wire n_970;
wire n_911;
wire n_1430;
wire n_513;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1534;
wire n_340;
wire n_1351;
wire n_1044;
wire n_1205;
wire n_346;
wire n_1209;
wire n_1552;
wire n_495;
wire n_602;
wire n_574;
wire n_1435;
wire n_879;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_1645;
wire n_490;
wire n_1327;
wire n_996;
wire n_921;
wire n_1684;
wire n_233;
wire n_572;
wire n_366;
wire n_815;
wire n_327;
wire n_1381;
wire n_1611;
wire n_1037;
wire n_1080;
wire n_1274;
wire n_1316;
wire n_426;
wire n_1438;
wire n_1082;
wire n_589;
wire n_716;
wire n_1630;
wire n_562;
wire n_1436;
wire n_952;
wire n_1229;
wire n_391;
wire n_701;
wire n_1437;
wire n_1023;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_238;
wire n_531;
wire n_890;
wire n_764;
wire n_1056;
wire n_1424;
wire n_162;
wire n_960;
wire n_222;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_634;
wire n_199;
wire n_1252;
wire n_348;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_1311;
wire n_1519;
wire n_256;
wire n_950;
wire n_1553;
wire n_380;
wire n_419;
wire n_1346;
wire n_444;
wire n_1299;
wire n_1060;
wire n_1141;
wire n_316;
wire n_389;
wire n_418;
wire n_248;
wire n_912;
wire n_315;
wire n_968;
wire n_451;
wire n_619;
wire n_408;
wire n_1386;
wire n_376;
wire n_967;
wire n_1442;
wire n_1139;
wire n_515;
wire n_351;
wire n_885;
wire n_397;
wire n_1432;
wire n_1357;
wire n_483;
wire n_683;
wire n_1632;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_1608;
wire n_983;
wire n_280;
wire n_1305;
wire n_873;
wire n_378;
wire n_1112;
wire n_762;
wire n_1283;
wire n_1644;
wire n_690;
wire n_583;
wire n_302;
wire n_1343;
wire n_1203;
wire n_1631;
wire n_821;
wire n_321;
wire n_1179;
wire n_621;
wire n_753;
wire n_455;
wire n_1048;
wire n_1288;
wire n_212;
wire n_385;
wire n_507;
wire n_1560;
wire n_1605;
wire n_330;
wire n_1228;
wire n_972;
wire n_692;
wire n_820;
wire n_1200;
wire n_1301;
wire n_1363;
wire n_1668;
wire n_1185;
wire n_991;
wire n_828;
wire n_779;
wire n_576;
wire n_1143;
wire n_1579;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_537;
wire n_945;
wire n_492;
wire n_1504;
wire n_943;
wire n_341;
wire n_250;
wire n_992;
wire n_543;
wire n_260;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_286;
wire n_1643;
wire n_883;
wire n_470;
wire n_325;
wire n_449;
wire n_1594;
wire n_1214;
wire n_1342;
wire n_1400;
wire n_900;
wire n_856;
wire n_918;
wire n_942;
wire n_189;
wire n_1147;
wire n_1557;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_540;
wire n_618;
wire n_896;
wire n_323;
wire n_195;
wire n_356;
wire n_894;
wire n_1636;
wire n_831;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1470;
wire n_1096;
wire n_234;
wire n_1575;
wire n_833;
wire n_1646;
wire n_225;
wire n_1307;
wire n_988;
wire n_814;
wire n_192;
wire n_1549;
wire n_1201;
wire n_1114;
wire n_655;
wire n_1616;
wire n_1446;
wire n_669;
wire n_472;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_387;
wire n_1149;
wire n_398;
wire n_1671;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_211;
wire n_1219;
wire n_1204;
wire n_178;
wire n_1035;
wire n_287;
wire n_555;
wire n_783;
wire n_1188;
wire n_661;
wire n_849;
wire n_336;
wire n_584;
wire n_681;
wire n_1638;
wire n_430;
wire n_510;
wire n_216;
wire n_311;
wire n_830;
wire n_1296;
wire n_1413;
wire n_801;
wire n_241;
wire n_875;
wire n_357;
wire n_1110;
wire n_1655;
wire n_445;
wire n_749;
wire n_1134;
wire n_1358;
wire n_717;
wire n_165;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_249;
wire n_304;
wire n_1338;
wire n_577;
wire n_1522;
wire n_1637;
wire n_1419;
wire n_338;
wire n_1653;
wire n_693;
wire n_1506;
wire n_836;
wire n_990;
wire n_1389;
wire n_975;
wire n_1256;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_306;
wire n_458;
wire n_770;
wire n_1375;
wire n_1102;
wire n_711;
wire n_1499;
wire n_1187;
wire n_1441;
wire n_1392;
wire n_1597;
wire n_1164;
wire n_1659;
wire n_489;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_1572;
wire n_876;
wire n_1516;
wire n_1190;
wire n_1685;
wire n_601;
wire n_917;
wire n_966;
wire n_253;
wire n_1116;
wire n_1661;
wire n_1212;
wire n_1541;
wire n_172;
wire n_206;
wire n_217;
wire n_726;
wire n_982;
wire n_1573;
wire n_1453;
wire n_818;
wire n_861;
wire n_1183;
wire n_1658;
wire n_899;
wire n_1253;
wire n_210;
wire n_774;
wire n_1628;
wire n_1335;
wire n_1514;
wire n_1059;
wire n_1345;
wire n_176;
wire n_1133;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_527;
wire n_1168;
wire n_707;
wire n_937;
wire n_1427;
wire n_393;
wire n_487;
wire n_1584;
wire n_665;
wire n_1440;
wire n_177;
wire n_421;
wire n_1356;
wire n_910;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1302;
wire n_205;
wire n_1136;
wire n_1313;
wire n_1491;
wire n_754;
wire n_1496;
wire n_179;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_735;
wire n_232;
wire n_1109;
wire n_895;
wire n_1310;
wire n_202;
wire n_427;
wire n_1399;
wire n_1543;
wire n_791;
wire n_732;
wire n_1533;
wire n_193;
wire n_808;
wire n_797;
wire n_1025;
wire n_500;
wire n_1067;
wire n_435;
wire n_159;
wire n_766;
wire n_1457;
wire n_541;
wire n_538;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_594;
wire n_200;
wire n_1291;
wire n_1297;
wire n_1155;
wire n_1418;
wire n_1524;
wire n_1485;
wire n_1011;
wire n_1184;
wire n_985;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_1352;
wire n_626;
wire n_1650;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_1170;
wire n_305;
wire n_676;
wire n_294;
wire n_318;
wire n_653;
wire n_642;
wire n_1602;
wire n_194;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_268;
wire n_664;
wire n_503;
wire n_235;
wire n_1372;
wire n_605;
wire n_1273;
wire n_353;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_1282;
wire n_1318;
wire n_780;
wire n_998;
wire n_1454;
wire n_467;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_501;
wire n_823;
wire n_245;
wire n_725;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_672;
wire n_581;
wire n_382;
wire n_554;
wire n_1625;
wire n_898;
wire n_1013;
wire n_1452;
wire n_718;
wire n_265;
wire n_1120;
wire n_719;
wire n_443;
wire n_198;
wire n_714;
wire n_1683;
wire n_909;
wire n_1497;
wire n_1530;
wire n_997;
wire n_932;
wire n_612;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_508;
wire n_506;
wire n_1320;
wire n_1663;
wire n_737;
wire n_986;
wire n_509;
wire n_1317;
wire n_1518;
wire n_1281;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_209;
wire n_1564;
wire n_1613;
wire n_733;
wire n_1489;
wire n_1376;
wire n_941;
wire n_981;
wire n_1569;
wire n_867;
wire n_186;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_298;
wire n_518;
wire n_505;
wire n_282;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1620;
wire n_381;
wire n_220;
wire n_390;
wire n_1330;
wire n_481;
wire n_1675;
wire n_1554;
wire n_769;
wire n_1046;
wire n_271;
wire n_934;
wire n_1618;
wire n_826;
wire n_886;
wire n_1221;
wire n_654;
wire n_1172;
wire n_167;
wire n_379;
wire n_428;
wire n_1341;
wire n_570;
wire n_1641;
wire n_1361;
wire n_853;
wire n_377;
wire n_751;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_392;
wire n_158;
wire n_704;
wire n_787;
wire n_961;
wire n_771;
wire n_276;
wire n_1225;
wire n_1520;
wire n_169;
wire n_522;
wire n_1287;
wire n_1262;
wire n_400;
wire n_930;
wire n_181;
wire n_1411;
wire n_221;
wire n_622;
wire n_1577;
wire n_1087;
wire n_386;
wire n_994;
wire n_848;
wire n_1550;
wire n_1498;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1567;
wire n_1247;
wire n_922;
wire n_816;
wire n_1648;
wire n_591;
wire n_1536;
wire n_1344;
wire n_313;
wire n_631;
wire n_479;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_432;
wire n_839;
wire n_1210;
wire n_1364;
wire n_328;
wire n_1250;
wire n_369;
wire n_871;
wire n_685;
wire n_598;
wire n_608;
wire n_928;
wire n_1367;
wire n_1460;
wire n_772;
wire n_1555;
wire n_499;
wire n_1589;
wire n_517;
wire n_402;
wire n_413;
wire n_1086;
wire n_796;
wire n_1619;
wire n_236;
wire n_1502;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_903;
wire n_1525;
wire n_740;
wire n_203;
wire n_384;
wire n_1404;
wire n_1315;
wire n_277;
wire n_1061;
wire n_333;
wire n_1298;
wire n_1652;
wire n_462;
wire n_1193;
wire n_1676;
wire n_1255;
wire n_258;
wire n_1113;
wire n_1226;
wire n_722;
wire n_1277;
wire n_188;
wire n_844;
wire n_201;
wire n_471;
wire n_852;
wire n_1487;
wire n_1028;
wire n_1601;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_1546;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_1627;
wire n_1245;
wire n_846;
wire n_1673;
wire n_465;
wire n_362;
wire n_1321;
wire n_170;
wire n_161;
wire n_273;
wire n_585;
wire n_270;
wire n_616;
wire n_745;
wire n_1654;
wire n_1103;
wire n_648;
wire n_1379;
wire n_312;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_494;
wire n_641;
wire n_730;
wire n_1325;
wire n_1595;
wire n_354;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_695;
wire n_180;
wire n_656;
wire n_1606;
wire n_1220;
wire n_1540;
wire n_229;
wire n_437;
wire n_1642;
wire n_403;
wire n_453;
wire n_1130;
wire n_720;
wire n_1526;
wire n_863;
wire n_805;
wire n_1604;
wire n_1275;
wire n_712;
wire n_246;
wire n_1583;
wire n_1042;
wire n_1402;
wire n_269;
wire n_285;
wire n_412;
wire n_1493;
wire n_657;
wire n_644;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_1621;
wire n_251;
wire n_160;
wire n_566;
wire n_565;
wire n_1448;
wire n_1507;
wire n_1398;
wire n_597;
wire n_1181;
wire n_1505;
wire n_1634;
wire n_1196;
wire n_651;
wire n_1340;
wire n_334;
wire n_811;
wire n_1558;
wire n_807;
wire n_835;
wire n_175;
wire n_666;
wire n_262;
wire n_1433;
wire n_1254;
wire n_1026;
wire n_1234;
wire n_319;
wire n_364;
wire n_1138;
wire n_927;
wire n_1089;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_242;
wire n_1681;
wire n_1018;
wire n_438;
wire n_713;
wire n_904;
wire n_1588;
wire n_1622;
wire n_166;
wire n_1180;
wire n_1271;
wire n_533;
wire n_1542;
wire n_1251;
wire n_278;

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_101),
.Y(n_155)
);

CKINVDCx5p33_ASAP7_75t_R g156 ( 
.A(n_40),
.Y(n_156)
);

CKINVDCx5p33_ASAP7_75t_R g157 ( 
.A(n_66),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_110),
.Y(n_158)
);

CKINVDCx16_ASAP7_75t_R g159 ( 
.A(n_77),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_82),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_70),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_116),
.Y(n_162)
);

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_86),
.Y(n_163)
);

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_93),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_91),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_117),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g167 ( 
.A(n_122),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_23),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_62),
.Y(n_169)
);

INVxp67_ASAP7_75t_L g170 ( 
.A(n_42),
.Y(n_170)
);

BUFx2_ASAP7_75t_L g171 ( 
.A(n_51),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_106),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_145),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_32),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_13),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_126),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_130),
.Y(n_177)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_27),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_80),
.Y(n_179)
);

BUFx3_ASAP7_75t_L g180 ( 
.A(n_1),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_40),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_69),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_19),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_99),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_123),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_78),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_8),
.Y(n_187)
);

BUFx3_ASAP7_75t_L g188 ( 
.A(n_79),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_137),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_121),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_151),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_143),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_100),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_76),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_132),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_64),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_141),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_127),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_153),
.Y(n_199)
);

BUFx8_ASAP7_75t_SL g200 ( 
.A(n_83),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_27),
.Y(n_201)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_49),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_22),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_134),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_13),
.Y(n_205)
);

BUFx3_ASAP7_75t_L g206 ( 
.A(n_103),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_52),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_55),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_3),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_3),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_2),
.Y(n_211)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_128),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_21),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_14),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_2),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_87),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_63),
.Y(n_217)
);

INVx1_ASAP7_75t_SL g218 ( 
.A(n_73),
.Y(n_218)
);

INVx1_ASAP7_75t_SL g219 ( 
.A(n_50),
.Y(n_219)
);

BUFx2_ASAP7_75t_SL g220 ( 
.A(n_98),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_120),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_1),
.Y(n_222)
);

BUFx10_ASAP7_75t_L g223 ( 
.A(n_41),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_95),
.Y(n_224)
);

BUFx6f_ASAP7_75t_L g225 ( 
.A(n_25),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_4),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_148),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_21),
.Y(n_228)
);

BUFx10_ASAP7_75t_L g229 ( 
.A(n_44),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_6),
.Y(n_230)
);

BUFx3_ASAP7_75t_L g231 ( 
.A(n_5),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_74),
.Y(n_232)
);

BUFx3_ASAP7_75t_L g233 ( 
.A(n_94),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_71),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_112),
.Y(n_235)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_5),
.Y(n_236)
);

HB1xp67_ASAP7_75t_L g237 ( 
.A(n_129),
.Y(n_237)
);

INVx2_ASAP7_75t_SL g238 ( 
.A(n_68),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_56),
.Y(n_239)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_142),
.Y(n_240)
);

BUFx8_ASAP7_75t_SL g241 ( 
.A(n_60),
.Y(n_241)
);

INVx1_ASAP7_75t_SL g242 ( 
.A(n_119),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_113),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_18),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_4),
.Y(n_245)
);

CKINVDCx16_ASAP7_75t_R g246 ( 
.A(n_81),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_37),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_31),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_38),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_111),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_125),
.Y(n_251)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_23),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_14),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_24),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_17),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_11),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_57),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_154),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_31),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_7),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_138),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_139),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_85),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_46),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_30),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_19),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_17),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_65),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_105),
.Y(n_269)
);

BUFx5_ASAP7_75t_L g270 ( 
.A(n_140),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_88),
.Y(n_271)
);

BUFx3_ASAP7_75t_L g272 ( 
.A(n_150),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_47),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_24),
.Y(n_274)
);

CKINVDCx16_ASAP7_75t_R g275 ( 
.A(n_96),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_75),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_46),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_131),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_67),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_135),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_38),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_59),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_146),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_84),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_58),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_18),
.Y(n_286)
);

BUFx3_ASAP7_75t_L g287 ( 
.A(n_147),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_92),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_108),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_104),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_25),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_7),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_53),
.Y(n_293)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_42),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_43),
.Y(n_295)
);

BUFx3_ASAP7_75t_L g296 ( 
.A(n_11),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_34),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_47),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_107),
.Y(n_299)
);

INVx2_ASAP7_75t_SL g300 ( 
.A(n_16),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_72),
.Y(n_301)
);

BUFx2_ASAP7_75t_SL g302 ( 
.A(n_29),
.Y(n_302)
);

INVx3_ASAP7_75t_L g303 ( 
.A(n_118),
.Y(n_303)
);

INVx1_ASAP7_75t_SL g304 ( 
.A(n_35),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_9),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_225),
.Y(n_306)
);

INVxp67_ASAP7_75t_SL g307 ( 
.A(n_237),
.Y(n_307)
);

INVxp33_ASAP7_75t_SL g308 ( 
.A(n_156),
.Y(n_308)
);

INVxp33_ASAP7_75t_L g309 ( 
.A(n_174),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_225),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_225),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_200),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_225),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_225),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_178),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_178),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_236),
.Y(n_317)
);

INVxp67_ASAP7_75t_SL g318 ( 
.A(n_171),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_236),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_252),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_252),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_241),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_294),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_294),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_180),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_180),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_231),
.Y(n_327)
);

INVxp67_ASAP7_75t_L g328 ( 
.A(n_223),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_195),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_231),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g331 ( 
.A(n_155),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_296),
.Y(n_332)
);

INVxp33_ASAP7_75t_L g333 ( 
.A(n_201),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_296),
.Y(n_334)
);

CKINVDCx20_ASAP7_75t_R g335 ( 
.A(n_176),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_214),
.Y(n_336)
);

INVxp67_ASAP7_75t_SL g337 ( 
.A(n_188),
.Y(n_337)
);

HB1xp67_ASAP7_75t_L g338 ( 
.A(n_156),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_197),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_198),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_222),
.Y(n_341)
);

INVxp33_ASAP7_75t_L g342 ( 
.A(n_228),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_248),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_249),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_199),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_254),
.Y(n_346)
);

CKINVDCx20_ASAP7_75t_R g347 ( 
.A(n_177),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_256),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_267),
.Y(n_349)
);

CKINVDCx20_ASAP7_75t_R g350 ( 
.A(n_192),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_273),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_281),
.Y(n_352)
);

INVx2_ASAP7_75t_SL g353 ( 
.A(n_223),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_300),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_216),
.Y(n_355)
);

INVx3_ASAP7_75t_L g356 ( 
.A(n_188),
.Y(n_356)
);

INVx2_ASAP7_75t_L g357 ( 
.A(n_270),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_300),
.Y(n_358)
);

INVx2_ASAP7_75t_L g359 ( 
.A(n_270),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_202),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_217),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_224),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_202),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_212),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_212),
.Y(n_365)
);

CKINVDCx20_ASAP7_75t_R g366 ( 
.A(n_227),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_240),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_240),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_158),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_160),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_165),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_169),
.Y(n_372)
);

CKINVDCx20_ASAP7_75t_R g373 ( 
.A(n_278),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_172),
.Y(n_374)
);

BUFx3_ASAP7_75t_L g375 ( 
.A(n_206),
.Y(n_375)
);

AOI22xp5_ASAP7_75t_L g376 ( 
.A1(n_307),
.A2(n_245),
.B1(n_295),
.B2(n_297),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_SL g377 ( 
.A(n_353),
.B(n_159),
.Y(n_377)
);

AND2x2_ASAP7_75t_L g378 ( 
.A(n_337),
.B(n_303),
.Y(n_378)
);

HB1xp67_ASAP7_75t_L g379 ( 
.A(n_338),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_306),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_356),
.B(n_238),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_329),
.Y(n_382)
);

CKINVDCx20_ASAP7_75t_R g383 ( 
.A(n_331),
.Y(n_383)
);

INVxp67_ASAP7_75t_L g384 ( 
.A(n_375),
.Y(n_384)
);

AND2x2_ASAP7_75t_L g385 ( 
.A(n_356),
.B(n_303),
.Y(n_385)
);

CKINVDCx20_ASAP7_75t_R g386 ( 
.A(n_335),
.Y(n_386)
);

CKINVDCx20_ASAP7_75t_R g387 ( 
.A(n_347),
.Y(n_387)
);

AND2x4_ASAP7_75t_L g388 ( 
.A(n_356),
.B(n_206),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_306),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_339),
.Y(n_390)
);

INVx2_ASAP7_75t_L g391 ( 
.A(n_310),
.Y(n_391)
);

BUFx6f_ASAP7_75t_L g392 ( 
.A(n_357),
.Y(n_392)
);

BUFx3_ASAP7_75t_L g393 ( 
.A(n_375),
.Y(n_393)
);

NOR2xp33_ASAP7_75t_L g394 ( 
.A(n_340),
.B(n_246),
.Y(n_394)
);

BUFx2_ASAP7_75t_L g395 ( 
.A(n_328),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_310),
.Y(n_396)
);

AND2x2_ASAP7_75t_L g397 ( 
.A(n_369),
.B(n_303),
.Y(n_397)
);

BUFx6f_ASAP7_75t_L g398 ( 
.A(n_357),
.Y(n_398)
);

INVx2_ASAP7_75t_L g399 ( 
.A(n_311),
.Y(n_399)
);

BUFx6f_ASAP7_75t_L g400 ( 
.A(n_359),
.Y(n_400)
);

BUFx6f_ASAP7_75t_L g401 ( 
.A(n_359),
.Y(n_401)
);

INVx3_ASAP7_75t_L g402 ( 
.A(n_311),
.Y(n_402)
);

CKINVDCx20_ASAP7_75t_R g403 ( 
.A(n_350),
.Y(n_403)
);

AOI22xp5_ASAP7_75t_L g404 ( 
.A1(n_318),
.A2(n_266),
.B1(n_298),
.B2(n_297),
.Y(n_404)
);

AND2x4_ASAP7_75t_L g405 ( 
.A(n_369),
.B(n_233),
.Y(n_405)
);

AND2x4_ASAP7_75t_L g406 ( 
.A(n_370),
.B(n_233),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_313),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_313),
.Y(n_408)
);

BUFx8_ASAP7_75t_L g409 ( 
.A(n_353),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_314),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_345),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_314),
.Y(n_412)
);

AND2x2_ASAP7_75t_L g413 ( 
.A(n_370),
.B(n_272),
.Y(n_413)
);

AND2x2_ASAP7_75t_L g414 ( 
.A(n_371),
.B(n_272),
.Y(n_414)
);

NOR2xp33_ASAP7_75t_L g415 ( 
.A(n_355),
.B(n_275),
.Y(n_415)
);

INVx2_ASAP7_75t_L g416 ( 
.A(n_360),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_360),
.Y(n_417)
);

CKINVDCx16_ASAP7_75t_R g418 ( 
.A(n_366),
.Y(n_418)
);

BUFx6f_ASAP7_75t_L g419 ( 
.A(n_363),
.Y(n_419)
);

BUFx2_ASAP7_75t_L g420 ( 
.A(n_361),
.Y(n_420)
);

BUFx8_ASAP7_75t_L g421 ( 
.A(n_325),
.Y(n_421)
);

BUFx2_ASAP7_75t_L g422 ( 
.A(n_362),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_371),
.B(n_238),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_363),
.Y(n_424)
);

AND2x2_ASAP7_75t_L g425 ( 
.A(n_372),
.B(n_287),
.Y(n_425)
);

BUFx6f_ASAP7_75t_L g426 ( 
.A(n_364),
.Y(n_426)
);

INVx3_ASAP7_75t_L g427 ( 
.A(n_364),
.Y(n_427)
);

NOR2xp33_ASAP7_75t_L g428 ( 
.A(n_308),
.B(n_218),
.Y(n_428)
);

INVx2_ASAP7_75t_L g429 ( 
.A(n_365),
.Y(n_429)
);

BUFx3_ASAP7_75t_L g430 ( 
.A(n_325),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_365),
.Y(n_431)
);

NOR2xp67_ASAP7_75t_L g432 ( 
.A(n_367),
.B(n_173),
.Y(n_432)
);

HB1xp67_ASAP7_75t_L g433 ( 
.A(n_326),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_372),
.B(n_157),
.Y(n_434)
);

INVx2_ASAP7_75t_L g435 ( 
.A(n_367),
.Y(n_435)
);

INVx2_ASAP7_75t_L g436 ( 
.A(n_368),
.Y(n_436)
);

CKINVDCx5p33_ASAP7_75t_R g437 ( 
.A(n_312),
.Y(n_437)
);

INVx2_ASAP7_75t_L g438 ( 
.A(n_368),
.Y(n_438)
);

AND2x4_ASAP7_75t_L g439 ( 
.A(n_374),
.B(n_287),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_378),
.B(n_374),
.Y(n_440)
);

INVxp67_ASAP7_75t_L g441 ( 
.A(n_428),
.Y(n_441)
);

INVx2_ASAP7_75t_L g442 ( 
.A(n_391),
.Y(n_442)
);

BUFx10_ASAP7_75t_L g443 ( 
.A(n_394),
.Y(n_443)
);

INVx2_ASAP7_75t_L g444 ( 
.A(n_391),
.Y(n_444)
);

AOI22xp33_ASAP7_75t_L g445 ( 
.A1(n_378),
.A2(n_388),
.B1(n_385),
.B2(n_397),
.Y(n_445)
);

AO21x2_ASAP7_75t_L g446 ( 
.A1(n_381),
.A2(n_434),
.B(n_184),
.Y(n_446)
);

INVx2_ASAP7_75t_L g447 ( 
.A(n_391),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_380),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_380),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_389),
.Y(n_450)
);

AOI22xp5_ASAP7_75t_L g451 ( 
.A1(n_415),
.A2(n_283),
.B1(n_373),
.B2(n_322),
.Y(n_451)
);

INVxp33_ASAP7_75t_SL g452 ( 
.A(n_404),
.Y(n_452)
);

AND2x2_ASAP7_75t_SL g453 ( 
.A(n_388),
.B(n_167),
.Y(n_453)
);

INVx2_ASAP7_75t_SL g454 ( 
.A(n_393),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_389),
.Y(n_455)
);

INVx2_ASAP7_75t_L g456 ( 
.A(n_399),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_L g457 ( 
.A(n_378),
.B(n_219),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_388),
.B(n_242),
.Y(n_458)
);

AND2x2_ASAP7_75t_L g459 ( 
.A(n_430),
.B(n_326),
.Y(n_459)
);

AND2x2_ASAP7_75t_L g460 ( 
.A(n_430),
.B(n_327),
.Y(n_460)
);

BUFx10_ASAP7_75t_L g461 ( 
.A(n_437),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_388),
.B(n_385),
.Y(n_462)
);

OR2x6_ASAP7_75t_L g463 ( 
.A(n_420),
.B(n_302),
.Y(n_463)
);

INVx2_ASAP7_75t_L g464 ( 
.A(n_399),
.Y(n_464)
);

INVx5_ASAP7_75t_L g465 ( 
.A(n_392),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_396),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_396),
.Y(n_467)
);

XOR2xp5_ASAP7_75t_L g468 ( 
.A(n_376),
.B(n_168),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_407),
.Y(n_469)
);

INVx2_ASAP7_75t_L g470 ( 
.A(n_399),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_408),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_SL g472 ( 
.A(n_377),
.B(n_157),
.Y(n_472)
);

INVx3_ASAP7_75t_L g473 ( 
.A(n_392),
.Y(n_473)
);

INVx4_ASAP7_75t_L g474 ( 
.A(n_392),
.Y(n_474)
);

INVx3_ASAP7_75t_L g475 ( 
.A(n_392),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_385),
.B(n_384),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_408),
.Y(n_477)
);

INVx2_ASAP7_75t_L g478 ( 
.A(n_410),
.Y(n_478)
);

INVx2_ASAP7_75t_L g479 ( 
.A(n_410),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_L g480 ( 
.A(n_384),
.B(n_232),
.Y(n_480)
);

NAND2xp33_ASAP7_75t_SL g481 ( 
.A(n_395),
.B(n_168),
.Y(n_481)
);

BUFx8_ASAP7_75t_SL g482 ( 
.A(n_383),
.Y(n_482)
);

INVx2_ASAP7_75t_L g483 ( 
.A(n_412),
.Y(n_483)
);

INVx3_ASAP7_75t_L g484 ( 
.A(n_392),
.Y(n_484)
);

CKINVDCx5p33_ASAP7_75t_R g485 ( 
.A(n_409),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_L g486 ( 
.A(n_393),
.B(n_235),
.Y(n_486)
);

INVxp67_ASAP7_75t_L g487 ( 
.A(n_395),
.Y(n_487)
);

INVx8_ASAP7_75t_L g488 ( 
.A(n_382),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_SL g489 ( 
.A(n_409),
.B(n_161),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_L g490 ( 
.A(n_393),
.B(n_239),
.Y(n_490)
);

INVx2_ASAP7_75t_L g491 ( 
.A(n_412),
.Y(n_491)
);

AO21x2_ASAP7_75t_L g492 ( 
.A1(n_381),
.A2(n_185),
.B(n_182),
.Y(n_492)
);

HB1xp67_ASAP7_75t_L g493 ( 
.A(n_379),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_405),
.B(n_243),
.Y(n_494)
);

NOR2xp33_ASAP7_75t_L g495 ( 
.A(n_390),
.B(n_309),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_402),
.Y(n_496)
);

AND2x2_ASAP7_75t_L g497 ( 
.A(n_430),
.B(n_327),
.Y(n_497)
);

NOR2xp33_ASAP7_75t_L g498 ( 
.A(n_411),
.B(n_333),
.Y(n_498)
);

BUFx6f_ASAP7_75t_L g499 ( 
.A(n_392),
.Y(n_499)
);

INVx2_ASAP7_75t_L g500 ( 
.A(n_402),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_SL g501 ( 
.A(n_409),
.B(n_161),
.Y(n_501)
);

CKINVDCx5p33_ASAP7_75t_R g502 ( 
.A(n_409),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_402),
.Y(n_503)
);

INVxp33_ASAP7_75t_L g504 ( 
.A(n_379),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_402),
.Y(n_505)
);

AND3x2_ASAP7_75t_L g506 ( 
.A(n_420),
.B(n_170),
.C(n_189),
.Y(n_506)
);

NAND3xp33_ASAP7_75t_L g507 ( 
.A(n_434),
.B(n_332),
.C(n_330),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_L g508 ( 
.A(n_405),
.B(n_250),
.Y(n_508)
);

INVxp67_ASAP7_75t_L g509 ( 
.A(n_433),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_417),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_417),
.Y(n_511)
);

INVx2_ASAP7_75t_L g512 ( 
.A(n_416),
.Y(n_512)
);

INVxp67_ASAP7_75t_SL g513 ( 
.A(n_392),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_424),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_SL g515 ( 
.A(n_422),
.B(n_421),
.Y(n_515)
);

OR2x2_ASAP7_75t_L g516 ( 
.A(n_404),
.B(n_330),
.Y(n_516)
);

INVx2_ASAP7_75t_L g517 ( 
.A(n_416),
.Y(n_517)
);

AND2x2_ASAP7_75t_L g518 ( 
.A(n_413),
.B(n_332),
.Y(n_518)
);

OAI22xp5_ASAP7_75t_L g519 ( 
.A1(n_376),
.A2(n_253),
.B1(n_247),
.B2(n_244),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_433),
.Y(n_520)
);

NOR2xp33_ASAP7_75t_L g521 ( 
.A(n_422),
.B(n_342),
.Y(n_521)
);

INVx2_ASAP7_75t_SL g522 ( 
.A(n_413),
.Y(n_522)
);

INVx2_ASAP7_75t_SL g523 ( 
.A(n_413),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_424),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_SL g525 ( 
.A(n_421),
.B(n_162),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_SL g526 ( 
.A(n_421),
.B(n_162),
.Y(n_526)
);

BUFx3_ASAP7_75t_L g527 ( 
.A(n_405),
.Y(n_527)
);

AOI22xp33_ASAP7_75t_L g528 ( 
.A1(n_397),
.A2(n_220),
.B1(n_346),
.B2(n_344),
.Y(n_528)
);

BUFx10_ASAP7_75t_L g529 ( 
.A(n_405),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_431),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_L g531 ( 
.A(n_406),
.B(n_251),
.Y(n_531)
);

INVx2_ASAP7_75t_L g532 ( 
.A(n_416),
.Y(n_532)
);

INVx2_ASAP7_75t_L g533 ( 
.A(n_429),
.Y(n_533)
);

NOR2xp67_ASAP7_75t_L g534 ( 
.A(n_423),
.B(n_257),
.Y(n_534)
);

INVx2_ASAP7_75t_L g535 ( 
.A(n_429),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_431),
.Y(n_536)
);

INVx2_ASAP7_75t_L g537 ( 
.A(n_429),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_398),
.Y(n_538)
);

INVx3_ASAP7_75t_L g539 ( 
.A(n_398),
.Y(n_539)
);

AND2x2_ASAP7_75t_L g540 ( 
.A(n_414),
.B(n_334),
.Y(n_540)
);

AOI22xp5_ASAP7_75t_L g541 ( 
.A1(n_406),
.A2(n_261),
.B1(n_193),
.B2(n_186),
.Y(n_541)
);

NOR2xp33_ASAP7_75t_L g542 ( 
.A(n_406),
.B(n_334),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_SL g543 ( 
.A(n_421),
.B(n_163),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_398),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_398),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_398),
.Y(n_546)
);

INVx2_ASAP7_75t_L g547 ( 
.A(n_435),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_398),
.Y(n_548)
);

INVx2_ASAP7_75t_L g549 ( 
.A(n_435),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_398),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_400),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_400),
.Y(n_552)
);

INVx2_ASAP7_75t_L g553 ( 
.A(n_435),
.Y(n_553)
);

CKINVDCx5p33_ASAP7_75t_R g554 ( 
.A(n_418),
.Y(n_554)
);

NOR2xp33_ASAP7_75t_L g555 ( 
.A(n_406),
.B(n_354),
.Y(n_555)
);

INVx2_ASAP7_75t_L g556 ( 
.A(n_436),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_SL g557 ( 
.A(n_439),
.B(n_163),
.Y(n_557)
);

INVx2_ASAP7_75t_L g558 ( 
.A(n_436),
.Y(n_558)
);

INVx2_ASAP7_75t_L g559 ( 
.A(n_436),
.Y(n_559)
);

INVx2_ASAP7_75t_L g560 ( 
.A(n_438),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_400),
.Y(n_561)
);

AO22x2_ASAP7_75t_L g562 ( 
.A1(n_397),
.A2(n_304),
.B1(n_190),
.B2(n_301),
.Y(n_562)
);

INVx2_ASAP7_75t_L g563 ( 
.A(n_438),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_400),
.Y(n_564)
);

INVx3_ASAP7_75t_L g565 ( 
.A(n_400),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_L g566 ( 
.A(n_439),
.B(n_258),
.Y(n_566)
);

INVx2_ASAP7_75t_L g567 ( 
.A(n_438),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_400),
.Y(n_568)
);

INVx4_ASAP7_75t_L g569 ( 
.A(n_400),
.Y(n_569)
);

CKINVDCx16_ASAP7_75t_R g570 ( 
.A(n_418),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_401),
.Y(n_571)
);

AND2x4_ASAP7_75t_L g572 ( 
.A(n_439),
.B(n_341),
.Y(n_572)
);

INVx2_ASAP7_75t_L g573 ( 
.A(n_401),
.Y(n_573)
);

NAND2xp33_ASAP7_75t_L g574 ( 
.A(n_401),
.B(n_167),
.Y(n_574)
);

BUFx2_ASAP7_75t_L g575 ( 
.A(n_386),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_L g576 ( 
.A(n_439),
.B(n_401),
.Y(n_576)
);

BUFx6f_ASAP7_75t_L g577 ( 
.A(n_401),
.Y(n_577)
);

CKINVDCx5p33_ASAP7_75t_R g578 ( 
.A(n_387),
.Y(n_578)
);

INVx2_ASAP7_75t_L g579 ( 
.A(n_401),
.Y(n_579)
);

CKINVDCx5p33_ASAP7_75t_R g580 ( 
.A(n_403),
.Y(n_580)
);

NOR2xp33_ASAP7_75t_L g581 ( 
.A(n_423),
.B(n_354),
.Y(n_581)
);

NAND2xp33_ASAP7_75t_SL g582 ( 
.A(n_414),
.B(n_175),
.Y(n_582)
);

INVx2_ASAP7_75t_L g583 ( 
.A(n_401),
.Y(n_583)
);

BUFx6f_ASAP7_75t_L g584 ( 
.A(n_419),
.Y(n_584)
);

NAND3xp33_ASAP7_75t_L g585 ( 
.A(n_414),
.B(n_343),
.C(n_349),
.Y(n_585)
);

INVx2_ASAP7_75t_L g586 ( 
.A(n_442),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_L g587 ( 
.A(n_445),
.B(n_427),
.Y(n_587)
);

INVx2_ASAP7_75t_L g588 ( 
.A(n_442),
.Y(n_588)
);

AO22x2_ASAP7_75t_L g589 ( 
.A1(n_468),
.A2(n_234),
.B1(n_221),
.B2(n_208),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_L g590 ( 
.A(n_476),
.B(n_427),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_SL g591 ( 
.A(n_453),
.B(n_167),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_L g592 ( 
.A(n_522),
.B(n_427),
.Y(n_592)
);

NOR2xp33_ASAP7_75t_L g593 ( 
.A(n_441),
.B(n_509),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_527),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_L g595 ( 
.A(n_522),
.B(n_427),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_L g596 ( 
.A(n_523),
.B(n_425),
.Y(n_596)
);

AOI22xp5_ASAP7_75t_L g597 ( 
.A1(n_523),
.A2(n_425),
.B1(n_164),
.B2(n_276),
.Y(n_597)
);

NOR2xp33_ASAP7_75t_L g598 ( 
.A(n_457),
.B(n_164),
.Y(n_598)
);

BUFx6f_ASAP7_75t_L g599 ( 
.A(n_527),
.Y(n_599)
);

NOR2xp33_ASAP7_75t_L g600 ( 
.A(n_520),
.B(n_166),
.Y(n_600)
);

AND2x2_ASAP7_75t_L g601 ( 
.A(n_521),
.B(n_425),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_510),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_SL g603 ( 
.A(n_453),
.B(n_167),
.Y(n_603)
);

BUFx3_ASAP7_75t_L g604 ( 
.A(n_454),
.Y(n_604)
);

INVx2_ASAP7_75t_SL g605 ( 
.A(n_518),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_L g606 ( 
.A(n_440),
.B(n_419),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_SL g607 ( 
.A(n_462),
.B(n_167),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_SL g608 ( 
.A(n_576),
.B(n_270),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_L g609 ( 
.A(n_446),
.B(n_419),
.Y(n_609)
);

NAND2xp33_ASAP7_75t_L g610 ( 
.A(n_454),
.B(n_458),
.Y(n_610)
);

INVx2_ASAP7_75t_L g611 ( 
.A(n_444),
.Y(n_611)
);

OR2x2_ASAP7_75t_L g612 ( 
.A(n_493),
.B(n_348),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_L g613 ( 
.A(n_446),
.B(n_419),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_SL g614 ( 
.A(n_529),
.B(n_270),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_SL g615 ( 
.A(n_529),
.B(n_270),
.Y(n_615)
);

INVx2_ASAP7_75t_L g616 ( 
.A(n_444),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_SL g617 ( 
.A(n_529),
.B(n_270),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_L g618 ( 
.A(n_446),
.B(n_419),
.Y(n_618)
);

AND2x2_ASAP7_75t_L g619 ( 
.A(n_495),
.B(n_358),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_L g620 ( 
.A(n_542),
.B(n_419),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_510),
.Y(n_621)
);

NOR3xp33_ASAP7_75t_L g622 ( 
.A(n_498),
.B(n_358),
.C(n_336),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_L g623 ( 
.A(n_511),
.B(n_419),
.Y(n_623)
);

INVx4_ASAP7_75t_L g624 ( 
.A(n_584),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_L g625 ( 
.A(n_511),
.B(n_426),
.Y(n_625)
);

INVx2_ASAP7_75t_L g626 ( 
.A(n_447),
.Y(n_626)
);

NOR2xp33_ASAP7_75t_SL g627 ( 
.A(n_461),
.B(n_166),
.Y(n_627)
);

INVx2_ASAP7_75t_L g628 ( 
.A(n_447),
.Y(n_628)
);

O2A1O1Ixp33_ASAP7_75t_L g629 ( 
.A1(n_581),
.A2(n_336),
.B(n_352),
.C(n_351),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_L g630 ( 
.A(n_514),
.B(n_426),
.Y(n_630)
);

INVx2_ASAP7_75t_L g631 ( 
.A(n_456),
.Y(n_631)
);

INVx2_ASAP7_75t_L g632 ( 
.A(n_456),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_L g633 ( 
.A(n_524),
.B(n_530),
.Y(n_633)
);

NOR2xp33_ASAP7_75t_L g634 ( 
.A(n_516),
.B(n_487),
.Y(n_634)
);

INVx2_ASAP7_75t_L g635 ( 
.A(n_464),
.Y(n_635)
);

INVx2_ASAP7_75t_L g636 ( 
.A(n_464),
.Y(n_636)
);

INVx2_ASAP7_75t_L g637 ( 
.A(n_470),
.Y(n_637)
);

NOR2xp33_ASAP7_75t_L g638 ( 
.A(n_516),
.B(n_179),
.Y(n_638)
);

NOR2xp33_ASAP7_75t_L g639 ( 
.A(n_472),
.B(n_179),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_L g640 ( 
.A(n_524),
.B(n_530),
.Y(n_640)
);

INVx2_ASAP7_75t_L g641 ( 
.A(n_470),
.Y(n_641)
);

INVx2_ASAP7_75t_SL g642 ( 
.A(n_518),
.Y(n_642)
);

INVx2_ASAP7_75t_L g643 ( 
.A(n_512),
.Y(n_643)
);

INVx2_ASAP7_75t_L g644 ( 
.A(n_512),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_SL g645 ( 
.A(n_572),
.B(n_270),
.Y(n_645)
);

NAND2x1_ASAP7_75t_L g646 ( 
.A(n_474),
.B(n_426),
.Y(n_646)
);

INVx8_ASAP7_75t_L g647 ( 
.A(n_488),
.Y(n_647)
);

BUFx6f_ASAP7_75t_L g648 ( 
.A(n_572),
.Y(n_648)
);

NAND2x1_ASAP7_75t_L g649 ( 
.A(n_474),
.B(n_426),
.Y(n_649)
);

BUFx12f_ASAP7_75t_SL g650 ( 
.A(n_463),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_L g651 ( 
.A(n_536),
.B(n_426),
.Y(n_651)
);

AOI22xp5_ASAP7_75t_L g652 ( 
.A1(n_572),
.A2(n_276),
.B1(n_193),
.B2(n_261),
.Y(n_652)
);

INVx2_ASAP7_75t_L g653 ( 
.A(n_517),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_L g654 ( 
.A(n_536),
.B(n_426),
.Y(n_654)
);

INVxp67_ASAP7_75t_L g655 ( 
.A(n_481),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_459),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_459),
.Y(n_657)
);

INVxp67_ASAP7_75t_SL g658 ( 
.A(n_499),
.Y(n_658)
);

NOR2xp33_ASAP7_75t_L g659 ( 
.A(n_541),
.B(n_186),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_L g660 ( 
.A(n_448),
.B(n_426),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_460),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_460),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_SL g663 ( 
.A(n_534),
.B(n_262),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_L g664 ( 
.A(n_448),
.B(n_432),
.Y(n_664)
);

HB1xp67_ASAP7_75t_L g665 ( 
.A(n_575),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_L g666 ( 
.A(n_449),
.B(n_450),
.Y(n_666)
);

AO221x1_ASAP7_75t_L g667 ( 
.A1(n_562),
.A2(n_207),
.B1(n_299),
.B2(n_191),
.C(n_194),
.Y(n_667)
);

AOI22xp33_ASAP7_75t_L g668 ( 
.A1(n_562),
.A2(n_270),
.B1(n_289),
.B2(n_290),
.Y(n_668)
);

OAI22xp5_ASAP7_75t_L g669 ( 
.A1(n_494),
.A2(n_196),
.B1(n_293),
.B2(n_204),
.Y(n_669)
);

BUFx6f_ASAP7_75t_L g670 ( 
.A(n_499),
.Y(n_670)
);

NOR2xp33_ASAP7_75t_L g671 ( 
.A(n_480),
.B(n_262),
.Y(n_671)
);

NOR2xp33_ASAP7_75t_L g672 ( 
.A(n_557),
.B(n_263),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_L g673 ( 
.A(n_449),
.B(n_432),
.Y(n_673)
);

AOI22xp5_ASAP7_75t_L g674 ( 
.A1(n_508),
.A2(n_280),
.B1(n_268),
.B2(n_288),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_497),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_L g676 ( 
.A(n_450),
.B(n_263),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_L g677 ( 
.A(n_455),
.B(n_268),
.Y(n_677)
);

INVxp67_ASAP7_75t_L g678 ( 
.A(n_582),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_SL g679 ( 
.A(n_496),
.B(n_269),
.Y(n_679)
);

AND2x2_ASAP7_75t_L g680 ( 
.A(n_504),
.B(n_229),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_497),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_455),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_SL g683 ( 
.A(n_496),
.B(n_269),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_466),
.B(n_271),
.Y(n_684)
);

INVxp67_ASAP7_75t_L g685 ( 
.A(n_555),
.Y(n_685)
);

NOR2xp33_ASAP7_75t_L g686 ( 
.A(n_531),
.B(n_271),
.Y(n_686)
);

NAND2x1_ASAP7_75t_L g687 ( 
.A(n_474),
.B(n_569),
.Y(n_687)
);

INVx4_ASAP7_75t_L g688 ( 
.A(n_584),
.Y(n_688)
);

NOR2xp33_ASAP7_75t_SL g689 ( 
.A(n_461),
.B(n_279),
.Y(n_689)
);

AND2x2_ASAP7_75t_L g690 ( 
.A(n_540),
.B(n_351),
.Y(n_690)
);

BUFx6f_ASAP7_75t_L g691 ( 
.A(n_499),
.Y(n_691)
);

OAI22xp5_ASAP7_75t_L g692 ( 
.A1(n_566),
.A2(n_282),
.B1(n_279),
.B2(n_280),
.Y(n_692)
);

BUFx6f_ASAP7_75t_L g693 ( 
.A(n_499),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_SL g694 ( 
.A(n_503),
.B(n_282),
.Y(n_694)
);

NOR2xp33_ASAP7_75t_L g695 ( 
.A(n_452),
.B(n_284),
.Y(n_695)
);

NOR2xp33_ASAP7_75t_L g696 ( 
.A(n_486),
.B(n_284),
.Y(n_696)
);

INVx2_ASAP7_75t_L g697 ( 
.A(n_517),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_L g698 ( 
.A(n_467),
.B(n_285),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_L g699 ( 
.A(n_467),
.B(n_285),
.Y(n_699)
);

NOR3xp33_ASAP7_75t_L g700 ( 
.A(n_519),
.B(n_352),
.C(n_203),
.Y(n_700)
);

HB1xp67_ASAP7_75t_L g701 ( 
.A(n_575),
.Y(n_701)
);

A2O1A1Ixp33_ASAP7_75t_L g702 ( 
.A1(n_469),
.A2(n_288),
.B(n_323),
.C(n_321),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_SL g703 ( 
.A(n_528),
.B(n_443),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_SL g704 ( 
.A(n_503),
.B(n_205),
.Y(n_704)
);

NOR2xp33_ASAP7_75t_L g705 ( 
.A(n_490),
.B(n_489),
.Y(n_705)
);

AND2x2_ASAP7_75t_L g706 ( 
.A(n_443),
.B(n_315),
.Y(n_706)
);

NOR2xp33_ASAP7_75t_L g707 ( 
.A(n_501),
.B(n_471),
.Y(n_707)
);

AOI22xp33_ASAP7_75t_L g708 ( 
.A1(n_562),
.A2(n_265),
.B1(n_183),
.B2(n_187),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_SL g709 ( 
.A(n_505),
.B(n_209),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_L g710 ( 
.A(n_471),
.B(n_210),
.Y(n_710)
);

INVx2_ASAP7_75t_L g711 ( 
.A(n_532),
.Y(n_711)
);

BUFx2_ASAP7_75t_L g712 ( 
.A(n_463),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_477),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_477),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_SL g715 ( 
.A(n_505),
.B(n_211),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_L g716 ( 
.A(n_513),
.B(n_213),
.Y(n_716)
);

INVx2_ASAP7_75t_L g717 ( 
.A(n_532),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_SL g718 ( 
.A(n_500),
.B(n_215),
.Y(n_718)
);

AND2x2_ASAP7_75t_L g719 ( 
.A(n_443),
.B(n_315),
.Y(n_719)
);

NOR2xp33_ASAP7_75t_L g720 ( 
.A(n_525),
.B(n_226),
.Y(n_720)
);

NOR3xp33_ASAP7_75t_L g721 ( 
.A(n_570),
.B(n_255),
.C(n_259),
.Y(n_721)
);

CKINVDCx5p33_ASAP7_75t_R g722 ( 
.A(n_482),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_478),
.Y(n_723)
);

CKINVDCx5p33_ASAP7_75t_R g724 ( 
.A(n_578),
.Y(n_724)
);

O2A1O1Ixp5_ASAP7_75t_L g725 ( 
.A1(n_473),
.A2(n_324),
.B(n_323),
.C(n_321),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_L g726 ( 
.A(n_478),
.B(n_305),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_SL g727 ( 
.A(n_500),
.B(n_277),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_SL g728 ( 
.A(n_573),
.B(n_277),
.Y(n_728)
);

OAI21xp5_ASAP7_75t_L g729 ( 
.A1(n_538),
.A2(n_324),
.B(n_320),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_SL g730 ( 
.A(n_573),
.B(n_579),
.Y(n_730)
);

INVx2_ASAP7_75t_L g731 ( 
.A(n_533),
.Y(n_731)
);

BUFx6f_ASAP7_75t_L g732 ( 
.A(n_499),
.Y(n_732)
);

NOR2xp33_ASAP7_75t_L g733 ( 
.A(n_526),
.B(n_181),
.Y(n_733)
);

AO22x2_ASAP7_75t_L g734 ( 
.A1(n_468),
.A2(n_320),
.B1(n_319),
.B2(n_317),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_479),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_L g736 ( 
.A(n_479),
.B(n_319),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_L g737 ( 
.A(n_483),
.B(n_317),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_L g738 ( 
.A(n_491),
.B(n_316),
.Y(n_738)
);

INVx3_ASAP7_75t_L g739 ( 
.A(n_533),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_SL g740 ( 
.A(n_579),
.B(n_265),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_535),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_535),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_SL g743 ( 
.A(n_583),
.B(n_266),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_537),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_SL g745 ( 
.A(n_583),
.B(n_298),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_L g746 ( 
.A(n_544),
.B(n_292),
.Y(n_746)
);

OR2x2_ASAP7_75t_L g747 ( 
.A(n_463),
.B(n_292),
.Y(n_747)
);

INVx2_ASAP7_75t_L g748 ( 
.A(n_739),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_L g749 ( 
.A(n_601),
.B(n_685),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_723),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_SL g751 ( 
.A(n_648),
.B(n_461),
.Y(n_751)
);

AND2x4_ASAP7_75t_L g752 ( 
.A(n_605),
.B(n_515),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_735),
.Y(n_753)
);

AND2x4_ASAP7_75t_L g754 ( 
.A(n_642),
.B(n_463),
.Y(n_754)
);

BUFx3_ASAP7_75t_L g755 ( 
.A(n_647),
.Y(n_755)
);

AND2x2_ASAP7_75t_L g756 ( 
.A(n_619),
.B(n_451),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_602),
.Y(n_757)
);

NOR2xp33_ASAP7_75t_L g758 ( 
.A(n_593),
.B(n_488),
.Y(n_758)
);

INVxp67_ASAP7_75t_L g759 ( 
.A(n_680),
.Y(n_759)
);

INVx5_ASAP7_75t_L g760 ( 
.A(n_670),
.Y(n_760)
);

AND2x2_ASAP7_75t_L g761 ( 
.A(n_706),
.B(n_580),
.Y(n_761)
);

INVx2_ASAP7_75t_L g762 ( 
.A(n_739),
.Y(n_762)
);

AOI22xp5_ASAP7_75t_L g763 ( 
.A1(n_705),
.A2(n_492),
.B1(n_543),
.B2(n_507),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_L g764 ( 
.A(n_598),
.B(n_492),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_L g765 ( 
.A(n_598),
.B(n_492),
.Y(n_765)
);

AOI22xp33_ASAP7_75t_L g766 ( 
.A1(n_668),
.A2(n_562),
.B1(n_585),
.B2(n_563),
.Y(n_766)
);

AOI22xp5_ASAP7_75t_L g767 ( 
.A1(n_705),
.A2(n_551),
.B1(n_552),
.B2(n_550),
.Y(n_767)
);

BUFx2_ASAP7_75t_L g768 ( 
.A(n_665),
.Y(n_768)
);

INVx2_ASAP7_75t_L g769 ( 
.A(n_586),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_621),
.Y(n_770)
);

BUFx2_ASAP7_75t_L g771 ( 
.A(n_701),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_SL g772 ( 
.A(n_648),
.B(n_544),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_L g773 ( 
.A(n_596),
.B(n_671),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_682),
.Y(n_774)
);

OR2x2_ASAP7_75t_L g775 ( 
.A(n_612),
.B(n_554),
.Y(n_775)
);

INVx2_ASAP7_75t_L g776 ( 
.A(n_588),
.Y(n_776)
);

INVx2_ASAP7_75t_L g777 ( 
.A(n_611),
.Y(n_777)
);

AND3x1_ASAP7_75t_L g778 ( 
.A(n_695),
.B(n_506),
.C(n_181),
.Y(n_778)
);

AOI22xp5_ASAP7_75t_L g779 ( 
.A1(n_707),
.A2(n_552),
.B1(n_561),
.B2(n_545),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_L g780 ( 
.A(n_671),
.B(n_545),
.Y(n_780)
);

BUFx6f_ASAP7_75t_L g781 ( 
.A(n_648),
.Y(n_781)
);

AND2x4_ASAP7_75t_L g782 ( 
.A(n_656),
.B(n_657),
.Y(n_782)
);

HB1xp67_ASAP7_75t_L g783 ( 
.A(n_719),
.Y(n_783)
);

NOR2xp33_ASAP7_75t_L g784 ( 
.A(n_593),
.B(n_488),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_L g785 ( 
.A(n_604),
.B(n_546),
.Y(n_785)
);

INVx2_ASAP7_75t_SL g786 ( 
.A(n_690),
.Y(n_786)
);

INVx3_ASAP7_75t_L g787 ( 
.A(n_599),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_L g788 ( 
.A(n_604),
.B(n_546),
.Y(n_788)
);

INVx2_ASAP7_75t_L g789 ( 
.A(n_616),
.Y(n_789)
);

BUFx6f_ASAP7_75t_L g790 ( 
.A(n_648),
.Y(n_790)
);

AOI22xp5_ASAP7_75t_L g791 ( 
.A1(n_707),
.A2(n_564),
.B1(n_550),
.B2(n_548),
.Y(n_791)
);

NAND2x1p5_ASAP7_75t_L g792 ( 
.A(n_599),
.B(n_473),
.Y(n_792)
);

INVx2_ASAP7_75t_L g793 ( 
.A(n_626),
.Y(n_793)
);

INVx2_ASAP7_75t_SL g794 ( 
.A(n_747),
.Y(n_794)
);

INVx3_ASAP7_75t_L g795 ( 
.A(n_599),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_SL g796 ( 
.A(n_599),
.B(n_548),
.Y(n_796)
);

AND2x4_ASAP7_75t_L g797 ( 
.A(n_661),
.B(n_662),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_L g798 ( 
.A(n_713),
.B(n_551),
.Y(n_798)
);

AND2x4_ASAP7_75t_L g799 ( 
.A(n_675),
.B(n_485),
.Y(n_799)
);

AND2x2_ASAP7_75t_L g800 ( 
.A(n_638),
.B(n_485),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_L g801 ( 
.A(n_714),
.B(n_561),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_L g802 ( 
.A(n_696),
.B(n_564),
.Y(n_802)
);

BUFx3_ASAP7_75t_L g803 ( 
.A(n_647),
.Y(n_803)
);

AOI22xp5_ASAP7_75t_L g804 ( 
.A1(n_610),
.A2(n_568),
.B1(n_571),
.B2(n_473),
.Y(n_804)
);

A2O1A1Ixp33_ASAP7_75t_L g805 ( 
.A1(n_638),
.A2(n_183),
.B(n_187),
.C(n_230),
.Y(n_805)
);

INVx5_ASAP7_75t_L g806 ( 
.A(n_670),
.Y(n_806)
);

INVx2_ASAP7_75t_L g807 ( 
.A(n_628),
.Y(n_807)
);

CKINVDCx5p33_ASAP7_75t_R g808 ( 
.A(n_722),
.Y(n_808)
);

OAI21xp5_ASAP7_75t_L g809 ( 
.A1(n_609),
.A2(n_571),
.B(n_568),
.Y(n_809)
);

INVx3_ASAP7_75t_L g810 ( 
.A(n_670),
.Y(n_810)
);

AOI21xp5_ASAP7_75t_L g811 ( 
.A1(n_606),
.A2(n_569),
.B(n_577),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_L g812 ( 
.A(n_696),
.B(n_475),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_SL g813 ( 
.A(n_587),
.B(n_475),
.Y(n_813)
);

OAI21xp5_ASAP7_75t_L g814 ( 
.A1(n_613),
.A2(n_484),
.B(n_539),
.Y(n_814)
);

AOI21xp5_ASAP7_75t_L g815 ( 
.A1(n_687),
.A2(n_569),
.B(n_577),
.Y(n_815)
);

INVx3_ASAP7_75t_L g816 ( 
.A(n_670),
.Y(n_816)
);

BUFx8_ASAP7_75t_L g817 ( 
.A(n_712),
.Y(n_817)
);

BUFx2_ASAP7_75t_L g818 ( 
.A(n_650),
.Y(n_818)
);

INVx2_ASAP7_75t_L g819 ( 
.A(n_631),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_SL g820 ( 
.A(n_590),
.B(n_475),
.Y(n_820)
);

INVx1_ASAP7_75t_L g821 ( 
.A(n_736),
.Y(n_821)
);

AOI22xp33_ASAP7_75t_L g822 ( 
.A1(n_668),
.A2(n_547),
.B1(n_537),
.B2(n_549),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_737),
.Y(n_823)
);

BUFx3_ASAP7_75t_L g824 ( 
.A(n_724),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_738),
.Y(n_825)
);

INVx8_ASAP7_75t_L g826 ( 
.A(n_691),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_L g827 ( 
.A(n_633),
.B(n_539),
.Y(n_827)
);

AND2x2_ASAP7_75t_L g828 ( 
.A(n_634),
.B(n_502),
.Y(n_828)
);

AND2x2_ASAP7_75t_SL g829 ( 
.A(n_708),
.B(n_574),
.Y(n_829)
);

AOI21xp5_ASAP7_75t_L g830 ( 
.A1(n_620),
.A2(n_577),
.B(n_565),
.Y(n_830)
);

INVx2_ASAP7_75t_L g831 ( 
.A(n_632),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_594),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_592),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_L g834 ( 
.A(n_640),
.B(n_539),
.Y(n_834)
);

INVx2_ASAP7_75t_L g835 ( 
.A(n_635),
.Y(n_835)
);

NOR3xp33_ASAP7_75t_SL g836 ( 
.A(n_695),
.B(n_230),
.C(n_260),
.Y(n_836)
);

OR2x2_ASAP7_75t_L g837 ( 
.A(n_634),
.B(n_502),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_SL g838 ( 
.A(n_618),
.B(n_484),
.Y(n_838)
);

INVx2_ASAP7_75t_L g839 ( 
.A(n_636),
.Y(n_839)
);

INVx2_ASAP7_75t_L g840 ( 
.A(n_637),
.Y(n_840)
);

CKINVDCx5p33_ASAP7_75t_R g841 ( 
.A(n_655),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_SL g842 ( 
.A(n_666),
.B(n_691),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_595),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_L g844 ( 
.A(n_686),
.B(n_565),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_681),
.Y(n_845)
);

AND2x4_ASAP7_75t_L g846 ( 
.A(n_678),
.B(n_484),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_L g847 ( 
.A(n_686),
.B(n_565),
.Y(n_847)
);

INVx1_ASAP7_75t_L g848 ( 
.A(n_741),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_742),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_SL g850 ( 
.A(n_691),
.B(n_577),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_L g851 ( 
.A(n_746),
.B(n_577),
.Y(n_851)
);

INVx2_ASAP7_75t_L g852 ( 
.A(n_641),
.Y(n_852)
);

INVxp67_ASAP7_75t_L g853 ( 
.A(n_600),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_744),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_L g855 ( 
.A(n_710),
.B(n_553),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_L g856 ( 
.A(n_716),
.B(n_553),
.Y(n_856)
);

INVx1_ASAP7_75t_L g857 ( 
.A(n_643),
.Y(n_857)
);

INVx2_ASAP7_75t_L g858 ( 
.A(n_644),
.Y(n_858)
);

INVx2_ASAP7_75t_L g859 ( 
.A(n_653),
.Y(n_859)
);

INVx2_ASAP7_75t_SL g860 ( 
.A(n_726),
.Y(n_860)
);

A2O1A1Ixp33_ASAP7_75t_L g861 ( 
.A1(n_659),
.A2(n_260),
.B(n_264),
.C(n_274),
.Y(n_861)
);

INVx3_ASAP7_75t_L g862 ( 
.A(n_691),
.Y(n_862)
);

AND2x4_ASAP7_75t_L g863 ( 
.A(n_727),
.B(n_559),
.Y(n_863)
);

AOI22xp33_ASAP7_75t_L g864 ( 
.A1(n_667),
.A2(n_556),
.B1(n_547),
.B2(n_567),
.Y(n_864)
);

INVx1_ASAP7_75t_L g865 ( 
.A(n_697),
.Y(n_865)
);

AND2x2_ASAP7_75t_SL g866 ( 
.A(n_708),
.B(n_574),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_711),
.Y(n_867)
);

CKINVDCx5p33_ASAP7_75t_R g868 ( 
.A(n_720),
.Y(n_868)
);

BUFx3_ASAP7_75t_L g869 ( 
.A(n_693),
.Y(n_869)
);

CKINVDCx20_ASAP7_75t_R g870 ( 
.A(n_703),
.Y(n_870)
);

CKINVDCx5p33_ASAP7_75t_R g871 ( 
.A(n_720),
.Y(n_871)
);

AOI22xp33_ASAP7_75t_SL g872 ( 
.A1(n_627),
.A2(n_274),
.B1(n_286),
.B2(n_291),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_SL g873 ( 
.A(n_693),
.B(n_584),
.Y(n_873)
);

AND3x1_ASAP7_75t_L g874 ( 
.A(n_659),
.B(n_700),
.C(n_721),
.Y(n_874)
);

AND2x4_ASAP7_75t_SL g875 ( 
.A(n_693),
.B(n_584),
.Y(n_875)
);

HB1xp67_ASAP7_75t_L g876 ( 
.A(n_645),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_L g877 ( 
.A(n_676),
.B(n_558),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_717),
.Y(n_878)
);

INVxp67_ASAP7_75t_L g879 ( 
.A(n_600),
.Y(n_879)
);

INVx2_ASAP7_75t_L g880 ( 
.A(n_731),
.Y(n_880)
);

INVx1_ASAP7_75t_L g881 ( 
.A(n_623),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_625),
.Y(n_882)
);

NAND2xp5_ASAP7_75t_SL g883 ( 
.A(n_693),
.B(n_732),
.Y(n_883)
);

AND2x2_ASAP7_75t_L g884 ( 
.A(n_733),
.B(n_286),
.Y(n_884)
);

OR2x6_ASAP7_75t_L g885 ( 
.A(n_734),
.B(n_559),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_630),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_651),
.Y(n_887)
);

INVx3_ASAP7_75t_L g888 ( 
.A(n_732),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_654),
.Y(n_889)
);

INVx2_ASAP7_75t_L g890 ( 
.A(n_730),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_L g891 ( 
.A(n_677),
.B(n_558),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_L g892 ( 
.A(n_684),
.B(n_556),
.Y(n_892)
);

INVx3_ASAP7_75t_L g893 ( 
.A(n_732),
.Y(n_893)
);

NAND2xp33_ASAP7_75t_L g894 ( 
.A(n_732),
.B(n_664),
.Y(n_894)
);

INVx1_ASAP7_75t_L g895 ( 
.A(n_660),
.Y(n_895)
);

INVx3_ASAP7_75t_L g896 ( 
.A(n_624),
.Y(n_896)
);

INVx2_ASAP7_75t_L g897 ( 
.A(n_730),
.Y(n_897)
);

AOI22xp33_ASAP7_75t_SL g898 ( 
.A1(n_689),
.A2(n_291),
.B1(n_567),
.B2(n_563),
.Y(n_898)
);

BUFx3_ASAP7_75t_L g899 ( 
.A(n_673),
.Y(n_899)
);

AOI22xp5_ASAP7_75t_L g900 ( 
.A1(n_704),
.A2(n_560),
.B1(n_549),
.B2(n_584),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_SL g901 ( 
.A(n_733),
.B(n_560),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_L g902 ( 
.A(n_698),
.B(n_465),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_L g903 ( 
.A(n_699),
.B(n_465),
.Y(n_903)
);

CKINVDCx20_ASAP7_75t_R g904 ( 
.A(n_727),
.Y(n_904)
);

OAI22xp5_ASAP7_75t_L g905 ( 
.A1(n_672),
.A2(n_465),
.B1(n_152),
.B2(n_149),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_645),
.Y(n_906)
);

HB1xp67_ASAP7_75t_L g907 ( 
.A(n_728),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_608),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_SL g909 ( 
.A(n_672),
.B(n_465),
.Y(n_909)
);

INVxp67_ASAP7_75t_L g910 ( 
.A(n_639),
.Y(n_910)
);

CKINVDCx16_ASAP7_75t_R g911 ( 
.A(n_652),
.Y(n_911)
);

CKINVDCx20_ASAP7_75t_R g912 ( 
.A(n_704),
.Y(n_912)
);

INVx2_ASAP7_75t_L g913 ( 
.A(n_725),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_SL g914 ( 
.A(n_614),
.B(n_465),
.Y(n_914)
);

INVx1_ASAP7_75t_L g915 ( 
.A(n_608),
.Y(n_915)
);

AOI22xp5_ASAP7_75t_L g916 ( 
.A1(n_709),
.A2(n_144),
.B1(n_136),
.B2(n_133),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_728),
.Y(n_917)
);

INVx2_ASAP7_75t_L g918 ( 
.A(n_624),
.Y(n_918)
);

HB1xp67_ASAP7_75t_L g919 ( 
.A(n_740),
.Y(n_919)
);

OR2x2_ASAP7_75t_SL g920 ( 
.A(n_589),
.B(n_0),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_740),
.Y(n_921)
);

AOI22xp5_ASAP7_75t_L g922 ( 
.A1(n_709),
.A2(n_124),
.B1(n_115),
.B2(n_114),
.Y(n_922)
);

AND2x4_ASAP7_75t_L g923 ( 
.A(n_715),
.B(n_109),
.Y(n_923)
);

O2A1O1Ixp5_ASAP7_75t_L g924 ( 
.A1(n_591),
.A2(n_102),
.B(n_97),
.C(n_90),
.Y(n_924)
);

INVx1_ASAP7_75t_L g925 ( 
.A(n_757),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_L g926 ( 
.A(n_773),
.B(n_639),
.Y(n_926)
);

NAND2xp5_ASAP7_75t_SL g927 ( 
.A(n_868),
.B(n_614),
.Y(n_927)
);

A2O1A1Ixp33_ASAP7_75t_L g928 ( 
.A1(n_910),
.A2(n_715),
.B(n_683),
.C(n_694),
.Y(n_928)
);

AND2x2_ASAP7_75t_L g929 ( 
.A(n_756),
.B(n_734),
.Y(n_929)
);

AND2x2_ASAP7_75t_L g930 ( 
.A(n_761),
.B(n_622),
.Y(n_930)
);

AOI21xp5_ASAP7_75t_L g931 ( 
.A1(n_760),
.A2(n_806),
.B(n_875),
.Y(n_931)
);

INVx1_ASAP7_75t_L g932 ( 
.A(n_770),
.Y(n_932)
);

BUFx12f_ASAP7_75t_L g933 ( 
.A(n_817),
.Y(n_933)
);

OR2x2_ASAP7_75t_L g934 ( 
.A(n_749),
.B(n_745),
.Y(n_934)
);

BUFx3_ASAP7_75t_L g935 ( 
.A(n_824),
.Y(n_935)
);

A2O1A1Ixp33_ASAP7_75t_L g936 ( 
.A1(n_763),
.A2(n_679),
.B(n_694),
.C(n_683),
.Y(n_936)
);

NAND2xp5_ASAP7_75t_L g937 ( 
.A(n_783),
.B(n_597),
.Y(n_937)
);

O2A1O1Ixp5_ASAP7_75t_L g938 ( 
.A1(n_764),
.A2(n_607),
.B(n_603),
.C(n_591),
.Y(n_938)
);

AND2x2_ASAP7_75t_L g939 ( 
.A(n_783),
.B(n_589),
.Y(n_939)
);

INVx3_ASAP7_75t_L g940 ( 
.A(n_781),
.Y(n_940)
);

AOI21xp5_ASAP7_75t_L g941 ( 
.A1(n_760),
.A2(n_688),
.B(n_658),
.Y(n_941)
);

HB1xp67_ASAP7_75t_L g942 ( 
.A(n_768),
.Y(n_942)
);

OAI22xp5_ASAP7_75t_L g943 ( 
.A1(n_871),
.A2(n_603),
.B1(n_674),
.B2(n_688),
.Y(n_943)
);

INVx1_ASAP7_75t_L g944 ( 
.A(n_774),
.Y(n_944)
);

NOR2xp33_ASAP7_75t_R g945 ( 
.A(n_808),
.B(n_89),
.Y(n_945)
);

NOR2xp33_ASAP7_75t_L g946 ( 
.A(n_853),
.B(n_679),
.Y(n_946)
);

OAI22xp5_ASAP7_75t_L g947 ( 
.A1(n_879),
.A2(n_607),
.B1(n_615),
.B2(n_617),
.Y(n_947)
);

AOI21xp5_ASAP7_75t_L g948 ( 
.A1(n_760),
.A2(n_806),
.B(n_875),
.Y(n_948)
);

INVx3_ASAP7_75t_L g949 ( 
.A(n_781),
.Y(n_949)
);

A2O1A1Ixp33_ASAP7_75t_SL g950 ( 
.A1(n_765),
.A2(n_729),
.B(n_669),
.C(n_629),
.Y(n_950)
);

INVx2_ASAP7_75t_L g951 ( 
.A(n_748),
.Y(n_951)
);

NOR2xp33_ASAP7_75t_L g952 ( 
.A(n_759),
.B(n_718),
.Y(n_952)
);

INVx2_ASAP7_75t_SL g953 ( 
.A(n_771),
.Y(n_953)
);

BUFx6f_ASAP7_75t_L g954 ( 
.A(n_826),
.Y(n_954)
);

BUFx3_ASAP7_75t_L g955 ( 
.A(n_824),
.Y(n_955)
);

BUFx2_ASAP7_75t_L g956 ( 
.A(n_904),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_SL g957 ( 
.A(n_906),
.B(n_617),
.Y(n_957)
);

O2A1O1Ixp33_ASAP7_75t_L g958 ( 
.A1(n_805),
.A2(n_702),
.B(n_743),
.C(n_745),
.Y(n_958)
);

NOR2xp33_ASAP7_75t_L g959 ( 
.A(n_786),
.B(n_692),
.Y(n_959)
);

AND2x2_ASAP7_75t_L g960 ( 
.A(n_884),
.B(n_589),
.Y(n_960)
);

NAND2xp5_ASAP7_75t_SL g961 ( 
.A(n_923),
.B(n_615),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_L g962 ( 
.A(n_833),
.B(n_743),
.Y(n_962)
);

OAI21xp5_ASAP7_75t_L g963 ( 
.A1(n_809),
.A2(n_649),
.B(n_646),
.Y(n_963)
);

OAI21x1_ASAP7_75t_SL g964 ( 
.A1(n_916),
.A2(n_61),
.B(n_54),
.Y(n_964)
);

INVx3_ASAP7_75t_L g965 ( 
.A(n_781),
.Y(n_965)
);

AND2x2_ASAP7_75t_L g966 ( 
.A(n_828),
.B(n_663),
.Y(n_966)
);

NAND2x1p5_ASAP7_75t_L g967 ( 
.A(n_790),
.B(n_6),
.Y(n_967)
);

O2A1O1Ixp5_ASAP7_75t_L g968 ( 
.A1(n_901),
.A2(n_9),
.B(n_10),
.C(n_12),
.Y(n_968)
);

HB1xp67_ASAP7_75t_L g969 ( 
.A(n_790),
.Y(n_969)
);

OAI21x1_ASAP7_75t_L g970 ( 
.A1(n_830),
.A2(n_10),
.B(n_12),
.Y(n_970)
);

BUFx6f_ASAP7_75t_L g971 ( 
.A(n_826),
.Y(n_971)
);

BUFx3_ASAP7_75t_L g972 ( 
.A(n_818),
.Y(n_972)
);

NAND2xp5_ASAP7_75t_SL g973 ( 
.A(n_923),
.B(n_15),
.Y(n_973)
);

NAND2xp5_ASAP7_75t_L g974 ( 
.A(n_843),
.B(n_15),
.Y(n_974)
);

O2A1O1Ixp33_ASAP7_75t_SL g975 ( 
.A1(n_861),
.A2(n_16),
.B(n_20),
.C(n_22),
.Y(n_975)
);

AOI21xp5_ASAP7_75t_L g976 ( 
.A1(n_760),
.A2(n_20),
.B(n_26),
.Y(n_976)
);

OR2x6_ASAP7_75t_SL g977 ( 
.A(n_841),
.B(n_26),
.Y(n_977)
);

INVx1_ASAP7_75t_L g978 ( 
.A(n_845),
.Y(n_978)
);

AOI221xp5_ASAP7_75t_L g979 ( 
.A1(n_861),
.A2(n_28),
.B1(n_29),
.B2(n_30),
.C(n_32),
.Y(n_979)
);

INVx4_ASAP7_75t_L g980 ( 
.A(n_790),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_SL g981 ( 
.A(n_790),
.B(n_28),
.Y(n_981)
);

AND2x6_ASAP7_75t_L g982 ( 
.A(n_908),
.B(n_33),
.Y(n_982)
);

INVx1_ASAP7_75t_L g983 ( 
.A(n_848),
.Y(n_983)
);

INVx3_ASAP7_75t_L g984 ( 
.A(n_826),
.Y(n_984)
);

NAND2xp5_ASAP7_75t_SL g985 ( 
.A(n_876),
.B(n_34),
.Y(n_985)
);

INVx2_ASAP7_75t_L g986 ( 
.A(n_748),
.Y(n_986)
);

A2O1A1Ixp33_ASAP7_75t_L g987 ( 
.A1(n_829),
.A2(n_35),
.B(n_36),
.C(n_37),
.Y(n_987)
);

NAND2xp5_ASAP7_75t_SL g988 ( 
.A(n_876),
.B(n_36),
.Y(n_988)
);

OR2x2_ASAP7_75t_L g989 ( 
.A(n_775),
.B(n_39),
.Y(n_989)
);

AOI21xp5_ASAP7_75t_L g990 ( 
.A1(n_806),
.A2(n_48),
.B(n_41),
.Y(n_990)
);

INVx1_ASAP7_75t_L g991 ( 
.A(n_849),
.Y(n_991)
);

A2O1A1Ixp33_ASAP7_75t_L g992 ( 
.A1(n_829),
.A2(n_39),
.B(n_43),
.C(n_45),
.Y(n_992)
);

NOR2xp33_ASAP7_75t_L g993 ( 
.A(n_837),
.B(n_45),
.Y(n_993)
);

AND2x2_ASAP7_75t_L g994 ( 
.A(n_800),
.B(n_48),
.Y(n_994)
);

NOR2xp33_ASAP7_75t_L g995 ( 
.A(n_758),
.B(n_784),
.Y(n_995)
);

AOI21xp5_ASAP7_75t_L g996 ( 
.A1(n_806),
.A2(n_896),
.B(n_838),
.Y(n_996)
);

O2A1O1Ixp33_ASAP7_75t_L g997 ( 
.A1(n_805),
.A2(n_907),
.B(n_919),
.C(n_917),
.Y(n_997)
);

NAND2x1p5_ASAP7_75t_L g998 ( 
.A(n_755),
.B(n_803),
.Y(n_998)
);

INVx5_ASAP7_75t_L g999 ( 
.A(n_896),
.Y(n_999)
);

NAND2xp5_ASAP7_75t_L g1000 ( 
.A(n_860),
.B(n_821),
.Y(n_1000)
);

AND2x2_ASAP7_75t_L g1001 ( 
.A(n_758),
.B(n_784),
.Y(n_1001)
);

BUFx3_ASAP7_75t_L g1002 ( 
.A(n_817),
.Y(n_1002)
);

AOI21xp5_ASAP7_75t_L g1003 ( 
.A1(n_838),
.A2(n_814),
.B(n_812),
.Y(n_1003)
);

INVx1_ASAP7_75t_SL g1004 ( 
.A(n_794),
.Y(n_1004)
);

A2O1A1Ixp33_ASAP7_75t_L g1005 ( 
.A1(n_866),
.A2(n_921),
.B(n_919),
.C(n_907),
.Y(n_1005)
);

INVx3_ASAP7_75t_L g1006 ( 
.A(n_787),
.Y(n_1006)
);

A2O1A1Ixp33_ASAP7_75t_L g1007 ( 
.A1(n_915),
.A2(n_866),
.B(n_823),
.C(n_825),
.Y(n_1007)
);

NOR2xp33_ASAP7_75t_L g1008 ( 
.A(n_870),
.B(n_904),
.Y(n_1008)
);

O2A1O1Ixp33_ASAP7_75t_L g1009 ( 
.A1(n_751),
.A2(n_901),
.B(n_885),
.C(n_832),
.Y(n_1009)
);

INVx3_ASAP7_75t_L g1010 ( 
.A(n_787),
.Y(n_1010)
);

NOR3xp33_ASAP7_75t_L g1011 ( 
.A(n_911),
.B(n_872),
.C(n_751),
.Y(n_1011)
);

INVx1_ASAP7_75t_L g1012 ( 
.A(n_854),
.Y(n_1012)
);

NAND2xp5_ASAP7_75t_L g1013 ( 
.A(n_899),
.B(n_881),
.Y(n_1013)
);

INVx1_ASAP7_75t_L g1014 ( 
.A(n_750),
.Y(n_1014)
);

OAI22xp5_ASAP7_75t_L g1015 ( 
.A1(n_780),
.A2(n_802),
.B1(n_844),
.B2(n_847),
.Y(n_1015)
);

AOI21xp5_ASAP7_75t_L g1016 ( 
.A1(n_811),
.A2(n_894),
.B(n_851),
.Y(n_1016)
);

INVx4_ASAP7_75t_L g1017 ( 
.A(n_755),
.Y(n_1017)
);

NAND2xp5_ASAP7_75t_L g1018 ( 
.A(n_882),
.B(n_886),
.Y(n_1018)
);

NAND2xp5_ASAP7_75t_L g1019 ( 
.A(n_887),
.B(n_889),
.Y(n_1019)
);

O2A1O1Ixp33_ASAP7_75t_L g1020 ( 
.A1(n_885),
.A2(n_905),
.B(n_753),
.C(n_836),
.Y(n_1020)
);

NOR2xp33_ASAP7_75t_L g1021 ( 
.A(n_912),
.B(n_885),
.Y(n_1021)
);

BUFx3_ASAP7_75t_L g1022 ( 
.A(n_803),
.Y(n_1022)
);

OR2x2_ASAP7_75t_L g1023 ( 
.A(n_782),
.B(n_797),
.Y(n_1023)
);

NAND3xp33_ASAP7_75t_SL g1024 ( 
.A(n_836),
.B(n_898),
.C(n_922),
.Y(n_1024)
);

NOR2xp33_ASAP7_75t_R g1025 ( 
.A(n_795),
.B(n_810),
.Y(n_1025)
);

INVx1_ASAP7_75t_L g1026 ( 
.A(n_782),
.Y(n_1026)
);

INVx3_ASAP7_75t_L g1027 ( 
.A(n_795),
.Y(n_1027)
);

INVx2_ASAP7_75t_L g1028 ( 
.A(n_762),
.Y(n_1028)
);

NAND2xp5_ASAP7_75t_L g1029 ( 
.A(n_895),
.B(n_797),
.Y(n_1029)
);

CKINVDCx14_ASAP7_75t_R g1030 ( 
.A(n_799),
.Y(n_1030)
);

BUFx2_ASAP7_75t_L g1031 ( 
.A(n_754),
.Y(n_1031)
);

OAI21xp33_ASAP7_75t_SL g1032 ( 
.A1(n_842),
.A2(n_855),
.B(n_766),
.Y(n_1032)
);

BUFx6f_ASAP7_75t_L g1033 ( 
.A(n_869),
.Y(n_1033)
);

AOI21xp5_ASAP7_75t_L g1034 ( 
.A1(n_856),
.A2(n_834),
.B(n_827),
.Y(n_1034)
);

A2O1A1Ixp33_ASAP7_75t_L g1035 ( 
.A1(n_752),
.A2(n_863),
.B(n_891),
.C(n_877),
.Y(n_1035)
);

NAND2xp5_ASAP7_75t_L g1036 ( 
.A(n_846),
.B(n_892),
.Y(n_1036)
);

INVxp67_ASAP7_75t_L g1037 ( 
.A(n_752),
.Y(n_1037)
);

INVx1_ASAP7_75t_L g1038 ( 
.A(n_769),
.Y(n_1038)
);

NAND2xp5_ASAP7_75t_L g1039 ( 
.A(n_766),
.B(n_788),
.Y(n_1039)
);

CKINVDCx20_ASAP7_75t_R g1040 ( 
.A(n_920),
.Y(n_1040)
);

BUFx2_ASAP7_75t_L g1041 ( 
.A(n_754),
.Y(n_1041)
);

AOI21xp5_ASAP7_75t_L g1042 ( 
.A1(n_902),
.A2(n_903),
.B(n_909),
.Y(n_1042)
);

O2A1O1Ixp33_ASAP7_75t_L g1043 ( 
.A1(n_842),
.A2(n_801),
.B(n_798),
.C(n_813),
.Y(n_1043)
);

OAI22xp5_ASAP7_75t_L g1044 ( 
.A1(n_767),
.A2(n_779),
.B1(n_791),
.B2(n_785),
.Y(n_1044)
);

NAND2xp5_ASAP7_75t_L g1045 ( 
.A(n_890),
.B(n_897),
.Y(n_1045)
);

AO22x1_ASAP7_75t_L g1046 ( 
.A1(n_799),
.A2(n_874),
.B1(n_878),
.B2(n_857),
.Y(n_1046)
);

INVx2_ASAP7_75t_L g1047 ( 
.A(n_769),
.Y(n_1047)
);

NAND2xp5_ASAP7_75t_L g1048 ( 
.A(n_890),
.B(n_897),
.Y(n_1048)
);

AOI21xp5_ASAP7_75t_L g1049 ( 
.A1(n_909),
.A2(n_815),
.B(n_820),
.Y(n_1049)
);

INVx2_ASAP7_75t_L g1050 ( 
.A(n_776),
.Y(n_1050)
);

INVx2_ASAP7_75t_L g1051 ( 
.A(n_776),
.Y(n_1051)
);

NOR2x1p5_ASAP7_75t_L g1052 ( 
.A(n_869),
.B(n_865),
.Y(n_1052)
);

NAND2xp5_ASAP7_75t_SL g1053 ( 
.A(n_918),
.B(n_840),
.Y(n_1053)
);

INVx2_ASAP7_75t_L g1054 ( 
.A(n_777),
.Y(n_1054)
);

INVx2_ASAP7_75t_L g1055 ( 
.A(n_777),
.Y(n_1055)
);

OAI21xp5_ASAP7_75t_L g1056 ( 
.A1(n_938),
.A2(n_813),
.B(n_820),
.Y(n_1056)
);

AO31x2_ASAP7_75t_L g1057 ( 
.A1(n_1005),
.A2(n_913),
.A3(n_918),
.B(n_789),
.Y(n_1057)
);

OAI22xp5_ASAP7_75t_L g1058 ( 
.A1(n_995),
.A2(n_792),
.B1(n_883),
.B2(n_914),
.Y(n_1058)
);

INVx1_ASAP7_75t_L g1059 ( 
.A(n_925),
.Y(n_1059)
);

INVxp67_ASAP7_75t_L g1060 ( 
.A(n_942),
.Y(n_1060)
);

OAI21xp5_ASAP7_75t_L g1061 ( 
.A1(n_938),
.A2(n_864),
.B(n_913),
.Y(n_1061)
);

INVx1_ASAP7_75t_L g1062 ( 
.A(n_932),
.Y(n_1062)
);

BUFx2_ASAP7_75t_L g1063 ( 
.A(n_942),
.Y(n_1063)
);

CKINVDCx11_ASAP7_75t_R g1064 ( 
.A(n_933),
.Y(n_1064)
);

AOI221x1_ASAP7_75t_L g1065 ( 
.A1(n_1024),
.A2(n_867),
.B1(n_862),
.B2(n_816),
.C(n_893),
.Y(n_1065)
);

BUFx10_ASAP7_75t_L g1066 ( 
.A(n_1008),
.Y(n_1066)
);

OAI22x1_ASAP7_75t_L g1067 ( 
.A1(n_973),
.A2(n_914),
.B1(n_778),
.B2(n_883),
.Y(n_1067)
);

AOI22xp5_ASAP7_75t_L g1068 ( 
.A1(n_929),
.A2(n_864),
.B1(n_789),
.B2(n_880),
.Y(n_1068)
);

HB1xp67_ASAP7_75t_L g1069 ( 
.A(n_953),
.Y(n_1069)
);

HB1xp67_ASAP7_75t_L g1070 ( 
.A(n_1023),
.Y(n_1070)
);

XOR2xp5_ASAP7_75t_L g1071 ( 
.A(n_1030),
.B(n_792),
.Y(n_1071)
);

NAND2xp5_ASAP7_75t_L g1072 ( 
.A(n_926),
.B(n_839),
.Y(n_1072)
);

NAND2xp5_ASAP7_75t_L g1073 ( 
.A(n_995),
.B(n_839),
.Y(n_1073)
);

O2A1O1Ixp5_ASAP7_75t_SL g1074 ( 
.A1(n_985),
.A2(n_796),
.B(n_873),
.C(n_850),
.Y(n_1074)
);

HB1xp67_ASAP7_75t_L g1075 ( 
.A(n_1004),
.Y(n_1075)
);

OAI21x1_ASAP7_75t_L g1076 ( 
.A1(n_1049),
.A2(n_796),
.B(n_772),
.Y(n_1076)
);

INVx4_ASAP7_75t_L g1077 ( 
.A(n_954),
.Y(n_1077)
);

AOI21xp5_ASAP7_75t_L g1078 ( 
.A1(n_1034),
.A2(n_850),
.B(n_873),
.Y(n_1078)
);

OAI21x1_ASAP7_75t_L g1079 ( 
.A1(n_1016),
.A2(n_772),
.B(n_804),
.Y(n_1079)
);

BUFx8_ASAP7_75t_SL g1080 ( 
.A(n_935),
.Y(n_1080)
);

INVx4_ASAP7_75t_L g1081 ( 
.A(n_954),
.Y(n_1081)
);

INVx6_ASAP7_75t_L g1082 ( 
.A(n_955),
.Y(n_1082)
);

A2O1A1Ixp33_ASAP7_75t_L g1083 ( 
.A1(n_936),
.A2(n_924),
.B(n_900),
.C(n_793),
.Y(n_1083)
);

NAND2xp5_ASAP7_75t_L g1084 ( 
.A(n_1001),
.B(n_793),
.Y(n_1084)
);

INVxp67_ASAP7_75t_L g1085 ( 
.A(n_956),
.Y(n_1085)
);

INVx1_ASAP7_75t_L g1086 ( 
.A(n_944),
.Y(n_1086)
);

OAI21x1_ASAP7_75t_L g1087 ( 
.A1(n_996),
.A2(n_822),
.B(n_840),
.Y(n_1087)
);

NOR2xp33_ASAP7_75t_L g1088 ( 
.A(n_1000),
.B(n_946),
.Y(n_1088)
);

NAND2xp5_ASAP7_75t_L g1089 ( 
.A(n_946),
.B(n_807),
.Y(n_1089)
);

CKINVDCx11_ASAP7_75t_R g1090 ( 
.A(n_977),
.Y(n_1090)
);

NAND2xp5_ASAP7_75t_L g1091 ( 
.A(n_1018),
.B(n_852),
.Y(n_1091)
);

OA21x2_ASAP7_75t_L g1092 ( 
.A1(n_1005),
.A2(n_822),
.B(n_880),
.Y(n_1092)
);

AOI221x1_ASAP7_75t_L g1093 ( 
.A1(n_1024),
.A2(n_810),
.B1(n_816),
.B2(n_888),
.C(n_893),
.Y(n_1093)
);

OAI21x1_ASAP7_75t_L g1094 ( 
.A1(n_1042),
.A2(n_819),
.B(n_831),
.Y(n_1094)
);

AOI21x1_ASAP7_75t_SL g1095 ( 
.A1(n_974),
.A2(n_888),
.B(n_831),
.Y(n_1095)
);

AND2x2_ASAP7_75t_L g1096 ( 
.A(n_930),
.B(n_939),
.Y(n_1096)
);

NAND2xp5_ASAP7_75t_L g1097 ( 
.A(n_1019),
.B(n_819),
.Y(n_1097)
);

O2A1O1Ixp5_ASAP7_75t_L g1098 ( 
.A1(n_1046),
.A2(n_927),
.B(n_1015),
.C(n_943),
.Y(n_1098)
);

A2O1A1Ixp33_ASAP7_75t_L g1099 ( 
.A1(n_928),
.A2(n_835),
.B(n_852),
.C(n_858),
.Y(n_1099)
);

AOI21xp5_ASAP7_75t_L g1100 ( 
.A1(n_1003),
.A2(n_835),
.B(n_858),
.Y(n_1100)
);

OAI21xp5_ASAP7_75t_L g1101 ( 
.A1(n_1007),
.A2(n_859),
.B(n_1032),
.Y(n_1101)
);

NAND3x1_ASAP7_75t_L g1102 ( 
.A(n_1011),
.B(n_993),
.C(n_1021),
.Y(n_1102)
);

XOR2xp5_ASAP7_75t_L g1103 ( 
.A(n_1040),
.B(n_859),
.Y(n_1103)
);

AND2x2_ASAP7_75t_L g1104 ( 
.A(n_960),
.B(n_966),
.Y(n_1104)
);

AOI21xp5_ASAP7_75t_L g1105 ( 
.A1(n_961),
.A2(n_999),
.B(n_1043),
.Y(n_1105)
);

NAND2xp5_ASAP7_75t_L g1106 ( 
.A(n_934),
.B(n_1029),
.Y(n_1106)
);

OAI22x1_ASAP7_75t_L g1107 ( 
.A1(n_973),
.A2(n_993),
.B1(n_1021),
.B2(n_988),
.Y(n_1107)
);

OAI21xp5_ASAP7_75t_L g1108 ( 
.A1(n_1035),
.A2(n_1044),
.B(n_958),
.Y(n_1108)
);

INVx4_ASAP7_75t_L g1109 ( 
.A(n_954),
.Y(n_1109)
);

A2O1A1Ixp33_ASAP7_75t_L g1110 ( 
.A1(n_997),
.A2(n_1009),
.B(n_952),
.C(n_959),
.Y(n_1110)
);

AOI21x1_ASAP7_75t_L g1111 ( 
.A1(n_947),
.A2(n_927),
.B(n_957),
.Y(n_1111)
);

OAI22xp5_ASAP7_75t_L g1112 ( 
.A1(n_1039),
.A2(n_1013),
.B1(n_961),
.B2(n_1037),
.Y(n_1112)
);

INVx1_ASAP7_75t_L g1113 ( 
.A(n_978),
.Y(n_1113)
);

BUFx6f_ASAP7_75t_L g1114 ( 
.A(n_971),
.Y(n_1114)
);

OAI21xp5_ASAP7_75t_SL g1115 ( 
.A1(n_979),
.A2(n_1011),
.B(n_992),
.Y(n_1115)
);

OAI21x1_ASAP7_75t_L g1116 ( 
.A1(n_963),
.A2(n_1045),
.B(n_1048),
.Y(n_1116)
);

INVx1_ASAP7_75t_L g1117 ( 
.A(n_983),
.Y(n_1117)
);

AOI21xp33_ASAP7_75t_L g1118 ( 
.A1(n_952),
.A2(n_959),
.B(n_937),
.Y(n_1118)
);

OAI21x1_ASAP7_75t_L g1119 ( 
.A1(n_970),
.A2(n_941),
.B(n_1053),
.Y(n_1119)
);

INVx1_ASAP7_75t_L g1120 ( 
.A(n_991),
.Y(n_1120)
);

OAI21xp5_ASAP7_75t_L g1121 ( 
.A1(n_950),
.A2(n_1020),
.B(n_1036),
.Y(n_1121)
);

OAI21xp5_ASAP7_75t_L g1122 ( 
.A1(n_950),
.A2(n_962),
.B(n_968),
.Y(n_1122)
);

INVxp67_ASAP7_75t_L g1123 ( 
.A(n_989),
.Y(n_1123)
);

AOI21xp5_ASAP7_75t_L g1124 ( 
.A1(n_999),
.A2(n_931),
.B(n_948),
.Y(n_1124)
);

OA21x2_ASAP7_75t_L g1125 ( 
.A1(n_968),
.A2(n_1053),
.B(n_987),
.Y(n_1125)
);

INVx1_ASAP7_75t_L g1126 ( 
.A(n_1012),
.Y(n_1126)
);

A2O1A1Ixp33_ASAP7_75t_L g1127 ( 
.A1(n_994),
.A2(n_992),
.B(n_987),
.C(n_1026),
.Y(n_1127)
);

BUFx6f_ASAP7_75t_L g1128 ( 
.A(n_971),
.Y(n_1128)
);

AOI221x1_ASAP7_75t_L g1129 ( 
.A1(n_964),
.A2(n_976),
.B1(n_990),
.B2(n_1014),
.C(n_1038),
.Y(n_1129)
);

AOI21xp5_ASAP7_75t_L g1130 ( 
.A1(n_1047),
.A2(n_1055),
.B(n_1054),
.Y(n_1130)
);

AOI21xp5_ASAP7_75t_L g1131 ( 
.A1(n_1050),
.A2(n_1051),
.B(n_969),
.Y(n_1131)
);

NAND2xp5_ASAP7_75t_L g1132 ( 
.A(n_1031),
.B(n_1041),
.Y(n_1132)
);

AO32x2_ASAP7_75t_L g1133 ( 
.A1(n_980),
.A2(n_975),
.A3(n_1017),
.B1(n_982),
.B2(n_981),
.Y(n_1133)
);

AOI21xp5_ASAP7_75t_L g1134 ( 
.A1(n_969),
.A2(n_1027),
.B(n_1006),
.Y(n_1134)
);

INVx3_ASAP7_75t_L g1135 ( 
.A(n_971),
.Y(n_1135)
);

AOI21xp5_ASAP7_75t_L g1136 ( 
.A1(n_1006),
.A2(n_1027),
.B(n_1010),
.Y(n_1136)
);

OAI21x1_ASAP7_75t_L g1137 ( 
.A1(n_951),
.A2(n_986),
.B(n_1028),
.Y(n_1137)
);

INVx1_ASAP7_75t_SL g1138 ( 
.A(n_972),
.Y(n_1138)
);

NOR2xp33_ASAP7_75t_L g1139 ( 
.A(n_1017),
.B(n_1022),
.Y(n_1139)
);

NAND2xp5_ASAP7_75t_L g1140 ( 
.A(n_1052),
.B(n_1033),
.Y(n_1140)
);

AOI21xp5_ASAP7_75t_L g1141 ( 
.A1(n_1010),
.A2(n_980),
.B(n_949),
.Y(n_1141)
);

NAND2xp5_ASAP7_75t_L g1142 ( 
.A(n_1033),
.B(n_940),
.Y(n_1142)
);

NAND2xp5_ASAP7_75t_L g1143 ( 
.A(n_1033),
.B(n_940),
.Y(n_1143)
);

NOR2xp67_ASAP7_75t_L g1144 ( 
.A(n_984),
.B(n_949),
.Y(n_1144)
);

NOR2xp33_ASAP7_75t_L g1145 ( 
.A(n_1033),
.B(n_998),
.Y(n_1145)
);

NAND2xp5_ASAP7_75t_SL g1146 ( 
.A(n_971),
.B(n_945),
.Y(n_1146)
);

NOR2xp33_ASAP7_75t_L g1147 ( 
.A(n_998),
.B(n_965),
.Y(n_1147)
);

INVx6_ASAP7_75t_SL g1148 ( 
.A(n_1002),
.Y(n_1148)
);

NAND2xp5_ASAP7_75t_L g1149 ( 
.A(n_965),
.B(n_982),
.Y(n_1149)
);

BUFx6f_ASAP7_75t_L g1150 ( 
.A(n_982),
.Y(n_1150)
);

AOI21xp5_ASAP7_75t_L g1151 ( 
.A1(n_975),
.A2(n_967),
.B(n_1025),
.Y(n_1151)
);

OR2x2_ASAP7_75t_L g1152 ( 
.A(n_967),
.B(n_945),
.Y(n_1152)
);

NAND2xp5_ASAP7_75t_L g1153 ( 
.A(n_982),
.B(n_1025),
.Y(n_1153)
);

AO31x2_ASAP7_75t_L g1154 ( 
.A1(n_982),
.A2(n_1005),
.A3(n_1007),
.B(n_1015),
.Y(n_1154)
);

BUFx3_ASAP7_75t_L g1155 ( 
.A(n_935),
.Y(n_1155)
);

NAND2xp5_ASAP7_75t_SL g1156 ( 
.A(n_926),
.B(n_868),
.Y(n_1156)
);

INVx1_ASAP7_75t_L g1157 ( 
.A(n_925),
.Y(n_1157)
);

AOI21xp5_ASAP7_75t_L g1158 ( 
.A1(n_1034),
.A2(n_1016),
.B(n_1015),
.Y(n_1158)
);

OAI21x1_ASAP7_75t_L g1159 ( 
.A1(n_1049),
.A2(n_1016),
.B(n_830),
.Y(n_1159)
);

AO31x2_ASAP7_75t_L g1160 ( 
.A1(n_1005),
.A2(n_1007),
.A3(n_1015),
.B(n_1042),
.Y(n_1160)
);

INVx1_ASAP7_75t_L g1161 ( 
.A(n_925),
.Y(n_1161)
);

NAND2xp5_ASAP7_75t_L g1162 ( 
.A(n_926),
.B(n_995),
.Y(n_1162)
);

INVx2_ASAP7_75t_L g1163 ( 
.A(n_1047),
.Y(n_1163)
);

INVx1_ASAP7_75t_L g1164 ( 
.A(n_925),
.Y(n_1164)
);

BUFx6f_ASAP7_75t_L g1165 ( 
.A(n_954),
.Y(n_1165)
);

AND2x4_ASAP7_75t_L g1166 ( 
.A(n_1026),
.B(n_1052),
.Y(n_1166)
);

AND2x2_ASAP7_75t_L g1167 ( 
.A(n_929),
.B(n_756),
.Y(n_1167)
);

AO21x1_ASAP7_75t_L g1168 ( 
.A1(n_995),
.A2(n_1009),
.B(n_1044),
.Y(n_1168)
);

AOI21xp5_ASAP7_75t_SL g1169 ( 
.A1(n_1035),
.A2(n_995),
.B(n_1007),
.Y(n_1169)
);

OAI21x1_ASAP7_75t_L g1170 ( 
.A1(n_1049),
.A2(n_1016),
.B(n_830),
.Y(n_1170)
);

INVx1_ASAP7_75t_L g1171 ( 
.A(n_925),
.Y(n_1171)
);

AND2x4_ASAP7_75t_L g1172 ( 
.A(n_1026),
.B(n_1052),
.Y(n_1172)
);

NAND2xp5_ASAP7_75t_L g1173 ( 
.A(n_926),
.B(n_995),
.Y(n_1173)
);

NAND2xp5_ASAP7_75t_L g1174 ( 
.A(n_926),
.B(n_995),
.Y(n_1174)
);

AO31x2_ASAP7_75t_L g1175 ( 
.A1(n_1005),
.A2(n_1007),
.A3(n_1015),
.B(n_1042),
.Y(n_1175)
);

BUFx6f_ASAP7_75t_SL g1176 ( 
.A(n_935),
.Y(n_1176)
);

OAI21xp5_ASAP7_75t_L g1177 ( 
.A1(n_938),
.A2(n_1007),
.B(n_1003),
.Y(n_1177)
);

CKINVDCx5p33_ASAP7_75t_R g1178 ( 
.A(n_933),
.Y(n_1178)
);

OAI21x1_ASAP7_75t_L g1179 ( 
.A1(n_1049),
.A2(n_1016),
.B(n_830),
.Y(n_1179)
);

NAND2xp5_ASAP7_75t_L g1180 ( 
.A(n_926),
.B(n_995),
.Y(n_1180)
);

INVx2_ASAP7_75t_L g1181 ( 
.A(n_1047),
.Y(n_1181)
);

INVx2_ASAP7_75t_L g1182 ( 
.A(n_1047),
.Y(n_1182)
);

A2O1A1Ixp33_ASAP7_75t_L g1183 ( 
.A1(n_926),
.A2(n_910),
.B(n_936),
.C(n_995),
.Y(n_1183)
);

AOI21xp5_ASAP7_75t_L g1184 ( 
.A1(n_1034),
.A2(n_1016),
.B(n_1015),
.Y(n_1184)
);

OAI21x1_ASAP7_75t_L g1185 ( 
.A1(n_1049),
.A2(n_1016),
.B(n_830),
.Y(n_1185)
);

AOI21xp5_ASAP7_75t_L g1186 ( 
.A1(n_1034),
.A2(n_1016),
.B(n_1015),
.Y(n_1186)
);

OAI21xp5_ASAP7_75t_L g1187 ( 
.A1(n_938),
.A2(n_1007),
.B(n_1003),
.Y(n_1187)
);

BUFx8_ASAP7_75t_L g1188 ( 
.A(n_1176),
.Y(n_1188)
);

NOR2xp67_ASAP7_75t_L g1189 ( 
.A(n_1075),
.B(n_1070),
.Y(n_1189)
);

OAI21x1_ASAP7_75t_L g1190 ( 
.A1(n_1119),
.A2(n_1100),
.B(n_1094),
.Y(n_1190)
);

AOI221xp5_ASAP7_75t_L g1191 ( 
.A1(n_1118),
.A2(n_1115),
.B1(n_1110),
.B2(n_1107),
.C(n_1108),
.Y(n_1191)
);

OA21x2_ASAP7_75t_L g1192 ( 
.A1(n_1177),
.A2(n_1187),
.B(n_1184),
.Y(n_1192)
);

OAI21x1_ASAP7_75t_L g1193 ( 
.A1(n_1159),
.A2(n_1179),
.B(n_1170),
.Y(n_1193)
);

NOR2xp33_ASAP7_75t_L g1194 ( 
.A(n_1162),
.B(n_1173),
.Y(n_1194)
);

NAND2xp5_ASAP7_75t_L g1195 ( 
.A(n_1174),
.B(n_1180),
.Y(n_1195)
);

BUFx2_ASAP7_75t_L g1196 ( 
.A(n_1063),
.Y(n_1196)
);

AOI22xp33_ASAP7_75t_L g1197 ( 
.A1(n_1168),
.A2(n_1108),
.B1(n_1167),
.B2(n_1088),
.Y(n_1197)
);

OAI22xp33_ASAP7_75t_L g1198 ( 
.A1(n_1115),
.A2(n_1106),
.B1(n_1123),
.B2(n_1073),
.Y(n_1198)
);

OAI21x1_ASAP7_75t_L g1199 ( 
.A1(n_1185),
.A2(n_1079),
.B(n_1076),
.Y(n_1199)
);

AND2x2_ASAP7_75t_L g1200 ( 
.A(n_1096),
.B(n_1104),
.Y(n_1200)
);

AO21x2_ASAP7_75t_L g1201 ( 
.A1(n_1122),
.A2(n_1187),
.B(n_1177),
.Y(n_1201)
);

BUFx2_ASAP7_75t_L g1202 ( 
.A(n_1069),
.Y(n_1202)
);

NOR2xp33_ASAP7_75t_L g1203 ( 
.A(n_1156),
.B(n_1085),
.Y(n_1203)
);

NOR3xp33_ASAP7_75t_L g1204 ( 
.A(n_1098),
.B(n_1183),
.C(n_1127),
.Y(n_1204)
);

OA21x2_ASAP7_75t_L g1205 ( 
.A1(n_1121),
.A2(n_1122),
.B(n_1065),
.Y(n_1205)
);

NOR2xp33_ASAP7_75t_L g1206 ( 
.A(n_1060),
.B(n_1112),
.Y(n_1206)
);

INVx2_ASAP7_75t_L g1207 ( 
.A(n_1137),
.Y(n_1207)
);

OAI21x1_ASAP7_75t_L g1208 ( 
.A1(n_1078),
.A2(n_1095),
.B(n_1087),
.Y(n_1208)
);

BUFx6f_ASAP7_75t_L g1209 ( 
.A(n_1114),
.Y(n_1209)
);

OAI21x1_ASAP7_75t_L g1210 ( 
.A1(n_1116),
.A2(n_1105),
.B(n_1056),
.Y(n_1210)
);

INVx1_ASAP7_75t_L g1211 ( 
.A(n_1062),
.Y(n_1211)
);

OAI21x1_ASAP7_75t_L g1212 ( 
.A1(n_1056),
.A2(n_1124),
.B(n_1061),
.Y(n_1212)
);

OR2x2_ASAP7_75t_L g1213 ( 
.A(n_1132),
.B(n_1089),
.Y(n_1213)
);

NAND2xp5_ASAP7_75t_L g1214 ( 
.A(n_1084),
.B(n_1072),
.Y(n_1214)
);

BUFx3_ASAP7_75t_L g1215 ( 
.A(n_1082),
.Y(n_1215)
);

BUFx2_ASAP7_75t_R g1216 ( 
.A(n_1080),
.Y(n_1216)
);

OAI21x1_ASAP7_75t_L g1217 ( 
.A1(n_1061),
.A2(n_1101),
.B(n_1111),
.Y(n_1217)
);

AO31x2_ASAP7_75t_L g1218 ( 
.A1(n_1093),
.A2(n_1083),
.A3(n_1129),
.B(n_1067),
.Y(n_1218)
);

INVxp67_ASAP7_75t_L g1219 ( 
.A(n_1086),
.Y(n_1219)
);

INVx2_ASAP7_75t_SL g1220 ( 
.A(n_1082),
.Y(n_1220)
);

AO21x2_ASAP7_75t_L g1221 ( 
.A1(n_1121),
.A2(n_1101),
.B(n_1169),
.Y(n_1221)
);

O2A1O1Ixp33_ASAP7_75t_L g1222 ( 
.A1(n_1099),
.A2(n_1058),
.B(n_1151),
.C(n_1091),
.Y(n_1222)
);

NOR2xp33_ASAP7_75t_L g1223 ( 
.A(n_1152),
.B(n_1066),
.Y(n_1223)
);

INVx2_ASAP7_75t_L g1224 ( 
.A(n_1057),
.Y(n_1224)
);

BUFx6f_ASAP7_75t_L g1225 ( 
.A(n_1114),
.Y(n_1225)
);

INVx1_ASAP7_75t_L g1226 ( 
.A(n_1113),
.Y(n_1226)
);

OR2x2_ASAP7_75t_L g1227 ( 
.A(n_1117),
.B(n_1120),
.Y(n_1227)
);

AND2x6_ASAP7_75t_L g1228 ( 
.A(n_1150),
.B(n_1068),
.Y(n_1228)
);

OR2x2_ASAP7_75t_L g1229 ( 
.A(n_1126),
.B(n_1157),
.Y(n_1229)
);

AOI211xp5_ASAP7_75t_L g1230 ( 
.A1(n_1138),
.A2(n_1102),
.B(n_1166),
.C(n_1172),
.Y(n_1230)
);

OAI21x1_ASAP7_75t_L g1231 ( 
.A1(n_1074),
.A2(n_1131),
.B(n_1149),
.Y(n_1231)
);

BUFx2_ASAP7_75t_L g1232 ( 
.A(n_1155),
.Y(n_1232)
);

OAI21x1_ASAP7_75t_L g1233 ( 
.A1(n_1136),
.A2(n_1130),
.B(n_1134),
.Y(n_1233)
);

AO21x2_ASAP7_75t_L g1234 ( 
.A1(n_1068),
.A2(n_1153),
.B(n_1141),
.Y(n_1234)
);

INVx1_ASAP7_75t_L g1235 ( 
.A(n_1161),
.Y(n_1235)
);

O2A1O1Ixp33_ASAP7_75t_L g1236 ( 
.A1(n_1097),
.A2(n_1146),
.B(n_1164),
.C(n_1171),
.Y(n_1236)
);

OAI21x1_ASAP7_75t_L g1237 ( 
.A1(n_1092),
.A2(n_1125),
.B(n_1181),
.Y(n_1237)
);

OAI21x1_ASAP7_75t_L g1238 ( 
.A1(n_1163),
.A2(n_1182),
.B(n_1142),
.Y(n_1238)
);

OAI22xp33_ASAP7_75t_L g1239 ( 
.A1(n_1150),
.A2(n_1140),
.B1(n_1138),
.B2(n_1143),
.Y(n_1239)
);

OAI22xp5_ASAP7_75t_L g1240 ( 
.A1(n_1103),
.A2(n_1071),
.B1(n_1139),
.B2(n_1150),
.Y(n_1240)
);

AO21x2_ASAP7_75t_L g1241 ( 
.A1(n_1144),
.A2(n_1057),
.B(n_1175),
.Y(n_1241)
);

AND2x4_ASAP7_75t_L g1242 ( 
.A(n_1135),
.B(n_1109),
.Y(n_1242)
);

BUFx3_ASAP7_75t_L g1243 ( 
.A(n_1114),
.Y(n_1243)
);

OAI21x1_ASAP7_75t_L g1244 ( 
.A1(n_1135),
.A2(n_1147),
.B(n_1145),
.Y(n_1244)
);

AO21x2_ASAP7_75t_L g1245 ( 
.A1(n_1057),
.A2(n_1175),
.B(n_1160),
.Y(n_1245)
);

OAI21x1_ASAP7_75t_L g1246 ( 
.A1(n_1160),
.A2(n_1175),
.B(n_1154),
.Y(n_1246)
);

O2A1O1Ixp33_ASAP7_75t_SL g1247 ( 
.A1(n_1133),
.A2(n_1154),
.B(n_1160),
.C(n_1081),
.Y(n_1247)
);

O2A1O1Ixp33_ASAP7_75t_L g1248 ( 
.A1(n_1133),
.A2(n_1154),
.B(n_1176),
.C(n_1090),
.Y(n_1248)
);

AO21x2_ASAP7_75t_L g1249 ( 
.A1(n_1133),
.A2(n_1077),
.B(n_1081),
.Y(n_1249)
);

OAI21xp5_ASAP7_75t_L g1250 ( 
.A1(n_1077),
.A2(n_1109),
.B(n_1178),
.Y(n_1250)
);

AOI22xp33_ASAP7_75t_SL g1251 ( 
.A1(n_1128),
.A2(n_1165),
.B1(n_1064),
.B2(n_1148),
.Y(n_1251)
);

NAND2x1p5_ASAP7_75t_L g1252 ( 
.A(n_1128),
.B(n_1165),
.Y(n_1252)
);

OAI21x1_ASAP7_75t_L g1253 ( 
.A1(n_1128),
.A2(n_1165),
.B(n_1148),
.Y(n_1253)
);

AOI22xp5_ASAP7_75t_L g1254 ( 
.A1(n_1156),
.A2(n_871),
.B1(n_868),
.B2(n_874),
.Y(n_1254)
);

AND2x4_ASAP7_75t_L g1255 ( 
.A(n_1166),
.B(n_1172),
.Y(n_1255)
);

INVx2_ASAP7_75t_L g1256 ( 
.A(n_1137),
.Y(n_1256)
);

OAI21xp5_ASAP7_75t_L g1257 ( 
.A1(n_1110),
.A2(n_910),
.B(n_926),
.Y(n_1257)
);

AOI21xp5_ASAP7_75t_L g1258 ( 
.A1(n_1158),
.A2(n_1186),
.B(n_1184),
.Y(n_1258)
);

AOI22xp33_ASAP7_75t_L g1259 ( 
.A1(n_1118),
.A2(n_979),
.B1(n_871),
.B2(n_868),
.Y(n_1259)
);

OAI21x1_ASAP7_75t_L g1260 ( 
.A1(n_1119),
.A2(n_1100),
.B(n_1094),
.Y(n_1260)
);

INVx1_ASAP7_75t_L g1261 ( 
.A(n_1059),
.Y(n_1261)
);

AOI21xp5_ASAP7_75t_L g1262 ( 
.A1(n_1158),
.A2(n_1186),
.B(n_1184),
.Y(n_1262)
);

NAND3xp33_ASAP7_75t_L g1263 ( 
.A(n_1110),
.B(n_871),
.C(n_868),
.Y(n_1263)
);

OAI21x1_ASAP7_75t_L g1264 ( 
.A1(n_1119),
.A2(n_1100),
.B(n_1094),
.Y(n_1264)
);

AND2x4_ASAP7_75t_L g1265 ( 
.A(n_1166),
.B(n_1172),
.Y(n_1265)
);

INVx1_ASAP7_75t_L g1266 ( 
.A(n_1059),
.Y(n_1266)
);

INVx2_ASAP7_75t_L g1267 ( 
.A(n_1137),
.Y(n_1267)
);

OAI22xp33_ASAP7_75t_L g1268 ( 
.A1(n_1115),
.A2(n_871),
.B1(n_868),
.B2(n_1162),
.Y(n_1268)
);

INVx1_ASAP7_75t_L g1269 ( 
.A(n_1059),
.Y(n_1269)
);

AND2x6_ASAP7_75t_L g1270 ( 
.A(n_1150),
.B(n_1068),
.Y(n_1270)
);

OAI21x1_ASAP7_75t_L g1271 ( 
.A1(n_1119),
.A2(n_1100),
.B(n_1094),
.Y(n_1271)
);

INVx1_ASAP7_75t_L g1272 ( 
.A(n_1059),
.Y(n_1272)
);

NOR2xp33_ASAP7_75t_L g1273 ( 
.A(n_1162),
.B(n_1173),
.Y(n_1273)
);

BUFx2_ASAP7_75t_L g1274 ( 
.A(n_1075),
.Y(n_1274)
);

OAI21x1_ASAP7_75t_SL g1275 ( 
.A1(n_1151),
.A2(n_1009),
.B(n_997),
.Y(n_1275)
);

NAND3xp33_ASAP7_75t_L g1276 ( 
.A(n_1110),
.B(n_871),
.C(n_868),
.Y(n_1276)
);

BUFx6f_ASAP7_75t_L g1277 ( 
.A(n_1114),
.Y(n_1277)
);

AOI21xp5_ASAP7_75t_L g1278 ( 
.A1(n_1158),
.A2(n_1186),
.B(n_1184),
.Y(n_1278)
);

NAND3xp33_ASAP7_75t_L g1279 ( 
.A(n_1110),
.B(n_871),
.C(n_868),
.Y(n_1279)
);

OAI21x1_ASAP7_75t_SL g1280 ( 
.A1(n_1151),
.A2(n_1009),
.B(n_997),
.Y(n_1280)
);

INVx2_ASAP7_75t_L g1281 ( 
.A(n_1137),
.Y(n_1281)
);

BUFx2_ASAP7_75t_SL g1282 ( 
.A(n_1176),
.Y(n_1282)
);

AO31x2_ASAP7_75t_L g1283 ( 
.A1(n_1168),
.A2(n_1065),
.A3(n_1093),
.B(n_1158),
.Y(n_1283)
);

OAI21x1_ASAP7_75t_L g1284 ( 
.A1(n_1119),
.A2(n_1100),
.B(n_1094),
.Y(n_1284)
);

OA21x2_ASAP7_75t_L g1285 ( 
.A1(n_1177),
.A2(n_1187),
.B(n_1184),
.Y(n_1285)
);

AND2x4_ASAP7_75t_L g1286 ( 
.A(n_1166),
.B(n_1172),
.Y(n_1286)
);

AOI221xp5_ASAP7_75t_L g1287 ( 
.A1(n_1118),
.A2(n_871),
.B1(n_868),
.B2(n_1115),
.C(n_695),
.Y(n_1287)
);

OAI21xp5_ASAP7_75t_L g1288 ( 
.A1(n_1110),
.A2(n_910),
.B(n_926),
.Y(n_1288)
);

BUFx3_ASAP7_75t_L g1289 ( 
.A(n_1082),
.Y(n_1289)
);

OAI21x1_ASAP7_75t_L g1290 ( 
.A1(n_1119),
.A2(n_1100),
.B(n_1094),
.Y(n_1290)
);

AND2x4_ASAP7_75t_L g1291 ( 
.A(n_1166),
.B(n_1172),
.Y(n_1291)
);

OAI21x1_ASAP7_75t_L g1292 ( 
.A1(n_1119),
.A2(n_1100),
.B(n_1094),
.Y(n_1292)
);

NAND2x1p5_ASAP7_75t_L g1293 ( 
.A(n_1150),
.B(n_999),
.Y(n_1293)
);

OAI21xp5_ASAP7_75t_L g1294 ( 
.A1(n_1110),
.A2(n_910),
.B(n_926),
.Y(n_1294)
);

CKINVDCx20_ASAP7_75t_R g1295 ( 
.A(n_1064),
.Y(n_1295)
);

AO31x2_ASAP7_75t_L g1296 ( 
.A1(n_1168),
.A2(n_1065),
.A3(n_1093),
.B(n_1158),
.Y(n_1296)
);

INVx1_ASAP7_75t_L g1297 ( 
.A(n_1059),
.Y(n_1297)
);

INVx1_ASAP7_75t_L g1298 ( 
.A(n_1059),
.Y(n_1298)
);

AND2x2_ASAP7_75t_L g1299 ( 
.A(n_1167),
.B(n_1096),
.Y(n_1299)
);

AOI21xp33_ASAP7_75t_L g1300 ( 
.A1(n_1108),
.A2(n_871),
.B(n_868),
.Y(n_1300)
);

BUFx3_ASAP7_75t_L g1301 ( 
.A(n_1082),
.Y(n_1301)
);

BUFx6f_ASAP7_75t_L g1302 ( 
.A(n_1114),
.Y(n_1302)
);

OAI21x1_ASAP7_75t_L g1303 ( 
.A1(n_1119),
.A2(n_1100),
.B(n_1094),
.Y(n_1303)
);

NAND2x1p5_ASAP7_75t_L g1304 ( 
.A(n_1150),
.B(n_999),
.Y(n_1304)
);

OAI22xp5_ASAP7_75t_L g1305 ( 
.A1(n_1162),
.A2(n_868),
.B1(n_871),
.B2(n_995),
.Y(n_1305)
);

AO32x2_ASAP7_75t_L g1306 ( 
.A1(n_1112),
.A2(n_1015),
.A3(n_1058),
.B1(n_1044),
.B2(n_943),
.Y(n_1306)
);

INVx1_ASAP7_75t_L g1307 ( 
.A(n_1059),
.Y(n_1307)
);

OA21x2_ASAP7_75t_L g1308 ( 
.A1(n_1210),
.A2(n_1260),
.B(n_1190),
.Y(n_1308)
);

AOI21xp5_ASAP7_75t_L g1309 ( 
.A1(n_1258),
.A2(n_1278),
.B(n_1262),
.Y(n_1309)
);

HB1xp67_ASAP7_75t_L g1310 ( 
.A(n_1196),
.Y(n_1310)
);

AOI21xp5_ASAP7_75t_SL g1311 ( 
.A1(n_1263),
.A2(n_1279),
.B(n_1276),
.Y(n_1311)
);

O2A1O1Ixp33_ASAP7_75t_L g1312 ( 
.A1(n_1300),
.A2(n_1268),
.B(n_1287),
.C(n_1288),
.Y(n_1312)
);

A2O1A1Ixp33_ASAP7_75t_L g1313 ( 
.A1(n_1287),
.A2(n_1300),
.B(n_1191),
.C(n_1204),
.Y(n_1313)
);

AOI221xp5_ASAP7_75t_L g1314 ( 
.A1(n_1191),
.A2(n_1259),
.B1(n_1268),
.B2(n_1204),
.C(n_1198),
.Y(n_1314)
);

AOI21xp5_ASAP7_75t_SL g1315 ( 
.A1(n_1257),
.A2(n_1294),
.B(n_1305),
.Y(n_1315)
);

OAI22xp5_ASAP7_75t_L g1316 ( 
.A1(n_1259),
.A2(n_1273),
.B1(n_1194),
.B2(n_1195),
.Y(n_1316)
);

INVxp67_ASAP7_75t_L g1317 ( 
.A(n_1274),
.Y(n_1317)
);

OAI22xp5_ASAP7_75t_L g1318 ( 
.A1(n_1194),
.A2(n_1273),
.B1(n_1195),
.B2(n_1197),
.Y(n_1318)
);

NAND2xp5_ASAP7_75t_L g1319 ( 
.A(n_1198),
.B(n_1197),
.Y(n_1319)
);

NOR2xp67_ASAP7_75t_L g1320 ( 
.A(n_1220),
.B(n_1223),
.Y(n_1320)
);

INVx2_ASAP7_75t_SL g1321 ( 
.A(n_1215),
.Y(n_1321)
);

AND2x2_ASAP7_75t_L g1322 ( 
.A(n_1200),
.B(n_1299),
.Y(n_1322)
);

AOI21xp5_ASAP7_75t_L g1323 ( 
.A1(n_1258),
.A2(n_1278),
.B(n_1262),
.Y(n_1323)
);

NAND2xp5_ASAP7_75t_L g1324 ( 
.A(n_1213),
.B(n_1214),
.Y(n_1324)
);

OAI22xp5_ASAP7_75t_L g1325 ( 
.A1(n_1254),
.A2(n_1219),
.B1(n_1230),
.B2(n_1206),
.Y(n_1325)
);

A2O1A1Ixp33_ASAP7_75t_L g1326 ( 
.A1(n_1248),
.A2(n_1206),
.B(n_1222),
.C(n_1236),
.Y(n_1326)
);

BUFx3_ASAP7_75t_L g1327 ( 
.A(n_1215),
.Y(n_1327)
);

CKINVDCx20_ASAP7_75t_R g1328 ( 
.A(n_1295),
.Y(n_1328)
);

A2O1A1Ixp33_ASAP7_75t_L g1329 ( 
.A1(n_1248),
.A2(n_1222),
.B(n_1236),
.C(n_1203),
.Y(n_1329)
);

AOI21xp5_ASAP7_75t_SL g1330 ( 
.A1(n_1221),
.A2(n_1293),
.B(n_1304),
.Y(n_1330)
);

CKINVDCx20_ASAP7_75t_R g1331 ( 
.A(n_1295),
.Y(n_1331)
);

OAI22xp5_ASAP7_75t_L g1332 ( 
.A1(n_1219),
.A2(n_1251),
.B1(n_1214),
.B2(n_1229),
.Y(n_1332)
);

OAI22xp5_ASAP7_75t_L g1333 ( 
.A1(n_1251),
.A2(n_1227),
.B1(n_1203),
.B2(n_1297),
.Y(n_1333)
);

CKINVDCx5p33_ASAP7_75t_R g1334 ( 
.A(n_1216),
.Y(n_1334)
);

OAI22xp5_ASAP7_75t_L g1335 ( 
.A1(n_1211),
.A2(n_1226),
.B1(n_1298),
.B2(n_1235),
.Y(n_1335)
);

O2A1O1Ixp5_ASAP7_75t_L g1336 ( 
.A1(n_1239),
.A2(n_1223),
.B(n_1224),
.C(n_1250),
.Y(n_1336)
);

NOR2xp67_ASAP7_75t_L g1337 ( 
.A(n_1189),
.B(n_1240),
.Y(n_1337)
);

BUFx6f_ASAP7_75t_L g1338 ( 
.A(n_1289),
.Y(n_1338)
);

OAI22xp5_ASAP7_75t_L g1339 ( 
.A1(n_1261),
.A2(n_1266),
.B1(n_1307),
.B2(n_1269),
.Y(n_1339)
);

CKINVDCx5p33_ASAP7_75t_R g1340 ( 
.A(n_1216),
.Y(n_1340)
);

OA22x2_ASAP7_75t_L g1341 ( 
.A1(n_1275),
.A2(n_1280),
.B1(n_1272),
.B2(n_1202),
.Y(n_1341)
);

AOI221x1_ASAP7_75t_SL g1342 ( 
.A1(n_1255),
.A2(n_1291),
.B1(n_1286),
.B2(n_1265),
.C(n_1306),
.Y(n_1342)
);

AOI21xp5_ASAP7_75t_SL g1343 ( 
.A1(n_1293),
.A2(n_1304),
.B(n_1192),
.Y(n_1343)
);

NAND2xp5_ASAP7_75t_L g1344 ( 
.A(n_1255),
.B(n_1291),
.Y(n_1344)
);

AND2x2_ASAP7_75t_L g1345 ( 
.A(n_1265),
.B(n_1286),
.Y(n_1345)
);

AOI221x1_ASAP7_75t_SL g1346 ( 
.A1(n_1306),
.A2(n_1242),
.B1(n_1224),
.B2(n_1188),
.C(n_1218),
.Y(n_1346)
);

INVx1_ASAP7_75t_SL g1347 ( 
.A(n_1232),
.Y(n_1347)
);

NAND2xp5_ASAP7_75t_L g1348 ( 
.A(n_1244),
.B(n_1228),
.Y(n_1348)
);

AND2x4_ASAP7_75t_L g1349 ( 
.A(n_1242),
.B(n_1243),
.Y(n_1349)
);

A2O1A1Ixp33_ASAP7_75t_L g1350 ( 
.A1(n_1217),
.A2(n_1212),
.B(n_1306),
.C(n_1246),
.Y(n_1350)
);

CKINVDCx16_ASAP7_75t_R g1351 ( 
.A(n_1289),
.Y(n_1351)
);

AND2x2_ASAP7_75t_L g1352 ( 
.A(n_1238),
.B(n_1243),
.Y(n_1352)
);

INVx1_ASAP7_75t_L g1353 ( 
.A(n_1237),
.Y(n_1353)
);

CKINVDCx5p33_ASAP7_75t_R g1354 ( 
.A(n_1188),
.Y(n_1354)
);

AOI21xp5_ASAP7_75t_L g1355 ( 
.A1(n_1192),
.A2(n_1285),
.B(n_1201),
.Y(n_1355)
);

OAI22xp5_ASAP7_75t_L g1356 ( 
.A1(n_1205),
.A2(n_1285),
.B1(n_1282),
.B2(n_1306),
.Y(n_1356)
);

AOI21xp5_ASAP7_75t_SL g1357 ( 
.A1(n_1301),
.A2(n_1234),
.B(n_1201),
.Y(n_1357)
);

O2A1O1Ixp33_ASAP7_75t_L g1358 ( 
.A1(n_1247),
.A2(n_1301),
.B(n_1267),
.C(n_1281),
.Y(n_1358)
);

CKINVDCx5p33_ASAP7_75t_R g1359 ( 
.A(n_1209),
.Y(n_1359)
);

OA21x2_ASAP7_75t_L g1360 ( 
.A1(n_1303),
.A2(n_1290),
.B(n_1271),
.Y(n_1360)
);

NAND2xp5_ASAP7_75t_L g1361 ( 
.A(n_1270),
.B(n_1205),
.Y(n_1361)
);

A2O1A1Ixp33_ASAP7_75t_L g1362 ( 
.A1(n_1231),
.A2(n_1233),
.B(n_1253),
.C(n_1208),
.Y(n_1362)
);

O2A1O1Ixp33_ASAP7_75t_L g1363 ( 
.A1(n_1207),
.A2(n_1256),
.B(n_1205),
.C(n_1252),
.Y(n_1363)
);

OAI22xp5_ASAP7_75t_L g1364 ( 
.A1(n_1252),
.A2(n_1302),
.B1(n_1277),
.B2(n_1209),
.Y(n_1364)
);

OA21x2_ASAP7_75t_L g1365 ( 
.A1(n_1264),
.A2(n_1284),
.B(n_1292),
.Y(n_1365)
);

A2O1A1Ixp33_ASAP7_75t_L g1366 ( 
.A1(n_1199),
.A2(n_1193),
.B(n_1218),
.C(n_1225),
.Y(n_1366)
);

AOI21x1_ASAP7_75t_SL g1367 ( 
.A1(n_1218),
.A2(n_1249),
.B(n_1296),
.Y(n_1367)
);

NAND2xp5_ASAP7_75t_L g1368 ( 
.A(n_1283),
.B(n_1296),
.Y(n_1368)
);

INVx1_ASAP7_75t_L g1369 ( 
.A(n_1241),
.Y(n_1369)
);

OAI22xp5_ASAP7_75t_L g1370 ( 
.A1(n_1225),
.A2(n_1277),
.B1(n_1302),
.B2(n_1283),
.Y(n_1370)
);

AOI221xp5_ASAP7_75t_L g1371 ( 
.A1(n_1245),
.A2(n_1118),
.B1(n_1287),
.B2(n_1191),
.C(n_1259),
.Y(n_1371)
);

AND2x2_ASAP7_75t_L g1372 ( 
.A(n_1302),
.B(n_1283),
.Y(n_1372)
);

NOR2x1_ASAP7_75t_SL g1373 ( 
.A(n_1283),
.B(n_1296),
.Y(n_1373)
);

CKINVDCx20_ASAP7_75t_R g1374 ( 
.A(n_1296),
.Y(n_1374)
);

O2A1O1Ixp33_ASAP7_75t_L g1375 ( 
.A1(n_1300),
.A2(n_1110),
.B(n_1268),
.C(n_1118),
.Y(n_1375)
);

BUFx2_ASAP7_75t_L g1376 ( 
.A(n_1196),
.Y(n_1376)
);

NAND2xp5_ASAP7_75t_L g1377 ( 
.A(n_1194),
.B(n_1273),
.Y(n_1377)
);

OR2x2_ASAP7_75t_L g1378 ( 
.A(n_1213),
.B(n_1299),
.Y(n_1378)
);

HB1xp67_ASAP7_75t_L g1379 ( 
.A(n_1196),
.Y(n_1379)
);

O2A1O1Ixp33_ASAP7_75t_L g1380 ( 
.A1(n_1300),
.A2(n_1110),
.B(n_1268),
.C(n_1118),
.Y(n_1380)
);

BUFx3_ASAP7_75t_L g1381 ( 
.A(n_1215),
.Y(n_1381)
);

AND2x2_ASAP7_75t_L g1382 ( 
.A(n_1200),
.B(n_1096),
.Y(n_1382)
);

A2O1A1Ixp33_ASAP7_75t_L g1383 ( 
.A1(n_1287),
.A2(n_1300),
.B(n_871),
.C(n_868),
.Y(n_1383)
);

INVx6_ASAP7_75t_L g1384 ( 
.A(n_1215),
.Y(n_1384)
);

OAI22xp5_ASAP7_75t_L g1385 ( 
.A1(n_1259),
.A2(n_871),
.B1(n_868),
.B2(n_1162),
.Y(n_1385)
);

O2A1O1Ixp33_ASAP7_75t_L g1386 ( 
.A1(n_1300),
.A2(n_1110),
.B(n_1268),
.C(n_1118),
.Y(n_1386)
);

OA21x2_ASAP7_75t_L g1387 ( 
.A1(n_1210),
.A2(n_1065),
.B(n_1093),
.Y(n_1387)
);

NAND2xp5_ASAP7_75t_L g1388 ( 
.A(n_1194),
.B(n_1273),
.Y(n_1388)
);

AND2x2_ASAP7_75t_L g1389 ( 
.A(n_1200),
.B(n_1096),
.Y(n_1389)
);

NAND2xp5_ASAP7_75t_L g1390 ( 
.A(n_1194),
.B(n_1273),
.Y(n_1390)
);

AOI21xp5_ASAP7_75t_L g1391 ( 
.A1(n_1258),
.A2(n_1108),
.B(n_1262),
.Y(n_1391)
);

HB1xp67_ASAP7_75t_L g1392 ( 
.A(n_1196),
.Y(n_1392)
);

O2A1O1Ixp5_ASAP7_75t_L g1393 ( 
.A1(n_1268),
.A2(n_1168),
.B(n_1108),
.C(n_995),
.Y(n_1393)
);

INVx2_ASAP7_75t_L g1394 ( 
.A(n_1353),
.Y(n_1394)
);

INVx4_ASAP7_75t_SL g1395 ( 
.A(n_1372),
.Y(n_1395)
);

OAI21xp5_ASAP7_75t_SL g1396 ( 
.A1(n_1314),
.A2(n_1313),
.B(n_1312),
.Y(n_1396)
);

OR2x2_ASAP7_75t_L g1397 ( 
.A(n_1368),
.B(n_1361),
.Y(n_1397)
);

HB1xp67_ASAP7_75t_L g1398 ( 
.A(n_1369),
.Y(n_1398)
);

AND2x2_ASAP7_75t_L g1399 ( 
.A(n_1373),
.B(n_1350),
.Y(n_1399)
);

INVx2_ASAP7_75t_L g1400 ( 
.A(n_1360),
.Y(n_1400)
);

AND2x2_ASAP7_75t_L g1401 ( 
.A(n_1356),
.B(n_1374),
.Y(n_1401)
);

INVx2_ASAP7_75t_SL g1402 ( 
.A(n_1352),
.Y(n_1402)
);

AND2x4_ASAP7_75t_L g1403 ( 
.A(n_1366),
.B(n_1362),
.Y(n_1403)
);

NAND3xp33_ASAP7_75t_L g1404 ( 
.A(n_1375),
.B(n_1380),
.C(n_1386),
.Y(n_1404)
);

OAI22xp5_ASAP7_75t_L g1405 ( 
.A1(n_1388),
.A2(n_1377),
.B1(n_1390),
.B2(n_1326),
.Y(n_1405)
);

HB1xp67_ASAP7_75t_L g1406 ( 
.A(n_1356),
.Y(n_1406)
);

OAI21x1_ASAP7_75t_L g1407 ( 
.A1(n_1309),
.A2(n_1323),
.B(n_1391),
.Y(n_1407)
);

OR2x2_ASAP7_75t_L g1408 ( 
.A(n_1355),
.B(n_1348),
.Y(n_1408)
);

NAND2xp5_ASAP7_75t_L g1409 ( 
.A(n_1318),
.B(n_1316),
.Y(n_1409)
);

INVx1_ASAP7_75t_L g1410 ( 
.A(n_1335),
.Y(n_1410)
);

INVxp67_ASAP7_75t_SL g1411 ( 
.A(n_1363),
.Y(n_1411)
);

AO21x2_ASAP7_75t_L g1412 ( 
.A1(n_1357),
.A2(n_1315),
.B(n_1329),
.Y(n_1412)
);

OA21x2_ASAP7_75t_L g1413 ( 
.A1(n_1393),
.A2(n_1371),
.B(n_1319),
.Y(n_1413)
);

INVx1_ASAP7_75t_L g1414 ( 
.A(n_1335),
.Y(n_1414)
);

INVx2_ASAP7_75t_L g1415 ( 
.A(n_1360),
.Y(n_1415)
);

OAI21x1_ASAP7_75t_L g1416 ( 
.A1(n_1367),
.A2(n_1365),
.B(n_1308),
.Y(n_1416)
);

AOI21x1_ASAP7_75t_L g1417 ( 
.A1(n_1365),
.A2(n_1308),
.B(n_1319),
.Y(n_1417)
);

INVx1_ASAP7_75t_L g1418 ( 
.A(n_1339),
.Y(n_1418)
);

INVx1_ASAP7_75t_L g1419 ( 
.A(n_1339),
.Y(n_1419)
);

HB1xp67_ASAP7_75t_L g1420 ( 
.A(n_1387),
.Y(n_1420)
);

AO21x2_ASAP7_75t_L g1421 ( 
.A1(n_1358),
.A2(n_1370),
.B(n_1332),
.Y(n_1421)
);

NAND3xp33_ASAP7_75t_L g1422 ( 
.A(n_1383),
.B(n_1385),
.C(n_1316),
.Y(n_1422)
);

AND2x2_ASAP7_75t_L g1423 ( 
.A(n_1382),
.B(n_1389),
.Y(n_1423)
);

AOI22xp33_ASAP7_75t_SL g1424 ( 
.A1(n_1333),
.A2(n_1332),
.B1(n_1318),
.B2(n_1325),
.Y(n_1424)
);

OA21x2_ASAP7_75t_L g1425 ( 
.A1(n_1336),
.A2(n_1370),
.B(n_1333),
.Y(n_1425)
);

AND2x2_ASAP7_75t_L g1426 ( 
.A(n_1341),
.B(n_1322),
.Y(n_1426)
);

INVxp67_ASAP7_75t_L g1427 ( 
.A(n_1310),
.Y(n_1427)
);

AO21x2_ASAP7_75t_L g1428 ( 
.A1(n_1343),
.A2(n_1330),
.B(n_1325),
.Y(n_1428)
);

INVx1_ASAP7_75t_L g1429 ( 
.A(n_1346),
.Y(n_1429)
);

INVx1_ASAP7_75t_L g1430 ( 
.A(n_1324),
.Y(n_1430)
);

OR2x2_ASAP7_75t_L g1431 ( 
.A(n_1378),
.B(n_1392),
.Y(n_1431)
);

INVx2_ASAP7_75t_SL g1432 ( 
.A(n_1379),
.Y(n_1432)
);

INVx1_ASAP7_75t_L g1433 ( 
.A(n_1342),
.Y(n_1433)
);

CKINVDCx5p33_ASAP7_75t_R g1434 ( 
.A(n_1334),
.Y(n_1434)
);

INVx1_ASAP7_75t_L g1435 ( 
.A(n_1364),
.Y(n_1435)
);

INVx2_ASAP7_75t_L g1436 ( 
.A(n_1376),
.Y(n_1436)
);

INVx3_ASAP7_75t_L g1437 ( 
.A(n_1349),
.Y(n_1437)
);

AND2x2_ASAP7_75t_L g1438 ( 
.A(n_1377),
.B(n_1390),
.Y(n_1438)
);

INVx1_ASAP7_75t_L g1439 ( 
.A(n_1317),
.Y(n_1439)
);

INVx2_ASAP7_75t_L g1440 ( 
.A(n_1359),
.Y(n_1440)
);

INVx1_ASAP7_75t_L g1441 ( 
.A(n_1320),
.Y(n_1441)
);

INVx1_ASAP7_75t_L g1442 ( 
.A(n_1311),
.Y(n_1442)
);

INVx1_ASAP7_75t_SL g1443 ( 
.A(n_1347),
.Y(n_1443)
);

OAI21xp5_ASAP7_75t_SL g1444 ( 
.A1(n_1396),
.A2(n_1385),
.B(n_1345),
.Y(n_1444)
);

AOI22xp33_ASAP7_75t_L g1445 ( 
.A1(n_1422),
.A2(n_1337),
.B1(n_1384),
.B2(n_1327),
.Y(n_1445)
);

BUFx2_ASAP7_75t_L g1446 ( 
.A(n_1395),
.Y(n_1446)
);

OA21x2_ASAP7_75t_L g1447 ( 
.A1(n_1416),
.A2(n_1344),
.B(n_1321),
.Y(n_1447)
);

AND2x2_ASAP7_75t_L g1448 ( 
.A(n_1401),
.B(n_1351),
.Y(n_1448)
);

INVx2_ASAP7_75t_L g1449 ( 
.A(n_1394),
.Y(n_1449)
);

HB1xp67_ASAP7_75t_L g1450 ( 
.A(n_1398),
.Y(n_1450)
);

NOR2x1_ASAP7_75t_R g1451 ( 
.A(n_1434),
.B(n_1340),
.Y(n_1451)
);

AND2x4_ASAP7_75t_L g1452 ( 
.A(n_1395),
.B(n_1402),
.Y(n_1452)
);

INVxp67_ASAP7_75t_L g1453 ( 
.A(n_1411),
.Y(n_1453)
);

INVxp67_ASAP7_75t_L g1454 ( 
.A(n_1411),
.Y(n_1454)
);

AOI22xp33_ASAP7_75t_L g1455 ( 
.A1(n_1422),
.A2(n_1384),
.B1(n_1381),
.B2(n_1338),
.Y(n_1455)
);

BUFx3_ASAP7_75t_L g1456 ( 
.A(n_1442),
.Y(n_1456)
);

INVx2_ASAP7_75t_L g1457 ( 
.A(n_1400),
.Y(n_1457)
);

OAI221xp5_ASAP7_75t_L g1458 ( 
.A1(n_1396),
.A2(n_1384),
.B1(n_1354),
.B2(n_1331),
.C(n_1328),
.Y(n_1458)
);

INVx2_ASAP7_75t_R g1459 ( 
.A(n_1435),
.Y(n_1459)
);

BUFx2_ASAP7_75t_L g1460 ( 
.A(n_1395),
.Y(n_1460)
);

HB1xp67_ASAP7_75t_L g1461 ( 
.A(n_1398),
.Y(n_1461)
);

INVx1_ASAP7_75t_SL g1462 ( 
.A(n_1443),
.Y(n_1462)
);

INVx2_ASAP7_75t_L g1463 ( 
.A(n_1400),
.Y(n_1463)
);

OR2x2_ASAP7_75t_L g1464 ( 
.A(n_1397),
.B(n_1408),
.Y(n_1464)
);

NOR4xp25_ASAP7_75t_SL g1465 ( 
.A(n_1424),
.B(n_1412),
.C(n_1441),
.D(n_1435),
.Y(n_1465)
);

OR2x2_ASAP7_75t_L g1466 ( 
.A(n_1397),
.B(n_1408),
.Y(n_1466)
);

BUFx3_ASAP7_75t_L g1467 ( 
.A(n_1441),
.Y(n_1467)
);

INVx2_ASAP7_75t_L g1468 ( 
.A(n_1400),
.Y(n_1468)
);

OAI221xp5_ASAP7_75t_L g1469 ( 
.A1(n_1424),
.A2(n_1404),
.B1(n_1409),
.B2(n_1413),
.C(n_1405),
.Y(n_1469)
);

BUFx2_ASAP7_75t_L g1470 ( 
.A(n_1446),
.Y(n_1470)
);

AND4x1_ASAP7_75t_L g1471 ( 
.A(n_1445),
.B(n_1404),
.C(n_1409),
.D(n_1433),
.Y(n_1471)
);

AND2x4_ASAP7_75t_L g1472 ( 
.A(n_1446),
.B(n_1428),
.Y(n_1472)
);

INVx1_ASAP7_75t_L g1473 ( 
.A(n_1449),
.Y(n_1473)
);

AOI22xp33_ASAP7_75t_SL g1474 ( 
.A1(n_1469),
.A2(n_1412),
.B1(n_1413),
.B2(n_1428),
.Y(n_1474)
);

INVx1_ASAP7_75t_SL g1475 ( 
.A(n_1462),
.Y(n_1475)
);

OAI332xp33_ASAP7_75t_L g1476 ( 
.A1(n_1469),
.A2(n_1405),
.A3(n_1433),
.B1(n_1429),
.B2(n_1443),
.B3(n_1439),
.C1(n_1418),
.C2(n_1414),
.Y(n_1476)
);

NOR2xp33_ASAP7_75t_R g1477 ( 
.A(n_1462),
.B(n_1437),
.Y(n_1477)
);

CKINVDCx16_ASAP7_75t_R g1478 ( 
.A(n_1448),
.Y(n_1478)
);

INVx5_ASAP7_75t_L g1479 ( 
.A(n_1460),
.Y(n_1479)
);

AOI21x1_ASAP7_75t_L g1480 ( 
.A1(n_1457),
.A2(n_1420),
.B(n_1417),
.Y(n_1480)
);

OAI211xp5_ASAP7_75t_L g1481 ( 
.A1(n_1465),
.A2(n_1425),
.B(n_1406),
.C(n_1413),
.Y(n_1481)
);

OAI221xp5_ASAP7_75t_L g1482 ( 
.A1(n_1444),
.A2(n_1425),
.B1(n_1413),
.B2(n_1408),
.C(n_1427),
.Y(n_1482)
);

INVx1_ASAP7_75t_L g1483 ( 
.A(n_1449),
.Y(n_1483)
);

INVx3_ASAP7_75t_L g1484 ( 
.A(n_1452),
.Y(n_1484)
);

INVx2_ASAP7_75t_L g1485 ( 
.A(n_1463),
.Y(n_1485)
);

NAND2xp5_ASAP7_75t_L g1486 ( 
.A(n_1464),
.B(n_1438),
.Y(n_1486)
);

NAND2xp5_ASAP7_75t_L g1487 ( 
.A(n_1466),
.B(n_1438),
.Y(n_1487)
);

OAI22xp5_ASAP7_75t_L g1488 ( 
.A1(n_1455),
.A2(n_1429),
.B1(n_1413),
.B2(n_1440),
.Y(n_1488)
);

AOI22xp33_ASAP7_75t_SL g1489 ( 
.A1(n_1458),
.A2(n_1412),
.B1(n_1413),
.B2(n_1428),
.Y(n_1489)
);

AOI221xp5_ASAP7_75t_L g1490 ( 
.A1(n_1453),
.A2(n_1427),
.B1(n_1406),
.B2(n_1439),
.C(n_1430),
.Y(n_1490)
);

AOI222xp33_ASAP7_75t_L g1491 ( 
.A1(n_1444),
.A2(n_1423),
.B1(n_1430),
.B2(n_1414),
.C1(n_1419),
.C2(n_1410),
.Y(n_1491)
);

INVxp67_ASAP7_75t_L g1492 ( 
.A(n_1467),
.Y(n_1492)
);

OAI211xp5_ASAP7_75t_SL g1493 ( 
.A1(n_1454),
.A2(n_1431),
.B(n_1436),
.C(n_1432),
.Y(n_1493)
);

HB1xp67_ASAP7_75t_L g1494 ( 
.A(n_1450),
.Y(n_1494)
);

NAND2xp5_ASAP7_75t_L g1495 ( 
.A(n_1466),
.B(n_1436),
.Y(n_1495)
);

AOI22xp33_ASAP7_75t_SL g1496 ( 
.A1(n_1458),
.A2(n_1412),
.B1(n_1428),
.B2(n_1421),
.Y(n_1496)
);

HB1xp67_ASAP7_75t_L g1497 ( 
.A(n_1450),
.Y(n_1497)
);

BUFx6f_ASAP7_75t_L g1498 ( 
.A(n_1456),
.Y(n_1498)
);

OAI221xp5_ASAP7_75t_L g1499 ( 
.A1(n_1454),
.A2(n_1425),
.B1(n_1436),
.B2(n_1432),
.C(n_1431),
.Y(n_1499)
);

OR2x2_ASAP7_75t_L g1500 ( 
.A(n_1494),
.B(n_1459),
.Y(n_1500)
);

NOR2xp33_ASAP7_75t_L g1501 ( 
.A(n_1471),
.B(n_1476),
.Y(n_1501)
);

AND2x2_ASAP7_75t_L g1502 ( 
.A(n_1484),
.B(n_1459),
.Y(n_1502)
);

INVx2_ASAP7_75t_SL g1503 ( 
.A(n_1479),
.Y(n_1503)
);

INVxp67_ASAP7_75t_SL g1504 ( 
.A(n_1497),
.Y(n_1504)
);

INVx1_ASAP7_75t_L g1505 ( 
.A(n_1473),
.Y(n_1505)
);

INVx1_ASAP7_75t_L g1506 ( 
.A(n_1473),
.Y(n_1506)
);

AND2x4_ASAP7_75t_L g1507 ( 
.A(n_1484),
.B(n_1460),
.Y(n_1507)
);

INVx2_ASAP7_75t_L g1508 ( 
.A(n_1480),
.Y(n_1508)
);

INVx2_ASAP7_75t_SL g1509 ( 
.A(n_1479),
.Y(n_1509)
);

INVx1_ASAP7_75t_L g1510 ( 
.A(n_1483),
.Y(n_1510)
);

BUFx3_ASAP7_75t_L g1511 ( 
.A(n_1498),
.Y(n_1511)
);

BUFx2_ASAP7_75t_L g1512 ( 
.A(n_1479),
.Y(n_1512)
);

INVx1_ASAP7_75t_SL g1513 ( 
.A(n_1470),
.Y(n_1513)
);

AND2x4_ASAP7_75t_L g1514 ( 
.A(n_1484),
.B(n_1452),
.Y(n_1514)
);

NAND2xp5_ASAP7_75t_L g1515 ( 
.A(n_1490),
.B(n_1461),
.Y(n_1515)
);

INVx3_ASAP7_75t_L g1516 ( 
.A(n_1479),
.Y(n_1516)
);

AO21x1_ASAP7_75t_L g1517 ( 
.A1(n_1488),
.A2(n_1403),
.B(n_1465),
.Y(n_1517)
);

OA21x2_ASAP7_75t_L g1518 ( 
.A1(n_1481),
.A2(n_1415),
.B(n_1468),
.Y(n_1518)
);

OA21x2_ASAP7_75t_L g1519 ( 
.A1(n_1499),
.A2(n_1399),
.B(n_1407),
.Y(n_1519)
);

NAND3xp33_ASAP7_75t_SL g1520 ( 
.A(n_1471),
.B(n_1448),
.C(n_1440),
.Y(n_1520)
);

OR2x2_ASAP7_75t_L g1521 ( 
.A(n_1485),
.B(n_1447),
.Y(n_1521)
);

AND2x2_ASAP7_75t_L g1522 ( 
.A(n_1514),
.B(n_1478),
.Y(n_1522)
);

INVx3_ASAP7_75t_L g1523 ( 
.A(n_1516),
.Y(n_1523)
);

AND2x2_ASAP7_75t_SL g1524 ( 
.A(n_1501),
.B(n_1478),
.Y(n_1524)
);

INVx1_ASAP7_75t_L g1525 ( 
.A(n_1505),
.Y(n_1525)
);

INVx1_ASAP7_75t_SL g1526 ( 
.A(n_1513),
.Y(n_1526)
);

INVx2_ASAP7_75t_L g1527 ( 
.A(n_1521),
.Y(n_1527)
);

OR2x2_ASAP7_75t_L g1528 ( 
.A(n_1515),
.B(n_1486),
.Y(n_1528)
);

AND2x2_ASAP7_75t_L g1529 ( 
.A(n_1514),
.B(n_1507),
.Y(n_1529)
);

NAND2xp5_ASAP7_75t_L g1530 ( 
.A(n_1501),
.B(n_1491),
.Y(n_1530)
);

NAND3xp33_ASAP7_75t_L g1531 ( 
.A(n_1518),
.B(n_1474),
.C(n_1496),
.Y(n_1531)
);

INVx1_ASAP7_75t_L g1532 ( 
.A(n_1505),
.Y(n_1532)
);

OR2x2_ASAP7_75t_L g1533 ( 
.A(n_1504),
.B(n_1487),
.Y(n_1533)
);

OAI31xp33_ASAP7_75t_L g1534 ( 
.A1(n_1520),
.A2(n_1482),
.A3(n_1493),
.B(n_1476),
.Y(n_1534)
);

AOI22xp33_ASAP7_75t_L g1535 ( 
.A1(n_1520),
.A2(n_1489),
.B1(n_1421),
.B2(n_1425),
.Y(n_1535)
);

OR2x2_ASAP7_75t_L g1536 ( 
.A(n_1504),
.B(n_1495),
.Y(n_1536)
);

AND2x2_ASAP7_75t_L g1537 ( 
.A(n_1507),
.B(n_1470),
.Y(n_1537)
);

NAND2xp5_ASAP7_75t_L g1538 ( 
.A(n_1513),
.B(n_1475),
.Y(n_1538)
);

NAND2xp5_ASAP7_75t_L g1539 ( 
.A(n_1511),
.B(n_1432),
.Y(n_1539)
);

OR2x2_ASAP7_75t_L g1540 ( 
.A(n_1518),
.B(n_1510),
.Y(n_1540)
);

OR2x2_ASAP7_75t_L g1541 ( 
.A(n_1518),
.B(n_1472),
.Y(n_1541)
);

HB1xp67_ASAP7_75t_L g1542 ( 
.A(n_1518),
.Y(n_1542)
);

INVx5_ASAP7_75t_L g1543 ( 
.A(n_1516),
.Y(n_1543)
);

AND2x2_ASAP7_75t_L g1544 ( 
.A(n_1507),
.B(n_1511),
.Y(n_1544)
);

AND2x2_ASAP7_75t_L g1545 ( 
.A(n_1507),
.B(n_1511),
.Y(n_1545)
);

INVx1_ASAP7_75t_L g1546 ( 
.A(n_1505),
.Y(n_1546)
);

NAND2xp33_ASAP7_75t_R g1547 ( 
.A(n_1512),
.B(n_1477),
.Y(n_1547)
);

OR2x2_ASAP7_75t_L g1548 ( 
.A(n_1518),
.B(n_1472),
.Y(n_1548)
);

AND2x2_ASAP7_75t_L g1549 ( 
.A(n_1511),
.B(n_1479),
.Y(n_1549)
);

NOR2xp33_ASAP7_75t_L g1550 ( 
.A(n_1517),
.B(n_1451),
.Y(n_1550)
);

INVx1_ASAP7_75t_L g1551 ( 
.A(n_1506),
.Y(n_1551)
);

NOR2xp33_ASAP7_75t_L g1552 ( 
.A(n_1517),
.B(n_1451),
.Y(n_1552)
);

OAI211xp5_ASAP7_75t_L g1553 ( 
.A1(n_1519),
.A2(n_1425),
.B(n_1492),
.C(n_1479),
.Y(n_1553)
);

INVx2_ASAP7_75t_L g1554 ( 
.A(n_1521),
.Y(n_1554)
);

AOI22xp33_ASAP7_75t_L g1555 ( 
.A1(n_1517),
.A2(n_1421),
.B1(n_1519),
.B2(n_1403),
.Y(n_1555)
);

INVxp67_ASAP7_75t_SL g1556 ( 
.A(n_1547),
.Y(n_1556)
);

INVx2_ASAP7_75t_L g1557 ( 
.A(n_1540),
.Y(n_1557)
);

INVx3_ASAP7_75t_SL g1558 ( 
.A(n_1524),
.Y(n_1558)
);

INVx1_ASAP7_75t_L g1559 ( 
.A(n_1525),
.Y(n_1559)
);

AND2x2_ASAP7_75t_L g1560 ( 
.A(n_1522),
.B(n_1512),
.Y(n_1560)
);

A2O1A1Ixp33_ASAP7_75t_L g1561 ( 
.A1(n_1550),
.A2(n_1512),
.B(n_1509),
.C(n_1503),
.Y(n_1561)
);

INVx1_ASAP7_75t_L g1562 ( 
.A(n_1525),
.Y(n_1562)
);

INVx1_ASAP7_75t_L g1563 ( 
.A(n_1532),
.Y(n_1563)
);

INVx1_ASAP7_75t_L g1564 ( 
.A(n_1532),
.Y(n_1564)
);

NOR2xp33_ASAP7_75t_L g1565 ( 
.A(n_1530),
.B(n_1423),
.Y(n_1565)
);

AND2x2_ASAP7_75t_L g1566 ( 
.A(n_1522),
.B(n_1503),
.Y(n_1566)
);

AND2x2_ASAP7_75t_L g1567 ( 
.A(n_1544),
.B(n_1509),
.Y(n_1567)
);

AND2x2_ASAP7_75t_L g1568 ( 
.A(n_1544),
.B(n_1509),
.Y(n_1568)
);

NAND2xp33_ASAP7_75t_L g1569 ( 
.A(n_1535),
.B(n_1498),
.Y(n_1569)
);

NOR2xp33_ASAP7_75t_L g1570 ( 
.A(n_1524),
.B(n_1552),
.Y(n_1570)
);

AOI22xp5_ASAP7_75t_L g1571 ( 
.A1(n_1524),
.A2(n_1421),
.B1(n_1519),
.B2(n_1518),
.Y(n_1571)
);

INVx1_ASAP7_75t_L g1572 ( 
.A(n_1546),
.Y(n_1572)
);

INVx1_ASAP7_75t_L g1573 ( 
.A(n_1546),
.Y(n_1573)
);

INVx1_ASAP7_75t_L g1574 ( 
.A(n_1551),
.Y(n_1574)
);

NAND2xp5_ASAP7_75t_L g1575 ( 
.A(n_1534),
.B(n_1467),
.Y(n_1575)
);

INVx2_ASAP7_75t_L g1576 ( 
.A(n_1540),
.Y(n_1576)
);

HB1xp67_ASAP7_75t_L g1577 ( 
.A(n_1526),
.Y(n_1577)
);

NAND2xp5_ASAP7_75t_L g1578 ( 
.A(n_1534),
.B(n_1423),
.Y(n_1578)
);

OR2x2_ASAP7_75t_L g1579 ( 
.A(n_1526),
.B(n_1500),
.Y(n_1579)
);

INVx1_ASAP7_75t_L g1580 ( 
.A(n_1551),
.Y(n_1580)
);

NOR2x1_ASAP7_75t_L g1581 ( 
.A(n_1531),
.B(n_1516),
.Y(n_1581)
);

NAND2x1_ASAP7_75t_L g1582 ( 
.A(n_1549),
.B(n_1516),
.Y(n_1582)
);

AND2x2_ASAP7_75t_L g1583 ( 
.A(n_1545),
.B(n_1516),
.Y(n_1583)
);

AND2x2_ASAP7_75t_L g1584 ( 
.A(n_1545),
.B(n_1502),
.Y(n_1584)
);

OR2x2_ASAP7_75t_L g1585 ( 
.A(n_1528),
.B(n_1533),
.Y(n_1585)
);

NAND2xp5_ASAP7_75t_L g1586 ( 
.A(n_1538),
.B(n_1426),
.Y(n_1586)
);

OR2x2_ASAP7_75t_L g1587 ( 
.A(n_1533),
.B(n_1519),
.Y(n_1587)
);

INVx1_ASAP7_75t_SL g1588 ( 
.A(n_1558),
.Y(n_1588)
);

INVx2_ASAP7_75t_SL g1589 ( 
.A(n_1582),
.Y(n_1589)
);

INVx1_ASAP7_75t_L g1590 ( 
.A(n_1577),
.Y(n_1590)
);

INVx2_ASAP7_75t_L g1591 ( 
.A(n_1557),
.Y(n_1591)
);

INVx2_ASAP7_75t_L g1592 ( 
.A(n_1557),
.Y(n_1592)
);

AO21x1_ASAP7_75t_L g1593 ( 
.A1(n_1570),
.A2(n_1542),
.B(n_1541),
.Y(n_1593)
);

NOR2x1_ASAP7_75t_L g1594 ( 
.A(n_1581),
.B(n_1531),
.Y(n_1594)
);

NAND2xp5_ASAP7_75t_L g1595 ( 
.A(n_1565),
.B(n_1536),
.Y(n_1595)
);

HB1xp67_ASAP7_75t_L g1596 ( 
.A(n_1579),
.Y(n_1596)
);

INVx1_ASAP7_75t_SL g1597 ( 
.A(n_1558),
.Y(n_1597)
);

AND2x2_ASAP7_75t_L g1598 ( 
.A(n_1556),
.B(n_1529),
.Y(n_1598)
);

OAI22xp5_ASAP7_75t_L g1599 ( 
.A1(n_1575),
.A2(n_1555),
.B1(n_1553),
.B2(n_1538),
.Y(n_1599)
);

OR2x2_ASAP7_75t_L g1600 ( 
.A(n_1585),
.B(n_1536),
.Y(n_1600)
);

INVx1_ASAP7_75t_L g1601 ( 
.A(n_1559),
.Y(n_1601)
);

HB1xp67_ASAP7_75t_L g1602 ( 
.A(n_1579),
.Y(n_1602)
);

INVx1_ASAP7_75t_SL g1603 ( 
.A(n_1560),
.Y(n_1603)
);

AND2x2_ASAP7_75t_L g1604 ( 
.A(n_1560),
.B(n_1549),
.Y(n_1604)
);

INVx2_ASAP7_75t_L g1605 ( 
.A(n_1576),
.Y(n_1605)
);

INVx2_ASAP7_75t_L g1606 ( 
.A(n_1576),
.Y(n_1606)
);

INVx2_ASAP7_75t_L g1607 ( 
.A(n_1584),
.Y(n_1607)
);

AND2x2_ASAP7_75t_L g1608 ( 
.A(n_1566),
.B(n_1537),
.Y(n_1608)
);

INVx1_ASAP7_75t_L g1609 ( 
.A(n_1562),
.Y(n_1609)
);

AND2x2_ASAP7_75t_L g1610 ( 
.A(n_1566),
.B(n_1567),
.Y(n_1610)
);

INVx3_ASAP7_75t_L g1611 ( 
.A(n_1584),
.Y(n_1611)
);

INVxp33_ASAP7_75t_L g1612 ( 
.A(n_1570),
.Y(n_1612)
);

INVx1_ASAP7_75t_L g1613 ( 
.A(n_1596),
.Y(n_1613)
);

AND2x2_ASAP7_75t_L g1614 ( 
.A(n_1610),
.B(n_1567),
.Y(n_1614)
);

OAI21xp5_ASAP7_75t_L g1615 ( 
.A1(n_1594),
.A2(n_1561),
.B(n_1569),
.Y(n_1615)
);

NOR2xp67_ASAP7_75t_SL g1616 ( 
.A(n_1590),
.B(n_1543),
.Y(n_1616)
);

AND2x2_ASAP7_75t_L g1617 ( 
.A(n_1610),
.B(n_1568),
.Y(n_1617)
);

OR2x2_ASAP7_75t_L g1618 ( 
.A(n_1603),
.B(n_1578),
.Y(n_1618)
);

INVx1_ASAP7_75t_L g1619 ( 
.A(n_1596),
.Y(n_1619)
);

INVx1_ASAP7_75t_L g1620 ( 
.A(n_1602),
.Y(n_1620)
);

NAND2xp5_ASAP7_75t_L g1621 ( 
.A(n_1588),
.B(n_1565),
.Y(n_1621)
);

HB1xp67_ASAP7_75t_L g1622 ( 
.A(n_1602),
.Y(n_1622)
);

NAND2xp5_ASAP7_75t_L g1623 ( 
.A(n_1590),
.B(n_1563),
.Y(n_1623)
);

INVx2_ASAP7_75t_L g1624 ( 
.A(n_1611),
.Y(n_1624)
);

INVx1_ASAP7_75t_SL g1625 ( 
.A(n_1588),
.Y(n_1625)
);

INVx2_ASAP7_75t_L g1626 ( 
.A(n_1611),
.Y(n_1626)
);

NAND3xp33_ASAP7_75t_L g1627 ( 
.A(n_1594),
.B(n_1569),
.C(n_1571),
.Y(n_1627)
);

OAI22xp5_ASAP7_75t_L g1628 ( 
.A1(n_1597),
.A2(n_1561),
.B1(n_1587),
.B2(n_1548),
.Y(n_1628)
);

AO32x1_ASAP7_75t_L g1629 ( 
.A1(n_1599),
.A2(n_1568),
.A3(n_1583),
.B1(n_1573),
.B2(n_1572),
.Y(n_1629)
);

OAI32xp33_ASAP7_75t_L g1630 ( 
.A1(n_1599),
.A2(n_1541),
.A3(n_1548),
.B1(n_1583),
.B2(n_1523),
.Y(n_1630)
);

AOI22xp5_ASAP7_75t_L g1631 ( 
.A1(n_1597),
.A2(n_1598),
.B1(n_1604),
.B2(n_1612),
.Y(n_1631)
);

NAND2xp5_ASAP7_75t_L g1632 ( 
.A(n_1622),
.B(n_1603),
.Y(n_1632)
);

OR2x2_ASAP7_75t_L g1633 ( 
.A(n_1625),
.B(n_1595),
.Y(n_1633)
);

NAND2xp5_ASAP7_75t_L g1634 ( 
.A(n_1625),
.B(n_1598),
.Y(n_1634)
);

INVx1_ASAP7_75t_L g1635 ( 
.A(n_1613),
.Y(n_1635)
);

INVx1_ASAP7_75t_L g1636 ( 
.A(n_1619),
.Y(n_1636)
);

CKINVDCx20_ASAP7_75t_R g1637 ( 
.A(n_1621),
.Y(n_1637)
);

AND2x2_ASAP7_75t_L g1638 ( 
.A(n_1614),
.B(n_1598),
.Y(n_1638)
);

NAND2xp5_ASAP7_75t_L g1639 ( 
.A(n_1631),
.B(n_1604),
.Y(n_1639)
);

NAND2x1_ASAP7_75t_L g1640 ( 
.A(n_1615),
.B(n_1589),
.Y(n_1640)
);

NOR2xp33_ASAP7_75t_L g1641 ( 
.A(n_1620),
.B(n_1595),
.Y(n_1641)
);

AND2x2_ASAP7_75t_L g1642 ( 
.A(n_1617),
.B(n_1608),
.Y(n_1642)
);

AOI22xp5_ASAP7_75t_L g1643 ( 
.A1(n_1627),
.A2(n_1615),
.B1(n_1628),
.B2(n_1608),
.Y(n_1643)
);

NAND4xp25_ASAP7_75t_L g1644 ( 
.A(n_1643),
.B(n_1618),
.C(n_1623),
.D(n_1628),
.Y(n_1644)
);

OAI211xp5_ASAP7_75t_L g1645 ( 
.A1(n_1640),
.A2(n_1630),
.B(n_1623),
.C(n_1629),
.Y(n_1645)
);

AOI22xp5_ASAP7_75t_L g1646 ( 
.A1(n_1637),
.A2(n_1593),
.B1(n_1607),
.B2(n_1611),
.Y(n_1646)
);

NOR3xp33_ASAP7_75t_SL g1647 ( 
.A(n_1634),
.B(n_1609),
.C(n_1601),
.Y(n_1647)
);

AOI221x1_ASAP7_75t_L g1648 ( 
.A1(n_1635),
.A2(n_1624),
.B1(n_1626),
.B2(n_1592),
.C(n_1606),
.Y(n_1648)
);

AND2x2_ASAP7_75t_L g1649 ( 
.A(n_1638),
.B(n_1607),
.Y(n_1649)
);

AOI31xp33_ASAP7_75t_L g1650 ( 
.A1(n_1633),
.A2(n_1593),
.A3(n_1589),
.B(n_1600),
.Y(n_1650)
);

OAI21xp5_ASAP7_75t_SL g1651 ( 
.A1(n_1639),
.A2(n_1641),
.B(n_1642),
.Y(n_1651)
);

AOI211x1_ASAP7_75t_L g1652 ( 
.A1(n_1632),
.A2(n_1616),
.B(n_1629),
.C(n_1609),
.Y(n_1652)
);

NAND2xp5_ASAP7_75t_L g1653 ( 
.A(n_1649),
.B(n_1632),
.Y(n_1653)
);

NAND2xp5_ASAP7_75t_L g1654 ( 
.A(n_1651),
.B(n_1636),
.Y(n_1654)
);

INVx1_ASAP7_75t_L g1655 ( 
.A(n_1648),
.Y(n_1655)
);

INVx1_ASAP7_75t_L g1656 ( 
.A(n_1650),
.Y(n_1656)
);

NAND3xp33_ASAP7_75t_L g1657 ( 
.A(n_1652),
.B(n_1605),
.C(n_1592),
.Y(n_1657)
);

HB1xp67_ASAP7_75t_L g1658 ( 
.A(n_1653),
.Y(n_1658)
);

INVxp67_ASAP7_75t_SL g1659 ( 
.A(n_1657),
.Y(n_1659)
);

NAND2xp5_ASAP7_75t_L g1660 ( 
.A(n_1656),
.B(n_1647),
.Y(n_1660)
);

INVxp67_ASAP7_75t_SL g1661 ( 
.A(n_1655),
.Y(n_1661)
);

NOR2xp67_ASAP7_75t_SL g1662 ( 
.A(n_1654),
.B(n_1645),
.Y(n_1662)
);

INVxp67_ASAP7_75t_L g1663 ( 
.A(n_1653),
.Y(n_1663)
);

AOI222xp33_ASAP7_75t_L g1664 ( 
.A1(n_1662),
.A2(n_1659),
.B1(n_1661),
.B2(n_1660),
.C1(n_1663),
.C2(n_1658),
.Y(n_1664)
);

XNOR2xp5_ASAP7_75t_L g1665 ( 
.A(n_1658),
.B(n_1644),
.Y(n_1665)
);

AOI22xp5_ASAP7_75t_L g1666 ( 
.A1(n_1662),
.A2(n_1646),
.B1(n_1607),
.B2(n_1611),
.Y(n_1666)
);

AOI221xp5_ASAP7_75t_L g1667 ( 
.A1(n_1662),
.A2(n_1601),
.B1(n_1606),
.B2(n_1605),
.C(n_1591),
.Y(n_1667)
);

NAND2xp33_ASAP7_75t_R g1668 ( 
.A(n_1660),
.B(n_1600),
.Y(n_1668)
);

AND2x2_ASAP7_75t_L g1669 ( 
.A(n_1666),
.B(n_1589),
.Y(n_1669)
);

NOR2xp33_ASAP7_75t_L g1670 ( 
.A(n_1665),
.B(n_1591),
.Y(n_1670)
);

CKINVDCx5p33_ASAP7_75t_R g1671 ( 
.A(n_1668),
.Y(n_1671)
);

INVx1_ASAP7_75t_L g1672 ( 
.A(n_1671),
.Y(n_1672)
);

OAI322xp33_ASAP7_75t_L g1673 ( 
.A1(n_1672),
.A2(n_1670),
.A3(n_1669),
.B1(n_1664),
.B2(n_1629),
.C1(n_1667),
.C2(n_1605),
.Y(n_1673)
);

NAND2x1_ASAP7_75t_L g1674 ( 
.A(n_1673),
.B(n_1591),
.Y(n_1674)
);

INVx1_ASAP7_75t_L g1675 ( 
.A(n_1674),
.Y(n_1675)
);

INVx1_ASAP7_75t_L g1676 ( 
.A(n_1675),
.Y(n_1676)
);

AO22x2_ASAP7_75t_L g1677 ( 
.A1(n_1676),
.A2(n_1592),
.B1(n_1606),
.B2(n_1580),
.Y(n_1677)
);

CKINVDCx20_ASAP7_75t_R g1678 ( 
.A(n_1676),
.Y(n_1678)
);

AOI21xp5_ASAP7_75t_L g1679 ( 
.A1(n_1678),
.A2(n_1564),
.B(n_1574),
.Y(n_1679)
);

AOI221xp5_ASAP7_75t_L g1680 ( 
.A1(n_1677),
.A2(n_1523),
.B1(n_1543),
.B2(n_1527),
.C(n_1554),
.Y(n_1680)
);

OAI21xp5_ASAP7_75t_SL g1681 ( 
.A1(n_1679),
.A2(n_1523),
.B(n_1586),
.Y(n_1681)
);

XNOR2xp5_ASAP7_75t_L g1682 ( 
.A(n_1680),
.B(n_1529),
.Y(n_1682)
);

AOI22xp5_ASAP7_75t_L g1683 ( 
.A1(n_1682),
.A2(n_1523),
.B1(n_1543),
.B2(n_1527),
.Y(n_1683)
);

INVx2_ASAP7_75t_L g1684 ( 
.A(n_1681),
.Y(n_1684)
);

A2O1A1Ixp33_ASAP7_75t_SL g1685 ( 
.A1(n_1684),
.A2(n_1527),
.B(n_1554),
.C(n_1508),
.Y(n_1685)
);

AOI211xp5_ASAP7_75t_L g1686 ( 
.A1(n_1685),
.A2(n_1683),
.B(n_1554),
.C(n_1539),
.Y(n_1686)
);


endmodule