module fake_jpeg_21839_n_330 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_330);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_330;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_260;
wire n_199;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_13),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_5),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_0),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_15),
.Y(n_21)
);

BUFx10_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_7),
.B(n_10),
.Y(n_23)
);

INVx11_ASAP7_75t_SL g24 ( 
.A(n_13),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_9),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_6),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

INVxp67_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_5),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_14),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_18),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_36),
.B(n_37),
.Y(n_63)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_18),
.Y(n_37)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_18),
.Y(n_38)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_38),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_18),
.Y(n_39)
);

INVx5_ASAP7_75t_L g47 ( 
.A(n_39),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_SL g40 ( 
.A(n_23),
.B(n_8),
.Y(n_40)
);

AND2x2_ASAP7_75t_L g51 ( 
.A(n_40),
.B(n_15),
.Y(n_51)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_18),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_41),
.B(n_43),
.Y(n_64)
);

INVx11_ASAP7_75t_L g42 ( 
.A(n_22),
.Y(n_42)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_42),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_23),
.B(n_8),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_29),
.Y(n_44)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_44),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_29),
.Y(n_45)
);

INVx5_ASAP7_75t_L g48 ( 
.A(n_45),
.Y(n_48)
);

INVx3_ASAP7_75t_SL g46 ( 
.A(n_29),
.Y(n_46)
);

INVx2_ASAP7_75t_SL g49 ( 
.A(n_46),
.Y(n_49)
);

INVx5_ASAP7_75t_L g50 ( 
.A(n_45),
.Y(n_50)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_50),
.Y(n_81)
);

AND2x2_ASAP7_75t_L g92 ( 
.A(n_51),
.B(n_14),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_45),
.Y(n_53)
);

INVx11_ASAP7_75t_L g70 ( 
.A(n_53),
.Y(n_70)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_45),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_55),
.B(n_56),
.Y(n_79)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

OR2x2_ASAP7_75t_SL g57 ( 
.A(n_40),
.B(n_31),
.Y(n_57)
);

OR2x2_ASAP7_75t_SL g71 ( 
.A(n_57),
.B(n_31),
.Y(n_71)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_44),
.Y(n_58)
);

INVx5_ASAP7_75t_L g107 ( 
.A(n_58),
.Y(n_107)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_42),
.Y(n_59)
);

INVx4_ASAP7_75t_SL g84 ( 
.A(n_59),
.Y(n_84)
);

HB1xp67_ASAP7_75t_L g60 ( 
.A(n_39),
.Y(n_60)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_60),
.Y(n_94)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_39),
.Y(n_61)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_61),
.Y(n_104)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_44),
.Y(n_65)
);

HB1xp67_ASAP7_75t_L g72 ( 
.A(n_65),
.Y(n_72)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_46),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_66),
.A2(n_46),
.B1(n_42),
.B2(n_38),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_43),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_67),
.Y(n_74)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_46),
.Y(n_68)
);

INVx1_ASAP7_75t_SL g80 ( 
.A(n_68),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_SL g69 ( 
.A(n_64),
.B(n_40),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_69),
.B(n_71),
.Y(n_115)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_52),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_73),
.B(n_77),
.Y(n_116)
);

BUFx12f_ASAP7_75t_L g75 ( 
.A(n_55),
.Y(n_75)
);

CKINVDCx14_ASAP7_75t_R g121 ( 
.A(n_75),
.Y(n_121)
);

O2A1O1Ixp33_ASAP7_75t_SL g76 ( 
.A1(n_63),
.A2(n_31),
.B(n_41),
.C(n_37),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_76),
.A2(n_97),
.B1(n_107),
.B2(n_84),
.Y(n_128)
);

BUFx8_ASAP7_75t_L g77 ( 
.A(n_47),
.Y(n_77)
);

CKINVDCx14_ASAP7_75t_R g137 ( 
.A(n_78),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_52),
.A2(n_46),
.B1(n_42),
.B2(n_27),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_82),
.A2(n_33),
.B1(n_20),
.B2(n_25),
.Y(n_134)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_58),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_83),
.B(n_86),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_51),
.B(n_21),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_85),
.B(n_87),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_57),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_62),
.B(n_21),
.Y(n_87)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_53),
.Y(n_88)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_88),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_54),
.B(n_17),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_89),
.B(n_90),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_54),
.B(n_17),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_47),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_91),
.B(n_92),
.Y(n_135)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_48),
.Y(n_93)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_93),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_49),
.A2(n_24),
.B1(n_27),
.B2(n_38),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_95),
.A2(n_98),
.B1(n_105),
.B2(n_106),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_59),
.B(n_26),
.Y(n_96)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_96),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_66),
.A2(n_38),
.B1(n_41),
.B2(n_37),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_49),
.A2(n_24),
.B1(n_30),
.B2(n_26),
.Y(n_98)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_48),
.Y(n_99)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_99),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_SL g100 ( 
.A(n_50),
.B(n_16),
.Y(n_100)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_100),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_51),
.B(n_30),
.Y(n_101)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_101),
.Y(n_127)
);

INVx1_ASAP7_75t_SL g102 ( 
.A(n_60),
.Y(n_102)
);

INVx4_ASAP7_75t_L g112 ( 
.A(n_102),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_51),
.B(n_28),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_103),
.B(n_25),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_49),
.A2(n_36),
.B1(n_20),
.B2(n_34),
.Y(n_105)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_48),
.Y(n_106)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_60),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_108),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_110),
.B(n_125),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_76),
.B(n_36),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_111),
.B(n_114),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_74),
.B(n_22),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_105),
.B(n_22),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_119),
.B(n_133),
.Y(n_142)
);

INVx8_ASAP7_75t_L g120 ( 
.A(n_75),
.Y(n_120)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_120),
.Y(n_148)
);

INVx4_ASAP7_75t_L g126 ( 
.A(n_102),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_126),
.B(n_130),
.Y(n_145)
);

OAI21xp33_ASAP7_75t_SL g157 ( 
.A1(n_128),
.A2(n_136),
.B(n_33),
.Y(n_157)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_75),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_L g131 ( 
.A1(n_71),
.A2(n_35),
.B1(n_34),
.B2(n_16),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_131),
.A2(n_138),
.B1(n_98),
.B2(n_95),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_92),
.B(n_22),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_134),
.A2(n_19),
.B1(n_106),
.B2(n_99),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_SL g136 ( 
.A1(n_107),
.A2(n_35),
.B1(n_28),
.B2(n_19),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_97),
.A2(n_80),
.B1(n_73),
.B2(n_84),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_L g139 ( 
.A1(n_111),
.A2(n_80),
.B(n_82),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_SL g178 ( 
.A1(n_139),
.A2(n_149),
.B(n_150),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_140),
.B(n_143),
.Y(n_194)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_114),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_116),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_144),
.B(n_146),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_129),
.B(n_79),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_129),
.B(n_94),
.Y(n_147)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_147),
.Y(n_172)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_138),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_112),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_120),
.B(n_81),
.Y(n_151)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_151),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_112),
.B(n_81),
.Y(n_152)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_152),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_126),
.B(n_93),
.Y(n_153)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_153),
.Y(n_199)
);

CKINVDCx16_ASAP7_75t_R g154 ( 
.A(n_123),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_SL g193 ( 
.A(n_154),
.B(n_164),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_155),
.A2(n_158),
.B1(n_169),
.B2(n_170),
.Y(n_173)
);

AO21x1_ASAP7_75t_L g156 ( 
.A1(n_137),
.A2(n_78),
.B(n_72),
.Y(n_156)
);

AOI21xp5_ASAP7_75t_L g191 ( 
.A1(n_156),
.A2(n_117),
.B(n_109),
.Y(n_191)
);

INVx1_ASAP7_75t_SL g190 ( 
.A(n_157),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_119),
.A2(n_83),
.B1(n_108),
.B2(n_70),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_115),
.B(n_104),
.C(n_77),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_159),
.B(n_165),
.C(n_109),
.Y(n_179)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_132),
.Y(n_160)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_160),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_110),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_161),
.Y(n_184)
);

INVxp33_ASAP7_75t_L g162 ( 
.A(n_123),
.Y(n_162)
);

INVxp67_ASAP7_75t_SL g175 ( 
.A(n_162),
.Y(n_175)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_128),
.Y(n_163)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_163),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_130),
.B(n_77),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_135),
.B(n_22),
.C(n_70),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_125),
.B(n_32),
.Y(n_166)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_166),
.Y(n_177)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_134),
.Y(n_167)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_167),
.Y(n_180)
);

NAND3xp33_ASAP7_75t_L g168 ( 
.A(n_127),
.B(n_9),
.C(n_14),
.Y(n_168)
);

NOR2xp67_ASAP7_75t_L g188 ( 
.A(n_168),
.B(n_124),
.Y(n_188)
);

AO22x1_ASAP7_75t_SL g169 ( 
.A1(n_122),
.A2(n_33),
.B1(n_22),
.B2(n_2),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_127),
.A2(n_33),
.B1(n_1),
.B2(n_2),
.Y(n_170)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_171),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_SL g227 ( 
.A1(n_179),
.A2(n_182),
.B(n_191),
.Y(n_227)
);

AND2x2_ASAP7_75t_SL g182 ( 
.A(n_142),
.B(n_133),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_142),
.B(n_135),
.C(n_113),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_183),
.B(n_189),
.C(n_204),
.Y(n_209)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_145),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_185),
.B(n_186),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_147),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g187 ( 
.A(n_141),
.B(n_124),
.Y(n_187)
);

XOR2xp5_ASAP7_75t_L g207 ( 
.A(n_187),
.B(n_139),
.Y(n_207)
);

INVxp67_ASAP7_75t_L g232 ( 
.A(n_188),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_143),
.B(n_113),
.C(n_117),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_SL g192 ( 
.A(n_141),
.B(n_7),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_192),
.B(n_6),
.Y(n_221)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_158),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_197),
.B(n_200),
.Y(n_218)
);

AOI21xp5_ASAP7_75t_L g198 ( 
.A1(n_156),
.A2(n_121),
.B(n_118),
.Y(n_198)
);

AOI21xp5_ASAP7_75t_L g211 ( 
.A1(n_198),
.A2(n_156),
.B(n_169),
.Y(n_211)
);

INVxp67_ASAP7_75t_L g200 ( 
.A(n_169),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_146),
.Y(n_202)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_202),
.Y(n_205)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_170),
.Y(n_203)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_203),
.Y(n_208)
);

XOR2xp5_ASAP7_75t_L g204 ( 
.A(n_165),
.B(n_123),
.Y(n_204)
);

XOR2xp5_ASAP7_75t_L g236 ( 
.A(n_207),
.B(n_212),
.Y(n_236)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_175),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_210),
.B(n_214),
.Y(n_246)
);

OAI21xp33_ASAP7_75t_SL g234 ( 
.A1(n_211),
.A2(n_226),
.B(n_192),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_SL g212 ( 
.A(n_194),
.B(n_140),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_176),
.A2(n_163),
.B1(n_149),
.B2(n_167),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_213),
.A2(n_228),
.B1(n_203),
.B2(n_173),
.Y(n_243)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_193),
.Y(n_214)
);

OR2x2_ASAP7_75t_L g215 ( 
.A(n_184),
.B(n_161),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_215),
.B(n_224),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_204),
.B(n_159),
.C(n_160),
.Y(n_216)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_216),
.B(n_219),
.Y(n_245)
);

XNOR2x1_ASAP7_75t_L g217 ( 
.A(n_178),
.B(n_144),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_SL g252 ( 
.A(n_217),
.B(n_222),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_179),
.B(n_150),
.C(n_155),
.Y(n_219)
);

AND2x2_ASAP7_75t_SL g220 ( 
.A(n_196),
.B(n_148),
.Y(n_220)
);

OAI21xp33_ASAP7_75t_L g239 ( 
.A1(n_220),
.A2(n_180),
.B(n_197),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_221),
.B(n_223),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_SL g222 ( 
.A(n_182),
.B(n_11),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_178),
.B(n_183),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_187),
.B(n_148),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_196),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_225),
.B(n_229),
.Y(n_250)
);

MAJx2_ASAP7_75t_L g226 ( 
.A(n_182),
.B(n_4),
.C(n_13),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_200),
.A2(n_118),
.B1(n_4),
.B2(n_11),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_189),
.Y(n_229)
);

INVxp67_ASAP7_75t_L g230 ( 
.A(n_191),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_230),
.B(n_231),
.Y(n_235)
);

CKINVDCx16_ASAP7_75t_R g231 ( 
.A(n_198),
.Y(n_231)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_206),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_233),
.B(n_238),
.Y(n_257)
);

XOR2xp5_ASAP7_75t_SL g270 ( 
.A(n_234),
.B(n_237),
.Y(n_270)
);

NAND2x1p5_ASAP7_75t_L g237 ( 
.A(n_217),
.B(n_176),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_218),
.Y(n_238)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_239),
.Y(n_256)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_220),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_240),
.B(n_241),
.Y(n_263)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_220),
.Y(n_241)
);

HB1xp67_ASAP7_75t_L g242 ( 
.A(n_208),
.Y(n_242)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_242),
.Y(n_262)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_243),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_L g244 ( 
.A1(n_230),
.A2(n_180),
.B1(n_190),
.B2(n_172),
.Y(n_244)
);

CKINVDCx16_ASAP7_75t_R g268 ( 
.A(n_244),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_227),
.A2(n_190),
.B1(n_172),
.B2(n_173),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_247),
.B(n_252),
.Y(n_271)
);

INVxp67_ASAP7_75t_L g249 ( 
.A(n_213),
.Y(n_249)
);

AOI21xp5_ASAP7_75t_L g258 ( 
.A1(n_249),
.A2(n_254),
.B(n_255),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_219),
.A2(n_185),
.B1(n_174),
.B2(n_195),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_251),
.B(n_212),
.C(n_209),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_215),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_222),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_SL g259 ( 
.A(n_237),
.B(n_223),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_259),
.B(n_269),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_SL g276 ( 
.A(n_260),
.B(n_253),
.Y(n_276)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_237),
.Y(n_261)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_261),
.Y(n_275)
);

AND2x2_ASAP7_75t_L g264 ( 
.A(n_236),
.B(n_216),
.Y(n_264)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_264),
.Y(n_279)
);

INVx1_ASAP7_75t_SL g265 ( 
.A(n_235),
.Y(n_265)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_265),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_245),
.B(n_209),
.C(n_207),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_267),
.B(n_273),
.C(n_274),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_236),
.B(n_245),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_L g288 ( 
.A(n_271),
.B(n_272),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_251),
.B(n_224),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_248),
.B(n_205),
.C(n_201),
.Y(n_273)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_253),
.B(n_221),
.Y(n_274)
);

OAI21xp5_ASAP7_75t_SL g297 ( 
.A1(n_276),
.A2(n_286),
.B(n_262),
.Y(n_297)
);

INVx13_ASAP7_75t_L g277 ( 
.A(n_265),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_277),
.B(n_281),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_L g278 ( 
.A1(n_268),
.A2(n_249),
.B1(n_243),
.B2(n_250),
.Y(n_278)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_278),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_SL g281 ( 
.A(n_273),
.B(n_199),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_256),
.A2(n_239),
.B1(n_232),
.B2(n_246),
.Y(n_282)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_282),
.Y(n_298)
);

FAx1_ASAP7_75t_L g283 ( 
.A(n_270),
.B(n_252),
.CI(n_226),
.CON(n_283),
.SN(n_283)
);

AOI22xp5_ASAP7_75t_SL g294 ( 
.A1(n_283),
.A2(n_275),
.B1(n_279),
.B2(n_286),
.Y(n_294)
);

CKINVDCx16_ASAP7_75t_R g285 ( 
.A(n_257),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_SL g303 ( 
.A(n_285),
.B(n_289),
.Y(n_303)
);

INVxp67_ASAP7_75t_L g286 ( 
.A(n_263),
.Y(n_286)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_258),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_266),
.A2(n_232),
.B1(n_181),
.B2(n_177),
.Y(n_290)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_290),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_SL g291 ( 
.A(n_283),
.B(n_270),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_291),
.B(n_292),
.C(n_296),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_288),
.B(n_260),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_SL g306 ( 
.A(n_294),
.B(n_282),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_L g295 ( 
.A(n_284),
.B(n_267),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_295),
.B(n_287),
.Y(n_305)
);

XOR2xp5_ASAP7_75t_L g296 ( 
.A(n_287),
.B(n_269),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_297),
.B(n_259),
.C(n_274),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_SL g301 ( 
.A(n_290),
.B(n_181),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_SL g309 ( 
.A(n_301),
.B(n_288),
.Y(n_309)
);

INVx1_ASAP7_75t_SL g302 ( 
.A(n_277),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_SL g308 ( 
.A(n_302),
.B(n_177),
.Y(n_308)
);

OAI21xp5_ASAP7_75t_L g304 ( 
.A1(n_303),
.A2(n_284),
.B(n_280),
.Y(n_304)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_304),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_305),
.B(n_310),
.C(n_311),
.Y(n_316)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_306),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_308),
.B(n_294),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_309),
.B(n_298),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_296),
.B(n_264),
.C(n_283),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_302),
.B(n_299),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_312),
.B(n_300),
.Y(n_313)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_313),
.Y(n_323)
);

XNOR2xp5_ASAP7_75t_L g315 ( 
.A(n_307),
.B(n_292),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_315),
.B(n_317),
.Y(n_320)
);

AOI21xp5_ASAP7_75t_SL g321 ( 
.A1(n_319),
.A2(n_293),
.B(n_308),
.Y(n_321)
);

OAI211xp5_ASAP7_75t_L g324 ( 
.A1(n_321),
.A2(n_322),
.B(n_317),
.C(n_11),
.Y(n_324)
);

AOI21xp5_ASAP7_75t_SL g322 ( 
.A1(n_314),
.A2(n_291),
.B(n_4),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_SL g326 ( 
.A(n_324),
.B(n_325),
.Y(n_326)
);

OAI21x1_ASAP7_75t_L g325 ( 
.A1(n_320),
.A2(n_318),
.B(n_316),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_326),
.B(n_323),
.Y(n_327)
);

OAI321xp33_ASAP7_75t_L g328 ( 
.A1(n_327),
.A2(n_12),
.A3(n_1),
.B1(n_2),
.B2(n_3),
.C(n_0),
.Y(n_328)
);

FAx1_ASAP7_75t_SL g329 ( 
.A(n_328),
.B(n_0),
.CI(n_1),
.CON(n_329),
.SN(n_329)
);

NAND2xp5_ASAP7_75t_SL g330 ( 
.A(n_329),
.B(n_12),
.Y(n_330)
);


endmodule