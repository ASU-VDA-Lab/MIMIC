module fake_jpeg_19209_n_213 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_213);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_213;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx12_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

INVx2_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_13),
.Y(n_18)
);

BUFx12_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_13),
.Y(n_20)
);

INVx3_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_3),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

INVxp67_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_14),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_4),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_21),
.Y(n_33)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_33),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_25),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_34),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_32),
.Y(n_35)
);

CKINVDCx16_ASAP7_75t_R g61 ( 
.A(n_35),
.Y(n_61)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_21),
.Y(n_36)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_36),
.Y(n_56)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_21),
.Y(n_37)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_37),
.Y(n_59)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_29),
.Y(n_38)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_38),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_25),
.Y(n_39)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_39),
.Y(n_49)
);

BUFx5_ASAP7_75t_L g40 ( 
.A(n_25),
.Y(n_40)
);

BUFx16f_ASAP7_75t_L g65 ( 
.A(n_40),
.Y(n_65)
);

BUFx5_ASAP7_75t_L g41 ( 
.A(n_16),
.Y(n_41)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_41),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_32),
.B(n_0),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_42),
.B(n_32),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_18),
.B(n_14),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_43),
.B(n_44),
.Y(n_47)
);

INVx1_ASAP7_75t_SL g44 ( 
.A(n_29),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_38),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_45),
.B(n_68),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_48),
.B(n_50),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_42),
.B(n_17),
.Y(n_50)
);

HAxp5_ASAP7_75t_SL g51 ( 
.A(n_44),
.B(n_16),
.CON(n_51),
.SN(n_51)
);

OR2x2_ASAP7_75t_L g94 ( 
.A(n_51),
.B(n_2),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g54 ( 
.A1(n_36),
.A2(n_17),
.B1(n_31),
.B2(n_22),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_54),
.A2(n_55),
.B1(n_45),
.B2(n_66),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_34),
.B(n_31),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_55),
.B(n_64),
.Y(n_72)
);

AND2x2_ASAP7_75t_SL g57 ( 
.A(n_34),
.B(n_27),
.Y(n_57)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_57),
.B(n_63),
.C(n_16),
.Y(n_80)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_39),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_58),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_33),
.A2(n_22),
.B1(n_24),
.B2(n_30),
.Y(n_60)
);

CKINVDCx16_ASAP7_75t_R g91 ( 
.A(n_60),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_37),
.A2(n_30),
.B1(n_18),
.B2(n_20),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_62),
.A2(n_19),
.B1(n_23),
.B2(n_26),
.Y(n_87)
);

AND2x2_ASAP7_75t_SL g63 ( 
.A(n_39),
.B(n_27),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_35),
.B(n_27),
.Y(n_64)
);

CKINVDCx12_ASAP7_75t_R g67 ( 
.A(n_41),
.Y(n_67)
);

CKINVDCx16_ASAP7_75t_R g95 ( 
.A(n_67),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_37),
.B(n_20),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_40),
.B(n_26),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_69),
.B(n_23),
.Y(n_74)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_52),
.Y(n_71)
);

INVx4_ASAP7_75t_L g112 ( 
.A(n_71),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_73),
.A2(n_9),
.B1(n_11),
.B2(n_15),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_74),
.B(n_89),
.Y(n_107)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_66),
.Y(n_75)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_75),
.Y(n_100)
);

O2A1O1Ixp33_ASAP7_75t_SL g76 ( 
.A1(n_51),
.A2(n_28),
.B(n_16),
.C(n_19),
.Y(n_76)
);

O2A1O1Ixp33_ASAP7_75t_L g111 ( 
.A1(n_76),
.A2(n_65),
.B(n_8),
.C(n_9),
.Y(n_111)
);

INVx5_ASAP7_75t_L g77 ( 
.A(n_46),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_77),
.Y(n_121)
);

AND2x2_ASAP7_75t_L g78 ( 
.A(n_50),
.B(n_48),
.Y(n_78)
);

OAI21xp5_ASAP7_75t_L g104 ( 
.A1(n_78),
.A2(n_82),
.B(n_92),
.Y(n_104)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_80),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_47),
.B(n_24),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_SL g122 ( 
.A(n_81),
.B(n_88),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_SL g82 ( 
.A1(n_57),
.A2(n_16),
.B(n_19),
.Y(n_82)
);

BUFx12_ASAP7_75t_L g83 ( 
.A(n_52),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_83),
.B(n_84),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_60),
.Y(n_84)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_54),
.Y(n_86)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_86),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_87),
.A2(n_90),
.B1(n_93),
.B2(n_94),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_64),
.B(n_26),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_57),
.B(n_0),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_53),
.A2(n_19),
.B1(n_23),
.B2(n_3),
.Y(n_90)
);

AND2x2_ASAP7_75t_L g92 ( 
.A(n_63),
.B(n_1),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_53),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_93)
);

INVx8_ASAP7_75t_L g96 ( 
.A(n_46),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_96),
.B(n_97),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_69),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_L g98 ( 
.A1(n_63),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_98),
.A2(n_99),
.B1(n_65),
.B2(n_89),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_L g99 ( 
.A1(n_56),
.A2(n_4),
.B1(n_5),
.B2(n_7),
.Y(n_99)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_85),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_102),
.B(n_119),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_86),
.A2(n_49),
.B1(n_58),
.B2(n_56),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_103),
.A2(n_106),
.B1(n_111),
.B2(n_114),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_91),
.A2(n_49),
.B1(n_59),
.B2(n_61),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_70),
.B(n_59),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_110),
.B(n_113),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_70),
.B(n_7),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_84),
.A2(n_65),
.B1(n_9),
.B2(n_8),
.Y(n_114)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_85),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_115),
.B(n_118),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_116),
.A2(n_72),
.B1(n_94),
.B2(n_97),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_78),
.B(n_11),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_117),
.B(n_78),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_79),
.B(n_15),
.Y(n_118)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_83),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_123),
.B(n_92),
.Y(n_142)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_100),
.Y(n_126)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_126),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_100),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_127),
.B(n_128),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_105),
.Y(n_128)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_121),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_129),
.B(n_135),
.Y(n_160)
);

OR2x2_ASAP7_75t_L g130 ( 
.A(n_101),
.B(n_76),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_L g154 ( 
.A1(n_130),
.A2(n_144),
.B(n_145),
.Y(n_154)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_103),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_131),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_132),
.A2(n_142),
.B1(n_112),
.B2(n_95),
.Y(n_162)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_120),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_133),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_122),
.B(n_83),
.Y(n_137)
);

INVxp67_ASAP7_75t_L g150 ( 
.A(n_137),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_109),
.B(n_80),
.C(n_72),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_138),
.B(n_141),
.C(n_143),
.Y(n_155)
);

AO22x1_ASAP7_75t_L g139 ( 
.A1(n_110),
.A2(n_73),
.B1(n_74),
.B2(n_76),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_139),
.B(n_140),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_120),
.Y(n_140)
);

XOR2xp5_ASAP7_75t_L g141 ( 
.A(n_104),
.B(n_107),
.Y(n_141)
);

XOR2xp5_ASAP7_75t_L g143 ( 
.A(n_104),
.B(n_82),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_108),
.A2(n_92),
.B1(n_75),
.B2(n_77),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_116),
.B(n_71),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_136),
.A2(n_109),
.B1(n_111),
.B2(n_113),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_147),
.A2(n_161),
.B1(n_132),
.B2(n_131),
.Y(n_169)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_124),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_148),
.B(n_152),
.Y(n_166)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_129),
.Y(n_152)
);

AOI21xp5_ASAP7_75t_L g153 ( 
.A1(n_130),
.A2(n_106),
.B(n_114),
.Y(n_153)
);

AND2x2_ASAP7_75t_L g175 ( 
.A(n_153),
.B(n_157),
.Y(n_175)
);

XNOR2x1_ASAP7_75t_SL g156 ( 
.A(n_143),
.B(n_141),
.Y(n_156)
);

OA21x2_ASAP7_75t_SL g167 ( 
.A1(n_156),
.A2(n_135),
.B(n_134),
.Y(n_167)
);

AOI21xp5_ASAP7_75t_L g157 ( 
.A1(n_133),
.A2(n_117),
.B(n_119),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_136),
.A2(n_107),
.B1(n_96),
.B2(n_102),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_162),
.B(n_128),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_163),
.B(n_164),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_155),
.B(n_138),
.C(n_139),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_155),
.B(n_139),
.C(n_134),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_L g180 ( 
.A1(n_165),
.A2(n_172),
.B(n_157),
.Y(n_180)
);

XNOR2x1_ASAP7_75t_L g181 ( 
.A(n_167),
.B(n_173),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_146),
.B(n_127),
.Y(n_168)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_168),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_169),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_149),
.B(n_125),
.Y(n_170)
);

BUFx24_ASAP7_75t_SL g184 ( 
.A(n_170),
.Y(n_184)
);

INVx1_ASAP7_75t_SL g171 ( 
.A(n_158),
.Y(n_171)
);

HB1xp67_ASAP7_75t_L g183 ( 
.A(n_171),
.Y(n_183)
);

NAND3xp33_ASAP7_75t_L g172 ( 
.A(n_156),
.B(n_126),
.C(n_144),
.Y(n_172)
);

XOR2xp5_ASAP7_75t_L g173 ( 
.A(n_146),
.B(n_112),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_150),
.B(n_121),
.Y(n_174)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_174),
.Y(n_187)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_160),
.Y(n_176)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_176),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g188 ( 
.A(n_180),
.B(n_164),
.Y(n_188)
);

AOI21xp5_ASAP7_75t_SL g182 ( 
.A1(n_168),
.A2(n_154),
.B(n_153),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g189 ( 
.A(n_182),
.B(n_185),
.Y(n_189)
);

AOI21xp5_ASAP7_75t_SL g185 ( 
.A1(n_175),
.A2(n_154),
.B(n_162),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g201 ( 
.A(n_188),
.B(n_194),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_186),
.B(n_150),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_190),
.B(n_191),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_177),
.B(n_165),
.C(n_173),
.Y(n_191)
);

AND2x4_ASAP7_75t_L g192 ( 
.A(n_181),
.B(n_175),
.Y(n_192)
);

INVxp33_ASAP7_75t_L g198 ( 
.A(n_192),
.Y(n_198)
);

AOI22xp33_ASAP7_75t_SL g193 ( 
.A1(n_187),
.A2(n_148),
.B1(n_151),
.B2(n_171),
.Y(n_193)
);

NAND4xp25_ASAP7_75t_L g199 ( 
.A(n_193),
.B(n_195),
.C(n_159),
.D(n_183),
.Y(n_199)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_183),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_178),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_188),
.B(n_179),
.C(n_169),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_197),
.B(n_200),
.C(n_161),
.Y(n_203)
);

AO21x1_ASAP7_75t_L g202 ( 
.A1(n_199),
.A2(n_193),
.B(n_166),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_189),
.B(n_147),
.C(n_175),
.Y(n_200)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_202),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_L g206 ( 
.A(n_203),
.B(n_204),
.Y(n_206)
);

HB1xp67_ASAP7_75t_L g204 ( 
.A(n_197),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_196),
.B(n_184),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_205),
.B(n_201),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_207),
.B(n_192),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_206),
.B(n_192),
.C(n_198),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_209),
.B(n_210),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_211),
.A2(n_208),
.B1(n_206),
.B2(n_198),
.Y(n_212)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_212),
.B(n_152),
.Y(n_213)
);


endmodule