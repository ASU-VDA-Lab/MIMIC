module real_jpeg_25004_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_80;
wire n_30;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_323;
wire n_166;
wire n_176;
wire n_215;
wire n_286;
wire n_312;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

INVxp67_ASAP7_75t_L g64 ( 
.A(n_0),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_0),
.B(n_67),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_0),
.B(n_27),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_0),
.B(n_141),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_0),
.B(n_17),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_0),
.B(n_33),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_0),
.B(n_52),
.Y(n_272)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_1),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_2),
.B(n_43),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_2),
.B(n_27),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_2),
.B(n_33),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_2),
.B(n_17),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_2),
.B(n_52),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_2),
.B(n_49),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_2),
.B(n_47),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_2),
.B(n_67),
.Y(n_266)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_3),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_4),
.B(n_47),
.Y(n_46)
);

INVxp67_ASAP7_75t_L g61 ( 
.A(n_4),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_4),
.B(n_67),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_4),
.B(n_229),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_4),
.B(n_33),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_4),
.B(n_52),
.Y(n_286)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_5),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_6),
.B(n_49),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_6),
.B(n_47),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_6),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_6),
.B(n_52),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_6),
.B(n_67),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_6),
.B(n_17),
.Y(n_265)
);

INVx8_ASAP7_75t_SL g28 ( 
.A(n_7),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_8),
.B(n_71),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_8),
.B(n_52),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_8),
.B(n_33),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_8),
.B(n_182),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_8),
.B(n_49),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_8),
.B(n_47),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_8),
.B(n_67),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_8),
.B(n_27),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_9),
.B(n_49),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_9),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_9),
.B(n_33),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_9),
.B(n_47),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_9),
.B(n_67),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_9),
.B(n_27),
.Y(n_241)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_10),
.Y(n_47)
);

CKINVDCx14_ASAP7_75t_R g25 ( 
.A(n_11),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_11),
.B(n_71),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_11),
.B(n_47),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_11),
.B(n_67),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_11),
.B(n_191),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_11),
.B(n_33),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_11),
.B(n_52),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_11),
.B(n_49),
.Y(n_271)
);

INVx13_ASAP7_75t_L g44 ( 
.A(n_12),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_13),
.B(n_33),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_13),
.B(n_52),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_13),
.B(n_49),
.Y(n_88)
);

CKINVDCx14_ASAP7_75t_R g113 ( 
.A(n_13),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_13),
.B(n_47),
.Y(n_144)
);

CKINVDCx14_ASAP7_75t_R g59 ( 
.A(n_14),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_14),
.B(n_71),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_14),
.B(n_160),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_14),
.B(n_33),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_14),
.B(n_52),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_14),
.B(n_49),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g253 ( 
.A(n_14),
.B(n_47),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_14),
.B(n_67),
.Y(n_287)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_15),
.Y(n_50)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_16),
.B(n_52),
.Y(n_83)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_17),
.Y(n_36)
);

INVx6_ASAP7_75t_L g161 ( 
.A(n_17),
.Y(n_161)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_17),
.Y(n_192)
);

INVx6_ASAP7_75t_L g230 ( 
.A(n_17),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_147),
.Y(n_18)
);

XOR2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_117),
.Y(n_19)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_78),
.C(n_90),
.Y(n_20)
);

XNOR2xp5_ASAP7_75t_L g323 ( 
.A(n_21),
.B(n_78),
.Y(n_323)
);

XNOR2xp5_ASAP7_75t_SL g21 ( 
.A(n_22),
.B(n_54),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_22),
.B(n_55),
.C(n_72),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_39),
.C(n_45),
.Y(n_22)
);

XOR2xp5_ASAP7_75t_L g316 ( 
.A(n_23),
.B(n_317),
.Y(n_316)
);

XNOR2xp5_ASAP7_75t_SL g23 ( 
.A(n_24),
.B(n_29),
.Y(n_23)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_24),
.B(n_30),
.C(n_37),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_26),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_26),
.B(n_59),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_26),
.B(n_61),
.Y(n_124)
);

CKINVDCx5p33_ASAP7_75t_R g26 ( 
.A(n_27),
.Y(n_26)
);

INVx8_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

AOI22xp5_ASAP7_75t_L g29 ( 
.A1(n_30),
.A2(n_35),
.B1(n_37),
.B2(n_38),
.Y(n_29)
);

CKINVDCx14_ASAP7_75t_R g38 ( 
.A(n_30),
.Y(n_38)
);

AOI22xp33_ASAP7_75t_L g81 ( 
.A1(n_30),
.A2(n_38),
.B1(n_82),
.B2(n_83),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_SL g131 ( 
.A(n_30),
.B(n_80),
.C(n_83),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_31),
.B(n_32),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_SL g35 ( 
.A(n_31),
.B(n_36),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_31),
.B(n_62),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_32),
.B(n_111),
.Y(n_110)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_35),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_35),
.A2(n_37),
.B1(n_40),
.B2(n_103),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_36),
.B(n_113),
.Y(n_112)
);

INVx3_ASAP7_75t_L g182 ( 
.A(n_36),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g39 ( 
.A(n_37),
.B(n_40),
.C(n_41),
.Y(n_39)
);

XNOR2xp5_ASAP7_75t_L g317 ( 
.A(n_39),
.B(n_45),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_40),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_41),
.A2(n_42),
.B1(n_101),
.B2(n_102),
.Y(n_100)
);

CKINVDCx16_ASAP7_75t_R g41 ( 
.A(n_42),
.Y(n_41)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx11_ASAP7_75t_L g71 ( 
.A(n_44),
.Y(n_71)
);

INVx8_ASAP7_75t_L g141 ( 
.A(n_44),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_44),
.B(n_177),
.Y(n_269)
);

BUFx24_ASAP7_75t_SL g325 ( 
.A(n_45),
.Y(n_325)
);

FAx1_ASAP7_75t_SL g45 ( 
.A(n_46),
.B(n_48),
.CI(n_51),
.CON(n_45),
.SN(n_45)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_46),
.B(n_48),
.C(n_51),
.Y(n_85)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_47),
.Y(n_65)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_49),
.Y(n_62)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx13_ASAP7_75t_L g178 ( 
.A(n_52),
.Y(n_178)
);

BUFx24_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

XNOR2xp5_ASAP7_75t_L g54 ( 
.A(n_55),
.B(n_72),
.Y(n_54)
);

MAJIxp5_ASAP7_75t_L g55 ( 
.A(n_56),
.B(n_66),
.C(n_70),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_56),
.A2(n_57),
.B1(n_105),
.B2(n_107),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_57),
.Y(n_56)
);

MAJIxp5_ASAP7_75t_L g57 ( 
.A(n_58),
.B(n_60),
.C(n_63),
.Y(n_57)
);

XNOR2xp5_ASAP7_75t_L g93 ( 
.A(n_58),
.B(n_63),
.Y(n_93)
);

XOR2xp5_ASAP7_75t_L g92 ( 
.A(n_60),
.B(n_93),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_61),
.B(n_62),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_62),
.B(n_64),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_64),
.B(n_65),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_66),
.A2(n_74),
.B1(n_75),
.B2(n_76),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_66),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_66),
.A2(n_70),
.B1(n_76),
.B2(n_106),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_66),
.B(n_75),
.C(n_77),
.Y(n_137)
);

BUFx12f_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx8_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_70),
.Y(n_106)
);

XOR2xp5_ASAP7_75t_L g72 ( 
.A(n_73),
.B(n_77),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_74),
.Y(n_75)
);

XOR2xp5_ASAP7_75t_L g78 ( 
.A(n_79),
.B(n_84),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_79),
.B(n_85),
.C(n_86),
.Y(n_134)
);

XOR2xp5_ASAP7_75t_L g79 ( 
.A(n_80),
.B(n_81),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_L g125 ( 
.A1(n_82),
.A2(n_83),
.B1(n_126),
.B2(n_127),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_83),
.Y(n_82)
);

XNOR2xp5_ASAP7_75t_L g84 ( 
.A(n_85),
.B(n_86),
.Y(n_84)
);

BUFx24_ASAP7_75t_SL g326 ( 
.A(n_86),
.Y(n_326)
);

FAx1_ASAP7_75t_SL g86 ( 
.A(n_87),
.B(n_88),
.CI(n_89),
.CON(n_86),
.SN(n_86)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_87),
.B(n_88),
.C(n_89),
.Y(n_130)
);

XNOR2xp5_ASAP7_75t_L g322 ( 
.A(n_90),
.B(n_323),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_104),
.C(n_108),
.Y(n_90)
);

XOR2xp5_ASAP7_75t_L g318 ( 
.A(n_91),
.B(n_319),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_92),
.B(n_94),
.C(n_100),
.Y(n_91)
);

XNOR2xp5_ASAP7_75t_L g301 ( 
.A(n_92),
.B(n_302),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_L g302 ( 
.A(n_94),
.B(n_100),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_97),
.C(n_98),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g282 ( 
.A1(n_95),
.A2(n_96),
.B1(n_98),
.B2(n_99),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_96),
.Y(n_95)
);

XOR2xp5_ASAP7_75t_L g281 ( 
.A(n_97),
.B(n_282),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_99),
.Y(n_98)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

XNOR2xp5_ASAP7_75t_L g319 ( 
.A(n_104),
.B(n_108),
.Y(n_319)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_105),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_109),
.B(n_115),
.C(n_116),
.Y(n_108)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_109),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_L g307 ( 
.A(n_109),
.B(n_308),
.Y(n_307)
);

FAx1_ASAP7_75t_SL g109 ( 
.A(n_110),
.B(n_112),
.CI(n_114),
.CON(n_109),
.SN(n_109)
);

XNOR2xp5_ASAP7_75t_L g308 ( 
.A(n_115),
.B(n_116),
.Y(n_308)
);

XNOR2xp5_ASAP7_75t_L g117 ( 
.A(n_118),
.B(n_119),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_120),
.A2(n_121),
.B1(n_132),
.B2(n_133),
.Y(n_119)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_122),
.A2(n_123),
.B1(n_128),
.B2(n_129),
.Y(n_121)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

XOR2xp5_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_125),
.Y(n_123)
);

CKINVDCx16_ASAP7_75t_R g127 ( 
.A(n_126),
.Y(n_127)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

XOR2xp5_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_131),
.Y(n_129)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_L g133 ( 
.A(n_134),
.B(n_135),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_136),
.A2(n_137),
.B1(n_138),
.B2(n_139),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

CKINVDCx16_ASAP7_75t_R g138 ( 
.A(n_139),
.Y(n_138)
);

XOR2xp5_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_142),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_143),
.A2(n_144),
.B1(n_145),
.B2(n_146),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_144),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_145),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_148),
.B(n_321),
.C(n_322),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_311),
.C(n_312),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_297),
.C(n_298),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_275),
.C(n_276),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_245),
.C(n_246),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_223),
.C(n_224),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_205),
.C(n_206),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_183),
.C(n_184),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_169),
.C(n_174),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_157),
.A2(n_158),
.B1(n_165),
.B2(n_166),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_157),
.B(n_167),
.C(n_168),
.Y(n_183)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_159),
.A2(n_162),
.B1(n_163),
.B2(n_164),
.Y(n_158)
);

CKINVDCx14_ASAP7_75t_R g164 ( 
.A(n_159),
.Y(n_164)
);

INVx5_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_162),
.B(n_164),
.Y(n_187)
);

CKINVDCx14_ASAP7_75t_R g162 ( 
.A(n_163),
.Y(n_162)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_SL g166 ( 
.A(n_167),
.B(n_168),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_170),
.B(n_172),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_170),
.A2(n_171),
.B1(n_172),
.B2(n_173),
.Y(n_175)
);

CKINVDCx16_ASAP7_75t_R g170 ( 
.A(n_171),
.Y(n_170)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_175),
.B(n_176),
.C(n_179),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_177),
.B(n_178),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_181),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_196),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_186),
.A2(n_187),
.B1(n_188),
.B2(n_189),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_186),
.B(n_189),
.C(n_196),
.Y(n_205)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_190),
.A2(n_193),
.B1(n_194),
.B2(n_195),
.Y(n_189)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_190),
.Y(n_195)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_193),
.B(n_195),
.Y(n_215)
);

CKINVDCx16_ASAP7_75t_R g193 ( 
.A(n_194),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_197),
.A2(n_198),
.B1(n_199),
.B2(n_204),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_197),
.Y(n_204)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_200),
.A2(n_201),
.B1(n_202),
.B2(n_203),
.Y(n_199)
);

CKINVDCx16_ASAP7_75t_R g203 ( 
.A(n_200),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_201),
.B(n_203),
.C(n_204),
.Y(n_208)
);

CKINVDCx14_ASAP7_75t_R g201 ( 
.A(n_202),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_SL g206 ( 
.A(n_207),
.B(n_214),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_209),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_208),
.B(n_209),
.C(n_214),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g209 ( 
.A(n_210),
.B(n_211),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_210),
.B(n_212),
.C(n_213),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_212),
.B(n_213),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_SL g214 ( 
.A(n_215),
.B(n_216),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_215),
.B(n_217),
.C(n_218),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g216 ( 
.A(n_217),
.B(n_218),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_219),
.A2(n_220),
.B1(n_221),
.B2(n_222),
.Y(n_218)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_219),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_220),
.B(n_222),
.Y(n_243)
);

CKINVDCx14_ASAP7_75t_R g220 ( 
.A(n_221),
.Y(n_220)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_225),
.B(n_239),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_225),
.B(n_240),
.C(n_244),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_SL g225 ( 
.A(n_226),
.B(n_235),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_227),
.B(n_234),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_227),
.B(n_234),
.C(n_235),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_228),
.A2(n_231),
.B1(n_232),
.B2(n_233),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_228),
.Y(n_233)
);

INVx5_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_231),
.B(n_233),
.Y(n_258)
);

CKINVDCx16_ASAP7_75t_R g231 ( 
.A(n_232),
.Y(n_231)
);

BUFx24_ASAP7_75t_SL g324 ( 
.A(n_235),
.Y(n_324)
);

FAx1_ASAP7_75t_SL g235 ( 
.A(n_236),
.B(n_237),
.CI(n_238),
.CON(n_235),
.SN(n_235)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_236),
.B(n_237),
.C(n_238),
.Y(n_260)
);

XOR2xp5_ASAP7_75t_L g239 ( 
.A(n_240),
.B(n_244),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_240),
.Y(n_262)
);

FAx1_ASAP7_75t_SL g240 ( 
.A(n_241),
.B(n_242),
.CI(n_243),
.CON(n_240),
.SN(n_240)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_247),
.B(n_261),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_248),
.A2(n_249),
.B1(n_250),
.B2(n_251),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_249),
.B(n_250),
.C(n_261),
.Y(n_275)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_SL g251 ( 
.A(n_252),
.B(n_256),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_252),
.B(n_257),
.C(n_260),
.Y(n_279)
);

BUFx24_ASAP7_75t_SL g328 ( 
.A(n_252),
.Y(n_328)
);

FAx1_ASAP7_75t_SL g252 ( 
.A(n_253),
.B(n_254),
.CI(n_255),
.CON(n_252),
.SN(n_252)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_253),
.B(n_254),
.C(n_255),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_257),
.A2(n_258),
.B1(n_259),
.B2(n_260),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

CKINVDCx16_ASAP7_75t_R g259 ( 
.A(n_260),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_SL g261 ( 
.A(n_262),
.B(n_263),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_262),
.B(n_268),
.C(n_273),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_264),
.A2(n_268),
.B1(n_273),
.B2(n_274),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_264),
.Y(n_273)
);

OAI21xp5_ASAP7_75t_L g264 ( 
.A1(n_265),
.A2(n_266),
.B(n_267),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_265),
.B(n_266),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g293 ( 
.A(n_267),
.B(n_294),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_267),
.B(n_294),
.C(n_295),
.Y(n_304)
);

CKINVDCx16_ASAP7_75t_R g274 ( 
.A(n_268),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_269),
.B(n_270),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_269),
.B(n_271),
.C(n_272),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_271),
.B(n_272),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_277),
.A2(n_278),
.B1(n_290),
.B2(n_296),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_277),
.B(n_291),
.C(n_292),
.Y(n_297)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_SL g278 ( 
.A(n_279),
.B(n_280),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_279),
.B(n_281),
.C(n_283),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_281),
.B(n_283),
.Y(n_280)
);

XOR2xp5_ASAP7_75t_L g283 ( 
.A(n_284),
.B(n_289),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_285),
.A2(n_286),
.B1(n_287),
.B2(n_288),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_285),
.B(n_288),
.C(n_289),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g285 ( 
.A(n_286),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_287),
.Y(n_288)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_290),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_SL g290 ( 
.A(n_291),
.B(n_292),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_293),
.B(n_295),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_299),
.A2(n_300),
.B1(n_309),
.B2(n_310),
.Y(n_298)
);

CKINVDCx14_ASAP7_75t_R g309 ( 
.A(n_299),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_300),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_SL g300 ( 
.A(n_301),
.B(n_303),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_301),
.B(n_303),
.C(n_309),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_L g303 ( 
.A(n_304),
.B(n_305),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_304),
.B(n_306),
.C(n_307),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_L g305 ( 
.A(n_306),
.B(n_307),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_L g312 ( 
.A(n_313),
.B(n_314),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_313),
.B(n_315),
.C(n_320),
.Y(n_321)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_315),
.A2(n_316),
.B1(n_318),
.B2(n_320),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_316),
.Y(n_315)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_318),
.Y(n_320)
);


endmodule