module real_aes_9121_n_102 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_102);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_102;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_742;
wire n_112;
wire n_364;
wire n_319;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_379;
wire n_374;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_564;
wire n_519;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_744;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_748;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_455;
wire n_310;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_527;
wire n_434;
wire n_505;
wire n_502;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_733;
wire n_552;
wire n_402;
wire n_602;
wire n_617;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_481;
wire n_148;
wire n_498;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_233;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_753;
wire n_314;
wire n_283;
wire n_252;
wire n_741;
wire n_249;
wire n_623;
wire n_721;
wire n_446;
wire n_221;
wire n_681;
wire n_156;
wire n_456;
wire n_359;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_479;
wire n_338;
wire n_442;
wire n_740;
wire n_371;
wire n_698;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_546;
wire n_151;
wire n_639;
wire n_587;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_241;
wire n_175;
wire n_687;
wire n_729;
wire n_646;
wire n_710;
wire n_650;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_554;
wire n_475;
wire n_264;
wire n_237;
wire n_668;
A2O1A1Ixp33_ASAP7_75t_SL g548 ( .A1(n_0), .A2(n_153), .B(n_549), .C(n_552), .Y(n_548) );
NAND2xp5_ASAP7_75t_L g553 ( .A(n_1), .B(n_493), .Y(n_553) );
INVx1_ASAP7_75t_L g109 ( .A(n_2), .Y(n_109) );
INVx1_ASAP7_75t_L g187 ( .A(n_3), .Y(n_187) );
NAND2xp5_ASAP7_75t_SL g527 ( .A(n_4), .B(n_145), .Y(n_527) );
AOI21xp5_ASAP7_75t_L g486 ( .A1(n_5), .A2(n_462), .B(n_487), .Y(n_486) );
AO21x2_ASAP7_75t_L g477 ( .A1(n_6), .A2(n_130), .B(n_478), .Y(n_477) );
AOI22xp33_ASAP7_75t_L g216 ( .A1(n_7), .A2(n_35), .B1(n_139), .B2(n_217), .Y(n_216) );
NAND2xp5_ASAP7_75t_L g156 ( .A(n_8), .B(n_130), .Y(n_156) );
AND2x6_ASAP7_75t_L g154 ( .A(n_9), .B(n_155), .Y(n_154) );
A2O1A1Ixp33_ASAP7_75t_L g451 ( .A1(n_10), .A2(n_154), .B(n_452), .C(n_454), .Y(n_451) );
NAND2xp5_ASAP7_75t_L g107 ( .A(n_11), .B(n_36), .Y(n_107) );
NOR2xp33_ASAP7_75t_L g438 ( .A(n_11), .B(n_36), .Y(n_438) );
INVx1_ASAP7_75t_L g135 ( .A(n_12), .Y(n_135) );
INVx1_ASAP7_75t_L g180 ( .A(n_13), .Y(n_180) );
NAND2xp5_ASAP7_75t_L g223 ( .A(n_14), .B(n_143), .Y(n_223) );
CKINVDCx20_ASAP7_75t_R g754 ( .A(n_15), .Y(n_754) );
NAND2xp5_ASAP7_75t_SL g483 ( .A(n_16), .B(n_145), .Y(n_483) );
NAND2xp5_ASAP7_75t_L g192 ( .A(n_17), .B(n_131), .Y(n_192) );
AO32x2_ASAP7_75t_L g214 ( .A1(n_18), .A2(n_130), .A3(n_160), .B1(n_171), .B2(n_215), .Y(n_214) );
NAND2xp5_ASAP7_75t_SL g227 ( .A(n_19), .B(n_139), .Y(n_227) );
NAND2xp5_ASAP7_75t_L g189 ( .A(n_20), .B(n_131), .Y(n_189) );
AOI22xp33_ASAP7_75t_L g218 ( .A1(n_21), .A2(n_54), .B1(n_139), .B2(n_217), .Y(n_218) );
AOI22xp33_ASAP7_75t_SL g239 ( .A1(n_22), .A2(n_81), .B1(n_139), .B2(n_143), .Y(n_239) );
NAND2xp5_ASAP7_75t_SL g209 ( .A(n_23), .B(n_139), .Y(n_209) );
A2O1A1Ixp33_ASAP7_75t_L g512 ( .A1(n_24), .A2(n_171), .B(n_452), .C(n_513), .Y(n_512) );
A2O1A1Ixp33_ASAP7_75t_L g480 ( .A1(n_25), .A2(n_171), .B(n_452), .C(n_481), .Y(n_480) );
BUFx6f_ASAP7_75t_L g147 ( .A(n_26), .Y(n_147) );
NAND2xp5_ASAP7_75t_L g172 ( .A(n_27), .B(n_173), .Y(n_172) );
AOI21xp5_ASAP7_75t_L g545 ( .A1(n_28), .A2(n_462), .B(n_546), .Y(n_545) );
NAND2xp5_ASAP7_75t_L g211 ( .A(n_29), .B(n_173), .Y(n_211) );
INVx2_ASAP7_75t_L g141 ( .A(n_30), .Y(n_141) );
A2O1A1Ixp33_ASAP7_75t_L g500 ( .A1(n_31), .A2(n_464), .B(n_472), .C(n_501), .Y(n_500) );
NAND2xp5_ASAP7_75t_SL g163 ( .A(n_32), .B(n_139), .Y(n_163) );
NAND2xp5_ASAP7_75t_L g229 ( .A(n_33), .B(n_173), .Y(n_229) );
NAND2xp5_ASAP7_75t_L g482 ( .A(n_34), .B(n_225), .Y(n_482) );
NAND2xp5_ASAP7_75t_L g510 ( .A(n_37), .B(n_511), .Y(n_510) );
CKINVDCx20_ASAP7_75t_R g458 ( .A(n_38), .Y(n_458) );
OAI22xp5_ASAP7_75t_L g115 ( .A1(n_39), .A2(n_78), .B1(n_116), .B2(n_117), .Y(n_115) );
CKINVDCx16_ASAP7_75t_R g117 ( .A(n_39), .Y(n_117) );
NAND2xp5_ASAP7_75t_L g470 ( .A(n_40), .B(n_145), .Y(n_470) );
AOI22xp33_ASAP7_75t_L g102 ( .A1(n_41), .A2(n_103), .B1(n_113), .B2(n_757), .Y(n_102) );
NAND2xp5_ASAP7_75t_L g479 ( .A(n_42), .B(n_462), .Y(n_479) );
OAI22xp5_ASAP7_75t_SL g744 ( .A1(n_43), .A2(n_79), .B1(n_433), .B2(n_745), .Y(n_744) );
CKINVDCx20_ASAP7_75t_R g745 ( .A(n_43), .Y(n_745) );
A2O1A1Ixp33_ASAP7_75t_L g463 ( .A1(n_44), .A2(n_464), .B(n_466), .C(n_472), .Y(n_463) );
NAND2xp5_ASAP7_75t_SL g138 ( .A(n_45), .B(n_139), .Y(n_138) );
INVx1_ASAP7_75t_L g550 ( .A(n_46), .Y(n_550) );
AOI22xp33_ASAP7_75t_L g237 ( .A1(n_47), .A2(n_90), .B1(n_217), .B2(n_238), .Y(n_237) );
INVx1_ASAP7_75t_L g467 ( .A(n_48), .Y(n_467) );
NAND2xp5_ASAP7_75t_SL g149 ( .A(n_49), .B(n_139), .Y(n_149) );
NAND2xp5_ASAP7_75t_L g182 ( .A(n_50), .B(n_139), .Y(n_182) );
NOR2xp33_ASAP7_75t_L g741 ( .A(n_51), .B(n_742), .Y(n_741) );
CKINVDCx20_ASAP7_75t_R g747 ( .A(n_51), .Y(n_747) );
NAND2xp5_ASAP7_75t_L g461 ( .A(n_52), .B(n_462), .Y(n_461) );
NAND2xp5_ASAP7_75t_L g150 ( .A(n_53), .B(n_151), .Y(n_150) );
AOI22xp33_ASAP7_75t_SL g196 ( .A1(n_55), .A2(n_59), .B1(n_139), .B2(n_143), .Y(n_196) );
CKINVDCx20_ASAP7_75t_R g518 ( .A(n_56), .Y(n_518) );
NAND2xp5_ASAP7_75t_SL g168 ( .A(n_57), .B(n_139), .Y(n_168) );
NAND2xp5_ASAP7_75t_SL g222 ( .A(n_58), .B(n_139), .Y(n_222) );
INVx1_ASAP7_75t_L g155 ( .A(n_60), .Y(n_155) );
NAND2xp5_ASAP7_75t_L g529 ( .A(n_61), .B(n_462), .Y(n_529) );
NAND2xp5_ASAP7_75t_L g492 ( .A(n_62), .B(n_493), .Y(n_492) );
A2O1A1Ixp33_ASAP7_75t_L g489 ( .A1(n_63), .A2(n_151), .B(n_183), .C(n_490), .Y(n_489) );
NAND2xp5_ASAP7_75t_L g188 ( .A(n_64), .B(n_139), .Y(n_188) );
INVx1_ASAP7_75t_L g134 ( .A(n_65), .Y(n_134) );
CKINVDCx20_ASAP7_75t_R g739 ( .A(n_66), .Y(n_739) );
NAND2xp5_ASAP7_75t_SL g503 ( .A(n_67), .B(n_145), .Y(n_503) );
AO32x2_ASAP7_75t_L g235 ( .A1(n_68), .A2(n_130), .A3(n_171), .B1(n_236), .B2(n_240), .Y(n_235) );
NAND2xp5_ASAP7_75t_L g455 ( .A(n_69), .B(n_146), .Y(n_455) );
INVx1_ASAP7_75t_L g166 ( .A(n_70), .Y(n_166) );
INVx1_ASAP7_75t_L g206 ( .A(n_71), .Y(n_206) );
CKINVDCx16_ASAP7_75t_R g547 ( .A(n_72), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g514 ( .A(n_73), .B(n_469), .Y(n_514) );
A2O1A1Ixp33_ASAP7_75t_L g524 ( .A1(n_74), .A2(n_452), .B(n_472), .C(n_525), .Y(n_524) );
NAND2xp5_ASAP7_75t_SL g207 ( .A(n_75), .B(n_143), .Y(n_207) );
CKINVDCx16_ASAP7_75t_R g488 ( .A(n_76), .Y(n_488) );
INVx1_ASAP7_75t_L g112 ( .A(n_77), .Y(n_112) );
CKINVDCx20_ASAP7_75t_R g116 ( .A(n_78), .Y(n_116) );
OAI22xp5_ASAP7_75t_SL g121 ( .A1(n_79), .A2(n_122), .B1(n_432), .B2(n_433), .Y(n_121) );
CKINVDCx20_ASAP7_75t_R g433 ( .A(n_79), .Y(n_433) );
NAND2xp5_ASAP7_75t_SL g515 ( .A(n_80), .B(n_468), .Y(n_515) );
NAND2xp5_ASAP7_75t_L g228 ( .A(n_82), .B(n_217), .Y(n_228) );
CKINVDCx20_ASAP7_75t_R g505 ( .A(n_83), .Y(n_505) );
NAND2xp5_ASAP7_75t_SL g210 ( .A(n_84), .B(n_143), .Y(n_210) );
INVx2_ASAP7_75t_L g132 ( .A(n_85), .Y(n_132) );
CKINVDCx20_ASAP7_75t_R g531 ( .A(n_86), .Y(n_531) );
NAND2xp5_ASAP7_75t_SL g456 ( .A(n_87), .B(n_170), .Y(n_456) );
NAND2xp5_ASAP7_75t_L g142 ( .A(n_88), .B(n_143), .Y(n_142) );
NAND3xp33_ASAP7_75t_SL g108 ( .A(n_89), .B(n_109), .C(n_110), .Y(n_108) );
OR2x2_ASAP7_75t_L g436 ( .A(n_89), .B(n_437), .Y(n_436) );
INVx2_ASAP7_75t_L g726 ( .A(n_89), .Y(n_726) );
OR2x2_ASAP7_75t_L g750 ( .A(n_89), .B(n_736), .Y(n_750) );
AOI22xp33_ASAP7_75t_L g195 ( .A1(n_91), .A2(n_101), .B1(n_143), .B2(n_144), .Y(n_195) );
NAND2xp5_ASAP7_75t_L g499 ( .A(n_92), .B(n_462), .Y(n_499) );
CKINVDCx20_ASAP7_75t_R g733 ( .A(n_93), .Y(n_733) );
INVx1_ASAP7_75t_L g502 ( .A(n_94), .Y(n_502) );
INVxp67_ASAP7_75t_L g491 ( .A(n_95), .Y(n_491) );
NAND2xp5_ASAP7_75t_L g164 ( .A(n_96), .B(n_143), .Y(n_164) );
NAND2xp5_ASAP7_75t_L g111 ( .A(n_97), .B(n_112), .Y(n_111) );
INVx1_ASAP7_75t_L g448 ( .A(n_98), .Y(n_448) );
INVx1_ASAP7_75t_L g526 ( .A(n_99), .Y(n_526) );
AND2x2_ASAP7_75t_L g474 ( .A(n_100), .B(n_173), .Y(n_474) );
INVx1_ASAP7_75t_L g103 ( .A(n_104), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_105), .Y(n_104) );
CKINVDCx20_ASAP7_75t_R g757 ( .A(n_105), .Y(n_757) );
CKINVDCx12_ASAP7_75t_R g105 ( .A(n_106), .Y(n_105) );
OR2x2_ASAP7_75t_L g106 ( .A(n_107), .B(n_108), .Y(n_106) );
AND2x2_ASAP7_75t_L g437 ( .A(n_109), .B(n_438), .Y(n_437) );
INVx1_ASAP7_75t_SL g110 ( .A(n_111), .Y(n_110) );
AO221x1_ASAP7_75t_L g113 ( .A1(n_114), .A2(n_737), .B1(n_740), .B2(n_751), .C(n_753), .Y(n_113) );
OAI222xp33_ASAP7_75t_SL g114 ( .A1(n_115), .A2(n_118), .B1(n_727), .B2(n_728), .C1(n_733), .C2(n_734), .Y(n_114) );
INVx1_ASAP7_75t_L g727 ( .A(n_115), .Y(n_727) );
INVxp67_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
OAI22xp5_ASAP7_75t_SL g119 ( .A1(n_120), .A2(n_434), .B1(n_439), .B2(n_723), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
OAI22xp5_ASAP7_75t_SL g729 ( .A1(n_121), .A2(n_730), .B1(n_731), .B2(n_732), .Y(n_729) );
INVx2_ASAP7_75t_L g432 ( .A(n_122), .Y(n_432) );
OAI22xp5_ASAP7_75t_L g742 ( .A1(n_122), .A2(n_432), .B1(n_743), .B2(n_744), .Y(n_742) );
NAND2x1p5_ASAP7_75t_L g122 ( .A(n_123), .B(n_356), .Y(n_122) );
AND2x2_ASAP7_75t_SL g123 ( .A(n_124), .B(n_314), .Y(n_123) );
NOR4xp25_ASAP7_75t_L g124 ( .A(n_125), .B(n_254), .C(n_290), .D(n_304), .Y(n_124) );
OAI221xp5_ASAP7_75t_SL g125 ( .A1(n_126), .A2(n_198), .B1(n_230), .B2(n_241), .C(n_245), .Y(n_125) );
NAND2xp5_ASAP7_75t_SL g388 ( .A(n_126), .B(n_389), .Y(n_388) );
OR2x2_ASAP7_75t_L g126 ( .A(n_127), .B(n_174), .Y(n_126) );
INVx1_ASAP7_75t_L g127 ( .A(n_128), .Y(n_127) );
AND2x2_ASAP7_75t_L g128 ( .A(n_129), .B(n_157), .Y(n_128) );
AND2x2_ASAP7_75t_L g251 ( .A(n_129), .B(n_158), .Y(n_251) );
INVx3_ASAP7_75t_L g259 ( .A(n_129), .Y(n_259) );
AND2x2_ASAP7_75t_L g313 ( .A(n_129), .B(n_177), .Y(n_313) );
NAND2xp5_ASAP7_75t_L g349 ( .A(n_129), .B(n_176), .Y(n_349) );
AND2x2_ASAP7_75t_L g407 ( .A(n_129), .B(n_269), .Y(n_407) );
OA21x2_ASAP7_75t_L g129 ( .A1(n_130), .A2(n_136), .B(n_156), .Y(n_129) );
INVx4_ASAP7_75t_L g197 ( .A(n_130), .Y(n_197) );
AOI21xp5_ASAP7_75t_L g478 ( .A1(n_130), .A2(n_479), .B(n_480), .Y(n_478) );
HB1xp67_ASAP7_75t_L g485 ( .A(n_130), .Y(n_485) );
BUFx6f_ASAP7_75t_L g130 ( .A(n_131), .Y(n_130) );
INVx1_ASAP7_75t_L g160 ( .A(n_131), .Y(n_160) );
AND2x2_ASAP7_75t_L g131 ( .A(n_132), .B(n_133), .Y(n_131) );
AND2x2_ASAP7_75t_SL g173 ( .A(n_132), .B(n_133), .Y(n_173) );
NAND2xp5_ASAP7_75t_L g133 ( .A(n_134), .B(n_135), .Y(n_133) );
OAI21xp5_ASAP7_75t_L g136 ( .A1(n_137), .A2(n_148), .B(n_154), .Y(n_136) );
AOI21xp5_ASAP7_75t_L g137 ( .A1(n_138), .A2(n_142), .B(n_145), .Y(n_137) );
INVx3_ASAP7_75t_L g205 ( .A(n_139), .Y(n_205) );
HB1xp67_ASAP7_75t_L g528 ( .A(n_139), .Y(n_528) );
BUFx6f_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
INVx1_ASAP7_75t_L g217 ( .A(n_140), .Y(n_217) );
BUFx3_ASAP7_75t_L g238 ( .A(n_140), .Y(n_238) );
AND2x6_ASAP7_75t_L g452 ( .A(n_140), .B(n_453), .Y(n_452) );
INVx2_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
INVx1_ASAP7_75t_L g144 ( .A(n_141), .Y(n_144) );
INVx1_ASAP7_75t_L g152 ( .A(n_141), .Y(n_152) );
INVx2_ASAP7_75t_L g181 ( .A(n_143), .Y(n_181) );
INVx3_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
INVx2_ASAP7_75t_L g153 ( .A(n_145), .Y(n_153) );
AOI21xp5_ASAP7_75t_L g162 ( .A1(n_145), .A2(n_163), .B(n_164), .Y(n_162) );
O2A1O1Ixp5_ASAP7_75t_SL g204 ( .A1(n_145), .A2(n_205), .B(n_206), .C(n_207), .Y(n_204) );
NOR2xp33_ASAP7_75t_L g490 ( .A(n_145), .B(n_491), .Y(n_490) );
INVx5_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
OAI22xp5_ASAP7_75t_SL g236 ( .A1(n_146), .A2(n_170), .B1(n_237), .B2(n_239), .Y(n_236) );
INVx3_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
BUFx6f_ASAP7_75t_L g170 ( .A(n_147), .Y(n_170) );
BUFx6f_ASAP7_75t_L g185 ( .A(n_147), .Y(n_185) );
INVx1_ASAP7_75t_L g225 ( .A(n_147), .Y(n_225) );
AND2x2_ASAP7_75t_L g450 ( .A(n_147), .B(n_152), .Y(n_450) );
INVx1_ASAP7_75t_L g453 ( .A(n_147), .Y(n_453) );
AOI21xp5_ASAP7_75t_L g148 ( .A1(n_149), .A2(n_150), .B(n_153), .Y(n_148) );
INVx2_ASAP7_75t_L g167 ( .A(n_151), .Y(n_167) );
INVx1_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
O2A1O1Ixp33_ASAP7_75t_L g186 ( .A1(n_153), .A2(n_167), .B(n_187), .C(n_188), .Y(n_186) );
OAI22xp5_ASAP7_75t_L g194 ( .A1(n_153), .A2(n_170), .B1(n_195), .B2(n_196), .Y(n_194) );
OAI22xp5_ASAP7_75t_L g215 ( .A1(n_153), .A2(n_170), .B1(n_216), .B2(n_218), .Y(n_215) );
BUFx3_ASAP7_75t_L g171 ( .A(n_154), .Y(n_171) );
OAI21xp5_ASAP7_75t_L g178 ( .A1(n_154), .A2(n_179), .B(n_186), .Y(n_178) );
OAI21xp5_ASAP7_75t_L g203 ( .A1(n_154), .A2(n_204), .B(n_208), .Y(n_203) );
OAI21xp5_ASAP7_75t_L g220 ( .A1(n_154), .A2(n_221), .B(n_226), .Y(n_220) );
NAND2x1p5_ASAP7_75t_L g449 ( .A(n_154), .B(n_450), .Y(n_449) );
AND2x4_ASAP7_75t_L g462 ( .A(n_154), .B(n_450), .Y(n_462) );
INVx4_ASAP7_75t_SL g473 ( .A(n_154), .Y(n_473) );
AND2x2_ASAP7_75t_L g242 ( .A(n_157), .B(n_243), .Y(n_242) );
AND2x2_ASAP7_75t_L g256 ( .A(n_157), .B(n_177), .Y(n_256) );
INVx2_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
NAND2xp5_ASAP7_75t_L g271 ( .A(n_158), .B(n_177), .Y(n_271) );
AND2x2_ASAP7_75t_L g283 ( .A(n_158), .B(n_259), .Y(n_283) );
OR2x2_ASAP7_75t_L g285 ( .A(n_158), .B(n_243), .Y(n_285) );
AND2x2_ASAP7_75t_L g320 ( .A(n_158), .B(n_243), .Y(n_320) );
HB1xp67_ASAP7_75t_L g365 ( .A(n_158), .Y(n_365) );
INVx1_ASAP7_75t_L g373 ( .A(n_158), .Y(n_373) );
OA21x2_ASAP7_75t_L g158 ( .A1(n_159), .A2(n_161), .B(n_172), .Y(n_158) );
OA21x2_ASAP7_75t_L g177 ( .A1(n_159), .A2(n_178), .B(n_189), .Y(n_177) );
INVx2_ASAP7_75t_L g159 ( .A(n_160), .Y(n_159) );
NOR2xp33_ASAP7_75t_L g457 ( .A(n_160), .B(n_458), .Y(n_457) );
OAI21xp5_ASAP7_75t_L g161 ( .A1(n_162), .A2(n_165), .B(n_171), .Y(n_161) );
O2A1O1Ixp5_ASAP7_75t_L g165 ( .A1(n_166), .A2(n_167), .B(n_168), .C(n_169), .Y(n_165) );
AOI21xp5_ASAP7_75t_L g513 ( .A1(n_167), .A2(n_514), .B(n_515), .Y(n_513) );
AOI21xp5_ASAP7_75t_L g226 ( .A1(n_169), .A2(n_227), .B(n_228), .Y(n_226) );
INVx2_ASAP7_75t_L g169 ( .A(n_170), .Y(n_169) );
INVx4_ASAP7_75t_L g551 ( .A(n_170), .Y(n_551) );
NAND3xp33_ASAP7_75t_L g193 ( .A(n_171), .B(n_194), .C(n_197), .Y(n_193) );
OA21x2_ASAP7_75t_L g202 ( .A1(n_173), .A2(n_203), .B(n_211), .Y(n_202) );
OA21x2_ASAP7_75t_L g219 ( .A1(n_173), .A2(n_220), .B(n_229), .Y(n_219) );
INVx2_ASAP7_75t_L g240 ( .A(n_173), .Y(n_240) );
AOI21xp5_ASAP7_75t_L g460 ( .A1(n_173), .A2(n_461), .B(n_463), .Y(n_460) );
AOI21xp5_ASAP7_75t_L g498 ( .A1(n_173), .A2(n_499), .B(n_500), .Y(n_498) );
INVx1_ASAP7_75t_L g519 ( .A(n_173), .Y(n_519) );
OAI221xp5_ASAP7_75t_L g290 ( .A1(n_174), .A2(n_291), .B1(n_295), .B2(n_299), .C(n_300), .Y(n_290) );
INVx1_ASAP7_75t_L g174 ( .A(n_175), .Y(n_174) );
AND2x2_ASAP7_75t_L g250 ( .A(n_175), .B(n_251), .Y(n_250) );
AND2x2_ASAP7_75t_L g175 ( .A(n_176), .B(n_190), .Y(n_175) );
INVx2_ASAP7_75t_L g249 ( .A(n_176), .Y(n_249) );
AND2x2_ASAP7_75t_L g302 ( .A(n_176), .B(n_303), .Y(n_302) );
AND2x2_ASAP7_75t_L g321 ( .A(n_176), .B(n_259), .Y(n_321) );
INVx2_ASAP7_75t_L g176 ( .A(n_177), .Y(n_176) );
AND2x2_ASAP7_75t_L g384 ( .A(n_177), .B(n_259), .Y(n_384) );
O2A1O1Ixp33_ASAP7_75t_L g179 ( .A1(n_180), .A2(n_181), .B(n_182), .C(n_183), .Y(n_179) );
AOI21xp5_ASAP7_75t_L g454 ( .A1(n_181), .A2(n_455), .B(n_456), .Y(n_454) );
AOI21xp5_ASAP7_75t_L g481 ( .A1(n_181), .A2(n_482), .B(n_483), .Y(n_481) );
O2A1O1Ixp33_ASAP7_75t_L g525 ( .A1(n_183), .A2(n_526), .B(n_527), .C(n_528), .Y(n_525) );
INVx1_ASAP7_75t_L g183 ( .A(n_184), .Y(n_183) );
AOI21xp5_ASAP7_75t_L g208 ( .A1(n_184), .A2(n_209), .B(n_210), .Y(n_208) );
INVx4_ASAP7_75t_L g184 ( .A(n_185), .Y(n_184) );
INVx2_ASAP7_75t_L g469 ( .A(n_185), .Y(n_469) );
AND2x2_ASAP7_75t_L g306 ( .A(n_190), .B(n_251), .Y(n_306) );
OAI322xp33_ASAP7_75t_L g374 ( .A1(n_190), .A2(n_330), .A3(n_375), .B1(n_377), .B2(n_380), .C1(n_382), .C2(n_386), .Y(n_374) );
INVx3_ASAP7_75t_L g190 ( .A(n_191), .Y(n_190) );
NOR2x1_ASAP7_75t_L g257 ( .A(n_191), .B(n_258), .Y(n_257) );
INVx2_ASAP7_75t_L g270 ( .A(n_191), .Y(n_270) );
AND2x2_ASAP7_75t_L g379 ( .A(n_191), .B(n_259), .Y(n_379) );
AND2x2_ASAP7_75t_L g411 ( .A(n_191), .B(n_283), .Y(n_411) );
OR2x2_ASAP7_75t_L g414 ( .A(n_191), .B(n_415), .Y(n_414) );
AND2x4_ASAP7_75t_L g191 ( .A(n_192), .B(n_193), .Y(n_191) );
INVx1_ASAP7_75t_L g244 ( .A(n_192), .Y(n_244) );
AO21x1_ASAP7_75t_L g243 ( .A1(n_194), .A2(n_197), .B(n_244), .Y(n_243) );
AO21x2_ASAP7_75t_L g446 ( .A1(n_197), .A2(n_447), .B(n_457), .Y(n_446) );
INVx3_ASAP7_75t_L g493 ( .A(n_197), .Y(n_493) );
NOR2xp33_ASAP7_75t_L g504 ( .A(n_197), .B(n_505), .Y(n_504) );
AO21x2_ASAP7_75t_L g522 ( .A1(n_197), .A2(n_523), .B(n_530), .Y(n_522) );
NOR2xp33_ASAP7_75t_L g530 ( .A(n_197), .B(n_531), .Y(n_530) );
INVx1_ASAP7_75t_L g198 ( .A(n_199), .Y(n_198) );
AND2x2_ASAP7_75t_L g199 ( .A(n_200), .B(n_212), .Y(n_199) );
INVx1_ASAP7_75t_L g427 ( .A(n_200), .Y(n_427) );
INVx1_ASAP7_75t_L g200 ( .A(n_201), .Y(n_200) );
OR2x2_ASAP7_75t_L g232 ( .A(n_201), .B(n_219), .Y(n_232) );
INVx2_ASAP7_75t_L g267 ( .A(n_201), .Y(n_267) );
INVx2_ASAP7_75t_L g201 ( .A(n_202), .Y(n_201) );
INVx2_ASAP7_75t_L g289 ( .A(n_202), .Y(n_289) );
HB1xp67_ASAP7_75t_L g297 ( .A(n_202), .Y(n_297) );
OR2x2_ASAP7_75t_L g421 ( .A(n_202), .B(n_422), .Y(n_421) );
AND2x2_ASAP7_75t_L g246 ( .A(n_212), .B(n_247), .Y(n_246) );
AND2x2_ASAP7_75t_L g286 ( .A(n_212), .B(n_287), .Y(n_286) );
AND2x2_ASAP7_75t_L g338 ( .A(n_212), .B(n_339), .Y(n_338) );
AND2x2_ASAP7_75t_L g212 ( .A(n_213), .B(n_219), .Y(n_212) );
AND2x2_ASAP7_75t_L g233 ( .A(n_213), .B(n_234), .Y(n_233) );
NOR2xp67_ASAP7_75t_L g293 ( .A(n_213), .B(n_294), .Y(n_293) );
AND2x2_ASAP7_75t_L g347 ( .A(n_213), .B(n_235), .Y(n_347) );
OR2x2_ASAP7_75t_L g355 ( .A(n_213), .B(n_289), .Y(n_355) );
INVx2_ASAP7_75t_L g213 ( .A(n_214), .Y(n_213) );
BUFx2_ASAP7_75t_L g264 ( .A(n_214), .Y(n_264) );
AND2x2_ASAP7_75t_L g274 ( .A(n_214), .B(n_275), .Y(n_274) );
AND2x2_ASAP7_75t_L g298 ( .A(n_214), .B(n_219), .Y(n_298) );
AND2x2_ASAP7_75t_L g362 ( .A(n_214), .B(n_235), .Y(n_362) );
NOR2xp33_ASAP7_75t_L g252 ( .A(n_219), .B(n_253), .Y(n_252) );
NAND2xp5_ASAP7_75t_L g266 ( .A(n_219), .B(n_267), .Y(n_266) );
INVx2_ASAP7_75t_L g275 ( .A(n_219), .Y(n_275) );
INVx1_ASAP7_75t_L g280 ( .A(n_219), .Y(n_280) );
AND2x2_ASAP7_75t_L g292 ( .A(n_219), .B(n_293), .Y(n_292) );
HB1xp67_ASAP7_75t_L g370 ( .A(n_219), .Y(n_370) );
INVx1_ASAP7_75t_L g422 ( .A(n_219), .Y(n_422) );
AOI21xp5_ASAP7_75t_L g221 ( .A1(n_222), .A2(n_223), .B(n_224), .Y(n_221) );
INVx1_ASAP7_75t_L g224 ( .A(n_225), .Y(n_224) );
NAND2xp5_ASAP7_75t_L g230 ( .A(n_231), .B(n_233), .Y(n_230) );
AND2x2_ASAP7_75t_L g399 ( .A(n_231), .B(n_308), .Y(n_399) );
INVx2_ASAP7_75t_SL g231 ( .A(n_232), .Y(n_231) );
AND2x2_ASAP7_75t_L g326 ( .A(n_233), .B(n_327), .Y(n_326) );
AND2x2_ASAP7_75t_L g425 ( .A(n_233), .B(n_360), .Y(n_425) );
INVx1_ASAP7_75t_L g247 ( .A(n_234), .Y(n_247) );
AND2x2_ASAP7_75t_L g273 ( .A(n_234), .B(n_267), .Y(n_273) );
BUFx2_ASAP7_75t_L g332 ( .A(n_234), .Y(n_332) );
INVx1_ASAP7_75t_L g234 ( .A(n_235), .Y(n_234) );
BUFx6f_ASAP7_75t_L g253 ( .A(n_235), .Y(n_253) );
INVx1_ASAP7_75t_L g263 ( .A(n_235), .Y(n_263) );
HB1xp67_ASAP7_75t_L g471 ( .A(n_238), .Y(n_471) );
INVx2_ASAP7_75t_L g552 ( .A(n_238), .Y(n_552) );
INVx1_ASAP7_75t_L g516 ( .A(n_240), .Y(n_516) );
NOR2xp67_ASAP7_75t_L g401 ( .A(n_241), .B(n_248), .Y(n_401) );
INVx2_ASAP7_75t_L g241 ( .A(n_242), .Y(n_241) );
AOI32xp33_ASAP7_75t_L g245 ( .A1(n_242), .A2(n_246), .A3(n_248), .B1(n_250), .B2(n_252), .Y(n_245) );
AND2x2_ASAP7_75t_L g385 ( .A(n_242), .B(n_258), .Y(n_385) );
AND2x2_ASAP7_75t_L g423 ( .A(n_242), .B(n_321), .Y(n_423) );
INVx1_ASAP7_75t_L g303 ( .A(n_243), .Y(n_303) );
NAND2xp5_ASAP7_75t_L g417 ( .A(n_247), .B(n_309), .Y(n_417) );
NAND2xp5_ASAP7_75t_L g282 ( .A(n_248), .B(n_283), .Y(n_282) );
NAND2xp5_ASAP7_75t_L g299 ( .A(n_248), .B(n_251), .Y(n_299) );
NAND2xp5_ASAP7_75t_SL g402 ( .A(n_248), .B(n_320), .Y(n_402) );
OR2x2_ASAP7_75t_L g416 ( .A(n_248), .B(n_285), .Y(n_416) );
INVx3_ASAP7_75t_L g248 ( .A(n_249), .Y(n_248) );
AND2x2_ASAP7_75t_L g343 ( .A(n_249), .B(n_251), .Y(n_343) );
OR2x2_ASAP7_75t_L g352 ( .A(n_249), .B(n_339), .Y(n_352) );
NAND2xp5_ASAP7_75t_L g324 ( .A(n_251), .B(n_302), .Y(n_324) );
INVx2_ASAP7_75t_L g339 ( .A(n_253), .Y(n_339) );
OR2x2_ASAP7_75t_L g354 ( .A(n_253), .B(n_355), .Y(n_354) );
AND2x2_ASAP7_75t_L g369 ( .A(n_253), .B(n_370), .Y(n_369) );
A2O1A1Ixp33_ASAP7_75t_L g426 ( .A1(n_253), .A2(n_346), .B(n_427), .C(n_428), .Y(n_426) );
OAI321xp33_ASAP7_75t_L g254 ( .A1(n_255), .A2(n_260), .A3(n_265), .B1(n_268), .B2(n_272), .C(n_276), .Y(n_254) );
INVx1_ASAP7_75t_L g367 ( .A(n_255), .Y(n_367) );
NAND2x1p5_ASAP7_75t_L g255 ( .A(n_256), .B(n_257), .Y(n_255) );
AND2x2_ASAP7_75t_L g378 ( .A(n_256), .B(n_379), .Y(n_378) );
INVx1_ASAP7_75t_L g330 ( .A(n_258), .Y(n_330) );
INVx2_ASAP7_75t_L g258 ( .A(n_259), .Y(n_258) );
NAND2xp5_ASAP7_75t_L g390 ( .A(n_259), .B(n_373), .Y(n_390) );
OAI221xp5_ASAP7_75t_L g397 ( .A1(n_260), .A2(n_398), .B1(n_400), .B2(n_402), .C(n_403), .Y(n_397) );
INVx1_ASAP7_75t_L g260 ( .A(n_261), .Y(n_260) );
AND2x2_ASAP7_75t_L g261 ( .A(n_262), .B(n_264), .Y(n_261) );
AND2x2_ASAP7_75t_L g335 ( .A(n_262), .B(n_309), .Y(n_335) );
HB1xp67_ASAP7_75t_L g262 ( .A(n_263), .Y(n_262) );
NAND2xp5_ASAP7_75t_L g288 ( .A(n_263), .B(n_289), .Y(n_288) );
INVx2_ASAP7_75t_L g308 ( .A(n_264), .Y(n_308) );
A2O1A1Ixp33_ASAP7_75t_L g350 ( .A1(n_265), .A2(n_306), .B(n_351), .C(n_353), .Y(n_350) );
INVx1_ASAP7_75t_L g265 ( .A(n_266), .Y(n_265) );
AND2x2_ASAP7_75t_L g317 ( .A(n_267), .B(n_274), .Y(n_317) );
BUFx2_ASAP7_75t_L g327 ( .A(n_267), .Y(n_327) );
INVx1_ASAP7_75t_L g342 ( .A(n_267), .Y(n_342) );
INVx1_ASAP7_75t_L g268 ( .A(n_269), .Y(n_268) );
NOR2xp33_ASAP7_75t_L g269 ( .A(n_270), .B(n_271), .Y(n_269) );
OR2x2_ASAP7_75t_L g348 ( .A(n_270), .B(n_349), .Y(n_348) );
INVx1_ASAP7_75t_L g431 ( .A(n_270), .Y(n_431) );
INVx1_ASAP7_75t_L g424 ( .A(n_271), .Y(n_424) );
NAND2xp5_ASAP7_75t_L g272 ( .A(n_273), .B(n_274), .Y(n_272) );
AND2x2_ASAP7_75t_L g277 ( .A(n_273), .B(n_278), .Y(n_277) );
AND2x2_ASAP7_75t_L g381 ( .A(n_273), .B(n_298), .Y(n_381) );
INVx1_ASAP7_75t_L g310 ( .A(n_274), .Y(n_310) );
AOI22xp5_ASAP7_75t_L g276 ( .A1(n_277), .A2(n_281), .B1(n_284), .B2(n_286), .Y(n_276) );
NAND2xp5_ASAP7_75t_L g393 ( .A(n_278), .B(n_394), .Y(n_393) );
INVxp67_ASAP7_75t_L g278 ( .A(n_279), .Y(n_278) );
AND2x4_ASAP7_75t_L g346 ( .A(n_279), .B(n_347), .Y(n_346) );
BUFx3_ASAP7_75t_L g279 ( .A(n_280), .Y(n_279) );
AND2x2_ASAP7_75t_SL g309 ( .A(n_280), .B(n_289), .Y(n_309) );
INVx1_ASAP7_75t_L g281 ( .A(n_282), .Y(n_281) );
AND2x2_ASAP7_75t_L g301 ( .A(n_283), .B(n_302), .Y(n_301) );
INVx1_ASAP7_75t_SL g284 ( .A(n_285), .Y(n_284) );
OR2x2_ASAP7_75t_L g311 ( .A(n_285), .B(n_312), .Y(n_311) );
INVx1_ASAP7_75t_SL g287 ( .A(n_288), .Y(n_287) );
OAI221xp5_ASAP7_75t_L g405 ( .A1(n_288), .A2(n_406), .B1(n_408), .B2(n_409), .C(n_410), .Y(n_405) );
INVx1_ASAP7_75t_L g294 ( .A(n_289), .Y(n_294) );
HB1xp67_ASAP7_75t_L g360 ( .A(n_289), .Y(n_360) );
INVx1_ASAP7_75t_SL g291 ( .A(n_292), .Y(n_291) );
NAND2xp5_ASAP7_75t_L g410 ( .A(n_292), .B(n_411), .Y(n_410) );
OAI21xp5_ASAP7_75t_L g300 ( .A1(n_293), .A2(n_298), .B(n_301), .Y(n_300) );
INVx1_ASAP7_75t_L g295 ( .A(n_296), .Y(n_295) );
NAND2xp5_ASAP7_75t_L g403 ( .A(n_296), .B(n_306), .Y(n_403) );
AND2x2_ASAP7_75t_L g296 ( .A(n_297), .B(n_298), .Y(n_296) );
INVx1_ASAP7_75t_L g372 ( .A(n_297), .Y(n_372) );
AND2x2_ASAP7_75t_L g331 ( .A(n_298), .B(n_332), .Y(n_331) );
INVx2_ASAP7_75t_L g420 ( .A(n_298), .Y(n_420) );
INVx1_ASAP7_75t_L g336 ( .A(n_301), .Y(n_336) );
INVx1_ASAP7_75t_L g391 ( .A(n_302), .Y(n_391) );
OAI22xp5_ASAP7_75t_L g304 ( .A1(n_305), .A2(n_307), .B1(n_310), .B2(n_311), .Y(n_304) );
INVx1_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
NAND2xp5_ASAP7_75t_L g307 ( .A(n_308), .B(n_309), .Y(n_307) );
NAND2xp5_ASAP7_75t_L g341 ( .A(n_308), .B(n_342), .Y(n_341) );
INVx2_ASAP7_75t_L g376 ( .A(n_309), .Y(n_376) );
NAND2xp5_ASAP7_75t_SL g413 ( .A(n_309), .B(n_347), .Y(n_413) );
OR2x2_ASAP7_75t_L g386 ( .A(n_310), .B(n_339), .Y(n_386) );
INVx1_ASAP7_75t_L g325 ( .A(n_311), .Y(n_325) );
INVx1_ASAP7_75t_SL g312 ( .A(n_313), .Y(n_312) );
NAND2xp5_ASAP7_75t_L g363 ( .A(n_313), .B(n_364), .Y(n_363) );
NOR3xp33_ASAP7_75t_L g314 ( .A(n_315), .B(n_333), .C(n_344), .Y(n_314) );
OAI211xp5_ASAP7_75t_L g315 ( .A1(n_316), .A2(n_318), .B(n_322), .C(n_328), .Y(n_315) );
INVxp67_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
AOI221xp5_ASAP7_75t_L g387 ( .A1(n_317), .A2(n_388), .B1(n_392), .B2(n_395), .C(n_397), .Y(n_387) );
INVx1_ASAP7_75t_SL g318 ( .A(n_319), .Y(n_318) );
AND2x2_ASAP7_75t_L g319 ( .A(n_320), .B(n_321), .Y(n_319) );
AND2x2_ASAP7_75t_L g329 ( .A(n_320), .B(n_330), .Y(n_329) );
AND2x2_ASAP7_75t_L g383 ( .A(n_320), .B(n_384), .Y(n_383) );
OAI211xp5_ASAP7_75t_L g368 ( .A1(n_321), .A2(n_369), .B(n_371), .C(n_373), .Y(n_368) );
INVx2_ASAP7_75t_L g415 ( .A(n_321), .Y(n_415) );
OAI21xp5_ASAP7_75t_SL g322 ( .A1(n_323), .A2(n_325), .B(n_326), .Y(n_322) );
INVx1_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
AND2x2_ASAP7_75t_L g394 ( .A(n_327), .B(n_347), .Y(n_394) );
NAND2xp5_ASAP7_75t_L g328 ( .A(n_329), .B(n_331), .Y(n_328) );
OAI21xp5_ASAP7_75t_SL g333 ( .A1(n_334), .A2(n_336), .B(n_337), .Y(n_333) );
INVxp67_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
OAI21xp5_ASAP7_75t_SL g337 ( .A1(n_338), .A2(n_340), .B(n_343), .Y(n_337) );
NAND2xp5_ASAP7_75t_L g366 ( .A(n_338), .B(n_367), .Y(n_366) );
INVxp67_ASAP7_75t_L g340 ( .A(n_341), .Y(n_340) );
NAND2xp5_ASAP7_75t_L g429 ( .A(n_343), .B(n_430), .Y(n_429) );
OAI21xp33_ASAP7_75t_L g344 ( .A1(n_345), .A2(n_348), .B(n_350), .Y(n_344) );
INVx1_ASAP7_75t_SL g345 ( .A(n_346), .Y(n_345) );
AND2x2_ASAP7_75t_L g371 ( .A(n_347), .B(n_372), .Y(n_371) );
INVx1_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
INVx1_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
AND4x1_ASAP7_75t_L g356 ( .A(n_357), .B(n_387), .C(n_404), .D(n_426), .Y(n_356) );
NOR2xp33_ASAP7_75t_L g357 ( .A(n_358), .B(n_374), .Y(n_357) );
OAI211xp5_ASAP7_75t_SL g358 ( .A1(n_359), .A2(n_363), .B(n_366), .C(n_368), .Y(n_358) );
OR2x2_ASAP7_75t_L g359 ( .A(n_360), .B(n_361), .Y(n_359) );
INVx1_ASAP7_75t_SL g361 ( .A(n_362), .Y(n_361) );
NAND2xp5_ASAP7_75t_L g375 ( .A(n_362), .B(n_376), .Y(n_375) );
INVx1_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
NOR2xp33_ASAP7_75t_L g395 ( .A(n_373), .B(n_396), .Y(n_395) );
INVx1_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
INVx1_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
NOR2xp33_ASAP7_75t_L g382 ( .A(n_383), .B(n_385), .Y(n_382) );
INVx1_ASAP7_75t_L g408 ( .A(n_383), .Y(n_408) );
INVx2_ASAP7_75t_SL g396 ( .A(n_384), .Y(n_396) );
OR2x2_ASAP7_75t_L g389 ( .A(n_390), .B(n_391), .Y(n_389) );
INVx1_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
INVx1_ASAP7_75t_L g409 ( .A(n_394), .Y(n_409) );
INVx1_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
INVx1_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
NOR2xp33_ASAP7_75t_SL g404 ( .A(n_405), .B(n_412), .Y(n_404) );
INVx1_ASAP7_75t_SL g406 ( .A(n_407), .Y(n_406) );
OAI221xp5_ASAP7_75t_SL g412 ( .A1(n_413), .A2(n_414), .B1(n_416), .B2(n_417), .C(n_418), .Y(n_412) );
AOI22xp5_ASAP7_75t_L g418 ( .A1(n_419), .A2(n_423), .B1(n_424), .B2(n_425), .Y(n_418) );
NAND2xp5_ASAP7_75t_SL g419 ( .A(n_420), .B(n_421), .Y(n_419) );
INVx1_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
INVx1_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
INVx2_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
INVx2_ASAP7_75t_L g730 ( .A(n_435), .Y(n_730) );
INVx1_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
OR2x2_ASAP7_75t_L g725 ( .A(n_437), .B(n_726), .Y(n_725) );
INVx2_ASAP7_75t_L g736 ( .A(n_437), .Y(n_736) );
INVx2_ASAP7_75t_L g731 ( .A(n_439), .Y(n_731) );
OR3x1_ASAP7_75t_L g439 ( .A(n_440), .B(n_621), .C(n_686), .Y(n_439) );
NAND4xp25_ASAP7_75t_SL g440 ( .A(n_441), .B(n_562), .C(n_588), .D(n_611), .Y(n_440) );
AOI221xp5_ASAP7_75t_L g441 ( .A1(n_442), .A2(n_494), .B1(n_532), .B2(n_539), .C(n_554), .Y(n_441) );
CKINVDCx14_ASAP7_75t_R g442 ( .A(n_443), .Y(n_442) );
OAI22xp5_ASAP7_75t_L g709 ( .A1(n_443), .A2(n_555), .B1(n_579), .B2(n_710), .Y(n_709) );
OR2x2_ASAP7_75t_L g443 ( .A(n_444), .B(n_475), .Y(n_443) );
INVx1_ASAP7_75t_SL g615 ( .A(n_444), .Y(n_615) );
OR2x2_ASAP7_75t_L g444 ( .A(n_445), .B(n_459), .Y(n_444) );
OR2x2_ASAP7_75t_L g537 ( .A(n_445), .B(n_538), .Y(n_537) );
AND2x2_ASAP7_75t_L g557 ( .A(n_445), .B(n_476), .Y(n_557) );
NAND2xp5_ASAP7_75t_L g570 ( .A(n_445), .B(n_484), .Y(n_570) );
AND2x2_ASAP7_75t_L g587 ( .A(n_445), .B(n_459), .Y(n_587) );
NAND2xp5_ASAP7_75t_L g609 ( .A(n_445), .B(n_535), .Y(n_609) );
NAND2xp5_ASAP7_75t_L g698 ( .A(n_445), .B(n_586), .Y(n_698) );
NOR2xp33_ASAP7_75t_L g708 ( .A(n_445), .B(n_475), .Y(n_708) );
AOI211xp5_ASAP7_75t_SL g719 ( .A1(n_445), .A2(n_625), .B(n_720), .C(n_721), .Y(n_719) );
INVx5_ASAP7_75t_SL g445 ( .A(n_446), .Y(n_445) );
NAND2xp5_ASAP7_75t_SL g591 ( .A(n_446), .B(n_476), .Y(n_591) );
AND2x2_ASAP7_75t_L g594 ( .A(n_446), .B(n_477), .Y(n_594) );
OR2x2_ASAP7_75t_L g639 ( .A(n_446), .B(n_476), .Y(n_639) );
NAND2xp5_ASAP7_75t_L g648 ( .A(n_446), .B(n_484), .Y(n_648) );
OAI21xp5_ASAP7_75t_L g447 ( .A1(n_448), .A2(n_449), .B(n_451), .Y(n_447) );
INVx5_ASAP7_75t_L g465 ( .A(n_452), .Y(n_465) );
INVx5_ASAP7_75t_SL g538 ( .A(n_459), .Y(n_538) );
AND2x2_ASAP7_75t_L g556 ( .A(n_459), .B(n_557), .Y(n_556) );
NOR2xp33_ASAP7_75t_L g638 ( .A(n_459), .B(n_639), .Y(n_638) );
AND2x2_ASAP7_75t_L g642 ( .A(n_459), .B(n_643), .Y(n_642) );
AND2x2_ASAP7_75t_L g674 ( .A(n_459), .B(n_484), .Y(n_674) );
OR2x2_ASAP7_75t_L g680 ( .A(n_459), .B(n_570), .Y(n_680) );
NAND2xp5_ASAP7_75t_L g689 ( .A(n_459), .B(n_630), .Y(n_689) );
OR2x6_ASAP7_75t_L g459 ( .A(n_460), .B(n_474), .Y(n_459) );
BUFx2_ASAP7_75t_L g511 ( .A(n_462), .Y(n_511) );
INVx2_ASAP7_75t_L g464 ( .A(n_465), .Y(n_464) );
O2A1O1Ixp33_ASAP7_75t_L g487 ( .A1(n_465), .A2(n_473), .B(n_488), .C(n_489), .Y(n_487) );
O2A1O1Ixp33_ASAP7_75t_SL g546 ( .A1(n_465), .A2(n_473), .B(n_547), .C(n_548), .Y(n_546) );
O2A1O1Ixp33_ASAP7_75t_L g466 ( .A1(n_467), .A2(n_468), .B(n_470), .C(n_471), .Y(n_466) );
O2A1O1Ixp33_ASAP7_75t_L g501 ( .A1(n_468), .A2(n_471), .B(n_502), .C(n_503), .Y(n_501) );
INVx2_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
INVx1_ASAP7_75t_L g472 ( .A(n_473), .Y(n_472) );
NAND2xp5_ASAP7_75t_L g475 ( .A(n_476), .B(n_484), .Y(n_475) );
AND2x2_ASAP7_75t_L g571 ( .A(n_476), .B(n_538), .Y(n_571) );
INVx1_ASAP7_75t_SL g584 ( .A(n_476), .Y(n_584) );
OR2x2_ASAP7_75t_L g619 ( .A(n_476), .B(n_620), .Y(n_619) );
OR2x2_ASAP7_75t_L g625 ( .A(n_476), .B(n_484), .Y(n_625) );
AND2x2_ASAP7_75t_L g683 ( .A(n_476), .B(n_535), .Y(n_683) );
INVx2_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
NAND2xp5_ASAP7_75t_L g610 ( .A(n_477), .B(n_538), .Y(n_610) );
INVx3_ASAP7_75t_L g535 ( .A(n_484), .Y(n_535) );
OR2x2_ASAP7_75t_L g576 ( .A(n_484), .B(n_538), .Y(n_576) );
AND2x2_ASAP7_75t_L g586 ( .A(n_484), .B(n_584), .Y(n_586) );
HB1xp67_ASAP7_75t_L g634 ( .A(n_484), .Y(n_634) );
AND2x2_ASAP7_75t_L g643 ( .A(n_484), .B(n_557), .Y(n_643) );
OA21x2_ASAP7_75t_L g484 ( .A1(n_485), .A2(n_486), .B(n_492), .Y(n_484) );
OA21x2_ASAP7_75t_L g544 ( .A1(n_493), .A2(n_545), .B(n_553), .Y(n_544) );
AOI221xp5_ASAP7_75t_L g659 ( .A1(n_494), .A2(n_660), .B1(n_662), .B2(n_664), .C(n_667), .Y(n_659) );
INVx2_ASAP7_75t_L g494 ( .A(n_495), .Y(n_494) );
OR2x2_ASAP7_75t_L g495 ( .A(n_496), .B(n_506), .Y(n_495) );
AND2x2_ASAP7_75t_L g633 ( .A(n_496), .B(n_614), .Y(n_633) );
NAND2xp5_ASAP7_75t_L g696 ( .A(n_496), .B(n_692), .Y(n_696) );
OR2x2_ASAP7_75t_L g717 ( .A(n_496), .B(n_718), .Y(n_717) );
NAND2xp5_ASAP7_75t_L g721 ( .A(n_496), .B(n_722), .Y(n_721) );
BUFx2_ASAP7_75t_L g496 ( .A(n_497), .Y(n_496) );
INVx5_ASAP7_75t_L g564 ( .A(n_497), .Y(n_564) );
AND2x2_ASAP7_75t_L g641 ( .A(n_497), .B(n_508), .Y(n_641) );
AND2x2_ASAP7_75t_L g702 ( .A(n_497), .B(n_581), .Y(n_702) );
AND2x2_ASAP7_75t_L g715 ( .A(n_497), .B(n_535), .Y(n_715) );
OR2x6_ASAP7_75t_L g497 ( .A(n_498), .B(n_504), .Y(n_497) );
NAND2xp5_ASAP7_75t_L g506 ( .A(n_507), .B(n_520), .Y(n_506) );
AND2x4_ASAP7_75t_L g542 ( .A(n_507), .B(n_543), .Y(n_542) );
AND2x2_ASAP7_75t_L g560 ( .A(n_507), .B(n_561), .Y(n_560) );
INVx2_ASAP7_75t_L g567 ( .A(n_507), .Y(n_567) );
AND2x2_ASAP7_75t_L g636 ( .A(n_507), .B(n_614), .Y(n_636) );
AND2x2_ASAP7_75t_L g646 ( .A(n_507), .B(n_564), .Y(n_646) );
HB1xp67_ASAP7_75t_L g654 ( .A(n_507), .Y(n_654) );
AND2x2_ASAP7_75t_L g666 ( .A(n_507), .B(n_544), .Y(n_666) );
NOR2xp33_ASAP7_75t_L g670 ( .A(n_507), .B(n_598), .Y(n_670) );
AND2x2_ASAP7_75t_L g707 ( .A(n_507), .B(n_702), .Y(n_707) );
NAND2xp5_ASAP7_75t_L g718 ( .A(n_507), .B(n_581), .Y(n_718) );
OR2x2_ASAP7_75t_L g720 ( .A(n_507), .B(n_656), .Y(n_720) );
INVx5_ASAP7_75t_L g507 ( .A(n_508), .Y(n_507) );
AND2x2_ASAP7_75t_L g606 ( .A(n_508), .B(n_607), .Y(n_606) );
AND2x2_ASAP7_75t_L g616 ( .A(n_508), .B(n_561), .Y(n_616) );
AND2x2_ASAP7_75t_L g628 ( .A(n_508), .B(n_544), .Y(n_628) );
HB1xp67_ASAP7_75t_L g658 ( .A(n_508), .Y(n_658) );
AND2x4_ASAP7_75t_L g692 ( .A(n_508), .B(n_543), .Y(n_692) );
OR2x6_ASAP7_75t_L g508 ( .A(n_509), .B(n_517), .Y(n_508) );
AOI21xp5_ASAP7_75t_SL g509 ( .A1(n_510), .A2(n_512), .B(n_516), .Y(n_509) );
NOR2xp33_ASAP7_75t_L g517 ( .A(n_518), .B(n_519), .Y(n_517) );
BUFx2_ASAP7_75t_L g541 ( .A(n_520), .Y(n_541) );
HB1xp67_ASAP7_75t_L g520 ( .A(n_521), .Y(n_520) );
INVx2_ASAP7_75t_L g581 ( .A(n_521), .Y(n_581) );
AND2x2_ASAP7_75t_L g614 ( .A(n_521), .B(n_544), .Y(n_614) );
INVx2_ASAP7_75t_L g521 ( .A(n_522), .Y(n_521) );
AND2x2_ASAP7_75t_L g561 ( .A(n_522), .B(n_544), .Y(n_561) );
BUFx2_ASAP7_75t_L g607 ( .A(n_522), .Y(n_607) );
NAND2xp5_ASAP7_75t_L g523 ( .A(n_524), .B(n_529), .Y(n_523) );
INVx1_ASAP7_75t_L g532 ( .A(n_533), .Y(n_532) );
NAND2xp5_ASAP7_75t_L g533 ( .A(n_534), .B(n_536), .Y(n_533) );
NAND2xp5_ASAP7_75t_L g694 ( .A(n_534), .B(n_615), .Y(n_694) );
INVx1_ASAP7_75t_L g534 ( .A(n_535), .Y(n_534) );
NAND2xp5_ASAP7_75t_L g558 ( .A(n_535), .B(n_557), .Y(n_558) );
NAND2xp5_ASAP7_75t_L g596 ( .A(n_535), .B(n_538), .Y(n_596) );
AND2x2_ASAP7_75t_L g651 ( .A(n_535), .B(n_587), .Y(n_651) );
AOI221xp5_ASAP7_75t_SL g588 ( .A1(n_536), .A2(n_589), .B1(n_597), .B2(n_599), .C(n_603), .Y(n_588) );
INVx2_ASAP7_75t_L g536 ( .A(n_537), .Y(n_536) );
OR2x2_ASAP7_75t_L g583 ( .A(n_537), .B(n_584), .Y(n_583) );
OR2x2_ASAP7_75t_L g624 ( .A(n_537), .B(n_625), .Y(n_624) );
OAI321xp33_ASAP7_75t_L g631 ( .A1(n_537), .A2(n_590), .A3(n_632), .B1(n_634), .B2(n_635), .C(n_637), .Y(n_631) );
NAND2xp5_ASAP7_75t_L g682 ( .A(n_538), .B(n_683), .Y(n_682) );
INVx1_ASAP7_75t_L g539 ( .A(n_540), .Y(n_539) );
NAND2xp5_ASAP7_75t_L g540 ( .A(n_541), .B(n_542), .Y(n_540) );
NAND2xp5_ASAP7_75t_L g710 ( .A(n_541), .B(n_692), .Y(n_710) );
AND2x2_ASAP7_75t_L g597 ( .A(n_542), .B(n_598), .Y(n_597) );
NAND2xp5_ASAP7_75t_L g600 ( .A(n_542), .B(n_601), .Y(n_600) );
HB1xp67_ASAP7_75t_L g573 ( .A(n_543), .Y(n_573) );
AND2x2_ASAP7_75t_L g580 ( .A(n_543), .B(n_581), .Y(n_580) );
NAND2xp5_ASAP7_75t_L g685 ( .A(n_543), .B(n_655), .Y(n_685) );
INVx1_ASAP7_75t_L g722 ( .A(n_543), .Y(n_722) );
INVx2_ASAP7_75t_L g543 ( .A(n_544), .Y(n_543) );
NOR2xp33_ASAP7_75t_L g549 ( .A(n_550), .B(n_551), .Y(n_549) );
AOI21xp5_ASAP7_75t_L g554 ( .A1(n_555), .A2(n_558), .B(n_559), .Y(n_554) );
INVx1_ASAP7_75t_SL g555 ( .A(n_556), .Y(n_555) );
A2O1A1Ixp33_ASAP7_75t_L g714 ( .A1(n_556), .A2(n_666), .B(n_715), .C(n_716), .Y(n_714) );
NAND2xp5_ASAP7_75t_L g574 ( .A(n_557), .B(n_575), .Y(n_574) );
NAND2xp5_ASAP7_75t_L g661 ( .A(n_557), .B(n_595), .Y(n_661) );
INVx1_ASAP7_75t_SL g559 ( .A(n_560), .Y(n_559) );
INVx1_ASAP7_75t_L g604 ( .A(n_561), .Y(n_604) );
NAND2xp5_ASAP7_75t_L g618 ( .A(n_561), .B(n_564), .Y(n_618) );
NOR2xp33_ASAP7_75t_L g627 ( .A(n_561), .B(n_628), .Y(n_627) );
NAND2xp5_ASAP7_75t_L g645 ( .A(n_561), .B(n_646), .Y(n_645) );
AOI22xp33_ASAP7_75t_L g562 ( .A1(n_563), .A2(n_565), .B1(n_577), .B2(n_582), .Y(n_562) );
HB1xp67_ASAP7_75t_L g563 ( .A(n_564), .Y(n_563) );
OR2x2_ASAP7_75t_L g578 ( .A(n_564), .B(n_579), .Y(n_578) );
AND2x2_ASAP7_75t_L g601 ( .A(n_564), .B(n_602), .Y(n_601) );
AND2x2_ASAP7_75t_L g613 ( .A(n_564), .B(n_614), .Y(n_613) );
NAND2xp5_ASAP7_75t_L g649 ( .A(n_564), .B(n_607), .Y(n_649) );
OR2x2_ASAP7_75t_L g656 ( .A(n_564), .B(n_581), .Y(n_656) );
NAND2xp5_ASAP7_75t_L g665 ( .A(n_564), .B(n_666), .Y(n_665) );
AND2x2_ASAP7_75t_L g706 ( .A(n_564), .B(n_692), .Y(n_706) );
OAI22xp33_ASAP7_75t_L g565 ( .A1(n_566), .A2(n_568), .B1(n_572), .B2(n_574), .Y(n_565) );
INVx1_ASAP7_75t_L g566 ( .A(n_567), .Y(n_566) );
AND2x2_ASAP7_75t_L g612 ( .A(n_567), .B(n_613), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g568 ( .A(n_569), .B(n_571), .Y(n_568) );
INVx1_ASAP7_75t_SL g569 ( .A(n_570), .Y(n_569) );
OAI22xp33_ASAP7_75t_L g652 ( .A1(n_570), .A2(n_585), .B1(n_653), .B2(n_657), .Y(n_652) );
INVx1_ASAP7_75t_L g700 ( .A(n_571), .Y(n_700) );
INVx1_ASAP7_75t_L g572 ( .A(n_573), .Y(n_572) );
AOI221xp5_ASAP7_75t_L g611 ( .A1(n_575), .A2(n_612), .B1(n_615), .B2(n_616), .C(n_617), .Y(n_611) );
INVx1_ASAP7_75t_L g575 ( .A(n_576), .Y(n_575) );
OR2x2_ASAP7_75t_L g590 ( .A(n_576), .B(n_591), .Y(n_590) );
INVx1_ASAP7_75t_L g577 ( .A(n_578), .Y(n_577) );
INVx1_ASAP7_75t_L g579 ( .A(n_580), .Y(n_579) );
NAND2xp5_ASAP7_75t_L g678 ( .A(n_580), .B(n_646), .Y(n_678) );
HB1xp67_ASAP7_75t_L g598 ( .A(n_581), .Y(n_598) );
INVx1_ASAP7_75t_L g602 ( .A(n_581), .Y(n_602) );
NAND2xp33_ASAP7_75t_L g582 ( .A(n_583), .B(n_585), .Y(n_582) );
NAND2xp5_ASAP7_75t_L g585 ( .A(n_586), .B(n_587), .Y(n_585) );
INVx1_ASAP7_75t_L g620 ( .A(n_587), .Y(n_620) );
AND2x2_ASAP7_75t_L g629 ( .A(n_587), .B(n_630), .Y(n_629) );
NAND2xp33_ASAP7_75t_L g589 ( .A(n_590), .B(n_592), .Y(n_589) );
INVx2_ASAP7_75t_SL g592 ( .A(n_593), .Y(n_592) );
AND2x4_ASAP7_75t_L g593 ( .A(n_594), .B(n_595), .Y(n_593) );
AND2x2_ASAP7_75t_L g673 ( .A(n_594), .B(n_674), .Y(n_673) );
INVx2_ASAP7_75t_L g595 ( .A(n_596), .Y(n_595) );
AOI221xp5_ASAP7_75t_L g622 ( .A1(n_597), .A2(n_623), .B1(n_626), .B2(n_629), .C(n_631), .Y(n_622) );
INVx1_ASAP7_75t_L g599 ( .A(n_600), .Y(n_599) );
NAND2xp5_ASAP7_75t_L g657 ( .A(n_601), .B(n_658), .Y(n_657) );
AOI21xp33_ASAP7_75t_SL g603 ( .A1(n_604), .A2(n_605), .B(n_608), .Y(n_603) );
INVx2_ASAP7_75t_L g605 ( .A(n_606), .Y(n_605) );
CKINVDCx16_ASAP7_75t_R g705 ( .A(n_608), .Y(n_705) );
OR2x2_ASAP7_75t_L g608 ( .A(n_609), .B(n_610), .Y(n_608) );
OR2x2_ASAP7_75t_L g647 ( .A(n_610), .B(n_648), .Y(n_647) );
INVx1_ASAP7_75t_SL g668 ( .A(n_613), .Y(n_668) );
NAND2xp5_ASAP7_75t_L g713 ( .A(n_613), .B(n_673), .Y(n_713) );
NAND2xp5_ASAP7_75t_L g637 ( .A(n_616), .B(n_638), .Y(n_637) );
NOR2xp33_ASAP7_75t_L g617 ( .A(n_618), .B(n_619), .Y(n_617) );
NAND4xp25_ASAP7_75t_L g621 ( .A(n_622), .B(n_640), .C(n_659), .D(n_672), .Y(n_621) );
INVx1_ASAP7_75t_SL g623 ( .A(n_624), .Y(n_623) );
INVx1_ASAP7_75t_SL g630 ( .A(n_625), .Y(n_630) );
INVxp67_ASAP7_75t_L g626 ( .A(n_627), .Y(n_626) );
INVx1_ASAP7_75t_L g632 ( .A(n_633), .Y(n_632) );
OR2x2_ASAP7_75t_L g663 ( .A(n_634), .B(n_639), .Y(n_663) );
INVxp67_ASAP7_75t_L g635 ( .A(n_636), .Y(n_635) );
AOI211xp5_ASAP7_75t_L g640 ( .A1(n_641), .A2(n_642), .B(n_644), .C(n_652), .Y(n_640) );
AOI211xp5_ASAP7_75t_L g711 ( .A1(n_642), .A2(n_684), .B(n_712), .C(n_719), .Y(n_711) );
INVx1_ASAP7_75t_SL g671 ( .A(n_643), .Y(n_671) );
OAI22xp5_ASAP7_75t_L g644 ( .A1(n_645), .A2(n_647), .B1(n_649), .B2(n_650), .Y(n_644) );
INVx1_ASAP7_75t_L g675 ( .A(n_649), .Y(n_675) );
INVx1_ASAP7_75t_L g650 ( .A(n_651), .Y(n_650) );
NAND2xp5_ASAP7_75t_L g653 ( .A(n_654), .B(n_655), .Y(n_653) );
NAND2xp5_ASAP7_75t_L g691 ( .A(n_655), .B(n_692), .Y(n_691) );
NAND2xp5_ASAP7_75t_L g699 ( .A(n_655), .B(n_666), .Y(n_699) );
INVx2_ASAP7_75t_SL g655 ( .A(n_656), .Y(n_655) );
INVx1_ASAP7_75t_L g660 ( .A(n_661), .Y(n_660) );
INVx1_ASAP7_75t_SL g662 ( .A(n_663), .Y(n_662) );
INVx1_ASAP7_75t_L g664 ( .A(n_665), .Y(n_664) );
INVx1_ASAP7_75t_L g676 ( .A(n_666), .Y(n_676) );
AOI21xp33_ASAP7_75t_L g667 ( .A1(n_668), .A2(n_669), .B(n_671), .Y(n_667) );
INVxp33_ASAP7_75t_L g669 ( .A(n_670), .Y(n_669) );
AOI322xp5_ASAP7_75t_L g672 ( .A1(n_673), .A2(n_675), .A3(n_676), .B1(n_677), .B2(n_679), .C1(n_681), .C2(n_684), .Y(n_672) );
INVxp67_ASAP7_75t_L g677 ( .A(n_678), .Y(n_677) );
INVx1_ASAP7_75t_L g679 ( .A(n_680), .Y(n_679) );
INVx1_ASAP7_75t_L g681 ( .A(n_682), .Y(n_681) );
INVx1_ASAP7_75t_L g684 ( .A(n_685), .Y(n_684) );
NAND3xp33_ASAP7_75t_SL g686 ( .A(n_687), .B(n_704), .C(n_711), .Y(n_686) );
AOI221xp5_ASAP7_75t_L g687 ( .A1(n_688), .A2(n_690), .B1(n_693), .B2(n_695), .C(n_697), .Y(n_687) );
INVx1_ASAP7_75t_L g688 ( .A(n_689), .Y(n_688) );
INVx1_ASAP7_75t_L g690 ( .A(n_691), .Y(n_690) );
INVx1_ASAP7_75t_SL g703 ( .A(n_692), .Y(n_703) );
INVx1_ASAP7_75t_L g693 ( .A(n_694), .Y(n_693) );
INVxp67_ASAP7_75t_L g695 ( .A(n_696), .Y(n_695) );
OAI22xp33_ASAP7_75t_L g697 ( .A1(n_698), .A2(n_699), .B1(n_700), .B2(n_701), .Y(n_697) );
NAND2xp5_ASAP7_75t_L g701 ( .A(n_702), .B(n_703), .Y(n_701) );
AOI221xp5_ASAP7_75t_L g704 ( .A1(n_705), .A2(n_706), .B1(n_707), .B2(n_708), .C(n_709), .Y(n_704) );
NAND2xp33_ASAP7_75t_L g712 ( .A(n_713), .B(n_714), .Y(n_712) );
INVxp67_ASAP7_75t_L g716 ( .A(n_717), .Y(n_716) );
INVx2_ASAP7_75t_L g723 ( .A(n_724), .Y(n_723) );
INVx2_ASAP7_75t_L g732 ( .A(n_724), .Y(n_732) );
INVx1_ASAP7_75t_L g724 ( .A(n_725), .Y(n_724) );
NOR2x2_ASAP7_75t_L g735 ( .A(n_726), .B(n_736), .Y(n_735) );
INVxp67_ASAP7_75t_L g728 ( .A(n_729), .Y(n_728) );
INVx2_ASAP7_75t_L g734 ( .A(n_735), .Y(n_734) );
BUFx2_ASAP7_75t_L g737 ( .A(n_738), .Y(n_737) );
INVx2_ASAP7_75t_SL g752 ( .A(n_738), .Y(n_752) );
INVx2_ASAP7_75t_L g738 ( .A(n_739), .Y(n_738) );
NOR3xp33_ASAP7_75t_L g740 ( .A(n_741), .B(n_746), .C(n_749), .Y(n_740) );
INVx1_ASAP7_75t_L g748 ( .A(n_742), .Y(n_748) );
INVx1_ASAP7_75t_L g743 ( .A(n_744), .Y(n_743) );
NOR2xp33_ASAP7_75t_L g746 ( .A(n_747), .B(n_748), .Y(n_746) );
INVx1_ASAP7_75t_SL g749 ( .A(n_750), .Y(n_749) );
INVx1_ASAP7_75t_SL g756 ( .A(n_750), .Y(n_756) );
BUFx3_ASAP7_75t_L g751 ( .A(n_752), .Y(n_751) );
NOR2xp33_ASAP7_75t_L g753 ( .A(n_754), .B(n_755), .Y(n_753) );
INVx1_ASAP7_75t_SL g755 ( .A(n_756), .Y(n_755) );
endmodule