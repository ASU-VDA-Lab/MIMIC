module fake_ariane_3102_n_3213 (n_8, n_56, n_60, n_24, n_7, n_22, n_43, n_1, n_49, n_6, n_13, n_20, n_27, n_48, n_29, n_64, n_17, n_4, n_41, n_50, n_38, n_55, n_2, n_62, n_47, n_18, n_32, n_28, n_37, n_58, n_65, n_9, n_51, n_45, n_11, n_34, n_26, n_3, n_46, n_14, n_0, n_52, n_36, n_33, n_44, n_19, n_30, n_39, n_40, n_59, n_31, n_42, n_57, n_16, n_63, n_5, n_12, n_15, n_53, n_21, n_23, n_61, n_35, n_10, n_54, n_25, n_3213);

input n_8;
input n_56;
input n_60;
input n_24;
input n_7;
input n_22;
input n_43;
input n_1;
input n_49;
input n_6;
input n_13;
input n_20;
input n_27;
input n_48;
input n_29;
input n_64;
input n_17;
input n_4;
input n_41;
input n_50;
input n_38;
input n_55;
input n_2;
input n_62;
input n_47;
input n_18;
input n_32;
input n_28;
input n_37;
input n_58;
input n_65;
input n_9;
input n_51;
input n_45;
input n_11;
input n_34;
input n_26;
input n_3;
input n_46;
input n_14;
input n_0;
input n_52;
input n_36;
input n_33;
input n_44;
input n_19;
input n_30;
input n_39;
input n_40;
input n_59;
input n_31;
input n_42;
input n_57;
input n_16;
input n_63;
input n_5;
input n_12;
input n_15;
input n_53;
input n_21;
input n_23;
input n_61;
input n_35;
input n_10;
input n_54;
input n_25;

output n_3213;

wire n_2752;
wire n_913;
wire n_1681;
wire n_2163;
wire n_1486;
wire n_1507;
wire n_1938;
wire n_589;
wire n_2484;
wire n_2866;
wire n_3153;
wire n_1174;
wire n_3152;
wire n_2346;
wire n_1469;
wire n_691;
wire n_1353;
wire n_3056;
wire n_2679;
wire n_1355;
wire n_2131;
wire n_2559;
wire n_2500;
wire n_2509;
wire n_423;
wire n_1383;
wire n_2182;
wire n_603;
wire n_373;
wire n_2135;
wire n_2680;
wire n_2334;
wire n_1250;
wire n_2030;
wire n_1169;
wire n_789;
wire n_3181;
wire n_850;
wire n_2993;
wire n_1916;
wire n_2879;
wire n_610;
wire n_245;
wire n_1713;
wire n_96;
wire n_319;
wire n_1436;
wire n_2407;
wire n_690;
wire n_2818;
wire n_416;
wire n_1109;
wire n_1430;
wire n_2537;
wire n_525;
wire n_187;
wire n_2002;
wire n_1463;
wire n_2243;
wire n_1238;
wire n_2694;
wire n_2011;
wire n_2729;
wire n_1515;
wire n_817;
wire n_1837;
wire n_924;
wire n_781;
wire n_2013;
wire n_2786;
wire n_1566;
wire n_2837;
wire n_189;
wire n_717;
wire n_72;
wire n_2006;
wire n_952;
wire n_864;
wire n_2446;
wire n_1096;
wire n_1379;
wire n_2436;
wire n_2376;
wire n_2367;
wire n_2671;
wire n_2790;
wire n_1706;
wire n_2207;
wire n_2461;
wire n_2702;
wire n_117;
wire n_524;
wire n_2731;
wire n_634;
wire n_1214;
wire n_1839;
wire n_1246;
wire n_1138;
wire n_214;
wire n_2042;
wire n_2123;
wire n_3198;
wire n_1853;
wire n_764;
wire n_1503;
wire n_2238;
wire n_2529;
wire n_2374;
wire n_462;
wire n_1196;
wire n_1181;
wire n_1999;
wire n_410;
wire n_2380;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_3154;
wire n_2646;
wire n_737;
wire n_137;
wire n_1298;
wire n_2653;
wire n_1745;
wire n_2873;
wire n_1366;
wire n_232;
wire n_2084;
wire n_3115;
wire n_568;
wire n_2278;
wire n_1088;
wire n_77;
wire n_1424;
wire n_766;
wire n_2976;
wire n_1835;
wire n_1457;
wire n_377;
wire n_2482;
wire n_1682;
wire n_2750;
wire n_1836;
wire n_520;
wire n_870;
wire n_2547;
wire n_1453;
wire n_279;
wire n_945;
wire n_958;
wire n_2554;
wire n_3145;
wire n_2248;
wire n_3063;
wire n_813;
wire n_419;
wire n_1985;
wire n_2288;
wire n_2621;
wire n_2908;
wire n_3081;
wire n_146;
wire n_270;
wire n_338;
wire n_995;
wire n_2579;
wire n_285;
wire n_1909;
wire n_2156;
wire n_1184;
wire n_1961;
wire n_202;
wire n_1535;
wire n_2960;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_2323;
wire n_1073;
wire n_2844;
wire n_239;
wire n_402;
wire n_1979;
wire n_1277;
wire n_2107;
wire n_1746;
wire n_829;
wire n_1761;
wire n_1062;
wire n_339;
wire n_738;
wire n_1690;
wire n_2221;
wire n_2807;
wire n_672;
wire n_740;
wire n_1283;
wire n_167;
wire n_2317;
wire n_2838;
wire n_1974;
wire n_2906;
wire n_1736;
wire n_1018;
wire n_2342;
wire n_2200;
wire n_2781;
wire n_259;
wire n_69;
wire n_2442;
wire n_2735;
wire n_953;
wire n_1364;
wire n_2390;
wire n_143;
wire n_1888;
wire n_1224;
wire n_2109;
wire n_1425;
wire n_2634;
wire n_2709;
wire n_625;
wire n_557;
wire n_2746;
wire n_2322;
wire n_1107;
wire n_2832;
wire n_1688;
wire n_989;
wire n_242;
wire n_645;
wire n_1944;
wire n_331;
wire n_559;
wire n_2233;
wire n_2370;
wire n_2663;
wire n_267;
wire n_495;
wire n_2914;
wire n_1988;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_1936;
wire n_2149;
wire n_2277;
wire n_200;
wire n_1428;
wire n_1284;
wire n_2878;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_2539;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_2782;
wire n_569;
wire n_2078;
wire n_1145;
wire n_971;
wire n_3144;
wire n_2359;
wire n_2201;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_2049;
wire n_1522;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_1404;
wire n_868;
wire n_2232;
wire n_1847;
wire n_2458;
wire n_2779;
wire n_3150;
wire n_2950;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_2227;
wire n_2301;
wire n_1539;
wire n_2859;
wire n_3121;
wire n_2847;
wire n_884;
wire n_1851;
wire n_2162;
wire n_3209;
wire n_3015;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_2192;
wire n_1676;
wire n_1085;
wire n_277;
wire n_2988;
wire n_1636;
wire n_432;
wire n_293;
wire n_823;
wire n_1900;
wire n_620;
wire n_93;
wire n_1074;
wire n_859;
wire n_1765;
wire n_108;
wire n_1889;
wire n_587;
wire n_1977;
wire n_693;
wire n_863;
wire n_2650;
wire n_303;
wire n_1254;
wire n_929;
wire n_3207;
wire n_2433;
wire n_206;
wire n_352;
wire n_899;
wire n_1703;
wire n_2332;
wire n_2391;
wire n_3073;
wire n_611;
wire n_1295;
wire n_2060;
wire n_1850;
wire n_238;
wire n_365;
wire n_2004;
wire n_3183;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_2571;
wire n_136;
wire n_334;
wire n_2427;
wire n_192;
wire n_2885;
wire n_661;
wire n_2098;
wire n_2616;
wire n_1751;
wire n_2874;
wire n_3003;
wire n_300;
wire n_533;
wire n_3049;
wire n_3136;
wire n_2867;
wire n_1917;
wire n_2456;
wire n_2769;
wire n_104;
wire n_1924;
wire n_438;
wire n_1560;
wire n_1654;
wire n_2341;
wire n_2899;
wire n_1548;
wire n_3066;
wire n_1811;
wire n_2045;
wire n_440;
wire n_3013;
wire n_273;
wire n_2575;
wire n_2722;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_1840;
wire n_2739;
wire n_376;
wire n_512;
wire n_1597;
wire n_2942;
wire n_1771;
wire n_2902;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_2685;
wire n_2061;
wire n_3164;
wire n_2094;
wire n_2512;
wire n_1354;
wire n_1790;
wire n_149;
wire n_1213;
wire n_2382;
wire n_2956;
wire n_237;
wire n_2043;
wire n_780;
wire n_2349;
wire n_1918;
wire n_2788;
wire n_1021;
wire n_1443;
wire n_3089;
wire n_491;
wire n_2595;
wire n_1465;
wire n_2686;
wire n_3084;
wire n_1949;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_2727;
wire n_942;
wire n_1437;
wire n_2077;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_2909;
wire n_209;
wire n_490;
wire n_1461;
wire n_2717;
wire n_3012;
wire n_1391;
wire n_2981;
wire n_1947;
wire n_225;
wire n_1599;
wire n_1876;
wire n_1006;
wire n_1830;
wire n_575;
wire n_546;
wire n_503;
wire n_2527;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_3126;
wire n_2759;
wire n_1245;
wire n_2743;
wire n_1669;
wire n_2969;
wire n_1675;
wire n_2466;
wire n_676;
wire n_2038;
wire n_2263;
wire n_2800;
wire n_2568;
wire n_2116;
wire n_2271;
wire n_2145;
wire n_2326;
wire n_1838;
wire n_1594;
wire n_680;
wire n_1935;
wire n_2806;
wire n_287;
wire n_3191;
wire n_1716;
wire n_302;
wire n_1872;
wire n_380;
wire n_1585;
wire n_2281;
wire n_1432;
wire n_94;
wire n_2245;
wire n_3119;
wire n_249;
wire n_1108;
wire n_355;
wire n_212;
wire n_123;
wire n_444;
wire n_851;
wire n_1590;
wire n_1351;
wire n_2216;
wire n_1274;
wire n_257;
wire n_2426;
wire n_652;
wire n_1819;
wire n_475;
wire n_135;
wire n_3095;
wire n_947;
wire n_2134;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_102;
wire n_2703;
wire n_182;
wire n_696;
wire n_1442;
wire n_2926;
wire n_482;
wire n_2620;
wire n_798;
wire n_577;
wire n_1833;
wire n_407;
wire n_1691;
wire n_916;
wire n_1386;
wire n_2810;
wire n_912;
wire n_1884;
wire n_460;
wire n_1555;
wire n_1842;
wire n_2499;
wire n_2549;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_2791;
wire n_555;
wire n_2683;
wire n_3212;
wire n_804;
wire n_1656;
wire n_1382;
wire n_3093;
wire n_2970;
wire n_3159;
wire n_966;
wire n_992;
wire n_955;
wire n_1182;
wire n_794;
wire n_2855;
wire n_78;
wire n_2166;
wire n_2848;
wire n_1692;
wire n_3192;
wire n_2611;
wire n_1562;
wire n_514;
wire n_2748;
wire n_418;
wire n_2185;
wire n_3029;
wire n_2398;
wire n_1376;
wire n_513;
wire n_288;
wire n_179;
wire n_1292;
wire n_1178;
wire n_1972;
wire n_2015;
wire n_2925;
wire n_1435;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_2202;
wire n_2072;
wire n_306;
wire n_2952;
wire n_2415;
wire n_2693;
wire n_2877;
wire n_92;
wire n_3120;
wire n_203;
wire n_2922;
wire n_436;
wire n_3000;
wire n_150;
wire n_2871;
wire n_2930;
wire n_3193;
wire n_324;
wire n_2745;
wire n_2087;
wire n_669;
wire n_931;
wire n_1491;
wire n_2628;
wire n_619;
wire n_437;
wire n_337;
wire n_274;
wire n_111;
wire n_967;
wire n_1083;
wire n_2161;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1787;
wire n_2462;
wire n_1389;
wire n_3172;
wire n_2155;
wire n_2659;
wire n_615;
wire n_1139;
wire n_2836;
wire n_76;
wire n_2439;
wire n_2864;
wire n_517;
wire n_1312;
wire n_1717;
wire n_1812;
wire n_824;
wire n_428;
wire n_159;
wire n_2172;
wire n_2601;
wire n_892;
wire n_1880;
wire n_959;
wire n_2365;
wire n_2257;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_2219;
wire n_3116;
wire n_1855;
wire n_2100;
wire n_2333;
wire n_3176;
wire n_144;
wire n_990;
wire n_1623;
wire n_1903;
wire n_867;
wire n_2147;
wire n_2435;
wire n_1226;
wire n_2224;
wire n_944;
wire n_749;
wire n_1932;
wire n_1780;
wire n_2825;
wire n_2888;
wire n_1970;
wire n_1920;
wire n_2083;
wire n_815;
wire n_542;
wire n_2167;
wire n_2293;
wire n_2753;
wire n_1340;
wire n_470;
wire n_2668;
wire n_1240;
wire n_2921;
wire n_3046;
wire n_1087;
wire n_2701;
wire n_2400;
wire n_3021;
wire n_632;
wire n_477;
wire n_650;
wire n_2388;
wire n_425;
wire n_2273;
wire n_2712;
wire n_1433;
wire n_1911;
wire n_2567;
wire n_2557;
wire n_2695;
wire n_2898;
wire n_1908;
wire n_1825;
wire n_1155;
wire n_2598;
wire n_1071;
wire n_2755;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1832;
wire n_2795;
wire n_2682;
wire n_1841;
wire n_1680;
wire n_2066;
wire n_2302;
wire n_2762;
wire n_964;
wire n_1627;
wire n_2220;
wire n_2954;
wire n_382;
wire n_3014;
wire n_489;
wire n_2294;
wire n_80;
wire n_2274;
wire n_2895;
wire n_2903;
wire n_251;
wire n_974;
wire n_506;
wire n_3127;
wire n_1731;
wire n_799;
wire n_1147;
wire n_2829;
wire n_2378;
wire n_397;
wire n_2467;
wire n_2768;
wire n_471;
wire n_351;
wire n_965;
wire n_1914;
wire n_155;
wire n_2253;
wire n_934;
wire n_2213;
wire n_1447;
wire n_2363;
wire n_1220;
wire n_356;
wire n_2019;
wire n_698;
wire n_2728;
wire n_2130;
wire n_1674;
wire n_2021;
wire n_2025;
wire n_3010;
wire n_2160;
wire n_1992;
wire n_124;
wire n_2924;
wire n_307;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_3052;
wire n_646;
wire n_2507;
wire n_2142;
wire n_1633;
wire n_404;
wire n_2625;
wire n_2896;
wire n_172;
wire n_1913;
wire n_2069;
wire n_2495;
wire n_3187;
wire n_1058;
wire n_2328;
wire n_347;
wire n_2434;
wire n_1042;
wire n_3170;
wire n_183;
wire n_1234;
wire n_2311;
wire n_479;
wire n_1578;
wire n_2261;
wire n_1455;
wire n_3147;
wire n_2287;
wire n_299;
wire n_836;
wire n_2223;
wire n_3082;
wire n_1279;
wire n_2473;
wire n_2144;
wire n_2511;
wire n_564;
wire n_133;
wire n_205;
wire n_66;
wire n_1029;
wire n_2649;
wire n_1247;
wire n_760;
wire n_522;
wire n_2438;
wire n_1568;
wire n_2919;
wire n_3210;
wire n_1483;
wire n_3108;
wire n_1363;
wire n_2681;
wire n_367;
wire n_1111;
wire n_970;
wire n_1689;
wire n_2535;
wire n_713;
wire n_1255;
wire n_2632;
wire n_1646;
wire n_598;
wire n_3031;
wire n_345;
wire n_2262;
wire n_3179;
wire n_2565;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_2980;
wire n_1728;
wire n_2335;
wire n_3078;
wire n_370;
wire n_706;
wire n_2120;
wire n_286;
wire n_2631;
wire n_1401;
wire n_1419;
wire n_3138;
wire n_1531;
wire n_776;
wire n_424;
wire n_2860;
wire n_2041;
wire n_2113;
wire n_1933;
wire n_1651;
wire n_3087;
wire n_85;
wire n_130;
wire n_2697;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_1817;
wire n_2404;
wire n_2168;
wire n_2757;
wire n_348;
wire n_552;
wire n_2312;
wire n_670;
wire n_2677;
wire n_1826;
wire n_3171;
wire n_379;
wire n_162;
wire n_138;
wire n_264;
wire n_2834;
wire n_2483;
wire n_441;
wire n_1951;
wire n_3185;
wire n_2490;
wire n_1032;
wire n_1217;
wire n_2558;
wire n_1496;
wire n_2996;
wire n_637;
wire n_1592;
wire n_2812;
wire n_73;
wire n_327;
wire n_2662;
wire n_1259;
wire n_2801;
wire n_1177;
wire n_3104;
wire n_3074;
wire n_2655;
wire n_1231;
wire n_2132;
wire n_980;
wire n_1618;
wire n_1869;
wire n_1743;
wire n_905;
wire n_2718;
wire n_207;
wire n_720;
wire n_926;
wire n_1943;
wire n_2687;
wire n_2296;
wire n_194;
wire n_1802;
wire n_2178;
wire n_2112;
wire n_2765;
wire n_1163;
wire n_2640;
wire n_3054;
wire n_2811;
wire n_3019;
wire n_186;
wire n_1795;
wire n_3200;
wire n_1384;
wire n_2237;
wire n_145;
wire n_2146;
wire n_2983;
wire n_1868;
wire n_1501;
wire n_2241;
wire n_2373;
wire n_1173;
wire n_2350;
wire n_1068;
wire n_1198;
wire n_2531;
wire n_1570;
wire n_2099;
wire n_487;
wire n_1518;
wire n_1456;
wire n_90;
wire n_1879;
wire n_1886;
wire n_1648;
wire n_2187;
wire n_1413;
wire n_2617;
wire n_2481;
wire n_2129;
wire n_855;
wire n_2327;
wire n_158;
wire n_808;
wire n_1365;
wire n_2476;
wire n_553;
wire n_2814;
wire n_2059;
wire n_2437;
wire n_2636;
wire n_1439;
wire n_814;
wire n_578;
wire n_2074;
wire n_1665;
wire n_1287;
wire n_2841;
wire n_405;
wire n_1611;
wire n_2122;
wire n_120;
wire n_2975;
wire n_2399;
wire n_320;
wire n_1414;
wire n_1134;
wire n_2067;
wire n_1484;
wire n_1901;
wire n_647;
wire n_2055;
wire n_2998;
wire n_2027;
wire n_2932;
wire n_1423;
wire n_2117;
wire n_481;
wire n_600;
wire n_1053;
wire n_1609;
wire n_3118;
wire n_2822;
wire n_1939;
wire n_2308;
wire n_2242;
wire n_1906;
wire n_529;
wire n_1899;
wire n_3039;
wire n_2195;
wire n_502;
wire n_2194;
wire n_2937;
wire n_218;
wire n_1467;
wire n_247;
wire n_1828;
wire n_2159;
wire n_1798;
wire n_3057;
wire n_1608;
wire n_1304;
wire n_1744;
wire n_3007;
wire n_2267;
wire n_1105;
wire n_547;
wire n_439;
wire n_604;
wire n_677;
wire n_3022;
wire n_478;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_2102;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_2286;
wire n_2023;
wire n_1278;
wire n_707;
wire n_129;
wire n_126;
wire n_983;
wire n_3036;
wire n_2783;
wire n_2599;
wire n_590;
wire n_727;
wire n_699;
wire n_301;
wire n_1726;
wire n_2075;
wire n_2523;
wire n_1945;
wire n_545;
wire n_2418;
wire n_1015;
wire n_1614;
wire n_1162;
wire n_536;
wire n_1377;
wire n_2031;
wire n_2496;
wire n_2118;
wire n_325;
wire n_1740;
wire n_1602;
wire n_688;
wire n_3139;
wire n_636;
wire n_2853;
wire n_427;
wire n_1098;
wire n_3009;
wire n_1490;
wire n_2338;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_3025;
wire n_3051;
wire n_3205;
wire n_2225;
wire n_986;
wire n_1104;
wire n_2802;
wire n_1963;
wire n_3035;
wire n_729;
wire n_887;
wire n_2057;
wire n_2218;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_2593;
wire n_163;
wire n_1693;
wire n_2125;
wire n_2716;
wire n_1132;
wire n_390;
wire n_1156;
wire n_2741;
wire n_501;
wire n_2184;
wire n_2714;
wire n_314;
wire n_1823;
wire n_2944;
wire n_2861;
wire n_2780;
wire n_3023;
wire n_1120;
wire n_1202;
wire n_627;
wire n_2254;
wire n_3130;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_2033;
wire n_2618;
wire n_233;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_2754;
wire n_2707;
wire n_2774;
wire n_2849;
wire n_1607;
wire n_1489;
wire n_2799;
wire n_1218;
wire n_2756;
wire n_2217;
wire n_221;
wire n_321;
wire n_86;
wire n_2226;
wire n_1586;
wire n_861;
wire n_2962;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1863;
wire n_1763;
wire n_1666;
wire n_1500;
wire n_616;
wire n_2214;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_2763;
wire n_3156;
wire n_2256;
wire n_1189;
wire n_1089;
wire n_281;
wire n_1859;
wire n_2660;
wire n_262;
wire n_1502;
wire n_3044;
wire n_1523;
wire n_2190;
wire n_1478;
wire n_2732;
wire n_1883;
wire n_2516;
wire n_2776;
wire n_2555;
wire n_1969;
wire n_2708;
wire n_735;
wire n_297;
wire n_3070;
wire n_1005;
wire n_527;
wire n_2379;
wire n_84;
wire n_1294;
wire n_2661;
wire n_1667;
wire n_845;
wire n_888;
wire n_2894;
wire n_2300;
wire n_2949;
wire n_1649;
wire n_2452;
wire n_1677;
wire n_2470;
wire n_1927;
wire n_1297;
wire n_2827;
wire n_178;
wire n_551;
wire n_417;
wire n_1708;
wire n_70;
wire n_343;
wire n_3085;
wire n_1222;
wire n_2284;
wire n_3005;
wire n_1844;
wire n_2283;
wire n_582;
wire n_2526;
wire n_1957;
wire n_1953;
wire n_2643;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_1919;
wire n_2994;
wire n_534;
wire n_2508;
wire n_1791;
wire n_3186;
wire n_2124;
wire n_1894;
wire n_1460;
wire n_1239;
wire n_2594;
wire n_278;
wire n_2266;
wire n_2449;
wire n_560;
wire n_890;
wire n_842;
wire n_148;
wire n_1898;
wire n_451;
wire n_745;
wire n_1741;
wire n_1572;
wire n_1907;
wire n_1793;
wire n_3180;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1975;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_2119;
wire n_2742;
wire n_769;
wire n_1797;
wire n_2366;
wire n_2493;
wire n_1753;
wire n_1990;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_1895;
wire n_2821;
wire n_2690;
wire n_3090;
wire n_2474;
wire n_2623;
wire n_982;
wire n_1800;
wire n_915;
wire n_215;
wire n_1075;
wire n_2008;
wire n_454;
wire n_298;
wire n_1331;
wire n_1890;
wire n_2904;
wire n_3064;
wire n_3199;
wire n_1529;
wire n_1227;
wire n_2127;
wire n_655;
wire n_2946;
wire n_3166;
wire n_3151;
wire n_1734;
wire n_1860;
wire n_3065;
wire n_403;
wire n_3016;
wire n_2785;
wire n_2460;
wire n_2840;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_3135;
wire n_657;
wire n_837;
wire n_812;
wire n_2448;
wire n_2211;
wire n_2292;
wire n_2480;
wire n_606;
wire n_951;
wire n_3024;
wire n_2772;
wire n_862;
wire n_1700;
wire n_2637;
wire n_659;
wire n_1332;
wire n_2306;
wire n_509;
wire n_1854;
wire n_666;
wire n_1747;
wire n_2071;
wire n_2424;
wire n_430;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_2414;
wire n_2893;
wire n_2959;
wire n_2082;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_3161;
wire n_3208;
wire n_2389;
wire n_1309;
wire n_999;
wire n_2280;
wire n_1766;
wire n_1338;
wire n_2978;
wire n_1342;
wire n_2737;
wire n_456;
wire n_1867;
wire n_852;
wire n_1394;
wire n_2916;
wire n_2576;
wire n_704;
wire n_2958;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_2696;
wire n_521;
wire n_2140;
wire n_873;
wire n_1301;
wire n_1748;
wire n_2157;
wire n_2468;
wire n_1243;
wire n_2171;
wire n_1966;
wire n_1400;
wire n_342;
wire n_2035;
wire n_2614;
wire n_1466;
wire n_1513;
wire n_1527;
wire n_2581;
wire n_358;
wire n_1783;
wire n_608;
wire n_2494;
wire n_1538;
wire n_2831;
wire n_2457;
wire n_2128;
wire n_3069;
wire n_2992;
wire n_1037;
wire n_1329;
wire n_317;
wire n_3197;
wire n_1993;
wire n_1545;
wire n_134;
wire n_2629;
wire n_1257;
wire n_1480;
wire n_1954;
wire n_1668;
wire n_1878;
wire n_2540;
wire n_1605;
wire n_1078;
wire n_3060;
wire n_266;
wire n_2486;
wire n_1897;
wire n_2984;
wire n_157;
wire n_2520;
wire n_2137;
wire n_1161;
wire n_2489;
wire n_811;
wire n_3097;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_2492;
wire n_2939;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_2337;
wire n_2265;
wire n_687;
wire n_2900;
wire n_797;
wire n_2026;
wire n_2912;
wire n_1786;
wire n_2627;
wire n_3173;
wire n_480;
wire n_1327;
wire n_1475;
wire n_211;
wire n_642;
wire n_2106;
wire n_1804;
wire n_97;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_2684;
wire n_3174;
wire n_2726;
wire n_602;
wire n_2622;
wire n_2272;
wire n_1757;
wire n_592;
wire n_3102;
wire n_1499;
wire n_854;
wire n_1318;
wire n_2091;
wire n_393;
wire n_1632;
wire n_1769;
wire n_474;
wire n_1929;
wire n_2264;
wire n_2691;
wire n_1950;
wire n_805;
wire n_2032;
wire n_2090;
wire n_2929;
wire n_3124;
wire n_295;
wire n_1658;
wire n_190;
wire n_2249;
wire n_1072;
wire n_695;
wire n_1526;
wire n_2991;
wire n_1305;
wire n_180;
wire n_730;
wire n_386;
wire n_1596;
wire n_2348;
wire n_2656;
wire n_1281;
wire n_516;
wire n_2364;
wire n_2574;
wire n_1997;
wire n_1137;
wire n_1873;
wire n_1258;
wire n_197;
wire n_640;
wire n_463;
wire n_1476;
wire n_1733;
wire n_1524;
wire n_1856;
wire n_2016;
wire n_2667;
wire n_2723;
wire n_2725;
wire n_2928;
wire n_943;
wire n_1118;
wire n_678;
wire n_2905;
wire n_2884;
wire n_651;
wire n_2850;
wire n_1874;
wire n_1293;
wire n_3167;
wire n_961;
wire n_469;
wire n_1046;
wire n_1807;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_2857;
wire n_1784;
wire n_3110;
wire n_771;
wire n_1321;
wire n_3050;
wire n_3157;
wire n_752;
wire n_2307;
wire n_71;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_2295;
wire n_2730;
wire n_283;
wire n_806;
wire n_3142;
wire n_1984;
wire n_1350;
wire n_3129;
wire n_1556;
wire n_649;
wire n_1561;
wire n_2412;
wire n_2720;
wire n_374;
wire n_3107;
wire n_1352;
wire n_2405;
wire n_2815;
wire n_1824;
wire n_643;
wire n_2606;
wire n_2700;
wire n_1492;
wire n_226;
wire n_2383;
wire n_2764;
wire n_1441;
wire n_1822;
wire n_682;
wire n_1616;
wire n_2633;
wire n_2416;
wire n_819;
wire n_2386;
wire n_2907;
wire n_1971;
wire n_2945;
wire n_586;
wire n_1324;
wire n_1429;
wire n_2064;
wire n_2353;
wire n_2528;
wire n_1778;
wire n_1776;
wire n_686;
wire n_605;
wire n_2936;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1759;
wire n_1829;
wire n_2325;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_2022;
wire n_1016;
wire n_2298;
wire n_1149;
wire n_1505;
wire n_2408;
wire n_2698;
wire n_2986;
wire n_2320;
wire n_3017;
wire n_979;
wire n_2570;
wire n_2329;
wire n_3140;
wire n_1642;
wire n_2417;
wire n_2789;
wire n_2525;
wire n_1815;
wire n_2813;
wire n_897;
wire n_2546;
wire n_949;
wire n_2454;
wire n_1493;
wire n_2890;
wire n_2911;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_2354;
wire n_198;
wire n_1864;
wire n_2760;
wire n_3086;
wire n_1887;
wire n_3165;
wire n_1208;
wire n_1987;
wire n_396;
wire n_2368;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_2352;
wire n_2502;
wire n_1256;
wire n_87;
wire n_714;
wire n_2170;
wire n_790;
wire n_2244;
wire n_2143;
wire n_2393;
wire n_354;
wire n_140;
wire n_725;
wire n_2377;
wire n_1577;
wire n_151;
wire n_1448;
wire n_2198;
wire n_1009;
wire n_230;
wire n_2652;
wire n_1133;
wire n_3067;
wire n_154;
wire n_883;
wire n_142;
wire n_473;
wire n_1852;
wire n_801;
wire n_1286;
wire n_2612;
wire n_818;
wire n_1685;
wire n_779;
wire n_2410;
wire n_2314;
wire n_2477;
wire n_2279;
wire n_3169;
wire n_594;
wire n_2222;
wire n_1995;
wire n_1877;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_1849;
wire n_2203;
wire n_2133;
wire n_2076;
wire n_833;
wire n_2943;
wire n_1426;
wire n_2250;
wire n_2497;
wire n_2247;
wire n_2230;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_75;
wire n_2001;
wire n_1047;
wire n_95;
wire n_2506;
wire n_1472;
wire n_2413;
wire n_1593;
wire n_2610;
wire n_1050;
wire n_2626;
wire n_566;
wire n_2158;
wire n_2578;
wire n_2607;
wire n_2285;
wire n_3184;
wire n_152;
wire n_2892;
wire n_169;
wire n_106;
wire n_1201;
wire n_1288;
wire n_173;
wire n_2605;
wire n_858;
wire n_2796;
wire n_1185;
wire n_2475;
wire n_2804;
wire n_2173;
wire n_2715;
wire n_3206;
wire n_335;
wire n_1035;
wire n_1143;
wire n_2665;
wire n_344;
wire n_2070;
wire n_2136;
wire n_426;
wire n_433;
wire n_3134;
wire n_398;
wire n_2771;
wire n_210;
wire n_2403;
wire n_1090;
wire n_2947;
wire n_1367;
wire n_2044;
wire n_253;
wire n_166;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_2619;
wire n_1565;
wire n_1192;
wire n_128;
wire n_224;
wire n_82;
wire n_894;
wire n_3098;
wire n_1380;
wire n_1624;
wire n_1801;
wire n_2854;
wire n_3055;
wire n_420;
wire n_1291;
wire n_562;
wire n_2020;
wire n_748;
wire n_2310;
wire n_510;
wire n_1045;
wire n_256;
wire n_3160;
wire n_1160;
wire n_2968;
wire n_1882;
wire n_1976;
wire n_1023;
wire n_2711;
wire n_1881;
wire n_2635;
wire n_2999;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_3043;
wire n_3190;
wire n_1958;
wire n_2747;
wire n_3027;
wire n_467;
wire n_1511;
wire n_2177;
wire n_2713;
wire n_1422;
wire n_2766;
wire n_1965;
wire n_644;
wire n_1197;
wire n_3011;
wire n_276;
wire n_2820;
wire n_2613;
wire n_497;
wire n_1165;
wire n_2934;
wire n_1641;
wire n_168;
wire n_81;
wire n_538;
wire n_2845;
wire n_1517;
wire n_2036;
wire n_576;
wire n_843;
wire n_511;
wire n_2647;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_2003;
wire n_2533;
wire n_2210;
wire n_1307;
wire n_1128;
wire n_3141;
wire n_2053;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_2343;
wire n_775;
wire n_3096;
wire n_667;
wire n_2419;
wire n_1049;
wire n_2330;
wire n_2826;
wire n_869;
wire n_141;
wire n_846;
wire n_1398;
wire n_1921;
wire n_2777;
wire n_2450;
wire n_2411;
wire n_1356;
wire n_1341;
wire n_2234;
wire n_2309;
wire n_3189;
wire n_1504;
wire n_1955;
wire n_2110;
wire n_2431;
wire n_1773;
wire n_3175;
wire n_1440;
wire n_2666;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_2935;
wire n_2401;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_2588;
wire n_2863;
wire n_2331;
wire n_935;
wire n_2886;
wire n_2478;
wire n_685;
wire n_911;
wire n_361;
wire n_89;
wire n_2658;
wire n_623;
wire n_2608;
wire n_2920;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_3006;
wire n_1948;
wire n_74;
wire n_2767;
wire n_810;
wire n_1290;
wire n_181;
wire n_1959;
wire n_617;
wire n_2396;
wire n_543;
wire n_1362;
wire n_1559;
wire n_2121;
wire n_3123;
wire n_2692;
wire n_236;
wire n_683;
wire n_601;
wire n_565;
wire n_628;
wire n_1300;
wire n_1960;
wire n_2068;
wire n_3117;
wire n_743;
wire n_1194;
wire n_2862;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_2553;
wire n_2645;
wire n_907;
wire n_2749;
wire n_1454;
wire n_2592;
wire n_660;
wire n_464;
wire n_2459;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_2566;
wire n_2751;
wire n_3113;
wire n_3101;
wire n_918;
wire n_1968;
wire n_107;
wire n_1885;
wire n_639;
wire n_452;
wire n_673;
wire n_2842;
wire n_2833;
wire n_2196;
wire n_1038;
wire n_2371;
wire n_1978;
wire n_414;
wire n_571;
wire n_1521;
wire n_1694;
wire n_1940;
wire n_284;
wire n_593;
wire n_3195;
wire n_3008;
wire n_1695;
wire n_2560;
wire n_1164;
wire n_2313;
wire n_609;
wire n_3077;
wire n_1193;
wire n_3048;
wire n_1345;
wire n_613;
wire n_3037;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_3062;
wire n_1774;
wire n_409;
wire n_171;
wire n_2963;
wire n_519;
wire n_384;
wire n_2609;
wire n_2561;
wire n_1166;
wire n_1056;
wire n_2007;
wire n_526;
wire n_1994;
wire n_1767;
wire n_1040;
wire n_674;
wire n_3131;
wire n_1158;
wire n_316;
wire n_3168;
wire n_125;
wire n_1973;
wire n_1444;
wire n_1803;
wire n_820;
wire n_1749;
wire n_872;
wire n_1653;
wire n_254;
wire n_2882;
wire n_2303;
wire n_2669;
wire n_1157;
wire n_1584;
wire n_234;
wire n_848;
wire n_1664;
wire n_280;
wire n_629;
wire n_1739;
wire n_161;
wire n_2642;
wire n_1814;
wire n_532;
wire n_2154;
wire n_2441;
wire n_2236;
wire n_1789;
wire n_763;
wire n_1986;
wire n_2174;
wire n_2688;
wire n_99;
wire n_540;
wire n_216;
wire n_692;
wire n_2624;
wire n_2054;
wire n_1857;
wire n_2315;
wire n_984;
wire n_1687;
wire n_2073;
wire n_223;
wire n_2150;
wire n_1552;
wire n_750;
wire n_2938;
wire n_834;
wire n_1612;
wire n_2498;
wire n_800;
wire n_2638;
wire n_2046;
wire n_1910;
wire n_1816;
wire n_2803;
wire n_1756;
wire n_2887;
wire n_1606;
wire n_2189;
wire n_395;
wire n_621;
wire n_2648;
wire n_1587;
wire n_213;
wire n_2093;
wire n_2340;
wire n_2018;
wire n_2672;
wire n_1772;
wire n_67;
wire n_2444;
wire n_2602;
wire n_1014;
wire n_724;
wire n_2204;
wire n_2931;
wire n_1427;
wire n_1481;
wire n_2040;
wire n_493;
wire n_1311;
wire n_2977;
wire n_3106;
wire n_2199;
wire n_2881;
wire n_1956;
wire n_1589;
wire n_114;
wire n_2151;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_2455;
wire n_827;
wire n_2600;
wire n_3092;
wire n_2231;
wire n_697;
wire n_2828;
wire n_622;
wire n_1626;
wire n_1962;
wire n_1335;
wire n_1715;
wire n_296;
wire n_2305;
wire n_880;
wire n_793;
wire n_2114;
wire n_2927;
wire n_1175;
wire n_2289;
wire n_132;
wire n_2530;
wire n_2299;
wire n_751;
wire n_1027;
wire n_1070;
wire n_2406;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_2883;
wire n_1221;
wire n_530;
wire n_1785;
wire n_792;
wire n_1262;
wire n_1942;
wire n_2180;
wire n_2951;
wire n_580;
wire n_1579;
wire n_494;
wire n_2809;
wire n_2181;
wire n_434;
wire n_2014;
wire n_975;
wire n_2974;
wire n_229;
wire n_394;
wire n_923;
wire n_1645;
wire n_1381;
wire n_1124;
wire n_2870;
wire n_1494;
wire n_932;
wire n_1893;
wire n_1183;
wire n_1326;
wire n_2889;
wire n_2276;
wire n_1805;
wire n_2282;
wire n_981;
wire n_2910;
wire n_2141;
wire n_1110;
wire n_1758;
wire n_2503;
wire n_2270;
wire n_243;
wire n_2443;
wire n_1407;
wire n_185;
wire n_2465;
wire n_1204;
wire n_2865;
wire n_1554;
wire n_994;
wire n_2428;
wire n_2972;
wire n_2586;
wire n_2989;
wire n_1360;
wire n_973;
wire n_3178;
wire n_2858;
wire n_268;
wire n_972;
wire n_2251;
wire n_2923;
wire n_3076;
wire n_164;
wire n_2843;
wire n_184;
wire n_856;
wire n_3100;
wire n_2572;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_2010;
wire n_1054;
wire n_508;
wire n_121;
wire n_118;
wire n_1679;
wire n_2872;
wire n_2126;
wire n_3109;
wire n_1952;
wire n_2425;
wire n_2394;
wire n_1858;
wire n_353;
wire n_3125;
wire n_1678;
wire n_2589;
wire n_1482;
wire n_1361;
wire n_2356;
wire n_1601;
wire n_1057;
wire n_191;
wire n_2487;
wire n_1834;
wire n_978;
wire n_1011;
wire n_1520;
wire n_2534;
wire n_2488;
wire n_1509;
wire n_828;
wire n_2941;
wire n_322;
wire n_1411;
wire n_1359;
wire n_3079;
wire n_558;
wire n_1721;
wire n_2564;
wire n_116;
wire n_2591;
wire n_653;
wire n_1445;
wire n_1317;
wire n_3034;
wire n_2050;
wire n_2197;
wire n_783;
wire n_2550;
wire n_556;
wire n_1127;
wire n_170;
wire n_1536;
wire n_3177;
wire n_1471;
wire n_2385;
wire n_160;
wire n_119;
wire n_2387;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_3091;
wire n_1024;
wire n_830;
wire n_176;
wire n_2291;
wire n_2816;
wire n_1980;
wire n_2518;
wire n_987;
wire n_936;
wire n_2510;
wire n_1620;
wire n_2501;
wire n_2542;
wire n_3105;
wire n_1385;
wire n_1525;
wire n_2793;
wire n_1998;
wire n_2165;
wire n_2675;
wire n_541;
wire n_499;
wire n_2604;
wire n_1775;
wire n_908;
wire n_788;
wire n_2639;
wire n_1036;
wire n_2169;
wire n_2985;
wire n_2603;
wire n_341;
wire n_1270;
wire n_109;
wire n_1167;
wire n_1272;
wire n_549;
wire n_2630;
wire n_591;
wire n_2794;
wire n_969;
wire n_2028;
wire n_919;
wire n_1663;
wire n_3114;
wire n_2901;
wire n_2092;
wire n_2175;
wire n_1625;
wire n_2086;
wire n_2817;
wire n_2773;
wire n_1926;
wire n_2402;
wire n_318;
wire n_1458;
wire n_103;
wire n_244;
wire n_679;
wire n_1630;
wire n_220;
wire n_3047;
wire n_663;
wire n_1720;
wire n_2409;
wire n_2966;
wire n_3163;
wire n_443;
wire n_2176;
wire n_1412;
wire n_3059;
wire n_1738;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_139;
wire n_2808;
wire n_2453;
wire n_2344;
wire n_1922;
wire n_1735;
wire n_1788;
wire n_391;
wire n_940;
wire n_2392;
wire n_1537;
wire n_2138;
wire n_3122;
wire n_3040;
wire n_2065;
wire n_2543;
wire n_2321;
wire n_1077;
wire n_2597;
wire n_607;
wire n_956;
wire n_445;
wire n_1930;
wire n_765;
wire n_1809;
wire n_2787;
wire n_1904;
wire n_1843;
wire n_122;
wire n_2000;
wire n_3133;
wire n_2805;
wire n_1268;
wire n_2676;
wire n_2758;
wire n_385;
wire n_3211;
wire n_2395;
wire n_917;
wire n_2868;
wire n_1271;
wire n_372;
wire n_2096;
wire n_2440;
wire n_2556;
wire n_2186;
wire n_1530;
wire n_2215;
wire n_2770;
wire n_631;
wire n_399;
wire n_1170;
wire n_2724;
wire n_2258;
wire n_1261;
wire n_2471;
wire n_702;
wire n_857;
wire n_898;
wire n_3042;
wire n_363;
wire n_968;
wire n_1067;
wire n_1235;
wire n_1323;
wire n_2584;
wire n_2375;
wire n_1462;
wire n_1937;
wire n_2012;
wire n_3182;
wire n_2967;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_3004;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_2039;
wire n_1755;
wire n_1285;
wire n_3111;
wire n_193;
wire n_733;
wire n_761;
wire n_2212;
wire n_731;
wire n_336;
wire n_1813;
wire n_315;
wire n_2268;
wire n_2997;
wire n_311;
wire n_1452;
wire n_2835;
wire n_1573;
wire n_2734;
wire n_668;
wire n_2569;
wire n_758;
wire n_2252;
wire n_2111;
wire n_2420;
wire n_2948;
wire n_3099;
wire n_1996;
wire n_1106;
wire n_2009;
wire n_153;
wire n_648;
wire n_784;
wire n_269;
wire n_816;
wire n_2897;
wire n_1322;
wire n_2583;
wire n_2918;
wire n_2987;
wire n_1473;
wire n_835;
wire n_3155;
wire n_446;
wire n_1076;
wire n_2024;
wire n_1348;
wire n_2651;
wire n_753;
wire n_2445;
wire n_2733;
wire n_1770;
wire n_701;
wire n_1003;
wire n_2469;
wire n_1125;
wire n_2103;
wire n_2358;
wire n_1710;
wire n_1865;
wire n_2522;
wire n_2641;
wire n_2463;
wire n_309;
wire n_1344;
wire n_115;
wire n_2355;
wire n_1390;
wire n_2699;
wire n_2580;
wire n_401;
wire n_485;
wire n_1792;
wire n_504;
wire n_2062;
wire n_483;
wire n_435;
wire n_3068;
wire n_1141;
wire n_1629;
wire n_291;
wire n_1640;
wire n_822;
wire n_1094;
wire n_2973;
wire n_840;
wire n_1459;
wire n_2153;
wire n_2324;
wire n_1510;
wire n_3002;
wire n_2710;
wire n_2505;
wire n_2139;
wire n_1099;
wire n_839;
wire n_79;
wire n_1754;
wire n_3146;
wire n_3038;
wire n_759;
wire n_567;
wire n_2397;
wire n_91;
wire n_2521;
wire n_240;
wire n_369;
wire n_1727;
wire n_2740;
wire n_2235;
wire n_1991;
wire n_1575;
wire n_2721;
wire n_1848;
wire n_1892;
wire n_1172;
wire n_3132;
wire n_2615;
wire n_614;
wire n_2775;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_2351;
wire n_188;
wire n_2260;
wire n_323;
wire n_550;
wire n_1315;
wire n_1660;
wire n_1902;
wire n_997;
wire n_635;
wire n_2206;
wire n_2784;
wire n_2541;
wire n_694;
wire n_1643;
wire n_1320;
wire n_3188;
wire n_3001;
wire n_1113;
wire n_2347;
wire n_248;
wire n_1152;
wire n_2657;
wire n_2990;
wire n_2447;
wire n_2538;
wire n_2034;
wire n_1845;
wire n_1934;
wire n_2101;
wire n_2577;
wire n_921;
wire n_2362;
wire n_1615;
wire n_1236;
wire n_228;
wire n_2104;
wire n_1265;
wire n_1576;
wire n_2105;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1806;
wire n_2552;
wire n_2372;
wire n_1409;
wire n_1148;
wire n_1684;
wire n_1588;
wire n_1673;
wire n_2422;
wire n_2704;
wire n_1334;
wire n_654;
wire n_2290;
wire n_2933;
wire n_2856;
wire n_2088;
wire n_1275;
wire n_3103;
wire n_488;
wire n_3018;
wire n_904;
wire n_505;
wire n_88;
wire n_2005;
wire n_2048;
wire n_1696;
wire n_498;
wire n_3028;
wire n_1875;
wire n_1059;
wire n_3148;
wire n_684;
wire n_2429;
wire n_2108;
wire n_2736;
wire n_1039;
wire n_2246;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_2339;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1831;
wire n_2532;
wire n_2191;
wire n_2971;
wire n_1497;
wire n_1866;
wire n_2472;
wire n_2664;
wire n_2705;
wire n_2056;
wire n_2852;
wire n_459;
wire n_1136;
wire n_2515;
wire n_1782;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_3203;
wire n_383;
wire n_838;
wire n_1558;
wire n_1941;
wire n_1316;
wire n_175;
wire n_2519;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_1915;
wire n_2360;
wire n_723;
wire n_1393;
wire n_2240;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_2846;
wire n_310;
wire n_1781;
wire n_709;
wire n_2917;
wire n_3137;
wire n_2544;
wire n_809;
wire n_3143;
wire n_3194;
wire n_2432;
wire n_2085;
wire n_3032;
wire n_1686;
wire n_1964;
wire n_235;
wire n_881;
wire n_1019;
wire n_1477;
wire n_1777;
wire n_2188;
wire n_1982;
wire n_2097;
wire n_662;
wire n_641;
wire n_2430;
wire n_2504;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_2297;
wire n_3094;
wire n_371;
wire n_199;
wire n_3020;
wire n_217;
wire n_2964;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_708;
wire n_308;
wire n_1223;
wire n_2545;
wire n_201;
wire n_1768;
wire n_2513;
wire n_2193;
wire n_2369;
wire n_572;
wire n_1199;
wire n_2957;
wire n_865;
wire n_1273;
wire n_1983;
wire n_2982;
wire n_1041;
wire n_2451;
wire n_2115;
wire n_2913;
wire n_993;
wire n_1862;
wire n_948;
wire n_2017;
wire n_922;
wire n_1004;
wire n_1810;
wire n_3061;
wire n_448;
wire n_2587;
wire n_1347;
wire n_2839;
wire n_860;
wire n_3072;
wire n_1043;
wire n_2961;
wire n_255;
wire n_2869;
wire n_450;
wire n_1923;
wire n_2955;
wire n_2670;
wire n_1764;
wire n_2674;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_3026;
wire n_2644;
wire n_902;
wire n_1031;
wire n_2979;
wire n_1723;
wire n_1638;
wire n_853;
wire n_3071;
wire n_716;
wire n_1571;
wire n_1698;
wire n_196;
wire n_1337;
wire n_774;
wire n_2148;
wire n_1946;
wire n_933;
wire n_3112;
wire n_2562;
wire n_596;
wire n_954;
wire n_2051;
wire n_1779;
wire n_1168;
wire n_1821;
wire n_219;
wire n_1310;
wire n_3196;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_2673;
wire n_252;
wire n_664;
wire n_1591;
wire n_2585;
wire n_2995;
wire n_1229;
wire n_1683;
wire n_2582;
wire n_2548;
wire n_68;
wire n_1896;
wire n_2164;
wire n_1732;
wire n_415;
wire n_2381;
wire n_2744;
wire n_1967;
wire n_2678;
wire n_2384;
wire n_2179;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_2052;
wire n_2485;
wire n_3149;
wire n_537;
wire n_1063;
wire n_991;
wire n_2183;
wire n_2205;
wire n_83;
wire n_2275;
wire n_389;
wire n_2563;
wire n_1724;
wire n_3088;
wire n_1670;
wire n_1707;
wire n_1799;
wire n_2080;
wire n_2058;
wire n_1126;
wire n_2761;
wire n_2357;
wire n_2029;
wire n_195;
wire n_1846;
wire n_1912;
wire n_938;
wire n_1891;
wire n_1328;
wire n_895;
wire n_110;
wire n_304;
wire n_2875;
wire n_1639;
wire n_583;
wire n_2209;
wire n_2421;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_1928;
wire n_98;
wire n_946;
wire n_757;
wire n_2047;
wire n_3058;
wire n_375;
wire n_113;
wire n_1655;
wire n_1818;
wire n_1146;
wire n_2792;
wire n_1634;
wire n_2596;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_2269;
wire n_472;
wire n_937;
wire n_1474;
wire n_2081;
wire n_2536;
wire n_2524;
wire n_265;
wire n_1583;
wire n_1604;
wire n_208;
wire n_1631;
wire n_1702;
wire n_156;
wire n_174;
wire n_275;
wire n_100;
wire n_3202;
wire n_1794;
wire n_1375;
wire n_3053;
wire n_147;
wire n_204;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_496;
wire n_2891;
wire n_2318;
wire n_1827;
wire n_3128;
wire n_866;
wire n_246;
wire n_925;
wire n_1752;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_2361;
wire n_1115;
wire n_2229;
wire n_2819;
wire n_2880;
wire n_3030;
wire n_3075;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_105;
wire n_1051;
wire n_2551;
wire n_719;
wire n_131;
wire n_263;
wire n_1102;
wire n_360;
wire n_2255;
wire n_1129;
wire n_1252;
wire n_2239;
wire n_3045;
wire n_250;
wire n_1464;
wire n_1296;
wire n_3158;
wire n_773;
wire n_2798;
wire n_2316;
wire n_165;
wire n_2464;
wire n_1010;
wire n_2830;
wire n_882;
wire n_2706;
wire n_2304;
wire n_1249;
wire n_101;
wire n_803;
wire n_1871;
wire n_2514;
wire n_329;
wire n_718;
wire n_1434;
wire n_340;
wire n_1905;
wire n_1569;
wire n_3201;
wire n_2573;
wire n_2940;
wire n_289;
wire n_112;
wire n_548;
wire n_2336;
wire n_523;
wire n_1662;
wire n_3162;
wire n_457;
wire n_1299;
wire n_1870;
wire n_177;
wire n_2063;
wire n_1925;
wire n_782;
wire n_364;
wire n_258;
wire n_2915;
wire n_3083;
wire n_431;
wire n_2654;
wire n_2491;
wire n_1861;
wire n_2079;
wire n_1228;
wire n_2319;
wire n_2152;
wire n_2517;
wire n_1931;
wire n_1244;
wire n_1796;
wire n_411;
wire n_484;
wire n_2259;
wire n_849;
wire n_2095;
wire n_2719;
wire n_2965;
wire n_2738;
wire n_1820;
wire n_2590;
wire n_2876;
wire n_2797;
wire n_357;
wire n_412;
wire n_1251;
wire n_1989;
wire n_3041;
wire n_447;
wire n_1421;
wire n_2208;
wire n_2689;
wire n_2423;
wire n_2778;
wire n_1762;
wire n_1233;
wire n_3080;
wire n_1808;
wire n_1574;
wire n_1672;
wire n_2228;
wire n_1635;
wire n_3033;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_2479;
wire n_3204;
wire n_886;
wire n_1069;
wire n_1981;
wire n_2824;
wire n_2037;
wire n_2953;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_2851;
wire n_2823;
wire n_127;
wire n_531;
wire n_2345;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_2089;
wire n_1487;
wire n_675;

INVx1_ASAP7_75t_L g66 ( 
.A(n_25),
.Y(n_66)
);

CKINVDCx5p33_ASAP7_75t_R g67 ( 
.A(n_21),
.Y(n_67)
);

CKINVDCx5p33_ASAP7_75t_R g68 ( 
.A(n_31),
.Y(n_68)
);

CKINVDCx5p33_ASAP7_75t_R g69 ( 
.A(n_15),
.Y(n_69)
);

CKINVDCx5p33_ASAP7_75t_R g70 ( 
.A(n_6),
.Y(n_70)
);

CKINVDCx5p33_ASAP7_75t_R g71 ( 
.A(n_54),
.Y(n_71)
);

INVx2_ASAP7_75t_SL g72 ( 
.A(n_9),
.Y(n_72)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_11),
.Y(n_73)
);

CKINVDCx5p33_ASAP7_75t_R g74 ( 
.A(n_14),
.Y(n_74)
);

CKINVDCx5p33_ASAP7_75t_R g75 ( 
.A(n_25),
.Y(n_75)
);

CKINVDCx5p33_ASAP7_75t_R g76 ( 
.A(n_57),
.Y(n_76)
);

INVx2_ASAP7_75t_SL g77 ( 
.A(n_29),
.Y(n_77)
);

CKINVDCx5p33_ASAP7_75t_R g78 ( 
.A(n_56),
.Y(n_78)
);

CKINVDCx5p33_ASAP7_75t_R g79 ( 
.A(n_50),
.Y(n_79)
);

CKINVDCx5p33_ASAP7_75t_R g80 ( 
.A(n_28),
.Y(n_80)
);

CKINVDCx5p33_ASAP7_75t_R g81 ( 
.A(n_60),
.Y(n_81)
);

BUFx10_ASAP7_75t_L g82 ( 
.A(n_42),
.Y(n_82)
);

CKINVDCx5p33_ASAP7_75t_R g83 ( 
.A(n_36),
.Y(n_83)
);

CKINVDCx5p33_ASAP7_75t_R g84 ( 
.A(n_8),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_12),
.Y(n_85)
);

CKINVDCx5p33_ASAP7_75t_R g86 ( 
.A(n_3),
.Y(n_86)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_30),
.Y(n_87)
);

CKINVDCx5p33_ASAP7_75t_R g88 ( 
.A(n_28),
.Y(n_88)
);

CKINVDCx5p33_ASAP7_75t_R g89 ( 
.A(n_38),
.Y(n_89)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_16),
.Y(n_90)
);

CKINVDCx5p33_ASAP7_75t_R g91 ( 
.A(n_8),
.Y(n_91)
);

CKINVDCx16_ASAP7_75t_R g92 ( 
.A(n_33),
.Y(n_92)
);

CKINVDCx5p33_ASAP7_75t_R g93 ( 
.A(n_27),
.Y(n_93)
);

CKINVDCx5p33_ASAP7_75t_R g94 ( 
.A(n_65),
.Y(n_94)
);

CKINVDCx5p33_ASAP7_75t_R g95 ( 
.A(n_44),
.Y(n_95)
);

INVxp67_ASAP7_75t_SL g96 ( 
.A(n_1),
.Y(n_96)
);

CKINVDCx5p33_ASAP7_75t_R g97 ( 
.A(n_39),
.Y(n_97)
);

BUFx10_ASAP7_75t_L g98 ( 
.A(n_6),
.Y(n_98)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_19),
.Y(n_99)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_20),
.Y(n_100)
);

BUFx2_ASAP7_75t_L g101 ( 
.A(n_31),
.Y(n_101)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_11),
.Y(n_102)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_64),
.Y(n_103)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_18),
.Y(n_104)
);

HB1xp67_ASAP7_75t_L g105 ( 
.A(n_17),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_36),
.Y(n_106)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_18),
.Y(n_107)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_23),
.Y(n_108)
);

CKINVDCx5p33_ASAP7_75t_R g109 ( 
.A(n_20),
.Y(n_109)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_44),
.Y(n_110)
);

CKINVDCx5p33_ASAP7_75t_R g111 ( 
.A(n_12),
.Y(n_111)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_62),
.Y(n_112)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_30),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_0),
.Y(n_114)
);

CKINVDCx5p33_ASAP7_75t_R g115 ( 
.A(n_46),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_33),
.Y(n_116)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_19),
.Y(n_117)
);

CKINVDCx5p33_ASAP7_75t_R g118 ( 
.A(n_52),
.Y(n_118)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_43),
.Y(n_119)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_43),
.Y(n_120)
);

CKINVDCx5p33_ASAP7_75t_R g121 ( 
.A(n_24),
.Y(n_121)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_47),
.Y(n_122)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_35),
.Y(n_123)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_24),
.Y(n_124)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_5),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_10),
.Y(n_126)
);

CKINVDCx5p33_ASAP7_75t_R g127 ( 
.A(n_35),
.Y(n_127)
);

CKINVDCx5p33_ASAP7_75t_R g128 ( 
.A(n_34),
.Y(n_128)
);

CKINVDCx5p33_ASAP7_75t_R g129 ( 
.A(n_53),
.Y(n_129)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_73),
.Y(n_130)
);

CKINVDCx5p33_ASAP7_75t_R g131 ( 
.A(n_76),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_73),
.Y(n_132)
);

CKINVDCx5p33_ASAP7_75t_R g133 ( 
.A(n_76),
.Y(n_133)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_73),
.Y(n_134)
);

INVxp67_ASAP7_75t_SL g135 ( 
.A(n_102),
.Y(n_135)
);

INVxp67_ASAP7_75t_SL g136 ( 
.A(n_102),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_102),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_119),
.Y(n_138)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_119),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_119),
.Y(n_140)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_106),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_116),
.Y(n_142)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_106),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_106),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_106),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_106),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_106),
.Y(n_147)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_106),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_114),
.Y(n_149)
);

BUFx3_ASAP7_75t_L g150 ( 
.A(n_103),
.Y(n_150)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_141),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g152 ( 
.A(n_141),
.Y(n_152)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_141),
.Y(n_153)
);

CKINVDCx6p67_ASAP7_75t_R g154 ( 
.A(n_150),
.Y(n_154)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_141),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_135),
.A2(n_92),
.B1(n_116),
.B2(n_101),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_143),
.Y(n_157)
);

OAI22x1_ASAP7_75t_L g158 ( 
.A1(n_135),
.A2(n_96),
.B1(n_101),
.B2(n_105),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_150),
.B(n_137),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_143),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_143),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_144),
.Y(n_162)
);

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_131),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g164 ( 
.A(n_141),
.Y(n_164)
);

AOI22x1_ASAP7_75t_SL g165 ( 
.A1(n_142),
.A2(n_96),
.B1(n_80),
.B2(n_79),
.Y(n_165)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_148),
.Y(n_166)
);

AND2x2_ASAP7_75t_SL g167 ( 
.A(n_148),
.B(n_114),
.Y(n_167)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_148),
.Y(n_168)
);

AND2x4_ASAP7_75t_L g169 ( 
.A(n_150),
.B(n_135),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_150),
.B(n_103),
.Y(n_170)
);

BUFx6f_ASAP7_75t_L g171 ( 
.A(n_148),
.Y(n_171)
);

BUFx6f_ASAP7_75t_L g172 ( 
.A(n_148),
.Y(n_172)
);

OA21x2_ASAP7_75t_L g173 ( 
.A1(n_137),
.A2(n_112),
.B(n_104),
.Y(n_173)
);

AND2x4_ASAP7_75t_L g174 ( 
.A(n_150),
.B(n_114),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_144),
.Y(n_175)
);

INVx2_ASAP7_75t_SL g176 ( 
.A(n_144),
.Y(n_176)
);

INVx2_ASAP7_75t_SL g177 ( 
.A(n_145),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_L g178 ( 
.A(n_142),
.B(n_105),
.Y(n_178)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_145),
.Y(n_179)
);

OAI21x1_ASAP7_75t_L g180 ( 
.A1(n_145),
.A2(n_112),
.B(n_104),
.Y(n_180)
);

INVx4_ASAP7_75t_L g181 ( 
.A(n_137),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_146),
.Y(n_182)
);

HB1xp67_ASAP7_75t_L g183 ( 
.A(n_131),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_133),
.B(n_114),
.Y(n_184)
);

HB1xp67_ASAP7_75t_L g185 ( 
.A(n_133),
.Y(n_185)
);

INVx6_ASAP7_75t_L g186 ( 
.A(n_174),
.Y(n_186)
);

NAND2xp33_ASAP7_75t_R g187 ( 
.A(n_163),
.B(n_101),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_157),
.Y(n_188)
);

INVxp67_ASAP7_75t_L g189 ( 
.A(n_183),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_163),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_163),
.Y(n_191)
);

INVxp67_ASAP7_75t_L g192 ( 
.A(n_183),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_157),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_178),
.Y(n_194)
);

INVxp67_ASAP7_75t_SL g195 ( 
.A(n_170),
.Y(n_195)
);

BUFx2_ASAP7_75t_L g196 ( 
.A(n_183),
.Y(n_196)
);

HB1xp67_ASAP7_75t_L g197 ( 
.A(n_169),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_178),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_157),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_157),
.Y(n_200)
);

OR2x2_ASAP7_75t_L g201 ( 
.A(n_156),
.B(n_92),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_178),
.Y(n_202)
);

BUFx2_ASAP7_75t_L g203 ( 
.A(n_185),
.Y(n_203)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_179),
.Y(n_204)
);

HB1xp67_ASAP7_75t_L g205 ( 
.A(n_169),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_178),
.Y(n_206)
);

BUFx10_ASAP7_75t_L g207 ( 
.A(n_169),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_160),
.Y(n_208)
);

INVx1_ASAP7_75t_SL g209 ( 
.A(n_185),
.Y(n_209)
);

BUFx3_ASAP7_75t_L g210 ( 
.A(n_154),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_178),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_160),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_160),
.Y(n_213)
);

CKINVDCx16_ASAP7_75t_R g214 ( 
.A(n_185),
.Y(n_214)
);

INVx3_ASAP7_75t_L g215 ( 
.A(n_181),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_156),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_156),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g218 ( 
.A(n_156),
.B(n_75),
.Y(n_218)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_179),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_160),
.Y(n_220)
);

BUFx10_ASAP7_75t_L g221 ( 
.A(n_169),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_165),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_165),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_165),
.Y(n_224)
);

NAND2xp33_ASAP7_75t_R g225 ( 
.A(n_165),
.B(n_75),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_158),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_158),
.Y(n_227)
);

BUFx2_ASAP7_75t_L g228 ( 
.A(n_158),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_158),
.Y(n_229)
);

CKINVDCx16_ASAP7_75t_R g230 ( 
.A(n_169),
.Y(n_230)
);

INVx2_ASAP7_75t_SL g231 ( 
.A(n_154),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_158),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_158),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_161),
.Y(n_234)
);

INVx3_ASAP7_75t_L g235 ( 
.A(n_181),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_169),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_169),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_R g238 ( 
.A(n_154),
.B(n_170),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_169),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_R g240 ( 
.A(n_154),
.B(n_78),
.Y(n_240)
);

AND2x4_ASAP7_75t_L g241 ( 
.A(n_169),
.B(n_136),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_169),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_170),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_170),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_159),
.B(n_136),
.Y(n_245)
);

BUFx10_ASAP7_75t_L g246 ( 
.A(n_167),
.Y(n_246)
);

INVx4_ASAP7_75t_L g247 ( 
.A(n_154),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_159),
.B(n_136),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_181),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_181),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_181),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_181),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_181),
.Y(n_253)
);

OR2x2_ASAP7_75t_L g254 ( 
.A(n_159),
.B(n_79),
.Y(n_254)
);

BUFx6f_ASAP7_75t_L g255 ( 
.A(n_152),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_161),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_181),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_181),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_159),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_174),
.Y(n_260)
);

NAND2xp33_ASAP7_75t_R g261 ( 
.A(n_173),
.B(n_80),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_174),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_174),
.Y(n_263)
);

AO21x2_ASAP7_75t_L g264 ( 
.A1(n_184),
.A2(n_149),
.B(n_147),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_174),
.Y(n_265)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_179),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_188),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_188),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_193),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_193),
.Y(n_270)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_204),
.Y(n_271)
);

INVx1_ASAP7_75t_SL g272 ( 
.A(n_209),
.Y(n_272)
);

BUFx2_ASAP7_75t_L g273 ( 
.A(n_230),
.Y(n_273)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_204),
.Y(n_274)
);

AND2x6_ASAP7_75t_L g275 ( 
.A(n_210),
.B(n_174),
.Y(n_275)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_204),
.Y(n_276)
);

BUFx2_ASAP7_75t_L g277 ( 
.A(n_230),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_199),
.Y(n_278)
);

BUFx2_ASAP7_75t_L g279 ( 
.A(n_196),
.Y(n_279)
);

OAI22xp33_ASAP7_75t_SL g280 ( 
.A1(n_216),
.A2(n_184),
.B1(n_77),
.B2(n_72),
.Y(n_280)
);

INVx3_ASAP7_75t_L g281 ( 
.A(n_246),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_243),
.B(n_167),
.Y(n_282)
);

BUFx3_ASAP7_75t_L g283 ( 
.A(n_207),
.Y(n_283)
);

INVx3_ASAP7_75t_L g284 ( 
.A(n_246),
.Y(n_284)
);

OAI22xp33_ASAP7_75t_L g285 ( 
.A1(n_187),
.A2(n_72),
.B1(n_77),
.B2(n_108),
.Y(n_285)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_219),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_199),
.Y(n_287)
);

AND2x4_ASAP7_75t_L g288 ( 
.A(n_197),
.B(n_174),
.Y(n_288)
);

BUFx6f_ASAP7_75t_L g289 ( 
.A(n_210),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_191),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_200),
.Y(n_291)
);

INVx2_ASAP7_75t_L g292 ( 
.A(n_219),
.Y(n_292)
);

INVx4_ASAP7_75t_L g293 ( 
.A(n_247),
.Y(n_293)
);

BUFx6f_ASAP7_75t_L g294 ( 
.A(n_210),
.Y(n_294)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_219),
.Y(n_295)
);

INVx2_ASAP7_75t_L g296 ( 
.A(n_266),
.Y(n_296)
);

AND2x4_ASAP7_75t_L g297 ( 
.A(n_197),
.B(n_174),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_200),
.Y(n_298)
);

INVx3_ASAP7_75t_L g299 ( 
.A(n_246),
.Y(n_299)
);

AND2x4_ASAP7_75t_L g300 ( 
.A(n_205),
.B(n_174),
.Y(n_300)
);

BUFx2_ASAP7_75t_L g301 ( 
.A(n_196),
.Y(n_301)
);

INVx1_ASAP7_75t_SL g302 ( 
.A(n_209),
.Y(n_302)
);

BUFx4f_ASAP7_75t_L g303 ( 
.A(n_231),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_208),
.Y(n_304)
);

BUFx3_ASAP7_75t_L g305 ( 
.A(n_207),
.Y(n_305)
);

INVx1_ASAP7_75t_SL g306 ( 
.A(n_203),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_208),
.Y(n_307)
);

AND2x2_ASAP7_75t_L g308 ( 
.A(n_205),
.B(n_167),
.Y(n_308)
);

INVx2_ASAP7_75t_L g309 ( 
.A(n_266),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_189),
.B(n_167),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_244),
.B(n_167),
.Y(n_311)
);

AND2x2_ASAP7_75t_L g312 ( 
.A(n_241),
.B(n_167),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_212),
.Y(n_313)
);

INVx2_ASAP7_75t_L g314 ( 
.A(n_266),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_213),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_189),
.B(n_192),
.Y(n_316)
);

AND2x4_ASAP7_75t_L g317 ( 
.A(n_241),
.B(n_228),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_213),
.Y(n_318)
);

INVx2_ASAP7_75t_L g319 ( 
.A(n_220),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_220),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_192),
.B(n_67),
.Y(n_321)
);

BUFx6f_ASAP7_75t_L g322 ( 
.A(n_247),
.Y(n_322)
);

INVx4_ASAP7_75t_L g323 ( 
.A(n_247),
.Y(n_323)
);

AOI22xp33_ASAP7_75t_L g324 ( 
.A1(n_228),
.A2(n_173),
.B1(n_98),
.B2(n_82),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_234),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_234),
.Y(n_326)
);

BUFx6f_ASAP7_75t_L g327 ( 
.A(n_246),
.Y(n_327)
);

INVx2_ASAP7_75t_L g328 ( 
.A(n_256),
.Y(n_328)
);

AND2x4_ASAP7_75t_L g329 ( 
.A(n_241),
.B(n_174),
.Y(n_329)
);

HB1xp67_ASAP7_75t_L g330 ( 
.A(n_214),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_190),
.Y(n_331)
);

AOI22xp33_ASAP7_75t_L g332 ( 
.A1(n_217),
.A2(n_201),
.B1(n_218),
.B2(n_227),
.Y(n_332)
);

AND2x4_ASAP7_75t_L g333 ( 
.A(n_241),
.B(n_180),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_259),
.B(n_68),
.Y(n_334)
);

INVx3_ASAP7_75t_L g335 ( 
.A(n_215),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_215),
.Y(n_336)
);

INVx2_ASAP7_75t_L g337 ( 
.A(n_215),
.Y(n_337)
);

AND2x4_ASAP7_75t_L g338 ( 
.A(n_236),
.B(n_180),
.Y(n_338)
);

INVx4_ASAP7_75t_L g339 ( 
.A(n_207),
.Y(n_339)
);

AND2x4_ASAP7_75t_L g340 ( 
.A(n_237),
.B(n_180),
.Y(n_340)
);

BUFx6f_ASAP7_75t_L g341 ( 
.A(n_255),
.Y(n_341)
);

INVx3_ASAP7_75t_L g342 ( 
.A(n_215),
.Y(n_342)
);

INVx4_ASAP7_75t_L g343 ( 
.A(n_207),
.Y(n_343)
);

AND2x4_ASAP7_75t_L g344 ( 
.A(n_239),
.B(n_180),
.Y(n_344)
);

INVx1_ASAP7_75t_SL g345 ( 
.A(n_203),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_195),
.B(n_173),
.Y(n_346)
);

INVx2_ASAP7_75t_L g347 ( 
.A(n_235),
.Y(n_347)
);

INVx2_ASAP7_75t_L g348 ( 
.A(n_235),
.Y(n_348)
);

INVx2_ASAP7_75t_L g349 ( 
.A(n_235),
.Y(n_349)
);

AND2x4_ASAP7_75t_L g350 ( 
.A(n_242),
.B(n_180),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_235),
.Y(n_351)
);

INVx2_ASAP7_75t_L g352 ( 
.A(n_186),
.Y(n_352)
);

NOR2xp33_ASAP7_75t_L g353 ( 
.A(n_254),
.B(n_214),
.Y(n_353)
);

AND2x6_ASAP7_75t_L g354 ( 
.A(n_238),
.B(n_153),
.Y(n_354)
);

AND2x6_ASAP7_75t_L g355 ( 
.A(n_255),
.B(n_153),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_221),
.Y(n_356)
);

NOR2x1p5_ASAP7_75t_L g357 ( 
.A(n_201),
.B(n_66),
.Y(n_357)
);

INVx4_ASAP7_75t_SL g358 ( 
.A(n_186),
.Y(n_358)
);

INVx2_ASAP7_75t_L g359 ( 
.A(n_186),
.Y(n_359)
);

INVx3_ASAP7_75t_L g360 ( 
.A(n_221),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_221),
.Y(n_361)
);

INVx2_ASAP7_75t_L g362 ( 
.A(n_186),
.Y(n_362)
);

BUFx6f_ASAP7_75t_L g363 ( 
.A(n_255),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_221),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_186),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_195),
.Y(n_366)
);

INVx2_ASAP7_75t_SL g367 ( 
.A(n_249),
.Y(n_367)
);

NAND2xp33_ASAP7_75t_SL g368 ( 
.A(n_240),
.B(n_72),
.Y(n_368)
);

INVx2_ASAP7_75t_L g369 ( 
.A(n_255),
.Y(n_369)
);

AOI22xp33_ASAP7_75t_L g370 ( 
.A1(n_218),
.A2(n_173),
.B1(n_82),
.B2(n_98),
.Y(n_370)
);

INVx2_ASAP7_75t_L g371 ( 
.A(n_255),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_245),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_245),
.Y(n_373)
);

INVxp67_ASAP7_75t_SL g374 ( 
.A(n_261),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_248),
.Y(n_375)
);

NAND2xp33_ASAP7_75t_L g376 ( 
.A(n_250),
.B(n_176),
.Y(n_376)
);

INVxp67_ASAP7_75t_L g377 ( 
.A(n_187),
.Y(n_377)
);

INVx2_ASAP7_75t_L g378 ( 
.A(n_255),
.Y(n_378)
);

AND2x4_ASAP7_75t_L g379 ( 
.A(n_260),
.B(n_180),
.Y(n_379)
);

NOR2xp33_ASAP7_75t_L g380 ( 
.A(n_254),
.B(n_69),
.Y(n_380)
);

AND2x2_ASAP7_75t_SL g381 ( 
.A(n_261),
.B(n_173),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_SL g382 ( 
.A(n_251),
.B(n_81),
.Y(n_382)
);

INVx2_ASAP7_75t_L g383 ( 
.A(n_264),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_248),
.Y(n_384)
);

INVx2_ASAP7_75t_L g385 ( 
.A(n_264),
.Y(n_385)
);

INVx2_ASAP7_75t_L g386 ( 
.A(n_264),
.Y(n_386)
);

INVx1_ASAP7_75t_SL g387 ( 
.A(n_194),
.Y(n_387)
);

INVxp67_ASAP7_75t_SL g388 ( 
.A(n_225),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_264),
.Y(n_389)
);

AND2x4_ASAP7_75t_L g390 ( 
.A(n_262),
.B(n_66),
.Y(n_390)
);

HB1xp67_ASAP7_75t_L g391 ( 
.A(n_263),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_252),
.Y(n_392)
);

AND2x4_ASAP7_75t_L g393 ( 
.A(n_265),
.B(n_85),
.Y(n_393)
);

AND2x2_ASAP7_75t_L g394 ( 
.A(n_226),
.B(n_173),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_253),
.Y(n_395)
);

INVx2_ASAP7_75t_L g396 ( 
.A(n_257),
.Y(n_396)
);

BUFx10_ASAP7_75t_L g397 ( 
.A(n_258),
.Y(n_397)
);

NAND2xp33_ASAP7_75t_SL g398 ( 
.A(n_229),
.B(n_77),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g399 ( 
.A(n_232),
.B(n_173),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_233),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_198),
.B(n_173),
.Y(n_401)
);

BUFx3_ASAP7_75t_L g402 ( 
.A(n_222),
.Y(n_402)
);

AND2x6_ASAP7_75t_L g403 ( 
.A(n_225),
.B(n_153),
.Y(n_403)
);

NAND3xp33_ASAP7_75t_L g404 ( 
.A(n_223),
.B(n_182),
.C(n_162),
.Y(n_404)
);

INVx2_ASAP7_75t_SL g405 ( 
.A(n_224),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_SL g406 ( 
.A(n_202),
.B(n_82),
.Y(n_406)
);

AOI22xp5_ASAP7_75t_L g407 ( 
.A1(n_206),
.A2(n_173),
.B1(n_97),
.B2(n_95),
.Y(n_407)
);

INVx2_ASAP7_75t_L g408 ( 
.A(n_211),
.Y(n_408)
);

INVx4_ASAP7_75t_L g409 ( 
.A(n_247),
.Y(n_409)
);

BUFx2_ASAP7_75t_L g410 ( 
.A(n_230),
.Y(n_410)
);

AND2x2_ASAP7_75t_L g411 ( 
.A(n_272),
.B(n_173),
.Y(n_411)
);

NOR3xp33_ASAP7_75t_L g412 ( 
.A(n_353),
.B(n_90),
.C(n_85),
.Y(n_412)
);

HB1xp67_ASAP7_75t_L g413 ( 
.A(n_317),
.Y(n_413)
);

INVx2_ASAP7_75t_L g414 ( 
.A(n_271),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_317),
.Y(n_415)
);

INVx2_ASAP7_75t_L g416 ( 
.A(n_271),
.Y(n_416)
);

INVx2_ASAP7_75t_L g417 ( 
.A(n_271),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_317),
.Y(n_418)
);

AOI22xp5_ASAP7_75t_L g419 ( 
.A1(n_317),
.A2(n_91),
.B1(n_74),
.B2(n_128),
.Y(n_419)
);

AO22x2_ASAP7_75t_L g420 ( 
.A1(n_374),
.A2(n_90),
.B1(n_87),
.B2(n_99),
.Y(n_420)
);

OAI22xp33_ASAP7_75t_L g421 ( 
.A1(n_407),
.A2(n_87),
.B1(n_99),
.B2(n_100),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_290),
.Y(n_422)
);

NAND2x1p5_ASAP7_75t_L g423 ( 
.A(n_283),
.B(n_130),
.Y(n_423)
);

A2O1A1Ixp33_ASAP7_75t_L g424 ( 
.A1(n_310),
.A2(n_100),
.B(n_107),
.C(n_108),
.Y(n_424)
);

INVxp67_ASAP7_75t_L g425 ( 
.A(n_272),
.Y(n_425)
);

BUFx8_ASAP7_75t_L g426 ( 
.A(n_279),
.Y(n_426)
);

AND2x4_ASAP7_75t_L g427 ( 
.A(n_358),
.B(n_329),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_329),
.Y(n_428)
);

INVxp67_ASAP7_75t_L g429 ( 
.A(n_302),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_329),
.Y(n_430)
);

BUFx6f_ASAP7_75t_L g431 ( 
.A(n_341),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_329),
.Y(n_432)
);

AO22x2_ASAP7_75t_L g433 ( 
.A1(n_400),
.A2(n_122),
.B1(n_107),
.B2(n_110),
.Y(n_433)
);

CKINVDCx16_ASAP7_75t_R g434 ( 
.A(n_330),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_316),
.B(n_110),
.Y(n_435)
);

INVxp67_ASAP7_75t_L g436 ( 
.A(n_302),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_267),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_267),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_268),
.Y(n_439)
);

INVx2_ASAP7_75t_L g440 ( 
.A(n_274),
.Y(n_440)
);

INVx2_ASAP7_75t_L g441 ( 
.A(n_274),
.Y(n_441)
);

INVxp67_ASAP7_75t_SL g442 ( 
.A(n_333),
.Y(n_442)
);

INVx4_ASAP7_75t_L g443 ( 
.A(n_358),
.Y(n_443)
);

AND2x4_ASAP7_75t_L g444 ( 
.A(n_358),
.B(n_113),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_269),
.Y(n_445)
);

AND2x2_ASAP7_75t_L g446 ( 
.A(n_306),
.B(n_82),
.Y(n_446)
);

AOI22xp5_ASAP7_75t_L g447 ( 
.A1(n_380),
.A2(n_88),
.B1(n_70),
.B2(n_127),
.Y(n_447)
);

INVxp67_ASAP7_75t_L g448 ( 
.A(n_279),
.Y(n_448)
);

INVx2_ASAP7_75t_L g449 ( 
.A(n_274),
.Y(n_449)
);

INVxp67_ASAP7_75t_L g450 ( 
.A(n_301),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_270),
.Y(n_451)
);

INVxp67_ASAP7_75t_L g452 ( 
.A(n_301),
.Y(n_452)
);

INVx2_ASAP7_75t_L g453 ( 
.A(n_276),
.Y(n_453)
);

AOI22xp33_ASAP7_75t_L g454 ( 
.A1(n_381),
.A2(n_82),
.B1(n_98),
.B2(n_113),
.Y(n_454)
);

INVxp67_ASAP7_75t_L g455 ( 
.A(n_306),
.Y(n_455)
);

BUFx6f_ASAP7_75t_L g456 ( 
.A(n_341),
.Y(n_456)
);

INVx4_ASAP7_75t_L g457 ( 
.A(n_358),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_366),
.B(n_117),
.Y(n_458)
);

INVx2_ASAP7_75t_L g459 ( 
.A(n_276),
.Y(n_459)
);

CKINVDCx5p33_ASAP7_75t_R g460 ( 
.A(n_331),
.Y(n_460)
);

AND2x2_ASAP7_75t_L g461 ( 
.A(n_345),
.B(n_98),
.Y(n_461)
);

INVx2_ASAP7_75t_L g462 ( 
.A(n_276),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_278),
.Y(n_463)
);

INVx2_ASAP7_75t_L g464 ( 
.A(n_286),
.Y(n_464)
);

BUFx4f_ASAP7_75t_L g465 ( 
.A(n_288),
.Y(n_465)
);

OR2x2_ASAP7_75t_L g466 ( 
.A(n_345),
.B(n_130),
.Y(n_466)
);

NAND2x1p5_ASAP7_75t_L g467 ( 
.A(n_283),
.B(n_130),
.Y(n_467)
);

NOR2xp33_ASAP7_75t_L g468 ( 
.A(n_377),
.B(n_83),
.Y(n_468)
);

INVx3_ASAP7_75t_L g469 ( 
.A(n_339),
.Y(n_469)
);

BUFx8_ASAP7_75t_L g470 ( 
.A(n_408),
.Y(n_470)
);

NAND2x1p5_ASAP7_75t_L g471 ( 
.A(n_283),
.B(n_132),
.Y(n_471)
);

INVx2_ASAP7_75t_L g472 ( 
.A(n_286),
.Y(n_472)
);

NAND2xp33_ASAP7_75t_L g473 ( 
.A(n_322),
.B(n_176),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_287),
.Y(n_474)
);

BUFx8_ASAP7_75t_L g475 ( 
.A(n_408),
.Y(n_475)
);

AOI22xp33_ASAP7_75t_L g476 ( 
.A1(n_381),
.A2(n_98),
.B1(n_122),
.B2(n_117),
.Y(n_476)
);

INVxp67_ASAP7_75t_L g477 ( 
.A(n_273),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_287),
.Y(n_478)
);

INVx2_ASAP7_75t_L g479 ( 
.A(n_286),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_291),
.Y(n_480)
);

AO22x2_ASAP7_75t_L g481 ( 
.A1(n_400),
.A2(n_120),
.B1(n_123),
.B2(n_124),
.Y(n_481)
);

AND2x2_ASAP7_75t_L g482 ( 
.A(n_387),
.B(n_132),
.Y(n_482)
);

INVx2_ASAP7_75t_L g483 ( 
.A(n_292),
.Y(n_483)
);

NAND2x1p5_ASAP7_75t_L g484 ( 
.A(n_305),
.B(n_132),
.Y(n_484)
);

INVxp67_ASAP7_75t_L g485 ( 
.A(n_273),
.Y(n_485)
);

INVx4_ASAP7_75t_L g486 ( 
.A(n_358),
.Y(n_486)
);

NOR2xp33_ASAP7_75t_L g487 ( 
.A(n_401),
.B(n_84),
.Y(n_487)
);

NOR2x1p5_ASAP7_75t_L g488 ( 
.A(n_408),
.B(n_120),
.Y(n_488)
);

OR2x2_ASAP7_75t_L g489 ( 
.A(n_387),
.B(n_134),
.Y(n_489)
);

NAND2x1p5_ASAP7_75t_L g490 ( 
.A(n_305),
.B(n_134),
.Y(n_490)
);

AOI22xp5_ASAP7_75t_L g491 ( 
.A1(n_407),
.A2(n_115),
.B1(n_89),
.B2(n_93),
.Y(n_491)
);

INVx2_ASAP7_75t_L g492 ( 
.A(n_292),
.Y(n_492)
);

AND2x2_ASAP7_75t_L g493 ( 
.A(n_357),
.B(n_134),
.Y(n_493)
);

AO22x2_ASAP7_75t_L g494 ( 
.A1(n_394),
.A2(n_123),
.B1(n_124),
.B2(n_125),
.Y(n_494)
);

AOI22xp5_ASAP7_75t_L g495 ( 
.A1(n_312),
.A2(n_111),
.B1(n_86),
.B2(n_121),
.Y(n_495)
);

INVxp67_ASAP7_75t_L g496 ( 
.A(n_277),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_L g497 ( 
.A(n_372),
.B(n_125),
.Y(n_497)
);

INVx2_ASAP7_75t_SL g498 ( 
.A(n_402),
.Y(n_498)
);

BUFx6f_ASAP7_75t_L g499 ( 
.A(n_341),
.Y(n_499)
);

NOR2xp33_ASAP7_75t_L g500 ( 
.A(n_277),
.B(n_109),
.Y(n_500)
);

AOI22xp5_ASAP7_75t_L g501 ( 
.A1(n_312),
.A2(n_71),
.B1(n_94),
.B2(n_118),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_L g502 ( 
.A(n_373),
.B(n_161),
.Y(n_502)
);

INVx2_ASAP7_75t_L g503 ( 
.A(n_292),
.Y(n_503)
);

INVx2_ASAP7_75t_L g504 ( 
.A(n_295),
.Y(n_504)
);

CKINVDCx5p33_ASAP7_75t_R g505 ( 
.A(n_402),
.Y(n_505)
);

INVx1_ASAP7_75t_SL g506 ( 
.A(n_410),
.Y(n_506)
);

INVx2_ASAP7_75t_SL g507 ( 
.A(n_402),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_298),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_298),
.Y(n_509)
);

AO22x2_ASAP7_75t_L g510 ( 
.A1(n_394),
.A2(n_332),
.B1(n_399),
.B2(n_404),
.Y(n_510)
);

AO22x2_ASAP7_75t_L g511 ( 
.A1(n_404),
.A2(n_140),
.B1(n_138),
.B2(n_139),
.Y(n_511)
);

AO22x2_ASAP7_75t_L g512 ( 
.A1(n_389),
.A2(n_140),
.B1(n_138),
.B2(n_139),
.Y(n_512)
);

AND2x4_ASAP7_75t_L g513 ( 
.A(n_305),
.B(n_138),
.Y(n_513)
);

AOI22xp5_ASAP7_75t_L g514 ( 
.A1(n_356),
.A2(n_129),
.B1(n_182),
.B2(n_162),
.Y(n_514)
);

CKINVDCx5p33_ASAP7_75t_R g515 ( 
.A(n_405),
.Y(n_515)
);

AND2x2_ASAP7_75t_L g516 ( 
.A(n_357),
.B(n_139),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_304),
.Y(n_517)
);

AO22x2_ASAP7_75t_L g518 ( 
.A1(n_389),
.A2(n_140),
.B1(n_137),
.B2(n_175),
.Y(n_518)
);

AOI22xp5_ASAP7_75t_L g519 ( 
.A1(n_356),
.A2(n_182),
.B1(n_162),
.B2(n_175),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_304),
.Y(n_520)
);

AO22x2_ASAP7_75t_L g521 ( 
.A1(n_383),
.A2(n_182),
.B1(n_175),
.B2(n_162),
.Y(n_521)
);

AOI22xp5_ASAP7_75t_L g522 ( 
.A1(n_361),
.A2(n_175),
.B1(n_177),
.B2(n_176),
.Y(n_522)
);

AO22x2_ASAP7_75t_L g523 ( 
.A1(n_383),
.A2(n_179),
.B1(n_2),
.B2(n_3),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_307),
.Y(n_524)
);

INVx2_ASAP7_75t_SL g525 ( 
.A(n_405),
.Y(n_525)
);

INVx2_ASAP7_75t_L g526 ( 
.A(n_295),
.Y(n_526)
);

BUFx2_ASAP7_75t_L g527 ( 
.A(n_410),
.Y(n_527)
);

AND2x4_ASAP7_75t_L g528 ( 
.A(n_288),
.B(n_179),
.Y(n_528)
);

AO22x2_ASAP7_75t_L g529 ( 
.A1(n_383),
.A2(n_179),
.B1(n_2),
.B2(n_4),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_307),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_L g531 ( 
.A(n_373),
.B(n_177),
.Y(n_531)
);

NOR2xp33_ASAP7_75t_L g532 ( 
.A(n_365),
.B(n_177),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_313),
.Y(n_533)
);

CKINVDCx5p33_ASAP7_75t_R g534 ( 
.A(n_388),
.Y(n_534)
);

NAND2x1p5_ASAP7_75t_L g535 ( 
.A(n_339),
.B(n_151),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_313),
.Y(n_536)
);

AND2x4_ASAP7_75t_L g537 ( 
.A(n_288),
.B(n_155),
.Y(n_537)
);

INVx2_ASAP7_75t_L g538 ( 
.A(n_296),
.Y(n_538)
);

BUFx2_ASAP7_75t_L g539 ( 
.A(n_391),
.Y(n_539)
);

INVx2_ASAP7_75t_L g540 ( 
.A(n_296),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_315),
.Y(n_541)
);

OAI22xp5_ASAP7_75t_L g542 ( 
.A1(n_333),
.A2(n_177),
.B1(n_176),
.B2(n_114),
.Y(n_542)
);

AND2x2_ASAP7_75t_L g543 ( 
.A(n_321),
.B(n_390),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_315),
.Y(n_544)
);

OAI221xp5_ASAP7_75t_L g545 ( 
.A1(n_370),
.A2(n_114),
.B1(n_126),
.B2(n_177),
.C(n_176),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_318),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_318),
.Y(n_547)
);

INVx2_ASAP7_75t_L g548 ( 
.A(n_296),
.Y(n_548)
);

AND2x4_ASAP7_75t_L g549 ( 
.A(n_288),
.B(n_168),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_SL g550 ( 
.A(n_322),
.B(n_333),
.Y(n_550)
);

AND2x4_ASAP7_75t_L g551 ( 
.A(n_297),
.B(n_300),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_320),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_320),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_325),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_L g555 ( 
.A(n_375),
.B(n_177),
.Y(n_555)
);

AND2x6_ASAP7_75t_L g556 ( 
.A(n_333),
.B(n_155),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_326),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_326),
.Y(n_558)
);

BUFx8_ASAP7_75t_L g559 ( 
.A(n_390),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_319),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_319),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_319),
.Y(n_562)
);

AND2x2_ASAP7_75t_L g563 ( 
.A(n_390),
.B(n_168),
.Y(n_563)
);

AND2x2_ASAP7_75t_L g564 ( 
.A(n_390),
.B(n_168),
.Y(n_564)
);

INVxp67_ASAP7_75t_L g565 ( 
.A(n_308),
.Y(n_565)
);

AND2x4_ASAP7_75t_L g566 ( 
.A(n_297),
.B(n_168),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_328),
.Y(n_567)
);

BUFx2_ASAP7_75t_L g568 ( 
.A(n_297),
.Y(n_568)
);

AO22x2_ASAP7_75t_L g569 ( 
.A1(n_385),
.A2(n_0),
.B1(n_4),
.B2(n_5),
.Y(n_569)
);

BUFx2_ASAP7_75t_L g570 ( 
.A(n_426),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_L g571 ( 
.A(n_543),
.B(n_375),
.Y(n_571)
);

NOR2xp33_ASAP7_75t_L g572 ( 
.A(n_448),
.B(n_365),
.Y(n_572)
);

A2O1A1Ixp33_ASAP7_75t_L g573 ( 
.A1(n_442),
.A2(n_487),
.B(n_424),
.C(n_412),
.Y(n_573)
);

AOI22xp5_ASAP7_75t_L g574 ( 
.A1(n_442),
.A2(n_285),
.B1(n_367),
.B2(n_392),
.Y(n_574)
);

NOR2xp33_ASAP7_75t_L g575 ( 
.A(n_448),
.B(n_384),
.Y(n_575)
);

AOI22xp33_ASAP7_75t_L g576 ( 
.A1(n_421),
.A2(n_280),
.B1(n_381),
.B2(n_393),
.Y(n_576)
);

HB1xp67_ASAP7_75t_L g577 ( 
.A(n_413),
.Y(n_577)
);

AOI21xp5_ASAP7_75t_L g578 ( 
.A1(n_473),
.A2(n_303),
.B(n_293),
.Y(n_578)
);

O2A1O1Ixp33_ASAP7_75t_L g579 ( 
.A1(n_435),
.A2(n_395),
.B(n_392),
.C(n_367),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_L g580 ( 
.A(n_565),
.B(n_384),
.Y(n_580)
);

INVx1_ASAP7_75t_SL g581 ( 
.A(n_434),
.Y(n_581)
);

OAI21xp5_ASAP7_75t_L g582 ( 
.A1(n_542),
.A2(n_346),
.B(n_282),
.Y(n_582)
);

NOR2xp33_ASAP7_75t_L g583 ( 
.A(n_450),
.B(n_339),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_L g584 ( 
.A(n_565),
.B(n_482),
.Y(n_584)
);

AOI21xp5_ASAP7_75t_L g585 ( 
.A1(n_550),
.A2(n_303),
.B(n_409),
.Y(n_585)
);

OAI22xp5_ASAP7_75t_L g586 ( 
.A1(n_465),
.A2(n_323),
.B1(n_293),
.B2(n_409),
.Y(n_586)
);

AOI21xp5_ASAP7_75t_L g587 ( 
.A1(n_550),
.A2(n_409),
.B(n_323),
.Y(n_587)
);

AOI21xp5_ASAP7_75t_L g588 ( 
.A1(n_502),
.A2(n_323),
.B(n_293),
.Y(n_588)
);

AOI21xp5_ASAP7_75t_L g589 ( 
.A1(n_531),
.A2(n_323),
.B(n_322),
.Y(n_589)
);

AOI21xp5_ASAP7_75t_L g590 ( 
.A1(n_555),
.A2(n_322),
.B(n_376),
.Y(n_590)
);

AND2x2_ASAP7_75t_L g591 ( 
.A(n_446),
.B(n_393),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_L g592 ( 
.A(n_425),
.B(n_393),
.Y(n_592)
);

NAND2x1p5_ASAP7_75t_L g593 ( 
.A(n_443),
.B(n_339),
.Y(n_593)
);

AOI22xp5_ASAP7_75t_L g594 ( 
.A1(n_455),
.A2(n_361),
.B1(n_364),
.B2(n_368),
.Y(n_594)
);

INVx2_ASAP7_75t_L g595 ( 
.A(n_414),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_SL g596 ( 
.A(n_469),
.B(n_322),
.Y(n_596)
);

INVx11_ASAP7_75t_L g597 ( 
.A(n_426),
.Y(n_597)
);

OAI321xp33_ASAP7_75t_L g598 ( 
.A1(n_454),
.A2(n_324),
.A3(n_406),
.B1(n_311),
.B2(n_396),
.C(n_114),
.Y(n_598)
);

AOI21xp5_ASAP7_75t_L g599 ( 
.A1(n_560),
.A2(n_294),
.B(n_289),
.Y(n_599)
);

INVx2_ASAP7_75t_L g600 ( 
.A(n_414),
.Y(n_600)
);

AND2x4_ASAP7_75t_L g601 ( 
.A(n_551),
.B(n_297),
.Y(n_601)
);

INVx2_ASAP7_75t_L g602 ( 
.A(n_416),
.Y(n_602)
);

INVx2_ASAP7_75t_L g603 ( 
.A(n_416),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_437),
.Y(n_604)
);

O2A1O1Ixp33_ASAP7_75t_L g605 ( 
.A1(n_412),
.A2(n_424),
.B(n_452),
.C(n_450),
.Y(n_605)
);

AOI21xp5_ASAP7_75t_L g606 ( 
.A1(n_561),
.A2(n_294),
.B(n_289),
.Y(n_606)
);

AOI21xp5_ASAP7_75t_L g607 ( 
.A1(n_562),
.A2(n_294),
.B(n_289),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_L g608 ( 
.A(n_425),
.B(n_300),
.Y(n_608)
);

A2O1A1Ixp33_ASAP7_75t_L g609 ( 
.A1(n_487),
.A2(n_340),
.B(n_344),
.C(n_350),
.Y(n_609)
);

AOI21xp5_ASAP7_75t_L g610 ( 
.A1(n_567),
.A2(n_369),
.B(n_371),
.Y(n_610)
);

OR2x2_ASAP7_75t_L g611 ( 
.A(n_452),
.B(n_300),
.Y(n_611)
);

A2O1A1Ixp33_ASAP7_75t_L g612 ( 
.A1(n_476),
.A2(n_340),
.B(n_344),
.C(n_350),
.Y(n_612)
);

NAND3xp33_ASAP7_75t_SL g613 ( 
.A(n_447),
.B(n_398),
.C(n_382),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_L g614 ( 
.A(n_429),
.B(n_436),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_L g615 ( 
.A(n_429),
.B(n_300),
.Y(n_615)
);

INVx2_ASAP7_75t_SL g616 ( 
.A(n_422),
.Y(n_616)
);

AOI21xp5_ASAP7_75t_L g617 ( 
.A1(n_438),
.A2(n_369),
.B(n_371),
.Y(n_617)
);

AOI21xp5_ASAP7_75t_L g618 ( 
.A1(n_439),
.A2(n_369),
.B(n_371),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_SL g619 ( 
.A(n_469),
.B(n_396),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_L g620 ( 
.A(n_436),
.B(n_308),
.Y(n_620)
);

OR2x2_ASAP7_75t_L g621 ( 
.A(n_506),
.B(n_352),
.Y(n_621)
);

AOI21xp5_ASAP7_75t_L g622 ( 
.A1(n_445),
.A2(n_378),
.B(n_341),
.Y(n_622)
);

OAI21xp5_ASAP7_75t_L g623 ( 
.A1(n_532),
.A2(n_336),
.B(n_351),
.Y(n_623)
);

NOR2xp33_ASAP7_75t_L g624 ( 
.A(n_477),
.B(n_343),
.Y(n_624)
);

INVx4_ASAP7_75t_L g625 ( 
.A(n_427),
.Y(n_625)
);

NAND2x1p5_ASAP7_75t_L g626 ( 
.A(n_443),
.B(n_457),
.Y(n_626)
);

INVx4_ASAP7_75t_L g627 ( 
.A(n_427),
.Y(n_627)
);

AOI21xp5_ASAP7_75t_L g628 ( 
.A1(n_451),
.A2(n_341),
.B(n_363),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_L g629 ( 
.A(n_413),
.B(n_352),
.Y(n_629)
);

OAI22xp5_ASAP7_75t_L g630 ( 
.A1(n_465),
.A2(n_343),
.B1(n_396),
.B2(n_338),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_SL g631 ( 
.A(n_431),
.B(n_281),
.Y(n_631)
);

BUFx6f_ASAP7_75t_L g632 ( 
.A(n_431),
.Y(n_632)
);

OAI22xp5_ASAP7_75t_L g633 ( 
.A1(n_463),
.A2(n_343),
.B1(n_344),
.B2(n_340),
.Y(n_633)
);

OAI22xp5_ASAP7_75t_L g634 ( 
.A1(n_474),
.A2(n_338),
.B1(n_350),
.B2(n_340),
.Y(n_634)
);

O2A1O1Ixp33_ASAP7_75t_L g635 ( 
.A1(n_497),
.A2(n_352),
.B(n_362),
.C(n_359),
.Y(n_635)
);

INVx2_ASAP7_75t_L g636 ( 
.A(n_417),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_478),
.Y(n_637)
);

NOR2xp33_ASAP7_75t_L g638 ( 
.A(n_477),
.B(n_359),
.Y(n_638)
);

A2O1A1Ixp33_ASAP7_75t_L g639 ( 
.A1(n_476),
.A2(n_344),
.B(n_338),
.C(n_350),
.Y(n_639)
);

INVx2_ASAP7_75t_L g640 ( 
.A(n_417),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_SL g641 ( 
.A(n_431),
.B(n_281),
.Y(n_641)
);

OAI22xp5_ASAP7_75t_L g642 ( 
.A1(n_480),
.A2(n_338),
.B1(n_360),
.B2(n_379),
.Y(n_642)
);

OR2x2_ASAP7_75t_L g643 ( 
.A(n_466),
.B(n_489),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_SL g644 ( 
.A(n_431),
.B(n_281),
.Y(n_644)
);

CKINVDCx10_ASAP7_75t_R g645 ( 
.A(n_460),
.Y(n_645)
);

AND2x2_ASAP7_75t_L g646 ( 
.A(n_461),
.B(n_527),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_508),
.Y(n_647)
);

NOR2xp33_ASAP7_75t_L g648 ( 
.A(n_485),
.B(n_359),
.Y(n_648)
);

HB1xp67_ASAP7_75t_L g649 ( 
.A(n_551),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_L g650 ( 
.A(n_551),
.B(n_362),
.Y(n_650)
);

OAI21xp5_ASAP7_75t_L g651 ( 
.A1(n_532),
.A2(n_336),
.B(n_351),
.Y(n_651)
);

A2O1A1Ixp33_ASAP7_75t_L g652 ( 
.A1(n_509),
.A2(n_379),
.B(n_337),
.C(n_347),
.Y(n_652)
);

NOR2xp33_ASAP7_75t_SL g653 ( 
.A(n_460),
.B(n_397),
.Y(n_653)
);

AOI21xp5_ASAP7_75t_L g654 ( 
.A1(n_517),
.A2(n_363),
.B(n_379),
.Y(n_654)
);

O2A1O1Ixp33_ASAP7_75t_L g655 ( 
.A1(n_485),
.A2(n_362),
.B(n_360),
.C(n_342),
.Y(n_655)
);

AOI21xp5_ASAP7_75t_L g656 ( 
.A1(n_520),
.A2(n_379),
.B(n_347),
.Y(n_656)
);

AOI21xp5_ASAP7_75t_L g657 ( 
.A1(n_524),
.A2(n_348),
.B(n_349),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_SL g658 ( 
.A(n_456),
.B(n_499),
.Y(n_658)
);

BUFx6f_ASAP7_75t_L g659 ( 
.A(n_456),
.Y(n_659)
);

AOI21xp5_ASAP7_75t_L g660 ( 
.A1(n_530),
.A2(n_347),
.B(n_337),
.Y(n_660)
);

AOI22xp33_ASAP7_75t_L g661 ( 
.A1(n_494),
.A2(n_403),
.B1(n_327),
.B2(n_386),
.Y(n_661)
);

BUFx2_ASAP7_75t_L g662 ( 
.A(n_559),
.Y(n_662)
);

O2A1O1Ixp33_ASAP7_75t_L g663 ( 
.A1(n_496),
.A2(n_360),
.B(n_335),
.C(n_342),
.Y(n_663)
);

INVxp67_ASAP7_75t_L g664 ( 
.A(n_539),
.Y(n_664)
);

AO21x1_ASAP7_75t_L g665 ( 
.A1(n_533),
.A2(n_386),
.B(n_385),
.Y(n_665)
);

CKINVDCx5p33_ASAP7_75t_R g666 ( 
.A(n_422),
.Y(n_666)
);

AOI21xp5_ASAP7_75t_L g667 ( 
.A1(n_536),
.A2(n_349),
.B(n_314),
.Y(n_667)
);

AO22x1_ASAP7_75t_L g668 ( 
.A1(n_559),
.A2(n_403),
.B1(n_275),
.B2(n_327),
.Y(n_668)
);

OAI22xp5_ASAP7_75t_L g669 ( 
.A1(n_541),
.A2(n_342),
.B1(n_335),
.B2(n_284),
.Y(n_669)
);

AOI21x1_ASAP7_75t_L g670 ( 
.A1(n_521),
.A2(n_309),
.B(n_314),
.Y(n_670)
);

OAI22xp5_ASAP7_75t_L g671 ( 
.A1(n_544),
.A2(n_342),
.B1(n_335),
.B2(n_284),
.Y(n_671)
);

OAI22xp5_ASAP7_75t_L g672 ( 
.A1(n_546),
.A2(n_335),
.B1(n_281),
.B2(n_284),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_L g673 ( 
.A(n_493),
.B(n_397),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_547),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_SL g675 ( 
.A(n_456),
.B(n_499),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_552),
.Y(n_676)
);

BUFx4f_ASAP7_75t_L g677 ( 
.A(n_415),
.Y(n_677)
);

AND2x2_ASAP7_75t_L g678 ( 
.A(n_516),
.B(n_397),
.Y(n_678)
);

OAI321xp33_ASAP7_75t_L g679 ( 
.A1(n_454),
.A2(n_126),
.A3(n_309),
.B1(n_314),
.B2(n_166),
.C(n_155),
.Y(n_679)
);

OAI22xp5_ASAP7_75t_L g680 ( 
.A1(n_553),
.A2(n_299),
.B1(n_284),
.B2(n_309),
.Y(n_680)
);

NOR2xp33_ASAP7_75t_L g681 ( 
.A(n_418),
.B(n_299),
.Y(n_681)
);

AOI22xp33_ASAP7_75t_SL g682 ( 
.A1(n_494),
.A2(n_275),
.B1(n_327),
.B2(n_403),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_554),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_568),
.B(n_386),
.Y(n_684)
);

A2O1A1Ixp33_ASAP7_75t_L g685 ( 
.A1(n_557),
.A2(n_299),
.B(n_168),
.C(n_153),
.Y(n_685)
);

INVx2_ASAP7_75t_L g686 ( 
.A(n_440),
.Y(n_686)
);

AOI21xp5_ASAP7_75t_L g687 ( 
.A1(n_558),
.A2(n_327),
.B(n_385),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_SL g688 ( 
.A(n_456),
.B(n_327),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_L g689 ( 
.A(n_411),
.B(n_403),
.Y(n_689)
);

OAI21xp5_ASAP7_75t_L g690 ( 
.A1(n_519),
.A2(n_354),
.B(n_275),
.Y(n_690)
);

AOI21x1_ASAP7_75t_L g691 ( 
.A1(n_521),
.A2(n_149),
.B(n_147),
.Y(n_691)
);

BUFx3_ASAP7_75t_L g692 ( 
.A(n_470),
.Y(n_692)
);

AOI22xp5_ASAP7_75t_L g693 ( 
.A1(n_500),
.A2(n_275),
.B1(n_403),
.B2(n_354),
.Y(n_693)
);

AOI21xp5_ASAP7_75t_L g694 ( 
.A1(n_499),
.A2(n_354),
.B(n_275),
.Y(n_694)
);

AOI21xp5_ASAP7_75t_L g695 ( 
.A1(n_499),
.A2(n_354),
.B(n_153),
.Y(n_695)
);

AOI21xp5_ASAP7_75t_L g696 ( 
.A1(n_440),
.A2(n_354),
.B(n_153),
.Y(n_696)
);

AND2x2_ASAP7_75t_L g697 ( 
.A(n_500),
.B(n_403),
.Y(n_697)
);

O2A1O1Ixp33_ASAP7_75t_L g698 ( 
.A1(n_468),
.A2(n_153),
.B(n_168),
.C(n_166),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_L g699 ( 
.A(n_428),
.B(n_403),
.Y(n_699)
);

AOI22xp5_ASAP7_75t_L g700 ( 
.A1(n_515),
.A2(n_354),
.B1(n_355),
.B2(n_126),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_512),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_512),
.Y(n_702)
);

BUFx2_ASAP7_75t_L g703 ( 
.A(n_470),
.Y(n_703)
);

O2A1O1Ixp33_ASAP7_75t_L g704 ( 
.A1(n_468),
.A2(n_458),
.B(n_513),
.C(n_430),
.Y(n_704)
);

INVx2_ASAP7_75t_L g705 ( 
.A(n_441),
.Y(n_705)
);

AOI21xp5_ASAP7_75t_L g706 ( 
.A1(n_441),
.A2(n_155),
.B(n_168),
.Y(n_706)
);

AOI22xp5_ASAP7_75t_L g707 ( 
.A1(n_515),
.A2(n_355),
.B1(n_126),
.B2(n_151),
.Y(n_707)
);

AOI21xp33_ASAP7_75t_L g708 ( 
.A1(n_545),
.A2(n_151),
.B(n_166),
.Y(n_708)
);

AOI21xp5_ASAP7_75t_L g709 ( 
.A1(n_449),
.A2(n_155),
.B(n_166),
.Y(n_709)
);

O2A1O1Ixp33_ASAP7_75t_L g710 ( 
.A1(n_513),
.A2(n_166),
.B(n_155),
.C(n_151),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_L g711 ( 
.A(n_432),
.B(n_355),
.Y(n_711)
);

INVx2_ASAP7_75t_L g712 ( 
.A(n_453),
.Y(n_712)
);

NOR2xp33_ASAP7_75t_L g713 ( 
.A(n_534),
.B(n_355),
.Y(n_713)
);

AND2x6_ASAP7_75t_L g714 ( 
.A(n_537),
.B(n_151),
.Y(n_714)
);

O2A1O1Ixp33_ASAP7_75t_L g715 ( 
.A1(n_488),
.A2(n_151),
.B(n_149),
.C(n_147),
.Y(n_715)
);

NOR2xp33_ASAP7_75t_L g716 ( 
.A(n_534),
.B(n_355),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_L g717 ( 
.A(n_528),
.B(n_355),
.Y(n_717)
);

INVx2_ASAP7_75t_L g718 ( 
.A(n_453),
.Y(n_718)
);

A2O1A1Ixp33_ASAP7_75t_L g719 ( 
.A1(n_491),
.A2(n_563),
.B(n_564),
.C(n_492),
.Y(n_719)
);

OAI22xp5_ASAP7_75t_L g720 ( 
.A1(n_423),
.A2(n_126),
.B1(n_355),
.B2(n_171),
.Y(n_720)
);

A2O1A1Ixp33_ASAP7_75t_L g721 ( 
.A1(n_459),
.A2(n_126),
.B(n_146),
.C(n_171),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_SL g722 ( 
.A(n_457),
.B(n_172),
.Y(n_722)
);

OAI21xp5_ASAP7_75t_L g723 ( 
.A1(n_522),
.A2(n_355),
.B(n_146),
.Y(n_723)
);

NOR2xp33_ASAP7_75t_L g724 ( 
.A(n_528),
.B(n_7),
.Y(n_724)
);

AOI22xp5_ASAP7_75t_L g725 ( 
.A1(n_505),
.A2(n_172),
.B1(n_171),
.B2(n_164),
.Y(n_725)
);

INVx3_ASAP7_75t_L g726 ( 
.A(n_486),
.Y(n_726)
);

INVx4_ASAP7_75t_L g727 ( 
.A(n_486),
.Y(n_727)
);

NAND3xp33_ASAP7_75t_L g728 ( 
.A(n_475),
.B(n_172),
.C(n_171),
.Y(n_728)
);

OAI21xp5_ASAP7_75t_L g729 ( 
.A1(n_514),
.A2(n_172),
.B(n_171),
.Y(n_729)
);

OAI21x1_ASAP7_75t_L g730 ( 
.A1(n_459),
.A2(n_503),
.B(n_462),
.Y(n_730)
);

AOI21xp5_ASAP7_75t_L g731 ( 
.A1(n_462),
.A2(n_172),
.B(n_171),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_L g732 ( 
.A(n_549),
.B(n_7),
.Y(n_732)
);

AOI22xp5_ASAP7_75t_L g733 ( 
.A1(n_505),
.A2(n_172),
.B1(n_171),
.B2(n_164),
.Y(n_733)
);

AOI21xp5_ASAP7_75t_L g734 ( 
.A1(n_464),
.A2(n_172),
.B(n_171),
.Y(n_734)
);

INVx2_ASAP7_75t_L g735 ( 
.A(n_464),
.Y(n_735)
);

NOR2x1_ASAP7_75t_L g736 ( 
.A(n_444),
.B(n_172),
.Y(n_736)
);

NOR2xp33_ASAP7_75t_L g737 ( 
.A(n_549),
.B(n_9),
.Y(n_737)
);

AOI21xp5_ASAP7_75t_L g738 ( 
.A1(n_472),
.A2(n_172),
.B(n_171),
.Y(n_738)
);

BUFx2_ASAP7_75t_L g739 ( 
.A(n_475),
.Y(n_739)
);

HB1xp67_ASAP7_75t_L g740 ( 
.A(n_537),
.Y(n_740)
);

AOI21xp5_ASAP7_75t_L g741 ( 
.A1(n_472),
.A2(n_172),
.B(n_171),
.Y(n_741)
);

AOI21xp5_ASAP7_75t_L g742 ( 
.A1(n_479),
.A2(n_172),
.B(n_171),
.Y(n_742)
);

INVx2_ASAP7_75t_L g743 ( 
.A(n_479),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_512),
.Y(n_744)
);

OAI22xp5_ASAP7_75t_L g745 ( 
.A1(n_423),
.A2(n_171),
.B1(n_164),
.B2(n_152),
.Y(n_745)
);

BUFx4f_ASAP7_75t_L g746 ( 
.A(n_498),
.Y(n_746)
);

AOI22xp5_ASAP7_75t_L g747 ( 
.A1(n_507),
.A2(n_172),
.B1(n_171),
.B2(n_164),
.Y(n_747)
);

INVx2_ASAP7_75t_L g748 ( 
.A(n_483),
.Y(n_748)
);

AND2x2_ASAP7_75t_L g749 ( 
.A(n_494),
.B(n_10),
.Y(n_749)
);

AOI21xp5_ASAP7_75t_L g750 ( 
.A1(n_483),
.A2(n_172),
.B(n_171),
.Y(n_750)
);

A2O1A1Ixp33_ASAP7_75t_L g751 ( 
.A1(n_504),
.A2(n_172),
.B(n_164),
.C(n_152),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_L g752 ( 
.A(n_566),
.B(n_13),
.Y(n_752)
);

AND2x2_ASAP7_75t_L g753 ( 
.A(n_646),
.B(n_420),
.Y(n_753)
);

NOR2xp33_ASAP7_75t_L g754 ( 
.A(n_649),
.B(n_566),
.Y(n_754)
);

NOR2xp33_ASAP7_75t_L g755 ( 
.A(n_649),
.B(n_537),
.Y(n_755)
);

INVx2_ASAP7_75t_L g756 ( 
.A(n_595),
.Y(n_756)
);

O2A1O1Ixp33_ASAP7_75t_L g757 ( 
.A1(n_573),
.A2(n_525),
.B(n_471),
.C(n_490),
.Y(n_757)
);

AOI21xp5_ASAP7_75t_L g758 ( 
.A1(n_578),
.A2(n_535),
.B(n_521),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_L g759 ( 
.A(n_643),
.B(n_420),
.Y(n_759)
);

O2A1O1Ixp33_ASAP7_75t_L g760 ( 
.A1(n_573),
.A2(n_605),
.B(n_613),
.C(n_579),
.Y(n_760)
);

INVx3_ASAP7_75t_L g761 ( 
.A(n_625),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_604),
.Y(n_762)
);

INVx4_ASAP7_75t_L g763 ( 
.A(n_597),
.Y(n_763)
);

INVx2_ASAP7_75t_L g764 ( 
.A(n_602),
.Y(n_764)
);

INVx1_ASAP7_75t_SL g765 ( 
.A(n_581),
.Y(n_765)
);

A2O1A1Ixp33_ASAP7_75t_L g766 ( 
.A1(n_704),
.A2(n_495),
.B(n_501),
.C(n_419),
.Y(n_766)
);

O2A1O1Ixp33_ASAP7_75t_L g767 ( 
.A1(n_575),
.A2(n_467),
.B(n_484),
.C(n_471),
.Y(n_767)
);

INVx2_ASAP7_75t_L g768 ( 
.A(n_603),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_637),
.Y(n_769)
);

INVx2_ASAP7_75t_SL g770 ( 
.A(n_645),
.Y(n_770)
);

AND2x2_ASAP7_75t_L g771 ( 
.A(n_591),
.B(n_420),
.Y(n_771)
);

HB1xp67_ASAP7_75t_L g772 ( 
.A(n_577),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_647),
.Y(n_773)
);

BUFx12f_ASAP7_75t_L g774 ( 
.A(n_666),
.Y(n_774)
);

INVx2_ASAP7_75t_L g775 ( 
.A(n_636),
.Y(n_775)
);

NAND3xp33_ASAP7_75t_L g776 ( 
.A(n_574),
.B(n_548),
.C(n_540),
.Y(n_776)
);

AOI21x1_ASAP7_75t_L g777 ( 
.A1(n_670),
.A2(n_518),
.B(n_511),
.Y(n_777)
);

NAND2x1p5_ASAP7_75t_L g778 ( 
.A(n_677),
.B(n_526),
.Y(n_778)
);

O2A1O1Ixp33_ASAP7_75t_L g779 ( 
.A1(n_575),
.A2(n_467),
.B(n_484),
.C(n_490),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_674),
.Y(n_780)
);

O2A1O1Ixp5_ASAP7_75t_L g781 ( 
.A1(n_582),
.A2(n_688),
.B(n_641),
.C(n_644),
.Y(n_781)
);

NOR2xp33_ASAP7_75t_L g782 ( 
.A(n_571),
.B(n_538),
.Y(n_782)
);

CKINVDCx5p33_ASAP7_75t_R g783 ( 
.A(n_692),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_L g784 ( 
.A(n_620),
.B(n_433),
.Y(n_784)
);

NOR2xp33_ASAP7_75t_L g785 ( 
.A(n_740),
.B(n_556),
.Y(n_785)
);

CKINVDCx5p33_ASAP7_75t_R g786 ( 
.A(n_692),
.Y(n_786)
);

NOR3xp33_ASAP7_75t_SL g787 ( 
.A(n_583),
.B(n_569),
.C(n_529),
.Y(n_787)
);

AOI22xp5_ASAP7_75t_L g788 ( 
.A1(n_678),
.A2(n_433),
.B1(n_481),
.B2(n_510),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_SL g789 ( 
.A(n_624),
.B(n_556),
.Y(n_789)
);

CKINVDCx5p33_ASAP7_75t_R g790 ( 
.A(n_570),
.Y(n_790)
);

AOI21xp5_ASAP7_75t_L g791 ( 
.A1(n_588),
.A2(n_529),
.B(n_523),
.Y(n_791)
);

AOI21xp5_ASAP7_75t_L g792 ( 
.A1(n_586),
.A2(n_529),
.B(n_523),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_SL g793 ( 
.A(n_624),
.B(n_556),
.Y(n_793)
);

A2O1A1Ixp33_ASAP7_75t_L g794 ( 
.A1(n_612),
.A2(n_511),
.B(n_510),
.C(n_481),
.Y(n_794)
);

CKINVDCx6p67_ASAP7_75t_R g795 ( 
.A(n_662),
.Y(n_795)
);

AOI22xp5_ASAP7_75t_L g796 ( 
.A1(n_576),
.A2(n_433),
.B1(n_481),
.B2(n_510),
.Y(n_796)
);

OAI22xp5_ASAP7_75t_L g797 ( 
.A1(n_609),
.A2(n_569),
.B1(n_523),
.B2(n_511),
.Y(n_797)
);

NOR2xp33_ASAP7_75t_L g798 ( 
.A(n_740),
.B(n_611),
.Y(n_798)
);

O2A1O1Ixp33_ASAP7_75t_L g799 ( 
.A1(n_609),
.A2(n_569),
.B(n_556),
.C(n_518),
.Y(n_799)
);

NOR2xp33_ASAP7_75t_L g800 ( 
.A(n_592),
.B(n_556),
.Y(n_800)
);

OAI22xp5_ASAP7_75t_L g801 ( 
.A1(n_612),
.A2(n_518),
.B1(n_15),
.B2(n_16),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_676),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_L g803 ( 
.A(n_584),
.B(n_14),
.Y(n_803)
);

O2A1O1Ixp33_ASAP7_75t_L g804 ( 
.A1(n_673),
.A2(n_17),
.B(n_21),
.C(n_22),
.Y(n_804)
);

AOI21xp5_ASAP7_75t_L g805 ( 
.A1(n_589),
.A2(n_164),
.B(n_152),
.Y(n_805)
);

BUFx2_ASAP7_75t_L g806 ( 
.A(n_664),
.Y(n_806)
);

INVx2_ASAP7_75t_L g807 ( 
.A(n_686),
.Y(n_807)
);

INVx6_ASAP7_75t_L g808 ( 
.A(n_625),
.Y(n_808)
);

BUFx12f_ASAP7_75t_L g809 ( 
.A(n_703),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_L g810 ( 
.A(n_608),
.B(n_22),
.Y(n_810)
);

OAI22xp5_ASAP7_75t_L g811 ( 
.A1(n_639),
.A2(n_23),
.B1(n_26),
.B2(n_27),
.Y(n_811)
);

AOI21xp5_ASAP7_75t_L g812 ( 
.A1(n_590),
.A2(n_164),
.B(n_152),
.Y(n_812)
);

AOI22xp5_ASAP7_75t_L g813 ( 
.A1(n_576),
.A2(n_164),
.B1(n_152),
.B2(n_32),
.Y(n_813)
);

AOI21xp5_ASAP7_75t_L g814 ( 
.A1(n_656),
.A2(n_164),
.B(n_152),
.Y(n_814)
);

AOI21xp5_ASAP7_75t_L g815 ( 
.A1(n_587),
.A2(n_654),
.B(n_585),
.Y(n_815)
);

O2A1O1Ixp33_ASAP7_75t_L g816 ( 
.A1(n_615),
.A2(n_26),
.B(n_29),
.C(n_34),
.Y(n_816)
);

CKINVDCx14_ASAP7_75t_R g817 ( 
.A(n_739),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_683),
.Y(n_818)
);

NOR2xp33_ASAP7_75t_L g819 ( 
.A(n_601),
.B(n_37),
.Y(n_819)
);

AOI21xp5_ASAP7_75t_L g820 ( 
.A1(n_694),
.A2(n_164),
.B(n_152),
.Y(n_820)
);

NOR2xp33_ASAP7_75t_L g821 ( 
.A(n_601),
.B(n_37),
.Y(n_821)
);

BUFx2_ASAP7_75t_L g822 ( 
.A(n_616),
.Y(n_822)
);

BUFx6f_ASAP7_75t_L g823 ( 
.A(n_627),
.Y(n_823)
);

NOR2xp33_ASAP7_75t_R g824 ( 
.A(n_653),
.B(n_63),
.Y(n_824)
);

NAND3xp33_ASAP7_75t_SL g825 ( 
.A(n_749),
.B(n_38),
.C(n_39),
.Y(n_825)
);

CKINVDCx5p33_ASAP7_75t_R g826 ( 
.A(n_614),
.Y(n_826)
);

AOI22xp5_ASAP7_75t_L g827 ( 
.A1(n_713),
.A2(n_164),
.B1(n_152),
.B2(n_42),
.Y(n_827)
);

AOI21xp5_ASAP7_75t_L g828 ( 
.A1(n_690),
.A2(n_164),
.B(n_152),
.Y(n_828)
);

AND2x2_ASAP7_75t_L g829 ( 
.A(n_724),
.B(n_40),
.Y(n_829)
);

NOR2xp33_ASAP7_75t_SL g830 ( 
.A(n_627),
.B(n_152),
.Y(n_830)
);

CKINVDCx14_ASAP7_75t_R g831 ( 
.A(n_746),
.Y(n_831)
);

A2O1A1Ixp33_ASAP7_75t_SL g832 ( 
.A1(n_583),
.A2(n_40),
.B(n_41),
.C(n_45),
.Y(n_832)
);

AOI22xp5_ASAP7_75t_L g833 ( 
.A1(n_713),
.A2(n_152),
.B1(n_45),
.B2(n_46),
.Y(n_833)
);

AOI21xp5_ASAP7_75t_L g834 ( 
.A1(n_634),
.A2(n_61),
.B(n_59),
.Y(n_834)
);

O2A1O1Ixp33_ASAP7_75t_L g835 ( 
.A1(n_719),
.A2(n_41),
.B(n_47),
.C(n_48),
.Y(n_835)
);

OAI22xp5_ASAP7_75t_L g836 ( 
.A1(n_693),
.A2(n_700),
.B1(n_580),
.B2(n_642),
.Y(n_836)
);

BUFx6f_ASAP7_75t_L g837 ( 
.A(n_632),
.Y(n_837)
);

AOI22xp5_ASAP7_75t_L g838 ( 
.A1(n_716),
.A2(n_48),
.B1(n_49),
.B2(n_50),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_L g839 ( 
.A(n_572),
.B(n_49),
.Y(n_839)
);

O2A1O1Ixp33_ASAP7_75t_L g840 ( 
.A1(n_572),
.A2(n_51),
.B(n_55),
.C(n_58),
.Y(n_840)
);

OAI22xp5_ASAP7_75t_L g841 ( 
.A1(n_633),
.A2(n_51),
.B1(n_594),
.B2(n_630),
.Y(n_841)
);

NOR2xp33_ASAP7_75t_SL g842 ( 
.A(n_677),
.B(n_716),
.Y(n_842)
);

NAND2xp33_ASAP7_75t_L g843 ( 
.A(n_714),
.B(n_593),
.Y(n_843)
);

AOI22xp33_ASAP7_75t_L g844 ( 
.A1(n_682),
.A2(n_661),
.B1(n_701),
.B2(n_702),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_L g845 ( 
.A(n_638),
.B(n_648),
.Y(n_845)
);

AND2x2_ASAP7_75t_L g846 ( 
.A(n_724),
.B(n_737),
.Y(n_846)
);

AOI21xp5_ASAP7_75t_L g847 ( 
.A1(n_596),
.A2(n_628),
.B(n_668),
.Y(n_847)
);

AOI21x1_ASAP7_75t_L g848 ( 
.A1(n_691),
.A2(n_687),
.B(n_688),
.Y(n_848)
);

NOR2xp33_ASAP7_75t_L g849 ( 
.A(n_650),
.B(n_577),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_L g850 ( 
.A(n_638),
.B(n_648),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_L g851 ( 
.A(n_621),
.B(n_737),
.Y(n_851)
);

BUFx12f_ASAP7_75t_L g852 ( 
.A(n_632),
.Y(n_852)
);

INVx2_ASAP7_75t_L g853 ( 
.A(n_705),
.Y(n_853)
);

O2A1O1Ixp33_ASAP7_75t_L g854 ( 
.A1(n_652),
.A2(n_752),
.B(n_732),
.C(n_663),
.Y(n_854)
);

INVxp67_ASAP7_75t_L g855 ( 
.A(n_629),
.Y(n_855)
);

BUFx4f_ASAP7_75t_SL g856 ( 
.A(n_714),
.Y(n_856)
);

HB1xp67_ASAP7_75t_L g857 ( 
.A(n_684),
.Y(n_857)
);

OR2x6_ASAP7_75t_L g858 ( 
.A(n_717),
.B(n_697),
.Y(n_858)
);

AND2x2_ASAP7_75t_L g859 ( 
.A(n_746),
.B(n_744),
.Y(n_859)
);

AND2x4_ASAP7_75t_L g860 ( 
.A(n_714),
.B(n_736),
.Y(n_860)
);

NOR2xp33_ASAP7_75t_L g861 ( 
.A(n_681),
.B(n_598),
.Y(n_861)
);

AOI21xp5_ASAP7_75t_L g862 ( 
.A1(n_617),
.A2(n_618),
.B(n_696),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_SL g863 ( 
.A(n_681),
.B(n_728),
.Y(n_863)
);

INVx3_ASAP7_75t_L g864 ( 
.A(n_727),
.Y(n_864)
);

BUFx12f_ASAP7_75t_L g865 ( 
.A(n_632),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_L g866 ( 
.A(n_714),
.B(n_712),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_L g867 ( 
.A(n_714),
.B(n_718),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_SL g868 ( 
.A(n_632),
.B(n_659),
.Y(n_868)
);

INVx8_ASAP7_75t_L g869 ( 
.A(n_659),
.Y(n_869)
);

AND2x2_ASAP7_75t_L g870 ( 
.A(n_735),
.B(n_600),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_L g871 ( 
.A(n_600),
.B(n_640),
.Y(n_871)
);

OR2x6_ASAP7_75t_L g872 ( 
.A(n_626),
.B(n_727),
.Y(n_872)
);

AOI21xp5_ASAP7_75t_L g873 ( 
.A1(n_622),
.A2(n_680),
.B(n_675),
.Y(n_873)
);

AND2x4_ASAP7_75t_L g874 ( 
.A(n_726),
.B(n_659),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_L g875 ( 
.A(n_743),
.B(n_748),
.Y(n_875)
);

INVx3_ASAP7_75t_L g876 ( 
.A(n_726),
.Y(n_876)
);

AOI21xp5_ASAP7_75t_L g877 ( 
.A1(n_658),
.A2(n_675),
.B(n_610),
.Y(n_877)
);

AND2x4_ASAP7_75t_L g878 ( 
.A(n_659),
.B(n_711),
.Y(n_878)
);

BUFx2_ASAP7_75t_L g879 ( 
.A(n_593),
.Y(n_879)
);

BUFx6f_ASAP7_75t_L g880 ( 
.A(n_626),
.Y(n_880)
);

AOI21xp5_ASAP7_75t_L g881 ( 
.A1(n_658),
.A2(n_679),
.B(n_672),
.Y(n_881)
);

AOI21xp5_ASAP7_75t_L g882 ( 
.A1(n_619),
.A2(n_667),
.B(n_722),
.Y(n_882)
);

HB1xp67_ASAP7_75t_L g883 ( 
.A(n_689),
.Y(n_883)
);

BUFx6f_ASAP7_75t_L g884 ( 
.A(n_730),
.Y(n_884)
);

AOI21xp5_ASAP7_75t_L g885 ( 
.A1(n_619),
.A2(n_722),
.B(n_623),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_SL g886 ( 
.A(n_655),
.B(n_707),
.Y(n_886)
);

AOI33xp33_ASAP7_75t_L g887 ( 
.A1(n_715),
.A2(n_635),
.A3(n_698),
.B1(n_710),
.B2(n_661),
.B3(n_733),
.Y(n_887)
);

NOR2xp33_ASAP7_75t_L g888 ( 
.A(n_699),
.B(n_669),
.Y(n_888)
);

AOI21xp5_ASAP7_75t_L g889 ( 
.A1(n_651),
.A2(n_644),
.B(n_641),
.Y(n_889)
);

AOI21xp5_ASAP7_75t_L g890 ( 
.A1(n_631),
.A2(n_695),
.B(n_671),
.Y(n_890)
);

CKINVDCx5p33_ASAP7_75t_R g891 ( 
.A(n_631),
.Y(n_891)
);

AND2x2_ASAP7_75t_L g892 ( 
.A(n_723),
.B(n_725),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_L g893 ( 
.A(n_657),
.B(n_660),
.Y(n_893)
);

AOI21xp33_ASAP7_75t_L g894 ( 
.A1(n_665),
.A2(n_747),
.B(n_720),
.Y(n_894)
);

NOR2xp33_ASAP7_75t_L g895 ( 
.A(n_685),
.B(n_599),
.Y(n_895)
);

AND2x4_ASAP7_75t_L g896 ( 
.A(n_606),
.B(n_607),
.Y(n_896)
);

BUFx10_ASAP7_75t_L g897 ( 
.A(n_721),
.Y(n_897)
);

AOI21xp5_ASAP7_75t_L g898 ( 
.A1(n_751),
.A2(n_729),
.B(n_750),
.Y(n_898)
);

BUFx6f_ASAP7_75t_L g899 ( 
.A(n_745),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_SL g900 ( 
.A(n_751),
.B(n_731),
.Y(n_900)
);

OAI22xp5_ASAP7_75t_L g901 ( 
.A1(n_706),
.A2(n_709),
.B1(n_734),
.B2(n_738),
.Y(n_901)
);

INVx2_ASAP7_75t_L g902 ( 
.A(n_721),
.Y(n_902)
);

NOR2xp33_ASAP7_75t_L g903 ( 
.A(n_708),
.B(n_741),
.Y(n_903)
);

INVx1_ASAP7_75t_L g904 ( 
.A(n_742),
.Y(n_904)
);

INVx4_ASAP7_75t_L g905 ( 
.A(n_597),
.Y(n_905)
);

OAI22xp5_ASAP7_75t_SL g906 ( 
.A1(n_666),
.A2(n_190),
.B1(n_217),
.B2(n_216),
.Y(n_906)
);

OAI22xp5_ASAP7_75t_L g907 ( 
.A1(n_609),
.A2(n_442),
.B1(n_217),
.B2(n_216),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_L g908 ( 
.A(n_643),
.B(n_272),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_L g909 ( 
.A(n_643),
.B(n_272),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_L g910 ( 
.A(n_643),
.B(n_272),
.Y(n_910)
);

AOI21xp5_ASAP7_75t_L g911 ( 
.A1(n_578),
.A2(n_303),
.B(n_231),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_604),
.Y(n_912)
);

AND2x2_ASAP7_75t_L g913 ( 
.A(n_646),
.B(n_408),
.Y(n_913)
);

NOR3xp33_ASAP7_75t_SL g914 ( 
.A(n_666),
.B(n_191),
.C(n_290),
.Y(n_914)
);

NOR2xp33_ASAP7_75t_R g915 ( 
.A(n_666),
.B(n_422),
.Y(n_915)
);

BUFx6f_ASAP7_75t_L g916 ( 
.A(n_625),
.Y(n_916)
);

BUFx12f_ASAP7_75t_L g917 ( 
.A(n_666),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_L g918 ( 
.A(n_643),
.B(n_272),
.Y(n_918)
);

BUFx6f_ASAP7_75t_L g919 ( 
.A(n_625),
.Y(n_919)
);

AOI21xp5_ASAP7_75t_L g920 ( 
.A1(n_578),
.A2(n_303),
.B(n_231),
.Y(n_920)
);

AOI21xp5_ASAP7_75t_L g921 ( 
.A1(n_578),
.A2(n_303),
.B(n_231),
.Y(n_921)
);

O2A1O1Ixp33_ASAP7_75t_L g922 ( 
.A1(n_573),
.A2(n_334),
.B(n_156),
.C(n_380),
.Y(n_922)
);

AOI22xp5_ASAP7_75t_L g923 ( 
.A1(n_591),
.A2(n_187),
.B1(n_217),
.B2(n_216),
.Y(n_923)
);

AOI21xp5_ASAP7_75t_L g924 ( 
.A1(n_578),
.A2(n_303),
.B(n_231),
.Y(n_924)
);

INVx1_ASAP7_75t_L g925 ( 
.A(n_604),
.Y(n_925)
);

NAND2xp33_ASAP7_75t_SL g926 ( 
.A(n_586),
.B(n_191),
.Y(n_926)
);

BUFx8_ASAP7_75t_L g927 ( 
.A(n_570),
.Y(n_927)
);

NOR2xp33_ASAP7_75t_L g928 ( 
.A(n_649),
.B(n_216),
.Y(n_928)
);

AND2x2_ASAP7_75t_L g929 ( 
.A(n_646),
.B(n_408),
.Y(n_929)
);

CKINVDCx20_ASAP7_75t_R g930 ( 
.A(n_666),
.Y(n_930)
);

NOR2xp67_ASAP7_75t_SL g931 ( 
.A(n_666),
.B(n_422),
.Y(n_931)
);

O2A1O1Ixp33_ASAP7_75t_L g932 ( 
.A1(n_573),
.A2(n_334),
.B(n_156),
.C(n_380),
.Y(n_932)
);

A2O1A1Ixp33_ASAP7_75t_L g933 ( 
.A1(n_573),
.A2(n_704),
.B(n_380),
.C(n_579),
.Y(n_933)
);

NOR2xp33_ASAP7_75t_R g934 ( 
.A(n_666),
.B(n_422),
.Y(n_934)
);

INVx2_ASAP7_75t_L g935 ( 
.A(n_595),
.Y(n_935)
);

OAI21x1_ASAP7_75t_L g936 ( 
.A1(n_628),
.A2(n_687),
.B(n_670),
.Y(n_936)
);

NOR2xp33_ASAP7_75t_L g937 ( 
.A(n_649),
.B(n_216),
.Y(n_937)
);

NOR2xp33_ASAP7_75t_L g938 ( 
.A(n_649),
.B(n_216),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_L g939 ( 
.A(n_643),
.B(n_272),
.Y(n_939)
);

AOI22xp5_ASAP7_75t_L g940 ( 
.A1(n_591),
.A2(n_187),
.B1(n_217),
.B2(n_216),
.Y(n_940)
);

AOI22xp33_ASAP7_75t_L g941 ( 
.A1(n_576),
.A2(n_216),
.B1(n_217),
.B2(n_421),
.Y(n_941)
);

INVx4_ASAP7_75t_L g942 ( 
.A(n_597),
.Y(n_942)
);

INVx2_ASAP7_75t_L g943 ( 
.A(n_595),
.Y(n_943)
);

OAI22xp5_ASAP7_75t_SL g944 ( 
.A1(n_666),
.A2(n_190),
.B1(n_217),
.B2(n_216),
.Y(n_944)
);

OAI22xp5_ASAP7_75t_L g945 ( 
.A1(n_609),
.A2(n_442),
.B1(n_217),
.B2(n_216),
.Y(n_945)
);

NOR2xp33_ASAP7_75t_SL g946 ( 
.A(n_666),
.B(n_290),
.Y(n_946)
);

INVx2_ASAP7_75t_L g947 ( 
.A(n_595),
.Y(n_947)
);

A2O1A1Ixp33_ASAP7_75t_SL g948 ( 
.A1(n_579),
.A2(n_334),
.B(n_380),
.C(n_353),
.Y(n_948)
);

BUFx6f_ASAP7_75t_L g949 ( 
.A(n_625),
.Y(n_949)
);

AOI21xp5_ASAP7_75t_L g950 ( 
.A1(n_578),
.A2(n_303),
.B(n_231),
.Y(n_950)
);

BUFx6f_ASAP7_75t_L g951 ( 
.A(n_625),
.Y(n_951)
);

OAI22xp5_ASAP7_75t_L g952 ( 
.A1(n_609),
.A2(n_442),
.B1(n_217),
.B2(n_216),
.Y(n_952)
);

INVx1_ASAP7_75t_L g953 ( 
.A(n_604),
.Y(n_953)
);

BUFx3_ASAP7_75t_L g954 ( 
.A(n_692),
.Y(n_954)
);

NAND2xp5_ASAP7_75t_L g955 ( 
.A(n_643),
.B(n_272),
.Y(n_955)
);

AND2x2_ASAP7_75t_L g956 ( 
.A(n_646),
.B(n_408),
.Y(n_956)
);

NOR2xp33_ASAP7_75t_L g957 ( 
.A(n_649),
.B(n_216),
.Y(n_957)
);

NAND3xp33_ASAP7_75t_SL g958 ( 
.A(n_605),
.B(n_191),
.C(n_190),
.Y(n_958)
);

INVx2_ASAP7_75t_L g959 ( 
.A(n_595),
.Y(n_959)
);

NAND2xp5_ASAP7_75t_L g960 ( 
.A(n_643),
.B(n_272),
.Y(n_960)
);

NOR2xp33_ASAP7_75t_L g961 ( 
.A(n_649),
.B(n_216),
.Y(n_961)
);

NOR2xp33_ASAP7_75t_L g962 ( 
.A(n_649),
.B(n_216),
.Y(n_962)
);

NAND2xp5_ASAP7_75t_L g963 ( 
.A(n_643),
.B(n_272),
.Y(n_963)
);

AOI21xp5_ASAP7_75t_L g964 ( 
.A1(n_578),
.A2(n_303),
.B(n_231),
.Y(n_964)
);

A2O1A1Ixp33_ASAP7_75t_L g965 ( 
.A1(n_573),
.A2(n_704),
.B(n_380),
.C(n_579),
.Y(n_965)
);

BUFx3_ASAP7_75t_L g966 ( 
.A(n_692),
.Y(n_966)
);

AOI21xp5_ASAP7_75t_L g967 ( 
.A1(n_578),
.A2(n_303),
.B(n_231),
.Y(n_967)
);

NOR2xp33_ASAP7_75t_R g968 ( 
.A(n_666),
.B(n_422),
.Y(n_968)
);

AND2x4_ASAP7_75t_L g969 ( 
.A(n_601),
.B(n_625),
.Y(n_969)
);

NOR3xp33_ASAP7_75t_SL g970 ( 
.A(n_666),
.B(n_191),
.C(n_290),
.Y(n_970)
);

A2O1A1Ixp33_ASAP7_75t_L g971 ( 
.A1(n_573),
.A2(n_704),
.B(n_380),
.C(n_579),
.Y(n_971)
);

NAND2xp5_ASAP7_75t_L g972 ( 
.A(n_643),
.B(n_272),
.Y(n_972)
);

OAI22xp5_ASAP7_75t_L g973 ( 
.A1(n_609),
.A2(n_442),
.B1(n_217),
.B2(n_216),
.Y(n_973)
);

NOR2xp33_ASAP7_75t_R g974 ( 
.A(n_666),
.B(n_422),
.Y(n_974)
);

NOR2xp33_ASAP7_75t_R g975 ( 
.A(n_666),
.B(n_422),
.Y(n_975)
);

BUFx6f_ASAP7_75t_L g976 ( 
.A(n_625),
.Y(n_976)
);

NOR2xp33_ASAP7_75t_L g977 ( 
.A(n_649),
.B(n_216),
.Y(n_977)
);

INVx2_ASAP7_75t_SL g978 ( 
.A(n_837),
.Y(n_978)
);

BUFx3_ASAP7_75t_L g979 ( 
.A(n_852),
.Y(n_979)
);

INVx1_ASAP7_75t_L g980 ( 
.A(n_762),
.Y(n_980)
);

OR2x6_ASAP7_75t_L g981 ( 
.A(n_799),
.B(n_792),
.Y(n_981)
);

BUFx6f_ASAP7_75t_L g982 ( 
.A(n_837),
.Y(n_982)
);

NAND2xp5_ASAP7_75t_L g983 ( 
.A(n_908),
.B(n_909),
.Y(n_983)
);

BUFx3_ASAP7_75t_L g984 ( 
.A(n_865),
.Y(n_984)
);

INVx6_ASAP7_75t_SL g985 ( 
.A(n_969),
.Y(n_985)
);

INVx1_ASAP7_75t_L g986 ( 
.A(n_769),
.Y(n_986)
);

INVx5_ASAP7_75t_L g987 ( 
.A(n_872),
.Y(n_987)
);

BUFx2_ASAP7_75t_L g988 ( 
.A(n_772),
.Y(n_988)
);

NAND2x1p5_ASAP7_75t_L g989 ( 
.A(n_789),
.B(n_793),
.Y(n_989)
);

BUFx3_ASAP7_75t_L g990 ( 
.A(n_954),
.Y(n_990)
);

BUFx3_ASAP7_75t_L g991 ( 
.A(n_966),
.Y(n_991)
);

INVx6_ASAP7_75t_L g992 ( 
.A(n_969),
.Y(n_992)
);

INVx1_ASAP7_75t_L g993 ( 
.A(n_773),
.Y(n_993)
);

INVxp67_ASAP7_75t_SL g994 ( 
.A(n_849),
.Y(n_994)
);

INVx6_ASAP7_75t_L g995 ( 
.A(n_808),
.Y(n_995)
);

CKINVDCx5p33_ASAP7_75t_R g996 ( 
.A(n_915),
.Y(n_996)
);

BUFx8_ASAP7_75t_L g997 ( 
.A(n_770),
.Y(n_997)
);

INVx2_ASAP7_75t_SL g998 ( 
.A(n_837),
.Y(n_998)
);

INVx1_ASAP7_75t_L g999 ( 
.A(n_780),
.Y(n_999)
);

CKINVDCx5p33_ASAP7_75t_R g1000 ( 
.A(n_915),
.Y(n_1000)
);

BUFx5_ASAP7_75t_L g1001 ( 
.A(n_897),
.Y(n_1001)
);

BUFx6f_ASAP7_75t_L g1002 ( 
.A(n_837),
.Y(n_1002)
);

INVx1_ASAP7_75t_L g1003 ( 
.A(n_802),
.Y(n_1003)
);

INVx1_ASAP7_75t_L g1004 ( 
.A(n_818),
.Y(n_1004)
);

BUFx2_ASAP7_75t_L g1005 ( 
.A(n_772),
.Y(n_1005)
);

INVx1_ASAP7_75t_SL g1006 ( 
.A(n_826),
.Y(n_1006)
);

NAND2xp5_ASAP7_75t_L g1007 ( 
.A(n_910),
.B(n_918),
.Y(n_1007)
);

CKINVDCx20_ASAP7_75t_R g1008 ( 
.A(n_930),
.Y(n_1008)
);

BUFx8_ASAP7_75t_L g1009 ( 
.A(n_774),
.Y(n_1009)
);

INVx1_ASAP7_75t_L g1010 ( 
.A(n_912),
.Y(n_1010)
);

INVx2_ASAP7_75t_SL g1011 ( 
.A(n_869),
.Y(n_1011)
);

NAND2xp5_ASAP7_75t_L g1012 ( 
.A(n_939),
.B(n_955),
.Y(n_1012)
);

AND2x2_ASAP7_75t_L g1013 ( 
.A(n_753),
.B(n_883),
.Y(n_1013)
);

AND2x2_ASAP7_75t_L g1014 ( 
.A(n_883),
.B(n_794),
.Y(n_1014)
);

BUFx2_ASAP7_75t_SL g1015 ( 
.A(n_763),
.Y(n_1015)
);

INVx1_ASAP7_75t_L g1016 ( 
.A(n_925),
.Y(n_1016)
);

AND2x2_ASAP7_75t_L g1017 ( 
.A(n_846),
.B(n_796),
.Y(n_1017)
);

INVx1_ASAP7_75t_L g1018 ( 
.A(n_953),
.Y(n_1018)
);

INVx2_ASAP7_75t_SL g1019 ( 
.A(n_869),
.Y(n_1019)
);

INVx4_ASAP7_75t_L g1020 ( 
.A(n_856),
.Y(n_1020)
);

INVx3_ASAP7_75t_L g1021 ( 
.A(n_878),
.Y(n_1021)
);

BUFx12f_ASAP7_75t_L g1022 ( 
.A(n_763),
.Y(n_1022)
);

CKINVDCx11_ASAP7_75t_R g1023 ( 
.A(n_917),
.Y(n_1023)
);

BUFx12f_ASAP7_75t_L g1024 ( 
.A(n_905),
.Y(n_1024)
);

INVx4_ASAP7_75t_L g1025 ( 
.A(n_856),
.Y(n_1025)
);

BUFx6f_ASAP7_75t_L g1026 ( 
.A(n_880),
.Y(n_1026)
);

INVx1_ASAP7_75t_L g1027 ( 
.A(n_756),
.Y(n_1027)
);

BUFx3_ASAP7_75t_L g1028 ( 
.A(n_809),
.Y(n_1028)
);

INVx5_ASAP7_75t_L g1029 ( 
.A(n_872),
.Y(n_1029)
);

BUFx6f_ASAP7_75t_SL g1030 ( 
.A(n_905),
.Y(n_1030)
);

NOR2xp33_ASAP7_75t_L g1031 ( 
.A(n_906),
.B(n_944),
.Y(n_1031)
);

NAND2xp5_ASAP7_75t_L g1032 ( 
.A(n_960),
.B(n_963),
.Y(n_1032)
);

INVx2_ASAP7_75t_SL g1033 ( 
.A(n_869),
.Y(n_1033)
);

BUFx2_ASAP7_75t_SL g1034 ( 
.A(n_942),
.Y(n_1034)
);

BUFx5_ASAP7_75t_L g1035 ( 
.A(n_897),
.Y(n_1035)
);

CKINVDCx6p67_ASAP7_75t_R g1036 ( 
.A(n_942),
.Y(n_1036)
);

INVx4_ASAP7_75t_L g1037 ( 
.A(n_872),
.Y(n_1037)
);

INVx2_ASAP7_75t_SL g1038 ( 
.A(n_874),
.Y(n_1038)
);

INVx3_ASAP7_75t_SL g1039 ( 
.A(n_783),
.Y(n_1039)
);

INVx1_ASAP7_75t_L g1040 ( 
.A(n_764),
.Y(n_1040)
);

INVx5_ASAP7_75t_L g1041 ( 
.A(n_880),
.Y(n_1041)
);

NAND2xp5_ASAP7_75t_L g1042 ( 
.A(n_972),
.B(n_845),
.Y(n_1042)
);

NAND2xp5_ASAP7_75t_L g1043 ( 
.A(n_850),
.B(n_851),
.Y(n_1043)
);

NAND2x1p5_ASAP7_75t_L g1044 ( 
.A(n_880),
.B(n_860),
.Y(n_1044)
);

BUFx2_ASAP7_75t_SL g1045 ( 
.A(n_913),
.Y(n_1045)
);

BUFx3_ASAP7_75t_L g1046 ( 
.A(n_808),
.Y(n_1046)
);

INVx1_ASAP7_75t_SL g1047 ( 
.A(n_934),
.Y(n_1047)
);

BUFx2_ASAP7_75t_L g1048 ( 
.A(n_896),
.Y(n_1048)
);

INVx5_ASAP7_75t_L g1049 ( 
.A(n_899),
.Y(n_1049)
);

INVx3_ASAP7_75t_L g1050 ( 
.A(n_858),
.Y(n_1050)
);

INVx1_ASAP7_75t_L g1051 ( 
.A(n_768),
.Y(n_1051)
);

CKINVDCx5p33_ASAP7_75t_R g1052 ( 
.A(n_934),
.Y(n_1052)
);

AND2x4_ASAP7_75t_L g1053 ( 
.A(n_858),
.B(n_859),
.Y(n_1053)
);

INVx1_ASAP7_75t_L g1054 ( 
.A(n_775),
.Y(n_1054)
);

BUFx10_ASAP7_75t_L g1055 ( 
.A(n_808),
.Y(n_1055)
);

INVx2_ASAP7_75t_SL g1056 ( 
.A(n_823),
.Y(n_1056)
);

INVx1_ASAP7_75t_L g1057 ( 
.A(n_807),
.Y(n_1057)
);

BUFx6f_ASAP7_75t_L g1058 ( 
.A(n_823),
.Y(n_1058)
);

INVx1_ASAP7_75t_L g1059 ( 
.A(n_853),
.Y(n_1059)
);

CKINVDCx5p33_ASAP7_75t_R g1060 ( 
.A(n_975),
.Y(n_1060)
);

CKINVDCx20_ASAP7_75t_R g1061 ( 
.A(n_927),
.Y(n_1061)
);

CKINVDCx6p67_ASAP7_75t_R g1062 ( 
.A(n_795),
.Y(n_1062)
);

CKINVDCx5p33_ASAP7_75t_R g1063 ( 
.A(n_975),
.Y(n_1063)
);

BUFx6f_ASAP7_75t_L g1064 ( 
.A(n_823),
.Y(n_1064)
);

BUFx6f_ASAP7_75t_L g1065 ( 
.A(n_916),
.Y(n_1065)
);

INVx1_ASAP7_75t_L g1066 ( 
.A(n_935),
.Y(n_1066)
);

BUFx3_ASAP7_75t_L g1067 ( 
.A(n_822),
.Y(n_1067)
);

INVx1_ASAP7_75t_L g1068 ( 
.A(n_943),
.Y(n_1068)
);

INVx3_ASAP7_75t_L g1069 ( 
.A(n_858),
.Y(n_1069)
);

INVx5_ASAP7_75t_L g1070 ( 
.A(n_899),
.Y(n_1070)
);

INVx3_ASAP7_75t_L g1071 ( 
.A(n_896),
.Y(n_1071)
);

NOR2xp33_ASAP7_75t_SL g1072 ( 
.A(n_946),
.B(n_931),
.Y(n_1072)
);

BUFx24_ASAP7_75t_L g1073 ( 
.A(n_787),
.Y(n_1073)
);

CKINVDCx16_ASAP7_75t_R g1074 ( 
.A(n_968),
.Y(n_1074)
);

INVx1_ASAP7_75t_SL g1075 ( 
.A(n_974),
.Y(n_1075)
);

BUFx2_ASAP7_75t_SL g1076 ( 
.A(n_929),
.Y(n_1076)
);

INVx1_ASAP7_75t_SL g1077 ( 
.A(n_765),
.Y(n_1077)
);

INVx1_ASAP7_75t_SL g1078 ( 
.A(n_806),
.Y(n_1078)
);

BUFx6f_ASAP7_75t_L g1079 ( 
.A(n_916),
.Y(n_1079)
);

NAND2xp5_ASAP7_75t_L g1080 ( 
.A(n_956),
.B(n_855),
.Y(n_1080)
);

BUFx2_ASAP7_75t_L g1081 ( 
.A(n_884),
.Y(n_1081)
);

AND2x2_ASAP7_75t_L g1082 ( 
.A(n_844),
.B(n_771),
.Y(n_1082)
);

BUFx2_ASAP7_75t_SL g1083 ( 
.A(n_916),
.Y(n_1083)
);

BUFx3_ASAP7_75t_L g1084 ( 
.A(n_916),
.Y(n_1084)
);

INVx5_ASAP7_75t_L g1085 ( 
.A(n_899),
.Y(n_1085)
);

BUFx2_ASAP7_75t_L g1086 ( 
.A(n_884),
.Y(n_1086)
);

AOI22xp33_ASAP7_75t_L g1087 ( 
.A1(n_941),
.A2(n_907),
.B1(n_945),
.B2(n_973),
.Y(n_1087)
);

NAND2x1p5_ASAP7_75t_L g1088 ( 
.A(n_868),
.B(n_758),
.Y(n_1088)
);

INVx1_ASAP7_75t_L g1089 ( 
.A(n_947),
.Y(n_1089)
);

BUFx6f_ASAP7_75t_L g1090 ( 
.A(n_919),
.Y(n_1090)
);

NAND2xp5_ASAP7_75t_L g1091 ( 
.A(n_855),
.B(n_928),
.Y(n_1091)
);

INVxp67_ASAP7_75t_SL g1092 ( 
.A(n_849),
.Y(n_1092)
);

NAND2x1p5_ASAP7_75t_L g1093 ( 
.A(n_919),
.B(n_949),
.Y(n_1093)
);

INVx5_ASAP7_75t_L g1094 ( 
.A(n_899),
.Y(n_1094)
);

NAND2xp5_ASAP7_75t_L g1095 ( 
.A(n_928),
.B(n_937),
.Y(n_1095)
);

BUFx3_ASAP7_75t_L g1096 ( 
.A(n_919),
.Y(n_1096)
);

BUFx2_ASAP7_75t_L g1097 ( 
.A(n_884),
.Y(n_1097)
);

INVx1_ASAP7_75t_SL g1098 ( 
.A(n_790),
.Y(n_1098)
);

BUFx6f_ASAP7_75t_L g1099 ( 
.A(n_949),
.Y(n_1099)
);

BUFx6f_ASAP7_75t_L g1100 ( 
.A(n_949),
.Y(n_1100)
);

NOR2xp33_ASAP7_75t_L g1101 ( 
.A(n_958),
.B(n_831),
.Y(n_1101)
);

BUFx2_ASAP7_75t_L g1102 ( 
.A(n_884),
.Y(n_1102)
);

CKINVDCx11_ASAP7_75t_R g1103 ( 
.A(n_951),
.Y(n_1103)
);

CKINVDCx14_ASAP7_75t_R g1104 ( 
.A(n_817),
.Y(n_1104)
);

BUFx3_ASAP7_75t_L g1105 ( 
.A(n_951),
.Y(n_1105)
);

BUFx2_ASAP7_75t_SL g1106 ( 
.A(n_951),
.Y(n_1106)
);

BUFx3_ASAP7_75t_L g1107 ( 
.A(n_951),
.Y(n_1107)
);

INVx2_ASAP7_75t_L g1108 ( 
.A(n_871),
.Y(n_1108)
);

CKINVDCx5p33_ASAP7_75t_R g1109 ( 
.A(n_914),
.Y(n_1109)
);

OR2x6_ASAP7_75t_L g1110 ( 
.A(n_797),
.B(n_791),
.Y(n_1110)
);

CKINVDCx20_ASAP7_75t_R g1111 ( 
.A(n_927),
.Y(n_1111)
);

NAND2x1p5_ASAP7_75t_L g1112 ( 
.A(n_976),
.B(n_761),
.Y(n_1112)
);

INVx3_ASAP7_75t_L g1113 ( 
.A(n_848),
.Y(n_1113)
);

BUFx12f_ASAP7_75t_L g1114 ( 
.A(n_786),
.Y(n_1114)
);

BUFx4f_ASAP7_75t_L g1115 ( 
.A(n_976),
.Y(n_1115)
);

BUFx12f_ASAP7_75t_L g1116 ( 
.A(n_976),
.Y(n_1116)
);

BUFx6f_ASAP7_75t_SL g1117 ( 
.A(n_976),
.Y(n_1117)
);

INVx1_ASAP7_75t_SL g1118 ( 
.A(n_824),
.Y(n_1118)
);

INVx2_ASAP7_75t_L g1119 ( 
.A(n_875),
.Y(n_1119)
);

AND2x2_ASAP7_75t_L g1120 ( 
.A(n_844),
.B(n_788),
.Y(n_1120)
);

BUFx2_ASAP7_75t_L g1121 ( 
.A(n_891),
.Y(n_1121)
);

INVx2_ASAP7_75t_L g1122 ( 
.A(n_870),
.Y(n_1122)
);

BUFx6f_ASAP7_75t_L g1123 ( 
.A(n_778),
.Y(n_1123)
);

BUFx3_ASAP7_75t_L g1124 ( 
.A(n_761),
.Y(n_1124)
);

AND2x4_ASAP7_75t_L g1125 ( 
.A(n_879),
.B(n_876),
.Y(n_1125)
);

INVx2_ASAP7_75t_SL g1126 ( 
.A(n_778),
.Y(n_1126)
);

INVxp67_ASAP7_75t_SL g1127 ( 
.A(n_782),
.Y(n_1127)
);

NAND2x1p5_ASAP7_75t_L g1128 ( 
.A(n_886),
.B(n_777),
.Y(n_1128)
);

BUFx4_ASAP7_75t_R g1129 ( 
.A(n_824),
.Y(n_1129)
);

INVx1_ASAP7_75t_L g1130 ( 
.A(n_959),
.Y(n_1130)
);

BUFx3_ASAP7_75t_L g1131 ( 
.A(n_864),
.Y(n_1131)
);

BUFx10_ASAP7_75t_L g1132 ( 
.A(n_754),
.Y(n_1132)
);

NAND2xp5_ASAP7_75t_L g1133 ( 
.A(n_937),
.B(n_938),
.Y(n_1133)
);

INVx2_ASAP7_75t_L g1134 ( 
.A(n_904),
.Y(n_1134)
);

INVx3_ASAP7_75t_L g1135 ( 
.A(n_876),
.Y(n_1135)
);

BUFx3_ASAP7_75t_L g1136 ( 
.A(n_864),
.Y(n_1136)
);

INVx5_ASAP7_75t_L g1137 ( 
.A(n_902),
.Y(n_1137)
);

BUFx3_ASAP7_75t_L g1138 ( 
.A(n_754),
.Y(n_1138)
);

BUFx8_ASAP7_75t_L g1139 ( 
.A(n_829),
.Y(n_1139)
);

AOI22xp33_ASAP7_75t_SL g1140 ( 
.A1(n_952),
.A2(n_801),
.B1(n_811),
.B2(n_861),
.Y(n_1140)
);

OR2x2_ASAP7_75t_L g1141 ( 
.A(n_759),
.B(n_784),
.Y(n_1141)
);

INVx5_ASAP7_75t_L g1142 ( 
.A(n_892),
.Y(n_1142)
);

BUFx3_ASAP7_75t_L g1143 ( 
.A(n_755),
.Y(n_1143)
);

INVx1_ASAP7_75t_SL g1144 ( 
.A(n_926),
.Y(n_1144)
);

INVxp67_ASAP7_75t_SL g1145 ( 
.A(n_782),
.Y(n_1145)
);

NOR2xp33_ASAP7_75t_L g1146 ( 
.A(n_819),
.B(n_821),
.Y(n_1146)
);

INVx5_ASAP7_75t_L g1147 ( 
.A(n_843),
.Y(n_1147)
);

INVx4_ASAP7_75t_L g1148 ( 
.A(n_857),
.Y(n_1148)
);

NOR2xp33_ASAP7_75t_L g1149 ( 
.A(n_819),
.B(n_821),
.Y(n_1149)
);

INVx3_ASAP7_75t_SL g1150 ( 
.A(n_863),
.Y(n_1150)
);

INVx1_ASAP7_75t_L g1151 ( 
.A(n_857),
.Y(n_1151)
);

BUFx3_ASAP7_75t_L g1152 ( 
.A(n_755),
.Y(n_1152)
);

BUFx2_ASAP7_75t_SL g1153 ( 
.A(n_838),
.Y(n_1153)
);

INVx1_ASAP7_75t_L g1154 ( 
.A(n_798),
.Y(n_1154)
);

NAND2x1p5_ASAP7_75t_L g1155 ( 
.A(n_785),
.B(n_800),
.Y(n_1155)
);

INVx3_ASAP7_75t_L g1156 ( 
.A(n_936),
.Y(n_1156)
);

BUFx6f_ASAP7_75t_L g1157 ( 
.A(n_866),
.Y(n_1157)
);

BUFx6f_ASAP7_75t_L g1158 ( 
.A(n_867),
.Y(n_1158)
);

BUFx2_ASAP7_75t_SL g1159 ( 
.A(n_923),
.Y(n_1159)
);

OAI22xp5_ASAP7_75t_L g1160 ( 
.A1(n_922),
.A2(n_932),
.B1(n_941),
.B2(n_965),
.Y(n_1160)
);

BUFx6f_ASAP7_75t_L g1161 ( 
.A(n_785),
.Y(n_1161)
);

INVx2_ASAP7_75t_SL g1162 ( 
.A(n_798),
.Y(n_1162)
);

CKINVDCx8_ASAP7_75t_R g1163 ( 
.A(n_938),
.Y(n_1163)
);

OAI22xp5_ASAP7_75t_L g1164 ( 
.A1(n_933),
.A2(n_971),
.B1(n_839),
.B2(n_766),
.Y(n_1164)
);

CKINVDCx5p33_ASAP7_75t_R g1165 ( 
.A(n_914),
.Y(n_1165)
);

AND2x2_ASAP7_75t_L g1166 ( 
.A(n_787),
.B(n_957),
.Y(n_1166)
);

BUFx6f_ASAP7_75t_L g1167 ( 
.A(n_800),
.Y(n_1167)
);

BUFx12f_ASAP7_75t_L g1168 ( 
.A(n_970),
.Y(n_1168)
);

INVx1_ASAP7_75t_L g1169 ( 
.A(n_776),
.Y(n_1169)
);

INVxp67_ASAP7_75t_SL g1170 ( 
.A(n_767),
.Y(n_1170)
);

BUFx6f_ASAP7_75t_L g1171 ( 
.A(n_900),
.Y(n_1171)
);

AOI22xp33_ASAP7_75t_SL g1172 ( 
.A1(n_861),
.A2(n_841),
.B1(n_977),
.B2(n_962),
.Y(n_1172)
);

BUFx6f_ASAP7_75t_L g1173 ( 
.A(n_893),
.Y(n_1173)
);

INVx1_ASAP7_75t_SL g1174 ( 
.A(n_957),
.Y(n_1174)
);

NOR2xp33_ASAP7_75t_L g1175 ( 
.A(n_961),
.B(n_962),
.Y(n_1175)
);

INVx1_ASAP7_75t_L g1176 ( 
.A(n_803),
.Y(n_1176)
);

INVx2_ASAP7_75t_L g1177 ( 
.A(n_781),
.Y(n_1177)
);

INVx1_ASAP7_75t_SL g1178 ( 
.A(n_961),
.Y(n_1178)
);

INVxp67_ASAP7_75t_SL g1179 ( 
.A(n_779),
.Y(n_1179)
);

CKINVDCx20_ASAP7_75t_R g1180 ( 
.A(n_970),
.Y(n_1180)
);

BUFx6f_ASAP7_75t_L g1181 ( 
.A(n_895),
.Y(n_1181)
);

NAND2x1p5_ASAP7_75t_L g1182 ( 
.A(n_888),
.B(n_847),
.Y(n_1182)
);

INVx5_ASAP7_75t_L g1183 ( 
.A(n_842),
.Y(n_1183)
);

BUFx2_ASAP7_75t_L g1184 ( 
.A(n_895),
.Y(n_1184)
);

BUFx6f_ASAP7_75t_L g1185 ( 
.A(n_903),
.Y(n_1185)
);

CKINVDCx5p33_ASAP7_75t_R g1186 ( 
.A(n_977),
.Y(n_1186)
);

INVx5_ASAP7_75t_L g1187 ( 
.A(n_757),
.Y(n_1187)
);

BUFx10_ASAP7_75t_L g1188 ( 
.A(n_903),
.Y(n_1188)
);

BUFx3_ASAP7_75t_L g1189 ( 
.A(n_810),
.Y(n_1189)
);

CKINVDCx5p33_ASAP7_75t_R g1190 ( 
.A(n_940),
.Y(n_1190)
);

INVx2_ASAP7_75t_L g1191 ( 
.A(n_781),
.Y(n_1191)
);

INVx1_ASAP7_75t_L g1192 ( 
.A(n_1134),
.Y(n_1192)
);

NAND2xp5_ASAP7_75t_L g1193 ( 
.A(n_994),
.B(n_760),
.Y(n_1193)
);

INVx1_ASAP7_75t_L g1194 ( 
.A(n_1134),
.Y(n_1194)
);

OR2x2_ASAP7_75t_L g1195 ( 
.A(n_1184),
.B(n_825),
.Y(n_1195)
);

OAI21xp5_ASAP7_75t_L g1196 ( 
.A1(n_1164),
.A2(n_835),
.B(n_948),
.Y(n_1196)
);

AOI22xp33_ASAP7_75t_L g1197 ( 
.A1(n_1159),
.A2(n_1140),
.B1(n_1087),
.B2(n_1120),
.Y(n_1197)
);

INVx1_ASAP7_75t_L g1198 ( 
.A(n_1184),
.Y(n_1198)
);

CKINVDCx5p33_ASAP7_75t_R g1199 ( 
.A(n_1022),
.Y(n_1199)
);

AO21x2_ASAP7_75t_L g1200 ( 
.A1(n_1169),
.A2(n_894),
.B(n_1177),
.Y(n_1200)
);

OAI21x1_ASAP7_75t_L g1201 ( 
.A1(n_1156),
.A2(n_815),
.B(n_873),
.Y(n_1201)
);

BUFx3_ASAP7_75t_L g1202 ( 
.A(n_990),
.Y(n_1202)
);

INVx1_ASAP7_75t_L g1203 ( 
.A(n_1181),
.Y(n_1203)
);

CKINVDCx5p33_ASAP7_75t_R g1204 ( 
.A(n_1022),
.Y(n_1204)
);

AOI22xp33_ASAP7_75t_L g1205 ( 
.A1(n_1120),
.A2(n_813),
.B1(n_836),
.B2(n_833),
.Y(n_1205)
);

AND2x4_ASAP7_75t_L g1206 ( 
.A(n_1071),
.B(n_877),
.Y(n_1206)
);

INVx6_ASAP7_75t_L g1207 ( 
.A(n_1024),
.Y(n_1207)
);

OAI21x1_ASAP7_75t_L g1208 ( 
.A1(n_1156),
.A2(n_862),
.B(n_890),
.Y(n_1208)
);

BUFx6f_ASAP7_75t_L g1209 ( 
.A(n_1049),
.Y(n_1209)
);

INVx1_ASAP7_75t_L g1210 ( 
.A(n_1181),
.Y(n_1210)
);

OAI211xp5_ASAP7_75t_L g1211 ( 
.A1(n_1172),
.A2(n_804),
.B(n_816),
.C(n_840),
.Y(n_1211)
);

OA21x2_ASAP7_75t_L g1212 ( 
.A1(n_1177),
.A2(n_889),
.B(n_885),
.Y(n_1212)
);

INVx1_ASAP7_75t_L g1213 ( 
.A(n_1181),
.Y(n_1213)
);

AND2x4_ASAP7_75t_L g1214 ( 
.A(n_1071),
.B(n_882),
.Y(n_1214)
);

AND2x2_ASAP7_75t_L g1215 ( 
.A(n_1185),
.B(n_1181),
.Y(n_1215)
);

AND2x2_ASAP7_75t_L g1216 ( 
.A(n_1185),
.B(n_881),
.Y(n_1216)
);

O2A1O1Ixp33_ASAP7_75t_SL g1217 ( 
.A1(n_1144),
.A2(n_832),
.B(n_827),
.C(n_854),
.Y(n_1217)
);

OA21x2_ASAP7_75t_L g1218 ( 
.A1(n_1191),
.A2(n_898),
.B(n_812),
.Y(n_1218)
);

AOI22xp5_ASAP7_75t_L g1219 ( 
.A1(n_1160),
.A2(n_830),
.B1(n_834),
.B2(n_901),
.Y(n_1219)
);

OAI22xp33_ASAP7_75t_SL g1220 ( 
.A1(n_1190),
.A2(n_828),
.B1(n_820),
.B2(n_814),
.Y(n_1220)
);

AOI21xp33_ASAP7_75t_L g1221 ( 
.A1(n_1170),
.A2(n_805),
.B(n_921),
.Y(n_1221)
);

OAI21x1_ASAP7_75t_L g1222 ( 
.A1(n_1113),
.A2(n_924),
.B(n_911),
.Y(n_1222)
);

AO31x2_ASAP7_75t_L g1223 ( 
.A1(n_1191),
.A2(n_1081),
.A3(n_1097),
.B(n_1086),
.Y(n_1223)
);

NAND2xp5_ASAP7_75t_L g1224 ( 
.A(n_1092),
.B(n_887),
.Y(n_1224)
);

AND2x4_ASAP7_75t_L g1225 ( 
.A(n_1142),
.B(n_920),
.Y(n_1225)
);

AOI22xp33_ASAP7_75t_SL g1226 ( 
.A1(n_1190),
.A2(n_967),
.B1(n_950),
.B2(n_964),
.Y(n_1226)
);

AND2x4_ASAP7_75t_L g1227 ( 
.A(n_1142),
.B(n_1048),
.Y(n_1227)
);

CKINVDCx6p67_ASAP7_75t_R g1228 ( 
.A(n_1039),
.Y(n_1228)
);

OAI21x1_ASAP7_75t_L g1229 ( 
.A1(n_1113),
.A2(n_1182),
.B(n_1088),
.Y(n_1229)
);

OA21x2_ASAP7_75t_L g1230 ( 
.A1(n_1048),
.A2(n_1086),
.B(n_1081),
.Y(n_1230)
);

OAI22xp5_ASAP7_75t_L g1231 ( 
.A1(n_1175),
.A2(n_1163),
.B1(n_1186),
.B2(n_1149),
.Y(n_1231)
);

AOI22xp33_ASAP7_75t_L g1232 ( 
.A1(n_1153),
.A2(n_1166),
.B1(n_981),
.B2(n_1110),
.Y(n_1232)
);

INVx1_ASAP7_75t_L g1233 ( 
.A(n_1185),
.Y(n_1233)
);

INVx4_ASAP7_75t_SL g1234 ( 
.A(n_1185),
.Y(n_1234)
);

INVx1_ASAP7_75t_L g1235 ( 
.A(n_1185),
.Y(n_1235)
);

NAND2xp5_ASAP7_75t_L g1236 ( 
.A(n_1042),
.B(n_1043),
.Y(n_1236)
);

NAND2xp5_ASAP7_75t_SL g1237 ( 
.A(n_1142),
.B(n_1183),
.Y(n_1237)
);

INVx1_ASAP7_75t_L g1238 ( 
.A(n_1173),
.Y(n_1238)
);

OAI21x1_ASAP7_75t_L g1239 ( 
.A1(n_1113),
.A2(n_1182),
.B(n_1088),
.Y(n_1239)
);

HB1xp67_ASAP7_75t_L g1240 ( 
.A(n_988),
.Y(n_1240)
);

OAI21x1_ASAP7_75t_L g1241 ( 
.A1(n_1182),
.A2(n_1088),
.B(n_1128),
.Y(n_1241)
);

AO21x2_ASAP7_75t_L g1242 ( 
.A1(n_1179),
.A2(n_1166),
.B(n_986),
.Y(n_1242)
);

BUFx6f_ASAP7_75t_L g1243 ( 
.A(n_1049),
.Y(n_1243)
);

INVx1_ASAP7_75t_L g1244 ( 
.A(n_1173),
.Y(n_1244)
);

OAI222xp33_ASAP7_75t_L g1245 ( 
.A1(n_1110),
.A2(n_1082),
.B1(n_981),
.B2(n_1163),
.C1(n_1133),
.C2(n_1095),
.Y(n_1245)
);

HB1xp67_ASAP7_75t_L g1246 ( 
.A(n_988),
.Y(n_1246)
);

NOR2x1_ASAP7_75t_SL g1247 ( 
.A(n_1147),
.B(n_1142),
.Y(n_1247)
);

INVxp67_ASAP7_75t_SL g1248 ( 
.A(n_1127),
.Y(n_1248)
);

INVx3_ASAP7_75t_L g1249 ( 
.A(n_1171),
.Y(n_1249)
);

AOI21xp5_ASAP7_75t_L g1250 ( 
.A1(n_1187),
.A2(n_1070),
.B(n_1049),
.Y(n_1250)
);

AOI21xp5_ASAP7_75t_L g1251 ( 
.A1(n_1187),
.A2(n_1070),
.B(n_1049),
.Y(n_1251)
);

BUFx2_ASAP7_75t_L g1252 ( 
.A(n_1142),
.Y(n_1252)
);

AOI21xp5_ASAP7_75t_L g1253 ( 
.A1(n_1187),
.A2(n_1070),
.B(n_1049),
.Y(n_1253)
);

INVx6_ASAP7_75t_L g1254 ( 
.A(n_1024),
.Y(n_1254)
);

AOI22x1_ASAP7_75t_L g1255 ( 
.A1(n_1186),
.A2(n_1109),
.B1(n_1165),
.B2(n_1052),
.Y(n_1255)
);

AND2x2_ASAP7_75t_L g1256 ( 
.A(n_1013),
.B(n_1005),
.Y(n_1256)
);

AND2x4_ASAP7_75t_L g1257 ( 
.A(n_1147),
.B(n_1050),
.Y(n_1257)
);

HB1xp67_ASAP7_75t_L g1258 ( 
.A(n_1005),
.Y(n_1258)
);

NAND2x1p5_ASAP7_75t_L g1259 ( 
.A(n_1147),
.B(n_1070),
.Y(n_1259)
);

AND2x4_ASAP7_75t_L g1260 ( 
.A(n_1147),
.B(n_1050),
.Y(n_1260)
);

INVx2_ASAP7_75t_L g1261 ( 
.A(n_1108),
.Y(n_1261)
);

BUFx2_ASAP7_75t_L g1262 ( 
.A(n_1148),
.Y(n_1262)
);

NAND2xp5_ASAP7_75t_L g1263 ( 
.A(n_1145),
.B(n_1154),
.Y(n_1263)
);

OAI21x1_ASAP7_75t_L g1264 ( 
.A1(n_989),
.A2(n_1044),
.B(n_1135),
.Y(n_1264)
);

NOR2xp33_ASAP7_75t_L g1265 ( 
.A(n_1174),
.B(n_1178),
.Y(n_1265)
);

INVx1_ASAP7_75t_SL g1266 ( 
.A(n_1045),
.Y(n_1266)
);

OA21x2_ASAP7_75t_L g1267 ( 
.A1(n_1097),
.A2(n_1102),
.B(n_993),
.Y(n_1267)
);

AO21x2_ASAP7_75t_L g1268 ( 
.A1(n_980),
.A2(n_1003),
.B(n_999),
.Y(n_1268)
);

INVx1_ASAP7_75t_L g1269 ( 
.A(n_1173),
.Y(n_1269)
);

NAND2x1p5_ASAP7_75t_L g1270 ( 
.A(n_1070),
.B(n_1085),
.Y(n_1270)
);

AOI22xp33_ASAP7_75t_SL g1271 ( 
.A1(n_1082),
.A2(n_1187),
.B1(n_981),
.B2(n_1014),
.Y(n_1271)
);

NAND2xp5_ASAP7_75t_L g1272 ( 
.A(n_1162),
.B(n_983),
.Y(n_1272)
);

NOR2x1_ASAP7_75t_L g1273 ( 
.A(n_1148),
.B(n_1189),
.Y(n_1273)
);

INVx1_ASAP7_75t_L g1274 ( 
.A(n_1173),
.Y(n_1274)
);

BUFx12f_ASAP7_75t_L g1275 ( 
.A(n_1023),
.Y(n_1275)
);

AO31x2_ASAP7_75t_L g1276 ( 
.A1(n_1102),
.A2(n_1119),
.A3(n_1016),
.B(n_1010),
.Y(n_1276)
);

INVx2_ASAP7_75t_L g1277 ( 
.A(n_1173),
.Y(n_1277)
);

AOI221xp5_ASAP7_75t_SL g1278 ( 
.A1(n_1031),
.A2(n_1146),
.B1(n_1078),
.B2(n_1180),
.C(n_1091),
.Y(n_1278)
);

INVx1_ASAP7_75t_L g1279 ( 
.A(n_1151),
.Y(n_1279)
);

AO21x2_ASAP7_75t_L g1280 ( 
.A1(n_1004),
.A2(n_1018),
.B(n_1176),
.Y(n_1280)
);

BUFx2_ASAP7_75t_L g1281 ( 
.A(n_1148),
.Y(n_1281)
);

INVx1_ASAP7_75t_L g1282 ( 
.A(n_1141),
.Y(n_1282)
);

INVx2_ASAP7_75t_L g1283 ( 
.A(n_1157),
.Y(n_1283)
);

INVx3_ASAP7_75t_L g1284 ( 
.A(n_1171),
.Y(n_1284)
);

INVx1_ASAP7_75t_L g1285 ( 
.A(n_1141),
.Y(n_1285)
);

INVx1_ASAP7_75t_L g1286 ( 
.A(n_1188),
.Y(n_1286)
);

INVx1_ASAP7_75t_L g1287 ( 
.A(n_1188),
.Y(n_1287)
);

AND2x4_ASAP7_75t_L g1288 ( 
.A(n_1050),
.B(n_1069),
.Y(n_1288)
);

AO21x2_ASAP7_75t_L g1289 ( 
.A1(n_1080),
.A2(n_1014),
.B(n_1027),
.Y(n_1289)
);

INVx2_ASAP7_75t_L g1290 ( 
.A(n_1157),
.Y(n_1290)
);

OAI21xp5_ASAP7_75t_L g1291 ( 
.A1(n_1189),
.A2(n_1118),
.B(n_1101),
.Y(n_1291)
);

INVx3_ASAP7_75t_L g1292 ( 
.A(n_1171),
.Y(n_1292)
);

OAI22xp33_ASAP7_75t_L g1293 ( 
.A1(n_981),
.A2(n_1110),
.B1(n_1187),
.B2(n_1150),
.Y(n_1293)
);

INVx2_ASAP7_75t_L g1294 ( 
.A(n_1157),
.Y(n_1294)
);

NOR2xp33_ASAP7_75t_SL g1295 ( 
.A(n_1183),
.B(n_1085),
.Y(n_1295)
);

AND2x2_ASAP7_75t_L g1296 ( 
.A(n_1013),
.B(n_1188),
.Y(n_1296)
);

INVx1_ASAP7_75t_L g1297 ( 
.A(n_1137),
.Y(n_1297)
);

INVx1_ASAP7_75t_L g1298 ( 
.A(n_1137),
.Y(n_1298)
);

INVx1_ASAP7_75t_L g1299 ( 
.A(n_1137),
.Y(n_1299)
);

OAI221xp5_ASAP7_75t_L g1300 ( 
.A1(n_1006),
.A2(n_1072),
.B1(n_1150),
.B2(n_1077),
.C(n_1110),
.Y(n_1300)
);

BUFx6f_ASAP7_75t_L g1301 ( 
.A(n_1085),
.Y(n_1301)
);

AO21x2_ASAP7_75t_L g1302 ( 
.A1(n_1040),
.A2(n_1068),
.B(n_1051),
.Y(n_1302)
);

AOI22xp33_ASAP7_75t_L g1303 ( 
.A1(n_1017),
.A2(n_1122),
.B1(n_1076),
.B2(n_1066),
.Y(n_1303)
);

INVx2_ASAP7_75t_SL g1304 ( 
.A(n_1085),
.Y(n_1304)
);

O2A1O1Ixp33_ASAP7_75t_SL g1305 ( 
.A1(n_1180),
.A2(n_1047),
.B(n_1075),
.C(n_1061),
.Y(n_1305)
);

INVx1_ASAP7_75t_L g1306 ( 
.A(n_1137),
.Y(n_1306)
);

AO21x2_ASAP7_75t_L g1307 ( 
.A1(n_1054),
.A2(n_1089),
.B(n_1130),
.Y(n_1307)
);

AOI21xp5_ASAP7_75t_L g1308 ( 
.A1(n_1085),
.A2(n_1094),
.B(n_1183),
.Y(n_1308)
);

INVx1_ASAP7_75t_L g1309 ( 
.A(n_1137),
.Y(n_1309)
);

OAI22xp5_ASAP7_75t_L g1310 ( 
.A1(n_1121),
.A2(n_1155),
.B1(n_1109),
.B2(n_1165),
.Y(n_1310)
);

INVx6_ASAP7_75t_L g1311 ( 
.A(n_1183),
.Y(n_1311)
);

INVx1_ASAP7_75t_L g1312 ( 
.A(n_1157),
.Y(n_1312)
);

OA21x2_ASAP7_75t_L g1313 ( 
.A1(n_1122),
.A2(n_1057),
.B(n_1059),
.Y(n_1313)
);

INVx2_ASAP7_75t_L g1314 ( 
.A(n_1157),
.Y(n_1314)
);

AND2x2_ASAP7_75t_L g1315 ( 
.A(n_1162),
.B(n_1017),
.Y(n_1315)
);

A2O1A1Ixp33_ASAP7_75t_L g1316 ( 
.A1(n_1094),
.A2(n_1129),
.B(n_1183),
.C(n_1138),
.Y(n_1316)
);

INVx1_ASAP7_75t_SL g1317 ( 
.A(n_1121),
.Y(n_1317)
);

INVx1_ASAP7_75t_L g1318 ( 
.A(n_1158),
.Y(n_1318)
);

OAI22xp5_ASAP7_75t_L g1319 ( 
.A1(n_1155),
.A2(n_1094),
.B1(n_1020),
.B2(n_1025),
.Y(n_1319)
);

INVx1_ASAP7_75t_SL g1320 ( 
.A(n_1094),
.Y(n_1320)
);

INVx2_ASAP7_75t_L g1321 ( 
.A(n_1158),
.Y(n_1321)
);

AO21x2_ASAP7_75t_L g1322 ( 
.A1(n_1007),
.A2(n_1012),
.B(n_1032),
.Y(n_1322)
);

OAI21xp5_ASAP7_75t_L g1323 ( 
.A1(n_1115),
.A2(n_1094),
.B(n_1112),
.Y(n_1323)
);

AND2x2_ASAP7_75t_L g1324 ( 
.A(n_1167),
.B(n_1161),
.Y(n_1324)
);

OA21x2_ASAP7_75t_L g1325 ( 
.A1(n_1053),
.A2(n_978),
.B(n_998),
.Y(n_1325)
);

AOI22xp5_ASAP7_75t_L g1326 ( 
.A1(n_1143),
.A2(n_1152),
.B1(n_1138),
.B2(n_1139),
.Y(n_1326)
);

BUFx3_ASAP7_75t_L g1327 ( 
.A(n_990),
.Y(n_1327)
);

AOI21xp33_ASAP7_75t_L g1328 ( 
.A1(n_1171),
.A2(n_1126),
.B(n_1158),
.Y(n_1328)
);

AOI22xp33_ASAP7_75t_L g1329 ( 
.A1(n_1167),
.A2(n_1053),
.B1(n_1143),
.B2(n_1152),
.Y(n_1329)
);

AND2x2_ASAP7_75t_L g1330 ( 
.A(n_1167),
.B(n_1161),
.Y(n_1330)
);

INVx4_ASAP7_75t_L g1331 ( 
.A(n_1001),
.Y(n_1331)
);

INVx1_ASAP7_75t_L g1332 ( 
.A(n_1158),
.Y(n_1332)
);

INVx2_ASAP7_75t_L g1333 ( 
.A(n_1158),
.Y(n_1333)
);

BUFx2_ASAP7_75t_R g1334 ( 
.A(n_1028),
.Y(n_1334)
);

INVx1_ASAP7_75t_L g1335 ( 
.A(n_1171),
.Y(n_1335)
);

OR2x6_ASAP7_75t_L g1336 ( 
.A(n_1037),
.B(n_1053),
.Y(n_1336)
);

AOI22xp33_ASAP7_75t_L g1337 ( 
.A1(n_1167),
.A2(n_1161),
.B1(n_1139),
.B2(n_1021),
.Y(n_1337)
);

BUFx3_ASAP7_75t_L g1338 ( 
.A(n_991),
.Y(n_1338)
);

OAI21x1_ASAP7_75t_L g1339 ( 
.A1(n_1093),
.A2(n_1112),
.B(n_1001),
.Y(n_1339)
);

BUFx3_ASAP7_75t_L g1340 ( 
.A(n_991),
.Y(n_1340)
);

NAND2xp33_ASAP7_75t_R g1341 ( 
.A(n_996),
.B(n_1000),
.Y(n_1341)
);

NOR2xp33_ASAP7_75t_L g1342 ( 
.A(n_1008),
.B(n_1098),
.Y(n_1342)
);

INVx2_ASAP7_75t_L g1343 ( 
.A(n_1167),
.Y(n_1343)
);

OAI21x1_ASAP7_75t_L g1344 ( 
.A1(n_1001),
.A2(n_1035),
.B(n_1073),
.Y(n_1344)
);

OAI21xp5_ASAP7_75t_L g1345 ( 
.A1(n_1115),
.A2(n_978),
.B(n_998),
.Y(n_1345)
);

INVx1_ASAP7_75t_SL g1346 ( 
.A(n_1067),
.Y(n_1346)
);

OAI21x1_ASAP7_75t_L g1347 ( 
.A1(n_1001),
.A2(n_1035),
.B(n_1073),
.Y(n_1347)
);

BUFx2_ASAP7_75t_L g1348 ( 
.A(n_1001),
.Y(n_1348)
);

INVx2_ASAP7_75t_L g1349 ( 
.A(n_1001),
.Y(n_1349)
);

OAI21x1_ASAP7_75t_L g1350 ( 
.A1(n_1001),
.A2(n_1035),
.B(n_982),
.Y(n_1350)
);

OAI21x1_ASAP7_75t_L g1351 ( 
.A1(n_1035),
.A2(n_982),
.B(n_1002),
.Y(n_1351)
);

NAND3xp33_ASAP7_75t_L g1352 ( 
.A(n_1139),
.B(n_1161),
.C(n_1103),
.Y(n_1352)
);

INVx2_ASAP7_75t_L g1353 ( 
.A(n_1035),
.Y(n_1353)
);

INVx1_ASAP7_75t_L g1354 ( 
.A(n_1268),
.Y(n_1354)
);

HB1xp67_ASAP7_75t_L g1355 ( 
.A(n_1240),
.Y(n_1355)
);

CKINVDCx11_ASAP7_75t_R g1356 ( 
.A(n_1275),
.Y(n_1356)
);

INVx1_ASAP7_75t_L g1357 ( 
.A(n_1268),
.Y(n_1357)
);

CKINVDCx16_ASAP7_75t_R g1358 ( 
.A(n_1275),
.Y(n_1358)
);

INVx2_ASAP7_75t_L g1359 ( 
.A(n_1192),
.Y(n_1359)
);

INVx2_ASAP7_75t_L g1360 ( 
.A(n_1192),
.Y(n_1360)
);

NOR2xp67_ASAP7_75t_L g1361 ( 
.A(n_1352),
.B(n_987),
.Y(n_1361)
);

BUFx3_ASAP7_75t_L g1362 ( 
.A(n_1325),
.Y(n_1362)
);

INVx2_ASAP7_75t_L g1363 ( 
.A(n_1194),
.Y(n_1363)
);

INVx1_ASAP7_75t_L g1364 ( 
.A(n_1268),
.Y(n_1364)
);

INVx2_ASAP7_75t_L g1365 ( 
.A(n_1194),
.Y(n_1365)
);

AND2x2_ASAP7_75t_L g1366 ( 
.A(n_1256),
.B(n_1035),
.Y(n_1366)
);

AND2x2_ASAP7_75t_L g1367 ( 
.A(n_1256),
.B(n_1161),
.Y(n_1367)
);

HB1xp67_ASAP7_75t_L g1368 ( 
.A(n_1246),
.Y(n_1368)
);

AND2x2_ASAP7_75t_L g1369 ( 
.A(n_1215),
.B(n_982),
.Y(n_1369)
);

INVx1_ASAP7_75t_L g1370 ( 
.A(n_1276),
.Y(n_1370)
);

AOI22xp33_ASAP7_75t_L g1371 ( 
.A1(n_1197),
.A2(n_1132),
.B1(n_992),
.B2(n_985),
.Y(n_1371)
);

INVx2_ASAP7_75t_L g1372 ( 
.A(n_1276),
.Y(n_1372)
);

BUFx6f_ASAP7_75t_L g1373 ( 
.A(n_1209),
.Y(n_1373)
);

INVx2_ASAP7_75t_L g1374 ( 
.A(n_1276),
.Y(n_1374)
);

INVx1_ASAP7_75t_L g1375 ( 
.A(n_1276),
.Y(n_1375)
);

INVx3_ASAP7_75t_L g1376 ( 
.A(n_1206),
.Y(n_1376)
);

INVx2_ASAP7_75t_L g1377 ( 
.A(n_1276),
.Y(n_1377)
);

INVx2_ASAP7_75t_L g1378 ( 
.A(n_1313),
.Y(n_1378)
);

INVx1_ASAP7_75t_L g1379 ( 
.A(n_1280),
.Y(n_1379)
);

INVx1_ASAP7_75t_L g1380 ( 
.A(n_1280),
.Y(n_1380)
);

INVx1_ASAP7_75t_L g1381 ( 
.A(n_1280),
.Y(n_1381)
);

OAI21x1_ASAP7_75t_L g1382 ( 
.A1(n_1201),
.A2(n_1002),
.B(n_1037),
.Y(n_1382)
);

BUFx2_ASAP7_75t_SL g1383 ( 
.A(n_1237),
.Y(n_1383)
);

OR2x2_ASAP7_75t_L g1384 ( 
.A(n_1198),
.B(n_1067),
.Y(n_1384)
);

BUFx3_ASAP7_75t_L g1385 ( 
.A(n_1325),
.Y(n_1385)
);

BUFx3_ASAP7_75t_L g1386 ( 
.A(n_1325),
.Y(n_1386)
);

HB1xp67_ASAP7_75t_L g1387 ( 
.A(n_1258),
.Y(n_1387)
);

INVx2_ASAP7_75t_L g1388 ( 
.A(n_1313),
.Y(n_1388)
);

INVx2_ASAP7_75t_L g1389 ( 
.A(n_1313),
.Y(n_1389)
);

BUFx3_ASAP7_75t_L g1390 ( 
.A(n_1325),
.Y(n_1390)
);

AND2x2_ASAP7_75t_L g1391 ( 
.A(n_1215),
.B(n_1002),
.Y(n_1391)
);

INVx2_ASAP7_75t_L g1392 ( 
.A(n_1313),
.Y(n_1392)
);

NOR2x1_ASAP7_75t_R g1393 ( 
.A(n_1207),
.B(n_1023),
.Y(n_1393)
);

INVx2_ASAP7_75t_L g1394 ( 
.A(n_1302),
.Y(n_1394)
);

INVx2_ASAP7_75t_L g1395 ( 
.A(n_1302),
.Y(n_1395)
);

OAI21x1_ASAP7_75t_L g1396 ( 
.A1(n_1201),
.A2(n_1002),
.B(n_1029),
.Y(n_1396)
);

HB1xp67_ASAP7_75t_L g1397 ( 
.A(n_1267),
.Y(n_1397)
);

INVx1_ASAP7_75t_L g1398 ( 
.A(n_1279),
.Y(n_1398)
);

INVx2_ASAP7_75t_SL g1399 ( 
.A(n_1267),
.Y(n_1399)
);

INVx3_ASAP7_75t_L g1400 ( 
.A(n_1206),
.Y(n_1400)
);

INVx2_ASAP7_75t_L g1401 ( 
.A(n_1302),
.Y(n_1401)
);

OAI21x1_ASAP7_75t_L g1402 ( 
.A1(n_1208),
.A2(n_1222),
.B(n_1241),
.Y(n_1402)
);

INVx2_ASAP7_75t_L g1403 ( 
.A(n_1307),
.Y(n_1403)
);

BUFx3_ASAP7_75t_L g1404 ( 
.A(n_1230),
.Y(n_1404)
);

AOI21x1_ASAP7_75t_L g1405 ( 
.A1(n_1250),
.A2(n_1125),
.B(n_1056),
.Y(n_1405)
);

INVx2_ASAP7_75t_L g1406 ( 
.A(n_1307),
.Y(n_1406)
);

INVx1_ASAP7_75t_L g1407 ( 
.A(n_1279),
.Y(n_1407)
);

INVx2_ASAP7_75t_L g1408 ( 
.A(n_1307),
.Y(n_1408)
);

INVx1_ASAP7_75t_L g1409 ( 
.A(n_1198),
.Y(n_1409)
);

INVx3_ASAP7_75t_L g1410 ( 
.A(n_1206),
.Y(n_1410)
);

AO21x2_ASAP7_75t_L g1411 ( 
.A1(n_1242),
.A2(n_1132),
.B(n_1029),
.Y(n_1411)
);

CKINVDCx20_ASAP7_75t_R g1412 ( 
.A(n_1228),
.Y(n_1412)
);

INVx1_ASAP7_75t_L g1413 ( 
.A(n_1289),
.Y(n_1413)
);

INVx2_ASAP7_75t_L g1414 ( 
.A(n_1261),
.Y(n_1414)
);

BUFx3_ASAP7_75t_L g1415 ( 
.A(n_1230),
.Y(n_1415)
);

BUFx3_ASAP7_75t_L g1416 ( 
.A(n_1230),
.Y(n_1416)
);

BUFx2_ASAP7_75t_L g1417 ( 
.A(n_1273),
.Y(n_1417)
);

BUFx3_ASAP7_75t_L g1418 ( 
.A(n_1230),
.Y(n_1418)
);

INVx1_ASAP7_75t_L g1419 ( 
.A(n_1289),
.Y(n_1419)
);

INVx1_ASAP7_75t_L g1420 ( 
.A(n_1289),
.Y(n_1420)
);

INVx2_ASAP7_75t_L g1421 ( 
.A(n_1261),
.Y(n_1421)
);

INVx3_ASAP7_75t_L g1422 ( 
.A(n_1206),
.Y(n_1422)
);

AO21x2_ASAP7_75t_L g1423 ( 
.A1(n_1242),
.A2(n_1200),
.B(n_1196),
.Y(n_1423)
);

AND2x2_ASAP7_75t_L g1424 ( 
.A(n_1212),
.B(n_1132),
.Y(n_1424)
);

AOI22xp33_ASAP7_75t_L g1425 ( 
.A1(n_1205),
.A2(n_992),
.B1(n_985),
.B2(n_1168),
.Y(n_1425)
);

HB1xp67_ASAP7_75t_L g1426 ( 
.A(n_1267),
.Y(n_1426)
);

OAI21x1_ASAP7_75t_L g1427 ( 
.A1(n_1208),
.A2(n_1029),
.B(n_987),
.Y(n_1427)
);

CKINVDCx6p67_ASAP7_75t_R g1428 ( 
.A(n_1228),
.Y(n_1428)
);

INVx2_ASAP7_75t_L g1429 ( 
.A(n_1212),
.Y(n_1429)
);

BUFx12f_ASAP7_75t_L g1430 ( 
.A(n_1199),
.Y(n_1430)
);

INVx2_ASAP7_75t_L g1431 ( 
.A(n_1212),
.Y(n_1431)
);

BUFx3_ASAP7_75t_L g1432 ( 
.A(n_1202),
.Y(n_1432)
);

INVxp67_ASAP7_75t_L g1433 ( 
.A(n_1242),
.Y(n_1433)
);

INVx1_ASAP7_75t_L g1434 ( 
.A(n_1233),
.Y(n_1434)
);

INVx2_ASAP7_75t_L g1435 ( 
.A(n_1212),
.Y(n_1435)
);

INVx1_ASAP7_75t_L g1436 ( 
.A(n_1233),
.Y(n_1436)
);

INVx1_ASAP7_75t_L g1437 ( 
.A(n_1235),
.Y(n_1437)
);

INVx1_ASAP7_75t_L g1438 ( 
.A(n_1235),
.Y(n_1438)
);

INVx2_ASAP7_75t_SL g1439 ( 
.A(n_1267),
.Y(n_1439)
);

INVx1_ASAP7_75t_L g1440 ( 
.A(n_1335),
.Y(n_1440)
);

NAND3xp33_ASAP7_75t_L g1441 ( 
.A(n_1211),
.B(n_1103),
.C(n_1065),
.Y(n_1441)
);

AOI221xp5_ASAP7_75t_L g1442 ( 
.A1(n_1278),
.A2(n_1028),
.B1(n_1104),
.B2(n_1111),
.C(n_1061),
.Y(n_1442)
);

HB1xp67_ASAP7_75t_L g1443 ( 
.A(n_1223),
.Y(n_1443)
);

INVx1_ASAP7_75t_L g1444 ( 
.A(n_1335),
.Y(n_1444)
);

AND2x4_ASAP7_75t_L g1445 ( 
.A(n_1252),
.B(n_1105),
.Y(n_1445)
);

INVx4_ASAP7_75t_L g1446 ( 
.A(n_1259),
.Y(n_1446)
);

BUFx2_ASAP7_75t_L g1447 ( 
.A(n_1273),
.Y(n_1447)
);

OR2x6_ASAP7_75t_L g1448 ( 
.A(n_1259),
.B(n_1025),
.Y(n_1448)
);

OA21x2_ASAP7_75t_L g1449 ( 
.A1(n_1229),
.A2(n_1038),
.B(n_1056),
.Y(n_1449)
);

INVx3_ASAP7_75t_L g1450 ( 
.A(n_1239),
.Y(n_1450)
);

INVx1_ASAP7_75t_L g1451 ( 
.A(n_1282),
.Y(n_1451)
);

AOI22xp5_ASAP7_75t_SL g1452 ( 
.A1(n_1266),
.A2(n_1111),
.B1(n_1008),
.B2(n_1063),
.Y(n_1452)
);

BUFx3_ASAP7_75t_L g1453 ( 
.A(n_1202),
.Y(n_1453)
);

INVx1_ASAP7_75t_L g1454 ( 
.A(n_1282),
.Y(n_1454)
);

AND2x2_ASAP7_75t_L g1455 ( 
.A(n_1203),
.B(n_1058),
.Y(n_1455)
);

INVx1_ASAP7_75t_L g1456 ( 
.A(n_1285),
.Y(n_1456)
);

AOI22xp33_ASAP7_75t_L g1457 ( 
.A1(n_1195),
.A2(n_992),
.B1(n_985),
.B2(n_1168),
.Y(n_1457)
);

INVx2_ASAP7_75t_L g1458 ( 
.A(n_1218),
.Y(n_1458)
);

INVx1_ASAP7_75t_L g1459 ( 
.A(n_1285),
.Y(n_1459)
);

HB1xp67_ASAP7_75t_L g1460 ( 
.A(n_1223),
.Y(n_1460)
);

INVx1_ASAP7_75t_L g1461 ( 
.A(n_1203),
.Y(n_1461)
);

AOI22xp33_ASAP7_75t_L g1462 ( 
.A1(n_1195),
.A2(n_992),
.B1(n_1114),
.B2(n_1020),
.Y(n_1462)
);

BUFx3_ASAP7_75t_L g1463 ( 
.A(n_1327),
.Y(n_1463)
);

INVx1_ASAP7_75t_L g1464 ( 
.A(n_1210),
.Y(n_1464)
);

HB1xp67_ASAP7_75t_L g1465 ( 
.A(n_1223),
.Y(n_1465)
);

OA21x2_ASAP7_75t_L g1466 ( 
.A1(n_1222),
.A2(n_1011),
.B(n_1033),
.Y(n_1466)
);

NAND2xp5_ASAP7_75t_L g1467 ( 
.A(n_1248),
.B(n_1136),
.Y(n_1467)
);

NAND2xp5_ASAP7_75t_L g1468 ( 
.A(n_1263),
.B(n_1136),
.Y(n_1468)
);

INVx1_ASAP7_75t_L g1469 ( 
.A(n_1210),
.Y(n_1469)
);

INVx2_ASAP7_75t_L g1470 ( 
.A(n_1218),
.Y(n_1470)
);

INVx1_ASAP7_75t_L g1471 ( 
.A(n_1213),
.Y(n_1471)
);

OAI22xp5_ASAP7_75t_L g1472 ( 
.A1(n_1224),
.A2(n_1025),
.B1(n_1020),
.B2(n_1074),
.Y(n_1472)
);

INVx1_ASAP7_75t_L g1473 ( 
.A(n_1213),
.Y(n_1473)
);

AND2x2_ASAP7_75t_L g1474 ( 
.A(n_1227),
.B(n_1079),
.Y(n_1474)
);

BUFx2_ASAP7_75t_L g1475 ( 
.A(n_1252),
.Y(n_1475)
);

AOI21x1_ASAP7_75t_L g1476 ( 
.A1(n_1251),
.A2(n_1253),
.B(n_1308),
.Y(n_1476)
);

INVx2_ASAP7_75t_L g1477 ( 
.A(n_1218),
.Y(n_1477)
);

INVx3_ASAP7_75t_L g1478 ( 
.A(n_1214),
.Y(n_1478)
);

INVx1_ASAP7_75t_L g1479 ( 
.A(n_1312),
.Y(n_1479)
);

AOI22xp5_ASAP7_75t_L g1480 ( 
.A1(n_1278),
.A2(n_995),
.B1(n_1114),
.B2(n_1030),
.Y(n_1480)
);

INVx2_ASAP7_75t_SL g1481 ( 
.A(n_1223),
.Y(n_1481)
);

BUFx3_ASAP7_75t_L g1482 ( 
.A(n_1327),
.Y(n_1482)
);

BUFx6f_ASAP7_75t_L g1483 ( 
.A(n_1209),
.Y(n_1483)
);

BUFx2_ASAP7_75t_L g1484 ( 
.A(n_1262),
.Y(n_1484)
);

INVx2_ASAP7_75t_L g1485 ( 
.A(n_1277),
.Y(n_1485)
);

AOI22xp33_ASAP7_75t_SL g1486 ( 
.A1(n_1300),
.A2(n_1123),
.B1(n_1117),
.B2(n_995),
.Y(n_1486)
);

INVx3_ASAP7_75t_L g1487 ( 
.A(n_1214),
.Y(n_1487)
);

CKINVDCx5p33_ASAP7_75t_R g1488 ( 
.A(n_1341),
.Y(n_1488)
);

INVx4_ASAP7_75t_SL g1489 ( 
.A(n_1311),
.Y(n_1489)
);

AOI21x1_ASAP7_75t_L g1490 ( 
.A1(n_1286),
.A2(n_1033),
.B(n_1019),
.Y(n_1490)
);

AND2x2_ASAP7_75t_L g1491 ( 
.A(n_1227),
.B(n_1079),
.Y(n_1491)
);

INVx1_ASAP7_75t_L g1492 ( 
.A(n_1312),
.Y(n_1492)
);

BUFx3_ASAP7_75t_L g1493 ( 
.A(n_1338),
.Y(n_1493)
);

OAI22xp33_ASAP7_75t_L g1494 ( 
.A1(n_1193),
.A2(n_995),
.B1(n_1046),
.B2(n_1062),
.Y(n_1494)
);

BUFx2_ASAP7_75t_L g1495 ( 
.A(n_1262),
.Y(n_1495)
);

INVx3_ASAP7_75t_L g1496 ( 
.A(n_1214),
.Y(n_1496)
);

NAND2xp5_ASAP7_75t_L g1497 ( 
.A(n_1322),
.B(n_1131),
.Y(n_1497)
);

INVx1_ASAP7_75t_L g1498 ( 
.A(n_1318),
.Y(n_1498)
);

INVx2_ASAP7_75t_L g1499 ( 
.A(n_1277),
.Y(n_1499)
);

INVx6_ASAP7_75t_L g1500 ( 
.A(n_1234),
.Y(n_1500)
);

OR2x6_ASAP7_75t_L g1501 ( 
.A(n_1259),
.B(n_1026),
.Y(n_1501)
);

INVx3_ASAP7_75t_L g1502 ( 
.A(n_1214),
.Y(n_1502)
);

BUFx2_ASAP7_75t_L g1503 ( 
.A(n_1281),
.Y(n_1503)
);

INVx3_ASAP7_75t_L g1504 ( 
.A(n_1331),
.Y(n_1504)
);

INVx2_ASAP7_75t_L g1505 ( 
.A(n_1238),
.Y(n_1505)
);

HB1xp67_ASAP7_75t_L g1506 ( 
.A(n_1223),
.Y(n_1506)
);

AOI22xp33_ASAP7_75t_SL g1507 ( 
.A1(n_1247),
.A2(n_1123),
.B1(n_1117),
.B2(n_995),
.Y(n_1507)
);

INVx1_ASAP7_75t_L g1508 ( 
.A(n_1318),
.Y(n_1508)
);

INVx1_ASAP7_75t_L g1509 ( 
.A(n_1332),
.Y(n_1509)
);

INVx2_ASAP7_75t_L g1510 ( 
.A(n_1238),
.Y(n_1510)
);

AND2x2_ASAP7_75t_L g1511 ( 
.A(n_1227),
.B(n_1216),
.Y(n_1511)
);

INVx1_ASAP7_75t_L g1512 ( 
.A(n_1332),
.Y(n_1512)
);

INVx2_ASAP7_75t_SL g1513 ( 
.A(n_1227),
.Y(n_1513)
);

BUFx3_ASAP7_75t_L g1514 ( 
.A(n_1338),
.Y(n_1514)
);

INVx1_ASAP7_75t_L g1515 ( 
.A(n_1409),
.Y(n_1515)
);

NAND2xp5_ASAP7_75t_L g1516 ( 
.A(n_1355),
.B(n_1317),
.Y(n_1516)
);

INVx1_ASAP7_75t_SL g1517 ( 
.A(n_1412),
.Y(n_1517)
);

CKINVDCx5p33_ASAP7_75t_R g1518 ( 
.A(n_1356),
.Y(n_1518)
);

AOI22xp5_ASAP7_75t_L g1519 ( 
.A1(n_1442),
.A2(n_1232),
.B1(n_1293),
.B2(n_1441),
.Y(n_1519)
);

OR2x6_ASAP7_75t_L g1520 ( 
.A(n_1361),
.B(n_1344),
.Y(n_1520)
);

OR2x6_ASAP7_75t_L g1521 ( 
.A(n_1361),
.B(n_1344),
.Y(n_1521)
);

OA21x2_ASAP7_75t_L g1522 ( 
.A1(n_1433),
.A2(n_1287),
.B(n_1286),
.Y(n_1522)
);

OR2x2_ASAP7_75t_L g1523 ( 
.A(n_1355),
.B(n_1315),
.Y(n_1523)
);

INVx1_ASAP7_75t_L g1524 ( 
.A(n_1409),
.Y(n_1524)
);

INVx1_ASAP7_75t_L g1525 ( 
.A(n_1398),
.Y(n_1525)
);

NAND2xp5_ASAP7_75t_L g1526 ( 
.A(n_1368),
.B(n_1317),
.Y(n_1526)
);

OR2x6_ASAP7_75t_L g1527 ( 
.A(n_1500),
.B(n_1347),
.Y(n_1527)
);

INVx1_ASAP7_75t_L g1528 ( 
.A(n_1398),
.Y(n_1528)
);

AO31x2_ASAP7_75t_L g1529 ( 
.A1(n_1379),
.A2(n_1247),
.A3(n_1298),
.B(n_1306),
.Y(n_1529)
);

NOR2xp33_ASAP7_75t_R g1530 ( 
.A(n_1356),
.B(n_1199),
.Y(n_1530)
);

NOR2xp33_ASAP7_75t_R g1531 ( 
.A(n_1358),
.B(n_1204),
.Y(n_1531)
);

OR2x6_ASAP7_75t_L g1532 ( 
.A(n_1500),
.B(n_1347),
.Y(n_1532)
);

NAND2xp5_ASAP7_75t_L g1533 ( 
.A(n_1368),
.B(n_1272),
.Y(n_1533)
);

HB1xp67_ASAP7_75t_L g1534 ( 
.A(n_1397),
.Y(n_1534)
);

NOR2xp33_ASAP7_75t_R g1535 ( 
.A(n_1358),
.B(n_1204),
.Y(n_1535)
);

NAND3xp33_ASAP7_75t_SL g1536 ( 
.A(n_1442),
.B(n_1231),
.C(n_1266),
.Y(n_1536)
);

NAND3xp33_ASAP7_75t_SL g1537 ( 
.A(n_1441),
.B(n_1326),
.C(n_1265),
.Y(n_1537)
);

INVx2_ASAP7_75t_L g1538 ( 
.A(n_1362),
.Y(n_1538)
);

CKINVDCx5p33_ASAP7_75t_R g1539 ( 
.A(n_1430),
.Y(n_1539)
);

O2A1O1Ixp33_ASAP7_75t_SL g1540 ( 
.A1(n_1412),
.A2(n_1346),
.B(n_1310),
.C(n_1342),
.Y(n_1540)
);

INVx1_ASAP7_75t_L g1541 ( 
.A(n_1407),
.Y(n_1541)
);

CKINVDCx11_ASAP7_75t_R g1542 ( 
.A(n_1430),
.Y(n_1542)
);

BUFx2_ASAP7_75t_L g1543 ( 
.A(n_1432),
.Y(n_1543)
);

OR2x2_ASAP7_75t_L g1544 ( 
.A(n_1387),
.B(n_1315),
.Y(n_1544)
);

BUFx12f_ASAP7_75t_L g1545 ( 
.A(n_1430),
.Y(n_1545)
);

INVx2_ASAP7_75t_L g1546 ( 
.A(n_1362),
.Y(n_1546)
);

CKINVDCx20_ASAP7_75t_R g1547 ( 
.A(n_1428),
.Y(n_1547)
);

NOR2xp67_ASAP7_75t_L g1548 ( 
.A(n_1399),
.B(n_1352),
.Y(n_1548)
);

CKINVDCx20_ASAP7_75t_R g1549 ( 
.A(n_1428),
.Y(n_1549)
);

CKINVDCx8_ASAP7_75t_R g1550 ( 
.A(n_1488),
.Y(n_1550)
);

HB1xp67_ASAP7_75t_L g1551 ( 
.A(n_1397),
.Y(n_1551)
);

AOI22xp33_ASAP7_75t_L g1552 ( 
.A1(n_1371),
.A2(n_1271),
.B1(n_1200),
.B2(n_1322),
.Y(n_1552)
);

BUFx6f_ASAP7_75t_L g1553 ( 
.A(n_1373),
.Y(n_1553)
);

INVx2_ASAP7_75t_L g1554 ( 
.A(n_1362),
.Y(n_1554)
);

AND2x2_ASAP7_75t_L g1555 ( 
.A(n_1511),
.B(n_1296),
.Y(n_1555)
);

OAI22xp5_ASAP7_75t_L g1556 ( 
.A1(n_1425),
.A2(n_1326),
.B1(n_1219),
.B2(n_1337),
.Y(n_1556)
);

OR2x2_ASAP7_75t_L g1557 ( 
.A(n_1387),
.B(n_1296),
.Y(n_1557)
);

NOR2x1_ASAP7_75t_L g1558 ( 
.A(n_1432),
.B(n_1340),
.Y(n_1558)
);

OAI21xp5_ASAP7_75t_SL g1559 ( 
.A1(n_1480),
.A2(n_1245),
.B(n_1219),
.Y(n_1559)
);

INVx1_ASAP7_75t_L g1560 ( 
.A(n_1407),
.Y(n_1560)
);

NOR2xp33_ASAP7_75t_R g1561 ( 
.A(n_1428),
.B(n_996),
.Y(n_1561)
);

INVx1_ASAP7_75t_L g1562 ( 
.A(n_1451),
.Y(n_1562)
);

NOR2x1p5_ASAP7_75t_L g1563 ( 
.A(n_1432),
.B(n_1062),
.Y(n_1563)
);

AND2x4_ASAP7_75t_L g1564 ( 
.A(n_1513),
.B(n_1287),
.Y(n_1564)
);

NOR2x1_ASAP7_75t_L g1565 ( 
.A(n_1453),
.B(n_1340),
.Y(n_1565)
);

INVx2_ASAP7_75t_L g1566 ( 
.A(n_1385),
.Y(n_1566)
);

AND2x2_ASAP7_75t_L g1567 ( 
.A(n_1511),
.B(n_1367),
.Y(n_1567)
);

INVx1_ASAP7_75t_L g1568 ( 
.A(n_1451),
.Y(n_1568)
);

NAND2xp5_ASAP7_75t_L g1569 ( 
.A(n_1468),
.B(n_1346),
.Y(n_1569)
);

INVx4_ASAP7_75t_SL g1570 ( 
.A(n_1500),
.Y(n_1570)
);

OR2x2_ASAP7_75t_L g1571 ( 
.A(n_1384),
.B(n_1343),
.Y(n_1571)
);

BUFx6f_ASAP7_75t_L g1572 ( 
.A(n_1373),
.Y(n_1572)
);

CKINVDCx16_ASAP7_75t_R g1573 ( 
.A(n_1452),
.Y(n_1573)
);

NOR2xp33_ASAP7_75t_L g1574 ( 
.A(n_1494),
.B(n_1236),
.Y(n_1574)
);

AO21x2_ASAP7_75t_L g1575 ( 
.A1(n_1379),
.A2(n_1200),
.B(n_1328),
.Y(n_1575)
);

INVx3_ASAP7_75t_L g1576 ( 
.A(n_1453),
.Y(n_1576)
);

INVx1_ASAP7_75t_L g1577 ( 
.A(n_1454),
.Y(n_1577)
);

AOI22xp33_ASAP7_75t_L g1578 ( 
.A1(n_1371),
.A2(n_1322),
.B1(n_1216),
.B2(n_1303),
.Y(n_1578)
);

BUFx2_ASAP7_75t_L g1579 ( 
.A(n_1453),
.Y(n_1579)
);

AOI22xp33_ASAP7_75t_L g1580 ( 
.A1(n_1423),
.A2(n_1291),
.B1(n_1255),
.B2(n_1311),
.Y(n_1580)
);

INVx1_ASAP7_75t_L g1581 ( 
.A(n_1454),
.Y(n_1581)
);

HB1xp67_ASAP7_75t_L g1582 ( 
.A(n_1426),
.Y(n_1582)
);

AND2x2_ASAP7_75t_SL g1583 ( 
.A(n_1449),
.B(n_1295),
.Y(n_1583)
);

NAND2xp33_ASAP7_75t_SL g1584 ( 
.A(n_1472),
.B(n_1000),
.Y(n_1584)
);

INVx1_ASAP7_75t_L g1585 ( 
.A(n_1456),
.Y(n_1585)
);

OR2x6_ASAP7_75t_L g1586 ( 
.A(n_1500),
.B(n_1336),
.Y(n_1586)
);

OAI21xp5_ASAP7_75t_SL g1587 ( 
.A1(n_1480),
.A2(n_1319),
.B(n_1316),
.Y(n_1587)
);

AND2x2_ASAP7_75t_L g1588 ( 
.A(n_1511),
.B(n_1324),
.Y(n_1588)
);

NAND2xp5_ASAP7_75t_L g1589 ( 
.A(n_1468),
.B(n_1281),
.Y(n_1589)
);

AND2x2_ASAP7_75t_L g1590 ( 
.A(n_1367),
.B(n_1324),
.Y(n_1590)
);

AND2x2_ASAP7_75t_L g1591 ( 
.A(n_1367),
.B(n_1330),
.Y(n_1591)
);

INVx2_ASAP7_75t_L g1592 ( 
.A(n_1385),
.Y(n_1592)
);

INVx4_ASAP7_75t_L g1593 ( 
.A(n_1448),
.Y(n_1593)
);

INVxp67_ASAP7_75t_L g1594 ( 
.A(n_1484),
.Y(n_1594)
);

NAND2xp5_ASAP7_75t_L g1595 ( 
.A(n_1456),
.B(n_1330),
.Y(n_1595)
);

NAND2xp5_ASAP7_75t_L g1596 ( 
.A(n_1459),
.B(n_1343),
.Y(n_1596)
);

AND2x2_ASAP7_75t_L g1597 ( 
.A(n_1369),
.B(n_1348),
.Y(n_1597)
);

NOR2xp33_ASAP7_75t_R g1598 ( 
.A(n_1463),
.B(n_997),
.Y(n_1598)
);

INVxp67_ASAP7_75t_L g1599 ( 
.A(n_1484),
.Y(n_1599)
);

AOI22xp33_ASAP7_75t_L g1600 ( 
.A1(n_1423),
.A2(n_1255),
.B1(n_1311),
.B2(n_1329),
.Y(n_1600)
);

NOR2x1p5_ASAP7_75t_L g1601 ( 
.A(n_1514),
.B(n_1036),
.Y(n_1601)
);

BUFx3_ASAP7_75t_L g1602 ( 
.A(n_1463),
.Y(n_1602)
);

AOI22xp33_ASAP7_75t_L g1603 ( 
.A1(n_1423),
.A2(n_1311),
.B1(n_1336),
.B2(n_1295),
.Y(n_1603)
);

NAND2xp5_ASAP7_75t_L g1604 ( 
.A(n_1459),
.B(n_1249),
.Y(n_1604)
);

INVx1_ASAP7_75t_L g1605 ( 
.A(n_1440),
.Y(n_1605)
);

INVx1_ASAP7_75t_L g1606 ( 
.A(n_1440),
.Y(n_1606)
);

NAND2xp5_ASAP7_75t_L g1607 ( 
.A(n_1467),
.B(n_1249),
.Y(n_1607)
);

INVx2_ASAP7_75t_L g1608 ( 
.A(n_1385),
.Y(n_1608)
);

OR2x6_ASAP7_75t_L g1609 ( 
.A(n_1500),
.B(n_1336),
.Y(n_1609)
);

INVx1_ASAP7_75t_L g1610 ( 
.A(n_1444),
.Y(n_1610)
);

NOR2xp33_ASAP7_75t_R g1611 ( 
.A(n_1500),
.B(n_1052),
.Y(n_1611)
);

INVxp67_ASAP7_75t_L g1612 ( 
.A(n_1484),
.Y(n_1612)
);

OR2x2_ASAP7_75t_L g1613 ( 
.A(n_1384),
.B(n_1244),
.Y(n_1613)
);

NAND2xp33_ASAP7_75t_R g1614 ( 
.A(n_1449),
.B(n_1475),
.Y(n_1614)
);

AND2x2_ASAP7_75t_L g1615 ( 
.A(n_1369),
.B(n_1348),
.Y(n_1615)
);

CKINVDCx5p33_ASAP7_75t_R g1616 ( 
.A(n_1452),
.Y(n_1616)
);

INVx5_ASAP7_75t_SL g1617 ( 
.A(n_1448),
.Y(n_1617)
);

INVxp67_ASAP7_75t_L g1618 ( 
.A(n_1495),
.Y(n_1618)
);

AND2x2_ASAP7_75t_L g1619 ( 
.A(n_1369),
.B(n_1391),
.Y(n_1619)
);

BUFx3_ASAP7_75t_L g1620 ( 
.A(n_1463),
.Y(n_1620)
);

OAI21x1_ASAP7_75t_L g1621 ( 
.A1(n_1476),
.A2(n_1351),
.B(n_1339),
.Y(n_1621)
);

CKINVDCx16_ASAP7_75t_R g1622 ( 
.A(n_1482),
.Y(n_1622)
);

OAI22xp5_ASAP7_75t_L g1623 ( 
.A1(n_1425),
.A2(n_1254),
.B1(n_1207),
.B2(n_1226),
.Y(n_1623)
);

CKINVDCx5p33_ASAP7_75t_R g1624 ( 
.A(n_1482),
.Y(n_1624)
);

INVx2_ASAP7_75t_L g1625 ( 
.A(n_1386),
.Y(n_1625)
);

INVx1_ASAP7_75t_SL g1626 ( 
.A(n_1482),
.Y(n_1626)
);

NAND2xp5_ASAP7_75t_SL g1627 ( 
.A(n_1494),
.B(n_1323),
.Y(n_1627)
);

AOI22xp33_ASAP7_75t_L g1628 ( 
.A1(n_1423),
.A2(n_1336),
.B1(n_1220),
.B2(n_1123),
.Y(n_1628)
);

INVx2_ASAP7_75t_L g1629 ( 
.A(n_1386),
.Y(n_1629)
);

AND2x2_ASAP7_75t_L g1630 ( 
.A(n_1391),
.B(n_1288),
.Y(n_1630)
);

INVx2_ASAP7_75t_L g1631 ( 
.A(n_1386),
.Y(n_1631)
);

INVx2_ASAP7_75t_SL g1632 ( 
.A(n_1493),
.Y(n_1632)
);

AND2x2_ASAP7_75t_L g1633 ( 
.A(n_1391),
.B(n_1288),
.Y(n_1633)
);

NAND2xp5_ASAP7_75t_L g1634 ( 
.A(n_1467),
.B(n_1249),
.Y(n_1634)
);

INVx1_ASAP7_75t_L g1635 ( 
.A(n_1444),
.Y(n_1635)
);

HB1xp67_ASAP7_75t_L g1636 ( 
.A(n_1426),
.Y(n_1636)
);

INVx2_ASAP7_75t_L g1637 ( 
.A(n_1390),
.Y(n_1637)
);

OAI22xp5_ASAP7_75t_L g1638 ( 
.A1(n_1462),
.A2(n_1472),
.B1(n_1457),
.B2(n_1448),
.Y(n_1638)
);

INVx1_ASAP7_75t_L g1639 ( 
.A(n_1359),
.Y(n_1639)
);

HB1xp67_ASAP7_75t_L g1640 ( 
.A(n_1399),
.Y(n_1640)
);

INVx1_ASAP7_75t_L g1641 ( 
.A(n_1359),
.Y(n_1641)
);

OR2x2_ASAP7_75t_L g1642 ( 
.A(n_1384),
.B(n_1244),
.Y(n_1642)
);

NAND2xp33_ASAP7_75t_R g1643 ( 
.A(n_1449),
.B(n_1336),
.Y(n_1643)
);

NOR2xp33_ASAP7_75t_R g1644 ( 
.A(n_1490),
.B(n_1060),
.Y(n_1644)
);

AO31x2_ASAP7_75t_L g1645 ( 
.A1(n_1380),
.A2(n_1299),
.A3(n_1297),
.B(n_1298),
.Y(n_1645)
);

INVx2_ASAP7_75t_L g1646 ( 
.A(n_1390),
.Y(n_1646)
);

NAND2xp5_ASAP7_75t_L g1647 ( 
.A(n_1497),
.B(n_1284),
.Y(n_1647)
);

HB1xp67_ASAP7_75t_L g1648 ( 
.A(n_1399),
.Y(n_1648)
);

INVx1_ASAP7_75t_L g1649 ( 
.A(n_1359),
.Y(n_1649)
);

NAND2xp33_ASAP7_75t_R g1650 ( 
.A(n_1449),
.B(n_1257),
.Y(n_1650)
);

INVx1_ASAP7_75t_L g1651 ( 
.A(n_1360),
.Y(n_1651)
);

NAND2xp33_ASAP7_75t_R g1652 ( 
.A(n_1449),
.B(n_1257),
.Y(n_1652)
);

INVx1_ASAP7_75t_L g1653 ( 
.A(n_1360),
.Y(n_1653)
);

AOI22xp5_ASAP7_75t_L g1654 ( 
.A1(n_1457),
.A2(n_1217),
.B1(n_1306),
.B2(n_1309),
.Y(n_1654)
);

AND2x4_ASAP7_75t_L g1655 ( 
.A(n_1513),
.B(n_1288),
.Y(n_1655)
);

OR2x2_ASAP7_75t_L g1656 ( 
.A(n_1497),
.B(n_1269),
.Y(n_1656)
);

AOI222xp33_ASAP7_75t_L g1657 ( 
.A1(n_1433),
.A2(n_1234),
.B1(n_1269),
.B2(n_1274),
.C1(n_1297),
.C2(n_1309),
.Y(n_1657)
);

NAND2xp33_ASAP7_75t_L g1658 ( 
.A(n_1373),
.B(n_1060),
.Y(n_1658)
);

INVx3_ASAP7_75t_L g1659 ( 
.A(n_1493),
.Y(n_1659)
);

CKINVDCx16_ASAP7_75t_R g1660 ( 
.A(n_1493),
.Y(n_1660)
);

INVx1_ASAP7_75t_L g1661 ( 
.A(n_1360),
.Y(n_1661)
);

OR2x2_ASAP7_75t_L g1662 ( 
.A(n_1495),
.B(n_1274),
.Y(n_1662)
);

NAND2xp5_ASAP7_75t_L g1663 ( 
.A(n_1514),
.B(n_1284),
.Y(n_1663)
);

INVx2_ASAP7_75t_L g1664 ( 
.A(n_1390),
.Y(n_1664)
);

INVx1_ASAP7_75t_SL g1665 ( 
.A(n_1514),
.Y(n_1665)
);

AOI21xp33_ASAP7_75t_L g1666 ( 
.A1(n_1481),
.A2(n_1299),
.B(n_1283),
.Y(n_1666)
);

HB1xp67_ASAP7_75t_L g1667 ( 
.A(n_1439),
.Y(n_1667)
);

INVx8_ASAP7_75t_L g1668 ( 
.A(n_1448),
.Y(n_1668)
);

CKINVDCx5p33_ASAP7_75t_R g1669 ( 
.A(n_1445),
.Y(n_1669)
);

NAND2xp5_ASAP7_75t_L g1670 ( 
.A(n_1434),
.B(n_1284),
.Y(n_1670)
);

INVx2_ASAP7_75t_SL g1671 ( 
.A(n_1445),
.Y(n_1671)
);

INVx2_ASAP7_75t_L g1672 ( 
.A(n_1414),
.Y(n_1672)
);

AO31x2_ASAP7_75t_L g1673 ( 
.A1(n_1380),
.A2(n_1314),
.A3(n_1321),
.B(n_1294),
.Y(n_1673)
);

CKINVDCx5p33_ASAP7_75t_R g1674 ( 
.A(n_1445),
.Y(n_1674)
);

CKINVDCx5p33_ASAP7_75t_R g1675 ( 
.A(n_1445),
.Y(n_1675)
);

NAND2xp5_ASAP7_75t_L g1676 ( 
.A(n_1434),
.B(n_1292),
.Y(n_1676)
);

INVx2_ASAP7_75t_L g1677 ( 
.A(n_1414),
.Y(n_1677)
);

HB1xp67_ASAP7_75t_L g1678 ( 
.A(n_1439),
.Y(n_1678)
);

NOR2xp33_ASAP7_75t_R g1679 ( 
.A(n_1490),
.B(n_1063),
.Y(n_1679)
);

AND2x2_ASAP7_75t_L g1680 ( 
.A(n_1474),
.B(n_1288),
.Y(n_1680)
);

OAI21xp33_ASAP7_75t_L g1681 ( 
.A1(n_1404),
.A2(n_1292),
.B(n_1220),
.Y(n_1681)
);

INVx1_ASAP7_75t_L g1682 ( 
.A(n_1363),
.Y(n_1682)
);

AND2x2_ASAP7_75t_L g1683 ( 
.A(n_1474),
.B(n_1234),
.Y(n_1683)
);

OR2x2_ASAP7_75t_SL g1684 ( 
.A(n_1393),
.B(n_1207),
.Y(n_1684)
);

NOR2xp33_ASAP7_75t_R g1685 ( 
.A(n_1446),
.B(n_1009),
.Y(n_1685)
);

HB1xp67_ASAP7_75t_L g1686 ( 
.A(n_1439),
.Y(n_1686)
);

INVx1_ASAP7_75t_L g1687 ( 
.A(n_1363),
.Y(n_1687)
);

AOI22xp33_ASAP7_75t_L g1688 ( 
.A1(n_1404),
.A2(n_1123),
.B1(n_1290),
.B2(n_1294),
.Y(n_1688)
);

NAND2xp33_ASAP7_75t_R g1689 ( 
.A(n_1475),
.B(n_1257),
.Y(n_1689)
);

INVx1_ASAP7_75t_L g1690 ( 
.A(n_1363),
.Y(n_1690)
);

NAND2xp33_ASAP7_75t_L g1691 ( 
.A(n_1373),
.B(n_1039),
.Y(n_1691)
);

BUFx2_ASAP7_75t_L g1692 ( 
.A(n_1495),
.Y(n_1692)
);

CKINVDCx11_ASAP7_75t_R g1693 ( 
.A(n_1393),
.Y(n_1693)
);

INVx2_ASAP7_75t_L g1694 ( 
.A(n_1414),
.Y(n_1694)
);

NOR2xp33_ASAP7_75t_R g1695 ( 
.A(n_1446),
.B(n_1009),
.Y(n_1695)
);

INVx1_ASAP7_75t_L g1696 ( 
.A(n_1365),
.Y(n_1696)
);

AOI222xp33_ASAP7_75t_L g1697 ( 
.A1(n_1404),
.A2(n_1234),
.B1(n_1283),
.B2(n_1321),
.C1(n_1290),
.C2(n_1314),
.Y(n_1697)
);

INVx2_ASAP7_75t_SL g1698 ( 
.A(n_1445),
.Y(n_1698)
);

INVx1_ASAP7_75t_L g1699 ( 
.A(n_1365),
.Y(n_1699)
);

HB1xp67_ASAP7_75t_L g1700 ( 
.A(n_1415),
.Y(n_1700)
);

AND2x4_ASAP7_75t_L g1701 ( 
.A(n_1513),
.B(n_1257),
.Y(n_1701)
);

BUFx3_ASAP7_75t_L g1702 ( 
.A(n_1455),
.Y(n_1702)
);

OAI22xp5_ASAP7_75t_L g1703 ( 
.A1(n_1462),
.A2(n_1254),
.B1(n_1207),
.B2(n_1115),
.Y(n_1703)
);

INVx1_ASAP7_75t_L g1704 ( 
.A(n_1365),
.Y(n_1704)
);

BUFx6f_ASAP7_75t_L g1705 ( 
.A(n_1373),
.Y(n_1705)
);

INVx4_ASAP7_75t_L g1706 ( 
.A(n_1448),
.Y(n_1706)
);

OR2x2_ASAP7_75t_L g1707 ( 
.A(n_1503),
.B(n_1333),
.Y(n_1707)
);

INVx1_ASAP7_75t_L g1708 ( 
.A(n_1436),
.Y(n_1708)
);

INVx1_ASAP7_75t_L g1709 ( 
.A(n_1436),
.Y(n_1709)
);

AND2x2_ASAP7_75t_L g1710 ( 
.A(n_1474),
.B(n_1349),
.Y(n_1710)
);

OR2x6_ASAP7_75t_L g1711 ( 
.A(n_1383),
.B(n_1270),
.Y(n_1711)
);

OR2x6_ASAP7_75t_L g1712 ( 
.A(n_1383),
.B(n_1270),
.Y(n_1712)
);

NOR3xp33_ASAP7_75t_SL g1713 ( 
.A(n_1437),
.B(n_1030),
.C(n_1009),
.Y(n_1713)
);

NOR2xp33_ASAP7_75t_L g1714 ( 
.A(n_1503),
.B(n_1305),
.Y(n_1714)
);

NAND2xp5_ASAP7_75t_L g1715 ( 
.A(n_1437),
.B(n_1292),
.Y(n_1715)
);

AO31x2_ASAP7_75t_L g1716 ( 
.A1(n_1381),
.A2(n_1333),
.A3(n_1353),
.B(n_1349),
.Y(n_1716)
);

AND2x2_ASAP7_75t_L g1717 ( 
.A(n_1491),
.B(n_1353),
.Y(n_1717)
);

NAND2xp5_ASAP7_75t_L g1718 ( 
.A(n_1438),
.B(n_1264),
.Y(n_1718)
);

AND2x2_ASAP7_75t_L g1719 ( 
.A(n_1491),
.B(n_1334),
.Y(n_1719)
);

OAI22xp33_ASAP7_75t_L g1720 ( 
.A1(n_1448),
.A2(n_1270),
.B1(n_1320),
.B2(n_1301),
.Y(n_1720)
);

CKINVDCx16_ASAP7_75t_R g1721 ( 
.A(n_1491),
.Y(n_1721)
);

BUFx3_ASAP7_75t_L g1722 ( 
.A(n_1455),
.Y(n_1722)
);

AND2x2_ASAP7_75t_L g1723 ( 
.A(n_1366),
.B(n_1351),
.Y(n_1723)
);

OR2x6_ASAP7_75t_L g1724 ( 
.A(n_1501),
.B(n_1260),
.Y(n_1724)
);

CKINVDCx5p33_ASAP7_75t_R g1725 ( 
.A(n_1503),
.Y(n_1725)
);

AND2x2_ASAP7_75t_L g1726 ( 
.A(n_1366),
.B(n_1350),
.Y(n_1726)
);

INVx1_ASAP7_75t_L g1727 ( 
.A(n_1438),
.Y(n_1727)
);

NOR2xp33_ASAP7_75t_L g1728 ( 
.A(n_1417),
.B(n_1254),
.Y(n_1728)
);

INVx2_ASAP7_75t_SL g1729 ( 
.A(n_1455),
.Y(n_1729)
);

AND2x4_ASAP7_75t_L g1730 ( 
.A(n_1489),
.B(n_1260),
.Y(n_1730)
);

AOI21xp5_ASAP7_75t_L g1731 ( 
.A1(n_1402),
.A2(n_1320),
.B(n_1225),
.Y(n_1731)
);

AO21x1_ASAP7_75t_L g1732 ( 
.A1(n_1424),
.A2(n_1331),
.B(n_1345),
.Y(n_1732)
);

INVx1_ASAP7_75t_L g1733 ( 
.A(n_1461),
.Y(n_1733)
);

INVx2_ASAP7_75t_L g1734 ( 
.A(n_1421),
.Y(n_1734)
);

INVx1_ASAP7_75t_L g1735 ( 
.A(n_1639),
.Y(n_1735)
);

NOR2xp33_ASAP7_75t_L g1736 ( 
.A(n_1550),
.B(n_1518),
.Y(n_1736)
);

INVx2_ASAP7_75t_SL g1737 ( 
.A(n_1662),
.Y(n_1737)
);

NOR2xp33_ASAP7_75t_L g1738 ( 
.A(n_1539),
.B(n_1693),
.Y(n_1738)
);

INVx2_ASAP7_75t_L g1739 ( 
.A(n_1645),
.Y(n_1739)
);

INVx1_ASAP7_75t_L g1740 ( 
.A(n_1641),
.Y(n_1740)
);

INVxp67_ASAP7_75t_L g1741 ( 
.A(n_1516),
.Y(n_1741)
);

INVx2_ASAP7_75t_L g1742 ( 
.A(n_1645),
.Y(n_1742)
);

OR2x2_ASAP7_75t_L g1743 ( 
.A(n_1523),
.B(n_1415),
.Y(n_1743)
);

INVx2_ASAP7_75t_L g1744 ( 
.A(n_1645),
.Y(n_1744)
);

BUFx2_ASAP7_75t_L g1745 ( 
.A(n_1684),
.Y(n_1745)
);

INVx1_ASAP7_75t_L g1746 ( 
.A(n_1649),
.Y(n_1746)
);

BUFx6f_ASAP7_75t_L g1747 ( 
.A(n_1542),
.Y(n_1747)
);

AOI22xp33_ASAP7_75t_SL g1748 ( 
.A1(n_1573),
.A2(n_1415),
.B1(n_1418),
.B2(n_1416),
.Y(n_1748)
);

INVx1_ASAP7_75t_L g1749 ( 
.A(n_1651),
.Y(n_1749)
);

AND2x2_ASAP7_75t_L g1750 ( 
.A(n_1721),
.B(n_1376),
.Y(n_1750)
);

INVx1_ASAP7_75t_L g1751 ( 
.A(n_1653),
.Y(n_1751)
);

OAI21xp5_ASAP7_75t_L g1752 ( 
.A1(n_1559),
.A2(n_1574),
.B(n_1536),
.Y(n_1752)
);

OA21x2_ASAP7_75t_L g1753 ( 
.A1(n_1681),
.A2(n_1395),
.B(n_1394),
.Y(n_1753)
);

INVx1_ASAP7_75t_L g1754 ( 
.A(n_1661),
.Y(n_1754)
);

AND2x2_ASAP7_75t_L g1755 ( 
.A(n_1567),
.B(n_1376),
.Y(n_1755)
);

INVx2_ASAP7_75t_L g1756 ( 
.A(n_1645),
.Y(n_1756)
);

AND2x2_ASAP7_75t_L g1757 ( 
.A(n_1726),
.B(n_1376),
.Y(n_1757)
);

INVx2_ASAP7_75t_L g1758 ( 
.A(n_1640),
.Y(n_1758)
);

INVx1_ASAP7_75t_L g1759 ( 
.A(n_1682),
.Y(n_1759)
);

INVx1_ASAP7_75t_L g1760 ( 
.A(n_1687),
.Y(n_1760)
);

BUFx4f_ASAP7_75t_L g1761 ( 
.A(n_1545),
.Y(n_1761)
);

INVxp67_ASAP7_75t_SL g1762 ( 
.A(n_1614),
.Y(n_1762)
);

NAND4xp25_ASAP7_75t_SL g1763 ( 
.A(n_1547),
.B(n_1366),
.C(n_1486),
.D(n_1507),
.Y(n_1763)
);

BUFx6f_ASAP7_75t_L g1764 ( 
.A(n_1553),
.Y(n_1764)
);

NAND2xp5_ASAP7_75t_L g1765 ( 
.A(n_1533),
.B(n_1461),
.Y(n_1765)
);

AND2x2_ASAP7_75t_L g1766 ( 
.A(n_1723),
.B(n_1376),
.Y(n_1766)
);

AND2x2_ASAP7_75t_L g1767 ( 
.A(n_1619),
.B(n_1555),
.Y(n_1767)
);

BUFx3_ASAP7_75t_L g1768 ( 
.A(n_1549),
.Y(n_1768)
);

AND2x2_ASAP7_75t_L g1769 ( 
.A(n_1588),
.B(n_1376),
.Y(n_1769)
);

HB1xp67_ASAP7_75t_L g1770 ( 
.A(n_1594),
.Y(n_1770)
);

AND2x2_ASAP7_75t_L g1771 ( 
.A(n_1692),
.B(n_1400),
.Y(n_1771)
);

INVx2_ASAP7_75t_L g1772 ( 
.A(n_1640),
.Y(n_1772)
);

AND2x2_ASAP7_75t_L g1773 ( 
.A(n_1630),
.B(n_1400),
.Y(n_1773)
);

INVx2_ASAP7_75t_SL g1774 ( 
.A(n_1707),
.Y(n_1774)
);

AND2x2_ASAP7_75t_L g1775 ( 
.A(n_1633),
.B(n_1400),
.Y(n_1775)
);

INVx2_ASAP7_75t_L g1776 ( 
.A(n_1648),
.Y(n_1776)
);

INVx1_ASAP7_75t_L g1777 ( 
.A(n_1690),
.Y(n_1777)
);

OAI22xp33_ASAP7_75t_L g1778 ( 
.A1(n_1519),
.A2(n_1418),
.B1(n_1416),
.B2(n_1446),
.Y(n_1778)
);

AND2x2_ASAP7_75t_L g1779 ( 
.A(n_1702),
.B(n_1400),
.Y(n_1779)
);

INVx1_ASAP7_75t_L g1780 ( 
.A(n_1696),
.Y(n_1780)
);

AND2x2_ASAP7_75t_L g1781 ( 
.A(n_1722),
.B(n_1400),
.Y(n_1781)
);

OAI221xp5_ASAP7_75t_L g1782 ( 
.A1(n_1580),
.A2(n_1418),
.B1(n_1416),
.B2(n_1486),
.C(n_1354),
.Y(n_1782)
);

INVx2_ASAP7_75t_L g1783 ( 
.A(n_1648),
.Y(n_1783)
);

OR2x6_ASAP7_75t_L g1784 ( 
.A(n_1520),
.B(n_1427),
.Y(n_1784)
);

INVx2_ASAP7_75t_L g1785 ( 
.A(n_1667),
.Y(n_1785)
);

NAND2xp5_ASAP7_75t_L g1786 ( 
.A(n_1574),
.B(n_1464),
.Y(n_1786)
);

AND2x4_ASAP7_75t_L g1787 ( 
.A(n_1570),
.B(n_1489),
.Y(n_1787)
);

NOR2x1_ASAP7_75t_SL g1788 ( 
.A(n_1711),
.B(n_1501),
.Y(n_1788)
);

INVx1_ASAP7_75t_L g1789 ( 
.A(n_1699),
.Y(n_1789)
);

INVx2_ASAP7_75t_L g1790 ( 
.A(n_1667),
.Y(n_1790)
);

INVx1_ASAP7_75t_L g1791 ( 
.A(n_1704),
.Y(n_1791)
);

BUFx3_ASAP7_75t_L g1792 ( 
.A(n_1624),
.Y(n_1792)
);

INVx1_ASAP7_75t_L g1793 ( 
.A(n_1605),
.Y(n_1793)
);

AND2x2_ASAP7_75t_L g1794 ( 
.A(n_1622),
.B(n_1410),
.Y(n_1794)
);

OR2x2_ASAP7_75t_L g1795 ( 
.A(n_1544),
.B(n_1505),
.Y(n_1795)
);

OR2x2_ASAP7_75t_L g1796 ( 
.A(n_1656),
.B(n_1505),
.Y(n_1796)
);

NAND2xp5_ASAP7_75t_L g1797 ( 
.A(n_1526),
.B(n_1464),
.Y(n_1797)
);

AND2x2_ASAP7_75t_L g1798 ( 
.A(n_1660),
.B(n_1410),
.Y(n_1798)
);

INVx2_ASAP7_75t_L g1799 ( 
.A(n_1678),
.Y(n_1799)
);

AND2x2_ASAP7_75t_L g1800 ( 
.A(n_1680),
.B(n_1410),
.Y(n_1800)
);

INVx1_ASAP7_75t_L g1801 ( 
.A(n_1606),
.Y(n_1801)
);

INVx1_ASAP7_75t_L g1802 ( 
.A(n_1610),
.Y(n_1802)
);

INVx4_ASAP7_75t_L g1803 ( 
.A(n_1711),
.Y(n_1803)
);

AND2x2_ASAP7_75t_L g1804 ( 
.A(n_1671),
.B(n_1410),
.Y(n_1804)
);

AND2x2_ASAP7_75t_L g1805 ( 
.A(n_1698),
.B(n_1410),
.Y(n_1805)
);

INVx2_ASAP7_75t_SL g1806 ( 
.A(n_1602),
.Y(n_1806)
);

NOR2x1p5_ASAP7_75t_L g1807 ( 
.A(n_1536),
.B(n_1422),
.Y(n_1807)
);

CKINVDCx14_ASAP7_75t_R g1808 ( 
.A(n_1530),
.Y(n_1808)
);

AND2x2_ASAP7_75t_L g1809 ( 
.A(n_1590),
.B(n_1422),
.Y(n_1809)
);

INVx1_ASAP7_75t_L g1810 ( 
.A(n_1635),
.Y(n_1810)
);

INVx2_ASAP7_75t_L g1811 ( 
.A(n_1678),
.Y(n_1811)
);

AND2x2_ASAP7_75t_L g1812 ( 
.A(n_1591),
.B(n_1422),
.Y(n_1812)
);

AND2x2_ASAP7_75t_L g1813 ( 
.A(n_1725),
.B(n_1422),
.Y(n_1813)
);

INVx2_ASAP7_75t_L g1814 ( 
.A(n_1686),
.Y(n_1814)
);

AND2x2_ASAP7_75t_L g1815 ( 
.A(n_1729),
.B(n_1422),
.Y(n_1815)
);

HB1xp67_ASAP7_75t_L g1816 ( 
.A(n_1594),
.Y(n_1816)
);

INVx1_ASAP7_75t_L g1817 ( 
.A(n_1708),
.Y(n_1817)
);

INVx2_ASAP7_75t_L g1818 ( 
.A(n_1686),
.Y(n_1818)
);

INVx2_ASAP7_75t_SL g1819 ( 
.A(n_1620),
.Y(n_1819)
);

AND2x2_ASAP7_75t_L g1820 ( 
.A(n_1655),
.B(n_1478),
.Y(n_1820)
);

INVx5_ASAP7_75t_SL g1821 ( 
.A(n_1711),
.Y(n_1821)
);

HB1xp67_ASAP7_75t_L g1822 ( 
.A(n_1599),
.Y(n_1822)
);

INVxp67_ASAP7_75t_SL g1823 ( 
.A(n_1614),
.Y(n_1823)
);

NOR2x1_ASAP7_75t_R g1824 ( 
.A(n_1616),
.B(n_1254),
.Y(n_1824)
);

HB1xp67_ASAP7_75t_L g1825 ( 
.A(n_1599),
.Y(n_1825)
);

AND2x4_ASAP7_75t_L g1826 ( 
.A(n_1570),
.B(n_1489),
.Y(n_1826)
);

NAND2xp5_ASAP7_75t_L g1827 ( 
.A(n_1589),
.B(n_1569),
.Y(n_1827)
);

INVx1_ASAP7_75t_L g1828 ( 
.A(n_1709),
.Y(n_1828)
);

AND2x2_ASAP7_75t_L g1829 ( 
.A(n_1655),
.B(n_1478),
.Y(n_1829)
);

OR2x2_ASAP7_75t_L g1830 ( 
.A(n_1557),
.B(n_1505),
.Y(n_1830)
);

OR2x2_ASAP7_75t_L g1831 ( 
.A(n_1595),
.B(n_1510),
.Y(n_1831)
);

INVxp67_ASAP7_75t_SL g1832 ( 
.A(n_1689),
.Y(n_1832)
);

AND2x2_ASAP7_75t_L g1833 ( 
.A(n_1543),
.B(n_1478),
.Y(n_1833)
);

AND2x4_ASAP7_75t_L g1834 ( 
.A(n_1570),
.B(n_1489),
.Y(n_1834)
);

AOI22xp33_ASAP7_75t_L g1835 ( 
.A1(n_1552),
.A2(n_1411),
.B1(n_1424),
.B2(n_1370),
.Y(n_1835)
);

INVx3_ASAP7_75t_L g1836 ( 
.A(n_1553),
.Y(n_1836)
);

INVx1_ASAP7_75t_L g1837 ( 
.A(n_1727),
.Y(n_1837)
);

BUFx2_ASAP7_75t_L g1838 ( 
.A(n_1644),
.Y(n_1838)
);

AND2x2_ASAP7_75t_L g1839 ( 
.A(n_1579),
.B(n_1478),
.Y(n_1839)
);

INVx1_ASAP7_75t_L g1840 ( 
.A(n_1733),
.Y(n_1840)
);

INVx2_ASAP7_75t_L g1841 ( 
.A(n_1673),
.Y(n_1841)
);

AND2x4_ASAP7_75t_L g1842 ( 
.A(n_1730),
.B(n_1489),
.Y(n_1842)
);

AND2x2_ASAP7_75t_L g1843 ( 
.A(n_1710),
.B(n_1478),
.Y(n_1843)
);

INVx1_ASAP7_75t_L g1844 ( 
.A(n_1525),
.Y(n_1844)
);

AND2x2_ASAP7_75t_L g1845 ( 
.A(n_1717),
.B(n_1487),
.Y(n_1845)
);

HB1xp67_ASAP7_75t_L g1846 ( 
.A(n_1612),
.Y(n_1846)
);

AND2x2_ASAP7_75t_L g1847 ( 
.A(n_1597),
.B(n_1487),
.Y(n_1847)
);

INVx1_ASAP7_75t_L g1848 ( 
.A(n_1528),
.Y(n_1848)
);

INVx1_ASAP7_75t_L g1849 ( 
.A(n_1541),
.Y(n_1849)
);

INVx1_ASAP7_75t_L g1850 ( 
.A(n_1560),
.Y(n_1850)
);

INVx1_ASAP7_75t_L g1851 ( 
.A(n_1515),
.Y(n_1851)
);

INVxp67_ASAP7_75t_SL g1852 ( 
.A(n_1689),
.Y(n_1852)
);

NOR2xp33_ASAP7_75t_L g1853 ( 
.A(n_1517),
.B(n_997),
.Y(n_1853)
);

AND2x2_ASAP7_75t_L g1854 ( 
.A(n_1615),
.B(n_1487),
.Y(n_1854)
);

BUFx3_ASAP7_75t_L g1855 ( 
.A(n_1719),
.Y(n_1855)
);

HB1xp67_ASAP7_75t_L g1856 ( 
.A(n_1612),
.Y(n_1856)
);

AND2x4_ASAP7_75t_L g1857 ( 
.A(n_1730),
.B(n_1489),
.Y(n_1857)
);

NOR2x1_ASAP7_75t_SL g1858 ( 
.A(n_1712),
.B(n_1501),
.Y(n_1858)
);

INVx1_ASAP7_75t_L g1859 ( 
.A(n_1524),
.Y(n_1859)
);

OAI21xp5_ASAP7_75t_L g1860 ( 
.A1(n_1537),
.A2(n_1424),
.B(n_1469),
.Y(n_1860)
);

AND2x2_ASAP7_75t_L g1861 ( 
.A(n_1564),
.B(n_1626),
.Y(n_1861)
);

NAND2xp5_ASAP7_75t_L g1862 ( 
.A(n_1647),
.B(n_1469),
.Y(n_1862)
);

NAND2xp5_ASAP7_75t_L g1863 ( 
.A(n_1714),
.B(n_1471),
.Y(n_1863)
);

BUFx3_ASAP7_75t_L g1864 ( 
.A(n_1632),
.Y(n_1864)
);

INVx2_ASAP7_75t_L g1865 ( 
.A(n_1673),
.Y(n_1865)
);

AND2x2_ASAP7_75t_L g1866 ( 
.A(n_1564),
.B(n_1487),
.Y(n_1866)
);

BUFx5_ASAP7_75t_L g1867 ( 
.A(n_1583),
.Y(n_1867)
);

HB1xp67_ASAP7_75t_L g1868 ( 
.A(n_1618),
.Y(n_1868)
);

AND2x4_ASAP7_75t_L g1869 ( 
.A(n_1527),
.B(n_1487),
.Y(n_1869)
);

INVx2_ASAP7_75t_L g1870 ( 
.A(n_1673),
.Y(n_1870)
);

INVx1_ASAP7_75t_L g1871 ( 
.A(n_1562),
.Y(n_1871)
);

INVx1_ASAP7_75t_L g1872 ( 
.A(n_1568),
.Y(n_1872)
);

AND2x2_ASAP7_75t_L g1873 ( 
.A(n_1665),
.B(n_1618),
.Y(n_1873)
);

INVx1_ASAP7_75t_L g1874 ( 
.A(n_1577),
.Y(n_1874)
);

BUFx6f_ASAP7_75t_L g1875 ( 
.A(n_1553),
.Y(n_1875)
);

INVx1_ASAP7_75t_L g1876 ( 
.A(n_1581),
.Y(n_1876)
);

INVx1_ASAP7_75t_L g1877 ( 
.A(n_1585),
.Y(n_1877)
);

AND2x2_ASAP7_75t_L g1878 ( 
.A(n_1701),
.B(n_1496),
.Y(n_1878)
);

NAND2xp5_ASAP7_75t_L g1879 ( 
.A(n_1714),
.B(n_1471),
.Y(n_1879)
);

BUFx3_ASAP7_75t_L g1880 ( 
.A(n_1728),
.Y(n_1880)
);

BUFx2_ASAP7_75t_L g1881 ( 
.A(n_1644),
.Y(n_1881)
);

OR2x2_ASAP7_75t_L g1882 ( 
.A(n_1571),
.B(n_1510),
.Y(n_1882)
);

NAND2xp5_ASAP7_75t_L g1883 ( 
.A(n_1604),
.B(n_1473),
.Y(n_1883)
);

AND2x2_ASAP7_75t_L g1884 ( 
.A(n_1701),
.B(n_1496),
.Y(n_1884)
);

INVx1_ASAP7_75t_L g1885 ( 
.A(n_1534),
.Y(n_1885)
);

HB1xp67_ASAP7_75t_L g1886 ( 
.A(n_1613),
.Y(n_1886)
);

NAND2xp5_ASAP7_75t_L g1887 ( 
.A(n_1607),
.B(n_1473),
.Y(n_1887)
);

INVx4_ASAP7_75t_L g1888 ( 
.A(n_1712),
.Y(n_1888)
);

INVx1_ASAP7_75t_L g1889 ( 
.A(n_1534),
.Y(n_1889)
);

HB1xp67_ASAP7_75t_L g1890 ( 
.A(n_1642),
.Y(n_1890)
);

INVx1_ASAP7_75t_L g1891 ( 
.A(n_1551),
.Y(n_1891)
);

INVx2_ASAP7_75t_L g1892 ( 
.A(n_1673),
.Y(n_1892)
);

AND2x2_ASAP7_75t_L g1893 ( 
.A(n_1700),
.B(n_1496),
.Y(n_1893)
);

NAND2xp5_ASAP7_75t_L g1894 ( 
.A(n_1634),
.B(n_1479),
.Y(n_1894)
);

AND2x2_ASAP7_75t_L g1895 ( 
.A(n_1700),
.B(n_1496),
.Y(n_1895)
);

BUFx12f_ASAP7_75t_L g1896 ( 
.A(n_1563),
.Y(n_1896)
);

INVx3_ASAP7_75t_L g1897 ( 
.A(n_1553),
.Y(n_1897)
);

NAND2xp5_ASAP7_75t_L g1898 ( 
.A(n_1596),
.B(n_1479),
.Y(n_1898)
);

AND2x4_ASAP7_75t_L g1899 ( 
.A(n_1527),
.B(n_1496),
.Y(n_1899)
);

NAND2xp5_ASAP7_75t_L g1900 ( 
.A(n_1551),
.B(n_1492),
.Y(n_1900)
);

INVx1_ASAP7_75t_L g1901 ( 
.A(n_1582),
.Y(n_1901)
);

OA21x2_ASAP7_75t_L g1902 ( 
.A1(n_1621),
.A2(n_1395),
.B(n_1394),
.Y(n_1902)
);

AND2x2_ASAP7_75t_L g1903 ( 
.A(n_1669),
.B(n_1674),
.Y(n_1903)
);

NAND2xp5_ASAP7_75t_L g1904 ( 
.A(n_1582),
.B(n_1492),
.Y(n_1904)
);

OR2x2_ASAP7_75t_L g1905 ( 
.A(n_1636),
.B(n_1510),
.Y(n_1905)
);

INVx1_ASAP7_75t_L g1906 ( 
.A(n_1636),
.Y(n_1906)
);

INVx2_ASAP7_75t_L g1907 ( 
.A(n_1716),
.Y(n_1907)
);

INVx5_ASAP7_75t_L g1908 ( 
.A(n_1520),
.Y(n_1908)
);

NAND2xp5_ASAP7_75t_L g1909 ( 
.A(n_1670),
.B(n_1498),
.Y(n_1909)
);

BUFx2_ASAP7_75t_L g1910 ( 
.A(n_1679),
.Y(n_1910)
);

INVx1_ASAP7_75t_L g1911 ( 
.A(n_1718),
.Y(n_1911)
);

AND2x2_ASAP7_75t_L g1912 ( 
.A(n_1675),
.B(n_1502),
.Y(n_1912)
);

INVx4_ASAP7_75t_L g1913 ( 
.A(n_1712),
.Y(n_1913)
);

INVx1_ASAP7_75t_L g1914 ( 
.A(n_1522),
.Y(n_1914)
);

INVx1_ASAP7_75t_L g1915 ( 
.A(n_1522),
.Y(n_1915)
);

INVx1_ASAP7_75t_L g1916 ( 
.A(n_1672),
.Y(n_1916)
);

INVx2_ASAP7_75t_SL g1917 ( 
.A(n_1576),
.Y(n_1917)
);

INVxp67_ASAP7_75t_L g1918 ( 
.A(n_1728),
.Y(n_1918)
);

AND2x2_ASAP7_75t_L g1919 ( 
.A(n_1576),
.B(n_1502),
.Y(n_1919)
);

INVx2_ASAP7_75t_L g1920 ( 
.A(n_1716),
.Y(n_1920)
);

INVx1_ASAP7_75t_L g1921 ( 
.A(n_1734),
.Y(n_1921)
);

INVx1_ASAP7_75t_L g1922 ( 
.A(n_1677),
.Y(n_1922)
);

AND2x2_ASAP7_75t_L g1923 ( 
.A(n_1659),
.B(n_1502),
.Y(n_1923)
);

HB1xp67_ASAP7_75t_L g1924 ( 
.A(n_1676),
.Y(n_1924)
);

INVx1_ASAP7_75t_L g1925 ( 
.A(n_1694),
.Y(n_1925)
);

HB1xp67_ASAP7_75t_L g1926 ( 
.A(n_1715),
.Y(n_1926)
);

INVx1_ASAP7_75t_L g1927 ( 
.A(n_1716),
.Y(n_1927)
);

AND2x2_ASAP7_75t_L g1928 ( 
.A(n_1659),
.B(n_1502),
.Y(n_1928)
);

AND2x4_ASAP7_75t_L g1929 ( 
.A(n_1527),
.B(n_1502),
.Y(n_1929)
);

NOR2xp33_ASAP7_75t_L g1930 ( 
.A(n_1537),
.B(n_997),
.Y(n_1930)
);

AND2x4_ASAP7_75t_L g1931 ( 
.A(n_1532),
.B(n_1475),
.Y(n_1931)
);

AND2x2_ASAP7_75t_L g1932 ( 
.A(n_1593),
.B(n_1417),
.Y(n_1932)
);

INVx2_ASAP7_75t_L g1933 ( 
.A(n_1716),
.Y(n_1933)
);

AOI22xp33_ASAP7_75t_L g1934 ( 
.A1(n_1552),
.A2(n_1411),
.B1(n_1370),
.B2(n_1375),
.Y(n_1934)
);

INVx1_ASAP7_75t_L g1935 ( 
.A(n_1529),
.Y(n_1935)
);

AND2x2_ASAP7_75t_L g1936 ( 
.A(n_1593),
.B(n_1417),
.Y(n_1936)
);

NAND2xp5_ASAP7_75t_L g1937 ( 
.A(n_1548),
.B(n_1498),
.Y(n_1937)
);

INVx1_ASAP7_75t_L g1938 ( 
.A(n_1529),
.Y(n_1938)
);

OAI222xp33_ASAP7_75t_L g1939 ( 
.A1(n_1578),
.A2(n_1389),
.B1(n_1388),
.B2(n_1378),
.C1(n_1392),
.C2(n_1420),
.Y(n_1939)
);

AND2x2_ASAP7_75t_L g1940 ( 
.A(n_1706),
.B(n_1724),
.Y(n_1940)
);

INVx1_ASAP7_75t_L g1941 ( 
.A(n_1529),
.Y(n_1941)
);

AND2x2_ASAP7_75t_L g1942 ( 
.A(n_1706),
.B(n_1447),
.Y(n_1942)
);

AND2x2_ASAP7_75t_L g1943 ( 
.A(n_1724),
.B(n_1572),
.Y(n_1943)
);

INVx1_ASAP7_75t_L g1944 ( 
.A(n_1529),
.Y(n_1944)
);

INVx1_ASAP7_75t_L g1945 ( 
.A(n_1538),
.Y(n_1945)
);

HB1xp67_ASAP7_75t_L g1946 ( 
.A(n_1546),
.Y(n_1946)
);

INVx2_ASAP7_75t_L g1947 ( 
.A(n_1554),
.Y(n_1947)
);

HB1xp67_ASAP7_75t_L g1948 ( 
.A(n_1566),
.Y(n_1948)
);

AND2x2_ASAP7_75t_L g1949 ( 
.A(n_1724),
.B(n_1447),
.Y(n_1949)
);

INVx2_ASAP7_75t_L g1950 ( 
.A(n_1841),
.Y(n_1950)
);

OAI22xp5_ASAP7_75t_L g1951 ( 
.A1(n_1752),
.A2(n_1580),
.B1(n_1654),
.B2(n_1627),
.Y(n_1951)
);

BUFx6f_ASAP7_75t_L g1952 ( 
.A(n_1747),
.Y(n_1952)
);

OAI21xp5_ASAP7_75t_L g1953 ( 
.A1(n_1860),
.A2(n_1540),
.B(n_1587),
.Y(n_1953)
);

OA21x2_ASAP7_75t_L g1954 ( 
.A1(n_1739),
.A2(n_1608),
.B(n_1592),
.Y(n_1954)
);

INVx1_ASAP7_75t_L g1955 ( 
.A(n_1793),
.Y(n_1955)
);

AOI21xp5_ASAP7_75t_L g1956 ( 
.A1(n_1763),
.A2(n_1858),
.B(n_1788),
.Y(n_1956)
);

AOI22xp33_ASAP7_75t_L g1957 ( 
.A1(n_1835),
.A2(n_1578),
.B1(n_1628),
.B2(n_1583),
.Y(n_1957)
);

BUFx3_ASAP7_75t_L g1958 ( 
.A(n_1747),
.Y(n_1958)
);

INVx8_ASAP7_75t_L g1959 ( 
.A(n_1747),
.Y(n_1959)
);

A2O1A1Ixp33_ASAP7_75t_L g1960 ( 
.A1(n_1832),
.A2(n_1600),
.B(n_1584),
.C(n_1623),
.Y(n_1960)
);

AOI21xp5_ASAP7_75t_L g1961 ( 
.A1(n_1788),
.A2(n_1658),
.B(n_1691),
.Y(n_1961)
);

A2O1A1Ixp33_ASAP7_75t_L g1962 ( 
.A1(n_1852),
.A2(n_1600),
.B(n_1628),
.C(n_1556),
.Y(n_1962)
);

OA21x2_ASAP7_75t_L g1963 ( 
.A1(n_1739),
.A2(n_1629),
.B(n_1625),
.Y(n_1963)
);

INVx2_ASAP7_75t_L g1964 ( 
.A(n_1841),
.Y(n_1964)
);

NAND4xp25_ASAP7_75t_L g1965 ( 
.A(n_1930),
.B(n_1657),
.C(n_1638),
.D(n_1663),
.Y(n_1965)
);

OAI21x1_ASAP7_75t_L g1966 ( 
.A1(n_1742),
.A2(n_1637),
.B(n_1631),
.Y(n_1966)
);

HB1xp67_ASAP7_75t_L g1967 ( 
.A(n_1911),
.Y(n_1967)
);

OA21x2_ASAP7_75t_L g1968 ( 
.A1(n_1742),
.A2(n_1664),
.B(n_1646),
.Y(n_1968)
);

AOI21xp5_ASAP7_75t_L g1969 ( 
.A1(n_1858),
.A2(n_1532),
.B(n_1720),
.Y(n_1969)
);

BUFx3_ASAP7_75t_L g1970 ( 
.A(n_1747),
.Y(n_1970)
);

AOI221xp5_ASAP7_75t_L g1971 ( 
.A1(n_1762),
.A2(n_1506),
.B1(n_1465),
.B2(n_1460),
.C(n_1443),
.Y(n_1971)
);

NOR2xp33_ASAP7_75t_L g1972 ( 
.A(n_1808),
.B(n_1732),
.Y(n_1972)
);

NAND2xp5_ASAP7_75t_SL g1973 ( 
.A(n_1838),
.B(n_1679),
.Y(n_1973)
);

OAI211xp5_ASAP7_75t_L g1974 ( 
.A1(n_1823),
.A2(n_1531),
.B(n_1535),
.C(n_1530),
.Y(n_1974)
);

INVx2_ASAP7_75t_L g1975 ( 
.A(n_1865),
.Y(n_1975)
);

INVxp67_ASAP7_75t_L g1976 ( 
.A(n_1824),
.Y(n_1976)
);

AND2x2_ASAP7_75t_L g1977 ( 
.A(n_1794),
.B(n_1558),
.Y(n_1977)
);

NOR2x1p5_ASAP7_75t_L g1978 ( 
.A(n_1747),
.B(n_1036),
.Y(n_1978)
);

AND2x4_ASAP7_75t_L g1979 ( 
.A(n_1842),
.B(n_1601),
.Y(n_1979)
);

AOI22xp5_ASAP7_75t_L g1980 ( 
.A1(n_1934),
.A2(n_1650),
.B1(n_1652),
.B2(n_1643),
.Y(n_1980)
);

INVx1_ASAP7_75t_L g1981 ( 
.A(n_1793),
.Y(n_1981)
);

BUFx3_ASAP7_75t_L g1982 ( 
.A(n_1768),
.Y(n_1982)
);

INVx1_ASAP7_75t_L g1983 ( 
.A(n_1801),
.Y(n_1983)
);

AO21x2_ASAP7_75t_L g1984 ( 
.A1(n_1914),
.A2(n_1357),
.B(n_1354),
.Y(n_1984)
);

INVx1_ASAP7_75t_L g1985 ( 
.A(n_1801),
.Y(n_1985)
);

NAND3xp33_ASAP7_75t_L g1986 ( 
.A(n_1782),
.B(n_1915),
.C(n_1914),
.Y(n_1986)
);

AND2x2_ASAP7_75t_L g1987 ( 
.A(n_1794),
.B(n_1798),
.Y(n_1987)
);

A2O1A1Ixp33_ASAP7_75t_L g1988 ( 
.A1(n_1807),
.A2(n_1713),
.B(n_1603),
.C(n_1731),
.Y(n_1988)
);

INVx1_ASAP7_75t_L g1989 ( 
.A(n_1802),
.Y(n_1989)
);

INVx1_ASAP7_75t_L g1990 ( 
.A(n_1802),
.Y(n_1990)
);

OA21x2_ASAP7_75t_L g1991 ( 
.A1(n_1744),
.A2(n_1364),
.B(n_1357),
.Y(n_1991)
);

OR2x2_ASAP7_75t_L g1992 ( 
.A(n_1886),
.B(n_1508),
.Y(n_1992)
);

OAI21x1_ASAP7_75t_L g1993 ( 
.A1(n_1744),
.A2(n_1731),
.B(n_1476),
.Y(n_1993)
);

INVx1_ASAP7_75t_L g1994 ( 
.A(n_1810),
.Y(n_1994)
);

INVx2_ASAP7_75t_L g1995 ( 
.A(n_1865),
.Y(n_1995)
);

INVx1_ASAP7_75t_L g1996 ( 
.A(n_1810),
.Y(n_1996)
);

INVx2_ASAP7_75t_L g1997 ( 
.A(n_1870),
.Y(n_1997)
);

AOI21xp5_ASAP7_75t_SL g1998 ( 
.A1(n_1807),
.A2(n_1521),
.B(n_1520),
.Y(n_1998)
);

INVx1_ASAP7_75t_L g1999 ( 
.A(n_1817),
.Y(n_1999)
);

INVx1_ASAP7_75t_L g2000 ( 
.A(n_1817),
.Y(n_2000)
);

OA21x2_ASAP7_75t_L g2001 ( 
.A1(n_1756),
.A2(n_1364),
.B(n_1381),
.Y(n_2001)
);

INVx1_ASAP7_75t_L g2002 ( 
.A(n_1828),
.Y(n_2002)
);

AOI22xp33_ASAP7_75t_L g2003 ( 
.A1(n_1867),
.A2(n_1748),
.B1(n_1753),
.B2(n_1778),
.Y(n_2003)
);

INVx1_ASAP7_75t_L g2004 ( 
.A(n_1828),
.Y(n_2004)
);

AO21x2_ASAP7_75t_L g2005 ( 
.A1(n_1915),
.A2(n_1666),
.B(n_1575),
.Y(n_2005)
);

AOI221xp5_ASAP7_75t_L g2006 ( 
.A1(n_1939),
.A2(n_1786),
.B1(n_1911),
.B2(n_1938),
.C(n_1935),
.Y(n_2006)
);

INVx1_ASAP7_75t_L g2007 ( 
.A(n_1837),
.Y(n_2007)
);

AND2x2_ASAP7_75t_L g2008 ( 
.A(n_1798),
.B(n_1565),
.Y(n_2008)
);

BUFx2_ASAP7_75t_L g2009 ( 
.A(n_1745),
.Y(n_2009)
);

AOI21xp5_ASAP7_75t_L g2010 ( 
.A1(n_1787),
.A2(n_1532),
.B(n_1720),
.Y(n_2010)
);

INVx4_ASAP7_75t_L g2011 ( 
.A(n_1761),
.Y(n_2011)
);

NAND2xp5_ASAP7_75t_L g2012 ( 
.A(n_1741),
.B(n_1508),
.Y(n_2012)
);

INVx1_ASAP7_75t_L g2013 ( 
.A(n_1837),
.Y(n_2013)
);

O2A1O1Ixp33_ASAP7_75t_L g2014 ( 
.A1(n_1863),
.A2(n_1465),
.B(n_1460),
.C(n_1443),
.Y(n_2014)
);

INVx4_ASAP7_75t_L g2015 ( 
.A(n_1761),
.Y(n_2015)
);

INVx1_ASAP7_75t_L g2016 ( 
.A(n_1840),
.Y(n_2016)
);

NAND4xp25_ASAP7_75t_L g2017 ( 
.A(n_1879),
.B(n_1447),
.C(n_1504),
.D(n_1697),
.Y(n_2017)
);

INVxp67_ASAP7_75t_L g2018 ( 
.A(n_1824),
.Y(n_2018)
);

AOI222xp33_ASAP7_75t_L g2019 ( 
.A1(n_1838),
.A2(n_1910),
.B1(n_1881),
.B2(n_1375),
.C1(n_1756),
.C2(n_1420),
.Y(n_2019)
);

INVx2_ASAP7_75t_L g2020 ( 
.A(n_1870),
.Y(n_2020)
);

OA21x2_ASAP7_75t_L g2021 ( 
.A1(n_1935),
.A2(n_1395),
.B(n_1394),
.Y(n_2021)
);

INVxp67_ASAP7_75t_L g2022 ( 
.A(n_1745),
.Y(n_2022)
);

INVx1_ASAP7_75t_L g2023 ( 
.A(n_1840),
.Y(n_2023)
);

INVx1_ASAP7_75t_L g2024 ( 
.A(n_1844),
.Y(n_2024)
);

A2O1A1Ixp33_ASAP7_75t_L g2025 ( 
.A1(n_1881),
.A2(n_1713),
.B(n_1603),
.C(n_1668),
.Y(n_2025)
);

HB1xp67_ASAP7_75t_L g2026 ( 
.A(n_1770),
.Y(n_2026)
);

AO21x2_ASAP7_75t_L g2027 ( 
.A1(n_1938),
.A2(n_1944),
.B(n_1941),
.Y(n_2027)
);

AOI21xp5_ASAP7_75t_L g2028 ( 
.A1(n_1787),
.A2(n_1521),
.B(n_1668),
.Y(n_2028)
);

INVx1_ASAP7_75t_L g2029 ( 
.A(n_1844),
.Y(n_2029)
);

AOI22xp33_ASAP7_75t_L g2030 ( 
.A1(n_1867),
.A2(n_1411),
.B1(n_1506),
.B2(n_1575),
.Y(n_2030)
);

NAND4xp25_ASAP7_75t_L g2031 ( 
.A(n_1885),
.B(n_1504),
.C(n_1703),
.D(n_1688),
.Y(n_2031)
);

INVx1_ASAP7_75t_L g2032 ( 
.A(n_1848),
.Y(n_2032)
);

AO21x2_ASAP7_75t_L g2033 ( 
.A1(n_1941),
.A2(n_1419),
.B(n_1413),
.Y(n_2033)
);

OAI21x1_ASAP7_75t_L g2034 ( 
.A1(n_1944),
.A2(n_1374),
.B(n_1372),
.Y(n_2034)
);

INVx2_ASAP7_75t_L g2035 ( 
.A(n_1892),
.Y(n_2035)
);

INVx1_ASAP7_75t_L g2036 ( 
.A(n_1848),
.Y(n_2036)
);

NAND2xp5_ASAP7_75t_L g2037 ( 
.A(n_1924),
.B(n_1509),
.Y(n_2037)
);

OAI211xp5_ASAP7_75t_L g2038 ( 
.A1(n_1910),
.A2(n_1531),
.B(n_1535),
.C(n_1561),
.Y(n_2038)
);

INVx1_ASAP7_75t_L g2039 ( 
.A(n_1849),
.Y(n_2039)
);

INVx1_ASAP7_75t_L g2040 ( 
.A(n_1849),
.Y(n_2040)
);

OR2x2_ASAP7_75t_L g2041 ( 
.A(n_1890),
.B(n_1509),
.Y(n_2041)
);

AOI22xp33_ASAP7_75t_L g2042 ( 
.A1(n_1867),
.A2(n_1411),
.B1(n_1374),
.B2(n_1377),
.Y(n_2042)
);

AOI22xp33_ASAP7_75t_SL g2043 ( 
.A1(n_1867),
.A2(n_1668),
.B1(n_1617),
.B2(n_1611),
.Y(n_2043)
);

INVx2_ASAP7_75t_L g2044 ( 
.A(n_1892),
.Y(n_2044)
);

A2O1A1Ixp33_ASAP7_75t_L g2045 ( 
.A1(n_1855),
.A2(n_1688),
.B(n_1481),
.C(n_1650),
.Y(n_2045)
);

INVx2_ASAP7_75t_L g2046 ( 
.A(n_1907),
.Y(n_2046)
);

AOI22xp33_ASAP7_75t_L g2047 ( 
.A1(n_1867),
.A2(n_1377),
.B1(n_1374),
.B2(n_1372),
.Y(n_2047)
);

INVx1_ASAP7_75t_L g2048 ( 
.A(n_1850),
.Y(n_2048)
);

INVx1_ASAP7_75t_L g2049 ( 
.A(n_1850),
.Y(n_2049)
);

AOI22xp33_ASAP7_75t_L g2050 ( 
.A1(n_1867),
.A2(n_1377),
.B1(n_1372),
.B2(n_1481),
.Y(n_2050)
);

AOI21xp5_ASAP7_75t_L g2051 ( 
.A1(n_1787),
.A2(n_1521),
.B(n_1586),
.Y(n_2051)
);

AND2x2_ASAP7_75t_L g2052 ( 
.A(n_1767),
.B(n_1683),
.Y(n_2052)
);

BUFx2_ASAP7_75t_L g2053 ( 
.A(n_1896),
.Y(n_2053)
);

NAND4xp25_ASAP7_75t_L g2054 ( 
.A(n_1885),
.B(n_1504),
.C(n_1512),
.D(n_1131),
.Y(n_2054)
);

NOR2xp33_ASAP7_75t_L g2055 ( 
.A(n_1768),
.B(n_1572),
.Y(n_2055)
);

INVx1_ASAP7_75t_L g2056 ( 
.A(n_1851),
.Y(n_2056)
);

NAND4xp25_ASAP7_75t_L g2057 ( 
.A(n_1889),
.B(n_1504),
.C(n_1512),
.D(n_1124),
.Y(n_2057)
);

BUFx3_ASAP7_75t_L g2058 ( 
.A(n_1761),
.Y(n_2058)
);

OAI221xp5_ASAP7_75t_L g2059 ( 
.A1(n_1784),
.A2(n_1652),
.B1(n_1643),
.B2(n_1419),
.C(n_1413),
.Y(n_2059)
);

A2O1A1Ixp33_ASAP7_75t_L g2060 ( 
.A1(n_1855),
.A2(n_1908),
.B(n_1826),
.C(n_1834),
.Y(n_2060)
);

INVx2_ASAP7_75t_L g2061 ( 
.A(n_1907),
.Y(n_2061)
);

INVx3_ASAP7_75t_L g2062 ( 
.A(n_1842),
.Y(n_2062)
);

NAND2xp5_ASAP7_75t_L g2063 ( 
.A(n_1926),
.B(n_1572),
.Y(n_2063)
);

AOI22xp5_ASAP7_75t_L g2064 ( 
.A1(n_1867),
.A2(n_1609),
.B1(n_1586),
.B2(n_1485),
.Y(n_2064)
);

OR2x2_ASAP7_75t_L g2065 ( 
.A(n_1827),
.B(n_1617),
.Y(n_2065)
);

BUFx2_ASAP7_75t_L g2066 ( 
.A(n_1896),
.Y(n_2066)
);

AND2x2_ASAP7_75t_L g2067 ( 
.A(n_1767),
.B(n_1617),
.Y(n_2067)
);

NAND2xp5_ASAP7_75t_L g2068 ( 
.A(n_1765),
.B(n_1572),
.Y(n_2068)
);

AOI22xp33_ASAP7_75t_SL g2069 ( 
.A1(n_1867),
.A2(n_1908),
.B1(n_1753),
.B2(n_1784),
.Y(n_2069)
);

INVx2_ASAP7_75t_SL g2070 ( 
.A(n_1792),
.Y(n_2070)
);

NAND2xp5_ASAP7_75t_SL g2071 ( 
.A(n_1787),
.B(n_1611),
.Y(n_2071)
);

NAND2xp5_ASAP7_75t_L g2072 ( 
.A(n_1797),
.B(n_1705),
.Y(n_2072)
);

INVx2_ASAP7_75t_L g2073 ( 
.A(n_1920),
.Y(n_2073)
);

INVxp67_ASAP7_75t_SL g2074 ( 
.A(n_1937),
.Y(n_2074)
);

INVx2_ASAP7_75t_L g2075 ( 
.A(n_1920),
.Y(n_2075)
);

OAI21x1_ASAP7_75t_L g2076 ( 
.A1(n_1933),
.A2(n_1402),
.B(n_1450),
.Y(n_2076)
);

INVx1_ASAP7_75t_L g2077 ( 
.A(n_1851),
.Y(n_2077)
);

INVx1_ASAP7_75t_L g2078 ( 
.A(n_1859),
.Y(n_2078)
);

AND2x4_ASAP7_75t_L g2079 ( 
.A(n_1842),
.B(n_1586),
.Y(n_2079)
);

INVx1_ASAP7_75t_SL g2080 ( 
.A(n_1792),
.Y(n_2080)
);

INVx2_ASAP7_75t_L g2081 ( 
.A(n_1933),
.Y(n_2081)
);

OAI21x1_ASAP7_75t_L g2082 ( 
.A1(n_1836),
.A2(n_1405),
.B(n_1402),
.Y(n_2082)
);

INVx1_ASAP7_75t_L g2083 ( 
.A(n_1859),
.Y(n_2083)
);

INVx2_ASAP7_75t_SL g2084 ( 
.A(n_1903),
.Y(n_2084)
);

AND2x4_ASAP7_75t_SL g2085 ( 
.A(n_1842),
.B(n_1609),
.Y(n_2085)
);

INVx2_ASAP7_75t_L g2086 ( 
.A(n_1902),
.Y(n_2086)
);

INVx1_ASAP7_75t_L g2087 ( 
.A(n_1871),
.Y(n_2087)
);

INVx2_ASAP7_75t_L g2088 ( 
.A(n_1902),
.Y(n_2088)
);

NAND2xp5_ASAP7_75t_L g2089 ( 
.A(n_1862),
.B(n_1705),
.Y(n_2089)
);

BUFx2_ASAP7_75t_L g2090 ( 
.A(n_1857),
.Y(n_2090)
);

AOI211xp5_ASAP7_75t_L g2091 ( 
.A1(n_1931),
.A2(n_1695),
.B(n_1685),
.C(n_1561),
.Y(n_2091)
);

NAND2xp5_ASAP7_75t_L g2092 ( 
.A(n_1887),
.B(n_1705),
.Y(n_2092)
);

AO21x2_ASAP7_75t_L g2093 ( 
.A1(n_1927),
.A2(n_1401),
.B(n_1406),
.Y(n_2093)
);

INVx1_ASAP7_75t_L g2094 ( 
.A(n_1871),
.Y(n_2094)
);

AOI22xp33_ASAP7_75t_SL g2095 ( 
.A1(n_1908),
.A2(n_1695),
.B1(n_1685),
.B2(n_1609),
.Y(n_2095)
);

INVx2_ASAP7_75t_L g2096 ( 
.A(n_1902),
.Y(n_2096)
);

INVxp67_ASAP7_75t_L g2097 ( 
.A(n_1806),
.Y(n_2097)
);

A2O1A1Ixp33_ASAP7_75t_L g2098 ( 
.A1(n_1908),
.A2(n_1427),
.B(n_1396),
.C(n_1507),
.Y(n_2098)
);

INVx1_ASAP7_75t_L g2099 ( 
.A(n_1872),
.Y(n_2099)
);

AO21x2_ASAP7_75t_L g2100 ( 
.A1(n_1927),
.A2(n_1401),
.B(n_1406),
.Y(n_2100)
);

INVx1_ASAP7_75t_L g2101 ( 
.A(n_1872),
.Y(n_2101)
);

A2O1A1Ixp33_ASAP7_75t_L g2102 ( 
.A1(n_1908),
.A2(n_1427),
.B(n_1396),
.C(n_1429),
.Y(n_2102)
);

AO31x2_ASAP7_75t_L g2103 ( 
.A1(n_1888),
.A2(n_1403),
.A3(n_1406),
.B(n_1401),
.Y(n_2103)
);

HB1xp67_ASAP7_75t_L g2104 ( 
.A(n_1816),
.Y(n_2104)
);

INVx1_ASAP7_75t_L g2105 ( 
.A(n_1874),
.Y(n_2105)
);

INVx1_ASAP7_75t_L g2106 ( 
.A(n_1874),
.Y(n_2106)
);

A2O1A1Ixp33_ASAP7_75t_L g2107 ( 
.A1(n_1908),
.A2(n_1396),
.B(n_1435),
.C(n_1431),
.Y(n_2107)
);

OR2x2_ASAP7_75t_L g2108 ( 
.A(n_1795),
.B(n_1705),
.Y(n_2108)
);

INVx3_ASAP7_75t_L g2109 ( 
.A(n_1857),
.Y(n_2109)
);

INVx2_ASAP7_75t_L g2110 ( 
.A(n_1902),
.Y(n_2110)
);

OA21x2_ASAP7_75t_L g2111 ( 
.A1(n_1758),
.A2(n_1403),
.B(n_1408),
.Y(n_2111)
);

INVx1_ASAP7_75t_L g2112 ( 
.A(n_1876),
.Y(n_2112)
);

AO21x2_ASAP7_75t_L g2113 ( 
.A1(n_1735),
.A2(n_1408),
.B(n_1403),
.Y(n_2113)
);

AOI211xp5_ASAP7_75t_L g2114 ( 
.A1(n_1931),
.A2(n_1598),
.B(n_1483),
.C(n_1373),
.Y(n_2114)
);

NAND2xp5_ASAP7_75t_L g2115 ( 
.A(n_1894),
.B(n_1429),
.Y(n_2115)
);

OAI22xp5_ASAP7_75t_L g2116 ( 
.A1(n_1918),
.A2(n_1483),
.B1(n_1373),
.B2(n_1446),
.Y(n_2116)
);

BUFx3_ASAP7_75t_L g2117 ( 
.A(n_1738),
.Y(n_2117)
);

BUFx3_ASAP7_75t_L g2118 ( 
.A(n_1736),
.Y(n_2118)
);

CKINVDCx6p67_ASAP7_75t_R g2119 ( 
.A(n_1864),
.Y(n_2119)
);

INVx1_ASAP7_75t_L g2120 ( 
.A(n_1876),
.Y(n_2120)
);

AOI22xp33_ASAP7_75t_L g2121 ( 
.A1(n_1753),
.A2(n_1431),
.B1(n_1435),
.B2(n_1429),
.Y(n_2121)
);

AOI21xp5_ASAP7_75t_L g2122 ( 
.A1(n_1826),
.A2(n_1501),
.B(n_1466),
.Y(n_2122)
);

HB1xp67_ASAP7_75t_L g2123 ( 
.A(n_1822),
.Y(n_2123)
);

AND2x2_ASAP7_75t_L g2124 ( 
.A(n_1750),
.B(n_1483),
.Y(n_2124)
);

INVxp67_ASAP7_75t_L g2125 ( 
.A(n_1806),
.Y(n_2125)
);

INVx1_ASAP7_75t_L g2126 ( 
.A(n_1877),
.Y(n_2126)
);

NAND2xp5_ASAP7_75t_L g2127 ( 
.A(n_1883),
.B(n_1431),
.Y(n_2127)
);

OAI22xp33_ASAP7_75t_L g2128 ( 
.A1(n_1888),
.A2(n_1446),
.B1(n_1301),
.B2(n_1243),
.Y(n_2128)
);

OR2x6_ASAP7_75t_L g2129 ( 
.A(n_1826),
.B(n_1501),
.Y(n_2129)
);

INVx1_ASAP7_75t_L g2130 ( 
.A(n_1877),
.Y(n_2130)
);

INVx1_ASAP7_75t_L g2131 ( 
.A(n_1898),
.Y(n_2131)
);

AOI21xp5_ASAP7_75t_L g2132 ( 
.A1(n_1826),
.A2(n_1834),
.B(n_1857),
.Y(n_2132)
);

AOI21xp5_ASAP7_75t_L g2133 ( 
.A1(n_1834),
.A2(n_1501),
.B(n_1466),
.Y(n_2133)
);

INVx2_ASAP7_75t_L g2134 ( 
.A(n_1905),
.Y(n_2134)
);

AND2x2_ASAP7_75t_L g2135 ( 
.A(n_1972),
.B(n_1931),
.Y(n_2135)
);

OAI22xp33_ASAP7_75t_L g2136 ( 
.A1(n_1980),
.A2(n_1784),
.B1(n_1888),
.B2(n_1803),
.Y(n_2136)
);

OAI33xp33_ASAP7_75t_L g2137 ( 
.A1(n_1951),
.A2(n_1906),
.A3(n_1901),
.B1(n_1891),
.B2(n_1889),
.B3(n_1900),
.Y(n_2137)
);

INVx1_ASAP7_75t_L g2138 ( 
.A(n_1955),
.Y(n_2138)
);

AND2x2_ASAP7_75t_L g2139 ( 
.A(n_1972),
.B(n_1931),
.Y(n_2139)
);

AND2x2_ASAP7_75t_L g2140 ( 
.A(n_2009),
.B(n_1750),
.Y(n_2140)
);

AND2x2_ASAP7_75t_L g2141 ( 
.A(n_2090),
.B(n_1861),
.Y(n_2141)
);

INVx1_ASAP7_75t_L g2142 ( 
.A(n_1981),
.Y(n_2142)
);

INVx2_ASAP7_75t_SL g2143 ( 
.A(n_1959),
.Y(n_2143)
);

AND2x2_ASAP7_75t_L g2144 ( 
.A(n_2062),
.B(n_1861),
.Y(n_2144)
);

HB1xp67_ASAP7_75t_L g2145 ( 
.A(n_2026),
.Y(n_2145)
);

OAI33xp33_ASAP7_75t_L g2146 ( 
.A1(n_2022),
.A2(n_1986),
.A3(n_2131),
.B1(n_1965),
.B2(n_2017),
.B3(n_2012),
.Y(n_2146)
);

AND2x2_ASAP7_75t_L g2147 ( 
.A(n_2062),
.B(n_1873),
.Y(n_2147)
);

AOI22xp33_ASAP7_75t_SL g2148 ( 
.A1(n_1953),
.A2(n_2059),
.B1(n_1753),
.B2(n_2074),
.Y(n_2148)
);

NAND2xp5_ASAP7_75t_L g2149 ( 
.A(n_2026),
.B(n_1825),
.Y(n_2149)
);

INVx1_ASAP7_75t_L g2150 ( 
.A(n_1983),
.Y(n_2150)
);

INVx1_ASAP7_75t_L g2151 ( 
.A(n_1985),
.Y(n_2151)
);

INVx3_ASAP7_75t_L g2152 ( 
.A(n_1952),
.Y(n_2152)
);

AO21x2_ASAP7_75t_L g2153 ( 
.A1(n_1960),
.A2(n_1901),
.B(n_1891),
.Y(n_2153)
);

AND2x2_ASAP7_75t_L g2154 ( 
.A(n_2109),
.B(n_1987),
.Y(n_2154)
);

INVx1_ASAP7_75t_L g2155 ( 
.A(n_1989),
.Y(n_2155)
);

INVx1_ASAP7_75t_L g2156 ( 
.A(n_1990),
.Y(n_2156)
);

AND2x2_ASAP7_75t_L g2157 ( 
.A(n_2109),
.B(n_1873),
.Y(n_2157)
);

INVxp33_ASAP7_75t_SL g2158 ( 
.A(n_2118),
.Y(n_2158)
);

AOI33xp33_ASAP7_75t_L g2159 ( 
.A1(n_2003),
.A2(n_1906),
.A3(n_1758),
.B1(n_1772),
.B2(n_1776),
.B3(n_1783),
.Y(n_2159)
);

AND2x2_ASAP7_75t_L g2160 ( 
.A(n_1979),
.B(n_1878),
.Y(n_2160)
);

OR2x2_ASAP7_75t_L g2161 ( 
.A(n_1992),
.B(n_1795),
.Y(n_2161)
);

OAI22xp5_ASAP7_75t_L g2162 ( 
.A1(n_1960),
.A2(n_1880),
.B1(n_1888),
.B2(n_1803),
.Y(n_2162)
);

INVx2_ASAP7_75t_L g2163 ( 
.A(n_2027),
.Y(n_2163)
);

AND2x4_ASAP7_75t_L g2164 ( 
.A(n_2060),
.B(n_2132),
.Y(n_2164)
);

NAND2xp5_ASAP7_75t_L g2165 ( 
.A(n_2104),
.B(n_1846),
.Y(n_2165)
);

CKINVDCx5p33_ASAP7_75t_R g2166 ( 
.A(n_1958),
.Y(n_2166)
);

AND2x2_ASAP7_75t_L g2167 ( 
.A(n_1979),
.B(n_1878),
.Y(n_2167)
);

INVx1_ASAP7_75t_L g2168 ( 
.A(n_1994),
.Y(n_2168)
);

INVx1_ASAP7_75t_L g2169 ( 
.A(n_1996),
.Y(n_2169)
);

OR2x2_ASAP7_75t_L g2170 ( 
.A(n_2041),
.B(n_1737),
.Y(n_2170)
);

INVx1_ASAP7_75t_SL g2171 ( 
.A(n_2118),
.Y(n_2171)
);

INVx2_ASAP7_75t_SL g2172 ( 
.A(n_1959),
.Y(n_2172)
);

AND2x4_ASAP7_75t_L g2173 ( 
.A(n_2060),
.B(n_1857),
.Y(n_2173)
);

CKINVDCx8_ASAP7_75t_R g2174 ( 
.A(n_1952),
.Y(n_2174)
);

INVx1_ASAP7_75t_L g2175 ( 
.A(n_1999),
.Y(n_2175)
);

AND2x2_ASAP7_75t_L g2176 ( 
.A(n_1979),
.B(n_1884),
.Y(n_2176)
);

INVx3_ASAP7_75t_L g2177 ( 
.A(n_1952),
.Y(n_2177)
);

AND2x4_ASAP7_75t_L g2178 ( 
.A(n_2079),
.B(n_1834),
.Y(n_2178)
);

INVx1_ASAP7_75t_L g2179 ( 
.A(n_2000),
.Y(n_2179)
);

INVx5_ASAP7_75t_L g2180 ( 
.A(n_2011),
.Y(n_2180)
);

AND2x2_ASAP7_75t_L g2181 ( 
.A(n_1977),
.B(n_1884),
.Y(n_2181)
);

AND2x2_ASAP7_75t_L g2182 ( 
.A(n_2008),
.B(n_1912),
.Y(n_2182)
);

AND2x2_ASAP7_75t_L g2183 ( 
.A(n_2067),
.B(n_1912),
.Y(n_2183)
);

AND2x2_ASAP7_75t_L g2184 ( 
.A(n_2119),
.B(n_1820),
.Y(n_2184)
);

INVx2_ASAP7_75t_L g2185 ( 
.A(n_2027),
.Y(n_2185)
);

BUFx3_ASAP7_75t_L g2186 ( 
.A(n_1959),
.Y(n_2186)
);

AND2x2_ASAP7_75t_L g2187 ( 
.A(n_2052),
.B(n_1820),
.Y(n_2187)
);

OR2x2_ASAP7_75t_L g2188 ( 
.A(n_2037),
.B(n_1737),
.Y(n_2188)
);

AND2x2_ASAP7_75t_L g2189 ( 
.A(n_1973),
.B(n_1829),
.Y(n_2189)
);

INVx1_ASAP7_75t_L g2190 ( 
.A(n_2002),
.Y(n_2190)
);

AND2x2_ASAP7_75t_L g2191 ( 
.A(n_1973),
.B(n_1829),
.Y(n_2191)
);

NAND2xp5_ASAP7_75t_L g2192 ( 
.A(n_2104),
.B(n_1856),
.Y(n_2192)
);

INVx4_ASAP7_75t_L g2193 ( 
.A(n_2011),
.Y(n_2193)
);

INVx5_ASAP7_75t_L g2194 ( 
.A(n_2011),
.Y(n_2194)
);

AND2x4_ASAP7_75t_L g2195 ( 
.A(n_2079),
.B(n_1869),
.Y(n_2195)
);

INVx1_ASAP7_75t_L g2196 ( 
.A(n_2004),
.Y(n_2196)
);

INVx2_ASAP7_75t_L g2197 ( 
.A(n_2113),
.Y(n_2197)
);

AND2x4_ASAP7_75t_L g2198 ( 
.A(n_2079),
.B(n_1869),
.Y(n_2198)
);

AO21x2_ASAP7_75t_L g2199 ( 
.A1(n_1962),
.A2(n_1740),
.B(n_1735),
.Y(n_2199)
);

NAND3xp33_ASAP7_75t_L g2200 ( 
.A(n_1962),
.B(n_1868),
.C(n_1776),
.Y(n_2200)
);

INVx1_ASAP7_75t_SL g2201 ( 
.A(n_1982),
.Y(n_2201)
);

INVx2_ASAP7_75t_L g2202 ( 
.A(n_2113),
.Y(n_2202)
);

INVx2_ASAP7_75t_L g2203 ( 
.A(n_2086),
.Y(n_2203)
);

AOI22xp33_ASAP7_75t_L g2204 ( 
.A1(n_1957),
.A2(n_1784),
.B1(n_1435),
.B2(n_1947),
.Y(n_2204)
);

AOI322xp5_ASAP7_75t_L g2205 ( 
.A1(n_2006),
.A2(n_1869),
.A3(n_1929),
.B1(n_1899),
.B2(n_1940),
.C1(n_1811),
.C2(n_1814),
.Y(n_2205)
);

INVx1_ASAP7_75t_L g2206 ( 
.A(n_2007),
.Y(n_2206)
);

AOI21xp5_ASAP7_75t_SL g2207 ( 
.A1(n_1988),
.A2(n_1913),
.B(n_1803),
.Y(n_2207)
);

AND2x4_ASAP7_75t_SL g2208 ( 
.A(n_1952),
.B(n_1903),
.Y(n_2208)
);

INVx1_ASAP7_75t_L g2209 ( 
.A(n_2013),
.Y(n_2209)
);

INVx1_ASAP7_75t_L g2210 ( 
.A(n_2016),
.Y(n_2210)
);

NAND2xp5_ASAP7_75t_L g2211 ( 
.A(n_2123),
.B(n_1909),
.Y(n_2211)
);

AND2x2_ASAP7_75t_L g2212 ( 
.A(n_2084),
.B(n_1813),
.Y(n_2212)
);

INVx1_ASAP7_75t_L g2213 ( 
.A(n_2023),
.Y(n_2213)
);

INVx1_ASAP7_75t_L g2214 ( 
.A(n_2024),
.Y(n_2214)
);

INVx1_ASAP7_75t_L g2215 ( 
.A(n_2029),
.Y(n_2215)
);

INVx2_ASAP7_75t_L g2216 ( 
.A(n_2086),
.Y(n_2216)
);

INVxp67_ASAP7_75t_SL g2217 ( 
.A(n_1982),
.Y(n_2217)
);

NAND2xp5_ASAP7_75t_L g2218 ( 
.A(n_2123),
.B(n_1772),
.Y(n_2218)
);

INVx1_ASAP7_75t_L g2219 ( 
.A(n_2032),
.Y(n_2219)
);

OAI221xp5_ASAP7_75t_L g2220 ( 
.A1(n_1957),
.A2(n_1784),
.B1(n_1947),
.B2(n_1743),
.C(n_1945),
.Y(n_2220)
);

INVx1_ASAP7_75t_L g2221 ( 
.A(n_2036),
.Y(n_2221)
);

OAI211xp5_ASAP7_75t_L g2222 ( 
.A1(n_1974),
.A2(n_1853),
.B(n_1897),
.C(n_1836),
.Y(n_2222)
);

AND2x2_ASAP7_75t_L g2223 ( 
.A(n_2124),
.B(n_1813),
.Y(n_2223)
);

INVx1_ASAP7_75t_L g2224 ( 
.A(n_2039),
.Y(n_2224)
);

INVx1_ASAP7_75t_L g2225 ( 
.A(n_2040),
.Y(n_2225)
);

NAND3x1_ASAP7_75t_L g2226 ( 
.A(n_1961),
.B(n_1943),
.C(n_1936),
.Y(n_2226)
);

OAI22xp5_ASAP7_75t_L g2227 ( 
.A1(n_1988),
.A2(n_1880),
.B1(n_1913),
.B2(n_1743),
.Y(n_2227)
);

INVx2_ASAP7_75t_L g2228 ( 
.A(n_2088),
.Y(n_2228)
);

AND2x2_ASAP7_75t_L g2229 ( 
.A(n_2097),
.B(n_1893),
.Y(n_2229)
);

OR2x2_ASAP7_75t_L g2230 ( 
.A(n_2134),
.B(n_1830),
.Y(n_2230)
);

BUFx2_ASAP7_75t_L g2231 ( 
.A(n_1958),
.Y(n_2231)
);

INVx1_ASAP7_75t_L g2232 ( 
.A(n_2048),
.Y(n_2232)
);

NAND2xp5_ASAP7_75t_L g2233 ( 
.A(n_1967),
.B(n_1783),
.Y(n_2233)
);

AOI31xp33_ASAP7_75t_L g2234 ( 
.A1(n_1976),
.A2(n_1819),
.A3(n_1936),
.B(n_1942),
.Y(n_2234)
);

INVx1_ASAP7_75t_L g2235 ( 
.A(n_2049),
.Y(n_2235)
);

NOR2xp33_ASAP7_75t_SL g2236 ( 
.A(n_2015),
.B(n_1913),
.Y(n_2236)
);

NAND2xp5_ASAP7_75t_L g2237 ( 
.A(n_1967),
.B(n_1785),
.Y(n_2237)
);

AND2x4_ASAP7_75t_L g2238 ( 
.A(n_1970),
.B(n_1869),
.Y(n_2238)
);

INVx4_ASAP7_75t_L g2239 ( 
.A(n_2015),
.Y(n_2239)
);

INVxp67_ASAP7_75t_SL g2240 ( 
.A(n_1970),
.Y(n_2240)
);

AOI22xp33_ASAP7_75t_SL g2241 ( 
.A1(n_1956),
.A2(n_1899),
.B1(n_1929),
.B2(n_1821),
.Y(n_2241)
);

AOI22xp33_ASAP7_75t_L g2242 ( 
.A1(n_2003),
.A2(n_1470),
.B1(n_1477),
.B2(n_1458),
.Y(n_2242)
);

NAND2xp5_ASAP7_75t_L g2243 ( 
.A(n_2056),
.B(n_2077),
.Y(n_2243)
);

INVx1_ASAP7_75t_L g2244 ( 
.A(n_2078),
.Y(n_2244)
);

INVx2_ASAP7_75t_L g2245 ( 
.A(n_2088),
.Y(n_2245)
);

NAND2xp5_ASAP7_75t_L g2246 ( 
.A(n_2083),
.B(n_1785),
.Y(n_2246)
);

INVx2_ASAP7_75t_L g2247 ( 
.A(n_2096),
.Y(n_2247)
);

AND2x2_ASAP7_75t_L g2248 ( 
.A(n_2125),
.B(n_1893),
.Y(n_2248)
);

AND2x2_ASAP7_75t_L g2249 ( 
.A(n_2071),
.B(n_2018),
.Y(n_2249)
);

INVxp67_ASAP7_75t_SL g2250 ( 
.A(n_2014),
.Y(n_2250)
);

INVx1_ASAP7_75t_L g2251 ( 
.A(n_2087),
.Y(n_2251)
);

INVx1_ASAP7_75t_L g2252 ( 
.A(n_2094),
.Y(n_2252)
);

AND2x4_ASAP7_75t_L g2253 ( 
.A(n_2071),
.B(n_1899),
.Y(n_2253)
);

AOI222xp33_ASAP7_75t_L g2254 ( 
.A1(n_2045),
.A2(n_1916),
.B1(n_1921),
.B2(n_1922),
.C1(n_1925),
.C2(n_1746),
.Y(n_2254)
);

OR2x2_ASAP7_75t_L g2255 ( 
.A(n_2134),
.B(n_1830),
.Y(n_2255)
);

INVx2_ASAP7_75t_L g2256 ( 
.A(n_2096),
.Y(n_2256)
);

AND2x2_ASAP7_75t_L g2257 ( 
.A(n_2055),
.B(n_1895),
.Y(n_2257)
);

OR2x2_ASAP7_75t_L g2258 ( 
.A(n_2099),
.B(n_1831),
.Y(n_2258)
);

INVx1_ASAP7_75t_L g2259 ( 
.A(n_2101),
.Y(n_2259)
);

INVxp67_ASAP7_75t_SL g2260 ( 
.A(n_2117),
.Y(n_2260)
);

OR2x2_ASAP7_75t_L g2261 ( 
.A(n_2105),
.B(n_2106),
.Y(n_2261)
);

OAI31xp33_ASAP7_75t_L g2262 ( 
.A1(n_2045),
.A2(n_1899),
.A3(n_1929),
.B(n_1940),
.Y(n_2262)
);

INVx1_ASAP7_75t_L g2263 ( 
.A(n_2112),
.Y(n_2263)
);

NAND3xp33_ASAP7_75t_L g2264 ( 
.A(n_2019),
.B(n_1799),
.C(n_1790),
.Y(n_2264)
);

AND2x2_ASAP7_75t_L g2265 ( 
.A(n_2055),
.B(n_1895),
.Y(n_2265)
);

AND2x2_ASAP7_75t_L g2266 ( 
.A(n_2114),
.B(n_1866),
.Y(n_2266)
);

INVx1_ASAP7_75t_L g2267 ( 
.A(n_2120),
.Y(n_2267)
);

NAND2xp5_ASAP7_75t_L g2268 ( 
.A(n_2126),
.B(n_2130),
.Y(n_2268)
);

AOI33xp33_ASAP7_75t_L g2269 ( 
.A1(n_2069),
.A2(n_1811),
.A3(n_1814),
.B1(n_1790),
.B2(n_1818),
.B3(n_1799),
.Y(n_2269)
);

INVx2_ASAP7_75t_L g2270 ( 
.A(n_2110),
.Y(n_2270)
);

AND2x2_ASAP7_75t_L g2271 ( 
.A(n_2053),
.B(n_1866),
.Y(n_2271)
);

OR2x2_ASAP7_75t_L g2272 ( 
.A(n_2031),
.B(n_2065),
.Y(n_2272)
);

AND2x2_ASAP7_75t_L g2273 ( 
.A(n_2066),
.B(n_1757),
.Y(n_2273)
);

AO21x2_ASAP7_75t_L g2274 ( 
.A1(n_2005),
.A2(n_1746),
.B(n_1740),
.Y(n_2274)
);

INVx2_ASAP7_75t_L g2275 ( 
.A(n_2110),
.Y(n_2275)
);

NOR2xp67_ASAP7_75t_L g2276 ( 
.A(n_2015),
.B(n_1949),
.Y(n_2276)
);

NOR2x1_ASAP7_75t_L g2277 ( 
.A(n_2117),
.B(n_1864),
.Y(n_2277)
);

INVx4_ASAP7_75t_L g2278 ( 
.A(n_2058),
.Y(n_2278)
);

INVx1_ASAP7_75t_L g2279 ( 
.A(n_1984),
.Y(n_2279)
);

INVx2_ASAP7_75t_L g2280 ( 
.A(n_2093),
.Y(n_2280)
);

NAND3xp33_ASAP7_75t_L g2281 ( 
.A(n_1971),
.B(n_1818),
.C(n_1904),
.Y(n_2281)
);

OR2x2_ASAP7_75t_L g2282 ( 
.A(n_2108),
.B(n_1831),
.Y(n_2282)
);

INVx2_ASAP7_75t_L g2283 ( 
.A(n_2093),
.Y(n_2283)
);

INVx1_ASAP7_75t_L g2284 ( 
.A(n_1984),
.Y(n_2284)
);

AND2x2_ASAP7_75t_L g2285 ( 
.A(n_2091),
.B(n_1757),
.Y(n_2285)
);

INVxp67_ASAP7_75t_SL g2286 ( 
.A(n_1993),
.Y(n_2286)
);

AO221x2_ASAP7_75t_L g2287 ( 
.A1(n_2116),
.A2(n_1821),
.B1(n_1819),
.B2(n_1917),
.C(n_1030),
.Y(n_2287)
);

HB1xp67_ASAP7_75t_L g2288 ( 
.A(n_2068),
.Y(n_2288)
);

INVx1_ASAP7_75t_L g2289 ( 
.A(n_2033),
.Y(n_2289)
);

AOI22xp5_ASAP7_75t_L g2290 ( 
.A1(n_2064),
.A2(n_1945),
.B1(n_1929),
.B2(n_1777),
.Y(n_2290)
);

HB1xp67_ASAP7_75t_L g2291 ( 
.A(n_2072),
.Y(n_2291)
);

AND2x2_ASAP7_75t_L g2292 ( 
.A(n_2164),
.B(n_2070),
.Y(n_2292)
);

INVx3_ASAP7_75t_L g2293 ( 
.A(n_2153),
.Y(n_2293)
);

AND2x4_ASAP7_75t_L g2294 ( 
.A(n_2173),
.B(n_2164),
.Y(n_2294)
);

INVx1_ASAP7_75t_L g2295 ( 
.A(n_2261),
.Y(n_2295)
);

NOR2xp33_ASAP7_75t_L g2296 ( 
.A(n_2158),
.B(n_2058),
.Y(n_2296)
);

INVx2_ASAP7_75t_SL g2297 ( 
.A(n_2208),
.Y(n_2297)
);

AOI22xp33_ASAP7_75t_L g2298 ( 
.A1(n_2199),
.A2(n_2042),
.B1(n_2030),
.B2(n_2050),
.Y(n_2298)
);

INVx1_ASAP7_75t_L g2299 ( 
.A(n_2138),
.Y(n_2299)
);

AND2x2_ASAP7_75t_L g2300 ( 
.A(n_2164),
.B(n_1978),
.Y(n_2300)
);

INVxp33_ASAP7_75t_L g2301 ( 
.A(n_2277),
.Y(n_2301)
);

INVx1_ASAP7_75t_L g2302 ( 
.A(n_2142),
.Y(n_2302)
);

BUFx3_ASAP7_75t_L g2303 ( 
.A(n_2158),
.Y(n_2303)
);

NAND2xp5_ASAP7_75t_L g2304 ( 
.A(n_2260),
.B(n_2080),
.Y(n_2304)
);

INVx1_ASAP7_75t_L g2305 ( 
.A(n_2150),
.Y(n_2305)
);

INVx2_ASAP7_75t_L g2306 ( 
.A(n_2199),
.Y(n_2306)
);

NOR2x1p5_ASAP7_75t_L g2307 ( 
.A(n_2217),
.B(n_2054),
.Y(n_2307)
);

NAND2xp5_ASAP7_75t_L g2308 ( 
.A(n_2171),
.B(n_2127),
.Y(n_2308)
);

INVx1_ASAP7_75t_L g2309 ( 
.A(n_2151),
.Y(n_2309)
);

INVx1_ASAP7_75t_L g2310 ( 
.A(n_2155),
.Y(n_2310)
);

INVx1_ASAP7_75t_L g2311 ( 
.A(n_2156),
.Y(n_2311)
);

AOI22xp33_ASAP7_75t_L g2312 ( 
.A1(n_2146),
.A2(n_2042),
.B1(n_2030),
.B2(n_2050),
.Y(n_2312)
);

AND2x2_ASAP7_75t_L g2313 ( 
.A(n_2182),
.B(n_1766),
.Y(n_2313)
);

INVxp67_ASAP7_75t_L g2314 ( 
.A(n_2249),
.Y(n_2314)
);

NAND2xp5_ASAP7_75t_L g2315 ( 
.A(n_2250),
.B(n_2115),
.Y(n_2315)
);

NOR3xp33_ASAP7_75t_SL g2316 ( 
.A(n_2166),
.B(n_2038),
.C(n_2025),
.Y(n_2316)
);

INVx2_ASAP7_75t_L g2317 ( 
.A(n_2274),
.Y(n_2317)
);

AND2x2_ASAP7_75t_L g2318 ( 
.A(n_2182),
.B(n_1766),
.Y(n_2318)
);

AOI22xp33_ASAP7_75t_L g2319 ( 
.A1(n_2153),
.A2(n_1969),
.B1(n_2129),
.B2(n_2005),
.Y(n_2319)
);

AND2x2_ASAP7_75t_L g2320 ( 
.A(n_2160),
.B(n_1917),
.Y(n_2320)
);

INVx8_ASAP7_75t_L g2321 ( 
.A(n_2180),
.Y(n_2321)
);

AND2x2_ASAP7_75t_L g2322 ( 
.A(n_2160),
.B(n_1919),
.Y(n_2322)
);

AND2x2_ASAP7_75t_L g2323 ( 
.A(n_2167),
.B(n_1919),
.Y(n_2323)
);

NOR2xp33_ASAP7_75t_L g2324 ( 
.A(n_2201),
.B(n_2057),
.Y(n_2324)
);

AND2x2_ASAP7_75t_L g2325 ( 
.A(n_2167),
.B(n_1923),
.Y(n_2325)
);

NAND2xp5_ASAP7_75t_L g2326 ( 
.A(n_2145),
.B(n_1749),
.Y(n_2326)
);

INVx1_ASAP7_75t_L g2327 ( 
.A(n_2168),
.Y(n_2327)
);

AND2x2_ASAP7_75t_L g2328 ( 
.A(n_2176),
.B(n_1923),
.Y(n_2328)
);

AND2x2_ASAP7_75t_L g2329 ( 
.A(n_2176),
.B(n_1928),
.Y(n_2329)
);

INVx1_ASAP7_75t_L g2330 ( 
.A(n_2169),
.Y(n_2330)
);

INVx1_ASAP7_75t_L g2331 ( 
.A(n_2175),
.Y(n_2331)
);

BUFx2_ASAP7_75t_L g2332 ( 
.A(n_2240),
.Y(n_2332)
);

NOR2xp33_ASAP7_75t_SL g2333 ( 
.A(n_2166),
.B(n_2025),
.Y(n_2333)
);

AND2x2_ASAP7_75t_L g2334 ( 
.A(n_2154),
.B(n_1928),
.Y(n_2334)
);

OR2x2_ASAP7_75t_L g2335 ( 
.A(n_2258),
.B(n_1905),
.Y(n_2335)
);

INVx2_ASAP7_75t_L g2336 ( 
.A(n_2274),
.Y(n_2336)
);

INVx1_ASAP7_75t_L g2337 ( 
.A(n_2179),
.Y(n_2337)
);

INVx1_ASAP7_75t_L g2338 ( 
.A(n_2190),
.Y(n_2338)
);

INVx1_ASAP7_75t_L g2339 ( 
.A(n_2196),
.Y(n_2339)
);

AND2x2_ASAP7_75t_L g2340 ( 
.A(n_2154),
.B(n_1800),
.Y(n_2340)
);

HB1xp67_ASAP7_75t_L g2341 ( 
.A(n_2231),
.Y(n_2341)
);

INVx1_ASAP7_75t_L g2342 ( 
.A(n_2206),
.Y(n_2342)
);

AND2x2_ASAP7_75t_L g2343 ( 
.A(n_2271),
.B(n_1800),
.Y(n_2343)
);

INVx3_ASAP7_75t_L g2344 ( 
.A(n_2173),
.Y(n_2344)
);

INVx1_ASAP7_75t_L g2345 ( 
.A(n_2209),
.Y(n_2345)
);

AND2x2_ASAP7_75t_L g2346 ( 
.A(n_2271),
.B(n_1833),
.Y(n_2346)
);

AND2x2_ASAP7_75t_L g2347 ( 
.A(n_2181),
.B(n_2208),
.Y(n_2347)
);

INVx2_ASAP7_75t_L g2348 ( 
.A(n_2197),
.Y(n_2348)
);

AND2x2_ASAP7_75t_L g2349 ( 
.A(n_2181),
.B(n_1833),
.Y(n_2349)
);

AND2x2_ASAP7_75t_L g2350 ( 
.A(n_2273),
.B(n_1839),
.Y(n_2350)
);

INVx1_ASAP7_75t_L g2351 ( 
.A(n_2210),
.Y(n_2351)
);

AND2x4_ASAP7_75t_L g2352 ( 
.A(n_2173),
.B(n_2129),
.Y(n_2352)
);

INVx1_ASAP7_75t_L g2353 ( 
.A(n_2213),
.Y(n_2353)
);

AND2x2_ASAP7_75t_L g2354 ( 
.A(n_2273),
.B(n_1839),
.Y(n_2354)
);

AND2x2_ASAP7_75t_L g2355 ( 
.A(n_2141),
.B(n_1773),
.Y(n_2355)
);

INVx1_ASAP7_75t_L g2356 ( 
.A(n_2214),
.Y(n_2356)
);

NOR2xp33_ASAP7_75t_L g2357 ( 
.A(n_2278),
.B(n_2193),
.Y(n_2357)
);

AND2x2_ASAP7_75t_L g2358 ( 
.A(n_2141),
.B(n_1773),
.Y(n_2358)
);

AND2x2_ASAP7_75t_L g2359 ( 
.A(n_2187),
.B(n_1775),
.Y(n_2359)
);

AND2x2_ASAP7_75t_L g2360 ( 
.A(n_2187),
.B(n_1775),
.Y(n_2360)
);

AND2x2_ASAP7_75t_L g2361 ( 
.A(n_2249),
.B(n_1755),
.Y(n_2361)
);

INVx1_ASAP7_75t_L g2362 ( 
.A(n_2215),
.Y(n_2362)
);

BUFx2_ASAP7_75t_L g2363 ( 
.A(n_2278),
.Y(n_2363)
);

OR2x2_ASAP7_75t_L g2364 ( 
.A(n_2211),
.B(n_1749),
.Y(n_2364)
);

NOR2xp67_ASAP7_75t_L g2365 ( 
.A(n_2180),
.B(n_2010),
.Y(n_2365)
);

INVx2_ASAP7_75t_L g2366 ( 
.A(n_2197),
.Y(n_2366)
);

INVx2_ASAP7_75t_L g2367 ( 
.A(n_2202),
.Y(n_2367)
);

INVx1_ASAP7_75t_L g2368 ( 
.A(n_2219),
.Y(n_2368)
);

INVx2_ASAP7_75t_L g2369 ( 
.A(n_2202),
.Y(n_2369)
);

OR2x2_ASAP7_75t_L g2370 ( 
.A(n_2243),
.B(n_1751),
.Y(n_2370)
);

AND2x2_ASAP7_75t_L g2371 ( 
.A(n_2147),
.B(n_1755),
.Y(n_2371)
);

AND2x2_ASAP7_75t_L g2372 ( 
.A(n_2147),
.B(n_1769),
.Y(n_2372)
);

INVx1_ASAP7_75t_L g2373 ( 
.A(n_2221),
.Y(n_2373)
);

NAND2xp5_ASAP7_75t_L g2374 ( 
.A(n_2212),
.B(n_2149),
.Y(n_2374)
);

INVx2_ASAP7_75t_L g2375 ( 
.A(n_2280),
.Y(n_2375)
);

AND2x2_ASAP7_75t_L g2376 ( 
.A(n_2157),
.B(n_1769),
.Y(n_2376)
);

AND2x2_ASAP7_75t_L g2377 ( 
.A(n_2157),
.B(n_1809),
.Y(n_2377)
);

AOI22xp33_ASAP7_75t_L g2378 ( 
.A1(n_2148),
.A2(n_2129),
.B1(n_2133),
.B2(n_2122),
.Y(n_2378)
);

INVxp67_ASAP7_75t_L g2379 ( 
.A(n_2236),
.Y(n_2379)
);

HB1xp67_ASAP7_75t_L g2380 ( 
.A(n_2224),
.Y(n_2380)
);

INVx1_ASAP7_75t_L g2381 ( 
.A(n_2225),
.Y(n_2381)
);

BUFx2_ASAP7_75t_SL g2382 ( 
.A(n_2180),
.Y(n_2382)
);

AND2x4_ASAP7_75t_L g2383 ( 
.A(n_2178),
.B(n_2102),
.Y(n_2383)
);

INVx2_ASAP7_75t_L g2384 ( 
.A(n_2280),
.Y(n_2384)
);

AND2x4_ASAP7_75t_L g2385 ( 
.A(n_2178),
.B(n_2276),
.Y(n_2385)
);

INVx1_ASAP7_75t_SL g2386 ( 
.A(n_2186),
.Y(n_2386)
);

BUFx2_ASAP7_75t_L g2387 ( 
.A(n_2278),
.Y(n_2387)
);

AND2x2_ASAP7_75t_L g2388 ( 
.A(n_2140),
.B(n_1809),
.Y(n_2388)
);

INVx1_ASAP7_75t_L g2389 ( 
.A(n_2232),
.Y(n_2389)
);

INVx1_ASAP7_75t_L g2390 ( 
.A(n_2235),
.Y(n_2390)
);

INVx2_ASAP7_75t_L g2391 ( 
.A(n_2283),
.Y(n_2391)
);

INVxp67_ASAP7_75t_L g2392 ( 
.A(n_2143),
.Y(n_2392)
);

AND2x2_ASAP7_75t_L g2393 ( 
.A(n_2140),
.B(n_1812),
.Y(n_2393)
);

INVx1_ASAP7_75t_L g2394 ( 
.A(n_2244),
.Y(n_2394)
);

AND2x2_ASAP7_75t_L g2395 ( 
.A(n_2184),
.B(n_1812),
.Y(n_2395)
);

INVx1_ASAP7_75t_L g2396 ( 
.A(n_2251),
.Y(n_2396)
);

INVx2_ASAP7_75t_L g2397 ( 
.A(n_2283),
.Y(n_2397)
);

AND2x2_ASAP7_75t_L g2398 ( 
.A(n_2184),
.B(n_1771),
.Y(n_2398)
);

OR2x2_ASAP7_75t_L g2399 ( 
.A(n_2268),
.B(n_1751),
.Y(n_2399)
);

AND2x2_ASAP7_75t_L g2400 ( 
.A(n_2144),
.B(n_2189),
.Y(n_2400)
);

OR2x2_ASAP7_75t_L g2401 ( 
.A(n_2246),
.B(n_1754),
.Y(n_2401)
);

INVx2_ASAP7_75t_SL g2402 ( 
.A(n_2180),
.Y(n_2402)
);

INVx1_ASAP7_75t_L g2403 ( 
.A(n_2252),
.Y(n_2403)
);

NAND2xp5_ASAP7_75t_SL g2404 ( 
.A(n_2162),
.B(n_2043),
.Y(n_2404)
);

NAND2xp5_ASAP7_75t_L g2405 ( 
.A(n_2212),
.B(n_1754),
.Y(n_2405)
);

INVx1_ASAP7_75t_L g2406 ( 
.A(n_2259),
.Y(n_2406)
);

AND2x2_ASAP7_75t_L g2407 ( 
.A(n_2144),
.B(n_2189),
.Y(n_2407)
);

NAND2xp5_ASAP7_75t_L g2408 ( 
.A(n_2165),
.B(n_1759),
.Y(n_2408)
);

AND2x2_ASAP7_75t_L g2409 ( 
.A(n_2191),
.B(n_1771),
.Y(n_2409)
);

NAND2xp5_ASAP7_75t_L g2410 ( 
.A(n_2192),
.B(n_1759),
.Y(n_2410)
);

HB1xp67_ASAP7_75t_L g2411 ( 
.A(n_2263),
.Y(n_2411)
);

OR2x2_ASAP7_75t_L g2412 ( 
.A(n_2218),
.B(n_1760),
.Y(n_2412)
);

INVx1_ASAP7_75t_L g2413 ( 
.A(n_2267),
.Y(n_2413)
);

NAND2x1p5_ASAP7_75t_L g2414 ( 
.A(n_2180),
.B(n_1993),
.Y(n_2414)
);

HB1xp67_ASAP7_75t_L g2415 ( 
.A(n_2288),
.Y(n_2415)
);

AND2x2_ASAP7_75t_L g2416 ( 
.A(n_2191),
.B(n_1804),
.Y(n_2416)
);

INVx2_ASAP7_75t_L g2417 ( 
.A(n_2163),
.Y(n_2417)
);

NAND3xp33_ASAP7_75t_L g2418 ( 
.A(n_2159),
.B(n_2098),
.C(n_2102),
.Y(n_2418)
);

NAND2xp5_ASAP7_75t_L g2419 ( 
.A(n_2159),
.B(n_1760),
.Y(n_2419)
);

AND2x4_ASAP7_75t_L g2420 ( 
.A(n_2178),
.B(n_2098),
.Y(n_2420)
);

INVx1_ASAP7_75t_L g2421 ( 
.A(n_2163),
.Y(n_2421)
);

AND2x2_ASAP7_75t_L g2422 ( 
.A(n_2238),
.B(n_1804),
.Y(n_2422)
);

OR2x2_ASAP7_75t_L g2423 ( 
.A(n_2233),
.B(n_1777),
.Y(n_2423)
);

INVx1_ASAP7_75t_L g2424 ( 
.A(n_2380),
.Y(n_2424)
);

INVx2_ASAP7_75t_L g2425 ( 
.A(n_2293),
.Y(n_2425)
);

OR2x2_ASAP7_75t_L g2426 ( 
.A(n_2314),
.B(n_2161),
.Y(n_2426)
);

INVx1_ASAP7_75t_L g2427 ( 
.A(n_2411),
.Y(n_2427)
);

NAND2xp5_ASAP7_75t_L g2428 ( 
.A(n_2332),
.B(n_2200),
.Y(n_2428)
);

HB1xp67_ASAP7_75t_L g2429 ( 
.A(n_2341),
.Y(n_2429)
);

AND2x4_ASAP7_75t_L g2430 ( 
.A(n_2294),
.B(n_2194),
.Y(n_2430)
);

NAND2xp5_ASAP7_75t_L g2431 ( 
.A(n_2332),
.B(n_2269),
.Y(n_2431)
);

NAND2xp5_ASAP7_75t_L g2432 ( 
.A(n_2415),
.B(n_2269),
.Y(n_2432)
);

INVx1_ASAP7_75t_L g2433 ( 
.A(n_2299),
.Y(n_2433)
);

INVx2_ASAP7_75t_SL g2434 ( 
.A(n_2321),
.Y(n_2434)
);

NAND2xp5_ASAP7_75t_L g2435 ( 
.A(n_2295),
.B(n_2229),
.Y(n_2435)
);

INVx1_ASAP7_75t_L g2436 ( 
.A(n_2299),
.Y(n_2436)
);

HB1xp67_ASAP7_75t_L g2437 ( 
.A(n_2304),
.Y(n_2437)
);

NAND2x1p5_ASAP7_75t_L g2438 ( 
.A(n_2293),
.B(n_2194),
.Y(n_2438)
);

INVx2_ASAP7_75t_SL g2439 ( 
.A(n_2321),
.Y(n_2439)
);

AND2x2_ASAP7_75t_L g2440 ( 
.A(n_2400),
.B(n_2285),
.Y(n_2440)
);

INVx3_ASAP7_75t_L g2441 ( 
.A(n_2293),
.Y(n_2441)
);

OR2x2_ASAP7_75t_L g2442 ( 
.A(n_2419),
.B(n_2237),
.Y(n_2442)
);

INVx1_ASAP7_75t_L g2443 ( 
.A(n_2302),
.Y(n_2443)
);

INVx2_ASAP7_75t_L g2444 ( 
.A(n_2306),
.Y(n_2444)
);

INVx2_ASAP7_75t_L g2445 ( 
.A(n_2306),
.Y(n_2445)
);

INVx1_ASAP7_75t_L g2446 ( 
.A(n_2302),
.Y(n_2446)
);

AND2x2_ASAP7_75t_L g2447 ( 
.A(n_2400),
.B(n_2285),
.Y(n_2447)
);

INVx2_ASAP7_75t_L g2448 ( 
.A(n_2317),
.Y(n_2448)
);

INVx1_ASAP7_75t_L g2449 ( 
.A(n_2305),
.Y(n_2449)
);

NOR2xp67_ASAP7_75t_SL g2450 ( 
.A(n_2303),
.B(n_2207),
.Y(n_2450)
);

NAND2xp5_ASAP7_75t_SL g2451 ( 
.A(n_2294),
.B(n_2174),
.Y(n_2451)
);

INVx1_ASAP7_75t_L g2452 ( 
.A(n_2305),
.Y(n_2452)
);

AND2x2_ASAP7_75t_L g2453 ( 
.A(n_2407),
.B(n_2186),
.Y(n_2453)
);

NOR2x1_ASAP7_75t_L g2454 ( 
.A(n_2303),
.B(n_2193),
.Y(n_2454)
);

INVx1_ASAP7_75t_L g2455 ( 
.A(n_2309),
.Y(n_2455)
);

OR2x2_ASAP7_75t_L g2456 ( 
.A(n_2315),
.B(n_2272),
.Y(n_2456)
);

INVx1_ASAP7_75t_L g2457 ( 
.A(n_2309),
.Y(n_2457)
);

INVxp67_ASAP7_75t_L g2458 ( 
.A(n_2296),
.Y(n_2458)
);

INVx2_ASAP7_75t_L g2459 ( 
.A(n_2317),
.Y(n_2459)
);

NAND2xp5_ASAP7_75t_L g2460 ( 
.A(n_2295),
.B(n_2229),
.Y(n_2460)
);

OR2x2_ASAP7_75t_L g2461 ( 
.A(n_2308),
.B(n_2188),
.Y(n_2461)
);

INVx1_ASAP7_75t_L g2462 ( 
.A(n_2310),
.Y(n_2462)
);

INVx2_ASAP7_75t_L g2463 ( 
.A(n_2336),
.Y(n_2463)
);

NOR2x1_ASAP7_75t_L g2464 ( 
.A(n_2363),
.B(n_2193),
.Y(n_2464)
);

INVxp67_ASAP7_75t_SL g2465 ( 
.A(n_2379),
.Y(n_2465)
);

OR2x2_ASAP7_75t_L g2466 ( 
.A(n_2370),
.B(n_2399),
.Y(n_2466)
);

AND2x2_ASAP7_75t_L g2467 ( 
.A(n_2407),
.B(n_2248),
.Y(n_2467)
);

AND2x2_ASAP7_75t_L g2468 ( 
.A(n_2347),
.B(n_2248),
.Y(n_2468)
);

AND2x2_ASAP7_75t_L g2469 ( 
.A(n_2347),
.B(n_2143),
.Y(n_2469)
);

INVx1_ASAP7_75t_L g2470 ( 
.A(n_2310),
.Y(n_2470)
);

INVx3_ASAP7_75t_L g2471 ( 
.A(n_2294),
.Y(n_2471)
);

AND2x4_ASAP7_75t_L g2472 ( 
.A(n_2294),
.B(n_2194),
.Y(n_2472)
);

OR2x2_ASAP7_75t_L g2473 ( 
.A(n_2370),
.B(n_2281),
.Y(n_2473)
);

INVx1_ASAP7_75t_L g2474 ( 
.A(n_2311),
.Y(n_2474)
);

INVxp67_ASAP7_75t_L g2475 ( 
.A(n_2357),
.Y(n_2475)
);

INVx2_ASAP7_75t_L g2476 ( 
.A(n_2336),
.Y(n_2476)
);

INVx4_ASAP7_75t_L g2477 ( 
.A(n_2321),
.Y(n_2477)
);

OAI32xp33_ASAP7_75t_L g2478 ( 
.A1(n_2301),
.A2(n_2418),
.A3(n_2344),
.B1(n_2312),
.B2(n_2227),
.Y(n_2478)
);

INVx1_ASAP7_75t_L g2479 ( 
.A(n_2311),
.Y(n_2479)
);

AND2x2_ASAP7_75t_L g2480 ( 
.A(n_2292),
.B(n_2172),
.Y(n_2480)
);

NAND2xp5_ASAP7_75t_L g2481 ( 
.A(n_2292),
.B(n_2239),
.Y(n_2481)
);

INVx1_ASAP7_75t_L g2482 ( 
.A(n_2327),
.Y(n_2482)
);

HB1xp67_ASAP7_75t_L g2483 ( 
.A(n_2363),
.Y(n_2483)
);

INVx2_ASAP7_75t_L g2484 ( 
.A(n_2344),
.Y(n_2484)
);

AND2x4_ASAP7_75t_L g2485 ( 
.A(n_2344),
.B(n_2194),
.Y(n_2485)
);

NAND2xp5_ASAP7_75t_L g2486 ( 
.A(n_2361),
.B(n_2374),
.Y(n_2486)
);

INVxp67_ASAP7_75t_L g2487 ( 
.A(n_2297),
.Y(n_2487)
);

NAND2xp5_ASAP7_75t_L g2488 ( 
.A(n_2361),
.B(n_2239),
.Y(n_2488)
);

INVx1_ASAP7_75t_L g2489 ( 
.A(n_2327),
.Y(n_2489)
);

INVx1_ASAP7_75t_L g2490 ( 
.A(n_2330),
.Y(n_2490)
);

AND2x2_ASAP7_75t_L g2491 ( 
.A(n_2300),
.B(n_2172),
.Y(n_2491)
);

INVx1_ASAP7_75t_L g2492 ( 
.A(n_2330),
.Y(n_2492)
);

AND2x2_ASAP7_75t_L g2493 ( 
.A(n_2300),
.B(n_2183),
.Y(n_2493)
);

INVx2_ASAP7_75t_L g2494 ( 
.A(n_2417),
.Y(n_2494)
);

OAI33xp33_ASAP7_75t_L g2495 ( 
.A1(n_2392),
.A2(n_2136),
.A3(n_2264),
.B1(n_2279),
.B2(n_2284),
.B3(n_2289),
.Y(n_2495)
);

INVx2_ASAP7_75t_L g2496 ( 
.A(n_2417),
.Y(n_2496)
);

INVx1_ASAP7_75t_L g2497 ( 
.A(n_2331),
.Y(n_2497)
);

NAND2xp5_ASAP7_75t_L g2498 ( 
.A(n_2386),
.B(n_2239),
.Y(n_2498)
);

AND2x2_ASAP7_75t_L g2499 ( 
.A(n_2355),
.B(n_2183),
.Y(n_2499)
);

AND2x4_ASAP7_75t_SL g2500 ( 
.A(n_2385),
.B(n_2238),
.Y(n_2500)
);

AND2x2_ASAP7_75t_L g2501 ( 
.A(n_2355),
.B(n_2152),
.Y(n_2501)
);

AND2x2_ASAP7_75t_L g2502 ( 
.A(n_2358),
.B(n_2152),
.Y(n_2502)
);

INVx2_ASAP7_75t_L g2503 ( 
.A(n_2348),
.Y(n_2503)
);

BUFx2_ASAP7_75t_L g2504 ( 
.A(n_2385),
.Y(n_2504)
);

NAND2xp5_ASAP7_75t_L g2505 ( 
.A(n_2387),
.B(n_2291),
.Y(n_2505)
);

OR2x6_ASAP7_75t_L g2506 ( 
.A(n_2321),
.B(n_2207),
.Y(n_2506)
);

INVx2_ASAP7_75t_L g2507 ( 
.A(n_2348),
.Y(n_2507)
);

HB1xp67_ASAP7_75t_L g2508 ( 
.A(n_2387),
.Y(n_2508)
);

INVx1_ASAP7_75t_L g2509 ( 
.A(n_2331),
.Y(n_2509)
);

OR2x2_ASAP7_75t_L g2510 ( 
.A(n_2405),
.B(n_2170),
.Y(n_2510)
);

NAND2xp5_ASAP7_75t_L g2511 ( 
.A(n_2337),
.B(n_2194),
.Y(n_2511)
);

AND2x2_ASAP7_75t_L g2512 ( 
.A(n_2358),
.B(n_2152),
.Y(n_2512)
);

HB1xp67_ASAP7_75t_L g2513 ( 
.A(n_2337),
.Y(n_2513)
);

INVx2_ASAP7_75t_L g2514 ( 
.A(n_2366),
.Y(n_2514)
);

INVx1_ASAP7_75t_L g2515 ( 
.A(n_2338),
.Y(n_2515)
);

INVx1_ASAP7_75t_L g2516 ( 
.A(n_2338),
.Y(n_2516)
);

INVx1_ASAP7_75t_L g2517 ( 
.A(n_2339),
.Y(n_2517)
);

INVx1_ASAP7_75t_L g2518 ( 
.A(n_2339),
.Y(n_2518)
);

OR2x2_ASAP7_75t_L g2519 ( 
.A(n_2399),
.B(n_2230),
.Y(n_2519)
);

OR2x2_ASAP7_75t_L g2520 ( 
.A(n_2364),
.B(n_2255),
.Y(n_2520)
);

AOI21xp33_ASAP7_75t_SL g2521 ( 
.A1(n_2297),
.A2(n_2234),
.B(n_2262),
.Y(n_2521)
);

AND2x2_ASAP7_75t_L g2522 ( 
.A(n_2343),
.B(n_2177),
.Y(n_2522)
);

OR2x2_ASAP7_75t_L g2523 ( 
.A(n_2408),
.B(n_2282),
.Y(n_2523)
);

NOR2xp33_ASAP7_75t_L g2524 ( 
.A(n_2385),
.B(n_2137),
.Y(n_2524)
);

OAI21xp5_ASAP7_75t_L g2525 ( 
.A1(n_2298),
.A2(n_2226),
.B(n_2205),
.Y(n_2525)
);

INVx2_ASAP7_75t_L g2526 ( 
.A(n_2366),
.Y(n_2526)
);

INVx2_ASAP7_75t_L g2527 ( 
.A(n_2367),
.Y(n_2527)
);

NAND2xp5_ASAP7_75t_L g2528 ( 
.A(n_2342),
.B(n_2177),
.Y(n_2528)
);

INVxp67_ASAP7_75t_L g2529 ( 
.A(n_2333),
.Y(n_2529)
);

AOI21xp33_ASAP7_75t_L g2530 ( 
.A1(n_2342),
.A2(n_2286),
.B(n_2185),
.Y(n_2530)
);

AND2x2_ASAP7_75t_L g2531 ( 
.A(n_2343),
.B(n_2177),
.Y(n_2531)
);

NAND2x1_ASAP7_75t_L g2532 ( 
.A(n_2385),
.B(n_2238),
.Y(n_2532)
);

AND2x2_ASAP7_75t_L g2533 ( 
.A(n_2395),
.B(n_2257),
.Y(n_2533)
);

NAND2xp5_ASAP7_75t_L g2534 ( 
.A(n_2345),
.B(n_2135),
.Y(n_2534)
);

INVx2_ASAP7_75t_L g2535 ( 
.A(n_2367),
.Y(n_2535)
);

INVx2_ASAP7_75t_L g2536 ( 
.A(n_2369),
.Y(n_2536)
);

AOI21xp5_ASAP7_75t_L g2537 ( 
.A1(n_2404),
.A2(n_2242),
.B(n_1998),
.Y(n_2537)
);

INVxp67_ASAP7_75t_SL g2538 ( 
.A(n_2414),
.Y(n_2538)
);

INVx2_ASAP7_75t_L g2539 ( 
.A(n_2369),
.Y(n_2539)
);

INVx1_ASAP7_75t_SL g2540 ( 
.A(n_2321),
.Y(n_2540)
);

NOR2x1p5_ASAP7_75t_L g2541 ( 
.A(n_2420),
.B(n_2253),
.Y(n_2541)
);

INVx1_ASAP7_75t_L g2542 ( 
.A(n_2345),
.Y(n_2542)
);

AND2x2_ASAP7_75t_L g2543 ( 
.A(n_2395),
.B(n_2257),
.Y(n_2543)
);

OR2x2_ASAP7_75t_L g2544 ( 
.A(n_2364),
.B(n_2326),
.Y(n_2544)
);

OA211x2_ASAP7_75t_L g2545 ( 
.A1(n_2324),
.A2(n_2242),
.B(n_2174),
.C(n_2226),
.Y(n_2545)
);

NAND4xp25_ASAP7_75t_L g2546 ( 
.A(n_2378),
.B(n_2222),
.C(n_2253),
.D(n_2266),
.Y(n_2546)
);

AND2x2_ASAP7_75t_L g2547 ( 
.A(n_2409),
.B(n_2265),
.Y(n_2547)
);

AND2x2_ASAP7_75t_L g2548 ( 
.A(n_2409),
.B(n_2265),
.Y(n_2548)
);

NAND2xp5_ASAP7_75t_L g2549 ( 
.A(n_2351),
.B(n_2135),
.Y(n_2549)
);

INVx2_ASAP7_75t_L g2550 ( 
.A(n_2441),
.Y(n_2550)
);

INVx1_ASAP7_75t_L g2551 ( 
.A(n_2513),
.Y(n_2551)
);

INVx1_ASAP7_75t_L g2552 ( 
.A(n_2429),
.Y(n_2552)
);

OR2x2_ASAP7_75t_L g2553 ( 
.A(n_2473),
.B(n_2412),
.Y(n_2553)
);

NOR2xp33_ASAP7_75t_L g2554 ( 
.A(n_2477),
.B(n_2402),
.Y(n_2554)
);

BUFx3_ASAP7_75t_L g2555 ( 
.A(n_2471),
.Y(n_2555)
);

AND2x2_ASAP7_75t_L g2556 ( 
.A(n_2499),
.B(n_2398),
.Y(n_2556)
);

AOI33xp33_ASAP7_75t_L g2557 ( 
.A1(n_2424),
.A2(n_2427),
.A3(n_2447),
.B1(n_2440),
.B2(n_2493),
.B3(n_2467),
.Y(n_2557)
);

AND2x4_ASAP7_75t_L g2558 ( 
.A(n_2471),
.B(n_2402),
.Y(n_2558)
);

BUFx12f_ASAP7_75t_L g2559 ( 
.A(n_2477),
.Y(n_2559)
);

OAI21xp33_ASAP7_75t_L g2560 ( 
.A1(n_2525),
.A2(n_2316),
.B(n_2410),
.Y(n_2560)
);

INVx1_ASAP7_75t_L g2561 ( 
.A(n_2466),
.Y(n_2561)
);

INVx4_ASAP7_75t_L g2562 ( 
.A(n_2477),
.Y(n_2562)
);

AND2x2_ASAP7_75t_L g2563 ( 
.A(n_2499),
.B(n_2493),
.Y(n_2563)
);

AND2x2_ASAP7_75t_L g2564 ( 
.A(n_2533),
.B(n_2398),
.Y(n_2564)
);

AND2x4_ASAP7_75t_L g2565 ( 
.A(n_2471),
.B(n_2388),
.Y(n_2565)
);

AND2x2_ASAP7_75t_L g2566 ( 
.A(n_2533),
.B(n_2388),
.Y(n_2566)
);

BUFx3_ASAP7_75t_L g2567 ( 
.A(n_2430),
.Y(n_2567)
);

INVx1_ASAP7_75t_L g2568 ( 
.A(n_2425),
.Y(n_2568)
);

AND2x2_ASAP7_75t_L g2569 ( 
.A(n_2543),
.B(n_2393),
.Y(n_2569)
);

INVx1_ASAP7_75t_L g2570 ( 
.A(n_2425),
.Y(n_2570)
);

AND2x4_ASAP7_75t_L g2571 ( 
.A(n_2541),
.B(n_2393),
.Y(n_2571)
);

INVx1_ASAP7_75t_SL g2572 ( 
.A(n_2453),
.Y(n_2572)
);

INVx6_ASAP7_75t_L g2573 ( 
.A(n_2430),
.Y(n_2573)
);

AND2x2_ASAP7_75t_L g2574 ( 
.A(n_2543),
.B(n_2547),
.Y(n_2574)
);

INVx1_ASAP7_75t_L g2575 ( 
.A(n_2466),
.Y(n_2575)
);

INVx2_ASAP7_75t_SL g2576 ( 
.A(n_2500),
.Y(n_2576)
);

INVx1_ASAP7_75t_L g2577 ( 
.A(n_2441),
.Y(n_2577)
);

OAI33xp33_ASAP7_75t_L g2578 ( 
.A1(n_2432),
.A2(n_2396),
.A3(n_2373),
.B1(n_2381),
.B2(n_2351),
.B3(n_2353),
.Y(n_2578)
);

OR2x6_ASAP7_75t_L g2579 ( 
.A(n_2484),
.B(n_2382),
.Y(n_2579)
);

INVx1_ASAP7_75t_L g2580 ( 
.A(n_2441),
.Y(n_2580)
);

NAND2xp5_ASAP7_75t_L g2581 ( 
.A(n_2465),
.B(n_2353),
.Y(n_2581)
);

HB1xp67_ASAP7_75t_L g2582 ( 
.A(n_2487),
.Y(n_2582)
);

NAND2xp5_ASAP7_75t_L g2583 ( 
.A(n_2467),
.B(n_2356),
.Y(n_2583)
);

INVx1_ASAP7_75t_SL g2584 ( 
.A(n_2453),
.Y(n_2584)
);

AND2x4_ASAP7_75t_L g2585 ( 
.A(n_2430),
.B(n_2352),
.Y(n_2585)
);

NAND2xp5_ASAP7_75t_L g2586 ( 
.A(n_2440),
.B(n_2356),
.Y(n_2586)
);

INVx2_ASAP7_75t_L g2587 ( 
.A(n_2504),
.Y(n_2587)
);

AND2x2_ASAP7_75t_L g2588 ( 
.A(n_2547),
.B(n_2320),
.Y(n_2588)
);

AND2x2_ASAP7_75t_L g2589 ( 
.A(n_2548),
.B(n_2320),
.Y(n_2589)
);

OR2x2_ASAP7_75t_L g2590 ( 
.A(n_2473),
.B(n_2412),
.Y(n_2590)
);

NAND2xp5_ASAP7_75t_L g2591 ( 
.A(n_2447),
.B(n_2362),
.Y(n_2591)
);

INVx1_ASAP7_75t_L g2592 ( 
.A(n_2448),
.Y(n_2592)
);

NOR2xp33_ASAP7_75t_L g2593 ( 
.A(n_2458),
.B(n_2352),
.Y(n_2593)
);

INVx3_ASAP7_75t_L g2594 ( 
.A(n_2532),
.Y(n_2594)
);

AND2x2_ASAP7_75t_L g2595 ( 
.A(n_2548),
.B(n_2346),
.Y(n_2595)
);

NAND2xp5_ASAP7_75t_L g2596 ( 
.A(n_2437),
.B(n_2362),
.Y(n_2596)
);

INVx1_ASAP7_75t_L g2597 ( 
.A(n_2519),
.Y(n_2597)
);

INVx1_ASAP7_75t_L g2598 ( 
.A(n_2519),
.Y(n_2598)
);

INVx1_ASAP7_75t_L g2599 ( 
.A(n_2448),
.Y(n_2599)
);

INVx1_ASAP7_75t_L g2600 ( 
.A(n_2459),
.Y(n_2600)
);

INVx2_ASAP7_75t_L g2601 ( 
.A(n_2468),
.Y(n_2601)
);

NAND2xp5_ASAP7_75t_L g2602 ( 
.A(n_2484),
.B(n_2368),
.Y(n_2602)
);

BUFx3_ASAP7_75t_L g2603 ( 
.A(n_2472),
.Y(n_2603)
);

INVx1_ASAP7_75t_SL g2604 ( 
.A(n_2500),
.Y(n_2604)
);

INVx1_ASAP7_75t_L g2605 ( 
.A(n_2459),
.Y(n_2605)
);

AND2x2_ASAP7_75t_L g2606 ( 
.A(n_2468),
.B(n_2346),
.Y(n_2606)
);

NAND2xp5_ASAP7_75t_L g2607 ( 
.A(n_2486),
.B(n_2368),
.Y(n_2607)
);

AND2x2_ASAP7_75t_L g2608 ( 
.A(n_2472),
.B(n_2416),
.Y(n_2608)
);

OR2x2_ASAP7_75t_L g2609 ( 
.A(n_2431),
.B(n_2373),
.Y(n_2609)
);

INVx3_ASAP7_75t_L g2610 ( 
.A(n_2472),
.Y(n_2610)
);

NAND2xp5_ASAP7_75t_L g2611 ( 
.A(n_2524),
.B(n_2381),
.Y(n_2611)
);

INVx1_ASAP7_75t_L g2612 ( 
.A(n_2463),
.Y(n_2612)
);

INVx1_ASAP7_75t_L g2613 ( 
.A(n_2463),
.Y(n_2613)
);

OR2x6_ASAP7_75t_L g2614 ( 
.A(n_2529),
.B(n_2382),
.Y(n_2614)
);

INVx1_ASAP7_75t_L g2615 ( 
.A(n_2476),
.Y(n_2615)
);

NAND2xp5_ASAP7_75t_L g2616 ( 
.A(n_2524),
.B(n_2389),
.Y(n_2616)
);

INVx2_ASAP7_75t_L g2617 ( 
.A(n_2444),
.Y(n_2617)
);

INVxp67_ASAP7_75t_L g2618 ( 
.A(n_2491),
.Y(n_2618)
);

AND2x2_ASAP7_75t_L g2619 ( 
.A(n_2480),
.B(n_2416),
.Y(n_2619)
);

INVx1_ASAP7_75t_L g2620 ( 
.A(n_2476),
.Y(n_2620)
);

XOR2xp5_ASAP7_75t_L g2621 ( 
.A(n_2456),
.B(n_1015),
.Y(n_2621)
);

AND2x2_ASAP7_75t_L g2622 ( 
.A(n_2480),
.B(n_2350),
.Y(n_2622)
);

INVx4_ASAP7_75t_L g2623 ( 
.A(n_2506),
.Y(n_2623)
);

HB1xp67_ASAP7_75t_L g2624 ( 
.A(n_2483),
.Y(n_2624)
);

AOI22xp33_ASAP7_75t_L g2625 ( 
.A1(n_2545),
.A2(n_2495),
.B1(n_2204),
.B2(n_2442),
.Y(n_2625)
);

AND2x2_ASAP7_75t_L g2626 ( 
.A(n_2491),
.B(n_2350),
.Y(n_2626)
);

INVx1_ASAP7_75t_L g2627 ( 
.A(n_2520),
.Y(n_2627)
);

BUFx2_ASAP7_75t_L g2628 ( 
.A(n_2428),
.Y(n_2628)
);

NOR3xp33_ASAP7_75t_L g2629 ( 
.A(n_2478),
.B(n_2421),
.C(n_2420),
.Y(n_2629)
);

INVx3_ASAP7_75t_L g2630 ( 
.A(n_2485),
.Y(n_2630)
);

AOI22xp33_ASAP7_75t_L g2631 ( 
.A1(n_2442),
.A2(n_2204),
.B1(n_2420),
.B2(n_2220),
.Y(n_2631)
);

AND2x2_ASAP7_75t_L g2632 ( 
.A(n_2469),
.B(n_2354),
.Y(n_2632)
);

INVx1_ASAP7_75t_L g2633 ( 
.A(n_2520),
.Y(n_2633)
);

BUFx3_ASAP7_75t_L g2634 ( 
.A(n_2498),
.Y(n_2634)
);

AND2x2_ASAP7_75t_L g2635 ( 
.A(n_2469),
.B(n_2501),
.Y(n_2635)
);

INVx2_ASAP7_75t_L g2636 ( 
.A(n_2444),
.Y(n_2636)
);

INVx2_ASAP7_75t_L g2637 ( 
.A(n_2445),
.Y(n_2637)
);

INVx2_ASAP7_75t_L g2638 ( 
.A(n_2445),
.Y(n_2638)
);

INVx1_ASAP7_75t_L g2639 ( 
.A(n_2508),
.Y(n_2639)
);

INVx1_ASAP7_75t_SL g2640 ( 
.A(n_2451),
.Y(n_2640)
);

INVx1_ASAP7_75t_SL g2641 ( 
.A(n_2451),
.Y(n_2641)
);

INVx1_ASAP7_75t_L g2642 ( 
.A(n_2433),
.Y(n_2642)
);

AND2x2_ASAP7_75t_L g2643 ( 
.A(n_2501),
.B(n_2354),
.Y(n_2643)
);

INVx1_ASAP7_75t_L g2644 ( 
.A(n_2436),
.Y(n_2644)
);

INVx2_ASAP7_75t_L g2645 ( 
.A(n_2502),
.Y(n_2645)
);

INVx2_ASAP7_75t_SL g2646 ( 
.A(n_2485),
.Y(n_2646)
);

AND2x2_ASAP7_75t_L g2647 ( 
.A(n_2502),
.B(n_2340),
.Y(n_2647)
);

AND2x2_ASAP7_75t_L g2648 ( 
.A(n_2512),
.B(n_2340),
.Y(n_2648)
);

BUFx3_ASAP7_75t_L g2649 ( 
.A(n_2434),
.Y(n_2649)
);

INVx1_ASAP7_75t_L g2650 ( 
.A(n_2443),
.Y(n_2650)
);

INVx1_ASAP7_75t_L g2651 ( 
.A(n_2446),
.Y(n_2651)
);

INVx2_ASAP7_75t_L g2652 ( 
.A(n_2512),
.Y(n_2652)
);

NAND2xp5_ASAP7_75t_L g2653 ( 
.A(n_2534),
.B(n_2389),
.Y(n_2653)
);

OR2x2_ASAP7_75t_L g2654 ( 
.A(n_2544),
.B(n_2390),
.Y(n_2654)
);

INVx1_ASAP7_75t_L g2655 ( 
.A(n_2449),
.Y(n_2655)
);

INVx1_ASAP7_75t_L g2656 ( 
.A(n_2452),
.Y(n_2656)
);

INVx2_ASAP7_75t_L g2657 ( 
.A(n_2522),
.Y(n_2657)
);

INVx3_ASAP7_75t_L g2658 ( 
.A(n_2485),
.Y(n_2658)
);

INVx1_ASAP7_75t_SL g2659 ( 
.A(n_2481),
.Y(n_2659)
);

AND2x2_ASAP7_75t_L g2660 ( 
.A(n_2522),
.B(n_2313),
.Y(n_2660)
);

INVx1_ASAP7_75t_L g2661 ( 
.A(n_2455),
.Y(n_2661)
);

INVx2_ASAP7_75t_L g2662 ( 
.A(n_2531),
.Y(n_2662)
);

INVx1_ASAP7_75t_L g2663 ( 
.A(n_2457),
.Y(n_2663)
);

INVx1_ASAP7_75t_L g2664 ( 
.A(n_2574),
.Y(n_2664)
);

NAND2xp5_ASAP7_75t_L g2665 ( 
.A(n_2563),
.B(n_2549),
.Y(n_2665)
);

INVx1_ASAP7_75t_L g2666 ( 
.A(n_2574),
.Y(n_2666)
);

INVx1_ASAP7_75t_L g2667 ( 
.A(n_2563),
.Y(n_2667)
);

INVx1_ASAP7_75t_L g2668 ( 
.A(n_2624),
.Y(n_2668)
);

OR2x2_ASAP7_75t_L g2669 ( 
.A(n_2601),
.B(n_2426),
.Y(n_2669)
);

AND2x2_ASAP7_75t_L g2670 ( 
.A(n_2635),
.B(n_2454),
.Y(n_2670)
);

INVx1_ASAP7_75t_L g2671 ( 
.A(n_2601),
.Y(n_2671)
);

NAND2xp5_ASAP7_75t_L g2672 ( 
.A(n_2606),
.B(n_2435),
.Y(n_2672)
);

OR2x2_ASAP7_75t_L g2673 ( 
.A(n_2553),
.B(n_2460),
.Y(n_2673)
);

NAND2xp5_ASAP7_75t_L g2674 ( 
.A(n_2606),
.B(n_2572),
.Y(n_2674)
);

NAND2xp5_ASAP7_75t_L g2675 ( 
.A(n_2584),
.B(n_2505),
.Y(n_2675)
);

AND2x2_ASAP7_75t_L g2676 ( 
.A(n_2635),
.B(n_2531),
.Y(n_2676)
);

INVx1_ASAP7_75t_L g2677 ( 
.A(n_2582),
.Y(n_2677)
);

INVx1_ASAP7_75t_L g2678 ( 
.A(n_2564),
.Y(n_2678)
);

INVx2_ASAP7_75t_L g2679 ( 
.A(n_2555),
.Y(n_2679)
);

NAND2xp5_ASAP7_75t_L g2680 ( 
.A(n_2564),
.B(n_2544),
.Y(n_2680)
);

INVx2_ASAP7_75t_L g2681 ( 
.A(n_2555),
.Y(n_2681)
);

INVx1_ASAP7_75t_L g2682 ( 
.A(n_2566),
.Y(n_2682)
);

OR2x2_ASAP7_75t_L g2683 ( 
.A(n_2553),
.B(n_2523),
.Y(n_2683)
);

AND2x2_ASAP7_75t_L g2684 ( 
.A(n_2632),
.B(n_2540),
.Y(n_2684)
);

AND2x2_ASAP7_75t_L g2685 ( 
.A(n_2632),
.B(n_2434),
.Y(n_2685)
);

OR2x4_ASAP7_75t_L g2686 ( 
.A(n_2593),
.B(n_2488),
.Y(n_2686)
);

INVx1_ASAP7_75t_L g2687 ( 
.A(n_2566),
.Y(n_2687)
);

INVx1_ASAP7_75t_SL g2688 ( 
.A(n_2640),
.Y(n_2688)
);

AND2x2_ASAP7_75t_L g2689 ( 
.A(n_2556),
.B(n_2439),
.Y(n_2689)
);

OR2x2_ASAP7_75t_L g2690 ( 
.A(n_2590),
.B(n_2510),
.Y(n_2690)
);

AND2x2_ASAP7_75t_L g2691 ( 
.A(n_2556),
.B(n_2439),
.Y(n_2691)
);

AND2x2_ASAP7_75t_L g2692 ( 
.A(n_2626),
.B(n_2475),
.Y(n_2692)
);

INVx1_ASAP7_75t_L g2693 ( 
.A(n_2569),
.Y(n_2693)
);

INVx1_ASAP7_75t_SL g2694 ( 
.A(n_2641),
.Y(n_2694)
);

INVxp67_ASAP7_75t_SL g2695 ( 
.A(n_2618),
.Y(n_2695)
);

AND2x2_ASAP7_75t_L g2696 ( 
.A(n_2626),
.B(n_2595),
.Y(n_2696)
);

NAND2xp5_ASAP7_75t_L g2697 ( 
.A(n_2595),
.B(n_2461),
.Y(n_2697)
);

OR2x2_ASAP7_75t_L g2698 ( 
.A(n_2590),
.B(n_2546),
.Y(n_2698)
);

INVx1_ASAP7_75t_SL g2699 ( 
.A(n_2604),
.Y(n_2699)
);

AND2x2_ASAP7_75t_L g2700 ( 
.A(n_2569),
.B(n_2506),
.Y(n_2700)
);

AOI21xp5_ASAP7_75t_L g2701 ( 
.A1(n_2560),
.A2(n_2537),
.B(n_2530),
.Y(n_2701)
);

AND2x2_ASAP7_75t_L g2702 ( 
.A(n_2622),
.B(n_2506),
.Y(n_2702)
);

HB1xp67_ASAP7_75t_L g2703 ( 
.A(n_2628),
.Y(n_2703)
);

HB1xp67_ASAP7_75t_L g2704 ( 
.A(n_2628),
.Y(n_2704)
);

NOR2x1_ASAP7_75t_L g2705 ( 
.A(n_2623),
.B(n_2506),
.Y(n_2705)
);

INVxp67_ASAP7_75t_SL g2706 ( 
.A(n_2594),
.Y(n_2706)
);

AND2x2_ASAP7_75t_L g2707 ( 
.A(n_2622),
.B(n_2521),
.Y(n_2707)
);

OR2x2_ASAP7_75t_L g2708 ( 
.A(n_2597),
.B(n_2528),
.Y(n_2708)
);

OR2x2_ASAP7_75t_L g2709 ( 
.A(n_2598),
.B(n_2335),
.Y(n_2709)
);

INVx1_ASAP7_75t_L g2710 ( 
.A(n_2575),
.Y(n_2710)
);

AND2x2_ASAP7_75t_L g2711 ( 
.A(n_2619),
.B(n_2313),
.Y(n_2711)
);

INVx1_ASAP7_75t_L g2712 ( 
.A(n_2575),
.Y(n_2712)
);

INVx1_ASAP7_75t_L g2713 ( 
.A(n_2654),
.Y(n_2713)
);

OR2x2_ASAP7_75t_L g2714 ( 
.A(n_2627),
.B(n_2335),
.Y(n_2714)
);

AOI22xp33_ASAP7_75t_L g2715 ( 
.A1(n_2629),
.A2(n_2496),
.B1(n_2503),
.B2(n_2494),
.Y(n_2715)
);

AND2x4_ASAP7_75t_L g2716 ( 
.A(n_2594),
.B(n_2464),
.Y(n_2716)
);

AND2x2_ASAP7_75t_L g2717 ( 
.A(n_2619),
.B(n_2318),
.Y(n_2717)
);

INVx1_ASAP7_75t_L g2718 ( 
.A(n_2654),
.Y(n_2718)
);

AND2x2_ASAP7_75t_L g2719 ( 
.A(n_2643),
.B(n_2588),
.Y(n_2719)
);

INVx1_ASAP7_75t_L g2720 ( 
.A(n_2587),
.Y(n_2720)
);

OR2x2_ASAP7_75t_L g2721 ( 
.A(n_2633),
.B(n_2586),
.Y(n_2721)
);

INVx1_ASAP7_75t_L g2722 ( 
.A(n_2587),
.Y(n_2722)
);

INVx1_ASAP7_75t_L g2723 ( 
.A(n_2639),
.Y(n_2723)
);

INVxp67_ASAP7_75t_L g2724 ( 
.A(n_2576),
.Y(n_2724)
);

OR2x2_ASAP7_75t_L g2725 ( 
.A(n_2591),
.B(n_2390),
.Y(n_2725)
);

INVx2_ASAP7_75t_L g2726 ( 
.A(n_2565),
.Y(n_2726)
);

OR2x6_ASAP7_75t_L g2727 ( 
.A(n_2623),
.B(n_2438),
.Y(n_2727)
);

NAND2xp5_ASAP7_75t_L g2728 ( 
.A(n_2588),
.B(n_2462),
.Y(n_2728)
);

INVx1_ASAP7_75t_L g2729 ( 
.A(n_2639),
.Y(n_2729)
);

AND2x2_ASAP7_75t_L g2730 ( 
.A(n_2643),
.B(n_2318),
.Y(n_2730)
);

INVx2_ASAP7_75t_L g2731 ( 
.A(n_2565),
.Y(n_2731)
);

NAND2xp5_ASAP7_75t_L g2732 ( 
.A(n_2589),
.B(n_2470),
.Y(n_2732)
);

AND2x2_ASAP7_75t_L g2733 ( 
.A(n_2589),
.B(n_2359),
.Y(n_2733)
);

NAND2xp5_ASAP7_75t_L g2734 ( 
.A(n_2645),
.B(n_2474),
.Y(n_2734)
);

INVx2_ASAP7_75t_SL g2735 ( 
.A(n_2573),
.Y(n_2735)
);

INVxp67_ASAP7_75t_L g2736 ( 
.A(n_2576),
.Y(n_2736)
);

INVx1_ASAP7_75t_L g2737 ( 
.A(n_2568),
.Y(n_2737)
);

AND2x2_ASAP7_75t_L g2738 ( 
.A(n_2660),
.B(n_2647),
.Y(n_2738)
);

HB1xp67_ASAP7_75t_L g2739 ( 
.A(n_2611),
.Y(n_2739)
);

AND2x2_ASAP7_75t_L g2740 ( 
.A(n_2660),
.B(n_2359),
.Y(n_2740)
);

AND2x2_ASAP7_75t_L g2741 ( 
.A(n_2647),
.B(n_2360),
.Y(n_2741)
);

INVx2_ASAP7_75t_L g2742 ( 
.A(n_2565),
.Y(n_2742)
);

OR2x2_ASAP7_75t_L g2743 ( 
.A(n_2561),
.B(n_2394),
.Y(n_2743)
);

NAND2xp5_ASAP7_75t_L g2744 ( 
.A(n_2645),
.B(n_2479),
.Y(n_2744)
);

NAND2xp5_ASAP7_75t_L g2745 ( 
.A(n_2652),
.B(n_2482),
.Y(n_2745)
);

NAND2x1p5_ASAP7_75t_L g2746 ( 
.A(n_2562),
.B(n_2450),
.Y(n_2746)
);

INVx1_ASAP7_75t_L g2747 ( 
.A(n_2568),
.Y(n_2747)
);

NAND2xp33_ASAP7_75t_SL g2748 ( 
.A(n_2616),
.B(n_2307),
.Y(n_2748)
);

OR2x2_ASAP7_75t_L g2749 ( 
.A(n_2583),
.B(n_2394),
.Y(n_2749)
);

NAND4xp25_ASAP7_75t_SL g2750 ( 
.A(n_2557),
.B(n_2319),
.C(n_2511),
.D(n_2490),
.Y(n_2750)
);

NAND2xp5_ASAP7_75t_L g2751 ( 
.A(n_2652),
.B(n_2489),
.Y(n_2751)
);

INVx1_ASAP7_75t_SL g2752 ( 
.A(n_2585),
.Y(n_2752)
);

INVx1_ASAP7_75t_L g2753 ( 
.A(n_2570),
.Y(n_2753)
);

INVx2_ASAP7_75t_SL g2754 ( 
.A(n_2573),
.Y(n_2754)
);

AND2x2_ASAP7_75t_L g2755 ( 
.A(n_2648),
.B(n_2608),
.Y(n_2755)
);

INVx1_ASAP7_75t_L g2756 ( 
.A(n_2696),
.Y(n_2756)
);

NAND2xp5_ASAP7_75t_SL g2757 ( 
.A(n_2703),
.B(n_2558),
.Y(n_2757)
);

OR2x2_ASAP7_75t_L g2758 ( 
.A(n_2683),
.B(n_2581),
.Y(n_2758)
);

AOI22xp5_ASAP7_75t_L g2759 ( 
.A1(n_2750),
.A2(n_2625),
.B1(n_2748),
.B2(n_2739),
.Y(n_2759)
);

OAI22xp5_ASAP7_75t_L g2760 ( 
.A1(n_2698),
.A2(n_2307),
.B1(n_2621),
.B2(n_2631),
.Y(n_2760)
);

OAI221xp5_ASAP7_75t_L g2761 ( 
.A1(n_2715),
.A2(n_2609),
.B1(n_2538),
.B2(n_2614),
.C(n_2594),
.Y(n_2761)
);

AND2x2_ASAP7_75t_L g2762 ( 
.A(n_2696),
.B(n_2608),
.Y(n_2762)
);

INVx1_ASAP7_75t_L g2763 ( 
.A(n_2703),
.Y(n_2763)
);

INVx1_ASAP7_75t_L g2764 ( 
.A(n_2704),
.Y(n_2764)
);

NAND2xp5_ASAP7_75t_L g2765 ( 
.A(n_2719),
.B(n_2657),
.Y(n_2765)
);

INVx1_ASAP7_75t_L g2766 ( 
.A(n_2704),
.Y(n_2766)
);

OAI221xp5_ASAP7_75t_L g2767 ( 
.A1(n_2715),
.A2(n_2609),
.B1(n_2614),
.B2(n_2596),
.C(n_2570),
.Y(n_2767)
);

OR2x2_ASAP7_75t_L g2768 ( 
.A(n_2690),
.B(n_2657),
.Y(n_2768)
);

INVx1_ASAP7_75t_L g2769 ( 
.A(n_2738),
.Y(n_2769)
);

NAND2xp5_ASAP7_75t_SL g2770 ( 
.A(n_2739),
.B(n_2558),
.Y(n_2770)
);

AOI22xp33_ASAP7_75t_L g2771 ( 
.A1(n_2748),
.A2(n_2701),
.B1(n_2707),
.B2(n_2578),
.Y(n_2771)
);

INVxp67_ASAP7_75t_L g2772 ( 
.A(n_2706),
.Y(n_2772)
);

OAI32xp33_ASAP7_75t_L g2773 ( 
.A1(n_2688),
.A2(n_2438),
.A3(n_2607),
.B1(n_2653),
.B2(n_2552),
.Y(n_2773)
);

OAI21xp5_ASAP7_75t_L g2774 ( 
.A1(n_2707),
.A2(n_2694),
.B(n_2738),
.Y(n_2774)
);

INVx1_ASAP7_75t_L g2775 ( 
.A(n_2719),
.Y(n_2775)
);

INVx1_ASAP7_75t_SL g2776 ( 
.A(n_2755),
.Y(n_2776)
);

INVx2_ASAP7_75t_L g2777 ( 
.A(n_2755),
.Y(n_2777)
);

OAI322xp33_ASAP7_75t_L g2778 ( 
.A1(n_2677),
.A2(n_2551),
.A3(n_2602),
.B1(n_2663),
.B2(n_2642),
.C1(n_2644),
.C2(n_2577),
.Y(n_2778)
);

OAI22xp5_ASAP7_75t_L g2779 ( 
.A1(n_2752),
.A2(n_2621),
.B1(n_2662),
.B2(n_2614),
.Y(n_2779)
);

AO221x1_ASAP7_75t_L g2780 ( 
.A1(n_2724),
.A2(n_2610),
.B1(n_2630),
.B2(n_2658),
.C(n_2662),
.Y(n_2780)
);

AOI22xp5_ASAP7_75t_L g2781 ( 
.A1(n_2699),
.A2(n_2571),
.B1(n_2676),
.B2(n_2713),
.Y(n_2781)
);

INVx1_ASAP7_75t_L g2782 ( 
.A(n_2711),
.Y(n_2782)
);

AOI211xp5_ASAP7_75t_L g2783 ( 
.A1(n_2673),
.A2(n_2551),
.B(n_2585),
.C(n_2659),
.Y(n_2783)
);

OAI21xp5_ASAP7_75t_L g2784 ( 
.A1(n_2676),
.A2(n_2585),
.B(n_2558),
.Y(n_2784)
);

INVxp67_ASAP7_75t_SL g2785 ( 
.A(n_2735),
.Y(n_2785)
);

INVx1_ASAP7_75t_L g2786 ( 
.A(n_2711),
.Y(n_2786)
);

INVx2_ASAP7_75t_L g2787 ( 
.A(n_2735),
.Y(n_2787)
);

NAND2xp5_ASAP7_75t_SL g2788 ( 
.A(n_2716),
.B(n_2610),
.Y(n_2788)
);

AOI21xp5_ASAP7_75t_SL g2789 ( 
.A1(n_2727),
.A2(n_2614),
.B(n_2623),
.Y(n_2789)
);

AND2x2_ASAP7_75t_L g2790 ( 
.A(n_2717),
.B(n_2648),
.Y(n_2790)
);

AND2x2_ASAP7_75t_L g2791 ( 
.A(n_2717),
.B(n_2571),
.Y(n_2791)
);

INVx1_ASAP7_75t_L g2792 ( 
.A(n_2674),
.Y(n_2792)
);

OAI211xp5_ASAP7_75t_L g2793 ( 
.A1(n_2695),
.A2(n_2562),
.B(n_2644),
.C(n_2642),
.Y(n_2793)
);

NOR2xp33_ASAP7_75t_SL g2794 ( 
.A(n_2692),
.B(n_2634),
.Y(n_2794)
);

INVx1_ASAP7_75t_L g2795 ( 
.A(n_2730),
.Y(n_2795)
);

INVx1_ASAP7_75t_L g2796 ( 
.A(n_2730),
.Y(n_2796)
);

AOI322xp5_ASAP7_75t_L g2797 ( 
.A1(n_2718),
.A2(n_2605),
.A3(n_2599),
.B1(n_2600),
.B2(n_2620),
.C1(n_2615),
.C2(n_2613),
.Y(n_2797)
);

INVx1_ASAP7_75t_L g2798 ( 
.A(n_2740),
.Y(n_2798)
);

INVx1_ASAP7_75t_L g2799 ( 
.A(n_2740),
.Y(n_2799)
);

INVxp67_ASAP7_75t_L g2800 ( 
.A(n_2754),
.Y(n_2800)
);

AND2x2_ASAP7_75t_L g2801 ( 
.A(n_2741),
.B(n_2571),
.Y(n_2801)
);

INVx2_ASAP7_75t_L g2802 ( 
.A(n_2741),
.Y(n_2802)
);

INVx2_ASAP7_75t_L g2803 ( 
.A(n_2733),
.Y(n_2803)
);

INVx1_ASAP7_75t_L g2804 ( 
.A(n_2733),
.Y(n_2804)
);

AND2x4_ASAP7_75t_L g2805 ( 
.A(n_2754),
.B(n_2567),
.Y(n_2805)
);

OAI322xp33_ASAP7_75t_L g2806 ( 
.A1(n_2720),
.A2(n_2663),
.A3(n_2580),
.B1(n_2577),
.B2(n_2656),
.C1(n_2655),
.C2(n_2651),
.Y(n_2806)
);

OAI21xp5_ASAP7_75t_L g2807 ( 
.A1(n_2670),
.A2(n_2646),
.B(n_2610),
.Y(n_2807)
);

INVx1_ASAP7_75t_SL g2808 ( 
.A(n_2692),
.Y(n_2808)
);

INVx1_ASAP7_75t_L g2809 ( 
.A(n_2669),
.Y(n_2809)
);

INVx1_ASAP7_75t_L g2810 ( 
.A(n_2664),
.Y(n_2810)
);

INVx1_ASAP7_75t_L g2811 ( 
.A(n_2666),
.Y(n_2811)
);

INVx1_ASAP7_75t_L g2812 ( 
.A(n_2667),
.Y(n_2812)
);

INVx1_ASAP7_75t_L g2813 ( 
.A(n_2678),
.Y(n_2813)
);

OR2x2_ASAP7_75t_L g2814 ( 
.A(n_2697),
.B(n_2634),
.Y(n_2814)
);

INVxp67_ASAP7_75t_SL g2815 ( 
.A(n_2679),
.Y(n_2815)
);

OR4x1_ASAP7_75t_L g2816 ( 
.A(n_2722),
.B(n_2646),
.C(n_2580),
.D(n_2650),
.Y(n_2816)
);

NAND2xp5_ASAP7_75t_L g2817 ( 
.A(n_2684),
.B(n_2689),
.Y(n_2817)
);

AOI21xp33_ASAP7_75t_L g2818 ( 
.A1(n_2743),
.A2(n_2612),
.B(n_2592),
.Y(n_2818)
);

INVx1_ASAP7_75t_L g2819 ( 
.A(n_2682),
.Y(n_2819)
);

INVx2_ASAP7_75t_L g2820 ( 
.A(n_2726),
.Y(n_2820)
);

INVx1_ASAP7_75t_L g2821 ( 
.A(n_2687),
.Y(n_2821)
);

NOR2xp33_ASAP7_75t_L g2822 ( 
.A(n_2736),
.B(n_2562),
.Y(n_2822)
);

INVx2_ASAP7_75t_L g2823 ( 
.A(n_2716),
.Y(n_2823)
);

HB1xp67_ASAP7_75t_L g2824 ( 
.A(n_2726),
.Y(n_2824)
);

INVx1_ASAP7_75t_L g2825 ( 
.A(n_2693),
.Y(n_2825)
);

INVx1_ASAP7_75t_L g2826 ( 
.A(n_2709),
.Y(n_2826)
);

OAI211xp5_ASAP7_75t_L g2827 ( 
.A1(n_2668),
.A2(n_2554),
.B(n_2661),
.C(n_2603),
.Y(n_2827)
);

OAI22xp5_ASAP7_75t_L g2828 ( 
.A1(n_2686),
.A2(n_2241),
.B1(n_2573),
.B2(n_2420),
.Y(n_2828)
);

OR2x2_ASAP7_75t_L g2829 ( 
.A(n_2680),
.B(n_2649),
.Y(n_2829)
);

OAI22xp5_ASAP7_75t_L g2830 ( 
.A1(n_2686),
.A2(n_2573),
.B1(n_2603),
.B2(n_2567),
.Y(n_2830)
);

INVx1_ASAP7_75t_L g2831 ( 
.A(n_2714),
.Y(n_2831)
);

INVx1_ASAP7_75t_L g2832 ( 
.A(n_2824),
.Y(n_2832)
);

NAND2xp33_ASAP7_75t_SL g2833 ( 
.A(n_2771),
.B(n_2731),
.Y(n_2833)
);

NOR2xp33_ASAP7_75t_L g2834 ( 
.A(n_2794),
.B(n_2731),
.Y(n_2834)
);

AND2x2_ASAP7_75t_L g2835 ( 
.A(n_2790),
.B(n_2689),
.Y(n_2835)
);

INVx1_ASAP7_75t_L g2836 ( 
.A(n_2824),
.Y(n_2836)
);

NAND2xp5_ASAP7_75t_L g2837 ( 
.A(n_2762),
.B(n_2684),
.Y(n_2837)
);

AND2x2_ASAP7_75t_L g2838 ( 
.A(n_2776),
.B(n_2691),
.Y(n_2838)
);

NOR2x1_ASAP7_75t_L g2839 ( 
.A(n_2789),
.B(n_2679),
.Y(n_2839)
);

NAND2xp5_ASAP7_75t_L g2840 ( 
.A(n_2808),
.B(n_2691),
.Y(n_2840)
);

INVx1_ASAP7_75t_L g2841 ( 
.A(n_2785),
.Y(n_2841)
);

INVxp67_ASAP7_75t_L g2842 ( 
.A(n_2785),
.Y(n_2842)
);

AND2x2_ASAP7_75t_L g2843 ( 
.A(n_2774),
.B(n_2791),
.Y(n_2843)
);

AND2x2_ASAP7_75t_L g2844 ( 
.A(n_2801),
.B(n_2685),
.Y(n_2844)
);

NAND2xp5_ASAP7_75t_L g2845 ( 
.A(n_2805),
.B(n_2685),
.Y(n_2845)
);

NAND2xp5_ASAP7_75t_L g2846 ( 
.A(n_2805),
.B(n_2681),
.Y(n_2846)
);

INVx1_ASAP7_75t_L g2847 ( 
.A(n_2768),
.Y(n_2847)
);

OR2x2_ASAP7_75t_L g2848 ( 
.A(n_2777),
.B(n_2765),
.Y(n_2848)
);

AND2x2_ASAP7_75t_L g2849 ( 
.A(n_2802),
.B(n_2670),
.Y(n_2849)
);

NAND2xp5_ASAP7_75t_L g2850 ( 
.A(n_2780),
.B(n_2681),
.Y(n_2850)
);

NAND2xp5_ASAP7_75t_L g2851 ( 
.A(n_2815),
.B(n_2742),
.Y(n_2851)
);

NAND2xp5_ASAP7_75t_L g2852 ( 
.A(n_2815),
.B(n_2742),
.Y(n_2852)
);

AND2x4_ASAP7_75t_L g2853 ( 
.A(n_2784),
.B(n_2700),
.Y(n_2853)
);

NAND2xp5_ASAP7_75t_L g2854 ( 
.A(n_2800),
.B(n_2672),
.Y(n_2854)
);

INVxp67_ASAP7_75t_SL g2855 ( 
.A(n_2757),
.Y(n_2855)
);

INVx1_ASAP7_75t_L g2856 ( 
.A(n_2756),
.Y(n_2856)
);

INVx1_ASAP7_75t_L g2857 ( 
.A(n_2769),
.Y(n_2857)
);

OR2x2_ASAP7_75t_L g2858 ( 
.A(n_2775),
.B(n_2721),
.Y(n_2858)
);

NOR2xp33_ASAP7_75t_L g2859 ( 
.A(n_2757),
.B(n_2559),
.Y(n_2859)
);

NAND2xp33_ASAP7_75t_SL g2860 ( 
.A(n_2771),
.B(n_2710),
.Y(n_2860)
);

INVx2_ASAP7_75t_L g2861 ( 
.A(n_2816),
.Y(n_2861)
);

NAND2xp5_ASAP7_75t_L g2862 ( 
.A(n_2800),
.B(n_2700),
.Y(n_2862)
);

NOR2xp33_ASAP7_75t_L g2863 ( 
.A(n_2817),
.B(n_2559),
.Y(n_2863)
);

HB1xp67_ASAP7_75t_L g2864 ( 
.A(n_2770),
.Y(n_2864)
);

INVx1_ASAP7_75t_L g2865 ( 
.A(n_2820),
.Y(n_2865)
);

INVx1_ASAP7_75t_L g2866 ( 
.A(n_2820),
.Y(n_2866)
);

OR2x2_ASAP7_75t_L g2867 ( 
.A(n_2803),
.B(n_2665),
.Y(n_2867)
);

BUFx2_ASAP7_75t_L g2868 ( 
.A(n_2807),
.Y(n_2868)
);

INVx1_ASAP7_75t_L g2869 ( 
.A(n_2787),
.Y(n_2869)
);

AND2x2_ASAP7_75t_L g2870 ( 
.A(n_2782),
.B(n_2786),
.Y(n_2870)
);

OR2x2_ASAP7_75t_L g2871 ( 
.A(n_2758),
.B(n_2728),
.Y(n_2871)
);

NAND2xp5_ASAP7_75t_L g2872 ( 
.A(n_2787),
.B(n_2702),
.Y(n_2872)
);

INVx1_ASAP7_75t_L g2873 ( 
.A(n_2795),
.Y(n_2873)
);

INVx1_ASAP7_75t_SL g2874 ( 
.A(n_2814),
.Y(n_2874)
);

INVx2_ASAP7_75t_L g2875 ( 
.A(n_2829),
.Y(n_2875)
);

INVx1_ASAP7_75t_L g2876 ( 
.A(n_2796),
.Y(n_2876)
);

AND2x2_ASAP7_75t_L g2877 ( 
.A(n_2798),
.B(n_2702),
.Y(n_2877)
);

INVx1_ASAP7_75t_L g2878 ( 
.A(n_2799),
.Y(n_2878)
);

INVx1_ASAP7_75t_L g2879 ( 
.A(n_2804),
.Y(n_2879)
);

INVx1_ASAP7_75t_L g2880 ( 
.A(n_2770),
.Y(n_2880)
);

NAND2xp5_ASAP7_75t_L g2881 ( 
.A(n_2809),
.B(n_2783),
.Y(n_2881)
);

INVx1_ASAP7_75t_L g2882 ( 
.A(n_2826),
.Y(n_2882)
);

INVx1_ASAP7_75t_L g2883 ( 
.A(n_2831),
.Y(n_2883)
);

NOR2x1_ASAP7_75t_L g2884 ( 
.A(n_2788),
.B(n_2727),
.Y(n_2884)
);

INVx1_ASAP7_75t_L g2885 ( 
.A(n_2763),
.Y(n_2885)
);

INVx2_ASAP7_75t_L g2886 ( 
.A(n_2823),
.Y(n_2886)
);

OR2x2_ASAP7_75t_L g2887 ( 
.A(n_2792),
.B(n_2732),
.Y(n_2887)
);

NAND2xp5_ASAP7_75t_L g2888 ( 
.A(n_2781),
.B(n_2671),
.Y(n_2888)
);

INVx1_ASAP7_75t_L g2889 ( 
.A(n_2764),
.Y(n_2889)
);

NOR2xp33_ASAP7_75t_L g2890 ( 
.A(n_2788),
.B(n_2649),
.Y(n_2890)
);

OAI33xp33_ASAP7_75t_L g2891 ( 
.A1(n_2760),
.A2(n_2729),
.A3(n_2723),
.B1(n_2712),
.B2(n_2747),
.B3(n_2753),
.Y(n_2891)
);

INVx1_ASAP7_75t_L g2892 ( 
.A(n_2766),
.Y(n_2892)
);

INVx1_ASAP7_75t_L g2893 ( 
.A(n_2772),
.Y(n_2893)
);

INVx1_ASAP7_75t_L g2894 ( 
.A(n_2772),
.Y(n_2894)
);

INVx1_ASAP7_75t_L g2895 ( 
.A(n_2793),
.Y(n_2895)
);

INVx1_ASAP7_75t_L g2896 ( 
.A(n_2793),
.Y(n_2896)
);

NOR2xp33_ASAP7_75t_R g2897 ( 
.A(n_2822),
.B(n_2675),
.Y(n_2897)
);

INVx1_ASAP7_75t_L g2898 ( 
.A(n_2810),
.Y(n_2898)
);

NAND2x1_ASAP7_75t_L g2899 ( 
.A(n_2830),
.B(n_2716),
.Y(n_2899)
);

AND2x2_ASAP7_75t_L g2900 ( 
.A(n_2779),
.B(n_2630),
.Y(n_2900)
);

NAND2x1_ASAP7_75t_L g2901 ( 
.A(n_2811),
.B(n_2727),
.Y(n_2901)
);

INVx2_ASAP7_75t_L g2902 ( 
.A(n_2864),
.Y(n_2902)
);

NAND2xp5_ASAP7_75t_L g2903 ( 
.A(n_2835),
.B(n_2822),
.Y(n_2903)
);

INVx2_ASAP7_75t_SL g2904 ( 
.A(n_2844),
.Y(n_2904)
);

AND2x2_ASAP7_75t_L g2905 ( 
.A(n_2843),
.B(n_2630),
.Y(n_2905)
);

INVx1_ASAP7_75t_L g2906 ( 
.A(n_2838),
.Y(n_2906)
);

AO22x1_ASAP7_75t_L g2907 ( 
.A1(n_2855),
.A2(n_2705),
.B1(n_2812),
.B2(n_2813),
.Y(n_2907)
);

NOR2xp33_ASAP7_75t_L g2908 ( 
.A(n_2842),
.B(n_2761),
.Y(n_2908)
);

INVxp67_ASAP7_75t_SL g2909 ( 
.A(n_2864),
.Y(n_2909)
);

NOR2xp33_ASAP7_75t_L g2910 ( 
.A(n_2842),
.B(n_2837),
.Y(n_2910)
);

AND2x2_ASAP7_75t_L g2911 ( 
.A(n_2849),
.B(n_2658),
.Y(n_2911)
);

AND2x2_ASAP7_75t_L g2912 ( 
.A(n_2877),
.B(n_2658),
.Y(n_2912)
);

O2A1O1Ixp33_ASAP7_75t_L g2913 ( 
.A1(n_2855),
.A2(n_2767),
.B(n_2773),
.C(n_2818),
.Y(n_2913)
);

INVx1_ASAP7_75t_L g2914 ( 
.A(n_2840),
.Y(n_2914)
);

INVx1_ASAP7_75t_L g2915 ( 
.A(n_2851),
.Y(n_2915)
);

NAND2xp5_ASAP7_75t_L g2916 ( 
.A(n_2874),
.B(n_2759),
.Y(n_2916)
);

INVx1_ASAP7_75t_L g2917 ( 
.A(n_2852),
.Y(n_2917)
);

OR2x2_ASAP7_75t_L g2918 ( 
.A(n_2848),
.B(n_2708),
.Y(n_2918)
);

OR2x2_ASAP7_75t_L g2919 ( 
.A(n_2858),
.B(n_2819),
.Y(n_2919)
);

AND2x2_ASAP7_75t_L g2920 ( 
.A(n_2875),
.B(n_2746),
.Y(n_2920)
);

NAND2xp5_ASAP7_75t_L g2921 ( 
.A(n_2834),
.B(n_2797),
.Y(n_2921)
);

INVx2_ASAP7_75t_L g2922 ( 
.A(n_2832),
.Y(n_2922)
);

NAND2xp5_ASAP7_75t_L g2923 ( 
.A(n_2834),
.B(n_2821),
.Y(n_2923)
);

INVx1_ASAP7_75t_L g2924 ( 
.A(n_2836),
.Y(n_2924)
);

INVx1_ASAP7_75t_L g2925 ( 
.A(n_2865),
.Y(n_2925)
);

NAND2x1_ASAP7_75t_L g2926 ( 
.A(n_2884),
.B(n_2579),
.Y(n_2926)
);

AND2x2_ASAP7_75t_L g2927 ( 
.A(n_2875),
.B(n_2746),
.Y(n_2927)
);

INVx1_ASAP7_75t_L g2928 ( 
.A(n_2866),
.Y(n_2928)
);

AND2x2_ASAP7_75t_L g2929 ( 
.A(n_2853),
.B(n_2825),
.Y(n_2929)
);

NAND2xp5_ASAP7_75t_L g2930 ( 
.A(n_2845),
.B(n_2734),
.Y(n_2930)
);

OR2x2_ASAP7_75t_L g2931 ( 
.A(n_2871),
.B(n_2725),
.Y(n_2931)
);

NAND2xp5_ASAP7_75t_L g2932 ( 
.A(n_2841),
.B(n_2744),
.Y(n_2932)
);

NOR2xp33_ASAP7_75t_L g2933 ( 
.A(n_2899),
.B(n_2778),
.Y(n_2933)
);

INVx1_ASAP7_75t_L g2934 ( 
.A(n_2846),
.Y(n_2934)
);

OAI211xp5_ASAP7_75t_L g2935 ( 
.A1(n_2860),
.A2(n_2827),
.B(n_2751),
.C(n_2745),
.Y(n_2935)
);

NAND2xp5_ASAP7_75t_L g2936 ( 
.A(n_2869),
.B(n_2749),
.Y(n_2936)
);

NAND2xp33_ASAP7_75t_R g2937 ( 
.A(n_2897),
.B(n_2737),
.Y(n_2937)
);

INVx1_ASAP7_75t_L g2938 ( 
.A(n_2867),
.Y(n_2938)
);

INVx1_ASAP7_75t_L g2939 ( 
.A(n_2847),
.Y(n_2939)
);

INVx2_ASAP7_75t_L g2940 ( 
.A(n_2853),
.Y(n_2940)
);

INVx2_ASAP7_75t_L g2941 ( 
.A(n_2880),
.Y(n_2941)
);

NOR2xp33_ASAP7_75t_L g2942 ( 
.A(n_2872),
.B(n_2827),
.Y(n_2942)
);

AND2x2_ASAP7_75t_L g2943 ( 
.A(n_2900),
.B(n_2579),
.Y(n_2943)
);

NOR2x1p5_ASAP7_75t_L g2944 ( 
.A(n_2901),
.B(n_2550),
.Y(n_2944)
);

NOR2xp33_ASAP7_75t_L g2945 ( 
.A(n_2862),
.B(n_2806),
.Y(n_2945)
);

INVx1_ASAP7_75t_L g2946 ( 
.A(n_2870),
.Y(n_2946)
);

AND2x2_ASAP7_75t_L g2947 ( 
.A(n_2839),
.B(n_2579),
.Y(n_2947)
);

NOR2xp33_ASAP7_75t_L g2948 ( 
.A(n_2891),
.B(n_2890),
.Y(n_2948)
);

INVx1_ASAP7_75t_L g2949 ( 
.A(n_2854),
.Y(n_2949)
);

INVxp33_ASAP7_75t_L g2950 ( 
.A(n_2897),
.Y(n_2950)
);

INVx1_ASAP7_75t_L g2951 ( 
.A(n_2886),
.Y(n_2951)
);

INVx1_ASAP7_75t_L g2952 ( 
.A(n_2886),
.Y(n_2952)
);

OR4x1_ASAP7_75t_L g2953 ( 
.A(n_2895),
.B(n_2497),
.C(n_2509),
.D(n_2492),
.Y(n_2953)
);

INVx1_ASAP7_75t_L g2954 ( 
.A(n_2888),
.Y(n_2954)
);

INVxp67_ASAP7_75t_SL g2955 ( 
.A(n_2890),
.Y(n_2955)
);

INVx1_ASAP7_75t_L g2956 ( 
.A(n_2887),
.Y(n_2956)
);

AND2x2_ASAP7_75t_L g2957 ( 
.A(n_2868),
.B(n_2856),
.Y(n_2957)
);

XNOR2xp5_ASAP7_75t_L g2958 ( 
.A(n_2881),
.B(n_2828),
.Y(n_2958)
);

NAND3xp33_ASAP7_75t_L g2959 ( 
.A(n_2860),
.B(n_2833),
.C(n_2896),
.Y(n_2959)
);

HB1xp67_ASAP7_75t_L g2960 ( 
.A(n_2850),
.Y(n_2960)
);

INVx1_ASAP7_75t_L g2961 ( 
.A(n_2857),
.Y(n_2961)
);

NOR3xp33_ASAP7_75t_L g2962 ( 
.A(n_2959),
.B(n_2833),
.C(n_2893),
.Y(n_2962)
);

INVx2_ASAP7_75t_L g2963 ( 
.A(n_2904),
.Y(n_2963)
);

AND2x2_ASAP7_75t_L g2964 ( 
.A(n_2905),
.B(n_2863),
.Y(n_2964)
);

NAND2xp33_ASAP7_75t_SL g2965 ( 
.A(n_2950),
.B(n_2861),
.Y(n_2965)
);

INVx2_ASAP7_75t_SL g2966 ( 
.A(n_2912),
.Y(n_2966)
);

INVx1_ASAP7_75t_L g2967 ( 
.A(n_2909),
.Y(n_2967)
);

O2A1O1Ixp33_ASAP7_75t_L g2968 ( 
.A1(n_2913),
.A2(n_2861),
.B(n_2891),
.C(n_2894),
.Y(n_2968)
);

NAND4xp25_ASAP7_75t_L g2969 ( 
.A(n_2933),
.B(n_2863),
.C(n_2859),
.D(n_2882),
.Y(n_2969)
);

NAND4xp25_ASAP7_75t_L g2970 ( 
.A(n_2945),
.B(n_2859),
.C(n_2883),
.D(n_2876),
.Y(n_2970)
);

NOR4xp25_ASAP7_75t_L g2971 ( 
.A(n_2935),
.B(n_2889),
.C(n_2892),
.D(n_2885),
.Y(n_2971)
);

INVx1_ASAP7_75t_L g2972 ( 
.A(n_2902),
.Y(n_2972)
);

OAI221xp5_ASAP7_75t_L g2973 ( 
.A1(n_2933),
.A2(n_2898),
.B1(n_2879),
.B2(n_2878),
.C(n_2873),
.Y(n_2973)
);

O2A1O1Ixp33_ASAP7_75t_L g2974 ( 
.A1(n_2902),
.A2(n_2550),
.B(n_2612),
.C(n_2592),
.Y(n_2974)
);

AND2x2_ASAP7_75t_L g2975 ( 
.A(n_2904),
.B(n_2579),
.Y(n_2975)
);

NAND3xp33_ASAP7_75t_L g2976 ( 
.A(n_2948),
.B(n_2615),
.C(n_2613),
.Y(n_2976)
);

NOR3x1_ASAP7_75t_L g2977 ( 
.A(n_2926),
.B(n_2516),
.C(n_2515),
.Y(n_2977)
);

INVx1_ASAP7_75t_L g2978 ( 
.A(n_2929),
.Y(n_2978)
);

OR2x2_ASAP7_75t_L g2979 ( 
.A(n_2940),
.B(n_2517),
.Y(n_2979)
);

INVx3_ASAP7_75t_L g2980 ( 
.A(n_2940),
.Y(n_2980)
);

AOI211x1_ASAP7_75t_L g2981 ( 
.A1(n_2907),
.A2(n_2542),
.B(n_2518),
.C(n_2403),
.Y(n_2981)
);

INVx1_ASAP7_75t_L g2982 ( 
.A(n_2929),
.Y(n_2982)
);

INVx2_ASAP7_75t_L g2983 ( 
.A(n_2918),
.Y(n_2983)
);

INVx1_ASAP7_75t_L g2984 ( 
.A(n_2957),
.Y(n_2984)
);

NOR2xp33_ASAP7_75t_L g2985 ( 
.A(n_2950),
.B(n_2617),
.Y(n_2985)
);

INVx1_ASAP7_75t_L g2986 ( 
.A(n_2957),
.Y(n_2986)
);

A2O1A1Ixp33_ASAP7_75t_SL g2987 ( 
.A1(n_2948),
.A2(n_2636),
.B(n_2637),
.C(n_2617),
.Y(n_2987)
);

INVx1_ASAP7_75t_L g2988 ( 
.A(n_2931),
.Y(n_2988)
);

NAND3xp33_ASAP7_75t_L g2989 ( 
.A(n_2942),
.B(n_2637),
.C(n_2636),
.Y(n_2989)
);

INVx2_ASAP7_75t_SL g2990 ( 
.A(n_2944),
.Y(n_2990)
);

INVx1_ASAP7_75t_L g2991 ( 
.A(n_2919),
.Y(n_2991)
);

INVx1_ASAP7_75t_L g2992 ( 
.A(n_2951),
.Y(n_2992)
);

AND3x2_ASAP7_75t_L g2993 ( 
.A(n_2947),
.B(n_2638),
.C(n_2383),
.Y(n_2993)
);

XNOR2x2_ASAP7_75t_L g2994 ( 
.A(n_2945),
.B(n_2638),
.Y(n_2994)
);

AOI21xp5_ASAP7_75t_L g2995 ( 
.A1(n_2921),
.A2(n_2496),
.B(n_2494),
.Y(n_2995)
);

NOR3xp33_ASAP7_75t_L g2996 ( 
.A(n_2916),
.B(n_2507),
.C(n_2503),
.Y(n_2996)
);

NOR2xp33_ASAP7_75t_L g2997 ( 
.A(n_2955),
.B(n_2396),
.Y(n_2997)
);

NAND2xp5_ASAP7_75t_L g2998 ( 
.A(n_2911),
.B(n_2403),
.Y(n_2998)
);

OAI21xp33_ASAP7_75t_SL g2999 ( 
.A1(n_2942),
.A2(n_2413),
.B(n_2406),
.Y(n_2999)
);

AOI21xp33_ASAP7_75t_L g3000 ( 
.A1(n_2937),
.A2(n_2952),
.B(n_2947),
.Y(n_3000)
);

NOR2xp33_ASAP7_75t_L g3001 ( 
.A(n_2954),
.B(n_2920),
.Y(n_3001)
);

NAND4xp25_ASAP7_75t_L g3002 ( 
.A(n_2910),
.B(n_2507),
.C(n_2526),
.D(n_2514),
.Y(n_3002)
);

INVx1_ASAP7_75t_L g3003 ( 
.A(n_2920),
.Y(n_3003)
);

NAND4xp25_ASAP7_75t_L g3004 ( 
.A(n_2910),
.B(n_2514),
.C(n_2527),
.D(n_2526),
.Y(n_3004)
);

AND2x2_ASAP7_75t_L g3005 ( 
.A(n_2943),
.B(n_2349),
.Y(n_3005)
);

NAND2xp5_ASAP7_75t_L g3006 ( 
.A(n_2927),
.B(n_2406),
.Y(n_3006)
);

AOI21xp5_ASAP7_75t_L g3007 ( 
.A1(n_2903),
.A2(n_2535),
.B(n_2527),
.Y(n_3007)
);

NOR2xp33_ASAP7_75t_L g3008 ( 
.A(n_2927),
.B(n_2413),
.Y(n_3008)
);

AND2x2_ASAP7_75t_L g3009 ( 
.A(n_2946),
.B(n_2349),
.Y(n_3009)
);

NAND4xp25_ASAP7_75t_L g3010 ( 
.A(n_2908),
.B(n_2535),
.C(n_2539),
.D(n_2536),
.Y(n_3010)
);

NOR2x1_ASAP7_75t_L g3011 ( 
.A(n_2938),
.B(n_1034),
.Y(n_3011)
);

NAND2xp33_ASAP7_75t_SL g3012 ( 
.A(n_2978),
.B(n_2941),
.Y(n_3012)
);

AOI221xp5_ASAP7_75t_L g3013 ( 
.A1(n_2987),
.A2(n_2960),
.B1(n_2953),
.B2(n_2908),
.C(n_2941),
.Y(n_3013)
);

OAI22xp5_ASAP7_75t_L g3014 ( 
.A1(n_2983),
.A2(n_2923),
.B1(n_2939),
.B2(n_2936),
.Y(n_3014)
);

NAND3xp33_ASAP7_75t_L g3015 ( 
.A(n_2962),
.B(n_2937),
.C(n_2958),
.Y(n_3015)
);

NOR3xp33_ASAP7_75t_L g3016 ( 
.A(n_3000),
.B(n_2917),
.C(n_2915),
.Y(n_3016)
);

AOI22xp5_ASAP7_75t_L g3017 ( 
.A1(n_3001),
.A2(n_2914),
.B1(n_2928),
.B2(n_2925),
.Y(n_3017)
);

AOI21xp5_ASAP7_75t_L g3018 ( 
.A1(n_2968),
.A2(n_2930),
.B(n_2932),
.Y(n_3018)
);

NAND4xp75_ASAP7_75t_L g3019 ( 
.A(n_2977),
.B(n_2906),
.C(n_2956),
.D(n_2934),
.Y(n_3019)
);

A2O1A1Ixp33_ASAP7_75t_L g3020 ( 
.A1(n_2976),
.A2(n_2922),
.B(n_2924),
.C(n_2961),
.Y(n_3020)
);

AOI211xp5_ASAP7_75t_SL g3021 ( 
.A1(n_2973),
.A2(n_2949),
.B(n_2922),
.C(n_2953),
.Y(n_3021)
);

NAND4xp25_ASAP7_75t_L g3022 ( 
.A(n_2969),
.B(n_2536),
.C(n_2539),
.D(n_2365),
.Y(n_3022)
);

AND2x2_ASAP7_75t_L g3023 ( 
.A(n_3005),
.B(n_2422),
.Y(n_3023)
);

AOI322xp5_ASAP7_75t_L g3024 ( 
.A1(n_2996),
.A2(n_2421),
.A3(n_2375),
.B1(n_2397),
.B2(n_2391),
.C1(n_2384),
.C2(n_2185),
.Y(n_3024)
);

INVx1_ASAP7_75t_L g3025 ( 
.A(n_2980),
.Y(n_3025)
);

NOR4xp25_ASAP7_75t_L g3026 ( 
.A(n_2976),
.B(n_2384),
.C(n_2391),
.D(n_2375),
.Y(n_3026)
);

AOI211xp5_ASAP7_75t_L g3027 ( 
.A1(n_2971),
.A2(n_2383),
.B(n_2365),
.C(n_2397),
.Y(n_3027)
);

NOR2x1_ASAP7_75t_L g3028 ( 
.A(n_2982),
.B(n_2253),
.Y(n_3028)
);

AND2x2_ASAP7_75t_L g3029 ( 
.A(n_3009),
.B(n_2422),
.Y(n_3029)
);

AOI22xp33_ASAP7_75t_L g3030 ( 
.A1(n_2994),
.A2(n_2203),
.B1(n_2228),
.B2(n_2216),
.Y(n_3030)
);

OAI21xp5_ASAP7_75t_L g3031 ( 
.A1(n_3007),
.A2(n_2414),
.B(n_2383),
.Y(n_3031)
);

AOI221x1_ASAP7_75t_SL g3032 ( 
.A1(n_2970),
.A2(n_2383),
.B1(n_2352),
.B2(n_2270),
.C(n_2275),
.Y(n_3032)
);

AOI221xp5_ASAP7_75t_L g3033 ( 
.A1(n_2989),
.A2(n_2414),
.B1(n_2203),
.B2(n_2247),
.C(n_2216),
.Y(n_3033)
);

INVx1_ASAP7_75t_L g3034 ( 
.A(n_2980),
.Y(n_3034)
);

NAND4xp25_ASAP7_75t_L g3035 ( 
.A(n_2988),
.B(n_2352),
.C(n_2139),
.D(n_979),
.Y(n_3035)
);

NAND2xp33_ASAP7_75t_L g3036 ( 
.A(n_2984),
.B(n_2423),
.Y(n_3036)
);

NOR2xp33_ASAP7_75t_R g3037 ( 
.A(n_2965),
.B(n_2372),
.Y(n_3037)
);

NAND2xp5_ASAP7_75t_L g3038 ( 
.A(n_2966),
.B(n_2372),
.Y(n_3038)
);

AND4x2_ASAP7_75t_L g3039 ( 
.A(n_3011),
.B(n_2287),
.C(n_2334),
.D(n_2322),
.Y(n_3039)
);

OAI21xp5_ASAP7_75t_SL g3040 ( 
.A1(n_2986),
.A2(n_2139),
.B(n_2266),
.Y(n_3040)
);

A2O1A1Ixp33_ASAP7_75t_L g3041 ( 
.A1(n_2989),
.A2(n_2228),
.B(n_2245),
.C(n_2247),
.Y(n_3041)
);

AOI221xp5_ASAP7_75t_L g3042 ( 
.A1(n_2995),
.A2(n_2245),
.B1(n_2256),
.B2(n_2270),
.C(n_2275),
.Y(n_3042)
);

OAI31xp33_ASAP7_75t_L g3043 ( 
.A1(n_3010),
.A2(n_2256),
.A3(n_2423),
.B(n_2401),
.Y(n_3043)
);

O2A1O1Ixp33_ASAP7_75t_L g3044 ( 
.A1(n_2990),
.A2(n_2401),
.B(n_2254),
.C(n_2107),
.Y(n_3044)
);

INVx1_ASAP7_75t_L g3045 ( 
.A(n_3003),
.Y(n_3045)
);

OAI211xp5_ASAP7_75t_L g3046 ( 
.A1(n_2972),
.A2(n_2334),
.B(n_2371),
.C(n_2376),
.Y(n_3046)
);

INVxp67_ASAP7_75t_L g3047 ( 
.A(n_2975),
.Y(n_3047)
);

AOI211xp5_ASAP7_75t_L g3048 ( 
.A1(n_2970),
.A2(n_2377),
.B(n_2376),
.C(n_2371),
.Y(n_3048)
);

OAI221xp5_ASAP7_75t_L g3049 ( 
.A1(n_2999),
.A2(n_2107),
.B1(n_2290),
.B2(n_2121),
.C(n_2377),
.Y(n_3049)
);

INVx1_ASAP7_75t_L g3050 ( 
.A(n_2963),
.Y(n_3050)
);

AOI211xp5_ASAP7_75t_L g3051 ( 
.A1(n_2967),
.A2(n_2329),
.B(n_2328),
.C(n_2325),
.Y(n_3051)
);

OAI22xp5_ASAP7_75t_L g3052 ( 
.A1(n_3017),
.A2(n_2991),
.B1(n_2979),
.B2(n_2992),
.Y(n_3052)
);

INVx2_ASAP7_75t_L g3053 ( 
.A(n_3023),
.Y(n_3053)
);

OAI311xp33_ASAP7_75t_L g3054 ( 
.A1(n_3013),
.A2(n_3010),
.A3(n_3004),
.B1(n_3002),
.C1(n_3006),
.Y(n_3054)
);

INVx2_ASAP7_75t_L g3055 ( 
.A(n_3029),
.Y(n_3055)
);

AOI221xp5_ASAP7_75t_L g3056 ( 
.A1(n_3013),
.A2(n_2974),
.B1(n_2985),
.B2(n_2981),
.C(n_3008),
.Y(n_3056)
);

OAI211xp5_ASAP7_75t_SL g3057 ( 
.A1(n_3021),
.A2(n_2998),
.B(n_2997),
.C(n_2964),
.Y(n_3057)
);

INVxp33_ASAP7_75t_SL g3058 ( 
.A(n_3014),
.Y(n_3058)
);

AOI22xp5_ASAP7_75t_L g3059 ( 
.A1(n_3015),
.A2(n_3025),
.B1(n_3034),
.B2(n_3012),
.Y(n_3059)
);

AOI221xp5_ASAP7_75t_L g3060 ( 
.A1(n_3026),
.A2(n_2993),
.B1(n_2121),
.B2(n_2329),
.C(n_2328),
.Y(n_3060)
);

AOI321xp33_ASAP7_75t_L g3061 ( 
.A1(n_3027),
.A2(n_2198),
.A3(n_2195),
.B1(n_2051),
.B2(n_979),
.C(n_984),
.Y(n_3061)
);

AOI22xp33_ASAP7_75t_L g3062 ( 
.A1(n_3042),
.A2(n_2287),
.B1(n_2195),
.B2(n_2198),
.Y(n_3062)
);

AOI322xp5_ASAP7_75t_L g3063 ( 
.A1(n_3030),
.A2(n_2047),
.A3(n_2195),
.B1(n_2198),
.B2(n_1975),
.C1(n_1995),
.C2(n_1997),
.Y(n_3063)
);

CKINVDCx14_ASAP7_75t_R g3064 ( 
.A(n_3037),
.Y(n_3064)
);

OAI211xp5_ASAP7_75t_SL g3065 ( 
.A1(n_3018),
.A2(n_2287),
.B(n_2095),
.C(n_2063),
.Y(n_3065)
);

NAND4xp25_ASAP7_75t_SL g3066 ( 
.A(n_3048),
.B(n_2325),
.C(n_2323),
.D(n_2322),
.Y(n_3066)
);

AOI221xp5_ASAP7_75t_L g3067 ( 
.A1(n_3032),
.A2(n_2323),
.B1(n_2020),
.B2(n_2081),
.C(n_2075),
.Y(n_3067)
);

A2O1A1Ixp33_ASAP7_75t_L g3068 ( 
.A1(n_3031),
.A2(n_2360),
.B(n_984),
.C(n_1950),
.Y(n_3068)
);

OAI21xp33_ASAP7_75t_L g3069 ( 
.A1(n_3035),
.A2(n_2223),
.B(n_2092),
.Y(n_3069)
);

OAI211xp5_ASAP7_75t_L g3070 ( 
.A1(n_3020),
.A2(n_3050),
.B(n_3045),
.C(n_3016),
.Y(n_3070)
);

NAND3xp33_ASAP7_75t_SL g3071 ( 
.A(n_3047),
.B(n_3024),
.C(n_3043),
.Y(n_3071)
);

OAI221xp5_ASAP7_75t_L g3072 ( 
.A1(n_3022),
.A2(n_1968),
.B1(n_1963),
.B2(n_1954),
.C(n_2028),
.Y(n_3072)
);

INVx1_ASAP7_75t_L g3073 ( 
.A(n_3038),
.Y(n_3073)
);

HB1xp67_ASAP7_75t_L g3074 ( 
.A(n_3028),
.Y(n_3074)
);

AND3x1_ASAP7_75t_L g3075 ( 
.A(n_3051),
.B(n_2223),
.C(n_1897),
.Y(n_3075)
);

NOR2xp33_ASAP7_75t_R g3076 ( 
.A(n_3036),
.B(n_1764),
.Y(n_3076)
);

AOI22xp5_ASAP7_75t_L g3077 ( 
.A1(n_3033),
.A2(n_3019),
.B1(n_3049),
.B2(n_3040),
.Y(n_3077)
);

AOI22xp5_ASAP7_75t_L g3078 ( 
.A1(n_3049),
.A2(n_3046),
.B1(n_3041),
.B2(n_3039),
.Y(n_3078)
);

AOI221xp5_ASAP7_75t_L g3079 ( 
.A1(n_3044),
.A2(n_1995),
.B1(n_2061),
.B2(n_2075),
.C(n_2046),
.Y(n_3079)
);

AOI221xp5_ASAP7_75t_L g3080 ( 
.A1(n_3013),
.A2(n_2081),
.B1(n_2061),
.B2(n_2046),
.C(n_1997),
.Y(n_3080)
);

AOI211xp5_ASAP7_75t_L g3081 ( 
.A1(n_3013),
.A2(n_2128),
.B(n_1764),
.C(n_1875),
.Y(n_3081)
);

OAI211xp5_ASAP7_75t_SL g3082 ( 
.A1(n_3013),
.A2(n_2089),
.B(n_2128),
.C(n_1836),
.Y(n_3082)
);

OAI222xp33_ASAP7_75t_L g3083 ( 
.A1(n_3028),
.A2(n_2020),
.B1(n_1950),
.B2(n_1964),
.C1(n_1975),
.C2(n_2073),
.Y(n_3083)
);

NAND2xp5_ASAP7_75t_L g3084 ( 
.A(n_3025),
.B(n_1964),
.Y(n_3084)
);

INVx1_ASAP7_75t_L g3085 ( 
.A(n_3025),
.Y(n_3085)
);

HB1xp67_ASAP7_75t_L g3086 ( 
.A(n_3037),
.Y(n_3086)
);

AOI211xp5_ASAP7_75t_L g3087 ( 
.A1(n_3054),
.A2(n_3056),
.B(n_3057),
.C(n_3052),
.Y(n_3087)
);

AO22x2_ASAP7_75t_L g3088 ( 
.A1(n_3070),
.A2(n_2035),
.B1(n_2073),
.B2(n_2044),
.Y(n_3088)
);

NOR2xp33_ASAP7_75t_L g3089 ( 
.A(n_3074),
.B(n_1954),
.Y(n_3089)
);

NAND3x1_ASAP7_75t_SL g3090 ( 
.A(n_3058),
.B(n_1942),
.C(n_1932),
.Y(n_3090)
);

INVx1_ASAP7_75t_L g3091 ( 
.A(n_3086),
.Y(n_3091)
);

OAI32xp33_ASAP7_75t_L g3092 ( 
.A1(n_3053),
.A2(n_1897),
.A3(n_2035),
.B1(n_2044),
.B2(n_1943),
.Y(n_3092)
);

INVx1_ASAP7_75t_L g3093 ( 
.A(n_3055),
.Y(n_3093)
);

NOR2xp33_ASAP7_75t_L g3094 ( 
.A(n_3064),
.B(n_1954),
.Y(n_3094)
);

INVx1_ASAP7_75t_L g3095 ( 
.A(n_3059),
.Y(n_3095)
);

NAND3x1_ASAP7_75t_SL g3096 ( 
.A(n_3060),
.B(n_1932),
.C(n_1949),
.Y(n_3096)
);

XNOR2xp5_ASAP7_75t_L g3097 ( 
.A(n_3078),
.B(n_2085),
.Y(n_3097)
);

AOI22xp5_ASAP7_75t_L g3098 ( 
.A1(n_3071),
.A2(n_1968),
.B1(n_1963),
.B2(n_1764),
.Y(n_3098)
);

OAI22xp5_ASAP7_75t_L g3099 ( 
.A1(n_3077),
.A2(n_1875),
.B1(n_1764),
.B2(n_1963),
.Y(n_3099)
);

INVx1_ASAP7_75t_L g3100 ( 
.A(n_3085),
.Y(n_3100)
);

CKINVDCx5p33_ASAP7_75t_R g3101 ( 
.A(n_3073),
.Y(n_3101)
);

AOI221xp5_ASAP7_75t_L g3102 ( 
.A1(n_3082),
.A2(n_1789),
.B1(n_1791),
.B2(n_1780),
.C(n_1875),
.Y(n_3102)
);

AND2x2_ASAP7_75t_L g3103 ( 
.A(n_3075),
.B(n_1774),
.Y(n_3103)
);

AOI22xp33_ASAP7_75t_L g3104 ( 
.A1(n_3072),
.A2(n_1968),
.B1(n_2111),
.B2(n_2033),
.Y(n_3104)
);

NOR3xp33_ASAP7_75t_L g3105 ( 
.A(n_3081),
.B(n_1966),
.C(n_2076),
.Y(n_3105)
);

AOI221xp5_ASAP7_75t_L g3106 ( 
.A1(n_3084),
.A2(n_1789),
.B1(n_1791),
.B2(n_1780),
.C(n_1875),
.Y(n_3106)
);

HB1xp67_ASAP7_75t_L g3107 ( 
.A(n_3076),
.Y(n_3107)
);

NOR2xp33_ASAP7_75t_L g3108 ( 
.A(n_3068),
.B(n_1966),
.Y(n_3108)
);

INVx1_ASAP7_75t_SL g3109 ( 
.A(n_3084),
.Y(n_3109)
);

NOR2x1p5_ASAP7_75t_L g3110 ( 
.A(n_3061),
.B(n_1764),
.Y(n_3110)
);

NAND2xp5_ASAP7_75t_L g3111 ( 
.A(n_3069),
.B(n_2076),
.Y(n_3111)
);

AOI22xp5_ASAP7_75t_L g3112 ( 
.A1(n_3065),
.A2(n_1875),
.B1(n_1774),
.B2(n_2085),
.Y(n_3112)
);

NAND3xp33_ASAP7_75t_SL g3113 ( 
.A(n_3087),
.B(n_3080),
.C(n_3063),
.Y(n_3113)
);

INVx1_ASAP7_75t_L g3114 ( 
.A(n_3088),
.Y(n_3114)
);

CKINVDCx5p33_ASAP7_75t_R g3115 ( 
.A(n_3101),
.Y(n_3115)
);

AND2x4_ASAP7_75t_L g3116 ( 
.A(n_3093),
.B(n_3062),
.Y(n_3116)
);

NAND3xp33_ASAP7_75t_SL g3117 ( 
.A(n_3109),
.B(n_3067),
.C(n_3079),
.Y(n_3117)
);

NOR2x1_ASAP7_75t_L g3118 ( 
.A(n_3095),
.B(n_3066),
.Y(n_3118)
);

AND2x2_ASAP7_75t_L g3119 ( 
.A(n_3110),
.B(n_3103),
.Y(n_3119)
);

NOR3xp33_ASAP7_75t_SL g3120 ( 
.A(n_3091),
.B(n_3083),
.C(n_1221),
.Y(n_3120)
);

OR2x2_ASAP7_75t_L g3121 ( 
.A(n_3100),
.B(n_1946),
.Y(n_3121)
);

NOR4xp75_ASAP7_75t_SL g3122 ( 
.A(n_3099),
.B(n_1821),
.C(n_2082),
.D(n_1847),
.Y(n_3122)
);

AOI21xp5_ASAP7_75t_L g3123 ( 
.A1(n_3107),
.A2(n_1948),
.B(n_2111),
.Y(n_3123)
);

NOR2x1_ASAP7_75t_L g3124 ( 
.A(n_3097),
.B(n_1046),
.Y(n_3124)
);

NOR2x1_ASAP7_75t_L g3125 ( 
.A(n_3094),
.B(n_1124),
.Y(n_3125)
);

NAND4xp75_ASAP7_75t_L g3126 ( 
.A(n_3098),
.B(n_1011),
.C(n_1019),
.D(n_2111),
.Y(n_3126)
);

NAND3xp33_ASAP7_75t_SL g3127 ( 
.A(n_3089),
.B(n_2047),
.C(n_1796),
.Y(n_3127)
);

NAND4xp75_ASAP7_75t_L g3128 ( 
.A(n_3112),
.B(n_1991),
.C(n_2001),
.D(n_2021),
.Y(n_3128)
);

NAND4xp75_ASAP7_75t_L g3129 ( 
.A(n_3108),
.B(n_1991),
.C(n_2001),
.D(n_2021),
.Y(n_3129)
);

NAND4xp75_ASAP7_75t_L g3130 ( 
.A(n_3102),
.B(n_1991),
.C(n_2001),
.D(n_2021),
.Y(n_3130)
);

NOR3xp33_ASAP7_75t_L g3131 ( 
.A(n_3096),
.B(n_2034),
.C(n_1096),
.Y(n_3131)
);

OAI211xp5_ASAP7_75t_L g3132 ( 
.A1(n_3111),
.A2(n_1781),
.B(n_1779),
.C(n_1805),
.Y(n_3132)
);

NAND2xp33_ASAP7_75t_L g3133 ( 
.A(n_3115),
.B(n_3118),
.Y(n_3133)
);

NAND2x1p5_ASAP7_75t_L g3134 ( 
.A(n_3116),
.B(n_3090),
.Y(n_3134)
);

INVx1_ASAP7_75t_L g3135 ( 
.A(n_3114),
.Y(n_3135)
);

INVx1_ASAP7_75t_SL g3136 ( 
.A(n_3116),
.Y(n_3136)
);

CKINVDCx5p33_ASAP7_75t_R g3137 ( 
.A(n_3113),
.Y(n_3137)
);

BUFx2_ASAP7_75t_L g3138 ( 
.A(n_3124),
.Y(n_3138)
);

NAND2x1p5_ASAP7_75t_L g3139 ( 
.A(n_3119),
.B(n_3088),
.Y(n_3139)
);

NAND2xp5_ASAP7_75t_L g3140 ( 
.A(n_3125),
.B(n_3105),
.Y(n_3140)
);

XNOR2xp5_ASAP7_75t_L g3141 ( 
.A(n_3117),
.B(n_3104),
.Y(n_3141)
);

BUFx2_ASAP7_75t_L g3142 ( 
.A(n_3121),
.Y(n_3142)
);

CKINVDCx16_ASAP7_75t_R g3143 ( 
.A(n_3127),
.Y(n_3143)
);

BUFx2_ASAP7_75t_L g3144 ( 
.A(n_3120),
.Y(n_3144)
);

INVx2_ASAP7_75t_L g3145 ( 
.A(n_3129),
.Y(n_3145)
);

CKINVDCx6p67_ASAP7_75t_R g3146 ( 
.A(n_3122),
.Y(n_3146)
);

CKINVDCx5p33_ASAP7_75t_R g3147 ( 
.A(n_3123),
.Y(n_3147)
);

NOR2x1_ASAP7_75t_L g3148 ( 
.A(n_3130),
.B(n_3092),
.Y(n_3148)
);

NOR4xp25_ASAP7_75t_SL g3149 ( 
.A(n_3131),
.B(n_3106),
.C(n_3126),
.D(n_3128),
.Y(n_3149)
);

NOR2xp67_ASAP7_75t_L g3150 ( 
.A(n_3132),
.B(n_1116),
.Y(n_3150)
);

NOR3xp33_ASAP7_75t_SL g3151 ( 
.A(n_3115),
.B(n_1821),
.C(n_1116),
.Y(n_3151)
);

NOR2xp33_ASAP7_75t_L g3152 ( 
.A(n_3136),
.B(n_1796),
.Y(n_3152)
);

AND3x1_ASAP7_75t_L g3153 ( 
.A(n_3145),
.B(n_1805),
.C(n_1779),
.Y(n_3153)
);

XNOR2x2_ASAP7_75t_L g3154 ( 
.A(n_3141),
.B(n_1781),
.Y(n_3154)
);

INVx1_ASAP7_75t_L g3155 ( 
.A(n_3134),
.Y(n_3155)
);

NAND3xp33_ASAP7_75t_L g3156 ( 
.A(n_3133),
.B(n_1090),
.C(n_1100),
.Y(n_3156)
);

AO22x2_ASAP7_75t_L g3157 ( 
.A1(n_3135),
.A2(n_3146),
.B1(n_3139),
.B2(n_3140),
.Y(n_3157)
);

AOI22x1_ASAP7_75t_L g3158 ( 
.A1(n_3137),
.A2(n_1854),
.B1(n_1847),
.B2(n_1815),
.Y(n_3158)
);

OAI22x1_ASAP7_75t_L g3159 ( 
.A1(n_3142),
.A2(n_1845),
.B1(n_1843),
.B2(n_1854),
.Y(n_3159)
);

OA22x2_ASAP7_75t_L g3160 ( 
.A1(n_3147),
.A2(n_1843),
.B1(n_1845),
.B2(n_1815),
.Y(n_3160)
);

INVx2_ASAP7_75t_L g3161 ( 
.A(n_3138),
.Y(n_3161)
);

OAI22xp5_ASAP7_75t_L g3162 ( 
.A1(n_3150),
.A2(n_3148),
.B1(n_3143),
.B2(n_3149),
.Y(n_3162)
);

NAND3xp33_ASAP7_75t_L g3163 ( 
.A(n_3144),
.B(n_1099),
.C(n_1100),
.Y(n_3163)
);

INVx1_ASAP7_75t_L g3164 ( 
.A(n_3150),
.Y(n_3164)
);

AOI22xp5_ASAP7_75t_L g3165 ( 
.A1(n_3151),
.A2(n_3149),
.B1(n_2100),
.B2(n_1117),
.Y(n_3165)
);

INVx1_ASAP7_75t_L g3166 ( 
.A(n_3136),
.Y(n_3166)
);

AO21x1_ASAP7_75t_L g3167 ( 
.A1(n_3134),
.A2(n_1331),
.B(n_1882),
.Y(n_3167)
);

INVx2_ASAP7_75t_L g3168 ( 
.A(n_3134),
.Y(n_3168)
);

HB1xp67_ASAP7_75t_L g3169 ( 
.A(n_3166),
.Y(n_3169)
);

INVx1_ASAP7_75t_L g3170 ( 
.A(n_3157),
.Y(n_3170)
);

HB1xp67_ASAP7_75t_L g3171 ( 
.A(n_3168),
.Y(n_3171)
);

INVx1_ASAP7_75t_L g3172 ( 
.A(n_3157),
.Y(n_3172)
);

AOI21xp33_ASAP7_75t_L g3173 ( 
.A1(n_3161),
.A2(n_2100),
.B(n_1925),
.Y(n_3173)
);

INVx1_ASAP7_75t_L g3174 ( 
.A(n_3154),
.Y(n_3174)
);

XOR2xp5_ASAP7_75t_L g3175 ( 
.A(n_3162),
.B(n_1083),
.Y(n_3175)
);

AND2x4_ASAP7_75t_L g3176 ( 
.A(n_3155),
.B(n_1084),
.Y(n_3176)
);

INVx2_ASAP7_75t_L g3177 ( 
.A(n_3153),
.Y(n_3177)
);

OAI22x1_ASAP7_75t_L g3178 ( 
.A1(n_3164),
.A2(n_1405),
.B1(n_1304),
.B2(n_1882),
.Y(n_3178)
);

OAI22xp5_ASAP7_75t_L g3179 ( 
.A1(n_3156),
.A2(n_1921),
.B1(n_1916),
.B2(n_1922),
.Y(n_3179)
);

NAND2xp5_ASAP7_75t_L g3180 ( 
.A(n_3152),
.B(n_2103),
.Y(n_3180)
);

XOR2xp5_ASAP7_75t_L g3181 ( 
.A(n_3165),
.B(n_1106),
.Y(n_3181)
);

OAI21xp5_ASAP7_75t_L g3182 ( 
.A1(n_3163),
.A2(n_2034),
.B(n_1382),
.Y(n_3182)
);

CKINVDCx20_ASAP7_75t_R g3183 ( 
.A(n_3167),
.Y(n_3183)
);

HB1xp67_ASAP7_75t_L g3184 ( 
.A(n_3160),
.Y(n_3184)
);

INVx3_ASAP7_75t_L g3185 ( 
.A(n_3170),
.Y(n_3185)
);

INVx1_ASAP7_75t_L g3186 ( 
.A(n_3171),
.Y(n_3186)
);

INVx1_ASAP7_75t_L g3187 ( 
.A(n_3169),
.Y(n_3187)
);

INVx1_ASAP7_75t_L g3188 ( 
.A(n_3172),
.Y(n_3188)
);

INVx1_ASAP7_75t_L g3189 ( 
.A(n_3174),
.Y(n_3189)
);

INVx1_ASAP7_75t_L g3190 ( 
.A(n_3184),
.Y(n_3190)
);

INVx2_ASAP7_75t_L g3191 ( 
.A(n_3183),
.Y(n_3191)
);

INVx2_ASAP7_75t_L g3192 ( 
.A(n_3176),
.Y(n_3192)
);

INVx1_ASAP7_75t_L g3193 ( 
.A(n_3177),
.Y(n_3193)
);

INVx1_ASAP7_75t_L g3194 ( 
.A(n_3176),
.Y(n_3194)
);

INVxp67_ASAP7_75t_L g3195 ( 
.A(n_3175),
.Y(n_3195)
);

OAI22xp5_ASAP7_75t_L g3196 ( 
.A1(n_3187),
.A2(n_3181),
.B1(n_3158),
.B2(n_3180),
.Y(n_3196)
);

AOI22xp5_ASAP7_75t_L g3197 ( 
.A1(n_3191),
.A2(n_3173),
.B1(n_3159),
.B2(n_3178),
.Y(n_3197)
);

OAI22x1_ASAP7_75t_L g3198 ( 
.A1(n_3186),
.A2(n_3182),
.B1(n_3179),
.B2(n_1041),
.Y(n_3198)
);

INVx1_ASAP7_75t_L g3199 ( 
.A(n_3185),
.Y(n_3199)
);

AO22x1_ASAP7_75t_L g3200 ( 
.A1(n_3190),
.A2(n_1107),
.B1(n_1105),
.B2(n_1096),
.Y(n_3200)
);

AOI22x1_ASAP7_75t_L g3201 ( 
.A1(n_3189),
.A2(n_3188),
.B1(n_3193),
.B2(n_3185),
.Y(n_3201)
);

AOI21xp33_ASAP7_75t_L g3202 ( 
.A1(n_3194),
.A2(n_1107),
.B(n_1084),
.Y(n_3202)
);

AOI21xp5_ASAP7_75t_L g3203 ( 
.A1(n_3199),
.A2(n_3195),
.B(n_3192),
.Y(n_3203)
);

OAI22xp5_ASAP7_75t_L g3204 ( 
.A1(n_3197),
.A2(n_3195),
.B1(n_1090),
.B2(n_1099),
.Y(n_3204)
);

OAI21xp5_ASAP7_75t_L g3205 ( 
.A1(n_3201),
.A2(n_1339),
.B(n_1382),
.Y(n_3205)
);

NAND5xp2_ASAP7_75t_L g3206 ( 
.A(n_3203),
.B(n_3196),
.C(n_3202),
.D(n_3200),
.E(n_3198),
.Y(n_3206)
);

OAI22xp5_ASAP7_75t_L g3207 ( 
.A1(n_3204),
.A2(n_1079),
.B1(n_1100),
.B2(n_1099),
.Y(n_3207)
);

AOI22xp33_ASAP7_75t_L g3208 ( 
.A1(n_3206),
.A2(n_3205),
.B1(n_1055),
.B2(n_1100),
.Y(n_3208)
);

AOI222xp33_ASAP7_75t_SL g3209 ( 
.A1(n_3207),
.A2(n_1504),
.B1(n_1450),
.B2(n_1055),
.C1(n_1485),
.C2(n_1499),
.Y(n_3209)
);

AOI22xp33_ASAP7_75t_L g3210 ( 
.A1(n_3208),
.A2(n_1055),
.B1(n_1058),
.B2(n_1100),
.Y(n_3210)
);

AOI22x1_ASAP7_75t_L g3211 ( 
.A1(n_3210),
.A2(n_3209),
.B1(n_1090),
.B2(n_1099),
.Y(n_3211)
);

AOI221xp5_ASAP7_75t_L g3212 ( 
.A1(n_3211),
.A2(n_1079),
.B1(n_1099),
.B2(n_1090),
.C(n_1058),
.Y(n_3212)
);

AOI211xp5_ASAP7_75t_L g3213 ( 
.A1(n_3212),
.A2(n_1090),
.B(n_1058),
.C(n_1064),
.Y(n_3213)
);


endmodule