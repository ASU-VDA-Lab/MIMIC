module fake_netlist_1_5391_n_47 (n_11, n_1, n_2, n_13, n_12, n_6, n_4, n_3, n_9, n_5, n_14, n_7, n_15, n_10, n_8, n_0, n_47);
input n_11;
input n_1;
input n_2;
input n_13;
input n_12;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_14;
input n_7;
input n_15;
input n_10;
input n_8;
input n_0;
output n_47;
wire n_45;
wire n_20;
wire n_38;
wire n_44;
wire n_36;
wire n_37;
wire n_34;
wire n_23;
wire n_28;
wire n_31;
wire n_22;
wire n_46;
wire n_25;
wire n_16;
wire n_26;
wire n_30;
wire n_33;
wire n_18;
wire n_32;
wire n_41;
wire n_35;
wire n_17;
wire n_42;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_43;
wire n_40;
wire n_27;
wire n_39;
BUFx6f_ASAP7_75t_L g16 ( .A(n_7), .Y(n_16) );
BUFx6f_ASAP7_75t_L g17 ( .A(n_6), .Y(n_17) );
AND2x2_ASAP7_75t_L g18 ( .A(n_13), .B(n_12), .Y(n_18) );
NAND2xp5_ASAP7_75t_SL g19 ( .A(n_14), .B(n_4), .Y(n_19) );
BUFx6f_ASAP7_75t_L g20 ( .A(n_3), .Y(n_20) );
OAI22xp5_ASAP7_75t_SL g21 ( .A1(n_9), .A2(n_6), .B1(n_2), .B2(n_5), .Y(n_21) );
AOI22xp5_ASAP7_75t_L g22 ( .A1(n_15), .A2(n_1), .B1(n_11), .B2(n_0), .Y(n_22) );
INVx2_ASAP7_75t_L g23 ( .A(n_16), .Y(n_23) );
AO22x1_ASAP7_75t_L g24 ( .A1(n_16), .A2(n_0), .B1(n_1), .B2(n_2), .Y(n_24) );
OR2x2_ASAP7_75t_L g25 ( .A(n_16), .B(n_3), .Y(n_25) );
NAND2xp5_ASAP7_75t_SL g26 ( .A(n_16), .B(n_4), .Y(n_26) );
OAI21xp5_ASAP7_75t_L g27 ( .A1(n_25), .A2(n_18), .B(n_19), .Y(n_27) );
OAI21x1_ASAP7_75t_L g28 ( .A1(n_23), .A2(n_22), .B(n_20), .Y(n_28) );
HB1xp67_ASAP7_75t_L g29 ( .A(n_28), .Y(n_29) );
AO21x2_ASAP7_75t_L g30 ( .A1(n_27), .A2(n_26), .B(n_24), .Y(n_30) );
OR2x2_ASAP7_75t_L g31 ( .A(n_30), .B(n_27), .Y(n_31) );
INVx1_ASAP7_75t_L g32 ( .A(n_29), .Y(n_32) );
OR2x2_ASAP7_75t_L g33 ( .A(n_31), .B(n_28), .Y(n_33) );
NAND2xp5_ASAP7_75t_L g34 ( .A(n_32), .B(n_30), .Y(n_34) );
AOI21xp5_ASAP7_75t_L g35 ( .A1(n_34), .A2(n_30), .B(n_26), .Y(n_35) );
INVx1_ASAP7_75t_L g36 ( .A(n_33), .Y(n_36) );
AOI22xp33_ASAP7_75t_SL g37 ( .A1(n_33), .A2(n_21), .B1(n_20), .B2(n_17), .Y(n_37) );
NAND3xp33_ASAP7_75t_L g38 ( .A(n_37), .B(n_17), .C(n_20), .Y(n_38) );
AOI21xp5_ASAP7_75t_L g39 ( .A1(n_35), .A2(n_17), .B(n_20), .Y(n_39) );
AOI211xp5_ASAP7_75t_SL g40 ( .A1(n_36), .A2(n_5), .B(n_7), .C(n_8), .Y(n_40) );
INVx2_ASAP7_75t_SL g41 ( .A(n_38), .Y(n_41) );
INVx2_ASAP7_75t_L g42 ( .A(n_40), .Y(n_42) );
NOR2x2_ASAP7_75t_L g43 ( .A(n_39), .B(n_8), .Y(n_43) );
OAI22x1_ASAP7_75t_SL g44 ( .A1(n_42), .A2(n_9), .B1(n_10), .B2(n_17), .Y(n_44) );
CKINVDCx5p33_ASAP7_75t_R g45 ( .A(n_41), .Y(n_45) );
AND3x4_ASAP7_75t_L g46 ( .A(n_44), .B(n_43), .C(n_10), .Y(n_46) );
OA21x2_ASAP7_75t_L g47 ( .A1(n_46), .A2(n_45), .B(n_44), .Y(n_47) );
endmodule