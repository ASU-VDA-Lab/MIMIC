module fake_jpeg_29418_n_60 (n_13, n_21, n_1, n_10, n_6, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_60);

input n_13;
input n_21;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_60;

wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_45;
wire n_23;
wire n_27;
wire n_55;
wire n_22;
wire n_47;
wire n_51;
wire n_40;
wire n_59;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_31;
wire n_25;
wire n_56;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_32;

INVx5_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

INVx8_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_26),
.B(n_0),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_28),
.B(n_29),
.Y(n_40)
);

INVxp67_ASAP7_75t_L g29 ( 
.A(n_24),
.Y(n_29)
);

AOI22xp33_ASAP7_75t_SL g30 ( 
.A1(n_26),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_30)
);

O2A1O1Ixp33_ASAP7_75t_L g42 ( 
.A1(n_30),
.A2(n_33),
.B(n_15),
.C(n_21),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_26),
.B(n_2),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_31),
.Y(n_36)
);

HB1xp67_ASAP7_75t_L g32 ( 
.A(n_25),
.Y(n_32)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_32),
.Y(n_35)
);

OAI22xp33_ASAP7_75t_SL g33 ( 
.A1(n_25),
.A2(n_13),
.B1(n_20),
.B2(n_19),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_27),
.B(n_3),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_34),
.Y(n_39)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_28),
.Y(n_37)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_37),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_29),
.B(n_23),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_38),
.B(n_42),
.Y(n_46)
);

INVx5_ASAP7_75t_L g41 ( 
.A(n_29),
.Y(n_41)
);

AND2x2_ASAP7_75t_L g44 ( 
.A(n_41),
.B(n_4),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_SL g43 ( 
.A1(n_42),
.A2(n_27),
.B1(n_22),
.B2(n_6),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_43),
.B(n_49),
.Y(n_54)
);

CKINVDCx14_ASAP7_75t_R g52 ( 
.A(n_44),
.Y(n_52)
);

MAJIxp5_ASAP7_75t_L g45 ( 
.A(n_38),
.B(n_11),
.C(n_17),
.Y(n_45)
);

MAJIxp5_ASAP7_75t_L g53 ( 
.A(n_45),
.B(n_47),
.C(n_44),
.Y(n_53)
);

OAI21xp5_ASAP7_75t_SL g47 ( 
.A1(n_40),
.A2(n_4),
.B(n_5),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g49 ( 
.A1(n_35),
.A2(n_9),
.B1(n_10),
.B2(n_16),
.Y(n_49)
);

AOI21xp5_ASAP7_75t_SL g50 ( 
.A1(n_46),
.A2(n_41),
.B(n_36),
.Y(n_50)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_50),
.Y(n_55)
);

XNOR2xp5_ASAP7_75t_L g51 ( 
.A(n_48),
.B(n_39),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_51),
.B(n_53),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g56 ( 
.A1(n_52),
.A2(n_5),
.B1(n_18),
.B2(n_45),
.Y(n_56)
);

HB1xp67_ASAP7_75t_L g58 ( 
.A(n_56),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_58),
.Y(n_59)
);

NOR4xp25_ASAP7_75t_L g60 ( 
.A(n_59),
.B(n_54),
.C(n_55),
.D(n_57),
.Y(n_60)
);


endmodule