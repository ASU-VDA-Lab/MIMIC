module fake_netlist_6_1457_n_1804 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_68, n_28, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_144, n_127, n_125, n_153, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_159, n_157, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_1804);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_68;
input n_28;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_144;
input n_127;
input n_125;
input n_153;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1804;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_168;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_783;
wire n_1738;
wire n_798;
wire n_188;
wire n_1575;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1691;
wire n_1688;
wire n_1009;
wire n_1743;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_1786;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_200;
wire n_447;
wire n_1803;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1704;
wire n_1078;
wire n_250;
wire n_544;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_616;
wire n_658;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1620;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1798;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_163;
wire n_1644;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_577;
wire n_166;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1762;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1697;
wire n_243;
wire n_979;
wire n_905;
wire n_1680;
wire n_175;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_530;
wire n_1563;
wire n_277;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_1760;
wire n_210;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_178;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_429;
wire n_1747;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1802;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_1801;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_697;
wire n_687;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_1709;
wire n_1757;
wire n_1796;
wire n_170;
wire n_1792;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_161;
wire n_462;
wire n_1052;
wire n_1033;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_297;
wire n_595;
wire n_627;
wire n_1767;
wire n_1779;
wire n_524;
wire n_1465;
wire n_342;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_1765;
wire n_353;
wire n_605;
wire n_1514;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_173;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_1788;
wire n_622;
wire n_1469;
wire n_1766;
wire n_1776;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_1771;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_899;
wire n_189;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1577;
wire n_1181;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_927;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_184;
wire n_552;
wire n_1358;
wire n_1388;
wire n_216;
wire n_912;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_527;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_211;
wire n_1483;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_1787;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1769;
wire n_1220;
wire n_556;
wire n_162;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1775;
wire n_1773;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_1745;
wire n_914;
wire n_759;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1580;
wire n_1425;
wire n_1267;
wire n_1281;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_177;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1594;
wire n_664;
wire n_171;
wire n_1764;
wire n_169;
wire n_1429;
wire n_1610;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_160;
wire n_186;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1024;
wire n_1768;
wire n_198;
wire n_179;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1639;
wire n_1623;
wire n_183;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1686;
wire n_167;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1262;
wire n_218;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_172;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1361;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_370;
wire n_1695;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_227;
wire n_1720;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_1795;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1489;
wire n_164;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_1782;
wire n_282;
wire n_1676;
wire n_833;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_1086;
wire n_1066;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_1758;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1794;
wire n_1236;
wire n_1559;
wire n_1725;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1746;
wire n_1325;
wire n_1002;
wire n_1741;
wire n_545;
wire n_489;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_187;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1800;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_566;
wire n_1023;
wire n_1118;
wire n_1076;
wire n_194;
wire n_1007;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1631;
wire n_591;
wire n_1377;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_180;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_181;
wire n_182;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_1729;
wire n_669;
wire n_176;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1785;
wire n_763;
wire n_1147;
wire n_360;
wire n_1754;
wire n_1506;
wire n_1652;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_174;
wire n_1173;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_185;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1525;
wire n_455;
wire n_1585;
wire n_363;
wire n_1799;
wire n_1090;
wire n_592;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_1789;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_404;
wire n_271;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_373;
wire n_1632;
wire n_257;
wire n_1557;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_207;
wire n_1089;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_339;
wire n_784;
wire n_434;
wire n_315;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_165;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_1259;
wire n_192;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

INVx1_ASAP7_75t_L g160 ( 
.A(n_120),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_112),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_119),
.Y(n_162)
);

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_113),
.Y(n_163)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_70),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_101),
.Y(n_165)
);

BUFx10_ASAP7_75t_L g166 ( 
.A(n_9),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_1),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_91),
.Y(n_168)
);

INVx3_ASAP7_75t_L g169 ( 
.A(n_103),
.Y(n_169)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_53),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_51),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_61),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_158),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_132),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_17),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_153),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_9),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_145),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_137),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_142),
.Y(n_180)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_17),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_10),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_43),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_69),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_18),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_12),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_16),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_136),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_131),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_32),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_40),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_159),
.Y(n_192)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_90),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_5),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_58),
.Y(n_195)
);

BUFx2_ASAP7_75t_L g196 ( 
.A(n_151),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_73),
.Y(n_197)
);

BUFx3_ASAP7_75t_L g198 ( 
.A(n_18),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_157),
.Y(n_199)
);

INVxp67_ASAP7_75t_L g200 ( 
.A(n_6),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_93),
.Y(n_201)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_99),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_21),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_114),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_111),
.Y(n_205)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_135),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_130),
.Y(n_207)
);

INVx1_ASAP7_75t_SL g208 ( 
.A(n_121),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_97),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_98),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_110),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_107),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_40),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_76),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_141),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_45),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_147),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_10),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_65),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_63),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_35),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_3),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_85),
.Y(n_223)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_29),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_118),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_64),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_102),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_127),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_106),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_116),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_47),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_28),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_125),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_154),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_139),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_105),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_8),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_11),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_25),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_72),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_46),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_115),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_56),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_19),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_27),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_81),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_44),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_129),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_84),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_60),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_2),
.Y(n_251)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_156),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_21),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_78),
.Y(n_254)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_67),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_2),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_149),
.Y(n_257)
);

BUFx6f_ASAP7_75t_L g258 ( 
.A(n_109),
.Y(n_258)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_117),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_29),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_79),
.Y(n_261)
);

CKINVDCx16_ASAP7_75t_R g262 ( 
.A(n_14),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_23),
.Y(n_263)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_51),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_52),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_14),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_144),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_148),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_133),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_33),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_49),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_25),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_5),
.Y(n_273)
);

BUFx10_ASAP7_75t_L g274 ( 
.A(n_32),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_94),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_60),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_11),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_56),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_87),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_20),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_52),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_134),
.Y(n_282)
);

INVx1_ASAP7_75t_SL g283 ( 
.A(n_46),
.Y(n_283)
);

BUFx10_ASAP7_75t_L g284 ( 
.A(n_53),
.Y(n_284)
);

INVx1_ASAP7_75t_SL g285 ( 
.A(n_71),
.Y(n_285)
);

CKINVDCx16_ASAP7_75t_R g286 ( 
.A(n_68),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_62),
.Y(n_287)
);

BUFx6f_ASAP7_75t_L g288 ( 
.A(n_22),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_12),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_66),
.Y(n_290)
);

BUFx3_ASAP7_75t_L g291 ( 
.A(n_50),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_138),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_150),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_19),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_8),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_45),
.Y(n_296)
);

INVx1_ASAP7_75t_SL g297 ( 
.A(n_49),
.Y(n_297)
);

BUFx6f_ASAP7_75t_L g298 ( 
.A(n_34),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_123),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_155),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g301 ( 
.A(n_20),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_77),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_48),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_4),
.Y(n_304)
);

INVx1_ASAP7_75t_SL g305 ( 
.A(n_74),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_48),
.Y(n_306)
);

INVx2_ASAP7_75t_L g307 ( 
.A(n_42),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_1),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_24),
.Y(n_309)
);

INVx1_ASAP7_75t_SL g310 ( 
.A(n_89),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_58),
.Y(n_311)
);

INVx1_ASAP7_75t_SL g312 ( 
.A(n_59),
.Y(n_312)
);

BUFx2_ASAP7_75t_L g313 ( 
.A(n_54),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_7),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_126),
.Y(n_315)
);

INVx1_ASAP7_75t_SL g316 ( 
.A(n_36),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_104),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_288),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_288),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_288),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_288),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_288),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_288),
.Y(n_323)
);

INVxp67_ASAP7_75t_SL g324 ( 
.A(n_196),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_298),
.Y(n_325)
);

BUFx2_ASAP7_75t_L g326 ( 
.A(n_313),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_298),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_161),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_298),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_298),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_163),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_298),
.Y(n_332)
);

INVx2_ASAP7_75t_L g333 ( 
.A(n_298),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_168),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_173),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_181),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_174),
.Y(n_337)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_214),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_196),
.B(n_0),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_181),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_181),
.Y(n_341)
);

CKINVDCx20_ASAP7_75t_R g342 ( 
.A(n_233),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_170),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_176),
.Y(n_344)
);

BUFx6f_ASAP7_75t_SL g345 ( 
.A(n_258),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_170),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_224),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_178),
.Y(n_348)
);

CKINVDCx20_ASAP7_75t_R g349 ( 
.A(n_235),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_179),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_224),
.Y(n_351)
);

INVxp67_ASAP7_75t_SL g352 ( 
.A(n_169),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_188),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_L g354 ( 
.A(n_160),
.B(n_0),
.Y(n_354)
);

NOR2xp67_ASAP7_75t_L g355 ( 
.A(n_169),
.B(n_3),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_264),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_264),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_189),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_192),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_307),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_197),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_307),
.Y(n_362)
);

INVxp67_ASAP7_75t_L g363 ( 
.A(n_313),
.Y(n_363)
);

CKINVDCx20_ASAP7_75t_R g364 ( 
.A(n_286),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_199),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_201),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_205),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_198),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_207),
.Y(n_369)
);

CKINVDCx20_ASAP7_75t_R g370 ( 
.A(n_286),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_198),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_210),
.Y(n_372)
);

CKINVDCx20_ASAP7_75t_R g373 ( 
.A(n_211),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_212),
.Y(n_374)
);

INVx1_ASAP7_75t_SL g375 ( 
.A(n_216),
.Y(n_375)
);

CKINVDCx20_ASAP7_75t_R g376 ( 
.A(n_219),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_223),
.Y(n_377)
);

INVxp67_ASAP7_75t_SL g378 ( 
.A(n_169),
.Y(n_378)
);

BUFx3_ASAP7_75t_L g379 ( 
.A(n_160),
.Y(n_379)
);

CKINVDCx20_ASAP7_75t_R g380 ( 
.A(n_225),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_226),
.Y(n_381)
);

NOR2xp33_ASAP7_75t_L g382 ( 
.A(n_162),
.B(n_4),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_198),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_291),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_230),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_234),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_236),
.Y(n_387)
);

NOR2xp67_ASAP7_75t_L g388 ( 
.A(n_169),
.B(n_6),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_291),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_240),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_291),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_167),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_167),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_318),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_352),
.B(n_242),
.Y(n_395)
);

OAI22xp5_ASAP7_75t_L g396 ( 
.A1(n_363),
.A2(n_262),
.B1(n_301),
.B2(n_244),
.Y(n_396)
);

INVx2_ASAP7_75t_L g397 ( 
.A(n_333),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_318),
.Y(n_398)
);

INVx2_ASAP7_75t_L g399 ( 
.A(n_333),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_319),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_378),
.B(n_317),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_368),
.B(n_246),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_368),
.B(n_371),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_371),
.B(n_248),
.Y(n_404)
);

INVx3_ASAP7_75t_L g405 ( 
.A(n_319),
.Y(n_405)
);

INVx2_ASAP7_75t_L g406 ( 
.A(n_320),
.Y(n_406)
);

AND2x2_ASAP7_75t_L g407 ( 
.A(n_383),
.B(n_164),
.Y(n_407)
);

INVx3_ASAP7_75t_L g408 ( 
.A(n_320),
.Y(n_408)
);

BUFx6f_ASAP7_75t_L g409 ( 
.A(n_321),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_321),
.Y(n_410)
);

BUFx6f_ASAP7_75t_L g411 ( 
.A(n_322),
.Y(n_411)
);

INVx2_ASAP7_75t_L g412 ( 
.A(n_322),
.Y(n_412)
);

INVx3_ASAP7_75t_L g413 ( 
.A(n_323),
.Y(n_413)
);

INVx2_ASAP7_75t_L g414 ( 
.A(n_323),
.Y(n_414)
);

BUFx2_ASAP7_75t_L g415 ( 
.A(n_364),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_383),
.B(n_257),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_325),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_325),
.Y(n_418)
);

INVx2_ASAP7_75t_L g419 ( 
.A(n_327),
.Y(n_419)
);

BUFx6f_ASAP7_75t_L g420 ( 
.A(n_327),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_373),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_329),
.Y(n_422)
);

INVx2_ASAP7_75t_L g423 ( 
.A(n_329),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_330),
.Y(n_424)
);

INVx2_ASAP7_75t_L g425 ( 
.A(n_330),
.Y(n_425)
);

INVx2_ASAP7_75t_L g426 ( 
.A(n_332),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_332),
.Y(n_427)
);

INVx6_ASAP7_75t_L g428 ( 
.A(n_379),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_392),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_392),
.Y(n_430)
);

BUFx6f_ASAP7_75t_L g431 ( 
.A(n_336),
.Y(n_431)
);

INVx2_ASAP7_75t_L g432 ( 
.A(n_336),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_376),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_393),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_393),
.Y(n_435)
);

INVx2_ASAP7_75t_L g436 ( 
.A(n_340),
.Y(n_436)
);

AND2x4_ASAP7_75t_L g437 ( 
.A(n_355),
.B(n_164),
.Y(n_437)
);

INVxp67_ASAP7_75t_L g438 ( 
.A(n_326),
.Y(n_438)
);

INVx2_ASAP7_75t_L g439 ( 
.A(n_340),
.Y(n_439)
);

NOR2xp33_ASAP7_75t_L g440 ( 
.A(n_339),
.B(n_262),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_L g441 ( 
.A(n_384),
.B(n_261),
.Y(n_441)
);

AND3x1_ASAP7_75t_L g442 ( 
.A(n_354),
.B(n_195),
.C(n_183),
.Y(n_442)
);

AND2x6_ASAP7_75t_L g443 ( 
.A(n_382),
.B(n_164),
.Y(n_443)
);

NAND2xp33_ASAP7_75t_R g444 ( 
.A(n_326),
.B(n_171),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_SL g445 ( 
.A(n_355),
.B(n_166),
.Y(n_445)
);

HB1xp67_ASAP7_75t_L g446 ( 
.A(n_384),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_341),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_341),
.Y(n_448)
);

NAND2xp33_ASAP7_75t_L g449 ( 
.A(n_389),
.B(n_258),
.Y(n_449)
);

HB1xp67_ASAP7_75t_L g450 ( 
.A(n_389),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_343),
.Y(n_451)
);

BUFx6f_ASAP7_75t_L g452 ( 
.A(n_343),
.Y(n_452)
);

BUFx6f_ASAP7_75t_L g453 ( 
.A(n_346),
.Y(n_453)
);

INVx2_ASAP7_75t_L g454 ( 
.A(n_346),
.Y(n_454)
);

INVx2_ASAP7_75t_L g455 ( 
.A(n_347),
.Y(n_455)
);

INVx2_ASAP7_75t_L g456 ( 
.A(n_347),
.Y(n_456)
);

BUFx6f_ASAP7_75t_L g457 ( 
.A(n_351),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_351),
.Y(n_458)
);

BUFx6f_ASAP7_75t_L g459 ( 
.A(n_356),
.Y(n_459)
);

INVx2_ASAP7_75t_L g460 ( 
.A(n_356),
.Y(n_460)
);

BUFx6f_ASAP7_75t_L g461 ( 
.A(n_357),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_357),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_360),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_360),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_362),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_394),
.Y(n_466)
);

INVxp67_ASAP7_75t_SL g467 ( 
.A(n_446),
.Y(n_467)
);

BUFx3_ASAP7_75t_L g468 ( 
.A(n_428),
.Y(n_468)
);

INVx2_ASAP7_75t_L g469 ( 
.A(n_406),
.Y(n_469)
);

INVx2_ASAP7_75t_L g470 ( 
.A(n_406),
.Y(n_470)
);

INVx3_ASAP7_75t_L g471 ( 
.A(n_409),
.Y(n_471)
);

NAND3xp33_ASAP7_75t_L g472 ( 
.A(n_440),
.B(n_442),
.C(n_437),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_394),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_398),
.Y(n_474)
);

NAND2xp33_ASAP7_75t_R g475 ( 
.A(n_415),
.B(n_328),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_398),
.Y(n_476)
);

INVx2_ASAP7_75t_L g477 ( 
.A(n_406),
.Y(n_477)
);

AND2x2_ASAP7_75t_L g478 ( 
.A(n_407),
.B(n_379),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_400),
.Y(n_479)
);

HB1xp67_ASAP7_75t_L g480 ( 
.A(n_438),
.Y(n_480)
);

AND2x4_ASAP7_75t_L g481 ( 
.A(n_437),
.B(n_388),
.Y(n_481)
);

NOR2xp33_ASAP7_75t_L g482 ( 
.A(n_395),
.B(n_331),
.Y(n_482)
);

INVx3_ASAP7_75t_L g483 ( 
.A(n_409),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_400),
.Y(n_484)
);

INVxp33_ASAP7_75t_L g485 ( 
.A(n_396),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_SL g486 ( 
.A(n_440),
.B(n_334),
.Y(n_486)
);

AOI22xp33_ASAP7_75t_L g487 ( 
.A1(n_443),
.A2(n_324),
.B1(n_238),
.B2(n_296),
.Y(n_487)
);

INVx2_ASAP7_75t_L g488 ( 
.A(n_406),
.Y(n_488)
);

INVxp33_ASAP7_75t_L g489 ( 
.A(n_396),
.Y(n_489)
);

INVx2_ASAP7_75t_L g490 ( 
.A(n_412),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_SL g491 ( 
.A(n_395),
.B(n_335),
.Y(n_491)
);

OR2x6_ASAP7_75t_L g492 ( 
.A(n_445),
.B(n_162),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_410),
.Y(n_493)
);

BUFx2_ASAP7_75t_L g494 ( 
.A(n_438),
.Y(n_494)
);

INVx2_ASAP7_75t_L g495 ( 
.A(n_412),
.Y(n_495)
);

INVx3_ASAP7_75t_L g496 ( 
.A(n_409),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_L g497 ( 
.A(n_401),
.B(n_337),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_410),
.Y(n_498)
);

OR2x2_ASAP7_75t_L g499 ( 
.A(n_402),
.B(n_375),
.Y(n_499)
);

AND2x6_ASAP7_75t_L g500 ( 
.A(n_437),
.B(n_258),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_L g501 ( 
.A(n_401),
.B(n_344),
.Y(n_501)
);

INVx4_ASAP7_75t_L g502 ( 
.A(n_409),
.Y(n_502)
);

INVx2_ASAP7_75t_L g503 ( 
.A(n_412),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_SL g504 ( 
.A(n_442),
.B(n_348),
.Y(n_504)
);

INVx3_ASAP7_75t_L g505 ( 
.A(n_409),
.Y(n_505)
);

NOR2xp33_ASAP7_75t_L g506 ( 
.A(n_402),
.B(n_350),
.Y(n_506)
);

INVx2_ASAP7_75t_L g507 ( 
.A(n_412),
.Y(n_507)
);

INVx3_ASAP7_75t_L g508 ( 
.A(n_409),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_L g509 ( 
.A(n_428),
.B(n_353),
.Y(n_509)
);

INVx2_ASAP7_75t_L g510 ( 
.A(n_414),
.Y(n_510)
);

NOR2xp33_ASAP7_75t_L g511 ( 
.A(n_404),
.B(n_358),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_417),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_417),
.Y(n_513)
);

AOI22xp5_ASAP7_75t_L g514 ( 
.A1(n_443),
.A2(n_276),
.B1(n_221),
.B2(n_314),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_428),
.B(n_359),
.Y(n_515)
);

CKINVDCx6p67_ASAP7_75t_R g516 ( 
.A(n_415),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_418),
.Y(n_517)
);

AND2x6_ASAP7_75t_L g518 ( 
.A(n_437),
.B(n_258),
.Y(n_518)
);

BUFx10_ASAP7_75t_L g519 ( 
.A(n_421),
.Y(n_519)
);

INVxp67_ASAP7_75t_L g520 ( 
.A(n_444),
.Y(n_520)
);

BUFx6f_ASAP7_75t_SL g521 ( 
.A(n_437),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_418),
.Y(n_522)
);

NAND2xp33_ASAP7_75t_L g523 ( 
.A(n_443),
.B(n_361),
.Y(n_523)
);

INVx2_ASAP7_75t_L g524 ( 
.A(n_414),
.Y(n_524)
);

AOI22xp5_ASAP7_75t_L g525 ( 
.A1(n_443),
.A2(n_311),
.B1(n_297),
.B2(n_283),
.Y(n_525)
);

BUFx3_ASAP7_75t_L g526 ( 
.A(n_428),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_L g527 ( 
.A(n_428),
.B(n_365),
.Y(n_527)
);

BUFx3_ASAP7_75t_L g528 ( 
.A(n_428),
.Y(n_528)
);

AND2x4_ASAP7_75t_L g529 ( 
.A(n_437),
.B(n_165),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_422),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_422),
.Y(n_531)
);

INVx3_ASAP7_75t_L g532 ( 
.A(n_409),
.Y(n_532)
);

INVxp33_ASAP7_75t_L g533 ( 
.A(n_415),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_L g534 ( 
.A(n_404),
.B(n_366),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_SL g535 ( 
.A(n_416),
.B(n_367),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_424),
.Y(n_536)
);

BUFx3_ASAP7_75t_L g537 ( 
.A(n_424),
.Y(n_537)
);

INVx3_ASAP7_75t_L g538 ( 
.A(n_409),
.Y(n_538)
);

AND2x4_ASAP7_75t_L g539 ( 
.A(n_407),
.B(n_165),
.Y(n_539)
);

NOR2xp33_ASAP7_75t_L g540 ( 
.A(n_416),
.B(n_369),
.Y(n_540)
);

NOR2xp33_ASAP7_75t_L g541 ( 
.A(n_441),
.B(n_372),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_L g542 ( 
.A(n_441),
.B(n_374),
.Y(n_542)
);

INVx2_ASAP7_75t_L g543 ( 
.A(n_414),
.Y(n_543)
);

AND2x2_ASAP7_75t_L g544 ( 
.A(n_407),
.B(n_391),
.Y(n_544)
);

OAI22xp33_ASAP7_75t_L g545 ( 
.A1(n_444),
.A2(n_312),
.B1(n_316),
.B2(n_247),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_SL g546 ( 
.A(n_445),
.B(n_377),
.Y(n_546)
);

AND3x1_ASAP7_75t_L g547 ( 
.A(n_446),
.B(n_195),
.C(n_183),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_427),
.Y(n_548)
);

BUFx10_ASAP7_75t_L g549 ( 
.A(n_421),
.Y(n_549)
);

NAND2xp33_ASAP7_75t_SL g550 ( 
.A(n_450),
.B(n_370),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_427),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_SL g552 ( 
.A(n_450),
.B(n_381),
.Y(n_552)
);

CKINVDCx6p67_ASAP7_75t_R g553 ( 
.A(n_443),
.Y(n_553)
);

AOI22xp33_ASAP7_75t_L g554 ( 
.A1(n_443),
.A2(n_296),
.B1(n_280),
.B2(n_281),
.Y(n_554)
);

INVx2_ASAP7_75t_L g555 ( 
.A(n_414),
.Y(n_555)
);

INVx2_ASAP7_75t_L g556 ( 
.A(n_419),
.Y(n_556)
);

INVx2_ASAP7_75t_SL g557 ( 
.A(n_443),
.Y(n_557)
);

AND2x4_ASAP7_75t_L g558 ( 
.A(n_429),
.B(n_172),
.Y(n_558)
);

INVx1_ASAP7_75t_SL g559 ( 
.A(n_433),
.Y(n_559)
);

BUFx6f_ASAP7_75t_L g560 ( 
.A(n_411),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_L g561 ( 
.A(n_443),
.B(n_385),
.Y(n_561)
);

INVx2_ASAP7_75t_L g562 ( 
.A(n_419),
.Y(n_562)
);

INVx6_ASAP7_75t_L g563 ( 
.A(n_411),
.Y(n_563)
);

INVx3_ASAP7_75t_L g564 ( 
.A(n_411),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_429),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_430),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_430),
.Y(n_567)
);

NOR2x1p5_ASAP7_75t_L g568 ( 
.A(n_403),
.B(n_238),
.Y(n_568)
);

INVx3_ASAP7_75t_L g569 ( 
.A(n_411),
.Y(n_569)
);

INVx1_ASAP7_75t_SL g570 ( 
.A(n_433),
.Y(n_570)
);

INVx2_ASAP7_75t_L g571 ( 
.A(n_419),
.Y(n_571)
);

NOR2xp33_ASAP7_75t_L g572 ( 
.A(n_403),
.B(n_386),
.Y(n_572)
);

BUFx3_ASAP7_75t_L g573 ( 
.A(n_434),
.Y(n_573)
);

BUFx6f_ASAP7_75t_L g574 ( 
.A(n_411),
.Y(n_574)
);

INVx2_ASAP7_75t_L g575 ( 
.A(n_419),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_SL g576 ( 
.A(n_434),
.B(n_387),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_435),
.Y(n_577)
);

INVx2_ASAP7_75t_L g578 ( 
.A(n_423),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_435),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_L g580 ( 
.A(n_443),
.B(n_390),
.Y(n_580)
);

INVx2_ASAP7_75t_L g581 ( 
.A(n_423),
.Y(n_581)
);

AOI22xp33_ASAP7_75t_L g582 ( 
.A1(n_443),
.A2(n_245),
.B1(n_294),
.B2(n_289),
.Y(n_582)
);

INVx3_ASAP7_75t_L g583 ( 
.A(n_411),
.Y(n_583)
);

INVx2_ASAP7_75t_L g584 ( 
.A(n_423),
.Y(n_584)
);

NAND2xp5_ASAP7_75t_SL g585 ( 
.A(n_465),
.B(n_380),
.Y(n_585)
);

BUFx6f_ASAP7_75t_L g586 ( 
.A(n_411),
.Y(n_586)
);

INVx2_ASAP7_75t_SL g587 ( 
.A(n_443),
.Y(n_587)
);

AO22x2_ASAP7_75t_L g588 ( 
.A1(n_451),
.A2(n_241),
.B1(n_245),
.B2(n_250),
.Y(n_588)
);

INVx4_ASAP7_75t_L g589 ( 
.A(n_411),
.Y(n_589)
);

INVx2_ASAP7_75t_L g590 ( 
.A(n_423),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_405),
.Y(n_591)
);

OR2x6_ASAP7_75t_L g592 ( 
.A(n_451),
.B(n_172),
.Y(n_592)
);

BUFx4f_ASAP7_75t_L g593 ( 
.A(n_420),
.Y(n_593)
);

INVx2_ASAP7_75t_L g594 ( 
.A(n_425),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_SL g595 ( 
.A(n_465),
.B(n_268),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_405),
.Y(n_596)
);

NOR2xp33_ASAP7_75t_L g597 ( 
.A(n_458),
.B(n_391),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_SL g598 ( 
.A(n_458),
.B(n_269),
.Y(n_598)
);

AND2x6_ASAP7_75t_L g599 ( 
.A(n_405),
.B(n_258),
.Y(n_599)
);

INVx2_ASAP7_75t_L g600 ( 
.A(n_425),
.Y(n_600)
);

INVx2_ASAP7_75t_L g601 ( 
.A(n_425),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_L g602 ( 
.A(n_405),
.B(n_208),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_405),
.Y(n_603)
);

INVx2_ASAP7_75t_L g604 ( 
.A(n_425),
.Y(n_604)
);

INVx3_ASAP7_75t_L g605 ( 
.A(n_420),
.Y(n_605)
);

HB1xp67_ASAP7_75t_L g606 ( 
.A(n_447),
.Y(n_606)
);

INVx2_ASAP7_75t_L g607 ( 
.A(n_426),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_408),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_408),
.Y(n_609)
);

INVxp67_ASAP7_75t_L g610 ( 
.A(n_462),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_L g611 ( 
.A(n_408),
.B(n_285),
.Y(n_611)
);

AND3x2_ASAP7_75t_L g612 ( 
.A(n_462),
.B(n_200),
.C(n_193),
.Y(n_612)
);

NOR2xp33_ASAP7_75t_L g613 ( 
.A(n_463),
.B(n_338),
.Y(n_613)
);

INVx2_ASAP7_75t_L g614 ( 
.A(n_426),
.Y(n_614)
);

AOI22xp33_ASAP7_75t_L g615 ( 
.A1(n_447),
.A2(n_260),
.B1(n_241),
.B2(n_250),
.Y(n_615)
);

A2O1A1Ixp33_ASAP7_75t_L g616 ( 
.A1(n_472),
.A2(n_193),
.B(n_202),
.C(n_206),
.Y(n_616)
);

AOI22xp5_ASAP7_75t_L g617 ( 
.A1(n_472),
.A2(n_349),
.B1(n_342),
.B2(n_310),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_L g618 ( 
.A(n_482),
.B(n_408),
.Y(n_618)
);

NAND2x1p5_ASAP7_75t_L g619 ( 
.A(n_557),
.B(n_180),
.Y(n_619)
);

NOR2xp67_ASAP7_75t_L g620 ( 
.A(n_520),
.B(n_448),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_606),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_L g622 ( 
.A(n_572),
.B(n_506),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_L g623 ( 
.A(n_511),
.B(n_408),
.Y(n_623)
);

INVx2_ASAP7_75t_L g624 ( 
.A(n_466),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_565),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_L g626 ( 
.A(n_540),
.B(n_413),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_SL g627 ( 
.A(n_557),
.B(n_258),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_L g628 ( 
.A(n_541),
.B(n_413),
.Y(n_628)
);

INVx2_ASAP7_75t_L g629 ( 
.A(n_466),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_565),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_L g631 ( 
.A(n_497),
.B(n_413),
.Y(n_631)
);

AOI22xp5_ASAP7_75t_L g632 ( 
.A1(n_504),
.A2(n_305),
.B1(n_279),
.B2(n_275),
.Y(n_632)
);

INVx1_ASAP7_75t_SL g633 ( 
.A(n_494),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_L g634 ( 
.A(n_501),
.B(n_413),
.Y(n_634)
);

NOR3xp33_ASAP7_75t_L g635 ( 
.A(n_545),
.B(n_177),
.C(n_175),
.Y(n_635)
);

BUFx6f_ASAP7_75t_L g636 ( 
.A(n_468),
.Y(n_636)
);

NOR2xp67_ASAP7_75t_L g637 ( 
.A(n_499),
.B(n_448),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_SL g638 ( 
.A(n_587),
.B(n_202),
.Y(n_638)
);

NOR2xp33_ASAP7_75t_L g639 ( 
.A(n_499),
.B(n_182),
.Y(n_639)
);

INVxp67_ASAP7_75t_L g640 ( 
.A(n_494),
.Y(n_640)
);

CKINVDCx5p33_ASAP7_75t_R g641 ( 
.A(n_475),
.Y(n_641)
);

INVx2_ASAP7_75t_SL g642 ( 
.A(n_568),
.Y(n_642)
);

AND2x2_ASAP7_75t_L g643 ( 
.A(n_467),
.B(n_463),
.Y(n_643)
);

INVx2_ASAP7_75t_L g644 ( 
.A(n_473),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_L g645 ( 
.A(n_481),
.B(n_534),
.Y(n_645)
);

NOR2xp33_ASAP7_75t_L g646 ( 
.A(n_542),
.B(n_185),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_L g647 ( 
.A(n_481),
.B(n_413),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_566),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_L g649 ( 
.A(n_481),
.B(n_573),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_566),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_L g651 ( 
.A(n_481),
.B(n_573),
.Y(n_651)
);

INVx3_ASAP7_75t_L g652 ( 
.A(n_573),
.Y(n_652)
);

NOR2xp33_ASAP7_75t_L g653 ( 
.A(n_486),
.B(n_186),
.Y(n_653)
);

INVx3_ASAP7_75t_R g654 ( 
.A(n_558),
.Y(n_654)
);

OAI22xp33_ASAP7_75t_SL g655 ( 
.A1(n_525),
.A2(n_229),
.B1(n_217),
.B2(n_315),
.Y(n_655)
);

NOR2xp33_ASAP7_75t_L g656 ( 
.A(n_491),
.B(n_187),
.Y(n_656)
);

INVx2_ASAP7_75t_L g657 ( 
.A(n_473),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_L g658 ( 
.A(n_544),
.B(n_452),
.Y(n_658)
);

O2A1O1Ixp5_ASAP7_75t_L g659 ( 
.A1(n_539),
.A2(n_259),
.B(n_255),
.C(n_252),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_L g660 ( 
.A(n_544),
.B(n_452),
.Y(n_660)
);

NAND2xp33_ASAP7_75t_SL g661 ( 
.A(n_485),
.B(n_489),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_SL g662 ( 
.A(n_587),
.B(n_206),
.Y(n_662)
);

AOI22xp5_ASAP7_75t_L g663 ( 
.A1(n_525),
.A2(n_292),
.B1(n_282),
.B2(n_293),
.Y(n_663)
);

INVx2_ASAP7_75t_L g664 ( 
.A(n_474),
.Y(n_664)
);

INVx2_ASAP7_75t_L g665 ( 
.A(n_474),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_L g666 ( 
.A(n_478),
.B(n_452),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_567),
.Y(n_667)
);

NOR2xp33_ASAP7_75t_L g668 ( 
.A(n_535),
.B(n_190),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_L g669 ( 
.A(n_478),
.B(n_452),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_L g670 ( 
.A(n_537),
.B(n_567),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_L g671 ( 
.A(n_537),
.B(n_452),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_L g672 ( 
.A(n_577),
.B(n_452),
.Y(n_672)
);

AND2x2_ASAP7_75t_L g673 ( 
.A(n_480),
.B(n_464),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_SL g674 ( 
.A(n_561),
.B(n_252),
.Y(n_674)
);

INVx2_ASAP7_75t_L g675 ( 
.A(n_476),
.Y(n_675)
);

OAI22xp33_ASAP7_75t_SL g676 ( 
.A1(n_514),
.A2(n_228),
.B1(n_229),
.B2(n_227),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_L g677 ( 
.A(n_577),
.B(n_452),
.Y(n_677)
);

AOI22xp33_ASAP7_75t_L g678 ( 
.A1(n_554),
.A2(n_260),
.B1(n_278),
.B2(n_280),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_L g679 ( 
.A(n_579),
.B(n_539),
.Y(n_679)
);

INVx3_ASAP7_75t_L g680 ( 
.A(n_521),
.Y(n_680)
);

AOI22xp33_ASAP7_75t_L g681 ( 
.A1(n_582),
.A2(n_278),
.B1(n_281),
.B2(n_289),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_579),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_L g683 ( 
.A(n_539),
.B(n_453),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_539),
.B(n_453),
.Y(n_684)
);

CKINVDCx14_ASAP7_75t_R g685 ( 
.A(n_516),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_SL g686 ( 
.A(n_580),
.B(n_300),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_SL g687 ( 
.A(n_529),
.B(n_302),
.Y(n_687)
);

AOI22xp5_ASAP7_75t_L g688 ( 
.A1(n_523),
.A2(n_217),
.B1(n_180),
.B2(n_184),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_L g689 ( 
.A(n_476),
.B(n_453),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_L g690 ( 
.A(n_479),
.B(n_453),
.Y(n_690)
);

NOR2xp33_ASAP7_75t_L g691 ( 
.A(n_552),
.B(n_191),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_479),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_L g693 ( 
.A(n_484),
.B(n_453),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_L g694 ( 
.A(n_484),
.B(n_453),
.Y(n_694)
);

INVx2_ASAP7_75t_L g695 ( 
.A(n_493),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_L g696 ( 
.A(n_493),
.B(n_498),
.Y(n_696)
);

NAND3xp33_ASAP7_75t_L g697 ( 
.A(n_514),
.B(n_218),
.C(n_194),
.Y(n_697)
);

INVx2_ASAP7_75t_L g698 ( 
.A(n_498),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_L g699 ( 
.A(n_512),
.B(n_453),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_SL g700 ( 
.A(n_529),
.B(n_461),
.Y(n_700)
);

NOR2xp33_ASAP7_75t_L g701 ( 
.A(n_610),
.B(n_203),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_512),
.Y(n_702)
);

INVx2_ASAP7_75t_L g703 ( 
.A(n_513),
.Y(n_703)
);

INVx2_ASAP7_75t_L g704 ( 
.A(n_513),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_SL g705 ( 
.A(n_529),
.B(n_453),
.Y(n_705)
);

INVx2_ASAP7_75t_L g706 ( 
.A(n_517),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_517),
.Y(n_707)
);

NOR3xp33_ASAP7_75t_L g708 ( 
.A(n_550),
.B(n_273),
.C(n_213),
.Y(n_708)
);

AND2x4_ASAP7_75t_L g709 ( 
.A(n_558),
.B(n_184),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_522),
.Y(n_710)
);

INVx2_ASAP7_75t_L g711 ( 
.A(n_522),
.Y(n_711)
);

INVx2_ASAP7_75t_SL g712 ( 
.A(n_568),
.Y(n_712)
);

INVx2_ASAP7_75t_L g713 ( 
.A(n_530),
.Y(n_713)
);

INVx2_ASAP7_75t_L g714 ( 
.A(n_530),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_L g715 ( 
.A(n_531),
.B(n_457),
.Y(n_715)
);

NOR2xp33_ASAP7_75t_L g716 ( 
.A(n_585),
.B(n_222),
.Y(n_716)
);

BUFx6f_ASAP7_75t_L g717 ( 
.A(n_468),
.Y(n_717)
);

BUFx3_ASAP7_75t_L g718 ( 
.A(n_558),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_L g719 ( 
.A(n_531),
.B(n_457),
.Y(n_719)
);

NAND2xp33_ASAP7_75t_L g720 ( 
.A(n_500),
.B(n_204),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_L g721 ( 
.A(n_536),
.B(n_457),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_L g722 ( 
.A(n_536),
.B(n_457),
.Y(n_722)
);

BUFx6f_ASAP7_75t_L g723 ( 
.A(n_468),
.Y(n_723)
);

NOR2xp33_ASAP7_75t_SL g724 ( 
.A(n_559),
.B(n_166),
.Y(n_724)
);

NAND2xp33_ASAP7_75t_L g725 ( 
.A(n_500),
.B(n_204),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_SL g726 ( 
.A(n_529),
.B(n_457),
.Y(n_726)
);

INVx6_ASAP7_75t_L g727 ( 
.A(n_558),
.Y(n_727)
);

INVx2_ASAP7_75t_SL g728 ( 
.A(n_576),
.Y(n_728)
);

HB1xp67_ASAP7_75t_L g729 ( 
.A(n_492),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_L g730 ( 
.A(n_548),
.B(n_457),
.Y(n_730)
);

INVxp67_ASAP7_75t_SL g731 ( 
.A(n_560),
.Y(n_731)
);

INVx2_ASAP7_75t_L g732 ( 
.A(n_548),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_L g733 ( 
.A(n_551),
.B(n_457),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_L g734 ( 
.A(n_551),
.B(n_457),
.Y(n_734)
);

INVx4_ASAP7_75t_L g735 ( 
.A(n_521),
.Y(n_735)
);

NOR2xp33_ASAP7_75t_L g736 ( 
.A(n_613),
.B(n_231),
.Y(n_736)
);

INVx2_ASAP7_75t_SL g737 ( 
.A(n_492),
.Y(n_737)
);

INVx3_ASAP7_75t_L g738 ( 
.A(n_521),
.Y(n_738)
);

BUFx5_ASAP7_75t_L g739 ( 
.A(n_500),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_591),
.Y(n_740)
);

NOR2xp33_ASAP7_75t_L g741 ( 
.A(n_546),
.B(n_232),
.Y(n_741)
);

AND2x4_ASAP7_75t_L g742 ( 
.A(n_592),
.B(n_209),
.Y(n_742)
);

NOR2xp67_ASAP7_75t_L g743 ( 
.A(n_509),
.B(n_454),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_L g744 ( 
.A(n_602),
.B(n_459),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_591),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_L g746 ( 
.A(n_611),
.B(n_459),
.Y(n_746)
);

AND2x2_ASAP7_75t_L g747 ( 
.A(n_533),
.B(n_166),
.Y(n_747)
);

OAI221xp5_ASAP7_75t_L g748 ( 
.A1(n_487),
.A2(n_266),
.B1(n_270),
.B2(n_294),
.C(n_287),
.Y(n_748)
);

INVx8_ASAP7_75t_L g749 ( 
.A(n_492),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_596),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_L g751 ( 
.A(n_515),
.B(n_459),
.Y(n_751)
);

INVx2_ASAP7_75t_L g752 ( 
.A(n_469),
.Y(n_752)
);

INVx2_ASAP7_75t_L g753 ( 
.A(n_469),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_L g754 ( 
.A(n_527),
.B(n_596),
.Y(n_754)
);

OAI22xp5_ASAP7_75t_L g755 ( 
.A1(n_553),
.A2(n_215),
.B1(n_220),
.B2(n_227),
.Y(n_755)
);

AND2x2_ASAP7_75t_L g756 ( 
.A(n_547),
.B(n_166),
.Y(n_756)
);

BUFx6f_ASAP7_75t_SL g757 ( 
.A(n_519),
.Y(n_757)
);

NOR2xp33_ASAP7_75t_L g758 ( 
.A(n_492),
.B(n_237),
.Y(n_758)
);

INVxp67_ASAP7_75t_L g759 ( 
.A(n_547),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_L g760 ( 
.A(n_603),
.B(n_459),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_L g761 ( 
.A(n_603),
.B(n_608),
.Y(n_761)
);

INVx2_ASAP7_75t_L g762 ( 
.A(n_470),
.Y(n_762)
);

AOI22xp33_ASAP7_75t_L g763 ( 
.A1(n_588),
.A2(n_266),
.B1(n_270),
.B2(n_287),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_L g764 ( 
.A(n_608),
.B(n_459),
.Y(n_764)
);

A2O1A1Ixp33_ASAP7_75t_L g765 ( 
.A1(n_609),
.A2(n_299),
.B(n_215),
.C(n_220),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_SL g766 ( 
.A(n_609),
.B(n_459),
.Y(n_766)
);

NOR2xp33_ASAP7_75t_L g767 ( 
.A(n_492),
.B(n_239),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_L g768 ( 
.A(n_526),
.B(n_459),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_597),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_L g770 ( 
.A(n_526),
.B(n_528),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_592),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_L g772 ( 
.A(n_526),
.B(n_459),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_592),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_SL g774 ( 
.A(n_528),
.B(n_461),
.Y(n_774)
);

INVx2_ASAP7_75t_L g775 ( 
.A(n_470),
.Y(n_775)
);

OAI22xp5_ASAP7_75t_L g776 ( 
.A1(n_592),
.A2(n_209),
.B1(n_228),
.B2(n_249),
.Y(n_776)
);

BUFx6f_ASAP7_75t_SL g777 ( 
.A(n_519),
.Y(n_777)
);

INVx1_ASAP7_75t_SL g778 ( 
.A(n_570),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_592),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_477),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_477),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_SL g782 ( 
.A(n_528),
.B(n_461),
.Y(n_782)
);

NOR2xp33_ASAP7_75t_L g783 ( 
.A(n_595),
.B(n_243),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_L g784 ( 
.A(n_505),
.B(n_461),
.Y(n_784)
);

INVx2_ASAP7_75t_L g785 ( 
.A(n_488),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_L g786 ( 
.A(n_505),
.B(n_461),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_624),
.Y(n_787)
);

AOI21xp5_ASAP7_75t_L g788 ( 
.A1(n_770),
.A2(n_593),
.B(n_589),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_L g789 ( 
.A(n_622),
.B(n_505),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_L g790 ( 
.A(n_769),
.B(n_646),
.Y(n_790)
);

NOR2xp33_ASAP7_75t_L g791 ( 
.A(n_759),
.B(n_598),
.Y(n_791)
);

AOI21xp5_ASAP7_75t_L g792 ( 
.A1(n_645),
.A2(n_593),
.B(n_589),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_L g793 ( 
.A(n_646),
.B(n_471),
.Y(n_793)
);

AOI21xp5_ASAP7_75t_L g794 ( 
.A1(n_751),
.A2(n_593),
.B(n_589),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_L g795 ( 
.A(n_620),
.B(n_471),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_624),
.Y(n_796)
);

OAI21xp33_ASAP7_75t_L g797 ( 
.A1(n_736),
.A2(n_615),
.B(n_253),
.Y(n_797)
);

OAI22xp5_ASAP7_75t_L g798 ( 
.A1(n_727),
.A2(n_737),
.B1(n_679),
.B2(n_718),
.Y(n_798)
);

INVx5_ASAP7_75t_L g799 ( 
.A(n_636),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_L g800 ( 
.A(n_637),
.B(n_471),
.Y(n_800)
);

AOI21xp5_ASAP7_75t_L g801 ( 
.A1(n_649),
.A2(n_589),
.B(n_502),
.Y(n_801)
);

AOI22xp33_ASAP7_75t_L g802 ( 
.A1(n_763),
.A2(n_588),
.B1(n_518),
.B2(n_500),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_SL g803 ( 
.A(n_739),
.B(n_471),
.Y(n_803)
);

O2A1O1Ixp33_ASAP7_75t_L g804 ( 
.A1(n_655),
.A2(n_267),
.B(n_290),
.C(n_299),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_L g805 ( 
.A(n_652),
.B(n_483),
.Y(n_805)
);

OAI21x1_ASAP7_75t_L g806 ( 
.A1(n_647),
.A2(n_483),
.B(n_496),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_L g807 ( 
.A(n_652),
.B(n_483),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_L g808 ( 
.A(n_625),
.B(n_496),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_SL g809 ( 
.A(n_739),
.B(n_496),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_L g810 ( 
.A(n_630),
.B(n_508),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_L g811 ( 
.A(n_648),
.B(n_508),
.Y(n_811)
);

AOI22xp5_ASAP7_75t_L g812 ( 
.A1(n_661),
.A2(n_500),
.B1(n_518),
.B2(n_516),
.Y(n_812)
);

CKINVDCx5p33_ASAP7_75t_R g813 ( 
.A(n_641),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_L g814 ( 
.A(n_650),
.B(n_508),
.Y(n_814)
);

BUFx8_ASAP7_75t_L g815 ( 
.A(n_757),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_L g816 ( 
.A(n_667),
.B(n_682),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_L g817 ( 
.A(n_692),
.B(n_508),
.Y(n_817)
);

INVx2_ASAP7_75t_L g818 ( 
.A(n_629),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_L g819 ( 
.A(n_702),
.B(n_707),
.Y(n_819)
);

AND2x2_ASAP7_75t_L g820 ( 
.A(n_639),
.B(n_519),
.Y(n_820)
);

INVx3_ASAP7_75t_L g821 ( 
.A(n_718),
.Y(n_821)
);

NOR2xp33_ASAP7_75t_L g822 ( 
.A(n_640),
.B(n_519),
.Y(n_822)
);

OAI21xp5_ASAP7_75t_L g823 ( 
.A1(n_616),
.A2(n_614),
.B(n_607),
.Y(n_823)
);

AOI21xp5_ASAP7_75t_L g824 ( 
.A1(n_651),
.A2(n_502),
.B(n_574),
.Y(n_824)
);

AO21x1_ASAP7_75t_L g825 ( 
.A1(n_676),
.A2(n_249),
.B(n_254),
.Y(n_825)
);

OAI21xp5_ASAP7_75t_L g826 ( 
.A1(n_674),
.A2(n_614),
.B(n_607),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_644),
.Y(n_827)
);

AO21x1_ASAP7_75t_L g828 ( 
.A1(n_688),
.A2(n_315),
.B(n_290),
.Y(n_828)
);

AOI21xp5_ASAP7_75t_L g829 ( 
.A1(n_666),
.A2(n_502),
.B(n_560),
.Y(n_829)
);

AOI21xp5_ASAP7_75t_L g830 ( 
.A1(n_669),
.A2(n_754),
.B(n_746),
.Y(n_830)
);

AND2x4_ASAP7_75t_L g831 ( 
.A(n_642),
.B(n_612),
.Y(n_831)
);

AOI21xp5_ASAP7_75t_L g832 ( 
.A1(n_744),
.A2(n_502),
.B(n_586),
.Y(n_832)
);

O2A1O1Ixp5_ASAP7_75t_L g833 ( 
.A1(n_686),
.A2(n_605),
.B(n_532),
.C(n_538),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_L g834 ( 
.A(n_710),
.B(n_643),
.Y(n_834)
);

INVx3_ASAP7_75t_L g835 ( 
.A(n_727),
.Y(n_835)
);

A2O1A1Ixp33_ASAP7_75t_L g836 ( 
.A1(n_758),
.A2(n_254),
.B(n_251),
.C(n_295),
.Y(n_836)
);

A2O1A1Ixp33_ASAP7_75t_L g837 ( 
.A1(n_758),
.A2(n_304),
.B(n_263),
.C(n_265),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_L g838 ( 
.A(n_696),
.B(n_532),
.Y(n_838)
);

NOR2xp33_ASAP7_75t_L g839 ( 
.A(n_736),
.B(n_639),
.Y(n_839)
);

AO21x1_ASAP7_75t_L g840 ( 
.A1(n_653),
.A2(n_686),
.B(n_618),
.Y(n_840)
);

A2O1A1Ixp33_ASAP7_75t_L g841 ( 
.A1(n_767),
.A2(n_306),
.B(n_271),
.C(n_272),
.Y(n_841)
);

OAI21xp5_ASAP7_75t_L g842 ( 
.A1(n_658),
.A2(n_488),
.B(n_604),
.Y(n_842)
);

OAI21xp5_ASAP7_75t_L g843 ( 
.A1(n_660),
.A2(n_490),
.B(n_604),
.Y(n_843)
);

INVx1_ASAP7_75t_SL g844 ( 
.A(n_633),
.Y(n_844)
);

OAI21xp5_ASAP7_75t_L g845 ( 
.A1(n_631),
.A2(n_490),
.B(n_601),
.Y(n_845)
);

NOR2xp33_ASAP7_75t_L g846 ( 
.A(n_621),
.B(n_549),
.Y(n_846)
);

AOI21xp5_ASAP7_75t_L g847 ( 
.A1(n_623),
.A2(n_560),
.B(n_574),
.Y(n_847)
);

AO21x1_ASAP7_75t_L g848 ( 
.A1(n_653),
.A2(n_449),
.B(n_594),
.Y(n_848)
);

BUFx2_ASAP7_75t_L g849 ( 
.A(n_778),
.Y(n_849)
);

AND2x2_ASAP7_75t_L g850 ( 
.A(n_673),
.B(n_549),
.Y(n_850)
);

AOI21xp5_ASAP7_75t_L g851 ( 
.A1(n_626),
.A2(n_560),
.B(n_574),
.Y(n_851)
);

INVx2_ASAP7_75t_L g852 ( 
.A(n_644),
.Y(n_852)
);

O2A1O1Ixp33_ASAP7_75t_SL g853 ( 
.A1(n_638),
.A2(n_578),
.B(n_601),
.C(n_600),
.Y(n_853)
);

AOI21xp5_ASAP7_75t_L g854 ( 
.A1(n_628),
.A2(n_560),
.B(n_574),
.Y(n_854)
);

OAI22xp5_ASAP7_75t_L g855 ( 
.A1(n_727),
.A2(n_588),
.B1(n_563),
.B2(n_538),
.Y(n_855)
);

AND2x2_ASAP7_75t_L g856 ( 
.A(n_747),
.B(n_549),
.Y(n_856)
);

OAI22xp5_ASAP7_75t_L g857 ( 
.A1(n_729),
.A2(n_588),
.B1(n_563),
.B2(n_538),
.Y(n_857)
);

AOI21xp5_ASAP7_75t_L g858 ( 
.A1(n_634),
.A2(n_574),
.B(n_586),
.Y(n_858)
);

OAI22xp5_ASAP7_75t_L g859 ( 
.A1(n_670),
.A2(n_563),
.B1(n_605),
.B2(n_532),
.Y(n_859)
);

INVx2_ASAP7_75t_L g860 ( 
.A(n_657),
.Y(n_860)
);

AOI21xp5_ASAP7_75t_L g861 ( 
.A1(n_683),
.A2(n_586),
.B(n_532),
.Y(n_861)
);

OAI21xp33_ASAP7_75t_L g862 ( 
.A1(n_716),
.A2(n_277),
.B(n_303),
.Y(n_862)
);

O2A1O1Ixp33_ASAP7_75t_L g863 ( 
.A1(n_748),
.A2(n_449),
.B(n_600),
.C(n_594),
.Y(n_863)
);

AOI21xp5_ASAP7_75t_L g864 ( 
.A1(n_684),
.A2(n_586),
.B(n_538),
.Y(n_864)
);

NOR2xp33_ASAP7_75t_SL g865 ( 
.A(n_757),
.B(n_549),
.Y(n_865)
);

NAND2x1_ASAP7_75t_L g866 ( 
.A(n_636),
.B(n_563),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_L g867 ( 
.A(n_657),
.B(n_564),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_L g868 ( 
.A(n_664),
.B(n_564),
.Y(n_868)
);

NAND2x1_ASAP7_75t_L g869 ( 
.A(n_636),
.B(n_564),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_664),
.Y(n_870)
);

NOR2xp33_ASAP7_75t_L g871 ( 
.A(n_697),
.B(n_256),
.Y(n_871)
);

AOI21x1_ASAP7_75t_L g872 ( 
.A1(n_774),
.A2(n_507),
.B(n_495),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_L g873 ( 
.A(n_665),
.B(n_564),
.Y(n_873)
);

AOI21xp33_ASAP7_75t_L g874 ( 
.A1(n_716),
.A2(n_308),
.B(n_309),
.Y(n_874)
);

OAI21xp33_ASAP7_75t_SL g875 ( 
.A1(n_665),
.A2(n_695),
.B(n_675),
.Y(n_875)
);

INVx1_ASAP7_75t_L g876 ( 
.A(n_675),
.Y(n_876)
);

BUFx4f_ASAP7_75t_L g877 ( 
.A(n_749),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_L g878 ( 
.A(n_695),
.B(n_569),
.Y(n_878)
);

AO21x2_ASAP7_75t_L g879 ( 
.A1(n_671),
.A2(n_555),
.B(n_503),
.Y(n_879)
);

INVx2_ASAP7_75t_L g880 ( 
.A(n_698),
.Y(n_880)
);

AND2x4_ASAP7_75t_L g881 ( 
.A(n_712),
.B(n_362),
.Y(n_881)
);

NOR2xp33_ASAP7_75t_SL g882 ( 
.A(n_777),
.B(n_274),
.Y(n_882)
);

INVx2_ASAP7_75t_L g883 ( 
.A(n_698),
.Y(n_883)
);

NOR2xp33_ASAP7_75t_SL g884 ( 
.A(n_777),
.B(n_735),
.Y(n_884)
);

INVx3_ASAP7_75t_L g885 ( 
.A(n_703),
.Y(n_885)
);

BUFx6f_ASAP7_75t_L g886 ( 
.A(n_636),
.Y(n_886)
);

HB1xp67_ASAP7_75t_L g887 ( 
.A(n_771),
.Y(n_887)
);

OAI22xp5_ASAP7_75t_L g888 ( 
.A1(n_619),
.A2(n_605),
.B1(n_569),
.B2(n_583),
.Y(n_888)
);

AOI21xp5_ASAP7_75t_L g889 ( 
.A1(n_731),
.A2(n_586),
.B(n_569),
.Y(n_889)
);

AOI21xp5_ASAP7_75t_L g890 ( 
.A1(n_768),
.A2(n_772),
.B(n_743),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_L g891 ( 
.A(n_703),
.B(n_569),
.Y(n_891)
);

INVx1_ASAP7_75t_L g892 ( 
.A(n_704),
.Y(n_892)
);

INVx3_ASAP7_75t_L g893 ( 
.A(n_704),
.Y(n_893)
);

INVx2_ASAP7_75t_L g894 ( 
.A(n_706),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_L g895 ( 
.A(n_706),
.B(n_583),
.Y(n_895)
);

NAND2xp5_ASAP7_75t_SL g896 ( 
.A(n_739),
.B(n_583),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_SL g897 ( 
.A(n_739),
.B(n_583),
.Y(n_897)
);

AOI21xp5_ASAP7_75t_L g898 ( 
.A1(n_700),
.A2(n_605),
.B(n_495),
.Y(n_898)
);

BUFx6f_ASAP7_75t_L g899 ( 
.A(n_717),
.Y(n_899)
);

NOR2xp33_ASAP7_75t_R g900 ( 
.A(n_685),
.B(n_680),
.Y(n_900)
);

INVx1_ASAP7_75t_L g901 ( 
.A(n_711),
.Y(n_901)
);

INVx1_ASAP7_75t_L g902 ( 
.A(n_711),
.Y(n_902)
);

OAI22xp5_ASAP7_75t_L g903 ( 
.A1(n_619),
.A2(n_510),
.B1(n_590),
.B2(n_584),
.Y(n_903)
);

INVx2_ASAP7_75t_L g904 ( 
.A(n_713),
.Y(n_904)
);

NOR3xp33_ASAP7_75t_L g905 ( 
.A(n_691),
.B(n_460),
.C(n_456),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_L g906 ( 
.A(n_713),
.B(n_500),
.Y(n_906)
);

AOI21xp5_ASAP7_75t_L g907 ( 
.A1(n_700),
.A2(n_510),
.B(n_590),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_SL g908 ( 
.A(n_739),
.B(n_728),
.Y(n_908)
);

BUFx2_ASAP7_75t_L g909 ( 
.A(n_617),
.Y(n_909)
);

AOI22x1_ASAP7_75t_L g910 ( 
.A1(n_714),
.A2(n_556),
.B1(n_581),
.B2(n_578),
.Y(n_910)
);

NAND2xp5_ASAP7_75t_L g911 ( 
.A(n_714),
.B(n_500),
.Y(n_911)
);

O2A1O1Ixp33_ASAP7_75t_SL g912 ( 
.A1(n_638),
.A2(n_503),
.B(n_575),
.C(n_571),
.Y(n_912)
);

AOI21xp5_ASAP7_75t_L g913 ( 
.A1(n_705),
.A2(n_556),
.B(n_581),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_L g914 ( 
.A(n_732),
.B(n_518),
.Y(n_914)
);

AND2x2_ASAP7_75t_L g915 ( 
.A(n_756),
.B(n_701),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_SL g916 ( 
.A(n_739),
.B(n_732),
.Y(n_916)
);

AOI21xp5_ASAP7_75t_L g917 ( 
.A1(n_705),
.A2(n_555),
.B(n_575),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_L g918 ( 
.A(n_709),
.B(n_518),
.Y(n_918)
);

NOR2xp33_ASAP7_75t_L g919 ( 
.A(n_691),
.B(n_524),
.Y(n_919)
);

AND2x2_ASAP7_75t_L g920 ( 
.A(n_701),
.B(n_274),
.Y(n_920)
);

NAND2xp5_ASAP7_75t_SL g921 ( 
.A(n_773),
.B(n_524),
.Y(n_921)
);

INVx2_ASAP7_75t_L g922 ( 
.A(n_752),
.Y(n_922)
);

AOI21xp5_ASAP7_75t_L g923 ( 
.A1(n_726),
.A2(n_571),
.B(n_562),
.Y(n_923)
);

NAND2xp5_ASAP7_75t_L g924 ( 
.A(n_709),
.B(n_518),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_L g925 ( 
.A(n_709),
.B(n_518),
.Y(n_925)
);

AOI21xp5_ASAP7_75t_L g926 ( 
.A1(n_726),
.A2(n_562),
.B(n_543),
.Y(n_926)
);

INVx2_ASAP7_75t_L g927 ( 
.A(n_752),
.Y(n_927)
);

AO21x1_ASAP7_75t_L g928 ( 
.A1(n_755),
.A2(n_426),
.B(n_460),
.Y(n_928)
);

OAI22xp5_ASAP7_75t_L g929 ( 
.A1(n_749),
.A2(n_454),
.B1(n_455),
.B2(n_456),
.Y(n_929)
);

HB1xp67_ASAP7_75t_L g930 ( 
.A(n_779),
.Y(n_930)
);

NAND2xp5_ASAP7_75t_L g931 ( 
.A(n_740),
.B(n_518),
.Y(n_931)
);

AOI21xp5_ASAP7_75t_L g932 ( 
.A1(n_774),
.A2(n_397),
.B(n_399),
.Y(n_932)
);

AOI21xp5_ASAP7_75t_L g933 ( 
.A1(n_782),
.A2(n_397),
.B(n_399),
.Y(n_933)
);

OAI21xp33_ASAP7_75t_L g934 ( 
.A1(n_656),
.A2(n_460),
.B(n_456),
.Y(n_934)
);

NAND2xp5_ASAP7_75t_L g935 ( 
.A(n_745),
.B(n_454),
.Y(n_935)
);

NOR2xp33_ASAP7_75t_R g936 ( 
.A(n_680),
.B(n_738),
.Y(n_936)
);

NAND2xp5_ASAP7_75t_L g937 ( 
.A(n_750),
.B(n_454),
.Y(n_937)
);

INVx2_ASAP7_75t_L g938 ( 
.A(n_753),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_SL g939 ( 
.A(n_738),
.B(n_461),
.Y(n_939)
);

INVx2_ASAP7_75t_L g940 ( 
.A(n_753),
.Y(n_940)
);

A2O1A1Ixp33_ASAP7_75t_L g941 ( 
.A1(n_767),
.A2(n_456),
.B(n_460),
.C(n_455),
.Y(n_941)
);

AOI21xp5_ASAP7_75t_L g942 ( 
.A1(n_782),
.A2(n_397),
.B(n_399),
.Y(n_942)
);

AND3x1_ASAP7_75t_SL g943 ( 
.A(n_724),
.B(n_274),
.C(n_284),
.Y(n_943)
);

NAND2xp5_ASAP7_75t_L g944 ( 
.A(n_668),
.B(n_455),
.Y(n_944)
);

OAI321xp33_ASAP7_75t_L g945 ( 
.A1(n_668),
.A2(n_741),
.A3(n_663),
.B1(n_763),
.B2(n_776),
.C(n_783),
.Y(n_945)
);

NAND2xp5_ASAP7_75t_L g946 ( 
.A(n_742),
.B(n_461),
.Y(n_946)
);

NOR2xp67_ASAP7_75t_L g947 ( 
.A(n_632),
.B(n_75),
.Y(n_947)
);

INVx2_ASAP7_75t_L g948 ( 
.A(n_762),
.Y(n_948)
);

AOI21xp5_ASAP7_75t_L g949 ( 
.A1(n_761),
.A2(n_399),
.B(n_426),
.Y(n_949)
);

NOR3xp33_ASAP7_75t_L g950 ( 
.A(n_741),
.B(n_439),
.C(n_436),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_L g951 ( 
.A(n_742),
.B(n_599),
.Y(n_951)
);

AOI21x1_ASAP7_75t_L g952 ( 
.A1(n_627),
.A2(n_439),
.B(n_436),
.Y(n_952)
);

NAND2xp5_ASAP7_75t_L g953 ( 
.A(n_742),
.B(n_599),
.Y(n_953)
);

OAI22xp5_ASAP7_75t_SL g954 ( 
.A1(n_783),
.A2(n_284),
.B1(n_274),
.B2(n_15),
.Y(n_954)
);

NAND2xp5_ASAP7_75t_SL g955 ( 
.A(n_717),
.B(n_431),
.Y(n_955)
);

OAI22xp5_ASAP7_75t_L g956 ( 
.A1(n_749),
.A2(n_681),
.B1(n_678),
.B2(n_717),
.Y(n_956)
);

AOI22xp5_ASAP7_75t_L g957 ( 
.A1(n_687),
.A2(n_599),
.B1(n_439),
.B2(n_436),
.Y(n_957)
);

INVx1_ASAP7_75t_L g958 ( 
.A(n_762),
.Y(n_958)
);

AOI22xp5_ASAP7_75t_L g959 ( 
.A1(n_687),
.A2(n_599),
.B1(n_439),
.B2(n_436),
.Y(n_959)
);

NAND2xp5_ASAP7_75t_L g960 ( 
.A(n_775),
.B(n_599),
.Y(n_960)
);

AOI21xp5_ASAP7_75t_L g961 ( 
.A1(n_784),
.A2(n_432),
.B(n_420),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_SL g962 ( 
.A(n_717),
.B(n_431),
.Y(n_962)
);

OAI21xp5_ASAP7_75t_L g963 ( 
.A1(n_662),
.A2(n_627),
.B(n_659),
.Y(n_963)
);

AOI21xp5_ASAP7_75t_L g964 ( 
.A1(n_786),
.A2(n_432),
.B(n_420),
.Y(n_964)
);

INVx1_ASAP7_75t_L g965 ( 
.A(n_775),
.Y(n_965)
);

AOI21xp5_ASAP7_75t_L g966 ( 
.A1(n_662),
.A2(n_432),
.B(n_420),
.Y(n_966)
);

OAI21xp5_ASAP7_75t_L g967 ( 
.A1(n_785),
.A2(n_599),
.B(n_432),
.Y(n_967)
);

NAND2xp5_ASAP7_75t_SL g968 ( 
.A(n_723),
.B(n_735),
.Y(n_968)
);

NAND2xp5_ASAP7_75t_L g969 ( 
.A(n_785),
.B(n_431),
.Y(n_969)
);

AOI21xp5_ASAP7_75t_L g970 ( 
.A1(n_723),
.A2(n_420),
.B(n_431),
.Y(n_970)
);

INVx2_ASAP7_75t_L g971 ( 
.A(n_780),
.Y(n_971)
);

AND2x2_ASAP7_75t_L g972 ( 
.A(n_635),
.B(n_284),
.Y(n_972)
);

BUFx2_ASAP7_75t_L g973 ( 
.A(n_765),
.Y(n_973)
);

INVx1_ASAP7_75t_L g974 ( 
.A(n_781),
.Y(n_974)
);

INVx1_ASAP7_75t_SL g975 ( 
.A(n_849),
.Y(n_975)
);

AOI21xp5_ASAP7_75t_L g976 ( 
.A1(n_830),
.A2(n_719),
.B(n_677),
.Y(n_976)
);

CKINVDCx5p33_ASAP7_75t_R g977 ( 
.A(n_813),
.Y(n_977)
);

O2A1O1Ixp33_ASAP7_75t_L g978 ( 
.A1(n_839),
.A2(n_722),
.B(n_672),
.C(n_689),
.Y(n_978)
);

INVx2_ASAP7_75t_L g979 ( 
.A(n_818),
.Y(n_979)
);

HB1xp67_ASAP7_75t_L g980 ( 
.A(n_844),
.Y(n_980)
);

A2O1A1Ixp33_ASAP7_75t_L g981 ( 
.A1(n_839),
.A2(n_694),
.B(n_699),
.C(n_693),
.Y(n_981)
);

INVx3_ASAP7_75t_SL g982 ( 
.A(n_831),
.Y(n_982)
);

AOI21xp5_ASAP7_75t_L g983 ( 
.A1(n_793),
.A2(n_730),
.B(n_721),
.Y(n_983)
);

A2O1A1Ixp33_ASAP7_75t_SL g984 ( 
.A1(n_871),
.A2(n_919),
.B(n_791),
.C(n_945),
.Y(n_984)
);

AOI21xp5_ASAP7_75t_L g985 ( 
.A1(n_944),
.A2(n_715),
.B(n_734),
.Y(n_985)
);

AOI21xp5_ASAP7_75t_L g986 ( 
.A1(n_792),
.A2(n_733),
.B(n_690),
.Y(n_986)
);

INVx6_ASAP7_75t_L g987 ( 
.A(n_815),
.Y(n_987)
);

A2O1A1Ixp33_ASAP7_75t_L g988 ( 
.A1(n_790),
.A2(n_708),
.B(n_764),
.C(n_760),
.Y(n_988)
);

AOI22xp5_ASAP7_75t_L g989 ( 
.A1(n_915),
.A2(n_723),
.B1(n_725),
.B2(n_720),
.Y(n_989)
);

AOI21xp5_ASAP7_75t_L g990 ( 
.A1(n_789),
.A2(n_723),
.B(n_766),
.Y(n_990)
);

OAI22xp5_ASAP7_75t_L g991 ( 
.A1(n_834),
.A2(n_681),
.B1(n_678),
.B2(n_654),
.Y(n_991)
);

AOI21xp5_ASAP7_75t_L g992 ( 
.A1(n_794),
.A2(n_766),
.B(n_420),
.Y(n_992)
);

NAND2xp5_ASAP7_75t_L g993 ( 
.A(n_820),
.B(n_431),
.Y(n_993)
);

AOI21xp5_ASAP7_75t_L g994 ( 
.A1(n_890),
.A2(n_420),
.B(n_431),
.Y(n_994)
);

OAI21xp5_ASAP7_75t_L g995 ( 
.A1(n_875),
.A2(n_345),
.B(n_431),
.Y(n_995)
);

NAND2xp5_ASAP7_75t_L g996 ( 
.A(n_816),
.B(n_431),
.Y(n_996)
);

INVx1_ASAP7_75t_L g997 ( 
.A(n_852),
.Y(n_997)
);

OAI21x1_ASAP7_75t_L g998 ( 
.A1(n_872),
.A2(n_100),
.B(n_152),
.Y(n_998)
);

OR2x6_ASAP7_75t_L g999 ( 
.A(n_850),
.B(n_284),
.Y(n_999)
);

INVx2_ASAP7_75t_L g1000 ( 
.A(n_852),
.Y(n_1000)
);

NAND2xp5_ASAP7_75t_SL g1001 ( 
.A(n_856),
.B(n_345),
.Y(n_1001)
);

A2O1A1Ixp33_ASAP7_75t_L g1002 ( 
.A1(n_791),
.A2(n_7),
.B(n_13),
.C(n_15),
.Y(n_1002)
);

AOI21xp5_ASAP7_75t_L g1003 ( 
.A1(n_832),
.A2(n_345),
.B(n_146),
.Y(n_1003)
);

AOI21xp5_ASAP7_75t_L g1004 ( 
.A1(n_829),
.A2(n_345),
.B(n_143),
.Y(n_1004)
);

NAND2x1p5_ASAP7_75t_L g1005 ( 
.A(n_799),
.B(n_140),
.Y(n_1005)
);

INVx1_ASAP7_75t_L g1006 ( 
.A(n_860),
.Y(n_1006)
);

AOI21xp5_ASAP7_75t_L g1007 ( 
.A1(n_847),
.A2(n_854),
.B(n_851),
.Y(n_1007)
);

INVx2_ASAP7_75t_L g1008 ( 
.A(n_860),
.Y(n_1008)
);

BUFx2_ASAP7_75t_L g1009 ( 
.A(n_831),
.Y(n_1009)
);

NOR2xp33_ASAP7_75t_L g1010 ( 
.A(n_909),
.B(n_13),
.Y(n_1010)
);

AOI21xp5_ASAP7_75t_L g1011 ( 
.A1(n_919),
.A2(n_128),
.B(n_124),
.Y(n_1011)
);

INVx1_ASAP7_75t_L g1012 ( 
.A(n_880),
.Y(n_1012)
);

INVx2_ASAP7_75t_L g1013 ( 
.A(n_880),
.Y(n_1013)
);

NAND2xp5_ASAP7_75t_SL g1014 ( 
.A(n_821),
.B(n_122),
.Y(n_1014)
);

OR2x2_ASAP7_75t_L g1015 ( 
.A(n_920),
.B(n_16),
.Y(n_1015)
);

NOR2xp33_ASAP7_75t_L g1016 ( 
.A(n_822),
.B(n_22),
.Y(n_1016)
);

INVx1_ASAP7_75t_L g1017 ( 
.A(n_883),
.Y(n_1017)
);

BUFx2_ASAP7_75t_SL g1018 ( 
.A(n_799),
.Y(n_1018)
);

AOI21xp5_ASAP7_75t_L g1019 ( 
.A1(n_858),
.A2(n_88),
.B(n_96),
.Y(n_1019)
);

INVx2_ASAP7_75t_L g1020 ( 
.A(n_883),
.Y(n_1020)
);

HB1xp67_ASAP7_75t_L g1021 ( 
.A(n_887),
.Y(n_1021)
);

INVx1_ASAP7_75t_L g1022 ( 
.A(n_787),
.Y(n_1022)
);

OAI22xp5_ASAP7_75t_L g1023 ( 
.A1(n_956),
.A2(n_108),
.B1(n_95),
.B2(n_92),
.Y(n_1023)
);

HB1xp67_ASAP7_75t_L g1024 ( 
.A(n_887),
.Y(n_1024)
);

A2O1A1Ixp33_ASAP7_75t_L g1025 ( 
.A1(n_871),
.A2(n_23),
.B(n_24),
.C(n_26),
.Y(n_1025)
);

OAI21xp33_ASAP7_75t_L g1026 ( 
.A1(n_874),
.A2(n_26),
.B(n_27),
.Y(n_1026)
);

AOI21xp5_ASAP7_75t_L g1027 ( 
.A1(n_824),
.A2(n_86),
.B(n_83),
.Y(n_1027)
);

AOI21xp5_ASAP7_75t_L g1028 ( 
.A1(n_838),
.A2(n_82),
.B(n_80),
.Y(n_1028)
);

AOI21xp5_ASAP7_75t_L g1029 ( 
.A1(n_788),
.A2(n_28),
.B(n_30),
.Y(n_1029)
);

NAND2xp5_ASAP7_75t_L g1030 ( 
.A(n_819),
.B(n_885),
.Y(n_1030)
);

INVx1_ASAP7_75t_L g1031 ( 
.A(n_796),
.Y(n_1031)
);

INVx2_ASAP7_75t_L g1032 ( 
.A(n_885),
.Y(n_1032)
);

NOR2xp33_ASAP7_75t_SL g1033 ( 
.A(n_865),
.B(n_30),
.Y(n_1033)
);

AOI21xp5_ASAP7_75t_L g1034 ( 
.A1(n_801),
.A2(n_31),
.B(n_33),
.Y(n_1034)
);

NAND2xp5_ASAP7_75t_L g1035 ( 
.A(n_893),
.B(n_31),
.Y(n_1035)
);

AOI22xp33_ASAP7_75t_L g1036 ( 
.A1(n_797),
.A2(n_34),
.B1(n_35),
.B2(n_36),
.Y(n_1036)
);

NAND2xp5_ASAP7_75t_L g1037 ( 
.A(n_893),
.B(n_37),
.Y(n_1037)
);

AOI22xp5_ASAP7_75t_L g1038 ( 
.A1(n_972),
.A2(n_59),
.B1(n_38),
.B2(n_39),
.Y(n_1038)
);

A2O1A1Ixp33_ASAP7_75t_L g1039 ( 
.A1(n_836),
.A2(n_37),
.B(n_38),
.C(n_39),
.Y(n_1039)
);

BUFx8_ASAP7_75t_L g1040 ( 
.A(n_881),
.Y(n_1040)
);

OAI22xp5_ASAP7_75t_L g1041 ( 
.A1(n_802),
.A2(n_41),
.B1(n_42),
.B2(n_43),
.Y(n_1041)
);

AOI21xp5_ASAP7_75t_L g1042 ( 
.A1(n_840),
.A2(n_41),
.B(n_44),
.Y(n_1042)
);

INVx2_ASAP7_75t_L g1043 ( 
.A(n_940),
.Y(n_1043)
);

NAND2xp5_ASAP7_75t_SL g1044 ( 
.A(n_821),
.B(n_47),
.Y(n_1044)
);

NOR2xp67_ASAP7_75t_SL g1045 ( 
.A(n_799),
.B(n_50),
.Y(n_1045)
);

NAND2xp5_ASAP7_75t_L g1046 ( 
.A(n_827),
.B(n_57),
.Y(n_1046)
);

AND2x2_ASAP7_75t_L g1047 ( 
.A(n_881),
.B(n_54),
.Y(n_1047)
);

OAI22xp5_ASAP7_75t_L g1048 ( 
.A1(n_802),
.A2(n_55),
.B1(n_57),
.B2(n_877),
.Y(n_1048)
);

INVx2_ASAP7_75t_L g1049 ( 
.A(n_940),
.Y(n_1049)
);

NAND2xp5_ASAP7_75t_SL g1050 ( 
.A(n_846),
.B(n_55),
.Y(n_1050)
);

NOR2xp33_ASAP7_75t_L g1051 ( 
.A(n_822),
.B(n_846),
.Y(n_1051)
);

INVx4_ASAP7_75t_L g1052 ( 
.A(n_799),
.Y(n_1052)
);

OAI21xp33_ASAP7_75t_L g1053 ( 
.A1(n_862),
.A2(n_882),
.B(n_836),
.Y(n_1053)
);

OAI22xp5_ASAP7_75t_L g1054 ( 
.A1(n_877),
.A2(n_902),
.B1(n_901),
.B2(n_892),
.Y(n_1054)
);

AOI21xp33_ASAP7_75t_L g1055 ( 
.A1(n_837),
.A2(n_841),
.B(n_798),
.Y(n_1055)
);

BUFx6f_ASAP7_75t_L g1056 ( 
.A(n_886),
.Y(n_1056)
);

NAND2xp5_ASAP7_75t_L g1057 ( 
.A(n_870),
.B(n_876),
.Y(n_1057)
);

NAND2xp5_ASAP7_75t_L g1058 ( 
.A(n_894),
.B(n_904),
.Y(n_1058)
);

NOR2xp33_ASAP7_75t_SL g1059 ( 
.A(n_884),
.B(n_815),
.Y(n_1059)
);

INVx3_ASAP7_75t_SL g1060 ( 
.A(n_886),
.Y(n_1060)
);

NAND2x1_ASAP7_75t_L g1061 ( 
.A(n_886),
.B(n_899),
.Y(n_1061)
);

NAND2xp5_ASAP7_75t_L g1062 ( 
.A(n_837),
.B(n_841),
.Y(n_1062)
);

INVx1_ASAP7_75t_L g1063 ( 
.A(n_971),
.Y(n_1063)
);

HB1xp67_ASAP7_75t_L g1064 ( 
.A(n_930),
.Y(n_1064)
);

OAI22xp5_ASAP7_75t_L g1065 ( 
.A1(n_855),
.A2(n_857),
.B1(n_800),
.B2(n_835),
.Y(n_1065)
);

NAND2x1p5_ASAP7_75t_L g1066 ( 
.A(n_886),
.B(n_899),
.Y(n_1066)
);

BUFx3_ASAP7_75t_L g1067 ( 
.A(n_930),
.Y(n_1067)
);

INVx2_ASAP7_75t_L g1068 ( 
.A(n_948),
.Y(n_1068)
);

INVx1_ASAP7_75t_L g1069 ( 
.A(n_971),
.Y(n_1069)
);

O2A1O1Ixp5_ASAP7_75t_SL g1070 ( 
.A1(n_921),
.A2(n_939),
.B(n_968),
.C(n_955),
.Y(n_1070)
);

NAND2xp5_ASAP7_75t_L g1071 ( 
.A(n_974),
.B(n_835),
.Y(n_1071)
);

BUFx2_ASAP7_75t_L g1072 ( 
.A(n_900),
.Y(n_1072)
);

NAND2xp5_ASAP7_75t_SL g1073 ( 
.A(n_936),
.B(n_812),
.Y(n_1073)
);

NAND2xp5_ASAP7_75t_L g1074 ( 
.A(n_948),
.B(n_922),
.Y(n_1074)
);

AOI21xp5_ASAP7_75t_L g1075 ( 
.A1(n_845),
.A2(n_963),
.B(n_795),
.Y(n_1075)
);

NAND2xp5_ASAP7_75t_L g1076 ( 
.A(n_927),
.B(n_938),
.Y(n_1076)
);

INVx2_ASAP7_75t_L g1077 ( 
.A(n_958),
.Y(n_1077)
);

INVx2_ASAP7_75t_SL g1078 ( 
.A(n_900),
.Y(n_1078)
);

NAND3xp33_ASAP7_75t_L g1079 ( 
.A(n_804),
.B(n_947),
.C(n_905),
.Y(n_1079)
);

NAND2xp5_ASAP7_75t_L g1080 ( 
.A(n_965),
.B(n_973),
.Y(n_1080)
);

NOR2xp33_ASAP7_75t_L g1081 ( 
.A(n_954),
.B(n_908),
.Y(n_1081)
);

NAND2xp5_ASAP7_75t_L g1082 ( 
.A(n_899),
.B(n_808),
.Y(n_1082)
);

HB1xp67_ASAP7_75t_L g1083 ( 
.A(n_936),
.Y(n_1083)
);

INVx1_ASAP7_75t_SL g1084 ( 
.A(n_899),
.Y(n_1084)
);

OA21x2_ASAP7_75t_L g1085 ( 
.A1(n_848),
.A2(n_941),
.B(n_806),
.Y(n_1085)
);

NAND2xp5_ASAP7_75t_L g1086 ( 
.A(n_810),
.B(n_811),
.Y(n_1086)
);

INVx1_ASAP7_75t_L g1087 ( 
.A(n_935),
.Y(n_1087)
);

INVx2_ASAP7_75t_L g1088 ( 
.A(n_910),
.Y(n_1088)
);

AOI22xp5_ASAP7_75t_L g1089 ( 
.A1(n_918),
.A2(n_925),
.B1(n_924),
.B2(n_908),
.Y(n_1089)
);

OAI22xp5_ASAP7_75t_L g1090 ( 
.A1(n_916),
.A2(n_946),
.B1(n_817),
.B2(n_814),
.Y(n_1090)
);

O2A1O1Ixp33_ASAP7_75t_L g1091 ( 
.A1(n_941),
.A2(n_921),
.B(n_937),
.C(n_929),
.Y(n_1091)
);

AND2x2_ASAP7_75t_L g1092 ( 
.A(n_950),
.B(n_825),
.Y(n_1092)
);

NAND2xp5_ASAP7_75t_L g1093 ( 
.A(n_867),
.B(n_868),
.Y(n_1093)
);

AO21x1_ASAP7_75t_L g1094 ( 
.A1(n_916),
.A2(n_939),
.B(n_859),
.Y(n_1094)
);

AND2x6_ASAP7_75t_L g1095 ( 
.A(n_951),
.B(n_953),
.Y(n_1095)
);

INVx4_ASAP7_75t_L g1096 ( 
.A(n_879),
.Y(n_1096)
);

INVx2_ASAP7_75t_L g1097 ( 
.A(n_873),
.Y(n_1097)
);

INVx3_ASAP7_75t_L g1098 ( 
.A(n_866),
.Y(n_1098)
);

AO21x1_ASAP7_75t_L g1099 ( 
.A1(n_968),
.A2(n_823),
.B(n_903),
.Y(n_1099)
);

NAND2xp5_ASAP7_75t_L g1100 ( 
.A(n_878),
.B(n_891),
.Y(n_1100)
);

AOI21xp5_ASAP7_75t_L g1101 ( 
.A1(n_842),
.A2(n_843),
.B(n_861),
.Y(n_1101)
);

NOR3xp33_ASAP7_75t_SL g1102 ( 
.A(n_943),
.B(n_888),
.C(n_934),
.Y(n_1102)
);

OR2x6_ASAP7_75t_L g1103 ( 
.A(n_906),
.B(n_914),
.Y(n_1103)
);

NAND2xp5_ASAP7_75t_L g1104 ( 
.A(n_895),
.B(n_805),
.Y(n_1104)
);

NOR3xp33_ASAP7_75t_SL g1105 ( 
.A(n_943),
.B(n_955),
.C(n_962),
.Y(n_1105)
);

OAI22xp5_ASAP7_75t_L g1106 ( 
.A1(n_807),
.A2(n_931),
.B1(n_911),
.B2(n_809),
.Y(n_1106)
);

NAND2xp5_ASAP7_75t_L g1107 ( 
.A(n_879),
.B(n_864),
.Y(n_1107)
);

INVx1_ASAP7_75t_SL g1108 ( 
.A(n_962),
.Y(n_1108)
);

BUFx6f_ASAP7_75t_L g1109 ( 
.A(n_869),
.Y(n_1109)
);

AND2x2_ASAP7_75t_L g1110 ( 
.A(n_957),
.B(n_959),
.Y(n_1110)
);

AOI21xp5_ASAP7_75t_L g1111 ( 
.A1(n_833),
.A2(n_889),
.B(n_969),
.Y(n_1111)
);

CKINVDCx16_ASAP7_75t_R g1112 ( 
.A(n_826),
.Y(n_1112)
);

AOI21xp5_ASAP7_75t_L g1113 ( 
.A1(n_853),
.A2(n_912),
.B(n_809),
.Y(n_1113)
);

CKINVDCx5p33_ASAP7_75t_R g1114 ( 
.A(n_970),
.Y(n_1114)
);

INVx2_ASAP7_75t_L g1115 ( 
.A(n_952),
.Y(n_1115)
);

INVx1_ASAP7_75t_L g1116 ( 
.A(n_863),
.Y(n_1116)
);

AO21x1_ASAP7_75t_L g1117 ( 
.A1(n_803),
.A2(n_897),
.B(n_896),
.Y(n_1117)
);

NAND2xp5_ASAP7_75t_L g1118 ( 
.A(n_907),
.B(n_917),
.Y(n_1118)
);

INVx2_ASAP7_75t_SL g1119 ( 
.A(n_803),
.Y(n_1119)
);

HB1xp67_ASAP7_75t_L g1120 ( 
.A(n_828),
.Y(n_1120)
);

BUFx2_ASAP7_75t_L g1121 ( 
.A(n_928),
.Y(n_1121)
);

BUFx3_ASAP7_75t_L g1122 ( 
.A(n_960),
.Y(n_1122)
);

OAI21xp5_ASAP7_75t_L g1123 ( 
.A1(n_913),
.A2(n_923),
.B(n_926),
.Y(n_1123)
);

OAI22xp5_ASAP7_75t_L g1124 ( 
.A1(n_896),
.A2(n_898),
.B1(n_967),
.B2(n_949),
.Y(n_1124)
);

AOI21xp5_ASAP7_75t_L g1125 ( 
.A1(n_853),
.A2(n_912),
.B(n_961),
.Y(n_1125)
);

AOI21xp5_ASAP7_75t_L g1126 ( 
.A1(n_964),
.A2(n_966),
.B(n_933),
.Y(n_1126)
);

AOI221xp5_ASAP7_75t_L g1127 ( 
.A1(n_1010),
.A2(n_932),
.B1(n_942),
.B2(n_984),
.C(n_1026),
.Y(n_1127)
);

NAND2xp5_ASAP7_75t_L g1128 ( 
.A(n_1051),
.B(n_1081),
.Y(n_1128)
);

AOI21xp5_ASAP7_75t_L g1129 ( 
.A1(n_1101),
.A2(n_1075),
.B(n_976),
.Y(n_1129)
);

INVx1_ASAP7_75t_L g1130 ( 
.A(n_1063),
.Y(n_1130)
);

AO31x2_ASAP7_75t_L g1131 ( 
.A1(n_1096),
.A2(n_1099),
.A3(n_1121),
.B(n_1094),
.Y(n_1131)
);

AOI22xp5_ASAP7_75t_L g1132 ( 
.A1(n_1016),
.A2(n_1050),
.B1(n_1053),
.B2(n_1038),
.Y(n_1132)
);

NAND2xp5_ASAP7_75t_L g1133 ( 
.A(n_1087),
.B(n_1030),
.Y(n_1133)
);

OAI21x1_ASAP7_75t_L g1134 ( 
.A1(n_994),
.A2(n_1007),
.B(n_1126),
.Y(n_1134)
);

INVx3_ASAP7_75t_L g1135 ( 
.A(n_1052),
.Y(n_1135)
);

INVx2_ASAP7_75t_SL g1136 ( 
.A(n_980),
.Y(n_1136)
);

INVxp67_ASAP7_75t_L g1137 ( 
.A(n_975),
.Y(n_1137)
);

NAND2xp5_ASAP7_75t_L g1138 ( 
.A(n_1097),
.B(n_1112),
.Y(n_1138)
);

NAND2xp5_ASAP7_75t_L g1139 ( 
.A(n_1080),
.B(n_1015),
.Y(n_1139)
);

INVx2_ASAP7_75t_L g1140 ( 
.A(n_979),
.Y(n_1140)
);

BUFx10_ASAP7_75t_L g1141 ( 
.A(n_977),
.Y(n_1141)
);

NOR2xp33_ASAP7_75t_L g1142 ( 
.A(n_1067),
.B(n_982),
.Y(n_1142)
);

OAI21xp5_ASAP7_75t_L g1143 ( 
.A1(n_1062),
.A2(n_988),
.B(n_1079),
.Y(n_1143)
);

O2A1O1Ixp33_ASAP7_75t_SL g1144 ( 
.A1(n_1039),
.A2(n_1055),
.B(n_1073),
.C(n_1014),
.Y(n_1144)
);

INVx1_ASAP7_75t_L g1145 ( 
.A(n_1069),
.Y(n_1145)
);

NOR2xp33_ASAP7_75t_L g1146 ( 
.A(n_982),
.B(n_1009),
.Y(n_1146)
);

NOR2xp33_ASAP7_75t_L g1147 ( 
.A(n_1021),
.B(n_1024),
.Y(n_1147)
);

AOI21xp5_ASAP7_75t_L g1148 ( 
.A1(n_1101),
.A2(n_976),
.B(n_1007),
.Y(n_1148)
);

OAI21xp5_ASAP7_75t_L g1149 ( 
.A1(n_981),
.A2(n_985),
.B(n_1091),
.Y(n_1149)
);

BUFx6f_ASAP7_75t_L g1150 ( 
.A(n_1060),
.Y(n_1150)
);

CKINVDCx5p33_ASAP7_75t_R g1151 ( 
.A(n_1072),
.Y(n_1151)
);

NAND2xp5_ASAP7_75t_L g1152 ( 
.A(n_991),
.B(n_1047),
.Y(n_1152)
);

BUFx3_ASAP7_75t_L g1153 ( 
.A(n_987),
.Y(n_1153)
);

OAI22x1_ASAP7_75t_L g1154 ( 
.A1(n_1044),
.A2(n_1064),
.B1(n_1120),
.B2(n_1001),
.Y(n_1154)
);

OAI22xp5_ASAP7_75t_L g1155 ( 
.A1(n_1065),
.A2(n_1114),
.B1(n_1054),
.B2(n_1071),
.Y(n_1155)
);

OA21x2_ASAP7_75t_L g1156 ( 
.A1(n_1107),
.A2(n_1125),
.B(n_1111),
.Y(n_1156)
);

A2O1A1Ixp33_ASAP7_75t_L g1157 ( 
.A1(n_1102),
.A2(n_1042),
.B(n_1105),
.C(n_1092),
.Y(n_1157)
);

AOI21xp5_ASAP7_75t_L g1158 ( 
.A1(n_985),
.A2(n_983),
.B(n_1111),
.Y(n_1158)
);

NOR2xp33_ASAP7_75t_L g1159 ( 
.A(n_1083),
.B(n_1078),
.Y(n_1159)
);

INVx1_ASAP7_75t_L g1160 ( 
.A(n_1022),
.Y(n_1160)
);

AND2x4_ASAP7_75t_L g1161 ( 
.A(n_1032),
.B(n_1031),
.Y(n_1161)
);

AOI21xp5_ASAP7_75t_SL g1162 ( 
.A1(n_1023),
.A2(n_978),
.B(n_1052),
.Y(n_1162)
);

BUFx6f_ASAP7_75t_L g1163 ( 
.A(n_1060),
.Y(n_1163)
);

O2A1O1Ixp5_ASAP7_75t_L g1164 ( 
.A1(n_1042),
.A2(n_1003),
.B(n_1004),
.C(n_1034),
.Y(n_1164)
);

OAI21xp5_ASAP7_75t_L g1165 ( 
.A1(n_1091),
.A2(n_1070),
.B(n_983),
.Y(n_1165)
);

AND2x2_ASAP7_75t_L g1166 ( 
.A(n_999),
.B(n_1033),
.Y(n_1166)
);

AO31x2_ASAP7_75t_L g1167 ( 
.A1(n_1096),
.A2(n_1125),
.A3(n_1124),
.B(n_1113),
.Y(n_1167)
);

BUFx2_ASAP7_75t_L g1168 ( 
.A(n_1040),
.Y(n_1168)
);

AOI21xp5_ASAP7_75t_L g1169 ( 
.A1(n_993),
.A2(n_986),
.B(n_1086),
.Y(n_1169)
);

AOI21xp5_ASAP7_75t_L g1170 ( 
.A1(n_986),
.A2(n_1118),
.B(n_1093),
.Y(n_1170)
);

NOR2xp33_ASAP7_75t_L g1171 ( 
.A(n_999),
.B(n_1040),
.Y(n_1171)
);

NOR2xp33_ASAP7_75t_L g1172 ( 
.A(n_999),
.B(n_1059),
.Y(n_1172)
);

AO31x2_ASAP7_75t_L g1173 ( 
.A1(n_1113),
.A2(n_1117),
.A3(n_1090),
.B(n_1126),
.Y(n_1173)
);

NAND3xp33_ASAP7_75t_L g1174 ( 
.A(n_1036),
.B(n_1025),
.C(n_1002),
.Y(n_1174)
);

AOI21xp5_ASAP7_75t_L g1175 ( 
.A1(n_1100),
.A2(n_1104),
.B(n_978),
.Y(n_1175)
);

O2A1O1Ixp33_ASAP7_75t_SL g1176 ( 
.A1(n_1048),
.A2(n_1041),
.B(n_1119),
.C(n_1035),
.Y(n_1176)
);

AO21x1_ASAP7_75t_L g1177 ( 
.A1(n_1029),
.A2(n_1034),
.B(n_1011),
.Y(n_1177)
);

AOI21xp5_ASAP7_75t_L g1178 ( 
.A1(n_1123),
.A2(n_990),
.B(n_1116),
.Y(n_1178)
);

AO32x2_ASAP7_75t_L g1179 ( 
.A1(n_1106),
.A2(n_1085),
.A3(n_1102),
.B1(n_1029),
.B2(n_1045),
.Y(n_1179)
);

INVxp33_ASAP7_75t_L g1180 ( 
.A(n_1046),
.Y(n_1180)
);

AOI21xp5_ASAP7_75t_L g1181 ( 
.A1(n_990),
.A2(n_996),
.B(n_1003),
.Y(n_1181)
);

AOI21xp5_ASAP7_75t_L g1182 ( 
.A1(n_1004),
.A2(n_992),
.B(n_1110),
.Y(n_1182)
);

NAND2x1p5_ASAP7_75t_L g1183 ( 
.A(n_1056),
.B(n_1061),
.Y(n_1183)
);

AOI21xp5_ASAP7_75t_L g1184 ( 
.A1(n_992),
.A2(n_1082),
.B(n_994),
.Y(n_1184)
);

AND2x4_ASAP7_75t_L g1185 ( 
.A(n_1077),
.B(n_1084),
.Y(n_1185)
);

AOI21xp5_ASAP7_75t_L g1186 ( 
.A1(n_995),
.A2(n_1027),
.B(n_1057),
.Y(n_1186)
);

AOI21xp5_ASAP7_75t_L g1187 ( 
.A1(n_1027),
.A2(n_989),
.B(n_1019),
.Y(n_1187)
);

INVx1_ASAP7_75t_L g1188 ( 
.A(n_997),
.Y(n_1188)
);

NAND2xp5_ASAP7_75t_L g1189 ( 
.A(n_1000),
.B(n_1020),
.Y(n_1189)
);

OAI21xp5_ASAP7_75t_L g1190 ( 
.A1(n_1089),
.A2(n_1037),
.B(n_1058),
.Y(n_1190)
);

NAND2xp5_ASAP7_75t_L g1191 ( 
.A(n_1008),
.B(n_1013),
.Y(n_1191)
);

AO31x2_ASAP7_75t_L g1192 ( 
.A1(n_1088),
.A2(n_1115),
.A3(n_1019),
.B(n_1011),
.Y(n_1192)
);

AO31x2_ASAP7_75t_L g1193 ( 
.A1(n_1028),
.A2(n_1012),
.A3(n_1017),
.B(n_1006),
.Y(n_1193)
);

NAND2xp5_ASAP7_75t_L g1194 ( 
.A(n_1122),
.B(n_1068),
.Y(n_1194)
);

AOI21xp5_ASAP7_75t_L g1195 ( 
.A1(n_1103),
.A2(n_1074),
.B(n_1085),
.Y(n_1195)
);

AOI22xp33_ASAP7_75t_L g1196 ( 
.A1(n_1095),
.A2(n_1103),
.B1(n_1108),
.B2(n_1049),
.Y(n_1196)
);

INVx1_ASAP7_75t_L g1197 ( 
.A(n_1043),
.Y(n_1197)
);

NAND2xp5_ASAP7_75t_L g1198 ( 
.A(n_1095),
.B(n_1076),
.Y(n_1198)
);

CKINVDCx6p67_ASAP7_75t_R g1199 ( 
.A(n_1056),
.Y(n_1199)
);

NOR2xp67_ASAP7_75t_L g1200 ( 
.A(n_1098),
.B(n_1109),
.Y(n_1200)
);

A2O1A1Ixp33_ASAP7_75t_L g1201 ( 
.A1(n_1028),
.A2(n_1098),
.B(n_998),
.C(n_1109),
.Y(n_1201)
);

NOR2xp33_ASAP7_75t_L g1202 ( 
.A(n_1056),
.B(n_987),
.Y(n_1202)
);

CKINVDCx11_ASAP7_75t_R g1203 ( 
.A(n_987),
.Y(n_1203)
);

NAND3xp33_ASAP7_75t_L g1204 ( 
.A(n_1103),
.B(n_1109),
.C(n_1095),
.Y(n_1204)
);

AOI21xp5_ASAP7_75t_L g1205 ( 
.A1(n_1066),
.A2(n_1018),
.B(n_1005),
.Y(n_1205)
);

A2O1A1Ixp33_ASAP7_75t_L g1206 ( 
.A1(n_1095),
.A2(n_1005),
.B(n_1066),
.C(n_839),
.Y(n_1206)
);

OAI22xp5_ASAP7_75t_L g1207 ( 
.A1(n_1095),
.A2(n_622),
.B1(n_839),
.B2(n_790),
.Y(n_1207)
);

BUFx12f_ASAP7_75t_L g1208 ( 
.A(n_987),
.Y(n_1208)
);

AO31x2_ASAP7_75t_L g1209 ( 
.A1(n_1096),
.A2(n_848),
.A3(n_1099),
.B(n_1121),
.Y(n_1209)
);

INVx3_ASAP7_75t_SL g1210 ( 
.A(n_977),
.Y(n_1210)
);

OAI21xp5_ASAP7_75t_L g1211 ( 
.A1(n_984),
.A2(n_839),
.B(n_622),
.Y(n_1211)
);

BUFx12f_ASAP7_75t_L g1212 ( 
.A(n_987),
.Y(n_1212)
);

INVx3_ASAP7_75t_L g1213 ( 
.A(n_1052),
.Y(n_1213)
);

NOR2x1_ASAP7_75t_R g1214 ( 
.A(n_987),
.B(n_421),
.Y(n_1214)
);

OAI21x1_ASAP7_75t_L g1215 ( 
.A1(n_994),
.A2(n_806),
.B(n_1007),
.Y(n_1215)
);

OAI21x1_ASAP7_75t_L g1216 ( 
.A1(n_994),
.A2(n_806),
.B(n_1007),
.Y(n_1216)
);

CKINVDCx5p33_ASAP7_75t_R g1217 ( 
.A(n_977),
.Y(n_1217)
);

AOI21xp5_ASAP7_75t_L g1218 ( 
.A1(n_1101),
.A2(n_622),
.B(n_1075),
.Y(n_1218)
);

NAND2xp5_ASAP7_75t_L g1219 ( 
.A(n_1051),
.B(n_622),
.Y(n_1219)
);

OA21x2_ASAP7_75t_L g1220 ( 
.A1(n_1075),
.A2(n_1107),
.B(n_1101),
.Y(n_1220)
);

NAND3xp33_ASAP7_75t_SL g1221 ( 
.A(n_984),
.B(n_622),
.C(n_839),
.Y(n_1221)
);

OAI21xp5_ASAP7_75t_L g1222 ( 
.A1(n_984),
.A2(n_839),
.B(n_622),
.Y(n_1222)
);

NAND2xp5_ASAP7_75t_L g1223 ( 
.A(n_1051),
.B(n_622),
.Y(n_1223)
);

OR2x2_ASAP7_75t_L g1224 ( 
.A(n_975),
.B(n_661),
.Y(n_1224)
);

NAND2xp5_ASAP7_75t_L g1225 ( 
.A(n_1051),
.B(n_622),
.Y(n_1225)
);

NAND2xp5_ASAP7_75t_L g1226 ( 
.A(n_1051),
.B(n_622),
.Y(n_1226)
);

NOR2xp33_ASAP7_75t_L g1227 ( 
.A(n_1051),
.B(n_622),
.Y(n_1227)
);

AOI221x1_ASAP7_75t_L g1228 ( 
.A1(n_1042),
.A2(n_839),
.B1(n_622),
.B2(n_1055),
.C(n_1029),
.Y(n_1228)
);

NAND2xp5_ASAP7_75t_L g1229 ( 
.A(n_1051),
.B(n_622),
.Y(n_1229)
);

AO31x2_ASAP7_75t_L g1230 ( 
.A1(n_1096),
.A2(n_848),
.A3(n_1099),
.B(n_1121),
.Y(n_1230)
);

OAI22xp5_ASAP7_75t_L g1231 ( 
.A1(n_1051),
.A2(n_622),
.B1(n_839),
.B2(n_790),
.Y(n_1231)
);

OR2x2_ASAP7_75t_L g1232 ( 
.A(n_975),
.B(n_661),
.Y(n_1232)
);

OAI21x1_ASAP7_75t_L g1233 ( 
.A1(n_994),
.A2(n_806),
.B(n_1007),
.Y(n_1233)
);

INVx1_ASAP7_75t_L g1234 ( 
.A(n_1063),
.Y(n_1234)
);

NAND3xp33_ASAP7_75t_SL g1235 ( 
.A(n_984),
.B(n_622),
.C(n_839),
.Y(n_1235)
);

INVxp67_ASAP7_75t_SL g1236 ( 
.A(n_1021),
.Y(n_1236)
);

OAI21x1_ASAP7_75t_L g1237 ( 
.A1(n_994),
.A2(n_806),
.B(n_1007),
.Y(n_1237)
);

AOI21xp5_ASAP7_75t_L g1238 ( 
.A1(n_1101),
.A2(n_622),
.B(n_1075),
.Y(n_1238)
);

AOI21xp5_ASAP7_75t_L g1239 ( 
.A1(n_1101),
.A2(n_622),
.B(n_1075),
.Y(n_1239)
);

BUFx4f_ASAP7_75t_SL g1240 ( 
.A(n_975),
.Y(n_1240)
);

AOI21xp5_ASAP7_75t_L g1241 ( 
.A1(n_1101),
.A2(n_622),
.B(n_1075),
.Y(n_1241)
);

AOI22xp5_ASAP7_75t_L g1242 ( 
.A1(n_1081),
.A2(n_839),
.B1(n_622),
.B2(n_1010),
.Y(n_1242)
);

OA21x2_ASAP7_75t_L g1243 ( 
.A1(n_1075),
.A2(n_1107),
.B(n_1101),
.Y(n_1243)
);

OAI21xp5_ASAP7_75t_L g1244 ( 
.A1(n_984),
.A2(n_839),
.B(n_622),
.Y(n_1244)
);

INVx1_ASAP7_75t_L g1245 ( 
.A(n_1063),
.Y(n_1245)
);

O2A1O1Ixp33_ASAP7_75t_L g1246 ( 
.A1(n_984),
.A2(n_622),
.B(n_839),
.C(n_736),
.Y(n_1246)
);

O2A1O1Ixp33_ASAP7_75t_SL g1247 ( 
.A1(n_984),
.A2(n_839),
.B(n_622),
.C(n_1062),
.Y(n_1247)
);

AND2x4_ASAP7_75t_L g1248 ( 
.A(n_1067),
.B(n_1009),
.Y(n_1248)
);

INVx1_ASAP7_75t_L g1249 ( 
.A(n_1063),
.Y(n_1249)
);

AOI21xp5_ASAP7_75t_L g1250 ( 
.A1(n_1101),
.A2(n_622),
.B(n_1075),
.Y(n_1250)
);

BUFx10_ASAP7_75t_L g1251 ( 
.A(n_977),
.Y(n_1251)
);

OAI21x1_ASAP7_75t_L g1252 ( 
.A1(n_994),
.A2(n_806),
.B(n_1007),
.Y(n_1252)
);

INVx1_ASAP7_75t_SL g1253 ( 
.A(n_975),
.Y(n_1253)
);

OAI21x1_ASAP7_75t_L g1254 ( 
.A1(n_994),
.A2(n_806),
.B(n_1007),
.Y(n_1254)
);

OAI22xp5_ASAP7_75t_L g1255 ( 
.A1(n_1051),
.A2(n_622),
.B1(n_839),
.B2(n_790),
.Y(n_1255)
);

AO31x2_ASAP7_75t_L g1256 ( 
.A1(n_1096),
.A2(n_848),
.A3(n_1099),
.B(n_1121),
.Y(n_1256)
);

AO32x2_ASAP7_75t_L g1257 ( 
.A1(n_1096),
.A2(n_1041),
.A3(n_1048),
.B1(n_857),
.B2(n_1065),
.Y(n_1257)
);

OAI21xp5_ASAP7_75t_SL g1258 ( 
.A1(n_1038),
.A2(n_839),
.B(n_622),
.Y(n_1258)
);

OAI22x1_ASAP7_75t_L g1259 ( 
.A1(n_1081),
.A2(n_839),
.B1(n_1051),
.B2(n_1016),
.Y(n_1259)
);

AO31x2_ASAP7_75t_L g1260 ( 
.A1(n_1096),
.A2(n_848),
.A3(n_1099),
.B(n_1121),
.Y(n_1260)
);

NOR2xp33_ASAP7_75t_L g1261 ( 
.A(n_1051),
.B(n_622),
.Y(n_1261)
);

OAI21x1_ASAP7_75t_L g1262 ( 
.A1(n_994),
.A2(n_806),
.B(n_1007),
.Y(n_1262)
);

AOI221xp5_ASAP7_75t_SL g1263 ( 
.A1(n_1041),
.A2(n_839),
.B1(n_1026),
.B2(n_1048),
.C(n_1036),
.Y(n_1263)
);

AO31x2_ASAP7_75t_L g1264 ( 
.A1(n_1096),
.A2(n_848),
.A3(n_1099),
.B(n_1121),
.Y(n_1264)
);

INVx2_ASAP7_75t_L g1265 ( 
.A(n_979),
.Y(n_1265)
);

O2A1O1Ixp33_ASAP7_75t_SL g1266 ( 
.A1(n_984),
.A2(n_839),
.B(n_622),
.C(n_1062),
.Y(n_1266)
);

INVx1_ASAP7_75t_L g1267 ( 
.A(n_1063),
.Y(n_1267)
);

A2O1A1Ixp33_ASAP7_75t_L g1268 ( 
.A1(n_984),
.A2(n_839),
.B(n_622),
.C(n_945),
.Y(n_1268)
);

INVxp67_ASAP7_75t_SL g1269 ( 
.A(n_1021),
.Y(n_1269)
);

OAI21x1_ASAP7_75t_L g1270 ( 
.A1(n_994),
.A2(n_806),
.B(n_1007),
.Y(n_1270)
);

INVx2_ASAP7_75t_L g1271 ( 
.A(n_979),
.Y(n_1271)
);

OAI21xp5_ASAP7_75t_L g1272 ( 
.A1(n_984),
.A2(n_839),
.B(n_622),
.Y(n_1272)
);

OAI21x1_ASAP7_75t_L g1273 ( 
.A1(n_994),
.A2(n_806),
.B(n_1007),
.Y(n_1273)
);

A2O1A1Ixp33_ASAP7_75t_L g1274 ( 
.A1(n_984),
.A2(n_839),
.B(n_622),
.C(n_945),
.Y(n_1274)
);

NAND2xp5_ASAP7_75t_L g1275 ( 
.A(n_1051),
.B(n_622),
.Y(n_1275)
);

INVx1_ASAP7_75t_SL g1276 ( 
.A(n_975),
.Y(n_1276)
);

NOR2xp33_ASAP7_75t_SL g1277 ( 
.A(n_1033),
.B(n_839),
.Y(n_1277)
);

OAI21xp33_ASAP7_75t_L g1278 ( 
.A1(n_1010),
.A2(n_839),
.B(n_622),
.Y(n_1278)
);

AOI22xp33_ASAP7_75t_L g1279 ( 
.A1(n_1227),
.A2(n_1261),
.B1(n_1278),
.B2(n_1242),
.Y(n_1279)
);

AOI22xp33_ASAP7_75t_SL g1280 ( 
.A1(n_1277),
.A2(n_1128),
.B1(n_1255),
.B2(n_1231),
.Y(n_1280)
);

AOI22xp33_ASAP7_75t_L g1281 ( 
.A1(n_1278),
.A2(n_1242),
.B1(n_1259),
.B2(n_1277),
.Y(n_1281)
);

AOI22xp33_ASAP7_75t_L g1282 ( 
.A1(n_1174),
.A2(n_1225),
.B1(n_1275),
.B2(n_1223),
.Y(n_1282)
);

CKINVDCx6p67_ASAP7_75t_R g1283 ( 
.A(n_1210),
.Y(n_1283)
);

INVx8_ASAP7_75t_L g1284 ( 
.A(n_1150),
.Y(n_1284)
);

CKINVDCx5p33_ASAP7_75t_R g1285 ( 
.A(n_1217),
.Y(n_1285)
);

AOI22xp33_ASAP7_75t_L g1286 ( 
.A1(n_1174),
.A2(n_1219),
.B1(n_1226),
.B2(n_1229),
.Y(n_1286)
);

CKINVDCx11_ASAP7_75t_R g1287 ( 
.A(n_1203),
.Y(n_1287)
);

CKINVDCx5p33_ASAP7_75t_R g1288 ( 
.A(n_1141),
.Y(n_1288)
);

AOI22xp33_ASAP7_75t_L g1289 ( 
.A1(n_1221),
.A2(n_1235),
.B1(n_1132),
.B2(n_1244),
.Y(n_1289)
);

AOI22xp33_ASAP7_75t_L g1290 ( 
.A1(n_1132),
.A2(n_1272),
.B1(n_1222),
.B2(n_1211),
.Y(n_1290)
);

NAND2xp5_ASAP7_75t_L g1291 ( 
.A(n_1139),
.B(n_1133),
.Y(n_1291)
);

NAND2xp5_ASAP7_75t_L g1292 ( 
.A(n_1138),
.B(n_1258),
.Y(n_1292)
);

AOI22xp33_ASAP7_75t_L g1293 ( 
.A1(n_1211),
.A2(n_1222),
.B1(n_1152),
.B2(n_1143),
.Y(n_1293)
);

INVx8_ASAP7_75t_L g1294 ( 
.A(n_1150),
.Y(n_1294)
);

INVx2_ASAP7_75t_SL g1295 ( 
.A(n_1141),
.Y(n_1295)
);

OAI22xp5_ASAP7_75t_L g1296 ( 
.A1(n_1258),
.A2(n_1268),
.B1(n_1274),
.B2(n_1180),
.Y(n_1296)
);

INVx6_ASAP7_75t_L g1297 ( 
.A(n_1163),
.Y(n_1297)
);

AOI22xp33_ASAP7_75t_L g1298 ( 
.A1(n_1207),
.A2(n_1149),
.B1(n_1155),
.B2(n_1166),
.Y(n_1298)
);

BUFx10_ASAP7_75t_L g1299 ( 
.A(n_1142),
.Y(n_1299)
);

OAI22xp5_ASAP7_75t_L g1300 ( 
.A1(n_1224),
.A2(n_1232),
.B1(n_1157),
.B2(n_1196),
.Y(n_1300)
);

AND2x2_ASAP7_75t_L g1301 ( 
.A(n_1248),
.B(n_1253),
.Y(n_1301)
);

AOI22xp33_ASAP7_75t_SL g1302 ( 
.A1(n_1172),
.A2(n_1171),
.B1(n_1240),
.B2(n_1149),
.Y(n_1302)
);

INVx1_ASAP7_75t_L g1303 ( 
.A(n_1130),
.Y(n_1303)
);

CKINVDCx20_ASAP7_75t_R g1304 ( 
.A(n_1151),
.Y(n_1304)
);

AOI22xp33_ASAP7_75t_L g1305 ( 
.A1(n_1177),
.A2(n_1127),
.B1(n_1154),
.B2(n_1263),
.Y(n_1305)
);

INVx6_ASAP7_75t_L g1306 ( 
.A(n_1163),
.Y(n_1306)
);

INVx1_ASAP7_75t_SL g1307 ( 
.A(n_1253),
.Y(n_1307)
);

BUFx6f_ASAP7_75t_L g1308 ( 
.A(n_1163),
.Y(n_1308)
);

CKINVDCx11_ASAP7_75t_R g1309 ( 
.A(n_1208),
.Y(n_1309)
);

INVx4_ASAP7_75t_L g1310 ( 
.A(n_1199),
.Y(n_1310)
);

AOI22xp33_ASAP7_75t_L g1311 ( 
.A1(n_1263),
.A2(n_1165),
.B1(n_1175),
.B2(n_1190),
.Y(n_1311)
);

INVx8_ASAP7_75t_L g1312 ( 
.A(n_1212),
.Y(n_1312)
);

BUFx6f_ASAP7_75t_L g1313 ( 
.A(n_1248),
.Y(n_1313)
);

INVx6_ASAP7_75t_L g1314 ( 
.A(n_1251),
.Y(n_1314)
);

OAI22xp33_ASAP7_75t_L g1315 ( 
.A1(n_1228),
.A2(n_1236),
.B1(n_1269),
.B2(n_1276),
.Y(n_1315)
);

AOI22xp33_ASAP7_75t_L g1316 ( 
.A1(n_1165),
.A2(n_1245),
.B1(n_1145),
.B2(n_1267),
.Y(n_1316)
);

AOI22xp5_ASAP7_75t_SL g1317 ( 
.A1(n_1159),
.A2(n_1168),
.B1(n_1146),
.B2(n_1276),
.Y(n_1317)
);

BUFx12f_ASAP7_75t_L g1318 ( 
.A(n_1251),
.Y(n_1318)
);

INVx1_ASAP7_75t_L g1319 ( 
.A(n_1234),
.Y(n_1319)
);

INVx1_ASAP7_75t_L g1320 ( 
.A(n_1249),
.Y(n_1320)
);

OAI21xp5_ASAP7_75t_SL g1321 ( 
.A1(n_1246),
.A2(n_1187),
.B(n_1206),
.Y(n_1321)
);

BUFx12f_ASAP7_75t_L g1322 ( 
.A(n_1136),
.Y(n_1322)
);

OAI22xp33_ASAP7_75t_L g1323 ( 
.A1(n_1194),
.A2(n_1188),
.B1(n_1137),
.B2(n_1197),
.Y(n_1323)
);

OAI21xp33_ASAP7_75t_L g1324 ( 
.A1(n_1147),
.A2(n_1241),
.B(n_1239),
.Y(n_1324)
);

NAND2xp5_ASAP7_75t_L g1325 ( 
.A(n_1247),
.B(n_1266),
.Y(n_1325)
);

BUFx6f_ASAP7_75t_L g1326 ( 
.A(n_1185),
.Y(n_1326)
);

BUFx12f_ASAP7_75t_L g1327 ( 
.A(n_1153),
.Y(n_1327)
);

INVx6_ASAP7_75t_L g1328 ( 
.A(n_1185),
.Y(n_1328)
);

AOI22xp33_ASAP7_75t_L g1329 ( 
.A1(n_1218),
.A2(n_1250),
.B1(n_1238),
.B2(n_1182),
.Y(n_1329)
);

AOI22xp33_ASAP7_75t_L g1330 ( 
.A1(n_1161),
.A2(n_1178),
.B1(n_1271),
.B2(n_1265),
.Y(n_1330)
);

AOI22xp5_ASAP7_75t_L g1331 ( 
.A1(n_1202),
.A2(n_1176),
.B1(n_1144),
.B2(n_1161),
.Y(n_1331)
);

CKINVDCx5p33_ASAP7_75t_R g1332 ( 
.A(n_1214),
.Y(n_1332)
);

INVx1_ASAP7_75t_L g1333 ( 
.A(n_1189),
.Y(n_1333)
);

OAI22xp5_ASAP7_75t_L g1334 ( 
.A1(n_1204),
.A2(n_1162),
.B1(n_1198),
.B2(n_1200),
.Y(n_1334)
);

AOI22xp33_ASAP7_75t_L g1335 ( 
.A1(n_1204),
.A2(n_1186),
.B1(n_1243),
.B2(n_1220),
.Y(n_1335)
);

BUFx6f_ASAP7_75t_L g1336 ( 
.A(n_1183),
.Y(n_1336)
);

BUFx12f_ASAP7_75t_SL g1337 ( 
.A(n_1200),
.Y(n_1337)
);

OAI22xp5_ASAP7_75t_L g1338 ( 
.A1(n_1191),
.A2(n_1201),
.B1(n_1213),
.B2(n_1135),
.Y(n_1338)
);

INVx1_ASAP7_75t_L g1339 ( 
.A(n_1193),
.Y(n_1339)
);

AOI22xp33_ASAP7_75t_L g1340 ( 
.A1(n_1220),
.A2(n_1243),
.B1(n_1129),
.B2(n_1148),
.Y(n_1340)
);

OAI22xp33_ASAP7_75t_L g1341 ( 
.A1(n_1257),
.A2(n_1169),
.B1(n_1170),
.B2(n_1156),
.Y(n_1341)
);

INVx1_ASAP7_75t_L g1342 ( 
.A(n_1131),
.Y(n_1342)
);

AOI22xp33_ASAP7_75t_L g1343 ( 
.A1(n_1158),
.A2(n_1156),
.B1(n_1195),
.B2(n_1184),
.Y(n_1343)
);

INVx1_ASAP7_75t_L g1344 ( 
.A(n_1131),
.Y(n_1344)
);

BUFx12f_ASAP7_75t_L g1345 ( 
.A(n_1205),
.Y(n_1345)
);

AOI22xp33_ASAP7_75t_L g1346 ( 
.A1(n_1181),
.A2(n_1257),
.B1(n_1134),
.B2(n_1262),
.Y(n_1346)
);

AOI22xp33_ASAP7_75t_L g1347 ( 
.A1(n_1257),
.A2(n_1273),
.B1(n_1233),
.B2(n_1237),
.Y(n_1347)
);

INVx1_ASAP7_75t_L g1348 ( 
.A(n_1131),
.Y(n_1348)
);

AOI22xp33_ASAP7_75t_L g1349 ( 
.A1(n_1215),
.A2(n_1216),
.B1(n_1254),
.B2(n_1252),
.Y(n_1349)
);

AOI22xp5_ASAP7_75t_L g1350 ( 
.A1(n_1270),
.A2(n_1164),
.B1(n_1179),
.B2(n_1260),
.Y(n_1350)
);

AOI22xp33_ASAP7_75t_L g1351 ( 
.A1(n_1179),
.A2(n_1173),
.B1(n_1264),
.B2(n_1209),
.Y(n_1351)
);

AOI22xp33_ASAP7_75t_L g1352 ( 
.A1(n_1179),
.A2(n_1173),
.B1(n_1264),
.B2(n_1209),
.Y(n_1352)
);

AOI22xp33_ASAP7_75t_L g1353 ( 
.A1(n_1173),
.A2(n_1230),
.B1(n_1260),
.B2(n_1256),
.Y(n_1353)
);

AOI22xp33_ASAP7_75t_L g1354 ( 
.A1(n_1209),
.A2(n_1230),
.B1(n_1256),
.B2(n_1260),
.Y(n_1354)
);

AOI22xp33_ASAP7_75t_SL g1355 ( 
.A1(n_1167),
.A2(n_1230),
.B1(n_1256),
.B2(n_1264),
.Y(n_1355)
);

AOI22xp33_ASAP7_75t_L g1356 ( 
.A1(n_1167),
.A2(n_839),
.B1(n_1261),
.B2(n_1227),
.Y(n_1356)
);

OAI22xp33_ASAP7_75t_L g1357 ( 
.A1(n_1167),
.A2(n_1242),
.B1(n_1128),
.B2(n_1277),
.Y(n_1357)
);

INVxp67_ASAP7_75t_L g1358 ( 
.A(n_1192),
.Y(n_1358)
);

AOI22xp33_ASAP7_75t_SL g1359 ( 
.A1(n_1277),
.A2(n_839),
.B1(n_622),
.B2(n_1128),
.Y(n_1359)
);

OAI21xp33_ASAP7_75t_L g1360 ( 
.A1(n_1242),
.A2(n_839),
.B(n_622),
.Y(n_1360)
);

AOI22xp33_ASAP7_75t_L g1361 ( 
.A1(n_1227),
.A2(n_839),
.B1(n_1261),
.B2(n_1278),
.Y(n_1361)
);

INVx1_ASAP7_75t_SL g1362 ( 
.A(n_1240),
.Y(n_1362)
);

INVx8_ASAP7_75t_L g1363 ( 
.A(n_1150),
.Y(n_1363)
);

OAI22xp5_ASAP7_75t_L g1364 ( 
.A1(n_1242),
.A2(n_622),
.B1(n_1261),
.B2(n_1227),
.Y(n_1364)
);

INVx6_ASAP7_75t_L g1365 ( 
.A(n_1150),
.Y(n_1365)
);

AOI22xp33_ASAP7_75t_L g1366 ( 
.A1(n_1227),
.A2(n_839),
.B1(n_1261),
.B2(n_1278),
.Y(n_1366)
);

BUFx4f_ASAP7_75t_SL g1367 ( 
.A(n_1208),
.Y(n_1367)
);

BUFx10_ASAP7_75t_L g1368 ( 
.A(n_1217),
.Y(n_1368)
);

OAI22xp5_ASAP7_75t_L g1369 ( 
.A1(n_1242),
.A2(n_622),
.B1(n_1261),
.B2(n_1227),
.Y(n_1369)
);

AOI22xp33_ASAP7_75t_SL g1370 ( 
.A1(n_1277),
.A2(n_839),
.B1(n_622),
.B2(n_1128),
.Y(n_1370)
);

INVx1_ASAP7_75t_SL g1371 ( 
.A(n_1240),
.Y(n_1371)
);

AOI22xp33_ASAP7_75t_L g1372 ( 
.A1(n_1227),
.A2(n_839),
.B1(n_1261),
.B2(n_1278),
.Y(n_1372)
);

BUFx10_ASAP7_75t_L g1373 ( 
.A(n_1217),
.Y(n_1373)
);

OAI22xp5_ASAP7_75t_L g1374 ( 
.A1(n_1242),
.A2(n_622),
.B1(n_1261),
.B2(n_1227),
.Y(n_1374)
);

INVx1_ASAP7_75t_L g1375 ( 
.A(n_1160),
.Y(n_1375)
);

INVx2_ASAP7_75t_L g1376 ( 
.A(n_1140),
.Y(n_1376)
);

BUFx12f_ASAP7_75t_L g1377 ( 
.A(n_1203),
.Y(n_1377)
);

INVx1_ASAP7_75t_L g1378 ( 
.A(n_1160),
.Y(n_1378)
);

CKINVDCx5p33_ASAP7_75t_R g1379 ( 
.A(n_1217),
.Y(n_1379)
);

INVx3_ASAP7_75t_L g1380 ( 
.A(n_1135),
.Y(n_1380)
);

CKINVDCx20_ASAP7_75t_R g1381 ( 
.A(n_1240),
.Y(n_1381)
);

INVx1_ASAP7_75t_L g1382 ( 
.A(n_1160),
.Y(n_1382)
);

CKINVDCx6p67_ASAP7_75t_R g1383 ( 
.A(n_1210),
.Y(n_1383)
);

OAI22xp5_ASAP7_75t_SL g1384 ( 
.A1(n_1128),
.A2(n_954),
.B1(n_1242),
.B2(n_1227),
.Y(n_1384)
);

AOI22xp33_ASAP7_75t_L g1385 ( 
.A1(n_1227),
.A2(n_839),
.B1(n_1261),
.B2(n_1278),
.Y(n_1385)
);

BUFx3_ASAP7_75t_L g1386 ( 
.A(n_1150),
.Y(n_1386)
);

BUFx4_ASAP7_75t_SL g1387 ( 
.A(n_1217),
.Y(n_1387)
);

NAND2xp5_ASAP7_75t_L g1388 ( 
.A(n_1227),
.B(n_1261),
.Y(n_1388)
);

BUFx12f_ASAP7_75t_L g1389 ( 
.A(n_1203),
.Y(n_1389)
);

AOI22xp33_ASAP7_75t_L g1390 ( 
.A1(n_1227),
.A2(n_839),
.B1(n_1261),
.B2(n_1278),
.Y(n_1390)
);

BUFx3_ASAP7_75t_L g1391 ( 
.A(n_1150),
.Y(n_1391)
);

AOI22xp5_ASAP7_75t_L g1392 ( 
.A1(n_1277),
.A2(n_839),
.B1(n_1242),
.B2(n_622),
.Y(n_1392)
);

OR2x2_ASAP7_75t_L g1393 ( 
.A(n_1139),
.B(n_1128),
.Y(n_1393)
);

CKINVDCx6p67_ASAP7_75t_R g1394 ( 
.A(n_1210),
.Y(n_1394)
);

BUFx3_ASAP7_75t_L g1395 ( 
.A(n_1150),
.Y(n_1395)
);

INVx1_ASAP7_75t_SL g1396 ( 
.A(n_1240),
.Y(n_1396)
);

INVxp67_ASAP7_75t_L g1397 ( 
.A(n_1147),
.Y(n_1397)
);

NAND2xp5_ASAP7_75t_L g1398 ( 
.A(n_1227),
.B(n_1261),
.Y(n_1398)
);

AOI22xp33_ASAP7_75t_L g1399 ( 
.A1(n_1227),
.A2(n_839),
.B1(n_1261),
.B2(n_1278),
.Y(n_1399)
);

CKINVDCx11_ASAP7_75t_R g1400 ( 
.A(n_1203),
.Y(n_1400)
);

AOI22xp33_ASAP7_75t_L g1401 ( 
.A1(n_1227),
.A2(n_839),
.B1(n_1261),
.B2(n_1278),
.Y(n_1401)
);

BUFx10_ASAP7_75t_L g1402 ( 
.A(n_1217),
.Y(n_1402)
);

INVx1_ASAP7_75t_L g1403 ( 
.A(n_1160),
.Y(n_1403)
);

INVx4_ASAP7_75t_L g1404 ( 
.A(n_1345),
.Y(n_1404)
);

INVx1_ASAP7_75t_L g1405 ( 
.A(n_1339),
.Y(n_1405)
);

OR2x6_ASAP7_75t_L g1406 ( 
.A(n_1321),
.B(n_1334),
.Y(n_1406)
);

INVx1_ASAP7_75t_L g1407 ( 
.A(n_1342),
.Y(n_1407)
);

INVx1_ASAP7_75t_L g1408 ( 
.A(n_1344),
.Y(n_1408)
);

HB1xp67_ASAP7_75t_SL g1409 ( 
.A(n_1386),
.Y(n_1409)
);

INVx2_ASAP7_75t_L g1410 ( 
.A(n_1348),
.Y(n_1410)
);

INVx1_ASAP7_75t_L g1411 ( 
.A(n_1358),
.Y(n_1411)
);

AO21x2_ASAP7_75t_L g1412 ( 
.A1(n_1341),
.A2(n_1350),
.B(n_1357),
.Y(n_1412)
);

NAND2xp5_ASAP7_75t_L g1413 ( 
.A(n_1282),
.B(n_1286),
.Y(n_1413)
);

INVx2_ASAP7_75t_L g1414 ( 
.A(n_1303),
.Y(n_1414)
);

INVx1_ASAP7_75t_L g1415 ( 
.A(n_1355),
.Y(n_1415)
);

BUFx3_ASAP7_75t_L g1416 ( 
.A(n_1314),
.Y(n_1416)
);

INVx1_ASAP7_75t_L g1417 ( 
.A(n_1354),
.Y(n_1417)
);

OA21x2_ASAP7_75t_L g1418 ( 
.A1(n_1343),
.A2(n_1329),
.B(n_1340),
.Y(n_1418)
);

AND2x2_ASAP7_75t_L g1419 ( 
.A(n_1356),
.B(n_1298),
.Y(n_1419)
);

AND2x2_ASAP7_75t_L g1420 ( 
.A(n_1353),
.B(n_1351),
.Y(n_1420)
);

INVx2_ASAP7_75t_L g1421 ( 
.A(n_1319),
.Y(n_1421)
);

INVx2_ASAP7_75t_L g1422 ( 
.A(n_1320),
.Y(n_1422)
);

AOI22xp33_ASAP7_75t_L g1423 ( 
.A1(n_1384),
.A2(n_1360),
.B1(n_1364),
.B2(n_1369),
.Y(n_1423)
);

INVx1_ASAP7_75t_L g1424 ( 
.A(n_1354),
.Y(n_1424)
);

INVx1_ASAP7_75t_L g1425 ( 
.A(n_1353),
.Y(n_1425)
);

INVx2_ASAP7_75t_L g1426 ( 
.A(n_1375),
.Y(n_1426)
);

INVx2_ASAP7_75t_L g1427 ( 
.A(n_1378),
.Y(n_1427)
);

BUFx12f_ASAP7_75t_L g1428 ( 
.A(n_1287),
.Y(n_1428)
);

INVx2_ASAP7_75t_L g1429 ( 
.A(n_1382),
.Y(n_1429)
);

AND2x2_ASAP7_75t_L g1430 ( 
.A(n_1356),
.B(n_1298),
.Y(n_1430)
);

HB1xp67_ASAP7_75t_L g1431 ( 
.A(n_1325),
.Y(n_1431)
);

BUFx3_ASAP7_75t_L g1432 ( 
.A(n_1314),
.Y(n_1432)
);

INVx2_ASAP7_75t_L g1433 ( 
.A(n_1403),
.Y(n_1433)
);

BUFx2_ASAP7_75t_L g1434 ( 
.A(n_1315),
.Y(n_1434)
);

INVx1_ASAP7_75t_L g1435 ( 
.A(n_1351),
.Y(n_1435)
);

INVx1_ASAP7_75t_L g1436 ( 
.A(n_1352),
.Y(n_1436)
);

OA21x2_ASAP7_75t_L g1437 ( 
.A1(n_1343),
.A2(n_1329),
.B(n_1340),
.Y(n_1437)
);

AOI22xp33_ASAP7_75t_SL g1438 ( 
.A1(n_1374),
.A2(n_1296),
.B1(n_1388),
.B2(n_1398),
.Y(n_1438)
);

INVx1_ASAP7_75t_L g1439 ( 
.A(n_1352),
.Y(n_1439)
);

INVx1_ASAP7_75t_L g1440 ( 
.A(n_1324),
.Y(n_1440)
);

AOI21xp5_ASAP7_75t_L g1441 ( 
.A1(n_1341),
.A2(n_1311),
.B(n_1335),
.Y(n_1441)
);

AND2x2_ASAP7_75t_L g1442 ( 
.A(n_1290),
.B(n_1293),
.Y(n_1442)
);

OAI21x1_ASAP7_75t_L g1443 ( 
.A1(n_1335),
.A2(n_1349),
.B(n_1347),
.Y(n_1443)
);

HB1xp67_ASAP7_75t_L g1444 ( 
.A(n_1315),
.Y(n_1444)
);

INVx1_ASAP7_75t_L g1445 ( 
.A(n_1316),
.Y(n_1445)
);

OAI21x1_ASAP7_75t_L g1446 ( 
.A1(n_1349),
.A2(n_1347),
.B(n_1346),
.Y(n_1446)
);

AND2x2_ASAP7_75t_L g1447 ( 
.A(n_1290),
.B(n_1293),
.Y(n_1447)
);

AND2x2_ASAP7_75t_L g1448 ( 
.A(n_1305),
.B(n_1289),
.Y(n_1448)
);

AND2x4_ASAP7_75t_L g1449 ( 
.A(n_1326),
.B(n_1376),
.Y(n_1449)
);

INVx1_ASAP7_75t_L g1450 ( 
.A(n_1316),
.Y(n_1450)
);

INVx1_ASAP7_75t_L g1451 ( 
.A(n_1311),
.Y(n_1451)
);

AOI21x1_ASAP7_75t_L g1452 ( 
.A1(n_1338),
.A2(n_1292),
.B(n_1300),
.Y(n_1452)
);

INVx1_ASAP7_75t_L g1453 ( 
.A(n_1333),
.Y(n_1453)
);

OA21x2_ASAP7_75t_L g1454 ( 
.A1(n_1346),
.A2(n_1305),
.B(n_1289),
.Y(n_1454)
);

HB1xp67_ASAP7_75t_L g1455 ( 
.A(n_1357),
.Y(n_1455)
);

OR2x2_ASAP7_75t_L g1456 ( 
.A(n_1281),
.B(n_1393),
.Y(n_1456)
);

OAI21x1_ASAP7_75t_L g1457 ( 
.A1(n_1330),
.A2(n_1331),
.B(n_1380),
.Y(n_1457)
);

NOR2x1_ASAP7_75t_R g1458 ( 
.A(n_1400),
.B(n_1377),
.Y(n_1458)
);

INVx2_ASAP7_75t_SL g1459 ( 
.A(n_1328),
.Y(n_1459)
);

OR2x2_ASAP7_75t_L g1460 ( 
.A(n_1279),
.B(n_1323),
.Y(n_1460)
);

AND2x2_ASAP7_75t_L g1461 ( 
.A(n_1280),
.B(n_1279),
.Y(n_1461)
);

INVx1_ASAP7_75t_L g1462 ( 
.A(n_1323),
.Y(n_1462)
);

NOR2xp33_ASAP7_75t_L g1463 ( 
.A(n_1397),
.B(n_1301),
.Y(n_1463)
);

AOI22xp33_ASAP7_75t_L g1464 ( 
.A1(n_1359),
.A2(n_1370),
.B1(n_1392),
.B2(n_1399),
.Y(n_1464)
);

INVx1_ASAP7_75t_SL g1465 ( 
.A(n_1307),
.Y(n_1465)
);

INVx1_ASAP7_75t_L g1466 ( 
.A(n_1291),
.Y(n_1466)
);

INVx2_ASAP7_75t_L g1467 ( 
.A(n_1328),
.Y(n_1467)
);

AND2x2_ASAP7_75t_L g1468 ( 
.A(n_1282),
.B(n_1286),
.Y(n_1468)
);

BUFx12f_ASAP7_75t_L g1469 ( 
.A(n_1309),
.Y(n_1469)
);

AND2x2_ASAP7_75t_L g1470 ( 
.A(n_1361),
.B(n_1385),
.Y(n_1470)
);

INVx1_ASAP7_75t_L g1471 ( 
.A(n_1336),
.Y(n_1471)
);

HB1xp67_ASAP7_75t_L g1472 ( 
.A(n_1313),
.Y(n_1472)
);

INVx2_ASAP7_75t_L g1473 ( 
.A(n_1308),
.Y(n_1473)
);

NAND2xp5_ASAP7_75t_L g1474 ( 
.A(n_1366),
.B(n_1372),
.Y(n_1474)
);

BUFx12f_ASAP7_75t_L g1475 ( 
.A(n_1285),
.Y(n_1475)
);

INVx1_ASAP7_75t_L g1476 ( 
.A(n_1372),
.Y(n_1476)
);

OA21x2_ASAP7_75t_L g1477 ( 
.A1(n_1385),
.A2(n_1390),
.B(n_1401),
.Y(n_1477)
);

BUFx3_ASAP7_75t_L g1478 ( 
.A(n_1299),
.Y(n_1478)
);

AO21x1_ASAP7_75t_SL g1479 ( 
.A1(n_1390),
.A2(n_1302),
.B(n_1337),
.Y(n_1479)
);

AO21x2_ASAP7_75t_L g1480 ( 
.A1(n_1317),
.A2(n_1297),
.B(n_1306),
.Y(n_1480)
);

NOR2x1_ASAP7_75t_R g1481 ( 
.A(n_1389),
.B(n_1318),
.Y(n_1481)
);

NAND2xp5_ASAP7_75t_L g1482 ( 
.A(n_1391),
.B(n_1395),
.Y(n_1482)
);

BUFx3_ASAP7_75t_L g1483 ( 
.A(n_1299),
.Y(n_1483)
);

INVx1_ASAP7_75t_L g1484 ( 
.A(n_1391),
.Y(n_1484)
);

AND2x4_ASAP7_75t_L g1485 ( 
.A(n_1295),
.B(n_1395),
.Y(n_1485)
);

CKINVDCx20_ASAP7_75t_R g1486 ( 
.A(n_1469),
.Y(n_1486)
);

INVx4_ASAP7_75t_L g1487 ( 
.A(n_1404),
.Y(n_1487)
);

OAI21xp5_ASAP7_75t_L g1488 ( 
.A1(n_1423),
.A2(n_1288),
.B(n_1304),
.Y(n_1488)
);

OAI221xp5_ASAP7_75t_L g1489 ( 
.A1(n_1438),
.A2(n_1396),
.B1(n_1362),
.B2(n_1371),
.C(n_1332),
.Y(n_1489)
);

AND2x4_ASAP7_75t_L g1490 ( 
.A(n_1416),
.B(n_1310),
.Y(n_1490)
);

AOI22xp5_ASAP7_75t_L g1491 ( 
.A1(n_1438),
.A2(n_1322),
.B1(n_1394),
.B2(n_1383),
.Y(n_1491)
);

AND2x4_ASAP7_75t_L g1492 ( 
.A(n_1414),
.B(n_1379),
.Y(n_1492)
);

AND2x2_ASAP7_75t_L g1493 ( 
.A(n_1463),
.B(n_1297),
.Y(n_1493)
);

OR2x2_ASAP7_75t_L g1494 ( 
.A(n_1456),
.B(n_1283),
.Y(n_1494)
);

O2A1O1Ixp33_ASAP7_75t_L g1495 ( 
.A1(n_1413),
.A2(n_1381),
.B(n_1294),
.C(n_1284),
.Y(n_1495)
);

O2A1O1Ixp33_ASAP7_75t_SL g1496 ( 
.A1(n_1413),
.A2(n_1312),
.B(n_1367),
.C(n_1363),
.Y(n_1496)
);

AOI221xp5_ASAP7_75t_L g1497 ( 
.A1(n_1461),
.A2(n_1464),
.B1(n_1468),
.B2(n_1448),
.C(n_1434),
.Y(n_1497)
);

OR2x6_ASAP7_75t_L g1498 ( 
.A(n_1406),
.B(n_1312),
.Y(n_1498)
);

OR2x2_ASAP7_75t_L g1499 ( 
.A(n_1456),
.B(n_1414),
.Y(n_1499)
);

OAI21xp5_ASAP7_75t_L g1500 ( 
.A1(n_1461),
.A2(n_1402),
.B(n_1373),
.Y(n_1500)
);

A2O1A1Ixp33_ASAP7_75t_L g1501 ( 
.A1(n_1441),
.A2(n_1284),
.B(n_1294),
.C(n_1363),
.Y(n_1501)
);

A2O1A1Ixp33_ASAP7_75t_L g1502 ( 
.A1(n_1441),
.A2(n_1294),
.B(n_1363),
.C(n_1312),
.Y(n_1502)
);

INVx1_ASAP7_75t_SL g1503 ( 
.A(n_1465),
.Y(n_1503)
);

NAND3xp33_ASAP7_75t_L g1504 ( 
.A(n_1460),
.B(n_1468),
.C(n_1440),
.Y(n_1504)
);

OR2x2_ASAP7_75t_SL g1505 ( 
.A(n_1460),
.B(n_1477),
.Y(n_1505)
);

NOR2xp33_ASAP7_75t_SL g1506 ( 
.A(n_1458),
.B(n_1367),
.Y(n_1506)
);

NAND2xp5_ASAP7_75t_L g1507 ( 
.A(n_1466),
.B(n_1365),
.Y(n_1507)
);

NAND2xp5_ASAP7_75t_L g1508 ( 
.A(n_1453),
.B(n_1440),
.Y(n_1508)
);

OA21x2_ASAP7_75t_L g1509 ( 
.A1(n_1446),
.A2(n_1365),
.B(n_1327),
.Y(n_1509)
);

NAND2x1_ASAP7_75t_L g1510 ( 
.A(n_1404),
.B(n_1387),
.Y(n_1510)
);

AND2x4_ASAP7_75t_L g1511 ( 
.A(n_1432),
.B(n_1368),
.Y(n_1511)
);

OAI22xp5_ASAP7_75t_L g1512 ( 
.A1(n_1406),
.A2(n_1368),
.B1(n_1373),
.B2(n_1402),
.Y(n_1512)
);

NOR2x1_ASAP7_75t_SL g1513 ( 
.A(n_1406),
.B(n_1480),
.Y(n_1513)
);

NOR2x1_ASAP7_75t_SL g1514 ( 
.A(n_1406),
.B(n_1480),
.Y(n_1514)
);

AND2x2_ASAP7_75t_L g1515 ( 
.A(n_1467),
.B(n_1449),
.Y(n_1515)
);

INVxp67_ASAP7_75t_L g1516 ( 
.A(n_1431),
.Y(n_1516)
);

AOI21xp5_ASAP7_75t_L g1517 ( 
.A1(n_1418),
.A2(n_1437),
.B(n_1406),
.Y(n_1517)
);

AOI221xp5_ASAP7_75t_L g1518 ( 
.A1(n_1448),
.A2(n_1434),
.B1(n_1455),
.B2(n_1442),
.C(n_1447),
.Y(n_1518)
);

AO21x2_ASAP7_75t_L g1519 ( 
.A1(n_1443),
.A2(n_1446),
.B(n_1412),
.Y(n_1519)
);

A2O1A1Ixp33_ASAP7_75t_L g1520 ( 
.A1(n_1419),
.A2(n_1430),
.B(n_1447),
.C(n_1442),
.Y(n_1520)
);

INVx2_ASAP7_75t_L g1521 ( 
.A(n_1421),
.Y(n_1521)
);

AO21x2_ASAP7_75t_L g1522 ( 
.A1(n_1443),
.A2(n_1446),
.B(n_1412),
.Y(n_1522)
);

OAI22xp5_ASAP7_75t_L g1523 ( 
.A1(n_1406),
.A2(n_1409),
.B1(n_1474),
.B2(n_1478),
.Y(n_1523)
);

AND2x2_ASAP7_75t_L g1524 ( 
.A(n_1449),
.B(n_1473),
.Y(n_1524)
);

AND2x2_ASAP7_75t_L g1525 ( 
.A(n_1449),
.B(n_1473),
.Y(n_1525)
);

AND2x4_ASAP7_75t_L g1526 ( 
.A(n_1421),
.B(n_1422),
.Y(n_1526)
);

NOR2xp33_ASAP7_75t_L g1527 ( 
.A(n_1452),
.B(n_1462),
.Y(n_1527)
);

HB1xp67_ASAP7_75t_L g1528 ( 
.A(n_1411),
.Y(n_1528)
);

A2O1A1Ixp33_ASAP7_75t_L g1529 ( 
.A1(n_1419),
.A2(n_1430),
.B(n_1444),
.C(n_1455),
.Y(n_1529)
);

OA21x2_ASAP7_75t_L g1530 ( 
.A1(n_1443),
.A2(n_1457),
.B(n_1407),
.Y(n_1530)
);

O2A1O1Ixp33_ASAP7_75t_L g1531 ( 
.A1(n_1474),
.A2(n_1444),
.B(n_1462),
.C(n_1476),
.Y(n_1531)
);

OAI21xp33_ASAP7_75t_L g1532 ( 
.A1(n_1452),
.A2(n_1470),
.B(n_1476),
.Y(n_1532)
);

AO22x2_ASAP7_75t_L g1533 ( 
.A1(n_1415),
.A2(n_1425),
.B1(n_1424),
.B2(n_1417),
.Y(n_1533)
);

AOI221xp5_ASAP7_75t_L g1534 ( 
.A1(n_1445),
.A2(n_1450),
.B1(n_1451),
.B2(n_1415),
.C(n_1424),
.Y(n_1534)
);

AND2x4_ASAP7_75t_L g1535 ( 
.A(n_1422),
.B(n_1426),
.Y(n_1535)
);

OA21x2_ASAP7_75t_L g1536 ( 
.A1(n_1457),
.A2(n_1408),
.B(n_1407),
.Y(n_1536)
);

AND2x2_ASAP7_75t_L g1537 ( 
.A(n_1472),
.B(n_1480),
.Y(n_1537)
);

OAI21xp5_ASAP7_75t_L g1538 ( 
.A1(n_1404),
.A2(n_1457),
.B(n_1477),
.Y(n_1538)
);

INVx2_ASAP7_75t_SL g1539 ( 
.A(n_1478),
.Y(n_1539)
);

INVx2_ASAP7_75t_L g1540 ( 
.A(n_1521),
.Y(n_1540)
);

HB1xp67_ASAP7_75t_L g1541 ( 
.A(n_1516),
.Y(n_1541)
);

INVx1_ASAP7_75t_SL g1542 ( 
.A(n_1503),
.Y(n_1542)
);

INVx2_ASAP7_75t_L g1543 ( 
.A(n_1536),
.Y(n_1543)
);

AND2x4_ASAP7_75t_L g1544 ( 
.A(n_1526),
.B(n_1410),
.Y(n_1544)
);

AND2x2_ASAP7_75t_L g1545 ( 
.A(n_1537),
.B(n_1420),
.Y(n_1545)
);

INVx1_ASAP7_75t_L g1546 ( 
.A(n_1535),
.Y(n_1546)
);

AND2x4_ASAP7_75t_L g1547 ( 
.A(n_1513),
.B(n_1410),
.Y(n_1547)
);

HB1xp67_ASAP7_75t_L g1548 ( 
.A(n_1516),
.Y(n_1548)
);

NOR2xp33_ASAP7_75t_L g1549 ( 
.A(n_1494),
.B(n_1404),
.Y(n_1549)
);

AOI22xp33_ASAP7_75t_L g1550 ( 
.A1(n_1497),
.A2(n_1479),
.B1(n_1518),
.B2(n_1504),
.Y(n_1550)
);

INVx2_ASAP7_75t_L g1551 ( 
.A(n_1536),
.Y(n_1551)
);

OR2x2_ASAP7_75t_L g1552 ( 
.A(n_1499),
.B(n_1412),
.Y(n_1552)
);

NAND2xp5_ASAP7_75t_L g1553 ( 
.A(n_1532),
.B(n_1427),
.Y(n_1553)
);

AOI22xp33_ASAP7_75t_L g1554 ( 
.A1(n_1491),
.A2(n_1479),
.B1(n_1477),
.B2(n_1451),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_1528),
.Y(n_1555)
);

AND2x4_ASAP7_75t_L g1556 ( 
.A(n_1514),
.B(n_1410),
.Y(n_1556)
);

AND2x2_ASAP7_75t_L g1557 ( 
.A(n_1524),
.B(n_1420),
.Y(n_1557)
);

AOI22xp33_ASAP7_75t_L g1558 ( 
.A1(n_1498),
.A2(n_1477),
.B1(n_1454),
.B2(n_1450),
.Y(n_1558)
);

NAND2xp5_ASAP7_75t_L g1559 ( 
.A(n_1527),
.B(n_1427),
.Y(n_1559)
);

OAI221xp5_ASAP7_75t_L g1560 ( 
.A1(n_1500),
.A2(n_1478),
.B1(n_1483),
.B2(n_1459),
.C(n_1445),
.Y(n_1560)
);

OR2x2_ASAP7_75t_L g1561 ( 
.A(n_1505),
.B(n_1412),
.Y(n_1561)
);

AND2x2_ASAP7_75t_L g1562 ( 
.A(n_1525),
.B(n_1420),
.Y(n_1562)
);

INVx2_ASAP7_75t_L g1563 ( 
.A(n_1530),
.Y(n_1563)
);

INVx1_ASAP7_75t_L g1564 ( 
.A(n_1508),
.Y(n_1564)
);

OR2x2_ASAP7_75t_L g1565 ( 
.A(n_1519),
.B(n_1435),
.Y(n_1565)
);

NAND2xp5_ASAP7_75t_L g1566 ( 
.A(n_1527),
.B(n_1429),
.Y(n_1566)
);

OR2x2_ASAP7_75t_L g1567 ( 
.A(n_1519),
.B(n_1436),
.Y(n_1567)
);

NOR2xp33_ASAP7_75t_L g1568 ( 
.A(n_1492),
.B(n_1483),
.Y(n_1568)
);

AND2x4_ASAP7_75t_L g1569 ( 
.A(n_1538),
.B(n_1433),
.Y(n_1569)
);

AOI22xp33_ASAP7_75t_L g1570 ( 
.A1(n_1550),
.A2(n_1477),
.B1(n_1454),
.B2(n_1498),
.Y(n_1570)
);

BUFx2_ASAP7_75t_L g1571 ( 
.A(n_1547),
.Y(n_1571)
);

NOR2xp67_ASAP7_75t_L g1572 ( 
.A(n_1561),
.B(n_1517),
.Y(n_1572)
);

AND2x2_ASAP7_75t_L g1573 ( 
.A(n_1545),
.B(n_1522),
.Y(n_1573)
);

OAI31xp33_ASAP7_75t_L g1574 ( 
.A1(n_1560),
.A2(n_1529),
.A3(n_1520),
.B(n_1523),
.Y(n_1574)
);

OAI221xp5_ASAP7_75t_L g1575 ( 
.A1(n_1554),
.A2(n_1520),
.B1(n_1529),
.B2(n_1488),
.C(n_1506),
.Y(n_1575)
);

OR2x2_ASAP7_75t_L g1576 ( 
.A(n_1565),
.B(n_1522),
.Y(n_1576)
);

OR2x2_ASAP7_75t_L g1577 ( 
.A(n_1565),
.B(n_1530),
.Y(n_1577)
);

NAND2xp5_ASAP7_75t_L g1578 ( 
.A(n_1564),
.B(n_1533),
.Y(n_1578)
);

AND2x2_ASAP7_75t_L g1579 ( 
.A(n_1545),
.B(n_1509),
.Y(n_1579)
);

INVx1_ASAP7_75t_L g1580 ( 
.A(n_1540),
.Y(n_1580)
);

INVx1_ASAP7_75t_L g1581 ( 
.A(n_1540),
.Y(n_1581)
);

AND2x2_ASAP7_75t_L g1582 ( 
.A(n_1546),
.B(n_1533),
.Y(n_1582)
);

NAND2xp5_ASAP7_75t_L g1583 ( 
.A(n_1564),
.B(n_1533),
.Y(n_1583)
);

OR2x2_ASAP7_75t_L g1584 ( 
.A(n_1567),
.B(n_1417),
.Y(n_1584)
);

NAND4xp25_ASAP7_75t_L g1585 ( 
.A(n_1558),
.B(n_1531),
.C(n_1534),
.D(n_1489),
.Y(n_1585)
);

AND2x4_ASAP7_75t_L g1586 ( 
.A(n_1547),
.B(n_1515),
.Y(n_1586)
);

AO21x2_ASAP7_75t_L g1587 ( 
.A1(n_1563),
.A2(n_1408),
.B(n_1405),
.Y(n_1587)
);

NAND2x1_ASAP7_75t_L g1588 ( 
.A(n_1556),
.B(n_1498),
.Y(n_1588)
);

OAI22xp5_ASAP7_75t_L g1589 ( 
.A1(n_1561),
.A2(n_1409),
.B1(n_1531),
.B2(n_1486),
.Y(n_1589)
);

BUFx3_ASAP7_75t_L g1590 ( 
.A(n_1556),
.Y(n_1590)
);

BUFx2_ASAP7_75t_L g1591 ( 
.A(n_1556),
.Y(n_1591)
);

INVx3_ASAP7_75t_L g1592 ( 
.A(n_1556),
.Y(n_1592)
);

OAI21xp33_ASAP7_75t_L g1593 ( 
.A1(n_1567),
.A2(n_1553),
.B(n_1559),
.Y(n_1593)
);

AND2x2_ASAP7_75t_L g1594 ( 
.A(n_1557),
.B(n_1562),
.Y(n_1594)
);

OAI321xp33_ASAP7_75t_L g1595 ( 
.A1(n_1566),
.A2(n_1512),
.A3(n_1502),
.B1(n_1495),
.B2(n_1501),
.C(n_1507),
.Y(n_1595)
);

AOI221xp5_ASAP7_75t_L g1596 ( 
.A1(n_1569),
.A2(n_1495),
.B1(n_1439),
.B2(n_1436),
.C(n_1502),
.Y(n_1596)
);

INVx3_ASAP7_75t_L g1597 ( 
.A(n_1590),
.Y(n_1597)
);

AND2x2_ASAP7_75t_L g1598 ( 
.A(n_1571),
.B(n_1569),
.Y(n_1598)
);

AND2x2_ASAP7_75t_L g1599 ( 
.A(n_1571),
.B(n_1569),
.Y(n_1599)
);

NAND2xp5_ASAP7_75t_L g1600 ( 
.A(n_1593),
.B(n_1541),
.Y(n_1600)
);

AND2x2_ASAP7_75t_L g1601 ( 
.A(n_1571),
.B(n_1569),
.Y(n_1601)
);

INVx1_ASAP7_75t_L g1602 ( 
.A(n_1580),
.Y(n_1602)
);

INVx1_ASAP7_75t_L g1603 ( 
.A(n_1580),
.Y(n_1603)
);

AND2x2_ASAP7_75t_L g1604 ( 
.A(n_1591),
.B(n_1563),
.Y(n_1604)
);

NAND2xp5_ASAP7_75t_L g1605 ( 
.A(n_1593),
.B(n_1548),
.Y(n_1605)
);

INVx2_ASAP7_75t_L g1606 ( 
.A(n_1587),
.Y(n_1606)
);

AND2x4_ASAP7_75t_L g1607 ( 
.A(n_1590),
.B(n_1543),
.Y(n_1607)
);

BUFx2_ASAP7_75t_L g1608 ( 
.A(n_1590),
.Y(n_1608)
);

AND2x4_ASAP7_75t_L g1609 ( 
.A(n_1590),
.B(n_1543),
.Y(n_1609)
);

NAND2xp5_ASAP7_75t_L g1610 ( 
.A(n_1578),
.B(n_1555),
.Y(n_1610)
);

HB1xp67_ASAP7_75t_L g1611 ( 
.A(n_1582),
.Y(n_1611)
);

AND2x2_ASAP7_75t_L g1612 ( 
.A(n_1591),
.B(n_1543),
.Y(n_1612)
);

INVx1_ASAP7_75t_L g1613 ( 
.A(n_1580),
.Y(n_1613)
);

OR2x2_ASAP7_75t_L g1614 ( 
.A(n_1577),
.B(n_1551),
.Y(n_1614)
);

AND2x2_ASAP7_75t_L g1615 ( 
.A(n_1591),
.B(n_1551),
.Y(n_1615)
);

NOR2xp33_ASAP7_75t_L g1616 ( 
.A(n_1585),
.B(n_1542),
.Y(n_1616)
);

NAND2xp5_ASAP7_75t_L g1617 ( 
.A(n_1578),
.B(n_1555),
.Y(n_1617)
);

INVx1_ASAP7_75t_SL g1618 ( 
.A(n_1584),
.Y(n_1618)
);

OR2x2_ASAP7_75t_L g1619 ( 
.A(n_1577),
.B(n_1551),
.Y(n_1619)
);

INVx1_ASAP7_75t_L g1620 ( 
.A(n_1581),
.Y(n_1620)
);

AOI22xp33_ASAP7_75t_L g1621 ( 
.A1(n_1585),
.A2(n_1454),
.B1(n_1486),
.B2(n_1428),
.Y(n_1621)
);

BUFx3_ASAP7_75t_L g1622 ( 
.A(n_1588),
.Y(n_1622)
);

HB1xp67_ASAP7_75t_L g1623 ( 
.A(n_1582),
.Y(n_1623)
);

INVx2_ASAP7_75t_L g1624 ( 
.A(n_1587),
.Y(n_1624)
);

OR2x2_ASAP7_75t_L g1625 ( 
.A(n_1584),
.B(n_1552),
.Y(n_1625)
);

NAND2x1_ASAP7_75t_L g1626 ( 
.A(n_1592),
.B(n_1544),
.Y(n_1626)
);

INVx1_ASAP7_75t_L g1627 ( 
.A(n_1611),
.Y(n_1627)
);

NAND2xp5_ASAP7_75t_L g1628 ( 
.A(n_1616),
.B(n_1583),
.Y(n_1628)
);

OR2x2_ASAP7_75t_L g1629 ( 
.A(n_1610),
.B(n_1584),
.Y(n_1629)
);

INVx2_ASAP7_75t_L g1630 ( 
.A(n_1614),
.Y(n_1630)
);

INVxp67_ASAP7_75t_L g1631 ( 
.A(n_1616),
.Y(n_1631)
);

NAND2xp5_ASAP7_75t_L g1632 ( 
.A(n_1621),
.B(n_1583),
.Y(n_1632)
);

INVx1_ASAP7_75t_L g1633 ( 
.A(n_1611),
.Y(n_1633)
);

NAND2xp5_ASAP7_75t_L g1634 ( 
.A(n_1621),
.B(n_1582),
.Y(n_1634)
);

NOR2xp33_ASAP7_75t_L g1635 ( 
.A(n_1600),
.B(n_1428),
.Y(n_1635)
);

INVx2_ASAP7_75t_SL g1636 ( 
.A(n_1608),
.Y(n_1636)
);

NOR2xp33_ASAP7_75t_L g1637 ( 
.A(n_1600),
.B(n_1428),
.Y(n_1637)
);

INVx2_ASAP7_75t_L g1638 ( 
.A(n_1614),
.Y(n_1638)
);

AND2x2_ASAP7_75t_L g1639 ( 
.A(n_1608),
.B(n_1586),
.Y(n_1639)
);

INVx1_ASAP7_75t_L g1640 ( 
.A(n_1623),
.Y(n_1640)
);

AND2x2_ASAP7_75t_L g1641 ( 
.A(n_1608),
.B(n_1586),
.Y(n_1641)
);

OR2x2_ASAP7_75t_L g1642 ( 
.A(n_1605),
.B(n_1594),
.Y(n_1642)
);

INVx1_ASAP7_75t_L g1643 ( 
.A(n_1623),
.Y(n_1643)
);

OR2x2_ASAP7_75t_L g1644 ( 
.A(n_1605),
.B(n_1594),
.Y(n_1644)
);

NAND2xp5_ASAP7_75t_L g1645 ( 
.A(n_1610),
.B(n_1594),
.Y(n_1645)
);

NAND2xp5_ASAP7_75t_L g1646 ( 
.A(n_1617),
.B(n_1573),
.Y(n_1646)
);

INVx1_ASAP7_75t_L g1647 ( 
.A(n_1602),
.Y(n_1647)
);

NAND2xp5_ASAP7_75t_L g1648 ( 
.A(n_1617),
.B(n_1573),
.Y(n_1648)
);

NAND2xp5_ASAP7_75t_L g1649 ( 
.A(n_1618),
.B(n_1573),
.Y(n_1649)
);

OR2x2_ASAP7_75t_L g1650 ( 
.A(n_1625),
.B(n_1589),
.Y(n_1650)
);

INVx1_ASAP7_75t_L g1651 ( 
.A(n_1602),
.Y(n_1651)
);

AND2x2_ASAP7_75t_L g1652 ( 
.A(n_1622),
.B(n_1586),
.Y(n_1652)
);

OR2x6_ASAP7_75t_L g1653 ( 
.A(n_1622),
.B(n_1510),
.Y(n_1653)
);

INVx2_ASAP7_75t_SL g1654 ( 
.A(n_1622),
.Y(n_1654)
);

INVx1_ASAP7_75t_L g1655 ( 
.A(n_1602),
.Y(n_1655)
);

NAND2x1_ASAP7_75t_L g1656 ( 
.A(n_1597),
.B(n_1592),
.Y(n_1656)
);

INVx1_ASAP7_75t_L g1657 ( 
.A(n_1603),
.Y(n_1657)
);

OR2x2_ASAP7_75t_L g1658 ( 
.A(n_1625),
.B(n_1589),
.Y(n_1658)
);

AOI22xp5_ASAP7_75t_L g1659 ( 
.A1(n_1598),
.A2(n_1575),
.B1(n_1570),
.B2(n_1596),
.Y(n_1659)
);

INVx1_ASAP7_75t_L g1660 ( 
.A(n_1603),
.Y(n_1660)
);

NAND2xp5_ASAP7_75t_L g1661 ( 
.A(n_1618),
.B(n_1579),
.Y(n_1661)
);

INVx2_ASAP7_75t_L g1662 ( 
.A(n_1614),
.Y(n_1662)
);

AND2x2_ASAP7_75t_L g1663 ( 
.A(n_1622),
.B(n_1586),
.Y(n_1663)
);

NOR2xp67_ASAP7_75t_L g1664 ( 
.A(n_1597),
.B(n_1469),
.Y(n_1664)
);

INVx1_ASAP7_75t_L g1665 ( 
.A(n_1603),
.Y(n_1665)
);

INVx2_ASAP7_75t_L g1666 ( 
.A(n_1614),
.Y(n_1666)
);

OR2x2_ASAP7_75t_L g1667 ( 
.A(n_1625),
.B(n_1576),
.Y(n_1667)
);

INVx1_ASAP7_75t_L g1668 ( 
.A(n_1613),
.Y(n_1668)
);

NAND2xp5_ASAP7_75t_L g1669 ( 
.A(n_1598),
.B(n_1579),
.Y(n_1669)
);

OR2x2_ASAP7_75t_L g1670 ( 
.A(n_1642),
.B(n_1576),
.Y(n_1670)
);

INVx2_ASAP7_75t_SL g1671 ( 
.A(n_1636),
.Y(n_1671)
);

INVx1_ASAP7_75t_L g1672 ( 
.A(n_1647),
.Y(n_1672)
);

NOR2xp33_ASAP7_75t_L g1673 ( 
.A(n_1635),
.B(n_1469),
.Y(n_1673)
);

NAND2xp5_ASAP7_75t_L g1674 ( 
.A(n_1631),
.B(n_1579),
.Y(n_1674)
);

INVx1_ASAP7_75t_L g1675 ( 
.A(n_1651),
.Y(n_1675)
);

NAND2xp33_ASAP7_75t_L g1676 ( 
.A(n_1659),
.B(n_1570),
.Y(n_1676)
);

INVx2_ASAP7_75t_SL g1677 ( 
.A(n_1636),
.Y(n_1677)
);

NAND4xp25_ASAP7_75t_L g1678 ( 
.A(n_1635),
.B(n_1574),
.C(n_1575),
.D(n_1596),
.Y(n_1678)
);

INVx2_ASAP7_75t_L g1679 ( 
.A(n_1630),
.Y(n_1679)
);

NOR3xp33_ASAP7_75t_SL g1680 ( 
.A(n_1637),
.B(n_1595),
.C(n_1574),
.Y(n_1680)
);

INVx2_ASAP7_75t_L g1681 ( 
.A(n_1630),
.Y(n_1681)
);

INVx2_ASAP7_75t_L g1682 ( 
.A(n_1638),
.Y(n_1682)
);

INVx1_ASAP7_75t_L g1683 ( 
.A(n_1655),
.Y(n_1683)
);

OR2x2_ASAP7_75t_L g1684 ( 
.A(n_1644),
.B(n_1576),
.Y(n_1684)
);

AND2x2_ASAP7_75t_L g1685 ( 
.A(n_1653),
.B(n_1597),
.Y(n_1685)
);

INVx2_ASAP7_75t_L g1686 ( 
.A(n_1638),
.Y(n_1686)
);

INVx1_ASAP7_75t_L g1687 ( 
.A(n_1657),
.Y(n_1687)
);

NAND2xp5_ASAP7_75t_L g1688 ( 
.A(n_1628),
.B(n_1598),
.Y(n_1688)
);

AND2x4_ASAP7_75t_L g1689 ( 
.A(n_1664),
.B(n_1597),
.Y(n_1689)
);

INVx1_ASAP7_75t_SL g1690 ( 
.A(n_1653),
.Y(n_1690)
);

INVx1_ASAP7_75t_L g1691 ( 
.A(n_1660),
.Y(n_1691)
);

NAND2xp5_ASAP7_75t_L g1692 ( 
.A(n_1632),
.B(n_1598),
.Y(n_1692)
);

NAND2xp5_ASAP7_75t_L g1693 ( 
.A(n_1637),
.B(n_1599),
.Y(n_1693)
);

INVx1_ASAP7_75t_L g1694 ( 
.A(n_1665),
.Y(n_1694)
);

AND2x2_ASAP7_75t_SL g1695 ( 
.A(n_1634),
.B(n_1487),
.Y(n_1695)
);

INVx1_ASAP7_75t_L g1696 ( 
.A(n_1668),
.Y(n_1696)
);

AO21x1_ASAP7_75t_L g1697 ( 
.A1(n_1650),
.A2(n_1601),
.B(n_1599),
.Y(n_1697)
);

OR2x6_ASAP7_75t_L g1698 ( 
.A(n_1653),
.B(n_1487),
.Y(n_1698)
);

NAND2xp5_ASAP7_75t_L g1699 ( 
.A(n_1645),
.B(n_1599),
.Y(n_1699)
);

AND2x2_ASAP7_75t_L g1700 ( 
.A(n_1653),
.B(n_1652),
.Y(n_1700)
);

NAND2xp5_ASAP7_75t_L g1701 ( 
.A(n_1627),
.B(n_1633),
.Y(n_1701)
);

INVx1_ASAP7_75t_SL g1702 ( 
.A(n_1658),
.Y(n_1702)
);

AND2x2_ASAP7_75t_L g1703 ( 
.A(n_1652),
.B(n_1663),
.Y(n_1703)
);

AOI221x1_ASAP7_75t_L g1704 ( 
.A1(n_1640),
.A2(n_1597),
.B1(n_1471),
.B2(n_1549),
.C(n_1484),
.Y(n_1704)
);

AND2x2_ASAP7_75t_L g1705 ( 
.A(n_1663),
.B(n_1597),
.Y(n_1705)
);

INVx1_ASAP7_75t_L g1706 ( 
.A(n_1672),
.Y(n_1706)
);

OAI22xp5_ASAP7_75t_L g1707 ( 
.A1(n_1680),
.A2(n_1702),
.B1(n_1695),
.B2(n_1692),
.Y(n_1707)
);

INVxp67_ASAP7_75t_L g1708 ( 
.A(n_1701),
.Y(n_1708)
);

INVx2_ASAP7_75t_L g1709 ( 
.A(n_1671),
.Y(n_1709)
);

INVx1_ASAP7_75t_L g1710 ( 
.A(n_1672),
.Y(n_1710)
);

AND2x2_ASAP7_75t_L g1711 ( 
.A(n_1703),
.B(n_1654),
.Y(n_1711)
);

OAI21xp5_ASAP7_75t_L g1712 ( 
.A1(n_1676),
.A2(n_1595),
.B(n_1654),
.Y(n_1712)
);

AOI21xp33_ASAP7_75t_SL g1713 ( 
.A1(n_1673),
.A2(n_1458),
.B(n_1481),
.Y(n_1713)
);

AOI22xp33_ASAP7_75t_L g1714 ( 
.A1(n_1676),
.A2(n_1641),
.B1(n_1639),
.B2(n_1643),
.Y(n_1714)
);

NOR2xp33_ASAP7_75t_L g1715 ( 
.A(n_1678),
.B(n_1481),
.Y(n_1715)
);

INVx1_ASAP7_75t_L g1716 ( 
.A(n_1675),
.Y(n_1716)
);

INVx1_ASAP7_75t_L g1717 ( 
.A(n_1675),
.Y(n_1717)
);

INVxp67_ASAP7_75t_L g1718 ( 
.A(n_1671),
.Y(n_1718)
);

INVx1_ASAP7_75t_L g1719 ( 
.A(n_1683),
.Y(n_1719)
);

INVx1_ASAP7_75t_L g1720 ( 
.A(n_1683),
.Y(n_1720)
);

INVx2_ASAP7_75t_L g1721 ( 
.A(n_1677),
.Y(n_1721)
);

INVx2_ASAP7_75t_L g1722 ( 
.A(n_1677),
.Y(n_1722)
);

AND2x2_ASAP7_75t_L g1723 ( 
.A(n_1703),
.B(n_1639),
.Y(n_1723)
);

INVx1_ASAP7_75t_L g1724 ( 
.A(n_1691),
.Y(n_1724)
);

AOI322xp5_ASAP7_75t_L g1725 ( 
.A1(n_1688),
.A2(n_1646),
.A3(n_1648),
.B1(n_1649),
.B2(n_1601),
.C1(n_1599),
.C2(n_1661),
.Y(n_1725)
);

INVx1_ASAP7_75t_SL g1726 ( 
.A(n_1695),
.Y(n_1726)
);

AND2x2_ASAP7_75t_L g1727 ( 
.A(n_1700),
.B(n_1641),
.Y(n_1727)
);

NAND2xp5_ASAP7_75t_L g1728 ( 
.A(n_1693),
.B(n_1629),
.Y(n_1728)
);

NOR2xp33_ASAP7_75t_L g1729 ( 
.A(n_1690),
.B(n_1475),
.Y(n_1729)
);

AOI22xp33_ASAP7_75t_SL g1730 ( 
.A1(n_1700),
.A2(n_1601),
.B1(n_1669),
.B2(n_1492),
.Y(n_1730)
);

AOI211xp5_ASAP7_75t_L g1731 ( 
.A1(n_1697),
.A2(n_1572),
.B(n_1501),
.C(n_1496),
.Y(n_1731)
);

INVx1_ASAP7_75t_L g1732 ( 
.A(n_1706),
.Y(n_1732)
);

INVxp67_ASAP7_75t_L g1733 ( 
.A(n_1715),
.Y(n_1733)
);

NOR2xp33_ASAP7_75t_L g1734 ( 
.A(n_1713),
.B(n_1475),
.Y(n_1734)
);

OAI21xp5_ASAP7_75t_L g1735 ( 
.A1(n_1712),
.A2(n_1704),
.B(n_1572),
.Y(n_1735)
);

OAI21xp5_ASAP7_75t_L g1736 ( 
.A1(n_1707),
.A2(n_1704),
.B(n_1674),
.Y(n_1736)
);

A2O1A1Ixp33_ASAP7_75t_L g1737 ( 
.A1(n_1714),
.A2(n_1689),
.B(n_1697),
.C(n_1685),
.Y(n_1737)
);

INVx1_ASAP7_75t_L g1738 ( 
.A(n_1706),
.Y(n_1738)
);

OR2x2_ASAP7_75t_L g1739 ( 
.A(n_1728),
.B(n_1699),
.Y(n_1739)
);

NOR2x1_ASAP7_75t_L g1740 ( 
.A(n_1709),
.B(n_1698),
.Y(n_1740)
);

AO22x1_ASAP7_75t_L g1741 ( 
.A1(n_1709),
.A2(n_1689),
.B1(n_1685),
.B2(n_1681),
.Y(n_1741)
);

OAI22xp33_ASAP7_75t_L g1742 ( 
.A1(n_1726),
.A2(n_1698),
.B1(n_1588),
.B2(n_1656),
.Y(n_1742)
);

NAND2xp5_ASAP7_75t_L g1743 ( 
.A(n_1718),
.B(n_1687),
.Y(n_1743)
);

NAND3xp33_ASAP7_75t_L g1744 ( 
.A(n_1708),
.B(n_1694),
.C(n_1691),
.Y(n_1744)
);

AOI221xp5_ASAP7_75t_L g1745 ( 
.A1(n_1721),
.A2(n_1722),
.B1(n_1710),
.B2(n_1719),
.C(n_1720),
.Y(n_1745)
);

INVx1_ASAP7_75t_SL g1746 ( 
.A(n_1711),
.Y(n_1746)
);

AND2x2_ASAP7_75t_L g1747 ( 
.A(n_1727),
.B(n_1689),
.Y(n_1747)
);

NOR2x1_ASAP7_75t_L g1748 ( 
.A(n_1721),
.B(n_1698),
.Y(n_1748)
);

INVx1_ASAP7_75t_L g1749 ( 
.A(n_1710),
.Y(n_1749)
);

AND2x2_ASAP7_75t_L g1750 ( 
.A(n_1727),
.B(n_1705),
.Y(n_1750)
);

INVx1_ASAP7_75t_L g1751 ( 
.A(n_1716),
.Y(n_1751)
);

INVx1_ASAP7_75t_L g1752 ( 
.A(n_1732),
.Y(n_1752)
);

INVx2_ASAP7_75t_L g1753 ( 
.A(n_1750),
.Y(n_1753)
);

AOI211xp5_ASAP7_75t_L g1754 ( 
.A1(n_1737),
.A2(n_1713),
.B(n_1729),
.C(n_1722),
.Y(n_1754)
);

OAI22xp33_ASAP7_75t_SL g1755 ( 
.A1(n_1735),
.A2(n_1698),
.B1(n_1719),
.B2(n_1717),
.Y(n_1755)
);

AOI21xp5_ASAP7_75t_SL g1756 ( 
.A1(n_1734),
.A2(n_1717),
.B(n_1716),
.Y(n_1756)
);

NAND2xp5_ASAP7_75t_L g1757 ( 
.A(n_1746),
.B(n_1720),
.Y(n_1757)
);

NAND2xp5_ASAP7_75t_L g1758 ( 
.A(n_1747),
.B(n_1711),
.Y(n_1758)
);

OR2x2_ASAP7_75t_L g1759 ( 
.A(n_1739),
.B(n_1743),
.Y(n_1759)
);

OAI211xp5_ASAP7_75t_L g1760 ( 
.A1(n_1736),
.A2(n_1725),
.B(n_1731),
.C(n_1730),
.Y(n_1760)
);

NAND2xp5_ASAP7_75t_L g1761 ( 
.A(n_1733),
.B(n_1723),
.Y(n_1761)
);

OAI22xp5_ASAP7_75t_L g1762 ( 
.A1(n_1736),
.A2(n_1731),
.B1(n_1723),
.B2(n_1588),
.Y(n_1762)
);

NOR4xp25_ASAP7_75t_L g1763 ( 
.A(n_1760),
.B(n_1745),
.C(n_1749),
.D(n_1738),
.Y(n_1763)
);

AND3x1_ASAP7_75t_L g1764 ( 
.A(n_1754),
.B(n_1753),
.C(n_1748),
.Y(n_1764)
);

NAND4xp25_ASAP7_75t_L g1765 ( 
.A(n_1761),
.B(n_1758),
.C(n_1756),
.D(n_1759),
.Y(n_1765)
);

NAND2xp5_ASAP7_75t_L g1766 ( 
.A(n_1757),
.B(n_1741),
.Y(n_1766)
);

OAI32xp33_ASAP7_75t_L g1767 ( 
.A1(n_1762),
.A2(n_1735),
.A3(n_1744),
.B1(n_1751),
.B2(n_1724),
.Y(n_1767)
);

INVx2_ASAP7_75t_L g1768 ( 
.A(n_1757),
.Y(n_1768)
);

INVx1_ASAP7_75t_L g1769 ( 
.A(n_1752),
.Y(n_1769)
);

NAND2xp33_ASAP7_75t_SL g1770 ( 
.A(n_1755),
.B(n_1724),
.Y(n_1770)
);

NAND3xp33_ASAP7_75t_SL g1771 ( 
.A(n_1760),
.B(n_1725),
.C(n_1740),
.Y(n_1771)
);

AOI21xp5_ASAP7_75t_L g1772 ( 
.A1(n_1756),
.A2(n_1742),
.B(n_1696),
.Y(n_1772)
);

AOI22xp33_ASAP7_75t_L g1773 ( 
.A1(n_1771),
.A2(n_1686),
.B1(n_1682),
.B2(n_1681),
.Y(n_1773)
);

A2O1A1Ixp33_ASAP7_75t_L g1774 ( 
.A1(n_1770),
.A2(n_1772),
.B(n_1766),
.C(n_1767),
.Y(n_1774)
);

AOI22xp5_ASAP7_75t_L g1775 ( 
.A1(n_1764),
.A2(n_1705),
.B1(n_1686),
.B2(n_1679),
.Y(n_1775)
);

NAND2xp5_ASAP7_75t_L g1776 ( 
.A(n_1763),
.B(n_1694),
.Y(n_1776)
);

NAND3xp33_ASAP7_75t_SL g1777 ( 
.A(n_1772),
.B(n_1768),
.C(n_1769),
.Y(n_1777)
);

AOI321xp33_ASAP7_75t_L g1778 ( 
.A1(n_1774),
.A2(n_1765),
.A3(n_1682),
.B1(n_1679),
.B2(n_1696),
.C(n_1684),
.Y(n_1778)
);

O2A1O1Ixp33_ASAP7_75t_L g1779 ( 
.A1(n_1776),
.A2(n_1684),
.B(n_1670),
.C(n_1662),
.Y(n_1779)
);

AOI221xp5_ASAP7_75t_L g1780 ( 
.A1(n_1777),
.A2(n_1662),
.B1(n_1666),
.B2(n_1670),
.C(n_1606),
.Y(n_1780)
);

NAND3xp33_ASAP7_75t_SL g1781 ( 
.A(n_1775),
.B(n_1629),
.C(n_1626),
.Y(n_1781)
);

OAI211xp5_ASAP7_75t_SL g1782 ( 
.A1(n_1773),
.A2(n_1666),
.B(n_1667),
.C(n_1496),
.Y(n_1782)
);

NAND2xp5_ASAP7_75t_L g1783 ( 
.A(n_1774),
.B(n_1601),
.Y(n_1783)
);

AOI22xp5_ASAP7_75t_L g1784 ( 
.A1(n_1783),
.A2(n_1511),
.B1(n_1475),
.B2(n_1483),
.Y(n_1784)
);

INVx1_ASAP7_75t_L g1785 ( 
.A(n_1778),
.Y(n_1785)
);

XNOR2x1_ASAP7_75t_L g1786 ( 
.A(n_1782),
.B(n_1511),
.Y(n_1786)
);

OAI22xp5_ASAP7_75t_L g1787 ( 
.A1(n_1780),
.A2(n_1667),
.B1(n_1626),
.B2(n_1619),
.Y(n_1787)
);

INVxp33_ASAP7_75t_SL g1788 ( 
.A(n_1781),
.Y(n_1788)
);

AND3x1_ASAP7_75t_L g1789 ( 
.A(n_1785),
.B(n_1779),
.C(n_1592),
.Y(n_1789)
);

AOI21xp5_ASAP7_75t_L g1790 ( 
.A1(n_1788),
.A2(n_1619),
.B(n_1613),
.Y(n_1790)
);

NOR3xp33_ASAP7_75t_L g1791 ( 
.A(n_1784),
.B(n_1568),
.C(n_1493),
.Y(n_1791)
);

OAI22xp5_ASAP7_75t_L g1792 ( 
.A1(n_1789),
.A2(n_1786),
.B1(n_1787),
.B2(n_1619),
.Y(n_1792)
);

INVx2_ASAP7_75t_L g1793 ( 
.A(n_1792),
.Y(n_1793)
);

AOI22xp5_ASAP7_75t_L g1794 ( 
.A1(n_1793),
.A2(n_1790),
.B1(n_1791),
.B2(n_1607),
.Y(n_1794)
);

XOR2xp5_ASAP7_75t_L g1795 ( 
.A(n_1793),
.B(n_1490),
.Y(n_1795)
);

BUFx2_ASAP7_75t_L g1796 ( 
.A(n_1795),
.Y(n_1796)
);

OAI22x1_ASAP7_75t_SL g1797 ( 
.A1(n_1794),
.A2(n_1539),
.B1(n_1620),
.B2(n_1613),
.Y(n_1797)
);

OAI22xp5_ASAP7_75t_L g1798 ( 
.A1(n_1796),
.A2(n_1619),
.B1(n_1626),
.B2(n_1615),
.Y(n_1798)
);

INVx1_ASAP7_75t_L g1799 ( 
.A(n_1797),
.Y(n_1799)
);

NAND2xp5_ASAP7_75t_SL g1800 ( 
.A(n_1799),
.B(n_1607),
.Y(n_1800)
);

NAND2xp5_ASAP7_75t_L g1801 ( 
.A(n_1800),
.B(n_1798),
.Y(n_1801)
);

XNOR2xp5_ASAP7_75t_L g1802 ( 
.A(n_1801),
.B(n_1490),
.Y(n_1802)
);

OAI221xp5_ASAP7_75t_R g1803 ( 
.A1(n_1802),
.A2(n_1612),
.B1(n_1615),
.B2(n_1604),
.C(n_1609),
.Y(n_1803)
);

AOI211xp5_ASAP7_75t_L g1804 ( 
.A1(n_1803),
.A2(n_1485),
.B(n_1482),
.C(n_1624),
.Y(n_1804)
);


endmodule