module fake_jpeg_17988_n_123 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_123);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_123;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_96;

INVx8_ASAP7_75t_L g14 ( 
.A(n_3),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_8),
.Y(n_15)
);

INVx2_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_SL g17 ( 
.A(n_13),
.B(n_4),
.Y(n_17)
);

INVx4_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

BUFx12_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_1),
.Y(n_21)
);

INVx6_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

INVx11_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

INVx6_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_16),
.B(n_24),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_SL g44 ( 
.A(n_28),
.B(n_29),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_24),
.B(n_0),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_16),
.B(n_0),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_SL g50 ( 
.A(n_30),
.B(n_32),
.Y(n_50)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_23),
.Y(n_31)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_31),
.Y(n_48)
);

AND2x2_ASAP7_75t_L g32 ( 
.A(n_17),
.B(n_2),
.Y(n_32)
);

NAND2x1_ASAP7_75t_SL g33 ( 
.A(n_18),
.B(n_2),
.Y(n_33)
);

OR2x2_ASAP7_75t_L g59 ( 
.A(n_33),
.B(n_19),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_21),
.B(n_3),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_34),
.B(n_35),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_21),
.B(n_4),
.Y(n_35)
);

INVx5_ASAP7_75t_L g36 ( 
.A(n_27),
.Y(n_36)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_36),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_L g37 ( 
.A1(n_22),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_L g42 ( 
.A1(n_37),
.A2(n_38),
.B1(n_14),
.B2(n_15),
.Y(n_42)
);

AO22x2_ASAP7_75t_L g38 ( 
.A1(n_27),
.A2(n_5),
.B1(n_7),
.B2(n_9),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_18),
.B(n_23),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_39),
.B(n_41),
.Y(n_47)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_22),
.Y(n_40)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_40),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_14),
.B(n_7),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_L g76 ( 
.A1(n_42),
.A2(n_19),
.B1(n_54),
.B2(n_49),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_34),
.B(n_15),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_43),
.B(n_45),
.Y(n_75)
);

INVx1_ASAP7_75t_SL g45 ( 
.A(n_33),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_35),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_49),
.B(n_61),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_38),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_51),
.Y(n_73)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_53),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g54 ( 
.A1(n_38),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_54),
.A2(n_36),
.B1(n_12),
.B2(n_26),
.Y(n_71)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_55),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_30),
.B(n_25),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_56),
.B(n_60),
.Y(n_70)
);

CKINVDCx14_ASAP7_75t_R g57 ( 
.A(n_29),
.Y(n_57)
);

INVx13_ASAP7_75t_L g80 ( 
.A(n_57),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_SL g58 ( 
.A(n_32),
.B(n_20),
.Y(n_58)
);

CKINVDCx16_ASAP7_75t_R g79 ( 
.A(n_58),
.Y(n_79)
);

OAI21xp5_ASAP7_75t_L g66 ( 
.A1(n_59),
.A2(n_64),
.B(n_31),
.Y(n_66)
);

INVx13_ASAP7_75t_L g60 ( 
.A(n_33),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_32),
.B(n_25),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_28),
.B(n_20),
.Y(n_62)
);

XNOR2xp5_ASAP7_75t_L g68 ( 
.A(n_62),
.B(n_38),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_38),
.A2(n_26),
.B1(n_19),
.B2(n_12),
.Y(n_63)
);

AOI21xp5_ASAP7_75t_L g72 ( 
.A1(n_63),
.A2(n_19),
.B(n_42),
.Y(n_72)
);

INVxp67_ASAP7_75t_L g64 ( 
.A(n_41),
.Y(n_64)
);

XNOR2xp5_ASAP7_75t_SL g82 ( 
.A(n_66),
.B(n_68),
.Y(n_82)
);

XOR2xp5_ASAP7_75t_L g67 ( 
.A(n_47),
.B(n_38),
.Y(n_67)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_67),
.B(n_77),
.C(n_44),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_71),
.A2(n_72),
.B1(n_76),
.B2(n_78),
.Y(n_86)
);

AOI21xp5_ASAP7_75t_L g77 ( 
.A1(n_45),
.A2(n_60),
.B(n_62),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_51),
.A2(n_55),
.B1(n_47),
.B2(n_46),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_78),
.B(n_46),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_83),
.B(n_88),
.Y(n_99)
);

XOR2xp5_ASAP7_75t_L g84 ( 
.A(n_77),
.B(n_56),
.Y(n_84)
);

XOR2xp5_ASAP7_75t_L g96 ( 
.A(n_84),
.B(n_87),
.Y(n_96)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_69),
.Y(n_85)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_85),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_69),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_74),
.B(n_44),
.Y(n_89)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_89),
.Y(n_101)
);

XOR2xp5_ASAP7_75t_L g90 ( 
.A(n_67),
.B(n_50),
.Y(n_90)
);

XOR2xp5_ASAP7_75t_L g102 ( 
.A(n_90),
.B(n_93),
.Y(n_102)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_75),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_91),
.Y(n_98)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_74),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_92),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_70),
.B(n_68),
.C(n_66),
.Y(n_93)
);

XOR2xp5_ASAP7_75t_L g94 ( 
.A(n_70),
.B(n_50),
.Y(n_94)
);

XOR2xp5_ASAP7_75t_L g104 ( 
.A(n_94),
.B(n_81),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_76),
.A2(n_64),
.B1(n_65),
.B2(n_53),
.Y(n_95)
);

AOI21xp5_ASAP7_75t_L g103 ( 
.A1(n_95),
.A2(n_65),
.B(n_73),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_L g107 ( 
.A1(n_103),
.A2(n_105),
.B(n_59),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_104),
.B(n_82),
.C(n_87),
.Y(n_110)
);

AOI21xp5_ASAP7_75t_L g105 ( 
.A1(n_84),
.A2(n_73),
.B(n_72),
.Y(n_105)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_97),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_106),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_107),
.A2(n_108),
.B1(n_110),
.B2(n_111),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_100),
.B(n_80),
.Y(n_108)
);

AOI21xp5_ASAP7_75t_L g109 ( 
.A1(n_96),
.A2(n_86),
.B(n_90),
.Y(n_109)
);

AOI21xp5_ASAP7_75t_L g116 ( 
.A1(n_109),
.A2(n_112),
.B(n_104),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_98),
.B(n_80),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_99),
.B(n_48),
.Y(n_112)
);

AOI21x1_ASAP7_75t_SL g115 ( 
.A1(n_107),
.A2(n_105),
.B(n_82),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_115),
.B(n_117),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_116),
.B(n_102),
.Y(n_118)
);

AOI322xp5_ASAP7_75t_L g117 ( 
.A1(n_110),
.A2(n_96),
.A3(n_93),
.B1(n_102),
.B2(n_101),
.C1(n_94),
.C2(n_81),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_L g122 ( 
.A1(n_118),
.A2(n_120),
.B(n_79),
.Y(n_122)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_113),
.Y(n_120)
);

AOI322xp5_ASAP7_75t_L g121 ( 
.A1(n_119),
.A2(n_114),
.A3(n_117),
.B1(n_71),
.B2(n_79),
.C1(n_52),
.C2(n_48),
.Y(n_121)
);

AOI31xp33_ASAP7_75t_L g123 ( 
.A1(n_121),
.A2(n_122),
.A3(n_120),
.B(n_52),
.Y(n_123)
);


endmodule