module real_jpeg_7086_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_80;
wire n_30;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_216;
wire n_202;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_288;
wire n_83;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_312;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

INVx8_ASAP7_75t_L g60 ( 
.A(n_0),
.Y(n_60)
);

AND2x2_ASAP7_75t_L g54 ( 
.A(n_1),
.B(n_55),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_1),
.B(n_73),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_1),
.B(n_114),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_1),
.B(n_139),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_1),
.B(n_205),
.Y(n_204)
);

AND2x2_ASAP7_75t_L g221 ( 
.A(n_1),
.B(n_222),
.Y(n_221)
);

AND2x2_ASAP7_75t_L g247 ( 
.A(n_1),
.B(n_248),
.Y(n_247)
);

AND2x2_ASAP7_75t_L g267 ( 
.A(n_1),
.B(n_268),
.Y(n_267)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_2),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_2),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_2),
.Y(n_129)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_3),
.Y(n_37)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_3),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g170 ( 
.A(n_3),
.Y(n_170)
);

AND2x2_ASAP7_75t_L g44 ( 
.A(n_4),
.B(n_45),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_4),
.B(n_65),
.Y(n_64)
);

AND2x2_ASAP7_75t_SL g89 ( 
.A(n_4),
.B(n_90),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_4),
.B(n_103),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_4),
.B(n_132),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_5),
.B(n_36),
.Y(n_35)
);

AND2x2_ASAP7_75t_L g49 ( 
.A(n_5),
.B(n_50),
.Y(n_49)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_5),
.B(n_77),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_5),
.B(n_100),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g61 ( 
.A(n_6),
.B(n_62),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_6),
.B(n_71),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_6),
.B(n_94),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_6),
.B(n_152),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_6),
.B(n_169),
.Y(n_168)
);

AND2x2_ASAP7_75t_L g240 ( 
.A(n_6),
.B(n_123),
.Y(n_240)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

INVx8_ASAP7_75t_L g51 ( 
.A(n_8),
.Y(n_51)
);

BUFx5_ASAP7_75t_L g123 ( 
.A(n_8),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_8),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_8),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g214 ( 
.A(n_8),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_9),
.B(n_87),
.Y(n_86)
);

AND2x2_ASAP7_75t_SL g180 ( 
.A(n_9),
.B(n_181),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_9),
.B(n_209),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_9),
.B(n_212),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_9),
.B(n_233),
.Y(n_232)
);

AND2x2_ASAP7_75t_L g246 ( 
.A(n_9),
.B(n_71),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_9),
.B(n_273),
.Y(n_272)
);

AND2x2_ASAP7_75t_L g122 ( 
.A(n_10),
.B(n_123),
.Y(n_122)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_11),
.Y(n_40)
);

BUFx5_ASAP7_75t_L g73 ( 
.A(n_11),
.Y(n_73)
);

INVx8_ASAP7_75t_L g84 ( 
.A(n_12),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g38 ( 
.A(n_13),
.B(n_39),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_13),
.B(n_129),
.Y(n_128)
);

AND2x2_ASAP7_75t_L g174 ( 
.A(n_13),
.B(n_175),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_13),
.B(n_201),
.Y(n_200)
);

AND2x2_ASAP7_75t_L g229 ( 
.A(n_13),
.B(n_230),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_SL g243 ( 
.A(n_13),
.B(n_244),
.Y(n_243)
);

AND2x2_ASAP7_75t_L g276 ( 
.A(n_13),
.B(n_30),
.Y(n_276)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

AND2x2_ASAP7_75t_L g56 ( 
.A(n_14),
.B(n_57),
.Y(n_56)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_14),
.B(n_82),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_14),
.B(n_106),
.Y(n_105)
);

AND2x2_ASAP7_75t_L g223 ( 
.A(n_14),
.B(n_224),
.Y(n_223)
);

AND2x2_ASAP7_75t_L g239 ( 
.A(n_14),
.B(n_134),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_15),
.B(n_134),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_15),
.B(n_137),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_15),
.B(n_148),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_16),
.B(n_118),
.Y(n_117)
);

AND2x2_ASAP7_75t_SL g131 ( 
.A(n_16),
.B(n_132),
.Y(n_131)
);

BUFx5_ASAP7_75t_L g62 ( 
.A(n_17),
.Y(n_62)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_17),
.Y(n_80)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_17),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_191),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_190),
.Y(n_19)
);

INVxp67_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_SL g21 ( 
.A(n_22),
.B(n_160),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_22),
.B(n_160),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_96),
.Y(n_22)
);

MAJIxp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_63),
.C(n_74),
.Y(n_23)
);

XNOR2xp5_ASAP7_75t_SL g162 ( 
.A(n_24),
.B(n_163),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_42),
.C(n_52),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_25),
.A2(n_26),
.B1(n_301),
.B2(n_302),
.Y(n_300)
);

INVx1_ASAP7_75t_SL g25 ( 
.A(n_26),
.Y(n_25)
);

XNOR2xp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_33),
.Y(n_26)
);

MAJx2_ASAP7_75t_L g141 ( 
.A(n_27),
.B(n_34),
.C(n_41),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_29),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_28),
.B(n_260),
.Y(n_259)
);

INVx5_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_32),
.Y(n_55)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_32),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g33 ( 
.A1(n_34),
.A2(n_35),
.B1(n_38),
.B2(n_41),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

BUFx5_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g120 ( 
.A(n_37),
.Y(n_120)
);

BUFx8_ASAP7_75t_L g134 ( 
.A(n_37),
.Y(n_134)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_38),
.Y(n_41)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_40),
.Y(n_107)
);

INVx5_ASAP7_75t_L g181 ( 
.A(n_40),
.Y(n_181)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

XNOR2xp5_ASAP7_75t_L g302 ( 
.A(n_43),
.B(n_53),
.Y(n_302)
);

AND2x2_ASAP7_75t_L g43 ( 
.A(n_44),
.B(n_49),
.Y(n_43)
);

XNOR2xp5_ASAP7_75t_L g291 ( 
.A(n_44),
.B(n_49),
.Y(n_291)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_46),
.Y(n_222)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx5_ASAP7_75t_L g203 ( 
.A(n_47),
.Y(n_203)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_51),
.Y(n_207)
);

BUFx6f_ASAP7_75t_L g225 ( 
.A(n_51),
.Y(n_225)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

MAJx2_ASAP7_75t_L g53 ( 
.A(n_54),
.B(n_56),
.C(n_61),
.Y(n_53)
);

XNOR2xp5_ASAP7_75t_L g288 ( 
.A(n_54),
.B(n_61),
.Y(n_288)
);

XOR2xp5_ASAP7_75t_L g287 ( 
.A(n_56),
.B(n_288),
.Y(n_287)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx6_ASAP7_75t_L g244 ( 
.A(n_58),
.Y(n_244)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g233 ( 
.A(n_59),
.Y(n_233)
);

BUFx6f_ASAP7_75t_L g270 ( 
.A(n_59),
.Y(n_270)
);

INVx11_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_60),
.Y(n_68)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_60),
.Y(n_95)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_60),
.Y(n_100)
);

INVx4_ASAP7_75t_SL g260 ( 
.A(n_62),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g163 ( 
.A(n_63),
.B(n_74),
.Y(n_163)
);

XOR2xp5_ASAP7_75t_L g63 ( 
.A(n_64),
.B(n_69),
.Y(n_63)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_64),
.B(n_70),
.C(n_72),
.Y(n_110)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

XNOR2xp5_ASAP7_75t_L g69 ( 
.A(n_70),
.B(n_72),
.Y(n_69)
);

INVx6_ASAP7_75t_L g104 ( 
.A(n_71),
.Y(n_104)
);

XNOR2xp5_ASAP7_75t_L g74 ( 
.A(n_75),
.B(n_85),
.Y(n_74)
);

XOR2xp5_ASAP7_75t_L g75 ( 
.A(n_76),
.B(n_81),
.Y(n_75)
);

MAJx2_ASAP7_75t_L g143 ( 
.A(n_76),
.B(n_81),
.C(n_144),
.Y(n_143)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_80),
.Y(n_91)
);

INVx5_ASAP7_75t_L g230 ( 
.A(n_80),
.Y(n_230)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

BUFx5_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_84),
.Y(n_140)
);

INVx6_ASAP7_75t_L g155 ( 
.A(n_84),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g178 ( 
.A(n_84),
.Y(n_178)
);

INVx3_ASAP7_75t_L g275 ( 
.A(n_84),
.Y(n_275)
);

INVx1_ASAP7_75t_SL g144 ( 
.A(n_85),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_86),
.B(n_89),
.C(n_92),
.Y(n_85)
);

XOR2xp5_ASAP7_75t_L g184 ( 
.A(n_86),
.B(n_185),
.Y(n_184)
);

INVx6_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_89),
.A2(n_92),
.B1(n_93),
.B2(n_186),
.Y(n_185)
);

INVx1_ASAP7_75t_SL g186 ( 
.A(n_89),
.Y(n_186)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

BUFx3_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

XOR2xp5_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_124),
.Y(n_96)
);

XNOR2xp5_ASAP7_75t_L g97 ( 
.A(n_98),
.B(n_108),
.Y(n_97)
);

XNOR2xp5_ASAP7_75t_SL g98 ( 
.A(n_99),
.B(n_101),
.Y(n_98)
);

XNOR2xp5_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_105),
.Y(n_101)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx6_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_109),
.A2(n_110),
.B1(n_111),
.B2(n_112),
.Y(n_108)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

XNOR2xp5_ASAP7_75t_L g112 ( 
.A(n_113),
.B(n_115),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_116),
.A2(n_117),
.B1(n_121),
.B2(n_122),
.Y(n_115)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx5_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

XOR2xp5_ASAP7_75t_L g124 ( 
.A(n_125),
.B(n_142),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_135),
.C(n_141),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_126),
.A2(n_127),
.B1(n_188),
.B2(n_189),
.Y(n_187)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

XNOR2xp5_ASAP7_75t_SL g127 ( 
.A(n_128),
.B(n_130),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_128),
.B(n_131),
.C(n_157),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_133),
.Y(n_130)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_133),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_L g182 ( 
.A1(n_135),
.A2(n_136),
.B(n_138),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g188 ( 
.A(n_135),
.B(n_141),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_136),
.B(n_138),
.Y(n_135)
);

INVx6_ASAP7_75t_SL g139 ( 
.A(n_140),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_L g142 ( 
.A1(n_143),
.A2(n_145),
.B1(n_158),
.B2(n_159),
.Y(n_142)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_143),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_145),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_L g145 ( 
.A(n_146),
.B(n_156),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_151),
.Y(n_146)
);

INVx4_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

INVx3_ASAP7_75t_L g209 ( 
.A(n_149),
.Y(n_209)
);

BUFx6f_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

BUFx5_ASAP7_75t_L g249 ( 
.A(n_150),
.Y(n_249)
);

INVx5_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

INVx3_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_161),
.B(n_164),
.C(n_187),
.Y(n_160)
);

INVxp67_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_SL g310 ( 
.A(n_162),
.B(n_311),
.Y(n_310)
);

XOR2xp5_ASAP7_75t_L g311 ( 
.A(n_164),
.B(n_187),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_165),
.B(n_182),
.C(n_183),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_SL g303 ( 
.A(n_165),
.B(n_304),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_173),
.C(n_179),
.Y(n_165)
);

XNOR2x1_ASAP7_75t_SL g283 ( 
.A(n_166),
.B(n_284),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_167),
.B(n_171),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_167),
.A2(n_168),
.B1(n_171),
.B2(n_172),
.Y(n_261)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

XNOR2x1_ASAP7_75t_SL g284 ( 
.A(n_174),
.B(n_180),
.Y(n_284)
);

INVx4_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

INVx3_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

INVx4_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

CKINVDCx14_ASAP7_75t_R g179 ( 
.A(n_180),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_182),
.A2(n_183),
.B1(n_184),
.B2(n_305),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_182),
.Y(n_305)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_188),
.Y(n_189)
);

AOI21x1_ASAP7_75t_L g191 ( 
.A1(n_192),
.A2(n_309),
.B(n_313),
.Y(n_191)
);

OAI21x1_ASAP7_75t_L g192 ( 
.A1(n_193),
.A2(n_296),
.B(n_308),
.Y(n_192)
);

AOI21xp5_ASAP7_75t_L g193 ( 
.A1(n_194),
.A2(n_280),
.B(n_295),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_L g194 ( 
.A1(n_195),
.A2(n_252),
.B(n_279),
.Y(n_194)
);

AOI21xp5_ASAP7_75t_L g195 ( 
.A1(n_196),
.A2(n_235),
.B(n_251),
.Y(n_195)
);

OAI21xp5_ASAP7_75t_L g196 ( 
.A1(n_197),
.A2(n_216),
.B(n_234),
.Y(n_196)
);

AOI21xp5_ASAP7_75t_L g197 ( 
.A1(n_198),
.A2(n_210),
.B(n_215),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_199),
.B(n_208),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_199),
.B(n_208),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_L g199 ( 
.A(n_200),
.B(n_204),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_200),
.B(n_211),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_200),
.B(n_204),
.Y(n_217)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

INVx3_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

INVx4_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

INVx4_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

INVx4_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_217),
.B(n_218),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_217),
.B(n_218),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_219),
.A2(n_220),
.B1(n_226),
.B2(n_227),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_219),
.B(n_229),
.C(n_231),
.Y(n_250)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_SL g220 ( 
.A(n_221),
.B(n_223),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_221),
.B(n_223),
.Y(n_241)
);

INVx8_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_228),
.A2(n_229),
.B1(n_231),
.B2(n_232),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_236),
.B(n_250),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_236),
.B(n_250),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_237),
.B(n_242),
.Y(n_236)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_238),
.B(n_241),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_238),
.B(n_241),
.C(n_254),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_239),
.B(n_240),
.Y(n_238)
);

AND2x2_ASAP7_75t_L g257 ( 
.A(n_239),
.B(n_240),
.Y(n_257)
);

INVxp67_ASAP7_75t_L g254 ( 
.A(n_242),
.Y(n_254)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_243),
.B(n_245),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_243),
.B(n_264),
.C(n_265),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_246),
.B(n_247),
.Y(n_245)
);

INVxp67_ASAP7_75t_L g264 ( 
.A(n_246),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_247),
.Y(n_265)
);

INVx8_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_253),
.B(n_255),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_253),
.B(n_255),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_256),
.B(n_262),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_256),
.B(n_263),
.C(n_266),
.Y(n_294)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_257),
.B(n_258),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_257),
.B(n_259),
.C(n_261),
.Y(n_285)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_259),
.B(n_261),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_263),
.B(n_266),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_L g266 ( 
.A(n_267),
.B(n_271),
.Y(n_266)
);

MAJx2_ASAP7_75t_L g293 ( 
.A(n_267),
.B(n_276),
.C(n_277),
.Y(n_293)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

INVx4_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_272),
.A2(n_276),
.B1(n_277),
.B2(n_278),
.Y(n_271)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_272),
.Y(n_277)
);

INVx6_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

INVx4_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

INVx1_ASAP7_75t_SL g278 ( 
.A(n_276),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_SL g280 ( 
.A(n_281),
.B(n_294),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_281),
.B(n_294),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_SL g281 ( 
.A(n_282),
.B(n_286),
.Y(n_281)
);

XOR2xp5_ASAP7_75t_L g282 ( 
.A(n_283),
.B(n_285),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_283),
.B(n_285),
.C(n_307),
.Y(n_306)
);

INVxp67_ASAP7_75t_L g307 ( 
.A(n_286),
.Y(n_307)
);

XOR2xp5_ASAP7_75t_L g286 ( 
.A(n_287),
.B(n_289),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_287),
.B(n_291),
.C(n_292),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_290),
.A2(n_291),
.B1(n_292),
.B2(n_293),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

INVx1_ASAP7_75t_SL g292 ( 
.A(n_293),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_SL g296 ( 
.A(n_297),
.B(n_306),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_297),
.B(n_306),
.Y(n_308)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_298),
.B(n_303),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_L g298 ( 
.A(n_299),
.B(n_300),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_299),
.B(n_300),
.C(n_303),
.Y(n_312)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_302),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_SL g309 ( 
.A(n_310),
.B(n_312),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_310),
.B(n_312),
.Y(n_313)
);


endmodule