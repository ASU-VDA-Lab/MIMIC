module fake_jpeg_9192_n_322 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_322);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_322;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_256;
wire n_221;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx5p33_ASAP7_75t_R g16 ( 
.A(n_10),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_14),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_7),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

INVx8_ASAP7_75t_SL g22 ( 
.A(n_1),
.Y(n_22)
);

INVxp67_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_1),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_6),
.Y(n_25)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_0),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_6),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_12),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_10),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_20),
.Y(n_34)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_34),
.Y(n_48)
);

CKINVDCx16_ASAP7_75t_R g35 ( 
.A(n_22),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_35),
.B(n_37),
.Y(n_61)
);

BUFx16f_ASAP7_75t_L g36 ( 
.A(n_22),
.Y(n_36)
);

INVx13_ASAP7_75t_L g49 ( 
.A(n_36),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_16),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_16),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_SL g46 ( 
.A(n_38),
.B(n_16),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_20),
.Y(n_39)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_39),
.Y(n_45)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_19),
.Y(n_40)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_40),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_20),
.Y(n_41)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_41),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_20),
.Y(n_42)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_42),
.Y(n_54)
);

INVxp67_ASAP7_75t_L g43 ( 
.A(n_23),
.Y(n_43)
);

CKINVDCx14_ASAP7_75t_R g58 ( 
.A(n_43),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_SL g76 ( 
.A(n_46),
.B(n_51),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_40),
.A2(n_32),
.B1(n_26),
.B2(n_17),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g65 ( 
.A1(n_47),
.A2(n_35),
.B1(n_26),
.B2(n_17),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_34),
.B(n_32),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_50),
.B(n_60),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_SL g51 ( 
.A(n_37),
.B(n_17),
.Y(n_51)
);

OR2x2_ASAP7_75t_L g52 ( 
.A(n_36),
.B(n_33),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_52),
.B(n_28),
.Y(n_80)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_36),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_53),
.B(n_55),
.Y(n_62)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_36),
.Y(n_55)
);

BUFx24_ASAP7_75t_L g57 ( 
.A(n_39),
.Y(n_57)
);

BUFx12f_ASAP7_75t_L g72 ( 
.A(n_57),
.Y(n_72)
);

OAI22xp33_ASAP7_75t_L g59 ( 
.A1(n_40),
.A2(n_26),
.B1(n_32),
.B2(n_31),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_59),
.A2(n_44),
.B1(n_48),
.B2(n_28),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_34),
.B(n_20),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_57),
.Y(n_63)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_63),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_L g108 ( 
.A1(n_65),
.A2(n_78),
.B1(n_45),
.B2(n_49),
.Y(n_108)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_51),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_66),
.B(n_69),
.Y(n_107)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_56),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_67),
.B(n_85),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_48),
.Y(n_68)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_68),
.Y(n_103)
);

INVx1_ASAP7_75t_SL g69 ( 
.A(n_60),
.Y(n_69)
);

CKINVDCx16_ASAP7_75t_R g70 ( 
.A(n_61),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_70),
.B(n_81),
.Y(n_110)
);

OA22x2_ASAP7_75t_L g71 ( 
.A1(n_56),
.A2(n_47),
.B1(n_45),
.B2(n_50),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_71),
.A2(n_75),
.B1(n_79),
.B2(n_87),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_48),
.Y(n_73)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_73),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g74 ( 
.A(n_50),
.B(n_39),
.C(n_38),
.Y(n_74)
);

AND2x2_ASAP7_75t_L g98 ( 
.A(n_74),
.B(n_80),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_60),
.A2(n_19),
.B1(n_21),
.B2(n_27),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_53),
.A2(n_25),
.B1(n_33),
.B2(n_18),
.Y(n_77)
);

OAI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_77),
.A2(n_84),
.B1(n_18),
.B2(n_29),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_44),
.A2(n_28),
.B1(n_24),
.B2(n_25),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_48),
.Y(n_81)
);

AND2x2_ASAP7_75t_L g82 ( 
.A(n_49),
.B(n_0),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_82),
.B(n_89),
.Y(n_99)
);

BUFx12f_ASAP7_75t_L g83 ( 
.A(n_57),
.Y(n_83)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_83),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_53),
.A2(n_25),
.B1(n_33),
.B2(n_18),
.Y(n_84)
);

CKINVDCx12_ASAP7_75t_R g85 ( 
.A(n_58),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_46),
.B(n_61),
.Y(n_86)
);

CKINVDCx16_ASAP7_75t_R g109 ( 
.A(n_86),
.Y(n_109)
);

OA22x2_ASAP7_75t_L g87 ( 
.A1(n_56),
.A2(n_34),
.B1(n_41),
.B2(n_42),
.Y(n_87)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_54),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_88),
.Y(n_93)
);

AND2x2_ASAP7_75t_L g89 ( 
.A(n_49),
.B(n_0),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_52),
.B(n_20),
.Y(n_90)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_90),
.Y(n_92)
);

CKINVDCx6p67_ASAP7_75t_R g91 ( 
.A(n_49),
.Y(n_91)
);

INVx4_ASAP7_75t_L g111 ( 
.A(n_91),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_64),
.A2(n_44),
.B1(n_54),
.B2(n_45),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_95),
.A2(n_114),
.B1(n_89),
.B2(n_58),
.Y(n_142)
);

BUFx3_ASAP7_75t_L g96 ( 
.A(n_91),
.Y(n_96)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_96),
.Y(n_123)
);

OR2x2_ASAP7_75t_L g97 ( 
.A(n_76),
.B(n_52),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_97),
.B(n_101),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_64),
.B(n_52),
.Y(n_101)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_87),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_104),
.B(n_106),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_105),
.A2(n_29),
.B1(n_24),
.B2(n_30),
.Y(n_145)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_87),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_L g128 ( 
.A1(n_108),
.A2(n_67),
.B1(n_81),
.B2(n_71),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_69),
.B(n_55),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_112),
.B(n_115),
.Y(n_126)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_87),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_113),
.B(n_117),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_71),
.A2(n_74),
.B1(n_78),
.B2(n_70),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_80),
.B(n_55),
.Y(n_115)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_62),
.Y(n_117)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_63),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_119),
.B(n_72),
.Y(n_127)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_110),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_120),
.B(n_122),
.Y(n_181)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_110),
.Y(n_122)
);

NAND2xp33_ASAP7_75t_SL g124 ( 
.A(n_114),
.B(n_71),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_SL g155 ( 
.A1(n_124),
.A2(n_131),
.B(n_138),
.Y(n_155)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_96),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_125),
.Y(n_179)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_127),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_L g178 ( 
.A1(n_128),
.A2(n_21),
.B1(n_19),
.B2(n_31),
.Y(n_178)
);

INVx13_ASAP7_75t_L g129 ( 
.A(n_111),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_SL g177 ( 
.A1(n_129),
.A2(n_137),
.B1(n_140),
.B2(n_94),
.Y(n_177)
);

AND2x6_ASAP7_75t_L g131 ( 
.A(n_98),
.B(n_91),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_101),
.B(n_76),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_132),
.B(n_133),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_SL g133 ( 
.A(n_97),
.B(n_107),
.Y(n_133)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_95),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_134),
.B(n_135),
.Y(n_159)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_112),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_102),
.A2(n_65),
.B1(n_75),
.B2(n_66),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_136),
.A2(n_141),
.B1(n_144),
.B2(n_145),
.Y(n_151)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_100),
.Y(n_137)
);

O2A1O1Ixp33_ASAP7_75t_L g138 ( 
.A1(n_102),
.A2(n_79),
.B(n_91),
.C(n_54),
.Y(n_138)
);

AND2x2_ASAP7_75t_SL g139 ( 
.A(n_99),
.B(n_82),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_L g158 ( 
.A1(n_139),
.A2(n_109),
.B(n_97),
.Y(n_158)
);

AOI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_104),
.A2(n_88),
.B1(n_82),
.B2(n_89),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_106),
.A2(n_42),
.B1(n_41),
.B2(n_68),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_L g150 ( 
.A(n_142),
.B(n_99),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_116),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_SL g173 ( 
.A1(n_143),
.A2(n_148),
.B(n_83),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_113),
.A2(n_73),
.B1(n_68),
.B2(n_30),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_98),
.A2(n_73),
.B1(n_29),
.B2(n_24),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_147),
.A2(n_30),
.B1(n_103),
.B2(n_100),
.Y(n_166)
);

AND2x6_ASAP7_75t_L g148 ( 
.A(n_98),
.B(n_85),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_107),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_149),
.B(n_118),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_L g198 ( 
.A(n_150),
.B(n_163),
.Y(n_198)
);

AOI21xp5_ASAP7_75t_L g152 ( 
.A1(n_120),
.A2(n_115),
.B(n_92),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_L g200 ( 
.A1(n_152),
.A2(n_158),
.B(n_160),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_139),
.B(n_92),
.C(n_117),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_156),
.B(n_168),
.C(n_169),
.Y(n_204)
);

INVx1_ASAP7_75t_SL g157 ( 
.A(n_126),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_157),
.B(n_173),
.Y(n_185)
);

AOI21xp5_ASAP7_75t_L g160 ( 
.A1(n_122),
.A2(n_109),
.B(n_111),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_138),
.A2(n_93),
.B1(n_118),
.B2(n_103),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_L g206 ( 
.A1(n_161),
.A2(n_164),
.B(n_182),
.Y(n_206)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_144),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_162),
.B(n_167),
.Y(n_208)
);

XOR2xp5_ASAP7_75t_SL g163 ( 
.A(n_139),
.B(n_15),
.Y(n_163)
);

AOI21xp5_ASAP7_75t_L g164 ( 
.A1(n_146),
.A2(n_93),
.B(n_57),
.Y(n_164)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_165),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_166),
.A2(n_170),
.B1(n_174),
.B2(n_129),
.Y(n_193)
);

INVxp67_ASAP7_75t_L g167 ( 
.A(n_141),
.Y(n_167)
);

XOR2xp5_ASAP7_75t_L g168 ( 
.A(n_142),
.B(n_57),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_139),
.B(n_57),
.C(n_83),
.Y(n_169)
);

OA21x2_ASAP7_75t_L g170 ( 
.A1(n_134),
.A2(n_31),
.B(n_21),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_146),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_171),
.B(n_175),
.Y(n_186)
);

INVxp67_ASAP7_75t_L g172 ( 
.A(n_138),
.Y(n_172)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_172),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_136),
.A2(n_94),
.B1(n_119),
.B2(n_31),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_130),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_130),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_176),
.B(n_180),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_177),
.A2(n_178),
.B1(n_129),
.B2(n_123),
.Y(n_191)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_126),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_L g182 ( 
.A1(n_121),
.A2(n_27),
.B(n_21),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_121),
.B(n_27),
.Y(n_183)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_183),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_165),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_184),
.B(n_187),
.Y(n_226)
);

INVxp67_ASAP7_75t_L g187 ( 
.A(n_161),
.Y(n_187)
);

BUFx3_ASAP7_75t_L g188 ( 
.A(n_153),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_188),
.Y(n_238)
);

INVxp67_ASAP7_75t_L g190 ( 
.A(n_164),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_190),
.B(n_213),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_L g235 ( 
.A1(n_191),
.A2(n_193),
.B1(n_208),
.B2(n_206),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_151),
.A2(n_124),
.B1(n_131),
.B2(n_135),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_194),
.A2(n_209),
.B1(n_162),
.B2(n_176),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_179),
.B(n_125),
.Y(n_195)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_195),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_179),
.B(n_123),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_SL g221 ( 
.A(n_196),
.B(n_197),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_153),
.B(n_137),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_154),
.B(n_132),
.Y(n_199)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_199),
.Y(n_217)
);

AND2x2_ASAP7_75t_L g202 ( 
.A(n_171),
.B(n_149),
.Y(n_202)
);

AOI21xp5_ASAP7_75t_SL g231 ( 
.A1(n_202),
.A2(n_160),
.B(n_158),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g203 ( 
.A(n_150),
.B(n_148),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_203),
.B(n_207),
.C(n_169),
.Y(n_230)
);

AND2x6_ASAP7_75t_L g205 ( 
.A(n_173),
.B(n_133),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_205),
.B(n_155),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_180),
.B(n_147),
.C(n_143),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_151),
.A2(n_145),
.B1(n_27),
.B2(n_19),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_159),
.A2(n_83),
.B1(n_72),
.B2(n_2),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_210),
.A2(n_175),
.B1(n_166),
.B2(n_163),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_181),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_SL g228 ( 
.A(n_211),
.B(n_154),
.Y(n_228)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_181),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_214),
.A2(n_219),
.B1(n_237),
.B2(n_213),
.Y(n_239)
);

CKINVDCx14_ASAP7_75t_R g248 ( 
.A(n_216),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_218),
.B(n_204),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_194),
.A2(n_155),
.B1(n_159),
.B2(n_157),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_199),
.B(n_157),
.Y(n_220)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_220),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_203),
.B(n_168),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_222),
.B(n_230),
.C(n_236),
.Y(n_241)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_186),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_223),
.B(n_227),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_210),
.B(n_152),
.Y(n_224)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_224),
.Y(n_254)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_186),
.Y(n_227)
);

OR2x2_ASAP7_75t_L g240 ( 
.A(n_228),
.B(n_202),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_187),
.A2(n_174),
.B1(n_170),
.B2(n_182),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_L g242 ( 
.A1(n_229),
.A2(n_234),
.B1(n_209),
.B2(n_206),
.Y(n_242)
);

AOI21x1_ASAP7_75t_L g256 ( 
.A1(n_231),
.A2(n_232),
.B(n_234),
.Y(n_256)
);

AND2x2_ASAP7_75t_L g232 ( 
.A(n_192),
.B(n_156),
.Y(n_232)
);

INVxp67_ASAP7_75t_L g233 ( 
.A(n_185),
.Y(n_233)
);

INVxp67_ASAP7_75t_L g246 ( 
.A(n_233),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_190),
.A2(n_170),
.B1(n_183),
.B2(n_72),
.Y(n_234)
);

CKINVDCx16_ASAP7_75t_R g252 ( 
.A(n_235),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_204),
.B(n_170),
.C(n_72),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_205),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_239),
.A2(n_249),
.B1(n_251),
.B2(n_253),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_SL g259 ( 
.A(n_240),
.B(n_257),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_242),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_L g243 ( 
.A1(n_233),
.A2(n_226),
.B1(n_215),
.B2(n_223),
.Y(n_243)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_243),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_230),
.B(n_198),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_245),
.B(n_258),
.C(n_236),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_L g247 ( 
.A1(n_229),
.A2(n_193),
.B1(n_200),
.B2(n_207),
.Y(n_247)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_247),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_219),
.A2(n_201),
.B1(n_212),
.B2(n_200),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_L g253 ( 
.A1(n_215),
.A2(n_201),
.B1(n_189),
.B2(n_212),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_237),
.A2(n_189),
.B1(n_202),
.B2(n_188),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_L g270 ( 
.A1(n_255),
.A2(n_15),
.B1(n_14),
.B2(n_13),
.Y(n_270)
);

AOI22xp33_ASAP7_75t_SL g266 ( 
.A1(n_256),
.A2(n_238),
.B1(n_232),
.B2(n_220),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_221),
.B(n_198),
.Y(n_257)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_222),
.B(n_15),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_262),
.B(n_268),
.C(n_269),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_252),
.A2(n_227),
.B1(n_214),
.B2(n_217),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_263),
.A2(n_265),
.B1(n_266),
.B2(n_248),
.Y(n_281)
);

OR2x2_ASAP7_75t_L g264 ( 
.A(n_255),
.B(n_216),
.Y(n_264)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_264),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_256),
.A2(n_217),
.B1(n_225),
.B2(n_231),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_241),
.B(n_232),
.C(n_4),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_241),
.B(n_3),
.C(n_4),
.Y(n_269)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_270),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_245),
.B(n_3),
.C(n_4),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_SL g277 ( 
.A(n_271),
.B(n_272),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_244),
.B(n_3),
.C(n_4),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_251),
.B(n_14),
.Y(n_273)
);

XOR2xp5_ASAP7_75t_L g278 ( 
.A(n_273),
.B(n_258),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g290 ( 
.A(n_278),
.B(n_273),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_SL g279 ( 
.A(n_261),
.B(n_246),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_279),
.B(n_280),
.Y(n_295)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_272),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_SL g296 ( 
.A(n_281),
.B(n_283),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_267),
.A2(n_239),
.B1(n_244),
.B2(n_250),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g299 ( 
.A1(n_282),
.A2(n_285),
.B1(n_8),
.B2(n_9),
.Y(n_299)
);

AO22x1_ASAP7_75t_L g283 ( 
.A1(n_265),
.A2(n_250),
.B1(n_253),
.B2(n_243),
.Y(n_283)
);

XOR2xp5_ASAP7_75t_L g284 ( 
.A(n_262),
.B(n_246),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_284),
.B(n_286),
.C(n_271),
.Y(n_291)
);

CKINVDCx14_ASAP7_75t_R g285 ( 
.A(n_259),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g286 ( 
.A(n_263),
.B(n_254),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_274),
.A2(n_254),
.B1(n_240),
.B2(n_13),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_288),
.A2(n_260),
.B1(n_264),
.B2(n_268),
.Y(n_289)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_289),
.Y(n_303)
);

XOR2xp5_ASAP7_75t_L g301 ( 
.A(n_290),
.B(n_291),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_286),
.B(n_269),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_292),
.B(n_299),
.Y(n_308)
);

XNOR2xp5_ASAP7_75t_L g293 ( 
.A(n_287),
.B(n_13),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_SL g304 ( 
.A(n_293),
.B(n_294),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_SL g294 ( 
.A1(n_288),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_284),
.B(n_5),
.C(n_6),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_297),
.B(n_298),
.C(n_300),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_287),
.B(n_5),
.C(n_7),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_281),
.B(n_8),
.C(n_9),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_300),
.B(n_282),
.Y(n_305)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_305),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_295),
.B(n_276),
.Y(n_306)
);

OAI21xp5_ASAP7_75t_SL g312 ( 
.A1(n_306),
.A2(n_307),
.B(n_298),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_291),
.B(n_275),
.C(n_278),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_L g310 ( 
.A1(n_303),
.A2(n_296),
.B1(n_283),
.B2(n_297),
.Y(n_310)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_310),
.Y(n_314)
);

OAI22xp5_ASAP7_75t_SL g311 ( 
.A1(n_308),
.A2(n_283),
.B1(n_296),
.B2(n_277),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_SL g315 ( 
.A(n_311),
.B(n_312),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_SL g313 ( 
.A1(n_302),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_315),
.B(n_309),
.Y(n_316)
);

OAI21xp5_ASAP7_75t_L g317 ( 
.A1(n_316),
.A2(n_302),
.B(n_314),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_317),
.B(n_311),
.C(n_301),
.Y(n_318)
);

AOI322xp5_ASAP7_75t_L g319 ( 
.A1(n_318),
.A2(n_301),
.A3(n_310),
.B1(n_304),
.B2(n_313),
.C1(n_12),
.C2(n_11),
.Y(n_319)
);

AOI21xp5_ASAP7_75t_L g320 ( 
.A1(n_319),
.A2(n_8),
.B(n_9),
.Y(n_320)
);

OAI21xp5_ASAP7_75t_L g321 ( 
.A1(n_320),
.A2(n_11),
.B(n_12),
.Y(n_321)
);

AOI21xp5_ASAP7_75t_L g322 ( 
.A1(n_321),
.A2(n_11),
.B(n_294),
.Y(n_322)
);


endmodule