module fake_ariane_1008_n_1528 (n_83, n_8, n_233, n_56, n_60, n_170, n_190, n_160, n_64, n_179, n_180, n_119, n_124, n_240, n_167, n_90, n_195, n_38, n_213, n_47, n_110, n_153, n_18, n_197, n_221, n_86, n_75, n_89, n_67, n_176, n_149, n_34, n_158, n_237, n_172, n_69, n_259, n_95, n_175, n_92, n_143, n_183, n_203, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_181, n_152, n_120, n_169, n_106, n_12, n_53, n_173, n_111, n_21, n_242, n_260, n_115, n_133, n_66, n_205, n_236, n_71, n_24, n_7, n_109, n_208, n_245, n_96, n_156, n_209, n_49, n_20, n_174, n_100, n_17, n_50, n_187, n_132, n_62, n_210, n_147, n_204, n_225, n_235, n_200, n_51, n_166, n_253, n_76, n_218, n_103, n_79, n_26, n_244, n_226, n_3, n_246, n_46, n_220, n_0, n_84, n_247, n_36, n_199, n_91, n_159, n_107, n_189, n_72, n_105, n_128, n_217, n_44, n_224, n_30, n_82, n_178, n_31, n_42, n_57, n_131, n_201, n_229, n_70, n_250, n_222, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_256, n_6, n_214, n_227, n_48, n_94, n_101, n_243, n_4, n_134, n_188, n_185, n_2, n_32, n_249, n_37, n_58, n_65, n_123, n_212, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_255, n_122, n_257, n_198, n_148, n_232, n_164, n_52, n_157, n_248, n_184, n_177, n_135, n_258, n_73, n_77, n_171, n_228, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_182, n_196, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_206, n_13, n_27, n_207, n_241, n_29, n_254, n_238, n_41, n_219, n_140, n_55, n_191, n_151, n_136, n_231, n_192, n_28, n_80, n_146, n_234, n_230, n_211, n_194, n_97, n_154, n_215, n_252, n_142, n_251, n_161, n_14, n_163, n_88, n_186, n_141, n_68, n_116, n_104, n_202, n_145, n_78, n_193, n_39, n_59, n_63, n_99, n_216, n_16, n_5, n_155, n_127, n_239, n_223, n_35, n_54, n_25, n_1528);

input n_83;
input n_8;
input n_233;
input n_56;
input n_60;
input n_170;
input n_190;
input n_160;
input n_64;
input n_179;
input n_180;
input n_119;
input n_124;
input n_240;
input n_167;
input n_90;
input n_195;
input n_38;
input n_213;
input n_47;
input n_110;
input n_153;
input n_18;
input n_197;
input n_221;
input n_86;
input n_75;
input n_89;
input n_67;
input n_176;
input n_149;
input n_34;
input n_158;
input n_237;
input n_172;
input n_69;
input n_259;
input n_95;
input n_175;
input n_92;
input n_143;
input n_183;
input n_203;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_181;
input n_152;
input n_120;
input n_169;
input n_106;
input n_12;
input n_53;
input n_173;
input n_111;
input n_21;
input n_242;
input n_260;
input n_115;
input n_133;
input n_66;
input n_205;
input n_236;
input n_71;
input n_24;
input n_7;
input n_109;
input n_208;
input n_245;
input n_96;
input n_156;
input n_209;
input n_49;
input n_20;
input n_174;
input n_100;
input n_17;
input n_50;
input n_187;
input n_132;
input n_62;
input n_210;
input n_147;
input n_204;
input n_225;
input n_235;
input n_200;
input n_51;
input n_166;
input n_253;
input n_76;
input n_218;
input n_103;
input n_79;
input n_26;
input n_244;
input n_226;
input n_3;
input n_246;
input n_46;
input n_220;
input n_0;
input n_84;
input n_247;
input n_36;
input n_199;
input n_91;
input n_159;
input n_107;
input n_189;
input n_72;
input n_105;
input n_128;
input n_217;
input n_44;
input n_224;
input n_30;
input n_82;
input n_178;
input n_31;
input n_42;
input n_57;
input n_131;
input n_201;
input n_229;
input n_70;
input n_250;
input n_222;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_256;
input n_6;
input n_214;
input n_227;
input n_48;
input n_94;
input n_101;
input n_243;
input n_4;
input n_134;
input n_188;
input n_185;
input n_2;
input n_32;
input n_249;
input n_37;
input n_58;
input n_65;
input n_123;
input n_212;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_255;
input n_122;
input n_257;
input n_198;
input n_148;
input n_232;
input n_164;
input n_52;
input n_157;
input n_248;
input n_184;
input n_177;
input n_135;
input n_258;
input n_73;
input n_77;
input n_171;
input n_228;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_182;
input n_196;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_206;
input n_13;
input n_27;
input n_207;
input n_241;
input n_29;
input n_254;
input n_238;
input n_41;
input n_219;
input n_140;
input n_55;
input n_191;
input n_151;
input n_136;
input n_231;
input n_192;
input n_28;
input n_80;
input n_146;
input n_234;
input n_230;
input n_211;
input n_194;
input n_97;
input n_154;
input n_215;
input n_252;
input n_142;
input n_251;
input n_161;
input n_14;
input n_163;
input n_88;
input n_186;
input n_141;
input n_68;
input n_116;
input n_104;
input n_202;
input n_145;
input n_78;
input n_193;
input n_39;
input n_59;
input n_63;
input n_99;
input n_216;
input n_16;
input n_5;
input n_155;
input n_127;
input n_239;
input n_223;
input n_35;
input n_54;
input n_25;

output n_1528;

wire n_913;
wire n_1486;
wire n_1507;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_1250;
wire n_1169;
wire n_789;
wire n_850;
wire n_610;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_1463;
wire n_1238;
wire n_1515;
wire n_817;
wire n_924;
wire n_781;
wire n_717;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_524;
wire n_1214;
wire n_634;
wire n_1246;
wire n_1138;
wire n_764;
wire n_1503;
wire n_462;
wire n_1196;
wire n_1181;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1366;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1457;
wire n_377;
wire n_520;
wire n_870;
wire n_1453;
wire n_279;
wire n_945;
wire n_958;
wire n_813;
wire n_419;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1184;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_1073;
wire n_402;
wire n_1277;
wire n_829;
wire n_1062;
wire n_339;
wire n_738;
wire n_672;
wire n_740;
wire n_1283;
wire n_1018;
wire n_953;
wire n_1364;
wire n_1224;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_989;
wire n_645;
wire n_331;
wire n_559;
wire n_267;
wire n_495;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1276;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1519;
wire n_1195;
wire n_1522;
wire n_518;
wire n_1207;
wire n_786;
wire n_1404;
wire n_868;
wire n_1314;
wire n_1512;
wire n_884;
wire n_1415;
wire n_1034;
wire n_1085;
wire n_277;
wire n_432;
wire n_293;
wire n_823;
wire n_620;
wire n_1074;
wire n_859;
wire n_587;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_352;
wire n_899;
wire n_611;
wire n_1295;
wire n_365;
wire n_1013;
wire n_1495;
wire n_334;
wire n_661;
wire n_300;
wire n_533;
wire n_438;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_376;
wire n_512;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1354;
wire n_1213;
wire n_780;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_942;
wire n_1437;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_490;
wire n_1461;
wire n_1391;
wire n_1006;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_676;
wire n_680;
wire n_287;
wire n_302;
wire n_380;
wire n_1432;
wire n_1108;
wire n_851;
wire n_355;
wire n_444;
wire n_1351;
wire n_1274;
wire n_652;
wire n_475;
wire n_947;
wire n_1260;
wire n_930;
wire n_1179;
wire n_468;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_407;
wire n_916;
wire n_1386;
wire n_912;
wire n_460;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_555;
wire n_804;
wire n_1382;
wire n_992;
wire n_966;
wire n_955;
wire n_1182;
wire n_794;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_288;
wire n_1292;
wire n_1178;
wire n_1435;
wire n_1026;
wire n_1506;
wire n_306;
wire n_436;
wire n_324;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_1083;
wire n_967;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_824;
wire n_428;
wire n_892;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1343;
wire n_563;
wire n_990;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_964;
wire n_382;
wire n_489;
wire n_974;
wire n_506;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_934;
wire n_1447;
wire n_1220;
wire n_356;
wire n_698;
wire n_307;
wire n_1209;
wire n_1020;
wire n_646;
wire n_404;
wire n_1058;
wire n_347;
wire n_1042;
wire n_1234;
wire n_479;
wire n_1455;
wire n_299;
wire n_836;
wire n_1279;
wire n_564;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_713;
wire n_1255;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_370;
wire n_706;
wire n_286;
wire n_1401;
wire n_1419;
wire n_776;
wire n_424;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_552;
wire n_348;
wire n_670;
wire n_379;
wire n_264;
wire n_441;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_905;
wire n_720;
wire n_926;
wire n_1163;
wire n_1384;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1413;
wire n_855;
wire n_808;
wire n_1365;
wire n_553;
wire n_1439;
wire n_814;
wire n_578;
wire n_1287;
wire n_405;
wire n_320;
wire n_1414;
wire n_1134;
wire n_1484;
wire n_647;
wire n_1423;
wire n_481;
wire n_600;
wire n_1053;
wire n_529;
wire n_502;
wire n_1467;
wire n_1304;
wire n_1105;
wire n_547;
wire n_439;
wire n_604;
wire n_677;
wire n_478;
wire n_703;
wire n_1349;
wire n_1061;
wire n_326;
wire n_681;
wire n_874;
wire n_1278;
wire n_707;
wire n_983;
wire n_590;
wire n_727;
wire n_699;
wire n_301;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_325;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1080;
wire n_920;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_729;
wire n_887;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_1402;
wire n_388;
wire n_957;
wire n_1242;
wire n_1489;
wire n_1218;
wire n_321;
wire n_861;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_281;
wire n_262;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_888;
wire n_845;
wire n_1297;
wire n_551;
wire n_417;
wire n_343;
wire n_1222;
wire n_582;
wire n_755;
wire n_1097;
wire n_1219;
wire n_710;
wire n_534;
wire n_1460;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_451;
wire n_745;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1388;
wire n_1266;
wire n_769;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_982;
wire n_915;
wire n_1075;
wire n_454;
wire n_298;
wire n_1331;
wire n_1227;
wire n_655;
wire n_403;
wire n_1007;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_659;
wire n_1332;
wire n_509;
wire n_666;
wire n_430;
wire n_1206;
wire n_722;
wire n_1508;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1338;
wire n_1342;
wire n_456;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_521;
wire n_873;
wire n_1301;
wire n_1243;
wire n_1400;
wire n_342;
wire n_1466;
wire n_1513;
wire n_1527;
wire n_358;
wire n_608;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1257;
wire n_1480;
wire n_1078;
wire n_266;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_1449;
wire n_687;
wire n_797;
wire n_480;
wire n_1327;
wire n_1475;
wire n_642;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_393;
wire n_474;
wire n_805;
wire n_295;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_730;
wire n_386;
wire n_1281;
wire n_516;
wire n_1137;
wire n_1258;
wire n_640;
wire n_463;
wire n_1476;
wire n_1524;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_726;
wire n_1123;
wire n_878;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_283;
wire n_806;
wire n_1350;
wire n_649;
wire n_374;
wire n_1352;
wire n_643;
wire n_1492;
wire n_1441;
wire n_682;
wire n_819;
wire n_586;
wire n_1324;
wire n_1429;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1208;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1448;
wire n_1009;
wire n_1133;
wire n_883;
wire n_473;
wire n_801;
wire n_1286;
wire n_818;
wire n_779;
wire n_594;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1438;
wire n_597;
wire n_1047;
wire n_1472;
wire n_1050;
wire n_566;
wire n_1201;
wire n_1288;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_426;
wire n_433;
wire n_398;
wire n_1090;
wire n_1367;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1192;
wire n_894;
wire n_1380;
wire n_420;
wire n_1291;
wire n_562;
wire n_748;
wire n_510;
wire n_1045;
wire n_1160;
wire n_1023;
wire n_988;
wire n_330;
wire n_914;
wire n_689;
wire n_400;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_467;
wire n_1511;
wire n_1422;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_538;
wire n_1517;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_1307;
wire n_1128;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1440;
wire n_1370;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1403;
wire n_1065;
wire n_453;
wire n_810;
wire n_1290;
wire n_617;
wire n_543;
wire n_1362;
wire n_601;
wire n_683;
wire n_565;
wire n_628;
wire n_1300;
wire n_743;
wire n_1194;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1135;
wire n_918;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_571;
wire n_414;
wire n_1521;
wire n_284;
wire n_593;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_409;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_526;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1444;
wire n_820;
wire n_872;
wire n_1157;
wire n_848;
wire n_280;
wire n_629;
wire n_532;
wire n_763;
wire n_540;
wire n_692;
wire n_984;
wire n_750;
wire n_834;
wire n_800;
wire n_395;
wire n_621;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_493;
wire n_1311;
wire n_1100;
wire n_585;
wire n_875;
wire n_827;
wire n_697;
wire n_622;
wire n_1335;
wire n_296;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_792;
wire n_1262;
wire n_580;
wire n_494;
wire n_434;
wire n_975;
wire n_394;
wire n_923;
wire n_1381;
wire n_1124;
wire n_1494;
wire n_932;
wire n_1183;
wire n_1326;
wire n_981;
wire n_1110;
wire n_1407;
wire n_1204;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1054;
wire n_508;
wire n_353;
wire n_1482;
wire n_1361;
wire n_1057;
wire n_978;
wire n_1011;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_653;
wire n_1445;
wire n_1317;
wire n_783;
wire n_556;
wire n_1127;
wire n_1471;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_987;
wire n_936;
wire n_1385;
wire n_1525;
wire n_541;
wire n_499;
wire n_788;
wire n_908;
wire n_1036;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_318;
wire n_1458;
wire n_679;
wire n_663;
wire n_443;
wire n_1412;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_391;
wire n_940;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_765;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_898;
wire n_857;
wire n_363;
wire n_968;
wire n_1067;
wire n_1323;
wire n_1235;
wire n_1462;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1093;
wire n_1285;
wire n_733;
wire n_761;
wire n_731;
wire n_336;
wire n_315;
wire n_311;
wire n_1452;
wire n_668;
wire n_758;
wire n_1106;
wire n_648;
wire n_784;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_1348;
wire n_753;
wire n_701;
wire n_1003;
wire n_1125;
wire n_309;
wire n_1344;
wire n_1390;
wire n_401;
wire n_485;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_291;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1510;
wire n_1099;
wire n_839;
wire n_759;
wire n_567;
wire n_369;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_323;
wire n_550;
wire n_1315;
wire n_997;
wire n_635;
wire n_694;
wire n_1320;
wire n_1113;
wire n_1152;
wire n_921;
wire n_1236;
wire n_1265;
wire n_1470;
wire n_671;
wire n_1409;
wire n_1148;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_498;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1289;
wire n_1497;
wire n_459;
wire n_1136;
wire n_458;
wire n_1190;
wire n_1144;
wire n_838;
wire n_383;
wire n_1316;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_709;
wire n_809;
wire n_881;
wire n_1019;
wire n_1477;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_1114;
wire n_1325;
wire n_708;
wire n_308;
wire n_1223;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1041;
wire n_993;
wire n_948;
wire n_922;
wire n_1004;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_450;
wire n_896;
wire n_1479;
wire n_902;
wire n_1031;
wire n_853;
wire n_716;
wire n_1337;
wire n_774;
wire n_933;
wire n_596;
wire n_954;
wire n_1168;
wire n_1310;
wire n_656;
wire n_492;
wire n_574;
wire n_664;
wire n_1229;
wire n_415;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1126;
wire n_938;
wire n_1328;
wire n_895;
wire n_304;
wire n_583;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_946;
wire n_757;
wire n_375;
wire n_1146;
wire n_1203;
wire n_998;
wire n_472;
wire n_937;
wire n_1474;
wire n_265;
wire n_275;
wire n_1375;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_496;
wire n_866;
wire n_925;
wire n_1313;
wire n_1001;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_1129;
wire n_1252;
wire n_1464;
wire n_1296;
wire n_773;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_329;
wire n_718;
wire n_1434;
wire n_340;
wire n_548;
wire n_289;
wire n_523;
wire n_457;
wire n_1299;
wire n_782;
wire n_364;
wire n_431;
wire n_1228;
wire n_1244;
wire n_484;
wire n_411;
wire n_849;
wire n_357;
wire n_412;
wire n_1251;
wire n_447;
wire n_1421;
wire n_1233;
wire n_893;
wire n_841;
wire n_886;
wire n_1069;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1374;
wire n_1451;
wire n_1487;
wire n_675;

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_155),
.Y(n_261)
);

INVx1_ASAP7_75t_SL g262 ( 
.A(n_175),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_55),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_19),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_104),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_214),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_95),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_123),
.Y(n_268)
);

INVx2_ASAP7_75t_SL g269 ( 
.A(n_254),
.Y(n_269)
);

BUFx8_ASAP7_75t_SL g270 ( 
.A(n_226),
.Y(n_270)
);

BUFx10_ASAP7_75t_L g271 ( 
.A(n_18),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_103),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_185),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_193),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_191),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_183),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_62),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_172),
.Y(n_278)
);

INVx1_ASAP7_75t_SL g279 ( 
.A(n_219),
.Y(n_279)
);

BUFx10_ASAP7_75t_L g280 ( 
.A(n_235),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_30),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_150),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_125),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_173),
.Y(n_284)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_105),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_174),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_142),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_108),
.Y(n_288)
);

INVx2_ASAP7_75t_SL g289 ( 
.A(n_143),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_229),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_257),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_2),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_9),
.Y(n_293)
);

BUFx6f_ASAP7_75t_L g294 ( 
.A(n_78),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_152),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_118),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_147),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_206),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_131),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_158),
.Y(n_300)
);

INVx2_ASAP7_75t_L g301 ( 
.A(n_19),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_115),
.Y(n_302)
);

INVx2_ASAP7_75t_SL g303 ( 
.A(n_163),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_188),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_107),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_208),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_195),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_92),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_196),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_168),
.Y(n_310)
);

INVx2_ASAP7_75t_L g311 ( 
.A(n_217),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_129),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_66),
.Y(n_313)
);

BUFx6f_ASAP7_75t_L g314 ( 
.A(n_170),
.Y(n_314)
);

HB1xp67_ASAP7_75t_L g315 ( 
.A(n_48),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_146),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_116),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_237),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g319 ( 
.A(n_194),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_200),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_132),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_41),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_149),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_18),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_209),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_81),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_241),
.Y(n_327)
);

INVx1_ASAP7_75t_SL g328 ( 
.A(n_100),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_47),
.Y(n_329)
);

CKINVDCx20_ASAP7_75t_R g330 ( 
.A(n_178),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_186),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_34),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_94),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_210),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_9),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_245),
.Y(n_336)
);

INVx3_ASAP7_75t_L g337 ( 
.A(n_130),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_49),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_205),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_164),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_128),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_251),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_23),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_169),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_114),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_11),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_44),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_134),
.Y(n_348)
);

BUFx5_ASAP7_75t_L g349 ( 
.A(n_25),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_41),
.Y(n_350)
);

INVx1_ASAP7_75t_SL g351 ( 
.A(n_180),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_203),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_223),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_162),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_247),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_153),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_61),
.Y(n_357)
);

BUFx10_ASAP7_75t_L g358 ( 
.A(n_80),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_145),
.Y(n_359)
);

BUFx6f_ASAP7_75t_L g360 ( 
.A(n_2),
.Y(n_360)
);

CKINVDCx14_ASAP7_75t_R g361 ( 
.A(n_59),
.Y(n_361)
);

BUFx2_ASAP7_75t_L g362 ( 
.A(n_62),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_1),
.Y(n_363)
);

HB1xp67_ASAP7_75t_L g364 ( 
.A(n_252),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_231),
.Y(n_365)
);

BUFx3_ASAP7_75t_L g366 ( 
.A(n_83),
.Y(n_366)
);

INVx2_ASAP7_75t_L g367 ( 
.A(n_165),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_236),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_133),
.Y(n_369)
);

BUFx3_ASAP7_75t_L g370 ( 
.A(n_136),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_69),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_22),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_73),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_76),
.Y(n_374)
);

INVx2_ASAP7_75t_L g375 ( 
.A(n_48),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_225),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_47),
.Y(n_377)
);

CKINVDCx16_ASAP7_75t_R g378 ( 
.A(n_181),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_151),
.Y(n_379)
);

CKINVDCx20_ASAP7_75t_R g380 ( 
.A(n_232),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_177),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_144),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_243),
.Y(n_383)
);

BUFx10_ASAP7_75t_L g384 ( 
.A(n_26),
.Y(n_384)
);

BUFx3_ASAP7_75t_L g385 ( 
.A(n_65),
.Y(n_385)
);

INVx2_ASAP7_75t_L g386 ( 
.A(n_65),
.Y(n_386)
);

INVx2_ASAP7_75t_L g387 ( 
.A(n_75),
.Y(n_387)
);

BUFx2_ASAP7_75t_L g388 ( 
.A(n_17),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_215),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_39),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_119),
.Y(n_391)
);

BUFx10_ASAP7_75t_L g392 ( 
.A(n_82),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_199),
.Y(n_393)
);

INVx2_ASAP7_75t_SL g394 ( 
.A(n_244),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_67),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_189),
.Y(n_396)
);

CKINVDCx16_ASAP7_75t_R g397 ( 
.A(n_171),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_141),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_15),
.Y(n_399)
);

BUFx3_ASAP7_75t_L g400 ( 
.A(n_230),
.Y(n_400)
);

CKINVDCx20_ASAP7_75t_R g401 ( 
.A(n_74),
.Y(n_401)
);

INVx2_ASAP7_75t_L g402 ( 
.A(n_160),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_76),
.Y(n_403)
);

CKINVDCx20_ASAP7_75t_R g404 ( 
.A(n_258),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_250),
.Y(n_405)
);

BUFx3_ASAP7_75t_L g406 ( 
.A(n_220),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_52),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_21),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_138),
.Y(n_409)
);

BUFx6f_ASAP7_75t_L g410 ( 
.A(n_97),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_56),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_166),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_57),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_85),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_33),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_113),
.Y(n_416)
);

INVx2_ASAP7_75t_SL g417 ( 
.A(n_86),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_101),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_135),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_218),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_51),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_11),
.Y(n_422)
);

INVx2_ASAP7_75t_L g423 ( 
.A(n_112),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_239),
.Y(n_424)
);

BUFx3_ASAP7_75t_L g425 ( 
.A(n_190),
.Y(n_425)
);

BUFx8_ASAP7_75t_SL g426 ( 
.A(n_227),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_7),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_12),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_216),
.Y(n_429)
);

CKINVDCx20_ASAP7_75t_R g430 ( 
.A(n_17),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_50),
.Y(n_431)
);

CKINVDCx5p33_ASAP7_75t_R g432 ( 
.A(n_16),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_102),
.Y(n_433)
);

NOR2xp33_ASAP7_75t_L g434 ( 
.A(n_364),
.B(n_0),
.Y(n_434)
);

CKINVDCx20_ASAP7_75t_R g435 ( 
.A(n_361),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_385),
.Y(n_436)
);

INVxp67_ASAP7_75t_SL g437 ( 
.A(n_385),
.Y(n_437)
);

BUFx2_ASAP7_75t_L g438 ( 
.A(n_362),
.Y(n_438)
);

CKINVDCx16_ASAP7_75t_R g439 ( 
.A(n_378),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_349),
.Y(n_440)
);

INVxp67_ASAP7_75t_L g441 ( 
.A(n_388),
.Y(n_441)
);

CKINVDCx20_ASAP7_75t_R g442 ( 
.A(n_291),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_349),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_397),
.Y(n_444)
);

CKINVDCx5p33_ASAP7_75t_R g445 ( 
.A(n_291),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_349),
.Y(n_446)
);

CKINVDCx20_ASAP7_75t_R g447 ( 
.A(n_319),
.Y(n_447)
);

CKINVDCx20_ASAP7_75t_R g448 ( 
.A(n_319),
.Y(n_448)
);

INVxp33_ASAP7_75t_SL g449 ( 
.A(n_315),
.Y(n_449)
);

INVxp67_ASAP7_75t_L g450 ( 
.A(n_271),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_349),
.Y(n_451)
);

CKINVDCx20_ASAP7_75t_R g452 ( 
.A(n_330),
.Y(n_452)
);

CKINVDCx20_ASAP7_75t_R g453 ( 
.A(n_330),
.Y(n_453)
);

CKINVDCx20_ASAP7_75t_R g454 ( 
.A(n_380),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_349),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_349),
.Y(n_456)
);

CKINVDCx5p33_ASAP7_75t_R g457 ( 
.A(n_380),
.Y(n_457)
);

HB1xp67_ASAP7_75t_L g458 ( 
.A(n_277),
.Y(n_458)
);

CKINVDCx5p33_ASAP7_75t_R g459 ( 
.A(n_404),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_349),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_263),
.Y(n_461)
);

CKINVDCx20_ASAP7_75t_R g462 ( 
.A(n_404),
.Y(n_462)
);

INVxp67_ASAP7_75t_SL g463 ( 
.A(n_294),
.Y(n_463)
);

HB1xp67_ASAP7_75t_L g464 ( 
.A(n_277),
.Y(n_464)
);

CKINVDCx20_ASAP7_75t_R g465 ( 
.A(n_401),
.Y(n_465)
);

CKINVDCx20_ASAP7_75t_R g466 ( 
.A(n_401),
.Y(n_466)
);

CKINVDCx5p33_ASAP7_75t_R g467 ( 
.A(n_280),
.Y(n_467)
);

CKINVDCx5p33_ASAP7_75t_R g468 ( 
.A(n_280),
.Y(n_468)
);

CKINVDCx20_ASAP7_75t_R g469 ( 
.A(n_430),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_L g470 ( 
.A(n_266),
.B(n_0),
.Y(n_470)
);

CKINVDCx5p33_ASAP7_75t_R g471 ( 
.A(n_280),
.Y(n_471)
);

INVxp67_ASAP7_75t_L g472 ( 
.A(n_271),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_313),
.Y(n_473)
);

INVx2_ASAP7_75t_L g474 ( 
.A(n_294),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_267),
.B(n_1),
.Y(n_475)
);

BUFx6f_ASAP7_75t_SL g476 ( 
.A(n_358),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_329),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_332),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_335),
.Y(n_479)
);

CKINVDCx20_ASAP7_75t_R g480 ( 
.A(n_430),
.Y(n_480)
);

CKINVDCx5p33_ASAP7_75t_R g481 ( 
.A(n_358),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_372),
.Y(n_482)
);

CKINVDCx5p33_ASAP7_75t_R g483 ( 
.A(n_358),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_377),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_399),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_422),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_301),
.Y(n_487)
);

CKINVDCx5p33_ASAP7_75t_R g488 ( 
.A(n_392),
.Y(n_488)
);

BUFx3_ASAP7_75t_L g489 ( 
.A(n_366),
.Y(n_489)
);

CKINVDCx5p33_ASAP7_75t_R g490 ( 
.A(n_392),
.Y(n_490)
);

CKINVDCx5p33_ASAP7_75t_R g491 ( 
.A(n_392),
.Y(n_491)
);

INVx1_ASAP7_75t_SL g492 ( 
.A(n_271),
.Y(n_492)
);

CKINVDCx5p33_ASAP7_75t_R g493 ( 
.A(n_261),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_301),
.Y(n_494)
);

CKINVDCx5p33_ASAP7_75t_R g495 ( 
.A(n_261),
.Y(n_495)
);

CKINVDCx5p33_ASAP7_75t_R g496 ( 
.A(n_268),
.Y(n_496)
);

NOR2xp33_ASAP7_75t_L g497 ( 
.A(n_337),
.B(n_3),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_375),
.Y(n_498)
);

INVxp67_ASAP7_75t_SL g499 ( 
.A(n_294),
.Y(n_499)
);

CKINVDCx5p33_ASAP7_75t_R g500 ( 
.A(n_268),
.Y(n_500)
);

CKINVDCx5p33_ASAP7_75t_R g501 ( 
.A(n_272),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_375),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_386),
.Y(n_503)
);

INVxp67_ASAP7_75t_L g504 ( 
.A(n_384),
.Y(n_504)
);

NOR2xp67_ASAP7_75t_L g505 ( 
.A(n_386),
.B(n_3),
.Y(n_505)
);

CKINVDCx5p33_ASAP7_75t_R g506 ( 
.A(n_272),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_L g507 ( 
.A(n_273),
.B(n_4),
.Y(n_507)
);

CKINVDCx5p33_ASAP7_75t_R g508 ( 
.A(n_274),
.Y(n_508)
);

CKINVDCx20_ASAP7_75t_R g509 ( 
.A(n_270),
.Y(n_509)
);

CKINVDCx20_ASAP7_75t_R g510 ( 
.A(n_426),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_387),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_387),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_294),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_294),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_360),
.Y(n_515)
);

CKINVDCx20_ASAP7_75t_R g516 ( 
.A(n_370),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_360),
.Y(n_517)
);

CKINVDCx20_ASAP7_75t_R g518 ( 
.A(n_370),
.Y(n_518)
);

HB1xp67_ASAP7_75t_L g519 ( 
.A(n_281),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_360),
.Y(n_520)
);

CKINVDCx16_ASAP7_75t_R g521 ( 
.A(n_439),
.Y(n_521)
);

AND2x2_ASAP7_75t_L g522 ( 
.A(n_437),
.B(n_384),
.Y(n_522)
);

INVx2_ASAP7_75t_L g523 ( 
.A(n_474),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_513),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_514),
.Y(n_525)
);

BUFx3_ASAP7_75t_L g526 ( 
.A(n_489),
.Y(n_526)
);

CKINVDCx5p33_ASAP7_75t_R g527 ( 
.A(n_509),
.Y(n_527)
);

CKINVDCx6p67_ASAP7_75t_R g528 ( 
.A(n_510),
.Y(n_528)
);

CKINVDCx5p33_ASAP7_75t_R g529 ( 
.A(n_445),
.Y(n_529)
);

INVx2_ASAP7_75t_L g530 ( 
.A(n_474),
.Y(n_530)
);

INVx2_ASAP7_75t_L g531 ( 
.A(n_440),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_515),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_517),
.Y(n_533)
);

CKINVDCx5p33_ASAP7_75t_R g534 ( 
.A(n_445),
.Y(n_534)
);

INVx2_ASAP7_75t_L g535 ( 
.A(n_443),
.Y(n_535)
);

BUFx2_ASAP7_75t_L g536 ( 
.A(n_444),
.Y(n_536)
);

NOR2xp33_ASAP7_75t_R g537 ( 
.A(n_493),
.B(n_433),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_520),
.Y(n_538)
);

BUFx6f_ASAP7_75t_L g539 ( 
.A(n_446),
.Y(n_539)
);

BUFx8_ASAP7_75t_L g540 ( 
.A(n_476),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_451),
.Y(n_541)
);

CKINVDCx5p33_ASAP7_75t_R g542 ( 
.A(n_457),
.Y(n_542)
);

CKINVDCx5p33_ASAP7_75t_R g543 ( 
.A(n_459),
.Y(n_543)
);

AND2x2_ASAP7_75t_L g544 ( 
.A(n_436),
.B(n_384),
.Y(n_544)
);

INVx2_ASAP7_75t_L g545 ( 
.A(n_455),
.Y(n_545)
);

INVx3_ASAP7_75t_L g546 ( 
.A(n_456),
.Y(n_546)
);

OA21x2_ASAP7_75t_L g547 ( 
.A1(n_460),
.A2(n_278),
.B(n_276),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_L g548 ( 
.A(n_463),
.B(n_284),
.Y(n_548)
);

BUFx8_ASAP7_75t_L g549 ( 
.A(n_476),
.Y(n_549)
);

NOR2xp33_ASAP7_75t_L g550 ( 
.A(n_493),
.B(n_337),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_499),
.Y(n_551)
);

OAI21x1_ASAP7_75t_L g552 ( 
.A1(n_470),
.A2(n_337),
.B(n_288),
.Y(n_552)
);

INVx4_ASAP7_75t_L g553 ( 
.A(n_476),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_497),
.Y(n_554)
);

BUFx6f_ASAP7_75t_L g555 ( 
.A(n_475),
.Y(n_555)
);

CKINVDCx5p33_ASAP7_75t_R g556 ( 
.A(n_459),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_487),
.Y(n_557)
);

XNOR2xp5_ASAP7_75t_L g558 ( 
.A(n_442),
.B(n_447),
.Y(n_558)
);

INVx3_ASAP7_75t_L g559 ( 
.A(n_489),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_494),
.Y(n_560)
);

CKINVDCx20_ASAP7_75t_R g561 ( 
.A(n_448),
.Y(n_561)
);

CKINVDCx5p33_ASAP7_75t_R g562 ( 
.A(n_452),
.Y(n_562)
);

NAND2xp33_ASAP7_75t_R g563 ( 
.A(n_444),
.B(n_281),
.Y(n_563)
);

INVx2_ASAP7_75t_L g564 ( 
.A(n_498),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_502),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_503),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_L g567 ( 
.A(n_461),
.B(n_287),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_511),
.Y(n_568)
);

NOR2xp33_ASAP7_75t_R g569 ( 
.A(n_495),
.B(n_496),
.Y(n_569)
);

AND2x2_ASAP7_75t_L g570 ( 
.A(n_473),
.B(n_360),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_512),
.Y(n_571)
);

CKINVDCx5p33_ASAP7_75t_R g572 ( 
.A(n_453),
.Y(n_572)
);

INVx2_ASAP7_75t_L g573 ( 
.A(n_477),
.Y(n_573)
);

CKINVDCx5p33_ASAP7_75t_R g574 ( 
.A(n_454),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_507),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_478),
.Y(n_576)
);

CKINVDCx5p33_ASAP7_75t_R g577 ( 
.A(n_462),
.Y(n_577)
);

CKINVDCx5p33_ASAP7_75t_R g578 ( 
.A(n_495),
.Y(n_578)
);

INVx3_ASAP7_75t_L g579 ( 
.A(n_479),
.Y(n_579)
);

CKINVDCx5p33_ASAP7_75t_R g580 ( 
.A(n_496),
.Y(n_580)
);

AND2x4_ASAP7_75t_L g581 ( 
.A(n_482),
.B(n_360),
.Y(n_581)
);

HB1xp67_ASAP7_75t_L g582 ( 
.A(n_492),
.Y(n_582)
);

INVx2_ASAP7_75t_L g583 ( 
.A(n_484),
.Y(n_583)
);

INVx2_ASAP7_75t_L g584 ( 
.A(n_485),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_486),
.Y(n_585)
);

AND2x2_ASAP7_75t_L g586 ( 
.A(n_467),
.B(n_350),
.Y(n_586)
);

CKINVDCx20_ASAP7_75t_R g587 ( 
.A(n_465),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_505),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_L g589 ( 
.A(n_467),
.B(n_300),
.Y(n_589)
);

CKINVDCx20_ASAP7_75t_R g590 ( 
.A(n_466),
.Y(n_590)
);

INVx4_ASAP7_75t_L g591 ( 
.A(n_559),
.Y(n_591)
);

INVx4_ASAP7_75t_SL g592 ( 
.A(n_539),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_531),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_L g594 ( 
.A(n_559),
.B(n_468),
.Y(n_594)
);

AOI22xp33_ASAP7_75t_L g595 ( 
.A1(n_575),
.A2(n_449),
.B1(n_434),
.B2(n_438),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_531),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_L g597 ( 
.A(n_559),
.B(n_468),
.Y(n_597)
);

AOI22xp33_ASAP7_75t_L g598 ( 
.A1(n_575),
.A2(n_449),
.B1(n_438),
.B2(n_441),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_531),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_SL g600 ( 
.A(n_537),
.B(n_500),
.Y(n_600)
);

OAI22xp5_ASAP7_75t_L g601 ( 
.A1(n_554),
.A2(n_501),
.B1(n_506),
.B2(n_500),
.Y(n_601)
);

BUFx6f_ASAP7_75t_L g602 ( 
.A(n_539),
.Y(n_602)
);

AO21x2_ASAP7_75t_L g603 ( 
.A1(n_552),
.A2(n_541),
.B(n_589),
.Y(n_603)
);

BUFx3_ASAP7_75t_L g604 ( 
.A(n_526),
.Y(n_604)
);

BUFx2_ASAP7_75t_L g605 ( 
.A(n_582),
.Y(n_605)
);

INVx4_ASAP7_75t_L g606 ( 
.A(n_559),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_535),
.Y(n_607)
);

BUFx6f_ASAP7_75t_L g608 ( 
.A(n_539),
.Y(n_608)
);

BUFx3_ASAP7_75t_L g609 ( 
.A(n_526),
.Y(n_609)
);

AND2x6_ASAP7_75t_L g610 ( 
.A(n_544),
.B(n_285),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_SL g611 ( 
.A(n_569),
.B(n_501),
.Y(n_611)
);

OAI221xp5_ASAP7_75t_L g612 ( 
.A1(n_554),
.A2(n_428),
.B1(n_431),
.B2(n_427),
.C(n_350),
.Y(n_612)
);

HB1xp67_ASAP7_75t_L g613 ( 
.A(n_529),
.Y(n_613)
);

INVx6_ASAP7_75t_L g614 ( 
.A(n_539),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_573),
.Y(n_615)
);

INVx5_ASAP7_75t_L g616 ( 
.A(n_539),
.Y(n_616)
);

INVx2_ASAP7_75t_L g617 ( 
.A(n_535),
.Y(n_617)
);

INVx2_ASAP7_75t_L g618 ( 
.A(n_535),
.Y(n_618)
);

OAI22xp33_ASAP7_75t_SL g619 ( 
.A1(n_578),
.A2(n_471),
.B1(n_483),
.B2(n_481),
.Y(n_619)
);

INVx3_ASAP7_75t_L g620 ( 
.A(n_539),
.Y(n_620)
);

OAI22xp33_ASAP7_75t_L g621 ( 
.A1(n_563),
.A2(n_472),
.B1(n_504),
.B2(n_450),
.Y(n_621)
);

INVx2_ASAP7_75t_SL g622 ( 
.A(n_526),
.Y(n_622)
);

AND2x2_ASAP7_75t_SL g623 ( 
.A(n_521),
.B(n_285),
.Y(n_623)
);

BUFx4f_ASAP7_75t_L g624 ( 
.A(n_555),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_545),
.Y(n_625)
);

BUFx6f_ASAP7_75t_L g626 ( 
.A(n_545),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_SL g627 ( 
.A(n_580),
.B(n_506),
.Y(n_627)
);

OR2x2_ASAP7_75t_L g628 ( 
.A(n_521),
.B(n_458),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_L g629 ( 
.A(n_550),
.B(n_471),
.Y(n_629)
);

NOR2xp33_ASAP7_75t_L g630 ( 
.A(n_551),
.B(n_508),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_545),
.Y(n_631)
);

OR2x2_ASAP7_75t_L g632 ( 
.A(n_536),
.B(n_464),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_SL g633 ( 
.A(n_586),
.B(n_508),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_L g634 ( 
.A(n_551),
.B(n_481),
.Y(n_634)
);

AOI22xp5_ASAP7_75t_SL g635 ( 
.A1(n_587),
.A2(n_469),
.B1(n_480),
.B2(n_435),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_L g636 ( 
.A(n_555),
.B(n_553),
.Y(n_636)
);

INVx2_ASAP7_75t_L g637 ( 
.A(n_523),
.Y(n_637)
);

BUFx2_ASAP7_75t_L g638 ( 
.A(n_536),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_541),
.Y(n_639)
);

NOR2xp33_ASAP7_75t_L g640 ( 
.A(n_555),
.B(n_488),
.Y(n_640)
);

OR2x2_ASAP7_75t_L g641 ( 
.A(n_522),
.B(n_519),
.Y(n_641)
);

AND2x2_ASAP7_75t_L g642 ( 
.A(n_579),
.B(n_488),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_546),
.Y(n_643)
);

INVx1_ASAP7_75t_SL g644 ( 
.A(n_590),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_L g645 ( 
.A(n_555),
.B(n_490),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_SL g646 ( 
.A(n_544),
.B(n_490),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_546),
.Y(n_647)
);

BUFx6f_ASAP7_75t_L g648 ( 
.A(n_546),
.Y(n_648)
);

AND2x6_ASAP7_75t_L g649 ( 
.A(n_555),
.B(n_311),
.Y(n_649)
);

CKINVDCx5p33_ASAP7_75t_R g650 ( 
.A(n_527),
.Y(n_650)
);

INVx2_ASAP7_75t_L g651 ( 
.A(n_523),
.Y(n_651)
);

AND2x2_ASAP7_75t_L g652 ( 
.A(n_579),
.B(n_491),
.Y(n_652)
);

INVx2_ASAP7_75t_L g653 ( 
.A(n_523),
.Y(n_653)
);

INVx3_ASAP7_75t_L g654 ( 
.A(n_546),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_L g655 ( 
.A(n_640),
.B(n_555),
.Y(n_655)
);

AND2x2_ASAP7_75t_L g656 ( 
.A(n_605),
.B(n_522),
.Y(n_656)
);

INVx2_ASAP7_75t_L g657 ( 
.A(n_617),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_L g658 ( 
.A(n_642),
.B(n_553),
.Y(n_658)
);

OR2x2_ASAP7_75t_L g659 ( 
.A(n_605),
.B(n_562),
.Y(n_659)
);

AOI22xp33_ASAP7_75t_L g660 ( 
.A1(n_623),
.A2(n_547),
.B1(n_588),
.B2(n_583),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_SL g661 ( 
.A(n_652),
.B(n_553),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_L g662 ( 
.A(n_652),
.B(n_491),
.Y(n_662)
);

INVx2_ASAP7_75t_SL g663 ( 
.A(n_624),
.Y(n_663)
);

AOI22xp5_ASAP7_75t_L g664 ( 
.A1(n_610),
.A2(n_579),
.B1(n_548),
.B2(n_576),
.Y(n_664)
);

BUFx3_ASAP7_75t_L g665 ( 
.A(n_604),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_639),
.Y(n_666)
);

INVx2_ASAP7_75t_L g667 ( 
.A(n_617),
.Y(n_667)
);

NAND2xp33_ASAP7_75t_L g668 ( 
.A(n_648),
.B(n_579),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_L g669 ( 
.A(n_629),
.B(n_630),
.Y(n_669)
);

INVx2_ASAP7_75t_L g670 ( 
.A(n_618),
.Y(n_670)
);

INVx2_ASAP7_75t_SL g671 ( 
.A(n_624),
.Y(n_671)
);

BUFx12f_ASAP7_75t_L g672 ( 
.A(n_650),
.Y(n_672)
);

INVx3_ASAP7_75t_L g673 ( 
.A(n_591),
.Y(n_673)
);

NOR2xp33_ASAP7_75t_L g674 ( 
.A(n_601),
.B(n_534),
.Y(n_674)
);

INVx2_ASAP7_75t_SL g675 ( 
.A(n_624),
.Y(n_675)
);

INVx2_ASAP7_75t_L g676 ( 
.A(n_618),
.Y(n_676)
);

BUFx6f_ASAP7_75t_L g677 ( 
.A(n_602),
.Y(n_677)
);

AND2x4_ASAP7_75t_L g678 ( 
.A(n_604),
.B(n_609),
.Y(n_678)
);

AND2x2_ASAP7_75t_L g679 ( 
.A(n_623),
.B(n_570),
.Y(n_679)
);

NAND2xp33_ASAP7_75t_L g680 ( 
.A(n_648),
.B(n_427),
.Y(n_680)
);

INVx2_ASAP7_75t_L g681 ( 
.A(n_637),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_SL g682 ( 
.A(n_621),
.B(n_542),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_L g683 ( 
.A(n_610),
.B(n_540),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_610),
.B(n_540),
.Y(n_684)
);

INVx2_ASAP7_75t_SL g685 ( 
.A(n_648),
.Y(n_685)
);

AND2x4_ASAP7_75t_L g686 ( 
.A(n_609),
.B(n_576),
.Y(n_686)
);

AND2x2_ASAP7_75t_L g687 ( 
.A(n_638),
.B(n_570),
.Y(n_687)
);

NOR2xp33_ASAP7_75t_L g688 ( 
.A(n_633),
.B(n_543),
.Y(n_688)
);

OAI22xp5_ASAP7_75t_L g689 ( 
.A1(n_645),
.A2(n_431),
.B1(n_432),
.B2(n_428),
.Y(n_689)
);

INVx2_ASAP7_75t_L g690 ( 
.A(n_637),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_L g691 ( 
.A(n_610),
.B(n_540),
.Y(n_691)
);

INVx2_ASAP7_75t_L g692 ( 
.A(n_651),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_L g693 ( 
.A(n_610),
.B(n_540),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_L g694 ( 
.A(n_610),
.B(n_549),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_SL g695 ( 
.A(n_634),
.B(n_556),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_L g696 ( 
.A(n_594),
.B(n_549),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_SL g697 ( 
.A(n_597),
.B(n_549),
.Y(n_697)
);

INVx2_ASAP7_75t_L g698 ( 
.A(n_651),
.Y(n_698)
);

INVx2_ASAP7_75t_L g699 ( 
.A(n_653),
.Y(n_699)
);

INVxp67_ASAP7_75t_L g700 ( 
.A(n_638),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_SL g701 ( 
.A(n_641),
.B(n_549),
.Y(n_701)
);

NAND2xp33_ASAP7_75t_L g702 ( 
.A(n_648),
.B(n_602),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_L g703 ( 
.A(n_639),
.B(n_548),
.Y(n_703)
);

NAND3xp33_ASAP7_75t_L g704 ( 
.A(n_595),
.B(n_585),
.C(n_567),
.Y(n_704)
);

CKINVDCx5p33_ASAP7_75t_R g705 ( 
.A(n_650),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_L g706 ( 
.A(n_654),
.B(n_585),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_593),
.Y(n_707)
);

INVx2_ASAP7_75t_SL g708 ( 
.A(n_648),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_L g709 ( 
.A(n_654),
.B(n_516),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_SL g710 ( 
.A(n_641),
.B(n_567),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_L g711 ( 
.A(n_622),
.B(n_518),
.Y(n_711)
);

AND2x2_ASAP7_75t_SL g712 ( 
.A(n_636),
.B(n_311),
.Y(n_712)
);

INVx2_ASAP7_75t_L g713 ( 
.A(n_653),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_593),
.Y(n_714)
);

INVx8_ASAP7_75t_L g715 ( 
.A(n_649),
.Y(n_715)
);

AOI221xp5_ASAP7_75t_L g716 ( 
.A1(n_598),
.A2(n_432),
.B1(n_264),
.B2(n_322),
.C(n_293),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_SL g717 ( 
.A(n_600),
.B(n_573),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_596),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_SL g719 ( 
.A(n_632),
.B(n_573),
.Y(n_719)
);

AND2x2_ASAP7_75t_L g720 ( 
.A(n_632),
.B(n_583),
.Y(n_720)
);

BUFx6f_ASAP7_75t_L g721 ( 
.A(n_602),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_SL g722 ( 
.A(n_611),
.B(n_583),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_SL g723 ( 
.A(n_627),
.B(n_584),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_SL g724 ( 
.A(n_622),
.B(n_584),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_L g725 ( 
.A(n_615),
.B(n_584),
.Y(n_725)
);

AOI22xp5_ASAP7_75t_L g726 ( 
.A1(n_646),
.A2(n_581),
.B1(n_269),
.B2(n_303),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_596),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_L g728 ( 
.A(n_643),
.B(n_588),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_643),
.Y(n_729)
);

NAND2xp33_ASAP7_75t_SL g730 ( 
.A(n_613),
.B(n_292),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_L g731 ( 
.A(n_647),
.B(n_581),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_SL g732 ( 
.A(n_619),
.B(n_274),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_SL g733 ( 
.A(n_628),
.B(n_275),
.Y(n_733)
);

INVx2_ASAP7_75t_L g734 ( 
.A(n_599),
.Y(n_734)
);

OAI22xp5_ASAP7_75t_L g735 ( 
.A1(n_612),
.A2(n_324),
.B1(n_343),
.B2(n_338),
.Y(n_735)
);

NOR2xp33_ASAP7_75t_R g736 ( 
.A(n_644),
.B(n_572),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_L g737 ( 
.A(n_647),
.B(n_581),
.Y(n_737)
);

AOI21xp5_ASAP7_75t_L g738 ( 
.A1(n_655),
.A2(n_606),
.B(n_591),
.Y(n_738)
);

AOI21xp5_ASAP7_75t_L g739 ( 
.A1(n_658),
.A2(n_606),
.B(n_620),
.Y(n_739)
);

NOR2xp33_ASAP7_75t_L g740 ( 
.A(n_669),
.B(n_574),
.Y(n_740)
);

AOI21xp33_ASAP7_75t_L g741 ( 
.A1(n_660),
.A2(n_603),
.B(n_599),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_L g742 ( 
.A(n_662),
.B(n_607),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_SL g743 ( 
.A(n_678),
.B(n_628),
.Y(n_743)
);

AOI21xp5_ASAP7_75t_L g744 ( 
.A1(n_703),
.A2(n_620),
.B(n_603),
.Y(n_744)
);

AOI21xp5_ASAP7_75t_L g745 ( 
.A1(n_673),
.A2(n_603),
.B(n_607),
.Y(n_745)
);

OAI21xp33_ASAP7_75t_L g746 ( 
.A1(n_674),
.A2(n_347),
.B(n_346),
.Y(n_746)
);

AO21x1_ASAP7_75t_L g747 ( 
.A1(n_666),
.A2(n_631),
.B(n_625),
.Y(n_747)
);

OAI21xp5_ASAP7_75t_L g748 ( 
.A1(n_666),
.A2(n_552),
.B(n_625),
.Y(n_748)
);

INVx4_ASAP7_75t_L g749 ( 
.A(n_715),
.Y(n_749)
);

NAND3xp33_ASAP7_75t_L g750 ( 
.A(n_700),
.B(n_705),
.C(n_716),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_L g751 ( 
.A(n_720),
.B(n_631),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_707),
.Y(n_752)
);

O2A1O1Ixp33_ASAP7_75t_L g753 ( 
.A1(n_710),
.A2(n_560),
.B(n_565),
.C(n_557),
.Y(n_753)
);

INVx4_ASAP7_75t_L g754 ( 
.A(n_715),
.Y(n_754)
);

AND2x2_ASAP7_75t_L g755 ( 
.A(n_656),
.B(n_577),
.Y(n_755)
);

BUFx12f_ASAP7_75t_L g756 ( 
.A(n_672),
.Y(n_756)
);

AOI21x1_ASAP7_75t_L g757 ( 
.A1(n_661),
.A2(n_547),
.B(n_525),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_L g758 ( 
.A(n_679),
.B(n_649),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_L g759 ( 
.A(n_679),
.B(n_649),
.Y(n_759)
);

AOI21x1_ASAP7_75t_L g760 ( 
.A1(n_725),
.A2(n_547),
.B(n_525),
.Y(n_760)
);

INVx2_ASAP7_75t_L g761 ( 
.A(n_681),
.Y(n_761)
);

OAI321xp33_ASAP7_75t_L g762 ( 
.A1(n_735),
.A2(n_568),
.A3(n_560),
.B1(n_565),
.B2(n_566),
.C(n_571),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_L g763 ( 
.A(n_686),
.B(n_687),
.Y(n_763)
);

NOR2xp33_ASAP7_75t_L g764 ( 
.A(n_659),
.B(n_561),
.Y(n_764)
);

INVx2_ASAP7_75t_L g765 ( 
.A(n_681),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_L g766 ( 
.A(n_686),
.B(n_649),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_L g767 ( 
.A(n_686),
.B(n_649),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_707),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_L g769 ( 
.A(n_687),
.B(n_626),
.Y(n_769)
);

AO32x1_ASAP7_75t_L g770 ( 
.A1(n_714),
.A2(n_533),
.A3(n_538),
.B1(n_532),
.B2(n_524),
.Y(n_770)
);

OAI21xp5_ASAP7_75t_L g771 ( 
.A1(n_714),
.A2(n_547),
.B(n_616),
.Y(n_771)
);

AOI21xp5_ASAP7_75t_L g772 ( 
.A1(n_702),
.A2(n_608),
.B(n_626),
.Y(n_772)
);

NOR2xp33_ASAP7_75t_L g773 ( 
.A(n_659),
.B(n_558),
.Y(n_773)
);

BUFx6f_ASAP7_75t_L g774 ( 
.A(n_677),
.Y(n_774)
);

OAI22xp5_ASAP7_75t_L g775 ( 
.A1(n_704),
.A2(n_363),
.B1(n_371),
.B2(n_357),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_L g776 ( 
.A(n_656),
.B(n_626),
.Y(n_776)
);

A2O1A1Ixp33_ASAP7_75t_L g777 ( 
.A1(n_664),
.A2(n_566),
.B(n_568),
.C(n_557),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_L g778 ( 
.A(n_711),
.B(n_571),
.Y(n_778)
);

INVx1_ASAP7_75t_SL g779 ( 
.A(n_736),
.Y(n_779)
);

O2A1O1Ixp33_ASAP7_75t_SL g780 ( 
.A1(n_685),
.A2(n_269),
.B(n_303),
.C(n_289),
.Y(n_780)
);

INVx2_ASAP7_75t_L g781 ( 
.A(n_690),
.Y(n_781)
);

NAND3xp33_ASAP7_75t_L g782 ( 
.A(n_705),
.B(n_558),
.C(n_635),
.Y(n_782)
);

AOI22xp33_ASAP7_75t_L g783 ( 
.A1(n_712),
.A2(n_528),
.B1(n_564),
.B2(n_614),
.Y(n_783)
);

AOI21xp5_ASAP7_75t_L g784 ( 
.A1(n_706),
.A2(n_616),
.B(n_424),
.Y(n_784)
);

AOI21x1_ASAP7_75t_L g785 ( 
.A1(n_724),
.A2(n_532),
.B(n_524),
.Y(n_785)
);

INVx3_ASAP7_75t_L g786 ( 
.A(n_678),
.Y(n_786)
);

AOI21xp5_ASAP7_75t_L g787 ( 
.A1(n_668),
.A2(n_708),
.B(n_685),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_L g788 ( 
.A(n_728),
.B(n_564),
.Y(n_788)
);

AOI21x1_ASAP7_75t_L g789 ( 
.A1(n_718),
.A2(n_538),
.B(n_533),
.Y(n_789)
);

A2O1A1Ixp33_ASAP7_75t_L g790 ( 
.A1(n_688),
.A2(n_302),
.B(n_308),
.C(n_307),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_SL g791 ( 
.A(n_678),
.B(n_616),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_718),
.Y(n_792)
);

OAI21xp33_ASAP7_75t_L g793 ( 
.A1(n_689),
.A2(n_374),
.B(n_373),
.Y(n_793)
);

AOI21x1_ASAP7_75t_L g794 ( 
.A1(n_727),
.A2(n_729),
.B(n_731),
.Y(n_794)
);

INVx4_ASAP7_75t_L g795 ( 
.A(n_715),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_L g796 ( 
.A(n_719),
.B(n_564),
.Y(n_796)
);

OAI22xp5_ASAP7_75t_L g797 ( 
.A1(n_727),
.A2(n_395),
.B1(n_403),
.B2(n_390),
.Y(n_797)
);

AOI21xp5_ASAP7_75t_L g798 ( 
.A1(n_668),
.A2(n_616),
.B(n_424),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_L g799 ( 
.A(n_709),
.B(n_614),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_L g800 ( 
.A(n_734),
.B(n_614),
.Y(n_800)
);

NOR2xp33_ASAP7_75t_L g801 ( 
.A(n_695),
.B(n_528),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_L g802 ( 
.A(n_734),
.B(n_614),
.Y(n_802)
);

O2A1O1Ixp33_ASAP7_75t_L g803 ( 
.A1(n_737),
.A2(n_309),
.B(n_316),
.C(n_312),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_SL g804 ( 
.A(n_665),
.B(n_663),
.Y(n_804)
);

AOI21xp5_ASAP7_75t_L g805 ( 
.A1(n_708),
.A2(n_429),
.B(n_275),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_L g806 ( 
.A(n_712),
.B(n_592),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_657),
.Y(n_807)
);

AOI21xp5_ASAP7_75t_L g808 ( 
.A1(n_663),
.A2(n_429),
.B(n_265),
.Y(n_808)
);

OR2x6_ASAP7_75t_L g809 ( 
.A(n_715),
.B(n_289),
.Y(n_809)
);

INVx2_ASAP7_75t_SL g810 ( 
.A(n_701),
.Y(n_810)
);

O2A1O1Ixp33_ASAP7_75t_L g811 ( 
.A1(n_723),
.A2(n_321),
.B(n_339),
.C(n_318),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_L g812 ( 
.A(n_696),
.B(n_592),
.Y(n_812)
);

AND2x2_ASAP7_75t_L g813 ( 
.A(n_733),
.B(n_407),
.Y(n_813)
);

NOR2xp33_ASAP7_75t_L g814 ( 
.A(n_682),
.B(n_408),
.Y(n_814)
);

OAI21xp5_ASAP7_75t_L g815 ( 
.A1(n_657),
.A2(n_670),
.B(n_667),
.Y(n_815)
);

OAI22xp5_ASAP7_75t_L g816 ( 
.A1(n_726),
.A2(n_675),
.B1(n_671),
.B2(n_677),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_L g817 ( 
.A(n_671),
.B(n_592),
.Y(n_817)
);

CKINVDCx8_ASAP7_75t_R g818 ( 
.A(n_677),
.Y(n_818)
);

O2A1O1Ixp33_ASAP7_75t_L g819 ( 
.A1(n_680),
.A2(n_352),
.B(n_368),
.C(n_340),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_SL g820 ( 
.A(n_675),
.B(n_411),
.Y(n_820)
);

OAI21xp5_ASAP7_75t_L g821 ( 
.A1(n_667),
.A2(n_376),
.B(n_369),
.Y(n_821)
);

OAI22xp5_ASAP7_75t_L g822 ( 
.A1(n_677),
.A2(n_415),
.B1(n_421),
.B2(n_413),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_L g823 ( 
.A(n_670),
.B(n_676),
.Y(n_823)
);

INVx2_ASAP7_75t_L g824 ( 
.A(n_690),
.Y(n_824)
);

OAI22xp5_ASAP7_75t_L g825 ( 
.A1(n_677),
.A2(n_379),
.B1(n_405),
.B2(n_398),
.Y(n_825)
);

INVx2_ASAP7_75t_L g826 ( 
.A(n_692),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_L g827 ( 
.A(n_676),
.B(n_722),
.Y(n_827)
);

BUFx3_ASAP7_75t_L g828 ( 
.A(n_756),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_L g829 ( 
.A(n_740),
.B(n_763),
.Y(n_829)
);

OAI21xp5_ASAP7_75t_L g830 ( 
.A1(n_744),
.A2(n_717),
.B(n_698),
.Y(n_830)
);

AOI21xp5_ASAP7_75t_L g831 ( 
.A1(n_738),
.A2(n_721),
.B(n_680),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_L g832 ( 
.A(n_752),
.B(n_692),
.Y(n_832)
);

O2A1O1Ixp5_ASAP7_75t_L g833 ( 
.A1(n_747),
.A2(n_697),
.B(n_732),
.C(n_730),
.Y(n_833)
);

OAI21x1_ASAP7_75t_L g834 ( 
.A1(n_745),
.A2(n_699),
.B(n_698),
.Y(n_834)
);

BUFx6f_ASAP7_75t_L g835 ( 
.A(n_818),
.Y(n_835)
);

AOI21xp5_ASAP7_75t_L g836 ( 
.A1(n_739),
.A2(n_721),
.B(n_684),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_768),
.Y(n_837)
);

BUFx6f_ASAP7_75t_L g838 ( 
.A(n_774),
.Y(n_838)
);

AND2x2_ASAP7_75t_L g839 ( 
.A(n_755),
.B(n_773),
.Y(n_839)
);

AO31x2_ASAP7_75t_L g840 ( 
.A1(n_777),
.A2(n_825),
.A3(n_812),
.B(n_816),
.Y(n_840)
);

AND2x2_ASAP7_75t_L g841 ( 
.A(n_764),
.B(n_699),
.Y(n_841)
);

AO31x2_ASAP7_75t_L g842 ( 
.A1(n_825),
.A2(n_713),
.A3(n_683),
.B(n_693),
.Y(n_842)
);

INVx3_ASAP7_75t_L g843 ( 
.A(n_749),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_L g844 ( 
.A(n_792),
.B(n_713),
.Y(n_844)
);

OAI21x1_ASAP7_75t_L g845 ( 
.A1(n_748),
.A2(n_760),
.B(n_789),
.Y(n_845)
);

INVx3_ASAP7_75t_L g846 ( 
.A(n_749),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_L g847 ( 
.A(n_751),
.B(n_721),
.Y(n_847)
);

AOI21xp33_ASAP7_75t_L g848 ( 
.A1(n_819),
.A2(n_694),
.B(n_691),
.Y(n_848)
);

AND2x2_ASAP7_75t_L g849 ( 
.A(n_743),
.B(n_530),
.Y(n_849)
);

AOI22xp5_ASAP7_75t_L g850 ( 
.A1(n_750),
.A2(n_730),
.B1(n_721),
.B2(n_417),
.Y(n_850)
);

OR2x6_ASAP7_75t_L g851 ( 
.A(n_782),
.B(n_721),
.Y(n_851)
);

OAI21xp5_ASAP7_75t_L g852 ( 
.A1(n_748),
.A2(n_420),
.B(n_394),
.Y(n_852)
);

OAI21x1_ASAP7_75t_L g853 ( 
.A1(n_772),
.A2(n_530),
.B(n_402),
.Y(n_853)
);

OAI22xp5_ASAP7_75t_L g854 ( 
.A1(n_742),
.A2(n_402),
.B1(n_423),
.B2(n_367),
.Y(n_854)
);

OAI21xp5_ASAP7_75t_L g855 ( 
.A1(n_741),
.A2(n_423),
.B(n_367),
.Y(n_855)
);

AO21x1_ASAP7_75t_L g856 ( 
.A1(n_816),
.A2(n_530),
.B(n_406),
.Y(n_856)
);

AOI21x1_ASAP7_75t_L g857 ( 
.A1(n_794),
.A2(n_785),
.B(n_757),
.Y(n_857)
);

BUFx2_ASAP7_75t_L g858 ( 
.A(n_779),
.Y(n_858)
);

AO21x1_ASAP7_75t_L g859 ( 
.A1(n_821),
.A2(n_406),
.B(n_400),
.Y(n_859)
);

NAND2x1p5_ASAP7_75t_L g860 ( 
.A(n_754),
.B(n_400),
.Y(n_860)
);

AOI21xp33_ASAP7_75t_L g861 ( 
.A1(n_803),
.A2(n_425),
.B(n_279),
.Y(n_861)
);

AOI22xp5_ASAP7_75t_L g862 ( 
.A1(n_746),
.A2(n_328),
.B1(n_351),
.B2(n_262),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_L g863 ( 
.A(n_776),
.B(n_425),
.Y(n_863)
);

BUFx2_ASAP7_75t_L g864 ( 
.A(n_786),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_L g865 ( 
.A(n_778),
.B(n_4),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_796),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_L g867 ( 
.A(n_769),
.B(n_5),
.Y(n_867)
);

OAI21x1_ASAP7_75t_L g868 ( 
.A1(n_815),
.A2(n_410),
.B(n_314),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_807),
.Y(n_869)
);

INVxp67_ASAP7_75t_L g870 ( 
.A(n_810),
.Y(n_870)
);

BUFx6f_ASAP7_75t_L g871 ( 
.A(n_774),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_L g872 ( 
.A(n_814),
.B(n_5),
.Y(n_872)
);

OAI21x1_ASAP7_75t_L g873 ( 
.A1(n_815),
.A2(n_410),
.B(n_314),
.Y(n_873)
);

AND2x2_ASAP7_75t_SL g874 ( 
.A(n_801),
.B(n_783),
.Y(n_874)
);

AOI21x1_ASAP7_75t_L g875 ( 
.A1(n_788),
.A2(n_410),
.B(n_314),
.Y(n_875)
);

OAI22xp5_ASAP7_75t_L g876 ( 
.A1(n_790),
.A2(n_283),
.B1(n_286),
.B2(n_282),
.Y(n_876)
);

INVx2_ASAP7_75t_L g877 ( 
.A(n_761),
.Y(n_877)
);

NOR2xp33_ASAP7_75t_L g878 ( 
.A(n_797),
.B(n_290),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_753),
.Y(n_879)
);

AOI21xp5_ASAP7_75t_L g880 ( 
.A1(n_787),
.A2(n_296),
.B(n_295),
.Y(n_880)
);

AOI21xp5_ASAP7_75t_L g881 ( 
.A1(n_799),
.A2(n_298),
.B(n_297),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_L g882 ( 
.A(n_765),
.B(n_6),
.Y(n_882)
);

INVxp67_ASAP7_75t_SL g883 ( 
.A(n_774),
.Y(n_883)
);

AO31x2_ASAP7_75t_L g884 ( 
.A1(n_823),
.A2(n_139),
.A3(n_260),
.B(n_259),
.Y(n_884)
);

INVx2_ASAP7_75t_L g885 ( 
.A(n_781),
.Y(n_885)
);

AOI21xp5_ASAP7_75t_L g886 ( 
.A1(n_784),
.A2(n_304),
.B(n_299),
.Y(n_886)
);

INVx2_ASAP7_75t_L g887 ( 
.A(n_824),
.Y(n_887)
);

AND2x2_ASAP7_75t_L g888 ( 
.A(n_813),
.B(n_797),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_826),
.Y(n_889)
);

AOI21xp5_ASAP7_75t_SL g890 ( 
.A1(n_795),
.A2(n_306),
.B(n_305),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_L g891 ( 
.A(n_758),
.B(n_6),
.Y(n_891)
);

INVx1_ASAP7_75t_L g892 ( 
.A(n_827),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_L g893 ( 
.A(n_759),
.B(n_7),
.Y(n_893)
);

A2O1A1Ixp33_ASAP7_75t_L g894 ( 
.A1(n_762),
.A2(n_419),
.B(n_418),
.C(n_416),
.Y(n_894)
);

OAI21x1_ASAP7_75t_L g895 ( 
.A1(n_771),
.A2(n_84),
.B(n_79),
.Y(n_895)
);

AND2x2_ASAP7_75t_L g896 ( 
.A(n_775),
.B(n_822),
.Y(n_896)
);

INVx2_ASAP7_75t_L g897 ( 
.A(n_800),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_L g898 ( 
.A(n_821),
.B(n_8),
.Y(n_898)
);

NAND2xp5_ASAP7_75t_L g899 ( 
.A(n_822),
.B(n_8),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_L g900 ( 
.A(n_802),
.B(n_10),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_L g901 ( 
.A(n_766),
.B(n_10),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_L g902 ( 
.A(n_767),
.B(n_12),
.Y(n_902)
);

AO31x2_ASAP7_75t_L g903 ( 
.A1(n_806),
.A2(n_137),
.A3(n_256),
.B(n_255),
.Y(n_903)
);

OAI22xp5_ASAP7_75t_L g904 ( 
.A1(n_809),
.A2(n_353),
.B1(n_412),
.B2(n_409),
.Y(n_904)
);

AO31x2_ASAP7_75t_L g905 ( 
.A1(n_741),
.A2(n_126),
.A3(n_253),
.B(n_249),
.Y(n_905)
);

BUFx2_ASAP7_75t_L g906 ( 
.A(n_809),
.Y(n_906)
);

OAI21x1_ASAP7_75t_L g907 ( 
.A1(n_771),
.A2(n_88),
.B(n_87),
.Y(n_907)
);

OAI21x1_ASAP7_75t_L g908 ( 
.A1(n_817),
.A2(n_90),
.B(n_89),
.Y(n_908)
);

AOI21xp5_ASAP7_75t_L g909 ( 
.A1(n_820),
.A2(n_317),
.B(n_310),
.Y(n_909)
);

OAI21x1_ASAP7_75t_SL g910 ( 
.A1(n_811),
.A2(n_13),
.B(n_14),
.Y(n_910)
);

AOI21xp5_ASAP7_75t_L g911 ( 
.A1(n_804),
.A2(n_323),
.B(n_320),
.Y(n_911)
);

OR2x6_ASAP7_75t_L g912 ( 
.A(n_835),
.B(n_851),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_L g913 ( 
.A(n_829),
.B(n_775),
.Y(n_913)
);

INVx1_ASAP7_75t_L g914 ( 
.A(n_837),
.Y(n_914)
);

BUFx2_ASAP7_75t_L g915 ( 
.A(n_858),
.Y(n_915)
);

AND2x4_ASAP7_75t_L g916 ( 
.A(n_835),
.B(n_791),
.Y(n_916)
);

INVx2_ASAP7_75t_L g917 ( 
.A(n_877),
.Y(n_917)
);

INVx2_ASAP7_75t_L g918 ( 
.A(n_885),
.Y(n_918)
);

INVx1_ASAP7_75t_L g919 ( 
.A(n_869),
.Y(n_919)
);

AND2x4_ASAP7_75t_L g920 ( 
.A(n_835),
.B(n_798),
.Y(n_920)
);

NAND2xp5_ASAP7_75t_L g921 ( 
.A(n_892),
.B(n_780),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_L g922 ( 
.A(n_896),
.B(n_866),
.Y(n_922)
);

OAI22xp5_ASAP7_75t_L g923 ( 
.A1(n_872),
.A2(n_793),
.B1(n_805),
.B2(n_808),
.Y(n_923)
);

INVx1_ASAP7_75t_L g924 ( 
.A(n_889),
.Y(n_924)
);

BUFx6f_ASAP7_75t_L g925 ( 
.A(n_838),
.Y(n_925)
);

OAI22xp5_ASAP7_75t_L g926 ( 
.A1(n_898),
.A2(n_865),
.B1(n_878),
.B2(n_899),
.Y(n_926)
);

NAND2xp5_ASAP7_75t_L g927 ( 
.A(n_847),
.B(n_13),
.Y(n_927)
);

O2A1O1Ixp5_ASAP7_75t_L g928 ( 
.A1(n_852),
.A2(n_770),
.B(n_15),
.C(n_16),
.Y(n_928)
);

OR2x2_ASAP7_75t_L g929 ( 
.A(n_839),
.B(n_14),
.Y(n_929)
);

INVx3_ASAP7_75t_L g930 ( 
.A(n_843),
.Y(n_930)
);

INVx2_ASAP7_75t_L g931 ( 
.A(n_887),
.Y(n_931)
);

INVx1_ASAP7_75t_L g932 ( 
.A(n_882),
.Y(n_932)
);

INVx1_ASAP7_75t_L g933 ( 
.A(n_882),
.Y(n_933)
);

BUFx6f_ASAP7_75t_L g934 ( 
.A(n_838),
.Y(n_934)
);

BUFx3_ASAP7_75t_L g935 ( 
.A(n_828),
.Y(n_935)
);

NAND2xp5_ASAP7_75t_L g936 ( 
.A(n_847),
.B(n_20),
.Y(n_936)
);

NAND2xp5_ASAP7_75t_L g937 ( 
.A(n_832),
.B(n_20),
.Y(n_937)
);

NAND2xp5_ASAP7_75t_L g938 ( 
.A(n_841),
.B(n_21),
.Y(n_938)
);

INVx1_ASAP7_75t_L g939 ( 
.A(n_832),
.Y(n_939)
);

INVx1_ASAP7_75t_L g940 ( 
.A(n_844),
.Y(n_940)
);

AO32x2_ASAP7_75t_L g941 ( 
.A1(n_854),
.A2(n_770),
.A3(n_23),
.B1(n_24),
.B2(n_25),
.Y(n_941)
);

INVx1_ASAP7_75t_SL g942 ( 
.A(n_864),
.Y(n_942)
);

OAI21xp33_ASAP7_75t_L g943 ( 
.A1(n_898),
.A2(n_326),
.B(n_325),
.Y(n_943)
);

NAND2xp5_ASAP7_75t_L g944 ( 
.A(n_897),
.B(n_22),
.Y(n_944)
);

INVx1_ASAP7_75t_SL g945 ( 
.A(n_906),
.Y(n_945)
);

INVx5_ASAP7_75t_L g946 ( 
.A(n_838),
.Y(n_946)
);

AOI221xp5_ASAP7_75t_L g947 ( 
.A1(n_888),
.A2(n_356),
.B1(n_414),
.B2(n_396),
.C(n_393),
.Y(n_947)
);

AOI22xp5_ASAP7_75t_L g948 ( 
.A1(n_874),
.A2(n_354),
.B1(n_391),
.B2(n_389),
.Y(n_948)
);

O2A1O1Ixp33_ASAP7_75t_L g949 ( 
.A1(n_852),
.A2(n_770),
.B(n_27),
.C(n_28),
.Y(n_949)
);

AOI22xp33_ASAP7_75t_L g950 ( 
.A1(n_862),
.A2(n_383),
.B1(n_382),
.B2(n_381),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_SL g951 ( 
.A(n_850),
.B(n_365),
.Y(n_951)
);

INVx2_ASAP7_75t_SL g952 ( 
.A(n_851),
.Y(n_952)
);

INVx5_ASAP7_75t_L g953 ( 
.A(n_871),
.Y(n_953)
);

AND2x2_ASAP7_75t_L g954 ( 
.A(n_870),
.B(n_26),
.Y(n_954)
);

AOI21xp33_ASAP7_75t_SL g955 ( 
.A1(n_904),
.A2(n_27),
.B(n_28),
.Y(n_955)
);

AND2x2_ASAP7_75t_L g956 ( 
.A(n_851),
.B(n_29),
.Y(n_956)
);

BUFx6f_ASAP7_75t_L g957 ( 
.A(n_871),
.Y(n_957)
);

NAND2xp5_ASAP7_75t_L g958 ( 
.A(n_879),
.B(n_29),
.Y(n_958)
);

BUFx8_ASAP7_75t_L g959 ( 
.A(n_871),
.Y(n_959)
);

INVx3_ASAP7_75t_L g960 ( 
.A(n_846),
.Y(n_960)
);

BUFx2_ASAP7_75t_L g961 ( 
.A(n_883),
.Y(n_961)
);

INVx2_ASAP7_75t_L g962 ( 
.A(n_849),
.Y(n_962)
);

INVx1_ASAP7_75t_L g963 ( 
.A(n_867),
.Y(n_963)
);

INVx1_ASAP7_75t_L g964 ( 
.A(n_867),
.Y(n_964)
);

INVx1_ASAP7_75t_L g965 ( 
.A(n_900),
.Y(n_965)
);

OR2x2_ASAP7_75t_L g966 ( 
.A(n_901),
.B(n_30),
.Y(n_966)
);

BUFx2_ASAP7_75t_L g967 ( 
.A(n_860),
.Y(n_967)
);

INVx1_ASAP7_75t_L g968 ( 
.A(n_900),
.Y(n_968)
);

INVx1_ASAP7_75t_L g969 ( 
.A(n_901),
.Y(n_969)
);

NAND2xp5_ASAP7_75t_L g970 ( 
.A(n_891),
.B(n_31),
.Y(n_970)
);

OR2x6_ASAP7_75t_SL g971 ( 
.A(n_876),
.B(n_854),
.Y(n_971)
);

BUFx8_ASAP7_75t_SL g972 ( 
.A(n_902),
.Y(n_972)
);

AOI221xp5_ASAP7_75t_L g973 ( 
.A1(n_876),
.A2(n_359),
.B1(n_355),
.B2(n_348),
.C(n_345),
.Y(n_973)
);

INVx2_ASAP7_75t_SL g974 ( 
.A(n_902),
.Y(n_974)
);

INVxp67_ASAP7_75t_SL g975 ( 
.A(n_891),
.Y(n_975)
);

CKINVDCx20_ASAP7_75t_R g976 ( 
.A(n_890),
.Y(n_976)
);

NOR2xp33_ASAP7_75t_L g977 ( 
.A(n_893),
.B(n_344),
.Y(n_977)
);

OA21x2_ASAP7_75t_L g978 ( 
.A1(n_845),
.A2(n_342),
.B(n_341),
.Y(n_978)
);

AND2x2_ASAP7_75t_L g979 ( 
.A(n_861),
.B(n_32),
.Y(n_979)
);

NAND2xp5_ASAP7_75t_L g980 ( 
.A(n_893),
.B(n_32),
.Y(n_980)
);

AOI22xp33_ASAP7_75t_L g981 ( 
.A1(n_861),
.A2(n_336),
.B1(n_334),
.B2(n_333),
.Y(n_981)
);

CKINVDCx5p33_ASAP7_75t_R g982 ( 
.A(n_911),
.Y(n_982)
);

BUFx4f_ASAP7_75t_L g983 ( 
.A(n_833),
.Y(n_983)
);

BUFx6f_ASAP7_75t_L g984 ( 
.A(n_908),
.Y(n_984)
);

AOI22xp33_ASAP7_75t_L g985 ( 
.A1(n_855),
.A2(n_331),
.B1(n_327),
.B2(n_35),
.Y(n_985)
);

INVx1_ASAP7_75t_L g986 ( 
.A(n_863),
.Y(n_986)
);

INVx4_ASAP7_75t_SL g987 ( 
.A(n_903),
.Y(n_987)
);

BUFx6f_ASAP7_75t_L g988 ( 
.A(n_895),
.Y(n_988)
);

OR2x6_ASAP7_75t_L g989 ( 
.A(n_910),
.B(n_33),
.Y(n_989)
);

A2O1A1Ixp33_ASAP7_75t_L g990 ( 
.A1(n_894),
.A2(n_34),
.B(n_35),
.C(n_36),
.Y(n_990)
);

BUFx3_ASAP7_75t_L g991 ( 
.A(n_863),
.Y(n_991)
);

INVxp67_ASAP7_75t_SL g992 ( 
.A(n_830),
.Y(n_992)
);

BUFx2_ASAP7_75t_L g993 ( 
.A(n_840),
.Y(n_993)
);

INVx1_ASAP7_75t_L g994 ( 
.A(n_830),
.Y(n_994)
);

AND2x2_ASAP7_75t_L g995 ( 
.A(n_909),
.B(n_36),
.Y(n_995)
);

OR2x2_ASAP7_75t_L g996 ( 
.A(n_840),
.B(n_37),
.Y(n_996)
);

BUFx6f_ASAP7_75t_L g997 ( 
.A(n_907),
.Y(n_997)
);

AOI21xp5_ASAP7_75t_L g998 ( 
.A1(n_836),
.A2(n_120),
.B(n_246),
.Y(n_998)
);

AOI21xp5_ASAP7_75t_L g999 ( 
.A1(n_831),
.A2(n_117),
.B(n_242),
.Y(n_999)
);

HB1xp67_ASAP7_75t_L g1000 ( 
.A(n_840),
.Y(n_1000)
);

INVx1_ASAP7_75t_L g1001 ( 
.A(n_834),
.Y(n_1001)
);

BUFx3_ASAP7_75t_L g1002 ( 
.A(n_903),
.Y(n_1002)
);

NAND2xp5_ASAP7_75t_SL g1003 ( 
.A(n_848),
.B(n_859),
.Y(n_1003)
);

INVx1_ASAP7_75t_L g1004 ( 
.A(n_884),
.Y(n_1004)
);

BUFx3_ASAP7_75t_L g1005 ( 
.A(n_903),
.Y(n_1005)
);

NAND2xp5_ASAP7_75t_L g1006 ( 
.A(n_855),
.B(n_37),
.Y(n_1006)
);

BUFx2_ASAP7_75t_SL g1007 ( 
.A(n_856),
.Y(n_1007)
);

HB1xp67_ASAP7_75t_L g1008 ( 
.A(n_842),
.Y(n_1008)
);

AND2x4_ASAP7_75t_L g1009 ( 
.A(n_842),
.B(n_248),
.Y(n_1009)
);

INVx1_ASAP7_75t_SL g1010 ( 
.A(n_915),
.Y(n_1010)
);

AOI22xp33_ASAP7_75t_L g1011 ( 
.A1(n_926),
.A2(n_848),
.B1(n_881),
.B2(n_886),
.Y(n_1011)
);

INVx1_ASAP7_75t_L g1012 ( 
.A(n_1000),
.Y(n_1012)
);

INVx2_ASAP7_75t_L g1013 ( 
.A(n_1004),
.Y(n_1013)
);

INVx1_ASAP7_75t_L g1014 ( 
.A(n_993),
.Y(n_1014)
);

INVx1_ASAP7_75t_L g1015 ( 
.A(n_1008),
.Y(n_1015)
);

CKINVDCx20_ASAP7_75t_R g1016 ( 
.A(n_935),
.Y(n_1016)
);

OAI21x1_ASAP7_75t_L g1017 ( 
.A1(n_1001),
.A2(n_873),
.B(n_868),
.Y(n_1017)
);

AOI22xp33_ASAP7_75t_L g1018 ( 
.A1(n_948),
.A2(n_880),
.B1(n_853),
.B2(n_905),
.Y(n_1018)
);

HB1xp67_ASAP7_75t_L g1019 ( 
.A(n_942),
.Y(n_1019)
);

BUFx6f_ASAP7_75t_L g1020 ( 
.A(n_925),
.Y(n_1020)
);

INVx2_ASAP7_75t_L g1021 ( 
.A(n_919),
.Y(n_1021)
);

INVx2_ASAP7_75t_L g1022 ( 
.A(n_924),
.Y(n_1022)
);

INVx3_ASAP7_75t_L g1023 ( 
.A(n_983),
.Y(n_1023)
);

BUFx8_ASAP7_75t_SL g1024 ( 
.A(n_976),
.Y(n_1024)
);

INVx2_ASAP7_75t_L g1025 ( 
.A(n_939),
.Y(n_1025)
);

AOI22xp33_ASAP7_75t_L g1026 ( 
.A1(n_948),
.A2(n_905),
.B1(n_842),
.B2(n_884),
.Y(n_1026)
);

INVx1_ASAP7_75t_L g1027 ( 
.A(n_994),
.Y(n_1027)
);

AOI22xp33_ASAP7_75t_L g1028 ( 
.A1(n_943),
.A2(n_905),
.B1(n_857),
.B2(n_875),
.Y(n_1028)
);

INVxp67_ASAP7_75t_L g1029 ( 
.A(n_929),
.Y(n_1029)
);

AND2x4_ASAP7_75t_L g1030 ( 
.A(n_912),
.B(n_91),
.Y(n_1030)
);

AOI22xp33_ASAP7_75t_L g1031 ( 
.A1(n_943),
.A2(n_38),
.B1(n_39),
.B2(n_40),
.Y(n_1031)
);

INVx1_ASAP7_75t_L g1032 ( 
.A(n_969),
.Y(n_1032)
);

INVx2_ASAP7_75t_L g1033 ( 
.A(n_940),
.Y(n_1033)
);

INVx1_ASAP7_75t_L g1034 ( 
.A(n_963),
.Y(n_1034)
);

INVx1_ASAP7_75t_L g1035 ( 
.A(n_964),
.Y(n_1035)
);

INVx1_ASAP7_75t_L g1036 ( 
.A(n_932),
.Y(n_1036)
);

AOI21x1_ASAP7_75t_L g1037 ( 
.A1(n_1003),
.A2(n_240),
.B(n_121),
.Y(n_1037)
);

INVx4_ASAP7_75t_L g1038 ( 
.A(n_946),
.Y(n_1038)
);

AND2x2_ASAP7_75t_L g1039 ( 
.A(n_996),
.B(n_922),
.Y(n_1039)
);

NAND2x1p5_ASAP7_75t_L g1040 ( 
.A(n_983),
.B(n_93),
.Y(n_1040)
);

OAI21x1_ASAP7_75t_L g1041 ( 
.A1(n_998),
.A2(n_122),
.B(n_234),
.Y(n_1041)
);

OAI21x1_ASAP7_75t_L g1042 ( 
.A1(n_999),
.A2(n_111),
.B(n_233),
.Y(n_1042)
);

INVx1_ASAP7_75t_L g1043 ( 
.A(n_933),
.Y(n_1043)
);

AOI21x1_ASAP7_75t_L g1044 ( 
.A1(n_978),
.A2(n_110),
.B(n_228),
.Y(n_1044)
);

INVx1_ASAP7_75t_L g1045 ( 
.A(n_992),
.Y(n_1045)
);

NOR2x1_ASAP7_75t_L g1046 ( 
.A(n_991),
.B(n_96),
.Y(n_1046)
);

INVx1_ASAP7_75t_L g1047 ( 
.A(n_965),
.Y(n_1047)
);

INVx3_ASAP7_75t_L g1048 ( 
.A(n_925),
.Y(n_1048)
);

INVx1_ASAP7_75t_L g1049 ( 
.A(n_968),
.Y(n_1049)
);

INVx1_ASAP7_75t_L g1050 ( 
.A(n_986),
.Y(n_1050)
);

OAI21x1_ASAP7_75t_L g1051 ( 
.A1(n_928),
.A2(n_109),
.B(n_224),
.Y(n_1051)
);

INVx1_ASAP7_75t_L g1052 ( 
.A(n_975),
.Y(n_1052)
);

HB1xp67_ASAP7_75t_L g1053 ( 
.A(n_942),
.Y(n_1053)
);

INVx1_ASAP7_75t_L g1054 ( 
.A(n_1002),
.Y(n_1054)
);

INVx1_ASAP7_75t_L g1055 ( 
.A(n_1005),
.Y(n_1055)
);

CKINVDCx11_ASAP7_75t_R g1056 ( 
.A(n_945),
.Y(n_1056)
);

AOI21x1_ASAP7_75t_L g1057 ( 
.A1(n_978),
.A2(n_238),
.B(n_106),
.Y(n_1057)
);

INVx4_ASAP7_75t_SL g1058 ( 
.A(n_1009),
.Y(n_1058)
);

AOI22xp33_ASAP7_75t_SL g1059 ( 
.A1(n_979),
.A2(n_38),
.B1(n_42),
.B2(n_43),
.Y(n_1059)
);

INVx2_ASAP7_75t_L g1060 ( 
.A(n_917),
.Y(n_1060)
);

INVx2_ASAP7_75t_L g1061 ( 
.A(n_918),
.Y(n_1061)
);

AND2x2_ASAP7_75t_L g1062 ( 
.A(n_922),
.B(n_42),
.Y(n_1062)
);

OAI21x1_ASAP7_75t_L g1063 ( 
.A1(n_949),
.A2(n_124),
.B(n_221),
.Y(n_1063)
);

INVx1_ASAP7_75t_L g1064 ( 
.A(n_1009),
.Y(n_1064)
);

AOI22xp33_ASAP7_75t_L g1065 ( 
.A1(n_962),
.A2(n_43),
.B1(n_44),
.B2(n_45),
.Y(n_1065)
);

AOI21x1_ASAP7_75t_L g1066 ( 
.A1(n_1006),
.A2(n_222),
.B(n_127),
.Y(n_1066)
);

OA21x2_ASAP7_75t_L g1067 ( 
.A1(n_921),
.A2(n_980),
.B(n_970),
.Y(n_1067)
);

AND2x2_ASAP7_75t_L g1068 ( 
.A(n_941),
.B(n_45),
.Y(n_1068)
);

INVx2_ASAP7_75t_L g1069 ( 
.A(n_931),
.Y(n_1069)
);

AND2x2_ASAP7_75t_L g1070 ( 
.A(n_941),
.B(n_46),
.Y(n_1070)
);

AOI22xp33_ASAP7_75t_L g1071 ( 
.A1(n_977),
.A2(n_46),
.B1(n_49),
.B2(n_50),
.Y(n_1071)
);

INVx1_ASAP7_75t_L g1072 ( 
.A(n_987),
.Y(n_1072)
);

AOI22xp33_ASAP7_75t_L g1073 ( 
.A1(n_913),
.A2(n_51),
.B1(n_52),
.B2(n_53),
.Y(n_1073)
);

AND2x2_ASAP7_75t_L g1074 ( 
.A(n_941),
.B(n_914),
.Y(n_1074)
);

OAI21x1_ASAP7_75t_L g1075 ( 
.A1(n_927),
.A2(n_140),
.B(n_213),
.Y(n_1075)
);

BUFx6f_ASAP7_75t_L g1076 ( 
.A(n_925),
.Y(n_1076)
);

INVx1_ASAP7_75t_SL g1077 ( 
.A(n_945),
.Y(n_1077)
);

OAI22xp5_ASAP7_75t_L g1078 ( 
.A1(n_971),
.A2(n_53),
.B1(n_54),
.B2(n_55),
.Y(n_1078)
);

INVx2_ASAP7_75t_L g1079 ( 
.A(n_987),
.Y(n_1079)
);

OA21x2_ASAP7_75t_L g1080 ( 
.A1(n_921),
.A2(n_54),
.B(n_56),
.Y(n_1080)
);

OAI21x1_ASAP7_75t_SL g1081 ( 
.A1(n_927),
.A2(n_57),
.B(n_58),
.Y(n_1081)
);

OR2x2_ASAP7_75t_L g1082 ( 
.A(n_936),
.B(n_58),
.Y(n_1082)
);

BUFx3_ASAP7_75t_L g1083 ( 
.A(n_959),
.Y(n_1083)
);

NAND2xp5_ASAP7_75t_L g1084 ( 
.A(n_938),
.B(n_59),
.Y(n_1084)
);

INVx2_ASAP7_75t_L g1085 ( 
.A(n_988),
.Y(n_1085)
);

INVx1_ASAP7_75t_SL g1086 ( 
.A(n_972),
.Y(n_1086)
);

INVx2_ASAP7_75t_L g1087 ( 
.A(n_988),
.Y(n_1087)
);

HB1xp67_ASAP7_75t_L g1088 ( 
.A(n_961),
.Y(n_1088)
);

CKINVDCx11_ASAP7_75t_R g1089 ( 
.A(n_934),
.Y(n_1089)
);

BUFx10_ASAP7_75t_L g1090 ( 
.A(n_934),
.Y(n_1090)
);

INVx2_ASAP7_75t_SL g1091 ( 
.A(n_946),
.Y(n_1091)
);

INVx3_ASAP7_75t_L g1092 ( 
.A(n_1085),
.Y(n_1092)
);

INVx1_ASAP7_75t_L g1093 ( 
.A(n_1027),
.Y(n_1093)
);

BUFx2_ASAP7_75t_L g1094 ( 
.A(n_1045),
.Y(n_1094)
);

INVx1_ASAP7_75t_L g1095 ( 
.A(n_1027),
.Y(n_1095)
);

OR2x6_ASAP7_75t_L g1096 ( 
.A(n_1064),
.B(n_1007),
.Y(n_1096)
);

NAND2x1p5_ASAP7_75t_L g1097 ( 
.A(n_1023),
.B(n_988),
.Y(n_1097)
);

HB1xp67_ASAP7_75t_L g1098 ( 
.A(n_1045),
.Y(n_1098)
);

HB1xp67_ASAP7_75t_L g1099 ( 
.A(n_1052),
.Y(n_1099)
);

HB1xp67_ASAP7_75t_L g1100 ( 
.A(n_1052),
.Y(n_1100)
);

HB1xp67_ASAP7_75t_L g1101 ( 
.A(n_1015),
.Y(n_1101)
);

AND2x2_ASAP7_75t_L g1102 ( 
.A(n_1074),
.B(n_974),
.Y(n_1102)
);

INVxp67_ASAP7_75t_L g1103 ( 
.A(n_1088),
.Y(n_1103)
);

INVx2_ASAP7_75t_L g1104 ( 
.A(n_1013),
.Y(n_1104)
);

OA21x2_ASAP7_75t_L g1105 ( 
.A1(n_1026),
.A2(n_970),
.B(n_980),
.Y(n_1105)
);

OA21x2_ASAP7_75t_L g1106 ( 
.A1(n_1017),
.A2(n_936),
.B(n_990),
.Y(n_1106)
);

NAND2xp5_ASAP7_75t_L g1107 ( 
.A(n_1039),
.B(n_958),
.Y(n_1107)
);

BUFx12f_ASAP7_75t_L g1108 ( 
.A(n_1089),
.Y(n_1108)
);

HB1xp67_ASAP7_75t_L g1109 ( 
.A(n_1015),
.Y(n_1109)
);

INVx2_ASAP7_75t_L g1110 ( 
.A(n_1025),
.Y(n_1110)
);

BUFx2_ASAP7_75t_L g1111 ( 
.A(n_1085),
.Y(n_1111)
);

AND2x2_ASAP7_75t_L g1112 ( 
.A(n_1074),
.B(n_956),
.Y(n_1112)
);

INVx2_ASAP7_75t_L g1113 ( 
.A(n_1025),
.Y(n_1113)
);

INVx2_ASAP7_75t_L g1114 ( 
.A(n_1033),
.Y(n_1114)
);

OAI21x1_ASAP7_75t_L g1115 ( 
.A1(n_1017),
.A2(n_923),
.B(n_958),
.Y(n_1115)
);

HB1xp67_ASAP7_75t_L g1116 ( 
.A(n_1012),
.Y(n_1116)
);

INVx2_ASAP7_75t_L g1117 ( 
.A(n_1087),
.Y(n_1117)
);

CKINVDCx5p33_ASAP7_75t_R g1118 ( 
.A(n_1024),
.Y(n_1118)
);

INVx1_ASAP7_75t_L g1119 ( 
.A(n_1050),
.Y(n_1119)
);

INVx2_ASAP7_75t_L g1120 ( 
.A(n_1087),
.Y(n_1120)
);

INVx1_ASAP7_75t_L g1121 ( 
.A(n_1050),
.Y(n_1121)
);

NAND2xp5_ASAP7_75t_L g1122 ( 
.A(n_1039),
.B(n_937),
.Y(n_1122)
);

AO21x2_ASAP7_75t_L g1123 ( 
.A1(n_1044),
.A2(n_955),
.B(n_937),
.Y(n_1123)
);

INVx2_ASAP7_75t_L g1124 ( 
.A(n_1012),
.Y(n_1124)
);

AOI21x1_ASAP7_75t_L g1125 ( 
.A1(n_1044),
.A2(n_1057),
.B(n_1037),
.Y(n_1125)
);

INVx1_ASAP7_75t_L g1126 ( 
.A(n_1036),
.Y(n_1126)
);

NAND2x1_ASAP7_75t_L g1127 ( 
.A(n_1023),
.B(n_984),
.Y(n_1127)
);

OA21x2_ASAP7_75t_L g1128 ( 
.A1(n_1028),
.A2(n_944),
.B(n_923),
.Y(n_1128)
);

INVx1_ASAP7_75t_L g1129 ( 
.A(n_1036),
.Y(n_1129)
);

INVx2_ASAP7_75t_L g1130 ( 
.A(n_1022),
.Y(n_1130)
);

INVx1_ASAP7_75t_L g1131 ( 
.A(n_1043),
.Y(n_1131)
);

INVx5_ASAP7_75t_SL g1132 ( 
.A(n_1030),
.Y(n_1132)
);

INVx2_ASAP7_75t_L g1133 ( 
.A(n_1022),
.Y(n_1133)
);

HB1xp67_ASAP7_75t_L g1134 ( 
.A(n_1014),
.Y(n_1134)
);

INVx1_ASAP7_75t_L g1135 ( 
.A(n_1043),
.Y(n_1135)
);

INVx2_ASAP7_75t_L g1136 ( 
.A(n_1021),
.Y(n_1136)
);

CKINVDCx5p33_ASAP7_75t_R g1137 ( 
.A(n_1016),
.Y(n_1137)
);

INVx2_ASAP7_75t_L g1138 ( 
.A(n_1014),
.Y(n_1138)
);

INVx2_ASAP7_75t_L g1139 ( 
.A(n_1032),
.Y(n_1139)
);

INVx3_ASAP7_75t_L g1140 ( 
.A(n_1023),
.Y(n_1140)
);

INVx1_ASAP7_75t_L g1141 ( 
.A(n_1032),
.Y(n_1141)
);

BUFx6f_ASAP7_75t_L g1142 ( 
.A(n_1040),
.Y(n_1142)
);

INVx2_ASAP7_75t_L g1143 ( 
.A(n_1034),
.Y(n_1143)
);

INVx1_ASAP7_75t_L g1144 ( 
.A(n_1034),
.Y(n_1144)
);

INVx2_ASAP7_75t_L g1145 ( 
.A(n_1035),
.Y(n_1145)
);

AOI21x1_ASAP7_75t_L g1146 ( 
.A1(n_1057),
.A2(n_920),
.B(n_989),
.Y(n_1146)
);

NAND2xp5_ASAP7_75t_L g1147 ( 
.A(n_1067),
.B(n_966),
.Y(n_1147)
);

INVx1_ASAP7_75t_L g1148 ( 
.A(n_1035),
.Y(n_1148)
);

HB1xp67_ASAP7_75t_L g1149 ( 
.A(n_1047),
.Y(n_1149)
);

OR2x2_ASAP7_75t_L g1150 ( 
.A(n_1147),
.B(n_1067),
.Y(n_1150)
);

AND2x2_ASAP7_75t_L g1151 ( 
.A(n_1112),
.B(n_1067),
.Y(n_1151)
);

INVx1_ASAP7_75t_L g1152 ( 
.A(n_1139),
.Y(n_1152)
);

INVx1_ASAP7_75t_L g1153 ( 
.A(n_1139),
.Y(n_1153)
);

NAND2xp5_ASAP7_75t_L g1154 ( 
.A(n_1147),
.B(n_1067),
.Y(n_1154)
);

AND2x4_ASAP7_75t_L g1155 ( 
.A(n_1096),
.B(n_1058),
.Y(n_1155)
);

AND2x2_ASAP7_75t_L g1156 ( 
.A(n_1112),
.B(n_1068),
.Y(n_1156)
);

AND2x2_ASAP7_75t_L g1157 ( 
.A(n_1112),
.B(n_1070),
.Y(n_1157)
);

INVx1_ASAP7_75t_L g1158 ( 
.A(n_1139),
.Y(n_1158)
);

INVx2_ASAP7_75t_L g1159 ( 
.A(n_1104),
.Y(n_1159)
);

NAND2xp5_ASAP7_75t_L g1160 ( 
.A(n_1099),
.B(n_1047),
.Y(n_1160)
);

AND2x4_ASAP7_75t_L g1161 ( 
.A(n_1096),
.B(n_1058),
.Y(n_1161)
);

AND2x4_ASAP7_75t_L g1162 ( 
.A(n_1096),
.B(n_1058),
.Y(n_1162)
);

AND2x2_ASAP7_75t_L g1163 ( 
.A(n_1102),
.B(n_1080),
.Y(n_1163)
);

INVx1_ASAP7_75t_L g1164 ( 
.A(n_1139),
.Y(n_1164)
);

INVx2_ASAP7_75t_SL g1165 ( 
.A(n_1138),
.Y(n_1165)
);

INVx2_ASAP7_75t_L g1166 ( 
.A(n_1104),
.Y(n_1166)
);

BUFx6f_ASAP7_75t_L g1167 ( 
.A(n_1142),
.Y(n_1167)
);

AOI21xp5_ASAP7_75t_SL g1168 ( 
.A1(n_1142),
.A2(n_1040),
.B(n_1080),
.Y(n_1168)
);

OA21x2_ASAP7_75t_L g1169 ( 
.A1(n_1115),
.A2(n_1055),
.B(n_1054),
.Y(n_1169)
);

AND2x4_ASAP7_75t_L g1170 ( 
.A(n_1096),
.B(n_1058),
.Y(n_1170)
);

INVx2_ASAP7_75t_L g1171 ( 
.A(n_1104),
.Y(n_1171)
);

AND2x2_ASAP7_75t_L g1172 ( 
.A(n_1102),
.B(n_1080),
.Y(n_1172)
);

INVx2_ASAP7_75t_L g1173 ( 
.A(n_1110),
.Y(n_1173)
);

OAI21xp5_ASAP7_75t_L g1174 ( 
.A1(n_1105),
.A2(n_1078),
.B(n_1031),
.Y(n_1174)
);

INVx1_ASAP7_75t_L g1175 ( 
.A(n_1143),
.Y(n_1175)
);

INVx4_ASAP7_75t_R g1176 ( 
.A(n_1132),
.Y(n_1176)
);

INVx1_ASAP7_75t_L g1177 ( 
.A(n_1143),
.Y(n_1177)
);

INVx1_ASAP7_75t_L g1178 ( 
.A(n_1143),
.Y(n_1178)
);

NAND2xp5_ASAP7_75t_L g1179 ( 
.A(n_1099),
.B(n_1049),
.Y(n_1179)
);

INVx1_ASAP7_75t_L g1180 ( 
.A(n_1145),
.Y(n_1180)
);

INVx1_ASAP7_75t_L g1181 ( 
.A(n_1145),
.Y(n_1181)
);

NAND2xp5_ASAP7_75t_L g1182 ( 
.A(n_1100),
.B(n_1049),
.Y(n_1182)
);

INVx1_ASAP7_75t_L g1183 ( 
.A(n_1145),
.Y(n_1183)
);

AND2x2_ASAP7_75t_L g1184 ( 
.A(n_1102),
.B(n_1080),
.Y(n_1184)
);

BUFx2_ASAP7_75t_L g1185 ( 
.A(n_1094),
.Y(n_1185)
);

AND2x2_ASAP7_75t_L g1186 ( 
.A(n_1119),
.B(n_1019),
.Y(n_1186)
);

INVx8_ASAP7_75t_L g1187 ( 
.A(n_1108),
.Y(n_1187)
);

AOI22xp33_ASAP7_75t_SL g1188 ( 
.A1(n_1105),
.A2(n_1062),
.B1(n_1081),
.B2(n_1064),
.Y(n_1188)
);

HB1xp67_ASAP7_75t_L g1189 ( 
.A(n_1103),
.Y(n_1189)
);

AND2x2_ASAP7_75t_L g1190 ( 
.A(n_1119),
.B(n_1053),
.Y(n_1190)
);

AND2x2_ASAP7_75t_L g1191 ( 
.A(n_1121),
.B(n_1062),
.Y(n_1191)
);

NOR2xp33_ASAP7_75t_L g1192 ( 
.A(n_1137),
.B(n_1056),
.Y(n_1192)
);

INVx1_ASAP7_75t_L g1193 ( 
.A(n_1093),
.Y(n_1193)
);

NAND2xp5_ASAP7_75t_L g1194 ( 
.A(n_1189),
.B(n_1103),
.Y(n_1194)
);

NAND2xp5_ASAP7_75t_L g1195 ( 
.A(n_1186),
.B(n_1100),
.Y(n_1195)
);

NAND2xp5_ASAP7_75t_L g1196 ( 
.A(n_1186),
.B(n_1107),
.Y(n_1196)
);

AND2x2_ASAP7_75t_L g1197 ( 
.A(n_1151),
.B(n_1094),
.Y(n_1197)
);

AOI21x1_ASAP7_75t_L g1198 ( 
.A1(n_1154),
.A2(n_1125),
.B(n_1146),
.Y(n_1198)
);

NOR2xp33_ASAP7_75t_R g1199 ( 
.A(n_1187),
.B(n_1118),
.Y(n_1199)
);

AND2x2_ASAP7_75t_L g1200 ( 
.A(n_1151),
.B(n_1094),
.Y(n_1200)
);

AND2x2_ASAP7_75t_L g1201 ( 
.A(n_1156),
.B(n_1149),
.Y(n_1201)
);

OAI221xp5_ASAP7_75t_L g1202 ( 
.A1(n_1174),
.A2(n_1059),
.B1(n_1084),
.B2(n_1071),
.C(n_1107),
.Y(n_1202)
);

NAND2xp5_ASAP7_75t_L g1203 ( 
.A(n_1190),
.B(n_1149),
.Y(n_1203)
);

INVxp67_ASAP7_75t_L g1204 ( 
.A(n_1190),
.Y(n_1204)
);

AND2x2_ASAP7_75t_L g1205 ( 
.A(n_1156),
.B(n_1098),
.Y(n_1205)
);

NAND3xp33_ASAP7_75t_L g1206 ( 
.A(n_1188),
.B(n_1105),
.C(n_1082),
.Y(n_1206)
);

NAND2xp5_ASAP7_75t_SL g1207 ( 
.A(n_1155),
.B(n_1132),
.Y(n_1207)
);

NAND2xp5_ASAP7_75t_SL g1208 ( 
.A(n_1155),
.B(n_1132),
.Y(n_1208)
);

AND2x2_ASAP7_75t_L g1209 ( 
.A(n_1157),
.B(n_1098),
.Y(n_1209)
);

AND2x2_ASAP7_75t_L g1210 ( 
.A(n_1157),
.B(n_1134),
.Y(n_1210)
);

AND2x2_ASAP7_75t_L g1211 ( 
.A(n_1163),
.B(n_1134),
.Y(n_1211)
);

AND2x2_ASAP7_75t_L g1212 ( 
.A(n_1163),
.B(n_1101),
.Y(n_1212)
);

NAND2xp5_ASAP7_75t_L g1213 ( 
.A(n_1191),
.B(n_1101),
.Y(n_1213)
);

AND2x2_ASAP7_75t_L g1214 ( 
.A(n_1172),
.B(n_1109),
.Y(n_1214)
);

AND2x2_ASAP7_75t_L g1215 ( 
.A(n_1172),
.B(n_1109),
.Y(n_1215)
);

NAND3xp33_ASAP7_75t_L g1216 ( 
.A(n_1154),
.B(n_1105),
.C(n_1082),
.Y(n_1216)
);

NAND2xp5_ASAP7_75t_L g1217 ( 
.A(n_1191),
.B(n_1116),
.Y(n_1217)
);

AND2x2_ASAP7_75t_L g1218 ( 
.A(n_1184),
.B(n_1116),
.Y(n_1218)
);

NAND2xp5_ASAP7_75t_L g1219 ( 
.A(n_1150),
.B(n_1122),
.Y(n_1219)
);

AND2x2_ASAP7_75t_L g1220 ( 
.A(n_1184),
.B(n_1121),
.Y(n_1220)
);

NAND3xp33_ASAP7_75t_L g1221 ( 
.A(n_1168),
.B(n_1011),
.C(n_1073),
.Y(n_1221)
);

NAND4xp25_ASAP7_75t_L g1222 ( 
.A(n_1185),
.B(n_1065),
.C(n_1086),
.D(n_995),
.Y(n_1222)
);

OAI221xp5_ASAP7_75t_L g1223 ( 
.A1(n_1168),
.A2(n_1122),
.B1(n_1029),
.B2(n_950),
.C(n_1128),
.Y(n_1223)
);

AND2x2_ASAP7_75t_L g1224 ( 
.A(n_1165),
.B(n_1126),
.Y(n_1224)
);

NAND4xp25_ASAP7_75t_L g1225 ( 
.A(n_1185),
.B(n_1010),
.C(n_954),
.D(n_947),
.Y(n_1225)
);

NOR2xp33_ASAP7_75t_L g1226 ( 
.A(n_1192),
.B(n_1108),
.Y(n_1226)
);

NAND2xp5_ASAP7_75t_L g1227 ( 
.A(n_1150),
.B(n_1126),
.Y(n_1227)
);

NAND2xp5_ASAP7_75t_L g1228 ( 
.A(n_1160),
.B(n_1129),
.Y(n_1228)
);

AND2x2_ASAP7_75t_L g1229 ( 
.A(n_1165),
.B(n_1129),
.Y(n_1229)
);

NAND2xp5_ASAP7_75t_L g1230 ( 
.A(n_1179),
.B(n_1131),
.Y(n_1230)
);

INVx2_ASAP7_75t_L g1231 ( 
.A(n_1159),
.Y(n_1231)
);

NAND2xp5_ASAP7_75t_SL g1232 ( 
.A(n_1155),
.B(n_1161),
.Y(n_1232)
);

NAND2xp5_ASAP7_75t_L g1233 ( 
.A(n_1179),
.B(n_1131),
.Y(n_1233)
);

AOI22xp33_ASAP7_75t_L g1234 ( 
.A1(n_1161),
.A2(n_1128),
.B1(n_1123),
.B2(n_1055),
.Y(n_1234)
);

NAND3xp33_ASAP7_75t_L g1235 ( 
.A(n_1182),
.B(n_1106),
.C(n_985),
.Y(n_1235)
);

OAI22xp5_ASAP7_75t_L g1236 ( 
.A1(n_1187),
.A2(n_1132),
.B1(n_1040),
.B2(n_989),
.Y(n_1236)
);

NAND2xp5_ASAP7_75t_L g1237 ( 
.A(n_1182),
.B(n_1135),
.Y(n_1237)
);

AND2x2_ASAP7_75t_L g1238 ( 
.A(n_1152),
.B(n_1153),
.Y(n_1238)
);

NAND2xp5_ASAP7_75t_L g1239 ( 
.A(n_1193),
.B(n_1141),
.Y(n_1239)
);

NAND2xp5_ASAP7_75t_L g1240 ( 
.A(n_1193),
.B(n_1141),
.Y(n_1240)
);

INVx1_ASAP7_75t_L g1241 ( 
.A(n_1152),
.Y(n_1241)
);

INVx1_ASAP7_75t_L g1242 ( 
.A(n_1241),
.Y(n_1242)
);

INVx1_ASAP7_75t_L g1243 ( 
.A(n_1241),
.Y(n_1243)
);

INVx1_ASAP7_75t_L g1244 ( 
.A(n_1238),
.Y(n_1244)
);

INVx1_ASAP7_75t_L g1245 ( 
.A(n_1238),
.Y(n_1245)
);

HB1xp67_ASAP7_75t_L g1246 ( 
.A(n_1212),
.Y(n_1246)
);

INVx3_ASAP7_75t_L g1247 ( 
.A(n_1198),
.Y(n_1247)
);

NAND2xp5_ASAP7_75t_L g1248 ( 
.A(n_1227),
.B(n_1153),
.Y(n_1248)
);

AND2x4_ASAP7_75t_L g1249 ( 
.A(n_1232),
.B(n_1161),
.Y(n_1249)
);

BUFx2_ASAP7_75t_L g1250 ( 
.A(n_1211),
.Y(n_1250)
);

NAND2xp5_ASAP7_75t_L g1251 ( 
.A(n_1219),
.B(n_1158),
.Y(n_1251)
);

INVx2_ASAP7_75t_L g1252 ( 
.A(n_1231),
.Y(n_1252)
);

AND2x2_ASAP7_75t_L g1253 ( 
.A(n_1197),
.B(n_1158),
.Y(n_1253)
);

NAND2xp5_ASAP7_75t_L g1254 ( 
.A(n_1216),
.B(n_1164),
.Y(n_1254)
);

HB1xp67_ASAP7_75t_L g1255 ( 
.A(n_1212),
.Y(n_1255)
);

AND2x2_ASAP7_75t_L g1256 ( 
.A(n_1197),
.B(n_1164),
.Y(n_1256)
);

NOR2x1_ASAP7_75t_L g1257 ( 
.A(n_1206),
.B(n_1161),
.Y(n_1257)
);

INVx2_ASAP7_75t_L g1258 ( 
.A(n_1231),
.Y(n_1258)
);

AND2x4_ASAP7_75t_SL g1259 ( 
.A(n_1201),
.B(n_1162),
.Y(n_1259)
);

OR2x2_ASAP7_75t_L g1260 ( 
.A(n_1203),
.B(n_1175),
.Y(n_1260)
);

INVx2_ASAP7_75t_SL g1261 ( 
.A(n_1224),
.Y(n_1261)
);

NAND2xp5_ASAP7_75t_L g1262 ( 
.A(n_1216),
.B(n_1175),
.Y(n_1262)
);

INVx1_ASAP7_75t_L g1263 ( 
.A(n_1224),
.Y(n_1263)
);

AND2x2_ASAP7_75t_L g1264 ( 
.A(n_1200),
.B(n_1177),
.Y(n_1264)
);

AND2x4_ASAP7_75t_SL g1265 ( 
.A(n_1201),
.B(n_1162),
.Y(n_1265)
);

INVxp67_ASAP7_75t_L g1266 ( 
.A(n_1206),
.Y(n_1266)
);

INVxp67_ASAP7_75t_SL g1267 ( 
.A(n_1198),
.Y(n_1267)
);

INVx1_ASAP7_75t_L g1268 ( 
.A(n_1229),
.Y(n_1268)
);

AND2x2_ASAP7_75t_L g1269 ( 
.A(n_1200),
.B(n_1177),
.Y(n_1269)
);

INVx1_ASAP7_75t_L g1270 ( 
.A(n_1229),
.Y(n_1270)
);

NAND2xp5_ASAP7_75t_L g1271 ( 
.A(n_1220),
.B(n_1228),
.Y(n_1271)
);

INVx3_ASAP7_75t_L g1272 ( 
.A(n_1220),
.Y(n_1272)
);

AND2x2_ASAP7_75t_L g1273 ( 
.A(n_1211),
.B(n_1178),
.Y(n_1273)
);

INVx2_ASAP7_75t_L g1274 ( 
.A(n_1214),
.Y(n_1274)
);

AND2x4_ASAP7_75t_L g1275 ( 
.A(n_1257),
.B(n_1207),
.Y(n_1275)
);

AND2x2_ASAP7_75t_L g1276 ( 
.A(n_1259),
.B(n_1214),
.Y(n_1276)
);

OR2x2_ASAP7_75t_L g1277 ( 
.A(n_1266),
.B(n_1195),
.Y(n_1277)
);

AND2x2_ASAP7_75t_L g1278 ( 
.A(n_1259),
.B(n_1215),
.Y(n_1278)
);

NAND2xp5_ASAP7_75t_SL g1279 ( 
.A(n_1257),
.B(n_1266),
.Y(n_1279)
);

INVx1_ASAP7_75t_L g1280 ( 
.A(n_1242),
.Y(n_1280)
);

AND2x4_ASAP7_75t_L g1281 ( 
.A(n_1249),
.B(n_1208),
.Y(n_1281)
);

INVx1_ASAP7_75t_L g1282 ( 
.A(n_1242),
.Y(n_1282)
);

AND2x2_ASAP7_75t_L g1283 ( 
.A(n_1265),
.B(n_1218),
.Y(n_1283)
);

INVx1_ASAP7_75t_L g1284 ( 
.A(n_1243),
.Y(n_1284)
);

AND2x2_ASAP7_75t_L g1285 ( 
.A(n_1265),
.B(n_1218),
.Y(n_1285)
);

OAI33xp33_ASAP7_75t_L g1286 ( 
.A1(n_1254),
.A2(n_1194),
.A3(n_1225),
.B1(n_1233),
.B2(n_1237),
.B3(n_1230),
.Y(n_1286)
);

AND2x2_ASAP7_75t_L g1287 ( 
.A(n_1265),
.B(n_1210),
.Y(n_1287)
);

NAND2xp5_ASAP7_75t_L g1288 ( 
.A(n_1271),
.B(n_1196),
.Y(n_1288)
);

INVx2_ASAP7_75t_L g1289 ( 
.A(n_1252),
.Y(n_1289)
);

INVx1_ASAP7_75t_L g1290 ( 
.A(n_1243),
.Y(n_1290)
);

INVx1_ASAP7_75t_L g1291 ( 
.A(n_1244),
.Y(n_1291)
);

NOR2xp33_ASAP7_75t_SL g1292 ( 
.A(n_1249),
.B(n_1108),
.Y(n_1292)
);

INVx1_ASAP7_75t_L g1293 ( 
.A(n_1244),
.Y(n_1293)
);

OR2x2_ASAP7_75t_L g1294 ( 
.A(n_1271),
.B(n_1260),
.Y(n_1294)
);

INVxp67_ASAP7_75t_SL g1295 ( 
.A(n_1254),
.Y(n_1295)
);

INVx1_ASAP7_75t_L g1296 ( 
.A(n_1245),
.Y(n_1296)
);

AND2x2_ASAP7_75t_L g1297 ( 
.A(n_1250),
.B(n_1272),
.Y(n_1297)
);

INVx2_ASAP7_75t_SL g1298 ( 
.A(n_1249),
.Y(n_1298)
);

INVx1_ASAP7_75t_L g1299 ( 
.A(n_1245),
.Y(n_1299)
);

INVxp67_ASAP7_75t_L g1300 ( 
.A(n_1262),
.Y(n_1300)
);

NAND2xp5_ASAP7_75t_L g1301 ( 
.A(n_1262),
.B(n_1205),
.Y(n_1301)
);

INVx1_ASAP7_75t_L g1302 ( 
.A(n_1260),
.Y(n_1302)
);

AND2x2_ASAP7_75t_L g1303 ( 
.A(n_1250),
.B(n_1210),
.Y(n_1303)
);

INVx1_ASAP7_75t_L g1304 ( 
.A(n_1248),
.Y(n_1304)
);

NOR2xp67_ASAP7_75t_L g1305 ( 
.A(n_1272),
.B(n_1108),
.Y(n_1305)
);

HB1xp67_ASAP7_75t_L g1306 ( 
.A(n_1300),
.Y(n_1306)
);

INVx1_ASAP7_75t_L g1307 ( 
.A(n_1280),
.Y(n_1307)
);

INVx2_ASAP7_75t_L g1308 ( 
.A(n_1289),
.Y(n_1308)
);

INVx1_ASAP7_75t_L g1309 ( 
.A(n_1280),
.Y(n_1309)
);

NOR2xp33_ASAP7_75t_L g1310 ( 
.A(n_1286),
.B(n_1226),
.Y(n_1310)
);

AND2x2_ASAP7_75t_L g1311 ( 
.A(n_1297),
.B(n_1272),
.Y(n_1311)
);

INVx1_ASAP7_75t_L g1312 ( 
.A(n_1282),
.Y(n_1312)
);

OR2x2_ASAP7_75t_L g1313 ( 
.A(n_1294),
.B(n_1277),
.Y(n_1313)
);

AND2x2_ASAP7_75t_L g1314 ( 
.A(n_1297),
.B(n_1272),
.Y(n_1314)
);

AND2x4_ASAP7_75t_L g1315 ( 
.A(n_1298),
.B(n_1249),
.Y(n_1315)
);

INVx1_ASAP7_75t_L g1316 ( 
.A(n_1282),
.Y(n_1316)
);

HB1xp67_ASAP7_75t_L g1317 ( 
.A(n_1277),
.Y(n_1317)
);

INVxp67_ASAP7_75t_SL g1318 ( 
.A(n_1279),
.Y(n_1318)
);

INVx1_ASAP7_75t_L g1319 ( 
.A(n_1284),
.Y(n_1319)
);

HB1xp67_ASAP7_75t_L g1320 ( 
.A(n_1302),
.Y(n_1320)
);

INVx1_ASAP7_75t_L g1321 ( 
.A(n_1284),
.Y(n_1321)
);

INVx1_ASAP7_75t_L g1322 ( 
.A(n_1290),
.Y(n_1322)
);

INVx2_ASAP7_75t_L g1323 ( 
.A(n_1289),
.Y(n_1323)
);

NOR2xp33_ASAP7_75t_SL g1324 ( 
.A(n_1292),
.B(n_1187),
.Y(n_1324)
);

INVx2_ASAP7_75t_L g1325 ( 
.A(n_1290),
.Y(n_1325)
);

INVxp67_ASAP7_75t_L g1326 ( 
.A(n_1295),
.Y(n_1326)
);

OR2x2_ASAP7_75t_L g1327 ( 
.A(n_1294),
.B(n_1251),
.Y(n_1327)
);

NAND2xp5_ASAP7_75t_L g1328 ( 
.A(n_1288),
.B(n_1261),
.Y(n_1328)
);

INVx1_ASAP7_75t_L g1329 ( 
.A(n_1291),
.Y(n_1329)
);

NAND2xp5_ASAP7_75t_L g1330 ( 
.A(n_1304),
.B(n_1303),
.Y(n_1330)
);

INVx1_ASAP7_75t_L g1331 ( 
.A(n_1291),
.Y(n_1331)
);

AND2x2_ASAP7_75t_L g1332 ( 
.A(n_1303),
.B(n_1261),
.Y(n_1332)
);

INVx1_ASAP7_75t_L g1333 ( 
.A(n_1293),
.Y(n_1333)
);

INVx1_ASAP7_75t_L g1334 ( 
.A(n_1293),
.Y(n_1334)
);

AND2x2_ASAP7_75t_L g1335 ( 
.A(n_1275),
.B(n_1261),
.Y(n_1335)
);

AND2x2_ASAP7_75t_L g1336 ( 
.A(n_1275),
.B(n_1246),
.Y(n_1336)
);

INVx1_ASAP7_75t_L g1337 ( 
.A(n_1296),
.Y(n_1337)
);

AND2x2_ASAP7_75t_L g1338 ( 
.A(n_1275),
.B(n_1255),
.Y(n_1338)
);

OAI21xp33_ASAP7_75t_L g1339 ( 
.A1(n_1318),
.A2(n_1304),
.B(n_1298),
.Y(n_1339)
);

INVx1_ASAP7_75t_SL g1340 ( 
.A(n_1317),
.Y(n_1340)
);

OR2x2_ASAP7_75t_L g1341 ( 
.A(n_1313),
.B(n_1330),
.Y(n_1341)
);

INVx1_ASAP7_75t_L g1342 ( 
.A(n_1320),
.Y(n_1342)
);

NOR2xp33_ASAP7_75t_L g1343 ( 
.A(n_1310),
.B(n_1137),
.Y(n_1343)
);

NOR2xp33_ASAP7_75t_L g1344 ( 
.A(n_1306),
.B(n_1281),
.Y(n_1344)
);

INVx1_ASAP7_75t_L g1345 ( 
.A(n_1307),
.Y(n_1345)
);

INVxp67_ASAP7_75t_L g1346 ( 
.A(n_1309),
.Y(n_1346)
);

INVx3_ASAP7_75t_L g1347 ( 
.A(n_1315),
.Y(n_1347)
);

INVx1_ASAP7_75t_L g1348 ( 
.A(n_1309),
.Y(n_1348)
);

BUFx3_ASAP7_75t_L g1349 ( 
.A(n_1315),
.Y(n_1349)
);

INVx1_ASAP7_75t_L g1350 ( 
.A(n_1312),
.Y(n_1350)
);

INVx1_ASAP7_75t_L g1351 ( 
.A(n_1312),
.Y(n_1351)
);

AND2x2_ASAP7_75t_L g1352 ( 
.A(n_1336),
.B(n_1287),
.Y(n_1352)
);

AOI22xp5_ASAP7_75t_L g1353 ( 
.A1(n_1326),
.A2(n_1222),
.B1(n_1221),
.B2(n_1223),
.Y(n_1353)
);

NOR2xp33_ASAP7_75t_L g1354 ( 
.A(n_1327),
.B(n_1336),
.Y(n_1354)
);

AND2x2_ASAP7_75t_L g1355 ( 
.A(n_1338),
.B(n_1332),
.Y(n_1355)
);

AOI22xp33_ASAP7_75t_L g1356 ( 
.A1(n_1308),
.A2(n_1222),
.B1(n_1202),
.B2(n_1221),
.Y(n_1356)
);

NAND2xp5_ASAP7_75t_L g1357 ( 
.A(n_1327),
.B(n_1301),
.Y(n_1357)
);

CKINVDCx5p33_ASAP7_75t_R g1358 ( 
.A(n_1315),
.Y(n_1358)
);

INVx3_ASAP7_75t_L g1359 ( 
.A(n_1335),
.Y(n_1359)
);

OR2x2_ASAP7_75t_L g1360 ( 
.A(n_1328),
.B(n_1316),
.Y(n_1360)
);

AND2x2_ASAP7_75t_L g1361 ( 
.A(n_1338),
.B(n_1287),
.Y(n_1361)
);

NOR2x1_ASAP7_75t_L g1362 ( 
.A(n_1335),
.B(n_1305),
.Y(n_1362)
);

AND2x2_ASAP7_75t_L g1363 ( 
.A(n_1311),
.B(n_1314),
.Y(n_1363)
);

OR2x2_ASAP7_75t_L g1364 ( 
.A(n_1316),
.B(n_1296),
.Y(n_1364)
);

OR2x2_ASAP7_75t_L g1365 ( 
.A(n_1319),
.B(n_1299),
.Y(n_1365)
);

AOI22xp5_ASAP7_75t_L g1366 ( 
.A1(n_1356),
.A2(n_1324),
.B1(n_1323),
.B2(n_1308),
.Y(n_1366)
);

AOI21xp33_ASAP7_75t_L g1367 ( 
.A1(n_1343),
.A2(n_1356),
.B(n_1340),
.Y(n_1367)
);

AOI221xp5_ASAP7_75t_SL g1368 ( 
.A1(n_1339),
.A2(n_1311),
.B1(n_1314),
.B2(n_1321),
.C(n_1319),
.Y(n_1368)
);

INVx1_ASAP7_75t_L g1369 ( 
.A(n_1345),
.Y(n_1369)
);

INVx1_ASAP7_75t_L g1370 ( 
.A(n_1348),
.Y(n_1370)
);

INVx2_ASAP7_75t_L g1371 ( 
.A(n_1349),
.Y(n_1371)
);

INVx1_ASAP7_75t_L g1372 ( 
.A(n_1350),
.Y(n_1372)
);

INVx1_ASAP7_75t_L g1373 ( 
.A(n_1351),
.Y(n_1373)
);

NOR2xp33_ASAP7_75t_R g1374 ( 
.A(n_1358),
.B(n_1187),
.Y(n_1374)
);

INVx1_ASAP7_75t_L g1375 ( 
.A(n_1346),
.Y(n_1375)
);

INVx1_ASAP7_75t_L g1376 ( 
.A(n_1346),
.Y(n_1376)
);

NOR3xp33_ASAP7_75t_L g1377 ( 
.A(n_1343),
.B(n_1267),
.C(n_1247),
.Y(n_1377)
);

INVx1_ASAP7_75t_SL g1378 ( 
.A(n_1349),
.Y(n_1378)
);

OAI21xp5_ASAP7_75t_L g1379 ( 
.A1(n_1353),
.A2(n_1322),
.B(n_1321),
.Y(n_1379)
);

A2O1A1Ixp33_ASAP7_75t_L g1380 ( 
.A1(n_1344),
.A2(n_1235),
.B(n_1325),
.C(n_1247),
.Y(n_1380)
);

INVx1_ASAP7_75t_L g1381 ( 
.A(n_1342),
.Y(n_1381)
);

OAI322xp33_ASAP7_75t_L g1382 ( 
.A1(n_1354),
.A2(n_1322),
.A3(n_1334),
.B1(n_1333),
.B2(n_1331),
.C1(n_1329),
.C2(n_1337),
.Y(n_1382)
);

HB1xp67_ASAP7_75t_L g1383 ( 
.A(n_1347),
.Y(n_1383)
);

INVx1_ASAP7_75t_L g1384 ( 
.A(n_1364),
.Y(n_1384)
);

AND2x2_ASAP7_75t_L g1385 ( 
.A(n_1355),
.B(n_1276),
.Y(n_1385)
);

AND2x2_ASAP7_75t_L g1386 ( 
.A(n_1352),
.B(n_1276),
.Y(n_1386)
);

O2A1O1Ixp33_ASAP7_75t_L g1387 ( 
.A1(n_1344),
.A2(n_1081),
.B(n_1247),
.C(n_1333),
.Y(n_1387)
);

OAI21xp33_ASAP7_75t_L g1388 ( 
.A1(n_1357),
.A2(n_1337),
.B(n_1334),
.Y(n_1388)
);

AOI322xp5_ASAP7_75t_L g1389 ( 
.A1(n_1362),
.A2(n_1323),
.A3(n_1308),
.B1(n_1234),
.B2(n_1247),
.C1(n_1205),
.C2(n_1209),
.Y(n_1389)
);

NAND2xp5_ASAP7_75t_SL g1390 ( 
.A(n_1347),
.B(n_1199),
.Y(n_1390)
);

INVxp67_ASAP7_75t_SL g1391 ( 
.A(n_1359),
.Y(n_1391)
);

INVx2_ASAP7_75t_SL g1392 ( 
.A(n_1359),
.Y(n_1392)
);

INVx1_ASAP7_75t_L g1393 ( 
.A(n_1365),
.Y(n_1393)
);

INVxp67_ASAP7_75t_L g1394 ( 
.A(n_1360),
.Y(n_1394)
);

AO21x1_ASAP7_75t_L g1395 ( 
.A1(n_1341),
.A2(n_1323),
.B(n_1299),
.Y(n_1395)
);

AND2x2_ASAP7_75t_L g1396 ( 
.A(n_1385),
.B(n_1386),
.Y(n_1396)
);

NAND2xp5_ASAP7_75t_L g1397 ( 
.A(n_1391),
.B(n_1363),
.Y(n_1397)
);

AOI22xp33_ASAP7_75t_L g1398 ( 
.A1(n_1379),
.A2(n_1367),
.B1(n_1395),
.B2(n_1377),
.Y(n_1398)
);

INVx1_ASAP7_75t_L g1399 ( 
.A(n_1383),
.Y(n_1399)
);

AOI22xp33_ASAP7_75t_R g1400 ( 
.A1(n_1394),
.A2(n_982),
.B1(n_1077),
.B2(n_1252),
.Y(n_1400)
);

NAND2xp5_ASAP7_75t_L g1401 ( 
.A(n_1391),
.B(n_1361),
.Y(n_1401)
);

INVx1_ASAP7_75t_L g1402 ( 
.A(n_1369),
.Y(n_1402)
);

AND2x2_ASAP7_75t_L g1403 ( 
.A(n_1378),
.B(n_1278),
.Y(n_1403)
);

INVx2_ASAP7_75t_L g1404 ( 
.A(n_1371),
.Y(n_1404)
);

INVx2_ASAP7_75t_L g1405 ( 
.A(n_1392),
.Y(n_1405)
);

NOR2xp33_ASAP7_75t_L g1406 ( 
.A(n_1382),
.B(n_1187),
.Y(n_1406)
);

NAND2xp5_ASAP7_75t_L g1407 ( 
.A(n_1384),
.B(n_1263),
.Y(n_1407)
);

INVx1_ASAP7_75t_L g1408 ( 
.A(n_1370),
.Y(n_1408)
);

NAND2xp5_ASAP7_75t_L g1409 ( 
.A(n_1393),
.B(n_1268),
.Y(n_1409)
);

OR2x2_ASAP7_75t_L g1410 ( 
.A(n_1381),
.B(n_1375),
.Y(n_1410)
);

INVx1_ASAP7_75t_L g1411 ( 
.A(n_1372),
.Y(n_1411)
);

INVx1_ASAP7_75t_L g1412 ( 
.A(n_1373),
.Y(n_1412)
);

INVx1_ASAP7_75t_L g1413 ( 
.A(n_1376),
.Y(n_1413)
);

INVxp67_ASAP7_75t_L g1414 ( 
.A(n_1366),
.Y(n_1414)
);

NAND2xp5_ASAP7_75t_L g1415 ( 
.A(n_1388),
.B(n_1268),
.Y(n_1415)
);

AOI221xp5_ASAP7_75t_L g1416 ( 
.A1(n_1380),
.A2(n_1251),
.B1(n_1248),
.B2(n_1236),
.C(n_973),
.Y(n_1416)
);

NAND2xp5_ASAP7_75t_L g1417 ( 
.A(n_1368),
.B(n_1270),
.Y(n_1417)
);

INVx1_ASAP7_75t_L g1418 ( 
.A(n_1387),
.Y(n_1418)
);

OR2x2_ASAP7_75t_L g1419 ( 
.A(n_1390),
.B(n_1274),
.Y(n_1419)
);

NOR3xp33_ASAP7_75t_SL g1420 ( 
.A(n_1387),
.B(n_1083),
.C(n_1213),
.Y(n_1420)
);

NOR2x1_ASAP7_75t_L g1421 ( 
.A(n_1374),
.B(n_1083),
.Y(n_1421)
);

INVx1_ASAP7_75t_L g1422 ( 
.A(n_1389),
.Y(n_1422)
);

NAND2x1_ASAP7_75t_SL g1423 ( 
.A(n_1383),
.B(n_1283),
.Y(n_1423)
);

NAND2xp5_ASAP7_75t_L g1424 ( 
.A(n_1391),
.B(n_1285),
.Y(n_1424)
);

OAI211xp5_ASAP7_75t_SL g1425 ( 
.A1(n_1398),
.A2(n_1274),
.B(n_1204),
.C(n_1217),
.Y(n_1425)
);

O2A1O1Ixp33_ASAP7_75t_L g1426 ( 
.A1(n_1422),
.A2(n_989),
.B(n_951),
.C(n_944),
.Y(n_1426)
);

AOI222xp33_ASAP7_75t_L g1427 ( 
.A1(n_1414),
.A2(n_981),
.B1(n_1252),
.B2(n_1258),
.C1(n_1063),
.C2(n_1046),
.Y(n_1427)
);

A2O1A1Ixp33_ASAP7_75t_L g1428 ( 
.A1(n_1406),
.A2(n_1063),
.B(n_1046),
.C(n_1115),
.Y(n_1428)
);

NAND4xp25_ASAP7_75t_SL g1429 ( 
.A(n_1401),
.B(n_1397),
.C(n_1396),
.D(n_1424),
.Y(n_1429)
);

AOI22xp5_ASAP7_75t_L g1430 ( 
.A1(n_1416),
.A2(n_1142),
.B1(n_1258),
.B2(n_1162),
.Y(n_1430)
);

NAND3xp33_ASAP7_75t_SL g1431 ( 
.A(n_1406),
.B(n_1038),
.C(n_967),
.Y(n_1431)
);

OAI322xp33_ASAP7_75t_L g1432 ( 
.A1(n_1418),
.A2(n_1239),
.A3(n_1240),
.B1(n_1148),
.B2(n_1144),
.C1(n_1273),
.C2(n_1095),
.Y(n_1432)
);

OAI211xp5_ASAP7_75t_L g1433 ( 
.A1(n_1423),
.A2(n_1405),
.B(n_1410),
.C(n_1413),
.Y(n_1433)
);

NAND4xp25_ASAP7_75t_L g1434 ( 
.A(n_1405),
.B(n_1269),
.C(n_1264),
.D(n_1256),
.Y(n_1434)
);

NAND4xp25_ASAP7_75t_L g1435 ( 
.A(n_1399),
.B(n_1269),
.C(n_1264),
.D(n_1256),
.Y(n_1435)
);

NAND3xp33_ASAP7_75t_SL g1436 ( 
.A(n_1420),
.B(n_1038),
.C(n_1018),
.Y(n_1436)
);

AOI21xp5_ASAP7_75t_L g1437 ( 
.A1(n_1421),
.A2(n_1417),
.B(n_1403),
.Y(n_1437)
);

AOI22xp5_ASAP7_75t_L g1438 ( 
.A1(n_1404),
.A2(n_1258),
.B1(n_1170),
.B2(n_1167),
.Y(n_1438)
);

NAND4xp25_ASAP7_75t_L g1439 ( 
.A(n_1402),
.B(n_1253),
.C(n_1140),
.D(n_1038),
.Y(n_1439)
);

AOI221xp5_ASAP7_75t_L g1440 ( 
.A1(n_1408),
.A2(n_1144),
.B1(n_1148),
.B2(n_1253),
.C(n_1095),
.Y(n_1440)
);

NAND3xp33_ASAP7_75t_L g1441 ( 
.A(n_1411),
.B(n_1076),
.C(n_1020),
.Y(n_1441)
);

INVx1_ASAP7_75t_L g1442 ( 
.A(n_1412),
.Y(n_1442)
);

NAND2xp5_ASAP7_75t_L g1443 ( 
.A(n_1407),
.B(n_60),
.Y(n_1443)
);

AOI221xp5_ASAP7_75t_L g1444 ( 
.A1(n_1415),
.A2(n_1167),
.B1(n_1183),
.B2(n_1181),
.C(n_1180),
.Y(n_1444)
);

AOI21xp5_ASAP7_75t_L g1445 ( 
.A1(n_1409),
.A2(n_1419),
.B(n_1400),
.Y(n_1445)
);

AOI21xp5_ASAP7_75t_L g1446 ( 
.A1(n_1398),
.A2(n_1127),
.B(n_1115),
.Y(n_1446)
);

A2O1A1Ixp33_ASAP7_75t_SL g1447 ( 
.A1(n_1398),
.A2(n_1140),
.B(n_960),
.C(n_930),
.Y(n_1447)
);

NAND2xp5_ASAP7_75t_L g1448 ( 
.A(n_1396),
.B(n_63),
.Y(n_1448)
);

NOR4xp25_ASAP7_75t_L g1449 ( 
.A(n_1433),
.B(n_64),
.C(n_66),
.D(n_67),
.Y(n_1449)
);

NOR3xp33_ASAP7_75t_L g1450 ( 
.A(n_1443),
.B(n_1066),
.C(n_1037),
.Y(n_1450)
);

AND2x4_ASAP7_75t_L g1451 ( 
.A(n_1442),
.B(n_1140),
.Y(n_1451)
);

NOR3x1_ASAP7_75t_L g1452 ( 
.A(n_1447),
.B(n_1448),
.C(n_1431),
.Y(n_1452)
);

NOR2x1_ASAP7_75t_L g1453 ( 
.A(n_1429),
.B(n_64),
.Y(n_1453)
);

NOR3xp33_ASAP7_75t_L g1454 ( 
.A(n_1426),
.B(n_1066),
.C(n_1075),
.Y(n_1454)
);

NOR3xp33_ASAP7_75t_L g1455 ( 
.A(n_1425),
.B(n_1075),
.C(n_1041),
.Y(n_1455)
);

NOR3xp33_ASAP7_75t_L g1456 ( 
.A(n_1436),
.B(n_1041),
.C(n_1042),
.Y(n_1456)
);

NAND2xp5_ASAP7_75t_SL g1457 ( 
.A(n_1437),
.B(n_1020),
.Y(n_1457)
);

INVx1_ASAP7_75t_L g1458 ( 
.A(n_1432),
.Y(n_1458)
);

NOR3xp33_ASAP7_75t_SL g1459 ( 
.A(n_1445),
.B(n_1428),
.C(n_1439),
.Y(n_1459)
);

AND2x2_ASAP7_75t_L g1460 ( 
.A(n_1440),
.B(n_68),
.Y(n_1460)
);

NAND3xp33_ASAP7_75t_L g1461 ( 
.A(n_1427),
.B(n_953),
.C(n_934),
.Y(n_1461)
);

AND2x2_ASAP7_75t_L g1462 ( 
.A(n_1444),
.B(n_70),
.Y(n_1462)
);

NOR2xp33_ASAP7_75t_L g1463 ( 
.A(n_1434),
.B(n_70),
.Y(n_1463)
);

NAND4xp25_ASAP7_75t_L g1464 ( 
.A(n_1446),
.B(n_960),
.C(n_930),
.D(n_1048),
.Y(n_1464)
);

NOR2xp33_ASAP7_75t_L g1465 ( 
.A(n_1435),
.B(n_71),
.Y(n_1465)
);

NAND4xp75_ASAP7_75t_L g1466 ( 
.A(n_1430),
.B(n_1091),
.C(n_1169),
.D(n_1106),
.Y(n_1466)
);

NOR3x1_ASAP7_75t_L g1467 ( 
.A(n_1441),
.B(n_1091),
.C(n_1051),
.Y(n_1467)
);

NAND2x1_ASAP7_75t_SL g1468 ( 
.A(n_1438),
.B(n_1048),
.Y(n_1468)
);

AOI22xp5_ASAP7_75t_L g1469 ( 
.A1(n_1433),
.A2(n_1106),
.B1(n_916),
.B2(n_920),
.Y(n_1469)
);

NOR2xp67_ASAP7_75t_L g1470 ( 
.A(n_1433),
.B(n_72),
.Y(n_1470)
);

INVx1_ASAP7_75t_L g1471 ( 
.A(n_1448),
.Y(n_1471)
);

AND2x2_ASAP7_75t_L g1472 ( 
.A(n_1448),
.B(n_74),
.Y(n_1472)
);

NAND2xp5_ASAP7_75t_L g1473 ( 
.A(n_1449),
.B(n_1472),
.Y(n_1473)
);

OAI22xp5_ASAP7_75t_L g1474 ( 
.A1(n_1470),
.A2(n_1097),
.B1(n_1138),
.B2(n_1124),
.Y(n_1474)
);

AOI21xp33_ASAP7_75t_L g1475 ( 
.A1(n_1453),
.A2(n_75),
.B(n_77),
.Y(n_1475)
);

NOR3xp33_ASAP7_75t_SL g1476 ( 
.A(n_1457),
.B(n_1176),
.C(n_953),
.Y(n_1476)
);

AOI211xp5_ASAP7_75t_SL g1477 ( 
.A1(n_1463),
.A2(n_1092),
.B(n_1176),
.C(n_1138),
.Y(n_1477)
);

OAI211xp5_ASAP7_75t_SL g1478 ( 
.A1(n_1459),
.A2(n_1124),
.B(n_1072),
.C(n_1092),
.Y(n_1478)
);

NAND3xp33_ASAP7_75t_L g1479 ( 
.A(n_1471),
.B(n_957),
.C(n_1076),
.Y(n_1479)
);

NOR2x1_ASAP7_75t_L g1480 ( 
.A(n_1465),
.B(n_912),
.Y(n_1480)
);

AOI32xp33_ASAP7_75t_L g1481 ( 
.A1(n_1458),
.A2(n_952),
.A3(n_1111),
.B1(n_1117),
.B2(n_1120),
.Y(n_1481)
);

NAND4xp25_ASAP7_75t_L g1482 ( 
.A(n_1452),
.B(n_1111),
.C(n_1092),
.D(n_1117),
.Y(n_1482)
);

NAND3xp33_ASAP7_75t_L g1483 ( 
.A(n_1462),
.B(n_1076),
.C(n_984),
.Y(n_1483)
);

NOR3xp33_ASAP7_75t_L g1484 ( 
.A(n_1461),
.B(n_1120),
.C(n_1054),
.Y(n_1484)
);

NAND4xp25_ASAP7_75t_L g1485 ( 
.A(n_1467),
.B(n_1469),
.C(n_1464),
.D(n_1456),
.Y(n_1485)
);

AOI211xp5_ASAP7_75t_SL g1486 ( 
.A1(n_1460),
.A2(n_1090),
.B(n_98),
.C(n_99),
.Y(n_1486)
);

NOR3xp33_ASAP7_75t_L g1487 ( 
.A(n_1454),
.B(n_1450),
.C(n_1455),
.Y(n_1487)
);

INVx1_ASAP7_75t_SL g1488 ( 
.A(n_1451),
.Y(n_1488)
);

INVx1_ASAP7_75t_L g1489 ( 
.A(n_1473),
.Y(n_1489)
);

AOI22xp5_ASAP7_75t_L g1490 ( 
.A1(n_1475),
.A2(n_1466),
.B1(n_1468),
.B2(n_997),
.Y(n_1490)
);

AOI22xp5_ASAP7_75t_L g1491 ( 
.A1(n_1487),
.A2(n_1079),
.B1(n_1061),
.B2(n_1069),
.Y(n_1491)
);

AOI22xp5_ASAP7_75t_L g1492 ( 
.A1(n_1480),
.A2(n_1079),
.B1(n_1061),
.B2(n_1069),
.Y(n_1492)
);

INVx1_ASAP7_75t_L g1493 ( 
.A(n_1488),
.Y(n_1493)
);

INVx1_ASAP7_75t_L g1494 ( 
.A(n_1474),
.Y(n_1494)
);

INVx1_ASAP7_75t_L g1495 ( 
.A(n_1479),
.Y(n_1495)
);

INVx2_ASAP7_75t_SL g1496 ( 
.A(n_1483),
.Y(n_1496)
);

INVx1_ASAP7_75t_L g1497 ( 
.A(n_1478),
.Y(n_1497)
);

INVx1_ASAP7_75t_L g1498 ( 
.A(n_1485),
.Y(n_1498)
);

NAND2xp5_ASAP7_75t_L g1499 ( 
.A(n_1486),
.B(n_1481),
.Y(n_1499)
);

INVx1_ASAP7_75t_L g1500 ( 
.A(n_1482),
.Y(n_1500)
);

AOI22xp5_ASAP7_75t_L g1501 ( 
.A1(n_1484),
.A2(n_1060),
.B1(n_1130),
.B2(n_1133),
.Y(n_1501)
);

AOI22xp5_ASAP7_75t_L g1502 ( 
.A1(n_1476),
.A2(n_1133),
.B1(n_1130),
.B2(n_1136),
.Y(n_1502)
);

INVx1_ASAP7_75t_L g1503 ( 
.A(n_1477),
.Y(n_1503)
);

HB1xp67_ASAP7_75t_L g1504 ( 
.A(n_1489),
.Y(n_1504)
);

AOI31xp33_ASAP7_75t_L g1505 ( 
.A1(n_1493),
.A2(n_148),
.A3(n_154),
.B(n_156),
.Y(n_1505)
);

NAND5xp2_ASAP7_75t_L g1506 ( 
.A(n_1498),
.B(n_157),
.C(n_159),
.D(n_161),
.E(n_167),
.Y(n_1506)
);

AND2x2_ASAP7_75t_L g1507 ( 
.A(n_1503),
.B(n_1173),
.Y(n_1507)
);

AND2x2_ASAP7_75t_L g1508 ( 
.A(n_1500),
.B(n_1171),
.Y(n_1508)
);

NAND2xp5_ASAP7_75t_L g1509 ( 
.A(n_1495),
.B(n_176),
.Y(n_1509)
);

NOR2xp33_ASAP7_75t_SL g1510 ( 
.A(n_1496),
.B(n_1166),
.Y(n_1510)
);

NAND2xp5_ASAP7_75t_L g1511 ( 
.A(n_1504),
.B(n_1497),
.Y(n_1511)
);

INVx1_ASAP7_75t_L g1512 ( 
.A(n_1509),
.Y(n_1512)
);

NOR3xp33_ASAP7_75t_L g1513 ( 
.A(n_1509),
.B(n_1499),
.C(n_1494),
.Y(n_1513)
);

NAND2xp5_ASAP7_75t_L g1514 ( 
.A(n_1505),
.B(n_1490),
.Y(n_1514)
);

INVxp67_ASAP7_75t_SL g1515 ( 
.A(n_1511),
.Y(n_1515)
);

AOI22xp5_ASAP7_75t_L g1516 ( 
.A1(n_1513),
.A2(n_1508),
.B1(n_1507),
.B2(n_1510),
.Y(n_1516)
);

OAI21x1_ASAP7_75t_L g1517 ( 
.A1(n_1515),
.A2(n_1514),
.B(n_1512),
.Y(n_1517)
);

OAI22x1_ASAP7_75t_L g1518 ( 
.A1(n_1516),
.A2(n_1506),
.B1(n_1491),
.B2(n_1492),
.Y(n_1518)
);

INVx1_ASAP7_75t_L g1519 ( 
.A(n_1517),
.Y(n_1519)
);

INVx1_ASAP7_75t_L g1520 ( 
.A(n_1518),
.Y(n_1520)
);

INVx2_ASAP7_75t_L g1521 ( 
.A(n_1519),
.Y(n_1521)
);

INVx1_ASAP7_75t_L g1522 ( 
.A(n_1520),
.Y(n_1522)
);

AOI21xp33_ASAP7_75t_L g1523 ( 
.A1(n_1521),
.A2(n_1502),
.B(n_1501),
.Y(n_1523)
);

AOI22x1_ASAP7_75t_L g1524 ( 
.A1(n_1522),
.A2(n_179),
.B1(n_182),
.B2(n_184),
.Y(n_1524)
);

AOI22x1_ASAP7_75t_L g1525 ( 
.A1(n_1524),
.A2(n_187),
.B1(n_192),
.B2(n_197),
.Y(n_1525)
);

AOI22xp33_ASAP7_75t_SL g1526 ( 
.A1(n_1525),
.A2(n_1523),
.B1(n_1114),
.B2(n_1113),
.Y(n_1526)
);

AOI221xp5_ASAP7_75t_L g1527 ( 
.A1(n_1526),
.A2(n_198),
.B1(n_201),
.B2(n_202),
.C(n_204),
.Y(n_1527)
);

AOI211xp5_ASAP7_75t_L g1528 ( 
.A1(n_1527),
.A2(n_207),
.B(n_211),
.C(n_212),
.Y(n_1528)
);


endmodule