module fake_netlist_1_3934_n_24 (n_9, n_10, n_4, n_2, n_12, n_11, n_6, n_7, n_1, n_8, n_3, n_5, n_0, n_24, n_27);
input n_9;
input n_10;
input n_4;
input n_2;
input n_12;
input n_11;
input n_6;
input n_7;
input n_1;
input n_8;
input n_3;
input n_5;
input n_0;
output n_24;
output n_27;
wire n_20;
wire n_12;
wire n_7;
wire n_1;
wire n_16;
wire n_22;
wire n_3;
wire n_19;
wire n_10;
wire n_25;
wire n_9;
wire n_13;
wire n_26;
wire n_11;
wire n_0;
wire n_4;
wire n_24;
wire n_6;
wire n_8;
wire n_15;
wire n_21;
wire n_2;
wire n_18;
wire n_17;
wire n_5;
wire n_14;
CKINVDCx16_ASAP7_75t_R g13 ( .A(n_0), .Y(n_13) );
NAND2xp5_ASAP7_75t_SL g14 ( .A(n_12), .B(n_4), .Y(n_14) );
NAND2xp5_ASAP7_75t_L g15 ( .A(n_0), .B(n_1), .Y(n_15) );
INVx1_ASAP7_75t_L g16 ( .A(n_9), .Y(n_16) );
INVx1_ASAP7_75t_L g17 ( .A(n_7), .Y(n_17) );
AOI22xp5_ASAP7_75t_L g18 ( .A1(n_13), .A2(n_15), .B1(n_16), .B2(n_17), .Y(n_18) );
AND2x2_ASAP7_75t_L g19 ( .A(n_14), .B(n_2), .Y(n_19) );
INVx1_ASAP7_75t_L g20 ( .A(n_19), .Y(n_20) );
AND2x2_ASAP7_75t_L g21 ( .A(n_20), .B(n_18), .Y(n_21) );
AND2x2_ASAP7_75t_L g22 ( .A(n_21), .B(n_14), .Y(n_22) );
AOI22xp33_ASAP7_75t_L g23 ( .A1(n_22), .A2(n_3), .B1(n_5), .B2(n_6), .Y(n_23) );
UNKNOWN g24 ( );
INVx1_ASAP7_75t_L g25 ( .A(n_24), .Y(n_25) );
CKINVDCx20_ASAP7_75t_R g26 ( .A(n_25), .Y(n_26) );
AOI22xp33_ASAP7_75t_L g27 ( .A1(n_26), .A2(n_8), .B1(n_10), .B2(n_11), .Y(n_27) );
endmodule