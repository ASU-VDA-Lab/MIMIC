module fake_jpeg_25073_n_222 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_222);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_222;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_121;
wire n_99;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx5_ASAP7_75t_L g16 ( 
.A(n_14),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_12),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

INVxp67_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_10),
.B(n_9),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_3),
.Y(n_23)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_10),
.Y(n_25)
);

INVx11_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_8),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_8),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_26),
.Y(n_34)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_34),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_26),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_35),
.Y(n_54)
);

CKINVDCx16_ASAP7_75t_R g36 ( 
.A(n_22),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_36),
.B(n_39),
.Y(n_49)
);

INVx5_ASAP7_75t_L g37 ( 
.A(n_33),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_37),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_26),
.Y(n_38)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_22),
.B(n_0),
.Y(n_39)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_33),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_40),
.B(n_41),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_33),
.B(n_0),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_24),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_42),
.Y(n_50)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_24),
.Y(n_43)
);

INVx5_ASAP7_75t_L g47 ( 
.A(n_43),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_SL g45 ( 
.A(n_36),
.B(n_25),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_SL g78 ( 
.A(n_45),
.B(n_46),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g46 ( 
.A(n_41),
.B(n_33),
.C(n_30),
.Y(n_46)
);

OR2x2_ASAP7_75t_L g48 ( 
.A(n_39),
.B(n_31),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_SL g85 ( 
.A(n_48),
.B(n_60),
.Y(n_85)
);

OR2x2_ASAP7_75t_SL g53 ( 
.A(n_40),
.B(n_25),
.Y(n_53)
);

A2O1A1Ixp33_ASAP7_75t_L g75 ( 
.A1(n_53),
.A2(n_32),
.B(n_27),
.C(n_29),
.Y(n_75)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_43),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_55),
.B(n_57),
.Y(n_63)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_43),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_37),
.A2(n_24),
.B1(n_30),
.B2(n_31),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_58),
.A2(n_28),
.B1(n_17),
.B2(n_16),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_L g59 ( 
.A1(n_42),
.A2(n_23),
.B1(n_18),
.B2(n_28),
.Y(n_59)
);

OAI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_59),
.A2(n_23),
.B1(n_17),
.B2(n_19),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_34),
.B(n_18),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_34),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_61),
.B(n_38),
.Y(n_71)
);

OAI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_62),
.A2(n_75),
.B1(n_79),
.B2(n_64),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_64),
.A2(n_68),
.B1(n_69),
.B2(n_84),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_44),
.Y(n_65)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_65),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_51),
.B(n_42),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_66),
.B(n_74),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g67 ( 
.A(n_60),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_67),
.B(n_72),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_53),
.A2(n_16),
.B1(n_20),
.B2(n_32),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_46),
.A2(n_29),
.B1(n_27),
.B2(n_21),
.Y(n_69)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_56),
.Y(n_70)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_70),
.Y(n_108)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_71),
.Y(n_99)
);

CKINVDCx16_ASAP7_75t_R g72 ( 
.A(n_51),
.Y(n_72)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_44),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_73),
.B(n_77),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_48),
.B(n_21),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_48),
.B(n_32),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_76),
.B(n_86),
.Y(n_90)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_54),
.Y(n_77)
);

CKINVDCx16_ASAP7_75t_R g79 ( 
.A(n_45),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_79),
.B(n_56),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_49),
.B(n_20),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_SL g107 ( 
.A(n_80),
.B(n_83),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_50),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_81),
.Y(n_89)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_56),
.Y(n_82)
);

BUFx12f_ASAP7_75t_L g105 ( 
.A(n_82),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_49),
.B(n_20),
.Y(n_83)
);

AOI21xp5_ASAP7_75t_SL g84 ( 
.A1(n_55),
.A2(n_29),
.B(n_27),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_57),
.B(n_21),
.Y(n_86)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_65),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_92),
.B(n_96),
.Y(n_116)
);

XOR2xp5_ASAP7_75t_L g93 ( 
.A(n_76),
.B(n_47),
.Y(n_93)
);

XOR2xp5_ASAP7_75t_L g127 ( 
.A(n_93),
.B(n_95),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_72),
.B(n_50),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_94),
.B(n_102),
.Y(n_113)
);

XOR2xp5_ASAP7_75t_L g95 ( 
.A(n_74),
.B(n_47),
.Y(n_95)
);

BUFx5_ASAP7_75t_L g96 ( 
.A(n_70),
.Y(n_96)
);

XOR2xp5_ASAP7_75t_L g98 ( 
.A(n_66),
.B(n_47),
.Y(n_98)
);

XOR2xp5_ASAP7_75t_L g134 ( 
.A(n_98),
.B(n_101),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_SL g115 ( 
.A(n_100),
.B(n_109),
.Y(n_115)
);

XOR2xp5_ASAP7_75t_L g101 ( 
.A(n_78),
.B(n_38),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_78),
.B(n_61),
.C(n_54),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_85),
.B(n_54),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_103),
.B(n_84),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_104),
.A2(n_85),
.B1(n_75),
.B2(n_69),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_81),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_106),
.B(n_111),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_80),
.B(n_15),
.Y(n_109)
);

BUFx5_ASAP7_75t_L g111 ( 
.A(n_82),
.Y(n_111)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_97),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_112),
.B(n_114),
.Y(n_147)
);

BUFx2_ASAP7_75t_L g118 ( 
.A(n_96),
.Y(n_118)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_118),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_119),
.B(n_126),
.Y(n_136)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_94),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_SL g151 ( 
.A(n_120),
.B(n_121),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_89),
.B(n_103),
.Y(n_121)
);

AND2x6_ASAP7_75t_L g122 ( 
.A(n_101),
.B(n_68),
.Y(n_122)
);

NOR3xp33_ASAP7_75t_L g146 ( 
.A(n_122),
.B(n_123),
.C(n_124),
.Y(n_146)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_88),
.Y(n_123)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_102),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_110),
.A2(n_86),
.B1(n_84),
.B2(n_71),
.Y(n_125)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_125),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_99),
.A2(n_63),
.B1(n_52),
.B2(n_77),
.Y(n_126)
);

A2O1A1Ixp33_ASAP7_75t_L g128 ( 
.A1(n_87),
.A2(n_63),
.B(n_2),
.C(n_3),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_L g145 ( 
.A1(n_128),
.A2(n_129),
.B(n_1),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_L g129 ( 
.A1(n_90),
.A2(n_73),
.B(n_2),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_87),
.A2(n_52),
.B1(n_65),
.B2(n_35),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_130),
.A2(n_131),
.B1(n_132),
.B2(n_92),
.Y(n_150)
);

INVxp67_ASAP7_75t_L g131 ( 
.A(n_107),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_110),
.A2(n_35),
.B1(n_2),
.B2(n_3),
.Y(n_132)
);

INVx4_ASAP7_75t_L g133 ( 
.A(n_105),
.Y(n_133)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_133),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_117),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_135),
.B(n_144),
.Y(n_167)
);

INVx5_ASAP7_75t_L g137 ( 
.A(n_118),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_137),
.B(n_148),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_134),
.B(n_98),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_138),
.B(n_140),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_134),
.B(n_95),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_127),
.B(n_93),
.C(n_90),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_141),
.B(n_129),
.C(n_124),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_119),
.B(n_99),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_L g168 ( 
.A1(n_145),
.A2(n_4),
.B(n_5),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_116),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_130),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_149),
.B(n_152),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_150),
.A2(n_112),
.B1(n_131),
.B2(n_91),
.Y(n_164)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_113),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_113),
.Y(n_153)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_153),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_115),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_SL g172 ( 
.A(n_154),
.B(n_15),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g155 ( 
.A(n_127),
.B(n_114),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_155),
.B(n_111),
.Y(n_169)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_125),
.Y(n_156)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_156),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_157),
.B(n_162),
.C(n_169),
.Y(n_178)
);

FAx1_ASAP7_75t_L g159 ( 
.A(n_142),
.B(n_122),
.CI(n_132),
.CON(n_159),
.SN(n_159)
);

OAI21xp5_ASAP7_75t_SL g181 ( 
.A1(n_159),
.A2(n_164),
.B(n_168),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_138),
.B(n_128),
.C(n_133),
.Y(n_162)
);

INVxp67_ASAP7_75t_L g163 ( 
.A(n_147),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_163),
.B(n_166),
.Y(n_176)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_151),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g170 ( 
.A1(n_150),
.A2(n_91),
.B1(n_108),
.B2(n_105),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_170),
.B(n_139),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_172),
.B(n_14),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_140),
.B(n_108),
.C(n_105),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_173),
.B(n_141),
.C(n_155),
.Y(n_182)
);

INVx2_ASAP7_75t_SL g174 ( 
.A(n_160),
.Y(n_174)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_174),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_167),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_175),
.B(n_177),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_165),
.B(n_158),
.Y(n_179)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_179),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_161),
.B(n_143),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_180),
.B(n_185),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_182),
.B(n_186),
.C(n_157),
.Y(n_193)
);

AOI21xp5_ASAP7_75t_L g183 ( 
.A1(n_163),
.A2(n_156),
.B(n_142),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_183),
.B(n_136),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_159),
.A2(n_149),
.B1(n_152),
.B2(n_153),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_184),
.A2(n_187),
.B1(n_136),
.B2(n_162),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_168),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_169),
.B(n_144),
.C(n_146),
.Y(n_186)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_188),
.Y(n_202)
);

AOI22xp33_ASAP7_75t_L g205 ( 
.A1(n_191),
.A2(n_137),
.B1(n_139),
.B2(n_143),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_193),
.B(n_195),
.C(n_178),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_182),
.B(n_171),
.Y(n_195)
);

OAI21x1_ASAP7_75t_L g196 ( 
.A1(n_176),
.A2(n_159),
.B(n_145),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_196),
.B(n_181),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_184),
.B(n_173),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_197),
.B(n_171),
.Y(n_204)
);

NOR2xp67_ASAP7_75t_L g198 ( 
.A(n_190),
.B(n_186),
.Y(n_198)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_198),
.Y(n_207)
);

AND2x2_ASAP7_75t_L g210 ( 
.A(n_199),
.B(n_4),
.Y(n_210)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_200),
.B(n_204),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_197),
.A2(n_183),
.B1(n_187),
.B2(n_181),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_201),
.B(n_205),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_SL g203 ( 
.A(n_189),
.B(n_174),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_203),
.Y(n_209)
);

AOI322xp5_ASAP7_75t_L g206 ( 
.A1(n_202),
.A2(n_188),
.A3(n_194),
.B1(n_195),
.B2(n_193),
.C1(n_178),
.C2(n_192),
.Y(n_206)
);

AO21x1_ASAP7_75t_L g215 ( 
.A1(n_206),
.A2(n_210),
.B(n_12),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_L g212 ( 
.A1(n_207),
.A2(n_202),
.B1(n_204),
.B2(n_201),
.Y(n_212)
);

AOI21xp5_ASAP7_75t_L g216 ( 
.A1(n_212),
.A2(n_213),
.B(n_215),
.Y(n_216)
);

AOI21xp5_ASAP7_75t_SL g213 ( 
.A1(n_211),
.A2(n_209),
.B(n_210),
.Y(n_213)
);

O2A1O1Ixp33_ASAP7_75t_SL g214 ( 
.A1(n_208),
.A2(n_200),
.B(n_6),
.C(n_7),
.Y(n_214)
);

AOI21xp5_ASAP7_75t_L g218 ( 
.A1(n_214),
.A2(n_5),
.B(n_7),
.Y(n_218)
);

AOI21xp5_ASAP7_75t_L g217 ( 
.A1(n_215),
.A2(n_208),
.B(n_6),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_217),
.B(n_218),
.C(n_5),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_216),
.A2(n_105),
.B1(n_7),
.B2(n_9),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_SL g221 ( 
.A(n_219),
.B(n_220),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_221),
.B(n_9),
.Y(n_222)
);


endmodule