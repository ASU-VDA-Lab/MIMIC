module fake_jpeg_3035_n_230 (n_13, n_21, n_53, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_51, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_52, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_230);

input n_13;
input n_21;
input n_53;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_51;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_52;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_230;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_228;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_76;
wire n_154;
wire n_127;
wire n_205;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_155;
wire n_207;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_223;
wire n_171;
wire n_119;
wire n_69;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_143;
wire n_202;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_91;
wire n_54;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_149;
wire n_157;
wire n_87;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx3_ASAP7_75t_L g54 ( 
.A(n_41),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_4),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_49),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_5),
.Y(n_57)
);

BUFx10_ASAP7_75t_L g58 ( 
.A(n_21),
.Y(n_58)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_16),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_28),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_34),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_7),
.Y(n_62)
);

CKINVDCx5p33_ASAP7_75t_R g63 ( 
.A(n_44),
.Y(n_63)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_13),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_16),
.Y(n_65)
);

BUFx5_ASAP7_75t_L g66 ( 
.A(n_2),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_9),
.Y(n_67)
);

BUFx5_ASAP7_75t_L g68 ( 
.A(n_0),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_47),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_20),
.Y(n_70)
);

BUFx12f_ASAP7_75t_L g71 ( 
.A(n_19),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_5),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_32),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_36),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_48),
.Y(n_75)
);

CKINVDCx5p33_ASAP7_75t_R g76 ( 
.A(n_17),
.Y(n_76)
);

INVx6_ASAP7_75t_L g77 ( 
.A(n_52),
.Y(n_77)
);

BUFx8_ASAP7_75t_L g78 ( 
.A(n_40),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_17),
.Y(n_79)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_29),
.Y(n_80)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_78),
.Y(n_81)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_81),
.Y(n_90)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_78),
.Y(n_82)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_82),
.Y(n_99)
);

BUFx5_ASAP7_75t_L g83 ( 
.A(n_78),
.Y(n_83)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_83),
.Y(n_97)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_74),
.Y(n_84)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_84),
.Y(n_101)
);

BUFx4f_ASAP7_75t_L g85 ( 
.A(n_56),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_85),
.Y(n_95)
);

INVx11_ASAP7_75t_L g86 ( 
.A(n_59),
.Y(n_86)
);

CKINVDCx16_ASAP7_75t_R g98 ( 
.A(n_86),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_76),
.B(n_0),
.Y(n_87)
);

OR2x2_ASAP7_75t_L g96 ( 
.A(n_87),
.B(n_88),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_54),
.B(n_53),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_85),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_89),
.B(n_91),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_84),
.B(n_79),
.Y(n_91)
);

INVx6_ASAP7_75t_L g92 ( 
.A(n_85),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_92),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_88),
.A2(n_57),
.B1(n_62),
.B2(n_67),
.Y(n_93)
);

AO22x1_ASAP7_75t_L g110 ( 
.A1(n_93),
.A2(n_70),
.B1(n_59),
.B2(n_71),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_84),
.B(n_65),
.Y(n_94)
);

CKINVDCx16_ASAP7_75t_R g102 ( 
.A(n_94),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_82),
.Y(n_100)
);

INVx4_ASAP7_75t_L g119 ( 
.A(n_100),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_96),
.A2(n_88),
.B1(n_57),
.B2(n_62),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_103),
.A2(n_104),
.B1(n_111),
.B2(n_64),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_96),
.A2(n_67),
.B1(n_70),
.B2(n_77),
.Y(n_104)
);

OAI21xp33_ASAP7_75t_L g105 ( 
.A1(n_89),
.A2(n_87),
.B(n_81),
.Y(n_105)
);

CKINVDCx14_ASAP7_75t_R g124 ( 
.A(n_105),
.Y(n_124)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_101),
.Y(n_107)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_107),
.Y(n_127)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_92),
.Y(n_108)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_108),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_93),
.B(n_85),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_109),
.B(n_113),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_110),
.A2(n_83),
.B1(n_108),
.B2(n_80),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_101),
.A2(n_77),
.B1(n_54),
.B2(n_60),
.Y(n_111)
);

AND2x2_ASAP7_75t_L g112 ( 
.A(n_95),
.B(n_85),
.Y(n_112)
);

CKINVDCx14_ASAP7_75t_R g132 ( 
.A(n_112),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_95),
.B(n_56),
.Y(n_113)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_100),
.Y(n_115)
);

BUFx3_ASAP7_75t_L g121 ( 
.A(n_115),
.Y(n_121)
);

CKINVDCx16_ASAP7_75t_R g116 ( 
.A(n_100),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_116),
.B(n_63),
.Y(n_141)
);

INVx1_ASAP7_75t_SL g117 ( 
.A(n_97),
.Y(n_117)
);

CKINVDCx16_ASAP7_75t_R g122 ( 
.A(n_117),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_L g118 ( 
.A1(n_95),
.A2(n_81),
.B1(n_86),
.B2(n_82),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_118),
.A2(n_112),
.B1(n_90),
.B2(n_98),
.Y(n_128)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_99),
.Y(n_120)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_120),
.Y(n_123)
);

XNOR2xp5_ASAP7_75t_L g125 ( 
.A(n_114),
.B(n_99),
.Y(n_125)
);

XOR2xp5_ASAP7_75t_L g158 ( 
.A(n_125),
.B(n_130),
.Y(n_158)
);

AO21x1_ASAP7_75t_L g126 ( 
.A1(n_109),
.A2(n_97),
.B(n_69),
.Y(n_126)
);

OR2x2_ASAP7_75t_L g165 ( 
.A(n_126),
.B(n_3),
.Y(n_165)
);

INVxp33_ASAP7_75t_L g166 ( 
.A(n_128),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_110),
.A2(n_59),
.B1(n_71),
.B2(n_64),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_129),
.A2(n_143),
.B1(n_50),
.B2(n_46),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_L g130 ( 
.A(n_113),
.B(n_73),
.Y(n_130)
);

OAI32xp33_ASAP7_75t_L g131 ( 
.A1(n_105),
.A2(n_73),
.A3(n_58),
.B1(n_86),
.B2(n_76),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_131),
.B(n_4),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_102),
.B(n_90),
.C(n_75),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_133),
.B(n_136),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_L g134 ( 
.A(n_117),
.B(n_60),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_134),
.B(n_51),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_135),
.A2(n_137),
.B1(n_140),
.B2(n_142),
.Y(n_153)
);

INVxp67_ASAP7_75t_L g136 ( 
.A(n_112),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_115),
.A2(n_71),
.B1(n_83),
.B2(n_72),
.Y(n_140)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_141),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_119),
.A2(n_55),
.B1(n_80),
.B2(n_61),
.Y(n_142)
);

OAI22xp33_ASAP7_75t_SL g143 ( 
.A1(n_106),
.A2(n_58),
.B1(n_66),
.B2(n_68),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_138),
.A2(n_106),
.B1(n_119),
.B2(n_58),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_145),
.A2(n_146),
.B1(n_151),
.B2(n_25),
.Y(n_183)
);

OA21x2_ASAP7_75t_L g146 ( 
.A1(n_124),
.A2(n_137),
.B(n_126),
.Y(n_146)
);

OA22x2_ASAP7_75t_L g148 ( 
.A1(n_136),
.A2(n_63),
.B1(n_68),
.B2(n_66),
.Y(n_148)
);

AO22x1_ASAP7_75t_SL g175 ( 
.A1(n_148),
.A2(n_153),
.B1(n_145),
.B2(n_146),
.Y(n_175)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_139),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_149),
.B(n_150),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_125),
.A2(n_45),
.B1(n_43),
.B2(n_42),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_152),
.A2(n_156),
.B1(n_6),
.B2(n_7),
.Y(n_170)
);

INVx11_ASAP7_75t_L g154 ( 
.A(n_122),
.Y(n_154)
);

INVx13_ASAP7_75t_L g171 ( 
.A(n_154),
.Y(n_171)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_127),
.Y(n_155)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_155),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_132),
.A2(n_39),
.B1(n_38),
.B2(n_37),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_130),
.B(n_1),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_157),
.B(n_159),
.Y(n_180)
);

INVx4_ASAP7_75t_L g159 ( 
.A(n_121),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_123),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_160),
.B(n_161),
.Y(n_187)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_123),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_SL g162 ( 
.A(n_133),
.B(n_1),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_162),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_134),
.B(n_2),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_SL g177 ( 
.A1(n_163),
.A2(n_165),
.B(n_167),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_SL g164 ( 
.A(n_121),
.B(n_3),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_164),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_170),
.B(n_173),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_166),
.A2(n_6),
.B1(n_8),
.B2(n_9),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_172),
.A2(n_175),
.B1(n_176),
.B2(n_183),
.Y(n_191)
);

AOI21xp5_ASAP7_75t_SL g173 ( 
.A1(n_167),
.A2(n_8),
.B(n_10),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_158),
.B(n_35),
.C(n_33),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_174),
.B(n_182),
.C(n_186),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_166),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_SL g178 ( 
.A1(n_144),
.A2(n_31),
.B(n_30),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_178),
.B(n_13),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_158),
.B(n_27),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_SL g195 ( 
.A(n_179),
.B(n_181),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g181 ( 
.A(n_146),
.B(n_26),
.Y(n_181)
);

XOR2xp5_ASAP7_75t_L g182 ( 
.A(n_152),
.B(n_147),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_156),
.B(n_11),
.C(n_12),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g205 ( 
.A(n_189),
.B(n_190),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_187),
.Y(n_190)
);

OAI32xp33_ASAP7_75t_L g192 ( 
.A1(n_180),
.A2(n_154),
.A3(n_165),
.B1(n_151),
.B2(n_148),
.Y(n_192)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_192),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_179),
.B(n_148),
.C(n_159),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_193),
.B(n_148),
.C(n_174),
.Y(n_203)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_185),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_194),
.B(n_196),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_SL g196 ( 
.A(n_169),
.B(n_14),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_184),
.B(n_14),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_SL g204 ( 
.A(n_198),
.B(n_186),
.Y(n_204)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_168),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_SL g207 ( 
.A(n_199),
.B(n_171),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_191),
.A2(n_175),
.B1(n_181),
.B2(n_182),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_200),
.A2(n_201),
.B1(n_15),
.B2(n_19),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_191),
.A2(n_175),
.B1(n_173),
.B2(n_177),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_197),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_L g213 ( 
.A1(n_202),
.A2(n_207),
.B1(n_195),
.B2(n_18),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g214 ( 
.A(n_203),
.B(n_15),
.Y(n_214)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_204),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_188),
.B(n_171),
.C(n_18),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_206),
.B(n_195),
.Y(n_211)
);

AOI21xp5_ASAP7_75t_L g210 ( 
.A1(n_209),
.A2(n_193),
.B(n_188),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_L g217 ( 
.A1(n_210),
.A2(n_213),
.B1(n_206),
.B2(n_205),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_211),
.B(n_203),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_214),
.B(n_216),
.Y(n_220)
);

XOR2xp5_ASAP7_75t_L g219 ( 
.A(n_215),
.B(n_208),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_L g216 ( 
.A(n_200),
.B(n_20),
.Y(n_216)
);

AOI21xp5_ASAP7_75t_SL g222 ( 
.A1(n_217),
.A2(n_218),
.B(n_211),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_219),
.A2(n_216),
.B1(n_212),
.B2(n_214),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_221),
.B(n_222),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_223),
.B(n_219),
.C(n_220),
.Y(n_224)
);

AOI31xp67_ASAP7_75t_L g225 ( 
.A1(n_224),
.A2(n_220),
.A3(n_22),
.B(n_23),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_225),
.B(n_21),
.Y(n_226)
);

AOI21xp5_ASAP7_75t_L g227 ( 
.A1(n_226),
.A2(n_22),
.B(n_23),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_227),
.B(n_24),
.C(n_25),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_228),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_229),
.B(n_24),
.Y(n_230)
);


endmodule