module fake_jpeg_29285_n_277 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_277);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_277;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_252;
wire n_251;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_272;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_258;
wire n_96;

INVx1_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

INVx11_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_15),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_17),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_17),
.Y(n_23)
);

BUFx2_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_16),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_5),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_5),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_9),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

INVx11_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_1),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_7),
.Y(n_34)
);

BUFx16f_ASAP7_75t_L g35 ( 
.A(n_0),
.Y(n_35)
);

CKINVDCx16_ASAP7_75t_R g36 ( 
.A(n_4),
.Y(n_36)
);

CKINVDCx14_ASAP7_75t_R g37 ( 
.A(n_5),
.Y(n_37)
);

BUFx5_ASAP7_75t_L g38 ( 
.A(n_9),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_7),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_10),
.Y(n_40)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_35),
.Y(n_41)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_41),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_24),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_42),
.B(n_47),
.Y(n_68)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_27),
.Y(n_43)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_43),
.Y(n_67)
);

BUFx10_ASAP7_75t_L g44 ( 
.A(n_35),
.Y(n_44)
);

BUFx10_ASAP7_75t_L g85 ( 
.A(n_44),
.Y(n_85)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_38),
.Y(n_45)
);

INVx8_ASAP7_75t_L g65 ( 
.A(n_45),
.Y(n_65)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_27),
.Y(n_46)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_46),
.Y(n_82)
);

BUFx12_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_19),
.Y(n_48)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_48),
.Y(n_75)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_49),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_24),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_50),
.B(n_51),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_24),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_24),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_52),
.B(n_58),
.Y(n_80)
);

INVx11_ASAP7_75t_L g53 ( 
.A(n_35),
.Y(n_53)
);

INVx5_ASAP7_75t_L g76 ( 
.A(n_53),
.Y(n_76)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_30),
.Y(n_54)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_54),
.Y(n_84)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_38),
.Y(n_55)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_55),
.Y(n_97)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_30),
.Y(n_56)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_56),
.Y(n_88)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_19),
.Y(n_57)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_57),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_26),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_40),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_59),
.Y(n_73)
);

AOI21xp5_ASAP7_75t_L g60 ( 
.A1(n_19),
.A2(n_0),
.B(n_1),
.Y(n_60)
);

A2O1A1Ixp33_ASAP7_75t_L g74 ( 
.A1(n_60),
.A2(n_36),
.B(n_37),
.C(n_39),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_40),
.Y(n_61)
);

BUFx12f_ASAP7_75t_L g78 ( 
.A(n_61),
.Y(n_78)
);

INVx13_ASAP7_75t_L g62 ( 
.A(n_37),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_62),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_26),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_63),
.B(n_23),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_40),
.Y(n_64)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_64),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_58),
.B(n_28),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_69),
.B(n_81),
.Y(n_107)
);

AND2x2_ASAP7_75t_L g70 ( 
.A(n_43),
.B(n_38),
.Y(n_70)
);

AND2x2_ASAP7_75t_L g104 ( 
.A(n_70),
.B(n_72),
.Y(n_104)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_48),
.Y(n_71)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_71),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g72 ( 
.A(n_57),
.B(n_40),
.C(n_39),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_74),
.B(n_87),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_63),
.B(n_28),
.Y(n_81)
);

HB1xp67_ASAP7_75t_L g83 ( 
.A(n_41),
.Y(n_83)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_83),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_46),
.B(n_33),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_54),
.B(n_33),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_89),
.B(n_92),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_56),
.B(n_29),
.Y(n_92)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_61),
.Y(n_93)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_93),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_60),
.B(n_29),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_94),
.B(n_21),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_SL g102 ( 
.A(n_95),
.B(n_98),
.Y(n_102)
);

AOI21xp33_ASAP7_75t_SL g96 ( 
.A1(n_49),
.A2(n_36),
.B(n_32),
.Y(n_96)
);

AND2x2_ASAP7_75t_SL g103 ( 
.A(n_96),
.B(n_45),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_44),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_L g99 ( 
.A1(n_96),
.A2(n_64),
.B1(n_59),
.B2(n_61),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_99),
.A2(n_49),
.B1(n_53),
.B2(n_73),
.Y(n_147)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_78),
.Y(n_100)
);

INVx4_ASAP7_75t_L g143 ( 
.A(n_100),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_103),
.A2(n_106),
.B1(n_117),
.B2(n_79),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_105),
.A2(n_126),
.B1(n_18),
.B2(n_31),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_72),
.A2(n_18),
.B1(n_50),
.B2(n_52),
.Y(n_106)
);

BUFx3_ASAP7_75t_L g108 ( 
.A(n_76),
.Y(n_108)
);

INVx3_ASAP7_75t_L g160 ( 
.A(n_108),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_80),
.B(n_21),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_109),
.B(n_111),
.Y(n_141)
);

HB1xp67_ASAP7_75t_L g110 ( 
.A(n_97),
.Y(n_110)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_110),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_77),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_67),
.B(n_25),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_112),
.B(n_114),
.Y(n_154)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_78),
.Y(n_113)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_113),
.Y(n_138)
);

CKINVDCx16_ASAP7_75t_R g114 ( 
.A(n_82),
.Y(n_114)
);

OAI22xp33_ASAP7_75t_L g117 ( 
.A1(n_91),
.A2(n_42),
.B1(n_51),
.B2(n_55),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_84),
.B(n_25),
.Y(n_119)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_119),
.Y(n_135)
);

INVx2_ASAP7_75t_SL g120 ( 
.A(n_79),
.Y(n_120)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_120),
.Y(n_150)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_71),
.Y(n_121)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_121),
.Y(n_145)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_78),
.Y(n_123)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_123),
.Y(n_155)
);

INVx4_ASAP7_75t_L g124 ( 
.A(n_66),
.Y(n_124)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_124),
.Y(n_157)
);

INVxp67_ASAP7_75t_L g125 ( 
.A(n_68),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_125),
.B(n_127),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_88),
.A2(n_31),
.B1(n_34),
.B2(n_49),
.Y(n_126)
);

CKINVDCx16_ASAP7_75t_R g127 ( 
.A(n_70),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_73),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_128),
.B(n_129),
.Y(n_134)
);

CKINVDCx16_ASAP7_75t_R g129 ( 
.A(n_85),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_75),
.B(n_44),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_130),
.B(n_131),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_85),
.Y(n_131)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_90),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_132),
.B(n_85),
.Y(n_144)
);

XOR2xp5_ASAP7_75t_L g137 ( 
.A(n_104),
.B(n_74),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_137),
.B(n_124),
.C(n_86),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_139),
.A2(n_23),
.B1(n_20),
.B2(n_2),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_SL g140 ( 
.A1(n_104),
.A2(n_66),
.B(n_97),
.Y(n_140)
);

AOI21xp5_ASAP7_75t_L g166 ( 
.A1(n_140),
.A2(n_146),
.B(n_120),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_142),
.A2(n_108),
.B1(n_113),
.B2(n_123),
.Y(n_164)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_144),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_SL g146 ( 
.A1(n_104),
.A2(n_86),
.B(n_34),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_147),
.A2(n_149),
.B1(n_153),
.B2(n_156),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_122),
.A2(n_105),
.B1(n_103),
.B2(n_101),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_101),
.B(n_103),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_151),
.B(n_44),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_117),
.A2(n_65),
.B1(n_76),
.B2(n_18),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_152),
.A2(n_2),
.B1(n_3),
.B2(n_6),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_125),
.A2(n_130),
.B1(n_107),
.B2(n_132),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_116),
.A2(n_121),
.B1(n_118),
.B2(n_128),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_116),
.A2(n_65),
.B1(n_20),
.B2(n_32),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_158),
.A2(n_159),
.B1(n_0),
.B2(n_1),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_115),
.A2(n_32),
.B1(n_20),
.B2(n_22),
.Y(n_159)
);

NOR3xp33_ASAP7_75t_L g161 ( 
.A(n_151),
.B(n_133),
.C(n_135),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_161),
.B(n_163),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_141),
.B(n_102),
.Y(n_162)
);

CKINVDCx14_ASAP7_75t_R g206 ( 
.A(n_162),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_164),
.A2(n_184),
.B1(n_185),
.B2(n_8),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_L g165 ( 
.A1(n_136),
.A2(n_120),
.B(n_62),
.Y(n_165)
);

AOI21xp5_ASAP7_75t_SL g191 ( 
.A1(n_165),
.A2(n_148),
.B(n_160),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_SL g188 ( 
.A1(n_166),
.A2(n_148),
.B(n_157),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_167),
.B(n_168),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_136),
.B(n_100),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_153),
.B(n_22),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_169),
.B(n_174),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_154),
.B(n_133),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_170),
.B(n_175),
.Y(n_192)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_144),
.Y(n_172)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_172),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_173),
.A2(n_180),
.B1(n_176),
.B2(n_165),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g174 ( 
.A(n_137),
.B(n_47),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_134),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_140),
.B(n_47),
.C(n_11),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_176),
.B(n_183),
.Y(n_189)
);

INVx13_ASAP7_75t_L g177 ( 
.A(n_160),
.Y(n_177)
);

INVxp33_ASAP7_75t_L g208 ( 
.A(n_177),
.Y(n_208)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_145),
.Y(n_179)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_179),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_L g199 ( 
.A1(n_180),
.A2(n_138),
.B1(n_143),
.B2(n_159),
.Y(n_199)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_134),
.Y(n_181)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_181),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_155),
.B(n_12),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_182),
.B(n_187),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g183 ( 
.A(n_146),
.B(n_47),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_L g185 ( 
.A1(n_142),
.A2(n_2),
.B1(n_3),
.B2(n_6),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_150),
.Y(n_186)
);

CKINVDCx16_ASAP7_75t_R g198 ( 
.A(n_186),
.Y(n_198)
);

INVx6_ASAP7_75t_SL g187 ( 
.A(n_150),
.Y(n_187)
);

INVxp67_ASAP7_75t_L g221 ( 
.A(n_188),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_SL g223 ( 
.A1(n_191),
.A2(n_204),
.B(n_173),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_SL g194 ( 
.A(n_169),
.B(n_152),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_194),
.B(n_184),
.Y(n_215)
);

OA21x2_ASAP7_75t_L g195 ( 
.A1(n_166),
.A2(n_147),
.B(n_138),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_195),
.B(n_199),
.Y(n_225)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_186),
.Y(n_200)
);

INVx1_ASAP7_75t_SL g210 ( 
.A(n_200),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_201),
.B(n_178),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_178),
.A2(n_158),
.B1(n_156),
.B2(n_143),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_203),
.A2(n_205),
.B1(n_8),
.B2(n_10),
.Y(n_226)
);

OAI21xp5_ASAP7_75t_SL g204 ( 
.A1(n_163),
.A2(n_3),
.B(n_6),
.Y(n_204)
);

NAND3xp33_ASAP7_75t_L g211 ( 
.A(n_206),
.B(n_167),
.C(n_168),
.Y(n_211)
);

NAND3xp33_ASAP7_75t_L g238 ( 
.A(n_211),
.B(n_212),
.C(n_216),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_SL g212 ( 
.A(n_192),
.B(n_181),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_197),
.Y(n_213)
);

INVxp67_ASAP7_75t_L g235 ( 
.A(n_213),
.Y(n_235)
);

OAI21xp5_ASAP7_75t_L g214 ( 
.A1(n_191),
.A2(n_172),
.B(n_171),
.Y(n_214)
);

OAI21xp5_ASAP7_75t_L g236 ( 
.A1(n_214),
.A2(n_224),
.B(n_195),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_215),
.A2(n_222),
.B1(n_226),
.B2(n_199),
.Y(n_230)
);

OA21x2_ASAP7_75t_SL g216 ( 
.A1(n_209),
.A2(n_174),
.B(n_183),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_200),
.Y(n_217)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_217),
.Y(n_231)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_196),
.Y(n_218)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_218),
.Y(n_232)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_196),
.Y(n_219)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_219),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_189),
.B(n_171),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_220),
.B(n_209),
.Y(n_233)
);

AOI21xp5_ASAP7_75t_L g234 ( 
.A1(n_223),
.A2(n_188),
.B(n_205),
.Y(n_234)
);

OAI21xp5_ASAP7_75t_L g224 ( 
.A1(n_195),
.A2(n_187),
.B(n_177),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_189),
.B(n_13),
.C(n_14),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_227),
.B(n_201),
.C(n_204),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_228),
.B(n_223),
.Y(n_246)
);

OAI21xp5_ASAP7_75t_SL g229 ( 
.A1(n_221),
.A2(n_193),
.B(n_202),
.Y(n_229)
);

AOI21xp5_ASAP7_75t_L g251 ( 
.A1(n_229),
.A2(n_239),
.B(n_240),
.Y(n_251)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_230),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g248 ( 
.A(n_233),
.B(n_225),
.Y(n_248)
);

OAI21xp5_ASAP7_75t_L g241 ( 
.A1(n_234),
.A2(n_224),
.B(n_225),
.Y(n_241)
);

INVxp67_ASAP7_75t_L g245 ( 
.A(n_236),
.Y(n_245)
);

AO221x1_ASAP7_75t_L g239 ( 
.A1(n_218),
.A2(n_202),
.B1(n_190),
.B2(n_208),
.C(n_198),
.Y(n_239)
);

OAI21xp5_ASAP7_75t_L g240 ( 
.A1(n_221),
.A2(n_207),
.B(n_190),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_241),
.B(n_242),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_SL g242 ( 
.A(n_233),
.B(n_220),
.Y(n_242)
);

HB1xp67_ASAP7_75t_L g243 ( 
.A(n_240),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_243),
.B(n_247),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_228),
.B(n_214),
.C(n_207),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_244),
.B(n_249),
.C(n_236),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_246),
.B(n_248),
.Y(n_252)
);

CKINVDCx16_ASAP7_75t_R g247 ( 
.A(n_232),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_235),
.B(n_227),
.C(n_217),
.Y(n_249)
);

OAI21xp5_ASAP7_75t_SL g253 ( 
.A1(n_245),
.A2(n_235),
.B(n_238),
.Y(n_253)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_253),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_254),
.B(n_252),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_251),
.B(n_213),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_256),
.B(n_258),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_250),
.A2(n_226),
.B1(n_203),
.B2(n_245),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_249),
.B(n_237),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_259),
.B(n_257),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_260),
.B(n_263),
.Y(n_268)
);

AOI322xp5_ASAP7_75t_L g261 ( 
.A1(n_255),
.A2(n_248),
.A3(n_244),
.B1(n_231),
.B2(n_210),
.C1(n_242),
.C2(n_219),
.Y(n_261)
);

INVxp67_ASAP7_75t_L g269 ( 
.A(n_261),
.Y(n_269)
);

OAI21xp5_ASAP7_75t_L g263 ( 
.A1(n_254),
.A2(n_210),
.B(n_198),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_265),
.B(n_194),
.Y(n_266)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_266),
.Y(n_273)
);

AOI21xp5_ASAP7_75t_SL g267 ( 
.A1(n_262),
.A2(n_255),
.B(n_15),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_267),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_264),
.B(n_14),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_270),
.B(n_16),
.C(n_261),
.Y(n_271)
);

AOI21xp5_ASAP7_75t_L g275 ( 
.A1(n_271),
.A2(n_269),
.B(n_268),
.Y(n_275)
);

INVxp33_ASAP7_75t_L g274 ( 
.A(n_273),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_274),
.B(n_275),
.C(n_272),
.Y(n_276)
);

XOR2xp5_ASAP7_75t_L g277 ( 
.A(n_276),
.B(n_267),
.Y(n_277)
);


endmodule