module real_jpeg_4260_n_19 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_16, n_15, n_13, n_19);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;

output n_19;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_95;
wire n_541;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_203;
wire n_198;
wire n_500;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_366;
wire n_332;
wire n_456;
wire n_259;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_538;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_216;
wire n_128;
wire n_202;
wire n_483;
wire n_367;
wire n_127;
wire n_365;
wire n_356;
wire n_423;
wire n_464;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_233;
wire n_73;
wire n_532;
wire n_348;
wire n_516;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_288;
wire n_525;
wire n_83;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_338;
wire n_175;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_372;
wire n_219;
wire n_470;
wire n_122;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_533;
wire n_289;
wire n_117;
wire n_193;
wire n_411;
wire n_382;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_25;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_215;
wire n_166;
wire n_176;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_412;
wire n_120;
wire n_155;
wire n_405;
wire n_319;
wire n_93;
wire n_487;
wire n_242;
wire n_493;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_531;
wire n_112;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_536;
wire n_148;
wire n_373;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_375;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_537;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_539;
wire n_512;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_534;
wire n_256;
wire n_520;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_343;
wire n_292;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_299;
wire n_243;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_540;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_530;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_438;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_447;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

AOI22xp33_ASAP7_75t_L g215 ( 
.A1(n_0),
.A2(n_134),
.B1(n_216),
.B2(n_217),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_0),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_L g233 ( 
.A1(n_0),
.A2(n_187),
.B1(n_194),
.B2(n_216),
.Y(n_233)
);

AOI22xp33_ASAP7_75t_SL g308 ( 
.A1(n_0),
.A2(n_216),
.B1(n_309),
.B2(n_311),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_L g436 ( 
.A1(n_0),
.A2(n_33),
.B1(n_140),
.B2(n_216),
.Y(n_436)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_1),
.A2(n_48),
.B1(n_52),
.B2(n_53),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_1),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g318 ( 
.A1(n_1),
.A2(n_53),
.B1(n_319),
.B2(n_322),
.Y(n_318)
);

OAI22xp33_ASAP7_75t_SL g394 ( 
.A1(n_1),
.A2(n_53),
.B1(n_174),
.B2(n_395),
.Y(n_394)
);

AOI22xp33_ASAP7_75t_SL g408 ( 
.A1(n_1),
.A2(n_53),
.B1(n_96),
.B2(n_409),
.Y(n_408)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_2),
.A2(n_95),
.B1(n_99),
.B2(n_101),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_2),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_2),
.A2(n_101),
.B1(n_131),
.B2(n_133),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_SL g145 ( 
.A1(n_2),
.A2(n_101),
.B1(n_138),
.B2(n_146),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g389 ( 
.A1(n_2),
.A2(n_101),
.B1(n_390),
.B2(n_391),
.Y(n_389)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_3),
.A2(n_88),
.B1(n_91),
.B2(n_92),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_3),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_3),
.A2(n_92),
.B1(n_138),
.B2(n_139),
.Y(n_137)
);

OAI22xp33_ASAP7_75t_SL g386 ( 
.A1(n_3),
.A2(n_92),
.B1(n_387),
.B2(n_388),
.Y(n_386)
);

OAI22xp5_ASAP7_75t_L g418 ( 
.A1(n_3),
.A2(n_92),
.B1(n_288),
.B2(n_419),
.Y(n_418)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_4),
.A2(n_171),
.B1(n_173),
.B2(n_174),
.Y(n_170)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_4),
.Y(n_173)
);

AOI22xp33_ASAP7_75t_L g206 ( 
.A1(n_4),
.A2(n_173),
.B1(n_207),
.B2(n_211),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_4),
.A2(n_90),
.B1(n_100),
.B2(n_173),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_L g368 ( 
.A1(n_4),
.A2(n_149),
.B1(n_173),
.B2(n_345),
.Y(n_368)
);

BUFx5_ASAP7_75t_L g199 ( 
.A(n_5),
.Y(n_199)
);

BUFx6f_ASAP7_75t_L g205 ( 
.A(n_5),
.Y(n_205)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_5),
.Y(n_229)
);

INVx8_ASAP7_75t_L g244 ( 
.A(n_5),
.Y(n_244)
);

BUFx6f_ASAP7_75t_L g284 ( 
.A(n_5),
.Y(n_284)
);

BUFx6f_ASAP7_75t_L g425 ( 
.A(n_5),
.Y(n_425)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_6),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_6),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_6),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_6),
.Y(n_52)
);

BUFx5_ASAP7_75t_L g58 ( 
.A(n_6),
.Y(n_58)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_6),
.Y(n_60)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_6),
.Y(n_151)
);

BUFx5_ASAP7_75t_L g339 ( 
.A(n_6),
.Y(n_339)
);

INVx3_ASAP7_75t_L g346 ( 
.A(n_6),
.Y(n_346)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

BUFx5_ASAP7_75t_L g36 ( 
.A(n_7),
.Y(n_36)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_7),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g342 ( 
.A(n_7),
.Y(n_342)
);

INVx3_ASAP7_75t_L g538 ( 
.A(n_8),
.Y(n_538)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_9),
.Y(n_112)
);

BUFx3_ASAP7_75t_L g121 ( 
.A(n_9),
.Y(n_121)
);

INVx8_ASAP7_75t_L g85 ( 
.A(n_10),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_11),
.Y(n_123)
);

BUFx3_ASAP7_75t_L g125 ( 
.A(n_11),
.Y(n_125)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_11),
.Y(n_192)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_12),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g541 ( 
.A(n_13),
.Y(n_541)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_14),
.A2(n_57),
.B1(n_59),
.B2(n_61),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_14),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_L g352 ( 
.A1(n_14),
.A2(n_61),
.B1(n_353),
.B2(n_357),
.Y(n_352)
);

OAI22xp5_ASAP7_75t_L g396 ( 
.A1(n_14),
.A2(n_61),
.B1(n_397),
.B2(n_399),
.Y(n_396)
);

OAI22xp5_ASAP7_75t_SL g447 ( 
.A1(n_14),
.A2(n_61),
.B1(n_311),
.B2(n_448),
.Y(n_447)
);

OAI22xp33_ASAP7_75t_SL g186 ( 
.A1(n_15),
.A2(n_187),
.B1(n_193),
.B2(n_194),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_15),
.Y(n_193)
);

AOI22xp33_ASAP7_75t_SL g255 ( 
.A1(n_15),
.A2(n_131),
.B1(n_193),
.B2(n_256),
.Y(n_255)
);

AOI22xp33_ASAP7_75t_L g371 ( 
.A1(n_15),
.A2(n_193),
.B1(n_343),
.B2(n_372),
.Y(n_371)
);

AOI22xp5_ASAP7_75t_L g411 ( 
.A1(n_15),
.A2(n_193),
.B1(n_412),
.B2(n_413),
.Y(n_411)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_16),
.Y(n_41)
);

AOI22xp33_ASAP7_75t_SL g164 ( 
.A1(n_17),
.A2(n_165),
.B1(n_167),
.B2(n_168),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_17),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_17),
.B(n_182),
.C(n_183),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g221 ( 
.A(n_17),
.B(n_78),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_17),
.B(n_228),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_17),
.B(n_129),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_17),
.B(n_270),
.Y(n_269)
);

AOI22xp33_ASAP7_75t_L g277 ( 
.A1(n_18),
.A2(n_278),
.B1(n_280),
.B2(n_281),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_18),
.Y(n_280)
);

AOI22xp33_ASAP7_75t_SL g375 ( 
.A1(n_18),
.A2(n_174),
.B1(n_280),
.B2(n_376),
.Y(n_375)
);

AOI22xp5_ASAP7_75t_L g403 ( 
.A1(n_18),
.A2(n_280),
.B1(n_286),
.B2(n_404),
.Y(n_403)
);

OAI22xp33_ASAP7_75t_L g461 ( 
.A1(n_18),
.A2(n_280),
.B1(n_339),
.B2(n_462),
.Y(n_461)
);

AOI21xp5_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_536),
.B(n_539),
.Y(n_19)
);

XNOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_154),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_152),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_SL g22 ( 
.A(n_23),
.B(n_144),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_23),
.B(n_144),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_136),
.C(n_141),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_SL g531 ( 
.A1(n_24),
.A2(n_25),
.B1(n_532),
.B2(n_533),
.Y(n_531)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

MAJIxp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_62),
.C(n_102),
.Y(n_25)
);

XNOR2xp5_ASAP7_75t_SL g523 ( 
.A(n_26),
.B(n_524),
.Y(n_523)
);

OAI22xp5_ASAP7_75t_SL g26 ( 
.A1(n_27),
.A2(n_47),
.B1(n_54),
.B2(n_56),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_27),
.A2(n_54),
.B1(n_56),
.B2(n_137),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_27),
.A2(n_54),
.B1(n_137),
.B2(n_145),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_SL g410 ( 
.A1(n_27),
.A2(n_367),
.B(n_411),
.Y(n_410)
);

OAI22xp5_ASAP7_75t_L g435 ( 
.A1(n_27),
.A2(n_37),
.B1(n_411),
.B2(n_436),
.Y(n_435)
);

OAI22xp5_ASAP7_75t_SL g508 ( 
.A1(n_27),
.A2(n_47),
.B1(n_54),
.B2(n_509),
.Y(n_508)
);

INVx2_ASAP7_75t_SL g27 ( 
.A(n_28),
.Y(n_27)
);

AOI21xp5_ASAP7_75t_L g364 ( 
.A1(n_28),
.A2(n_365),
.B(n_366),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_28),
.B(n_368),
.Y(n_463)
);

AND2x2_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_37),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_L g29 ( 
.A1(n_30),
.A2(n_32),
.B1(n_34),
.B2(n_35),
.Y(n_29)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx5_ASAP7_75t_L g38 ( 
.A(n_31),
.Y(n_38)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx4_ASAP7_75t_L g412 ( 
.A(n_33),
.Y(n_412)
);

INVx4_ASAP7_75t_L g140 ( 
.A(n_34),
.Y(n_140)
);

INVx2_ASAP7_75t_L g462 ( 
.A(n_34),
.Y(n_462)
);

INVx3_ASAP7_75t_SL g35 ( 
.A(n_36),
.Y(n_35)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_37),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_37),
.B(n_168),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_L g37 ( 
.A1(n_38),
.A2(n_39),
.B1(n_42),
.B2(n_44),
.Y(n_37)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx4_ASAP7_75t_L g287 ( 
.A(n_40),
.Y(n_287)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

BUFx5_ASAP7_75t_L g43 ( 
.A(n_41),
.Y(n_43)
);

INVx6_ASAP7_75t_L g71 ( 
.A(n_41),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g267 ( 
.A(n_41),
.Y(n_267)
);

BUFx6f_ASAP7_75t_L g373 ( 
.A(n_41),
.Y(n_373)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_42),
.Y(n_77)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g90 ( 
.A(n_43),
.Y(n_90)
);

INVx6_ASAP7_75t_L g337 ( 
.A(n_43),
.Y(n_337)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

OAI32xp33_ASAP7_75t_L g333 ( 
.A1(n_45),
.A2(n_334),
.A3(n_338),
.B1(n_340),
.B2(n_344),
.Y(n_333)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_52),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_L g473 ( 
.A1(n_54),
.A2(n_436),
.B(n_463),
.Y(n_473)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_55),
.B(n_368),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_55),
.B(n_461),
.Y(n_460)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g524 ( 
.A1(n_62),
.A2(n_102),
.B1(n_103),
.B2(n_525),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_62),
.Y(n_525)
);

OAI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_63),
.A2(n_87),
.B1(n_93),
.B2(n_94),
.Y(n_62)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_63),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g370 ( 
.A1(n_63),
.A2(n_93),
.B1(n_308),
.B2(n_371),
.Y(n_370)
);

OAI22xp5_ASAP7_75t_SL g402 ( 
.A1(n_63),
.A2(n_93),
.B1(n_403),
.B2(n_408),
.Y(n_402)
);

OAI22xp5_ASAP7_75t_SL g512 ( 
.A1(n_63),
.A2(n_87),
.B1(n_93),
.B2(n_513),
.Y(n_512)
);

OR2x2_ASAP7_75t_L g63 ( 
.A(n_64),
.B(n_78),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_L g64 ( 
.A1(n_65),
.A2(n_68),
.B1(n_72),
.B2(n_77),
.Y(n_64)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_66),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g293 ( 
.A(n_66),
.Y(n_293)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_67),
.Y(n_76)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_67),
.Y(n_297)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx5_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_71),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_71),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g271 ( 
.A(n_71),
.Y(n_271)
);

INVx2_ASAP7_75t_L g312 ( 
.A(n_71),
.Y(n_312)
);

BUFx6f_ASAP7_75t_L g407 ( 
.A(n_71),
.Y(n_407)
);

INVx1_ASAP7_75t_SL g72 ( 
.A(n_73),
.Y(n_72)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_77),
.Y(n_91)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_78),
.Y(n_93)
);

OAI21xp5_ASAP7_75t_SL g141 ( 
.A1(n_78),
.A2(n_142),
.B(n_143),
.Y(n_141)
);

AOI22x1_ASAP7_75t_L g437 ( 
.A1(n_78),
.A2(n_142),
.B1(n_314),
.B2(n_438),
.Y(n_437)
);

AOI22xp5_ASAP7_75t_SL g445 ( 
.A1(n_78),
.A2(n_142),
.B1(n_446),
.B2(n_447),
.Y(n_445)
);

AO22x2_ASAP7_75t_L g78 ( 
.A1(n_79),
.A2(n_80),
.B1(n_81),
.B2(n_86),
.Y(n_78)
);

INVx6_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVx3_ASAP7_75t_SL g81 ( 
.A(n_82),
.Y(n_81)
);

BUFx2_ASAP7_75t_L g400 ( 
.A(n_82),
.Y(n_400)
);

INVx8_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx6_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_84),
.Y(n_86)
);

INVx6_ASAP7_75t_L g109 ( 
.A(n_84),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_84),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g167 ( 
.A(n_84),
.Y(n_167)
);

INVx5_ASAP7_75t_L g290 ( 
.A(n_84),
.Y(n_290)
);

BUFx6f_ASAP7_75t_L g395 ( 
.A(n_84),
.Y(n_395)
);

INVx11_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_85),
.Y(n_117)
);

BUFx5_ASAP7_75t_L g176 ( 
.A(n_85),
.Y(n_176)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_85),
.Y(n_260)
);

BUFx6f_ASAP7_75t_L g398 ( 
.A(n_85),
.Y(n_398)
);

BUFx3_ASAP7_75t_L g166 ( 
.A(n_86),
.Y(n_166)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_93),
.B(n_273),
.Y(n_272)
);

OAI21xp5_ASAP7_75t_SL g307 ( 
.A1(n_93),
.A2(n_308),
.B(n_313),
.Y(n_307)
);

INVxp67_ASAP7_75t_L g143 ( 
.A(n_94),
.Y(n_143)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

INVx4_ASAP7_75t_SL g96 ( 
.A(n_97),
.Y(n_96)
);

INVx5_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

BUFx12f_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g510 ( 
.A1(n_102),
.A2(n_103),
.B1(n_511),
.B2(n_512),
.Y(n_510)
);

MAJIxp5_ASAP7_75t_L g519 ( 
.A(n_102),
.B(n_508),
.C(n_511),
.Y(n_519)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

AOI21xp5_ASAP7_75t_SL g103 ( 
.A1(n_104),
.A2(n_128),
.B(n_130),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_SL g163 ( 
.A1(n_104),
.A2(n_164),
.B(n_169),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_104),
.A2(n_128),
.B1(n_215),
.B2(n_255),
.Y(n_254)
);

OAI21xp5_ASAP7_75t_SL g304 ( 
.A1(n_104),
.A2(n_169),
.B(n_255),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_SL g429 ( 
.A1(n_104),
.A2(n_128),
.B1(n_375),
.B2(n_430),
.Y(n_429)
);

INVx2_ASAP7_75t_SL g104 ( 
.A(n_105),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_105),
.B(n_170),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g393 ( 
.A1(n_105),
.A2(n_129),
.B1(n_394),
.B2(n_396),
.Y(n_393)
);

AOI22xp5_ASAP7_75t_L g417 ( 
.A1(n_105),
.A2(n_129),
.B1(n_396),
.B2(n_418),
.Y(n_417)
);

AOI22xp5_ASAP7_75t_SL g451 ( 
.A1(n_105),
.A2(n_129),
.B1(n_418),
.B2(n_452),
.Y(n_451)
);

AND2x2_ASAP7_75t_L g105 ( 
.A(n_106),
.B(n_118),
.Y(n_105)
);

OAI22xp33_ASAP7_75t_L g106 ( 
.A1(n_107),
.A2(n_110),
.B1(n_113),
.B2(n_116),
.Y(n_106)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx5_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVx6_ASAP7_75t_L g135 ( 
.A(n_109),
.Y(n_135)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_109),
.Y(n_180)
);

INVx2_ASAP7_75t_L g421 ( 
.A(n_109),
.Y(n_421)
);

INVx4_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVx5_ASAP7_75t_L g115 ( 
.A(n_112),
.Y(n_115)
);

INVx4_ASAP7_75t_L g127 ( 
.A(n_112),
.Y(n_127)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx4_ASAP7_75t_L g218 ( 
.A(n_117),
.Y(n_218)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_118),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_SL g214 ( 
.A1(n_118),
.A2(n_215),
.B(n_219),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_119),
.A2(n_122),
.B1(n_124),
.B2(n_126),
.Y(n_118)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_120),
.Y(n_182)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

BUFx5_ASAP7_75t_L g183 ( 
.A(n_123),
.Y(n_183)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_123),
.Y(n_202)
);

BUFx6f_ASAP7_75t_L g281 ( 
.A(n_123),
.Y(n_281)
);

INVx2_ASAP7_75t_L g388 ( 
.A(n_123),
.Y(n_388)
);

BUFx6f_ASAP7_75t_L g390 ( 
.A(n_123),
.Y(n_390)
);

BUFx2_ASAP7_75t_L g322 ( 
.A(n_124),
.Y(n_322)
);

BUFx8_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

BUFx5_ASAP7_75t_L g279 ( 
.A(n_125),
.Y(n_279)
);

INVx2_ASAP7_75t_L g356 ( 
.A(n_125),
.Y(n_356)
);

INVx4_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_SL g374 ( 
.A1(n_128),
.A2(n_219),
.B(n_375),
.Y(n_374)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_129),
.B(n_170),
.Y(n_169)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_130),
.Y(n_452)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

NAND2xp33_ASAP7_75t_SL g294 ( 
.A(n_133),
.B(n_295),
.Y(n_294)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

INVx3_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

XOR2xp5_ASAP7_75t_L g533 ( 
.A(n_136),
.B(n_141),
.Y(n_533)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

AOI21xp5_ASAP7_75t_L g262 ( 
.A1(n_142),
.A2(n_263),
.B(n_272),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_142),
.B(n_314),
.Y(n_313)
);

AOI21xp5_ASAP7_75t_L g475 ( 
.A1(n_142),
.A2(n_272),
.B(n_476),
.Y(n_475)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

INVx3_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

INVx4_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

INVx2_ASAP7_75t_L g414 ( 
.A(n_151),
.Y(n_414)
);

INVxp67_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_SL g154 ( 
.A1(n_155),
.A2(n_530),
.B(n_535),
.Y(n_154)
);

AOI21xp5_ASAP7_75t_SL g155 ( 
.A1(n_156),
.A2(n_502),
.B(n_527),
.Y(n_155)
);

OAI311xp33_ASAP7_75t_L g156 ( 
.A1(n_157),
.A2(n_380),
.A3(n_478),
.B1(n_496),
.C1(n_501),
.Y(n_156)
);

AOI21x1_ASAP7_75t_L g157 ( 
.A1(n_158),
.A2(n_327),
.B(n_379),
.Y(n_157)
);

AO21x1_ASAP7_75t_L g158 ( 
.A1(n_159),
.A2(n_299),
.B(n_326),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_SL g159 ( 
.A1(n_160),
.A2(n_249),
.B(n_298),
.Y(n_159)
);

AOI21xp5_ASAP7_75t_L g160 ( 
.A1(n_161),
.A2(n_222),
.B(n_248),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_162),
.B(n_184),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_162),
.B(n_184),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_163),
.B(n_177),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_163),
.A2(n_177),
.B1(n_178),
.B2(n_246),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_163),
.Y(n_246)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

INVx11_ASAP7_75t_L g172 ( 
.A(n_167),
.Y(n_172)
);

AOI21xp5_ASAP7_75t_L g230 ( 
.A1(n_168),
.A2(n_197),
.B(n_203),
.Y(n_230)
);

OAI21xp33_ASAP7_75t_SL g263 ( 
.A1(n_168),
.A2(n_264),
.B(n_268),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_168),
.B(n_345),
.Y(n_344)
);

OAI21xp33_ASAP7_75t_SL g365 ( 
.A1(n_168),
.A2(n_344),
.B(n_345),
.Y(n_365)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

INVx5_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_181),
.Y(n_178)
);

HB1xp67_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_212),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_185),
.B(n_213),
.C(n_221),
.Y(n_250)
);

AOI21xp5_ASAP7_75t_L g185 ( 
.A1(n_186),
.A2(n_197),
.B(n_203),
.Y(n_185)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_186),
.Y(n_241)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

INVx6_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

BUFx6f_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

INVx5_ASAP7_75t_L g210 ( 
.A(n_191),
.Y(n_210)
);

BUFx6f_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

BUFx6f_ASAP7_75t_L g196 ( 
.A(n_192),
.Y(n_196)
);

BUFx3_ASAP7_75t_L g321 ( 
.A(n_192),
.Y(n_321)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_194),
.Y(n_226)
);

INVx4_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

INVx8_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

INVx4_ASAP7_75t_L g211 ( 
.A(n_196),
.Y(n_211)
);

INVx4_ASAP7_75t_L g392 ( 
.A(n_196),
.Y(n_392)
);

AOI22xp5_ASAP7_75t_L g348 ( 
.A1(n_197),
.A2(n_349),
.B1(n_350),
.B2(n_351),
.Y(n_348)
);

AOI22xp5_ASAP7_75t_L g385 ( 
.A1(n_197),
.A2(n_350),
.B1(n_386),
.B2(n_389),
.Y(n_385)
);

OAI21xp5_ASAP7_75t_SL g422 ( 
.A1(n_197),
.A2(n_389),
.B(n_423),
.Y(n_422)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_198),
.B(n_206),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_198),
.A2(n_240),
.B1(n_241),
.B2(n_242),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g317 ( 
.A1(n_198),
.A2(n_277),
.B1(n_318),
.B2(n_323),
.Y(n_317)
);

OAI22xp5_ASAP7_75t_SL g431 ( 
.A1(n_198),
.A2(n_352),
.B1(n_432),
.B2(n_433),
.Y(n_431)
);

OR2x2_ASAP7_75t_L g198 ( 
.A(n_199),
.B(n_200),
.Y(n_198)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_204),
.B(n_206),
.Y(n_203)
);

INVx4_ASAP7_75t_L g350 ( 
.A(n_204),
.Y(n_350)
);

INVx4_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

INVx3_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_213),
.A2(n_214),
.B1(n_220),
.B2(n_221),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

OAI21xp5_ASAP7_75t_L g222 ( 
.A1(n_223),
.A2(n_238),
.B(n_247),
.Y(n_222)
);

AOI21xp5_ASAP7_75t_L g223 ( 
.A1(n_224),
.A2(n_231),
.B(n_237),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_225),
.B(n_230),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_227),
.Y(n_225)
);

INVx3_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_229),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_232),
.B(n_236),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_232),
.B(n_236),
.Y(n_237)
);

AOI21xp5_ASAP7_75t_L g232 ( 
.A1(n_233),
.A2(n_234),
.B(n_235),
.Y(n_232)
);

INVxp67_ASAP7_75t_L g240 ( 
.A(n_233),
.Y(n_240)
);

AOI21xp5_ASAP7_75t_L g275 ( 
.A1(n_235),
.A2(n_276),
.B(n_282),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_239),
.B(n_245),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_239),
.B(n_245),
.Y(n_247)
);

INVx4_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_250),
.B(n_251),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_250),
.B(n_251),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_252),
.B(n_274),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_253),
.A2(n_254),
.B1(n_261),
.B2(n_262),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_254),
.B(n_261),
.C(n_274),
.Y(n_300)
);

INVx3_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

INVx5_ASAP7_75t_SL g257 ( 
.A(n_258),
.Y(n_257)
);

INVx4_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

INVx4_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

INVx2_ASAP7_75t_L g409 ( 
.A(n_264),
.Y(n_409)
);

INVx4_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

INVx3_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

INVx4_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

INVx2_ASAP7_75t_L g310 ( 
.A(n_267),
.Y(n_310)
);

BUFx6f_ASAP7_75t_L g343 ( 
.A(n_267),
.Y(n_343)
);

INVx3_ASAP7_75t_L g449 ( 
.A(n_267),
.Y(n_449)
);

INVxp33_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

AOI32xp33_ASAP7_75t_L g285 ( 
.A1(n_269),
.A2(n_286),
.A3(n_288),
.B1(n_291),
.B2(n_294),
.Y(n_285)
);

INVx6_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_273),
.Y(n_314)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_275),
.B(n_285),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_275),
.B(n_285),
.Y(n_305)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

INVx3_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

INVx3_ASAP7_75t_SL g282 ( 
.A(n_283),
.Y(n_282)
);

INVx4_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

BUFx6f_ASAP7_75t_L g324 ( 
.A(n_284),
.Y(n_324)
);

INVx8_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

INVx3_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

INVx4_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

INVx5_ASAP7_75t_L g377 ( 
.A(n_290),
.Y(n_377)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

BUFx2_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

INVx2_ASAP7_75t_L g296 ( 
.A(n_297),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_300),
.B(n_301),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_SL g326 ( 
.A(n_300),
.B(n_301),
.Y(n_326)
);

AOI22xp5_ASAP7_75t_L g301 ( 
.A1(n_302),
.A2(n_303),
.B1(n_306),
.B2(n_325),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_303),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_SL g303 ( 
.A(n_304),
.B(n_305),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_304),
.B(n_305),
.C(n_325),
.Y(n_328)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_306),
.Y(n_325)
);

XNOR2xp5_ASAP7_75t_SL g306 ( 
.A(n_307),
.B(n_315),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g359 ( 
.A(n_307),
.B(n_316),
.C(n_317),
.Y(n_359)
);

INVx3_ASAP7_75t_L g309 ( 
.A(n_310),
.Y(n_309)
);

INVx2_ASAP7_75t_L g311 ( 
.A(n_312),
.Y(n_311)
);

XOR2xp5_ASAP7_75t_L g315 ( 
.A(n_316),
.B(n_317),
.Y(n_315)
);

INVxp67_ASAP7_75t_L g349 ( 
.A(n_318),
.Y(n_349)
);

INVx1_ASAP7_75t_SL g319 ( 
.A(n_320),
.Y(n_319)
);

INVx3_ASAP7_75t_L g320 ( 
.A(n_321),
.Y(n_320)
);

INVx2_ASAP7_75t_L g358 ( 
.A(n_321),
.Y(n_358)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_321),
.Y(n_387)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_324),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_328),
.B(n_329),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_SL g379 ( 
.A(n_328),
.B(n_329),
.Y(n_379)
);

XNOR2xp5_ASAP7_75t_L g329 ( 
.A(n_330),
.B(n_362),
.Y(n_329)
);

AOI22xp5_ASAP7_75t_L g330 ( 
.A1(n_331),
.A2(n_359),
.B1(n_360),
.B2(n_361),
.Y(n_330)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_331),
.Y(n_360)
);

OAI22xp5_ASAP7_75t_L g331 ( 
.A1(n_332),
.A2(n_333),
.B1(n_347),
.B2(n_348),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_333),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_333),
.B(n_347),
.Y(n_474)
);

INVx2_ASAP7_75t_L g334 ( 
.A(n_335),
.Y(n_334)
);

INVx3_ASAP7_75t_L g335 ( 
.A(n_336),
.Y(n_335)
);

BUFx2_ASAP7_75t_L g336 ( 
.A(n_337),
.Y(n_336)
);

INVx3_ASAP7_75t_L g338 ( 
.A(n_339),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_341),
.B(n_343),
.Y(n_340)
);

INVx4_ASAP7_75t_L g341 ( 
.A(n_342),
.Y(n_341)
);

INVx6_ASAP7_75t_L g345 ( 
.A(n_346),
.Y(n_345)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_348),
.Y(n_347)
);

INVxp67_ASAP7_75t_L g351 ( 
.A(n_352),
.Y(n_351)
);

BUFx2_ASAP7_75t_L g353 ( 
.A(n_354),
.Y(n_353)
);

INVx2_ASAP7_75t_L g354 ( 
.A(n_355),
.Y(n_354)
);

INVx2_ASAP7_75t_L g355 ( 
.A(n_356),
.Y(n_355)
);

BUFx3_ASAP7_75t_L g357 ( 
.A(n_358),
.Y(n_357)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_359),
.Y(n_361)
);

MAJIxp5_ASAP7_75t_L g492 ( 
.A(n_359),
.B(n_360),
.C(n_362),
.Y(n_492)
);

AOI22xp5_ASAP7_75t_L g362 ( 
.A1(n_363),
.A2(n_364),
.B1(n_369),
.B2(n_378),
.Y(n_362)
);

MAJIxp5_ASAP7_75t_L g487 ( 
.A(n_363),
.B(n_370),
.C(n_374),
.Y(n_487)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_364),
.Y(n_363)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_367),
.Y(n_366)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_369),
.Y(n_378)
);

XNOR2xp5_ASAP7_75t_SL g369 ( 
.A(n_370),
.B(n_374),
.Y(n_369)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_371),
.Y(n_476)
);

INVx6_ASAP7_75t_SL g372 ( 
.A(n_373),
.Y(n_372)
);

BUFx3_ASAP7_75t_L g376 ( 
.A(n_377),
.Y(n_376)
);

NAND2xp33_ASAP7_75t_SL g380 ( 
.A(n_381),
.B(n_464),
.Y(n_380)
);

A2O1A1Ixp33_ASAP7_75t_SL g496 ( 
.A1(n_381),
.A2(n_464),
.B(n_497),
.C(n_500),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_382),
.B(n_439),
.Y(n_381)
);

OR2x2_ASAP7_75t_L g501 ( 
.A(n_382),
.B(n_439),
.Y(n_501)
);

MAJIxp5_ASAP7_75t_L g382 ( 
.A(n_383),
.B(n_415),
.C(n_427),
.Y(n_382)
);

FAx1_ASAP7_75t_SL g477 ( 
.A(n_383),
.B(n_415),
.CI(n_427),
.CON(n_477),
.SN(n_477)
);

XNOR2xp5_ASAP7_75t_L g383 ( 
.A(n_384),
.B(n_401),
.Y(n_383)
);

MAJIxp5_ASAP7_75t_L g440 ( 
.A(n_384),
.B(n_402),
.C(n_410),
.Y(n_440)
);

NOR2xp33_ASAP7_75t_L g384 ( 
.A(n_385),
.B(n_393),
.Y(n_384)
);

XOR2xp5_ASAP7_75t_L g470 ( 
.A(n_385),
.B(n_393),
.Y(n_470)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_386),
.Y(n_432)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_392),
.Y(n_391)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_394),
.Y(n_430)
);

INVx5_ASAP7_75t_L g397 ( 
.A(n_398),
.Y(n_397)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_400),
.Y(n_399)
);

XNOR2xp5_ASAP7_75t_L g401 ( 
.A(n_402),
.B(n_410),
.Y(n_401)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_403),
.Y(n_438)
);

INVx1_ASAP7_75t_SL g404 ( 
.A(n_405),
.Y(n_404)
);

INVx5_ASAP7_75t_L g405 ( 
.A(n_406),
.Y(n_405)
);

INVx3_ASAP7_75t_L g406 ( 
.A(n_407),
.Y(n_406)
);

INVxp67_ASAP7_75t_L g446 ( 
.A(n_408),
.Y(n_446)
);

BUFx6f_ASAP7_75t_L g413 ( 
.A(n_414),
.Y(n_413)
);

OAI22xp5_ASAP7_75t_SL g415 ( 
.A1(n_416),
.A2(n_417),
.B1(n_422),
.B2(n_426),
.Y(n_415)
);

INVxp67_ASAP7_75t_L g416 ( 
.A(n_417),
.Y(n_416)
);

NOR2xp33_ASAP7_75t_L g456 ( 
.A(n_417),
.B(n_422),
.Y(n_456)
);

INVx2_ASAP7_75t_L g419 ( 
.A(n_420),
.Y(n_419)
);

INVx2_ASAP7_75t_L g420 ( 
.A(n_421),
.Y(n_420)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_422),
.Y(n_426)
);

AOI22xp5_ASAP7_75t_L g457 ( 
.A1(n_422),
.A2(n_426),
.B1(n_458),
.B2(n_459),
.Y(n_457)
);

OAI21xp5_ASAP7_75t_L g505 ( 
.A1(n_422),
.A2(n_456),
.B(n_459),
.Y(n_505)
);

INVx2_ASAP7_75t_L g423 ( 
.A(n_424),
.Y(n_423)
);

INVx2_ASAP7_75t_L g424 ( 
.A(n_425),
.Y(n_424)
);

INVx3_ASAP7_75t_L g433 ( 
.A(n_425),
.Y(n_433)
);

MAJIxp5_ASAP7_75t_L g427 ( 
.A(n_428),
.B(n_434),
.C(n_437),
.Y(n_427)
);

XNOR2xp5_ASAP7_75t_L g467 ( 
.A(n_428),
.B(n_468),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_SL g428 ( 
.A(n_429),
.B(n_431),
.Y(n_428)
);

XOR2xp5_ASAP7_75t_L g486 ( 
.A(n_429),
.B(n_431),
.Y(n_486)
);

AOI22xp5_ASAP7_75t_SL g468 ( 
.A1(n_434),
.A2(n_435),
.B1(n_437),
.B2(n_469),
.Y(n_468)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_435),
.Y(n_434)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_437),
.Y(n_469)
);

XNOR2xp5_ASAP7_75t_L g439 ( 
.A(n_440),
.B(n_441),
.Y(n_439)
);

MAJIxp5_ASAP7_75t_L g515 ( 
.A(n_440),
.B(n_443),
.C(n_454),
.Y(n_515)
);

AOI22xp5_ASAP7_75t_L g441 ( 
.A1(n_442),
.A2(n_443),
.B1(n_454),
.B2(n_455),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_443),
.Y(n_442)
);

AOI21xp5_ASAP7_75t_L g443 ( 
.A1(n_444),
.A2(n_450),
.B(n_453),
.Y(n_443)
);

INVxp67_ASAP7_75t_L g444 ( 
.A(n_445),
.Y(n_444)
);

AND2x2_ASAP7_75t_L g453 ( 
.A(n_445),
.B(n_451),
.Y(n_453)
);

INVxp67_ASAP7_75t_L g513 ( 
.A(n_447),
.Y(n_513)
);

INVx2_ASAP7_75t_L g448 ( 
.A(n_449),
.Y(n_448)
);

INVxp67_ASAP7_75t_L g450 ( 
.A(n_451),
.Y(n_450)
);

FAx1_ASAP7_75t_SL g504 ( 
.A(n_453),
.B(n_505),
.CI(n_506),
.CON(n_504),
.SN(n_504)
);

MAJIxp5_ASAP7_75t_L g526 ( 
.A(n_453),
.B(n_505),
.C(n_506),
.Y(n_526)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_455),
.Y(n_454)
);

XNOR2xp5_ASAP7_75t_L g455 ( 
.A(n_456),
.B(n_457),
.Y(n_455)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_459),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_460),
.B(n_463),
.Y(n_459)
);

INVxp67_ASAP7_75t_L g509 ( 
.A(n_461),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_L g464 ( 
.A(n_465),
.B(n_477),
.Y(n_464)
);

NOR2xp33_ASAP7_75t_L g500 ( 
.A(n_465),
.B(n_477),
.Y(n_500)
);

MAJIxp5_ASAP7_75t_L g465 ( 
.A(n_466),
.B(n_470),
.C(n_471),
.Y(n_465)
);

AOI22xp5_ASAP7_75t_SL g489 ( 
.A1(n_466),
.A2(n_467),
.B1(n_470),
.B2(n_490),
.Y(n_489)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_467),
.Y(n_466)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_470),
.Y(n_490)
);

XNOR2xp5_ASAP7_75t_L g488 ( 
.A(n_471),
.B(n_489),
.Y(n_488)
);

MAJIxp5_ASAP7_75t_L g471 ( 
.A(n_472),
.B(n_474),
.C(n_475),
.Y(n_471)
);

OAI22xp5_ASAP7_75t_SL g483 ( 
.A1(n_472),
.A2(n_473),
.B1(n_475),
.B2(n_484),
.Y(n_483)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_473),
.Y(n_472)
);

XOR2xp5_ASAP7_75t_L g482 ( 
.A(n_474),
.B(n_483),
.Y(n_482)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_475),
.Y(n_484)
);

BUFx24_ASAP7_75t_SL g543 ( 
.A(n_477),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_SL g478 ( 
.A(n_479),
.B(n_491),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_480),
.Y(n_479)
);

OAI21xp5_ASAP7_75t_L g497 ( 
.A1(n_480),
.A2(n_498),
.B(n_499),
.Y(n_497)
);

NOR2x1_ASAP7_75t_L g480 ( 
.A(n_481),
.B(n_488),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_L g499 ( 
.A(n_481),
.B(n_488),
.Y(n_499)
);

MAJIxp5_ASAP7_75t_L g481 ( 
.A(n_482),
.B(n_485),
.C(n_487),
.Y(n_481)
);

XOR2xp5_ASAP7_75t_L g493 ( 
.A(n_482),
.B(n_494),
.Y(n_493)
);

AOI22xp5_ASAP7_75t_L g494 ( 
.A1(n_485),
.A2(n_486),
.B1(n_487),
.B2(n_495),
.Y(n_494)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_486),
.Y(n_485)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_487),
.Y(n_495)
);

OR2x2_ASAP7_75t_L g491 ( 
.A(n_492),
.B(n_493),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_L g498 ( 
.A(n_492),
.B(n_493),
.Y(n_498)
);

NOR2xp33_ASAP7_75t_L g502 ( 
.A(n_503),
.B(n_516),
.Y(n_502)
);

NOR2xp33_ASAP7_75t_SL g503 ( 
.A(n_504),
.B(n_515),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_L g528 ( 
.A(n_504),
.B(n_515),
.Y(n_528)
);

BUFx24_ASAP7_75t_SL g544 ( 
.A(n_504),
.Y(n_544)
);

AOI22xp5_ASAP7_75t_L g506 ( 
.A1(n_507),
.A2(n_508),
.B1(n_510),
.B2(n_514),
.Y(n_506)
);

AOI22xp5_ASAP7_75t_L g521 ( 
.A1(n_507),
.A2(n_508),
.B1(n_522),
.B2(n_523),
.Y(n_521)
);

MAJIxp5_ASAP7_75t_L g534 ( 
.A(n_507),
.B(n_518),
.C(n_522),
.Y(n_534)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_508),
.Y(n_507)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_510),
.Y(n_514)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_512),
.Y(n_511)
);

OAI21xp5_ASAP7_75t_L g527 ( 
.A1(n_516),
.A2(n_528),
.B(n_529),
.Y(n_527)
);

NOR2xp33_ASAP7_75t_SL g516 ( 
.A(n_517),
.B(n_526),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_L g529 ( 
.A(n_517),
.B(n_526),
.Y(n_529)
);

OAI22xp5_ASAP7_75t_L g517 ( 
.A1(n_518),
.A2(n_519),
.B1(n_520),
.B2(n_521),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_519),
.Y(n_518)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_521),
.Y(n_520)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_523),
.Y(n_522)
);

NOR2xp33_ASAP7_75t_L g530 ( 
.A(n_531),
.B(n_534),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_L g535 ( 
.A(n_531),
.B(n_534),
.Y(n_535)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_533),
.Y(n_532)
);

BUFx6f_ASAP7_75t_L g536 ( 
.A(n_537),
.Y(n_536)
);

BUFx6f_ASAP7_75t_L g540 ( 
.A(n_537),
.Y(n_540)
);

INVx13_ASAP7_75t_L g537 ( 
.A(n_538),
.Y(n_537)
);

NOR2xp33_ASAP7_75t_L g539 ( 
.A(n_540),
.B(n_541),
.Y(n_539)
);


endmodule