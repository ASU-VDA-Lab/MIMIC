module fake_aes_5933_n_512 (n_53, n_67, n_45, n_20, n_2, n_38, n_44, n_64, n_54, n_62, n_36, n_47, n_37, n_69, n_34, n_5, n_23, n_8, n_28, n_31, n_22, n_46, n_48, n_58, n_57, n_11, n_25, n_16, n_26, n_13, n_30, n_33, n_50, n_52, n_49, n_59, n_73, n_3, n_18, n_60, n_66, n_32, n_0, n_41, n_1, n_35, n_55, n_65, n_12, n_9, n_70, n_17, n_63, n_14, n_10, n_15, n_56, n_71, n_42, n_24, n_19, n_61, n_21, n_6, n_4, n_74, n_72, n_51, n_29, n_43, n_7, n_68, n_40, n_27, n_39, n_512, n_221);
input n_53;
input n_67;
input n_45;
input n_20;
input n_2;
input n_38;
input n_44;
input n_64;
input n_54;
input n_62;
input n_36;
input n_47;
input n_37;
input n_69;
input n_34;
input n_5;
input n_23;
input n_8;
input n_28;
input n_31;
input n_22;
input n_46;
input n_48;
input n_58;
input n_57;
input n_11;
input n_25;
input n_16;
input n_26;
input n_13;
input n_30;
input n_33;
input n_50;
input n_52;
input n_49;
input n_59;
input n_73;
input n_3;
input n_18;
input n_60;
input n_66;
input n_32;
input n_0;
input n_41;
input n_1;
input n_35;
input n_55;
input n_65;
input n_12;
input n_9;
input n_70;
input n_17;
input n_63;
input n_14;
input n_10;
input n_15;
input n_56;
input n_71;
input n_42;
input n_24;
input n_19;
input n_61;
input n_21;
input n_6;
input n_4;
input n_74;
input n_72;
input n_51;
input n_29;
input n_43;
input n_7;
input n_68;
input n_40;
input n_27;
input n_39;
output n_512;
output n_221;
wire n_117;
wire n_361;
wire n_185;
wire n_407;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_154;
wire n_328;
wire n_468;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_353;
wire n_206;
wire n_288;
wire n_383;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_462;
wire n_316;
wire n_211;
wire n_334;
wire n_389;
wire n_436;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_231;
wire n_452;
wire n_298;
wire n_411;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_366;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_324;
wire n_392;
wire n_279;
wire n_303;
wire n_437;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_244;
wire n_119;
wire n_141;
wire n_479;
wire n_97;
wire n_167;
wire n_447;
wire n_171;
wire n_196;
wire n_192;
wire n_502;
wire n_312;
wire n_455;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_367;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_293;
wire n_506;
wire n_393;
wire n_135;
wire n_247;
wire n_490;
wire n_381;
wire n_304;
wire n_399;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_307;
wire n_191;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_256;
wire n_77;
wire n_404;
wire n_369;
wire n_509;
wire n_172;
wire n_329;
wire n_251;
wire n_218;
wire n_507;
wire n_271;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_133;
wire n_149;
wire n_81;
wire n_214;
wire n_204;
wire n_430;
wire n_88;
wire n_450;
wire n_107;
wire n_403;
wire n_254;
wire n_262;
wire n_239;
wire n_439;
wire n_87;
wire n_379;
wire n_98;
wire n_276;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_446;
wire n_342;
wire n_423;
wire n_370;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_486;
wire n_245;
wire n_90;
wire n_357;
wire n_260;
wire n_78;
wire n_201;
wire n_197;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_265;
wire n_264;
wire n_200;
wire n_208;
wire n_126;
wire n_178;
wire n_118;
wire n_365;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_295;
wire n_143;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_75;
wire n_376;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_76;
wire n_435;
wire n_216;
wire n_147;
wire n_148;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_398;
wire n_445;
wire n_438;
wire n_134;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_225;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_121;
wire n_497;
wire n_339;
wire n_240;
wire n_378;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_335;
wire n_272;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_198;
wire n_169;
wire n_424;
wire n_156;
wire n_124;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_418;
wire n_493;
wire n_380;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_258;
wire n_253;
wire n_84;
wire n_266;
wire n_213;
wire n_182;
wire n_492;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_444;
wire n_176;
wire n_469;
wire n_123;
wire n_457;
wire n_223;
wire n_494;
wire n_480;
wire n_372;
wire n_453;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_425;
wire n_332;
wire n_414;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_132;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
CKINVDCx20_ASAP7_75t_R g75 ( .A(n_71), .Y(n_75) );
INVx2_ASAP7_75t_L g76 ( .A(n_16), .Y(n_76) );
INVx1_ASAP7_75t_L g77 ( .A(n_14), .Y(n_77) );
INVx1_ASAP7_75t_L g78 ( .A(n_39), .Y(n_78) );
INVx1_ASAP7_75t_L g79 ( .A(n_17), .Y(n_79) );
INVx1_ASAP7_75t_L g80 ( .A(n_66), .Y(n_80) );
INVxp33_ASAP7_75t_SL g81 ( .A(n_5), .Y(n_81) );
CKINVDCx5p33_ASAP7_75t_R g82 ( .A(n_53), .Y(n_82) );
INVx1_ASAP7_75t_L g83 ( .A(n_63), .Y(n_83) );
INVx1_ASAP7_75t_L g84 ( .A(n_29), .Y(n_84) );
INVxp67_ASAP7_75t_SL g85 ( .A(n_11), .Y(n_85) );
INVxp67_ASAP7_75t_L g86 ( .A(n_15), .Y(n_86) );
INVx1_ASAP7_75t_L g87 ( .A(n_45), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_24), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_27), .Y(n_89) );
INVx1_ASAP7_75t_L g90 ( .A(n_32), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_42), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_16), .Y(n_92) );
INVx1_ASAP7_75t_L g93 ( .A(n_56), .Y(n_93) );
INVxp67_ASAP7_75t_L g94 ( .A(n_18), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_69), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_57), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_43), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_15), .Y(n_98) );
INVxp33_ASAP7_75t_SL g99 ( .A(n_54), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_21), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_40), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_12), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_19), .Y(n_103) );
INVxp67_ASAP7_75t_SL g104 ( .A(n_30), .Y(n_104) );
CKINVDCx14_ASAP7_75t_R g105 ( .A(n_9), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_6), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_4), .Y(n_107) );
BUFx6f_ASAP7_75t_L g108 ( .A(n_23), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_31), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_14), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_70), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_79), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_79), .Y(n_113) );
INVx2_ASAP7_75t_L g114 ( .A(n_80), .Y(n_114) );
CKINVDCx5p33_ASAP7_75t_R g115 ( .A(n_105), .Y(n_115) );
NAND2xp5_ASAP7_75t_L g116 ( .A(n_86), .B(n_0), .Y(n_116) );
INVx2_ASAP7_75t_L g117 ( .A(n_108), .Y(n_117) );
INVx2_ASAP7_75t_L g118 ( .A(n_108), .Y(n_118) );
INVx2_ASAP7_75t_L g119 ( .A(n_108), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_80), .Y(n_120) );
CKINVDCx5p33_ASAP7_75t_R g121 ( .A(n_105), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_83), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_83), .Y(n_123) );
CKINVDCx5p33_ASAP7_75t_R g124 ( .A(n_75), .Y(n_124) );
HB1xp67_ASAP7_75t_L g125 ( .A(n_76), .Y(n_125) );
INVx2_ASAP7_75t_SL g126 ( .A(n_84), .Y(n_126) );
CKINVDCx5p33_ASAP7_75t_R g127 ( .A(n_75), .Y(n_127) );
BUFx6f_ASAP7_75t_L g128 ( .A(n_108), .Y(n_128) );
CKINVDCx5p33_ASAP7_75t_R g129 ( .A(n_82), .Y(n_129) );
CKINVDCx5p33_ASAP7_75t_R g130 ( .A(n_82), .Y(n_130) );
CKINVDCx20_ASAP7_75t_R g131 ( .A(n_77), .Y(n_131) );
CKINVDCx5p33_ASAP7_75t_R g132 ( .A(n_99), .Y(n_132) );
INVx2_ASAP7_75t_SL g133 ( .A(n_112), .Y(n_133) );
INVx2_ASAP7_75t_L g134 ( .A(n_128), .Y(n_134) );
BUFx6f_ASAP7_75t_L g135 ( .A(n_128), .Y(n_135) );
NAND2xp5_ASAP7_75t_SL g136 ( .A(n_115), .B(n_94), .Y(n_136) );
OR2x2_ASAP7_75t_L g137 ( .A(n_125), .B(n_85), .Y(n_137) );
INVx2_ASAP7_75t_SL g138 ( .A(n_112), .Y(n_138) );
INVx3_ASAP7_75t_L g139 ( .A(n_114), .Y(n_139) );
INVx2_ASAP7_75t_L g140 ( .A(n_128), .Y(n_140) );
OR2x6_ASAP7_75t_L g141 ( .A(n_116), .B(n_76), .Y(n_141) );
INVxp67_ASAP7_75t_L g142 ( .A(n_129), .Y(n_142) );
INVx4_ASAP7_75t_SL g143 ( .A(n_128), .Y(n_143) );
INVx3_ASAP7_75t_L g144 ( .A(n_114), .Y(n_144) );
AND2x4_ASAP7_75t_L g145 ( .A(n_126), .B(n_92), .Y(n_145) );
BUFx3_ASAP7_75t_L g146 ( .A(n_126), .Y(n_146) );
AND2x4_ASAP7_75t_L g147 ( .A(n_113), .B(n_98), .Y(n_147) );
INVx1_ASAP7_75t_L g148 ( .A(n_113), .Y(n_148) );
INVx1_ASAP7_75t_L g149 ( .A(n_120), .Y(n_149) );
INVx1_ASAP7_75t_L g150 ( .A(n_120), .Y(n_150) );
INVx2_ASAP7_75t_L g151 ( .A(n_128), .Y(n_151) );
INVx1_ASAP7_75t_L g152 ( .A(n_122), .Y(n_152) );
INVx3_ASAP7_75t_R g153 ( .A(n_117), .Y(n_153) );
INVxp67_ASAP7_75t_L g154 ( .A(n_130), .Y(n_154) );
NAND2xp5_ASAP7_75t_L g155 ( .A(n_122), .B(n_78), .Y(n_155) );
AOI22xp33_ASAP7_75t_L g156 ( .A1(n_141), .A2(n_123), .B1(n_81), .B2(n_99), .Y(n_156) );
BUFx2_ASAP7_75t_L g157 ( .A(n_141), .Y(n_157) );
INVxp67_ASAP7_75t_SL g158 ( .A(n_133), .Y(n_158) );
INVx2_ASAP7_75t_L g159 ( .A(n_139), .Y(n_159) );
AND2x6_ASAP7_75t_L g160 ( .A(n_145), .B(n_84), .Y(n_160) );
NOR2xp67_ASAP7_75t_L g161 ( .A(n_139), .B(n_123), .Y(n_161) );
INVx1_ASAP7_75t_L g162 ( .A(n_148), .Y(n_162) );
NOR2xp33_ASAP7_75t_L g163 ( .A(n_136), .B(n_132), .Y(n_163) );
BUFx3_ASAP7_75t_L g164 ( .A(n_146), .Y(n_164) );
INVx2_ASAP7_75t_L g165 ( .A(n_139), .Y(n_165) );
INVx2_ASAP7_75t_L g166 ( .A(n_139), .Y(n_166) );
BUFx6f_ASAP7_75t_L g167 ( .A(n_133), .Y(n_167) );
INVx2_ASAP7_75t_L g168 ( .A(n_144), .Y(n_168) );
BUFx2_ASAP7_75t_L g169 ( .A(n_141), .Y(n_169) );
NOR2xp33_ASAP7_75t_SL g170 ( .A(n_133), .B(n_104), .Y(n_170) );
INVx2_ASAP7_75t_SL g171 ( .A(n_141), .Y(n_171) );
INVx3_ASAP7_75t_L g172 ( .A(n_144), .Y(n_172) );
INVx1_ASAP7_75t_L g173 ( .A(n_148), .Y(n_173) );
AND2x4_ASAP7_75t_SL g174 ( .A(n_141), .B(n_147), .Y(n_174) );
OR2x6_ASAP7_75t_L g175 ( .A(n_142), .B(n_154), .Y(n_175) );
NAND2xp5_ASAP7_75t_L g176 ( .A(n_145), .B(n_121), .Y(n_176) );
INVxp67_ASAP7_75t_L g177 ( .A(n_142), .Y(n_177) );
NAND2xp5_ASAP7_75t_L g178 ( .A(n_145), .B(n_111), .Y(n_178) );
NAND2xp33_ASAP7_75t_R g179 ( .A(n_137), .B(n_124), .Y(n_179) );
BUFx4f_ASAP7_75t_L g180 ( .A(n_149), .Y(n_180) );
NOR2xp33_ASAP7_75t_R g181 ( .A(n_154), .B(n_127), .Y(n_181) );
AND2x2_ASAP7_75t_L g182 ( .A(n_147), .B(n_102), .Y(n_182) );
INVx1_ASAP7_75t_L g183 ( .A(n_149), .Y(n_183) );
NAND2x1p5_ASAP7_75t_L g184 ( .A(n_150), .B(n_111), .Y(n_184) );
BUFx3_ASAP7_75t_L g185 ( .A(n_146), .Y(n_185) );
NOR2xp33_ASAP7_75t_L g186 ( .A(n_176), .B(n_145), .Y(n_186) );
AND2x4_ASAP7_75t_L g187 ( .A(n_174), .B(n_147), .Y(n_187) );
BUFx6f_ASAP7_75t_L g188 ( .A(n_167), .Y(n_188) );
OR2x2_ASAP7_75t_L g189 ( .A(n_175), .B(n_137), .Y(n_189) );
INVx2_ASAP7_75t_L g190 ( .A(n_162), .Y(n_190) );
AOI21x1_ASAP7_75t_SL g191 ( .A1(n_178), .A2(n_155), .B(n_147), .Y(n_191) );
CKINVDCx5p33_ASAP7_75t_R g192 ( .A(n_181), .Y(n_192) );
INVx1_ASAP7_75t_L g193 ( .A(n_162), .Y(n_193) );
NOR2xp33_ASAP7_75t_L g194 ( .A(n_177), .B(n_131), .Y(n_194) );
AOI22xp33_ASAP7_75t_L g195 ( .A1(n_160), .A2(n_152), .B1(n_150), .B2(n_138), .Y(n_195) );
A2O1A1Ixp33_ASAP7_75t_L g196 ( .A1(n_173), .A2(n_152), .B(n_138), .C(n_155), .Y(n_196) );
INVx3_ASAP7_75t_L g197 ( .A(n_180), .Y(n_197) );
INVx1_ASAP7_75t_L g198 ( .A(n_173), .Y(n_198) );
AND2x4_ASAP7_75t_L g199 ( .A(n_174), .B(n_146), .Y(n_199) );
AOI22xp33_ASAP7_75t_L g200 ( .A1(n_160), .A2(n_138), .B1(n_144), .B2(n_81), .Y(n_200) );
BUFx3_ASAP7_75t_L g201 ( .A(n_180), .Y(n_201) );
HB1xp67_ASAP7_75t_L g202 ( .A(n_174), .Y(n_202) );
INVx4_ASAP7_75t_L g203 ( .A(n_180), .Y(n_203) );
INVx2_ASAP7_75t_L g204 ( .A(n_183), .Y(n_204) );
INVx3_ASAP7_75t_L g205 ( .A(n_180), .Y(n_205) );
BUFx3_ASAP7_75t_L g206 ( .A(n_164), .Y(n_206) );
BUFx6f_ASAP7_75t_L g207 ( .A(n_167), .Y(n_207) );
INVx2_ASAP7_75t_L g208 ( .A(n_183), .Y(n_208) );
A2O1A1Ixp33_ASAP7_75t_L g209 ( .A1(n_161), .A2(n_144), .B(n_106), .C(n_107), .Y(n_209) );
INVx2_ASAP7_75t_L g210 ( .A(n_167), .Y(n_210) );
AOI21xp5_ASAP7_75t_L g211 ( .A1(n_158), .A2(n_87), .B(n_90), .Y(n_211) );
BUFx12f_ASAP7_75t_L g212 ( .A(n_175), .Y(n_212) );
INVx2_ASAP7_75t_L g213 ( .A(n_167), .Y(n_213) );
INVx2_ASAP7_75t_L g214 ( .A(n_167), .Y(n_214) );
INVx1_ASAP7_75t_L g215 ( .A(n_159), .Y(n_215) );
OAI22xp33_ASAP7_75t_L g216 ( .A1(n_212), .A2(n_175), .B1(n_179), .B2(n_169), .Y(n_216) );
AOI221xp5_ASAP7_75t_L g217 ( .A1(n_194), .A2(n_156), .B1(n_182), .B2(n_163), .C(n_169), .Y(n_217) );
AOI22xp33_ASAP7_75t_SL g218 ( .A1(n_212), .A2(n_175), .B1(n_157), .B2(n_171), .Y(n_218) );
AOI22xp33_ASAP7_75t_L g219 ( .A1(n_189), .A2(n_157), .B1(n_160), .B2(n_171), .Y(n_219) );
AOI22xp33_ASAP7_75t_L g220 ( .A1(n_189), .A2(n_160), .B1(n_175), .B2(n_182), .Y(n_220) );
UNKNOWN g221 ( );
OAI22xp33_ASAP7_75t_L g222 ( .A1(n_212), .A2(n_184), .B1(n_170), .B2(n_161), .Y(n_222) );
A2O1A1Ixp33_ASAP7_75t_L g223 ( .A1(n_186), .A2(n_172), .B(n_159), .C(n_168), .Y(n_223) );
AOI22xp33_ASAP7_75t_L g224 ( .A1(n_187), .A2(n_160), .B1(n_184), .B2(n_172), .Y(n_224) );
OAI21xp5_ASAP7_75t_L g225 ( .A1(n_196), .A2(n_184), .B(n_159), .Y(n_225) );
CKINVDCx8_ASAP7_75t_R g226 ( .A(n_192), .Y(n_226) );
INVx2_ASAP7_75t_L g227 ( .A(n_190), .Y(n_227) );
CKINVDCx11_ASAP7_75t_R g228 ( .A(n_187), .Y(n_228) );
OAI22xp33_ASAP7_75t_L g229 ( .A1(n_203), .A2(n_170), .B1(n_164), .B2(n_185), .Y(n_229) );
NAND3xp33_ASAP7_75t_L g230 ( .A(n_186), .B(n_209), .C(n_200), .Y(n_230) );
AND2x2_ASAP7_75t_L g231 ( .A(n_190), .B(n_172), .Y(n_231) );
CKINVDCx14_ASAP7_75t_R g232 ( .A(n_187), .Y(n_232) );
AOI22xp33_ASAP7_75t_L g233 ( .A1(n_187), .A2(n_160), .B1(n_172), .B2(n_185), .Y(n_233) );
INVx1_ASAP7_75t_L g234 ( .A(n_193), .Y(n_234) );
AOI221xp5_ASAP7_75t_L g235 ( .A1(n_193), .A2(n_110), .B1(n_168), .B2(n_165), .C(n_166), .Y(n_235) );
OR2x2_ASAP7_75t_L g236 ( .A(n_190), .B(n_165), .Y(n_236) );
AOI221xp5_ASAP7_75t_L g237 ( .A1(n_198), .A2(n_165), .B1(n_168), .B2(n_166), .C(n_89), .Y(n_237) );
AOI21xp5_ASAP7_75t_L g238 ( .A1(n_198), .A2(n_167), .B(n_185), .Y(n_238) );
NAND2xp5_ASAP7_75t_L g239 ( .A(n_204), .B(n_160), .Y(n_239) );
INVx2_ASAP7_75t_L g240 ( .A(n_204), .Y(n_240) );
INVx1_ASAP7_75t_L g241 ( .A(n_227), .Y(n_241) );
AO21x1_ASAP7_75t_L g242 ( .A1(n_225), .A2(n_204), .B(n_208), .Y(n_242) );
BUFx6f_ASAP7_75t_L g243 ( .A(n_227), .Y(n_243) );
OAI221xp5_ASAP7_75t_SL g244 ( .A1(n_217), .A2(n_195), .B1(n_211), .B2(n_208), .C(n_93), .Y(n_244) );
AOI221xp5_ASAP7_75t_L g245 ( .A1(n_230), .A2(n_211), .B1(n_208), .B2(n_202), .C(n_215), .Y(n_245) );
OAI211xp5_ASAP7_75t_L g246 ( .A1(n_220), .A2(n_195), .B(n_202), .C(n_95), .Y(n_246) );
AND2x4_ASAP7_75t_L g247 ( .A(n_234), .B(n_203), .Y(n_247) );
INVx1_ASAP7_75t_L g248 ( .A(n_240), .Y(n_248) );
INVx1_ASAP7_75t_L g249 ( .A(n_240), .Y(n_249) );
INVx2_ASAP7_75t_L g250 ( .A(n_236), .Y(n_250) );
OAI22xp5_ASAP7_75t_L g251 ( .A1(n_224), .A2(n_203), .B1(n_199), .B2(n_201), .Y(n_251) );
AND2x2_ASAP7_75t_L g252 ( .A(n_234), .B(n_215), .Y(n_252) );
AOI22xp33_ASAP7_75t_SL g253 ( .A1(n_232), .A2(n_203), .B1(n_160), .B2(n_201), .Y(n_253) );
INVx1_ASAP7_75t_L g254 ( .A(n_236), .Y(n_254) );
AO21x2_ASAP7_75t_L g255 ( .A1(n_223), .A2(n_214), .B(n_213), .Y(n_255) );
INVx1_ASAP7_75t_L g256 ( .A(n_231), .Y(n_256) );
AOI22xp33_ASAP7_75t_L g257 ( .A1(n_221), .A2(n_199), .B1(n_197), .B2(n_205), .Y(n_257) );
AOI22xp33_ASAP7_75t_L g258 ( .A1(n_216), .A2(n_199), .B1(n_197), .B2(n_205), .Y(n_258) );
OAI21xp5_ASAP7_75t_L g259 ( .A1(n_238), .A2(n_214), .B(n_213), .Y(n_259) );
BUFx3_ASAP7_75t_L g260 ( .A(n_228), .Y(n_260) );
INVx1_ASAP7_75t_L g261 ( .A(n_231), .Y(n_261) );
AO21x2_ASAP7_75t_L g262 ( .A1(n_242), .A2(n_222), .B(n_229), .Y(n_262) );
INVx1_ASAP7_75t_L g263 ( .A(n_241), .Y(n_263) );
AOI22xp33_ASAP7_75t_L g264 ( .A1(n_260), .A2(n_228), .B1(n_218), .B2(n_235), .Y(n_264) );
AO21x2_ASAP7_75t_L g265 ( .A1(n_242), .A2(n_239), .B(n_88), .Y(n_265) );
INVxp67_ASAP7_75t_L g266 ( .A(n_252), .Y(n_266) );
INVx2_ASAP7_75t_SL g267 ( .A(n_250), .Y(n_267) );
HB1xp67_ASAP7_75t_L g268 ( .A(n_243), .Y(n_268) );
BUFx2_ASAP7_75t_L g269 ( .A(n_250), .Y(n_269) );
AND2x6_ASAP7_75t_SL g270 ( .A(n_260), .B(n_226), .Y(n_270) );
OAI221xp5_ASAP7_75t_L g271 ( .A1(n_244), .A2(n_219), .B1(n_233), .B2(n_237), .C(n_226), .Y(n_271) );
INVx3_ASAP7_75t_L g272 ( .A(n_243), .Y(n_272) );
AOI22xp5_ASAP7_75t_L g273 ( .A1(n_257), .A2(n_199), .B1(n_197), .B2(n_205), .Y(n_273) );
OAI33xp33_ASAP7_75t_L g274 ( .A1(n_254), .A2(n_91), .A3(n_96), .B1(n_97), .B2(n_100), .B3(n_101), .Y(n_274) );
AO21x2_ASAP7_75t_L g275 ( .A1(n_259), .A2(n_103), .B(n_109), .Y(n_275) );
INVxp67_ASAP7_75t_SL g276 ( .A(n_250), .Y(n_276) );
INVx2_ASAP7_75t_L g277 ( .A(n_243), .Y(n_277) );
INVx1_ASAP7_75t_L g278 ( .A(n_241), .Y(n_278) );
INVx1_ASAP7_75t_L g279 ( .A(n_248), .Y(n_279) );
INVx2_ASAP7_75t_L g280 ( .A(n_243), .Y(n_280) );
INVxp67_ASAP7_75t_L g281 ( .A(n_252), .Y(n_281) );
INVx1_ASAP7_75t_L g282 ( .A(n_263), .Y(n_282) );
NAND2xp5_ASAP7_75t_L g283 ( .A(n_266), .B(n_254), .Y(n_283) );
INVx4_ASAP7_75t_L g284 ( .A(n_270), .Y(n_284) );
NOR3xp33_ASAP7_75t_L g285 ( .A(n_274), .B(n_246), .C(n_260), .Y(n_285) );
OR2x2_ASAP7_75t_L g286 ( .A(n_269), .B(n_248), .Y(n_286) );
OR2x2_ASAP7_75t_L g287 ( .A(n_269), .B(n_249), .Y(n_287) );
INVx2_ASAP7_75t_L g288 ( .A(n_263), .Y(n_288) );
AOI33xp33_ASAP7_75t_L g289 ( .A1(n_264), .A2(n_258), .A3(n_261), .B1(n_256), .B2(n_253), .B3(n_117), .Y(n_289) );
NAND2xp5_ASAP7_75t_L g290 ( .A(n_266), .B(n_261), .Y(n_290) );
INVx1_ASAP7_75t_L g291 ( .A(n_278), .Y(n_291) );
OR2x2_ASAP7_75t_L g292 ( .A(n_267), .B(n_249), .Y(n_292) );
INVx1_ASAP7_75t_L g293 ( .A(n_278), .Y(n_293) );
AND2x2_ASAP7_75t_L g294 ( .A(n_267), .B(n_243), .Y(n_294) );
INVx1_ASAP7_75t_L g295 ( .A(n_279), .Y(n_295) );
HB1xp67_ASAP7_75t_L g296 ( .A(n_267), .Y(n_296) );
AND2x2_ASAP7_75t_L g297 ( .A(n_276), .B(n_243), .Y(n_297) );
INVx1_ASAP7_75t_L g298 ( .A(n_279), .Y(n_298) );
INVx1_ASAP7_75t_L g299 ( .A(n_281), .Y(n_299) );
INVx1_ASAP7_75t_L g300 ( .A(n_281), .Y(n_300) );
INVx1_ASAP7_75t_L g301 ( .A(n_276), .Y(n_301) );
AND2x2_ASAP7_75t_L g302 ( .A(n_268), .B(n_256), .Y(n_302) );
AND2x4_ASAP7_75t_L g303 ( .A(n_272), .B(n_255), .Y(n_303) );
AOI21xp5_ASAP7_75t_L g304 ( .A1(n_268), .A2(n_259), .B(n_245), .Y(n_304) );
INVx2_ASAP7_75t_L g305 ( .A(n_277), .Y(n_305) );
NAND2x1p5_ASAP7_75t_L g306 ( .A(n_272), .B(n_247), .Y(n_306) );
INVx1_ASAP7_75t_L g307 ( .A(n_277), .Y(n_307) );
HB1xp67_ASAP7_75t_L g308 ( .A(n_280), .Y(n_308) );
AND2x2_ASAP7_75t_L g309 ( .A(n_265), .B(n_247), .Y(n_309) );
INVx1_ASAP7_75t_L g310 ( .A(n_282), .Y(n_310) );
OAI21xp33_ASAP7_75t_SL g311 ( .A1(n_292), .A2(n_273), .B(n_264), .Y(n_311) );
AOI22xp33_ASAP7_75t_L g312 ( .A1(n_285), .A2(n_271), .B1(n_274), .B2(n_273), .Y(n_312) );
INVx1_ASAP7_75t_L g313 ( .A(n_282), .Y(n_313) );
AND2x2_ASAP7_75t_L g314 ( .A(n_309), .B(n_262), .Y(n_314) );
NAND3xp33_ASAP7_75t_L g315 ( .A(n_289), .B(n_108), .C(n_128), .Y(n_315) );
AOI22xp33_ASAP7_75t_L g316 ( .A1(n_284), .A2(n_271), .B1(n_247), .B2(n_262), .Y(n_316) );
AND2x2_ASAP7_75t_L g317 ( .A(n_309), .B(n_262), .Y(n_317) );
HB1xp67_ASAP7_75t_L g318 ( .A(n_296), .Y(n_318) );
INVx1_ASAP7_75t_L g319 ( .A(n_291), .Y(n_319) );
AND2x4_ASAP7_75t_SL g320 ( .A(n_284), .B(n_247), .Y(n_320) );
NAND2xp5_ASAP7_75t_L g321 ( .A(n_299), .B(n_275), .Y(n_321) );
AND2x2_ASAP7_75t_L g322 ( .A(n_297), .B(n_262), .Y(n_322) );
INVx1_ASAP7_75t_L g323 ( .A(n_291), .Y(n_323) );
INVx1_ASAP7_75t_L g324 ( .A(n_293), .Y(n_324) );
INVx1_ASAP7_75t_L g325 ( .A(n_293), .Y(n_325) );
INVx3_ASAP7_75t_L g326 ( .A(n_303), .Y(n_326) );
INVx1_ASAP7_75t_L g327 ( .A(n_295), .Y(n_327) );
OR2x2_ASAP7_75t_L g328 ( .A(n_286), .B(n_275), .Y(n_328) );
INVx1_ASAP7_75t_L g329 ( .A(n_295), .Y(n_329) );
NAND2xp5_ASAP7_75t_L g330 ( .A(n_300), .B(n_275), .Y(n_330) );
AND2x2_ASAP7_75t_L g331 ( .A(n_297), .B(n_288), .Y(n_331) );
OR2x2_ASAP7_75t_L g332 ( .A(n_286), .B(n_287), .Y(n_332) );
INVx1_ASAP7_75t_SL g333 ( .A(n_287), .Y(n_333) );
OAI21xp5_ASAP7_75t_SL g334 ( .A1(n_306), .A2(n_270), .B(n_251), .Y(n_334) );
NAND2xp5_ASAP7_75t_L g335 ( .A(n_283), .B(n_275), .Y(n_335) );
INVx1_ASAP7_75t_L g336 ( .A(n_288), .Y(n_336) );
HB1xp67_ASAP7_75t_L g337 ( .A(n_292), .Y(n_337) );
AND2x2_ASAP7_75t_L g338 ( .A(n_294), .B(n_265), .Y(n_338) );
HB1xp67_ASAP7_75t_L g339 ( .A(n_301), .Y(n_339) );
BUFx3_ASAP7_75t_L g340 ( .A(n_306), .Y(n_340) );
INVx1_ASAP7_75t_L g341 ( .A(n_298), .Y(n_341) );
AND4x1_ASAP7_75t_L g342 ( .A(n_284), .B(n_0), .C(n_1), .D(n_2), .Y(n_342) );
AND2x2_ASAP7_75t_L g343 ( .A(n_294), .B(n_265), .Y(n_343) );
NAND2xp33_ASAP7_75t_L g344 ( .A(n_301), .B(n_272), .Y(n_344) );
BUFx2_ASAP7_75t_L g345 ( .A(n_308), .Y(n_345) );
INVx1_ASAP7_75t_SL g346 ( .A(n_306), .Y(n_346) );
INVx1_ASAP7_75t_L g347 ( .A(n_307), .Y(n_347) );
INVx2_ASAP7_75t_L g348 ( .A(n_305), .Y(n_348) );
INVxp67_ASAP7_75t_L g349 ( .A(n_290), .Y(n_349) );
AND2x2_ASAP7_75t_L g350 ( .A(n_307), .B(n_265), .Y(n_350) );
AND2x2_ASAP7_75t_L g351 ( .A(n_305), .B(n_277), .Y(n_351) );
INVxp67_ASAP7_75t_L g352 ( .A(n_318), .Y(n_352) );
NAND2xp5_ASAP7_75t_L g353 ( .A(n_349), .B(n_302), .Y(n_353) );
AND2x4_ASAP7_75t_SL g354 ( .A(n_337), .B(n_302), .Y(n_354) );
AOI22xp33_ASAP7_75t_SL g355 ( .A1(n_311), .A2(n_303), .B1(n_272), .B2(n_304), .Y(n_355) );
AOI21xp33_ASAP7_75t_L g356 ( .A1(n_311), .A2(n_334), .B(n_330), .Y(n_356) );
AND2x2_ASAP7_75t_L g357 ( .A(n_333), .B(n_303), .Y(n_357) );
OR2x2_ASAP7_75t_L g358 ( .A(n_332), .B(n_280), .Y(n_358) );
OAI21xp5_ASAP7_75t_L g359 ( .A1(n_315), .A2(n_117), .B(n_118), .Y(n_359) );
NAND2xp5_ASAP7_75t_L g360 ( .A(n_332), .B(n_272), .Y(n_360) );
INVx2_ASAP7_75t_L g361 ( .A(n_345), .Y(n_361) );
INVx1_ASAP7_75t_SL g362 ( .A(n_320), .Y(n_362) );
AND2x2_ASAP7_75t_L g363 ( .A(n_331), .B(n_280), .Y(n_363) );
INVx1_ASAP7_75t_L g364 ( .A(n_310), .Y(n_364) );
NAND2xp5_ASAP7_75t_L g365 ( .A(n_331), .B(n_255), .Y(n_365) );
AND2x4_ASAP7_75t_L g366 ( .A(n_326), .B(n_255), .Y(n_366) );
INVx2_ASAP7_75t_SL g367 ( .A(n_320), .Y(n_367) );
AOI22xp5_ASAP7_75t_L g368 ( .A1(n_312), .A2(n_255), .B1(n_197), .B2(n_205), .Y(n_368) );
AOI21xp5_ASAP7_75t_L g369 ( .A1(n_315), .A2(n_214), .B(n_213), .Y(n_369) );
INVx2_ASAP7_75t_L g370 ( .A(n_345), .Y(n_370) );
INVx1_ASAP7_75t_L g371 ( .A(n_310), .Y(n_371) );
AOI222xp33_ASAP7_75t_L g372 ( .A1(n_314), .A2(n_118), .B1(n_119), .B2(n_3), .C1(n_4), .C2(n_5), .Y(n_372) );
AOI22xp5_ASAP7_75t_L g373 ( .A1(n_316), .A2(n_201), .B1(n_191), .B2(n_118), .Y(n_373) );
INVxp67_ASAP7_75t_L g374 ( .A(n_339), .Y(n_374) );
NOR2x1p5_ASAP7_75t_SL g375 ( .A(n_328), .B(n_119), .Y(n_375) );
INVxp67_ASAP7_75t_L g376 ( .A(n_328), .Y(n_376) );
NAND2xp5_ASAP7_75t_L g377 ( .A(n_341), .B(n_1), .Y(n_377) );
NAND2x1p5_ASAP7_75t_L g378 ( .A(n_342), .B(n_206), .Y(n_378) );
NAND2xp5_ASAP7_75t_L g379 ( .A(n_341), .B(n_2), .Y(n_379) );
AND2x2_ASAP7_75t_L g380 ( .A(n_314), .B(n_3), .Y(n_380) );
INVx1_ASAP7_75t_L g381 ( .A(n_313), .Y(n_381) );
INVx1_ASAP7_75t_L g382 ( .A(n_313), .Y(n_382) );
NOR3xp33_ASAP7_75t_L g383 ( .A(n_321), .B(n_119), .C(n_166), .Y(n_383) );
AOI22xp5_ASAP7_75t_L g384 ( .A1(n_338), .A2(n_191), .B1(n_206), .B2(n_210), .Y(n_384) );
AOI32xp33_ASAP7_75t_L g385 ( .A1(n_344), .A2(n_6), .A3(n_7), .B1(n_8), .B2(n_9), .Y(n_385) );
INVxp67_ASAP7_75t_L g386 ( .A(n_347), .Y(n_386) );
NAND2xp5_ASAP7_75t_L g387 ( .A(n_319), .B(n_7), .Y(n_387) );
NOR2x1_ASAP7_75t_L g388 ( .A(n_340), .B(n_206), .Y(n_388) );
OAI22xp5_ASAP7_75t_L g389 ( .A1(n_340), .A2(n_346), .B1(n_335), .B2(n_327), .Y(n_389) );
OR2x2_ASAP7_75t_L g390 ( .A(n_336), .B(n_8), .Y(n_390) );
AOI22xp5_ASAP7_75t_L g391 ( .A1(n_338), .A2(n_210), .B1(n_207), .B2(n_188), .Y(n_391) );
AOI22xp5_ASAP7_75t_L g392 ( .A1(n_343), .A2(n_210), .B1(n_207), .B2(n_188), .Y(n_392) );
AND2x2_ASAP7_75t_L g393 ( .A(n_317), .B(n_10), .Y(n_393) );
INVx1_ASAP7_75t_SL g394 ( .A(n_351), .Y(n_394) );
INVx1_ASAP7_75t_L g395 ( .A(n_319), .Y(n_395) );
INVx1_ASAP7_75t_L g396 ( .A(n_323), .Y(n_396) );
AND2x2_ASAP7_75t_L g397 ( .A(n_317), .B(n_10), .Y(n_397) );
INVx1_ASAP7_75t_L g398 ( .A(n_323), .Y(n_398) );
A2O1A1Ixp33_ASAP7_75t_L g399 ( .A1(n_342), .A2(n_11), .B(n_12), .C(n_13), .Y(n_399) );
OAI21xp33_ASAP7_75t_L g400 ( .A1(n_322), .A2(n_151), .B(n_140), .Y(n_400) );
AOI33xp33_ASAP7_75t_L g401 ( .A1(n_322), .A2(n_13), .A3(n_151), .B1(n_140), .B2(n_134), .B3(n_26), .Y(n_401) );
AND2x2_ASAP7_75t_L g402 ( .A(n_357), .B(n_326), .Y(n_402) );
INVx1_ASAP7_75t_L g403 ( .A(n_364), .Y(n_403) );
NOR3xp33_ASAP7_75t_SL g404 ( .A(n_399), .B(n_329), .C(n_327), .Y(n_404) );
AO21x1_ASAP7_75t_L g405 ( .A1(n_356), .A2(n_324), .B(n_325), .Y(n_405) );
NAND2xp5_ASAP7_75t_L g406 ( .A(n_380), .B(n_324), .Y(n_406) );
XNOR2x2_ASAP7_75t_L g407 ( .A(n_362), .B(n_347), .Y(n_407) );
INVx2_ASAP7_75t_L g408 ( .A(n_371), .Y(n_408) );
NAND2xp5_ASAP7_75t_L g409 ( .A(n_393), .B(n_325), .Y(n_409) );
NAND2xp5_ASAP7_75t_L g410 ( .A(n_397), .B(n_329), .Y(n_410) );
INVx1_ASAP7_75t_L g411 ( .A(n_381), .Y(n_411) );
INVx2_ASAP7_75t_SL g412 ( .A(n_354), .Y(n_412) );
INVx1_ASAP7_75t_L g413 ( .A(n_382), .Y(n_413) );
INVx1_ASAP7_75t_L g414 ( .A(n_395), .Y(n_414) );
INVx1_ASAP7_75t_L g415 ( .A(n_396), .Y(n_415) );
INVxp67_ASAP7_75t_L g416 ( .A(n_361), .Y(n_416) );
XNOR2xp5_ASAP7_75t_L g417 ( .A(n_367), .B(n_343), .Y(n_417) );
INVx1_ASAP7_75t_L g418 ( .A(n_398), .Y(n_418) );
INVx1_ASAP7_75t_L g419 ( .A(n_374), .Y(n_419) );
INVx1_ASAP7_75t_L g420 ( .A(n_386), .Y(n_420) );
OAI21xp33_ASAP7_75t_L g421 ( .A1(n_355), .A2(n_326), .B(n_350), .Y(n_421) );
INVxp67_ASAP7_75t_SL g422 ( .A(n_370), .Y(n_422) );
OAI21xp5_ASAP7_75t_L g423 ( .A1(n_383), .A2(n_336), .B(n_350), .Y(n_423) );
NOR2xp33_ASAP7_75t_L g424 ( .A(n_352), .B(n_326), .Y(n_424) );
XNOR2x2_ASAP7_75t_L g425 ( .A(n_389), .B(n_351), .Y(n_425) );
INVx2_ASAP7_75t_L g426 ( .A(n_363), .Y(n_426) );
INVx1_ASAP7_75t_L g427 ( .A(n_353), .Y(n_427) );
AND2x2_ASAP7_75t_L g428 ( .A(n_394), .B(n_348), .Y(n_428) );
OR2x2_ASAP7_75t_L g429 ( .A(n_376), .B(n_348), .Y(n_429) );
NOR2xp33_ASAP7_75t_L g430 ( .A(n_377), .B(n_20), .Y(n_430) );
INVx1_ASAP7_75t_L g431 ( .A(n_358), .Y(n_431) );
NOR2x1_ASAP7_75t_L g432 ( .A(n_388), .B(n_164), .Y(n_432) );
INVx1_ASAP7_75t_L g433 ( .A(n_360), .Y(n_433) );
INVx2_ASAP7_75t_L g434 ( .A(n_365), .Y(n_434) );
AO22x1_ASAP7_75t_L g435 ( .A1(n_366), .A2(n_359), .B1(n_379), .B2(n_387), .Y(n_435) );
NAND2xp5_ASAP7_75t_L g436 ( .A(n_368), .B(n_22), .Y(n_436) );
INVx1_ASAP7_75t_L g437 ( .A(n_390), .Y(n_437) );
INVx1_ASAP7_75t_L g438 ( .A(n_375), .Y(n_438) );
NAND2xp5_ASAP7_75t_SL g439 ( .A(n_400), .B(n_207), .Y(n_439) );
INVx2_ASAP7_75t_L g440 ( .A(n_366), .Y(n_440) );
INVx1_ASAP7_75t_SL g441 ( .A(n_378), .Y(n_441) );
INVx1_ASAP7_75t_L g442 ( .A(n_384), .Y(n_442) );
INVx1_ASAP7_75t_L g443 ( .A(n_384), .Y(n_443) );
INVx1_ASAP7_75t_L g444 ( .A(n_392), .Y(n_444) );
AOI22xp5_ASAP7_75t_L g445 ( .A1(n_405), .A2(n_372), .B1(n_373), .B2(n_368), .Y(n_445) );
INVx1_ASAP7_75t_L g446 ( .A(n_420), .Y(n_446) );
NOR3xp33_ASAP7_75t_L g447 ( .A(n_435), .B(n_385), .C(n_401), .Y(n_447) );
OAI21xp33_ASAP7_75t_L g448 ( .A1(n_421), .A2(n_373), .B(n_392), .Y(n_448) );
NOR2x1_ASAP7_75t_L g449 ( .A(n_441), .B(n_369), .Y(n_449) );
AO22x2_ASAP7_75t_L g450 ( .A1(n_419), .A2(n_391), .B1(n_151), .B2(n_140), .Y(n_450) );
INVx1_ASAP7_75t_L g451 ( .A(n_408), .Y(n_451) );
INVx1_ASAP7_75t_L g452 ( .A(n_408), .Y(n_452) );
OAI21xp5_ASAP7_75t_SL g453 ( .A1(n_412), .A2(n_207), .B(n_188), .Y(n_453) );
NAND2xp5_ASAP7_75t_L g454 ( .A(n_433), .B(n_25), .Y(n_454) );
INVx1_ASAP7_75t_L g455 ( .A(n_403), .Y(n_455) );
AOI22xp33_ASAP7_75t_L g456 ( .A1(n_442), .A2(n_135), .B1(n_188), .B2(n_207), .Y(n_456) );
INVx1_ASAP7_75t_L g457 ( .A(n_411), .Y(n_457) );
INVx1_ASAP7_75t_L g458 ( .A(n_413), .Y(n_458) );
AOI21x1_ASAP7_75t_L g459 ( .A1(n_439), .A2(n_134), .B(n_33), .Y(n_459) );
NOR3x1_ASAP7_75t_L g460 ( .A(n_425), .B(n_427), .C(n_407), .Y(n_460) );
NAND2xp5_ASAP7_75t_L g461 ( .A(n_444), .B(n_28), .Y(n_461) );
AOI22xp5_ASAP7_75t_L g462 ( .A1(n_424), .A2(n_134), .B1(n_135), .B2(n_188), .Y(n_462) );
INVx1_ASAP7_75t_L g463 ( .A(n_414), .Y(n_463) );
NOR2xp33_ASAP7_75t_L g464 ( .A(n_424), .B(n_34), .Y(n_464) );
OAI22xp5_ASAP7_75t_SL g465 ( .A1(n_417), .A2(n_35), .B1(n_36), .B2(n_37), .Y(n_465) );
NOR2x1_ASAP7_75t_L g466 ( .A(n_438), .B(n_207), .Y(n_466) );
NAND2xp5_ASAP7_75t_L g467 ( .A(n_437), .B(n_38), .Y(n_467) );
AOI21xp5_ASAP7_75t_L g468 ( .A1(n_439), .A2(n_207), .B(n_188), .Y(n_468) );
XOR2xp5_ASAP7_75t_L g469 ( .A(n_406), .B(n_41), .Y(n_469) );
INVx1_ASAP7_75t_L g470 ( .A(n_415), .Y(n_470) );
INVx1_ASAP7_75t_L g471 ( .A(n_418), .Y(n_471) );
INVx1_ASAP7_75t_L g472 ( .A(n_431), .Y(n_472) );
INVx1_ASAP7_75t_L g473 ( .A(n_429), .Y(n_473) );
NAND2xp5_ASAP7_75t_L g474 ( .A(n_446), .B(n_443), .Y(n_474) );
INVx1_ASAP7_75t_L g475 ( .A(n_455), .Y(n_475) );
NAND2xp33_ASAP7_75t_SL g476 ( .A(n_460), .B(n_404), .Y(n_476) );
INVx1_ASAP7_75t_L g477 ( .A(n_457), .Y(n_477) );
INVx2_ASAP7_75t_SL g478 ( .A(n_473), .Y(n_478) );
AOI222xp33_ASAP7_75t_L g479 ( .A1(n_448), .A2(n_472), .B1(n_409), .B2(n_410), .C1(n_471), .C2(n_463), .Y(n_479) );
AOI322xp5_ASAP7_75t_L g480 ( .A1(n_447), .A2(n_404), .A3(n_426), .B1(n_402), .B2(n_422), .C1(n_434), .C2(n_416), .Y(n_480) );
OAI21xp5_ASAP7_75t_L g481 ( .A1(n_445), .A2(n_423), .B(n_416), .Y(n_481) );
AOI22xp5_ASAP7_75t_L g482 ( .A1(n_445), .A2(n_440), .B1(n_434), .B2(n_422), .Y(n_482) );
OAI21xp5_ASAP7_75t_L g483 ( .A1(n_453), .A2(n_432), .B(n_430), .Y(n_483) );
INVx1_ASAP7_75t_L g484 ( .A(n_458), .Y(n_484) );
NOR2xp33_ASAP7_75t_L g485 ( .A(n_470), .B(n_426), .Y(n_485) );
INVx1_ASAP7_75t_SL g486 ( .A(n_469), .Y(n_486) );
NAND2xp5_ASAP7_75t_L g487 ( .A(n_451), .B(n_428), .Y(n_487) );
NOR2xp33_ASAP7_75t_R g488 ( .A(n_459), .B(n_430), .Y(n_488) );
AOI31xp33_ASAP7_75t_L g489 ( .A1(n_449), .A2(n_436), .A3(n_440), .B(n_47), .Y(n_489) );
NOR2x1_ASAP7_75t_SL g490 ( .A(n_452), .B(n_188), .Y(n_490) );
AOI22xp5_ASAP7_75t_L g491 ( .A1(n_465), .A2(n_135), .B1(n_143), .B2(n_48), .Y(n_491) );
OAI21xp5_ASAP7_75t_L g492 ( .A1(n_466), .A2(n_44), .B(n_46), .Y(n_492) );
OAI211xp5_ASAP7_75t_SL g493 ( .A1(n_467), .A2(n_49), .B(n_50), .C(n_51), .Y(n_493) );
OAI221xp5_ASAP7_75t_L g494 ( .A1(n_464), .A2(n_135), .B1(n_55), .B2(n_58), .C(n_59), .Y(n_494) );
NOR3xp33_ASAP7_75t_L g495 ( .A(n_461), .B(n_52), .C(n_60), .Y(n_495) );
AOI22xp5_ASAP7_75t_L g496 ( .A1(n_450), .A2(n_454), .B1(n_462), .B2(n_456), .Y(n_496) );
OAI211xp5_ASAP7_75t_SL g497 ( .A1(n_468), .A2(n_61), .B(n_62), .C(n_64), .Y(n_497) );
NAND4xp75_ASAP7_75t_L g498 ( .A(n_450), .B(n_65), .C(n_67), .D(n_68), .Y(n_498) );
OAI22xp5_ASAP7_75t_L g499 ( .A1(n_445), .A2(n_135), .B1(n_73), .B2(n_74), .Y(n_499) );
AOI22xp33_ASAP7_75t_R g500 ( .A1(n_488), .A2(n_486), .B1(n_476), .B2(n_480), .Y(n_500) );
BUFx2_ASAP7_75t_L g501 ( .A(n_481), .Y(n_501) );
OAI322xp33_ASAP7_75t_L g502 ( .A1(n_482), .A2(n_474), .A3(n_478), .B1(n_484), .B2(n_475), .C1(n_477), .C2(n_485), .Y(n_502) );
NAND3x1_ASAP7_75t_L g503 ( .A(n_483), .B(n_491), .C(n_496), .Y(n_503) );
INVxp67_ASAP7_75t_SL g504 ( .A(n_499), .Y(n_504) );
NOR3xp33_ASAP7_75t_L g505 ( .A(n_501), .B(n_489), .C(n_494), .Y(n_505) );
NAND3xp33_ASAP7_75t_L g506 ( .A(n_500), .B(n_479), .C(n_495), .Y(n_506) );
NAND5xp2_ASAP7_75t_L g507 ( .A(n_504), .B(n_492), .C(n_488), .D(n_485), .E(n_498), .Y(n_507) );
INVx1_ASAP7_75t_SL g508 ( .A(n_506), .Y(n_508) );
OAI322xp33_ASAP7_75t_L g509 ( .A1(n_505), .A2(n_504), .A3(n_503), .B1(n_502), .B2(n_487), .C1(n_490), .C2(n_493), .Y(n_509) );
AND3x4_ASAP7_75t_L g510 ( .A(n_509), .B(n_507), .C(n_497), .Y(n_510) );
AOI322xp5_ASAP7_75t_L g511 ( .A1(n_510), .A2(n_72), .A3(n_135), .B1(n_143), .B2(n_153), .C1(n_508), .C2(n_501), .Y(n_511) );
AOI21xp5_ASAP7_75t_L g512 ( .A1(n_511), .A2(n_153), .B(n_143), .Y(n_512) );
endmodule