module fake_jpeg_7760_n_231 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_231);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_231;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_96;

BUFx12f_ASAP7_75t_L g15 ( 
.A(n_13),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

BUFx5_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_10),
.B(n_0),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_11),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_9),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_10),
.Y(n_27)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_7),
.B(n_11),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_17),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_31),
.B(n_32),
.Y(n_47)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_17),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_33),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_15),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_34),
.B(n_35),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_15),
.Y(n_35)
);

AOI22xp5_ASAP7_75t_L g36 ( 
.A1(n_28),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_SL g42 ( 
.A1(n_36),
.A2(n_20),
.B1(n_18),
.B2(n_16),
.Y(n_42)
);

INVx11_ASAP7_75t_L g37 ( 
.A(n_22),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_37),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_15),
.Y(n_38)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_38),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_15),
.Y(n_39)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_39),
.Y(n_57)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_17),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_40),
.B(n_41),
.Y(n_51)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_19),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_42),
.A2(n_46),
.B1(n_52),
.B2(n_61),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_L g46 ( 
.A1(n_37),
.A2(n_28),
.B1(n_20),
.B2(n_18),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_33),
.Y(n_49)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_49),
.Y(n_63)
);

AOI21xp33_ASAP7_75t_L g50 ( 
.A1(n_36),
.A2(n_23),
.B(n_30),
.Y(n_50)
);

A2O1A1Ixp33_ASAP7_75t_L g81 ( 
.A1(n_50),
.A2(n_25),
.B(n_19),
.C(n_21),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_L g52 ( 
.A1(n_37),
.A2(n_28),
.B1(n_41),
.B2(n_32),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_37),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_53),
.B(n_56),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_36),
.B(n_30),
.Y(n_54)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_54),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_34),
.B(n_23),
.Y(n_55)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_55),
.Y(n_68)
);

CKINVDCx16_ASAP7_75t_R g56 ( 
.A(n_32),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_34),
.B(n_24),
.Y(n_58)
);

XNOR2xp5_ASAP7_75t_L g66 ( 
.A(n_58),
.B(n_41),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_35),
.B(n_20),
.Y(n_59)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_59),
.Y(n_70)
);

BUFx4f_ASAP7_75t_SL g60 ( 
.A(n_33),
.Y(n_60)
);

CKINVDCx16_ASAP7_75t_R g79 ( 
.A(n_60),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_41),
.A2(n_27),
.B1(n_26),
.B2(n_25),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_35),
.B(n_29),
.Y(n_62)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_62),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_61),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_65),
.B(n_76),
.Y(n_86)
);

AND2x2_ASAP7_75t_L g85 ( 
.A(n_66),
.B(n_58),
.Y(n_85)
);

OAI21xp5_ASAP7_75t_L g67 ( 
.A1(n_54),
.A2(n_16),
.B(n_40),
.Y(n_67)
);

AOI21xp5_ASAP7_75t_SL g103 ( 
.A1(n_67),
.A2(n_55),
.B(n_47),
.Y(n_103)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_45),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_69),
.Y(n_91)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_59),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_73),
.B(n_62),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g74 ( 
.A(n_51),
.Y(n_74)
);

CKINVDCx16_ASAP7_75t_R g89 ( 
.A(n_74),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_58),
.Y(n_76)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_49),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_77),
.B(n_82),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_43),
.A2(n_29),
.B1(n_27),
.B2(n_26),
.Y(n_78)
);

INVxp67_ASAP7_75t_L g99 ( 
.A(n_78),
.Y(n_99)
);

BUFx2_ASAP7_75t_L g80 ( 
.A(n_45),
.Y(n_80)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_80),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_SL g100 ( 
.A(n_81),
.B(n_42),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_L g82 ( 
.A1(n_50),
.A2(n_40),
.B1(n_31),
.B2(n_19),
.Y(n_82)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_80),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_85),
.B(n_93),
.Y(n_105)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_87),
.Y(n_108)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_72),
.Y(n_88)
);

XNOR2xp5_ASAP7_75t_L g90 ( 
.A(n_66),
.B(n_48),
.Y(n_90)
);

XNOR2xp5_ASAP7_75t_L g122 ( 
.A(n_90),
.B(n_98),
.Y(n_122)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_80),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_92),
.B(n_94),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_64),
.B(n_67),
.Y(n_93)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_72),
.Y(n_94)
);

AND2x2_ASAP7_75t_SL g95 ( 
.A(n_64),
.B(n_57),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_95),
.B(n_97),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_74),
.B(n_42),
.Y(n_97)
);

XNOR2xp5_ASAP7_75t_L g98 ( 
.A(n_81),
.B(n_48),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_100),
.A2(n_65),
.B1(n_68),
.B2(n_76),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_71),
.B(n_51),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_101),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_71),
.B(n_47),
.Y(n_102)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_102),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_103),
.A2(n_68),
.B1(n_73),
.B2(n_70),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_L g135 ( 
.A1(n_104),
.A2(n_113),
.B(n_83),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_106),
.B(n_98),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_97),
.A2(n_75),
.B1(n_52),
.B2(n_46),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_107),
.A2(n_117),
.B1(n_63),
.B2(n_45),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_86),
.A2(n_99),
.B1(n_75),
.B2(n_96),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_L g130 ( 
.A1(n_109),
.A2(n_89),
.B1(n_103),
.B2(n_85),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_87),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_110),
.B(n_114),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_100),
.A2(n_70),
.B1(n_56),
.B2(n_43),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_112),
.A2(n_120),
.B1(n_124),
.B2(n_92),
.Y(n_129)
);

AOI21xp5_ASAP7_75t_L g113 ( 
.A1(n_99),
.A2(n_60),
.B(n_79),
.Y(n_113)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_95),
.Y(n_114)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_95),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_115),
.B(n_121),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_93),
.A2(n_53),
.B1(n_43),
.B2(n_44),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_88),
.A2(n_43),
.B1(n_57),
.B2(n_44),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_95),
.Y(n_121)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_84),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_123),
.B(n_49),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_94),
.A2(n_57),
.B1(n_44),
.B2(n_31),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_122),
.B(n_90),
.C(n_85),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_125),
.B(n_122),
.C(n_105),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_126),
.B(n_127),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_104),
.B(n_89),
.Y(n_127)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_123),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_128),
.B(n_133),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_130),
.A2(n_132),
.B1(n_140),
.B2(n_127),
.Y(n_157)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_118),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_131),
.B(n_134),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_SL g132 ( 
.A1(n_114),
.A2(n_69),
.B1(n_63),
.B2(n_77),
.Y(n_132)
);

AOI21xp5_ASAP7_75t_L g133 ( 
.A1(n_115),
.A2(n_79),
.B(n_60),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_120),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_135),
.B(n_139),
.Y(n_160)
);

INVxp67_ASAP7_75t_L g137 ( 
.A(n_113),
.Y(n_137)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_137),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_119),
.B(n_83),
.Y(n_139)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_141),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_L g142 ( 
.A1(n_119),
.A2(n_21),
.B(n_24),
.Y(n_142)
);

XOR2xp5_ASAP7_75t_L g148 ( 
.A(n_142),
.B(n_107),
.Y(n_148)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_124),
.Y(n_143)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_143),
.Y(n_154)
);

HB1xp67_ASAP7_75t_L g144 ( 
.A(n_117),
.Y(n_144)
);

INVx3_ASAP7_75t_L g159 ( 
.A(n_144),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_112),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_145),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_147),
.B(n_148),
.C(n_150),
.Y(n_167)
);

XOR2xp5_ASAP7_75t_L g150 ( 
.A(n_125),
.B(n_105),
.Y(n_150)
);

XOR2xp5_ASAP7_75t_L g153 ( 
.A(n_126),
.B(n_121),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_153),
.B(n_156),
.C(n_164),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_139),
.B(n_108),
.C(n_111),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_157),
.A2(n_161),
.B1(n_162),
.B2(n_131),
.Y(n_177)
);

AOI322xp5_ASAP7_75t_L g158 ( 
.A1(n_135),
.A2(n_108),
.A3(n_116),
.B1(n_111),
.B2(n_60),
.C1(n_39),
.C2(n_33),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_SL g178 ( 
.A(n_158),
.B(n_140),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_145),
.A2(n_116),
.B1(n_91),
.B2(n_60),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_130),
.A2(n_91),
.B1(n_45),
.B2(n_39),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_138),
.B(n_39),
.C(n_33),
.Y(n_164)
);

OAI321xp33_ASAP7_75t_L g165 ( 
.A1(n_144),
.A2(n_24),
.A3(n_22),
.B1(n_39),
.B2(n_38),
.C(n_21),
.Y(n_165)
);

AO21x1_ASAP7_75t_L g183 ( 
.A1(n_165),
.A2(n_21),
.B(n_24),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_138),
.B(n_38),
.C(n_91),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_166),
.B(n_141),
.C(n_133),
.Y(n_176)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_155),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_168),
.B(n_169),
.Y(n_195)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_155),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_163),
.B(n_136),
.Y(n_171)
);

AOI321xp33_ASAP7_75t_L g172 ( 
.A1(n_153),
.A2(n_136),
.A3(n_142),
.B1(n_143),
.B2(n_129),
.C(n_134),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g187 ( 
.A(n_172),
.B(n_178),
.Y(n_187)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_161),
.Y(n_173)
);

AOI21xp5_ASAP7_75t_L g189 ( 
.A1(n_173),
.A2(n_174),
.B(n_179),
.Y(n_189)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_166),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_154),
.B(n_149),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_175),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_176),
.B(n_147),
.C(n_164),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_177),
.A2(n_183),
.B1(n_21),
.B2(n_22),
.Y(n_192)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_152),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_160),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_180),
.A2(n_182),
.B1(n_8),
.B2(n_13),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_160),
.Y(n_181)
);

INVx3_ASAP7_75t_L g197 ( 
.A(n_181),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_SL g182 ( 
.A(n_149),
.B(n_128),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_151),
.B(n_22),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_L g188 ( 
.A(n_184),
.B(n_171),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_168),
.A2(n_157),
.B1(n_159),
.B2(n_162),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_L g208 ( 
.A1(n_185),
.A2(n_186),
.B1(n_194),
.B2(n_178),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_169),
.A2(n_159),
.B1(n_146),
.B2(n_148),
.Y(n_186)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_188),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g190 ( 
.A(n_167),
.B(n_150),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_190),
.B(n_191),
.C(n_193),
.Y(n_199)
);

CKINVDCx16_ASAP7_75t_R g202 ( 
.A(n_192),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g193 ( 
.A(n_167),
.B(n_38),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_173),
.A2(n_7),
.B1(n_13),
.B2(n_12),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_196),
.B(n_183),
.Y(n_200)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_200),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g201 ( 
.A(n_187),
.B(n_170),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_201),
.B(n_204),
.C(n_205),
.Y(n_216)
);

OAI31xp33_ASAP7_75t_L g203 ( 
.A1(n_195),
.A2(n_180),
.A3(n_179),
.B(n_172),
.Y(n_203)
);

OR2x2_ASAP7_75t_L g215 ( 
.A(n_203),
.B(n_6),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_187),
.B(n_186),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_191),
.B(n_170),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_198),
.B(n_176),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g210 ( 
.A(n_206),
.B(n_208),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_202),
.A2(n_185),
.B1(n_197),
.B2(n_189),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_209),
.B(n_213),
.Y(n_221)
);

A2O1A1Ixp33_ASAP7_75t_SL g212 ( 
.A1(n_203),
.A2(n_197),
.B(n_207),
.C(n_204),
.Y(n_212)
);

NAND4xp25_ASAP7_75t_SL g213 ( 
.A(n_199),
.B(n_1),
.C(n_2),
.D(n_3),
.Y(n_213)
);

AOI21xp33_ASAP7_75t_L g214 ( 
.A1(n_199),
.A2(n_6),
.B(n_12),
.Y(n_214)
);

OAI21xp5_ASAP7_75t_SL g218 ( 
.A1(n_214),
.A2(n_215),
.B(n_14),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_SL g217 ( 
.A(n_215),
.B(n_6),
.Y(n_217)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_217),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_218),
.B(n_14),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_SL g219 ( 
.A(n_210),
.B(n_9),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_219),
.B(n_211),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_216),
.B(n_1),
.C(n_3),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_223),
.B(n_224),
.Y(n_227)
);

OAI21xp5_ASAP7_75t_SL g225 ( 
.A1(n_221),
.A2(n_212),
.B(n_216),
.Y(n_225)
);

MAJx2_ASAP7_75t_L g226 ( 
.A(n_222),
.B(n_212),
.C(n_220),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_226),
.B(n_228),
.C(n_3),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_225),
.B(n_212),
.C(n_3),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_229),
.B(n_227),
.C(n_4),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_230),
.B(n_4),
.Y(n_231)
);


endmodule