module fake_jpeg_29027_n_84 (n_13, n_21, n_1, n_10, n_23, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_26, n_9, n_5, n_11, n_17, n_25, n_2, n_12, n_8, n_15, n_7, n_84);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_84;

wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_57;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_44;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_35;
wire n_48;
wire n_46;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;

INVx4_ASAP7_75t_L g27 ( 
.A(n_18),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_5),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_17),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_23),
.Y(n_30)
);

BUFx16f_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_24),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_21),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_16),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_28),
.B(n_0),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_35),
.B(n_37),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_28),
.B(n_0),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_36),
.B(n_2),
.Y(n_51)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_33),
.Y(n_37)
);

AND2x2_ASAP7_75t_L g38 ( 
.A(n_31),
.B(n_1),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_38),
.B(n_40),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g39 ( 
.A1(n_31),
.A2(n_27),
.B1(n_29),
.B2(n_34),
.Y(n_39)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_39),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_31),
.Y(n_40)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_27),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_41),
.B(n_29),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_SL g42 ( 
.A(n_38),
.B(n_30),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_SL g55 ( 
.A(n_42),
.B(n_44),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_SL g44 ( 
.A(n_41),
.B(n_32),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_SL g45 ( 
.A(n_39),
.B(n_33),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_45),
.B(n_50),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_SL g47 ( 
.A(n_36),
.B(n_1),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_SL g56 ( 
.A(n_47),
.B(n_51),
.Y(n_56)
);

AND2x2_ASAP7_75t_L g52 ( 
.A(n_49),
.B(n_34),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_36),
.B(n_2),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_52),
.B(n_60),
.Y(n_68)
);

CKINVDCx16_ASAP7_75t_R g53 ( 
.A(n_48),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_53),
.B(n_54),
.Y(n_63)
);

INVxp67_ASAP7_75t_L g54 ( 
.A(n_46),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g57 ( 
.A1(n_48),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_57),
.A2(n_58),
.B1(n_59),
.B2(n_12),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g58 ( 
.A1(n_47),
.A2(n_4),
.B1(n_6),
.B2(n_7),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_L g59 ( 
.A1(n_43),
.A2(n_6),
.B1(n_8),
.B2(n_9),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_47),
.B(n_10),
.Y(n_60)
);

INVxp67_ASAP7_75t_L g62 ( 
.A(n_52),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_62),
.B(n_65),
.Y(n_72)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_61),
.Y(n_64)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_64),
.Y(n_75)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_59),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_55),
.B(n_11),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_66),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_56),
.B(n_26),
.Y(n_67)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_67),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g76 ( 
.A1(n_69),
.A2(n_14),
.B1(n_15),
.B2(n_19),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_SL g70 ( 
.A(n_56),
.B(n_25),
.Y(n_70)
);

NOR2xp67_ASAP7_75t_SL g74 ( 
.A(n_70),
.B(n_13),
.Y(n_74)
);

XNOR2xp5_ASAP7_75t_L g78 ( 
.A(n_74),
.B(n_76),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_75),
.B(n_68),
.C(n_63),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_77),
.A2(n_71),
.B1(n_62),
.B2(n_73),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_79),
.B(n_78),
.C(n_72),
.Y(n_80)
);

INVxp67_ASAP7_75t_L g81 ( 
.A(n_80),
.Y(n_81)
);

INVxp67_ASAP7_75t_L g82 ( 
.A(n_81),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_82),
.B(n_20),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_83),
.B(n_22),
.Y(n_84)
);


endmodule