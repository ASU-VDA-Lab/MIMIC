module real_aes_5063_n_77 (n_17, n_28, n_76, n_56, n_34, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_43, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_44, n_7, n_4, n_6, n_12, n_68, n_69, n_46, n_59, n_25, n_73, n_48, n_37, n_70, n_50, n_26, n_13, n_24, n_2, n_55, n_62, n_67, n_33, n_14, n_11, n_16, n_39, n_5, n_45, n_60, n_38, n_0, n_63, n_1, n_53, n_36, n_77);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_43;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_44;
input n_7;
input n_4;
input n_6;
input n_12;
input n_68;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_48;
input n_37;
input n_70;
input n_50;
input n_26;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_67;
input n_33;
input n_14;
input n_11;
input n_16;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_0;
input n_63;
input n_1;
input n_53;
input n_36;
output n_77;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_90;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_518;
wire n_254;
wire n_207;
wire n_580;
wire n_577;
wire n_469;
wire n_83;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_322;
wire n_328;
wire n_318;
wire n_355;
wire n_239;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_319;
wire n_421;
wire n_364;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_376;
wire n_549;
wire n_571;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_560;
wire n_260;
wire n_594;
wire n_97;
wire n_186;
wire n_138;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_235;
wire n_399;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_92;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_94;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_98;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_82;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_517;
wire n_174;
wire n_570;
wire n_530;
wire n_104;
wire n_535;
wire n_211;
wire n_281;
wire n_496;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_178;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_504;
wire n_455;
wire n_164;
wire n_231;
wire n_102;
wire n_547;
wire n_634;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_80;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_367;
wire n_267;
wire n_218;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_339;
wire n_398;
wire n_89;
wire n_277;
wire n_609;
wire n_425;
wire n_331;
wire n_93;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_323;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_654;
wire n_527;
wire n_434;
wire n_502;
wire n_505;
wire n_600;
wire n_250;
wire n_85;
wire n_605;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_87;
wire n_171;
wire n_78;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_96;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_95;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_533;
wire n_366;
wire n_346;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_622;
wire n_470;
wire n_81;
wire n_133;
wire n_494;
wire n_377;
wire n_273;
wire n_114;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_643;
wire n_486;
wire n_411;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_88;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_633;
wire n_520;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_249;
wire n_623;
wire n_446;
wire n_221;
wire n_156;
wire n_359;
wire n_456;
wire n_312;
wire n_266;
wire n_183;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_371;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_99;
wire n_440;
wire n_525;
wire n_644;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_79;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_566;
wire n_474;
wire n_170;
wire n_86;
wire n_375;
wire n_597;
wire n_640;
wire n_340;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_646;
wire n_650;
wire n_105;
wire n_84;
wire n_393;
wire n_294;
wire n_258;
wire n_652;
wire n_206;
wire n_307;
wire n_500;
wire n_601;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_91;
INVx1_ASAP7_75t_L g342 ( .A(n_0), .Y(n_342) );
AOI22xp5_ASAP7_75t_L g241 ( .A1(n_1), .A2(n_16), .B1(n_227), .B2(n_242), .Y(n_241) );
AOI22xp5_ASAP7_75t_L g84 ( .A1(n_2), .A2(n_10), .B1(n_85), .B2(n_109), .Y(n_84) );
INVx2_ASAP7_75t_L g302 ( .A(n_3), .Y(n_302) );
INVx1_ASAP7_75t_SL g367 ( .A(n_4), .Y(n_367) );
AOI22xp33_ASAP7_75t_L g140 ( .A1(n_5), .A2(n_67), .B1(n_141), .B2(n_143), .Y(n_140) );
AOI22xp33_ASAP7_75t_L g129 ( .A1(n_6), .A2(n_43), .B1(n_130), .B2(n_134), .Y(n_129) );
HB1xp67_ASAP7_75t_L g190 ( .A(n_7), .Y(n_190) );
NAND2xp5_ASAP7_75t_L g332 ( .A(n_8), .B(n_333), .Y(n_332) );
NAND2xp5_ASAP7_75t_L g352 ( .A(n_9), .B(n_353), .Y(n_352) );
INVx1_ASAP7_75t_L g106 ( .A(n_11), .Y(n_106) );
NOR2xp33_ASAP7_75t_L g115 ( .A(n_11), .B(n_56), .Y(n_115) );
INVxp67_ASAP7_75t_L g150 ( .A(n_11), .Y(n_150) );
INVx1_ASAP7_75t_L g196 ( .A(n_12), .Y(n_196) );
AOI22xp33_ASAP7_75t_L g347 ( .A1(n_12), .A2(n_42), .B1(n_348), .B2(n_349), .Y(n_347) );
NAND2xp5_ASAP7_75t_L g123 ( .A(n_13), .B(n_124), .Y(n_123) );
OA21x2_ASAP7_75t_L g253 ( .A1(n_14), .A2(n_54), .B(n_254), .Y(n_253) );
OA21x2_ASAP7_75t_L g257 ( .A1(n_14), .A2(n_54), .B(n_254), .Y(n_257) );
NAND2xp5_ASAP7_75t_SL g102 ( .A(n_15), .B(n_91), .Y(n_102) );
NOR2xp33_ASAP7_75t_L g313 ( .A(n_17), .B(n_243), .Y(n_313) );
AOI22xp33_ASAP7_75t_L g162 ( .A1(n_18), .A2(n_64), .B1(n_163), .B2(n_169), .Y(n_162) );
INVx2_ASAP7_75t_L g284 ( .A(n_19), .Y(n_284) );
AOI22xp5_ASAP7_75t_L g292 ( .A1(n_20), .A2(n_61), .B1(n_293), .B2(n_295), .Y(n_292) );
AOI22xp5_ASAP7_75t_L g244 ( .A1(n_21), .A2(n_25), .B1(n_245), .B2(n_247), .Y(n_244) );
BUFx3_ASAP7_75t_L g204 ( .A(n_22), .Y(n_204) );
O2A1O1Ixp5_ASAP7_75t_L g276 ( .A1(n_23), .A2(n_223), .B(n_277), .C(n_281), .Y(n_276) );
AOI22xp33_ASAP7_75t_L g297 ( .A1(n_24), .A2(n_48), .B1(n_278), .B2(n_298), .Y(n_297) );
CKINVDCx5p33_ASAP7_75t_R g389 ( .A(n_26), .Y(n_389) );
BUFx6f_ASAP7_75t_L g91 ( .A(n_27), .Y(n_91) );
AOI22xp33_ASAP7_75t_L g171 ( .A1(n_28), .A2(n_53), .B1(n_172), .B2(n_175), .Y(n_171) );
AOI22xp5_ASAP7_75t_L g355 ( .A1(n_29), .A2(n_62), .B1(n_356), .B2(n_359), .Y(n_355) );
INVx1_ASAP7_75t_L g270 ( .A(n_30), .Y(n_270) );
AOI22xp5_ASAP7_75t_L g152 ( .A1(n_31), .A2(n_47), .B1(n_153), .B2(n_158), .Y(n_152) );
INVx1_ASAP7_75t_L g92 ( .A(n_32), .Y(n_92) );
NAND2xp5_ASAP7_75t_L g147 ( .A(n_32), .B(n_55), .Y(n_147) );
NAND2xp5_ASAP7_75t_L g337 ( .A(n_33), .B(n_266), .Y(n_337) );
CKINVDCx5p33_ASAP7_75t_R g185 ( .A(n_34), .Y(n_185) );
INVx2_ASAP7_75t_L g282 ( .A(n_35), .Y(n_282) );
CKINVDCx5p33_ASAP7_75t_R g390 ( .A(n_36), .Y(n_390) );
INVx2_ASAP7_75t_L g312 ( .A(n_37), .Y(n_312) );
NAND2xp5_ASAP7_75t_L g334 ( .A(n_38), .B(n_335), .Y(n_334) );
INVx1_ASAP7_75t_SL g370 ( .A(n_39), .Y(n_370) );
INVx1_ASAP7_75t_L g385 ( .A(n_40), .Y(n_385) );
INVx1_ASAP7_75t_L g254 ( .A(n_41), .Y(n_254) );
HB1xp67_ASAP7_75t_L g215 ( .A(n_44), .Y(n_215) );
AND2x4_ASAP7_75t_L g219 ( .A(n_44), .B(n_213), .Y(n_219) );
AND2x4_ASAP7_75t_L g274 ( .A(n_44), .B(n_213), .Y(n_274) );
INVx1_ASAP7_75t_L g374 ( .A(n_45), .Y(n_374) );
BUFx6f_ASAP7_75t_L g224 ( .A(n_46), .Y(n_224) );
NOR2xp33_ASAP7_75t_L g317 ( .A(n_49), .B(n_318), .Y(n_317) );
OA22x2_ASAP7_75t_L g96 ( .A1(n_50), .A2(n_56), .B1(n_91), .B2(n_95), .Y(n_96) );
INVx1_ASAP7_75t_L g122 ( .A(n_50), .Y(n_122) );
OAI22xp5_ASAP7_75t_L g645 ( .A1(n_51), .A2(n_80), .B1(n_81), .B2(n_646), .Y(n_645) );
CKINVDCx5p33_ASAP7_75t_R g646 ( .A(n_51), .Y(n_646) );
CKINVDCx5p33_ASAP7_75t_R g192 ( .A(n_52), .Y(n_192) );
INVx1_ASAP7_75t_L g108 ( .A(n_55), .Y(n_108) );
NAND2xp5_ASAP7_75t_L g118 ( .A(n_55), .B(n_119), .Y(n_118) );
HB1xp67_ASAP7_75t_L g207 ( .A(n_55), .Y(n_207) );
OAI21xp33_ASAP7_75t_L g138 ( .A1(n_56), .A2(n_60), .B(n_139), .Y(n_138) );
CKINVDCx5p33_ASAP7_75t_R g380 ( .A(n_57), .Y(n_380) );
CKINVDCx5p33_ASAP7_75t_R g268 ( .A(n_58), .Y(n_268) );
NOR2xp33_ASAP7_75t_L g372 ( .A(n_59), .B(n_248), .Y(n_372) );
INVx1_ASAP7_75t_L g94 ( .A(n_60), .Y(n_94) );
NOR2xp33_ASAP7_75t_L g116 ( .A(n_60), .B(n_74), .Y(n_116) );
BUFx6f_ASAP7_75t_L g228 ( .A(n_63), .Y(n_228) );
BUFx5_ASAP7_75t_L g246 ( .A(n_63), .Y(n_246) );
INVx1_ASAP7_75t_L g280 ( .A(n_63), .Y(n_280) );
NOR2xp33_ASAP7_75t_L g368 ( .A(n_65), .B(n_318), .Y(n_368) );
HB1xp67_ASAP7_75t_L g640 ( .A(n_65), .Y(n_640) );
INVx2_ASAP7_75t_L g315 ( .A(n_66), .Y(n_315) );
INVx1_ASAP7_75t_L g322 ( .A(n_68), .Y(n_322) );
INVx2_ASAP7_75t_L g392 ( .A(n_69), .Y(n_392) );
INVx2_ASAP7_75t_SL g213 ( .A(n_70), .Y(n_213) );
AOI22xp5_ASAP7_75t_L g177 ( .A1(n_71), .A2(n_75), .B1(n_178), .B2(n_181), .Y(n_177) );
NAND2xp5_ASAP7_75t_SL g328 ( .A(n_72), .B(n_329), .Y(n_328) );
HB1xp67_ASAP7_75t_L g195 ( .A(n_73), .Y(n_195) );
NAND2xp5_ASAP7_75t_L g100 ( .A(n_74), .B(n_101), .Y(n_100) );
AO32x2_ASAP7_75t_L g239 ( .A1(n_76), .A2(n_218), .A3(n_240), .B1(n_251), .B2(n_255), .Y(n_239) );
AO22x2_ASAP7_75t_L g397 ( .A1(n_76), .A2(n_240), .B1(n_398), .B2(n_400), .Y(n_397) );
AOI221xp5_ASAP7_75t_L g77 ( .A1(n_78), .A2(n_199), .B1(n_216), .B2(n_229), .C(n_638), .Y(n_77) );
XNOR2xp5_ASAP7_75t_L g78 ( .A(n_79), .B(n_186), .Y(n_78) );
OAI22xp5_ASAP7_75t_L g79 ( .A1(n_80), .A2(n_81), .B1(n_183), .B2(n_184), .Y(n_79) );
OAI22xp5_ASAP7_75t_L g639 ( .A1(n_80), .A2(n_81), .B1(n_640), .B2(n_641), .Y(n_639) );
INVx1_ASAP7_75t_L g80 ( .A(n_81), .Y(n_80) );
HB1xp67_ASAP7_75t_L g81 ( .A(n_82), .Y(n_81) );
NOR2x1_ASAP7_75t_L g82 ( .A(n_83), .B(n_151), .Y(n_82) );
NAND4xp25_ASAP7_75t_L g83 ( .A(n_84), .B(n_123), .C(n_129), .D(n_140), .Y(n_83) );
INVx2_ASAP7_75t_L g85 ( .A(n_86), .Y(n_85) );
INVx3_ASAP7_75t_L g86 ( .A(n_87), .Y(n_86) );
AND2x2_ASAP7_75t_L g87 ( .A(n_88), .B(n_97), .Y(n_87) );
AND2x2_ASAP7_75t_L g142 ( .A(n_88), .B(n_133), .Y(n_142) );
AND2x4_ASAP7_75t_L g154 ( .A(n_88), .B(n_155), .Y(n_154) );
AND2x2_ASAP7_75t_L g182 ( .A(n_88), .B(n_167), .Y(n_182) );
AND2x2_ASAP7_75t_L g88 ( .A(n_89), .B(n_96), .Y(n_88) );
INVx1_ASAP7_75t_L g128 ( .A(n_89), .Y(n_128) );
NAND2xp5_ASAP7_75t_L g89 ( .A(n_90), .B(n_93), .Y(n_89) );
NAND2xp33_ASAP7_75t_L g90 ( .A(n_91), .B(n_92), .Y(n_90) );
INVx2_ASAP7_75t_L g95 ( .A(n_91), .Y(n_95) );
INVx3_ASAP7_75t_L g101 ( .A(n_91), .Y(n_101) );
NAND2xp33_ASAP7_75t_L g107 ( .A(n_91), .B(n_108), .Y(n_107) );
HB1xp67_ASAP7_75t_L g113 ( .A(n_91), .Y(n_113) );
INVx1_ASAP7_75t_L g139 ( .A(n_91), .Y(n_139) );
NAND2xp5_ASAP7_75t_L g121 ( .A(n_92), .B(n_122), .Y(n_121) );
INVxp67_ASAP7_75t_L g208 ( .A(n_92), .Y(n_208) );
NAND2xp5_ASAP7_75t_L g93 ( .A(n_94), .B(n_95), .Y(n_93) );
OAI21xp5_ASAP7_75t_L g149 ( .A1(n_94), .A2(n_139), .B(n_150), .Y(n_149) );
AND2x2_ASAP7_75t_L g127 ( .A(n_96), .B(n_128), .Y(n_127) );
AND2x2_ASAP7_75t_L g148 ( .A(n_96), .B(n_149), .Y(n_148) );
INVx1_ASAP7_75t_L g166 ( .A(n_96), .Y(n_166) );
AND2x4_ASAP7_75t_L g126 ( .A(n_97), .B(n_127), .Y(n_126) );
AND2x4_ASAP7_75t_L g136 ( .A(n_97), .B(n_137), .Y(n_136) );
AND2x2_ASAP7_75t_L g176 ( .A(n_97), .B(n_165), .Y(n_176) );
AND2x4_ASAP7_75t_L g97 ( .A(n_98), .B(n_103), .Y(n_97) );
INVx2_ASAP7_75t_L g98 ( .A(n_99), .Y(n_98) );
AND2x4_ASAP7_75t_L g133 ( .A(n_99), .B(n_103), .Y(n_133) );
AND2x2_ASAP7_75t_L g145 ( .A(n_99), .B(n_146), .Y(n_145) );
OR2x2_ASAP7_75t_L g156 ( .A(n_99), .B(n_157), .Y(n_156) );
AND2x4_ASAP7_75t_L g167 ( .A(n_99), .B(n_168), .Y(n_167) );
AND2x4_ASAP7_75t_L g99 ( .A(n_100), .B(n_102), .Y(n_99) );
NAND2xp5_ASAP7_75t_L g105 ( .A(n_101), .B(n_106), .Y(n_105) );
INVxp67_ASAP7_75t_L g119 ( .A(n_101), .Y(n_119) );
NAND3xp33_ASAP7_75t_L g117 ( .A(n_102), .B(n_118), .C(n_120), .Y(n_117) );
INVx1_ASAP7_75t_L g103 ( .A(n_104), .Y(n_103) );
INVx1_ASAP7_75t_L g157 ( .A(n_104), .Y(n_157) );
AND2x2_ASAP7_75t_L g104 ( .A(n_105), .B(n_107), .Y(n_104) );
INVx1_ASAP7_75t_L g109 ( .A(n_110), .Y(n_109) );
BUFx6f_ASAP7_75t_L g110 ( .A(n_111), .Y(n_110) );
AO21x2_ASAP7_75t_L g111 ( .A1(n_112), .A2(n_114), .B(n_117), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_113), .Y(n_112) );
NAND2xp5_ASAP7_75t_L g146 ( .A(n_113), .B(n_147), .Y(n_146) );
NAND2xp5_ASAP7_75t_L g114 ( .A(n_115), .B(n_116), .Y(n_114) );
NAND2xp5_ASAP7_75t_L g120 ( .A(n_119), .B(n_121), .Y(n_120) );
AND2x2_ASAP7_75t_L g137 ( .A(n_120), .B(n_138), .Y(n_137) );
HB1xp67_ASAP7_75t_L g209 ( .A(n_122), .Y(n_209) );
INVx3_ASAP7_75t_L g124 ( .A(n_125), .Y(n_124) );
INVx2_ASAP7_75t_L g125 ( .A(n_126), .Y(n_125) );
AND2x4_ASAP7_75t_L g132 ( .A(n_127), .B(n_133), .Y(n_132) );
AND2x4_ASAP7_75t_L g165 ( .A(n_128), .B(n_166), .Y(n_165) );
INVx2_ASAP7_75t_L g130 ( .A(n_131), .Y(n_130) );
INVx1_ASAP7_75t_L g131 ( .A(n_132), .Y(n_131) );
AND2x4_ASAP7_75t_L g174 ( .A(n_133), .B(n_165), .Y(n_174) );
INVx3_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
INVx3_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
AND2x4_ASAP7_75t_L g160 ( .A(n_137), .B(n_161), .Y(n_160) );
AND2x4_ASAP7_75t_L g180 ( .A(n_137), .B(n_167), .Y(n_180) );
BUFx6f_ASAP7_75t_L g141 ( .A(n_142), .Y(n_141) );
BUFx2_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
AND2x4_ASAP7_75t_L g144 ( .A(n_145), .B(n_148), .Y(n_144) );
HB1xp67_ASAP7_75t_L g205 ( .A(n_147), .Y(n_205) );
NAND4xp25_ASAP7_75t_L g151 ( .A(n_152), .B(n_162), .C(n_171), .D(n_177), .Y(n_151) );
BUFx6f_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
INVx2_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
INVx2_ASAP7_75t_L g161 ( .A(n_156), .Y(n_161) );
INVx1_ASAP7_75t_L g168 ( .A(n_157), .Y(n_168) );
INVx3_ASAP7_75t_L g158 ( .A(n_159), .Y(n_158) );
INVx6_ASAP7_75t_L g159 ( .A(n_160), .Y(n_159) );
AND2x4_ASAP7_75t_L g170 ( .A(n_161), .B(n_165), .Y(n_170) );
BUFx12f_ASAP7_75t_L g163 ( .A(n_164), .Y(n_163) );
AND2x4_ASAP7_75t_L g164 ( .A(n_165), .B(n_167), .Y(n_164) );
BUFx6f_ASAP7_75t_L g169 ( .A(n_170), .Y(n_169) );
INVx1_ASAP7_75t_L g172 ( .A(n_173), .Y(n_172) );
INVx3_ASAP7_75t_L g173 ( .A(n_174), .Y(n_173) );
BUFx6f_ASAP7_75t_L g175 ( .A(n_176), .Y(n_175) );
INVx2_ASAP7_75t_L g178 ( .A(n_179), .Y(n_178) );
INVx8_ASAP7_75t_L g179 ( .A(n_180), .Y(n_179) );
BUFx6f_ASAP7_75t_L g181 ( .A(n_182), .Y(n_181) );
CKINVDCx5p33_ASAP7_75t_R g183 ( .A(n_184), .Y(n_183) );
HB1xp67_ASAP7_75t_L g184 ( .A(n_185), .Y(n_184) );
OAI22xp5_ASAP7_75t_L g186 ( .A1(n_187), .A2(n_188), .B1(n_193), .B2(n_194), .Y(n_186) );
CKINVDCx20_ASAP7_75t_R g187 ( .A(n_188), .Y(n_187) );
OAI22xp5_ASAP7_75t_L g188 ( .A1(n_189), .A2(n_190), .B1(n_191), .B2(n_192), .Y(n_188) );
CKINVDCx5p33_ASAP7_75t_R g189 ( .A(n_190), .Y(n_189) );
CKINVDCx5p33_ASAP7_75t_R g191 ( .A(n_192), .Y(n_191) );
CKINVDCx20_ASAP7_75t_R g193 ( .A(n_194), .Y(n_193) );
AOI22xp5_ASAP7_75t_L g194 ( .A1(n_195), .A2(n_196), .B1(n_197), .B2(n_198), .Y(n_194) );
CKINVDCx5p33_ASAP7_75t_R g198 ( .A(n_195), .Y(n_198) );
CKINVDCx20_ASAP7_75t_R g197 ( .A(n_196), .Y(n_197) );
BUFx2_ASAP7_75t_L g199 ( .A(n_200), .Y(n_199) );
CKINVDCx5p33_ASAP7_75t_R g200 ( .A(n_201), .Y(n_200) );
NAND2xp5_ASAP7_75t_L g201 ( .A(n_202), .B(n_210), .Y(n_201) );
INVxp67_ASAP7_75t_SL g202 ( .A(n_203), .Y(n_202) );
AND2x2_ASAP7_75t_L g643 ( .A(n_203), .B(n_210), .Y(n_643) );
AOI211xp5_ASAP7_75t_L g203 ( .A1(n_204), .A2(n_205), .B(n_206), .C(n_209), .Y(n_203) );
NOR2xp33_ASAP7_75t_L g206 ( .A(n_207), .B(n_208), .Y(n_206) );
NOR2xp33_ASAP7_75t_L g210 ( .A(n_211), .B(n_214), .Y(n_210) );
OR2x2_ASAP7_75t_L g648 ( .A(n_211), .B(n_215), .Y(n_648) );
INVx1_ASAP7_75t_L g651 ( .A(n_211), .Y(n_651) );
NAND2xp5_ASAP7_75t_L g652 ( .A(n_211), .B(n_214), .Y(n_652) );
HB1xp67_ASAP7_75t_L g211 ( .A(n_212), .Y(n_211) );
HB1xp67_ASAP7_75t_L g212 ( .A(n_213), .Y(n_212) );
INVx1_ASAP7_75t_L g214 ( .A(n_215), .Y(n_214) );
BUFx2_ASAP7_75t_L g216 ( .A(n_217), .Y(n_216) );
AND2x2_ASAP7_75t_L g217 ( .A(n_218), .B(n_220), .Y(n_217) );
BUFx6f_ASAP7_75t_L g218 ( .A(n_219), .Y(n_218) );
AND2x2_ASAP7_75t_L g287 ( .A(n_219), .B(n_288), .Y(n_287) );
INVx3_ASAP7_75t_L g320 ( .A(n_219), .Y(n_320) );
AND2x2_ASAP7_75t_L g398 ( .A(n_219), .B(n_399), .Y(n_398) );
OA21x2_ASAP7_75t_L g650 ( .A1(n_220), .A2(n_651), .B(n_652), .Y(n_650) );
NOR2xp33_ASAP7_75t_L g220 ( .A(n_221), .B(n_225), .Y(n_220) );
HB1xp67_ASAP7_75t_L g221 ( .A(n_222), .Y(n_221) );
NOR2xp33_ASAP7_75t_L g387 ( .A(n_222), .B(n_273), .Y(n_387) );
INVx4_ASAP7_75t_L g222 ( .A(n_223), .Y(n_222) );
OAI22xp5_ASAP7_75t_L g240 ( .A1(n_223), .A2(n_241), .B1(n_244), .B2(n_249), .Y(n_240) );
AOI21xp5_ASAP7_75t_L g331 ( .A1(n_223), .A2(n_332), .B(n_334), .Y(n_331) );
BUFx6f_ASAP7_75t_L g223 ( .A(n_224), .Y(n_223) );
BUFx6f_ASAP7_75t_L g250 ( .A(n_224), .Y(n_250) );
INVx4_ASAP7_75t_L g267 ( .A(n_224), .Y(n_267) );
INVx3_ASAP7_75t_L g300 ( .A(n_224), .Y(n_300) );
INVx1_ASAP7_75t_L g361 ( .A(n_224), .Y(n_361) );
HB1xp67_ASAP7_75t_L g225 ( .A(n_226), .Y(n_225) );
INVx1_ASAP7_75t_L g226 ( .A(n_227), .Y(n_226) );
INVx2_ASAP7_75t_L g272 ( .A(n_227), .Y(n_272) );
INVxp67_ASAP7_75t_SL g359 ( .A(n_227), .Y(n_359) );
INVx2_ASAP7_75t_L g227 ( .A(n_228), .Y(n_227) );
INVx6_ASAP7_75t_L g243 ( .A(n_228), .Y(n_243) );
INVx3_ASAP7_75t_L g248 ( .A(n_228), .Y(n_248) );
INVx2_ASAP7_75t_L g358 ( .A(n_228), .Y(n_358) );
INVx1_ASAP7_75t_L g229 ( .A(n_230), .Y(n_229) );
HB1xp67_ASAP7_75t_L g230 ( .A(n_231), .Y(n_230) );
INVxp67_ASAP7_75t_SL g231 ( .A(n_232), .Y(n_231) );
OR2x2_ASAP7_75t_L g232 ( .A(n_233), .B(n_543), .Y(n_232) );
NAND4xp25_ASAP7_75t_L g233 ( .A(n_234), .B(n_439), .C(n_486), .D(n_518), .Y(n_233) );
NOR2xp33_ASAP7_75t_L g234 ( .A(n_235), .B(n_423), .Y(n_234) );
NAND2xp5_ASAP7_75t_L g235 ( .A(n_236), .B(n_393), .Y(n_235) );
OAI21xp33_ASAP7_75t_SL g236 ( .A1(n_237), .A2(n_303), .B(n_325), .Y(n_236) );
AND2x4_ASAP7_75t_L g237 ( .A(n_238), .B(n_258), .Y(n_237) );
INVx1_ASAP7_75t_L g438 ( .A(n_238), .Y(n_438) );
AND2x2_ASAP7_75t_SL g443 ( .A(n_238), .B(n_307), .Y(n_443) );
AND2x2_ASAP7_75t_L g522 ( .A(n_238), .B(n_416), .Y(n_522) );
OR2x2_ASAP7_75t_L g546 ( .A(n_238), .B(n_547), .Y(n_546) );
AND2x2_ASAP7_75t_L g564 ( .A(n_238), .B(n_446), .Y(n_564) );
AND2x2_ASAP7_75t_L g586 ( .A(n_238), .B(n_587), .Y(n_586) );
INVx2_ASAP7_75t_L g602 ( .A(n_238), .Y(n_602) );
BUFx8_ASAP7_75t_L g238 ( .A(n_239), .Y(n_238) );
INVx2_ASAP7_75t_L g470 ( .A(n_239), .Y(n_470) );
AND2x2_ASAP7_75t_L g618 ( .A(n_239), .B(n_469), .Y(n_618) );
NAND2xp5_ASAP7_75t_L g281 ( .A(n_242), .B(n_282), .Y(n_281) );
INVx2_ASAP7_75t_SL g242 ( .A(n_243), .Y(n_242) );
INVx2_ASAP7_75t_L g264 ( .A(n_243), .Y(n_264) );
INVx1_ASAP7_75t_L g298 ( .A(n_243), .Y(n_298) );
INVx2_ASAP7_75t_L g343 ( .A(n_243), .Y(n_343) );
OAI22xp33_ASAP7_75t_L g388 ( .A1(n_245), .A2(n_343), .B1(n_389), .B2(n_390), .Y(n_388) );
INVx2_ASAP7_75t_L g245 ( .A(n_246), .Y(n_245) );
INVx2_ASAP7_75t_L g335 ( .A(n_246), .Y(n_335) );
INVx1_ASAP7_75t_L g339 ( .A(n_246), .Y(n_339) );
INVx2_ASAP7_75t_L g348 ( .A(n_246), .Y(n_348) );
INVx2_ASAP7_75t_L g371 ( .A(n_246), .Y(n_371) );
INVx1_ASAP7_75t_L g366 ( .A(n_247), .Y(n_366) );
INVx2_ASAP7_75t_L g247 ( .A(n_248), .Y(n_247) );
INVx2_ASAP7_75t_L g295 ( .A(n_248), .Y(n_295) );
INVx1_ASAP7_75t_L g333 ( .A(n_248), .Y(n_333) );
INVx1_ASAP7_75t_L g349 ( .A(n_248), .Y(n_349) );
INVx1_ASAP7_75t_L g249 ( .A(n_250), .Y(n_249) );
INVx1_ASAP7_75t_L g296 ( .A(n_250), .Y(n_296) );
A2O1A1Ixp33_ASAP7_75t_L g314 ( .A1(n_250), .A2(n_315), .B(n_316), .C(n_317), .Y(n_314) );
NAND2xp5_ASAP7_75t_SL g350 ( .A(n_250), .B(n_351), .Y(n_350) );
A2O1A1Ixp33_ASAP7_75t_L g365 ( .A1(n_250), .A2(n_366), .B(n_367), .C(n_368), .Y(n_365) );
AO31x2_ASAP7_75t_L g260 ( .A1(n_251), .A2(n_261), .A3(n_275), .B(n_283), .Y(n_260) );
INVx2_ASAP7_75t_L g400 ( .A(n_251), .Y(n_400) );
BUFx3_ASAP7_75t_L g251 ( .A(n_252), .Y(n_251) );
NOR2xp33_ASAP7_75t_L g283 ( .A(n_252), .B(n_284), .Y(n_283) );
NOR2xp33_ASAP7_75t_L g301 ( .A(n_252), .B(n_302), .Y(n_301) );
INVx3_ASAP7_75t_L g329 ( .A(n_252), .Y(n_329) );
INVx2_ASAP7_75t_L g252 ( .A(n_253), .Y(n_252) );
INVx4_ASAP7_75t_L g290 ( .A(n_253), .Y(n_290) );
BUFx3_ASAP7_75t_L g411 ( .A(n_253), .Y(n_411) );
INVxp67_ASAP7_75t_L g376 ( .A(n_255), .Y(n_376) );
INVx1_ASAP7_75t_L g255 ( .A(n_256), .Y(n_255) );
NOR2xp33_ASAP7_75t_L g391 ( .A(n_256), .B(n_392), .Y(n_391) );
INVx1_ASAP7_75t_L g256 ( .A(n_257), .Y(n_256) );
NOR2xp33_ASAP7_75t_L g319 ( .A(n_257), .B(n_320), .Y(n_319) );
INVx1_ASAP7_75t_L g323 ( .A(n_257), .Y(n_323) );
NOR2xp33_ASAP7_75t_L g344 ( .A(n_257), .B(n_320), .Y(n_344) );
NOR2xp67_ASAP7_75t_L g351 ( .A(n_257), .B(n_320), .Y(n_351) );
BUFx3_ASAP7_75t_L g353 ( .A(n_257), .Y(n_353) );
INVx1_ASAP7_75t_L g399 ( .A(n_257), .Y(n_399) );
AND2x2_ASAP7_75t_L g526 ( .A(n_258), .B(n_527), .Y(n_526) );
AND2x2_ASAP7_75t_L g607 ( .A(n_258), .B(n_463), .Y(n_607) );
INVxp67_ASAP7_75t_SL g623 ( .A(n_258), .Y(n_623) );
AND2x2_ASAP7_75t_L g258 ( .A(n_259), .B(n_285), .Y(n_258) );
INVx1_ASAP7_75t_L g483 ( .A(n_259), .Y(n_483) );
INVx2_ASAP7_75t_SL g580 ( .A(n_259), .Y(n_580) );
NAND2xp5_ASAP7_75t_L g593 ( .A(n_259), .B(n_470), .Y(n_593) );
INVx2_ASAP7_75t_L g259 ( .A(n_260), .Y(n_259) );
INVx1_ASAP7_75t_L g324 ( .A(n_260), .Y(n_324) );
OR2x2_ASAP7_75t_L g403 ( .A(n_260), .B(n_404), .Y(n_403) );
AND2x2_ASAP7_75t_L g416 ( .A(n_260), .B(n_308), .Y(n_416) );
AND2x2_ASAP7_75t_L g446 ( .A(n_260), .B(n_401), .Y(n_446) );
NAND2xp5_ASAP7_75t_L g499 ( .A(n_260), .B(n_404), .Y(n_499) );
AOI221x1_ASAP7_75t_L g261 ( .A1(n_262), .A2(n_265), .B1(n_269), .B2(n_271), .C(n_273), .Y(n_261) );
INVx1_ASAP7_75t_L g262 ( .A(n_263), .Y(n_262) );
INVx1_ASAP7_75t_L g263 ( .A(n_264), .Y(n_263) );
AND2x2_ASAP7_75t_L g265 ( .A(n_266), .B(n_268), .Y(n_265) );
AND2x2_ASAP7_75t_L g269 ( .A(n_266), .B(n_270), .Y(n_269) );
INVx2_ASAP7_75t_L g266 ( .A(n_267), .Y(n_266) );
NOR2xp33_ASAP7_75t_L g341 ( .A(n_267), .B(n_342), .Y(n_341) );
INVx1_ASAP7_75t_L g271 ( .A(n_272), .Y(n_271) );
NOR2xp33_ASAP7_75t_L g381 ( .A(n_273), .B(n_299), .Y(n_381) );
NOR3xp33_ASAP7_75t_L g384 ( .A(n_273), .B(n_299), .C(n_385), .Y(n_384) );
INVx4_ASAP7_75t_L g273 ( .A(n_274), .Y(n_273) );
INVx1_ASAP7_75t_L g275 ( .A(n_276), .Y(n_275) );
INVx3_ASAP7_75t_L g277 ( .A(n_278), .Y(n_277) );
INVx2_ASAP7_75t_L g278 ( .A(n_279), .Y(n_278) );
INVx1_ASAP7_75t_L g318 ( .A(n_279), .Y(n_318) );
INVx2_ASAP7_75t_L g279 ( .A(n_280), .Y(n_279) );
INVx2_ASAP7_75t_L g294 ( .A(n_280), .Y(n_294) );
HB1xp67_ASAP7_75t_L g429 ( .A(n_285), .Y(n_429) );
INVx2_ASAP7_75t_L g462 ( .A(n_285), .Y(n_462) );
AND2x2_ASAP7_75t_L g629 ( .A(n_285), .B(n_401), .Y(n_629) );
INVx1_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
INVx1_ASAP7_75t_L g306 ( .A(n_286), .Y(n_306) );
INVx1_ASAP7_75t_L g404 ( .A(n_286), .Y(n_404) );
AOI21x1_ASAP7_75t_L g286 ( .A1(n_287), .A2(n_291), .B(n_301), .Y(n_286) );
INVx2_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
NOR2xp33_ASAP7_75t_L g364 ( .A(n_289), .B(n_320), .Y(n_364) );
INVx2_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
OAI22xp5_ASAP7_75t_L g291 ( .A1(n_292), .A2(n_296), .B1(n_297), .B2(n_299), .Y(n_291) );
INVx2_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
INVx2_ASAP7_75t_L g316 ( .A(n_294), .Y(n_316) );
INVx1_ASAP7_75t_L g311 ( .A(n_298), .Y(n_311) );
INVx3_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
A2O1A1Ixp33_ASAP7_75t_L g310 ( .A1(n_300), .A2(n_311), .B(n_312), .C(n_313), .Y(n_310) );
A2O1A1Ixp33_ASAP7_75t_L g369 ( .A1(n_300), .A2(n_370), .B(n_371), .C(n_372), .Y(n_369) );
INVx2_ASAP7_75t_L g551 ( .A(n_303), .Y(n_551) );
AND2x2_ASAP7_75t_L g303 ( .A(n_304), .B(n_307), .Y(n_303) );
NAND2x1p5_ASAP7_75t_L g415 ( .A(n_304), .B(n_416), .Y(n_415) );
NAND2xp5_ASAP7_75t_L g501 ( .A(n_304), .B(n_396), .Y(n_501) );
INVx4_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
HB1xp67_ASAP7_75t_SL g441 ( .A(n_305), .Y(n_441) );
AND2x2_ASAP7_75t_L g560 ( .A(n_305), .B(n_446), .Y(n_560) );
AND2x2_ASAP7_75t_L g573 ( .A(n_305), .B(n_307), .Y(n_573) );
INVx2_ASAP7_75t_L g576 ( .A(n_305), .Y(n_576) );
BUFx3_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
INVx1_ASAP7_75t_L g469 ( .A(n_306), .Y(n_469) );
INVx2_ASAP7_75t_L g547 ( .A(n_307), .Y(n_547) );
AND2x4_ASAP7_75t_L g307 ( .A(n_308), .B(n_324), .Y(n_307) );
INVx2_ASAP7_75t_L g401 ( .A(n_308), .Y(n_401) );
INVx1_ASAP7_75t_L g464 ( .A(n_308), .Y(n_464) );
BUFx3_ASAP7_75t_L g482 ( .A(n_308), .Y(n_482) );
AND2x4_ASAP7_75t_L g527 ( .A(n_308), .B(n_470), .Y(n_527) );
INVx3_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
AO31x2_ASAP7_75t_L g309 ( .A1(n_310), .A2(n_314), .A3(n_319), .B(n_321), .Y(n_309) );
NOR2xp67_ASAP7_75t_L g379 ( .A(n_316), .B(n_380), .Y(n_379) );
NOR2xp33_ASAP7_75t_L g321 ( .A(n_322), .B(n_323), .Y(n_321) );
NOR2xp33_ASAP7_75t_SL g373 ( .A(n_323), .B(n_374), .Y(n_373) );
AND2x2_ASAP7_75t_L g325 ( .A(n_326), .B(n_362), .Y(n_325) );
AND2x2_ASAP7_75t_L g589 ( .A(n_326), .B(n_421), .Y(n_589) );
AND2x2_ASAP7_75t_L g326 ( .A(n_327), .B(n_345), .Y(n_326) );
INVx2_ASAP7_75t_L g413 ( .A(n_327), .Y(n_413) );
INVx1_ASAP7_75t_L g436 ( .A(n_327), .Y(n_436) );
AND2x2_ASAP7_75t_L g452 ( .A(n_327), .B(n_453), .Y(n_452) );
INVx1_ASAP7_75t_L g515 ( .A(n_327), .Y(n_515) );
HB1xp67_ASAP7_75t_L g626 ( .A(n_327), .Y(n_626) );
AND2x4_ASAP7_75t_L g327 ( .A(n_328), .B(n_330), .Y(n_327) );
OAI21xp5_ASAP7_75t_L g330 ( .A1(n_331), .A2(n_336), .B(n_344), .Y(n_330) );
OAI21xp5_ASAP7_75t_L g336 ( .A1(n_337), .A2(n_338), .B(n_340), .Y(n_336) );
INVx1_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
NAND2xp5_ASAP7_75t_L g340 ( .A(n_341), .B(n_343), .Y(n_340) );
AND2x2_ASAP7_75t_L g412 ( .A(n_345), .B(n_413), .Y(n_412) );
INVx1_ASAP7_75t_L g432 ( .A(n_345), .Y(n_432) );
INVx2_ASAP7_75t_L g450 ( .A(n_345), .Y(n_450) );
INVx1_ASAP7_75t_L g474 ( .A(n_345), .Y(n_474) );
NAND2x1p5_ASAP7_75t_L g345 ( .A(n_346), .B(n_354), .Y(n_345) );
AND2x2_ASAP7_75t_SL g420 ( .A(n_346), .B(n_354), .Y(n_420) );
OA21x2_ASAP7_75t_L g346 ( .A1(n_347), .A2(n_350), .B(n_352), .Y(n_346) );
NAND2xp5_ASAP7_75t_L g360 ( .A(n_351), .B(n_361), .Y(n_360) );
OR2x2_ASAP7_75t_L g354 ( .A(n_355), .B(n_360), .Y(n_354) );
INVx1_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
INVx2_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
INVx1_ASAP7_75t_L g383 ( .A(n_358), .Y(n_383) );
INVx1_ASAP7_75t_L g500 ( .A(n_362), .Y(n_500) );
AND2x2_ASAP7_75t_L g549 ( .A(n_362), .B(n_550), .Y(n_549) );
AND2x2_ASAP7_75t_L g637 ( .A(n_362), .B(n_412), .Y(n_637) );
AND2x2_ASAP7_75t_L g362 ( .A(n_363), .B(n_375), .Y(n_362) );
OR2x2_ASAP7_75t_L g408 ( .A(n_363), .B(n_409), .Y(n_408) );
INVx2_ASAP7_75t_L g422 ( .A(n_363), .Y(n_422) );
INVx2_ASAP7_75t_L g453 ( .A(n_363), .Y(n_453) );
HB1xp67_ASAP7_75t_L g479 ( .A(n_363), .Y(n_479) );
INVx1_ASAP7_75t_L g513 ( .A(n_363), .Y(n_513) );
INVx1_ASAP7_75t_L g559 ( .A(n_363), .Y(n_559) );
AO31x2_ASAP7_75t_L g363 ( .A1(n_364), .A2(n_365), .A3(n_369), .B(n_373), .Y(n_363) );
INVx1_ASAP7_75t_L g654 ( .A(n_367), .Y(n_654) );
OR2x2_ASAP7_75t_L g458 ( .A(n_375), .B(n_413), .Y(n_458) );
AND2x2_ASAP7_75t_L g514 ( .A(n_375), .B(n_515), .Y(n_514) );
AND2x2_ASAP7_75t_L g582 ( .A(n_375), .B(n_583), .Y(n_582) );
AND2x2_ASAP7_75t_L g605 ( .A(n_375), .B(n_450), .Y(n_605) );
AO21x2_ASAP7_75t_L g375 ( .A1(n_376), .A2(n_377), .B(n_391), .Y(n_375) );
AO21x2_ASAP7_75t_L g409 ( .A1(n_377), .A2(n_391), .B(n_410), .Y(n_409) );
NAND2xp5_ASAP7_75t_L g377 ( .A(n_378), .B(n_386), .Y(n_377) );
AOI22xp5_ASAP7_75t_L g378 ( .A1(n_379), .A2(n_381), .B1(n_382), .B2(n_384), .Y(n_378) );
INVx1_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
NAND2xp5_ASAP7_75t_L g386 ( .A(n_387), .B(n_388), .Y(n_386) );
AOI22xp33_ASAP7_75t_SL g393 ( .A1(n_394), .A2(n_405), .B1(n_414), .B2(n_417), .Y(n_393) );
NOR2xp33_ASAP7_75t_L g394 ( .A(n_395), .B(n_402), .Y(n_394) );
OAI221xp5_ASAP7_75t_L g599 ( .A1(n_395), .A2(n_535), .B1(n_600), .B2(n_603), .C(n_606), .Y(n_599) );
INVx4_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
AND2x4_ASAP7_75t_L g541 ( .A(n_396), .B(n_542), .Y(n_541) );
NOR2xp33_ASAP7_75t_L g622 ( .A(n_396), .B(n_623), .Y(n_622) );
AND2x4_ASAP7_75t_L g396 ( .A(n_397), .B(n_401), .Y(n_396) );
INVx1_ASAP7_75t_L g426 ( .A(n_397), .Y(n_426) );
INVx1_ASAP7_75t_L g465 ( .A(n_397), .Y(n_465) );
AND2x4_ASAP7_75t_L g493 ( .A(n_397), .B(n_482), .Y(n_493) );
AND2x2_ASAP7_75t_L g517 ( .A(n_402), .B(n_481), .Y(n_517) );
INVx2_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
INVx2_ASAP7_75t_L g542 ( .A(n_403), .Y(n_542) );
HB1xp67_ASAP7_75t_L g494 ( .A(n_404), .Y(n_494) );
INVx2_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
NAND2xp67_ASAP7_75t_L g406 ( .A(n_407), .B(n_412), .Y(n_406) );
INVx2_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
OR2x2_ASAP7_75t_L g508 ( .A(n_408), .B(n_473), .Y(n_508) );
AND2x2_ASAP7_75t_L g421 ( .A(n_409), .B(n_422), .Y(n_421) );
INVx2_ASAP7_75t_L g451 ( .A(n_409), .Y(n_451) );
BUFx2_ASAP7_75t_L g485 ( .A(n_409), .Y(n_485) );
INVx3_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
AND2x2_ASAP7_75t_L g529 ( .A(n_412), .B(n_530), .Y(n_529) );
NAND2xp5_ASAP7_75t_L g539 ( .A(n_412), .B(n_485), .Y(n_539) );
AND2x2_ASAP7_75t_L g590 ( .A(n_412), .B(n_484), .Y(n_590) );
AND2x2_ASAP7_75t_L g613 ( .A(n_412), .B(n_503), .Y(n_613) );
INVx3_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
AND2x2_ASAP7_75t_L g425 ( .A(n_416), .B(n_426), .Y(n_425) );
INVx2_ASAP7_75t_L g467 ( .A(n_416), .Y(n_467) );
INVx2_ASAP7_75t_L g533 ( .A(n_416), .Y(n_533) );
AOI22xp5_ASAP7_75t_L g606 ( .A1(n_417), .A2(n_607), .B1(n_608), .B2(n_609), .Y(n_606) );
INVx2_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
NAND2x1p5_ASAP7_75t_L g418 ( .A(n_419), .B(n_421), .Y(n_418) );
NAND2xp5_ASAP7_75t_L g502 ( .A(n_419), .B(n_503), .Y(n_502) );
INVx1_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
AND2x2_ASAP7_75t_L g558 ( .A(n_420), .B(n_436), .Y(n_558) );
INVx2_ASAP7_75t_L g583 ( .A(n_420), .Y(n_583) );
AND2x2_ASAP7_75t_L g616 ( .A(n_420), .B(n_436), .Y(n_616) );
AND2x4_ASAP7_75t_L g428 ( .A(n_421), .B(n_429), .Y(n_428) );
INVx2_ASAP7_75t_L g555 ( .A(n_421), .Y(n_555) );
INVxp67_ASAP7_75t_SL g457 ( .A(n_422), .Y(n_457) );
HB1xp67_ASAP7_75t_L g562 ( .A(n_422), .Y(n_562) );
OAI32xp33_ASAP7_75t_L g423 ( .A1(n_424), .A2(n_427), .A3(n_430), .B1(n_433), .B2(n_437), .Y(n_423) );
OAI22xp33_ASAP7_75t_L g632 ( .A1(n_424), .A2(n_633), .B1(n_634), .B2(n_636), .Y(n_632) );
INVx2_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
INVx1_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
NAND2xp5_ASAP7_75t_L g433 ( .A(n_428), .B(n_434), .Y(n_433) );
INVx1_ASAP7_75t_L g532 ( .A(n_429), .Y(n_532) );
INVx1_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
AOI311xp33_ASAP7_75t_L g518 ( .A1(n_431), .A2(n_519), .A3(n_520), .B(n_523), .C(n_534), .Y(n_518) );
BUFx3_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
AND2x2_ASAP7_75t_L g511 ( .A(n_432), .B(n_512), .Y(n_511) );
INVx2_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
NAND5xp2_ASAP7_75t_L g477 ( .A(n_435), .B(n_478), .C(n_480), .D(n_483), .E(n_484), .Y(n_477) );
INVx1_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
INVx1_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
NOR3xp33_ASAP7_75t_L g439 ( .A(n_440), .B(n_454), .C(n_476), .Y(n_439) );
AOI31xp33_ASAP7_75t_L g440 ( .A1(n_441), .A2(n_442), .A3(n_444), .B(n_447), .Y(n_440) );
INVx2_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
INVx1_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
HB1xp67_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
AND2x2_ASAP7_75t_L g601 ( .A(n_446), .B(n_602), .Y(n_601) );
AND2x2_ASAP7_75t_L g617 ( .A(n_446), .B(n_618), .Y(n_617) );
AND2x2_ASAP7_75t_L g635 ( .A(n_446), .B(n_462), .Y(n_635) );
INVx1_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
AND2x2_ASAP7_75t_L g448 ( .A(n_449), .B(n_452), .Y(n_448) );
AND2x4_ASAP7_75t_L g624 ( .A(n_449), .B(n_625), .Y(n_624) );
AND2x2_ASAP7_75t_L g449 ( .A(n_450), .B(n_451), .Y(n_449) );
HB1xp67_ASAP7_75t_L g537 ( .A(n_450), .Y(n_537) );
BUFx2_ASAP7_75t_L g550 ( .A(n_450), .Y(n_550) );
AND2x4_ASAP7_75t_L g503 ( .A(n_451), .B(n_504), .Y(n_503) );
OR2x2_ASAP7_75t_L g563 ( .A(n_451), .B(n_515), .Y(n_563) );
AND2x2_ASAP7_75t_L g604 ( .A(n_452), .B(n_605), .Y(n_604) );
AND2x2_ASAP7_75t_L g610 ( .A(n_452), .B(n_474), .Y(n_610) );
INVx1_ASAP7_75t_L g504 ( .A(n_453), .Y(n_504) );
OAI22xp5_ASAP7_75t_L g454 ( .A1(n_455), .A2(n_459), .B1(n_466), .B2(n_471), .Y(n_454) );
HB1xp67_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
INVx2_ASAP7_75t_L g490 ( .A(n_456), .Y(n_490) );
OAI322xp33_ASAP7_75t_L g495 ( .A1(n_456), .A2(n_496), .A3(n_497), .B1(n_500), .B2(n_501), .C1(n_502), .C2(n_505), .Y(n_495) );
OR2x6_ASAP7_75t_L g456 ( .A(n_457), .B(n_458), .Y(n_456) );
INVxp67_ASAP7_75t_L g475 ( .A(n_458), .Y(n_475) );
INVxp67_ASAP7_75t_SL g538 ( .A(n_458), .Y(n_538) );
INVx1_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
AND2x2_ASAP7_75t_L g460 ( .A(n_461), .B(n_463), .Y(n_460) );
INVx1_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
BUFx3_ASAP7_75t_L g521 ( .A(n_462), .Y(n_521) );
AND2x2_ASAP7_75t_L g608 ( .A(n_462), .B(n_481), .Y(n_608) );
INVx1_ASAP7_75t_L g496 ( .A(n_463), .Y(n_496) );
AND2x4_ASAP7_75t_SL g463 ( .A(n_464), .B(n_465), .Y(n_463) );
OR2x2_ASAP7_75t_L g466 ( .A(n_467), .B(n_468), .Y(n_466) );
INVx1_ASAP7_75t_L g506 ( .A(n_468), .Y(n_506) );
NAND2xp5_ASAP7_75t_L g468 ( .A(n_469), .B(n_470), .Y(n_468) );
AND2x2_ASAP7_75t_L g579 ( .A(n_470), .B(n_580), .Y(n_579) );
INVx3_ASAP7_75t_L g471 ( .A(n_472), .Y(n_471) );
AND2x4_ASAP7_75t_L g472 ( .A(n_473), .B(n_475), .Y(n_472) );
AND2x2_ASAP7_75t_L g478 ( .A(n_473), .B(n_479), .Y(n_478) );
INVx1_ASAP7_75t_L g489 ( .A(n_473), .Y(n_489) );
INVx2_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
INVxp67_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
INVx1_ASAP7_75t_L g480 ( .A(n_481), .Y(n_480) );
NOR2xp33_ASAP7_75t_L g575 ( .A(n_481), .B(n_576), .Y(n_575) );
INVx2_ASAP7_75t_SL g481 ( .A(n_482), .Y(n_481) );
INVx2_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
AOI211xp5_ASAP7_75t_L g486 ( .A1(n_487), .A2(n_491), .B(n_495), .C(n_507), .Y(n_486) );
AND2x4_ASAP7_75t_L g487 ( .A(n_488), .B(n_490), .Y(n_487) );
INVxp67_ASAP7_75t_L g488 ( .A(n_489), .Y(n_488) );
INVx1_ASAP7_75t_L g491 ( .A(n_492), .Y(n_491) );
NAND2xp5_ASAP7_75t_L g492 ( .A(n_493), .B(n_494), .Y(n_492) );
OR2x2_ASAP7_75t_L g620 ( .A(n_494), .B(n_593), .Y(n_620) );
OAI211xp5_ASAP7_75t_L g611 ( .A1(n_496), .A2(n_612), .B(n_614), .C(n_621), .Y(n_611) );
INVx2_ASAP7_75t_L g497 ( .A(n_498), .Y(n_497) );
INVx1_ASAP7_75t_L g498 ( .A(n_499), .Y(n_498) );
INVx1_ASAP7_75t_L g587 ( .A(n_499), .Y(n_587) );
INVx1_ASAP7_75t_L g519 ( .A(n_503), .Y(n_519) );
AND2x2_ASAP7_75t_L g569 ( .A(n_503), .B(n_550), .Y(n_569) );
AND2x4_ASAP7_75t_L g596 ( .A(n_503), .B(n_597), .Y(n_596) );
AND2x2_ASAP7_75t_L g615 ( .A(n_503), .B(n_616), .Y(n_615) );
INVx1_ASAP7_75t_L g505 ( .A(n_506), .Y(n_505) );
AOI21xp33_ASAP7_75t_L g507 ( .A1(n_508), .A2(n_509), .B(n_516), .Y(n_507) );
INVx2_ASAP7_75t_L g509 ( .A(n_510), .Y(n_509) );
AND2x4_ASAP7_75t_L g510 ( .A(n_511), .B(n_514), .Y(n_510) );
INVxp67_ASAP7_75t_L g530 ( .A(n_512), .Y(n_530) );
HB1xp67_ASAP7_75t_L g572 ( .A(n_512), .Y(n_572) );
AND2x2_ASAP7_75t_L g631 ( .A(n_512), .B(n_626), .Y(n_631) );
INVx2_ASAP7_75t_L g512 ( .A(n_513), .Y(n_512) );
INVx1_ASAP7_75t_L g524 ( .A(n_514), .Y(n_524) );
AND2x2_ASAP7_75t_L g567 ( .A(n_515), .B(n_559), .Y(n_567) );
INVx1_ASAP7_75t_L g597 ( .A(n_515), .Y(n_597) );
INVx2_ASAP7_75t_L g516 ( .A(n_517), .Y(n_516) );
AND2x2_ASAP7_75t_L g520 ( .A(n_521), .B(n_522), .Y(n_520) );
OAI22xp5_ASAP7_75t_L g523 ( .A1(n_524), .A2(n_525), .B1(n_528), .B2(n_531), .Y(n_523) );
INVx2_ASAP7_75t_SL g525 ( .A(n_526), .Y(n_525) );
INVx1_ASAP7_75t_L g528 ( .A(n_529), .Y(n_528) );
OR2x2_ASAP7_75t_L g531 ( .A(n_532), .B(n_533), .Y(n_531) );
AOI21xp5_ASAP7_75t_L g534 ( .A1(n_535), .A2(n_539), .B(n_540), .Y(n_534) );
INVx1_ASAP7_75t_L g535 ( .A(n_536), .Y(n_535) );
AND2x4_ASAP7_75t_L g536 ( .A(n_537), .B(n_538), .Y(n_536) );
INVx1_ASAP7_75t_L g595 ( .A(n_537), .Y(n_595) );
INVx1_ASAP7_75t_L g540 ( .A(n_541), .Y(n_540) );
NAND2xp5_ASAP7_75t_L g543 ( .A(n_544), .B(n_598), .Y(n_543) );
NOR3xp33_ASAP7_75t_L g544 ( .A(n_545), .B(n_565), .C(n_584), .Y(n_544) );
OAI221xp5_ASAP7_75t_L g545 ( .A1(n_546), .A2(n_548), .B1(n_551), .B2(n_552), .C(n_556), .Y(n_545) );
OAI211xp5_ASAP7_75t_L g565 ( .A1(n_546), .A2(n_566), .B(n_568), .C(n_574), .Y(n_565) );
INVx1_ASAP7_75t_L g548 ( .A(n_549), .Y(n_548) );
INVx1_ASAP7_75t_L g554 ( .A(n_550), .Y(n_554) );
INVxp67_ASAP7_75t_SL g552 ( .A(n_553), .Y(n_552) );
NOR2x1p5_ASAP7_75t_L g553 ( .A(n_554), .B(n_555), .Y(n_553) );
AOI22xp5_ASAP7_75t_L g556 ( .A1(n_557), .A2(n_560), .B1(n_561), .B2(n_564), .Y(n_556) );
AND2x2_ASAP7_75t_L g557 ( .A(n_558), .B(n_559), .Y(n_557) );
NAND2xp5_ASAP7_75t_L g571 ( .A(n_558), .B(n_572), .Y(n_571) );
NOR2xp67_ASAP7_75t_L g561 ( .A(n_562), .B(n_563), .Y(n_561) );
INVx1_ASAP7_75t_L g566 ( .A(n_567), .Y(n_566) );
AND2x4_ASAP7_75t_L g581 ( .A(n_567), .B(n_582), .Y(n_581) );
OAI21xp33_ASAP7_75t_L g568 ( .A1(n_569), .A2(n_570), .B(n_573), .Y(n_568) );
INVx2_ASAP7_75t_L g570 ( .A(n_571), .Y(n_570) );
OAI21xp33_ASAP7_75t_L g574 ( .A1(n_575), .A2(n_577), .B(n_581), .Y(n_574) );
INVx1_ASAP7_75t_L g577 ( .A(n_578), .Y(n_577) );
NAND2xp5_ASAP7_75t_L g627 ( .A(n_578), .B(n_628), .Y(n_627) );
INVx1_ASAP7_75t_L g578 ( .A(n_579), .Y(n_578) );
OAI22xp33_ASAP7_75t_SL g584 ( .A1(n_585), .A2(n_588), .B1(n_591), .B2(n_594), .Y(n_584) );
INVx2_ASAP7_75t_L g585 ( .A(n_586), .Y(n_585) );
NOR2xp33_ASAP7_75t_L g588 ( .A(n_589), .B(n_590), .Y(n_588) );
AOI22xp5_ASAP7_75t_L g614 ( .A1(n_590), .A2(n_615), .B1(n_617), .B2(n_619), .Y(n_614) );
INVx1_ASAP7_75t_L g591 ( .A(n_592), .Y(n_591) );
INVxp67_ASAP7_75t_SL g592 ( .A(n_593), .Y(n_592) );
NAND2xp5_ASAP7_75t_L g594 ( .A(n_595), .B(n_596), .Y(n_594) );
NOR3xp33_ASAP7_75t_L g598 ( .A(n_599), .B(n_611), .C(n_632), .Y(n_598) );
INVx2_ASAP7_75t_L g600 ( .A(n_601), .Y(n_600) );
INVx1_ASAP7_75t_L g603 ( .A(n_604), .Y(n_603) );
AND2x4_ASAP7_75t_L g630 ( .A(n_605), .B(n_631), .Y(n_630) );
BUFx2_ASAP7_75t_L g609 ( .A(n_610), .Y(n_609) );
INVx2_ASAP7_75t_L g612 ( .A(n_613), .Y(n_612) );
INVx2_ASAP7_75t_L g633 ( .A(n_615), .Y(n_633) );
INVx2_ASAP7_75t_L g619 ( .A(n_620), .Y(n_619) );
AOI22xp5_ASAP7_75t_L g621 ( .A1(n_622), .A2(n_624), .B1(n_627), .B2(n_630), .Y(n_621) );
INVx1_ASAP7_75t_L g625 ( .A(n_626), .Y(n_625) );
INVx1_ASAP7_75t_L g628 ( .A(n_629), .Y(n_628) );
INVx1_ASAP7_75t_L g634 ( .A(n_635), .Y(n_634) );
INVx2_ASAP7_75t_L g636 ( .A(n_637), .Y(n_636) );
OAI222xp33_ASAP7_75t_L g638 ( .A1(n_639), .A2(n_642), .B1(n_644), .B2(n_647), .C1(n_649), .C2(n_653), .Y(n_638) );
CKINVDCx20_ASAP7_75t_R g641 ( .A(n_640), .Y(n_641) );
INVx1_ASAP7_75t_SL g642 ( .A(n_643), .Y(n_642) );
INVx1_ASAP7_75t_L g644 ( .A(n_645), .Y(n_644) );
BUFx2_ASAP7_75t_L g647 ( .A(n_648), .Y(n_647) );
BUFx2_ASAP7_75t_L g649 ( .A(n_650), .Y(n_649) );
CKINVDCx20_ASAP7_75t_R g653 ( .A(n_654), .Y(n_653) );
endmodule