module real_jpeg_8254_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_68;
wire n_146;
wire n_83;
wire n_78;
wire n_166;
wire n_176;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_64;
wire n_177;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_197;
wire n_40;
wire n_173;
wire n_105;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_200;
wire n_48;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_188;
wire n_139;
wire n_142;
wire n_175;
wire n_178;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_136;
wire n_44;
wire n_28;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_160;
wire n_172;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_165;
wire n_134;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_192;
wire n_198;
wire n_100;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_117;
wire n_193;
wire n_99;
wire n_86;
wire n_150;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_70;
wire n_30;
wire n_158;
wire n_149;
wire n_144;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_185;
wire n_55;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_202;
wire n_167;
wire n_179;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_181;
wire n_85;
wire n_101;
wire n_182;
wire n_96;
wire n_89;

BUFx24_ASAP7_75t_L g66 ( 
.A(n_0),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_L g55 ( 
.A1(n_1),
.A2(n_38),
.B1(n_39),
.B2(n_56),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_1),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_1),
.A2(n_56),
.B1(n_60),
.B2(n_69),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_L g96 ( 
.A1(n_1),
.A2(n_56),
.B1(n_65),
.B2(n_66),
.Y(n_96)
);

OAI22xp33_ASAP7_75t_SL g144 ( 
.A1(n_1),
.A2(n_26),
.B1(n_27),
.B2(n_56),
.Y(n_144)
);

INVx2_ASAP7_75t_SL g62 ( 
.A(n_2),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g64 ( 
.A1(n_2),
.A2(n_62),
.B1(n_65),
.B2(n_66),
.Y(n_64)
);

AOI21xp33_ASAP7_75t_L g101 ( 
.A1(n_2),
.A2(n_10),
.B(n_66),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_L g37 ( 
.A1(n_3),
.A2(n_38),
.B1(n_39),
.B2(n_40),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_3),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_3),
.A2(n_26),
.B1(n_27),
.B2(n_40),
.Y(n_118)
);

BUFx10_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

BUFx10_ASAP7_75t_L g44 ( 
.A(n_6),
.Y(n_44)
);

BUFx6f_ASAP7_75t_SL g79 ( 
.A(n_7),
.Y(n_79)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_8),
.Y(n_39)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_9),
.A2(n_65),
.B1(n_66),
.B2(n_86),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_9),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_9),
.A2(n_26),
.B1(n_27),
.B2(n_86),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_L g171 ( 
.A1(n_9),
.A2(n_38),
.B1(n_39),
.B2(n_86),
.Y(n_171)
);

OAI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_10),
.A2(n_60),
.B1(n_68),
.B2(n_69),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_10),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_10),
.B(n_72),
.Y(n_116)
);

A2O1A1O1Ixp25_ASAP7_75t_L g127 ( 
.A1(n_10),
.A2(n_38),
.B(n_42),
.C(n_128),
.D(n_129),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_10),
.B(n_38),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_10),
.B(n_81),
.Y(n_137)
);

OAI21xp33_ASAP7_75t_L g159 ( 
.A1(n_10),
.A2(n_24),
.B(n_143),
.Y(n_159)
);

A2O1A1O1Ixp25_ASAP7_75t_L g172 ( 
.A1(n_10),
.A2(n_65),
.B(n_77),
.C(n_95),
.D(n_173),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_10),
.B(n_65),
.Y(n_173)
);

BUFx2_ASAP7_75t_L g61 ( 
.A(n_11),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_SL g47 ( 
.A1(n_12),
.A2(n_38),
.B1(n_39),
.B2(n_48),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_12),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_12),
.A2(n_26),
.B1(n_27),
.B2(n_48),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g31 ( 
.A1(n_13),
.A2(n_26),
.B1(n_27),
.B2(n_32),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_13),
.Y(n_32)
);

AOI22xp5_ASAP7_75t_L g34 ( 
.A1(n_14),
.A2(n_26),
.B1(n_27),
.B2(n_35),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_14),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_15),
.A2(n_65),
.B1(n_66),
.B2(n_83),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_15),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_15),
.A2(n_60),
.B1(n_69),
.B2(n_83),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_15),
.A2(n_38),
.B1(n_39),
.B2(n_83),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_SL g149 ( 
.A1(n_15),
.A2(n_26),
.B1(n_27),
.B2(n_83),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_121),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_119),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_19),
.Y(n_18)
);

AND2x2_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_105),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_20),
.B(n_105),
.Y(n_120)
);

XNOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_87),
.Y(n_20)
);

XNOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_50),
.Y(n_21)
);

XOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_36),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_31),
.B1(n_33),
.B2(n_34),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_24),
.A2(n_31),
.B1(n_33),
.B2(n_103),
.Y(n_102)
);

OAI21xp5_ASAP7_75t_SL g141 ( 
.A1(n_24),
.A2(n_142),
.B(n_143),
.Y(n_141)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_25),
.A2(n_30),
.B1(n_104),
.B2(n_118),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_25),
.A2(n_30),
.B1(n_148),
.B2(n_150),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_25),
.B(n_144),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_SL g25 ( 
.A(n_26),
.B(n_30),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_L g46 ( 
.A1(n_26),
.A2(n_27),
.B1(n_43),
.B2(n_44),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_SL g132 ( 
.A(n_26),
.B(n_43),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_SL g160 ( 
.A(n_26),
.B(n_161),
.Y(n_160)
);

CKINVDCx16_ASAP7_75t_R g26 ( 
.A(n_27),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_27),
.A2(n_45),
.B1(n_132),
.B2(n_133),
.Y(n_131)
);

BUFx8_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

BUFx24_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

CKINVDCx16_ASAP7_75t_R g33 ( 
.A(n_30),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_30),
.B(n_144),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_L g156 ( 
.A1(n_33),
.A2(n_149),
.B(n_157),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_33),
.B(n_68),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_SL g180 ( 
.A1(n_33),
.A2(n_157),
.B(n_181),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_L g36 ( 
.A1(n_37),
.A2(n_41),
.B1(n_47),
.B2(n_49),
.Y(n_36)
);

OAI21xp5_ASAP7_75t_L g52 ( 
.A1(n_37),
.A2(n_49),
.B(n_53),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_38),
.A2(n_39),
.B1(n_78),
.B2(n_79),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_SL g179 ( 
.A(n_38),
.B(n_78),
.Y(n_179)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

O2A1O1Ixp33_ASAP7_75t_L g42 ( 
.A1(n_39),
.A2(n_43),
.B(n_45),
.C(n_46),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_39),
.B(n_43),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g177 ( 
.A1(n_39),
.A2(n_80),
.B1(n_178),
.B2(n_179),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_L g170 ( 
.A1(n_41),
.A2(n_49),
.B1(n_140),
.B2(n_171),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_SL g192 ( 
.A1(n_41),
.A2(n_171),
.B(n_193),
.Y(n_192)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_42),
.B(n_54),
.Y(n_53)
);

CKINVDCx16_ASAP7_75t_R g43 ( 
.A(n_44),
.Y(n_43)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_46),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_49),
.B(n_55),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_L g139 ( 
.A1(n_49),
.A2(n_53),
.B(n_140),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_SL g155 ( 
.A(n_49),
.B(n_68),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g50 ( 
.A(n_51),
.B(n_57),
.C(n_74),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_51),
.A2(n_52),
.B1(n_74),
.B2(n_75),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_52),
.Y(n_51)
);

INVxp67_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

XOR2xp5_ASAP7_75t_L g106 ( 
.A(n_57),
.B(n_107),
.Y(n_106)
);

AOI21xp5_ASAP7_75t_L g57 ( 
.A1(n_58),
.A2(n_67),
.B(n_70),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_58),
.B(n_73),
.Y(n_91)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

A2O1A1Ixp33_ASAP7_75t_L g59 ( 
.A1(n_60),
.A2(n_62),
.B(n_63),
.C(n_64),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_60),
.B(n_62),
.Y(n_63)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_60),
.Y(n_69)
);

A2O1A1Ixp33_ASAP7_75t_L g100 ( 
.A1(n_60),
.A2(n_62),
.B(n_68),
.C(n_101),
.Y(n_100)
);

BUFx2_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_64),
.Y(n_72)
);

OAI21xp33_ASAP7_75t_L g89 ( 
.A1(n_64),
.A2(n_90),
.B(n_91),
.Y(n_89)
);

INVx8_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

O2A1O1Ixp33_ASAP7_75t_SL g77 ( 
.A1(n_66),
.A2(n_78),
.B(n_80),
.C(n_81),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_66),
.B(n_78),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_71),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_72),
.B(n_73),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_75),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_76),
.A2(n_82),
.B1(n_84),
.B2(n_85),
.Y(n_75)
);

OAI21xp5_ASAP7_75t_L g93 ( 
.A1(n_76),
.A2(n_85),
.B(n_94),
.Y(n_93)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_77),
.B(n_115),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_79),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_81),
.Y(n_84)
);

OAI21xp5_ASAP7_75t_L g113 ( 
.A1(n_82),
.A2(n_84),
.B(n_114),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_84),
.B(n_96),
.Y(n_95)
);

XOR2xp5_ASAP7_75t_L g87 ( 
.A(n_88),
.B(n_98),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_89),
.A2(n_92),
.B1(n_93),
.B2(n_97),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_89),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_93),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_95),
.Y(n_94)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_96),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_102),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_99),
.A2(n_100),
.B1(n_102),
.B2(n_109),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_100),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_102),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_104),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_106),
.B(n_108),
.C(n_110),
.Y(n_105)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_106),
.B(n_200),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_L g200 ( 
.A1(n_108),
.A2(n_110),
.B1(n_111),
.B2(n_201),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_108),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_111),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_112),
.B(n_116),
.C(n_117),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_112),
.A2(n_113),
.B1(n_188),
.B2(n_189),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_113),
.Y(n_112)
);

XOR2xp5_ASAP7_75t_L g188 ( 
.A(n_116),
.B(n_117),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_118),
.Y(n_181)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

AOI21xp5_ASAP7_75t_L g121 ( 
.A1(n_122),
.A2(n_197),
.B(n_202),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_SL g122 ( 
.A1(n_123),
.A2(n_184),
.B(n_196),
.Y(n_122)
);

AOI21xp5_ASAP7_75t_L g123 ( 
.A1(n_124),
.A2(n_165),
.B(n_183),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_SL g124 ( 
.A1(n_125),
.A2(n_145),
.B(n_164),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_134),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_126),
.B(n_134),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_SL g126 ( 
.A(n_127),
.B(n_130),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_127),
.A2(n_130),
.B1(n_131),
.B2(n_152),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_127),
.Y(n_152)
);

INVxp67_ASAP7_75t_L g133 ( 
.A(n_128),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_129),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_131),
.Y(n_130)
);

XNOR2xp5_ASAP7_75t_L g134 ( 
.A(n_135),
.B(n_141),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_136),
.A2(n_137),
.B1(n_138),
.B2(n_139),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_136),
.B(n_139),
.C(n_141),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_137),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_139),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_142),
.Y(n_150)
);

AOI21xp5_ASAP7_75t_L g145 ( 
.A1(n_146),
.A2(n_153),
.B(n_163),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_151),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_SL g163 ( 
.A(n_147),
.B(n_151),
.Y(n_163)
);

CKINVDCx16_ASAP7_75t_R g148 ( 
.A(n_149),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_SL g153 ( 
.A1(n_154),
.A2(n_158),
.B(n_162),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_156),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_155),
.B(n_156),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_159),
.B(n_160),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_167),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_SL g183 ( 
.A(n_166),
.B(n_167),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_168),
.A2(n_169),
.B1(n_176),
.B2(n_182),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_170),
.A2(n_172),
.B1(n_174),
.B2(n_175),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_170),
.Y(n_175)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_172),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_172),
.B(n_175),
.C(n_182),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_173),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_176),
.Y(n_182)
);

XOR2xp5_ASAP7_75t_L g176 ( 
.A(n_177),
.B(n_180),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_177),
.B(n_180),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_186),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_185),
.B(n_186),
.Y(n_196)
);

XOR2xp5_ASAP7_75t_L g186 ( 
.A(n_187),
.B(n_190),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_187),
.B(n_192),
.C(n_194),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_188),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_191),
.A2(n_192),
.B1(n_194),
.B2(n_195),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_191),
.Y(n_194)
);

CKINVDCx16_ASAP7_75t_R g195 ( 
.A(n_192),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_199),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_SL g202 ( 
.A(n_198),
.B(n_199),
.Y(n_202)
);


endmodule