module real_jpeg_33930_n_9 (n_79, n_77, n_5, n_4, n_8, n_0, n_1, n_73, n_74, n_2, n_75, n_78, n_6, n_72, n_7, n_3, n_76, n_9);

input n_79;
input n_77;
input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_73;
input n_74;
input n_2;
input n_75;
input n_78;
input n_6;
input n_72;
input n_7;
input n_3;
input n_76;

output n_9;

wire n_54;
wire n_37;
wire n_38;
wire n_35;
wire n_29;
wire n_49;
wire n_10;
wire n_68;
wire n_64;
wire n_11;
wire n_47;
wire n_22;
wire n_40;
wire n_27;
wire n_56;
wire n_48;
wire n_13;
wire n_65;
wire n_33;
wire n_67;
wire n_66;
wire n_28;
wire n_44;
wire n_62;
wire n_45;
wire n_42;
wire n_18;
wire n_39;
wire n_26;
wire n_19;
wire n_17;
wire n_21;
wire n_50;
wire n_69;
wire n_31;
wire n_23;
wire n_51;
wire n_14;
wire n_61;
wire n_70;
wire n_41;
wire n_32;
wire n_20;
wire n_30;
wire n_15;
wire n_43;
wire n_57;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_12;
wire n_24;
wire n_34;
wire n_60;
wire n_46;
wire n_59;
wire n_25;
wire n_53;
wire n_36;
wire n_16;

INVx1_ASAP7_75t_L g54 ( 
.A(n_0),
.Y(n_54)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_1),
.Y(n_56)
);

AOI221xp5_ASAP7_75t_L g38 ( 
.A1(n_2),
.A2(n_5),
.B1(n_39),
.B2(n_43),
.C(n_46),
.Y(n_38)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_2),
.Y(n_48)
);

OAI22xp33_ASAP7_75t_SL g10 ( 
.A1(n_3),
.A2(n_11),
.B1(n_12),
.B2(n_19),
.Y(n_10)
);

INVx1_ASAP7_75t_L g11 ( 
.A(n_3),
.Y(n_11)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_4),
.Y(n_37)
);

MAJIxp5_ASAP7_75t_L g49 ( 
.A(n_5),
.B(n_39),
.C(n_43),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_SL g64 ( 
.A(n_6),
.B(n_65),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_6),
.B(n_65),
.Y(n_70)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_7),
.B(n_24),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_8),
.B(n_41),
.Y(n_40)
);

XNOR2xp5_ASAP7_75t_L g9 ( 
.A(n_10),
.B(n_20),
.Y(n_9)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_14),
.Y(n_12)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_14),
.B(n_53),
.Y(n_52)
);

INVx2_ASAP7_75t_L g14 ( 
.A(n_15),
.Y(n_14)
);

INVx3_ASAP7_75t_L g15 ( 
.A(n_16),
.Y(n_15)
);

INVx5_ASAP7_75t_L g16 ( 
.A(n_17),
.Y(n_16)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_17),
.Y(n_69)
);

INVx8_ASAP7_75t_L g17 ( 
.A(n_18),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_18),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_18),
.Y(n_45)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_18),
.Y(n_61)
);

OAI21xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_64),
.B(n_70),
.Y(n_20)
);

AOI21xp5_ASAP7_75t_SL g21 ( 
.A1(n_22),
.A2(n_29),
.B(n_62),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_SL g22 ( 
.A(n_23),
.B(n_28),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_26),
.Y(n_24)
);

HB1xp67_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_27),
.B(n_42),
.Y(n_41)
);

MAJIxp5_ASAP7_75t_L g29 ( 
.A(n_30),
.B(n_56),
.C(n_57),
.Y(n_29)
);

AOI21xp5_ASAP7_75t_SL g30 ( 
.A1(n_31),
.A2(n_50),
.B(n_55),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_L g31 ( 
.A1(n_32),
.A2(n_38),
.B1(n_48),
.B2(n_49),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_34),
.B(n_35),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_SL g46 ( 
.A(n_40),
.B(n_47),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_43),
.Y(n_47)
);

AND2x2_ASAP7_75t_L g43 ( 
.A(n_44),
.B(n_76),
.Y(n_43)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g50 ( 
.A(n_51),
.B(n_54),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_51),
.B(n_54),
.Y(n_55)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_59),
.B(n_60),
.Y(n_58)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVxp67_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

NOR2x1_ASAP7_75t_L g65 ( 
.A(n_66),
.B(n_67),
.Y(n_65)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_72),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_73),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_74),
.Y(n_34)
);

INVxp67_ASAP7_75t_L g42 ( 
.A(n_75),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_77),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_78),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_79),
.Y(n_66)
);


endmodule