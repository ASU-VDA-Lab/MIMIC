module fake_jpeg_28634_n_147 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_39, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_147);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_39;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_147;

wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_138;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g41 ( 
.A(n_9),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_23),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_29),
.Y(n_43)
);

CKINVDCx14_ASAP7_75t_R g44 ( 
.A(n_19),
.Y(n_44)
);

BUFx12_ASAP7_75t_L g45 ( 
.A(n_8),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_1),
.Y(n_46)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_27),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_40),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_24),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_5),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_28),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_6),
.Y(n_52)
);

BUFx16f_ASAP7_75t_L g53 ( 
.A(n_7),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_37),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_14),
.Y(n_55)
);

BUFx10_ASAP7_75t_L g56 ( 
.A(n_5),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_38),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_3),
.B(n_33),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_47),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_59),
.Y(n_71)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_47),
.Y(n_60)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_60),
.Y(n_74)
);

BUFx16f_ASAP7_75t_L g61 ( 
.A(n_53),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_61),
.B(n_65),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_56),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_62),
.B(n_63),
.Y(n_82)
);

INVx4_ASAP7_75t_SL g63 ( 
.A(n_53),
.Y(n_63)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_56),
.Y(n_64)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_64),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_56),
.Y(n_65)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_42),
.Y(n_66)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_66),
.Y(n_81)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_41),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_67),
.B(n_48),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_66),
.B(n_50),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_69),
.B(n_75),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_SL g70 ( 
.A(n_61),
.B(n_58),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_70),
.B(n_73),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_60),
.B(n_46),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_59),
.B(n_44),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_76),
.B(n_80),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_63),
.B(n_58),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_77),
.B(n_78),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_SL g78 ( 
.A(n_64),
.B(n_51),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_L g79 ( 
.A1(n_60),
.A2(n_44),
.B1(n_55),
.B2(n_54),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_79),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_67),
.B(n_52),
.Y(n_80)
);

INVx13_ASAP7_75t_L g83 ( 
.A(n_81),
.Y(n_83)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_83),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_L g84 ( 
.A1(n_82),
.A2(n_57),
.B(n_49),
.Y(n_84)
);

OR2x2_ASAP7_75t_L g118 ( 
.A(n_84),
.B(n_21),
.Y(n_118)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_81),
.Y(n_85)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_85),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_72),
.B(n_43),
.C(n_45),
.Y(n_86)
);

OAI21xp5_ASAP7_75t_SL g105 ( 
.A1(n_86),
.A2(n_92),
.B(n_4),
.Y(n_105)
);

INVx1_ASAP7_75t_SL g87 ( 
.A(n_68),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_87),
.B(n_94),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_79),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_89),
.B(n_3),
.Y(n_103)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_68),
.Y(n_91)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_91),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_74),
.B(n_45),
.C(n_22),
.Y(n_92)
);

INVx1_ASAP7_75t_SL g94 ( 
.A(n_71),
.Y(n_94)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_71),
.Y(n_96)
);

INVx1_ASAP7_75t_SL g117 ( 
.A(n_96),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_97),
.A2(n_16),
.B1(n_17),
.B2(n_18),
.Y(n_112)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_82),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_98),
.B(n_4),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_77),
.B(n_0),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_99),
.B(n_2),
.Y(n_102)
);

BUFx3_ASAP7_75t_L g100 ( 
.A(n_68),
.Y(n_100)
);

BUFx5_ASAP7_75t_L g101 ( 
.A(n_100),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_102),
.B(n_105),
.Y(n_131)
);

CKINVDCx14_ASAP7_75t_R g124 ( 
.A(n_103),
.Y(n_124)
);

BUFx3_ASAP7_75t_L g104 ( 
.A(n_83),
.Y(n_104)
);

INVx1_ASAP7_75t_SL g121 ( 
.A(n_104),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_107),
.B(n_109),
.Y(n_132)
);

AOI21xp5_ASAP7_75t_L g108 ( 
.A1(n_98),
.A2(n_10),
.B(n_11),
.Y(n_108)
);

INVxp67_ASAP7_75t_L g128 ( 
.A(n_108),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_93),
.B(n_12),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_SL g110 ( 
.A(n_93),
.B(n_13),
.C(n_15),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_110),
.A2(n_26),
.B1(n_30),
.B2(n_31),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_90),
.B(n_95),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_111),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_112),
.A2(n_116),
.B1(n_120),
.B2(n_32),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_90),
.B(n_20),
.Y(n_114)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_114),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_88),
.B(n_39),
.Y(n_116)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_118),
.Y(n_130)
);

HAxp5_ASAP7_75t_SL g120 ( 
.A(n_98),
.B(n_25),
.CON(n_120),
.SN(n_120)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_123),
.B(n_126),
.Y(n_133)
);

BUFx2_ASAP7_75t_L g126 ( 
.A(n_101),
.Y(n_126)
);

INVxp33_ASAP7_75t_L g127 ( 
.A(n_106),
.Y(n_127)
);

INVxp67_ASAP7_75t_L g135 ( 
.A(n_127),
.Y(n_135)
);

NAND3xp33_ASAP7_75t_L g137 ( 
.A(n_129),
.B(n_34),
.C(n_35),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_125),
.A2(n_117),
.B1(n_113),
.B2(n_118),
.Y(n_134)
);

FAx1_ASAP7_75t_SL g139 ( 
.A(n_134),
.B(n_136),
.CI(n_137),
.CON(n_139),
.SN(n_139)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_124),
.A2(n_119),
.B1(n_115),
.B2(n_120),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_135),
.B(n_128),
.C(n_131),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_138),
.B(n_140),
.Y(n_141)
);

AOI21xp5_ASAP7_75t_SL g140 ( 
.A1(n_133),
.A2(n_130),
.B(n_124),
.Y(n_140)
);

HB1xp67_ASAP7_75t_L g142 ( 
.A(n_141),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_SL g143 ( 
.A1(n_142),
.A2(n_126),
.B1(n_122),
.B2(n_121),
.Y(n_143)
);

OR2x2_ASAP7_75t_L g144 ( 
.A(n_143),
.B(n_104),
.Y(n_144)
);

CKINVDCx5p33_ASAP7_75t_R g145 ( 
.A(n_144),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_L g146 ( 
.A(n_145),
.B(n_139),
.Y(n_146)
);

FAx1_ASAP7_75t_SL g147 ( 
.A(n_146),
.B(n_132),
.CI(n_36),
.CON(n_147),
.SN(n_147)
);


endmodule