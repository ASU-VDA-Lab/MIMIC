module real_jpeg_23449_n_14 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_2, n_13, n_6, n_7, n_3, n_10, n_9, n_14);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_2;
input n_13;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_14;

wire n_108;
wire n_54;
wire n_37;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_78;
wire n_83;
wire n_104;
wire n_64;
wire n_47;
wire n_22;
wire n_87;
wire n_105;
wire n_40;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_113;
wire n_120;
wire n_93;
wire n_95;
wire n_65;
wire n_33;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_66;
wire n_28;
wire n_44;
wire n_62;
wire n_121;
wire n_106;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_77;
wire n_109;
wire n_39;
wire n_94;
wire n_26;
wire n_19;
wire n_118;
wire n_17;
wire n_116;
wire n_21;
wire n_50;
wire n_69;
wire n_31;
wire n_72;
wire n_100;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_117;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_30;
wire n_15;
wire n_103;
wire n_43;
wire n_57;
wire n_84;
wire n_82;
wire n_111;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_25;
wire n_53;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_101;
wire n_96;
wire n_89;
wire n_16;

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_0),
.B(n_105),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_1),
.B(n_60),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_1),
.B(n_26),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_1),
.B(n_35),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_2),
.Y(n_86)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_3),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_4),
.B(n_95),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_4),
.B(n_26),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

INVx8_ASAP7_75t_SL g118 ( 
.A(n_6),
.Y(n_118)
);

BUFx12f_ASAP7_75t_L g70 ( 
.A(n_7),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_8),
.B(n_26),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_8),
.B(n_13),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_8),
.B(n_35),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_8),
.B(n_32),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_8),
.B(n_70),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_9),
.B(n_22),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_9),
.B(n_26),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_9),
.B(n_35),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_9),
.B(n_32),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_10),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_11),
.B(n_32),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_11),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_11),
.B(n_26),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_11),
.B(n_70),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_11),
.B(n_84),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_11),
.B(n_117),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_12),
.B(n_35),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_12),
.B(n_26),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_12),
.B(n_50),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_12),
.B(n_32),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_12),
.B(n_70),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_12),
.B(n_84),
.Y(n_119)
);

INVx6_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_13),
.Y(n_51)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_13),
.Y(n_61)
);

INVx6_ASAP7_75t_L g96 ( 
.A(n_13),
.Y(n_96)
);

XNOR2xp5_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_98),
.Y(n_14)
);

MAJIxp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_75),
.C(n_76),
.Y(n_15)
);

MAJIxp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_52),
.C(n_53),
.Y(n_16)
);

MAJIxp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_37),
.C(n_42),
.Y(n_17)
);

AOI22xp5_ASAP7_75t_SL g18 ( 
.A1(n_19),
.A2(n_20),
.B1(n_29),
.B2(n_30),
.Y(n_18)
);

MAJIxp5_ASAP7_75t_L g52 ( 
.A(n_19),
.B(n_31),
.C(n_34),
.Y(n_52)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

OAI22xp5_ASAP7_75t_SL g20 ( 
.A1(n_21),
.A2(n_24),
.B1(n_25),
.B2(n_28),
.Y(n_20)
);

CKINVDCx14_ASAP7_75t_R g28 ( 
.A(n_21),
.Y(n_28)
);

INVx5_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

INVx8_ASAP7_75t_L g105 ( 
.A(n_23),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_24),
.B(n_28),
.Y(n_56)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

XNOR2xp5_ASAP7_75t_SL g30 ( 
.A(n_31),
.B(n_34),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx13_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

BUFx24_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_SL g37 ( 
.A(n_38),
.B(n_40),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_SL g43 ( 
.A1(n_38),
.A2(n_39),
.B1(n_40),
.B2(n_41),
.Y(n_43)
);

CKINVDCx16_ASAP7_75t_R g38 ( 
.A(n_39),
.Y(n_38)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

MAJIxp5_ASAP7_75t_L g42 ( 
.A(n_43),
.B(n_44),
.C(n_47),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_45),
.B(n_46),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_48),
.B(n_49),
.Y(n_47)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

XNOR2xp5_ASAP7_75t_L g53 ( 
.A(n_54),
.B(n_65),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g54 ( 
.A1(n_55),
.A2(n_56),
.B1(n_57),
.B2(n_58),
.Y(n_54)
);

MAJIxp5_ASAP7_75t_L g75 ( 
.A(n_55),
.B(n_58),
.C(n_65),
.Y(n_75)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_59),
.A2(n_62),
.B1(n_63),
.B2(n_64),
.Y(n_58)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_59),
.Y(n_64)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_62),
.B(n_64),
.Y(n_88)
);

CKINVDCx14_ASAP7_75t_R g62 ( 
.A(n_63),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g65 ( 
.A1(n_66),
.A2(n_67),
.B1(n_68),
.B2(n_74),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_66),
.Y(n_74)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g68 ( 
.A1(n_69),
.A2(n_71),
.B1(n_72),
.B2(n_73),
.Y(n_68)
);

CKINVDCx16_ASAP7_75t_R g73 ( 
.A(n_69),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g78 ( 
.A(n_71),
.B(n_73),
.C(n_74),
.Y(n_78)
);

CKINVDCx14_ASAP7_75t_R g71 ( 
.A(n_72),
.Y(n_71)
);

XNOR2xp5_ASAP7_75t_SL g76 ( 
.A(n_77),
.B(n_87),
.Y(n_76)
);

XNOR2xp5_ASAP7_75t_L g77 ( 
.A(n_78),
.B(n_79),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_78),
.B(n_79),
.C(n_87),
.Y(n_99)
);

XNOR2xp5_ASAP7_75t_L g79 ( 
.A(n_80),
.B(n_81),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_80),
.B(n_82),
.C(n_83),
.Y(n_109)
);

XNOR2xp5_ASAP7_75t_L g81 ( 
.A(n_82),
.B(n_83),
.Y(n_81)
);

BUFx12f_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

BUFx12f_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

XNOR2xp5_ASAP7_75t_SL g87 ( 
.A(n_88),
.B(n_89),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_88),
.B(n_90),
.C(n_91),
.Y(n_121)
);

XNOR2xp5_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_91),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_92),
.A2(n_93),
.B1(n_94),
.B2(n_97),
.Y(n_91)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_92),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_93),
.B(n_97),
.Y(n_120)
);

CKINVDCx14_ASAP7_75t_R g93 ( 
.A(n_94),
.Y(n_93)
);

INVx5_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

XOR2xp5_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_100),
.Y(n_98)
);

XOR2xp5_ASAP7_75t_L g100 ( 
.A(n_101),
.B(n_114),
.Y(n_100)
);

XNOR2xp5_ASAP7_75t_SL g101 ( 
.A(n_102),
.B(n_110),
.Y(n_101)
);

XNOR2xp5_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_109),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_104),
.A2(n_106),
.B1(n_107),
.B2(n_108),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_104),
.Y(n_108)
);

CKINVDCx16_ASAP7_75t_R g106 ( 
.A(n_107),
.Y(n_106)
);

BUFx24_ASAP7_75t_SL g124 ( 
.A(n_110),
.Y(n_124)
);

FAx1_ASAP7_75t_SL g110 ( 
.A(n_111),
.B(n_112),
.CI(n_113),
.CON(n_110),
.SN(n_110)
);

XOR2xp5_ASAP7_75t_L g114 ( 
.A(n_115),
.B(n_121),
.Y(n_114)
);

BUFx24_ASAP7_75t_SL g122 ( 
.A(n_115),
.Y(n_122)
);

FAx1_ASAP7_75t_SL g115 ( 
.A(n_116),
.B(n_119),
.CI(n_120),
.CON(n_115),
.SN(n_115)
);

INVx8_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);


endmodule