module fake_jpeg_12002_n_145 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_145);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_145;

wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_38;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_37;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_138;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx4f_ASAP7_75t_SL g37 ( 
.A(n_14),
.Y(n_37)
);

BUFx5_ASAP7_75t_L g38 ( 
.A(n_0),
.Y(n_38)
);

BUFx5_ASAP7_75t_L g39 ( 
.A(n_12),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_36),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_2),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_33),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_28),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_22),
.Y(n_44)
);

BUFx16f_ASAP7_75t_L g45 ( 
.A(n_26),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_18),
.Y(n_46)
);

BUFx5_ASAP7_75t_L g47 ( 
.A(n_19),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_2),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_35),
.Y(n_49)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_3),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_1),
.Y(n_51)
);

BUFx12_ASAP7_75t_L g52 ( 
.A(n_34),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_23),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_13),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_20),
.Y(n_55)
);

BUFx5_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_56),
.Y(n_75)
);

INVx13_ASAP7_75t_L g57 ( 
.A(n_37),
.Y(n_57)
);

HB1xp67_ASAP7_75t_L g70 ( 
.A(n_57),
.Y(n_70)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_50),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_58),
.Y(n_77)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_38),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_59),
.B(n_60),
.Y(n_73)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_41),
.Y(n_60)
);

INVx3_ASAP7_75t_SL g61 ( 
.A(n_51),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_61),
.B(n_64),
.Y(n_72)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_38),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_62),
.B(n_63),
.Y(n_79)
);

BUFx5_ASAP7_75t_L g63 ( 
.A(n_39),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_44),
.B(n_0),
.Y(n_64)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_50),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_65),
.B(n_48),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_59),
.A2(n_48),
.B1(n_51),
.B2(n_42),
.Y(n_66)
);

CKINVDCx16_ASAP7_75t_R g81 ( 
.A(n_66),
.Y(n_81)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_61),
.Y(n_67)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_67),
.Y(n_85)
);

NAND2xp33_ASAP7_75t_SL g87 ( 
.A(n_68),
.B(n_52),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_62),
.A2(n_42),
.B1(n_54),
.B2(n_40),
.Y(n_69)
);

OAI32xp33_ASAP7_75t_L g86 ( 
.A1(n_69),
.A2(n_45),
.A3(n_52),
.B1(n_47),
.B2(n_6),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_57),
.A2(n_43),
.B1(n_55),
.B2(n_53),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_L g94 ( 
.A1(n_71),
.A2(n_74),
.B1(n_52),
.B2(n_4),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_56),
.A2(n_49),
.B1(n_46),
.B2(n_37),
.Y(n_74)
);

INVx6_ASAP7_75t_L g76 ( 
.A(n_61),
.Y(n_76)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_76),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_59),
.A2(n_37),
.B1(n_47),
.B2(n_45),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_78),
.B(n_4),
.Y(n_96)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_71),
.Y(n_82)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_82),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_72),
.B(n_1),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_83),
.B(n_84),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_70),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_86),
.B(n_91),
.Y(n_113)
);

AOI21xp5_ASAP7_75t_L g98 ( 
.A1(n_87),
.A2(n_96),
.B(n_75),
.Y(n_98)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_73),
.Y(n_88)
);

HB1xp67_ASAP7_75t_L g110 ( 
.A(n_88),
.Y(n_110)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_77),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_89),
.B(n_90),
.Y(n_101)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_77),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_74),
.Y(n_91)
);

HB1xp67_ASAP7_75t_L g92 ( 
.A(n_67),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_92),
.B(n_93),
.Y(n_102)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_69),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_94),
.B(n_95),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_68),
.B(n_3),
.Y(n_95)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_76),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_97),
.B(n_75),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_L g121 ( 
.A1(n_98),
.A2(n_111),
.B(n_114),
.Y(n_121)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_85),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_104),
.B(n_107),
.Y(n_125)
);

AO22x1_ASAP7_75t_SL g105 ( 
.A1(n_87),
.A2(n_86),
.B1(n_81),
.B2(n_94),
.Y(n_105)
);

A2O1A1Ixp33_ASAP7_75t_SL g119 ( 
.A1(n_105),
.A2(n_114),
.B(n_10),
.C(n_11),
.Y(n_119)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_106),
.Y(n_120)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_85),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_80),
.B(n_79),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_108),
.B(n_109),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_80),
.B(n_5),
.Y(n_109)
);

OAI21xp5_ASAP7_75t_L g111 ( 
.A1(n_87),
.A2(n_5),
.B(n_6),
.Y(n_111)
);

AND2x2_ASAP7_75t_L g112 ( 
.A(n_95),
.B(n_7),
.Y(n_112)
);

XNOR2xp5_ASAP7_75t_L g118 ( 
.A(n_112),
.B(n_116),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_81),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_L g115 ( 
.A1(n_93),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_115),
.A2(n_103),
.B1(n_99),
.B2(n_100),
.Y(n_128)
);

XOR2xp5_ASAP7_75t_L g116 ( 
.A(n_87),
.B(n_30),
.Y(n_116)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_101),
.Y(n_117)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_117),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_119),
.A2(n_123),
.B1(n_124),
.B2(n_126),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_121),
.B(n_122),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_110),
.B(n_11),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_113),
.A2(n_15),
.B1(n_16),
.B2(n_17),
.Y(n_123)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_104),
.Y(n_124)
);

CKINVDCx16_ASAP7_75t_R g126 ( 
.A(n_102),
.Y(n_126)
);

NOR4xp25_ASAP7_75t_L g131 ( 
.A(n_128),
.B(n_105),
.C(n_115),
.D(n_112),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_131),
.A2(n_133),
.B1(n_119),
.B2(n_118),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_120),
.A2(n_105),
.B1(n_107),
.B2(n_25),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_129),
.B(n_127),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_134),
.B(n_135),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_133),
.A2(n_120),
.B1(n_119),
.B2(n_125),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_136),
.B(n_130),
.Y(n_138)
);

AOI21xp5_ASAP7_75t_SL g139 ( 
.A1(n_138),
.A2(n_132),
.B(n_119),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_139),
.A2(n_135),
.B1(n_137),
.B2(n_27),
.Y(n_140)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_140),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_141),
.B(n_21),
.C(n_24),
.Y(n_142)
);

INVxp67_ASAP7_75t_L g143 ( 
.A(n_142),
.Y(n_143)
);

OA21x2_ASAP7_75t_SL g144 ( 
.A1(n_143),
.A2(n_29),
.B(n_31),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_SL g145 ( 
.A(n_144),
.B(n_32),
.Y(n_145)
);


endmodule