module fake_jpeg_31642_n_320 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_320);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_320;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_12),
.B(n_3),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_0),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_9),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_15),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_12),
.Y(n_23)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_12),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_15),
.Y(n_26)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

HB1xp67_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

BUFx8_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

INVx11_ASAP7_75t_SL g33 ( 
.A(n_0),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_28),
.Y(n_34)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_34),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_22),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_35),
.Y(n_57)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_28),
.Y(n_36)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_36),
.Y(n_55)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_33),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_37),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_22),
.Y(n_38)
);

BUFx2_ASAP7_75t_L g47 ( 
.A(n_38),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_22),
.Y(n_39)
);

BUFx2_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

INVx2_ASAP7_75t_SL g40 ( 
.A(n_33),
.Y(n_40)
);

CKINVDCx16_ASAP7_75t_R g46 ( 
.A(n_40),
.Y(n_46)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_22),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_41),
.B(n_42),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_29),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_18),
.B(n_0),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_43),
.B(n_18),
.Y(n_45)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_29),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_44),
.B(n_32),
.Y(n_52)
);

AND2x2_ASAP7_75t_L g82 ( 
.A(n_45),
.B(n_52),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_34),
.A2(n_24),
.B1(n_27),
.B2(n_21),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_48),
.A2(n_40),
.B1(n_19),
.B2(n_39),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_L g49 ( 
.A(n_36),
.B(n_43),
.C(n_44),
.Y(n_49)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_49),
.B(n_29),
.C(n_31),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_40),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_51),
.B(n_37),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_40),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_53),
.B(n_54),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_SL g54 ( 
.A(n_37),
.B(n_20),
.Y(n_54)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_55),
.Y(n_60)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_60),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_55),
.A2(n_24),
.B1(n_27),
.B2(n_17),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_61),
.A2(n_66),
.B1(n_59),
.B2(n_32),
.Y(n_111)
);

AOI21xp33_ASAP7_75t_L g62 ( 
.A1(n_45),
.A2(n_17),
.B(n_30),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_62),
.B(n_65),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_49),
.A2(n_41),
.B1(n_42),
.B2(n_38),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_63),
.A2(n_83),
.B1(n_86),
.B2(n_59),
.Y(n_113)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_55),
.Y(n_64)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_64),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_54),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_48),
.A2(n_24),
.B1(n_27),
.B2(n_30),
.Y(n_66)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_58),
.Y(n_68)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_68),
.Y(n_123)
);

HB1xp67_ASAP7_75t_L g69 ( 
.A(n_58),
.Y(n_69)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_69),
.Y(n_120)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_58),
.Y(n_70)
);

CKINVDCx16_ASAP7_75t_R g101 ( 
.A(n_70),
.Y(n_101)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_50),
.Y(n_71)
);

INVx1_ASAP7_75t_SL g115 ( 
.A(n_71),
.Y(n_115)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_50),
.Y(n_72)
);

AND2x2_ASAP7_75t_L g109 ( 
.A(n_72),
.B(n_74),
.Y(n_109)
);

INVxp67_ASAP7_75t_L g73 ( 
.A(n_52),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_73),
.B(n_84),
.Y(n_112)
);

O2A1O1Ixp33_ASAP7_75t_L g75 ( 
.A1(n_51),
.A2(n_19),
.B(n_26),
.C(n_20),
.Y(n_75)
);

O2A1O1Ixp33_ASAP7_75t_L g100 ( 
.A1(n_75),
.A2(n_26),
.B(n_59),
.C(n_37),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_76),
.B(n_80),
.Y(n_105)
);

XNOR2xp5_ASAP7_75t_L g103 ( 
.A(n_77),
.B(n_90),
.Y(n_103)
);

BUFx3_ASAP7_75t_L g78 ( 
.A(n_57),
.Y(n_78)
);

INVx5_ASAP7_75t_L g106 ( 
.A(n_78),
.Y(n_106)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_47),
.Y(n_79)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_79),
.Y(n_122)
);

AO22x1_ASAP7_75t_SL g80 ( 
.A1(n_49),
.A2(n_39),
.B1(n_42),
.B2(n_38),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_45),
.A2(n_35),
.B1(n_39),
.B2(n_25),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_L g107 ( 
.A1(n_81),
.A2(n_85),
.B1(n_26),
.B2(n_56),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_47),
.A2(n_35),
.B1(n_29),
.B2(n_31),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_53),
.B(n_23),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_57),
.A2(n_25),
.B1(n_23),
.B2(n_20),
.Y(n_85)
);

OA22x2_ASAP7_75t_L g86 ( 
.A1(n_46),
.A2(n_32),
.B1(n_16),
.B2(n_17),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_57),
.A2(n_21),
.B1(n_31),
.B2(n_16),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_87),
.A2(n_95),
.B1(n_32),
.B2(n_37),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_57),
.Y(n_88)
);

INVx11_ASAP7_75t_L g119 ( 
.A(n_88),
.Y(n_119)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_47),
.Y(n_89)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_89),
.Y(n_108)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_46),
.B(n_32),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_51),
.B(n_19),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_91),
.B(n_92),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_47),
.B(n_23),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_56),
.B(n_25),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_93),
.B(n_59),
.Y(n_118)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_56),
.Y(n_94)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_94),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_56),
.A2(n_21),
.B1(n_30),
.B2(n_16),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_91),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_97),
.B(n_98),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_75),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_100),
.B(n_118),
.Y(n_146)
);

AOI21xp5_ASAP7_75t_L g102 ( 
.A1(n_73),
.A2(n_0),
.B(n_1),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g133 ( 
.A(n_102),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_107),
.A2(n_111),
.B1(n_124),
.B2(n_126),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_110),
.A2(n_113),
.B1(n_116),
.B2(n_121),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_77),
.A2(n_59),
.B1(n_32),
.B2(n_8),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_82),
.A2(n_59),
.B1(n_15),
.B2(n_14),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_71),
.A2(n_14),
.B1(n_13),
.B2(n_11),
.Y(n_124)
);

AND2x4_ASAP7_75t_SL g125 ( 
.A(n_82),
.B(n_1),
.Y(n_125)
);

AND2x2_ASAP7_75t_L g136 ( 
.A(n_125),
.B(n_90),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_72),
.A2(n_14),
.B1(n_13),
.B2(n_11),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_100),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_127),
.B(n_147),
.Y(n_165)
);

INVx13_ASAP7_75t_L g129 ( 
.A(n_104),
.Y(n_129)
);

INVxp67_ASAP7_75t_L g184 ( 
.A(n_129),
.Y(n_184)
);

BUFx3_ASAP7_75t_L g130 ( 
.A(n_106),
.Y(n_130)
);

BUFx5_ASAP7_75t_L g164 ( 
.A(n_130),
.Y(n_164)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_99),
.Y(n_131)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_131),
.Y(n_159)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_99),
.Y(n_132)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_132),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_97),
.B(n_67),
.Y(n_134)
);

CKINVDCx14_ASAP7_75t_R g156 ( 
.A(n_134),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_115),
.B(n_112),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_135),
.B(n_138),
.Y(n_182)
);

AND2x2_ASAP7_75t_L g172 ( 
.A(n_136),
.B(n_144),
.Y(n_172)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_122),
.Y(n_137)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_137),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_114),
.B(n_82),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_SL g139 ( 
.A(n_96),
.B(n_63),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_139),
.B(n_145),
.C(n_103),
.Y(n_161)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_117),
.Y(n_140)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_140),
.Y(n_171)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_117),
.Y(n_142)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_142),
.Y(n_177)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_123),
.Y(n_143)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_143),
.Y(n_180)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_123),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_103),
.B(n_65),
.C(n_64),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_SL g147 ( 
.A(n_112),
.B(n_92),
.Y(n_147)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_122),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_148),
.B(n_150),
.Y(n_155)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_120),
.Y(n_149)
);

AND2x2_ASAP7_75t_L g174 ( 
.A(n_149),
.B(n_108),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_114),
.B(n_80),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_SL g152 ( 
.A(n_96),
.B(n_93),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_152),
.B(n_153),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_115),
.B(n_76),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_141),
.A2(n_105),
.B1(n_98),
.B2(n_109),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_154),
.A2(n_166),
.B1(n_173),
.B2(n_179),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_L g157 ( 
.A1(n_133),
.A2(n_102),
.B(n_109),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_L g187 ( 
.A1(n_157),
.A2(n_178),
.B(n_183),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_128),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_158),
.B(n_160),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_128),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_161),
.B(n_125),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_141),
.A2(n_109),
.B1(n_105),
.B2(n_113),
.Y(n_166)
);

AND2x6_ASAP7_75t_L g167 ( 
.A(n_139),
.B(n_80),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_167),
.B(n_169),
.Y(n_188)
);

CKINVDCx12_ASAP7_75t_R g168 ( 
.A(n_135),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_168),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_146),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_146),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_170),
.B(n_176),
.Y(n_206)
);

OAI21xp33_ASAP7_75t_SL g173 ( 
.A1(n_138),
.A2(n_151),
.B(n_127),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_174),
.B(n_140),
.Y(n_195)
);

NAND2x1_ASAP7_75t_L g175 ( 
.A(n_153),
.B(n_121),
.Y(n_175)
);

OAI21xp33_ASAP7_75t_L g190 ( 
.A1(n_175),
.A2(n_152),
.B(n_165),
.Y(n_190)
);

AOI32xp33_ASAP7_75t_L g176 ( 
.A1(n_134),
.A2(n_125),
.A3(n_118),
.B1(n_116),
.B2(n_124),
.Y(n_176)
);

AND2x2_ASAP7_75t_L g178 ( 
.A(n_136),
.B(n_86),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_150),
.A2(n_110),
.B1(n_125),
.B2(n_100),
.Y(n_179)
);

AOI22xp33_ASAP7_75t_L g181 ( 
.A1(n_151),
.A2(n_95),
.B1(n_87),
.B2(n_60),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_181),
.A2(n_147),
.B1(n_101),
.B2(n_142),
.Y(n_189)
);

AND2x2_ASAP7_75t_L g183 ( 
.A(n_136),
.B(n_86),
.Y(n_183)
);

XOR2xp5_ASAP7_75t_L g186 ( 
.A(n_161),
.B(n_145),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_186),
.B(n_193),
.C(n_197),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_189),
.A2(n_196),
.B1(n_204),
.B2(n_208),
.Y(n_228)
);

AND2x2_ASAP7_75t_L g220 ( 
.A(n_190),
.B(n_215),
.Y(n_220)
);

AND2x2_ASAP7_75t_SL g191 ( 
.A(n_169),
.B(n_132),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_191),
.B(n_183),
.Y(n_217)
);

INVxp33_ASAP7_75t_SL g194 ( 
.A(n_156),
.Y(n_194)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_194),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_195),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_170),
.A2(n_131),
.B1(n_144),
.B2(n_143),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_182),
.B(n_149),
.C(n_101),
.Y(n_197)
);

INVx6_ASAP7_75t_L g199 ( 
.A(n_164),
.Y(n_199)
);

INVx3_ASAP7_75t_L g225 ( 
.A(n_199),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_155),
.B(n_126),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_200),
.B(n_202),
.Y(n_233)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_159),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g203 ( 
.A(n_182),
.B(n_90),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_203),
.B(n_180),
.C(n_177),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_154),
.A2(n_148),
.B1(n_137),
.B2(n_68),
.Y(n_204)
);

AO22x1_ASAP7_75t_L g205 ( 
.A1(n_179),
.A2(n_86),
.B1(n_129),
.B2(n_83),
.Y(n_205)
);

AOI22x1_ASAP7_75t_L g230 ( 
.A1(n_205),
.A2(n_175),
.B1(n_183),
.B2(n_172),
.Y(n_230)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_159),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_207),
.B(n_209),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_157),
.A2(n_70),
.B1(n_130),
.B2(n_88),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_185),
.B(n_120),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_167),
.A2(n_130),
.B1(n_88),
.B2(n_119),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_210),
.A2(n_174),
.B1(n_184),
.B2(n_177),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_184),
.B(n_129),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_211),
.B(n_212),
.Y(n_226)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_162),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_162),
.Y(n_213)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_213),
.Y(n_227)
);

OAI21xp5_ASAP7_75t_L g214 ( 
.A1(n_178),
.A2(n_106),
.B(n_79),
.Y(n_214)
);

OAI21xp5_ASAP7_75t_L g236 ( 
.A1(n_214),
.A2(n_174),
.B(n_171),
.Y(n_236)
);

AND2x4_ASAP7_75t_L g215 ( 
.A(n_178),
.B(n_108),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_198),
.B(n_164),
.Y(n_216)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_216),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_SL g259 ( 
.A(n_217),
.B(n_89),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_SL g219 ( 
.A(n_201),
.B(n_171),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_219),
.B(n_231),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_186),
.B(n_172),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_223),
.B(n_229),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_193),
.B(n_172),
.Y(n_229)
);

AOI22xp33_ASAP7_75t_L g247 ( 
.A1(n_230),
.A2(n_215),
.B1(n_192),
.B2(n_191),
.Y(n_247)
);

HB1xp67_ASAP7_75t_L g231 ( 
.A(n_199),
.Y(n_231)
);

XOR2xp5_ASAP7_75t_L g257 ( 
.A(n_232),
.B(n_234),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_187),
.B(n_175),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_L g258 ( 
.A1(n_235),
.A2(n_215),
.B1(n_190),
.B2(n_119),
.Y(n_258)
);

A2O1A1Ixp33_ASAP7_75t_SL g244 ( 
.A1(n_236),
.A2(n_214),
.B(n_205),
.C(n_215),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_197),
.B(n_180),
.C(n_163),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_237),
.B(n_238),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_187),
.B(n_163),
.Y(n_238)
);

OR2x2_ASAP7_75t_L g239 ( 
.A(n_200),
.B(n_94),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_239),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_221),
.A2(n_206),
.B1(n_188),
.B2(n_210),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_240),
.B(n_245),
.Y(n_274)
);

AOI21x1_ASAP7_75t_L g272 ( 
.A1(n_244),
.A2(n_1),
.B(n_2),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_218),
.B(n_203),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_247),
.A2(n_228),
.B1(n_222),
.B2(n_230),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_218),
.B(n_192),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_248),
.B(n_255),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_226),
.A2(n_204),
.B1(n_191),
.B2(n_208),
.Y(n_249)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_249),
.Y(n_262)
);

INVxp67_ASAP7_75t_L g251 ( 
.A(n_220),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_251),
.B(n_234),
.Y(n_268)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_233),
.Y(n_252)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_252),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_239),
.B(n_198),
.Y(n_253)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_253),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_224),
.B(n_195),
.Y(n_254)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_254),
.Y(n_276)
);

HB1xp67_ASAP7_75t_L g255 ( 
.A(n_225),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_227),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_256),
.B(n_258),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_259),
.B(n_2),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_260),
.A2(n_251),
.B1(n_244),
.B2(n_247),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_242),
.B(n_257),
.C(n_237),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_264),
.B(n_270),
.C(n_271),
.Y(n_284)
);

MAJx2_ASAP7_75t_L g266 ( 
.A(n_257),
.B(n_220),
.C(n_232),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_266),
.B(n_259),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_241),
.B(n_225),
.Y(n_267)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_267),
.Y(n_278)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_268),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_243),
.B(n_238),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_269),
.B(n_7),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_250),
.B(n_223),
.C(n_229),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_250),
.B(n_78),
.C(n_13),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g281 ( 
.A(n_272),
.B(n_275),
.Y(n_281)
);

XOR2xp5_ASAP7_75t_L g293 ( 
.A(n_277),
.B(n_270),
.Y(n_293)
);

OR2x2_ASAP7_75t_L g279 ( 
.A(n_273),
.B(n_246),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_279),
.A2(n_280),
.B1(n_283),
.B2(n_3),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_276),
.A2(n_244),
.B1(n_9),
.B2(n_4),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_282),
.B(n_285),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_262),
.A2(n_244),
.B1(n_9),
.B2(n_4),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_265),
.B(n_261),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_SL g294 ( 
.A(n_286),
.B(n_290),
.Y(n_294)
);

BUFx24_ASAP7_75t_SL g287 ( 
.A(n_263),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_287),
.B(n_289),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_272),
.Y(n_289)
);

BUFx24_ASAP7_75t_SL g290 ( 
.A(n_274),
.Y(n_290)
);

AOI21xp5_ASAP7_75t_L g291 ( 
.A1(n_279),
.A2(n_264),
.B(n_268),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_288),
.A2(n_260),
.B1(n_275),
.B2(n_266),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_292),
.B(n_299),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_L g303 ( 
.A(n_293),
.B(n_296),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_L g296 ( 
.A(n_284),
.B(n_271),
.Y(n_296)
);

BUFx6f_ASAP7_75t_L g298 ( 
.A(n_289),
.Y(n_298)
);

INVx11_ASAP7_75t_L g307 ( 
.A(n_298),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_SL g299 ( 
.A(n_278),
.B(n_2),
.Y(n_299)
);

AOI322xp5_ASAP7_75t_L g302 ( 
.A1(n_300),
.A2(n_3),
.A3(n_5),
.B1(n_6),
.B2(n_7),
.C1(n_281),
.C2(n_298),
.Y(n_302)
);

OA21x2_ASAP7_75t_SL g301 ( 
.A1(n_297),
.A2(n_281),
.B(n_5),
.Y(n_301)
);

AOI31xp67_ASAP7_75t_L g310 ( 
.A1(n_301),
.A2(n_308),
.A3(n_307),
.B(n_304),
.Y(n_310)
);

CKINVDCx16_ASAP7_75t_R g311 ( 
.A(n_302),
.Y(n_311)
);

OAI21xp5_ASAP7_75t_L g304 ( 
.A1(n_292),
.A2(n_3),
.B(n_5),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_304),
.B(n_306),
.Y(n_312)
);

AOI322xp5_ASAP7_75t_L g306 ( 
.A1(n_294),
.A2(n_5),
.A3(n_6),
.B1(n_7),
.B2(n_296),
.C1(n_295),
.C2(n_293),
.Y(n_306)
);

OAI21x1_ASAP7_75t_L g308 ( 
.A1(n_291),
.A2(n_6),
.B(n_7),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_307),
.B(n_6),
.Y(n_309)
);

INVxp67_ASAP7_75t_L g314 ( 
.A(n_309),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_310),
.B(n_313),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_305),
.B(n_303),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_314),
.B(n_311),
.Y(n_316)
);

XOR2xp5_ASAP7_75t_L g318 ( 
.A(n_316),
.B(n_317),
.Y(n_318)
);

AOI21xp5_ASAP7_75t_L g317 ( 
.A1(n_315),
.A2(n_312),
.B(n_305),
.Y(n_317)
);

BUFx24_ASAP7_75t_SL g319 ( 
.A(n_318),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_L g320 ( 
.A(n_319),
.B(n_309),
.Y(n_320)
);


endmodule