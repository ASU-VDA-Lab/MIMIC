module real_jpeg_1109_n_7 (n_5, n_4, n_40, n_0, n_43, n_1, n_41, n_2, n_45, n_6, n_42, n_44, n_3, n_7);

input n_5;
input n_4;
input n_40;
input n_0;
input n_43;
input n_1;
input n_41;
input n_2;
input n_45;
input n_6;
input n_42;
input n_44;
input n_3;

output n_7;

wire n_17;
wire n_8;
wire n_37;
wire n_21;
wire n_33;
wire n_35;
wire n_29;
wire n_10;
wire n_31;
wire n_9;
wire n_12;
wire n_24;
wire n_34;
wire n_28;
wire n_23;
wire n_11;
wire n_14;
wire n_25;
wire n_22;
wire n_18;
wire n_36;
wire n_27;
wire n_26;
wire n_20;
wire n_19;
wire n_32;
wire n_30;
wire n_16;
wire n_15;
wire n_13;

OAI21xp5_ASAP7_75t_SL g20 ( 
.A1(n_0),
.A2(n_21),
.B(n_25),
.Y(n_20)
);

BUFx16f_ASAP7_75t_L g10 ( 
.A(n_1),
.Y(n_10)
);

INVx3_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

BUFx4f_ASAP7_75t_SL g24 ( 
.A(n_1),
.Y(n_24)
);

AND2x2_ASAP7_75t_L g21 ( 
.A(n_2),
.B(n_22),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_3),
.Y(n_33)
);

MAJIxp5_ASAP7_75t_L g13 ( 
.A(n_4),
.B(n_14),
.C(n_30),
.Y(n_13)
);

AO22x1_ASAP7_75t_L g14 ( 
.A1(n_5),
.A2(n_15),
.B1(n_19),
.B2(n_29),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_5),
.Y(n_28)
);

FAx1_ASAP7_75t_SL g7 ( 
.A(n_6),
.B(n_8),
.CI(n_11),
.CON(n_7),
.SN(n_7)
);

NOR2xp33_ASAP7_75t_L g8 ( 
.A(n_9),
.B(n_10),
.Y(n_8)
);

HB1xp67_ASAP7_75t_L g11 ( 
.A(n_12),
.Y(n_11)
);

MAJIxp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_33),
.C(n_34),
.Y(n_12)
);

NOR2xp33_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_17),
.Y(n_15)
);

INVx5_ASAP7_75t_L g17 ( 
.A(n_18),
.Y(n_17)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_18),
.Y(n_32)
);

INVx6_ASAP7_75t_SL g37 ( 
.A(n_18),
.Y(n_37)
);

NAND3xp33_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_27),
.C(n_28),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_20),
.B(n_27),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_21),
.B(n_25),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_24),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_24),
.B(n_26),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_31),
.B(n_32),
.Y(n_30)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_36),
.B(n_37),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g9 ( 
.A(n_40),
.Y(n_9)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_41),
.Y(n_16)
);

CKINVDCx16_ASAP7_75t_R g23 ( 
.A(n_42),
.Y(n_23)
);

CKINVDCx16_ASAP7_75t_R g26 ( 
.A(n_43),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_44),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_45),
.Y(n_36)
);


endmodule