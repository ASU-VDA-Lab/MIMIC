module fake_jpeg_28395_n_224 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_224);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_224;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_171;
wire n_119;
wire n_23;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_212;
wire n_131;
wire n_56;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_96;

BUFx10_ASAP7_75t_L g15 ( 
.A(n_13),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_8),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_10),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

BUFx10_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_13),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_4),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_10),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_6),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_9),
.Y(n_26)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_10),
.Y(n_28)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_9),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_8),
.Y(n_31)
);

MAJIxp5_ASAP7_75t_L g32 ( 
.A(n_18),
.B(n_0),
.C(n_1),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_32),
.B(n_34),
.Y(n_58)
);

INVx11_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_33),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_18),
.B(n_0),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_18),
.Y(n_35)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_35),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_16),
.B(n_1),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_36),
.B(n_37),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_16),
.B(n_1),
.Y(n_37)
);

INVx4_ASAP7_75t_SL g38 ( 
.A(n_15),
.Y(n_38)
);

CKINVDCx16_ASAP7_75t_R g57 ( 
.A(n_38),
.Y(n_57)
);

OR2x2_ASAP7_75t_SL g39 ( 
.A(n_16),
.B(n_2),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_SL g56 ( 
.A1(n_39),
.A2(n_22),
.B1(n_30),
.B2(n_24),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_15),
.Y(n_40)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_40),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g41 ( 
.A(n_17),
.B(n_2),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g47 ( 
.A(n_41),
.B(n_22),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_27),
.Y(n_42)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_42),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_41),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_46),
.B(n_47),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_38),
.A2(n_29),
.B1(n_27),
.B2(n_30),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_48),
.A2(n_53),
.B1(n_29),
.B2(n_27),
.Y(n_64)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_50),
.B(n_56),
.Y(n_66)
);

BUFx4f_ASAP7_75t_SL g51 ( 
.A(n_38),
.Y(n_51)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_51),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_37),
.B(n_22),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_52),
.B(n_54),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_38),
.A2(n_29),
.B1(n_27),
.B2(n_30),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_32),
.B(n_20),
.Y(n_54)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_42),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_55),
.B(n_42),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_39),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_59),
.B(n_60),
.Y(n_72)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_34),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_32),
.B(n_20),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_62),
.B(n_20),
.Y(n_70)
);

BUFx10_ASAP7_75t_L g63 ( 
.A(n_33),
.Y(n_63)
);

INVxp67_ASAP7_75t_L g71 ( 
.A(n_63),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_64),
.A2(n_43),
.B1(n_26),
.B2(n_25),
.Y(n_96)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_61),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_67),
.B(n_76),
.Y(n_86)
);

NAND2xp33_ASAP7_75t_SL g68 ( 
.A(n_54),
.B(n_39),
.Y(n_68)
);

AND2x2_ASAP7_75t_L g87 ( 
.A(n_68),
.B(n_70),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_60),
.B(n_25),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_73),
.B(n_81),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_62),
.B(n_35),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_75),
.B(n_78),
.Y(n_89)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_44),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_59),
.A2(n_29),
.B1(n_31),
.B2(n_24),
.Y(n_77)
);

INVxp67_ASAP7_75t_L g105 ( 
.A(n_77),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_58),
.B(n_56),
.Y(n_78)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_44),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_79),
.B(n_80),
.Y(n_93)
);

INVxp67_ASAP7_75t_L g80 ( 
.A(n_51),
.Y(n_80)
);

NAND3xp33_ASAP7_75t_L g81 ( 
.A(n_49),
.B(n_2),
.C(n_3),
.Y(n_81)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_61),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_82),
.B(n_61),
.Y(n_95)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_83),
.Y(n_94)
);

OAI32xp33_ASAP7_75t_L g84 ( 
.A1(n_70),
.A2(n_46),
.A3(n_47),
.B1(n_52),
.B2(n_50),
.Y(n_84)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_84),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_75),
.A2(n_43),
.B1(n_45),
.B2(n_55),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_85),
.A2(n_92),
.B1(n_100),
.B2(n_20),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_69),
.B(n_51),
.C(n_57),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_88),
.B(n_98),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_83),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_90),
.Y(n_115)
);

AND2x2_ASAP7_75t_L g91 ( 
.A(n_78),
.B(n_35),
.Y(n_91)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_91),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_69),
.A2(n_43),
.B1(n_45),
.B2(n_33),
.Y(n_92)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_95),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_96),
.A2(n_64),
.B1(n_74),
.B2(n_71),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_65),
.B(n_73),
.Y(n_98)
);

HB1xp67_ASAP7_75t_L g99 ( 
.A(n_76),
.Y(n_99)
);

CKINVDCx16_ASAP7_75t_R g108 ( 
.A(n_99),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_66),
.A2(n_57),
.B1(n_35),
.B2(n_49),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_65),
.B(n_17),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_101),
.B(n_104),
.Y(n_112)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_77),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_102),
.B(n_103),
.Y(n_109)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_72),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_66),
.B(n_51),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_107),
.A2(n_111),
.B1(n_119),
.B2(n_120),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_102),
.A2(n_105),
.B1(n_89),
.B2(n_88),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_90),
.B(n_74),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_SL g141 ( 
.A(n_113),
.B(n_114),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_103),
.B(n_79),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_89),
.B(n_72),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_117),
.B(n_123),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_104),
.A2(n_68),
.B1(n_67),
.B2(n_82),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_94),
.A2(n_82),
.B1(n_42),
.B2(n_63),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_94),
.A2(n_63),
.B1(n_40),
.B2(n_19),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_121),
.A2(n_122),
.B1(n_126),
.B2(n_107),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_85),
.A2(n_63),
.B1(n_40),
.B2(n_19),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_87),
.B(n_81),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_124),
.B(n_95),
.Y(n_140)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_86),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_125),
.B(n_108),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_98),
.A2(n_92),
.B1(n_84),
.B2(n_97),
.Y(n_126)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_120),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_127),
.B(n_132),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_117),
.B(n_101),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_128),
.B(n_130),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_L g129 ( 
.A1(n_116),
.A2(n_87),
.B(n_91),
.Y(n_129)
);

AOI21xp5_ASAP7_75t_L g162 ( 
.A1(n_129),
.A2(n_110),
.B(n_123),
.Y(n_162)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_109),
.Y(n_130)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_121),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_115),
.B(n_87),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_134),
.B(n_135),
.Y(n_155)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_122),
.Y(n_135)
);

CKINVDCx14_ASAP7_75t_R g136 ( 
.A(n_112),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_136),
.B(n_139),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_116),
.A2(n_91),
.B1(n_100),
.B2(n_86),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_137),
.A2(n_140),
.B1(n_126),
.B2(n_110),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_138),
.A2(n_135),
.B1(n_132),
.B2(n_127),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_115),
.B(n_97),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_L g142 ( 
.A(n_106),
.B(n_93),
.Y(n_142)
);

XOR2xp5_ASAP7_75t_L g151 ( 
.A(n_142),
.B(n_144),
.Y(n_151)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_112),
.Y(n_143)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_143),
.Y(n_158)
);

XOR2xp5_ASAP7_75t_L g144 ( 
.A(n_106),
.B(n_93),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_125),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_145),
.B(n_118),
.Y(n_160)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_146),
.Y(n_152)
);

INVxp67_ASAP7_75t_L g148 ( 
.A(n_141),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_148),
.B(n_154),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_144),
.B(n_111),
.C(n_119),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_149),
.B(n_19),
.C(n_40),
.Y(n_174)
);

INVxp67_ASAP7_75t_L g154 ( 
.A(n_133),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_156),
.B(n_163),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_157),
.A2(n_129),
.B1(n_142),
.B2(n_131),
.Y(n_166)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_145),
.Y(n_159)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_159),
.Y(n_170)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_160),
.Y(n_172)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_134),
.Y(n_161)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_161),
.Y(n_173)
);

XOR2xp5_ASAP7_75t_L g176 ( 
.A(n_162),
.B(n_20),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_137),
.A2(n_118),
.B1(n_124),
.B2(n_31),
.Y(n_163)
);

AOI21xp5_ASAP7_75t_L g164 ( 
.A1(n_133),
.A2(n_3),
.B(n_4),
.Y(n_164)
);

O2A1O1Ixp33_ASAP7_75t_L g168 ( 
.A1(n_164),
.A2(n_17),
.B(n_28),
.C(n_26),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_154),
.A2(n_157),
.B1(n_138),
.B2(n_147),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_165),
.B(n_166),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_152),
.A2(n_131),
.B1(n_31),
.B2(n_28),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_167),
.B(n_171),
.Y(n_190)
);

AOI22xp33_ASAP7_75t_L g180 ( 
.A1(n_168),
.A2(n_23),
.B1(n_21),
.B2(n_153),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_147),
.A2(n_24),
.B1(n_28),
.B2(n_26),
.Y(n_171)
);

XOR2xp5_ASAP7_75t_L g181 ( 
.A(n_174),
.B(n_176),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_152),
.A2(n_25),
.B1(n_23),
.B2(n_21),
.Y(n_177)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_177),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_151),
.B(n_19),
.C(n_20),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_178),
.B(n_160),
.C(n_155),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g179 ( 
.A(n_151),
.B(n_20),
.Y(n_179)
);

XOR2xp5_ASAP7_75t_L g183 ( 
.A(n_179),
.B(n_149),
.Y(n_183)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_180),
.Y(n_197)
);

NOR3xp33_ASAP7_75t_SL g182 ( 
.A(n_175),
.B(n_148),
.C(n_162),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_182),
.B(n_187),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_L g198 ( 
.A(n_183),
.B(n_184),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_179),
.B(n_156),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_186),
.B(n_174),
.C(n_178),
.Y(n_194)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_171),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_173),
.A2(n_158),
.B1(n_164),
.B2(n_163),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_188),
.B(n_189),
.Y(n_196)
);

AOI21xp5_ASAP7_75t_L g189 ( 
.A1(n_169),
.A2(n_155),
.B(n_150),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_185),
.A2(n_172),
.B1(n_170),
.B2(n_165),
.Y(n_192)
);

OR2x2_ASAP7_75t_L g204 ( 
.A(n_192),
.B(n_195),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_194),
.B(n_199),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_SL g195 ( 
.A(n_190),
.B(n_168),
.Y(n_195)
);

HB1xp67_ASAP7_75t_L g199 ( 
.A(n_184),
.Y(n_199)
);

BUFx24_ASAP7_75t_SL g200 ( 
.A(n_183),
.Y(n_200)
);

NAND3xp33_ASAP7_75t_L g205 ( 
.A(n_200),
.B(n_14),
.C(n_186),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_SL g201 ( 
.A1(n_193),
.A2(n_188),
.B(n_182),
.Y(n_201)
);

AOI21xp5_ASAP7_75t_L g212 ( 
.A1(n_201),
.A2(n_7),
.B(n_8),
.Y(n_212)
);

AOI31xp33_ASAP7_75t_L g203 ( 
.A1(n_196),
.A2(n_169),
.A3(n_191),
.B(n_176),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_203),
.B(n_205),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_197),
.A2(n_181),
.B1(n_23),
.B2(n_21),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_L g209 ( 
.A1(n_206),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_209)
);

NAND3xp33_ASAP7_75t_L g207 ( 
.A(n_199),
.B(n_181),
.C(n_14),
.Y(n_207)
);

OAI21xp5_ASAP7_75t_L g208 ( 
.A1(n_207),
.A2(n_3),
.B(n_4),
.Y(n_208)
);

AO21x1_ASAP7_75t_L g214 ( 
.A1(n_208),
.A2(n_212),
.B(n_7),
.Y(n_214)
);

AND2x2_ASAP7_75t_L g216 ( 
.A(n_209),
.B(n_11),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_204),
.B(n_198),
.Y(n_211)
);

AOI21xp5_ASAP7_75t_L g217 ( 
.A1(n_211),
.A2(n_213),
.B(n_11),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_202),
.B(n_19),
.Y(n_213)
);

AOI21xp5_ASAP7_75t_SL g220 ( 
.A1(n_214),
.A2(n_12),
.B(n_15),
.Y(n_220)
);

FAx1_ASAP7_75t_SL g215 ( 
.A(n_210),
.B(n_207),
.CI(n_12),
.CON(n_215),
.SN(n_215)
);

XNOR2xp5_ASAP7_75t_L g218 ( 
.A(n_215),
.B(n_217),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_216),
.B(n_11),
.C(n_12),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_219),
.B(n_15),
.C(n_218),
.Y(n_221)
);

INVxp33_ASAP7_75t_L g222 ( 
.A(n_220),
.Y(n_222)
);

OAI21xp5_ASAP7_75t_L g223 ( 
.A1(n_221),
.A2(n_15),
.B(n_222),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_223),
.B(n_15),
.Y(n_224)
);


endmodule