module fake_jpeg_24691_n_322 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_322);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_322;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_145;
wire n_18;
wire n_20;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_3),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_2),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_16),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_10),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_1),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_8),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_28),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_SL g50 ( 
.A(n_35),
.B(n_39),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_28),
.Y(n_36)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_36),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_28),
.Y(n_37)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_37),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_19),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_38),
.B(n_44),
.Y(n_45)
);

AND2x2_ASAP7_75t_L g39 ( 
.A(n_28),
.B(n_0),
.Y(n_39)
);

BUFx10_ASAP7_75t_L g40 ( 
.A(n_28),
.Y(n_40)
);

INVx1_ASAP7_75t_SL g61 ( 
.A(n_40),
.Y(n_61)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_26),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_41),
.B(n_0),
.Y(n_69)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_29),
.Y(n_42)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_42),
.Y(n_48)
);

BUFx5_ASAP7_75t_L g43 ( 
.A(n_33),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g67 ( 
.A(n_43),
.Y(n_67)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_33),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_43),
.Y(n_46)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_46),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_L g47 ( 
.A(n_35),
.B(n_29),
.C(n_33),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_47),
.B(n_60),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_SL g49 ( 
.A1(n_39),
.A2(n_29),
.B1(n_34),
.B2(n_26),
.Y(n_49)
);

OAI22x1_ASAP7_75t_L g86 ( 
.A1(n_49),
.A2(n_57),
.B1(n_58),
.B2(n_63),
.Y(n_86)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_43),
.Y(n_51)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_51),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_38),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_52),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_38),
.B(n_27),
.Y(n_53)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_53),
.Y(n_89)
);

NOR2x1_ASAP7_75t_L g55 ( 
.A(n_39),
.B(n_29),
.Y(n_55)
);

OR2x2_ASAP7_75t_L g87 ( 
.A(n_55),
.B(n_62),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_39),
.B(n_17),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_56),
.B(n_23),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g57 ( 
.A1(n_41),
.A2(n_44),
.B1(n_39),
.B2(n_26),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_41),
.A2(n_29),
.B1(n_34),
.B2(n_31),
.Y(n_58)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_36),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_42),
.B(n_21),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_44),
.A2(n_34),
.B1(n_21),
.B2(n_32),
.Y(n_63)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_36),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_64),
.B(n_66),
.Y(n_83)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_36),
.Y(n_65)
);

INVx6_ASAP7_75t_L g84 ( 
.A(n_65),
.Y(n_84)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_37),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_44),
.A2(n_32),
.B1(n_31),
.B2(n_23),
.Y(n_68)
);

CKINVDCx16_ASAP7_75t_R g85 ( 
.A(n_68),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_69),
.B(n_27),
.Y(n_93)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_59),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_71),
.B(n_75),
.Y(n_100)
);

INVx6_ASAP7_75t_SL g73 ( 
.A(n_67),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_73),
.B(n_76),
.Y(n_98)
);

XOR2xp5_ASAP7_75t_L g122 ( 
.A(n_74),
.B(n_22),
.Y(n_122)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_59),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_52),
.Y(n_76)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_59),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_77),
.B(n_79),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_56),
.B(n_40),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_78),
.B(n_82),
.Y(n_107)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_67),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_45),
.B(n_53),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_81),
.B(n_92),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_50),
.B(n_45),
.Y(n_82)
);

INVx5_ASAP7_75t_L g90 ( 
.A(n_54),
.Y(n_90)
);

INVx4_ASAP7_75t_L g97 ( 
.A(n_90),
.Y(n_97)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_67),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_91),
.B(n_61),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_62),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_93),
.B(n_19),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_50),
.B(n_55),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_94),
.B(n_57),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_67),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_95),
.Y(n_118)
);

OR2x2_ASAP7_75t_L g96 ( 
.A(n_70),
.B(n_55),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_96),
.B(n_112),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_70),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_99),
.Y(n_125)
);

BUFx3_ASAP7_75t_L g101 ( 
.A(n_73),
.Y(n_101)
);

INVx4_ASAP7_75t_L g145 ( 
.A(n_101),
.Y(n_145)
);

AOI21xp5_ASAP7_75t_SL g103 ( 
.A1(n_94),
.A2(n_69),
.B(n_49),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_SL g124 ( 
.A1(n_103),
.A2(n_86),
.B(n_92),
.Y(n_124)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_83),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_104),
.B(n_106),
.Y(n_131)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_72),
.Y(n_106)
);

OAI21xp33_ASAP7_75t_L g152 ( 
.A1(n_108),
.A2(n_0),
.B(n_1),
.Y(n_152)
);

OA22x2_ASAP7_75t_L g109 ( 
.A1(n_85),
.A2(n_40),
.B1(n_61),
.B2(n_47),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_109),
.A2(n_110),
.B1(n_54),
.B2(n_71),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_86),
.A2(n_48),
.B1(n_42),
.B2(n_35),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_111),
.B(n_113),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_78),
.B(n_48),
.Y(n_112)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_84),
.Y(n_113)
);

INVx13_ASAP7_75t_L g114 ( 
.A(n_91),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_114),
.B(n_116),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_89),
.B(n_51),
.Y(n_115)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_115),
.Y(n_128)
);

INVx13_ASAP7_75t_L g116 ( 
.A(n_95),
.Y(n_116)
);

CKINVDCx14_ASAP7_75t_R g133 ( 
.A(n_117),
.Y(n_133)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_84),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_119),
.B(n_120),
.Y(n_140)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_74),
.Y(n_120)
);

AND2x2_ASAP7_75t_SL g121 ( 
.A(n_82),
.B(n_40),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_L g127 ( 
.A1(n_121),
.A2(n_87),
.B(n_88),
.Y(n_127)
);

XNOR2xp5_ASAP7_75t_L g149 ( 
.A(n_122),
.B(n_22),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_76),
.B(n_40),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_123),
.B(n_88),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_SL g180 ( 
.A1(n_124),
.A2(n_109),
.B(n_65),
.Y(n_180)
);

AOI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_97),
.A2(n_90),
.B1(n_80),
.B2(n_51),
.Y(n_126)
);

INVxp67_ASAP7_75t_L g167 ( 
.A(n_126),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_L g159 ( 
.A1(n_127),
.A2(n_121),
.B(n_96),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_105),
.B(n_89),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_129),
.B(n_138),
.Y(n_181)
);

INVxp67_ASAP7_75t_L g132 ( 
.A(n_102),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_132),
.B(n_142),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_134),
.A2(n_150),
.B1(n_106),
.B2(n_64),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_99),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_135),
.Y(n_154)
);

A2O1A1O1Ixp25_ASAP7_75t_L g139 ( 
.A1(n_103),
.A2(n_87),
.B(n_40),
.C(n_37),
.D(n_22),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_139),
.B(n_109),
.C(n_104),
.Y(n_172)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_101),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_141),
.B(n_151),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_98),
.B(n_123),
.Y(n_142)
);

XNOR2xp5_ASAP7_75t_SL g143 ( 
.A(n_110),
.B(n_40),
.Y(n_143)
);

XOR2xp5_ASAP7_75t_L g179 ( 
.A(n_143),
.B(n_149),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_98),
.B(n_79),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_144),
.B(n_146),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_105),
.B(n_80),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_107),
.B(n_46),
.Y(n_147)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_147),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_107),
.B(n_46),
.Y(n_148)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_148),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_108),
.A2(n_54),
.B1(n_66),
.B2(n_77),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_115),
.B(n_75),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_152),
.B(n_2),
.Y(n_156)
);

AOI22xp33_ASAP7_75t_SL g153 ( 
.A1(n_145),
.A2(n_97),
.B1(n_113),
.B2(n_119),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_153),
.A2(n_60),
.B1(n_118),
.B2(n_25),
.Y(n_208)
);

NAND2xp67_ASAP7_75t_SL g193 ( 
.A(n_156),
.B(n_176),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_157),
.B(n_169),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_124),
.A2(n_130),
.B1(n_148),
.B2(n_147),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_158),
.A2(n_168),
.B1(n_174),
.B2(n_180),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_SL g205 ( 
.A(n_159),
.B(n_111),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_125),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_161),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_L g163 ( 
.A1(n_127),
.A2(n_121),
.B(n_96),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_163),
.B(n_166),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_125),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_164),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_135),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_165),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_145),
.B(n_114),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_130),
.A2(n_112),
.B1(n_109),
.B2(n_120),
.Y(n_168)
);

INVxp67_ASAP7_75t_L g169 ( 
.A(n_137),
.Y(n_169)
);

FAx1_ASAP7_75t_SL g170 ( 
.A(n_138),
.B(n_121),
.CI(n_122),
.CON(n_170),
.SN(n_170)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_170),
.B(n_172),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_134),
.A2(n_150),
.B1(n_143),
.B2(n_139),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_140),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_175),
.B(n_128),
.Y(n_192)
);

NOR2x1_ASAP7_75t_L g176 ( 
.A(n_129),
.B(n_109),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_141),
.B(n_114),
.Y(n_177)
);

CKINVDCx16_ASAP7_75t_R g209 ( 
.A(n_177),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_137),
.B(n_100),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_178),
.Y(n_184)
);

HB1xp67_ASAP7_75t_L g182 ( 
.A(n_151),
.Y(n_182)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_182),
.Y(n_186)
);

INVxp67_ASAP7_75t_L g183 ( 
.A(n_144),
.Y(n_183)
);

INVxp33_ASAP7_75t_SL g191 ( 
.A(n_183),
.Y(n_191)
);

AND2x2_ASAP7_75t_L g187 ( 
.A(n_176),
.B(n_149),
.Y(n_187)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_187),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_179),
.B(n_142),
.C(n_140),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_189),
.B(n_197),
.C(n_206),
.Y(n_211)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_160),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_190),
.B(n_196),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_192),
.Y(n_228)
);

XOR2x2_ASAP7_75t_L g194 ( 
.A(n_176),
.B(n_146),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_SL g230 ( 
.A(n_194),
.B(n_24),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_181),
.B(n_128),
.Y(n_195)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_195),
.Y(n_233)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_181),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_179),
.B(n_131),
.C(n_133),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_173),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_198),
.B(n_203),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_155),
.B(n_131),
.Y(n_199)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_199),
.Y(n_234)
);

NOR2xp67_ASAP7_75t_L g201 ( 
.A(n_170),
.B(n_136),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_SL g225 ( 
.A(n_201),
.B(n_30),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_155),
.B(n_136),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_205),
.B(n_156),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_171),
.B(n_95),
.C(n_37),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_L g223 ( 
.A1(n_208),
.A2(n_167),
.B1(n_183),
.B2(n_169),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_204),
.A2(n_167),
.B1(n_158),
.B2(n_168),
.Y(n_212)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_212),
.Y(n_239)
);

INVxp67_ASAP7_75t_L g214 ( 
.A(n_191),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_214),
.B(n_218),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_189),
.B(n_171),
.C(n_163),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_215),
.B(n_216),
.C(n_220),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_197),
.B(n_159),
.C(n_170),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_194),
.A2(n_180),
.B1(n_174),
.B2(n_157),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_217),
.A2(n_18),
.B1(n_17),
.B2(n_20),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_185),
.B(n_154),
.Y(n_218)
);

OAI21xp5_ASAP7_75t_L g219 ( 
.A1(n_210),
.A2(n_161),
.B(n_154),
.Y(n_219)
);

AOI21xp5_ASAP7_75t_L g251 ( 
.A1(n_219),
.A2(n_25),
.B(n_18),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_207),
.B(n_172),
.C(n_162),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_205),
.B(n_175),
.C(n_165),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_221),
.B(n_224),
.C(n_226),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g236 ( 
.A(n_222),
.B(n_230),
.Y(n_236)
);

AOI322xp5_ASAP7_75t_L g244 ( 
.A1(n_223),
.A2(n_193),
.A3(n_187),
.B1(n_184),
.B2(n_190),
.C1(n_186),
.C2(n_198),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_196),
.B(n_164),
.C(n_118),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_225),
.B(n_20),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_200),
.B(n_118),
.C(n_116),
.Y(n_226)
);

HB1xp67_ASAP7_75t_L g229 ( 
.A(n_188),
.Y(n_229)
);

INVx1_ASAP7_75t_SL g238 ( 
.A(n_229),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_SL g231 ( 
.A(n_200),
.B(n_24),
.Y(n_231)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_231),
.B(n_206),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_202),
.B(n_116),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_235),
.B(n_209),
.Y(n_245)
);

OAI21xp5_ASAP7_75t_SL g242 ( 
.A1(n_213),
.A2(n_192),
.B(n_193),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_242),
.B(n_222),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_243),
.B(n_247),
.Y(n_264)
);

BUFx24_ASAP7_75t_SL g271 ( 
.A(n_244),
.Y(n_271)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_245),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_211),
.B(n_195),
.C(n_203),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_246),
.B(n_250),
.C(n_255),
.Y(n_262)
);

OAI322xp33_ASAP7_75t_L g247 ( 
.A1(n_232),
.A2(n_199),
.A3(n_187),
.B1(n_184),
.B2(n_186),
.C1(n_208),
.C2(n_30),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_SL g259 ( 
.A(n_248),
.B(n_251),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_SL g249 ( 
.A(n_216),
.B(n_24),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_249),
.B(n_231),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_211),
.B(n_215),
.C(n_221),
.Y(n_250)
);

BUFx12_ASAP7_75t_L g252 ( 
.A(n_214),
.Y(n_252)
);

INVx11_ASAP7_75t_L g266 ( 
.A(n_252),
.Y(n_266)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_253),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_224),
.B(n_4),
.Y(n_254)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_254),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_220),
.B(n_5),
.C(n_6),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_230),
.B(n_5),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_256),
.B(n_226),
.C(n_228),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_257),
.B(n_241),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_SL g273 ( 
.A(n_258),
.B(n_261),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_SL g261 ( 
.A(n_246),
.B(n_227),
.Y(n_261)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_240),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_263),
.B(n_238),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_265),
.B(n_241),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_252),
.B(n_233),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_SL g274 ( 
.A(n_267),
.B(n_270),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_250),
.B(n_234),
.Y(n_269)
);

XOR2xp5_ASAP7_75t_L g280 ( 
.A(n_269),
.B(n_236),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_252),
.B(n_5),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_275),
.B(n_277),
.Y(n_292)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_276),
.Y(n_291)
);

AND2x2_ASAP7_75t_SL g278 ( 
.A(n_263),
.B(n_243),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_278),
.B(n_279),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_SL g279 ( 
.A(n_259),
.B(n_239),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_280),
.B(n_272),
.C(n_257),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_268),
.B(n_238),
.Y(n_281)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_281),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_260),
.B(n_253),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_SL g293 ( 
.A(n_282),
.B(n_284),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_262),
.B(n_237),
.C(n_249),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_283),
.B(n_256),
.C(n_264),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_266),
.B(n_255),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_265),
.B(n_237),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g295 ( 
.A(n_285),
.B(n_286),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_L g286 ( 
.A(n_262),
.B(n_236),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_287),
.B(n_288),
.C(n_289),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_283),
.B(n_269),
.C(n_264),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_278),
.B(n_273),
.C(n_280),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_290),
.B(n_297),
.C(n_7),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_275),
.B(n_266),
.C(n_271),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_SL g298 ( 
.A(n_274),
.B(n_7),
.Y(n_298)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_298),
.Y(n_302)
);

XOR2xp5_ASAP7_75t_L g314 ( 
.A(n_300),
.B(n_303),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_288),
.B(n_7),
.C(n_8),
.Y(n_301)
);

AOI21xp5_ASAP7_75t_L g313 ( 
.A1(n_301),
.A2(n_304),
.B(n_12),
.Y(n_313)
);

XOR2xp5_ASAP7_75t_L g303 ( 
.A(n_292),
.B(n_294),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_291),
.B(n_8),
.Y(n_304)
);

XOR2xp5_ASAP7_75t_L g305 ( 
.A(n_295),
.B(n_9),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_305),
.B(n_306),
.Y(n_308)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_293),
.Y(n_306)
);

AOI21x1_ASAP7_75t_L g307 ( 
.A1(n_296),
.A2(n_9),
.B(n_10),
.Y(n_307)
);

OA21x2_ASAP7_75t_L g309 ( 
.A1(n_307),
.A2(n_9),
.B(n_11),
.Y(n_309)
);

AOI21xp5_ASAP7_75t_L g316 ( 
.A1(n_309),
.A2(n_310),
.B(n_312),
.Y(n_316)
);

OAI21xp5_ASAP7_75t_SL g310 ( 
.A1(n_299),
.A2(n_287),
.B(n_12),
.Y(n_310)
);

AOI322xp5_ASAP7_75t_L g311 ( 
.A1(n_305),
.A2(n_11),
.A3(n_12),
.B1(n_13),
.B2(n_14),
.C1(n_15),
.C2(n_16),
.Y(n_311)
);

AOI322xp5_ASAP7_75t_L g315 ( 
.A1(n_311),
.A2(n_313),
.A3(n_302),
.B1(n_14),
.B2(n_15),
.C1(n_16),
.C2(n_13),
.Y(n_315)
);

INVxp67_ASAP7_75t_L g312 ( 
.A(n_303),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_315),
.B(n_317),
.C(n_309),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_314),
.B(n_13),
.C(n_14),
.Y(n_317)
);

INVxp67_ASAP7_75t_L g318 ( 
.A(n_308),
.Y(n_318)
);

INVxp67_ASAP7_75t_L g320 ( 
.A(n_318),
.Y(n_320)
);

OAI21xp5_ASAP7_75t_SL g321 ( 
.A1(n_319),
.A2(n_316),
.B(n_15),
.Y(n_321)
);

XNOR2xp5_ASAP7_75t_L g322 ( 
.A(n_321),
.B(n_320),
.Y(n_322)
);


endmodule