module fake_jpeg_25478_n_94 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_94);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_94;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_57;
wire n_21;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;

BUFx10_ASAP7_75t_L g11 ( 
.A(n_0),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_9),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_0),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_L g14 ( 
.A(n_6),
.B(n_8),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_9),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_10),
.Y(n_16)
);

BUFx10_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_6),
.Y(n_18)
);

BUFx12_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

BUFx10_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_8),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_3),
.Y(n_22)
);

AND2x2_ASAP7_75t_SL g23 ( 
.A(n_11),
.B(n_0),
.Y(n_23)
);

AOI21xp5_ASAP7_75t_L g35 ( 
.A1(n_23),
.A2(n_1),
.B(n_11),
.Y(n_35)
);

INVx2_ASAP7_75t_SL g24 ( 
.A(n_11),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_24),
.B(n_29),
.Y(n_37)
);

INVx6_ASAP7_75t_L g25 ( 
.A(n_17),
.Y(n_25)
);

BUFx2_ASAP7_75t_L g34 ( 
.A(n_25),
.Y(n_34)
);

INVx8_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_26),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_19),
.Y(n_27)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_27),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_14),
.B(n_1),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_28),
.B(n_30),
.Y(n_39)
);

INVx5_ASAP7_75t_L g29 ( 
.A(n_17),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_17),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_SL g31 ( 
.A(n_28),
.B(n_14),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_SL g46 ( 
.A(n_31),
.B(n_38),
.Y(n_46)
);

AOI21xp5_ASAP7_75t_SL g33 ( 
.A1(n_23),
.A2(n_13),
.B(n_15),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_33),
.B(n_40),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_35),
.B(n_17),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_23),
.B(n_22),
.Y(n_38)
);

CKINVDCx16_ASAP7_75t_R g40 ( 
.A(n_23),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_27),
.B(n_16),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_41),
.B(n_12),
.Y(n_48)
);

AOI21xp5_ASAP7_75t_L g43 ( 
.A1(n_35),
.A2(n_11),
.B(n_17),
.Y(n_43)
);

AOI21xp5_ASAP7_75t_SL g60 ( 
.A1(n_43),
.A2(n_45),
.B(n_20),
.Y(n_60)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_34),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_44),
.B(n_47),
.Y(n_59)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_34),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_48),
.B(n_16),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g49 ( 
.A1(n_39),
.A2(n_25),
.B1(n_18),
.B2(n_12),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_49),
.B(n_50),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g50 ( 
.A1(n_32),
.A2(n_25),
.B1(n_30),
.B2(n_29),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_51),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_SL g53 ( 
.A(n_46),
.B(n_33),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_SL g67 ( 
.A(n_53),
.B(n_55),
.Y(n_67)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_50),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_54),
.B(n_58),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_45),
.B(n_17),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_44),
.Y(n_58)
);

OAI21xp5_ASAP7_75t_SL g65 ( 
.A1(n_60),
.A2(n_47),
.B(n_24),
.Y(n_65)
);

INVxp67_ASAP7_75t_L g61 ( 
.A(n_43),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_61),
.B(n_42),
.Y(n_62)
);

INVxp67_ASAP7_75t_L g76 ( 
.A(n_62),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_59),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_63),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_65),
.B(n_68),
.Y(n_75)
);

MAJIxp5_ASAP7_75t_L g66 ( 
.A(n_57),
.B(n_26),
.C(n_36),
.Y(n_66)
);

MAJIxp5_ASAP7_75t_L g73 ( 
.A(n_66),
.B(n_70),
.C(n_19),
.Y(n_73)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_56),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_56),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_69),
.B(n_13),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g70 ( 
.A(n_61),
.B(n_26),
.C(n_36),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_66),
.A2(n_60),
.B1(n_52),
.B2(n_24),
.Y(n_72)
);

XNOR2xp5_ASAP7_75t_L g80 ( 
.A(n_73),
.B(n_20),
.Y(n_80)
);

NOR2x1_ASAP7_75t_L g74 ( 
.A(n_64),
.B(n_21),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_74),
.B(n_77),
.Y(n_81)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_70),
.Y(n_78)
);

A2O1A1O1Ixp25_ASAP7_75t_L g79 ( 
.A1(n_72),
.A2(n_67),
.B(n_20),
.C(n_19),
.D(n_15),
.Y(n_79)
);

XOR2xp5_ASAP7_75t_L g85 ( 
.A(n_79),
.B(n_75),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_80),
.B(n_82),
.C(n_83),
.Y(n_84)
);

XNOR2xp5_ASAP7_75t_SL g82 ( 
.A(n_73),
.B(n_20),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_78),
.B(n_2),
.C(n_3),
.Y(n_83)
);

XNOR2xp5_ASAP7_75t_L g88 ( 
.A(n_85),
.B(n_86),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_81),
.B(n_71),
.C(n_76),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_81),
.A2(n_76),
.B1(n_74),
.B2(n_4),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_SL g89 ( 
.A1(n_87),
.A2(n_2),
.B(n_5),
.Y(n_89)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_89),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_85),
.B(n_10),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_90),
.B(n_84),
.C(n_7),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_91),
.B(n_88),
.Y(n_93)
);

OAI21xp5_ASAP7_75t_L g94 ( 
.A1(n_93),
.A2(n_92),
.B(n_1),
.Y(n_94)
);


endmodule