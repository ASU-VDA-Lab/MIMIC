module fake_jpeg_28523_n_68 (n_13, n_21, n_1, n_10, n_23, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_68);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_68;

wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_27;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_40;
wire n_59;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_65;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_62;
wire n_31;
wire n_25;
wire n_56;
wire n_67;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_32;
wire n_66;

INVx1_ASAP7_75t_L g25 ( 
.A(n_22),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_15),
.B(n_6),
.Y(n_26)
);

INVx6_ASAP7_75t_SL g27 ( 
.A(n_14),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_24),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

INVx11_ASAP7_75t_L g30 ( 
.A(n_20),
.Y(n_30)
);

BUFx16f_ASAP7_75t_L g31 ( 
.A(n_23),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_26),
.B(n_0),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_32),
.B(n_35),
.Y(n_45)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_29),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_33),
.B(n_37),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_31),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_34),
.Y(n_39)
);

INVx5_ASAP7_75t_L g35 ( 
.A(n_31),
.Y(n_35)
);

OAI22xp33_ASAP7_75t_SL g36 ( 
.A1(n_28),
.A2(n_9),
.B1(n_19),
.B2(n_18),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_L g42 ( 
.A1(n_36),
.A2(n_28),
.B1(n_30),
.B2(n_25),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_26),
.B(n_29),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_31),
.Y(n_38)
);

FAx1_ASAP7_75t_SL g41 ( 
.A(n_38),
.B(n_27),
.CI(n_30),
.CON(n_41),
.SN(n_41)
);

AO21x2_ASAP7_75t_SL g40 ( 
.A1(n_33),
.A2(n_31),
.B(n_27),
.Y(n_40)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_40),
.Y(n_51)
);

AOI21xp5_ASAP7_75t_L g47 ( 
.A1(n_41),
.A2(n_42),
.B(n_46),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g44 ( 
.A1(n_34),
.A2(n_28),
.B1(n_25),
.B2(n_10),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_L g52 ( 
.A1(n_44),
.A2(n_35),
.B1(n_2),
.B2(n_3),
.Y(n_52)
);

MAJIxp5_ASAP7_75t_L g46 ( 
.A(n_38),
.B(n_17),
.C(n_16),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_45),
.B(n_0),
.Y(n_48)
);

XNOR2xp5_ASAP7_75t_L g57 ( 
.A(n_48),
.B(n_53),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_SL g49 ( 
.A(n_43),
.B(n_41),
.Y(n_49)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_49),
.Y(n_60)
);

INVxp67_ASAP7_75t_L g50 ( 
.A(n_44),
.Y(n_50)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_50),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g56 ( 
.A1(n_52),
.A2(n_54),
.B1(n_40),
.B2(n_3),
.Y(n_56)
);

AOI21xp5_ASAP7_75t_L g53 ( 
.A1(n_41),
.A2(n_1),
.B(n_2),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g54 ( 
.A1(n_40),
.A2(n_21),
.B1(n_13),
.B2(n_12),
.Y(n_54)
);

MAJIxp5_ASAP7_75t_L g55 ( 
.A(n_47),
.B(n_39),
.C(n_46),
.Y(n_55)
);

MAJIxp5_ASAP7_75t_L g63 ( 
.A(n_55),
.B(n_58),
.C(n_1),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_56),
.A2(n_50),
.B1(n_4),
.B2(n_5),
.Y(n_61)
);

XOR2xp5_ASAP7_75t_L g58 ( 
.A(n_51),
.B(n_40),
.Y(n_58)
);

XNOR2xp5_ASAP7_75t_L g65 ( 
.A(n_61),
.B(n_62),
.Y(n_65)
);

OAI221xp5_ASAP7_75t_L g62 ( 
.A1(n_60),
.A2(n_11),
.B1(n_4),
.B2(n_6),
.C(n_7),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_L g64 ( 
.A1(n_63),
.A2(n_57),
.B1(n_55),
.B2(n_59),
.Y(n_64)
);

AOI21xp5_ASAP7_75t_L g66 ( 
.A1(n_64),
.A2(n_58),
.B(n_7),
.Y(n_66)
);

OAI21xp5_ASAP7_75t_L g67 ( 
.A1(n_66),
.A2(n_65),
.B(n_8),
.Y(n_67)
);

XNOR2xp5_ASAP7_75t_L g68 ( 
.A(n_67),
.B(n_8),
.Y(n_68)
);


endmodule