module real_aes_6610_n_103 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_103);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_103;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_555;
wire n_421;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_545;
wire n_556;
wire n_341;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_537;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_564;
wire n_519;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_744;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_178;
wire n_409;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_504;
wire n_455;
wire n_310;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_417;
wire n_363;
wire n_449;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_505;
wire n_434;
wire n_502;
wire n_527;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_552;
wire n_402;
wire n_617;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_735;
wire n_728;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_420;
wire n_336;
wire n_349;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_741;
wire n_283;
wire n_314;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_740;
wire n_371;
wire n_698;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_639;
wire n_587;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
INVx1_ASAP7_75t_L g112 ( .A(n_0), .Y(n_112) );
INVx1_ASAP7_75t_L g536 ( .A(n_1), .Y(n_536) );
INVx1_ASAP7_75t_L g157 ( .A(n_2), .Y(n_157) );
AOI22xp33_ASAP7_75t_L g505 ( .A1(n_3), .A2(n_38), .B1(n_182), .B2(n_482), .Y(n_505) );
AOI21xp33_ASAP7_75t_L g189 ( .A1(n_4), .A2(n_173), .B(n_190), .Y(n_189) );
NAND2xp5_ASAP7_75t_L g548 ( .A(n_5), .B(n_171), .Y(n_548) );
AND2x6_ASAP7_75t_L g150 ( .A(n_6), .B(n_151), .Y(n_150) );
AOI21xp5_ASAP7_75t_L g259 ( .A1(n_7), .A2(n_260), .B(n_261), .Y(n_259) );
NAND2xp5_ASAP7_75t_L g109 ( .A(n_8), .B(n_39), .Y(n_109) );
NOR2xp33_ASAP7_75t_L g124 ( .A(n_8), .B(n_39), .Y(n_124) );
INVx1_ASAP7_75t_L g195 ( .A(n_9), .Y(n_195) );
NAND2xp5_ASAP7_75t_L g251 ( .A(n_10), .B(n_252), .Y(n_251) );
INVx1_ASAP7_75t_L g142 ( .A(n_11), .Y(n_142) );
NAND2xp5_ASAP7_75t_L g491 ( .A(n_12), .B(n_163), .Y(n_491) );
INVx1_ASAP7_75t_L g266 ( .A(n_13), .Y(n_266) );
INVx1_ASAP7_75t_L g530 ( .A(n_14), .Y(n_530) );
NAND2xp5_ASAP7_75t_L g519 ( .A(n_15), .B(n_138), .Y(n_519) );
AO32x2_ASAP7_75t_L g503 ( .A1(n_16), .A2(n_137), .A3(n_171), .B1(n_484), .B2(n_504), .Y(n_503) );
NAND2xp5_ASAP7_75t_SL g494 ( .A(n_17), .B(n_182), .Y(n_494) );
NAND2xp5_ASAP7_75t_L g240 ( .A(n_18), .B(n_178), .Y(n_240) );
NAND2xp5_ASAP7_75t_L g538 ( .A(n_19), .B(n_138), .Y(n_538) );
AOI22xp33_ASAP7_75t_L g507 ( .A1(n_20), .A2(n_50), .B1(n_182), .B2(n_482), .Y(n_507) );
NAND2xp5_ASAP7_75t_SL g223 ( .A(n_21), .B(n_173), .Y(n_223) );
AOI22xp5_ASAP7_75t_L g737 ( .A1(n_22), .A2(n_98), .B1(n_738), .B2(n_739), .Y(n_737) );
INVx1_ASAP7_75t_L g739 ( .A(n_22), .Y(n_739) );
AOI22xp33_ASAP7_75t_SL g483 ( .A1(n_23), .A2(n_76), .B1(n_163), .B2(n_182), .Y(n_483) );
NAND2xp5_ASAP7_75t_SL g473 ( .A(n_24), .B(n_182), .Y(n_473) );
NAND2xp5_ASAP7_75t_L g184 ( .A(n_25), .B(n_185), .Y(n_184) );
A2O1A1Ixp33_ASAP7_75t_L g263 ( .A1(n_26), .A2(n_264), .B(n_265), .C(n_267), .Y(n_263) );
BUFx6f_ASAP7_75t_L g149 ( .A(n_27), .Y(n_149) );
NAND2xp5_ASAP7_75t_L g557 ( .A(n_28), .B(n_168), .Y(n_557) );
NAND2xp5_ASAP7_75t_L g160 ( .A(n_29), .B(n_161), .Y(n_160) );
NAND2xp5_ASAP7_75t_L g444 ( .A(n_30), .B(n_119), .Y(n_444) );
OAI22xp5_ASAP7_75t_SL g127 ( .A1(n_31), .A2(n_88), .B1(n_128), .B2(n_129), .Y(n_127) );
CKINVDCx20_ASAP7_75t_R g128 ( .A(n_31), .Y(n_128) );
INVx1_ASAP7_75t_L g210 ( .A(n_32), .Y(n_210) );
NAND2xp5_ASAP7_75t_L g475 ( .A(n_33), .B(n_168), .Y(n_475) );
INVx2_ASAP7_75t_L g148 ( .A(n_34), .Y(n_148) );
NAND2xp5_ASAP7_75t_SL g552 ( .A(n_35), .B(n_182), .Y(n_552) );
NAND2xp5_ASAP7_75t_L g496 ( .A(n_36), .B(n_168), .Y(n_496) );
A2O1A1Ixp33_ASAP7_75t_L g224 ( .A1(n_37), .A2(n_150), .B(n_153), .C(n_225), .Y(n_224) );
INVx1_ASAP7_75t_L g208 ( .A(n_40), .Y(n_208) );
NAND2xp5_ASAP7_75t_SL g239 ( .A(n_41), .B(n_161), .Y(n_239) );
AOI22xp33_ASAP7_75t_L g103 ( .A1(n_42), .A2(n_104), .B1(n_117), .B2(n_746), .Y(n_103) );
NAND2xp5_ASAP7_75t_SL g543 ( .A(n_43), .B(n_182), .Y(n_543) );
AOI22xp33_ASAP7_75t_L g481 ( .A1(n_44), .A2(n_86), .B1(n_230), .B2(n_482), .Y(n_481) );
NAND2xp5_ASAP7_75t_SL g546 ( .A(n_45), .B(n_182), .Y(n_546) );
NAND2xp5_ASAP7_75t_L g531 ( .A(n_46), .B(n_182), .Y(n_531) );
CKINVDCx16_ASAP7_75t_R g211 ( .A(n_47), .Y(n_211) );
NAND2xp5_ASAP7_75t_L g547 ( .A(n_48), .B(n_535), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g254 ( .A(n_49), .B(n_173), .Y(n_254) );
AOI22xp33_ASAP7_75t_SL g523 ( .A1(n_51), .A2(n_61), .B1(n_163), .B2(n_182), .Y(n_523) );
OAI22xp5_ASAP7_75t_SL g735 ( .A1(n_52), .A2(n_736), .B1(n_737), .B2(n_740), .Y(n_735) );
CKINVDCx20_ASAP7_75t_R g740 ( .A(n_52), .Y(n_740) );
AOI22xp5_ASAP7_75t_L g205 ( .A1(n_53), .A2(n_153), .B1(n_163), .B2(n_206), .Y(n_205) );
CKINVDCx20_ASAP7_75t_R g233 ( .A(n_54), .Y(n_233) );
NAND2xp5_ASAP7_75t_SL g490 ( .A(n_55), .B(n_182), .Y(n_490) );
CKINVDCx16_ASAP7_75t_R g144 ( .A(n_56), .Y(n_144) );
NAND2xp5_ASAP7_75t_SL g556 ( .A(n_57), .B(n_182), .Y(n_556) );
A2O1A1Ixp33_ASAP7_75t_L g192 ( .A1(n_58), .A2(n_181), .B(n_193), .C(n_194), .Y(n_192) );
CKINVDCx20_ASAP7_75t_R g243 ( .A(n_59), .Y(n_243) );
INVx1_ASAP7_75t_L g191 ( .A(n_60), .Y(n_191) );
INVx1_ASAP7_75t_L g151 ( .A(n_62), .Y(n_151) );
NAND2xp5_ASAP7_75t_L g537 ( .A(n_63), .B(n_182), .Y(n_537) );
INVx1_ASAP7_75t_L g141 ( .A(n_64), .Y(n_141) );
CKINVDCx20_ASAP7_75t_R g447 ( .A(n_65), .Y(n_447) );
AO32x2_ASAP7_75t_L g479 ( .A1(n_66), .A2(n_171), .A3(n_246), .B1(n_480), .B2(n_484), .Y(n_479) );
INVx1_ASAP7_75t_L g555 ( .A(n_67), .Y(n_555) );
INVx1_ASAP7_75t_L g470 ( .A(n_68), .Y(n_470) );
AOI22xp33_ASAP7_75t_L g125 ( .A1(n_69), .A2(n_126), .B1(n_442), .B2(n_443), .Y(n_125) );
CKINVDCx20_ASAP7_75t_R g442 ( .A(n_69), .Y(n_442) );
A2O1A1Ixp33_ASAP7_75t_SL g177 ( .A1(n_70), .A2(n_178), .B(n_179), .C(n_181), .Y(n_177) );
INVxp67_ASAP7_75t_L g180 ( .A(n_71), .Y(n_180) );
NAND2xp5_ASAP7_75t_SL g471 ( .A(n_72), .B(n_163), .Y(n_471) );
INVx1_ASAP7_75t_L g116 ( .A(n_73), .Y(n_116) );
CKINVDCx20_ASAP7_75t_R g213 ( .A(n_74), .Y(n_213) );
INVx1_ASAP7_75t_L g236 ( .A(n_75), .Y(n_236) );
A2O1A1Ixp33_ASAP7_75t_L g237 ( .A1(n_77), .A2(n_150), .B(n_153), .C(n_238), .Y(n_237) );
NAND2xp5_ASAP7_75t_L g495 ( .A(n_78), .B(n_482), .Y(n_495) );
NAND2xp5_ASAP7_75t_SL g474 ( .A(n_79), .B(n_163), .Y(n_474) );
NAND2xp5_ASAP7_75t_SL g226 ( .A(n_80), .B(n_158), .Y(n_226) );
INVx2_ASAP7_75t_L g139 ( .A(n_81), .Y(n_139) );
NAND2xp5_ASAP7_75t_L g227 ( .A(n_82), .B(n_178), .Y(n_227) );
NAND2xp5_ASAP7_75t_L g544 ( .A(n_83), .B(n_163), .Y(n_544) );
A2O1A1Ixp33_ASAP7_75t_L g152 ( .A1(n_84), .A2(n_150), .B(n_153), .C(n_156), .Y(n_152) );
INVx2_ASAP7_75t_L g113 ( .A(n_85), .Y(n_113) );
OR2x2_ASAP7_75t_L g121 ( .A(n_85), .B(n_122), .Y(n_121) );
OR2x2_ASAP7_75t_L g453 ( .A(n_85), .B(n_123), .Y(n_453) );
AOI22xp33_ASAP7_75t_L g522 ( .A1(n_87), .A2(n_102), .B1(n_163), .B2(n_164), .Y(n_522) );
CKINVDCx20_ASAP7_75t_R g129 ( .A(n_88), .Y(n_129) );
NAND2xp5_ASAP7_75t_L g196 ( .A(n_89), .B(n_168), .Y(n_196) );
CKINVDCx20_ASAP7_75t_R g166 ( .A(n_90), .Y(n_166) );
A2O1A1Ixp33_ASAP7_75t_L g248 ( .A1(n_91), .A2(n_150), .B(n_153), .C(n_249), .Y(n_248) );
CKINVDCx20_ASAP7_75t_R g256 ( .A(n_92), .Y(n_256) );
INVx1_ASAP7_75t_L g176 ( .A(n_93), .Y(n_176) );
CKINVDCx16_ASAP7_75t_R g262 ( .A(n_94), .Y(n_262) );
NAND2xp5_ASAP7_75t_SL g250 ( .A(n_95), .B(n_158), .Y(n_250) );
NAND2xp5_ASAP7_75t_L g553 ( .A(n_96), .B(n_163), .Y(n_553) );
NAND2xp5_ASAP7_75t_L g268 ( .A(n_97), .B(n_171), .Y(n_268) );
CKINVDCx20_ASAP7_75t_R g738 ( .A(n_98), .Y(n_738) );
NAND2xp5_ASAP7_75t_L g115 ( .A(n_99), .B(n_116), .Y(n_115) );
AOI21xp5_ASAP7_75t_L g172 ( .A1(n_100), .A2(n_173), .B(n_174), .Y(n_172) );
AOI222xp33_ASAP7_75t_L g449 ( .A1(n_101), .A2(n_450), .B1(n_734), .B2(n_735), .C1(n_741), .C2(n_744), .Y(n_449) );
INVx1_ASAP7_75t_SL g104 ( .A(n_105), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_106), .Y(n_105) );
INVx1_ASAP7_75t_SL g746 ( .A(n_106), .Y(n_746) );
CKINVDCx9p33_ASAP7_75t_R g106 ( .A(n_107), .Y(n_106) );
NAND2xp5_ASAP7_75t_L g107 ( .A(n_108), .B(n_110), .Y(n_107) );
CKINVDCx20_ASAP7_75t_R g108 ( .A(n_109), .Y(n_108) );
CKINVDCx14_ASAP7_75t_R g110 ( .A(n_111), .Y(n_110) );
NAND3xp33_ASAP7_75t_SL g111 ( .A(n_112), .B(n_113), .C(n_114), .Y(n_111) );
AND2x2_ASAP7_75t_L g123 ( .A(n_112), .B(n_124), .Y(n_123) );
OR2x2_ASAP7_75t_L g457 ( .A(n_113), .B(n_123), .Y(n_457) );
NOR2x2_ASAP7_75t_L g743 ( .A(n_113), .B(n_122), .Y(n_743) );
INVx1_ASAP7_75t_SL g114 ( .A(n_115), .Y(n_114) );
AO21x1_ASAP7_75t_SL g117 ( .A1(n_118), .A2(n_445), .B(n_448), .Y(n_117) );
OAI21xp5_ASAP7_75t_L g118 ( .A1(n_119), .A2(n_125), .B(n_444), .Y(n_118) );
CKINVDCx20_ASAP7_75t_R g119 ( .A(n_120), .Y(n_119) );
HB1xp67_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
INVx2_ASAP7_75t_L g122 ( .A(n_123), .Y(n_122) );
INVx1_ASAP7_75t_L g443 ( .A(n_126), .Y(n_443) );
XNOR2xp5_ASAP7_75t_L g126 ( .A(n_127), .B(n_130), .Y(n_126) );
INVx1_ASAP7_75t_L g454 ( .A(n_130), .Y(n_454) );
OAI22xp5_ASAP7_75t_SL g744 ( .A1(n_130), .A2(n_455), .B1(n_459), .B2(n_745), .Y(n_744) );
NAND2x1_ASAP7_75t_L g130 ( .A(n_131), .B(n_358), .Y(n_130) );
NOR5xp2_ASAP7_75t_L g131 ( .A(n_132), .B(n_281), .C(n_313), .D(n_328), .E(n_345), .Y(n_131) );
A2O1A1Ixp33_ASAP7_75t_L g132 ( .A1(n_133), .A2(n_197), .B(n_218), .C(n_269), .Y(n_132) );
NAND2xp5_ASAP7_75t_L g133 ( .A(n_134), .B(n_169), .Y(n_133) );
NAND2xp5_ASAP7_75t_L g380 ( .A(n_134), .B(n_381), .Y(n_380) );
NAND2xp5_ASAP7_75t_L g396 ( .A(n_134), .B(n_333), .Y(n_396) );
INVx1_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
NAND2xp5_ASAP7_75t_L g277 ( .A(n_135), .B(n_278), .Y(n_277) );
NAND2xp5_ASAP7_75t_L g282 ( .A(n_135), .B(n_215), .Y(n_282) );
AND2x2_ASAP7_75t_L g323 ( .A(n_135), .B(n_324), .Y(n_323) );
NAND2xp5_ASAP7_75t_L g327 ( .A(n_135), .B(n_292), .Y(n_327) );
OR2x2_ASAP7_75t_L g364 ( .A(n_135), .B(n_203), .Y(n_364) );
INVx3_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
AND2x2_ASAP7_75t_L g202 ( .A(n_136), .B(n_203), .Y(n_202) );
INVx3_ASAP7_75t_L g272 ( .A(n_136), .Y(n_272) );
OR2x2_ASAP7_75t_L g435 ( .A(n_136), .B(n_275), .Y(n_435) );
AO21x2_ASAP7_75t_L g136 ( .A1(n_137), .A2(n_143), .B(n_165), .Y(n_136) );
AO21x2_ASAP7_75t_L g203 ( .A1(n_137), .A2(n_204), .B(n_212), .Y(n_203) );
NOR2xp33_ASAP7_75t_L g212 ( .A(n_137), .B(n_213), .Y(n_212) );
INVx2_ASAP7_75t_L g231 ( .A(n_137), .Y(n_231) );
INVx1_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
BUFx6f_ASAP7_75t_L g171 ( .A(n_138), .Y(n_171) );
AND2x2_ASAP7_75t_L g138 ( .A(n_139), .B(n_140), .Y(n_138) );
AND2x2_ASAP7_75t_SL g168 ( .A(n_139), .B(n_140), .Y(n_168) );
NAND2xp5_ASAP7_75t_L g140 ( .A(n_141), .B(n_142), .Y(n_140) );
OAI21xp5_ASAP7_75t_L g143 ( .A1(n_144), .A2(n_145), .B(n_152), .Y(n_143) );
OAI22xp33_ASAP7_75t_L g204 ( .A1(n_145), .A2(n_183), .B1(n_205), .B2(n_211), .Y(n_204) );
OAI21xp5_ASAP7_75t_L g235 ( .A1(n_145), .A2(n_236), .B(n_237), .Y(n_235) );
NAND2x1p5_ASAP7_75t_L g145 ( .A(n_146), .B(n_150), .Y(n_145) );
AND2x4_ASAP7_75t_L g173 ( .A(n_146), .B(n_150), .Y(n_173) );
AND2x2_ASAP7_75t_L g146 ( .A(n_147), .B(n_149), .Y(n_146) );
INVx1_ASAP7_75t_L g535 ( .A(n_147), .Y(n_535) );
INVx1_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
INVx2_ASAP7_75t_L g154 ( .A(n_148), .Y(n_154) );
INVx1_ASAP7_75t_L g164 ( .A(n_148), .Y(n_164) );
INVx1_ASAP7_75t_L g155 ( .A(n_149), .Y(n_155) );
INVx3_ASAP7_75t_L g159 ( .A(n_149), .Y(n_159) );
BUFx6f_ASAP7_75t_L g161 ( .A(n_149), .Y(n_161) );
INVx1_ASAP7_75t_L g178 ( .A(n_149), .Y(n_178) );
BUFx6f_ASAP7_75t_L g207 ( .A(n_149), .Y(n_207) );
INVx4_ASAP7_75t_SL g183 ( .A(n_150), .Y(n_183) );
OAI21xp5_ASAP7_75t_L g468 ( .A1(n_150), .A2(n_469), .B(n_472), .Y(n_468) );
BUFx3_ASAP7_75t_L g484 ( .A(n_150), .Y(n_484) );
OAI21xp5_ASAP7_75t_L g488 ( .A1(n_150), .A2(n_489), .B(n_493), .Y(n_488) );
OAI21xp5_ASAP7_75t_L g528 ( .A1(n_150), .A2(n_529), .B(n_533), .Y(n_528) );
OAI21xp5_ASAP7_75t_L g541 ( .A1(n_150), .A2(n_542), .B(n_545), .Y(n_541) );
INVx5_ASAP7_75t_L g175 ( .A(n_153), .Y(n_175) );
AND2x6_ASAP7_75t_L g153 ( .A(n_154), .B(n_155), .Y(n_153) );
BUFx6f_ASAP7_75t_L g182 ( .A(n_154), .Y(n_182) );
BUFx3_ASAP7_75t_L g230 ( .A(n_154), .Y(n_230) );
INVx1_ASAP7_75t_L g482 ( .A(n_154), .Y(n_482) );
O2A1O1Ixp33_ASAP7_75t_L g156 ( .A1(n_157), .A2(n_158), .B(n_160), .C(n_162), .Y(n_156) );
O2A1O1Ixp5_ASAP7_75t_SL g469 ( .A1(n_158), .A2(n_181), .B(n_470), .C(n_471), .Y(n_469) );
INVx2_ASAP7_75t_L g506 ( .A(n_158), .Y(n_506) );
AOI21xp5_ASAP7_75t_L g542 ( .A1(n_158), .A2(n_543), .B(n_544), .Y(n_542) );
AOI21xp5_ASAP7_75t_L g551 ( .A1(n_158), .A2(n_552), .B(n_553), .Y(n_551) );
INVx5_ASAP7_75t_L g158 ( .A(n_159), .Y(n_158) );
NOR2xp33_ASAP7_75t_L g179 ( .A(n_159), .B(n_180), .Y(n_179) );
NOR2xp33_ASAP7_75t_L g194 ( .A(n_159), .B(n_195), .Y(n_194) );
OAI22xp5_ASAP7_75t_SL g480 ( .A1(n_159), .A2(n_161), .B1(n_481), .B2(n_483), .Y(n_480) );
INVx2_ASAP7_75t_L g193 ( .A(n_161), .Y(n_193) );
INVx4_ASAP7_75t_L g252 ( .A(n_161), .Y(n_252) );
OAI22xp5_ASAP7_75t_L g504 ( .A1(n_161), .A2(n_505), .B1(n_506), .B2(n_507), .Y(n_504) );
OAI22xp5_ASAP7_75t_L g521 ( .A1(n_161), .A2(n_506), .B1(n_522), .B2(n_523), .Y(n_521) );
O2A1O1Ixp33_ASAP7_75t_L g529 ( .A1(n_162), .A2(n_530), .B(n_531), .C(n_532), .Y(n_529) );
INVx2_ASAP7_75t_L g162 ( .A(n_163), .Y(n_162) );
INVx3_ASAP7_75t_L g163 ( .A(n_164), .Y(n_163) );
NOR2xp33_ASAP7_75t_L g165 ( .A(n_166), .B(n_167), .Y(n_165) );
NOR2xp33_ASAP7_75t_L g242 ( .A(n_167), .B(n_243), .Y(n_242) );
NOR2xp33_ASAP7_75t_L g255 ( .A(n_167), .B(n_256), .Y(n_255) );
INVx1_ASAP7_75t_L g167 ( .A(n_168), .Y(n_167) );
INVx2_ASAP7_75t_L g246 ( .A(n_168), .Y(n_246) );
OA21x2_ASAP7_75t_L g258 ( .A1(n_168), .A2(n_259), .B(n_268), .Y(n_258) );
OA21x2_ASAP7_75t_L g467 ( .A1(n_168), .A2(n_468), .B(n_475), .Y(n_467) );
OA21x2_ASAP7_75t_L g487 ( .A1(n_168), .A2(n_488), .B(n_496), .Y(n_487) );
AOI22xp5_ASAP7_75t_L g337 ( .A1(n_169), .A2(n_338), .B1(n_339), .B2(n_342), .Y(n_337) );
NAND2xp5_ASAP7_75t_L g421 ( .A(n_169), .B(n_272), .Y(n_421) );
AND2x2_ASAP7_75t_L g169 ( .A(n_170), .B(n_187), .Y(n_169) );
AND2x2_ASAP7_75t_L g217 ( .A(n_170), .B(n_203), .Y(n_217) );
AND2x2_ASAP7_75t_L g274 ( .A(n_170), .B(n_275), .Y(n_274) );
INVx1_ASAP7_75t_L g279 ( .A(n_170), .Y(n_279) );
INVx3_ASAP7_75t_L g292 ( .A(n_170), .Y(n_292) );
OR2x2_ASAP7_75t_L g312 ( .A(n_170), .B(n_275), .Y(n_312) );
AND2x2_ASAP7_75t_L g331 ( .A(n_170), .B(n_188), .Y(n_331) );
BUFx2_ASAP7_75t_L g363 ( .A(n_170), .Y(n_363) );
OA21x2_ASAP7_75t_L g170 ( .A1(n_171), .A2(n_172), .B(n_184), .Y(n_170) );
INVx4_ASAP7_75t_L g186 ( .A(n_171), .Y(n_186) );
OA21x2_ASAP7_75t_L g540 ( .A1(n_171), .A2(n_541), .B(n_548), .Y(n_540) );
BUFx2_ASAP7_75t_L g260 ( .A(n_173), .Y(n_260) );
O2A1O1Ixp33_ASAP7_75t_L g174 ( .A1(n_175), .A2(n_176), .B(n_177), .C(n_183), .Y(n_174) );
O2A1O1Ixp33_ASAP7_75t_L g190 ( .A1(n_175), .A2(n_183), .B(n_191), .C(n_192), .Y(n_190) );
O2A1O1Ixp33_ASAP7_75t_L g261 ( .A1(n_175), .A2(n_183), .B(n_262), .C(n_263), .Y(n_261) );
INVx1_ASAP7_75t_L g492 ( .A(n_178), .Y(n_492) );
INVx3_ASAP7_75t_L g181 ( .A(n_182), .Y(n_181) );
HB1xp67_ASAP7_75t_L g253 ( .A(n_182), .Y(n_253) );
OA21x2_ASAP7_75t_L g188 ( .A1(n_185), .A2(n_189), .B(n_196), .Y(n_188) );
INVx3_ASAP7_75t_L g185 ( .A(n_186), .Y(n_185) );
NOR2xp33_ASAP7_75t_SL g232 ( .A(n_186), .B(n_233), .Y(n_232) );
NAND3xp33_ASAP7_75t_L g520 ( .A(n_186), .B(n_484), .C(n_521), .Y(n_520) );
AO21x1_ASAP7_75t_L g610 ( .A1(n_186), .A2(n_521), .B(n_611), .Y(n_610) );
AND2x4_ASAP7_75t_L g278 ( .A(n_187), .B(n_279), .Y(n_278) );
INVx1_ASAP7_75t_SL g187 ( .A(n_188), .Y(n_187) );
BUFx2_ASAP7_75t_L g201 ( .A(n_188), .Y(n_201) );
INVx2_ASAP7_75t_L g216 ( .A(n_188), .Y(n_216) );
OR2x2_ASAP7_75t_L g294 ( .A(n_188), .B(n_275), .Y(n_294) );
AND2x2_ASAP7_75t_L g324 ( .A(n_188), .B(n_203), .Y(n_324) );
AND2x2_ASAP7_75t_L g341 ( .A(n_188), .B(n_272), .Y(n_341) );
AND2x2_ASAP7_75t_L g381 ( .A(n_188), .B(n_292), .Y(n_381) );
AND2x2_ASAP7_75t_SL g417 ( .A(n_188), .B(n_217), .Y(n_417) );
AOI21xp5_ASAP7_75t_L g493 ( .A1(n_193), .A2(n_494), .B(n_495), .Y(n_493) );
O2A1O1Ixp5_ASAP7_75t_L g554 ( .A1(n_193), .A2(n_534), .B(n_555), .C(n_556), .Y(n_554) );
INVx1_ASAP7_75t_L g197 ( .A(n_198), .Y(n_197) );
NAND2xp33_ASAP7_75t_SL g198 ( .A(n_199), .B(n_214), .Y(n_198) );
NAND2xp5_ASAP7_75t_L g199 ( .A(n_200), .B(n_202), .Y(n_199) );
NOR2xp33_ASAP7_75t_L g395 ( .A(n_200), .B(n_396), .Y(n_395) );
INVx1_ASAP7_75t_SL g200 ( .A(n_201), .Y(n_200) );
OAI21xp33_ASAP7_75t_L g355 ( .A1(n_201), .A2(n_217), .B(n_356), .Y(n_355) );
NOR2xp33_ASAP7_75t_L g411 ( .A(n_201), .B(n_203), .Y(n_411) );
AND2x2_ASAP7_75t_L g347 ( .A(n_202), .B(n_348), .Y(n_347) );
INVx3_ASAP7_75t_L g275 ( .A(n_203), .Y(n_275) );
HB1xp67_ASAP7_75t_L g373 ( .A(n_203), .Y(n_373) );
OAI22xp5_ASAP7_75t_SL g206 ( .A1(n_207), .A2(n_208), .B1(n_209), .B2(n_210), .Y(n_206) );
INVx2_ASAP7_75t_L g209 ( .A(n_207), .Y(n_209) );
INVx4_ASAP7_75t_L g264 ( .A(n_207), .Y(n_264) );
NOR2xp33_ASAP7_75t_L g440 ( .A(n_214), .B(n_272), .Y(n_440) );
INVx2_ASAP7_75t_L g214 ( .A(n_215), .Y(n_214) );
AOI22xp33_ASAP7_75t_L g382 ( .A1(n_215), .A2(n_383), .B1(n_384), .B2(n_389), .Y(n_382) );
AND2x2_ASAP7_75t_L g215 ( .A(n_216), .B(n_217), .Y(n_215) );
AND2x2_ASAP7_75t_L g273 ( .A(n_216), .B(n_274), .Y(n_273) );
OR2x2_ASAP7_75t_L g311 ( .A(n_216), .B(n_312), .Y(n_311) );
INVx1_ASAP7_75t_SL g348 ( .A(n_216), .Y(n_348) );
NAND2xp5_ASAP7_75t_L g340 ( .A(n_217), .B(n_341), .Y(n_340) );
INVx1_ASAP7_75t_L g402 ( .A(n_217), .Y(n_402) );
CKINVDCx16_ASAP7_75t_R g218 ( .A(n_219), .Y(n_218) );
AND2x2_ASAP7_75t_L g219 ( .A(n_220), .B(n_244), .Y(n_219) );
INVx4_ASAP7_75t_L g288 ( .A(n_220), .Y(n_288) );
AND2x2_ASAP7_75t_L g366 ( .A(n_220), .B(n_333), .Y(n_366) );
AND2x2_ASAP7_75t_L g220 ( .A(n_221), .B(n_234), .Y(n_220) );
INVx3_ASAP7_75t_L g285 ( .A(n_221), .Y(n_285) );
AND2x2_ASAP7_75t_L g299 ( .A(n_221), .B(n_300), .Y(n_299) );
INVx1_ASAP7_75t_L g303 ( .A(n_221), .Y(n_303) );
INVx2_ASAP7_75t_L g317 ( .A(n_221), .Y(n_317) );
NAND2xp5_ASAP7_75t_L g332 ( .A(n_221), .B(n_333), .Y(n_332) );
AND2x2_ASAP7_75t_L g374 ( .A(n_221), .B(n_369), .Y(n_374) );
AND2x2_ASAP7_75t_L g439 ( .A(n_221), .B(n_409), .Y(n_439) );
OR2x6_ASAP7_75t_L g221 ( .A(n_222), .B(n_232), .Y(n_221) );
AOI21xp5_ASAP7_75t_SL g222 ( .A1(n_223), .A2(n_224), .B(n_231), .Y(n_222) );
AOI21xp5_ASAP7_75t_L g225 ( .A1(n_226), .A2(n_227), .B(n_228), .Y(n_225) );
AOI21xp5_ASAP7_75t_L g238 ( .A1(n_228), .A2(n_239), .B(n_240), .Y(n_238) );
INVx2_ASAP7_75t_L g228 ( .A(n_229), .Y(n_228) );
INVx2_ASAP7_75t_L g229 ( .A(n_230), .Y(n_229) );
INVx1_ASAP7_75t_L g267 ( .A(n_230), .Y(n_267) );
INVx1_ASAP7_75t_L g241 ( .A(n_231), .Y(n_241) );
OA21x2_ASAP7_75t_L g527 ( .A1(n_231), .A2(n_528), .B(n_538), .Y(n_527) );
OA21x2_ASAP7_75t_L g549 ( .A1(n_231), .A2(n_550), .B(n_557), .Y(n_549) );
AND2x2_ASAP7_75t_L g280 ( .A(n_234), .B(n_258), .Y(n_280) );
INVx2_ASAP7_75t_L g300 ( .A(n_234), .Y(n_300) );
AO21x2_ASAP7_75t_L g234 ( .A1(n_235), .A2(n_241), .B(n_242), .Y(n_234) );
INVx1_ASAP7_75t_L g305 ( .A(n_244), .Y(n_305) );
AND2x2_ASAP7_75t_L g351 ( .A(n_244), .B(n_299), .Y(n_351) );
AND2x2_ASAP7_75t_L g244 ( .A(n_245), .B(n_257), .Y(n_244) );
INVx2_ASAP7_75t_L g290 ( .A(n_245), .Y(n_290) );
INVx1_ASAP7_75t_L g298 ( .A(n_245), .Y(n_298) );
AND2x2_ASAP7_75t_L g316 ( .A(n_245), .B(n_317), .Y(n_316) );
NAND2xp5_ASAP7_75t_L g354 ( .A(n_245), .B(n_300), .Y(n_354) );
AO21x2_ASAP7_75t_L g245 ( .A1(n_246), .A2(n_247), .B(n_255), .Y(n_245) );
NAND2xp5_ASAP7_75t_L g247 ( .A(n_248), .B(n_254), .Y(n_247) );
AOI21xp5_ASAP7_75t_L g249 ( .A1(n_250), .A2(n_251), .B(n_253), .Y(n_249) );
AND2x2_ASAP7_75t_L g333 ( .A(n_257), .B(n_290), .Y(n_333) );
INVx1_ASAP7_75t_L g257 ( .A(n_258), .Y(n_257) );
INVx2_ASAP7_75t_L g286 ( .A(n_258), .Y(n_286) );
AND2x2_ASAP7_75t_L g369 ( .A(n_258), .B(n_300), .Y(n_369) );
NOR2xp33_ASAP7_75t_L g265 ( .A(n_264), .B(n_266), .Y(n_265) );
AOI21xp5_ASAP7_75t_L g472 ( .A1(n_264), .A2(n_473), .B(n_474), .Y(n_472) );
INVx1_ASAP7_75t_L g532 ( .A(n_264), .Y(n_532) );
OAI21xp5_ASAP7_75t_SL g269 ( .A1(n_270), .A2(n_276), .B(n_280), .Y(n_269) );
INVx1_ASAP7_75t_SL g314 ( .A(n_270), .Y(n_314) );
AND2x2_ASAP7_75t_L g270 ( .A(n_271), .B(n_273), .Y(n_270) );
NAND2xp5_ASAP7_75t_L g371 ( .A(n_271), .B(n_278), .Y(n_371) );
INVx1_ASAP7_75t_SL g271 ( .A(n_272), .Y(n_271) );
AND2x2_ASAP7_75t_L g320 ( .A(n_272), .B(n_275), .Y(n_320) );
AND2x2_ASAP7_75t_L g349 ( .A(n_272), .B(n_293), .Y(n_349) );
OR2x2_ASAP7_75t_L g352 ( .A(n_272), .B(n_312), .Y(n_352) );
AOI222xp33_ASAP7_75t_L g416 ( .A1(n_273), .A2(n_365), .B1(n_417), .B2(n_418), .C1(n_420), .C2(n_422), .Y(n_416) );
BUFx2_ASAP7_75t_L g330 ( .A(n_275), .Y(n_330) );
INVx1_ASAP7_75t_L g276 ( .A(n_277), .Y(n_276) );
AND2x2_ASAP7_75t_L g319 ( .A(n_278), .B(n_320), .Y(n_319) );
INVx3_ASAP7_75t_SL g336 ( .A(n_278), .Y(n_336) );
NAND2xp5_ASAP7_75t_L g390 ( .A(n_278), .B(n_330), .Y(n_390) );
AND2x2_ASAP7_75t_L g325 ( .A(n_280), .B(n_285), .Y(n_325) );
INVx1_ASAP7_75t_L g344 ( .A(n_280), .Y(n_344) );
OAI221xp5_ASAP7_75t_SL g281 ( .A1(n_282), .A2(n_283), .B1(n_287), .B2(n_291), .C(n_295), .Y(n_281) );
OR2x2_ASAP7_75t_L g353 ( .A(n_283), .B(n_354), .Y(n_353) );
INVx1_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
AND2x2_ASAP7_75t_L g284 ( .A(n_285), .B(n_286), .Y(n_284) );
AND2x2_ASAP7_75t_L g338 ( .A(n_285), .B(n_308), .Y(n_338) );
NAND2xp5_ASAP7_75t_L g378 ( .A(n_285), .B(n_298), .Y(n_378) );
AND2x2_ASAP7_75t_L g383 ( .A(n_285), .B(n_333), .Y(n_383) );
HB1xp67_ASAP7_75t_L g393 ( .A(n_285), .Y(n_393) );
NAND2x1_ASAP7_75t_SL g404 ( .A(n_285), .B(n_405), .Y(n_404) );
OR2x2_ASAP7_75t_L g289 ( .A(n_286), .B(n_290), .Y(n_289) );
INVx2_ASAP7_75t_L g309 ( .A(n_286), .Y(n_309) );
NAND2xp5_ASAP7_75t_L g335 ( .A(n_286), .B(n_304), .Y(n_335) );
INVx1_ASAP7_75t_L g401 ( .A(n_286), .Y(n_401) );
INVx1_ASAP7_75t_L g376 ( .A(n_287), .Y(n_376) );
OR2x2_ASAP7_75t_L g287 ( .A(n_288), .B(n_289), .Y(n_287) );
INVx1_ASAP7_75t_L g388 ( .A(n_288), .Y(n_388) );
NOR2xp67_ASAP7_75t_L g400 ( .A(n_288), .B(n_401), .Y(n_400) );
INVx2_ASAP7_75t_L g405 ( .A(n_289), .Y(n_405) );
NOR2xp33_ASAP7_75t_L g412 ( .A(n_289), .B(n_413), .Y(n_412) );
AND2x2_ASAP7_75t_L g308 ( .A(n_290), .B(n_309), .Y(n_308) );
NAND2xp5_ASAP7_75t_L g321 ( .A(n_290), .B(n_300), .Y(n_321) );
INVx1_ASAP7_75t_L g387 ( .A(n_290), .Y(n_387) );
INVx1_ASAP7_75t_L g408 ( .A(n_291), .Y(n_408) );
NAND2xp5_ASAP7_75t_L g291 ( .A(n_292), .B(n_293), .Y(n_291) );
INVx1_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
OAI21xp5_ASAP7_75t_SL g295 ( .A1(n_296), .A2(n_301), .B(n_310), .Y(n_295) );
AND2x2_ASAP7_75t_L g296 ( .A(n_297), .B(n_299), .Y(n_296) );
AND2x2_ASAP7_75t_L g441 ( .A(n_297), .B(n_374), .Y(n_441) );
INVx1_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
AND2x2_ASAP7_75t_L g409 ( .A(n_298), .B(n_369), .Y(n_409) );
AOI32xp33_ASAP7_75t_L g322 ( .A1(n_299), .A2(n_305), .A3(n_323), .B1(n_325), .B2(n_326), .Y(n_322) );
AOI322xp5_ASAP7_75t_L g424 ( .A1(n_299), .A2(n_331), .A3(n_414), .B1(n_425), .B2(n_426), .C1(n_427), .C2(n_429), .Y(n_424) );
INVx2_ASAP7_75t_L g304 ( .A(n_300), .Y(n_304) );
INVx1_ASAP7_75t_L g414 ( .A(n_300), .Y(n_414) );
OAI22xp5_ASAP7_75t_L g301 ( .A1(n_302), .A2(n_305), .B1(n_306), .B2(n_307), .Y(n_301) );
NAND2xp5_ASAP7_75t_L g357 ( .A(n_302), .B(n_308), .Y(n_357) );
AND2x2_ASAP7_75t_L g302 ( .A(n_303), .B(n_304), .Y(n_302) );
NAND2xp5_ASAP7_75t_L g419 ( .A(n_303), .B(n_369), .Y(n_419) );
INVx1_ASAP7_75t_L g306 ( .A(n_304), .Y(n_306) );
NAND2xp5_ASAP7_75t_L g423 ( .A(n_304), .B(n_333), .Y(n_423) );
INVx1_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
INVx1_ASAP7_75t_SL g310 ( .A(n_311), .Y(n_310) );
NOR2xp33_ASAP7_75t_L g406 ( .A(n_312), .B(n_407), .Y(n_406) );
OAI221xp5_ASAP7_75t_SL g313 ( .A1(n_314), .A2(n_315), .B1(n_318), .B2(n_321), .C(n_322), .Y(n_313) );
OR2x2_ASAP7_75t_L g334 ( .A(n_315), .B(n_335), .Y(n_334) );
OR2x2_ASAP7_75t_L g343 ( .A(n_315), .B(n_344), .Y(n_343) );
INVx1_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
AND2x2_ASAP7_75t_L g368 ( .A(n_316), .B(n_369), .Y(n_368) );
INVx2_ASAP7_75t_L g318 ( .A(n_319), .Y(n_318) );
AND2x2_ASAP7_75t_L g372 ( .A(n_326), .B(n_373), .Y(n_372) );
INVx1_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
OAI221xp5_ASAP7_75t_L g328 ( .A1(n_329), .A2(n_332), .B1(n_334), .B2(n_336), .C(n_337), .Y(n_328) );
NAND2xp5_ASAP7_75t_L g329 ( .A(n_330), .B(n_331), .Y(n_329) );
AOI22xp5_ASAP7_75t_L g360 ( .A1(n_330), .A2(n_361), .B1(n_365), .B2(n_366), .Y(n_360) );
NAND2xp5_ASAP7_75t_L g431 ( .A(n_331), .B(n_432), .Y(n_431) );
INVx1_ASAP7_75t_L g436 ( .A(n_331), .Y(n_436) );
INVx1_ASAP7_75t_L g430 ( .A(n_333), .Y(n_430) );
INVx1_ASAP7_75t_SL g365 ( .A(n_334), .Y(n_365) );
NOR2xp33_ASAP7_75t_L g426 ( .A(n_336), .B(n_364), .Y(n_426) );
INVx1_ASAP7_75t_L g339 ( .A(n_340), .Y(n_339) );
NAND2xp5_ASAP7_75t_L g399 ( .A(n_341), .B(n_400), .Y(n_399) );
INVx1_ASAP7_75t_SL g407 ( .A(n_341), .Y(n_407) );
INVx1_ASAP7_75t_SL g342 ( .A(n_343), .Y(n_342) );
OAI221xp5_ASAP7_75t_SL g345 ( .A1(n_346), .A2(n_350), .B1(n_352), .B2(n_353), .C(n_355), .Y(n_345) );
NOR2xp33_ASAP7_75t_SL g346 ( .A(n_347), .B(n_349), .Y(n_346) );
AOI22xp5_ASAP7_75t_L g410 ( .A1(n_347), .A2(n_365), .B1(n_411), .B2(n_412), .Y(n_410) );
CKINVDCx14_ASAP7_75t_R g350 ( .A(n_351), .Y(n_350) );
OAI21xp33_ASAP7_75t_L g429 ( .A1(n_352), .A2(n_430), .B(n_431), .Y(n_429) );
INVx1_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
NOR3xp33_ASAP7_75t_SL g358 ( .A(n_359), .B(n_391), .C(n_415), .Y(n_358) );
NAND4xp25_ASAP7_75t_L g359 ( .A(n_360), .B(n_367), .C(n_375), .D(n_382), .Y(n_359) );
INVx1_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
OR2x2_ASAP7_75t_L g362 ( .A(n_363), .B(n_364), .Y(n_362) );
INVx1_ASAP7_75t_L g438 ( .A(n_363), .Y(n_438) );
INVx3_ASAP7_75t_SL g432 ( .A(n_364), .Y(n_432) );
OR2x2_ASAP7_75t_L g437 ( .A(n_364), .B(n_438), .Y(n_437) );
AOI22xp5_ASAP7_75t_L g367 ( .A1(n_368), .A2(n_370), .B1(n_372), .B2(n_374), .Y(n_367) );
NAND2xp5_ASAP7_75t_L g428 ( .A(n_369), .B(n_387), .Y(n_428) );
INVxp67_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
OAI21xp5_ASAP7_75t_SL g375 ( .A1(n_376), .A2(n_377), .B(n_379), .Y(n_375) );
INVxp67_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
INVx1_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
INVx1_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
NAND2xp5_ASAP7_75t_L g385 ( .A(n_386), .B(n_388), .Y(n_385) );
INVxp67_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
INVx1_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
OAI211xp5_ASAP7_75t_SL g391 ( .A1(n_392), .A2(n_394), .B(n_397), .C(n_410), .Y(n_391) );
INVx1_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
INVx1_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
INVx1_ASAP7_75t_L g425 ( .A(n_396), .Y(n_425) );
AOI222xp33_ASAP7_75t_L g397 ( .A1(n_398), .A2(n_402), .B1(n_403), .B2(n_406), .C1(n_408), .C2(n_409), .Y(n_397) );
INVxp67_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
INVx1_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
NAND4xp25_ASAP7_75t_SL g434 ( .A(n_407), .B(n_435), .C(n_436), .D(n_437), .Y(n_434) );
INVx1_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
NAND3xp33_ASAP7_75t_SL g415 ( .A(n_416), .B(n_424), .C(n_433), .Y(n_415) );
INVx1_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
INVx1_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
INVx1_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
INVx1_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
AOI22xp33_ASAP7_75t_L g433 ( .A1(n_434), .A2(n_439), .B1(n_440), .B2(n_441), .Y(n_433) );
AOI21xp33_ASAP7_75t_L g448 ( .A1(n_444), .A2(n_445), .B(n_449), .Y(n_448) );
INVx2_ASAP7_75t_SL g445 ( .A(n_446), .Y(n_445) );
INVx2_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
OAI22xp5_ASAP7_75t_L g450 ( .A1(n_451), .A2(n_454), .B1(n_455), .B2(n_458), .Y(n_450) );
INVx2_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
INVx2_ASAP7_75t_L g745 ( .A(n_452), .Y(n_745) );
INVx1_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
INVx2_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
INVx1_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
INVx1_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
OR2x2_ASAP7_75t_L g459 ( .A(n_460), .B(n_655), .Y(n_459) );
NAND3xp33_ASAP7_75t_L g460 ( .A(n_461), .B(n_604), .C(n_646), .Y(n_460) );
AOI211xp5_ASAP7_75t_L g461 ( .A1(n_462), .A2(n_513), .B(n_558), .C(n_580), .Y(n_461) );
OAI211xp5_ASAP7_75t_SL g462 ( .A1(n_463), .A2(n_476), .B(n_497), .C(n_508), .Y(n_462) );
INVxp67_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
NAND2xp5_ASAP7_75t_L g561 ( .A(n_464), .B(n_562), .Y(n_561) );
AND2x2_ASAP7_75t_L g667 ( .A(n_464), .B(n_584), .Y(n_667) );
BUFx2_ASAP7_75t_L g464 ( .A(n_465), .Y(n_464) );
AND2x2_ASAP7_75t_L g569 ( .A(n_465), .B(n_500), .Y(n_569) );
NAND2xp5_ASAP7_75t_L g686 ( .A(n_465), .B(n_487), .Y(n_686) );
INVx1_ASAP7_75t_L g704 ( .A(n_465), .Y(n_704) );
AND2x2_ASAP7_75t_L g713 ( .A(n_465), .B(n_601), .Y(n_713) );
INVx2_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
OR2x2_ASAP7_75t_L g596 ( .A(n_466), .B(n_487), .Y(n_596) );
AND2x2_ASAP7_75t_L g654 ( .A(n_466), .B(n_601), .Y(n_654) );
INVx1_ASAP7_75t_L g698 ( .A(n_466), .Y(n_698) );
INVx2_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
OR2x2_ASAP7_75t_L g575 ( .A(n_467), .B(n_576), .Y(n_575) );
INVx2_ASAP7_75t_L g583 ( .A(n_467), .Y(n_583) );
HB1xp67_ASAP7_75t_L g623 ( .A(n_467), .Y(n_623) );
INVxp67_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
NAND2xp5_ASAP7_75t_L g477 ( .A(n_478), .B(n_485), .Y(n_477) );
AND2x2_ASAP7_75t_L g562 ( .A(n_478), .B(n_563), .Y(n_562) );
INVx2_ASAP7_75t_L g595 ( .A(n_478), .Y(n_595) );
OR2x2_ASAP7_75t_L g721 ( .A(n_478), .B(n_722), .Y(n_721) );
NOR2xp33_ASAP7_75t_L g725 ( .A(n_478), .B(n_487), .Y(n_725) );
BUFx6f_ASAP7_75t_L g478 ( .A(n_479), .Y(n_478) );
INVx1_ASAP7_75t_L g500 ( .A(n_479), .Y(n_500) );
INVx1_ASAP7_75t_L g511 ( .A(n_479), .Y(n_511) );
AND2x2_ASAP7_75t_L g584 ( .A(n_479), .B(n_502), .Y(n_584) );
AND2x2_ASAP7_75t_L g624 ( .A(n_479), .B(n_503), .Y(n_624) );
OAI21xp5_ASAP7_75t_L g550 ( .A1(n_484), .A2(n_551), .B(n_554), .Y(n_550) );
INVxp67_ASAP7_75t_L g666 ( .A(n_485), .Y(n_666) );
AND2x4_ASAP7_75t_L g691 ( .A(n_485), .B(n_584), .Y(n_691) );
BUFx3_ASAP7_75t_L g485 ( .A(n_486), .Y(n_485) );
AND2x2_ASAP7_75t_SL g582 ( .A(n_486), .B(n_583), .Y(n_582) );
INVx1_ASAP7_75t_L g486 ( .A(n_487), .Y(n_486) );
AND2x2_ASAP7_75t_L g501 ( .A(n_487), .B(n_502), .Y(n_501) );
AND2x2_ASAP7_75t_L g570 ( .A(n_487), .B(n_503), .Y(n_570) );
INVx1_ASAP7_75t_L g576 ( .A(n_487), .Y(n_576) );
INVx2_ASAP7_75t_L g602 ( .A(n_487), .Y(n_602) );
AND2x2_ASAP7_75t_L g618 ( .A(n_487), .B(n_619), .Y(n_618) );
AOI21xp5_ASAP7_75t_L g489 ( .A1(n_490), .A2(n_491), .B(n_492), .Y(n_489) );
INVx1_ASAP7_75t_L g497 ( .A(n_498), .Y(n_497) );
NAND2xp5_ASAP7_75t_L g606 ( .A(n_498), .B(n_607), .Y(n_606) );
AND2x2_ASAP7_75t_L g498 ( .A(n_499), .B(n_501), .Y(n_498) );
INVx1_ASAP7_75t_L g499 ( .A(n_500), .Y(n_499) );
BUFx2_ASAP7_75t_L g573 ( .A(n_500), .Y(n_573) );
AND2x2_ASAP7_75t_L g681 ( .A(n_500), .B(n_502), .Y(n_681) );
AND2x2_ASAP7_75t_L g598 ( .A(n_501), .B(n_583), .Y(n_598) );
AND2x2_ASAP7_75t_L g697 ( .A(n_501), .B(n_698), .Y(n_697) );
NOR2xp67_ASAP7_75t_L g619 ( .A(n_502), .B(n_620), .Y(n_619) );
OR2x2_ASAP7_75t_L g722 ( .A(n_502), .B(n_583), .Y(n_722) );
INVx2_ASAP7_75t_L g502 ( .A(n_503), .Y(n_502) );
BUFx2_ASAP7_75t_L g512 ( .A(n_503), .Y(n_512) );
AND2x2_ASAP7_75t_L g601 ( .A(n_503), .B(n_602), .Y(n_601) );
O2A1O1Ixp33_ASAP7_75t_L g533 ( .A1(n_506), .A2(n_534), .B(n_536), .C(n_537), .Y(n_533) );
AOI21xp5_ASAP7_75t_L g545 ( .A1(n_506), .A2(n_546), .B(n_547), .Y(n_545) );
INVx1_ASAP7_75t_L g508 ( .A(n_509), .Y(n_508) );
AND2x2_ASAP7_75t_L g509 ( .A(n_510), .B(n_512), .Y(n_509) );
AND2x2_ASAP7_75t_L g647 ( .A(n_510), .B(n_582), .Y(n_647) );
HB1xp67_ASAP7_75t_L g510 ( .A(n_511), .Y(n_510) );
NAND2xp5_ASAP7_75t_L g632 ( .A(n_511), .B(n_583), .Y(n_632) );
INVx2_ASAP7_75t_L g631 ( .A(n_512), .Y(n_631) );
OAI222xp33_ASAP7_75t_L g635 ( .A1(n_512), .A2(n_575), .B1(n_636), .B2(n_638), .C1(n_639), .C2(n_642), .Y(n_635) );
INVx1_ASAP7_75t_L g513 ( .A(n_514), .Y(n_513) );
NAND2xp5_ASAP7_75t_L g514 ( .A(n_515), .B(n_524), .Y(n_514) );
INVx1_ASAP7_75t_L g515 ( .A(n_516), .Y(n_515) );
INVx1_ASAP7_75t_L g516 ( .A(n_517), .Y(n_516) );
INVx2_ASAP7_75t_L g560 ( .A(n_517), .Y(n_560) );
OR2x2_ASAP7_75t_L g671 ( .A(n_517), .B(n_672), .Y(n_671) );
INVx2_ASAP7_75t_L g517 ( .A(n_518), .Y(n_517) );
INVx3_ASAP7_75t_L g593 ( .A(n_518), .Y(n_593) );
NOR2x1_ASAP7_75t_L g644 ( .A(n_518), .B(n_645), .Y(n_644) );
AND2x2_ASAP7_75t_L g650 ( .A(n_518), .B(n_564), .Y(n_650) );
AND2x4_ASAP7_75t_L g518 ( .A(n_519), .B(n_520), .Y(n_518) );
INVx1_ASAP7_75t_L g611 ( .A(n_519), .Y(n_611) );
AOI22xp5_ASAP7_75t_L g652 ( .A1(n_524), .A2(n_614), .B1(n_653), .B2(n_654), .Y(n_652) );
AND2x2_ASAP7_75t_L g524 ( .A(n_525), .B(n_539), .Y(n_524) );
INVx3_ASAP7_75t_L g586 ( .A(n_525), .Y(n_586) );
OR2x2_ASAP7_75t_L g719 ( .A(n_525), .B(n_595), .Y(n_719) );
INVx2_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
AND2x2_ASAP7_75t_L g592 ( .A(n_526), .B(n_593), .Y(n_592) );
AND2x2_ASAP7_75t_L g608 ( .A(n_526), .B(n_609), .Y(n_608) );
AND2x2_ASAP7_75t_L g616 ( .A(n_526), .B(n_564), .Y(n_616) );
NAND2xp5_ASAP7_75t_L g672 ( .A(n_526), .B(n_540), .Y(n_672) );
INVx2_ASAP7_75t_L g526 ( .A(n_527), .Y(n_526) );
AND2x2_ASAP7_75t_L g563 ( .A(n_527), .B(n_564), .Y(n_563) );
AND2x2_ASAP7_75t_L g567 ( .A(n_527), .B(n_540), .Y(n_567) );
AND2x2_ASAP7_75t_L g643 ( .A(n_527), .B(n_590), .Y(n_643) );
NAND2xp5_ASAP7_75t_L g683 ( .A(n_527), .B(n_549), .Y(n_683) );
INVx2_ASAP7_75t_L g534 ( .A(n_535), .Y(n_534) );
NAND2xp5_ASAP7_75t_L g585 ( .A(n_539), .B(n_586), .Y(n_585) );
AND2x2_ASAP7_75t_L g599 ( .A(n_539), .B(n_560), .Y(n_599) );
AND2x2_ASAP7_75t_L g603 ( .A(n_539), .B(n_593), .Y(n_603) );
AND2x2_ASAP7_75t_L g539 ( .A(n_540), .B(n_549), .Y(n_539) );
INVx3_ASAP7_75t_L g564 ( .A(n_540), .Y(n_564) );
AND2x2_ASAP7_75t_L g589 ( .A(n_540), .B(n_590), .Y(n_589) );
AND2x2_ASAP7_75t_L g724 ( .A(n_540), .B(n_707), .Y(n_724) );
HB1xp67_ASAP7_75t_L g578 ( .A(n_549), .Y(n_578) );
INVx2_ASAP7_75t_L g590 ( .A(n_549), .Y(n_590) );
AND2x2_ASAP7_75t_L g634 ( .A(n_549), .B(n_610), .Y(n_634) );
INVx1_ASAP7_75t_L g677 ( .A(n_549), .Y(n_677) );
OR2x2_ASAP7_75t_L g708 ( .A(n_549), .B(n_610), .Y(n_708) );
AND2x2_ASAP7_75t_L g728 ( .A(n_549), .B(n_564), .Y(n_728) );
OAI21xp5_ASAP7_75t_L g558 ( .A1(n_559), .A2(n_561), .B(n_565), .Y(n_558) );
INVx1_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
AND2x2_ASAP7_75t_L g566 ( .A(n_560), .B(n_567), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g693 ( .A(n_560), .B(n_694), .Y(n_693) );
INVx1_ASAP7_75t_L g685 ( .A(n_562), .Y(n_685) );
INVx2_ASAP7_75t_SL g579 ( .A(n_563), .Y(n_579) );
AND2x2_ASAP7_75t_L g699 ( .A(n_563), .B(n_593), .Y(n_699) );
INVx2_ASAP7_75t_L g645 ( .A(n_564), .Y(n_645) );
NAND2xp5_ASAP7_75t_L g676 ( .A(n_564), .B(n_677), .Y(n_676) );
AOI22xp5_ASAP7_75t_L g565 ( .A1(n_566), .A2(n_568), .B1(n_571), .B2(n_577), .Y(n_565) );
NAND2xp5_ASAP7_75t_L g711 ( .A(n_567), .B(n_712), .Y(n_711) );
INVx1_ASAP7_75t_SL g733 ( .A(n_567), .Y(n_733) );
AND2x2_ASAP7_75t_L g568 ( .A(n_569), .B(n_570), .Y(n_568) );
INVx1_ASAP7_75t_L g658 ( .A(n_569), .Y(n_658) );
NAND2xp5_ASAP7_75t_L g670 ( .A(n_569), .B(n_601), .Y(n_670) );
NOR2xp33_ASAP7_75t_L g657 ( .A(n_570), .B(n_658), .Y(n_657) );
AND2x2_ASAP7_75t_L g674 ( .A(n_570), .B(n_623), .Y(n_674) );
INVx2_ASAP7_75t_L g730 ( .A(n_570), .Y(n_730) );
INVx1_ASAP7_75t_L g571 ( .A(n_572), .Y(n_571) );
NAND2xp5_ASAP7_75t_L g572 ( .A(n_573), .B(n_574), .Y(n_572) );
AND2x2_ASAP7_75t_L g600 ( .A(n_573), .B(n_601), .Y(n_600) );
NAND2xp5_ASAP7_75t_L g651 ( .A(n_573), .B(n_618), .Y(n_651) );
INVx2_ASAP7_75t_L g574 ( .A(n_575), .Y(n_574) );
NOR2xp33_ASAP7_75t_L g653 ( .A(n_575), .B(n_595), .Y(n_653) );
NOR2xp33_ASAP7_75t_L g577 ( .A(n_578), .B(n_579), .Y(n_577) );
INVx1_ASAP7_75t_L g712 ( .A(n_578), .Y(n_712) );
O2A1O1Ixp33_ASAP7_75t_SL g662 ( .A1(n_579), .A2(n_663), .B(n_665), .C(n_668), .Y(n_662) );
OR2x2_ASAP7_75t_L g689 ( .A(n_579), .B(n_593), .Y(n_689) );
OAI221xp5_ASAP7_75t_SL g580 ( .A1(n_581), .A2(n_585), .B1(n_587), .B2(n_594), .C(n_597), .Y(n_580) );
NAND2xp5_ASAP7_75t_SL g581 ( .A(n_582), .B(n_584), .Y(n_581) );
NAND2xp5_ASAP7_75t_L g638 ( .A(n_582), .B(n_631), .Y(n_638) );
AND2x2_ASAP7_75t_L g680 ( .A(n_582), .B(n_681), .Y(n_680) );
INVx2_ASAP7_75t_L g716 ( .A(n_582), .Y(n_716) );
HB1xp67_ASAP7_75t_L g607 ( .A(n_583), .Y(n_607) );
INVx1_ASAP7_75t_L g620 ( .A(n_583), .Y(n_620) );
NOR2xp67_ASAP7_75t_L g640 ( .A(n_586), .B(n_641), .Y(n_640) );
INVxp67_ASAP7_75t_L g694 ( .A(n_586), .Y(n_694) );
NAND2xp5_ASAP7_75t_SL g710 ( .A(n_586), .B(n_634), .Y(n_710) );
INVx2_ASAP7_75t_L g696 ( .A(n_587), .Y(n_696) );
OR2x2_ASAP7_75t_L g587 ( .A(n_588), .B(n_591), .Y(n_587) );
INVx1_ASAP7_75t_L g588 ( .A(n_589), .Y(n_588) );
AND2x2_ASAP7_75t_L g637 ( .A(n_589), .B(n_608), .Y(n_637) );
O2A1O1Ixp33_ASAP7_75t_L g646 ( .A1(n_589), .A2(n_605), .B(n_647), .C(n_648), .Y(n_646) );
AND2x2_ASAP7_75t_L g615 ( .A(n_590), .B(n_610), .Y(n_615) );
INVx1_ASAP7_75t_L g591 ( .A(n_592), .Y(n_591) );
NOR2xp33_ASAP7_75t_L g692 ( .A(n_594), .B(n_693), .Y(n_692) );
OR2x2_ASAP7_75t_L g594 ( .A(n_595), .B(n_596), .Y(n_594) );
OR2x2_ASAP7_75t_L g663 ( .A(n_595), .B(n_664), .Y(n_663) );
AOI22xp5_ASAP7_75t_L g597 ( .A1(n_598), .A2(n_599), .B1(n_600), .B2(n_603), .Y(n_597) );
INVx1_ASAP7_75t_L g717 ( .A(n_599), .Y(n_717) );
INVx1_ASAP7_75t_L g664 ( .A(n_601), .Y(n_664) );
INVx1_ASAP7_75t_L g715 ( .A(n_603), .Y(n_715) );
AOI211xp5_ASAP7_75t_SL g604 ( .A1(n_605), .A2(n_608), .B(n_612), .C(n_635), .Y(n_604) );
INVx1_ASAP7_75t_L g605 ( .A(n_606), .Y(n_605) );
OR2x2_ASAP7_75t_L g627 ( .A(n_607), .B(n_628), .Y(n_627) );
INVx1_ASAP7_75t_L g678 ( .A(n_608), .Y(n_678) );
AND2x2_ASAP7_75t_L g727 ( .A(n_608), .B(n_728), .Y(n_727) );
INVx1_ASAP7_75t_L g609 ( .A(n_610), .Y(n_609) );
OAI21xp33_ASAP7_75t_L g612 ( .A1(n_613), .A2(n_617), .B(n_625), .Y(n_612) );
INVx1_ASAP7_75t_SL g613 ( .A(n_614), .Y(n_613) );
AND2x2_ASAP7_75t_L g614 ( .A(n_615), .B(n_616), .Y(n_614) );
INVx2_ASAP7_75t_L g641 ( .A(n_615), .Y(n_641) );
NAND2xp5_ASAP7_75t_L g660 ( .A(n_615), .B(n_661), .Y(n_660) );
AND2x2_ASAP7_75t_L g633 ( .A(n_616), .B(n_634), .Y(n_633) );
INVx2_ASAP7_75t_L g709 ( .A(n_616), .Y(n_709) );
OAI32xp33_ASAP7_75t_L g720 ( .A1(n_616), .A2(n_668), .A3(n_675), .B1(n_716), .B2(n_721), .Y(n_720) );
NOR2xp33_ASAP7_75t_SL g617 ( .A(n_618), .B(n_621), .Y(n_617) );
INVx1_ASAP7_75t_SL g688 ( .A(n_618), .Y(n_688) );
AND2x2_ASAP7_75t_L g621 ( .A(n_622), .B(n_624), .Y(n_621) );
INVx1_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
INVx1_ASAP7_75t_SL g628 ( .A(n_624), .Y(n_628) );
OAI21xp33_ASAP7_75t_L g625 ( .A1(n_626), .A2(n_629), .B(n_633), .Y(n_625) );
INVx1_ASAP7_75t_L g626 ( .A(n_627), .Y(n_626) );
OAI22xp33_ASAP7_75t_L g700 ( .A1(n_627), .A2(n_675), .B1(n_701), .B2(n_703), .Y(n_700) );
INVx1_ASAP7_75t_L g629 ( .A(n_630), .Y(n_629) );
OR2x2_ASAP7_75t_L g630 ( .A(n_631), .B(n_632), .Y(n_630) );
NAND2xp5_ASAP7_75t_L g703 ( .A(n_631), .B(n_704), .Y(n_703) );
INVx1_ASAP7_75t_L g668 ( .A(n_634), .Y(n_668) );
INVx1_ASAP7_75t_L g636 ( .A(n_637), .Y(n_636) );
INVx1_ASAP7_75t_L g639 ( .A(n_640), .Y(n_639) );
NAND2x1p5_ASAP7_75t_L g642 ( .A(n_643), .B(n_644), .Y(n_642) );
INVx1_ASAP7_75t_L g661 ( .A(n_645), .Y(n_661) );
OAI21xp5_ASAP7_75t_L g648 ( .A1(n_649), .A2(n_651), .B(n_652), .Y(n_648) );
INVx1_ASAP7_75t_L g649 ( .A(n_650), .Y(n_649) );
AOI221xp5_ASAP7_75t_L g695 ( .A1(n_654), .A2(n_696), .B1(n_697), .B2(n_699), .C(n_700), .Y(n_695) );
NAND5xp2_ASAP7_75t_L g655 ( .A(n_656), .B(n_679), .C(n_695), .D(n_705), .E(n_723), .Y(n_655) );
AOI211xp5_ASAP7_75t_SL g656 ( .A1(n_657), .A2(n_659), .B(n_662), .C(n_669), .Y(n_656) );
INVx1_ASAP7_75t_L g659 ( .A(n_660), .Y(n_659) );
INVx1_ASAP7_75t_L g726 ( .A(n_663), .Y(n_726) );
NAND2xp5_ASAP7_75t_L g665 ( .A(n_666), .B(n_667), .Y(n_665) );
OAI22xp33_ASAP7_75t_L g669 ( .A1(n_670), .A2(n_671), .B1(n_673), .B2(n_675), .Y(n_669) );
INVx1_ASAP7_75t_SL g702 ( .A(n_672), .Y(n_702) );
INVx1_ASAP7_75t_L g673 ( .A(n_674), .Y(n_673) );
OAI322xp33_ASAP7_75t_L g684 ( .A1(n_675), .A2(n_685), .A3(n_686), .B1(n_687), .B2(n_688), .C1(n_689), .C2(n_690), .Y(n_684) );
OR2x2_ASAP7_75t_L g675 ( .A(n_676), .B(n_678), .Y(n_675) );
INVx1_ASAP7_75t_L g687 ( .A(n_677), .Y(n_687) );
NAND2xp5_ASAP7_75t_L g701 ( .A(n_677), .B(n_702), .Y(n_701) );
AOI211xp5_ASAP7_75t_SL g679 ( .A1(n_680), .A2(n_682), .B(n_684), .C(n_692), .Y(n_679) );
INVx1_ASAP7_75t_L g682 ( .A(n_683), .Y(n_682) );
OAI22xp33_ASAP7_75t_L g714 ( .A1(n_688), .A2(n_715), .B1(n_716), .B2(n_717), .Y(n_714) );
INVx1_ASAP7_75t_SL g690 ( .A(n_691), .Y(n_690) );
INVx1_ASAP7_75t_L g731 ( .A(n_698), .Y(n_731) );
AOI221xp5_ASAP7_75t_L g705 ( .A1(n_706), .A2(n_713), .B1(n_714), .B2(n_718), .C(n_720), .Y(n_705) );
OAI211xp5_ASAP7_75t_SL g706 ( .A1(n_707), .A2(n_709), .B(n_710), .C(n_711), .Y(n_706) );
INVx1_ASAP7_75t_SL g707 ( .A(n_708), .Y(n_707) );
OR2x2_ASAP7_75t_L g732 ( .A(n_708), .B(n_733), .Y(n_732) );
INVx1_ASAP7_75t_L g718 ( .A(n_719), .Y(n_718) );
AOI221xp5_ASAP7_75t_L g723 ( .A1(n_724), .A2(n_725), .B1(n_726), .B2(n_727), .C(n_729), .Y(n_723) );
AOI21xp33_ASAP7_75t_SL g729 ( .A1(n_730), .A2(n_731), .B(n_732), .Y(n_729) );
CKINVDCx16_ASAP7_75t_R g734 ( .A(n_735), .Y(n_734) );
INVx1_ASAP7_75t_L g736 ( .A(n_737), .Y(n_736) );
INVx1_ASAP7_75t_SL g741 ( .A(n_742), .Y(n_741) );
INVx2_ASAP7_75t_L g742 ( .A(n_743), .Y(n_742) );
endmodule