module fake_jpeg_395_n_234 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_51, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_52, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_234);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_51;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_52;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_234;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_182;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_155;
wire n_207;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_223;
wire n_171;
wire n_119;
wire n_69;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_143;
wire n_202;
wire n_75;
wire n_122;
wire n_233;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_232;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_149;
wire n_157;
wire n_87;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g53 ( 
.A(n_26),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_0),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_14),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_0),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_15),
.Y(n_57)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_45),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_49),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_30),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_28),
.Y(n_61)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_34),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_8),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_17),
.Y(n_64)
);

INVx11_ASAP7_75t_L g65 ( 
.A(n_29),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_13),
.Y(n_66)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_9),
.Y(n_67)
);

INVx5_ASAP7_75t_L g68 ( 
.A(n_32),
.Y(n_68)
);

BUFx12f_ASAP7_75t_L g69 ( 
.A(n_6),
.Y(n_69)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_43),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_16),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_10),
.Y(n_72)
);

BUFx5_ASAP7_75t_L g73 ( 
.A(n_9),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_33),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_42),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_31),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_4),
.Y(n_77)
);

BUFx3_ASAP7_75t_L g78 ( 
.A(n_41),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_20),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_74),
.Y(n_80)
);

INVx8_ASAP7_75t_L g93 ( 
.A(n_80),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_61),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_81),
.B(n_79),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_74),
.Y(n_82)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_82),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_75),
.Y(n_83)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_83),
.Y(n_90)
);

BUFx10_ASAP7_75t_L g84 ( 
.A(n_69),
.Y(n_84)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_84),
.Y(n_98)
);

INVx5_ASAP7_75t_SL g85 ( 
.A(n_57),
.Y(n_85)
);

OR2x2_ASAP7_75t_L g99 ( 
.A(n_85),
.B(n_67),
.Y(n_99)
);

INVx8_ASAP7_75t_L g86 ( 
.A(n_69),
.Y(n_86)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_86),
.Y(n_91)
);

INVx8_ASAP7_75t_L g87 ( 
.A(n_69),
.Y(n_87)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_87),
.Y(n_96)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_58),
.Y(n_88)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_88),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_89),
.B(n_53),
.Y(n_110)
);

A2O1A1Ixp33_ASAP7_75t_L g94 ( 
.A1(n_88),
.A2(n_63),
.B(n_71),
.C(n_56),
.Y(n_94)
);

A2O1A1Ixp33_ASAP7_75t_L g120 ( 
.A1(n_94),
.A2(n_60),
.B(n_84),
.C(n_73),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_80),
.B(n_54),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_95),
.B(n_100),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_82),
.B(n_64),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_97),
.B(n_101),
.Y(n_111)
);

CKINVDCx14_ASAP7_75t_R g105 ( 
.A(n_99),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_83),
.B(n_76),
.Y(n_100)
);

OR2x2_ASAP7_75t_L g101 ( 
.A(n_85),
.B(n_55),
.Y(n_101)
);

INVx5_ASAP7_75t_L g103 ( 
.A(n_93),
.Y(n_103)
);

INVx3_ASAP7_75t_L g131 ( 
.A(n_103),
.Y(n_131)
);

INVx3_ASAP7_75t_SL g104 ( 
.A(n_98),
.Y(n_104)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_104),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_99),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_106),
.B(n_107),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_101),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_94),
.A2(n_66),
.B1(n_57),
.B2(n_72),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_108),
.A2(n_112),
.B1(n_118),
.B2(n_121),
.Y(n_141)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_90),
.Y(n_109)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_109),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_110),
.B(n_68),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_91),
.A2(n_55),
.B1(n_67),
.B2(n_87),
.Y(n_112)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_102),
.Y(n_114)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_114),
.Y(n_137)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_92),
.Y(n_115)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_115),
.Y(n_138)
);

AND2x2_ASAP7_75t_L g116 ( 
.A(n_98),
.B(n_86),
.Y(n_116)
);

XNOR2xp5_ASAP7_75t_L g140 ( 
.A(n_116),
.B(n_119),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_91),
.B(n_59),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_117),
.B(n_120),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_L g118 ( 
.A1(n_90),
.A2(n_77),
.B1(n_66),
.B2(n_72),
.Y(n_118)
);

AND2x2_ASAP7_75t_L g119 ( 
.A(n_96),
.B(n_70),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_102),
.A2(n_77),
.B1(n_75),
.B2(n_78),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_96),
.B(n_78),
.Y(n_122)
);

XNOR2xp5_ASAP7_75t_L g145 ( 
.A(n_122),
.B(n_18),
.Y(n_145)
);

AND2x6_ASAP7_75t_L g123 ( 
.A(n_120),
.B(n_24),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_123),
.B(n_126),
.Y(n_160)
);

NAND2x1_ASAP7_75t_SL g125 ( 
.A(n_105),
.B(n_84),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_L g158 ( 
.A1(n_125),
.A2(n_127),
.B(n_1),
.Y(n_158)
);

NAND2x1_ASAP7_75t_SL g127 ( 
.A(n_111),
.B(n_84),
.Y(n_127)
);

INVx13_ASAP7_75t_L g128 ( 
.A(n_104),
.Y(n_128)
);

CKINVDCx16_ASAP7_75t_R g152 ( 
.A(n_128),
.Y(n_152)
);

AND2x6_ASAP7_75t_L g129 ( 
.A(n_113),
.B(n_22),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_129),
.B(n_132),
.Y(n_161)
);

CKINVDCx12_ASAP7_75t_R g132 ( 
.A(n_116),
.Y(n_132)
);

INVx3_ASAP7_75t_L g133 ( 
.A(n_103),
.Y(n_133)
);

INVx3_ASAP7_75t_SL g157 ( 
.A(n_133),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_SL g136 ( 
.A1(n_112),
.A2(n_65),
.B(n_2),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_L g154 ( 
.A(n_136),
.B(n_145),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_119),
.B(n_93),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_139),
.B(n_142),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_114),
.B(n_62),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_121),
.A2(n_62),
.B1(n_65),
.B2(n_3),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_143),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_167)
);

O2A1O1Ixp33_ASAP7_75t_L g144 ( 
.A1(n_118),
.A2(n_19),
.B(n_51),
.C(n_50),
.Y(n_144)
);

AO21x2_ASAP7_75t_L g163 ( 
.A1(n_144),
.A2(n_48),
.B(n_47),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_L g146 ( 
.A(n_140),
.B(n_124),
.Y(n_146)
);

XOR2xp5_ASAP7_75t_L g188 ( 
.A(n_146),
.B(n_148),
.Y(n_188)
);

INVxp67_ASAP7_75t_L g147 ( 
.A(n_142),
.Y(n_147)
);

INVxp67_ASAP7_75t_L g178 ( 
.A(n_147),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g148 ( 
.A(n_127),
.B(n_52),
.Y(n_148)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_137),
.Y(n_149)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_149),
.Y(n_173)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_138),
.Y(n_150)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_150),
.Y(n_176)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_134),
.Y(n_153)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_153),
.Y(n_179)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_130),
.Y(n_155)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_155),
.Y(n_185)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_139),
.Y(n_156)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_156),
.Y(n_186)
);

CKINVDCx14_ASAP7_75t_R g177 ( 
.A(n_158),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_135),
.B(n_126),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_SL g184 ( 
.A(n_159),
.B(n_162),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_131),
.B(n_1),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_163),
.B(n_27),
.Y(n_190)
);

OAI22xp33_ASAP7_75t_L g164 ( 
.A1(n_141),
.A2(n_36),
.B1(n_44),
.B2(n_40),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_164),
.A2(n_167),
.B1(n_12),
.B2(n_13),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_125),
.B(n_144),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_165),
.B(n_169),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_128),
.B(n_2),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_SL g187 ( 
.A(n_166),
.B(n_46),
.Y(n_187)
);

AOI21xp5_ASAP7_75t_L g168 ( 
.A1(n_135),
.A2(n_5),
.B(n_6),
.Y(n_168)
);

AOI21xp5_ASAP7_75t_L g172 ( 
.A1(n_168),
.A2(n_7),
.B(n_11),
.Y(n_172)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_137),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_124),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g180 ( 
.A(n_170),
.B(n_11),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_147),
.A2(n_7),
.B1(n_8),
.B2(n_10),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_171),
.A2(n_182),
.B1(n_183),
.B2(n_190),
.Y(n_194)
);

INVxp67_ASAP7_75t_L g193 ( 
.A(n_172),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_151),
.B(n_23),
.Y(n_174)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_174),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_180),
.B(n_187),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_146),
.B(n_25),
.Y(n_181)
);

XOR2x2_ASAP7_75t_SL g196 ( 
.A(n_181),
.B(n_148),
.Y(n_196)
);

OAI22x1_ASAP7_75t_L g182 ( 
.A1(n_163),
.A2(n_21),
.B1(n_39),
.B2(n_38),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_SL g189 ( 
.A(n_161),
.B(n_12),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_189),
.B(n_191),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_157),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_L g192 ( 
.A(n_188),
.B(n_154),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_192),
.B(n_196),
.C(n_188),
.Y(n_211)
);

OAI21xp5_ASAP7_75t_SL g199 ( 
.A1(n_175),
.A2(n_160),
.B(n_163),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_199),
.B(n_203),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_184),
.B(n_157),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_200),
.B(n_202),
.Y(n_210)
);

INVx8_ASAP7_75t_L g201 ( 
.A(n_177),
.Y(n_201)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_201),
.Y(n_206)
);

INVxp67_ASAP7_75t_L g202 ( 
.A(n_173),
.Y(n_202)
);

CKINVDCx16_ASAP7_75t_R g203 ( 
.A(n_174),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_186),
.B(n_152),
.Y(n_204)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_204),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_201),
.A2(n_178),
.B1(n_164),
.B2(n_171),
.Y(n_205)
);

BUFx2_ASAP7_75t_L g219 ( 
.A(n_205),
.Y(n_219)
);

HB1xp67_ASAP7_75t_L g207 ( 
.A(n_202),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_207),
.B(n_209),
.Y(n_218)
);

NOR2xp67_ASAP7_75t_SL g208 ( 
.A(n_198),
.B(n_163),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_208),
.B(n_211),
.C(n_213),
.Y(n_215)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_197),
.Y(n_209)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_196),
.B(n_181),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_212),
.B(n_178),
.C(n_193),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_L g224 ( 
.A1(n_216),
.A2(n_217),
.B(n_221),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_213),
.B(n_193),
.C(n_182),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_210),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_220),
.A2(n_207),
.B1(n_194),
.B2(n_185),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_SL g221 ( 
.A(n_214),
.B(n_206),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_222),
.Y(n_227)
);

FAx1_ASAP7_75t_SL g223 ( 
.A(n_215),
.B(n_195),
.CI(n_172),
.CON(n_223),
.SN(n_223)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_223),
.B(n_225),
.Y(n_226)
);

CKINVDCx16_ASAP7_75t_R g225 ( 
.A(n_218),
.Y(n_225)
);

OAI21xp5_ASAP7_75t_SL g228 ( 
.A1(n_226),
.A2(n_224),
.B(n_225),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_228),
.B(n_219),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_229),
.B(n_227),
.Y(n_230)
);

A2O1A1O1Ixp25_ASAP7_75t_L g231 ( 
.A1(n_230),
.A2(n_179),
.B(n_176),
.C(n_183),
.D(n_35),
.Y(n_231)
);

INVxp67_ASAP7_75t_L g232 ( 
.A(n_231),
.Y(n_232)
);

NAND3xp33_ASAP7_75t_L g233 ( 
.A(n_232),
.B(n_37),
.C(n_15),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_233),
.B(n_14),
.Y(n_234)
);


endmodule