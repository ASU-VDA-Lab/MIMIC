module fake_jpeg_21133_n_172 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_172);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_172;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g46 ( 
.A(n_41),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_37),
.Y(n_47)
);

INVx13_ASAP7_75t_L g48 ( 
.A(n_42),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_13),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_10),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_9),
.Y(n_51)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_39),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_33),
.Y(n_53)
);

INVx1_ASAP7_75t_SL g54 ( 
.A(n_5),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_28),
.Y(n_55)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_44),
.Y(n_56)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_8),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_19),
.Y(n_58)
);

HB1xp67_ASAP7_75t_L g59 ( 
.A(n_24),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_11),
.Y(n_60)
);

INVxp33_ASAP7_75t_L g61 ( 
.A(n_31),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_0),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_9),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_21),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_1),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_14),
.Y(n_66)
);

BUFx8_ASAP7_75t_L g67 ( 
.A(n_6),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_26),
.Y(n_68)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_12),
.Y(n_69)
);

BUFx16f_ASAP7_75t_L g70 ( 
.A(n_40),
.Y(n_70)
);

INVx13_ASAP7_75t_L g71 ( 
.A(n_22),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_43),
.Y(n_72)
);

BUFx12f_ASAP7_75t_L g73 ( 
.A(n_7),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_35),
.Y(n_74)
);

INVx8_ASAP7_75t_L g75 ( 
.A(n_17),
.Y(n_75)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_25),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_47),
.Y(n_77)
);

INVx5_ASAP7_75t_L g87 ( 
.A(n_77),
.Y(n_87)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_67),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_78),
.B(n_81),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_61),
.B(n_0),
.Y(n_79)
);

OR2x2_ASAP7_75t_L g85 ( 
.A(n_79),
.B(n_84),
.Y(n_85)
);

BUFx5_ASAP7_75t_L g80 ( 
.A(n_47),
.Y(n_80)
);

AND2x2_ASAP7_75t_SL g89 ( 
.A(n_80),
.B(n_49),
.Y(n_89)
);

BUFx3_ASAP7_75t_L g81 ( 
.A(n_70),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_49),
.Y(n_82)
);

INVx5_ASAP7_75t_L g90 ( 
.A(n_82),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_76),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_83),
.A2(n_54),
.B1(n_51),
.B2(n_65),
.Y(n_94)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_67),
.Y(n_84)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_79),
.Y(n_86)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_86),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_89),
.B(n_74),
.Y(n_101)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_77),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_91),
.B(n_70),
.Y(n_107)
);

BUFx2_ASAP7_75t_R g92 ( 
.A(n_79),
.Y(n_92)
);

OR2x2_ASAP7_75t_L g104 ( 
.A(n_92),
.B(n_95),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_L g93 ( 
.A1(n_77),
.A2(n_56),
.B1(n_61),
.B2(n_57),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_93),
.A2(n_94),
.B1(n_69),
.B2(n_75),
.Y(n_106)
);

HAxp5_ASAP7_75t_SL g95 ( 
.A(n_79),
.B(n_59),
.CON(n_95),
.SN(n_95)
);

BUFx2_ASAP7_75t_L g96 ( 
.A(n_87),
.Y(n_96)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_96),
.Y(n_125)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_87),
.Y(n_97)
);

BUFx2_ASAP7_75t_SL g112 ( 
.A(n_97),
.Y(n_112)
);

CKINVDCx14_ASAP7_75t_R g98 ( 
.A(n_88),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_98),
.B(n_101),
.Y(n_117)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_89),
.Y(n_99)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_99),
.Y(n_109)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_90),
.Y(n_100)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_100),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_85),
.B(n_62),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_102),
.B(n_108),
.Y(n_119)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_90),
.Y(n_103)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_103),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_106),
.A2(n_55),
.B1(n_58),
.B2(n_64),
.Y(n_123)
);

CKINVDCx16_ASAP7_75t_R g116 ( 
.A(n_107),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_85),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_L g110 ( 
.A1(n_103),
.A2(n_93),
.B1(n_95),
.B2(n_52),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_110),
.A2(n_114),
.B1(n_126),
.B2(n_73),
.Y(n_137)
);

INVxp67_ASAP7_75t_L g111 ( 
.A(n_104),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_111),
.B(n_113),
.Y(n_128)
);

INVxp67_ASAP7_75t_L g113 ( 
.A(n_104),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_98),
.A2(n_60),
.B1(n_50),
.B2(n_72),
.Y(n_114)
);

XOR2xp5_ASAP7_75t_L g115 ( 
.A(n_105),
.B(n_59),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_115),
.B(n_121),
.Y(n_134)
);

CKINVDCx16_ASAP7_75t_R g121 ( 
.A(n_96),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_108),
.B(n_46),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_122),
.A2(n_123),
.B1(n_68),
.B2(n_63),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_L g124 ( 
.A(n_102),
.B(n_48),
.Y(n_124)
);

AOI21xp5_ASAP7_75t_L g140 ( 
.A1(n_124),
.A2(n_119),
.B(n_116),
.Y(n_140)
);

AO22x1_ASAP7_75t_SL g126 ( 
.A1(n_108),
.A2(n_74),
.B1(n_71),
.B2(n_66),
.Y(n_126)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_118),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_127),
.B(n_129),
.Y(n_150)
);

INVx5_ASAP7_75t_L g130 ( 
.A(n_112),
.Y(n_130)
);

INVxp67_ASAP7_75t_L g141 ( 
.A(n_130),
.Y(n_141)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_112),
.Y(n_131)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_131),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_117),
.A2(n_53),
.B1(n_63),
.B2(n_73),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_132),
.A2(n_139),
.B1(n_8),
.B2(n_15),
.Y(n_145)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_125),
.Y(n_133)
);

INVxp67_ASAP7_75t_L g146 ( 
.A(n_133),
.Y(n_146)
);

INVx4_ASAP7_75t_L g135 ( 
.A(n_120),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_135),
.Y(n_142)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_126),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_136),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_137),
.A2(n_138),
.B1(n_140),
.B2(n_7),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_109),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_110),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_143),
.B(n_145),
.Y(n_153)
);

AOI21xp5_ASAP7_75t_L g147 ( 
.A1(n_128),
.A2(n_16),
.B(n_18),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_L g151 ( 
.A1(n_147),
.A2(n_29),
.B(n_30),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_134),
.A2(n_20),
.B1(n_23),
.B2(n_27),
.Y(n_149)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_149),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_L g158 ( 
.A(n_151),
.B(n_152),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_L g152 ( 
.A1(n_148),
.A2(n_134),
.B(n_135),
.Y(n_152)
);

XOR2xp5_ASAP7_75t_L g154 ( 
.A(n_150),
.B(n_130),
.Y(n_154)
);

XOR2xp5_ASAP7_75t_L g157 ( 
.A(n_154),
.B(n_142),
.Y(n_157)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_144),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_156),
.Y(n_159)
);

INVxp67_ASAP7_75t_L g160 ( 
.A(n_157),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_160),
.B(n_158),
.C(n_155),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_SL g162 ( 
.A1(n_161),
.A2(n_159),
.B(n_153),
.Y(n_162)
);

CKINVDCx16_ASAP7_75t_R g163 ( 
.A(n_162),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_L g164 ( 
.A(n_163),
.B(n_153),
.Y(n_164)
);

INVxp67_ASAP7_75t_L g165 ( 
.A(n_164),
.Y(n_165)
);

AO21x1_ASAP7_75t_L g166 ( 
.A1(n_165),
.A2(n_141),
.B(n_146),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_SL g167 ( 
.A1(n_166),
.A2(n_141),
.B(n_146),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_167),
.B(n_32),
.C(n_34),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_168),
.B(n_36),
.Y(n_169)
);

BUFx24_ASAP7_75t_SL g170 ( 
.A(n_169),
.Y(n_170)
);

XOR2xp5_ASAP7_75t_L g171 ( 
.A(n_170),
.B(n_38),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_171),
.B(n_45),
.Y(n_172)
);


endmodule