module fake_jpeg_1660_n_541 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_541);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_541;

wire n_529;
wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_349;
wire n_21;
wire n_288;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_511;
wire n_486;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_419;
wire n_378;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_11),
.B(n_8),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_17),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

INVxp67_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_2),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_5),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_1),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_6),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_12),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_2),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_8),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_6),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_9),
.Y(n_38)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_15),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_5),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_12),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_10),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_15),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_3),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_7),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_1),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_7),
.Y(n_47)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_10),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_2),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_13),
.Y(n_50)
);

INVx8_ASAP7_75t_SL g51 ( 
.A(n_7),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_7),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_10),
.Y(n_53)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_11),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_0),
.Y(n_55)
);

BUFx5_ASAP7_75t_L g56 ( 
.A(n_2),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_4),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_22),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_58),
.Y(n_137)
);

INVx11_ASAP7_75t_L g59 ( 
.A(n_33),
.Y(n_59)
);

INVx11_ASAP7_75t_L g132 ( 
.A(n_59),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_22),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g141 ( 
.A(n_60),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_39),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_61),
.B(n_66),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_21),
.B(n_17),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_62),
.B(n_65),
.Y(n_129)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_33),
.Y(n_63)
);

INVx4_ASAP7_75t_SL g169 ( 
.A(n_63),
.Y(n_169)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_29),
.Y(n_64)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_64),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_21),
.B(n_29),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_25),
.Y(n_66)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_22),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g152 ( 
.A(n_67),
.Y(n_152)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_23),
.Y(n_68)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_68),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_37),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g166 ( 
.A(n_69),
.Y(n_166)
);

INVx1_ASAP7_75t_SL g70 ( 
.A(n_51),
.Y(n_70)
);

AND2x2_ASAP7_75t_L g191 ( 
.A(n_70),
.B(n_116),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_20),
.B(n_18),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_71),
.B(n_75),
.Y(n_134)
);

BUFx12f_ASAP7_75t_L g72 ( 
.A(n_54),
.Y(n_72)
);

INVx8_ASAP7_75t_L g172 ( 
.A(n_72),
.Y(n_172)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_25),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_73),
.B(n_77),
.Y(n_145)
);

INVx13_ASAP7_75t_L g74 ( 
.A(n_51),
.Y(n_74)
);

INVx13_ASAP7_75t_L g193 ( 
.A(n_74),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_20),
.B(n_36),
.Y(n_75)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_56),
.Y(n_76)
);

INVx3_ASAP7_75t_L g133 ( 
.A(n_76),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_39),
.Y(n_77)
);

INVx8_ASAP7_75t_L g78 ( 
.A(n_33),
.Y(n_78)
);

INVx5_ASAP7_75t_L g178 ( 
.A(n_78),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_36),
.B(n_57),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_79),
.B(n_110),
.Y(n_138)
);

INVx8_ASAP7_75t_L g80 ( 
.A(n_33),
.Y(n_80)
);

INVx5_ASAP7_75t_L g209 ( 
.A(n_80),
.Y(n_209)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_37),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g167 ( 
.A(n_81),
.Y(n_167)
);

INVx8_ASAP7_75t_L g82 ( 
.A(n_33),
.Y(n_82)
);

BUFx2_ASAP7_75t_L g162 ( 
.A(n_82),
.Y(n_162)
);

BUFx5_ASAP7_75t_L g83 ( 
.A(n_56),
.Y(n_83)
);

INVx4_ASAP7_75t_L g160 ( 
.A(n_83),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_37),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g175 ( 
.A(n_84),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_39),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_85),
.B(n_86),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_19),
.Y(n_86)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_35),
.Y(n_87)
);

INVx3_ASAP7_75t_L g150 ( 
.A(n_87),
.Y(n_150)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_23),
.Y(n_88)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_88),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_19),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_89),
.B(n_94),
.Y(n_151)
);

BUFx12f_ASAP7_75t_L g90 ( 
.A(n_54),
.Y(n_90)
);

INVx8_ASAP7_75t_L g198 ( 
.A(n_90),
.Y(n_198)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_45),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g192 ( 
.A(n_91),
.Y(n_192)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_35),
.Y(n_92)
);

INVx3_ASAP7_75t_L g156 ( 
.A(n_92),
.Y(n_156)
);

BUFx12f_ASAP7_75t_L g93 ( 
.A(n_54),
.Y(n_93)
);

INVx4_ASAP7_75t_L g181 ( 
.A(n_93),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_19),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_45),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g196 ( 
.A(n_95),
.Y(n_196)
);

INVx8_ASAP7_75t_L g96 ( 
.A(n_35),
.Y(n_96)
);

BUFx2_ASAP7_75t_L g170 ( 
.A(n_96),
.Y(n_170)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_48),
.Y(n_97)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_97),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_43),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_98),
.B(n_119),
.Y(n_155)
);

INVx13_ASAP7_75t_L g99 ( 
.A(n_24),
.Y(n_99)
);

CKINVDCx16_ASAP7_75t_R g184 ( 
.A(n_99),
.Y(n_184)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_48),
.Y(n_100)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_100),
.Y(n_189)
);

INVx5_ASAP7_75t_L g101 ( 
.A(n_35),
.Y(n_101)
);

BUFx3_ASAP7_75t_L g157 ( 
.A(n_101),
.Y(n_157)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_35),
.Y(n_102)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_102),
.Y(n_190)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_45),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g208 ( 
.A(n_103),
.Y(n_208)
);

INVx8_ASAP7_75t_L g104 ( 
.A(n_38),
.Y(n_104)
);

BUFx2_ASAP7_75t_L g185 ( 
.A(n_104),
.Y(n_185)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_38),
.Y(n_105)
);

INVx3_ASAP7_75t_L g173 ( 
.A(n_105),
.Y(n_173)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_38),
.Y(n_106)
);

INVx3_ASAP7_75t_L g174 ( 
.A(n_106),
.Y(n_174)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_38),
.Y(n_107)
);

INVx3_ASAP7_75t_L g188 ( 
.A(n_107),
.Y(n_188)
);

BUFx12_ASAP7_75t_L g108 ( 
.A(n_38),
.Y(n_108)
);

BUFx2_ASAP7_75t_L g194 ( 
.A(n_108),
.Y(n_194)
);

BUFx12f_ASAP7_75t_L g109 ( 
.A(n_52),
.Y(n_109)
);

INVx4_ASAP7_75t_L g195 ( 
.A(n_109),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_27),
.B(n_17),
.Y(n_110)
);

BUFx12f_ASAP7_75t_L g111 ( 
.A(n_52),
.Y(n_111)
);

INVx3_ASAP7_75t_L g207 ( 
.A(n_111),
.Y(n_207)
);

BUFx3_ASAP7_75t_L g112 ( 
.A(n_52),
.Y(n_112)
);

INVx6_ASAP7_75t_L g158 ( 
.A(n_112),
.Y(n_158)
);

BUFx3_ASAP7_75t_L g113 ( 
.A(n_55),
.Y(n_113)
);

INVx6_ASAP7_75t_L g177 ( 
.A(n_113),
.Y(n_177)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_44),
.Y(n_114)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_114),
.Y(n_204)
);

INVx4_ASAP7_75t_L g115 ( 
.A(n_44),
.Y(n_115)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_115),
.Y(n_206)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_44),
.Y(n_116)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_44),
.Y(n_117)
);

AND2x2_ASAP7_75t_L g199 ( 
.A(n_117),
.B(n_118),
.Y(n_199)
);

INVx1_ASAP7_75t_SL g118 ( 
.A(n_44),
.Y(n_118)
);

BUFx3_ASAP7_75t_L g119 ( 
.A(n_55),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_43),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_120),
.B(n_125),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_27),
.B(n_18),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_121),
.B(n_122),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_30),
.B(n_18),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_55),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_123),
.Y(n_143)
);

INVx11_ASAP7_75t_L g124 ( 
.A(n_30),
.Y(n_124)
);

AOI21xp33_ASAP7_75t_L g130 ( 
.A1(n_124),
.A2(n_53),
.B(n_49),
.Y(n_130)
);

BUFx3_ASAP7_75t_L g125 ( 
.A(n_43),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_67),
.A2(n_50),
.B1(n_57),
.B2(n_28),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_127),
.A2(n_131),
.B1(n_142),
.B2(n_144),
.Y(n_215)
);

AOI21xp5_ASAP7_75t_L g251 ( 
.A1(n_130),
.A2(n_140),
.B(n_168),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_125),
.A2(n_50),
.B1(n_26),
.B2(n_47),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_L g136 ( 
.A1(n_58),
.A2(n_26),
.B1(n_28),
.B2(n_47),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_136),
.A2(n_139),
.B1(n_154),
.B2(n_163),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_60),
.A2(n_50),
.B1(n_53),
.B2(n_49),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_76),
.A2(n_42),
.B1(n_41),
.B2(n_40),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_SL g218 ( 
.A1(n_140),
.A2(n_159),
.B1(n_168),
.B2(n_197),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_69),
.A2(n_46),
.B1(n_34),
.B2(n_32),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_81),
.A2(n_46),
.B1(n_34),
.B2(n_32),
.Y(n_144)
);

AND2x2_ASAP7_75t_SL g148 ( 
.A(n_118),
.B(n_42),
.Y(n_148)
);

CKINVDCx14_ASAP7_75t_R g253 ( 
.A(n_148),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_84),
.A2(n_41),
.B1(n_40),
.B2(n_31),
.Y(n_154)
);

AOI22xp33_ASAP7_75t_SL g159 ( 
.A1(n_72),
.A2(n_31),
.B1(n_3),
.B2(n_4),
.Y(n_159)
);

AOI22xp33_ASAP7_75t_L g163 ( 
.A1(n_91),
.A2(n_0),
.B1(n_3),
.B2(n_4),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_63),
.B(n_16),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_SL g237 ( 
.A(n_164),
.B(n_165),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_70),
.B(n_16),
.Y(n_165)
);

AOI22xp33_ASAP7_75t_SL g168 ( 
.A1(n_72),
.A2(n_0),
.B1(n_3),
.B2(n_4),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_87),
.B(n_16),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_SL g254 ( 
.A(n_171),
.B(n_176),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_92),
.B(n_15),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_117),
.B(n_14),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_179),
.B(n_184),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_SL g180 ( 
.A(n_115),
.B(n_14),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_180),
.B(n_187),
.Y(n_283)
);

OAI22xp33_ASAP7_75t_SL g182 ( 
.A1(n_95),
.A2(n_13),
.B1(n_6),
.B2(n_8),
.Y(n_182)
);

AOI22xp33_ASAP7_75t_L g242 ( 
.A1(n_182),
.A2(n_183),
.B1(n_141),
.B2(n_175),
.Y(n_242)
);

OAI22xp33_ASAP7_75t_SL g183 ( 
.A1(n_103),
.A2(n_5),
.B1(n_6),
.B2(n_8),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_101),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_186),
.B(n_169),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_90),
.B(n_5),
.Y(n_187)
);

AOI22xp33_ASAP7_75t_SL g197 ( 
.A1(n_90),
.A2(n_93),
.B1(n_59),
.B2(n_111),
.Y(n_197)
);

AOI22xp33_ASAP7_75t_SL g200 ( 
.A1(n_93),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_200)
);

AOI22xp33_ASAP7_75t_SL g244 ( 
.A1(n_200),
.A2(n_203),
.B1(n_205),
.B2(n_210),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_123),
.A2(n_9),
.B1(n_119),
.B2(n_113),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_201),
.A2(n_202),
.B1(n_211),
.B2(n_210),
.Y(n_233)
);

AOI22xp33_ASAP7_75t_L g202 ( 
.A1(n_124),
.A2(n_112),
.B1(n_109),
.B2(n_111),
.Y(n_202)
);

AOI22xp33_ASAP7_75t_SL g203 ( 
.A1(n_109),
.A2(n_96),
.B1(n_78),
.B2(n_80),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_82),
.A2(n_104),
.B1(n_108),
.B2(n_99),
.Y(n_205)
);

AOI22xp33_ASAP7_75t_SL g210 ( 
.A1(n_108),
.A2(n_76),
.B1(n_48),
.B2(n_23),
.Y(n_210)
);

AOI22xp33_ASAP7_75t_SL g211 ( 
.A1(n_74),
.A2(n_76),
.B1(n_48),
.B2(n_23),
.Y(n_211)
);

AOI22xp33_ASAP7_75t_SL g259 ( 
.A1(n_211),
.A2(n_160),
.B1(n_194),
.B2(n_181),
.Y(n_259)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_153),
.Y(n_212)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_212),
.Y(n_285)
);

INVxp67_ASAP7_75t_L g213 ( 
.A(n_191),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_213),
.B(n_222),
.Y(n_291)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_151),
.Y(n_214)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_214),
.Y(n_286)
);

INVx3_ASAP7_75t_L g216 ( 
.A(n_178),
.Y(n_216)
);

INVx3_ASAP7_75t_L g327 ( 
.A(n_216),
.Y(n_327)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_146),
.Y(n_217)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_217),
.Y(n_288)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_152),
.Y(n_219)
);

INVx2_ASAP7_75t_L g312 ( 
.A(n_219),
.Y(n_312)
);

AND2x2_ASAP7_75t_L g221 ( 
.A(n_191),
.B(n_199),
.Y(n_221)
);

CKINVDCx16_ASAP7_75t_R g306 ( 
.A(n_221),
.Y(n_306)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_152),
.Y(n_223)
);

INVx2_ASAP7_75t_L g315 ( 
.A(n_223),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_138),
.B(n_134),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_SL g298 ( 
.A(n_224),
.B(n_238),
.Y(n_298)
);

CKINVDCx16_ASAP7_75t_R g326 ( 
.A(n_225),
.Y(n_326)
);

INVx4_ASAP7_75t_L g226 ( 
.A(n_178),
.Y(n_226)
);

INVx5_ASAP7_75t_L g289 ( 
.A(n_226),
.Y(n_289)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_150),
.Y(n_227)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_227),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_129),
.B(n_149),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_228),
.B(n_236),
.Y(n_299)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_135),
.Y(n_229)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_229),
.Y(n_302)
);

INVx3_ASAP7_75t_SL g230 ( 
.A(n_169),
.Y(n_230)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_230),
.Y(n_319)
);

BUFx2_ASAP7_75t_L g231 ( 
.A(n_172),
.Y(n_231)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_231),
.Y(n_325)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_150),
.Y(n_232)
);

BUFx6f_ASAP7_75t_L g297 ( 
.A(n_232),
.Y(n_297)
);

AOI22xp33_ASAP7_75t_SL g313 ( 
.A1(n_233),
.A2(n_248),
.B1(n_259),
.B2(n_268),
.Y(n_313)
);

INVx6_ASAP7_75t_L g234 ( 
.A(n_137),
.Y(n_234)
);

BUFx6f_ASAP7_75t_L g317 ( 
.A(n_234),
.Y(n_317)
);

INVx3_ASAP7_75t_L g235 ( 
.A(n_209),
.Y(n_235)
);

INVx13_ASAP7_75t_L g329 ( 
.A(n_235),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_145),
.B(n_161),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_148),
.B(n_144),
.Y(n_238)
);

INVx8_ASAP7_75t_L g239 ( 
.A(n_158),
.Y(n_239)
);

INVx13_ASAP7_75t_L g335 ( 
.A(n_239),
.Y(n_335)
);

AND2x2_ASAP7_75t_L g240 ( 
.A(n_148),
.B(n_199),
.Y(n_240)
);

CKINVDCx12_ASAP7_75t_R g300 ( 
.A(n_240),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_201),
.A2(n_139),
.B1(n_154),
.B2(n_143),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_241),
.A2(n_277),
.B1(n_220),
.B2(n_233),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_L g296 ( 
.A1(n_242),
.A2(n_215),
.B1(n_213),
.B2(n_221),
.Y(n_296)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_155),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_243),
.B(n_249),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_128),
.B(n_189),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_SL g301 ( 
.A(n_245),
.B(n_251),
.Y(n_301)
);

INVx6_ASAP7_75t_L g246 ( 
.A(n_137),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_246),
.Y(n_287)
);

INVx4_ASAP7_75t_L g247 ( 
.A(n_209),
.Y(n_247)
);

INVx13_ASAP7_75t_L g321 ( 
.A(n_247),
.Y(n_321)
);

INVx1_ASAP7_75t_SL g248 ( 
.A(n_193),
.Y(n_248)
);

AND2x2_ASAP7_75t_L g249 ( 
.A(n_133),
.B(n_147),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_126),
.B(n_133),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_250),
.B(n_252),
.Y(n_305)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_156),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_190),
.B(n_206),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_SL g311 ( 
.A(n_255),
.B(n_269),
.Y(n_311)
);

OAI21xp5_ASAP7_75t_SL g256 ( 
.A1(n_200),
.A2(n_126),
.B(n_159),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_256),
.B(n_257),
.Y(n_307)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_156),
.Y(n_257)
);

INVx5_ASAP7_75t_L g258 ( 
.A(n_172),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_258),
.Y(n_314)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_173),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_260),
.B(n_261),
.Y(n_308)
);

INVx3_ASAP7_75t_L g261 ( 
.A(n_198),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_162),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_262),
.B(n_263),
.Y(n_309)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_204),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_173),
.B(n_188),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_264),
.B(n_266),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_174),
.B(n_188),
.C(n_194),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_265),
.B(n_276),
.C(n_249),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_174),
.B(n_181),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_162),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_267),
.B(n_270),
.Y(n_323)
);

BUFx6f_ASAP7_75t_L g268 ( 
.A(n_141),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_170),
.B(n_185),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_170),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_185),
.B(n_192),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_271),
.B(n_272),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_157),
.B(n_207),
.Y(n_272)
);

BUFx6f_ASAP7_75t_L g273 ( 
.A(n_166),
.Y(n_273)
);

AOI22xp33_ASAP7_75t_SL g328 ( 
.A1(n_273),
.A2(n_279),
.B1(n_280),
.B2(n_282),
.Y(n_328)
);

AOI21xp5_ASAP7_75t_L g274 ( 
.A1(n_197),
.A2(n_203),
.B(n_160),
.Y(n_274)
);

A2O1A1Ixp33_ASAP7_75t_SL g284 ( 
.A1(n_274),
.A2(n_193),
.B(n_132),
.C(n_196),
.Y(n_284)
);

INVx4_ASAP7_75t_L g275 ( 
.A(n_198),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_275),
.B(n_278),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_207),
.B(n_157),
.C(n_195),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_166),
.A2(n_192),
.B1(n_196),
.B2(n_167),
.Y(n_277)
);

INVx5_ASAP7_75t_L g278 ( 
.A(n_158),
.Y(n_278)
);

INVx5_ASAP7_75t_L g279 ( 
.A(n_177),
.Y(n_279)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_167),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_195),
.B(n_177),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_SL g316 ( 
.A1(n_281),
.A2(n_230),
.B1(n_248),
.B2(n_216),
.Y(n_316)
);

BUFx6f_ASAP7_75t_L g282 ( 
.A(n_175),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_SL g367 ( 
.A1(n_284),
.A2(n_300),
.B1(n_314),
.B2(n_331),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_253),
.B(n_208),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_290),
.B(n_294),
.Y(n_337)
);

FAx1_ASAP7_75t_SL g292 ( 
.A(n_240),
.B(n_132),
.CI(n_208),
.CON(n_292),
.SN(n_292)
);

NOR2xp33_ASAP7_75t_SL g341 ( 
.A(n_292),
.B(n_226),
.Y(n_341)
);

OAI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_251),
.A2(n_215),
.B1(n_218),
.B2(n_244),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_L g338 ( 
.A1(n_293),
.A2(n_296),
.B1(n_303),
.B2(n_310),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_283),
.B(n_254),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_SL g310 ( 
.A1(n_274),
.A2(n_241),
.B1(n_220),
.B2(n_221),
.Y(n_310)
);

OAI21xp5_ASAP7_75t_SL g339 ( 
.A1(n_316),
.A2(n_322),
.B(n_258),
.Y(n_339)
);

AND2x2_ASAP7_75t_L g353 ( 
.A(n_320),
.B(n_324),
.Y(n_353)
);

AOI22xp5_ASAP7_75t_SL g322 ( 
.A1(n_237),
.A2(n_277),
.B1(n_279),
.B2(n_278),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_265),
.B(n_276),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_324),
.B(n_333),
.Y(n_340)
);

OAI22xp5_ASAP7_75t_SL g330 ( 
.A1(n_219),
.A2(n_223),
.B1(n_280),
.B2(n_246),
.Y(n_330)
);

AOI22xp5_ASAP7_75t_L g364 ( 
.A1(n_330),
.A2(n_331),
.B1(n_287),
.B2(n_312),
.Y(n_364)
);

OAI22xp5_ASAP7_75t_SL g331 ( 
.A1(n_234),
.A2(n_282),
.B1(n_273),
.B2(n_268),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_227),
.B(n_252),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_232),
.B(n_257),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_336),
.B(n_235),
.Y(n_346)
);

INVxp67_ASAP7_75t_L g380 ( 
.A(n_339),
.Y(n_380)
);

NOR2xp33_ASAP7_75t_L g407 ( 
.A(n_341),
.B(n_348),
.Y(n_407)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_333),
.Y(n_342)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_342),
.Y(n_386)
);

CKINVDCx16_ASAP7_75t_R g343 ( 
.A(n_318),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_SL g382 ( 
.A(n_343),
.B(n_352),
.Y(n_382)
);

INVx2_ASAP7_75t_L g344 ( 
.A(n_312),
.Y(n_344)
);

INVxp67_ASAP7_75t_L g388 ( 
.A(n_344),
.Y(n_388)
);

INVx5_ASAP7_75t_L g345 ( 
.A(n_317),
.Y(n_345)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_345),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_346),
.B(n_350),
.Y(n_391)
);

OAI22xp5_ASAP7_75t_SL g347 ( 
.A1(n_303),
.A2(n_239),
.B1(n_260),
.B2(n_247),
.Y(n_347)
);

AOI22xp5_ASAP7_75t_L g410 ( 
.A1(n_347),
.A2(n_356),
.B1(n_362),
.B2(n_341),
.Y(n_410)
);

CKINVDCx20_ASAP7_75t_R g348 ( 
.A(n_297),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_L g349 ( 
.A(n_326),
.B(n_261),
.Y(n_349)
);

NAND3xp33_ASAP7_75t_L g385 ( 
.A(n_349),
.B(n_358),
.C(n_359),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_SL g350 ( 
.A(n_298),
.B(n_231),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_298),
.B(n_275),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_351),
.B(n_354),
.Y(n_400)
);

CKINVDCx16_ASAP7_75t_R g352 ( 
.A(n_323),
.Y(n_352)
);

MAJIxp5_ASAP7_75t_L g384 ( 
.A(n_353),
.B(n_334),
.C(n_314),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_311),
.B(n_310),
.Y(n_354)
);

INVxp67_ASAP7_75t_SL g355 ( 
.A(n_319),
.Y(n_355)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_355),
.Y(n_403)
);

OAI22xp5_ASAP7_75t_SL g356 ( 
.A1(n_301),
.A2(n_293),
.B1(n_307),
.B2(n_313),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_311),
.B(n_332),
.Y(n_357)
);

XNOR2xp5_ASAP7_75t_L g401 ( 
.A(n_357),
.B(n_360),
.Y(n_401)
);

NOR2xp33_ASAP7_75t_L g358 ( 
.A(n_326),
.B(n_299),
.Y(n_358)
);

NOR2xp33_ASAP7_75t_L g359 ( 
.A(n_286),
.B(n_288),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_SL g360 ( 
.A(n_294),
.B(n_301),
.Y(n_360)
);

NOR2xp33_ASAP7_75t_L g361 ( 
.A(n_286),
.B(n_288),
.Y(n_361)
);

NOR2xp33_ASAP7_75t_SL g379 ( 
.A(n_361),
.B(n_363),
.Y(n_379)
);

OAI22xp5_ASAP7_75t_SL g362 ( 
.A1(n_296),
.A2(n_322),
.B1(n_306),
.B2(n_290),
.Y(n_362)
);

NOR2xp33_ASAP7_75t_L g363 ( 
.A(n_304),
.B(n_302),
.Y(n_363)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_364),
.Y(n_383)
);

OAI21xp5_ASAP7_75t_SL g365 ( 
.A1(n_305),
.A2(n_316),
.B(n_306),
.Y(n_365)
);

OAI21xp5_ASAP7_75t_L g390 ( 
.A1(n_365),
.A2(n_374),
.B(n_377),
.Y(n_390)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_336),
.Y(n_366)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_366),
.Y(n_394)
);

A2O1A1Ixp33_ASAP7_75t_SL g399 ( 
.A1(n_367),
.A2(n_375),
.B(n_335),
.C(n_329),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_320),
.B(n_308),
.Y(n_368)
);

XNOR2xp5_ASAP7_75t_L g405 ( 
.A(n_368),
.B(n_329),
.Y(n_405)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_285),
.Y(n_369)
);

AND2x2_ASAP7_75t_L g393 ( 
.A(n_369),
.B(n_370),
.Y(n_393)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_285),
.Y(n_370)
);

CKINVDCx16_ASAP7_75t_R g371 ( 
.A(n_309),
.Y(n_371)
);

CKINVDCx20_ASAP7_75t_R g392 ( 
.A(n_371),
.Y(n_392)
);

CKINVDCx20_ASAP7_75t_R g372 ( 
.A(n_297),
.Y(n_372)
);

OAI22xp5_ASAP7_75t_L g398 ( 
.A1(n_372),
.A2(n_373),
.B1(n_376),
.B2(n_289),
.Y(n_398)
);

BUFx2_ASAP7_75t_L g373 ( 
.A(n_319),
.Y(n_373)
);

NOR2xp33_ASAP7_75t_L g374 ( 
.A(n_302),
.B(n_291),
.Y(n_374)
);

OA22x2_ASAP7_75t_L g375 ( 
.A1(n_284),
.A2(n_328),
.B1(n_295),
.B2(n_315),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_315),
.Y(n_376)
);

NOR2xp33_ASAP7_75t_L g377 ( 
.A(n_295),
.B(n_325),
.Y(n_377)
);

OAI22xp5_ASAP7_75t_SL g381 ( 
.A1(n_338),
.A2(n_284),
.B1(n_300),
.B2(n_287),
.Y(n_381)
);

AOI22xp5_ASAP7_75t_L g434 ( 
.A1(n_381),
.A2(n_387),
.B1(n_404),
.B2(n_410),
.Y(n_434)
);

MAJIxp5_ASAP7_75t_L g414 ( 
.A(n_384),
.B(n_389),
.C(n_397),
.Y(n_414)
);

OAI22xp5_ASAP7_75t_SL g387 ( 
.A1(n_338),
.A2(n_284),
.B1(n_292),
.B2(n_317),
.Y(n_387)
);

MAJIxp5_ASAP7_75t_L g389 ( 
.A(n_353),
.B(n_327),
.C(n_325),
.Y(n_389)
);

OAI21xp5_ASAP7_75t_L g395 ( 
.A1(n_354),
.A2(n_284),
.B(n_292),
.Y(n_395)
);

OAI21xp5_ASAP7_75t_L g429 ( 
.A1(n_395),
.A2(n_396),
.B(n_399),
.Y(n_429)
);

OAI21xp5_ASAP7_75t_L g396 ( 
.A1(n_365),
.A2(n_327),
.B(n_297),
.Y(n_396)
);

XOR2xp5_ASAP7_75t_L g397 ( 
.A(n_353),
.B(n_330),
.Y(n_397)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_398),
.Y(n_411)
);

AOI21xp5_ASAP7_75t_L g402 ( 
.A1(n_339),
.A2(n_329),
.B(n_321),
.Y(n_402)
);

AOI21xp5_ASAP7_75t_L g436 ( 
.A1(n_402),
.A2(n_409),
.B(n_375),
.Y(n_436)
);

OAI22xp5_ASAP7_75t_SL g404 ( 
.A1(n_340),
.A2(n_360),
.B1(n_368),
.B2(n_342),
.Y(n_404)
);

XOR2xp5_ASAP7_75t_L g417 ( 
.A(n_405),
.B(n_346),
.Y(n_417)
);

MAJIxp5_ASAP7_75t_L g406 ( 
.A(n_340),
.B(n_321),
.C(n_317),
.Y(n_406)
);

MAJIxp5_ASAP7_75t_L g421 ( 
.A(n_406),
.B(n_373),
.C(n_377),
.Y(n_421)
);

OAI21xp5_ASAP7_75t_L g408 ( 
.A1(n_356),
.A2(n_335),
.B(n_289),
.Y(n_408)
);

INVxp67_ASAP7_75t_L g438 ( 
.A(n_408),
.Y(n_438)
);

AOI21xp5_ASAP7_75t_L g409 ( 
.A1(n_362),
.A2(n_335),
.B(n_349),
.Y(n_409)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_393),
.Y(n_412)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_412),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_391),
.B(n_366),
.Y(n_413)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_413),
.Y(n_441)
);

BUFx12_ASAP7_75t_L g415 ( 
.A(n_388),
.Y(n_415)
);

HB1xp67_ASAP7_75t_L g450 ( 
.A(n_415),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_SL g416 ( 
.A(n_394),
.B(n_351),
.Y(n_416)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_416),
.Y(n_447)
);

XNOR2xp5_ASAP7_75t_SL g440 ( 
.A(n_417),
.B(n_404),
.Y(n_440)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_393),
.Y(n_418)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_418),
.Y(n_449)
);

NAND3xp33_ASAP7_75t_L g419 ( 
.A(n_382),
.B(n_357),
.C(n_374),
.Y(n_419)
);

NOR2xp33_ASAP7_75t_L g459 ( 
.A(n_419),
.B(n_425),
.Y(n_459)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_393),
.Y(n_420)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_420),
.Y(n_451)
);

MAJIxp5_ASAP7_75t_L g448 ( 
.A(n_421),
.B(n_424),
.C(n_389),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_391),
.B(n_350),
.Y(n_422)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_422),
.Y(n_452)
);

NOR2xp33_ASAP7_75t_SL g423 ( 
.A(n_392),
.B(n_358),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_SL g454 ( 
.A(n_423),
.B(n_428),
.Y(n_454)
);

MAJIxp5_ASAP7_75t_L g424 ( 
.A(n_405),
.B(n_337),
.C(n_343),
.Y(n_424)
);

BUFx12f_ASAP7_75t_L g425 ( 
.A(n_399),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_394),
.Y(n_426)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_426),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_386),
.B(n_337),
.Y(n_427)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_427),
.Y(n_453)
);

NOR2xp33_ASAP7_75t_L g428 ( 
.A(n_379),
.B(n_352),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_400),
.B(n_361),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_430),
.B(n_433),
.Y(n_442)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_403),
.Y(n_431)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_431),
.Y(n_460)
);

NOR2xp33_ASAP7_75t_L g432 ( 
.A(n_401),
.B(n_371),
.Y(n_432)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_432),
.Y(n_464)
);

INVx13_ASAP7_75t_L g433 ( 
.A(n_399),
.Y(n_433)
);

AOI22xp5_ASAP7_75t_L g435 ( 
.A1(n_387),
.A2(n_347),
.B1(n_364),
.B2(n_367),
.Y(n_435)
);

OAI22xp5_ASAP7_75t_SL g458 ( 
.A1(n_435),
.A2(n_409),
.B1(n_395),
.B2(n_380),
.Y(n_458)
);

OAI21xp5_ASAP7_75t_L g455 ( 
.A1(n_436),
.A2(n_429),
.B(n_402),
.Y(n_455)
);

NOR2xp33_ASAP7_75t_L g437 ( 
.A(n_401),
.B(n_359),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_L g446 ( 
.A(n_437),
.B(n_439),
.Y(n_446)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_383),
.Y(n_439)
);

XNOR2xp5_ASAP7_75t_L g468 ( 
.A(n_440),
.B(n_457),
.Y(n_468)
);

AOI22xp5_ASAP7_75t_L g443 ( 
.A1(n_434),
.A2(n_408),
.B1(n_410),
.B2(n_381),
.Y(n_443)
);

OAI22xp5_ASAP7_75t_L g475 ( 
.A1(n_443),
.A2(n_444),
.B1(n_436),
.B2(n_435),
.Y(n_475)
);

AOI22xp5_ASAP7_75t_SL g444 ( 
.A1(n_438),
.A2(n_380),
.B1(n_399),
.B2(n_383),
.Y(n_444)
);

MAJIxp5_ASAP7_75t_L g466 ( 
.A(n_448),
.B(n_461),
.C(n_421),
.Y(n_466)
);

AOI21xp5_ASAP7_75t_L g482 ( 
.A1(n_455),
.A2(n_407),
.B(n_433),
.Y(n_482)
);

XNOR2xp5_ASAP7_75t_L g457 ( 
.A(n_424),
.B(n_384),
.Y(n_457)
);

AOI22xp5_ASAP7_75t_L g479 ( 
.A1(n_458),
.A2(n_396),
.B1(n_399),
.B2(n_411),
.Y(n_479)
);

MAJIxp5_ASAP7_75t_L g461 ( 
.A(n_414),
.B(n_397),
.C(n_406),
.Y(n_461)
);

XNOR2xp5_ASAP7_75t_SL g462 ( 
.A(n_417),
.B(n_390),
.Y(n_462)
);

XNOR2xp5_ASAP7_75t_L g474 ( 
.A(n_462),
.B(n_463),
.Y(n_474)
);

XNOR2xp5_ASAP7_75t_L g463 ( 
.A(n_414),
.B(n_390),
.Y(n_463)
);

OAI322xp33_ASAP7_75t_L g465 ( 
.A1(n_464),
.A2(n_385),
.A3(n_423),
.B1(n_446),
.B2(n_427),
.C1(n_462),
.C2(n_454),
.Y(n_465)
);

NOR2xp33_ASAP7_75t_SL g492 ( 
.A(n_465),
.B(n_471),
.Y(n_492)
);

XNOR2xp5_ASAP7_75t_L g485 ( 
.A(n_466),
.B(n_484),
.Y(n_485)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_445),
.Y(n_467)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_467),
.Y(n_486)
);

BUFx2_ASAP7_75t_L g469 ( 
.A(n_450),
.Y(n_469)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_469),
.Y(n_488)
);

AOI21xp5_ASAP7_75t_SL g470 ( 
.A1(n_442),
.A2(n_429),
.B(n_438),
.Y(n_470)
);

AOI21xp5_ASAP7_75t_L g489 ( 
.A1(n_470),
.A2(n_455),
.B(n_459),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_SL g471 ( 
.A(n_463),
.B(n_363),
.Y(n_471)
);

MAJIxp5_ASAP7_75t_L g472 ( 
.A(n_461),
.B(n_412),
.C(n_418),
.Y(n_472)
);

MAJIxp5_ASAP7_75t_L g495 ( 
.A(n_472),
.B(n_478),
.C(n_481),
.Y(n_495)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_460),
.Y(n_473)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_473),
.Y(n_496)
);

AND2x2_ASAP7_75t_L g491 ( 
.A(n_475),
.B(n_482),
.Y(n_491)
);

OAI32xp33_ASAP7_75t_L g476 ( 
.A1(n_442),
.A2(n_439),
.A3(n_413),
.B1(n_400),
.B2(n_430),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_L g487 ( 
.A(n_476),
.B(n_477),
.Y(n_487)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_449),
.Y(n_477)
);

MAJIxp5_ASAP7_75t_L g478 ( 
.A(n_448),
.B(n_420),
.C(n_434),
.Y(n_478)
);

OAI22xp5_ASAP7_75t_SL g493 ( 
.A1(n_479),
.A2(n_444),
.B1(n_425),
.B2(n_433),
.Y(n_493)
);

CKINVDCx20_ASAP7_75t_R g480 ( 
.A(n_446),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_L g498 ( 
.A(n_480),
.B(n_483),
.Y(n_498)
);

MAJIxp5_ASAP7_75t_L g481 ( 
.A(n_457),
.B(n_422),
.C(n_426),
.Y(n_481)
);

OAI22xp5_ASAP7_75t_SL g483 ( 
.A1(n_443),
.A2(n_425),
.B1(n_411),
.B2(n_416),
.Y(n_483)
);

MAJIxp5_ASAP7_75t_L g484 ( 
.A(n_440),
.B(n_431),
.C(n_369),
.Y(n_484)
);

OAI21xp5_ASAP7_75t_L g504 ( 
.A1(n_489),
.A2(n_498),
.B(n_487),
.Y(n_504)
);

XNOR2xp5_ASAP7_75t_L g490 ( 
.A(n_466),
.B(n_458),
.Y(n_490)
);

XNOR2xp5_ASAP7_75t_L g506 ( 
.A(n_490),
.B(n_493),
.Y(n_506)
);

OAI22xp5_ASAP7_75t_SL g494 ( 
.A1(n_479),
.A2(n_441),
.B1(n_453),
.B2(n_452),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_L g508 ( 
.A(n_494),
.B(n_483),
.Y(n_508)
);

NOR2x1_ASAP7_75t_L g497 ( 
.A(n_484),
.B(n_447),
.Y(n_497)
);

NOR3xp33_ASAP7_75t_L g501 ( 
.A(n_497),
.B(n_478),
.C(n_472),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_L g499 ( 
.A(n_476),
.B(n_441),
.Y(n_499)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_499),
.Y(n_507)
);

AOI221xp5_ASAP7_75t_L g500 ( 
.A1(n_497),
.A2(n_451),
.B1(n_453),
.B2(n_481),
.C(n_452),
.Y(n_500)
);

NOR2x1_ASAP7_75t_L g517 ( 
.A(n_500),
.B(n_473),
.Y(n_517)
);

AOI21x1_ASAP7_75t_L g512 ( 
.A1(n_501),
.A2(n_504),
.B(n_498),
.Y(n_512)
);

OAI21xp5_ASAP7_75t_SL g502 ( 
.A1(n_489),
.A2(n_470),
.B(n_482),
.Y(n_502)
);

NOR3xp33_ASAP7_75t_L g520 ( 
.A(n_502),
.B(n_509),
.C(n_511),
.Y(n_520)
);

MAJIxp5_ASAP7_75t_L g503 ( 
.A(n_485),
.B(n_468),
.C(n_474),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_SL g521 ( 
.A(n_503),
.B(n_505),
.Y(n_521)
);

MAJIxp5_ASAP7_75t_L g505 ( 
.A(n_485),
.B(n_495),
.C(n_490),
.Y(n_505)
);

NOR2xp33_ASAP7_75t_L g519 ( 
.A(n_508),
.B(n_510),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_L g509 ( 
.A(n_486),
.B(n_469),
.Y(n_509)
);

XNOR2xp5_ASAP7_75t_L g510 ( 
.A(n_495),
.B(n_468),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_L g511 ( 
.A(n_488),
.B(n_494),
.Y(n_511)
);

O2A1O1Ixp33_ASAP7_75t_L g526 ( 
.A1(n_512),
.A2(n_513),
.B(n_375),
.C(n_415),
.Y(n_526)
);

O2A1O1Ixp33_ASAP7_75t_SL g513 ( 
.A1(n_507),
.A2(n_487),
.B(n_499),
.C(n_491),
.Y(n_513)
);

XOR2xp5_ASAP7_75t_SL g514 ( 
.A(n_502),
.B(n_491),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_L g524 ( 
.A(n_514),
.B(n_516),
.Y(n_524)
);

OAI22xp5_ASAP7_75t_SL g515 ( 
.A1(n_504),
.A2(n_491),
.B1(n_492),
.B2(n_496),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_SL g528 ( 
.A(n_515),
.B(n_518),
.Y(n_528)
);

MAJIxp5_ASAP7_75t_L g516 ( 
.A(n_505),
.B(n_474),
.C(n_493),
.Y(n_516)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_517),
.Y(n_529)
);

MAJIxp5_ASAP7_75t_L g518 ( 
.A(n_506),
.B(n_378),
.C(n_388),
.Y(n_518)
);

OAI21x1_ASAP7_75t_L g522 ( 
.A1(n_517),
.A2(n_506),
.B(n_456),
.Y(n_522)
);

AOI21xp5_ASAP7_75t_L g530 ( 
.A1(n_522),
.A2(n_525),
.B(n_526),
.Y(n_530)
);

MAJIxp5_ASAP7_75t_L g523 ( 
.A(n_521),
.B(n_510),
.C(n_503),
.Y(n_523)
);

MAJIxp5_ASAP7_75t_L g534 ( 
.A(n_523),
.B(n_527),
.C(n_522),
.Y(n_534)
);

AOI21xp5_ASAP7_75t_SL g525 ( 
.A1(n_519),
.A2(n_425),
.B(n_370),
.Y(n_525)
);

MAJIxp5_ASAP7_75t_L g527 ( 
.A(n_516),
.B(n_378),
.C(n_348),
.Y(n_527)
);

INVxp67_ASAP7_75t_L g531 ( 
.A(n_524),
.Y(n_531)
);

NOR2xp33_ASAP7_75t_L g537 ( 
.A(n_531),
.B(n_534),
.Y(n_537)
);

OAI21xp5_ASAP7_75t_SL g532 ( 
.A1(n_528),
.A2(n_520),
.B(n_514),
.Y(n_532)
);

AOI21xp5_ASAP7_75t_L g535 ( 
.A1(n_532),
.A2(n_533),
.B(n_530),
.Y(n_535)
);

AOI21xp5_ASAP7_75t_L g533 ( 
.A1(n_529),
.A2(n_518),
.B(n_513),
.Y(n_533)
);

MAJIxp5_ASAP7_75t_L g539 ( 
.A(n_535),
.B(n_536),
.C(n_372),
.Y(n_539)
);

INVxp67_ASAP7_75t_L g536 ( 
.A(n_534),
.Y(n_536)
);

BUFx24_ASAP7_75t_SL g538 ( 
.A(n_537),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_L g540 ( 
.A(n_538),
.B(n_539),
.Y(n_540)
);

XNOR2xp5_ASAP7_75t_L g541 ( 
.A(n_540),
.B(n_415),
.Y(n_541)
);


endmodule