module real_aes_15592_n_103 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_103);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_103;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_887;
wire n_187;
wire n_436;
wire n_599;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_830;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_800;
wire n_778;
wire n_522;
wire n_838;
wire n_485;
wire n_822;
wire n_846;
wire n_222;
wire n_750;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_254;
wire n_207;
wire n_878;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_841;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_421;
wire n_555;
wire n_364;
wire n_329;
wire n_766;
wire n_852;
wire n_132;
wire n_857;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_865;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_884;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_886;
wire n_594;
wire n_856;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_889;
wire n_704;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_870;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_564;
wire n_519;
wire n_815;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_883;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_578;
wire n_528;
wire n_372;
wire n_202;
wire n_892;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_824;
wire n_467;
wire n_875;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_559;
wire n_466;
wire n_636;
wire n_872;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_840;
wire n_570;
wire n_675;
wire n_530;
wire n_835;
wire n_104;
wire n_535;
wire n_732;
wire n_834;
wire n_882;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_755;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_746;
wire n_178;
wire n_409;
wire n_860;
wire n_781;
wire n_748;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_874;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_812;
wire n_817;
wire n_443;
wire n_565;
wire n_782;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_885;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_722;
wire n_745;
wire n_867;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_879;
wire n_331;
wire n_182;
wire n_449;
wire n_363;
wire n_417;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_876;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_527;
wire n_502;
wire n_434;
wire n_505;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_733;
wire n_402;
wire n_552;
wire n_617;
wire n_602;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_880;
wire n_807;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_832;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_859;
wire n_695;
wire n_685;
wire n_881;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_869;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_848;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_188;
wire n_891;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_853;
wire n_810;
wire n_843;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_649;
wire n_193;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_397;
wire n_749;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_851;
wire n_133;
wire n_494;
wire n_711;
wire n_864;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_845;
wire n_850;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_847;
wire n_779;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_765;
wire n_826;
wire n_159;
wire n_108;
wire n_648;
wire n_373;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_831;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_827;
wire n_809;
wire n_482;
wire n_633;
wire n_520;
wire n_679;
wire n_149;
wire n_472;
wire n_866;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_858;
wire n_873;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_753;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_456;
wire n_359;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_861;
wire n_705;
wire n_180;
wire n_212;
wire n_575;
wire n_210;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_541;
wire n_224;
wire n_839;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_863;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_836;
wire n_888;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_890;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_837;
wire n_871;
wire n_474;
wire n_829;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_844;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_601;
wire n_307;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_854;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_877;
wire n_802;
wire n_868;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_842;
wire n_259;
wire n_143;
wire n_849;
wire n_192;
wire n_554;
wire n_475;
wire n_264;
wire n_855;
wire n_798;
wire n_237;
wire n_668;
wire n_797;
wire n_862;
AND2x4_ASAP7_75t_L g104 ( .A(n_0), .B(n_105), .Y(n_104) );
AOI22xp33_ASAP7_75t_L g646 ( .A1(n_1), .A2(n_34), .B1(n_127), .B2(n_177), .Y(n_646) );
AOI22xp5_ASAP7_75t_L g526 ( .A1(n_2), .A2(n_94), .B1(n_527), .B2(n_528), .Y(n_526) );
INVx1_ASAP7_75t_L g527 ( .A(n_2), .Y(n_527) );
OAI22xp5_ASAP7_75t_L g524 ( .A1(n_3), .A2(n_525), .B1(n_526), .B2(n_529), .Y(n_524) );
CKINVDCx5p33_ASAP7_75t_R g529 ( .A(n_3), .Y(n_529) );
AOI22xp5_ASAP7_75t_L g587 ( .A1(n_4), .A2(n_11), .B1(n_554), .B2(n_588), .Y(n_587) );
INVx1_ASAP7_75t_L g105 ( .A(n_5), .Y(n_105) );
CKINVDCx5p33_ASAP7_75t_R g600 ( .A(n_6), .Y(n_600) );
AOI22xp5_ASAP7_75t_L g573 ( .A1(n_7), .A2(n_12), .B1(n_574), .B2(n_575), .Y(n_573) );
OR2x2_ASAP7_75t_L g512 ( .A(n_8), .B(n_30), .Y(n_512) );
BUFx6f_ASAP7_75t_L g128 ( .A(n_9), .Y(n_128) );
CKINVDCx5p33_ASAP7_75t_R g591 ( .A(n_10), .Y(n_591) );
NAND2xp5_ASAP7_75t_SL g141 ( .A(n_13), .B(n_142), .Y(n_141) );
AOI22xp5_ASAP7_75t_L g553 ( .A1(n_14), .A2(n_100), .B1(n_221), .B2(n_554), .Y(n_553) );
AOI22xp33_ASAP7_75t_L g584 ( .A1(n_15), .A2(n_31), .B1(n_585), .B2(n_586), .Y(n_584) );
NAND2xp5_ASAP7_75t_SL g601 ( .A(n_16), .B(n_142), .Y(n_601) );
OAI21x1_ASAP7_75t_L g122 ( .A1(n_17), .A2(n_47), .B(n_123), .Y(n_122) );
NAND2xp5_ASAP7_75t_L g235 ( .A(n_18), .B(n_236), .Y(n_235) );
AOI22xp33_ASAP7_75t_L g882 ( .A1(n_19), .A2(n_58), .B1(n_883), .B2(n_887), .Y(n_882) );
CKINVDCx5p33_ASAP7_75t_R g559 ( .A(n_20), .Y(n_559) );
AOI22xp33_ASAP7_75t_L g647 ( .A1(n_21), .A2(n_38), .B1(n_197), .B2(n_226), .Y(n_647) );
CKINVDCx5p33_ASAP7_75t_R g191 ( .A(n_22), .Y(n_191) );
AOI22xp33_ASAP7_75t_L g564 ( .A1(n_23), .A2(n_44), .B1(n_197), .B2(n_554), .Y(n_564) );
CKINVDCx5p33_ASAP7_75t_R g633 ( .A(n_24), .Y(n_633) );
NAND2xp5_ASAP7_75t_L g603 ( .A(n_25), .B(n_585), .Y(n_603) );
NAND2xp5_ASAP7_75t_SL g234 ( .A(n_26), .B(n_171), .Y(n_234) );
CKINVDCx5p33_ASAP7_75t_R g613 ( .A(n_27), .Y(n_613) );
NAND2xp5_ASAP7_75t_L g119 ( .A(n_28), .B(n_120), .Y(n_119) );
CKINVDCx5p33_ASAP7_75t_R g220 ( .A(n_29), .Y(n_220) );
AOI22xp5_ASAP7_75t_L g628 ( .A1(n_32), .A2(n_84), .B1(n_127), .B2(n_629), .Y(n_628) );
AOI22xp33_ASAP7_75t_L g576 ( .A1(n_33), .A2(n_37), .B1(n_127), .B2(n_577), .Y(n_576) );
AOI22xp33_ASAP7_75t_L g555 ( .A1(n_35), .A2(n_51), .B1(n_554), .B2(n_556), .Y(n_555) );
CKINVDCx5p33_ASAP7_75t_R g196 ( .A(n_36), .Y(n_196) );
CKINVDCx20_ASAP7_75t_R g521 ( .A(n_39), .Y(n_521) );
NAND2xp5_ASAP7_75t_SL g210 ( .A(n_40), .B(n_142), .Y(n_210) );
INVx2_ASAP7_75t_L g505 ( .A(n_41), .Y(n_505) );
NAND2xp5_ASAP7_75t_L g231 ( .A(n_42), .B(n_214), .Y(n_231) );
INVx1_ASAP7_75t_L g510 ( .A(n_43), .Y(n_510) );
BUFx3_ASAP7_75t_L g877 ( .A(n_43), .Y(n_877) );
OAI22x1_ASAP7_75t_SL g495 ( .A1(n_45), .A2(n_496), .B1(n_497), .B2(n_500), .Y(n_495) );
CKINVDCx5p33_ASAP7_75t_R g500 ( .A(n_45), .Y(n_500) );
NAND2xp5_ASAP7_75t_L g238 ( .A(n_46), .B(n_160), .Y(n_238) );
AND2x2_ASAP7_75t_L g199 ( .A(n_48), .B(n_160), .Y(n_199) );
NAND2xp5_ASAP7_75t_L g156 ( .A(n_49), .B(n_157), .Y(n_156) );
OAI22xp5_ASAP7_75t_L g497 ( .A1(n_50), .A2(n_80), .B1(n_498), .B2(n_499), .Y(n_497) );
INVxp67_ASAP7_75t_L g498 ( .A(n_50), .Y(n_498) );
NAND2xp5_ASAP7_75t_SL g170 ( .A(n_52), .B(n_171), .Y(n_170) );
NAND2xp5_ASAP7_75t_L g225 ( .A(n_53), .B(n_226), .Y(n_225) );
AOI22xp33_ASAP7_75t_L g563 ( .A1(n_54), .A2(n_71), .B1(n_226), .B2(n_556), .Y(n_563) );
AOI22xp33_ASAP7_75t_L g611 ( .A1(n_55), .A2(n_74), .B1(n_127), .B2(n_577), .Y(n_611) );
NAND2xp5_ASAP7_75t_L g175 ( .A(n_56), .B(n_176), .Y(n_175) );
A2O1A1Ixp33_ASAP7_75t_L g189 ( .A1(n_57), .A2(n_131), .B(n_140), .C(n_190), .Y(n_189) );
AOI22xp5_ASAP7_75t_L g107 ( .A1(n_58), .A2(n_108), .B1(n_501), .B2(n_502), .Y(n_107) );
INVx1_ASAP7_75t_L g502 ( .A(n_58), .Y(n_502) );
AOI22xp5_ASAP7_75t_L g610 ( .A1(n_59), .A2(n_96), .B1(n_554), .B2(n_575), .Y(n_610) );
INVx1_ASAP7_75t_L g123 ( .A(n_60), .Y(n_123) );
AND2x4_ASAP7_75t_L g145 ( .A(n_61), .B(n_146), .Y(n_145) );
AOI22xp33_ASAP7_75t_L g261 ( .A1(n_62), .A2(n_63), .B1(n_197), .B2(n_262), .Y(n_261) );
NAND2xp5_ASAP7_75t_L g227 ( .A(n_64), .B(n_120), .Y(n_227) );
NAND2xp5_ASAP7_75t_L g159 ( .A(n_65), .B(n_160), .Y(n_159) );
CKINVDCx5p33_ASAP7_75t_R g198 ( .A(n_66), .Y(n_198) );
NAND2xp5_ASAP7_75t_SL g213 ( .A(n_67), .B(n_197), .Y(n_213) );
INVx1_ASAP7_75t_L g146 ( .A(n_68), .Y(n_146) );
CKINVDCx5p33_ASAP7_75t_R g264 ( .A(n_69), .Y(n_264) );
NAND2xp5_ASAP7_75t_L g215 ( .A(n_70), .B(n_120), .Y(n_215) );
NAND2xp5_ASAP7_75t_L g169 ( .A(n_72), .B(n_127), .Y(n_169) );
NAND3xp33_ASAP7_75t_L g232 ( .A(n_73), .B(n_177), .C(n_214), .Y(n_232) );
NAND2xp5_ASAP7_75t_L g126 ( .A(n_75), .B(n_127), .Y(n_126) );
INVx2_ASAP7_75t_L g133 ( .A(n_76), .Y(n_133) );
NAND2xp5_ASAP7_75t_SL g152 ( .A(n_77), .B(n_153), .Y(n_152) );
NAND2xp5_ASAP7_75t_SL g224 ( .A(n_78), .B(n_142), .Y(n_224) );
NAND2xp5_ASAP7_75t_L g135 ( .A(n_79), .B(n_136), .Y(n_135) );
INVx1_ASAP7_75t_L g499 ( .A(n_80), .Y(n_499) );
XNOR2x1_ASAP7_75t_L g537 ( .A(n_80), .B(n_538), .Y(n_537) );
AOI22xp33_ASAP7_75t_L g630 ( .A1(n_81), .A2(n_97), .B1(n_140), .B2(n_197), .Y(n_630) );
CKINVDCx5p33_ASAP7_75t_R g568 ( .A(n_82), .Y(n_568) );
CKINVDCx5p33_ASAP7_75t_R g650 ( .A(n_83), .Y(n_650) );
AOI22xp33_ASAP7_75t_L g258 ( .A1(n_85), .A2(n_90), .B1(n_171), .B2(n_259), .Y(n_258) );
NAND2xp5_ASAP7_75t_L g222 ( .A(n_86), .B(n_142), .Y(n_222) );
NAND2xp33_ASAP7_75t_SL g158 ( .A(n_87), .B(n_130), .Y(n_158) );
NAND2xp5_ASAP7_75t_L g208 ( .A(n_88), .B(n_209), .Y(n_208) );
NAND2xp5_ASAP7_75t_SL g606 ( .A(n_89), .B(n_120), .Y(n_606) );
CKINVDCx5p33_ASAP7_75t_R g581 ( .A(n_91), .Y(n_581) );
NOR2xp33_ASAP7_75t_L g508 ( .A(n_92), .B(n_509), .Y(n_508) );
INVx1_ASAP7_75t_L g536 ( .A(n_92), .Y(n_536) );
NAND2xp33_ASAP7_75t_L g604 ( .A(n_93), .B(n_142), .Y(n_604) );
INVx1_ASAP7_75t_L g528 ( .A(n_94), .Y(n_528) );
NAND2xp33_ASAP7_75t_L g129 ( .A(n_95), .B(n_130), .Y(n_129) );
NAND2xp5_ASAP7_75t_L g180 ( .A(n_98), .B(n_160), .Y(n_180) );
NAND3xp33_ASAP7_75t_L g154 ( .A(n_99), .B(n_130), .C(n_153), .Y(n_154) );
NAND2xp5_ASAP7_75t_L g212 ( .A(n_101), .B(n_127), .Y(n_212) );
NAND2xp5_ASAP7_75t_SL g174 ( .A(n_102), .B(n_171), .Y(n_174) );
AOI21xp5_ASAP7_75t_L g103 ( .A1(n_104), .A2(n_106), .B(n_522), .Y(n_103) );
NAND2xp5_ASAP7_75t_SL g880 ( .A(n_104), .B(n_881), .Y(n_880) );
INVx2_ASAP7_75t_SL g890 ( .A(n_104), .Y(n_890) );
OAI22x1_ASAP7_75t_L g106 ( .A1(n_107), .A2(n_503), .B1(n_513), .B2(n_515), .Y(n_106) );
INVx2_ASAP7_75t_L g501 ( .A(n_108), .Y(n_501) );
XNOR2x1_ASAP7_75t_L g108 ( .A(n_109), .B(n_495), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_110), .Y(n_109) );
INVx2_ASAP7_75t_L g538 ( .A(n_110), .Y(n_538) );
NAND4xp75_ASAP7_75t_L g110 ( .A(n_111), .B(n_341), .C(n_414), .D(n_473), .Y(n_110) );
AND2x2_ASAP7_75t_L g111 ( .A(n_112), .B(n_297), .Y(n_111) );
NOR2xp33_ASAP7_75t_L g112 ( .A(n_113), .B(n_267), .Y(n_112) );
OAI221xp5_ASAP7_75t_L g113 ( .A1(n_114), .A2(n_200), .B1(n_239), .B2(n_244), .C(n_248), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_115), .Y(n_114) );
OAI21xp33_ASAP7_75t_SL g248 ( .A1(n_115), .A2(n_249), .B(n_253), .Y(n_248) );
AND2x2_ASAP7_75t_L g115 ( .A(n_116), .B(n_163), .Y(n_115) );
AND2x2_ASAP7_75t_L g294 ( .A(n_116), .B(n_251), .Y(n_294) );
NAND2xp5_ASAP7_75t_L g367 ( .A(n_116), .B(n_305), .Y(n_367) );
AND2x2_ASAP7_75t_L g116 ( .A(n_117), .B(n_147), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
BUFx2_ASAP7_75t_L g250 ( .A(n_118), .Y(n_250) );
INVx4_ASAP7_75t_L g273 ( .A(n_118), .Y(n_273) );
AND2x2_ASAP7_75t_L g301 ( .A(n_118), .B(n_164), .Y(n_301) );
OR2x2_ASAP7_75t_L g463 ( .A(n_118), .B(n_247), .Y(n_463) );
AND2x4_ASAP7_75t_L g118 ( .A(n_119), .B(n_124), .Y(n_118) );
INVx2_ASAP7_75t_L g648 ( .A(n_120), .Y(n_648) );
INVx4_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
AND2x4_ASAP7_75t_SL g143 ( .A(n_121), .B(n_144), .Y(n_143) );
INVx1_ASAP7_75t_SL g149 ( .A(n_121), .Y(n_149) );
INVx2_ASAP7_75t_L g205 ( .A(n_121), .Y(n_205) );
BUFx3_ASAP7_75t_L g589 ( .A(n_121), .Y(n_589) );
NOR2xp33_ASAP7_75t_L g590 ( .A(n_121), .B(n_591), .Y(n_590) );
INVx2_ASAP7_75t_SL g597 ( .A(n_121), .Y(n_597) );
NOR2xp33_ASAP7_75t_L g612 ( .A(n_121), .B(n_613), .Y(n_612) );
NOR2xp33_ASAP7_75t_L g649 ( .A(n_121), .B(n_650), .Y(n_649) );
BUFx6f_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
INVx2_ASAP7_75t_L g162 ( .A(n_122), .Y(n_162) );
OAI21x1_ASAP7_75t_L g124 ( .A1(n_125), .A2(n_134), .B(n_143), .Y(n_124) );
AOI21xp5_ASAP7_75t_L g125 ( .A1(n_126), .A2(n_129), .B(n_131), .Y(n_125) );
OAI22xp33_ASAP7_75t_L g195 ( .A1(n_127), .A2(n_196), .B1(n_197), .B2(n_198), .Y(n_195) );
INVx1_ASAP7_75t_L g556 ( .A(n_127), .Y(n_556) );
INVx1_ASAP7_75t_L g575 ( .A(n_127), .Y(n_575) );
INVx4_ASAP7_75t_L g577 ( .A(n_127), .Y(n_577) );
INVx3_ASAP7_75t_L g127 ( .A(n_128), .Y(n_127) );
BUFx6f_ASAP7_75t_L g130 ( .A(n_128), .Y(n_130) );
INVx1_ASAP7_75t_L g140 ( .A(n_128), .Y(n_140) );
BUFx6f_ASAP7_75t_L g142 ( .A(n_128), .Y(n_142) );
INVx1_ASAP7_75t_L g157 ( .A(n_128), .Y(n_157) );
INVx1_ASAP7_75t_L g172 ( .A(n_128), .Y(n_172) );
BUFx6f_ASAP7_75t_L g177 ( .A(n_128), .Y(n_177) );
INVx2_ASAP7_75t_L g192 ( .A(n_128), .Y(n_192) );
BUFx6f_ASAP7_75t_L g197 ( .A(n_128), .Y(n_197) );
INVx1_ASAP7_75t_L g209 ( .A(n_128), .Y(n_209) );
INVx1_ASAP7_75t_L g262 ( .A(n_128), .Y(n_262) );
INVx2_ASAP7_75t_L g226 ( .A(n_130), .Y(n_226) );
INVx1_ASAP7_75t_L g585 ( .A(n_130), .Y(n_585) );
AOI21xp5_ASAP7_75t_L g155 ( .A1(n_131), .A2(n_156), .B(n_158), .Y(n_155) );
AOI21xp5_ASAP7_75t_L g168 ( .A1(n_131), .A2(n_169), .B(n_170), .Y(n_168) );
AOI21xp5_ASAP7_75t_L g207 ( .A1(n_131), .A2(n_208), .B(n_210), .Y(n_207) );
BUFx4f_ASAP7_75t_L g131 ( .A(n_132), .Y(n_131) );
INVx1_ASAP7_75t_L g132 ( .A(n_133), .Y(n_132) );
INVx2_ASAP7_75t_L g138 ( .A(n_133), .Y(n_138) );
INVx1_ASAP7_75t_L g153 ( .A(n_133), .Y(n_153) );
BUFx8_ASAP7_75t_L g214 ( .A(n_133), .Y(n_214) );
OAI22xp5_ASAP7_75t_L g134 ( .A1(n_135), .A2(n_137), .B1(n_139), .B2(n_141), .Y(n_134) );
AOI21xp5_ASAP7_75t_L g223 ( .A1(n_136), .A2(n_224), .B(n_225), .Y(n_223) );
INVx2_ASAP7_75t_SL g136 ( .A(n_137), .Y(n_136) );
INVx2_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
BUFx3_ASAP7_75t_L g179 ( .A(n_138), .Y(n_179) );
INVx1_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
OAI21xp5_ASAP7_75t_L g151 ( .A1(n_142), .A2(n_152), .B(n_154), .Y(n_151) );
INVx1_ASAP7_75t_L g236 ( .A(n_142), .Y(n_236) );
INVx3_ASAP7_75t_L g554 ( .A(n_142), .Y(n_554) );
OAI21x1_ASAP7_75t_L g150 ( .A1(n_144), .A2(n_151), .B(n_155), .Y(n_150) );
OAI21x1_ASAP7_75t_L g167 ( .A1(n_144), .A2(n_168), .B(n_173), .Y(n_167) );
OAI21x1_ASAP7_75t_L g206 ( .A1(n_144), .A2(n_207), .B(n_211), .Y(n_206) );
OAI21x1_ASAP7_75t_L g218 ( .A1(n_144), .A2(n_219), .B(n_223), .Y(n_218) );
OAI21x1_ASAP7_75t_L g229 ( .A1(n_144), .A2(n_230), .B(n_233), .Y(n_229) );
BUFx10_ASAP7_75t_L g144 ( .A(n_145), .Y(n_144) );
BUFx10_ASAP7_75t_L g187 ( .A(n_145), .Y(n_187) );
INVx1_ASAP7_75t_L g566 ( .A(n_145), .Y(n_566) );
INVx2_ASAP7_75t_L g276 ( .A(n_147), .Y(n_276) );
HB1xp67_ASAP7_75t_L g302 ( .A(n_147), .Y(n_302) );
INVx1_ASAP7_75t_L g312 ( .A(n_147), .Y(n_312) );
INVx2_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
INVx1_ASAP7_75t_L g247 ( .A(n_148), .Y(n_247) );
AND2x2_ASAP7_75t_L g403 ( .A(n_148), .B(n_182), .Y(n_403) );
OAI21x1_ASAP7_75t_L g148 ( .A1(n_149), .A2(n_150), .B(n_159), .Y(n_148) );
INVx1_ASAP7_75t_L g237 ( .A(n_153), .Y(n_237) );
INVx1_ASAP7_75t_SL g578 ( .A(n_153), .Y(n_578) );
INVx1_ASAP7_75t_L g631 ( .A(n_153), .Y(n_631) );
INVx1_ASAP7_75t_L g586 ( .A(n_157), .Y(n_586) );
INVx2_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
INVx2_ASAP7_75t_L g166 ( .A(n_161), .Y(n_166) );
NOR2xp33_ASAP7_75t_L g558 ( .A(n_161), .B(n_559), .Y(n_558) );
NOR2xp33_ASAP7_75t_L g567 ( .A(n_161), .B(n_568), .Y(n_567) );
INVx2_ASAP7_75t_L g161 ( .A(n_162), .Y(n_161) );
INVx2_ASAP7_75t_L g185 ( .A(n_162), .Y(n_185) );
INVx2_ASAP7_75t_L g265 ( .A(n_162), .Y(n_265) );
INVx2_ASAP7_75t_L g360 ( .A(n_163), .Y(n_360) );
AND2x2_ASAP7_75t_L g364 ( .A(n_163), .B(n_276), .Y(n_364) );
NAND2xp5_ASAP7_75t_L g493 ( .A(n_163), .B(n_395), .Y(n_493) );
AND2x2_ASAP7_75t_L g163 ( .A(n_164), .B(n_181), .Y(n_163) );
INVx2_ASAP7_75t_L g327 ( .A(n_164), .Y(n_327) );
AND2x2_ASAP7_75t_L g421 ( .A(n_164), .B(n_287), .Y(n_421) );
AND2x2_ASAP7_75t_L g472 ( .A(n_164), .B(n_273), .Y(n_472) );
INVx2_ASAP7_75t_L g164 ( .A(n_165), .Y(n_164) );
INVx1_ASAP7_75t_L g246 ( .A(n_165), .Y(n_246) );
OAI21x1_ASAP7_75t_L g165 ( .A1(n_166), .A2(n_167), .B(n_180), .Y(n_165) );
OAI21xp5_ASAP7_75t_L g217 ( .A1(n_166), .A2(n_218), .B(n_227), .Y(n_217) );
OAI21x1_ASAP7_75t_L g243 ( .A1(n_166), .A2(n_218), .B(n_227), .Y(n_243) );
OAI21xp33_ASAP7_75t_SL g252 ( .A1(n_166), .A2(n_167), .B(n_180), .Y(n_252) );
INVx1_ASAP7_75t_L g574 ( .A(n_171), .Y(n_574) );
INVx2_ASAP7_75t_L g171 ( .A(n_172), .Y(n_171) );
AOI21xp5_ASAP7_75t_L g173 ( .A1(n_174), .A2(n_175), .B(n_178), .Y(n_173) );
INVx2_ASAP7_75t_L g176 ( .A(n_177), .Y(n_176) );
INVx2_ASAP7_75t_L g178 ( .A(n_179), .Y(n_178) );
INVx2_ASAP7_75t_L g194 ( .A(n_179), .Y(n_194) );
AND2x2_ASAP7_75t_L g251 ( .A(n_181), .B(n_252), .Y(n_251) );
INVx1_ASAP7_75t_L g181 ( .A(n_182), .Y(n_181) );
INVx2_ASAP7_75t_L g275 ( .A(n_182), .Y(n_275) );
AOI21x1_ASAP7_75t_L g182 ( .A1(n_183), .A2(n_188), .B(n_199), .Y(n_182) );
NOR2xp67_ASAP7_75t_SL g183 ( .A(n_184), .B(n_186), .Y(n_183) );
INVx2_ASAP7_75t_L g557 ( .A(n_184), .Y(n_557) );
INVx2_ASAP7_75t_L g184 ( .A(n_185), .Y(n_184) );
AO31x2_ASAP7_75t_L g256 ( .A1(n_185), .A2(n_187), .A3(n_257), .B(n_263), .Y(n_256) );
NOR2xp33_ASAP7_75t_SL g580 ( .A(n_185), .B(n_581), .Y(n_580) );
NOR2xp33_ASAP7_75t_L g632 ( .A(n_185), .B(n_633), .Y(n_632) );
INVx1_ASAP7_75t_L g551 ( .A(n_186), .Y(n_551) );
INVx2_ASAP7_75t_L g186 ( .A(n_187), .Y(n_186) );
AO31x2_ASAP7_75t_L g571 ( .A1(n_187), .A2(n_572), .A3(n_579), .B(n_580), .Y(n_571) );
AO31x2_ASAP7_75t_L g582 ( .A1(n_187), .A2(n_583), .A3(n_589), .B(n_590), .Y(n_582) );
AO31x2_ASAP7_75t_L g644 ( .A1(n_187), .A2(n_645), .A3(n_648), .B(n_649), .Y(n_644) );
NAND2xp5_ASAP7_75t_L g188 ( .A(n_189), .B(n_193), .Y(n_188) );
NOR2xp33_ASAP7_75t_L g190 ( .A(n_191), .B(n_192), .Y(n_190) );
INVx2_ASAP7_75t_SL g629 ( .A(n_192), .Y(n_629) );
NAND2xp5_ASAP7_75t_L g193 ( .A(n_194), .B(n_195), .Y(n_193) );
OAI22xp5_ASAP7_75t_L g257 ( .A1(n_194), .A2(n_258), .B1(n_260), .B2(n_261), .Y(n_257) );
OAI22xp5_ASAP7_75t_L g552 ( .A1(n_194), .A2(n_260), .B1(n_553), .B2(n_555), .Y(n_552) );
OAI22xp5_ASAP7_75t_L g562 ( .A1(n_194), .A2(n_260), .B1(n_563), .B2(n_564), .Y(n_562) );
OAI22xp5_ASAP7_75t_L g583 ( .A1(n_194), .A2(n_260), .B1(n_584), .B2(n_587), .Y(n_583) );
OAI22xp5_ASAP7_75t_L g645 ( .A1(n_194), .A2(n_260), .B1(n_646), .B2(n_647), .Y(n_645) );
OAI21xp5_ASAP7_75t_L g230 ( .A1(n_197), .A2(n_231), .B(n_232), .Y(n_230) );
INVx2_ASAP7_75t_L g259 ( .A(n_197), .Y(n_259) );
INVx1_ASAP7_75t_L g200 ( .A(n_201), .Y(n_200) );
AND2x2_ASAP7_75t_L g201 ( .A(n_202), .B(n_216), .Y(n_201) );
INVx2_ASAP7_75t_L g240 ( .A(n_202), .Y(n_240) );
AND2x2_ASAP7_75t_L g404 ( .A(n_202), .B(n_254), .Y(n_404) );
NAND2xp5_ASAP7_75t_L g411 ( .A(n_202), .B(n_412), .Y(n_411) );
NAND2xp5_ASAP7_75t_L g434 ( .A(n_202), .B(n_425), .Y(n_434) );
OR2x2_ASAP7_75t_L g457 ( .A(n_202), .B(n_316), .Y(n_457) );
INVx3_ASAP7_75t_L g202 ( .A(n_203), .Y(n_202) );
NOR2xp67_ASAP7_75t_L g340 ( .A(n_203), .B(n_283), .Y(n_340) );
AND2x2_ASAP7_75t_L g446 ( .A(n_203), .B(n_255), .Y(n_446) );
BUFx3_ASAP7_75t_L g203 ( .A(n_204), .Y(n_203) );
INVx1_ASAP7_75t_L g280 ( .A(n_204), .Y(n_280) );
OAI21x1_ASAP7_75t_L g204 ( .A1(n_205), .A2(n_206), .B(n_215), .Y(n_204) );
OA21x2_ASAP7_75t_L g228 ( .A1(n_205), .A2(n_229), .B(n_238), .Y(n_228) );
OAI21x1_ASAP7_75t_L g255 ( .A1(n_205), .A2(n_229), .B(n_238), .Y(n_255) );
OAI21x1_ASAP7_75t_L g292 ( .A1(n_205), .A2(n_206), .B(n_215), .Y(n_292) );
INVx2_ASAP7_75t_L g221 ( .A(n_209), .Y(n_221) );
AOI21xp5_ASAP7_75t_L g211 ( .A1(n_212), .A2(n_213), .B(n_214), .Y(n_211) );
O2A1O1Ixp5_ASAP7_75t_L g219 ( .A1(n_214), .A2(n_220), .B(n_221), .C(n_222), .Y(n_219) );
INVx6_ASAP7_75t_L g260 ( .A(n_214), .Y(n_260) );
O2A1O1Ixp5_ASAP7_75t_L g599 ( .A1(n_214), .A2(n_577), .B(n_600), .C(n_601), .Y(n_599) );
AND2x2_ASAP7_75t_L g333 ( .A(n_216), .B(n_278), .Y(n_333) );
NAND2xp5_ASAP7_75t_L g369 ( .A(n_216), .B(n_370), .Y(n_369) );
NAND2xp5_ASAP7_75t_L g397 ( .A(n_216), .B(n_389), .Y(n_397) );
AND2x2_ASAP7_75t_L g216 ( .A(n_217), .B(n_228), .Y(n_216) );
AND2x2_ASAP7_75t_L g309 ( .A(n_217), .B(n_255), .Y(n_309) );
INVx1_ASAP7_75t_L g453 ( .A(n_217), .Y(n_453) );
AND2x2_ASAP7_75t_L g241 ( .A(n_228), .B(n_242), .Y(n_241) );
OR2x2_ASAP7_75t_L g316 ( .A(n_228), .B(n_256), .Y(n_316) );
NAND2xp5_ASAP7_75t_L g374 ( .A(n_228), .B(n_256), .Y(n_374) );
AOI21x1_ASAP7_75t_L g233 ( .A1(n_234), .A2(n_235), .B(n_237), .Y(n_233) );
NAND2xp5_ASAP7_75t_L g239 ( .A(n_240), .B(n_241), .Y(n_239) );
NAND2xp5_ASAP7_75t_L g356 ( .A(n_240), .B(n_357), .Y(n_356) );
AND2x4_ASAP7_75t_L g479 ( .A(n_240), .B(n_282), .Y(n_479) );
AND2x2_ASAP7_75t_L g409 ( .A(n_241), .B(n_410), .Y(n_409) );
INVxp67_ASAP7_75t_SL g266 ( .A(n_242), .Y(n_266) );
AND2x2_ASAP7_75t_L g290 ( .A(n_242), .B(n_291), .Y(n_290) );
BUFx3_ASAP7_75t_L g296 ( .A(n_242), .Y(n_296) );
INVxp67_ASAP7_75t_SL g332 ( .A(n_242), .Y(n_332) );
INVx1_ASAP7_75t_L g357 ( .A(n_242), .Y(n_357) );
AND2x2_ASAP7_75t_L g363 ( .A(n_242), .B(n_255), .Y(n_363) );
INVx1_ASAP7_75t_L g444 ( .A(n_242), .Y(n_444) );
INVx3_ASAP7_75t_L g242 ( .A(n_243), .Y(n_242) );
INVx1_ASAP7_75t_L g244 ( .A(n_245), .Y(n_244) );
AND2x2_ASAP7_75t_L g286 ( .A(n_245), .B(n_287), .Y(n_286) );
AOI32xp33_ASAP7_75t_SL g418 ( .A1(n_245), .A2(n_310), .A3(n_419), .B1(n_421), .B2(n_422), .Y(n_418) );
AND2x2_ASAP7_75t_L g245 ( .A(n_246), .B(n_247), .Y(n_245) );
INVx2_ASAP7_75t_L g271 ( .A(n_246), .Y(n_271) );
OR2x2_ASAP7_75t_L g320 ( .A(n_246), .B(n_276), .Y(n_320) );
HB1xp67_ASAP7_75t_L g324 ( .A(n_247), .Y(n_324) );
INVxp67_ASAP7_75t_L g350 ( .A(n_247), .Y(n_350) );
OR2x2_ASAP7_75t_L g452 ( .A(n_247), .B(n_453), .Y(n_452) );
AND2x2_ASAP7_75t_L g249 ( .A(n_250), .B(n_251), .Y(n_249) );
OR3x2_ASAP7_75t_L g317 ( .A(n_250), .B(n_318), .C(n_320), .Y(n_317) );
INVx1_ASAP7_75t_L g423 ( .A(n_250), .Y(n_423) );
AND2x2_ASAP7_75t_L g351 ( .A(n_251), .B(n_352), .Y(n_351) );
INVx1_ASAP7_75t_L g407 ( .A(n_251), .Y(n_407) );
NAND2xp5_ASAP7_75t_L g413 ( .A(n_251), .B(n_302), .Y(n_413) );
BUFx2_ASAP7_75t_L g306 ( .A(n_252), .Y(n_306) );
AND2x2_ASAP7_75t_L g253 ( .A(n_254), .B(n_266), .Y(n_253) );
NAND2xp5_ASAP7_75t_L g289 ( .A(n_254), .B(n_290), .Y(n_289) );
HB1xp67_ASAP7_75t_L g486 ( .A(n_254), .Y(n_486) );
AND2x2_ASAP7_75t_L g254 ( .A(n_255), .B(n_256), .Y(n_254) );
INVx1_ASAP7_75t_L g283 ( .A(n_255), .Y(n_283) );
INVx1_ASAP7_75t_L g425 ( .A(n_255), .Y(n_425) );
INVx1_ASAP7_75t_L g284 ( .A(n_256), .Y(n_284) );
HB1xp67_ASAP7_75t_L g330 ( .A(n_256), .Y(n_330) );
OR2x2_ASAP7_75t_L g371 ( .A(n_256), .B(n_292), .Y(n_371) );
AND2x2_ASAP7_75t_L g389 ( .A(n_256), .B(n_292), .Y(n_389) );
AND2x2_ASAP7_75t_L g410 ( .A(n_256), .B(n_280), .Y(n_410) );
OAI22xp5_ASAP7_75t_L g572 ( .A1(n_260), .A2(n_573), .B1(n_576), .B2(n_578), .Y(n_572) );
AOI21xp5_ASAP7_75t_L g602 ( .A1(n_260), .A2(n_603), .B(n_604), .Y(n_602) );
OAI22xp5_ASAP7_75t_L g609 ( .A1(n_260), .A2(n_578), .B1(n_610), .B2(n_611), .Y(n_609) );
OAI22xp5_ASAP7_75t_L g627 ( .A1(n_260), .A2(n_628), .B1(n_630), .B2(n_631), .Y(n_627) );
INVx1_ASAP7_75t_L g588 ( .A(n_262), .Y(n_588) );
NOR2xp33_ASAP7_75t_L g263 ( .A(n_264), .B(n_265), .Y(n_263) );
BUFx2_ASAP7_75t_L g579 ( .A(n_265), .Y(n_579) );
BUFx2_ASAP7_75t_L g478 ( .A(n_266), .Y(n_478) );
NAND3xp33_ASAP7_75t_L g267 ( .A(n_268), .B(n_285), .C(n_293), .Y(n_267) );
NAND2xp5_ASAP7_75t_L g268 ( .A(n_269), .B(n_277), .Y(n_268) );
INVx3_ASAP7_75t_L g400 ( .A(n_269), .Y(n_400) );
AND2x4_ASAP7_75t_L g269 ( .A(n_270), .B(n_274), .Y(n_269) );
AND2x2_ASAP7_75t_L g270 ( .A(n_271), .B(n_272), .Y(n_270) );
AND2x2_ASAP7_75t_L g430 ( .A(n_271), .B(n_386), .Y(n_430) );
INVx1_ASAP7_75t_L g352 ( .A(n_272), .Y(n_352) );
NAND2xp5_ASAP7_75t_SL g385 ( .A(n_272), .B(n_386), .Y(n_385) );
AND2x2_ASAP7_75t_L g437 ( .A(n_272), .B(n_276), .Y(n_437) );
INVx2_ASAP7_75t_L g272 ( .A(n_273), .Y(n_272) );
OR2x2_ASAP7_75t_L g311 ( .A(n_273), .B(n_312), .Y(n_311) );
NAND2x1_ASAP7_75t_L g326 ( .A(n_273), .B(n_327), .Y(n_326) );
BUFx2_ASAP7_75t_L g395 ( .A(n_273), .Y(n_395) );
NAND2xp33_ASAP7_75t_R g378 ( .A(n_274), .B(n_301), .Y(n_378) );
AND2x2_ASAP7_75t_L g394 ( .A(n_274), .B(n_395), .Y(n_394) );
INVx1_ASAP7_75t_L g460 ( .A(n_274), .Y(n_460) );
AND2x2_ASAP7_75t_L g274 ( .A(n_275), .B(n_276), .Y(n_274) );
INVx2_ASAP7_75t_L g287 ( .A(n_275), .Y(n_287) );
INVx1_ASAP7_75t_L g319 ( .A(n_275), .Y(n_319) );
INVx2_ASAP7_75t_L g386 ( .A(n_275), .Y(n_386) );
NAND2xp5_ASAP7_75t_L g471 ( .A(n_276), .B(n_472), .Y(n_471) );
NOR2xp33_ASAP7_75t_L g277 ( .A(n_278), .B(n_281), .Y(n_277) );
INVx2_ASAP7_75t_L g278 ( .A(n_279), .Y(n_278) );
AND2x2_ASAP7_75t_L g308 ( .A(n_279), .B(n_309), .Y(n_308) );
BUFx2_ASAP7_75t_L g279 ( .A(n_280), .Y(n_279) );
INVx2_ASAP7_75t_L g281 ( .A(n_282), .Y(n_281) );
AND2x2_ASAP7_75t_L g295 ( .A(n_282), .B(n_296), .Y(n_295) );
AND2x4_ASAP7_75t_L g466 ( .A(n_282), .B(n_357), .Y(n_466) );
AND2x4_ASAP7_75t_L g282 ( .A(n_283), .B(n_284), .Y(n_282) );
AND2x2_ASAP7_75t_L g347 ( .A(n_284), .B(n_292), .Y(n_347) );
NAND2xp5_ASAP7_75t_L g285 ( .A(n_286), .B(n_288), .Y(n_285) );
INVx1_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
AND2x2_ASAP7_75t_L g314 ( .A(n_290), .B(n_315), .Y(n_314) );
INVx1_ASAP7_75t_L g417 ( .A(n_291), .Y(n_417) );
INVx1_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
NAND2xp5_ASAP7_75t_L g293 ( .A(n_294), .B(n_295), .Y(n_293) );
INVx2_ASAP7_75t_L g475 ( .A(n_294), .Y(n_475) );
INVx1_ASAP7_75t_L g303 ( .A(n_295), .Y(n_303) );
NAND2xp5_ASAP7_75t_L g339 ( .A(n_296), .B(n_340), .Y(n_339) );
OR2x2_ASAP7_75t_L g373 ( .A(n_296), .B(n_374), .Y(n_373) );
INVx2_ASAP7_75t_L g420 ( .A(n_296), .Y(n_420) );
NAND2xp5_ASAP7_75t_SL g469 ( .A(n_296), .B(n_370), .Y(n_469) );
NOR3xp33_ASAP7_75t_L g297 ( .A(n_298), .B(n_304), .C(n_321), .Y(n_297) );
NOR2xp33_ASAP7_75t_L g298 ( .A(n_299), .B(n_303), .Y(n_298) );
INVx3_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
AND2x2_ASAP7_75t_L g300 ( .A(n_301), .B(n_302), .Y(n_300) );
AND2x2_ASAP7_75t_L g335 ( .A(n_301), .B(n_336), .Y(n_335) );
INVx1_ASAP7_75t_L g428 ( .A(n_301), .Y(n_428) );
OAI22xp5_ASAP7_75t_L g304 ( .A1(n_305), .A2(n_307), .B1(n_313), .B2(n_317), .Y(n_304) );
NAND3x2_ASAP7_75t_L g447 ( .A(n_305), .B(n_448), .C(n_449), .Y(n_447) );
INVx2_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
NAND2xp5_ASAP7_75t_L g307 ( .A(n_308), .B(n_310), .Y(n_307) );
NAND2x1_ASAP7_75t_L g387 ( .A(n_309), .B(n_388), .Y(n_387) );
INVx1_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
OR2x2_ASAP7_75t_L g359 ( .A(n_311), .B(n_360), .Y(n_359) );
INVx1_ASAP7_75t_L g431 ( .A(n_311), .Y(n_431) );
INVxp67_ASAP7_75t_SL g313 ( .A(n_314), .Y(n_313) );
AND2x4_ASAP7_75t_L g483 ( .A(n_315), .B(n_416), .Y(n_483) );
INVx2_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
INVx1_ASAP7_75t_L g345 ( .A(n_316), .Y(n_345) );
NOR2x1p5_ASAP7_75t_SL g392 ( .A(n_318), .B(n_320), .Y(n_392) );
INVx1_ASAP7_75t_L g318 ( .A(n_319), .Y(n_318) );
INVx1_ASAP7_75t_L g336 ( .A(n_319), .Y(n_336) );
HB1xp67_ASAP7_75t_L g438 ( .A(n_319), .Y(n_438) );
OAI22xp33_ASAP7_75t_SL g321 ( .A1(n_322), .A2(n_328), .B1(n_334), .B2(n_337), .Y(n_321) );
NAND2xp5_ASAP7_75t_L g322 ( .A(n_323), .B(n_325), .Y(n_322) );
INVx1_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
OR2x2_ASAP7_75t_L g481 ( .A(n_324), .B(n_428), .Y(n_481) );
INVxp67_ASAP7_75t_SL g325 ( .A(n_326), .Y(n_325) );
OR2x6_ASAP7_75t_L g401 ( .A(n_326), .B(n_402), .Y(n_401) );
NOR2xp33_ASAP7_75t_SL g328 ( .A(n_329), .B(n_333), .Y(n_328) );
NOR2xp33_ASAP7_75t_L g329 ( .A(n_330), .B(n_331), .Y(n_329) );
INVx1_ASAP7_75t_L g383 ( .A(n_330), .Y(n_383) );
INVx1_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
INVx1_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
AOI22xp5_ASAP7_75t_L g450 ( .A1(n_335), .A2(n_451), .B1(n_456), .B2(n_458), .Y(n_450) );
AOI22xp5_ASAP7_75t_L g485 ( .A1(n_335), .A2(n_429), .B1(n_486), .B2(n_487), .Y(n_485) );
NAND2xp5_ASAP7_75t_L g490 ( .A(n_335), .B(n_483), .Y(n_490) );
INVx1_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
INVx1_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
NOR2x1_ASAP7_75t_L g341 ( .A(n_342), .B(n_375), .Y(n_341) );
NAND3xp33_ASAP7_75t_SL g342 ( .A(n_343), .B(n_353), .C(n_365), .Y(n_342) );
AO21x1_ASAP7_75t_L g343 ( .A1(n_344), .A2(n_346), .B(n_348), .Y(n_343) );
INVx1_ASAP7_75t_L g445 ( .A(n_344), .Y(n_445) );
INVx1_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
INVx1_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
NAND2x1p5_ASAP7_75t_L g348 ( .A(n_349), .B(n_351), .Y(n_348) );
AOI32xp33_ASAP7_75t_L g465 ( .A1(n_349), .A2(n_466), .A3(n_467), .B1(n_468), .B2(n_470), .Y(n_465) );
BUFx2_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
BUFx2_ASAP7_75t_L g448 ( .A(n_352), .Y(n_448) );
AOI22xp5_ASAP7_75t_L g353 ( .A1(n_354), .A2(n_358), .B1(n_361), .B2(n_364), .Y(n_353) );
INVxp67_ASAP7_75t_SL g354 ( .A(n_355), .Y(n_354) );
HB1xp67_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
INVx1_ASAP7_75t_L g381 ( .A(n_357), .Y(n_381) );
NAND2xp5_ASAP7_75t_L g390 ( .A(n_357), .B(n_389), .Y(n_390) );
AOI22xp33_ASAP7_75t_SL g365 ( .A1(n_358), .A2(n_366), .B1(n_368), .B2(n_372), .Y(n_365) );
INVx1_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
OR2x2_ASAP7_75t_L g462 ( .A(n_360), .B(n_463), .Y(n_462) );
INVx1_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
OAI322xp33_ASAP7_75t_L g474 ( .A1(n_362), .A2(n_455), .A3(n_475), .B1(n_476), .B2(n_480), .C1(n_481), .C2(n_482), .Y(n_474) );
INVx2_ASAP7_75t_SL g362 ( .A(n_363), .Y(n_362) );
AND2x2_ASAP7_75t_L g494 ( .A(n_363), .B(n_383), .Y(n_494) );
INVx1_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
INVx1_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
INVx1_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
INVx1_ASAP7_75t_L g455 ( .A(n_371), .Y(n_455) );
NAND2xp5_ASAP7_75t_L g435 ( .A(n_372), .B(n_436), .Y(n_435) );
INVx2_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
INVx1_ASAP7_75t_L g412 ( .A(n_374), .Y(n_412) );
NAND2xp5_ASAP7_75t_L g375 ( .A(n_376), .B(n_398), .Y(n_375) );
AOI211xp5_ASAP7_75t_L g376 ( .A1(n_377), .A2(n_379), .B(n_384), .C(n_393), .Y(n_376) );
INVxp67_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
INVx1_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
NAND2xp5_ASAP7_75t_L g380 ( .A(n_381), .B(n_382), .Y(n_380) );
INVx1_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
OAI22xp33_ASAP7_75t_L g384 ( .A1(n_385), .A2(n_387), .B1(n_390), .B2(n_391), .Y(n_384) );
INVx1_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
NAND2xp5_ASAP7_75t_L g442 ( .A(n_389), .B(n_443), .Y(n_442) );
NAND2xp5_ASAP7_75t_L g488 ( .A(n_389), .B(n_425), .Y(n_488) );
INVx1_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
AND2x2_ASAP7_75t_L g393 ( .A(n_394), .B(n_396), .Y(n_393) );
INVxp67_ASAP7_75t_SL g396 ( .A(n_397), .Y(n_396) );
AOI21xp5_ASAP7_75t_L g398 ( .A1(n_399), .A2(n_404), .B(n_405), .Y(n_398) );
NAND2x1_ASAP7_75t_L g399 ( .A(n_400), .B(n_401), .Y(n_399) );
NOR2x1_ASAP7_75t_SL g427 ( .A(n_402), .B(n_428), .Y(n_427) );
INVx1_ASAP7_75t_L g449 ( .A(n_402), .Y(n_449) );
INVx2_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
INVx2_ASAP7_75t_L g464 ( .A(n_404), .Y(n_464) );
OAI22xp5_ASAP7_75t_L g405 ( .A1(n_406), .A2(n_408), .B1(n_411), .B2(n_413), .Y(n_405) );
HB1xp67_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
INVx1_ASAP7_75t_L g467 ( .A(n_407), .Y(n_467) );
INVx1_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
NOR3x1_ASAP7_75t_L g414 ( .A(n_415), .B(n_439), .C(n_461), .Y(n_414) );
OAI211xp5_ASAP7_75t_L g415 ( .A1(n_416), .A2(n_418), .B(n_426), .C(n_435), .Y(n_415) );
INVx1_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
INVxp67_ASAP7_75t_SL g419 ( .A(n_420), .Y(n_419) );
OR2x2_ASAP7_75t_L g433 ( .A(n_420), .B(n_434), .Y(n_433) );
NAND2xp5_ASAP7_75t_L g459 ( .A(n_421), .B(n_423), .Y(n_459) );
NOR2xp33_ASAP7_75t_L g422 ( .A(n_423), .B(n_424), .Y(n_422) );
INVx2_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
OAI21xp5_ASAP7_75t_SL g426 ( .A1(n_427), .A2(n_429), .B(n_432), .Y(n_426) );
AND2x2_ASAP7_75t_L g429 ( .A(n_430), .B(n_431), .Y(n_429) );
INVxp67_ASAP7_75t_L g480 ( .A(n_430), .Y(n_480) );
INVx1_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
AND2x2_ASAP7_75t_L g436 ( .A(n_437), .B(n_438), .Y(n_436) );
OAI21xp5_ASAP7_75t_L g439 ( .A1(n_440), .A2(n_447), .B(n_450), .Y(n_439) );
NOR3xp33_ASAP7_75t_L g440 ( .A(n_441), .B(n_445), .C(n_446), .Y(n_440) );
INVx1_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
INVx1_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
NOR2xp33_ASAP7_75t_L g451 ( .A(n_452), .B(n_454), .Y(n_451) );
INVx1_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
INVx2_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
NAND2xp5_ASAP7_75t_SL g458 ( .A(n_459), .B(n_460), .Y(n_458) );
OAI21xp5_ASAP7_75t_SL g461 ( .A1(n_462), .A2(n_464), .B(n_465), .Y(n_461) );
INVx1_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
INVx1_ASAP7_75t_L g470 ( .A(n_471), .Y(n_470) );
NOR3xp33_ASAP7_75t_L g473 ( .A(n_474), .B(n_484), .C(n_489), .Y(n_473) );
NAND2x1p5_ASAP7_75t_L g476 ( .A(n_477), .B(n_479), .Y(n_476) );
INVx1_ASAP7_75t_L g477 ( .A(n_478), .Y(n_477) );
INVx2_ASAP7_75t_L g482 ( .A(n_483), .Y(n_482) );
INVx1_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
INVx1_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
NAND2xp33_ASAP7_75t_SL g489 ( .A(n_490), .B(n_491), .Y(n_489) );
NAND2xp5_ASAP7_75t_L g491 ( .A(n_492), .B(n_494), .Y(n_491) );
INVx1_ASAP7_75t_L g492 ( .A(n_493), .Y(n_492) );
INVx1_ASAP7_75t_L g496 ( .A(n_497), .Y(n_496) );
CKINVDCx5p33_ASAP7_75t_R g503 ( .A(n_504), .Y(n_503) );
AND2x2_ASAP7_75t_L g504 ( .A(n_505), .B(n_506), .Y(n_504) );
INVx3_ASAP7_75t_L g514 ( .A(n_505), .Y(n_514) );
NOR2xp33_ASAP7_75t_L g891 ( .A(n_505), .B(n_892), .Y(n_891) );
INVx5_ASAP7_75t_L g506 ( .A(n_507), .Y(n_506) );
INVx4_ASAP7_75t_L g520 ( .A(n_507), .Y(n_520) );
CKINVDCx8_ASAP7_75t_R g886 ( .A(n_507), .Y(n_886) );
INVx3_ASAP7_75t_L g892 ( .A(n_507), .Y(n_892) );
AND2x6_ASAP7_75t_SL g507 ( .A(n_508), .B(n_511), .Y(n_507) );
INVx1_ASAP7_75t_L g509 ( .A(n_510), .Y(n_509) );
INVx1_ASAP7_75t_L g511 ( .A(n_512), .Y(n_511) );
NOR2x1_ASAP7_75t_L g876 ( .A(n_512), .B(n_877), .Y(n_876) );
BUFx8_ASAP7_75t_SL g513 ( .A(n_514), .Y(n_513) );
BUFx2_ASAP7_75t_L g881 ( .A(n_514), .Y(n_881) );
INVxp67_ASAP7_75t_SL g515 ( .A(n_516), .Y(n_515) );
NOR2xp67_ASAP7_75t_SL g516 ( .A(n_517), .B(n_521), .Y(n_516) );
CKINVDCx5p33_ASAP7_75t_R g517 ( .A(n_518), .Y(n_517) );
INVx4_ASAP7_75t_L g518 ( .A(n_519), .Y(n_518) );
BUFx12f_ASAP7_75t_L g519 ( .A(n_520), .Y(n_519) );
OAI21xp33_ASAP7_75t_L g522 ( .A1(n_523), .A2(n_873), .B(n_882), .Y(n_522) );
AOI22xp5_ASAP7_75t_L g523 ( .A1(n_524), .A2(n_530), .B1(n_871), .B2(n_872), .Y(n_523) );
INVx1_ASAP7_75t_L g871 ( .A(n_524), .Y(n_871) );
INVx1_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
INVx1_ASAP7_75t_L g872 ( .A(n_530), .Y(n_872) );
AOI21x1_ASAP7_75t_L g530 ( .A1(n_531), .A2(n_537), .B(n_539), .Y(n_530) );
CKINVDCx5p33_ASAP7_75t_R g531 ( .A(n_532), .Y(n_531) );
INVx8_ASAP7_75t_L g532 ( .A(n_533), .Y(n_532) );
BUFx12f_ASAP7_75t_L g533 ( .A(n_534), .Y(n_533) );
CKINVDCx5p33_ASAP7_75t_R g534 ( .A(n_535), .Y(n_534) );
BUFx8_ASAP7_75t_SL g541 ( .A(n_535), .Y(n_541) );
AND2x2_ASAP7_75t_L g879 ( .A(n_535), .B(n_876), .Y(n_879) );
INVx2_ASAP7_75t_L g535 ( .A(n_536), .Y(n_535) );
NOR2x1_ASAP7_75t_L g539 ( .A(n_540), .B(n_542), .Y(n_539) );
CKINVDCx5p33_ASAP7_75t_R g540 ( .A(n_541), .Y(n_540) );
AND3x4_ASAP7_75t_L g542 ( .A(n_543), .B(n_768), .C(n_846), .Y(n_542) );
NOR2x1_ASAP7_75t_L g543 ( .A(n_544), .B(n_711), .Y(n_543) );
NAND3xp33_ASAP7_75t_L g544 ( .A(n_545), .B(n_658), .C(n_681), .Y(n_544) );
AOI221x1_ASAP7_75t_L g545 ( .A1(n_546), .A2(n_592), .B1(n_614), .B2(n_623), .C(n_634), .Y(n_545) );
AND2x2_ASAP7_75t_L g546 ( .A(n_547), .B(n_569), .Y(n_546) );
AND2x4_ASAP7_75t_L g748 ( .A(n_547), .B(n_749), .Y(n_748) );
INVx2_ASAP7_75t_L g547 ( .A(n_548), .Y(n_547) );
OR2x2_ASAP7_75t_L g548 ( .A(n_549), .B(n_560), .Y(n_548) );
INVx2_ASAP7_75t_L g707 ( .A(n_549), .Y(n_707) );
INVx1_ASAP7_75t_L g734 ( .A(n_549), .Y(n_734) );
INVx2_ASAP7_75t_L g549 ( .A(n_550), .Y(n_549) );
INVx2_ASAP7_75t_L g617 ( .A(n_550), .Y(n_617) );
AND2x4_ASAP7_75t_L g685 ( .A(n_550), .B(n_618), .Y(n_685) );
AO31x2_ASAP7_75t_L g550 ( .A1(n_551), .A2(n_552), .A3(n_557), .B(n_558), .Y(n_550) );
AO31x2_ASAP7_75t_L g608 ( .A1(n_551), .A2(n_579), .A3(n_609), .B(n_612), .Y(n_608) );
AO31x2_ASAP7_75t_L g561 ( .A1(n_557), .A2(n_562), .A3(n_565), .B(n_567), .Y(n_561) );
INVx1_ASAP7_75t_L g767 ( .A(n_560), .Y(n_767) );
INVx2_ASAP7_75t_L g560 ( .A(n_561), .Y(n_560) );
INVx2_ASAP7_75t_L g618 ( .A(n_561), .Y(n_618) );
AND2x4_ASAP7_75t_L g656 ( .A(n_561), .B(n_657), .Y(n_656) );
OR2x2_ASAP7_75t_L g676 ( .A(n_561), .B(n_582), .Y(n_676) );
HB1xp67_ASAP7_75t_L g728 ( .A(n_561), .Y(n_728) );
INVx1_ASAP7_75t_L g821 ( .A(n_561), .Y(n_821) );
AND2x2_ASAP7_75t_L g867 ( .A(n_561), .B(n_571), .Y(n_867) );
AO31x2_ASAP7_75t_L g626 ( .A1(n_565), .A2(n_589), .A3(n_627), .B(n_632), .Y(n_626) );
INVx2_ASAP7_75t_SL g565 ( .A(n_566), .Y(n_565) );
INVx2_ASAP7_75t_SL g605 ( .A(n_566), .Y(n_605) );
INVx2_ASAP7_75t_L g569 ( .A(n_570), .Y(n_569) );
NAND2xp5_ASAP7_75t_L g732 ( .A(n_570), .B(n_733), .Y(n_732) );
NAND2x1_ASAP7_75t_L g737 ( .A(n_570), .B(n_738), .Y(n_737) );
AND2x2_ASAP7_75t_L g861 ( .A(n_570), .B(n_759), .Y(n_861) );
NAND2xp5_ASAP7_75t_L g865 ( .A(n_570), .B(n_815), .Y(n_865) );
AND2x2_ASAP7_75t_L g570 ( .A(n_571), .B(n_582), .Y(n_570) );
INVx4_ASAP7_75t_SL g620 ( .A(n_571), .Y(n_620) );
NAND2xp5_ASAP7_75t_L g669 ( .A(n_571), .B(n_622), .Y(n_669) );
BUFx2_ASAP7_75t_L g753 ( .A(n_571), .Y(n_753) );
NAND2xp5_ASAP7_75t_L g820 ( .A(n_571), .B(n_821), .Y(n_820) );
INVx1_ASAP7_75t_L g622 ( .A(n_582), .Y(n_622) );
INVx2_ASAP7_75t_L g657 ( .A(n_582), .Y(n_657) );
AND2x2_ASAP7_75t_L g659 ( .A(n_582), .B(n_617), .Y(n_659) );
INVx1_ASAP7_75t_L g684 ( .A(n_582), .Y(n_684) );
HB1xp67_ASAP7_75t_L g775 ( .A(n_582), .Y(n_775) );
NAND2xp5_ASAP7_75t_L g798 ( .A(n_582), .B(n_767), .Y(n_798) );
INVxp67_ASAP7_75t_L g592 ( .A(n_593), .Y(n_592) );
INVxp67_ASAP7_75t_SL g593 ( .A(n_594), .Y(n_593) );
AND2x2_ASAP7_75t_L g842 ( .A(n_594), .B(n_843), .Y(n_842) );
AND2x2_ASAP7_75t_L g594 ( .A(n_595), .B(n_607), .Y(n_594) );
AND2x4_ASAP7_75t_L g638 ( .A(n_595), .B(n_639), .Y(n_638) );
AND2x2_ASAP7_75t_L g699 ( .A(n_595), .B(n_643), .Y(n_699) );
INVx2_ASAP7_75t_L g595 ( .A(n_596), .Y(n_595) );
BUFx2_ASAP7_75t_L g785 ( .A(n_596), .Y(n_785) );
OAI21x1_ASAP7_75t_L g596 ( .A1(n_597), .A2(n_598), .B(n_606), .Y(n_596) );
OAI21x1_ASAP7_75t_L g672 ( .A1(n_597), .A2(n_598), .B(n_606), .Y(n_672) );
OAI21x1_ASAP7_75t_L g598 ( .A1(n_599), .A2(n_602), .B(n_605), .Y(n_598) );
AND2x4_ASAP7_75t_L g697 ( .A(n_607), .B(n_626), .Y(n_697) );
INVx3_ASAP7_75t_L g720 ( .A(n_607), .Y(n_720) );
INVx2_ASAP7_75t_L g741 ( .A(n_607), .Y(n_741) );
NAND2xp5_ASAP7_75t_L g829 ( .A(n_607), .B(n_830), .Y(n_829) );
NAND2xp5_ASAP7_75t_L g835 ( .A(n_607), .B(n_642), .Y(n_835) );
INVx3_ASAP7_75t_L g607 ( .A(n_608), .Y(n_607) );
AND2x2_ASAP7_75t_L g625 ( .A(n_608), .B(n_626), .Y(n_625) );
BUFx2_ASAP7_75t_L g637 ( .A(n_608), .Y(n_637) );
AND2x2_ASAP7_75t_L g714 ( .A(n_608), .B(n_639), .Y(n_714) );
INVx1_ASAP7_75t_L g614 ( .A(n_615), .Y(n_614) );
NAND2xp5_ASAP7_75t_L g615 ( .A(n_616), .B(n_619), .Y(n_615) );
AND2x2_ASAP7_75t_L g616 ( .A(n_617), .B(n_618), .Y(n_616) );
INVx3_ASAP7_75t_L g692 ( .A(n_617), .Y(n_692) );
AND2x2_ASAP7_75t_L g727 ( .A(n_617), .B(n_728), .Y(n_727) );
AND2x2_ASAP7_75t_L g796 ( .A(n_617), .B(n_620), .Y(n_796) );
NAND2xp5_ASAP7_75t_L g693 ( .A(n_618), .B(n_620), .Y(n_693) );
NAND2xp5_ASAP7_75t_SL g758 ( .A(n_619), .B(n_759), .Y(n_758) );
AND2x4_ASAP7_75t_L g619 ( .A(n_620), .B(n_621), .Y(n_619) );
INVx2_ASAP7_75t_L g655 ( .A(n_620), .Y(n_655) );
AND2x2_ASAP7_75t_L g683 ( .A(n_620), .B(n_684), .Y(n_683) );
OR2x2_ASAP7_75t_L g701 ( .A(n_620), .B(n_702), .Y(n_701) );
INVx1_ASAP7_75t_L g743 ( .A(n_620), .Y(n_743) );
NAND2xp5_ASAP7_75t_L g766 ( .A(n_620), .B(n_767), .Y(n_766) );
INVx1_ASAP7_75t_L g804 ( .A(n_620), .Y(n_804) );
INVx1_ASAP7_75t_L g621 ( .A(n_622), .Y(n_621) );
INVx2_ASAP7_75t_L g623 ( .A(n_624), .Y(n_623) );
INVx1_ASAP7_75t_SL g624 ( .A(n_625), .Y(n_624) );
NAND2xp5_ASAP7_75t_L g670 ( .A(n_625), .B(n_671), .Y(n_670) );
AND2x4_ASAP7_75t_SL g678 ( .A(n_625), .B(n_679), .Y(n_678) );
AND2x2_ASAP7_75t_L g757 ( .A(n_625), .B(n_641), .Y(n_757) );
HB1xp67_ASAP7_75t_L g792 ( .A(n_625), .Y(n_792) );
INVx2_ASAP7_75t_L g809 ( .A(n_625), .Y(n_809) );
INVx2_ASAP7_75t_L g639 ( .A(n_626), .Y(n_639) );
OR2x2_ASAP7_75t_L g689 ( .A(n_626), .B(n_680), .Y(n_689) );
INVx1_ASAP7_75t_L g710 ( .A(n_626), .Y(n_710) );
BUFx2_ASAP7_75t_L g725 ( .A(n_626), .Y(n_725) );
OR2x2_ASAP7_75t_L g794 ( .A(n_626), .B(n_644), .Y(n_794) );
AOI21xp5_ASAP7_75t_SL g634 ( .A1(n_635), .A2(n_640), .B(n_652), .Y(n_634) );
O2A1O1Ixp33_ASAP7_75t_L g760 ( .A1(n_635), .A2(n_716), .B(n_761), .C(n_764), .Y(n_760) );
INVx1_ASAP7_75t_L g635 ( .A(n_636), .Y(n_635) );
AND2x2_ASAP7_75t_L g660 ( .A(n_636), .B(n_661), .Y(n_660) );
AOI22xp5_ASAP7_75t_L g859 ( .A1(n_636), .A2(n_694), .B1(n_860), .B2(n_861), .Y(n_859) );
AND2x4_ASAP7_75t_L g636 ( .A(n_637), .B(n_638), .Y(n_636) );
INVx1_ASAP7_75t_L g651 ( .A(n_638), .Y(n_651) );
AND2x4_ASAP7_75t_L g779 ( .A(n_638), .B(n_688), .Y(n_779) );
NAND2xp5_ASAP7_75t_L g833 ( .A(n_638), .B(n_834), .Y(n_833) );
OR2x2_ASAP7_75t_L g640 ( .A(n_641), .B(n_651), .Y(n_640) );
INVx1_ASAP7_75t_L g661 ( .A(n_641), .Y(n_661) );
INVx1_ASAP7_75t_L g641 ( .A(n_642), .Y(n_641) );
AND2x4_ASAP7_75t_L g679 ( .A(n_642), .B(n_680), .Y(n_679) );
INVx2_ASAP7_75t_L g642 ( .A(n_643), .Y(n_642) );
NAND2xp5_ASAP7_75t_L g722 ( .A(n_643), .B(n_672), .Y(n_722) );
INVx2_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
AND2x2_ASAP7_75t_L g671 ( .A(n_644), .B(n_672), .Y(n_671) );
INVx1_ASAP7_75t_L g688 ( .A(n_644), .Y(n_688) );
HB1xp67_ASAP7_75t_L g763 ( .A(n_644), .Y(n_763) );
INVx2_ASAP7_75t_L g652 ( .A(n_653), .Y(n_652) );
AND2x4_ASAP7_75t_L g653 ( .A(n_654), .B(n_656), .Y(n_653) );
AND2x2_ASAP7_75t_L g674 ( .A(n_654), .B(n_675), .Y(n_674) );
INVx2_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
NAND2xp5_ASAP7_75t_L g773 ( .A(n_655), .B(n_734), .Y(n_773) );
INVx2_ASAP7_75t_L g665 ( .A(n_656), .Y(n_665) );
AND2x2_ASAP7_75t_L g742 ( .A(n_656), .B(n_743), .Y(n_742) );
NAND2x1p5_ASAP7_75t_L g787 ( .A(n_656), .B(n_706), .Y(n_787) );
AND2x2_ASAP7_75t_L g824 ( .A(n_656), .B(n_796), .Y(n_824) );
AOI21xp5_ASAP7_75t_L g658 ( .A1(n_659), .A2(n_660), .B(n_662), .Y(n_658) );
OAI22xp5_ASAP7_75t_L g662 ( .A1(n_663), .A2(n_670), .B1(n_673), .B2(n_677), .Y(n_662) );
NOR2x1_ASAP7_75t_L g663 ( .A(n_664), .B(n_666), .Y(n_663) );
INVx1_ASAP7_75t_L g664 ( .A(n_665), .Y(n_664) );
INVx1_ASAP7_75t_L g868 ( .A(n_665), .Y(n_868) );
INVx1_ASAP7_75t_L g666 ( .A(n_667), .Y(n_666) );
INVx1_ASAP7_75t_L g667 ( .A(n_668), .Y(n_667) );
INVx1_ASAP7_75t_L g668 ( .A(n_669), .Y(n_668) );
INVx1_ASAP7_75t_L g708 ( .A(n_671), .Y(n_708) );
AND2x2_ASAP7_75t_L g735 ( .A(n_671), .B(n_720), .Y(n_735) );
NAND2xp5_ASAP7_75t_L g805 ( .A(n_671), .B(n_714), .Y(n_805) );
AND2x4_ASAP7_75t_L g851 ( .A(n_671), .B(n_697), .Y(n_851) );
INVx1_ASAP7_75t_L g680 ( .A(n_672), .Y(n_680) );
INVx1_ASAP7_75t_L g673 ( .A(n_674), .Y(n_673) );
AND2x4_ASAP7_75t_L g857 ( .A(n_675), .B(n_753), .Y(n_857) );
INVx2_ASAP7_75t_L g675 ( .A(n_676), .Y(n_675) );
OR2x2_ASAP7_75t_L g790 ( .A(n_676), .B(n_791), .Y(n_790) );
OR2x2_ASAP7_75t_L g818 ( .A(n_676), .B(n_692), .Y(n_818) );
NAND2xp5_ASAP7_75t_L g849 ( .A(n_677), .B(n_850), .Y(n_849) );
INVx3_ASAP7_75t_L g677 ( .A(n_678), .Y(n_677) );
AND2x2_ASAP7_75t_L g799 ( .A(n_679), .B(n_800), .Y(n_799) );
AOI221xp5_ASAP7_75t_L g681 ( .A1(n_682), .A2(n_686), .B1(n_690), .B2(n_694), .C(n_700), .Y(n_681) );
AND2x2_ASAP7_75t_L g682 ( .A(n_683), .B(n_685), .Y(n_682) );
INVx1_ASAP7_75t_L g716 ( .A(n_683), .Y(n_716) );
AND2x2_ASAP7_75t_L g840 ( .A(n_683), .B(n_706), .Y(n_840) );
HB1xp67_ASAP7_75t_L g704 ( .A(n_684), .Y(n_704) );
INVx3_ASAP7_75t_L g702 ( .A(n_685), .Y(n_702) );
NAND2xp5_ASAP7_75t_L g751 ( .A(n_685), .B(n_752), .Y(n_751) );
AND2x4_ASAP7_75t_L g774 ( .A(n_685), .B(n_775), .Y(n_774) );
NOR2xp67_ASAP7_75t_SL g686 ( .A(n_687), .B(n_689), .Y(n_686) );
AND2x2_ASAP7_75t_L g713 ( .A(n_687), .B(n_714), .Y(n_713) );
NAND2xp5_ASAP7_75t_L g782 ( .A(n_687), .B(n_720), .Y(n_782) );
AOI322xp5_ASAP7_75t_L g788 ( .A1(n_687), .A2(n_774), .A3(n_789), .B1(n_792), .B2(n_793), .C1(n_795), .C2(n_799), .Y(n_788) );
INVx2_ASAP7_75t_L g687 ( .A(n_688), .Y(n_687) );
AND2x2_ASAP7_75t_L g730 ( .A(n_688), .B(n_697), .Y(n_730) );
NOR2xp33_ASAP7_75t_L g740 ( .A(n_689), .B(n_741), .Y(n_740) );
NOR2x1_ASAP7_75t_L g838 ( .A(n_689), .B(n_839), .Y(n_838) );
AOI22xp5_ASAP7_75t_L g831 ( .A1(n_690), .A2(n_832), .B1(n_836), .B2(n_840), .Y(n_831) );
INVx1_ASAP7_75t_L g690 ( .A(n_691), .Y(n_690) );
OR2x2_ASAP7_75t_L g691 ( .A(n_692), .B(n_693), .Y(n_691) );
INVx4_ASAP7_75t_L g815 ( .A(n_692), .Y(n_815) );
OR2x2_ASAP7_75t_L g845 ( .A(n_692), .B(n_820), .Y(n_845) );
INVx1_ASAP7_75t_L g694 ( .A(n_695), .Y(n_694) );
OR2x2_ASAP7_75t_L g695 ( .A(n_696), .B(n_698), .Y(n_695) );
INVx2_ASAP7_75t_SL g696 ( .A(n_697), .Y(n_696) );
INVx1_ASAP7_75t_L g858 ( .A(n_697), .Y(n_858) );
NOR2xp33_ASAP7_75t_L g745 ( .A(n_698), .B(n_724), .Y(n_745) );
INVx1_ASAP7_75t_L g698 ( .A(n_699), .Y(n_698) );
AOI211x1_ASAP7_75t_L g700 ( .A1(n_701), .A2(n_703), .B(n_708), .C(n_709), .Y(n_700) );
INVx2_ASAP7_75t_L g738 ( .A(n_702), .Y(n_738) );
NAND2xp5_ASAP7_75t_L g703 ( .A(n_704), .B(n_705), .Y(n_703) );
INVx1_ASAP7_75t_L g705 ( .A(n_706), .Y(n_705) );
INVx2_ASAP7_75t_L g765 ( .A(n_706), .Y(n_765) );
NAND2x1_ASAP7_75t_L g856 ( .A(n_706), .B(n_857), .Y(n_856) );
INVx3_ASAP7_75t_L g706 ( .A(n_707), .Y(n_706) );
AND2x2_ASAP7_75t_L g762 ( .A(n_707), .B(n_763), .Y(n_762) );
INVx1_ASAP7_75t_L g827 ( .A(n_709), .Y(n_827) );
BUFx2_ASAP7_75t_L g709 ( .A(n_710), .Y(n_709) );
NAND3xp33_ASAP7_75t_L g711 ( .A(n_712), .B(n_729), .C(n_744), .Y(n_711) );
OAI211xp5_ASAP7_75t_L g712 ( .A1(n_713), .A2(n_715), .B(n_717), .C(n_727), .Y(n_712) );
INVx1_ASAP7_75t_L g726 ( .A(n_713), .Y(n_726) );
NAND2xp5_ASAP7_75t_L g754 ( .A(n_714), .B(n_755), .Y(n_754) );
AND2x2_ASAP7_75t_L g784 ( .A(n_714), .B(n_785), .Y(n_784) );
NAND2xp33_ASAP7_75t_L g807 ( .A(n_714), .B(n_755), .Y(n_807) );
HB1xp67_ASAP7_75t_L g715 ( .A(n_716), .Y(n_715) );
NAND2xp5_ASAP7_75t_L g717 ( .A(n_718), .B(n_726), .Y(n_717) );
INVx1_ASAP7_75t_L g853 ( .A(n_718), .Y(n_853) );
NAND2x1p5_ASAP7_75t_L g718 ( .A(n_719), .B(n_723), .Y(n_718) );
AND2x4_ASAP7_75t_L g719 ( .A(n_720), .B(n_721), .Y(n_719) );
INVx2_ASAP7_75t_L g800 ( .A(n_720), .Y(n_800) );
INVx1_ASAP7_75t_L g721 ( .A(n_722), .Y(n_721) );
INVx1_ASAP7_75t_L g755 ( .A(n_722), .Y(n_755) );
INVxp67_ASAP7_75t_SL g830 ( .A(n_722), .Y(n_830) );
INVx1_ASAP7_75t_L g723 ( .A(n_724), .Y(n_723) );
INVx1_ASAP7_75t_L g724 ( .A(n_725), .Y(n_724) );
INVx1_ASAP7_75t_L g759 ( .A(n_728), .Y(n_759) );
AOI221xp5_ASAP7_75t_L g729 ( .A1(n_730), .A2(n_731), .B1(n_735), .B2(n_736), .C(n_739), .Y(n_729) );
INVxp67_ASAP7_75t_SL g731 ( .A(n_732), .Y(n_731) );
HB1xp67_ASAP7_75t_L g733 ( .A(n_734), .Y(n_733) );
INVx1_ASAP7_75t_L g791 ( .A(n_734), .Y(n_791) );
INVx1_ASAP7_75t_L g736 ( .A(n_737), .Y(n_736) );
AND2x2_ASAP7_75t_L g739 ( .A(n_740), .B(n_742), .Y(n_739) );
INVx1_ASAP7_75t_L g777 ( .A(n_741), .Y(n_777) );
NOR2x1p5_ASAP7_75t_L g793 ( .A(n_741), .B(n_794), .Y(n_793) );
AOI21xp5_ASAP7_75t_L g780 ( .A1(n_742), .A2(n_781), .B(n_783), .Y(n_780) );
INVx1_ASAP7_75t_L g749 ( .A(n_743), .Y(n_749) );
AOI211xp5_ASAP7_75t_L g744 ( .A1(n_745), .A2(n_746), .B(n_750), .C(n_760), .Y(n_744) );
INVx1_ASAP7_75t_L g746 ( .A(n_747), .Y(n_746) );
INVx1_ASAP7_75t_L g747 ( .A(n_748), .Y(n_747) );
OAI22xp5_ASAP7_75t_L g750 ( .A1(n_751), .A2(n_754), .B1(n_756), .B2(n_758), .Y(n_750) );
INVx1_ASAP7_75t_L g752 ( .A(n_753), .Y(n_752) );
INVx1_ASAP7_75t_L g756 ( .A(n_757), .Y(n_756) );
INVx1_ASAP7_75t_L g761 ( .A(n_762), .Y(n_761) );
INVx1_ASAP7_75t_L g839 ( .A(n_763), .Y(n_839) );
OR2x2_ASAP7_75t_L g764 ( .A(n_765), .B(n_766), .Y(n_764) );
NOR3xp33_ASAP7_75t_L g768 ( .A(n_769), .B(n_801), .C(n_822), .Y(n_768) );
NAND3xp33_ASAP7_75t_SL g769 ( .A(n_770), .B(n_780), .C(n_788), .Y(n_769) );
OAI21xp33_ASAP7_75t_L g770 ( .A1(n_771), .A2(n_774), .B(n_776), .Y(n_770) );
INVxp67_ASAP7_75t_SL g771 ( .A(n_772), .Y(n_771) );
HB1xp67_ASAP7_75t_L g772 ( .A(n_773), .Y(n_772) );
NOR2xp33_ASAP7_75t_L g776 ( .A(n_777), .B(n_778), .Y(n_776) );
AND2x2_ASAP7_75t_L g870 ( .A(n_777), .B(n_838), .Y(n_870) );
INVx2_ASAP7_75t_L g778 ( .A(n_779), .Y(n_778) );
OAI21xp5_ASAP7_75t_L g816 ( .A1(n_779), .A2(n_817), .B(n_819), .Y(n_816) );
INVxp67_ASAP7_75t_SL g781 ( .A(n_782), .Y(n_781) );
AND2x2_ASAP7_75t_L g783 ( .A(n_784), .B(n_786), .Y(n_783) );
OR2x2_ASAP7_75t_L g808 ( .A(n_785), .B(n_809), .Y(n_808) );
INVx2_ASAP7_75t_L g786 ( .A(n_787), .Y(n_786) );
INVx2_ASAP7_75t_L g789 ( .A(n_790), .Y(n_789) );
INVx1_ASAP7_75t_L g843 ( .A(n_794), .Y(n_843) );
AND2x2_ASAP7_75t_L g795 ( .A(n_796), .B(n_797), .Y(n_795) );
HB1xp67_ASAP7_75t_L g860 ( .A(n_797), .Y(n_860) );
INVx1_ASAP7_75t_L g797 ( .A(n_798), .Y(n_797) );
OR2x2_ASAP7_75t_L g803 ( .A(n_798), .B(n_804), .Y(n_803) );
INVx1_ASAP7_75t_L g813 ( .A(n_798), .Y(n_813) );
OAI221xp5_ASAP7_75t_L g801 ( .A1(n_802), .A2(n_805), .B1(n_806), .B2(n_810), .C(n_816), .Y(n_801) );
OAI21xp5_ASAP7_75t_L g847 ( .A1(n_802), .A2(n_848), .B(n_852), .Y(n_847) );
BUFx2_ASAP7_75t_L g802 ( .A(n_803), .Y(n_802) );
AOI32xp33_ASAP7_75t_L g841 ( .A1(n_804), .A2(n_815), .A3(n_842), .B1(n_843), .B2(n_844), .Y(n_841) );
AND2x2_ASAP7_75t_SL g806 ( .A(n_807), .B(n_808), .Y(n_806) );
INVx1_ASAP7_75t_L g810 ( .A(n_811), .Y(n_810) );
INVx1_ASAP7_75t_L g811 ( .A(n_812), .Y(n_811) );
NAND2xp5_ASAP7_75t_L g812 ( .A(n_813), .B(n_814), .Y(n_812) );
INVx1_ASAP7_75t_L g814 ( .A(n_815), .Y(n_814) );
NAND2xp5_ASAP7_75t_L g852 ( .A(n_817), .B(n_853), .Y(n_852) );
INVx1_ASAP7_75t_L g817 ( .A(n_818), .Y(n_817) );
INVx1_ASAP7_75t_L g819 ( .A(n_820), .Y(n_819) );
OAI211xp5_ASAP7_75t_SL g822 ( .A1(n_823), .A2(n_825), .B(n_831), .C(n_841), .Y(n_822) );
INVx2_ASAP7_75t_L g823 ( .A(n_824), .Y(n_823) );
INVx1_ASAP7_75t_L g825 ( .A(n_826), .Y(n_825) );
AND2x4_ASAP7_75t_L g826 ( .A(n_827), .B(n_828), .Y(n_826) );
INVx1_ASAP7_75t_L g828 ( .A(n_829), .Y(n_828) );
INVx1_ASAP7_75t_L g832 ( .A(n_833), .Y(n_832) );
INVx1_ASAP7_75t_L g834 ( .A(n_835), .Y(n_834) );
INVx1_ASAP7_75t_L g836 ( .A(n_837), .Y(n_836) );
INVx1_ASAP7_75t_L g837 ( .A(n_838), .Y(n_837) );
INVx1_ASAP7_75t_L g844 ( .A(n_845), .Y(n_844) );
NOR3xp33_ASAP7_75t_L g846 ( .A(n_847), .B(n_854), .C(n_862), .Y(n_846) );
INVxp33_ASAP7_75t_L g848 ( .A(n_849), .Y(n_848) );
INVx1_ASAP7_75t_L g850 ( .A(n_851), .Y(n_850) );
OAI21xp33_ASAP7_75t_SL g854 ( .A1(n_855), .A2(n_858), .B(n_859), .Y(n_854) );
HB1xp67_ASAP7_75t_L g855 ( .A(n_856), .Y(n_855) );
AOI21xp5_ASAP7_75t_L g862 ( .A1(n_863), .A2(n_866), .B(n_869), .Y(n_862) );
INVxp67_ASAP7_75t_L g863 ( .A(n_864), .Y(n_863) );
INVx1_ASAP7_75t_L g864 ( .A(n_865), .Y(n_864) );
NOR2xp33_ASAP7_75t_SL g866 ( .A(n_867), .B(n_868), .Y(n_866) );
INVx2_ASAP7_75t_L g869 ( .A(n_870), .Y(n_869) );
BUFx4f_ASAP7_75t_SL g873 ( .A(n_874), .Y(n_873) );
OR2x2_ASAP7_75t_L g874 ( .A(n_875), .B(n_878), .Y(n_874) );
BUFx2_ASAP7_75t_L g875 ( .A(n_876), .Y(n_875) );
OR2x2_ASAP7_75t_L g878 ( .A(n_879), .B(n_880), .Y(n_878) );
AND2x2_ASAP7_75t_L g883 ( .A(n_879), .B(n_884), .Y(n_883) );
NOR2xp33_ASAP7_75t_L g884 ( .A(n_880), .B(n_885), .Y(n_884) );
INVx3_ASAP7_75t_L g885 ( .A(n_886), .Y(n_885) );
BUFx3_ASAP7_75t_L g887 ( .A(n_888), .Y(n_887) );
OR2x4_ASAP7_75t_L g888 ( .A(n_889), .B(n_891), .Y(n_888) );
BUFx2_ASAP7_75t_L g889 ( .A(n_890), .Y(n_889) );
endmodule