module fake_jpeg_20450_n_308 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_308);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_308;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_208;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_14),
.Y(n_19)
);

INVx3_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_3),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_16),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_13),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_4),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_9),
.Y(n_31)
);

INVx11_ASAP7_75t_L g32 ( 
.A(n_8),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_15),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_9),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_SL g35 ( 
.A(n_19),
.B(n_7),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_35),
.B(n_36),
.Y(n_53)
);

CKINVDCx16_ASAP7_75t_R g36 ( 
.A(n_23),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_27),
.Y(n_37)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_37),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_27),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_38),
.Y(n_57)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_27),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_39),
.Y(n_52)
);

INVx5_ASAP7_75t_L g40 ( 
.A(n_21),
.Y(n_40)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_40),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_21),
.B(n_16),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_41),
.B(n_30),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_23),
.Y(n_42)
);

OA22x2_ASAP7_75t_L g61 ( 
.A1(n_42),
.A2(n_19),
.B1(n_33),
.B2(n_31),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_27),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_43),
.Y(n_60)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_40),
.Y(n_44)
);

INVx5_ASAP7_75t_L g84 ( 
.A(n_44),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_L g45 ( 
.A1(n_41),
.A2(n_20),
.B1(n_34),
.B2(n_23),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_45),
.A2(n_54),
.B1(n_25),
.B2(n_34),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g46 ( 
.A(n_41),
.B(n_26),
.C(n_21),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_46),
.B(n_62),
.Y(n_67)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_38),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_49),
.Y(n_86)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_40),
.Y(n_50)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_50),
.Y(n_69)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_38),
.Y(n_51)
);

INVx6_ASAP7_75t_L g75 ( 
.A(n_51),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g54 ( 
.A1(n_37),
.A2(n_39),
.B1(n_42),
.B2(n_36),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_40),
.A2(n_32),
.B1(n_20),
.B2(n_29),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_55),
.A2(n_32),
.B1(n_20),
.B2(n_25),
.Y(n_83)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_38),
.Y(n_56)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_56),
.Y(n_90)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_38),
.Y(n_58)
);

INVx6_ASAP7_75t_L g92 ( 
.A(n_58),
.Y(n_92)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_40),
.Y(n_59)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_59),
.Y(n_76)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_61),
.Y(n_94)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_43),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_63),
.B(n_64),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_35),
.B(n_33),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_35),
.B(n_31),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_65),
.B(n_30),
.Y(n_71)
);

INVx13_ASAP7_75t_L g66 ( 
.A(n_60),
.Y(n_66)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_66),
.Y(n_112)
);

INVx5_ASAP7_75t_L g70 ( 
.A(n_44),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_70),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_SL g109 ( 
.A(n_71),
.B(n_72),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_53),
.B(n_42),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_52),
.A2(n_39),
.B1(n_37),
.B2(n_42),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_73),
.A2(n_74),
.B1(n_56),
.B2(n_49),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_52),
.A2(n_46),
.B1(n_39),
.B2(n_37),
.Y(n_74)
);

INVx11_ASAP7_75t_L g77 ( 
.A(n_60),
.Y(n_77)
);

INVx4_ASAP7_75t_SL g102 ( 
.A(n_77),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_61),
.B(n_36),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_SL g113 ( 
.A(n_78),
.B(n_81),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_61),
.B(n_43),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_79),
.B(n_91),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_61),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_80),
.B(n_85),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_54),
.B(n_22),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_82),
.B(n_24),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_83),
.A2(n_32),
.B1(n_34),
.B2(n_17),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_50),
.B(n_22),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_59),
.B(n_28),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_87),
.B(n_88),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_48),
.B(n_28),
.Y(n_88)
);

HB1xp67_ASAP7_75t_L g89 ( 
.A(n_47),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_89),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_48),
.B(n_43),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_47),
.B(n_29),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_93),
.B(n_26),
.Y(n_114)
);

AOI21xp5_ASAP7_75t_L g95 ( 
.A1(n_67),
.A2(n_62),
.B(n_58),
.Y(n_95)
);

OAI21xp5_ASAP7_75t_SL g150 ( 
.A1(n_95),
.A2(n_106),
.B(n_118),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_94),
.A2(n_80),
.B1(n_78),
.B2(n_72),
.Y(n_96)
);

OAI21xp5_ASAP7_75t_L g138 ( 
.A1(n_96),
.A2(n_116),
.B(n_68),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_L g98 ( 
.A(n_67),
.B(n_17),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_98),
.B(n_119),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_99),
.A2(n_103),
.B1(n_107),
.B2(n_108),
.Y(n_134)
);

OAI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_94),
.A2(n_51),
.B1(n_25),
.B2(n_29),
.Y(n_103)
);

OAI22x1_ASAP7_75t_L g140 ( 
.A1(n_104),
.A2(n_66),
.B1(n_77),
.B2(n_26),
.Y(n_140)
);

INVxp67_ASAP7_75t_L g105 ( 
.A(n_93),
.Y(n_105)
);

CKINVDCx16_ASAP7_75t_R g127 ( 
.A(n_105),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_SL g106 ( 
.A1(n_79),
.A2(n_26),
.B(n_21),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_81),
.A2(n_43),
.B1(n_57),
.B2(n_60),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_91),
.A2(n_57),
.B1(n_60),
.B2(n_24),
.Y(n_108)
);

OAI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_74),
.A2(n_24),
.B1(n_18),
.B2(n_21),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_110),
.A2(n_117),
.B1(n_92),
.B2(n_75),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_114),
.B(n_86),
.Y(n_132)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_69),
.Y(n_115)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_115),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_82),
.A2(n_92),
.B1(n_75),
.B2(n_88),
.Y(n_116)
);

AND2x2_ASAP7_75t_L g118 ( 
.A(n_73),
.B(n_26),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_90),
.Y(n_119)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_85),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_120),
.B(n_100),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_SL g124 ( 
.A(n_109),
.B(n_68),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_SL g161 ( 
.A(n_124),
.B(n_147),
.Y(n_161)
);

INVx5_ASAP7_75t_L g125 ( 
.A(n_121),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_125),
.B(n_131),
.Y(n_176)
);

CKINVDCx14_ASAP7_75t_R g182 ( 
.A(n_126),
.Y(n_182)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_121),
.Y(n_128)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_128),
.Y(n_159)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_121),
.Y(n_129)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_129),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_101),
.A2(n_92),
.B1(n_75),
.B2(n_90),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_130),
.A2(n_148),
.B1(n_18),
.B2(n_1),
.Y(n_175)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_115),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_132),
.B(n_133),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_101),
.B(n_87),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_135),
.A2(n_117),
.B1(n_107),
.B2(n_111),
.Y(n_167)
);

INVx3_ASAP7_75t_L g136 ( 
.A(n_111),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_136),
.B(n_149),
.Y(n_178)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_99),
.Y(n_137)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_137),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_L g181 ( 
.A1(n_138),
.A2(n_18),
.B(n_9),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_97),
.B(n_86),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_139),
.B(n_145),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_SL g155 ( 
.A1(n_140),
.A2(n_118),
.B(n_119),
.Y(n_155)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_108),
.Y(n_141)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_141),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_112),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_142),
.B(n_146),
.Y(n_153)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_95),
.Y(n_143)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_143),
.Y(n_183)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_112),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_144),
.B(n_151),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_97),
.B(n_86),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_109),
.B(n_71),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_SL g147 ( 
.A(n_100),
.B(n_69),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_96),
.A2(n_76),
.B1(n_84),
.B2(n_70),
.Y(n_148)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_115),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_98),
.B(n_76),
.Y(n_151)
);

OA21x2_ASAP7_75t_L g152 ( 
.A1(n_143),
.A2(n_116),
.B(n_118),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_152),
.B(n_158),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_139),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_154),
.B(n_160),
.Y(n_209)
);

OAI21xp5_ASAP7_75t_SL g188 ( 
.A1(n_155),
.A2(n_156),
.B(n_166),
.Y(n_188)
);

AOI21xp5_ASAP7_75t_L g156 ( 
.A1(n_150),
.A2(n_138),
.B(n_148),
.Y(n_156)
);

OA21x2_ASAP7_75t_L g158 ( 
.A1(n_137),
.A2(n_118),
.B(n_110),
.Y(n_158)
);

INVxp67_ASAP7_75t_L g160 ( 
.A(n_130),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_145),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_162),
.B(n_171),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g164 ( 
.A(n_151),
.B(n_106),
.Y(n_164)
);

XOR2xp5_ASAP7_75t_L g186 ( 
.A(n_164),
.B(n_134),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_SL g166 ( 
.A1(n_150),
.A2(n_113),
.B(n_114),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_167),
.A2(n_170),
.B1(n_149),
.B2(n_131),
.Y(n_198)
);

AOI21xp5_ASAP7_75t_L g168 ( 
.A1(n_140),
.A2(n_113),
.B(n_102),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_SL g196 ( 
.A1(n_168),
.A2(n_174),
.B(n_136),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_142),
.B(n_102),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_169),
.B(n_172),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_141),
.A2(n_102),
.B1(n_84),
.B2(n_70),
.Y(n_170)
);

CKINVDCx16_ASAP7_75t_R g171 ( 
.A(n_144),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_133),
.B(n_132),
.Y(n_172)
);

A2O1A1O1Ixp25_ASAP7_75t_L g174 ( 
.A1(n_123),
.A2(n_24),
.B(n_18),
.C(n_77),
.D(n_66),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_175),
.A2(n_135),
.B1(n_129),
.B2(n_125),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_128),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_SL g189 ( 
.A(n_177),
.B(n_161),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_L g203 ( 
.A1(n_181),
.A2(n_168),
.B(n_156),
.Y(n_203)
);

AOI21xp5_ASAP7_75t_L g185 ( 
.A1(n_155),
.A2(n_127),
.B(n_134),
.Y(n_185)
);

INVxp67_ASAP7_75t_L g219 ( 
.A(n_185),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_SL g218 ( 
.A(n_186),
.B(n_204),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_187),
.A2(n_170),
.B1(n_179),
.B2(n_180),
.Y(n_215)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_189),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g190 ( 
.A(n_164),
.B(n_166),
.Y(n_190)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_190),
.B(n_210),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_153),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_193),
.B(n_195),
.Y(n_214)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_178),
.Y(n_194)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_194),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_153),
.Y(n_195)
);

AOI21xp5_ASAP7_75t_L g230 ( 
.A1(n_196),
.A2(n_207),
.B(n_174),
.Y(n_230)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_169),
.Y(n_197)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_197),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_L g233 ( 
.A1(n_198),
.A2(n_205),
.B1(n_158),
.B2(n_171),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_172),
.B(n_122),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_199),
.B(n_200),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_SL g200 ( 
.A(n_161),
.B(n_122),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_165),
.Y(n_201)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_201),
.Y(n_232)
);

AOI21xp5_ASAP7_75t_L g202 ( 
.A1(n_183),
.A2(n_0),
.B(n_1),
.Y(n_202)
);

INVxp67_ASAP7_75t_L g224 ( 
.A(n_202),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_203),
.A2(n_154),
.B1(n_162),
.B2(n_152),
.Y(n_213)
);

AOI322xp5_ASAP7_75t_L g204 ( 
.A1(n_181),
.A2(n_7),
.A3(n_15),
.B1(n_2),
.B2(n_3),
.C1(n_4),
.C2(n_5),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_167),
.A2(n_10),
.B1(n_15),
.B2(n_3),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_157),
.B(n_10),
.C(n_14),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_206),
.B(n_182),
.C(n_152),
.Y(n_220)
);

A2O1A1Ixp33_ASAP7_75t_L g207 ( 
.A1(n_157),
.A2(n_10),
.B(n_14),
.C(n_4),
.Y(n_207)
);

AOI21xp5_ASAP7_75t_L g208 ( 
.A1(n_183),
.A2(n_0),
.B(n_1),
.Y(n_208)
);

INVxp67_ASAP7_75t_L g227 ( 
.A(n_208),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g210 ( 
.A(n_163),
.B(n_5),
.Y(n_210)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_213),
.B(n_231),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_L g237 ( 
.A1(n_215),
.A2(n_222),
.B1(n_226),
.B2(n_230),
.Y(n_237)
);

BUFx6f_ASAP7_75t_L g216 ( 
.A(n_193),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_216),
.B(n_220),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_187),
.A2(n_179),
.B1(n_180),
.B2(n_165),
.Y(n_222)
);

NOR2x1_ASAP7_75t_L g223 ( 
.A(n_189),
.B(n_195),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_223),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_190),
.B(n_163),
.C(n_152),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_225),
.B(n_188),
.C(n_196),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_191),
.A2(n_158),
.B1(n_177),
.B2(n_175),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_184),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_228),
.B(n_200),
.Y(n_238)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_188),
.B(n_158),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_233),
.A2(n_197),
.B1(n_209),
.B2(n_191),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_SL g234 ( 
.A(n_186),
.B(n_203),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_SL g248 ( 
.A(n_234),
.B(n_210),
.Y(n_248)
);

BUFx12_ASAP7_75t_L g236 ( 
.A(n_216),
.Y(n_236)
);

HB1xp67_ASAP7_75t_L g265 ( 
.A(n_236),
.Y(n_265)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_238),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_SL g239 ( 
.A(n_211),
.B(n_206),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_239),
.B(n_240),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_214),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_217),
.B(n_192),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_241),
.B(n_242),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_229),
.B(n_192),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_243),
.B(n_244),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_221),
.B(n_185),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_245),
.B(n_252),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_L g246 ( 
.A1(n_224),
.A2(n_205),
.B1(n_198),
.B2(n_209),
.Y(n_246)
);

BUFx2_ASAP7_75t_L g256 ( 
.A(n_246),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_225),
.B(n_199),
.C(n_201),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_247),
.B(n_220),
.C(n_234),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_248),
.B(n_253),
.Y(n_260)
);

AOI21xp5_ASAP7_75t_L g249 ( 
.A1(n_219),
.A2(n_194),
.B(n_207),
.Y(n_249)
);

OAI21xp5_ASAP7_75t_SL g254 ( 
.A1(n_249),
.A2(n_224),
.B(n_227),
.Y(n_254)
);

HB1xp67_ASAP7_75t_L g252 ( 
.A(n_213),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_232),
.B(n_208),
.Y(n_253)
);

MAJx2_ASAP7_75t_L g276 ( 
.A(n_254),
.B(n_249),
.C(n_250),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_SL g274 ( 
.A(n_261),
.B(n_259),
.Y(n_274)
);

AOI22xp33_ASAP7_75t_SL g262 ( 
.A1(n_235),
.A2(n_212),
.B1(n_219),
.B2(n_227),
.Y(n_262)
);

INVxp67_ASAP7_75t_L g270 ( 
.A(n_262),
.Y(n_270)
);

FAx1_ASAP7_75t_SL g263 ( 
.A(n_248),
.B(n_223),
.CI(n_221),
.CON(n_263),
.SN(n_263)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_263),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_247),
.B(n_218),
.C(n_231),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_266),
.B(n_268),
.Y(n_281)
);

OAI21xp5_ASAP7_75t_SL g267 ( 
.A1(n_251),
.A2(n_202),
.B(n_226),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_267),
.B(n_245),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_243),
.B(n_218),
.C(n_222),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_268),
.B(n_244),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_SL g283 ( 
.A(n_269),
.B(n_274),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_255),
.B(n_236),
.Y(n_271)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_271),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_258),
.B(n_236),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_273),
.B(n_176),
.Y(n_287)
);

XOR2xp5_ASAP7_75t_L g275 ( 
.A(n_266),
.B(n_250),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_275),
.B(n_277),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_276),
.A2(n_262),
.B1(n_260),
.B2(n_259),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_264),
.A2(n_237),
.B1(n_241),
.B2(n_253),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_SL g278 ( 
.A(n_260),
.B(n_261),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_SL g291 ( 
.A(n_278),
.B(n_173),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_279),
.B(n_280),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_263),
.A2(n_173),
.B1(n_159),
.B2(n_242),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_272),
.B(n_257),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_284),
.B(n_285),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_281),
.B(n_256),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_287),
.B(n_288),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_270),
.B(n_256),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_L g297 ( 
.A1(n_290),
.A2(n_0),
.B1(n_6),
.B2(n_11),
.Y(n_297)
);

OAI21xp5_ASAP7_75t_L g294 ( 
.A1(n_291),
.A2(n_278),
.B(n_265),
.Y(n_294)
);

OAI21xp33_ASAP7_75t_L g293 ( 
.A1(n_286),
.A2(n_276),
.B(n_270),
.Y(n_293)
);

AOI322xp5_ASAP7_75t_L g301 ( 
.A1(n_293),
.A2(n_294),
.A3(n_0),
.B1(n_6),
.B2(n_12),
.C1(n_16),
.C2(n_296),
.Y(n_301)
);

OAI21xp5_ASAP7_75t_SL g295 ( 
.A1(n_283),
.A2(n_159),
.B(n_5),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_SL g300 ( 
.A(n_295),
.B(n_298),
.Y(n_300)
);

AND2x2_ASAP7_75t_L g302 ( 
.A(n_297),
.B(n_12),
.Y(n_302)
);

OAI21xp5_ASAP7_75t_SL g298 ( 
.A1(n_282),
.A2(n_6),
.B(n_11),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_L g299 ( 
.A1(n_292),
.A2(n_289),
.B1(n_287),
.B2(n_290),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_SL g304 ( 
.A1(n_299),
.A2(n_301),
.B1(n_302),
.B2(n_300),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_SL g303 ( 
.A(n_293),
.B(n_12),
.Y(n_303)
);

HB1xp67_ASAP7_75t_L g305 ( 
.A(n_303),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_304),
.Y(n_306)
);

HB1xp67_ASAP7_75t_L g307 ( 
.A(n_306),
.Y(n_307)
);

XOR2xp5_ASAP7_75t_L g308 ( 
.A(n_307),
.B(n_305),
.Y(n_308)
);


endmodule