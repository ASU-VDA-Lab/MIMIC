module fake_jpeg_12592_n_275 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_275);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_275;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_272;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_125;
wire n_80;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_140;
wire n_82;
wire n_128;
wire n_100;
wire n_258;
wire n_96;

INVxp67_ASAP7_75t_L g15 ( 
.A(n_2),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_13),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_8),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_11),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_14),
.Y(n_22)
);

INVx1_ASAP7_75t_SL g23 ( 
.A(n_3),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_7),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_2),
.Y(n_26)
);

INVx1_ASAP7_75t_SL g27 ( 
.A(n_6),
.Y(n_27)
);

BUFx16f_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_2),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_6),
.Y(n_31)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_5),
.Y(n_33)
);

BUFx2_ASAP7_75t_L g34 ( 
.A(n_9),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_14),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_6),
.Y(n_36)
);

BUFx5_ASAP7_75t_L g37 ( 
.A(n_10),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_16),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_38),
.B(n_46),
.Y(n_63)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_30),
.Y(n_39)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_39),
.Y(n_69)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_28),
.Y(n_40)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_40),
.Y(n_67)
);

INVx11_ASAP7_75t_L g41 ( 
.A(n_28),
.Y(n_41)
);

CKINVDCx16_ASAP7_75t_R g79 ( 
.A(n_41),
.Y(n_79)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_21),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_42),
.Y(n_80)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_28),
.Y(n_43)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_43),
.Y(n_85)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_32),
.Y(n_44)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_44),
.Y(n_61)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_20),
.Y(n_45)
);

INVx5_ASAP7_75t_L g68 ( 
.A(n_45),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_16),
.Y(n_46)
);

INVx11_ASAP7_75t_L g47 ( 
.A(n_28),
.Y(n_47)
);

INVx1_ASAP7_75t_SL g81 ( 
.A(n_47),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_27),
.B(n_23),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_48),
.B(n_52),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_21),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_49),
.Y(n_97)
);

INVx11_ASAP7_75t_L g50 ( 
.A(n_20),
.Y(n_50)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_50),
.Y(n_64)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_21),
.Y(n_51)
);

INVx8_ASAP7_75t_L g72 ( 
.A(n_51),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_18),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_18),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_53),
.B(n_54),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_27),
.B(n_1),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_22),
.Y(n_55)
);

INVx8_ASAP7_75t_L g73 ( 
.A(n_55),
.Y(n_73)
);

BUFx5_ASAP7_75t_L g56 ( 
.A(n_37),
.Y(n_56)
);

BUFx12f_ASAP7_75t_L g65 ( 
.A(n_56),
.Y(n_65)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_37),
.Y(n_57)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_57),
.Y(n_92)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_32),
.Y(n_58)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_58),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_23),
.B(n_1),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_SL g66 ( 
.A(n_59),
.B(n_15),
.Y(n_66)
);

BUFx5_ASAP7_75t_L g60 ( 
.A(n_22),
.Y(n_60)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_60),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_66),
.B(n_88),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_54),
.A2(n_25),
.B1(n_22),
.B2(n_34),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_70),
.A2(n_103),
.B1(n_33),
.B2(n_19),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_L g71 ( 
.A1(n_42),
.A2(n_34),
.B1(n_23),
.B2(n_32),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_71),
.A2(n_82),
.B1(n_49),
.B2(n_56),
.Y(n_125)
);

AND2x2_ASAP7_75t_L g74 ( 
.A(n_48),
.B(n_25),
.Y(n_74)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_74),
.B(n_75),
.Y(n_106)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_59),
.B(n_34),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_39),
.Y(n_76)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_76),
.Y(n_110)
);

AND2x2_ASAP7_75t_SL g77 ( 
.A(n_44),
.B(n_40),
.Y(n_77)
);

AND2x2_ASAP7_75t_L g115 ( 
.A(n_77),
.B(n_57),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_45),
.A2(n_19),
.B1(n_33),
.B2(n_36),
.Y(n_82)
);

INVx5_ASAP7_75t_L g83 ( 
.A(n_57),
.Y(n_83)
);

INVx4_ASAP7_75t_L g111 ( 
.A(n_83),
.Y(n_111)
);

CKINVDCx12_ASAP7_75t_R g84 ( 
.A(n_41),
.Y(n_84)
);

OR2x2_ASAP7_75t_L g123 ( 
.A(n_84),
.B(n_99),
.Y(n_123)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_43),
.Y(n_87)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_87),
.Y(n_112)
);

OR2x2_ASAP7_75t_L g88 ( 
.A(n_38),
.B(n_30),
.Y(n_88)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_58),
.Y(n_89)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_89),
.Y(n_135)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_47),
.Y(n_90)
);

INVx4_ASAP7_75t_L g131 ( 
.A(n_90),
.Y(n_131)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_58),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_91),
.B(n_93),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_SL g93 ( 
.A(n_46),
.B(n_35),
.Y(n_93)
);

OA22x2_ASAP7_75t_L g94 ( 
.A1(n_55),
.A2(n_29),
.B1(n_24),
.B2(n_26),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_94),
.B(n_17),
.C(n_26),
.Y(n_113)
);

BUFx2_ASAP7_75t_L g95 ( 
.A(n_45),
.Y(n_95)
);

BUFx3_ASAP7_75t_L g104 ( 
.A(n_95),
.Y(n_104)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_42),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_96),
.B(n_49),
.Y(n_126)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_51),
.Y(n_98)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_98),
.Y(n_120)
);

OR2x2_ASAP7_75t_SL g99 ( 
.A(n_52),
.B(n_53),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_51),
.B(n_35),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_101),
.B(n_17),
.Y(n_108)
);

BUFx12_ASAP7_75t_L g102 ( 
.A(n_50),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g118 ( 
.A(n_102),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_55),
.A2(n_19),
.B1(n_33),
.B2(n_31),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_63),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_105),
.B(n_109),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_62),
.B(n_86),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_107),
.B(n_122),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_108),
.B(n_119),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_88),
.Y(n_109)
);

AND2x2_ASAP7_75t_L g153 ( 
.A(n_113),
.B(n_115),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g158 ( 
.A1(n_117),
.A2(n_129),
.B1(n_73),
.B2(n_97),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_86),
.B(n_31),
.Y(n_119)
);

OR2x2_ASAP7_75t_SL g121 ( 
.A(n_74),
.B(n_57),
.Y(n_121)
);

OR2x2_ASAP7_75t_L g145 ( 
.A(n_121),
.B(n_92),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_69),
.B(n_36),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_75),
.B(n_29),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_124),
.B(n_132),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_125),
.A2(n_136),
.B1(n_92),
.B2(n_73),
.Y(n_156)
);

INVxp67_ASAP7_75t_L g154 ( 
.A(n_126),
.Y(n_154)
);

AOI22xp33_ASAP7_75t_SL g127 ( 
.A1(n_95),
.A2(n_24),
.B1(n_60),
.B2(n_4),
.Y(n_127)
);

CKINVDCx16_ASAP7_75t_R g162 ( 
.A(n_127),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_94),
.B(n_1),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_128),
.B(n_4),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_77),
.A2(n_94),
.B1(n_72),
.B2(n_80),
.Y(n_129)
);

AND2x2_ASAP7_75t_L g130 ( 
.A(n_61),
.B(n_3),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_130),
.B(n_79),
.C(n_81),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_67),
.B(n_13),
.Y(n_132)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_78),
.Y(n_133)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_133),
.Y(n_142)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_80),
.Y(n_134)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_134),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_71),
.A2(n_4),
.B1(n_5),
.B2(n_7),
.Y(n_136)
);

AOI21xp33_ASAP7_75t_L g137 ( 
.A1(n_106),
.A2(n_82),
.B(n_65),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_SL g191 ( 
.A(n_137),
.B(n_143),
.Y(n_191)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_120),
.Y(n_140)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_140),
.Y(n_182)
);

INVx4_ASAP7_75t_L g141 ( 
.A(n_104),
.Y(n_141)
);

BUFx2_ASAP7_75t_L g177 ( 
.A(n_141),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_SL g143 ( 
.A(n_107),
.B(n_12),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_120),
.Y(n_144)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_144),
.Y(n_185)
);

AND2x2_ASAP7_75t_L g193 ( 
.A(n_145),
.B(n_65),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_SL g146 ( 
.A(n_114),
.B(n_11),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_146),
.B(n_151),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g171 ( 
.A(n_148),
.B(n_130),
.Y(n_171)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_110),
.Y(n_149)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_149),
.Y(n_189)
);

INVxp67_ASAP7_75t_SL g150 ( 
.A(n_104),
.Y(n_150)
);

CKINVDCx14_ASAP7_75t_R g188 ( 
.A(n_150),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_116),
.B(n_85),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_133),
.Y(n_152)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_152),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_123),
.B(n_68),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_155),
.B(n_157),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_156),
.A2(n_64),
.B1(n_131),
.B2(n_111),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_158),
.A2(n_165),
.B1(n_136),
.B2(n_130),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_123),
.B(n_5),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_159),
.B(n_164),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_122),
.B(n_72),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_161),
.B(n_118),
.Y(n_181)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_135),
.Y(n_163)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_163),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_112),
.B(n_106),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_129),
.A2(n_97),
.B1(n_100),
.B2(n_64),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_134),
.Y(n_166)
);

INVx2_ASAP7_75t_SL g196 ( 
.A(n_166),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_106),
.B(n_8),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_167),
.B(n_65),
.Y(n_176)
);

AOI21xp5_ASAP7_75t_L g169 ( 
.A1(n_145),
.A2(n_115),
.B(n_156),
.Y(n_169)
);

AOI21xp5_ASAP7_75t_L g208 ( 
.A1(n_169),
.A2(n_153),
.B(n_147),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_139),
.B(n_115),
.C(n_121),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_L g218 ( 
.A(n_170),
.B(n_144),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_SL g205 ( 
.A(n_171),
.B(n_153),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_161),
.A2(n_128),
.B1(n_117),
.B2(n_113),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_172),
.B(n_178),
.Y(n_200)
);

INVxp67_ASAP7_75t_L g209 ( 
.A(n_174),
.Y(n_209)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_175),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_SL g214 ( 
.A(n_176),
.B(n_186),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_139),
.A2(n_131),
.B1(n_118),
.B2(n_111),
.Y(n_178)
);

INVxp67_ASAP7_75t_L g180 ( 
.A(n_140),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_180),
.B(n_149),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_181),
.B(n_183),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_154),
.B(n_9),
.Y(n_183)
);

BUFx5_ASAP7_75t_L g184 ( 
.A(n_138),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_184),
.B(n_152),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_146),
.B(n_9),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_154),
.B(n_10),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_187),
.B(n_194),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_SL g203 ( 
.A1(n_193),
.A2(n_138),
.B(n_166),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_157),
.A2(n_10),
.B1(n_102),
.B2(n_158),
.Y(n_194)
);

AOI22xp33_ASAP7_75t_SL g198 ( 
.A1(n_177),
.A2(n_162),
.B1(n_141),
.B2(n_165),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_L g225 ( 
.A1(n_198),
.A2(n_209),
.B1(n_188),
.B2(n_177),
.Y(n_225)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_192),
.Y(n_199)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_199),
.Y(n_229)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_192),
.Y(n_201)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_201),
.Y(n_233)
);

INVxp67_ASAP7_75t_L g231 ( 
.A(n_203),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_181),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_204),
.B(n_210),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g232 ( 
.A(n_205),
.B(n_175),
.Y(n_232)
);

OAI21xp5_ASAP7_75t_SL g207 ( 
.A1(n_169),
.A2(n_153),
.B(n_148),
.Y(n_207)
);

OAI21xp5_ASAP7_75t_L g234 ( 
.A1(n_207),
.A2(n_208),
.B(n_194),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_211),
.B(n_212),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_172),
.B(n_160),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_189),
.Y(n_213)
);

AND2x2_ASAP7_75t_L g222 ( 
.A(n_213),
.B(n_195),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_190),
.B(n_143),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_SL g220 ( 
.A(n_215),
.B(n_217),
.Y(n_220)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_171),
.B(n_168),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_216),
.B(n_218),
.C(n_170),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_179),
.B(n_163),
.Y(n_217)
);

NOR3xp33_ASAP7_75t_SL g221 ( 
.A(n_212),
.B(n_193),
.C(n_187),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_SL g244 ( 
.A(n_221),
.B(n_228),
.Y(n_244)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_222),
.Y(n_240)
);

XNOR2x1_ASAP7_75t_L g236 ( 
.A(n_223),
.B(n_227),
.Y(n_236)
);

INVxp67_ASAP7_75t_L g245 ( 
.A(n_225),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_197),
.A2(n_193),
.B1(n_191),
.B2(n_178),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_L g246 ( 
.A1(n_226),
.A2(n_208),
.B1(n_209),
.B2(n_213),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_205),
.B(n_183),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_218),
.B(n_173),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_202),
.B(n_182),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_SL g242 ( 
.A(n_230),
.B(n_235),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_232),
.B(n_216),
.Y(n_239)
);

A2O1A1O1Ixp25_ASAP7_75t_L g238 ( 
.A1(n_234),
.A2(n_207),
.B(n_200),
.C(n_206),
.D(n_202),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_SL g235 ( 
.A(n_214),
.B(n_180),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_232),
.A2(n_197),
.B1(n_200),
.B2(n_204),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_237),
.A2(n_231),
.B1(n_224),
.B2(n_244),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_SL g253 ( 
.A(n_238),
.B(n_241),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_239),
.B(n_246),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_220),
.B(n_206),
.Y(n_241)
);

BUFx12f_ASAP7_75t_SL g243 ( 
.A(n_226),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_243),
.Y(n_250)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_240),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_247),
.B(n_248),
.Y(n_256)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_242),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_245),
.B(n_219),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_SL g260 ( 
.A(n_249),
.B(n_251),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_245),
.B(n_233),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_252),
.A2(n_238),
.B1(n_221),
.B2(n_229),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_236),
.B(n_223),
.C(n_228),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_255),
.B(n_236),
.C(n_227),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_250),
.B(n_237),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_257),
.B(n_259),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_SL g266 ( 
.A(n_258),
.B(n_262),
.Y(n_266)
);

AOI21xp5_ASAP7_75t_L g259 ( 
.A1(n_253),
.A2(n_231),
.B(n_243),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_261),
.B(n_255),
.C(n_199),
.Y(n_267)
);

AOI21xp5_ASAP7_75t_L g262 ( 
.A1(n_254),
.A2(n_203),
.B(n_222),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_256),
.A2(n_252),
.B1(n_249),
.B2(n_251),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_264),
.B(n_267),
.C(n_260),
.Y(n_268)
);

NOR2x1_ASAP7_75t_L g265 ( 
.A(n_260),
.B(n_254),
.Y(n_265)
);

OAI21xp5_ASAP7_75t_SL g269 ( 
.A1(n_265),
.A2(n_201),
.B(n_196),
.Y(n_269)
);

AOI21xp5_ASAP7_75t_L g272 ( 
.A1(n_268),
.A2(n_269),
.B(n_265),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_263),
.A2(n_196),
.B1(n_185),
.B2(n_142),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_270),
.B(n_196),
.C(n_266),
.Y(n_271)
);

AO21x1_ASAP7_75t_L g273 ( 
.A1(n_271),
.A2(n_272),
.B(n_267),
.Y(n_273)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_273),
.B(n_184),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_274),
.B(n_142),
.Y(n_275)
);


endmodule