module fake_jpeg_28262_n_171 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_171);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_171;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_1),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_13),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_2),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_7),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

INVx5_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_SL g22 ( 
.A(n_0),
.B(n_3),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_2),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

CKINVDCx14_ASAP7_75t_R g26 ( 
.A(n_5),
.Y(n_26)
);

INVx13_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_6),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_3),
.Y(n_30)
);

INVx11_ASAP7_75t_L g31 ( 
.A(n_23),
.Y(n_31)
);

INVx5_ASAP7_75t_L g48 ( 
.A(n_31),
.Y(n_48)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_23),
.Y(n_32)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_23),
.Y(n_33)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_33),
.Y(n_53)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_23),
.Y(n_34)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_34),
.Y(n_54)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_29),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_35),
.B(n_40),
.Y(n_45)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_29),
.Y(n_36)
);

INVx2_ASAP7_75t_SL g41 ( 
.A(n_36),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_22),
.B(n_0),
.Y(n_37)
);

OR2x2_ASAP7_75t_L g42 ( 
.A(n_37),
.B(n_22),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_29),
.Y(n_38)
);

INVx11_ASAP7_75t_L g44 ( 
.A(n_38),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_29),
.Y(n_39)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_39),
.Y(n_47)
);

BUFx5_ASAP7_75t_L g40 ( 
.A(n_27),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_42),
.B(n_46),
.Y(n_67)
);

OR2x2_ASAP7_75t_L g46 ( 
.A(n_37),
.B(n_15),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_32),
.B(n_15),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_49),
.B(n_52),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_L g50 ( 
.A1(n_36),
.A2(n_21),
.B1(n_27),
.B2(n_24),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_50),
.A2(n_21),
.B1(n_20),
.B2(n_30),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_40),
.B(n_19),
.Y(n_51)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_51),
.Y(n_66)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_34),
.Y(n_52)
);

OR2x2_ASAP7_75t_L g55 ( 
.A(n_40),
.B(n_18),
.Y(n_55)
);

INVx1_ASAP7_75t_SL g70 ( 
.A(n_55),
.Y(n_70)
);

AO22x2_ASAP7_75t_L g56 ( 
.A1(n_49),
.A2(n_35),
.B1(n_39),
.B2(n_31),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_56),
.A2(n_58),
.B1(n_65),
.B2(n_69),
.Y(n_82)
);

OAI22xp33_ASAP7_75t_L g58 ( 
.A1(n_54),
.A2(n_36),
.B1(n_34),
.B2(n_39),
.Y(n_58)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_44),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_59),
.B(n_60),
.Y(n_80)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_54),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_45),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_61),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_55),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_SL g85 ( 
.A(n_62),
.B(n_63),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_46),
.B(n_28),
.Y(n_63)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_43),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_64),
.B(n_68),
.Y(n_84)
);

AO22x1_ASAP7_75t_SL g65 ( 
.A1(n_41),
.A2(n_39),
.B1(n_38),
.B2(n_31),
.Y(n_65)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_55),
.Y(n_68)
);

INVxp67_ASAP7_75t_L g71 ( 
.A(n_41),
.Y(n_71)
);

INVxp67_ASAP7_75t_L g94 ( 
.A(n_71),
.Y(n_94)
);

INVxp67_ASAP7_75t_L g72 ( 
.A(n_41),
.Y(n_72)
);

INVxp67_ASAP7_75t_L g95 ( 
.A(n_72),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_43),
.A2(n_20),
.B1(n_18),
.B2(n_30),
.Y(n_73)
);

AND2x2_ASAP7_75t_L g93 ( 
.A(n_73),
.B(n_16),
.Y(n_93)
);

CKINVDCx14_ASAP7_75t_R g74 ( 
.A(n_53),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g96 ( 
.A(n_74),
.B(n_48),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_46),
.B(n_28),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g87 ( 
.A(n_75),
.B(n_76),
.Y(n_87)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_47),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_65),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_77),
.B(n_86),
.Y(n_109)
);

OAI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_56),
.A2(n_44),
.B1(n_24),
.B2(n_19),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_78),
.A2(n_89),
.B1(n_90),
.B2(n_72),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_57),
.B(n_70),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_79),
.B(n_81),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_70),
.B(n_42),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_67),
.B(n_42),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_83),
.B(n_91),
.Y(n_105)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_65),
.Y(n_86)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_56),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_88),
.B(n_96),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_56),
.A2(n_47),
.B1(n_52),
.B2(n_53),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_73),
.A2(n_16),
.B1(n_26),
.B2(n_17),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_64),
.B(n_69),
.Y(n_91)
);

CKINVDCx14_ASAP7_75t_R g106 ( 
.A(n_93),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_92),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_98),
.Y(n_124)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_80),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_99),
.B(n_100),
.Y(n_126)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_84),
.Y(n_100)
);

XOR2xp5_ASAP7_75t_L g101 ( 
.A(n_79),
.B(n_66),
.Y(n_101)
);

A2O1A1O1Ixp25_ASAP7_75t_L g117 ( 
.A1(n_101),
.A2(n_85),
.B(n_82),
.C(n_17),
.D(n_94),
.Y(n_117)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_89),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_102),
.B(n_104),
.Y(n_116)
);

OAI22x1_ASAP7_75t_SL g103 ( 
.A1(n_88),
.A2(n_58),
.B1(n_35),
.B2(n_33),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_103),
.A2(n_93),
.B1(n_95),
.B2(n_94),
.Y(n_115)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_91),
.Y(n_104)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_82),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_107),
.B(n_113),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_81),
.B(n_83),
.Y(n_108)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_108),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_77),
.B(n_71),
.Y(n_110)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_110),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_87),
.B(n_60),
.Y(n_112)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_112),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_L g114 ( 
.A1(n_111),
.A2(n_86),
.B(n_93),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_114),
.B(n_123),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_115),
.A2(n_113),
.B1(n_99),
.B2(n_100),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_117),
.A2(n_106),
.B1(n_103),
.B2(n_104),
.Y(n_134)
);

AOI21xp5_ASAP7_75t_SL g118 ( 
.A1(n_109),
.A2(n_95),
.B(n_33),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_118),
.B(n_125),
.Y(n_131)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_110),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_105),
.Y(n_125)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_105),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_127),
.B(n_128),
.Y(n_138)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_97),
.Y(n_128)
);

OAI21xp33_ASAP7_75t_L g129 ( 
.A1(n_121),
.A2(n_108),
.B(n_97),
.Y(n_129)
);

XOR2xp5_ASAP7_75t_L g149 ( 
.A(n_129),
.B(n_2),
.Y(n_149)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_126),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_130),
.B(n_136),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_120),
.B(n_101),
.C(n_107),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_132),
.B(n_139),
.C(n_118),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_134),
.A2(n_135),
.B1(n_140),
.B2(n_115),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_SL g136 ( 
.A(n_126),
.B(n_11),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_116),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_137),
.B(n_25),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_120),
.B(n_38),
.C(n_48),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_119),
.A2(n_59),
.B1(n_17),
.B2(n_25),
.Y(n_140)
);

AOI321xp33_ASAP7_75t_L g141 ( 
.A1(n_129),
.A2(n_114),
.A3(n_117),
.B1(n_122),
.B2(n_121),
.C(n_124),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_L g151 ( 
.A(n_141),
.B(n_148),
.Y(n_151)
);

CKINVDCx6p67_ASAP7_75t_R g142 ( 
.A(n_139),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_142),
.B(n_144),
.Y(n_153)
);

OR2x2_ASAP7_75t_L g150 ( 
.A(n_143),
.B(n_140),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_145),
.B(n_4),
.C(n_6),
.Y(n_156)
);

OA21x2_ASAP7_75t_SL g147 ( 
.A1(n_133),
.A2(n_132),
.B(n_131),
.Y(n_147)
);

OAI31xp33_ASAP7_75t_L g155 ( 
.A1(n_147),
.A2(n_149),
.A3(n_145),
.B(n_148),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_L g148 ( 
.A(n_134),
.B(n_1),
.Y(n_148)
);

XNOR2xp5_ASAP7_75t_L g154 ( 
.A(n_149),
.B(n_3),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_150),
.A2(n_142),
.B1(n_9),
.B2(n_10),
.Y(n_158)
);

AOI21xp5_ASAP7_75t_SL g152 ( 
.A1(n_146),
.A2(n_138),
.B(n_4),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_152),
.B(n_154),
.Y(n_157)
);

AOI21xp5_ASAP7_75t_L g160 ( 
.A1(n_155),
.A2(n_151),
.B(n_153),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_156),
.B(n_8),
.C(n_9),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_158),
.B(n_159),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_153),
.B(n_142),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_160),
.B(n_161),
.C(n_14),
.Y(n_164)
);

OAI21x1_ASAP7_75t_SL g163 ( 
.A1(n_158),
.A2(n_150),
.B(n_12),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_163),
.B(n_165),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_164),
.B(n_161),
.C(n_14),
.Y(n_166)
);

AOI21xp5_ASAP7_75t_L g165 ( 
.A1(n_157),
.A2(n_10),
.B(n_13),
.Y(n_165)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_166),
.Y(n_168)
);

BUFx24_ASAP7_75t_SL g169 ( 
.A(n_167),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_169),
.B(n_162),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_L g171 ( 
.A(n_170),
.B(n_168),
.Y(n_171)
);


endmodule