module fake_ariane_786_n_1827 (n_83, n_8, n_56, n_60, n_170, n_160, n_64, n_119, n_124, n_167, n_90, n_38, n_47, n_110, n_153, n_18, n_86, n_75, n_89, n_67, n_176, n_149, n_34, n_158, n_172, n_69, n_95, n_175, n_92, n_143, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_152, n_120, n_169, n_106, n_12, n_53, n_173, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_156, n_49, n_20, n_174, n_100, n_17, n_50, n_132, n_62, n_147, n_51, n_166, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_159, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_148, n_164, n_52, n_157, n_135, n_73, n_77, n_171, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_151, n_136, n_28, n_80, n_146, n_97, n_154, n_142, n_161, n_14, n_163, n_88, n_141, n_68, n_116, n_104, n_145, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_1827);

input n_83;
input n_8;
input n_56;
input n_60;
input n_170;
input n_160;
input n_64;
input n_119;
input n_124;
input n_167;
input n_90;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_176;
input n_149;
input n_34;
input n_158;
input n_172;
input n_69;
input n_95;
input n_175;
input n_92;
input n_143;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_152;
input n_120;
input n_169;
input n_106;
input n_12;
input n_53;
input n_173;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_156;
input n_49;
input n_20;
input n_174;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_147;
input n_51;
input n_166;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_159;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_164;
input n_52;
input n_157;
input n_135;
input n_73;
input n_77;
input n_171;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_151;
input n_136;
input n_28;
input n_80;
input n_146;
input n_97;
input n_154;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_1827;

wire n_913;
wire n_1681;
wire n_1486;
wire n_1507;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_1250;
wire n_1169;
wire n_789;
wire n_850;
wire n_610;
wire n_245;
wire n_1713;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_187;
wire n_1463;
wire n_1238;
wire n_1515;
wire n_817;
wire n_924;
wire n_781;
wire n_1566;
wire n_189;
wire n_717;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_1706;
wire n_524;
wire n_634;
wire n_1214;
wire n_1246;
wire n_1138;
wire n_214;
wire n_764;
wire n_1503;
wire n_462;
wire n_1196;
wire n_1181;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1745;
wire n_1366;
wire n_232;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1457;
wire n_377;
wire n_1682;
wire n_520;
wire n_870;
wire n_1453;
wire n_279;
wire n_958;
wire n_945;
wire n_813;
wire n_419;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1184;
wire n_202;
wire n_1535;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_1277;
wire n_1746;
wire n_829;
wire n_1761;
wire n_1062;
wire n_339;
wire n_738;
wire n_1690;
wire n_672;
wire n_740;
wire n_1283;
wire n_1736;
wire n_1018;
wire n_259;
wire n_953;
wire n_1364;
wire n_1224;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_1688;
wire n_989;
wire n_242;
wire n_645;
wire n_331;
wire n_559;
wire n_267;
wire n_495;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_200;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_1522;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_1404;
wire n_868;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_1676;
wire n_1085;
wire n_277;
wire n_1636;
wire n_432;
wire n_293;
wire n_823;
wire n_620;
wire n_1074;
wire n_859;
wire n_1765;
wire n_587;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_206;
wire n_352;
wire n_899;
wire n_1703;
wire n_611;
wire n_1295;
wire n_365;
wire n_238;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_334;
wire n_192;
wire n_661;
wire n_1751;
wire n_300;
wire n_533;
wire n_438;
wire n_1560;
wire n_1654;
wire n_1548;
wire n_1811;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_376;
wire n_512;
wire n_1597;
wire n_1771;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1354;
wire n_1790;
wire n_1213;
wire n_237;
wire n_780;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_490;
wire n_209;
wire n_1461;
wire n_1391;
wire n_225;
wire n_1599;
wire n_1006;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_1594;
wire n_680;
wire n_287;
wire n_1716;
wire n_302;
wire n_380;
wire n_1585;
wire n_1432;
wire n_249;
wire n_1108;
wire n_355;
wire n_212;
wire n_444;
wire n_851;
wire n_1590;
wire n_1351;
wire n_1274;
wire n_257;
wire n_652;
wire n_1819;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_182;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_407;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_460;
wire n_1555;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_966;
wire n_992;
wire n_955;
wire n_1182;
wire n_794;
wire n_1692;
wire n_1562;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_288;
wire n_179;
wire n_1292;
wire n_1178;
wire n_1435;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_306;
wire n_203;
wire n_436;
wire n_324;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_437;
wire n_337;
wire n_274;
wire n_967;
wire n_1083;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1787;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_1717;
wire n_1812;
wire n_824;
wire n_428;
wire n_892;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_990;
wire n_1623;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_1780;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1825;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1680;
wire n_964;
wire n_1627;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_1731;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_934;
wire n_1447;
wire n_1220;
wire n_356;
wire n_698;
wire n_1674;
wire n_307;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_1633;
wire n_404;
wire n_1058;
wire n_347;
wire n_1042;
wire n_183;
wire n_1234;
wire n_479;
wire n_1578;
wire n_1455;
wire n_299;
wire n_836;
wire n_1279;
wire n_564;
wire n_205;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_1689;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_1728;
wire n_370;
wire n_706;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_1817;
wire n_348;
wire n_552;
wire n_670;
wire n_1826;
wire n_379;
wire n_264;
wire n_441;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_1618;
wire n_1743;
wire n_905;
wire n_207;
wire n_720;
wire n_926;
wire n_194;
wire n_1802;
wire n_1163;
wire n_186;
wire n_1795;
wire n_1384;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1648;
wire n_1413;
wire n_855;
wire n_808;
wire n_1365;
wire n_553;
wire n_1439;
wire n_814;
wire n_578;
wire n_1665;
wire n_1287;
wire n_405;
wire n_1611;
wire n_320;
wire n_1414;
wire n_1134;
wire n_1484;
wire n_647;
wire n_1423;
wire n_481;
wire n_600;
wire n_1053;
wire n_1609;
wire n_529;
wire n_502;
wire n_218;
wire n_1467;
wire n_247;
wire n_1798;
wire n_1304;
wire n_1608;
wire n_1744;
wire n_1105;
wire n_547;
wire n_439;
wire n_604;
wire n_677;
wire n_478;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_1278;
wire n_707;
wire n_983;
wire n_590;
wire n_727;
wire n_699;
wire n_301;
wire n_1726;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_325;
wire n_1740;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_729;
wire n_887;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_1693;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1823;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_233;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_321;
wire n_221;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1763;
wire n_1666;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_281;
wire n_262;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_1667;
wire n_845;
wire n_888;
wire n_1649;
wire n_1677;
wire n_1297;
wire n_178;
wire n_551;
wire n_417;
wire n_1708;
wire n_343;
wire n_1222;
wire n_582;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_534;
wire n_1791;
wire n_1460;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_451;
wire n_745;
wire n_1741;
wire n_1572;
wire n_1793;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_769;
wire n_1797;
wire n_1753;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_982;
wire n_1800;
wire n_915;
wire n_215;
wire n_1075;
wire n_454;
wire n_298;
wire n_1331;
wire n_1529;
wire n_1227;
wire n_655;
wire n_1734;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_1700;
wire n_659;
wire n_1332;
wire n_509;
wire n_666;
wire n_1747;
wire n_430;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1766;
wire n_1338;
wire n_1342;
wire n_456;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_521;
wire n_873;
wire n_1301;
wire n_1748;
wire n_1243;
wire n_1400;
wire n_342;
wire n_1466;
wire n_1513;
wire n_1527;
wire n_358;
wire n_1783;
wire n_608;
wire n_1538;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1668;
wire n_1605;
wire n_1078;
wire n_266;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_687;
wire n_797;
wire n_1786;
wire n_480;
wire n_1327;
wire n_1475;
wire n_211;
wire n_642;
wire n_1804;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_1757;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_393;
wire n_1632;
wire n_1769;
wire n_474;
wire n_805;
wire n_295;
wire n_1658;
wire n_190;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_180;
wire n_730;
wire n_386;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1137;
wire n_1258;
wire n_197;
wire n_640;
wire n_463;
wire n_1476;
wire n_1524;
wire n_1733;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_1807;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_1784;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_283;
wire n_806;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_1824;
wire n_643;
wire n_1492;
wire n_226;
wire n_1441;
wire n_1822;
wire n_682;
wire n_1616;
wire n_819;
wire n_586;
wire n_1324;
wire n_1429;
wire n_1778;
wire n_1776;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1759;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_1815;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_198;
wire n_1208;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1577;
wire n_1448;
wire n_1009;
wire n_230;
wire n_1133;
wire n_883;
wire n_473;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_594;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_1201;
wire n_1288;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_426;
wire n_433;
wire n_398;
wire n_210;
wire n_1090;
wire n_1367;
wire n_253;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_224;
wire n_894;
wire n_1380;
wire n_1624;
wire n_1801;
wire n_420;
wire n_1291;
wire n_562;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1023;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_467;
wire n_1511;
wire n_1422;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_1641;
wire n_538;
wire n_1517;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_1307;
wire n_1128;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1773;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_810;
wire n_1290;
wire n_181;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_236;
wire n_683;
wire n_601;
wire n_565;
wire n_628;
wire n_1300;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_414;
wire n_571;
wire n_1521;
wire n_1694;
wire n_284;
wire n_593;
wire n_1695;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_1774;
wire n_409;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_526;
wire n_1767;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1444;
wire n_1803;
wire n_820;
wire n_1749;
wire n_872;
wire n_1653;
wire n_254;
wire n_1157;
wire n_1584;
wire n_234;
wire n_848;
wire n_1664;
wire n_280;
wire n_629;
wire n_1739;
wire n_1814;
wire n_532;
wire n_1789;
wire n_763;
wire n_540;
wire n_216;
wire n_692;
wire n_984;
wire n_1687;
wire n_223;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_1816;
wire n_1756;
wire n_1606;
wire n_395;
wire n_621;
wire n_1587;
wire n_213;
wire n_1772;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_493;
wire n_1311;
wire n_1589;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_697;
wire n_622;
wire n_1626;
wire n_1335;
wire n_1715;
wire n_296;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_1785;
wire n_792;
wire n_1262;
wire n_580;
wire n_1579;
wire n_494;
wire n_434;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1183;
wire n_1326;
wire n_1805;
wire n_981;
wire n_1110;
wire n_1758;
wire n_243;
wire n_1407;
wire n_185;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_184;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_1054;
wire n_508;
wire n_1679;
wire n_353;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_191;
wire n_978;
wire n_1011;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_1721;
wire n_653;
wire n_1445;
wire n_1317;
wire n_783;
wire n_556;
wire n_1127;
wire n_1536;
wire n_1471;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_541;
wire n_499;
wire n_1775;
wire n_788;
wire n_908;
wire n_1036;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_1663;
wire n_1625;
wire n_318;
wire n_1458;
wire n_244;
wire n_679;
wire n_1630;
wire n_220;
wire n_663;
wire n_1720;
wire n_443;
wire n_1412;
wire n_1738;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_1735;
wire n_1788;
wire n_391;
wire n_940;
wire n_1537;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_765;
wire n_1809;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_1530;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_857;
wire n_898;
wire n_363;
wire n_968;
wire n_1067;
wire n_1235;
wire n_1323;
wire n_1462;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_1755;
wire n_1285;
wire n_193;
wire n_733;
wire n_761;
wire n_731;
wire n_336;
wire n_1813;
wire n_315;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_1106;
wire n_648;
wire n_784;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_1348;
wire n_753;
wire n_1770;
wire n_701;
wire n_1003;
wire n_1125;
wire n_1710;
wire n_309;
wire n_1344;
wire n_1390;
wire n_401;
wire n_485;
wire n_1792;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_291;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1510;
wire n_1099;
wire n_839;
wire n_1754;
wire n_759;
wire n_567;
wire n_240;
wire n_369;
wire n_1727;
wire n_1575;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_188;
wire n_323;
wire n_550;
wire n_1315;
wire n_1660;
wire n_997;
wire n_635;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_248;
wire n_1152;
wire n_921;
wire n_1615;
wire n_1236;
wire n_228;
wire n_1265;
wire n_1576;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1806;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1684;
wire n_1673;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_1696;
wire n_498;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1497;
wire n_459;
wire n_1136;
wire n_1782;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_383;
wire n_838;
wire n_1558;
wire n_1316;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_1781;
wire n_709;
wire n_809;
wire n_1686;
wire n_235;
wire n_881;
wire n_1019;
wire n_1477;
wire n_1777;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_199;
wire n_217;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_708;
wire n_308;
wire n_1223;
wire n_201;
wire n_1768;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1041;
wire n_993;
wire n_948;
wire n_922;
wire n_1004;
wire n_1810;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_1764;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_196;
wire n_1337;
wire n_774;
wire n_933;
wire n_1779;
wire n_596;
wire n_954;
wire n_1168;
wire n_1821;
wire n_219;
wire n_1310;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_252;
wire n_664;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_1732;
wire n_415;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1724;
wire n_1670;
wire n_1799;
wire n_1707;
wire n_1126;
wire n_195;
wire n_938;
wire n_1328;
wire n_895;
wire n_304;
wire n_1639;
wire n_583;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_946;
wire n_757;
wire n_375;
wire n_1655;
wire n_1818;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_472;
wire n_937;
wire n_1474;
wire n_265;
wire n_1583;
wire n_1604;
wire n_208;
wire n_1631;
wire n_1702;
wire n_275;
wire n_1794;
wire n_1375;
wire n_204;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_496;
wire n_866;
wire n_246;
wire n_925;
wire n_1752;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_1129;
wire n_1252;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_329;
wire n_718;
wire n_1434;
wire n_340;
wire n_1569;
wire n_548;
wire n_289;
wire n_523;
wire n_1662;
wire n_457;
wire n_1299;
wire n_177;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1228;
wire n_1244;
wire n_1796;
wire n_411;
wire n_484;
wire n_849;
wire n_1820;
wire n_357;
wire n_412;
wire n_1251;
wire n_447;
wire n_1421;
wire n_1762;
wire n_1233;
wire n_1808;
wire n_1574;
wire n_1672;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_1487;
wire n_675;

INVx2_ASAP7_75t_SL g177 ( 
.A(n_164),
.Y(n_177)
);

BUFx3_ASAP7_75t_L g178 ( 
.A(n_18),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_170),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_105),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_7),
.Y(n_181)
);

BUFx10_ASAP7_75t_L g182 ( 
.A(n_18),
.Y(n_182)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_108),
.Y(n_183)
);

BUFx2_ASAP7_75t_SL g184 ( 
.A(n_140),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_47),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_86),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_37),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_129),
.Y(n_188)
);

BUFx2_ASAP7_75t_L g189 ( 
.A(n_63),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_152),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_73),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_121),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_119),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_77),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_35),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_147),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_91),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_132),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_2),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_53),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_131),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_156),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_17),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_3),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_120),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_116),
.Y(n_206)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_57),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_53),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_166),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_59),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_47),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_146),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_128),
.Y(n_213)
);

BUFx6f_ASAP7_75t_L g214 ( 
.A(n_61),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_25),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_63),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_36),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_42),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_138),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_52),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_30),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_15),
.Y(n_222)
);

INVxp67_ASAP7_75t_L g223 ( 
.A(n_13),
.Y(n_223)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_159),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_58),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_27),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_0),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_117),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_58),
.Y(n_229)
);

INVxp67_ASAP7_75t_L g230 ( 
.A(n_126),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_122),
.Y(n_231)
);

BUFx3_ASAP7_75t_L g232 ( 
.A(n_22),
.Y(n_232)
);

BUFx10_ASAP7_75t_L g233 ( 
.A(n_57),
.Y(n_233)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_78),
.Y(n_234)
);

BUFx10_ASAP7_75t_L g235 ( 
.A(n_127),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_95),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_98),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_34),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_79),
.Y(n_239)
);

HB1xp67_ASAP7_75t_L g240 ( 
.A(n_88),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_148),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_27),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_52),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_49),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_9),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_55),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_110),
.Y(n_247)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_74),
.Y(n_248)
);

CKINVDCx16_ASAP7_75t_R g249 ( 
.A(n_64),
.Y(n_249)
);

BUFx3_ASAP7_75t_L g250 ( 
.A(n_134),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_85),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_115),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_145),
.Y(n_253)
);

CKINVDCx11_ASAP7_75t_R g254 ( 
.A(n_2),
.Y(n_254)
);

INVx1_ASAP7_75t_SL g255 ( 
.A(n_45),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_37),
.Y(n_256)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_112),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_167),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_14),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_174),
.Y(n_260)
);

HB1xp67_ASAP7_75t_L g261 ( 
.A(n_113),
.Y(n_261)
);

CKINVDCx16_ASAP7_75t_R g262 ( 
.A(n_62),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_141),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_102),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_8),
.Y(n_265)
);

CKINVDCx16_ASAP7_75t_R g266 ( 
.A(n_64),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_35),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_153),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_12),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_109),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_125),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_36),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_161),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_94),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_59),
.Y(n_275)
);

BUFx3_ASAP7_75t_L g276 ( 
.A(n_19),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_13),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_118),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_123),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_33),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_4),
.Y(n_281)
);

BUFx8_ASAP7_75t_SL g282 ( 
.A(n_143),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_130),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_43),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_3),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_55),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_54),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_154),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_81),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_34),
.Y(n_290)
);

HB1xp67_ASAP7_75t_L g291 ( 
.A(n_114),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_60),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_46),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_80),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_103),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g296 ( 
.A(n_162),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_144),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g298 ( 
.A(n_71),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_14),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_163),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_30),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_43),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_136),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_87),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_93),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_51),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_60),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_7),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_33),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_32),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_83),
.Y(n_311)
);

HB1xp67_ASAP7_75t_L g312 ( 
.A(n_54),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_44),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_50),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_44),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_10),
.Y(n_316)
);

INVx2_ASAP7_75t_L g317 ( 
.A(n_65),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_17),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_48),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_96),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_84),
.Y(n_321)
);

INVx3_ASAP7_75t_L g322 ( 
.A(n_62),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_16),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_151),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_111),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_46),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_160),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_0),
.Y(n_328)
);

CKINVDCx20_ASAP7_75t_R g329 ( 
.A(n_69),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_107),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_26),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g332 ( 
.A(n_68),
.Y(n_332)
);

INVx1_ASAP7_75t_SL g333 ( 
.A(n_22),
.Y(n_333)
);

INVx2_ASAP7_75t_L g334 ( 
.A(n_104),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_157),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_48),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_5),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_32),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_90),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_124),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_139),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_9),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_6),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_8),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_176),
.Y(n_345)
);

CKINVDCx20_ASAP7_75t_R g346 ( 
.A(n_42),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_89),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_169),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_4),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_50),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_67),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_20),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_254),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_282),
.Y(n_354)
);

INVxp67_ASAP7_75t_SL g355 ( 
.A(n_322),
.Y(n_355)
);

NOR2xp33_ASAP7_75t_R g356 ( 
.A(n_201),
.B(n_175),
.Y(n_356)
);

INVxp67_ASAP7_75t_L g357 ( 
.A(n_189),
.Y(n_357)
);

NOR2xp67_ASAP7_75t_L g358 ( 
.A(n_322),
.B(n_1),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_322),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_247),
.Y(n_360)
);

CKINVDCx20_ASAP7_75t_R g361 ( 
.A(n_252),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_296),
.Y(n_362)
);

CKINVDCx20_ASAP7_75t_R g363 ( 
.A(n_298),
.Y(n_363)
);

CKINVDCx20_ASAP7_75t_R g364 ( 
.A(n_329),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_332),
.Y(n_365)
);

BUFx3_ASAP7_75t_L g366 ( 
.A(n_250),
.Y(n_366)
);

INVxp67_ASAP7_75t_L g367 ( 
.A(n_189),
.Y(n_367)
);

CKINVDCx20_ASAP7_75t_R g368 ( 
.A(n_281),
.Y(n_368)
);

HB1xp67_ASAP7_75t_L g369 ( 
.A(n_249),
.Y(n_369)
);

INVxp67_ASAP7_75t_L g370 ( 
.A(n_312),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_322),
.Y(n_371)
);

INVx2_ASAP7_75t_L g372 ( 
.A(n_214),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_249),
.Y(n_373)
);

INVx2_ASAP7_75t_L g374 ( 
.A(n_214),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_180),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_180),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_262),
.Y(n_377)
);

NOR2xp33_ASAP7_75t_L g378 ( 
.A(n_186),
.B(n_191),
.Y(n_378)
);

NOR2xp33_ASAP7_75t_L g379 ( 
.A(n_186),
.B(n_1),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_191),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_262),
.Y(n_381)
);

AND2x4_ASAP7_75t_L g382 ( 
.A(n_178),
.B(n_5),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_266),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_266),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_181),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_206),
.Y(n_386)
);

CKINVDCx20_ASAP7_75t_R g387 ( 
.A(n_346),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_206),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_187),
.Y(n_389)
);

CKINVDCx20_ASAP7_75t_R g390 ( 
.A(n_250),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_212),
.Y(n_391)
);

CKINVDCx20_ASAP7_75t_R g392 ( 
.A(n_250),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_195),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_212),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_219),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_219),
.Y(n_396)
);

NOR2xp67_ASAP7_75t_L g397 ( 
.A(n_317),
.B(n_6),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_228),
.Y(n_398)
);

CKINVDCx20_ASAP7_75t_R g399 ( 
.A(n_235),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_228),
.Y(n_400)
);

CKINVDCx20_ASAP7_75t_R g401 ( 
.A(n_235),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_240),
.B(n_10),
.Y(n_402)
);

CKINVDCx20_ASAP7_75t_R g403 ( 
.A(n_235),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_231),
.Y(n_404)
);

CKINVDCx20_ASAP7_75t_R g405 ( 
.A(n_235),
.Y(n_405)
);

BUFx2_ASAP7_75t_L g406 ( 
.A(n_178),
.Y(n_406)
);

BUFx6f_ASAP7_75t_L g407 ( 
.A(n_214),
.Y(n_407)
);

CKINVDCx20_ASAP7_75t_R g408 ( 
.A(n_182),
.Y(n_408)
);

NOR2xp67_ASAP7_75t_L g409 ( 
.A(n_317),
.B(n_11),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_261),
.B(n_11),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_199),
.Y(n_411)
);

INVxp67_ASAP7_75t_L g412 ( 
.A(n_185),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_231),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_251),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_203),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_211),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_251),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_258),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_215),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_216),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_217),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_258),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_264),
.Y(n_423)
);

CKINVDCx16_ASAP7_75t_R g424 ( 
.A(n_182),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_218),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_220),
.Y(n_426)
);

CKINVDCx20_ASAP7_75t_R g427 ( 
.A(n_182),
.Y(n_427)
);

NOR2xp33_ASAP7_75t_L g428 ( 
.A(n_264),
.B(n_12),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_270),
.Y(n_429)
);

INVxp33_ASAP7_75t_L g430 ( 
.A(n_185),
.Y(n_430)
);

INVxp33_ASAP7_75t_SL g431 ( 
.A(n_222),
.Y(n_431)
);

CKINVDCx14_ASAP7_75t_R g432 ( 
.A(n_182),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_270),
.Y(n_433)
);

CKINVDCx20_ASAP7_75t_R g434 ( 
.A(n_233),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_271),
.Y(n_435)
);

INVx1_ASAP7_75t_SL g436 ( 
.A(n_255),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_271),
.Y(n_437)
);

INVxp67_ASAP7_75t_L g438 ( 
.A(n_200),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_273),
.Y(n_439)
);

CKINVDCx5p33_ASAP7_75t_R g440 ( 
.A(n_225),
.Y(n_440)
);

OA21x2_ASAP7_75t_L g441 ( 
.A1(n_372),
.A2(n_274),
.B(n_273),
.Y(n_441)
);

INVx3_ASAP7_75t_L g442 ( 
.A(n_407),
.Y(n_442)
);

BUFx6f_ASAP7_75t_L g443 ( 
.A(n_407),
.Y(n_443)
);

AOI22xp5_ASAP7_75t_L g444 ( 
.A1(n_436),
.A2(n_357),
.B1(n_367),
.B2(n_399),
.Y(n_444)
);

INVxp67_ASAP7_75t_L g445 ( 
.A(n_369),
.Y(n_445)
);

BUFx6f_ASAP7_75t_L g446 ( 
.A(n_407),
.Y(n_446)
);

INVx2_ASAP7_75t_L g447 ( 
.A(n_407),
.Y(n_447)
);

AND2x2_ASAP7_75t_L g448 ( 
.A(n_406),
.B(n_178),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_359),
.Y(n_449)
);

BUFx6f_ASAP7_75t_L g450 ( 
.A(n_407),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_359),
.Y(n_451)
);

AND2x2_ASAP7_75t_L g452 ( 
.A(n_406),
.B(n_232),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_371),
.Y(n_453)
);

BUFx6f_ASAP7_75t_L g454 ( 
.A(n_372),
.Y(n_454)
);

NOR2xp33_ASAP7_75t_L g455 ( 
.A(n_355),
.B(n_291),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_371),
.B(n_274),
.Y(n_456)
);

CKINVDCx20_ASAP7_75t_R g457 ( 
.A(n_368),
.Y(n_457)
);

INVx2_ASAP7_75t_L g458 ( 
.A(n_374),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_378),
.B(n_366),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_375),
.Y(n_460)
);

INVx3_ASAP7_75t_L g461 ( 
.A(n_374),
.Y(n_461)
);

BUFx2_ASAP7_75t_L g462 ( 
.A(n_373),
.Y(n_462)
);

INVx2_ASAP7_75t_L g463 ( 
.A(n_375),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_376),
.Y(n_464)
);

INVx2_ASAP7_75t_L g465 ( 
.A(n_376),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_L g466 ( 
.A(n_366),
.B(n_278),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_L g467 ( 
.A(n_380),
.B(n_386),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_L g468 ( 
.A(n_380),
.B(n_278),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_386),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_388),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_SL g471 ( 
.A(n_424),
.B(n_233),
.Y(n_471)
);

HB1xp67_ASAP7_75t_L g472 ( 
.A(n_377),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_388),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_391),
.Y(n_474)
);

NOR2xp33_ASAP7_75t_L g475 ( 
.A(n_431),
.B(n_230),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_391),
.Y(n_476)
);

INVx2_ASAP7_75t_L g477 ( 
.A(n_394),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_L g478 ( 
.A(n_394),
.B(n_294),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_395),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_L g480 ( 
.A(n_395),
.B(n_294),
.Y(n_480)
);

BUFx6f_ASAP7_75t_L g481 ( 
.A(n_382),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_396),
.Y(n_482)
);

NOR2xp33_ASAP7_75t_L g483 ( 
.A(n_385),
.B(n_300),
.Y(n_483)
);

NAND2x1p5_ASAP7_75t_L g484 ( 
.A(n_382),
.B(n_300),
.Y(n_484)
);

BUFx6f_ASAP7_75t_L g485 ( 
.A(n_382),
.Y(n_485)
);

INVx4_ASAP7_75t_L g486 ( 
.A(n_382),
.Y(n_486)
);

INVx2_ASAP7_75t_L g487 ( 
.A(n_396),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_398),
.Y(n_488)
);

AND2x2_ASAP7_75t_L g489 ( 
.A(n_430),
.B(n_232),
.Y(n_489)
);

HB1xp67_ASAP7_75t_L g490 ( 
.A(n_381),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_L g491 ( 
.A(n_398),
.B(n_305),
.Y(n_491)
);

BUFx3_ASAP7_75t_L g492 ( 
.A(n_400),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_400),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_404),
.B(n_305),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_L g495 ( 
.A(n_404),
.B(n_320),
.Y(n_495)
);

HB1xp67_ASAP7_75t_L g496 ( 
.A(n_383),
.Y(n_496)
);

INVx3_ASAP7_75t_L g497 ( 
.A(n_413),
.Y(n_497)
);

INVx2_ASAP7_75t_L g498 ( 
.A(n_413),
.Y(n_498)
);

NAND2xp33_ASAP7_75t_L g499 ( 
.A(n_389),
.B(n_214),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_414),
.Y(n_500)
);

INVx2_ASAP7_75t_L g501 ( 
.A(n_414),
.Y(n_501)
);

BUFx6f_ASAP7_75t_L g502 ( 
.A(n_417),
.Y(n_502)
);

BUFx6f_ASAP7_75t_L g503 ( 
.A(n_417),
.Y(n_503)
);

AND2x4_ASAP7_75t_L g504 ( 
.A(n_418),
.B(n_422),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_418),
.Y(n_505)
);

AND2x4_ASAP7_75t_L g506 ( 
.A(n_422),
.B(n_232),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_L g507 ( 
.A(n_423),
.B(n_320),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_423),
.Y(n_508)
);

BUFx6f_ASAP7_75t_L g509 ( 
.A(n_429),
.Y(n_509)
);

INVx5_ASAP7_75t_L g510 ( 
.A(n_358),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_429),
.Y(n_511)
);

NOR2xp33_ASAP7_75t_L g512 ( 
.A(n_393),
.B(n_321),
.Y(n_512)
);

NOR2xp33_ASAP7_75t_L g513 ( 
.A(n_411),
.B(n_321),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_433),
.Y(n_514)
);

BUFx8_ASAP7_75t_L g515 ( 
.A(n_432),
.Y(n_515)
);

BUFx6f_ASAP7_75t_L g516 ( 
.A(n_433),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_435),
.Y(n_517)
);

NOR2xp33_ASAP7_75t_L g518 ( 
.A(n_459),
.B(n_415),
.Y(n_518)
);

INVx2_ASAP7_75t_L g519 ( 
.A(n_458),
.Y(n_519)
);

AOI22xp33_ASAP7_75t_L g520 ( 
.A1(n_455),
.A2(n_402),
.B1(n_410),
.B2(n_379),
.Y(n_520)
);

OR2x6_ASAP7_75t_L g521 ( 
.A(n_484),
.B(n_397),
.Y(n_521)
);

XNOR2xp5_ASAP7_75t_L g522 ( 
.A(n_444),
.B(n_387),
.Y(n_522)
);

AOI22xp33_ASAP7_75t_L g523 ( 
.A1(n_484),
.A2(n_428),
.B1(n_409),
.B2(n_370),
.Y(n_523)
);

INVx2_ASAP7_75t_L g524 ( 
.A(n_458),
.Y(n_524)
);

BUFx2_ASAP7_75t_L g525 ( 
.A(n_445),
.Y(n_525)
);

XNOR2xp5_ASAP7_75t_L g526 ( 
.A(n_444),
.B(n_361),
.Y(n_526)
);

CKINVDCx20_ASAP7_75t_R g527 ( 
.A(n_457),
.Y(n_527)
);

OR2x6_ASAP7_75t_L g528 ( 
.A(n_484),
.B(n_412),
.Y(n_528)
);

INVx2_ASAP7_75t_L g529 ( 
.A(n_458),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_502),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_L g531 ( 
.A(n_459),
.B(n_504),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_SL g532 ( 
.A(n_475),
.B(n_416),
.Y(n_532)
);

INVx2_ASAP7_75t_L g533 ( 
.A(n_461),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_502),
.Y(n_534)
);

INVx2_ASAP7_75t_L g535 ( 
.A(n_461),
.Y(n_535)
);

BUFx3_ASAP7_75t_L g536 ( 
.A(n_515),
.Y(n_536)
);

INVxp67_ASAP7_75t_L g537 ( 
.A(n_462),
.Y(n_537)
);

INVxp67_ASAP7_75t_SL g538 ( 
.A(n_481),
.Y(n_538)
);

INVx2_ASAP7_75t_L g539 ( 
.A(n_461),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_502),
.Y(n_540)
);

INVx2_ASAP7_75t_L g541 ( 
.A(n_461),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_L g542 ( 
.A(n_504),
.B(n_483),
.Y(n_542)
);

NOR2xp33_ASAP7_75t_L g543 ( 
.A(n_512),
.B(n_513),
.Y(n_543)
);

AOI22xp33_ASAP7_75t_L g544 ( 
.A1(n_484),
.A2(n_392),
.B1(n_390),
.B2(n_435),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_L g545 ( 
.A(n_504),
.B(n_437),
.Y(n_545)
);

INVxp33_ASAP7_75t_L g546 ( 
.A(n_472),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_L g547 ( 
.A(n_504),
.B(n_437),
.Y(n_547)
);

AND2x2_ASAP7_75t_L g548 ( 
.A(n_489),
.B(n_439),
.Y(n_548)
);

NAND2xp33_ASAP7_75t_L g549 ( 
.A(n_481),
.B(n_356),
.Y(n_549)
);

INVx6_ASAP7_75t_L g550 ( 
.A(n_486),
.Y(n_550)
);

INVxp33_ASAP7_75t_L g551 ( 
.A(n_472),
.Y(n_551)
);

INVx2_ASAP7_75t_L g552 ( 
.A(n_502),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_L g553 ( 
.A(n_492),
.B(n_439),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_L g554 ( 
.A(n_492),
.B(n_419),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_L g555 ( 
.A(n_492),
.B(n_420),
.Y(n_555)
);

INVx2_ASAP7_75t_L g556 ( 
.A(n_502),
.Y(n_556)
);

AOI22xp33_ASAP7_75t_L g557 ( 
.A1(n_441),
.A2(n_401),
.B1(n_403),
.B2(n_405),
.Y(n_557)
);

CKINVDCx6p67_ASAP7_75t_R g558 ( 
.A(n_462),
.Y(n_558)
);

AOI22xp5_ASAP7_75t_L g559 ( 
.A1(n_445),
.A2(n_333),
.B1(n_223),
.B2(n_259),
.Y(n_559)
);

NOR2xp33_ASAP7_75t_L g560 ( 
.A(n_471),
.B(n_421),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_L g561 ( 
.A(n_497),
.B(n_425),
.Y(n_561)
);

AOI22xp33_ASAP7_75t_L g562 ( 
.A1(n_441),
.A2(n_317),
.B1(n_207),
.B2(n_314),
.Y(n_562)
);

INVx2_ASAP7_75t_L g563 ( 
.A(n_502),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_L g564 ( 
.A(n_497),
.B(n_426),
.Y(n_564)
);

NAND3xp33_ASAP7_75t_L g565 ( 
.A(n_481),
.B(n_440),
.C(n_384),
.Y(n_565)
);

INVx2_ASAP7_75t_L g566 ( 
.A(n_503),
.Y(n_566)
);

BUFx6f_ASAP7_75t_L g567 ( 
.A(n_503),
.Y(n_567)
);

INVx2_ASAP7_75t_L g568 ( 
.A(n_503),
.Y(n_568)
);

AND3x2_ASAP7_75t_L g569 ( 
.A(n_490),
.B(n_496),
.C(n_489),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_L g570 ( 
.A(n_497),
.B(n_438),
.Y(n_570)
);

NOR2xp33_ASAP7_75t_SL g571 ( 
.A(n_515),
.B(n_354),
.Y(n_571)
);

INVx4_ASAP7_75t_L g572 ( 
.A(n_481),
.Y(n_572)
);

AND2x2_ASAP7_75t_L g573 ( 
.A(n_467),
.B(n_448),
.Y(n_573)
);

INVx2_ASAP7_75t_L g574 ( 
.A(n_503),
.Y(n_574)
);

NOR2xp33_ASAP7_75t_SL g575 ( 
.A(n_515),
.B(n_360),
.Y(n_575)
);

INVx4_ASAP7_75t_L g576 ( 
.A(n_481),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_L g577 ( 
.A(n_497),
.B(n_276),
.Y(n_577)
);

INVx3_ASAP7_75t_L g578 ( 
.A(n_503),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_SL g579 ( 
.A(n_481),
.B(n_353),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_503),
.Y(n_580)
);

INVx2_ASAP7_75t_L g581 ( 
.A(n_509),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_509),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_509),
.Y(n_583)
);

INVx2_ASAP7_75t_SL g584 ( 
.A(n_485),
.Y(n_584)
);

INVx4_ASAP7_75t_L g585 ( 
.A(n_485),
.Y(n_585)
);

INVx3_ASAP7_75t_L g586 ( 
.A(n_509),
.Y(n_586)
);

AND2x2_ASAP7_75t_L g587 ( 
.A(n_467),
.B(n_448),
.Y(n_587)
);

AOI22xp5_ASAP7_75t_L g588 ( 
.A1(n_506),
.A2(n_243),
.B1(n_352),
.B2(n_269),
.Y(n_588)
);

AOI22xp5_ASAP7_75t_L g589 ( 
.A1(n_506),
.A2(n_293),
.B1(n_265),
.B2(n_229),
.Y(n_589)
);

OAI22xp5_ASAP7_75t_L g590 ( 
.A1(n_485),
.A2(n_302),
.B1(n_227),
.B2(n_226),
.Y(n_590)
);

OAI21xp33_ASAP7_75t_SL g591 ( 
.A1(n_486),
.A2(n_204),
.B(n_200),
.Y(n_591)
);

INVx2_ASAP7_75t_L g592 ( 
.A(n_509),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_SL g593 ( 
.A(n_485),
.B(n_362),
.Y(n_593)
);

INVxp67_ASAP7_75t_SL g594 ( 
.A(n_485),
.Y(n_594)
);

BUFx6f_ASAP7_75t_L g595 ( 
.A(n_509),
.Y(n_595)
);

BUFx2_ASAP7_75t_L g596 ( 
.A(n_490),
.Y(n_596)
);

NAND3xp33_ASAP7_75t_L g597 ( 
.A(n_485),
.B(n_244),
.C(n_242),
.Y(n_597)
);

NAND2xp33_ASAP7_75t_L g598 ( 
.A(n_516),
.B(n_214),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_516),
.Y(n_599)
);

BUFx2_ASAP7_75t_L g600 ( 
.A(n_496),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_516),
.Y(n_601)
);

AND2x2_ASAP7_75t_L g602 ( 
.A(n_452),
.B(n_233),
.Y(n_602)
);

INVx2_ASAP7_75t_L g603 ( 
.A(n_516),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_516),
.Y(n_604)
);

INVx6_ASAP7_75t_L g605 ( 
.A(n_486),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_L g606 ( 
.A(n_486),
.B(n_276),
.Y(n_606)
);

INVx2_ASAP7_75t_SL g607 ( 
.A(n_452),
.Y(n_607)
);

INVx2_ASAP7_75t_L g608 ( 
.A(n_516),
.Y(n_608)
);

BUFx6f_ASAP7_75t_L g609 ( 
.A(n_454),
.Y(n_609)
);

BUFx3_ASAP7_75t_L g610 ( 
.A(n_515),
.Y(n_610)
);

CKINVDCx5p33_ASAP7_75t_R g611 ( 
.A(n_510),
.Y(n_611)
);

INVx3_ASAP7_75t_L g612 ( 
.A(n_463),
.Y(n_612)
);

INVx4_ASAP7_75t_L g613 ( 
.A(n_510),
.Y(n_613)
);

INVx2_ASAP7_75t_L g614 ( 
.A(n_454),
.Y(n_614)
);

AND2x2_ASAP7_75t_SL g615 ( 
.A(n_441),
.B(n_183),
.Y(n_615)
);

AND2x6_ASAP7_75t_L g616 ( 
.A(n_449),
.B(n_183),
.Y(n_616)
);

INVx2_ASAP7_75t_SL g617 ( 
.A(n_506),
.Y(n_617)
);

NAND2xp33_ASAP7_75t_SL g618 ( 
.A(n_460),
.B(n_408),
.Y(n_618)
);

AOI22xp33_ASAP7_75t_L g619 ( 
.A1(n_441),
.A2(n_506),
.B1(n_466),
.B2(n_460),
.Y(n_619)
);

BUFx6f_ASAP7_75t_L g620 ( 
.A(n_454),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_451),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_451),
.Y(n_622)
);

AOI22xp5_ASAP7_75t_L g623 ( 
.A1(n_463),
.A2(n_306),
.B1(n_310),
.B2(n_309),
.Y(n_623)
);

NOR2xp33_ASAP7_75t_R g624 ( 
.A(n_499),
.B(n_365),
.Y(n_624)
);

INVx4_ASAP7_75t_L g625 ( 
.A(n_510),
.Y(n_625)
);

INVx2_ASAP7_75t_L g626 ( 
.A(n_454),
.Y(n_626)
);

INVx4_ASAP7_75t_L g627 ( 
.A(n_510),
.Y(n_627)
);

OAI22xp33_ASAP7_75t_L g628 ( 
.A1(n_468),
.A2(n_286),
.B1(n_245),
.B2(n_256),
.Y(n_628)
);

NOR2xp33_ASAP7_75t_L g629 ( 
.A(n_464),
.B(n_469),
.Y(n_629)
);

INVx2_ASAP7_75t_L g630 ( 
.A(n_454),
.Y(n_630)
);

NOR2xp33_ASAP7_75t_L g631 ( 
.A(n_464),
.B(n_434),
.Y(n_631)
);

BUFx6f_ASAP7_75t_SL g632 ( 
.A(n_469),
.Y(n_632)
);

INVx2_ASAP7_75t_L g633 ( 
.A(n_454),
.Y(n_633)
);

NAND3xp33_ASAP7_75t_L g634 ( 
.A(n_466),
.B(n_275),
.C(n_267),
.Y(n_634)
);

INVx2_ASAP7_75t_L g635 ( 
.A(n_463),
.Y(n_635)
);

INVx3_ASAP7_75t_L g636 ( 
.A(n_465),
.Y(n_636)
);

CKINVDCx16_ASAP7_75t_R g637 ( 
.A(n_470),
.Y(n_637)
);

INVx2_ASAP7_75t_SL g638 ( 
.A(n_510),
.Y(n_638)
);

INVx5_ASAP7_75t_L g639 ( 
.A(n_443),
.Y(n_639)
);

AOI22xp5_ASAP7_75t_L g640 ( 
.A1(n_465),
.A2(n_308),
.B1(n_277),
.B2(n_349),
.Y(n_640)
);

AND2x6_ASAP7_75t_L g641 ( 
.A(n_453),
.B(n_183),
.Y(n_641)
);

INVx2_ASAP7_75t_L g642 ( 
.A(n_465),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_SL g643 ( 
.A(n_470),
.B(n_233),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_453),
.Y(n_644)
);

AOI22xp33_ASAP7_75t_L g645 ( 
.A1(n_441),
.A2(n_207),
.B1(n_350),
.B2(n_326),
.Y(n_645)
);

INVx2_ASAP7_75t_L g646 ( 
.A(n_477),
.Y(n_646)
);

INVx3_ASAP7_75t_L g647 ( 
.A(n_477),
.Y(n_647)
);

INVx1_ASAP7_75t_SL g648 ( 
.A(n_468),
.Y(n_648)
);

AOI22xp33_ASAP7_75t_L g649 ( 
.A1(n_473),
.A2(n_285),
.B1(n_350),
.B2(n_326),
.Y(n_649)
);

BUFx3_ASAP7_75t_L g650 ( 
.A(n_473),
.Y(n_650)
);

BUFx2_ASAP7_75t_L g651 ( 
.A(n_474),
.Y(n_651)
);

NOR2x1p5_ASAP7_75t_L g652 ( 
.A(n_478),
.B(n_204),
.Y(n_652)
);

INVx1_ASAP7_75t_SL g653 ( 
.A(n_478),
.Y(n_653)
);

INVx2_ASAP7_75t_L g654 ( 
.A(n_477),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_L g655 ( 
.A(n_474),
.B(n_276),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_487),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_L g657 ( 
.A(n_476),
.B(n_324),
.Y(n_657)
);

INVx2_ASAP7_75t_L g658 ( 
.A(n_487),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_487),
.Y(n_659)
);

NOR3xp33_ASAP7_75t_L g660 ( 
.A(n_480),
.B(n_210),
.C(n_208),
.Y(n_660)
);

INVx1_ASAP7_75t_SL g661 ( 
.A(n_480),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_SL g662 ( 
.A(n_476),
.B(n_280),
.Y(n_662)
);

NOR2xp33_ASAP7_75t_L g663 ( 
.A(n_479),
.B(n_427),
.Y(n_663)
);

HB1xp67_ASAP7_75t_L g664 ( 
.A(n_498),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_SL g665 ( 
.A(n_479),
.B(n_482),
.Y(n_665)
);

NOR2xp33_ASAP7_75t_SL g666 ( 
.A(n_510),
.B(n_363),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_L g667 ( 
.A(n_482),
.B(n_488),
.Y(n_667)
);

OR2x6_ASAP7_75t_L g668 ( 
.A(n_491),
.B(n_208),
.Y(n_668)
);

INVx2_ASAP7_75t_L g669 ( 
.A(n_498),
.Y(n_669)
);

HB1xp67_ASAP7_75t_L g670 ( 
.A(n_525),
.Y(n_670)
);

INVx3_ASAP7_75t_L g671 ( 
.A(n_572),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_SL g672 ( 
.A(n_543),
.B(n_510),
.Y(n_672)
);

AOI22xp33_ASAP7_75t_L g673 ( 
.A1(n_668),
.A2(n_517),
.B1(n_514),
.B2(n_511),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_L g674 ( 
.A(n_648),
.B(n_488),
.Y(n_674)
);

INVx2_ASAP7_75t_L g675 ( 
.A(n_519),
.Y(n_675)
);

INVx2_ASAP7_75t_SL g676 ( 
.A(n_525),
.Y(n_676)
);

BUFx6f_ASAP7_75t_L g677 ( 
.A(n_567),
.Y(n_677)
);

AOI22xp5_ASAP7_75t_L g678 ( 
.A1(n_528),
.A2(n_517),
.B1(n_514),
.B2(n_511),
.Y(n_678)
);

AOI22xp33_ASAP7_75t_L g679 ( 
.A1(n_668),
.A2(n_508),
.B1(n_493),
.B2(n_505),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_SL g680 ( 
.A(n_572),
.B(n_493),
.Y(n_680)
);

BUFx8_ASAP7_75t_L g681 ( 
.A(n_632),
.Y(n_681)
);

INVx3_ASAP7_75t_L g682 ( 
.A(n_572),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_L g683 ( 
.A(n_653),
.B(n_500),
.Y(n_683)
);

OAI22xp5_ASAP7_75t_L g684 ( 
.A1(n_528),
.A2(n_508),
.B1(n_500),
.B2(n_505),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_SL g685 ( 
.A(n_576),
.B(n_498),
.Y(n_685)
);

OAI221xp5_ASAP7_75t_L g686 ( 
.A1(n_520),
.A2(n_272),
.B1(n_210),
.B2(n_319),
.C(n_314),
.Y(n_686)
);

INVx2_ASAP7_75t_L g687 ( 
.A(n_519),
.Y(n_687)
);

INVxp67_ASAP7_75t_L g688 ( 
.A(n_596),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_L g689 ( 
.A(n_661),
.B(n_501),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_621),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_SL g691 ( 
.A(n_576),
.B(n_501),
.Y(n_691)
);

INVxp33_ASAP7_75t_L g692 ( 
.A(n_522),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_621),
.Y(n_693)
);

NOR2xp67_ASAP7_75t_L g694 ( 
.A(n_537),
.B(n_501),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_L g695 ( 
.A(n_518),
.B(n_491),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_622),
.Y(n_696)
);

NAND2xp33_ASAP7_75t_L g697 ( 
.A(n_584),
.B(n_214),
.Y(n_697)
);

INVx2_ASAP7_75t_L g698 ( 
.A(n_524),
.Y(n_698)
);

INVx2_ASAP7_75t_L g699 ( 
.A(n_524),
.Y(n_699)
);

INVx2_ASAP7_75t_L g700 ( 
.A(n_529),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_L g701 ( 
.A(n_542),
.B(n_494),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_622),
.Y(n_702)
);

AND2x2_ASAP7_75t_L g703 ( 
.A(n_637),
.B(n_364),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_644),
.Y(n_704)
);

INVx2_ASAP7_75t_L g705 ( 
.A(n_529),
.Y(n_705)
);

INVxp67_ASAP7_75t_L g706 ( 
.A(n_596),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_644),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_SL g708 ( 
.A(n_576),
.B(n_585),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_L g709 ( 
.A(n_531),
.B(n_494),
.Y(n_709)
);

O2A1O1Ixp5_ASAP7_75t_L g710 ( 
.A1(n_665),
.A2(n_456),
.B(n_495),
.C(n_507),
.Y(n_710)
);

NOR2xp33_ASAP7_75t_L g711 ( 
.A(n_546),
.B(n_495),
.Y(n_711)
);

NOR2xp33_ASAP7_75t_L g712 ( 
.A(n_551),
.B(n_507),
.Y(n_712)
);

INVxp67_ASAP7_75t_SL g713 ( 
.A(n_584),
.Y(n_713)
);

OAI22xp33_ASAP7_75t_L g714 ( 
.A1(n_528),
.A2(n_456),
.B1(n_221),
.B2(n_238),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_L g715 ( 
.A(n_573),
.B(n_324),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_650),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_SL g717 ( 
.A(n_585),
.B(n_330),
.Y(n_717)
);

INVx2_ASAP7_75t_L g718 ( 
.A(n_635),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_L g719 ( 
.A(n_573),
.B(n_330),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_L g720 ( 
.A(n_587),
.B(n_340),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_650),
.Y(n_721)
);

INVx2_ASAP7_75t_L g722 ( 
.A(n_635),
.Y(n_722)
);

NOR2xp33_ASAP7_75t_L g723 ( 
.A(n_532),
.B(n_284),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_L g724 ( 
.A(n_587),
.B(n_340),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_L g725 ( 
.A(n_548),
.B(n_341),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_L g726 ( 
.A(n_548),
.B(n_341),
.Y(n_726)
);

AOI22xp5_ASAP7_75t_L g727 ( 
.A1(n_528),
.A2(n_347),
.B1(n_351),
.B2(n_177),
.Y(n_727)
);

INVxp67_ASAP7_75t_SL g728 ( 
.A(n_538),
.Y(n_728)
);

INVx2_ASAP7_75t_L g729 ( 
.A(n_642),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_L g730 ( 
.A(n_651),
.B(n_347),
.Y(n_730)
);

BUFx3_ASAP7_75t_L g731 ( 
.A(n_536),
.Y(n_731)
);

A2O1A1Ixp33_ASAP7_75t_L g732 ( 
.A1(n_591),
.A2(n_246),
.B(n_292),
.C(n_287),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_SL g733 ( 
.A(n_585),
.B(n_351),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_664),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_L g735 ( 
.A(n_651),
.B(n_221),
.Y(n_735)
);

INVx3_ASAP7_75t_L g736 ( 
.A(n_550),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_SL g737 ( 
.A(n_637),
.B(n_177),
.Y(n_737)
);

NAND2xp33_ASAP7_75t_L g738 ( 
.A(n_616),
.B(n_290),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_L g739 ( 
.A(n_570),
.B(n_238),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_SL g740 ( 
.A(n_567),
.B(n_595),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_L g741 ( 
.A(n_602),
.B(n_246),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_667),
.Y(n_742)
);

NAND2xp33_ASAP7_75t_L g743 ( 
.A(n_616),
.B(n_299),
.Y(n_743)
);

INVx2_ASAP7_75t_L g744 ( 
.A(n_642),
.Y(n_744)
);

AND2x2_ASAP7_75t_L g745 ( 
.A(n_600),
.B(n_272),
.Y(n_745)
);

AOI22xp5_ASAP7_75t_L g746 ( 
.A1(n_521),
.A2(n_184),
.B1(n_295),
.B2(n_237),
.Y(n_746)
);

AOI22xp33_ASAP7_75t_L g747 ( 
.A1(n_668),
.A2(n_184),
.B1(n_224),
.B2(n_334),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_L g748 ( 
.A(n_602),
.B(n_545),
.Y(n_748)
);

INVx2_ASAP7_75t_L g749 ( 
.A(n_646),
.Y(n_749)
);

AND2x2_ASAP7_75t_SL g750 ( 
.A(n_544),
.B(n_224),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_SL g751 ( 
.A(n_567),
.B(n_224),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_L g752 ( 
.A(n_547),
.B(n_285),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_656),
.Y(n_753)
);

BUFx5_ASAP7_75t_L g754 ( 
.A(n_615),
.Y(n_754)
);

INVx2_ASAP7_75t_L g755 ( 
.A(n_646),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_SL g756 ( 
.A(n_567),
.B(n_257),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_L g757 ( 
.A(n_617),
.B(n_287),
.Y(n_757)
);

NAND3xp33_ASAP7_75t_L g758 ( 
.A(n_631),
.B(n_342),
.C(n_328),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_L g759 ( 
.A(n_617),
.B(n_292),
.Y(n_759)
);

NAND2xp33_ASAP7_75t_L g760 ( 
.A(n_616),
.B(n_641),
.Y(n_760)
);

INVx2_ASAP7_75t_L g761 ( 
.A(n_654),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_L g762 ( 
.A(n_561),
.B(n_301),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_656),
.Y(n_763)
);

INVx3_ASAP7_75t_L g764 ( 
.A(n_550),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_SL g765 ( 
.A(n_567),
.B(n_257),
.Y(n_765)
);

AOI221xp5_ASAP7_75t_L g766 ( 
.A1(n_559),
.A2(n_319),
.B1(n_323),
.B2(n_313),
.C(n_301),
.Y(n_766)
);

AOI22xp33_ASAP7_75t_L g767 ( 
.A1(n_668),
.A2(n_334),
.B1(n_257),
.B2(n_323),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_L g768 ( 
.A(n_564),
.B(n_607),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_L g769 ( 
.A(n_607),
.B(n_313),
.Y(n_769)
);

O2A1O1Ixp33_ASAP7_75t_L g770 ( 
.A1(n_591),
.A2(n_442),
.B(n_334),
.C(n_234),
.Y(n_770)
);

NOR2xp67_ASAP7_75t_SL g771 ( 
.A(n_550),
.B(n_605),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_L g772 ( 
.A(n_629),
.B(n_307),
.Y(n_772)
);

OAI22x1_ASAP7_75t_R g773 ( 
.A1(n_527),
.A2(n_315),
.B1(n_316),
.B2(n_318),
.Y(n_773)
);

NOR2xp33_ASAP7_75t_L g774 ( 
.A(n_663),
.B(n_554),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_SL g775 ( 
.A(n_595),
.B(n_234),
.Y(n_775)
);

NOR2xp33_ASAP7_75t_SL g776 ( 
.A(n_575),
.B(n_331),
.Y(n_776)
);

INVxp67_ASAP7_75t_L g777 ( 
.A(n_600),
.Y(n_777)
);

O2A1O1Ixp5_ASAP7_75t_L g778 ( 
.A1(n_594),
.A2(n_442),
.B(n_447),
.C(n_248),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_659),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_659),
.Y(n_780)
);

INVx2_ASAP7_75t_L g781 ( 
.A(n_654),
.Y(n_781)
);

NOR2xp67_ASAP7_75t_L g782 ( 
.A(n_536),
.B(n_442),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_L g783 ( 
.A(n_555),
.B(n_336),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_L g784 ( 
.A(n_553),
.B(n_337),
.Y(n_784)
);

INVx2_ASAP7_75t_L g785 ( 
.A(n_658),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_SL g786 ( 
.A(n_595),
.B(n_248),
.Y(n_786)
);

AOI22xp33_ASAP7_75t_L g787 ( 
.A1(n_615),
.A2(n_338),
.B1(n_343),
.B2(n_344),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_SL g788 ( 
.A(n_595),
.B(n_443),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_L g789 ( 
.A(n_652),
.B(n_179),
.Y(n_789)
);

NOR3xp33_ASAP7_75t_L g790 ( 
.A(n_628),
.B(n_442),
.C(n_205),
.Y(n_790)
);

NAND3xp33_ASAP7_75t_L g791 ( 
.A(n_559),
.B(n_268),
.C(n_190),
.Y(n_791)
);

INVx2_ASAP7_75t_SL g792 ( 
.A(n_569),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_L g793 ( 
.A(n_652),
.B(n_188),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_SL g794 ( 
.A(n_595),
.B(n_615),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_L g795 ( 
.A(n_523),
.B(n_550),
.Y(n_795)
);

AOI22xp5_ASAP7_75t_SL g796 ( 
.A1(n_522),
.A2(n_335),
.B1(n_196),
.B2(n_194),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_612),
.Y(n_797)
);

INVx2_ASAP7_75t_L g798 ( 
.A(n_658),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_612),
.Y(n_799)
);

INVx2_ASAP7_75t_SL g800 ( 
.A(n_605),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_612),
.Y(n_801)
);

O2A1O1Ixp33_ASAP7_75t_L g802 ( 
.A1(n_657),
.A2(n_447),
.B(n_16),
.C(n_19),
.Y(n_802)
);

NOR2xp33_ASAP7_75t_L g803 ( 
.A(n_560),
.B(n_192),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_SL g804 ( 
.A(n_619),
.B(n_443),
.Y(n_804)
);

INVx2_ASAP7_75t_L g805 ( 
.A(n_669),
.Y(n_805)
);

CKINVDCx5p33_ASAP7_75t_R g806 ( 
.A(n_527),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_636),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_SL g808 ( 
.A(n_636),
.B(n_443),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_SL g809 ( 
.A(n_636),
.B(n_443),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_L g810 ( 
.A(n_605),
.B(n_193),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_SL g811 ( 
.A(n_647),
.B(n_443),
.Y(n_811)
);

INVx2_ASAP7_75t_L g812 ( 
.A(n_669),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_L g813 ( 
.A(n_605),
.B(n_647),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_L g814 ( 
.A(n_647),
.B(n_197),
.Y(n_814)
);

AND2x4_ASAP7_75t_L g815 ( 
.A(n_610),
.B(n_15),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_L g816 ( 
.A(n_521),
.B(n_549),
.Y(n_816)
);

NOR2xp33_ASAP7_75t_L g817 ( 
.A(n_593),
.B(n_198),
.Y(n_817)
);

AND2x4_ASAP7_75t_SL g818 ( 
.A(n_558),
.B(n_447),
.Y(n_818)
);

AOI22xp5_ASAP7_75t_L g819 ( 
.A1(n_521),
.A2(n_288),
.B1(n_209),
.B2(n_348),
.Y(n_819)
);

O2A1O1Ixp33_ASAP7_75t_L g820 ( 
.A1(n_660),
.A2(n_20),
.B(n_21),
.C(n_23),
.Y(n_820)
);

NAND2x1p5_ASAP7_75t_L g821 ( 
.A(n_610),
.B(n_446),
.Y(n_821)
);

AOI22xp33_ASAP7_75t_L g822 ( 
.A1(n_521),
.A2(n_289),
.B1(n_213),
.B2(n_345),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_L g823 ( 
.A(n_549),
.B(n_283),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_L g824 ( 
.A(n_655),
.B(n_297),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_SL g825 ( 
.A(n_578),
.B(n_450),
.Y(n_825)
);

INVx2_ASAP7_75t_L g826 ( 
.A(n_533),
.Y(n_826)
);

NAND2xp33_ASAP7_75t_L g827 ( 
.A(n_616),
.B(n_279),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_533),
.Y(n_828)
);

INVx2_ASAP7_75t_L g829 ( 
.A(n_535),
.Y(n_829)
);

O2A1O1Ixp33_ASAP7_75t_L g830 ( 
.A1(n_577),
.A2(n_21),
.B(n_23),
.C(n_24),
.Y(n_830)
);

NOR3xp33_ASAP7_75t_L g831 ( 
.A(n_579),
.B(n_202),
.C(n_236),
.Y(n_831)
);

AND2x4_ASAP7_75t_L g832 ( 
.A(n_565),
.B(n_24),
.Y(n_832)
);

AOI22xp5_ASAP7_75t_L g833 ( 
.A1(n_632),
.A2(n_304),
.B1(n_241),
.B2(n_339),
.Y(n_833)
);

INVx2_ASAP7_75t_L g834 ( 
.A(n_535),
.Y(n_834)
);

INVx2_ASAP7_75t_L g835 ( 
.A(n_539),
.Y(n_835)
);

AND2x4_ASAP7_75t_L g836 ( 
.A(n_634),
.B(n_25),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_539),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_L g838 ( 
.A(n_588),
.B(n_303),
.Y(n_838)
);

INVx2_ASAP7_75t_L g839 ( 
.A(n_541),
.Y(n_839)
);

NOR2xp33_ASAP7_75t_L g840 ( 
.A(n_643),
.B(n_662),
.Y(n_840)
);

AOI22xp33_ASAP7_75t_L g841 ( 
.A1(n_750),
.A2(n_645),
.B1(n_562),
.B2(n_641),
.Y(n_841)
);

AOI21xp5_ASAP7_75t_L g842 ( 
.A1(n_709),
.A2(n_606),
.B(n_530),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_L g843 ( 
.A(n_695),
.B(n_588),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_L g844 ( 
.A(n_774),
.B(n_589),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_L g845 ( 
.A(n_711),
.B(n_589),
.Y(n_845)
);

NOR2xp67_ASAP7_75t_L g846 ( 
.A(n_712),
.B(n_526),
.Y(n_846)
);

BUFx12f_ASAP7_75t_L g847 ( 
.A(n_806),
.Y(n_847)
);

OAI21xp33_ASAP7_75t_L g848 ( 
.A1(n_803),
.A2(n_623),
.B(n_640),
.Y(n_848)
);

HB1xp67_ASAP7_75t_L g849 ( 
.A(n_670),
.Y(n_849)
);

INVx1_ASAP7_75t_SL g850 ( 
.A(n_676),
.Y(n_850)
);

INVx2_ASAP7_75t_L g851 ( 
.A(n_675),
.Y(n_851)
);

INVx2_ASAP7_75t_L g852 ( 
.A(n_675),
.Y(n_852)
);

NAND2xp5_ASAP7_75t_SL g853 ( 
.A(n_815),
.B(n_624),
.Y(n_853)
);

INVx2_ASAP7_75t_L g854 ( 
.A(n_687),
.Y(n_854)
);

NOR2xp33_ASAP7_75t_L g855 ( 
.A(n_701),
.B(n_666),
.Y(n_855)
);

OAI21xp33_ASAP7_75t_L g856 ( 
.A1(n_772),
.A2(n_640),
.B(n_623),
.Y(n_856)
);

O2A1O1Ixp33_ASAP7_75t_SL g857 ( 
.A1(n_672),
.A2(n_534),
.B(n_540),
.C(n_604),
.Y(n_857)
);

OAI21xp5_ASAP7_75t_L g858 ( 
.A1(n_778),
.A2(n_710),
.B(n_672),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_L g859 ( 
.A(n_742),
.B(n_557),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_L g860 ( 
.A(n_689),
.B(n_590),
.Y(n_860)
);

NAND2x1_ASAP7_75t_L g861 ( 
.A(n_771),
.B(n_578),
.Y(n_861)
);

NAND2xp33_ASAP7_75t_L g862 ( 
.A(n_754),
.B(n_800),
.Y(n_862)
);

AOI21xp5_ASAP7_75t_L g863 ( 
.A1(n_813),
.A2(n_583),
.B(n_540),
.Y(n_863)
);

AND2x2_ASAP7_75t_L g864 ( 
.A(n_745),
.B(n_558),
.Y(n_864)
);

AOI21xp5_ASAP7_75t_L g865 ( 
.A1(n_740),
.A2(n_599),
.B(n_580),
.Y(n_865)
);

AOI21xp5_ASAP7_75t_L g866 ( 
.A1(n_740),
.A2(n_599),
.B(n_580),
.Y(n_866)
);

NOR2xp33_ASAP7_75t_L g867 ( 
.A(n_748),
.B(n_632),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_L g868 ( 
.A(n_674),
.B(n_683),
.Y(n_868)
);

BUFx2_ASAP7_75t_L g869 ( 
.A(n_703),
.Y(n_869)
);

AOI21x1_ASAP7_75t_L g870 ( 
.A1(n_804),
.A2(n_601),
.B(n_530),
.Y(n_870)
);

O2A1O1Ixp33_ASAP7_75t_L g871 ( 
.A1(n_732),
.A2(n_586),
.B(n_578),
.C(n_534),
.Y(n_871)
);

OAI22xp5_ASAP7_75t_L g872 ( 
.A1(n_678),
.A2(n_597),
.B1(n_586),
.B2(n_601),
.Y(n_872)
);

INVx1_ASAP7_75t_L g873 ( 
.A(n_690),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_SL g874 ( 
.A(n_815),
.B(n_571),
.Y(n_874)
);

AOI21xp5_ASAP7_75t_L g875 ( 
.A1(n_708),
.A2(n_604),
.B(n_582),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_L g876 ( 
.A(n_768),
.B(n_649),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_SL g877 ( 
.A(n_754),
.B(n_586),
.Y(n_877)
);

AO21x2_ASAP7_75t_L g878 ( 
.A1(n_804),
.A2(n_583),
.B(n_582),
.Y(n_878)
);

AOI21xp5_ASAP7_75t_L g879 ( 
.A1(n_708),
.A2(n_592),
.B(n_566),
.Y(n_879)
);

NOR2xp33_ASAP7_75t_L g880 ( 
.A(n_737),
.B(n_618),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_L g881 ( 
.A(n_715),
.B(n_616),
.Y(n_881)
);

OAI22xp5_ASAP7_75t_L g882 ( 
.A1(n_693),
.A2(n_581),
.B1(n_563),
.B2(n_566),
.Y(n_882)
);

BUFx6f_ASAP7_75t_L g883 ( 
.A(n_677),
.Y(n_883)
);

AOI22xp5_ASAP7_75t_L g884 ( 
.A1(n_754),
.A2(n_616),
.B1(n_641),
.B2(n_592),
.Y(n_884)
);

O2A1O1Ixp5_ASAP7_75t_L g885 ( 
.A1(n_680),
.A2(n_762),
.B(n_733),
.C(n_717),
.Y(n_885)
);

HB1xp67_ASAP7_75t_L g886 ( 
.A(n_688),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_SL g887 ( 
.A(n_754),
.B(n_816),
.Y(n_887)
);

AOI21xp5_ASAP7_75t_L g888 ( 
.A1(n_685),
.A2(n_556),
.B(n_563),
.Y(n_888)
);

AOI21xp5_ASAP7_75t_L g889 ( 
.A1(n_685),
.A2(n_691),
.B(n_810),
.Y(n_889)
);

AND2x2_ASAP7_75t_L g890 ( 
.A(n_706),
.B(n_541),
.Y(n_890)
);

BUFx8_ASAP7_75t_SL g891 ( 
.A(n_815),
.Y(n_891)
);

OAI22xp5_ASAP7_75t_L g892 ( 
.A1(n_696),
.A2(n_704),
.B1(n_707),
.B2(n_702),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_L g893 ( 
.A(n_719),
.B(n_616),
.Y(n_893)
);

AO21x1_ASAP7_75t_L g894 ( 
.A1(n_794),
.A2(n_684),
.B(n_775),
.Y(n_894)
);

AOI21xp5_ASAP7_75t_L g895 ( 
.A1(n_691),
.A2(n_680),
.B(n_825),
.Y(n_895)
);

NAND2xp5_ASAP7_75t_L g896 ( 
.A(n_720),
.B(n_641),
.Y(n_896)
);

NOR3xp33_ASAP7_75t_L g897 ( 
.A(n_686),
.B(n_598),
.C(n_552),
.Y(n_897)
);

AOI21xp5_ASAP7_75t_L g898 ( 
.A1(n_825),
.A2(n_556),
.B(n_568),
.Y(n_898)
);

NAND2xp5_ASAP7_75t_L g899 ( 
.A(n_724),
.B(n_641),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_L g900 ( 
.A(n_750),
.B(n_641),
.Y(n_900)
);

INVx1_ASAP7_75t_L g901 ( 
.A(n_734),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_L g902 ( 
.A(n_730),
.B(n_641),
.Y(n_902)
);

INVx1_ASAP7_75t_L g903 ( 
.A(n_753),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_L g904 ( 
.A(n_741),
.B(n_552),
.Y(n_904)
);

BUFx8_ASAP7_75t_L g905 ( 
.A(n_792),
.Y(n_905)
);

AOI21xp5_ASAP7_75t_L g906 ( 
.A1(n_713),
.A2(n_603),
.B(n_581),
.Y(n_906)
);

BUFx6f_ASAP7_75t_L g907 ( 
.A(n_677),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_763),
.Y(n_908)
);

INVx1_ASAP7_75t_L g909 ( 
.A(n_779),
.Y(n_909)
);

AO21x1_ASAP7_75t_L g910 ( 
.A1(n_794),
.A2(n_574),
.B(n_603),
.Y(n_910)
);

NAND2xp5_ASAP7_75t_SL g911 ( 
.A(n_754),
.B(n_568),
.Y(n_911)
);

NOR2xp67_ASAP7_75t_L g912 ( 
.A(n_777),
.B(n_574),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_SL g913 ( 
.A(n_754),
.B(n_608),
.Y(n_913)
);

INVx1_ASAP7_75t_SL g914 ( 
.A(n_818),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_L g915 ( 
.A(n_694),
.B(n_608),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_780),
.Y(n_916)
);

INVx4_ASAP7_75t_L g917 ( 
.A(n_731),
.Y(n_917)
);

INVx1_ASAP7_75t_L g918 ( 
.A(n_828),
.Y(n_918)
);

OAI21xp5_ASAP7_75t_L g919 ( 
.A1(n_826),
.A2(n_626),
.B(n_614),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_L g920 ( 
.A(n_673),
.B(n_679),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_837),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_L g922 ( 
.A(n_725),
.B(n_611),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_826),
.Y(n_923)
);

OAI22xp5_ASAP7_75t_L g924 ( 
.A1(n_800),
.A2(n_795),
.B1(n_736),
.B2(n_764),
.Y(n_924)
);

INVx3_ASAP7_75t_L g925 ( 
.A(n_736),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_SL g926 ( 
.A(n_754),
.B(n_611),
.Y(n_926)
);

A2O1A1Ixp33_ASAP7_75t_L g927 ( 
.A1(n_723),
.A2(n_638),
.B(n_633),
.C(n_630),
.Y(n_927)
);

BUFx12f_ASAP7_75t_L g928 ( 
.A(n_681),
.Y(n_928)
);

AOI21xp5_ASAP7_75t_L g929 ( 
.A1(n_808),
.A2(n_638),
.B(n_626),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_L g930 ( 
.A(n_726),
.B(n_633),
.Y(n_930)
);

OR2x2_ASAP7_75t_L g931 ( 
.A(n_735),
.B(n_614),
.Y(n_931)
);

O2A1O1Ixp33_ASAP7_75t_SL g932 ( 
.A1(n_732),
.A2(n_630),
.B(n_639),
.C(n_29),
.Y(n_932)
);

O2A1O1Ixp5_ASAP7_75t_L g933 ( 
.A1(n_717),
.A2(n_613),
.B(n_627),
.C(n_625),
.Y(n_933)
);

OR2x6_ASAP7_75t_L g934 ( 
.A(n_731),
.B(n_613),
.Y(n_934)
);

NAND3xp33_ASAP7_75t_L g935 ( 
.A(n_787),
.B(n_598),
.C(n_609),
.Y(n_935)
);

NOR2xp33_ASAP7_75t_L g936 ( 
.A(n_737),
.B(n_613),
.Y(n_936)
);

AOI21xp5_ASAP7_75t_L g937 ( 
.A1(n_808),
.A2(n_811),
.B(n_809),
.Y(n_937)
);

INVx1_ASAP7_75t_L g938 ( 
.A(n_829),
.Y(n_938)
);

INVx2_ASAP7_75t_L g939 ( 
.A(n_698),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_L g940 ( 
.A(n_783),
.B(n_620),
.Y(n_940)
);

AO21x1_ASAP7_75t_L g941 ( 
.A1(n_775),
.A2(n_627),
.B(n_625),
.Y(n_941)
);

AOI21xp5_ASAP7_75t_L g942 ( 
.A1(n_809),
.A2(n_620),
.B(n_609),
.Y(n_942)
);

AOI21xp5_ASAP7_75t_L g943 ( 
.A1(n_811),
.A2(n_620),
.B(n_609),
.Y(n_943)
);

NOR3xp33_ASAP7_75t_L g944 ( 
.A(n_758),
.B(n_627),
.C(n_625),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_L g945 ( 
.A(n_767),
.B(n_620),
.Y(n_945)
);

OAI22xp5_ASAP7_75t_L g946 ( 
.A1(n_736),
.A2(n_620),
.B1(n_609),
.B2(n_639),
.Y(n_946)
);

AOI21xp5_ASAP7_75t_L g947 ( 
.A1(n_823),
.A2(n_609),
.B(n_639),
.Y(n_947)
);

NAND2x1p5_ASAP7_75t_L g948 ( 
.A(n_764),
.B(n_639),
.Y(n_948)
);

AOI21xp5_ASAP7_75t_L g949 ( 
.A1(n_728),
.A2(n_639),
.B(n_311),
.Y(n_949)
);

INVx1_ASAP7_75t_L g950 ( 
.A(n_829),
.Y(n_950)
);

NOR2xp33_ASAP7_75t_L g951 ( 
.A(n_838),
.B(n_26),
.Y(n_951)
);

INVx1_ASAP7_75t_L g952 ( 
.A(n_834),
.Y(n_952)
);

NAND2xp5_ASAP7_75t_L g953 ( 
.A(n_716),
.B(n_639),
.Y(n_953)
);

O2A1O1Ixp33_ASAP7_75t_L g954 ( 
.A1(n_784),
.A2(n_28),
.B(n_29),
.C(n_31),
.Y(n_954)
);

NAND2xp5_ASAP7_75t_SL g955 ( 
.A(n_714),
.B(n_263),
.Y(n_955)
);

AOI21xp5_ASAP7_75t_L g956 ( 
.A1(n_797),
.A2(n_801),
.B(n_799),
.Y(n_956)
);

AOI21xp33_ASAP7_75t_L g957 ( 
.A1(n_747),
.A2(n_239),
.B(n_253),
.Y(n_957)
);

AOI21xp5_ASAP7_75t_L g958 ( 
.A1(n_807),
.A2(n_327),
.B(n_325),
.Y(n_958)
);

NAND2xp5_ASAP7_75t_SL g959 ( 
.A(n_671),
.B(n_450),
.Y(n_959)
);

NAND2xp5_ASAP7_75t_SL g960 ( 
.A(n_746),
.B(n_260),
.Y(n_960)
);

INVx3_ASAP7_75t_L g961 ( 
.A(n_764),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_L g962 ( 
.A(n_721),
.B(n_739),
.Y(n_962)
);

OAI21xp5_ASAP7_75t_L g963 ( 
.A1(n_834),
.A2(n_450),
.B(n_446),
.Y(n_963)
);

NOR2xp33_ASAP7_75t_L g964 ( 
.A(n_840),
.B(n_28),
.Y(n_964)
);

NAND2xp5_ASAP7_75t_L g965 ( 
.A(n_757),
.B(n_31),
.Y(n_965)
);

O2A1O1Ixp33_ASAP7_75t_L g966 ( 
.A1(n_820),
.A2(n_38),
.B(n_39),
.C(n_40),
.Y(n_966)
);

AOI21xp5_ASAP7_75t_L g967 ( 
.A1(n_788),
.A2(n_450),
.B(n_446),
.Y(n_967)
);

NAND2xp5_ASAP7_75t_L g968 ( 
.A(n_759),
.B(n_38),
.Y(n_968)
);

NAND2xp33_ASAP7_75t_L g969 ( 
.A(n_671),
.B(n_450),
.Y(n_969)
);

AOI22xp5_ASAP7_75t_L g970 ( 
.A1(n_727),
.A2(n_450),
.B1(n_446),
.B2(n_41),
.Y(n_970)
);

AOI21xp5_ASAP7_75t_L g971 ( 
.A1(n_788),
.A2(n_446),
.B(n_99),
.Y(n_971)
);

AND2x2_ASAP7_75t_L g972 ( 
.A(n_796),
.B(n_39),
.Y(n_972)
);

NAND2xp5_ASAP7_75t_L g973 ( 
.A(n_752),
.B(n_40),
.Y(n_973)
);

AND2x2_ASAP7_75t_L g974 ( 
.A(n_818),
.B(n_41),
.Y(n_974)
);

INVxp67_ASAP7_75t_L g975 ( 
.A(n_776),
.Y(n_975)
);

INVx4_ASAP7_75t_L g976 ( 
.A(n_671),
.Y(n_976)
);

NAND2xp5_ASAP7_75t_SL g977 ( 
.A(n_682),
.B(n_446),
.Y(n_977)
);

OAI22xp5_ASAP7_75t_L g978 ( 
.A1(n_682),
.A2(n_45),
.B1(n_49),
.B2(n_51),
.Y(n_978)
);

AOI21xp5_ASAP7_75t_L g979 ( 
.A1(n_814),
.A2(n_106),
.B(n_172),
.Y(n_979)
);

NAND2xp5_ASAP7_75t_SL g980 ( 
.A(n_682),
.B(n_56),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_L g981 ( 
.A(n_769),
.B(n_56),
.Y(n_981)
);

AOI21xp5_ASAP7_75t_L g982 ( 
.A1(n_824),
.A2(n_133),
.B(n_171),
.Y(n_982)
);

NAND2xp5_ASAP7_75t_SL g983 ( 
.A(n_677),
.B(n_61),
.Y(n_983)
);

NAND2xp5_ASAP7_75t_L g984 ( 
.A(n_817),
.B(n_65),
.Y(n_984)
);

AOI21xp5_ASAP7_75t_L g985 ( 
.A1(n_835),
.A2(n_66),
.B(n_70),
.Y(n_985)
);

OAI21xp5_ASAP7_75t_L g986 ( 
.A1(n_835),
.A2(n_72),
.B(n_75),
.Y(n_986)
);

NAND2xp5_ASAP7_75t_L g987 ( 
.A(n_832),
.B(n_76),
.Y(n_987)
);

NAND2xp5_ASAP7_75t_L g988 ( 
.A(n_832),
.B(n_82),
.Y(n_988)
);

OAI22xp33_ASAP7_75t_SL g989 ( 
.A1(n_836),
.A2(n_92),
.B1(n_97),
.B2(n_100),
.Y(n_989)
);

BUFx6f_ASAP7_75t_L g990 ( 
.A(n_677),
.Y(n_990)
);

A2O1A1Ixp33_ASAP7_75t_L g991 ( 
.A1(n_766),
.A2(n_770),
.B(n_832),
.C(n_836),
.Y(n_991)
);

OAI21xp33_ASAP7_75t_L g992 ( 
.A1(n_789),
.A2(n_101),
.B(n_135),
.Y(n_992)
);

AOI21xp5_ASAP7_75t_L g993 ( 
.A1(n_839),
.A2(n_137),
.B(n_142),
.Y(n_993)
);

NAND2xp5_ASAP7_75t_L g994 ( 
.A(n_819),
.B(n_149),
.Y(n_994)
);

INVx2_ASAP7_75t_L g995 ( 
.A(n_699),
.Y(n_995)
);

AOI21xp5_ASAP7_75t_L g996 ( 
.A1(n_839),
.A2(n_150),
.B(n_155),
.Y(n_996)
);

NAND2xp5_ASAP7_75t_L g997 ( 
.A(n_793),
.B(n_158),
.Y(n_997)
);

INVx1_ASAP7_75t_L g998 ( 
.A(n_718),
.Y(n_998)
);

NAND2xp5_ASAP7_75t_SL g999 ( 
.A(n_790),
.B(n_165),
.Y(n_999)
);

INVx3_ASAP7_75t_L g1000 ( 
.A(n_821),
.Y(n_1000)
);

NOR3xp33_ASAP7_75t_L g1001 ( 
.A(n_791),
.B(n_168),
.C(n_173),
.Y(n_1001)
);

AOI21xp5_ASAP7_75t_L g1002 ( 
.A1(n_760),
.A2(n_755),
.B(n_812),
.Y(n_1002)
);

NOR2xp33_ASAP7_75t_L g1003 ( 
.A(n_733),
.B(n_836),
.Y(n_1003)
);

AOI21xp5_ASAP7_75t_L g1004 ( 
.A1(n_760),
.A2(n_761),
.B(n_812),
.Y(n_1004)
);

NAND2x1p5_ASAP7_75t_L g1005 ( 
.A(n_782),
.B(n_761),
.Y(n_1005)
);

NAND2xp5_ASAP7_75t_L g1006 ( 
.A(n_718),
.B(n_749),
.Y(n_1006)
);

AOI21xp5_ASAP7_75t_L g1007 ( 
.A1(n_722),
.A2(n_755),
.B(n_798),
.Y(n_1007)
);

NOR2xp33_ASAP7_75t_SL g1008 ( 
.A(n_692),
.B(n_821),
.Y(n_1008)
);

O2A1O1Ixp33_ASAP7_75t_L g1009 ( 
.A1(n_830),
.A2(n_802),
.B(n_743),
.C(n_738),
.Y(n_1009)
);

AOI22xp5_ASAP7_75t_L g1010 ( 
.A1(n_822),
.A2(n_743),
.B1(n_738),
.B2(n_833),
.Y(n_1010)
);

OAI22xp5_ASAP7_75t_L g1011 ( 
.A1(n_722),
.A2(n_749),
.B1(n_785),
.B2(n_798),
.Y(n_1011)
);

INVx1_ASAP7_75t_L g1012 ( 
.A(n_729),
.Y(n_1012)
);

INVx1_ASAP7_75t_L g1013 ( 
.A(n_729),
.Y(n_1013)
);

BUFx12f_ASAP7_75t_L g1014 ( 
.A(n_773),
.Y(n_1014)
);

AOI21xp5_ASAP7_75t_L g1015 ( 
.A1(n_744),
.A2(n_781),
.B(n_805),
.Y(n_1015)
);

AOI21xp5_ASAP7_75t_L g1016 ( 
.A1(n_744),
.A2(n_781),
.B(n_805),
.Y(n_1016)
);

AOI21xp5_ASAP7_75t_L g1017 ( 
.A1(n_785),
.A2(n_827),
.B(n_700),
.Y(n_1017)
);

NAND2xp5_ASAP7_75t_L g1018 ( 
.A(n_700),
.B(n_705),
.Y(n_1018)
);

OAI22xp5_ASAP7_75t_L g1019 ( 
.A1(n_705),
.A2(n_831),
.B1(n_751),
.B2(n_756),
.Y(n_1019)
);

AOI21xp5_ASAP7_75t_L g1020 ( 
.A1(n_827),
.A2(n_697),
.B(n_751),
.Y(n_1020)
);

A2O1A1Ixp33_ASAP7_75t_L g1021 ( 
.A1(n_697),
.A2(n_756),
.B(n_765),
.C(n_786),
.Y(n_1021)
);

OAI21xp33_ASAP7_75t_L g1022 ( 
.A1(n_765),
.A2(n_543),
.B(n_695),
.Y(n_1022)
);

INVx1_ASAP7_75t_SL g1023 ( 
.A(n_786),
.Y(n_1023)
);

AOI21xp5_ASAP7_75t_L g1024 ( 
.A1(n_709),
.A2(n_549),
.B(n_672),
.Y(n_1024)
);

OAI22xp5_ASAP7_75t_L g1025 ( 
.A1(n_695),
.A2(n_543),
.B1(n_701),
.B2(n_709),
.Y(n_1025)
);

O2A1O1Ixp33_ASAP7_75t_L g1026 ( 
.A1(n_695),
.A2(n_543),
.B(n_774),
.C(n_542),
.Y(n_1026)
);

NAND2xp5_ASAP7_75t_L g1027 ( 
.A(n_695),
.B(n_543),
.Y(n_1027)
);

BUFx6f_ASAP7_75t_SL g1028 ( 
.A(n_917),
.Y(n_1028)
);

BUFx3_ASAP7_75t_L g1029 ( 
.A(n_847),
.Y(n_1029)
);

NOR2xp33_ASAP7_75t_R g1030 ( 
.A(n_928),
.B(n_1014),
.Y(n_1030)
);

OAI22xp5_ASAP7_75t_L g1031 ( 
.A1(n_1027),
.A2(n_1025),
.B1(n_844),
.B2(n_843),
.Y(n_1031)
);

NAND2xp5_ASAP7_75t_L g1032 ( 
.A(n_868),
.B(n_1026),
.Y(n_1032)
);

INVx2_ASAP7_75t_SL g1033 ( 
.A(n_905),
.Y(n_1033)
);

INVx1_ASAP7_75t_L g1034 ( 
.A(n_901),
.Y(n_1034)
);

BUFx6f_ASAP7_75t_L g1035 ( 
.A(n_883),
.Y(n_1035)
);

AOI22xp5_ASAP7_75t_L g1036 ( 
.A1(n_848),
.A2(n_964),
.B1(n_845),
.B2(n_864),
.Y(n_1036)
);

OAI22xp5_ASAP7_75t_L g1037 ( 
.A1(n_964),
.A2(n_856),
.B1(n_991),
.B2(n_984),
.Y(n_1037)
);

AOI22xp33_ASAP7_75t_L g1038 ( 
.A1(n_846),
.A2(n_1003),
.B1(n_859),
.B2(n_869),
.Y(n_1038)
);

NAND2xp5_ASAP7_75t_SL g1039 ( 
.A(n_850),
.B(n_867),
.Y(n_1039)
);

NAND2xp5_ASAP7_75t_L g1040 ( 
.A(n_855),
.B(n_1022),
.Y(n_1040)
);

BUFx4f_ASAP7_75t_L g1041 ( 
.A(n_974),
.Y(n_1041)
);

NOR2xp33_ASAP7_75t_L g1042 ( 
.A(n_886),
.B(n_849),
.Y(n_1042)
);

INVx1_ASAP7_75t_L g1043 ( 
.A(n_873),
.Y(n_1043)
);

INVx1_ASAP7_75t_L g1044 ( 
.A(n_903),
.Y(n_1044)
);

NAND2xp5_ASAP7_75t_L g1045 ( 
.A(n_867),
.B(n_855),
.Y(n_1045)
);

OR2x6_ASAP7_75t_L g1046 ( 
.A(n_874),
.B(n_853),
.Y(n_1046)
);

INVx4_ASAP7_75t_L g1047 ( 
.A(n_917),
.Y(n_1047)
);

NAND2xp5_ASAP7_75t_SL g1048 ( 
.A(n_886),
.B(n_880),
.Y(n_1048)
);

AOI22xp5_ASAP7_75t_L g1049 ( 
.A1(n_951),
.A2(n_880),
.B1(n_1003),
.B2(n_920),
.Y(n_1049)
);

INVx4_ASAP7_75t_L g1050 ( 
.A(n_934),
.Y(n_1050)
);

NAND2xp5_ASAP7_75t_L g1051 ( 
.A(n_975),
.B(n_876),
.Y(n_1051)
);

NAND2xp5_ASAP7_75t_L g1052 ( 
.A(n_975),
.B(n_890),
.Y(n_1052)
);

BUFx12f_ASAP7_75t_L g1053 ( 
.A(n_905),
.Y(n_1053)
);

NAND2xp5_ASAP7_75t_L g1054 ( 
.A(n_962),
.B(n_908),
.Y(n_1054)
);

AOI21xp5_ASAP7_75t_L g1055 ( 
.A1(n_969),
.A2(n_1024),
.B(n_889),
.Y(n_1055)
);

NOR2x1_ASAP7_75t_L g1056 ( 
.A(n_934),
.B(n_912),
.Y(n_1056)
);

BUFx3_ASAP7_75t_L g1057 ( 
.A(n_891),
.Y(n_1057)
);

O2A1O1Ixp33_ASAP7_75t_L g1058 ( 
.A1(n_951),
.A2(n_966),
.B(n_973),
.C(n_980),
.Y(n_1058)
);

BUFx6f_ASAP7_75t_L g1059 ( 
.A(n_883),
.Y(n_1059)
);

OAI21xp5_ASAP7_75t_L g1060 ( 
.A1(n_842),
.A2(n_858),
.B(n_885),
.Y(n_1060)
);

INVx2_ASAP7_75t_L g1061 ( 
.A(n_851),
.Y(n_1061)
);

INVx4_ASAP7_75t_L g1062 ( 
.A(n_934),
.Y(n_1062)
);

BUFx2_ASAP7_75t_L g1063 ( 
.A(n_849),
.Y(n_1063)
);

O2A1O1Ixp5_ASAP7_75t_L g1064 ( 
.A1(n_999),
.A2(n_885),
.B(n_968),
.C(n_965),
.Y(n_1064)
);

AOI21xp5_ASAP7_75t_L g1065 ( 
.A1(n_940),
.A2(n_862),
.B(n_922),
.Y(n_1065)
);

BUFx2_ASAP7_75t_L g1066 ( 
.A(n_972),
.Y(n_1066)
);

AOI21xp5_ASAP7_75t_L g1067 ( 
.A1(n_877),
.A2(n_857),
.B(n_937),
.Y(n_1067)
);

NAND2x1p5_ASAP7_75t_L g1068 ( 
.A(n_1000),
.B(n_914),
.Y(n_1068)
);

INVx2_ASAP7_75t_L g1069 ( 
.A(n_852),
.Y(n_1069)
);

CKINVDCx8_ASAP7_75t_R g1070 ( 
.A(n_883),
.Y(n_1070)
);

INVx1_ASAP7_75t_L g1071 ( 
.A(n_909),
.Y(n_1071)
);

AND2x4_ASAP7_75t_L g1072 ( 
.A(n_916),
.B(n_1000),
.Y(n_1072)
);

NOR2xp33_ASAP7_75t_L g1073 ( 
.A(n_1008),
.B(n_860),
.Y(n_1073)
);

A2O1A1Ixp33_ASAP7_75t_L g1074 ( 
.A1(n_1010),
.A2(n_1009),
.B(n_994),
.C(n_987),
.Y(n_1074)
);

NOR2x1_ASAP7_75t_R g1075 ( 
.A(n_960),
.B(n_983),
.Y(n_1075)
);

A2O1A1Ixp33_ASAP7_75t_L g1076 ( 
.A1(n_988),
.A2(n_896),
.B(n_881),
.C(n_893),
.Y(n_1076)
);

O2A1O1Ixp33_ASAP7_75t_L g1077 ( 
.A1(n_980),
.A2(n_981),
.B(n_983),
.C(n_978),
.Y(n_1077)
);

BUFx2_ASAP7_75t_L g1078 ( 
.A(n_883),
.Y(n_1078)
);

NOR2xp67_ASAP7_75t_L g1079 ( 
.A(n_936),
.B(n_925),
.Y(n_1079)
);

O2A1O1Ixp5_ASAP7_75t_L g1080 ( 
.A1(n_999),
.A2(n_927),
.B(n_997),
.C(n_926),
.Y(n_1080)
);

INVx5_ASAP7_75t_L g1081 ( 
.A(n_907),
.Y(n_1081)
);

AOI22xp5_ASAP7_75t_L g1082 ( 
.A1(n_936),
.A2(n_892),
.B1(n_955),
.B2(n_902),
.Y(n_1082)
);

AND2x4_ASAP7_75t_L g1083 ( 
.A(n_907),
.B(n_990),
.Y(n_1083)
);

BUFx6f_ASAP7_75t_L g1084 ( 
.A(n_907),
.Y(n_1084)
);

INVx1_ASAP7_75t_L g1085 ( 
.A(n_918),
.Y(n_1085)
);

NAND2xp5_ASAP7_75t_L g1086 ( 
.A(n_931),
.B(n_904),
.Y(n_1086)
);

AOI21xp5_ASAP7_75t_L g1087 ( 
.A1(n_877),
.A2(n_977),
.B(n_959),
.Y(n_1087)
);

NOR2xp33_ASAP7_75t_R g1088 ( 
.A(n_990),
.B(n_925),
.Y(n_1088)
);

NAND2xp5_ASAP7_75t_SL g1089 ( 
.A(n_976),
.B(n_990),
.Y(n_1089)
);

NAND2xp5_ASAP7_75t_SL g1090 ( 
.A(n_976),
.B(n_990),
.Y(n_1090)
);

NOR2xp33_ASAP7_75t_R g1091 ( 
.A(n_961),
.B(n_870),
.Y(n_1091)
);

NAND2xp5_ASAP7_75t_SL g1092 ( 
.A(n_961),
.B(n_899),
.Y(n_1092)
);

AND2x4_ASAP7_75t_L g1093 ( 
.A(n_921),
.B(n_884),
.Y(n_1093)
);

NAND2xp5_ASAP7_75t_L g1094 ( 
.A(n_923),
.B(n_938),
.Y(n_1094)
);

AND2x2_ASAP7_75t_SL g1095 ( 
.A(n_841),
.B(n_1001),
.Y(n_1095)
);

OAI22xp5_ASAP7_75t_L g1096 ( 
.A1(n_841),
.A2(n_970),
.B1(n_930),
.B2(n_900),
.Y(n_1096)
);

NOR2xp33_ASAP7_75t_L g1097 ( 
.A(n_887),
.B(n_1023),
.Y(n_1097)
);

AOI21xp5_ASAP7_75t_L g1098 ( 
.A1(n_959),
.A2(n_977),
.B(n_1002),
.Y(n_1098)
);

INVxp67_ASAP7_75t_L g1099 ( 
.A(n_950),
.Y(n_1099)
);

O2A1O1Ixp5_ASAP7_75t_L g1100 ( 
.A1(n_924),
.A2(n_894),
.B(n_947),
.C(n_872),
.Y(n_1100)
);

NAND2xp5_ASAP7_75t_L g1101 ( 
.A(n_952),
.B(n_998),
.Y(n_1101)
);

NOR2xp33_ASAP7_75t_L g1102 ( 
.A(n_887),
.B(n_957),
.Y(n_1102)
);

O2A1O1Ixp5_ASAP7_75t_L g1103 ( 
.A1(n_1020),
.A2(n_913),
.B(n_911),
.C(n_910),
.Y(n_1103)
);

AOI22xp5_ASAP7_75t_L g1104 ( 
.A1(n_897),
.A2(n_1001),
.B1(n_1019),
.B2(n_989),
.Y(n_1104)
);

INVx1_ASAP7_75t_L g1105 ( 
.A(n_1012),
.Y(n_1105)
);

INVx1_ASAP7_75t_L g1106 ( 
.A(n_1013),
.Y(n_1106)
);

BUFx4f_ASAP7_75t_L g1107 ( 
.A(n_1005),
.Y(n_1107)
);

NOR2xp33_ASAP7_75t_L g1108 ( 
.A(n_915),
.B(n_854),
.Y(n_1108)
);

INVx1_ASAP7_75t_L g1109 ( 
.A(n_939),
.Y(n_1109)
);

A2O1A1Ixp33_ASAP7_75t_L g1110 ( 
.A1(n_992),
.A2(n_954),
.B(n_871),
.C(n_895),
.Y(n_1110)
);

AOI21xp5_ASAP7_75t_L g1111 ( 
.A1(n_1004),
.A2(n_942),
.B(n_943),
.Y(n_1111)
);

NAND2xp5_ASAP7_75t_SL g1112 ( 
.A(n_897),
.B(n_958),
.Y(n_1112)
);

O2A1O1Ixp33_ASAP7_75t_L g1113 ( 
.A1(n_932),
.A2(n_956),
.B(n_882),
.C(n_911),
.Y(n_1113)
);

AOI21xp5_ASAP7_75t_L g1114 ( 
.A1(n_861),
.A2(n_879),
.B(n_863),
.Y(n_1114)
);

INVx8_ASAP7_75t_L g1115 ( 
.A(n_948),
.Y(n_1115)
);

AOI21xp5_ASAP7_75t_L g1116 ( 
.A1(n_913),
.A2(n_898),
.B(n_865),
.Y(n_1116)
);

NOR2xp33_ASAP7_75t_R g1117 ( 
.A(n_953),
.B(n_945),
.Y(n_1117)
);

NAND2xp5_ASAP7_75t_L g1118 ( 
.A(n_995),
.B(n_1006),
.Y(n_1118)
);

INVx1_ASAP7_75t_L g1119 ( 
.A(n_1018),
.Y(n_1119)
);

CKINVDCx5p33_ASAP7_75t_R g1120 ( 
.A(n_982),
.Y(n_1120)
);

OAI22xp5_ASAP7_75t_L g1121 ( 
.A1(n_935),
.A2(n_986),
.B1(n_948),
.B2(n_946),
.Y(n_1121)
);

O2A1O1Ixp33_ASAP7_75t_SL g1122 ( 
.A1(n_1021),
.A2(n_875),
.B(n_979),
.C(n_866),
.Y(n_1122)
);

A2O1A1Ixp33_ASAP7_75t_L g1123 ( 
.A1(n_1017),
.A2(n_888),
.B(n_906),
.C(n_944),
.Y(n_1123)
);

INVx3_ASAP7_75t_L g1124 ( 
.A(n_1005),
.Y(n_1124)
);

BUFx2_ASAP7_75t_L g1125 ( 
.A(n_878),
.Y(n_1125)
);

NAND2xp5_ASAP7_75t_L g1126 ( 
.A(n_1007),
.B(n_1016),
.Y(n_1126)
);

NOR3xp33_ASAP7_75t_SL g1127 ( 
.A(n_971),
.B(n_949),
.C(n_929),
.Y(n_1127)
);

AOI22xp5_ASAP7_75t_L g1128 ( 
.A1(n_944),
.A2(n_878),
.B1(n_1011),
.B2(n_941),
.Y(n_1128)
);

OAI22xp5_ASAP7_75t_L g1129 ( 
.A1(n_1015),
.A2(n_963),
.B1(n_919),
.B2(n_967),
.Y(n_1129)
);

AOI21xp5_ASAP7_75t_L g1130 ( 
.A1(n_933),
.A2(n_985),
.B(n_993),
.Y(n_1130)
);

AOI21xp5_ASAP7_75t_L g1131 ( 
.A1(n_933),
.A2(n_996),
.B(n_1025),
.Y(n_1131)
);

OAI22xp5_ASAP7_75t_L g1132 ( 
.A1(n_1027),
.A2(n_1025),
.B1(n_844),
.B2(n_843),
.Y(n_1132)
);

NAND2xp5_ASAP7_75t_SL g1133 ( 
.A(n_850),
.B(n_637),
.Y(n_1133)
);

NAND2xp5_ASAP7_75t_L g1134 ( 
.A(n_1027),
.B(n_1025),
.Y(n_1134)
);

AOI22xp33_ASAP7_75t_L g1135 ( 
.A1(n_846),
.A2(n_750),
.B1(n_848),
.B2(n_544),
.Y(n_1135)
);

INVx1_ASAP7_75t_L g1136 ( 
.A(n_901),
.Y(n_1136)
);

BUFx2_ASAP7_75t_L g1137 ( 
.A(n_849),
.Y(n_1137)
);

NAND2xp5_ASAP7_75t_SL g1138 ( 
.A(n_850),
.B(n_637),
.Y(n_1138)
);

NAND2xp5_ASAP7_75t_L g1139 ( 
.A(n_1027),
.B(n_1025),
.Y(n_1139)
);

INVx2_ASAP7_75t_L g1140 ( 
.A(n_851),
.Y(n_1140)
);

AOI22xp5_ASAP7_75t_L g1141 ( 
.A1(n_848),
.A2(n_543),
.B1(n_844),
.B2(n_803),
.Y(n_1141)
);

NAND2xp5_ASAP7_75t_L g1142 ( 
.A(n_1027),
.B(n_1025),
.Y(n_1142)
);

BUFx6f_ASAP7_75t_L g1143 ( 
.A(n_883),
.Y(n_1143)
);

AND2x2_ASAP7_75t_L g1144 ( 
.A(n_864),
.B(n_846),
.Y(n_1144)
);

NAND2xp5_ASAP7_75t_L g1145 ( 
.A(n_1027),
.B(n_1025),
.Y(n_1145)
);

AOI21xp5_ASAP7_75t_L g1146 ( 
.A1(n_1025),
.A2(n_1027),
.B(n_549),
.Y(n_1146)
);

NOR3xp33_ASAP7_75t_L g1147 ( 
.A(n_844),
.B(n_543),
.C(n_848),
.Y(n_1147)
);

OR2x2_ASAP7_75t_L g1148 ( 
.A(n_844),
.B(n_525),
.Y(n_1148)
);

NAND2xp5_ASAP7_75t_L g1149 ( 
.A(n_1027),
.B(n_1025),
.Y(n_1149)
);

BUFx8_ASAP7_75t_L g1150 ( 
.A(n_1014),
.Y(n_1150)
);

O2A1O1Ixp5_ASAP7_75t_L g1151 ( 
.A1(n_984),
.A2(n_543),
.B(n_964),
.C(n_999),
.Y(n_1151)
);

AOI21xp5_ASAP7_75t_L g1152 ( 
.A1(n_1025),
.A2(n_1027),
.B(n_549),
.Y(n_1152)
);

A2O1A1Ixp33_ASAP7_75t_L g1153 ( 
.A1(n_848),
.A2(n_1026),
.B(n_844),
.C(n_964),
.Y(n_1153)
);

NAND2xp5_ASAP7_75t_SL g1154 ( 
.A(n_850),
.B(n_637),
.Y(n_1154)
);

INVx2_ASAP7_75t_L g1155 ( 
.A(n_851),
.Y(n_1155)
);

NAND2xp5_ASAP7_75t_L g1156 ( 
.A(n_1027),
.B(n_1025),
.Y(n_1156)
);

NOR2xp33_ASAP7_75t_L g1157 ( 
.A(n_1027),
.B(n_543),
.Y(n_1157)
);

O2A1O1Ixp33_ASAP7_75t_L g1158 ( 
.A1(n_1027),
.A2(n_543),
.B(n_844),
.C(n_1026),
.Y(n_1158)
);

INVx2_ASAP7_75t_SL g1159 ( 
.A(n_847),
.Y(n_1159)
);

CKINVDCx5p33_ASAP7_75t_R g1160 ( 
.A(n_1014),
.Y(n_1160)
);

INVx3_ASAP7_75t_L g1161 ( 
.A(n_976),
.Y(n_1161)
);

BUFx3_ASAP7_75t_L g1162 ( 
.A(n_847),
.Y(n_1162)
);

OAI22xp5_ASAP7_75t_SL g1163 ( 
.A1(n_1014),
.A2(n_527),
.B1(n_844),
.B2(n_543),
.Y(n_1163)
);

O2A1O1Ixp33_ASAP7_75t_L g1164 ( 
.A1(n_1027),
.A2(n_543),
.B(n_844),
.C(n_1026),
.Y(n_1164)
);

AO32x1_ASAP7_75t_L g1165 ( 
.A1(n_978),
.A2(n_1019),
.A3(n_924),
.B1(n_872),
.B2(n_892),
.Y(n_1165)
);

CKINVDCx5p33_ASAP7_75t_R g1166 ( 
.A(n_1014),
.Y(n_1166)
);

NAND2xp5_ASAP7_75t_L g1167 ( 
.A(n_1027),
.B(n_1025),
.Y(n_1167)
);

NAND2xp5_ASAP7_75t_SL g1168 ( 
.A(n_850),
.B(n_637),
.Y(n_1168)
);

INVx2_ASAP7_75t_L g1169 ( 
.A(n_851),
.Y(n_1169)
);

AOI21xp5_ASAP7_75t_L g1170 ( 
.A1(n_1025),
.A2(n_1027),
.B(n_549),
.Y(n_1170)
);

NAND2xp5_ASAP7_75t_L g1171 ( 
.A(n_1027),
.B(n_1025),
.Y(n_1171)
);

INVx2_ASAP7_75t_L g1172 ( 
.A(n_851),
.Y(n_1172)
);

AOI21xp5_ASAP7_75t_L g1173 ( 
.A1(n_1025),
.A2(n_1027),
.B(n_549),
.Y(n_1173)
);

AOI21xp5_ASAP7_75t_L g1174 ( 
.A1(n_1025),
.A2(n_1027),
.B(n_549),
.Y(n_1174)
);

INVx2_ASAP7_75t_L g1175 ( 
.A(n_851),
.Y(n_1175)
);

AOI21xp5_ASAP7_75t_L g1176 ( 
.A1(n_1025),
.A2(n_1027),
.B(n_549),
.Y(n_1176)
);

BUFx8_ASAP7_75t_L g1177 ( 
.A(n_1014),
.Y(n_1177)
);

AOI21xp5_ASAP7_75t_L g1178 ( 
.A1(n_1025),
.A2(n_1027),
.B(n_549),
.Y(n_1178)
);

OAI21xp33_ASAP7_75t_SL g1179 ( 
.A1(n_964),
.A2(n_844),
.B(n_843),
.Y(n_1179)
);

INVx2_ASAP7_75t_L g1180 ( 
.A(n_851),
.Y(n_1180)
);

OAI21x1_ASAP7_75t_L g1181 ( 
.A1(n_1055),
.A2(n_1114),
.B(n_1111),
.Y(n_1181)
);

BUFx3_ASAP7_75t_L g1182 ( 
.A(n_1063),
.Y(n_1182)
);

AOI21xp5_ASAP7_75t_L g1183 ( 
.A1(n_1134),
.A2(n_1156),
.B(n_1149),
.Y(n_1183)
);

INVx3_ASAP7_75t_L g1184 ( 
.A(n_1070),
.Y(n_1184)
);

CKINVDCx5p33_ASAP7_75t_R g1185 ( 
.A(n_1150),
.Y(n_1185)
);

NAND2xp5_ASAP7_75t_L g1186 ( 
.A(n_1139),
.B(n_1142),
.Y(n_1186)
);

INVx1_ASAP7_75t_L g1187 ( 
.A(n_1034),
.Y(n_1187)
);

BUFx2_ASAP7_75t_L g1188 ( 
.A(n_1137),
.Y(n_1188)
);

BUFx2_ASAP7_75t_L g1189 ( 
.A(n_1041),
.Y(n_1189)
);

AOI221xp5_ASAP7_75t_L g1190 ( 
.A1(n_1157),
.A2(n_1132),
.B1(n_1031),
.B2(n_1147),
.C(n_1164),
.Y(n_1190)
);

NOR2xp33_ASAP7_75t_L g1191 ( 
.A(n_1167),
.B(n_1171),
.Y(n_1191)
);

INVx1_ASAP7_75t_L g1192 ( 
.A(n_1136),
.Y(n_1192)
);

NOR2xp33_ASAP7_75t_L g1193 ( 
.A(n_1139),
.B(n_1142),
.Y(n_1193)
);

AOI21xp5_ASAP7_75t_L g1194 ( 
.A1(n_1145),
.A2(n_1132),
.B(n_1031),
.Y(n_1194)
);

AOI21xp5_ASAP7_75t_L g1195 ( 
.A1(n_1145),
.A2(n_1141),
.B(n_1153),
.Y(n_1195)
);

NAND2xp5_ASAP7_75t_L g1196 ( 
.A(n_1032),
.B(n_1158),
.Y(n_1196)
);

OAI22xp5_ASAP7_75t_L g1197 ( 
.A1(n_1036),
.A2(n_1049),
.B1(n_1037),
.B2(n_1095),
.Y(n_1197)
);

NAND2xp5_ASAP7_75t_SL g1198 ( 
.A(n_1045),
.B(n_1179),
.Y(n_1198)
);

AO31x2_ASAP7_75t_L g1199 ( 
.A1(n_1125),
.A2(n_1037),
.A3(n_1074),
.B(n_1121),
.Y(n_1199)
);

AOI21xp5_ASAP7_75t_L g1200 ( 
.A1(n_1146),
.A2(n_1170),
.B(n_1152),
.Y(n_1200)
);

NAND2xp5_ASAP7_75t_L g1201 ( 
.A(n_1073),
.B(n_1086),
.Y(n_1201)
);

NOR2xp33_ASAP7_75t_SL g1202 ( 
.A(n_1163),
.B(n_1075),
.Y(n_1202)
);

AND2x4_ASAP7_75t_L g1203 ( 
.A(n_1050),
.B(n_1062),
.Y(n_1203)
);

O2A1O1Ixp33_ASAP7_75t_SL g1204 ( 
.A1(n_1058),
.A2(n_1112),
.B(n_1089),
.C(n_1090),
.Y(n_1204)
);

INVx3_ASAP7_75t_SL g1205 ( 
.A(n_1160),
.Y(n_1205)
);

AOI21xp5_ASAP7_75t_L g1206 ( 
.A1(n_1173),
.A2(n_1174),
.B(n_1178),
.Y(n_1206)
);

OAI21xp5_ASAP7_75t_L g1207 ( 
.A1(n_1151),
.A2(n_1176),
.B(n_1104),
.Y(n_1207)
);

OAI21x1_ASAP7_75t_L g1208 ( 
.A1(n_1116),
.A2(n_1098),
.B(n_1067),
.Y(n_1208)
);

CKINVDCx16_ASAP7_75t_R g1209 ( 
.A(n_1030),
.Y(n_1209)
);

AOI21xp5_ASAP7_75t_L g1210 ( 
.A1(n_1131),
.A2(n_1065),
.B(n_1122),
.Y(n_1210)
);

NAND2xp5_ASAP7_75t_SL g1211 ( 
.A(n_1148),
.B(n_1042),
.Y(n_1211)
);

AOI21xp5_ASAP7_75t_L g1212 ( 
.A1(n_1130),
.A2(n_1060),
.B(n_1121),
.Y(n_1212)
);

BUFx6f_ASAP7_75t_L g1213 ( 
.A(n_1081),
.Y(n_1213)
);

A2O1A1Ixp33_ASAP7_75t_L g1214 ( 
.A1(n_1077),
.A2(n_1102),
.B(n_1064),
.C(n_1135),
.Y(n_1214)
);

O2A1O1Ixp33_ASAP7_75t_L g1215 ( 
.A1(n_1048),
.A2(n_1110),
.B(n_1040),
.C(n_1168),
.Y(n_1215)
);

AOI21xp5_ASAP7_75t_L g1216 ( 
.A1(n_1060),
.A2(n_1120),
.B(n_1123),
.Y(n_1216)
);

NOR2xp33_ASAP7_75t_L g1217 ( 
.A(n_1039),
.B(n_1144),
.Y(n_1217)
);

NAND2x1p5_ASAP7_75t_L g1218 ( 
.A(n_1107),
.B(n_1050),
.Y(n_1218)
);

BUFx3_ASAP7_75t_L g1219 ( 
.A(n_1053),
.Y(n_1219)
);

A2O1A1Ixp33_ASAP7_75t_L g1220 ( 
.A1(n_1082),
.A2(n_1040),
.B(n_1080),
.C(n_1097),
.Y(n_1220)
);

HB1xp67_ASAP7_75t_L g1221 ( 
.A(n_1052),
.Y(n_1221)
);

O2A1O1Ixp33_ASAP7_75t_SL g1222 ( 
.A1(n_1092),
.A2(n_1076),
.B(n_1054),
.C(n_1161),
.Y(n_1222)
);

AND2x4_ASAP7_75t_L g1223 ( 
.A(n_1062),
.B(n_1046),
.Y(n_1223)
);

OAI21x1_ASAP7_75t_L g1224 ( 
.A1(n_1103),
.A2(n_1126),
.B(n_1129),
.Y(n_1224)
);

BUFx3_ASAP7_75t_L g1225 ( 
.A(n_1057),
.Y(n_1225)
);

BUFx3_ASAP7_75t_L g1226 ( 
.A(n_1029),
.Y(n_1226)
);

INVx2_ASAP7_75t_L g1227 ( 
.A(n_1061),
.Y(n_1227)
);

AO21x2_ASAP7_75t_L g1228 ( 
.A1(n_1128),
.A2(n_1091),
.B(n_1117),
.Y(n_1228)
);

NAND2xp5_ASAP7_75t_L g1229 ( 
.A(n_1051),
.B(n_1119),
.Y(n_1229)
);

AOI21xp5_ASAP7_75t_L g1230 ( 
.A1(n_1165),
.A2(n_1113),
.B(n_1129),
.Y(n_1230)
);

BUFx10_ASAP7_75t_L g1231 ( 
.A(n_1166),
.Y(n_1231)
);

NAND2xp33_ASAP7_75t_L g1232 ( 
.A(n_1088),
.B(n_1161),
.Y(n_1232)
);

O2A1O1Ixp33_ASAP7_75t_SL g1233 ( 
.A1(n_1087),
.A2(n_1043),
.B(n_1044),
.C(n_1071),
.Y(n_1233)
);

NOR3xp33_ASAP7_75t_L g1234 ( 
.A(n_1133),
.B(n_1154),
.C(n_1138),
.Y(n_1234)
);

NAND2xp5_ASAP7_75t_L g1235 ( 
.A(n_1093),
.B(n_1118),
.Y(n_1235)
);

O2A1O1Ixp33_ASAP7_75t_L g1236 ( 
.A1(n_1100),
.A2(n_1046),
.B(n_1033),
.C(n_1085),
.Y(n_1236)
);

AO31x2_ASAP7_75t_L g1237 ( 
.A1(n_1096),
.A2(n_1108),
.A3(n_1118),
.B(n_1101),
.Y(n_1237)
);

AO31x2_ASAP7_75t_L g1238 ( 
.A1(n_1096),
.A2(n_1101),
.A3(n_1094),
.B(n_1105),
.Y(n_1238)
);

BUFx8_ASAP7_75t_SL g1239 ( 
.A(n_1162),
.Y(n_1239)
);

INVx3_ASAP7_75t_L g1240 ( 
.A(n_1115),
.Y(n_1240)
);

INVx1_ASAP7_75t_L g1241 ( 
.A(n_1106),
.Y(n_1241)
);

AOI21xp5_ASAP7_75t_L g1242 ( 
.A1(n_1165),
.A2(n_1093),
.B(n_1079),
.Y(n_1242)
);

AOI21xp5_ASAP7_75t_L g1243 ( 
.A1(n_1165),
.A2(n_1083),
.B(n_1081),
.Y(n_1243)
);

AOI21xp5_ASAP7_75t_L g1244 ( 
.A1(n_1083),
.A2(n_1081),
.B(n_1094),
.Y(n_1244)
);

NAND2xp33_ASAP7_75t_L g1245 ( 
.A(n_1081),
.B(n_1035),
.Y(n_1245)
);

A2O1A1Ixp33_ASAP7_75t_L g1246 ( 
.A1(n_1107),
.A2(n_1072),
.B(n_1099),
.C(n_1056),
.Y(n_1246)
);

O2A1O1Ixp33_ASAP7_75t_SL g1247 ( 
.A1(n_1124),
.A2(n_1159),
.B(n_1109),
.C(n_1172),
.Y(n_1247)
);

OAI21xp5_ASAP7_75t_L g1248 ( 
.A1(n_1127),
.A2(n_1072),
.B(n_1038),
.Y(n_1248)
);

INVx1_ASAP7_75t_L g1249 ( 
.A(n_1069),
.Y(n_1249)
);

INVx2_ASAP7_75t_L g1250 ( 
.A(n_1140),
.Y(n_1250)
);

INVx1_ASAP7_75t_SL g1251 ( 
.A(n_1078),
.Y(n_1251)
);

AND2x4_ASAP7_75t_L g1252 ( 
.A(n_1046),
.B(n_1047),
.Y(n_1252)
);

AOI21xp5_ASAP7_75t_L g1253 ( 
.A1(n_1115),
.A2(n_1035),
.B(n_1059),
.Y(n_1253)
);

AOI21xp5_ASAP7_75t_L g1254 ( 
.A1(n_1115),
.A2(n_1035),
.B(n_1059),
.Y(n_1254)
);

BUFx12f_ASAP7_75t_L g1255 ( 
.A(n_1150),
.Y(n_1255)
);

OAI21xp5_ASAP7_75t_L g1256 ( 
.A1(n_1155),
.A2(n_1180),
.B(n_1169),
.Y(n_1256)
);

INVx1_ASAP7_75t_L g1257 ( 
.A(n_1175),
.Y(n_1257)
);

AO31x2_ASAP7_75t_L g1258 ( 
.A1(n_1066),
.A2(n_1047),
.A3(n_1068),
.B(n_1059),
.Y(n_1258)
);

CKINVDCx20_ASAP7_75t_R g1259 ( 
.A(n_1177),
.Y(n_1259)
);

AOI21xp5_ASAP7_75t_L g1260 ( 
.A1(n_1084),
.A2(n_1143),
.B(n_1028),
.Y(n_1260)
);

AOI22xp5_ASAP7_75t_L g1261 ( 
.A1(n_1028),
.A2(n_1177),
.B1(n_1084),
.B2(n_1143),
.Y(n_1261)
);

AO21x1_ASAP7_75t_L g1262 ( 
.A1(n_1037),
.A2(n_1141),
.B(n_1147),
.Y(n_1262)
);

O2A1O1Ixp5_ASAP7_75t_L g1263 ( 
.A1(n_1151),
.A2(n_1037),
.B(n_999),
.C(n_1153),
.Y(n_1263)
);

OAI21x1_ASAP7_75t_L g1264 ( 
.A1(n_1055),
.A2(n_1114),
.B(n_1111),
.Y(n_1264)
);

AOI21xp5_ASAP7_75t_L g1265 ( 
.A1(n_1134),
.A2(n_1156),
.B(n_1149),
.Y(n_1265)
);

OAI21xp5_ASAP7_75t_L g1266 ( 
.A1(n_1141),
.A2(n_1179),
.B(n_1153),
.Y(n_1266)
);

CKINVDCx20_ASAP7_75t_R g1267 ( 
.A(n_1150),
.Y(n_1267)
);

AOI21xp5_ASAP7_75t_L g1268 ( 
.A1(n_1139),
.A2(n_1145),
.B(n_1142),
.Y(n_1268)
);

AOI21xp5_ASAP7_75t_L g1269 ( 
.A1(n_1134),
.A2(n_1156),
.B(n_1149),
.Y(n_1269)
);

AO21x2_ASAP7_75t_L g1270 ( 
.A1(n_1128),
.A2(n_1060),
.B(n_1091),
.Y(n_1270)
);

AOI21xp5_ASAP7_75t_L g1271 ( 
.A1(n_1134),
.A2(n_1156),
.B(n_1149),
.Y(n_1271)
);

OAI21x1_ASAP7_75t_L g1272 ( 
.A1(n_1055),
.A2(n_1114),
.B(n_1111),
.Y(n_1272)
);

NAND2xp5_ASAP7_75t_L g1273 ( 
.A(n_1139),
.B(n_1142),
.Y(n_1273)
);

BUFx6f_ASAP7_75t_L g1274 ( 
.A(n_1070),
.Y(n_1274)
);

INVx2_ASAP7_75t_L g1275 ( 
.A(n_1061),
.Y(n_1275)
);

NAND2xp5_ASAP7_75t_L g1276 ( 
.A(n_1139),
.B(n_1142),
.Y(n_1276)
);

NAND2xp5_ASAP7_75t_L g1277 ( 
.A(n_1139),
.B(n_1142),
.Y(n_1277)
);

AOI21xp5_ASAP7_75t_L g1278 ( 
.A1(n_1134),
.A2(n_1156),
.B(n_1149),
.Y(n_1278)
);

INVx2_ASAP7_75t_SL g1279 ( 
.A(n_1041),
.Y(n_1279)
);

BUFx2_ASAP7_75t_L g1280 ( 
.A(n_1063),
.Y(n_1280)
);

OAI21x1_ASAP7_75t_L g1281 ( 
.A1(n_1055),
.A2(n_1114),
.B(n_1111),
.Y(n_1281)
);

BUFx12f_ASAP7_75t_L g1282 ( 
.A(n_1150),
.Y(n_1282)
);

AOI21xp5_ASAP7_75t_L g1283 ( 
.A1(n_1134),
.A2(n_1156),
.B(n_1149),
.Y(n_1283)
);

AOI21xp5_ASAP7_75t_L g1284 ( 
.A1(n_1134),
.A2(n_1156),
.B(n_1149),
.Y(n_1284)
);

NAND2xp5_ASAP7_75t_L g1285 ( 
.A(n_1139),
.B(n_1142),
.Y(n_1285)
);

CKINVDCx11_ASAP7_75t_R g1286 ( 
.A(n_1053),
.Y(n_1286)
);

AO21x1_ASAP7_75t_L g1287 ( 
.A1(n_1037),
.A2(n_1141),
.B(n_1147),
.Y(n_1287)
);

OAI21x1_ASAP7_75t_L g1288 ( 
.A1(n_1055),
.A2(n_1114),
.B(n_1111),
.Y(n_1288)
);

NOR2xp33_ASAP7_75t_L g1289 ( 
.A(n_1157),
.B(n_543),
.Y(n_1289)
);

A2O1A1Ixp33_ASAP7_75t_L g1290 ( 
.A1(n_1141),
.A2(n_848),
.B(n_1179),
.C(n_1026),
.Y(n_1290)
);

AOI21xp5_ASAP7_75t_L g1291 ( 
.A1(n_1134),
.A2(n_1156),
.B(n_1149),
.Y(n_1291)
);

OAI22x1_ASAP7_75t_L g1292 ( 
.A1(n_1049),
.A2(n_1036),
.B1(n_526),
.B2(n_522),
.Y(n_1292)
);

INVx3_ASAP7_75t_L g1293 ( 
.A(n_1070),
.Y(n_1293)
);

BUFx3_ASAP7_75t_L g1294 ( 
.A(n_1063),
.Y(n_1294)
);

AOI21xp5_ASAP7_75t_L g1295 ( 
.A1(n_1134),
.A2(n_1156),
.B(n_1149),
.Y(n_1295)
);

AOI21xp5_ASAP7_75t_L g1296 ( 
.A1(n_1134),
.A2(n_1156),
.B(n_1149),
.Y(n_1296)
);

BUFx10_ASAP7_75t_L g1297 ( 
.A(n_1160),
.Y(n_1297)
);

NAND3xp33_ASAP7_75t_L g1298 ( 
.A(n_1141),
.B(n_543),
.C(n_1147),
.Y(n_1298)
);

OAI21xp5_ASAP7_75t_L g1299 ( 
.A1(n_1141),
.A2(n_1179),
.B(n_1153),
.Y(n_1299)
);

AO32x2_ASAP7_75t_L g1300 ( 
.A1(n_1037),
.A2(n_1031),
.A3(n_1132),
.B1(n_1096),
.B2(n_1121),
.Y(n_1300)
);

AOI21xp5_ASAP7_75t_L g1301 ( 
.A1(n_1134),
.A2(n_1156),
.B(n_1149),
.Y(n_1301)
);

INVx1_ASAP7_75t_L g1302 ( 
.A(n_1034),
.Y(n_1302)
);

INVx8_ASAP7_75t_L g1303 ( 
.A(n_1053),
.Y(n_1303)
);

OAI21x1_ASAP7_75t_L g1304 ( 
.A1(n_1055),
.A2(n_1114),
.B(n_1111),
.Y(n_1304)
);

INVx2_ASAP7_75t_L g1305 ( 
.A(n_1061),
.Y(n_1305)
);

OAI21x1_ASAP7_75t_L g1306 ( 
.A1(n_1055),
.A2(n_1114),
.B(n_1111),
.Y(n_1306)
);

INVx1_ASAP7_75t_L g1307 ( 
.A(n_1034),
.Y(n_1307)
);

NAND3xp33_ASAP7_75t_L g1308 ( 
.A(n_1141),
.B(n_543),
.C(n_1147),
.Y(n_1308)
);

O2A1O1Ixp33_ASAP7_75t_SL g1309 ( 
.A1(n_1153),
.A2(n_1134),
.B(n_1156),
.C(n_1149),
.Y(n_1309)
);

INVx2_ASAP7_75t_L g1310 ( 
.A(n_1061),
.Y(n_1310)
);

INVx5_ASAP7_75t_L g1311 ( 
.A(n_1115),
.Y(n_1311)
);

AOI21xp5_ASAP7_75t_L g1312 ( 
.A1(n_1134),
.A2(n_1156),
.B(n_1149),
.Y(n_1312)
);

OAI21x1_ASAP7_75t_L g1313 ( 
.A1(n_1055),
.A2(n_1114),
.B(n_1111),
.Y(n_1313)
);

NAND2xp5_ASAP7_75t_L g1314 ( 
.A(n_1139),
.B(n_1142),
.Y(n_1314)
);

NOR2xp33_ASAP7_75t_L g1315 ( 
.A(n_1157),
.B(n_543),
.Y(n_1315)
);

OAI21x1_ASAP7_75t_L g1316 ( 
.A1(n_1055),
.A2(n_1114),
.B(n_1111),
.Y(n_1316)
);

INVx3_ASAP7_75t_L g1317 ( 
.A(n_1070),
.Y(n_1317)
);

INVx2_ASAP7_75t_L g1318 ( 
.A(n_1061),
.Y(n_1318)
);

AOI21xp5_ASAP7_75t_L g1319 ( 
.A1(n_1139),
.A2(n_1145),
.B(n_1142),
.Y(n_1319)
);

INVx3_ASAP7_75t_L g1320 ( 
.A(n_1070),
.Y(n_1320)
);

INVx1_ASAP7_75t_L g1321 ( 
.A(n_1034),
.Y(n_1321)
);

AOI21xp5_ASAP7_75t_L g1322 ( 
.A1(n_1139),
.A2(n_1145),
.B(n_1142),
.Y(n_1322)
);

AOI21xp5_ASAP7_75t_L g1323 ( 
.A1(n_1139),
.A2(n_1145),
.B(n_1142),
.Y(n_1323)
);

AOI21x1_ASAP7_75t_L g1324 ( 
.A1(n_1037),
.A2(n_1131),
.B(n_1055),
.Y(n_1324)
);

AO31x2_ASAP7_75t_L g1325 ( 
.A1(n_1125),
.A2(n_910),
.A3(n_1037),
.B(n_894),
.Y(n_1325)
);

NAND2xp5_ASAP7_75t_L g1326 ( 
.A(n_1139),
.B(n_1142),
.Y(n_1326)
);

NAND2xp5_ASAP7_75t_L g1327 ( 
.A(n_1139),
.B(n_1142),
.Y(n_1327)
);

INVx1_ASAP7_75t_SL g1328 ( 
.A(n_1063),
.Y(n_1328)
);

HB1xp67_ASAP7_75t_L g1329 ( 
.A(n_1063),
.Y(n_1329)
);

A2O1A1Ixp33_ASAP7_75t_L g1330 ( 
.A1(n_1141),
.A2(n_848),
.B(n_1179),
.C(n_1026),
.Y(n_1330)
);

INVx1_ASAP7_75t_L g1331 ( 
.A(n_1034),
.Y(n_1331)
);

INVx2_ASAP7_75t_L g1332 ( 
.A(n_1061),
.Y(n_1332)
);

INVx4_ASAP7_75t_L g1333 ( 
.A(n_1274),
.Y(n_1333)
);

AOI22xp33_ASAP7_75t_SL g1334 ( 
.A1(n_1197),
.A2(n_1202),
.B1(n_1315),
.B2(n_1289),
.Y(n_1334)
);

BUFx4f_ASAP7_75t_L g1335 ( 
.A(n_1282),
.Y(n_1335)
);

INVx4_ASAP7_75t_L g1336 ( 
.A(n_1274),
.Y(n_1336)
);

AOI22xp33_ASAP7_75t_L g1337 ( 
.A1(n_1292),
.A2(n_1197),
.B1(n_1190),
.B2(n_1202),
.Y(n_1337)
);

AOI22xp33_ASAP7_75t_L g1338 ( 
.A1(n_1190),
.A2(n_1193),
.B1(n_1299),
.B2(n_1266),
.Y(n_1338)
);

CKINVDCx11_ASAP7_75t_R g1339 ( 
.A(n_1259),
.Y(n_1339)
);

AOI22xp5_ASAP7_75t_SL g1340 ( 
.A1(n_1267),
.A2(n_1209),
.B1(n_1201),
.B2(n_1217),
.Y(n_1340)
);

BUFx4f_ASAP7_75t_SL g1341 ( 
.A(n_1205),
.Y(n_1341)
);

CKINVDCx5p33_ASAP7_75t_R g1342 ( 
.A(n_1286),
.Y(n_1342)
);

INVx1_ASAP7_75t_L g1343 ( 
.A(n_1187),
.Y(n_1343)
);

INVx1_ASAP7_75t_L g1344 ( 
.A(n_1192),
.Y(n_1344)
);

CKINVDCx11_ASAP7_75t_R g1345 ( 
.A(n_1231),
.Y(n_1345)
);

CKINVDCx5p33_ASAP7_75t_R g1346 ( 
.A(n_1185),
.Y(n_1346)
);

CKINVDCx11_ASAP7_75t_R g1347 ( 
.A(n_1231),
.Y(n_1347)
);

INVx6_ASAP7_75t_L g1348 ( 
.A(n_1297),
.Y(n_1348)
);

OAI22xp33_ASAP7_75t_L g1349 ( 
.A1(n_1266),
.A2(n_1299),
.B1(n_1201),
.B2(n_1298),
.Y(n_1349)
);

AOI22xp33_ASAP7_75t_SL g1350 ( 
.A1(n_1191),
.A2(n_1308),
.B1(n_1195),
.B2(n_1196),
.Y(n_1350)
);

BUFx3_ASAP7_75t_L g1351 ( 
.A(n_1226),
.Y(n_1351)
);

AOI22xp33_ASAP7_75t_SL g1352 ( 
.A1(n_1196),
.A2(n_1194),
.B1(n_1285),
.B2(n_1277),
.Y(n_1352)
);

NAND2xp5_ASAP7_75t_L g1353 ( 
.A(n_1268),
.B(n_1319),
.Y(n_1353)
);

INVx3_ASAP7_75t_SL g1354 ( 
.A(n_1303),
.Y(n_1354)
);

INVxp67_ASAP7_75t_L g1355 ( 
.A(n_1188),
.Y(n_1355)
);

NAND2xp5_ASAP7_75t_L g1356 ( 
.A(n_1268),
.B(n_1319),
.Y(n_1356)
);

AOI22xp33_ASAP7_75t_SL g1357 ( 
.A1(n_1194),
.A2(n_1314),
.B1(n_1285),
.B2(n_1277),
.Y(n_1357)
);

INVx2_ASAP7_75t_SL g1358 ( 
.A(n_1303),
.Y(n_1358)
);

AOI22xp5_ASAP7_75t_L g1359 ( 
.A1(n_1234),
.A2(n_1198),
.B1(n_1262),
.B2(n_1287),
.Y(n_1359)
);

AOI22xp33_ASAP7_75t_L g1360 ( 
.A1(n_1250),
.A2(n_1332),
.B1(n_1318),
.B2(n_1310),
.Y(n_1360)
);

INVx2_ASAP7_75t_L g1361 ( 
.A(n_1275),
.Y(n_1361)
);

CKINVDCx11_ASAP7_75t_R g1362 ( 
.A(n_1219),
.Y(n_1362)
);

CKINVDCx9p33_ASAP7_75t_R g1363 ( 
.A(n_1189),
.Y(n_1363)
);

CKINVDCx20_ASAP7_75t_R g1364 ( 
.A(n_1239),
.Y(n_1364)
);

BUFx8_ASAP7_75t_L g1365 ( 
.A(n_1280),
.Y(n_1365)
);

OAI22xp5_ASAP7_75t_L g1366 ( 
.A1(n_1186),
.A2(n_1326),
.B1(n_1273),
.B2(n_1327),
.Y(n_1366)
);

INVx1_ASAP7_75t_SL g1367 ( 
.A(n_1328),
.Y(n_1367)
);

OAI21xp33_ASAP7_75t_L g1368 ( 
.A1(n_1290),
.A2(n_1330),
.B(n_1295),
.Y(n_1368)
);

AOI22xp33_ASAP7_75t_L g1369 ( 
.A1(n_1305),
.A2(n_1235),
.B1(n_1248),
.B2(n_1257),
.Y(n_1369)
);

INVx11_ASAP7_75t_L g1370 ( 
.A(n_1225),
.Y(n_1370)
);

NAND2xp5_ASAP7_75t_L g1371 ( 
.A(n_1322),
.B(n_1323),
.Y(n_1371)
);

OAI22xp5_ASAP7_75t_L g1372 ( 
.A1(n_1186),
.A2(n_1327),
.B1(n_1314),
.B2(n_1273),
.Y(n_1372)
);

AOI22xp33_ASAP7_75t_L g1373 ( 
.A1(n_1235),
.A2(n_1248),
.B1(n_1249),
.B2(n_1221),
.Y(n_1373)
);

OAI21xp33_ASAP7_75t_L g1374 ( 
.A1(n_1183),
.A2(n_1284),
.B(n_1278),
.Y(n_1374)
);

CKINVDCx11_ASAP7_75t_R g1375 ( 
.A(n_1328),
.Y(n_1375)
);

NAND2xp5_ASAP7_75t_L g1376 ( 
.A(n_1322),
.B(n_1323),
.Y(n_1376)
);

BUFx2_ASAP7_75t_SL g1377 ( 
.A(n_1279),
.Y(n_1377)
);

AOI22xp33_ASAP7_75t_L g1378 ( 
.A1(n_1229),
.A2(n_1228),
.B1(n_1326),
.B2(n_1276),
.Y(n_1378)
);

OAI22xp5_ASAP7_75t_L g1379 ( 
.A1(n_1276),
.A2(n_1271),
.B1(n_1283),
.B2(n_1269),
.Y(n_1379)
);

INVx6_ASAP7_75t_L g1380 ( 
.A(n_1311),
.Y(n_1380)
);

BUFx12f_ASAP7_75t_L g1381 ( 
.A(n_1213),
.Y(n_1381)
);

OAI21xp5_ASAP7_75t_L g1382 ( 
.A1(n_1263),
.A2(n_1214),
.B(n_1220),
.Y(n_1382)
);

OAI22xp5_ASAP7_75t_L g1383 ( 
.A1(n_1265),
.A2(n_1301),
.B1(n_1296),
.B2(n_1312),
.Y(n_1383)
);

BUFx8_ASAP7_75t_SL g1384 ( 
.A(n_1294),
.Y(n_1384)
);

BUFx12f_ASAP7_75t_L g1385 ( 
.A(n_1218),
.Y(n_1385)
);

CKINVDCx5p33_ASAP7_75t_R g1386 ( 
.A(n_1329),
.Y(n_1386)
);

OAI22xp5_ASAP7_75t_L g1387 ( 
.A1(n_1291),
.A2(n_1211),
.B1(n_1216),
.B2(n_1207),
.Y(n_1387)
);

NAND2xp5_ASAP7_75t_L g1388 ( 
.A(n_1309),
.B(n_1229),
.Y(n_1388)
);

BUFx12f_ASAP7_75t_L g1389 ( 
.A(n_1218),
.Y(n_1389)
);

INVx6_ASAP7_75t_L g1390 ( 
.A(n_1311),
.Y(n_1390)
);

INVx4_ASAP7_75t_L g1391 ( 
.A(n_1184),
.Y(n_1391)
);

OAI22xp33_ASAP7_75t_L g1392 ( 
.A1(n_1261),
.A2(n_1242),
.B1(n_1184),
.B2(n_1293),
.Y(n_1392)
);

INVx4_ASAP7_75t_L g1393 ( 
.A(n_1293),
.Y(n_1393)
);

CKINVDCx5p33_ASAP7_75t_R g1394 ( 
.A(n_1251),
.Y(n_1394)
);

OAI22xp5_ASAP7_75t_L g1395 ( 
.A1(n_1207),
.A2(n_1212),
.B1(n_1230),
.B2(n_1300),
.Y(n_1395)
);

AOI22xp33_ASAP7_75t_L g1396 ( 
.A1(n_1228),
.A2(n_1256),
.B1(n_1223),
.B2(n_1270),
.Y(n_1396)
);

OAI22xp5_ASAP7_75t_L g1397 ( 
.A1(n_1300),
.A2(n_1215),
.B1(n_1321),
.B2(n_1307),
.Y(n_1397)
);

BUFx10_ASAP7_75t_L g1398 ( 
.A(n_1252),
.Y(n_1398)
);

AND2x2_ASAP7_75t_L g1399 ( 
.A(n_1251),
.B(n_1317),
.Y(n_1399)
);

BUFx10_ASAP7_75t_L g1400 ( 
.A(n_1252),
.Y(n_1400)
);

BUFx6f_ASAP7_75t_SL g1401 ( 
.A(n_1203),
.Y(n_1401)
);

BUFx4f_ASAP7_75t_L g1402 ( 
.A(n_1317),
.Y(n_1402)
);

CKINVDCx11_ASAP7_75t_R g1403 ( 
.A(n_1223),
.Y(n_1403)
);

OR2x2_ASAP7_75t_L g1404 ( 
.A(n_1302),
.B(n_1331),
.Y(n_1404)
);

AOI22xp33_ASAP7_75t_SL g1405 ( 
.A1(n_1270),
.A2(n_1242),
.B1(n_1300),
.B2(n_1241),
.Y(n_1405)
);

BUFx6f_ASAP7_75t_L g1406 ( 
.A(n_1320),
.Y(n_1406)
);

INVx1_ASAP7_75t_L g1407 ( 
.A(n_1233),
.Y(n_1407)
);

OAI22xp33_ASAP7_75t_L g1408 ( 
.A1(n_1311),
.A2(n_1243),
.B1(n_1244),
.B2(n_1240),
.Y(n_1408)
);

INVx1_ASAP7_75t_L g1409 ( 
.A(n_1256),
.Y(n_1409)
);

BUFx3_ASAP7_75t_L g1410 ( 
.A(n_1258),
.Y(n_1410)
);

INVx6_ASAP7_75t_L g1411 ( 
.A(n_1203),
.Y(n_1411)
);

INVx4_ASAP7_75t_L g1412 ( 
.A(n_1240),
.Y(n_1412)
);

OAI21xp33_ASAP7_75t_L g1413 ( 
.A1(n_1324),
.A2(n_1236),
.B(n_1210),
.Y(n_1413)
);

INVx6_ASAP7_75t_L g1414 ( 
.A(n_1232),
.Y(n_1414)
);

BUFx8_ASAP7_75t_L g1415 ( 
.A(n_1260),
.Y(n_1415)
);

AOI22xp33_ASAP7_75t_L g1416 ( 
.A1(n_1245),
.A2(n_1253),
.B1(n_1254),
.B2(n_1224),
.Y(n_1416)
);

OAI22xp5_ASAP7_75t_L g1417 ( 
.A1(n_1246),
.A2(n_1206),
.B1(n_1200),
.B2(n_1199),
.Y(n_1417)
);

AOI22xp33_ASAP7_75t_L g1418 ( 
.A1(n_1200),
.A2(n_1206),
.B1(n_1247),
.B2(n_1199),
.Y(n_1418)
);

CKINVDCx5p33_ASAP7_75t_R g1419 ( 
.A(n_1204),
.Y(n_1419)
);

INVx3_ASAP7_75t_L g1420 ( 
.A(n_1238),
.Y(n_1420)
);

INVx6_ASAP7_75t_L g1421 ( 
.A(n_1222),
.Y(n_1421)
);

BUFx6f_ASAP7_75t_L g1422 ( 
.A(n_1208),
.Y(n_1422)
);

AOI22xp33_ASAP7_75t_L g1423 ( 
.A1(n_1199),
.A2(n_1237),
.B1(n_1181),
.B2(n_1264),
.Y(n_1423)
);

BUFx8_ASAP7_75t_L g1424 ( 
.A(n_1237),
.Y(n_1424)
);

BUFx12f_ASAP7_75t_L g1425 ( 
.A(n_1325),
.Y(n_1425)
);

OAI22xp33_ASAP7_75t_L g1426 ( 
.A1(n_1325),
.A2(n_1272),
.B1(n_1281),
.B2(n_1288),
.Y(n_1426)
);

AOI22xp33_ASAP7_75t_L g1427 ( 
.A1(n_1304),
.A2(n_1306),
.B1(n_1313),
.B2(n_1316),
.Y(n_1427)
);

INVx1_ASAP7_75t_L g1428 ( 
.A(n_1187),
.Y(n_1428)
);

AOI22xp33_ASAP7_75t_L g1429 ( 
.A1(n_1292),
.A2(n_750),
.B1(n_848),
.B2(n_1135),
.Y(n_1429)
);

AOI22xp5_ASAP7_75t_L g1430 ( 
.A1(n_1289),
.A2(n_1315),
.B1(n_543),
.B2(n_1157),
.Y(n_1430)
);

INVx3_ASAP7_75t_L g1431 ( 
.A(n_1213),
.Y(n_1431)
);

AOI22xp33_ASAP7_75t_L g1432 ( 
.A1(n_1292),
.A2(n_750),
.B1(n_848),
.B2(n_1135),
.Y(n_1432)
);

BUFx8_ASAP7_75t_L g1433 ( 
.A(n_1255),
.Y(n_1433)
);

AOI22xp5_ASAP7_75t_L g1434 ( 
.A1(n_1289),
.A2(n_1315),
.B1(n_543),
.B2(n_1157),
.Y(n_1434)
);

BUFx10_ASAP7_75t_L g1435 ( 
.A(n_1185),
.Y(n_1435)
);

AOI22xp33_ASAP7_75t_L g1436 ( 
.A1(n_1292),
.A2(n_750),
.B1(n_848),
.B2(n_1135),
.Y(n_1436)
);

INVx1_ASAP7_75t_L g1437 ( 
.A(n_1187),
.Y(n_1437)
);

CKINVDCx6p67_ASAP7_75t_R g1438 ( 
.A(n_1255),
.Y(n_1438)
);

AOI22xp33_ASAP7_75t_SL g1439 ( 
.A1(n_1197),
.A2(n_1095),
.B1(n_750),
.B2(n_1037),
.Y(n_1439)
);

NAND2xp5_ASAP7_75t_L g1440 ( 
.A(n_1193),
.B(n_1268),
.Y(n_1440)
);

CKINVDCx11_ASAP7_75t_R g1441 ( 
.A(n_1259),
.Y(n_1441)
);

AOI22xp33_ASAP7_75t_L g1442 ( 
.A1(n_1292),
.A2(n_750),
.B1(n_848),
.B2(n_1135),
.Y(n_1442)
);

HB1xp67_ASAP7_75t_L g1443 ( 
.A(n_1329),
.Y(n_1443)
);

INVx2_ASAP7_75t_L g1444 ( 
.A(n_1227),
.Y(n_1444)
);

BUFx2_ASAP7_75t_L g1445 ( 
.A(n_1182),
.Y(n_1445)
);

OAI21xp33_ASAP7_75t_L g1446 ( 
.A1(n_1289),
.A2(n_1315),
.B(n_543),
.Y(n_1446)
);

CKINVDCx20_ASAP7_75t_R g1447 ( 
.A(n_1259),
.Y(n_1447)
);

AOI22xp33_ASAP7_75t_L g1448 ( 
.A1(n_1292),
.A2(n_750),
.B1(n_848),
.B2(n_1135),
.Y(n_1448)
);

CKINVDCx20_ASAP7_75t_R g1449 ( 
.A(n_1259),
.Y(n_1449)
);

BUFx12f_ASAP7_75t_L g1450 ( 
.A(n_1286),
.Y(n_1450)
);

BUFx6f_ASAP7_75t_SL g1451 ( 
.A(n_1231),
.Y(n_1451)
);

CKINVDCx11_ASAP7_75t_R g1452 ( 
.A(n_1259),
.Y(n_1452)
);

OAI22xp33_ASAP7_75t_L g1453 ( 
.A1(n_1202),
.A2(n_1141),
.B1(n_844),
.B2(n_1036),
.Y(n_1453)
);

INVx1_ASAP7_75t_L g1454 ( 
.A(n_1440),
.Y(n_1454)
);

INVx1_ASAP7_75t_L g1455 ( 
.A(n_1440),
.Y(n_1455)
);

BUFx4f_ASAP7_75t_L g1456 ( 
.A(n_1414),
.Y(n_1456)
);

INVx2_ASAP7_75t_SL g1457 ( 
.A(n_1443),
.Y(n_1457)
);

INVx1_ASAP7_75t_L g1458 ( 
.A(n_1409),
.Y(n_1458)
);

INVx1_ASAP7_75t_L g1459 ( 
.A(n_1420),
.Y(n_1459)
);

INVx1_ASAP7_75t_L g1460 ( 
.A(n_1353),
.Y(n_1460)
);

AO21x2_ASAP7_75t_L g1461 ( 
.A1(n_1426),
.A2(n_1413),
.B(n_1374),
.Y(n_1461)
);

HB1xp67_ASAP7_75t_L g1462 ( 
.A(n_1367),
.Y(n_1462)
);

AND2x2_ASAP7_75t_L g1463 ( 
.A(n_1405),
.B(n_1343),
.Y(n_1463)
);

BUFx2_ASAP7_75t_L g1464 ( 
.A(n_1422),
.Y(n_1464)
);

AND2x2_ASAP7_75t_L g1465 ( 
.A(n_1405),
.B(n_1344),
.Y(n_1465)
);

AOI221xp5_ASAP7_75t_L g1466 ( 
.A1(n_1446),
.A2(n_1349),
.B1(n_1453),
.B2(n_1337),
.C(n_1338),
.Y(n_1466)
);

INVx1_ASAP7_75t_L g1467 ( 
.A(n_1353),
.Y(n_1467)
);

INVx1_ASAP7_75t_L g1468 ( 
.A(n_1356),
.Y(n_1468)
);

OR2x6_ASAP7_75t_L g1469 ( 
.A(n_1410),
.B(n_1425),
.Y(n_1469)
);

INVx2_ASAP7_75t_SL g1470 ( 
.A(n_1414),
.Y(n_1470)
);

INVx1_ASAP7_75t_L g1471 ( 
.A(n_1371),
.Y(n_1471)
);

INVx1_ASAP7_75t_L g1472 ( 
.A(n_1371),
.Y(n_1472)
);

OAI21x1_ASAP7_75t_L g1473 ( 
.A1(n_1383),
.A2(n_1427),
.B(n_1417),
.Y(n_1473)
);

BUFx8_ASAP7_75t_L g1474 ( 
.A(n_1451),
.Y(n_1474)
);

NOR2xp33_ASAP7_75t_L g1475 ( 
.A(n_1430),
.B(n_1434),
.Y(n_1475)
);

OAI21x1_ASAP7_75t_L g1476 ( 
.A1(n_1383),
.A2(n_1417),
.B(n_1418),
.Y(n_1476)
);

OAI21xp5_ASAP7_75t_L g1477 ( 
.A1(n_1334),
.A2(n_1350),
.B(n_1382),
.Y(n_1477)
);

HB1xp67_ASAP7_75t_L g1478 ( 
.A(n_1355),
.Y(n_1478)
);

OR2x2_ASAP7_75t_L g1479 ( 
.A(n_1395),
.B(n_1376),
.Y(n_1479)
);

AOI22xp33_ASAP7_75t_SL g1480 ( 
.A1(n_1424),
.A2(n_1382),
.B1(n_1421),
.B2(n_1340),
.Y(n_1480)
);

INVx1_ASAP7_75t_L g1481 ( 
.A(n_1428),
.Y(n_1481)
);

BUFx3_ASAP7_75t_L g1482 ( 
.A(n_1415),
.Y(n_1482)
);

BUFx2_ASAP7_75t_L g1483 ( 
.A(n_1424),
.Y(n_1483)
);

HB1xp67_ASAP7_75t_L g1484 ( 
.A(n_1404),
.Y(n_1484)
);

INVxp67_ASAP7_75t_SL g1485 ( 
.A(n_1388),
.Y(n_1485)
);

CKINVDCx20_ASAP7_75t_R g1486 ( 
.A(n_1447),
.Y(n_1486)
);

INVx1_ASAP7_75t_L g1487 ( 
.A(n_1437),
.Y(n_1487)
);

NAND2xp5_ASAP7_75t_L g1488 ( 
.A(n_1366),
.B(n_1372),
.Y(n_1488)
);

OR2x2_ASAP7_75t_L g1489 ( 
.A(n_1395),
.B(n_1366),
.Y(n_1489)
);

BUFx3_ASAP7_75t_L g1490 ( 
.A(n_1415),
.Y(n_1490)
);

INVx3_ASAP7_75t_L g1491 ( 
.A(n_1407),
.Y(n_1491)
);

INVx1_ASAP7_75t_L g1492 ( 
.A(n_1379),
.Y(n_1492)
);

AOI22xp33_ASAP7_75t_L g1493 ( 
.A1(n_1439),
.A2(n_1432),
.B1(n_1429),
.B2(n_1436),
.Y(n_1493)
);

INVx1_ASAP7_75t_L g1494 ( 
.A(n_1379),
.Y(n_1494)
);

INVx1_ASAP7_75t_L g1495 ( 
.A(n_1397),
.Y(n_1495)
);

OAI21x1_ASAP7_75t_L g1496 ( 
.A1(n_1423),
.A2(n_1387),
.B(n_1416),
.Y(n_1496)
);

INVx1_ASAP7_75t_L g1497 ( 
.A(n_1397),
.Y(n_1497)
);

INVx2_ASAP7_75t_SL g1498 ( 
.A(n_1414),
.Y(n_1498)
);

BUFx3_ASAP7_75t_L g1499 ( 
.A(n_1445),
.Y(n_1499)
);

INVx2_ASAP7_75t_SL g1500 ( 
.A(n_1411),
.Y(n_1500)
);

OAI21x1_ASAP7_75t_L g1501 ( 
.A1(n_1387),
.A2(n_1388),
.B(n_1368),
.Y(n_1501)
);

INVx2_ASAP7_75t_L g1502 ( 
.A(n_1361),
.Y(n_1502)
);

INVx2_ASAP7_75t_L g1503 ( 
.A(n_1444),
.Y(n_1503)
);

INVx1_ASAP7_75t_L g1504 ( 
.A(n_1372),
.Y(n_1504)
);

AND2x2_ASAP7_75t_L g1505 ( 
.A(n_1352),
.B(n_1357),
.Y(n_1505)
);

AND2x2_ASAP7_75t_L g1506 ( 
.A(n_1352),
.B(n_1357),
.Y(n_1506)
);

AOI22xp33_ASAP7_75t_L g1507 ( 
.A1(n_1439),
.A2(n_1448),
.B1(n_1442),
.B2(n_1334),
.Y(n_1507)
);

INVx1_ASAP7_75t_L g1508 ( 
.A(n_1378),
.Y(n_1508)
);

INVx1_ASAP7_75t_L g1509 ( 
.A(n_1359),
.Y(n_1509)
);

AND2x2_ASAP7_75t_L g1510 ( 
.A(n_1399),
.B(n_1396),
.Y(n_1510)
);

INVx1_ASAP7_75t_L g1511 ( 
.A(n_1408),
.Y(n_1511)
);

OAI21xp33_ASAP7_75t_SL g1512 ( 
.A1(n_1373),
.A2(n_1369),
.B(n_1419),
.Y(n_1512)
);

NAND2xp5_ASAP7_75t_L g1513 ( 
.A(n_1394),
.B(n_1386),
.Y(n_1513)
);

BUFx2_ASAP7_75t_L g1514 ( 
.A(n_1365),
.Y(n_1514)
);

INVx2_ASAP7_75t_SL g1515 ( 
.A(n_1411),
.Y(n_1515)
);

INVx1_ASAP7_75t_SL g1516 ( 
.A(n_1375),
.Y(n_1516)
);

OA21x2_ASAP7_75t_L g1517 ( 
.A1(n_1360),
.A2(n_1392),
.B(n_1380),
.Y(n_1517)
);

INVx3_ASAP7_75t_L g1518 ( 
.A(n_1412),
.Y(n_1518)
);

NOR2xp33_ASAP7_75t_L g1519 ( 
.A(n_1449),
.B(n_1393),
.Y(n_1519)
);

NAND2xp5_ASAP7_75t_L g1520 ( 
.A(n_1406),
.B(n_1393),
.Y(n_1520)
);

AOI21xp5_ASAP7_75t_L g1521 ( 
.A1(n_1412),
.A2(n_1402),
.B(n_1431),
.Y(n_1521)
);

AND2x2_ASAP7_75t_L g1522 ( 
.A(n_1391),
.B(n_1403),
.Y(n_1522)
);

INVx1_ASAP7_75t_L g1523 ( 
.A(n_1398),
.Y(n_1523)
);

INVx2_ASAP7_75t_L g1524 ( 
.A(n_1411),
.Y(n_1524)
);

INVx1_ASAP7_75t_L g1525 ( 
.A(n_1400),
.Y(n_1525)
);

AND2x2_ASAP7_75t_L g1526 ( 
.A(n_1391),
.B(n_1406),
.Y(n_1526)
);

INVx1_ASAP7_75t_L g1527 ( 
.A(n_1380),
.Y(n_1527)
);

OAI21x1_ASAP7_75t_L g1528 ( 
.A1(n_1390),
.A2(n_1401),
.B(n_1363),
.Y(n_1528)
);

BUFx3_ASAP7_75t_L g1529 ( 
.A(n_1381),
.Y(n_1529)
);

INVx1_ASAP7_75t_L g1530 ( 
.A(n_1333),
.Y(n_1530)
);

INVx1_ASAP7_75t_L g1531 ( 
.A(n_1336),
.Y(n_1531)
);

INVx1_ASAP7_75t_L g1532 ( 
.A(n_1377),
.Y(n_1532)
);

BUFx3_ASAP7_75t_L g1533 ( 
.A(n_1365),
.Y(n_1533)
);

INVx1_ASAP7_75t_L g1534 ( 
.A(n_1385),
.Y(n_1534)
);

INVx1_ASAP7_75t_L g1535 ( 
.A(n_1389),
.Y(n_1535)
);

OAI21x1_ASAP7_75t_L g1536 ( 
.A1(n_1402),
.A2(n_1451),
.B(n_1348),
.Y(n_1536)
);

O2A1O1Ixp33_ASAP7_75t_L g1537 ( 
.A1(n_1354),
.A2(n_1358),
.B(n_1351),
.C(n_1364),
.Y(n_1537)
);

OA21x2_ASAP7_75t_L g1538 ( 
.A1(n_1501),
.A2(n_1346),
.B(n_1342),
.Y(n_1538)
);

AO21x2_ASAP7_75t_L g1539 ( 
.A1(n_1508),
.A2(n_1384),
.B(n_1362),
.Y(n_1539)
);

NOR2xp33_ASAP7_75t_L g1540 ( 
.A(n_1475),
.B(n_1341),
.Y(n_1540)
);

OA21x2_ASAP7_75t_L g1541 ( 
.A1(n_1501),
.A2(n_1345),
.B(n_1347),
.Y(n_1541)
);

AND2x2_ASAP7_75t_L g1542 ( 
.A(n_1499),
.B(n_1335),
.Y(n_1542)
);

AO32x2_ASAP7_75t_L g1543 ( 
.A1(n_1457),
.A2(n_1470),
.A3(n_1498),
.B1(n_1515),
.B2(n_1500),
.Y(n_1543)
);

CKINVDCx5p33_ASAP7_75t_R g1544 ( 
.A(n_1486),
.Y(n_1544)
);

A2O1A1Ixp33_ASAP7_75t_L g1545 ( 
.A1(n_1477),
.A2(n_1450),
.B(n_1438),
.C(n_1433),
.Y(n_1545)
);

AOI21xp33_ASAP7_75t_L g1546 ( 
.A1(n_1512),
.A2(n_1433),
.B(n_1370),
.Y(n_1546)
);

OR2x2_ASAP7_75t_L g1547 ( 
.A(n_1484),
.B(n_1339),
.Y(n_1547)
);

NAND2xp5_ASAP7_75t_L g1548 ( 
.A(n_1454),
.B(n_1435),
.Y(n_1548)
);

HB1xp67_ASAP7_75t_SL g1549 ( 
.A(n_1474),
.Y(n_1549)
);

INVxp67_ASAP7_75t_L g1550 ( 
.A(n_1462),
.Y(n_1550)
);

O2A1O1Ixp33_ASAP7_75t_SL g1551 ( 
.A1(n_1466),
.A2(n_1441),
.B(n_1452),
.C(n_1488),
.Y(n_1551)
);

NAND2xp5_ASAP7_75t_L g1552 ( 
.A(n_1455),
.B(n_1504),
.Y(n_1552)
);

OAI21xp5_ASAP7_75t_L g1553 ( 
.A1(n_1505),
.A2(n_1506),
.B(n_1512),
.Y(n_1553)
);

AND2x4_ASAP7_75t_L g1554 ( 
.A(n_1528),
.B(n_1510),
.Y(n_1554)
);

OAI21xp5_ASAP7_75t_L g1555 ( 
.A1(n_1505),
.A2(n_1506),
.B(n_1507),
.Y(n_1555)
);

HB1xp67_ASAP7_75t_L g1556 ( 
.A(n_1478),
.Y(n_1556)
);

AOI221xp5_ASAP7_75t_L g1557 ( 
.A1(n_1495),
.A2(n_1497),
.B1(n_1489),
.B2(n_1509),
.C(n_1504),
.Y(n_1557)
);

OAI22xp5_ASAP7_75t_L g1558 ( 
.A1(n_1493),
.A2(n_1509),
.B1(n_1479),
.B2(n_1480),
.Y(n_1558)
);

OAI22xp5_ASAP7_75t_L g1559 ( 
.A1(n_1479),
.A2(n_1456),
.B1(n_1492),
.B2(n_1494),
.Y(n_1559)
);

OR2x6_ASAP7_75t_L g1560 ( 
.A(n_1469),
.B(n_1483),
.Y(n_1560)
);

AOI22xp33_ASAP7_75t_L g1561 ( 
.A1(n_1510),
.A2(n_1463),
.B1(n_1465),
.B2(n_1497),
.Y(n_1561)
);

NOR2xp33_ASAP7_75t_L g1562 ( 
.A(n_1516),
.B(n_1519),
.Y(n_1562)
);

A2O1A1Ixp33_ASAP7_75t_L g1563 ( 
.A1(n_1463),
.A2(n_1465),
.B(n_1511),
.C(n_1476),
.Y(n_1563)
);

AOI221xp5_ASAP7_75t_L g1564 ( 
.A1(n_1492),
.A2(n_1494),
.B1(n_1511),
.B2(n_1485),
.C(n_1481),
.Y(n_1564)
);

NAND2xp5_ASAP7_75t_L g1565 ( 
.A(n_1460),
.B(n_1467),
.Y(n_1565)
);

O2A1O1Ixp33_ASAP7_75t_SL g1566 ( 
.A1(n_1532),
.A2(n_1537),
.B(n_1513),
.C(n_1520),
.Y(n_1566)
);

AND2x4_ASAP7_75t_L g1567 ( 
.A(n_1482),
.B(n_1490),
.Y(n_1567)
);

AND2x4_ASAP7_75t_L g1568 ( 
.A(n_1482),
.B(n_1490),
.Y(n_1568)
);

NAND2x1_ASAP7_75t_L g1569 ( 
.A(n_1518),
.B(n_1491),
.Y(n_1569)
);

O2A1O1Ixp33_ASAP7_75t_SL g1570 ( 
.A1(n_1532),
.A2(n_1521),
.B(n_1531),
.C(n_1530),
.Y(n_1570)
);

AND2x2_ASAP7_75t_L g1571 ( 
.A(n_1522),
.B(n_1526),
.Y(n_1571)
);

NAND3xp33_ASAP7_75t_L g1572 ( 
.A(n_1460),
.B(n_1471),
.C(n_1472),
.Y(n_1572)
);

NOR2xp33_ASAP7_75t_L g1573 ( 
.A(n_1514),
.B(n_1533),
.Y(n_1573)
);

OAI21xp5_ASAP7_75t_L g1574 ( 
.A1(n_1476),
.A2(n_1496),
.B(n_1473),
.Y(n_1574)
);

AO32x2_ASAP7_75t_L g1575 ( 
.A1(n_1500),
.A2(n_1515),
.A3(n_1487),
.B1(n_1503),
.B2(n_1502),
.Y(n_1575)
);

AND2x6_ASAP7_75t_L g1576 ( 
.A(n_1524),
.B(n_1527),
.Y(n_1576)
);

INVx2_ASAP7_75t_L g1577 ( 
.A(n_1575),
.Y(n_1577)
);

HB1xp67_ASAP7_75t_L g1578 ( 
.A(n_1565),
.Y(n_1578)
);

BUFx2_ASAP7_75t_L g1579 ( 
.A(n_1543),
.Y(n_1579)
);

AOI22xp33_ASAP7_75t_SL g1580 ( 
.A1(n_1553),
.A2(n_1461),
.B1(n_1517),
.B2(n_1496),
.Y(n_1580)
);

AOI222xp33_ASAP7_75t_L g1581 ( 
.A1(n_1555),
.A2(n_1474),
.B1(n_1514),
.B2(n_1534),
.C1(n_1535),
.C2(n_1533),
.Y(n_1581)
);

INVx2_ASAP7_75t_L g1582 ( 
.A(n_1575),
.Y(n_1582)
);

AOI22xp33_ASAP7_75t_L g1583 ( 
.A1(n_1553),
.A2(n_1517),
.B1(n_1461),
.B2(n_1458),
.Y(n_1583)
);

INVx3_ASAP7_75t_L g1584 ( 
.A(n_1569),
.Y(n_1584)
);

BUFx2_ASAP7_75t_L g1585 ( 
.A(n_1543),
.Y(n_1585)
);

NOR2xp33_ASAP7_75t_L g1586 ( 
.A(n_1566),
.B(n_1531),
.Y(n_1586)
);

INVx2_ASAP7_75t_L g1587 ( 
.A(n_1575),
.Y(n_1587)
);

NAND2xp5_ASAP7_75t_L g1588 ( 
.A(n_1572),
.B(n_1557),
.Y(n_1588)
);

AND2x4_ASAP7_75t_L g1589 ( 
.A(n_1576),
.B(n_1459),
.Y(n_1589)
);

NAND2xp5_ASAP7_75t_L g1590 ( 
.A(n_1557),
.B(n_1468),
.Y(n_1590)
);

INVx1_ASAP7_75t_L g1591 ( 
.A(n_1552),
.Y(n_1591)
);

AND2x2_ASAP7_75t_L g1592 ( 
.A(n_1574),
.B(n_1473),
.Y(n_1592)
);

AND2x2_ASAP7_75t_L g1593 ( 
.A(n_1574),
.B(n_1491),
.Y(n_1593)
);

INVx3_ASAP7_75t_L g1594 ( 
.A(n_1538),
.Y(n_1594)
);

OR2x6_ASAP7_75t_SL g1595 ( 
.A(n_1559),
.B(n_1523),
.Y(n_1595)
);

AOI22xp5_ASAP7_75t_L g1596 ( 
.A1(n_1558),
.A2(n_1534),
.B1(n_1535),
.B2(n_1525),
.Y(n_1596)
);

AND2x2_ASAP7_75t_L g1597 ( 
.A(n_1543),
.B(n_1464),
.Y(n_1597)
);

AND2x2_ASAP7_75t_L g1598 ( 
.A(n_1579),
.B(n_1559),
.Y(n_1598)
);

AND2x2_ASAP7_75t_L g1599 ( 
.A(n_1579),
.B(n_1538),
.Y(n_1599)
);

BUFx3_ASAP7_75t_L g1600 ( 
.A(n_1595),
.Y(n_1600)
);

INVx1_ASAP7_75t_L g1601 ( 
.A(n_1578),
.Y(n_1601)
);

INVx2_ASAP7_75t_L g1602 ( 
.A(n_1577),
.Y(n_1602)
);

AND2x2_ASAP7_75t_L g1603 ( 
.A(n_1579),
.B(n_1541),
.Y(n_1603)
);

AND2x2_ASAP7_75t_L g1604 ( 
.A(n_1585),
.B(n_1541),
.Y(n_1604)
);

NAND2xp5_ASAP7_75t_L g1605 ( 
.A(n_1588),
.B(n_1564),
.Y(n_1605)
);

BUFx3_ASAP7_75t_L g1606 ( 
.A(n_1595),
.Y(n_1606)
);

INVx4_ASAP7_75t_L g1607 ( 
.A(n_1584),
.Y(n_1607)
);

AOI221xp5_ASAP7_75t_L g1608 ( 
.A1(n_1588),
.A2(n_1558),
.B1(n_1551),
.B2(n_1546),
.C(n_1563),
.Y(n_1608)
);

NAND2xp5_ASAP7_75t_L g1609 ( 
.A(n_1590),
.B(n_1550),
.Y(n_1609)
);

AND2x2_ASAP7_75t_L g1610 ( 
.A(n_1585),
.B(n_1571),
.Y(n_1610)
);

AOI22xp33_ASAP7_75t_L g1611 ( 
.A1(n_1596),
.A2(n_1546),
.B1(n_1561),
.B2(n_1539),
.Y(n_1611)
);

AOI22xp33_ASAP7_75t_L g1612 ( 
.A1(n_1596),
.A2(n_1539),
.B1(n_1554),
.B2(n_1560),
.Y(n_1612)
);

AND2x2_ASAP7_75t_L g1613 ( 
.A(n_1592),
.B(n_1548),
.Y(n_1613)
);

AND2x2_ASAP7_75t_L g1614 ( 
.A(n_1592),
.B(n_1548),
.Y(n_1614)
);

HB1xp67_ASAP7_75t_L g1615 ( 
.A(n_1577),
.Y(n_1615)
);

NAND2xp5_ASAP7_75t_L g1616 ( 
.A(n_1590),
.B(n_1556),
.Y(n_1616)
);

INVx2_ASAP7_75t_L g1617 ( 
.A(n_1577),
.Y(n_1617)
);

OAI31xp33_ASAP7_75t_SL g1618 ( 
.A1(n_1580),
.A2(n_1573),
.A3(n_1540),
.B(n_1542),
.Y(n_1618)
);

HB1xp67_ASAP7_75t_L g1619 ( 
.A(n_1582),
.Y(n_1619)
);

INVx2_ASAP7_75t_L g1620 ( 
.A(n_1582),
.Y(n_1620)
);

INVxp67_ASAP7_75t_L g1621 ( 
.A(n_1586),
.Y(n_1621)
);

BUFx2_ASAP7_75t_L g1622 ( 
.A(n_1595),
.Y(n_1622)
);

NAND3xp33_ASAP7_75t_L g1623 ( 
.A(n_1580),
.B(n_1545),
.C(n_1474),
.Y(n_1623)
);

AND2x2_ASAP7_75t_L g1624 ( 
.A(n_1598),
.B(n_1597),
.Y(n_1624)
);

INVx1_ASAP7_75t_L g1625 ( 
.A(n_1615),
.Y(n_1625)
);

AND2x2_ASAP7_75t_L g1626 ( 
.A(n_1598),
.B(n_1597),
.Y(n_1626)
);

INVx2_ASAP7_75t_L g1627 ( 
.A(n_1602),
.Y(n_1627)
);

OR2x2_ASAP7_75t_L g1628 ( 
.A(n_1605),
.B(n_1582),
.Y(n_1628)
);

INVx3_ASAP7_75t_L g1629 ( 
.A(n_1600),
.Y(n_1629)
);

INVx1_ASAP7_75t_SL g1630 ( 
.A(n_1622),
.Y(n_1630)
);

AND2x2_ASAP7_75t_L g1631 ( 
.A(n_1598),
.B(n_1597),
.Y(n_1631)
);

HB1xp67_ASAP7_75t_L g1632 ( 
.A(n_1615),
.Y(n_1632)
);

INVx1_ASAP7_75t_L g1633 ( 
.A(n_1619),
.Y(n_1633)
);

HB1xp67_ASAP7_75t_L g1634 ( 
.A(n_1619),
.Y(n_1634)
);

AND2x2_ASAP7_75t_L g1635 ( 
.A(n_1598),
.B(n_1622),
.Y(n_1635)
);

AND2x2_ASAP7_75t_L g1636 ( 
.A(n_1622),
.B(n_1593),
.Y(n_1636)
);

AND2x4_ASAP7_75t_L g1637 ( 
.A(n_1607),
.B(n_1589),
.Y(n_1637)
);

NAND2xp5_ASAP7_75t_L g1638 ( 
.A(n_1605),
.B(n_1591),
.Y(n_1638)
);

AND2x2_ASAP7_75t_L g1639 ( 
.A(n_1600),
.B(n_1593),
.Y(n_1639)
);

OR2x2_ASAP7_75t_L g1640 ( 
.A(n_1605),
.B(n_1582),
.Y(n_1640)
);

AND2x2_ASAP7_75t_L g1641 ( 
.A(n_1600),
.B(n_1593),
.Y(n_1641)
);

AND2x2_ASAP7_75t_L g1642 ( 
.A(n_1600),
.B(n_1587),
.Y(n_1642)
);

AND2x2_ASAP7_75t_L g1643 ( 
.A(n_1606),
.B(n_1587),
.Y(n_1643)
);

NAND2xp5_ASAP7_75t_L g1644 ( 
.A(n_1616),
.B(n_1601),
.Y(n_1644)
);

NOR4xp25_ASAP7_75t_SL g1645 ( 
.A(n_1608),
.B(n_1544),
.C(n_1570),
.D(n_1549),
.Y(n_1645)
);

OR2x2_ASAP7_75t_L g1646 ( 
.A(n_1617),
.B(n_1620),
.Y(n_1646)
);

NAND2xp5_ASAP7_75t_L g1647 ( 
.A(n_1616),
.B(n_1591),
.Y(n_1647)
);

NOR3xp33_ASAP7_75t_L g1648 ( 
.A(n_1608),
.B(n_1586),
.C(n_1594),
.Y(n_1648)
);

INVx2_ASAP7_75t_L g1649 ( 
.A(n_1646),
.Y(n_1649)
);

INVx2_ASAP7_75t_L g1650 ( 
.A(n_1646),
.Y(n_1650)
);

INVx1_ASAP7_75t_L g1651 ( 
.A(n_1632),
.Y(n_1651)
);

AOI22xp33_ASAP7_75t_L g1652 ( 
.A1(n_1648),
.A2(n_1608),
.B1(n_1623),
.B2(n_1583),
.Y(n_1652)
);

INVxp67_ASAP7_75t_SL g1653 ( 
.A(n_1648),
.Y(n_1653)
);

INVxp67_ASAP7_75t_SL g1654 ( 
.A(n_1628),
.Y(n_1654)
);

AND2x2_ASAP7_75t_L g1655 ( 
.A(n_1635),
.B(n_1606),
.Y(n_1655)
);

AND2x2_ASAP7_75t_L g1656 ( 
.A(n_1635),
.B(n_1606),
.Y(n_1656)
);

INVx2_ASAP7_75t_L g1657 ( 
.A(n_1646),
.Y(n_1657)
);

INVx1_ASAP7_75t_L g1658 ( 
.A(n_1632),
.Y(n_1658)
);

INVx1_ASAP7_75t_L g1659 ( 
.A(n_1634),
.Y(n_1659)
);

OR2x2_ASAP7_75t_L g1660 ( 
.A(n_1628),
.B(n_1616),
.Y(n_1660)
);

NOR2xp33_ASAP7_75t_L g1661 ( 
.A(n_1638),
.B(n_1621),
.Y(n_1661)
);

INVx1_ASAP7_75t_L g1662 ( 
.A(n_1634),
.Y(n_1662)
);

INVx1_ASAP7_75t_L g1663 ( 
.A(n_1625),
.Y(n_1663)
);

INVx2_ASAP7_75t_L g1664 ( 
.A(n_1627),
.Y(n_1664)
);

AND2x2_ASAP7_75t_L g1665 ( 
.A(n_1635),
.B(n_1606),
.Y(n_1665)
);

BUFx2_ASAP7_75t_SL g1666 ( 
.A(n_1629),
.Y(n_1666)
);

INVx2_ASAP7_75t_L g1667 ( 
.A(n_1627),
.Y(n_1667)
);

NAND2xp5_ASAP7_75t_L g1668 ( 
.A(n_1638),
.B(n_1628),
.Y(n_1668)
);

INVx2_ASAP7_75t_SL g1669 ( 
.A(n_1629),
.Y(n_1669)
);

OR2x2_ASAP7_75t_L g1670 ( 
.A(n_1640),
.B(n_1609),
.Y(n_1670)
);

OR2x2_ASAP7_75t_L g1671 ( 
.A(n_1640),
.B(n_1609),
.Y(n_1671)
);

NAND2xp5_ASAP7_75t_L g1672 ( 
.A(n_1640),
.B(n_1621),
.Y(n_1672)
);

HB1xp67_ASAP7_75t_L g1673 ( 
.A(n_1642),
.Y(n_1673)
);

AND2x2_ASAP7_75t_L g1674 ( 
.A(n_1624),
.B(n_1610),
.Y(n_1674)
);

INVx1_ASAP7_75t_L g1675 ( 
.A(n_1625),
.Y(n_1675)
);

INVxp67_ASAP7_75t_L g1676 ( 
.A(n_1630),
.Y(n_1676)
);

INVx1_ASAP7_75t_L g1677 ( 
.A(n_1625),
.Y(n_1677)
);

OR2x2_ASAP7_75t_L g1678 ( 
.A(n_1647),
.B(n_1609),
.Y(n_1678)
);

HB1xp67_ASAP7_75t_L g1679 ( 
.A(n_1642),
.Y(n_1679)
);

INVx1_ASAP7_75t_L g1680 ( 
.A(n_1633),
.Y(n_1680)
);

INVx1_ASAP7_75t_L g1681 ( 
.A(n_1633),
.Y(n_1681)
);

INVx3_ASAP7_75t_L g1682 ( 
.A(n_1637),
.Y(n_1682)
);

AND2x2_ASAP7_75t_L g1683 ( 
.A(n_1624),
.B(n_1610),
.Y(n_1683)
);

NAND2xp5_ASAP7_75t_L g1684 ( 
.A(n_1647),
.B(n_1601),
.Y(n_1684)
);

AND2x2_ASAP7_75t_L g1685 ( 
.A(n_1624),
.B(n_1610),
.Y(n_1685)
);

INVx1_ASAP7_75t_L g1686 ( 
.A(n_1633),
.Y(n_1686)
);

OR2x2_ASAP7_75t_L g1687 ( 
.A(n_1644),
.B(n_1601),
.Y(n_1687)
);

AND2x4_ASAP7_75t_SL g1688 ( 
.A(n_1629),
.B(n_1567),
.Y(n_1688)
);

OR2x6_ASAP7_75t_L g1689 ( 
.A(n_1629),
.B(n_1623),
.Y(n_1689)
);

NAND2x1_ASAP7_75t_L g1690 ( 
.A(n_1629),
.B(n_1607),
.Y(n_1690)
);

INVx1_ASAP7_75t_L g1691 ( 
.A(n_1651),
.Y(n_1691)
);

NAND2xp5_ASAP7_75t_L g1692 ( 
.A(n_1653),
.B(n_1661),
.Y(n_1692)
);

NAND2xp5_ASAP7_75t_L g1693 ( 
.A(n_1653),
.B(n_1630),
.Y(n_1693)
);

INVx1_ASAP7_75t_L g1694 ( 
.A(n_1651),
.Y(n_1694)
);

INVx1_ASAP7_75t_L g1695 ( 
.A(n_1658),
.Y(n_1695)
);

HB1xp67_ASAP7_75t_L g1696 ( 
.A(n_1676),
.Y(n_1696)
);

INVx1_ASAP7_75t_SL g1697 ( 
.A(n_1655),
.Y(n_1697)
);

AND2x2_ASAP7_75t_L g1698 ( 
.A(n_1655),
.B(n_1636),
.Y(n_1698)
);

OR2x2_ASAP7_75t_L g1699 ( 
.A(n_1668),
.B(n_1644),
.Y(n_1699)
);

AND2x2_ASAP7_75t_L g1700 ( 
.A(n_1656),
.B(n_1665),
.Y(n_1700)
);

AND2x2_ASAP7_75t_L g1701 ( 
.A(n_1656),
.B(n_1636),
.Y(n_1701)
);

NAND2x1_ASAP7_75t_L g1702 ( 
.A(n_1689),
.B(n_1636),
.Y(n_1702)
);

NAND2xp5_ASAP7_75t_L g1703 ( 
.A(n_1672),
.B(n_1613),
.Y(n_1703)
);

OR2x2_ASAP7_75t_L g1704 ( 
.A(n_1668),
.B(n_1626),
.Y(n_1704)
);

INVx1_ASAP7_75t_L g1705 ( 
.A(n_1658),
.Y(n_1705)
);

INVx2_ASAP7_75t_L g1706 ( 
.A(n_1664),
.Y(n_1706)
);

NAND2xp5_ASAP7_75t_L g1707 ( 
.A(n_1672),
.B(n_1613),
.Y(n_1707)
);

INVx1_ASAP7_75t_L g1708 ( 
.A(n_1659),
.Y(n_1708)
);

AND2x2_ASAP7_75t_L g1709 ( 
.A(n_1665),
.B(n_1639),
.Y(n_1709)
);

NOR2xp33_ASAP7_75t_L g1710 ( 
.A(n_1676),
.B(n_1547),
.Y(n_1710)
);

AND2x2_ASAP7_75t_L g1711 ( 
.A(n_1689),
.B(n_1639),
.Y(n_1711)
);

OR2x2_ASAP7_75t_L g1712 ( 
.A(n_1670),
.B(n_1626),
.Y(n_1712)
);

AOI221x1_ASAP7_75t_L g1713 ( 
.A1(n_1659),
.A2(n_1623),
.B1(n_1603),
.B2(n_1604),
.C(n_1562),
.Y(n_1713)
);

NAND2xp5_ASAP7_75t_L g1714 ( 
.A(n_1654),
.B(n_1613),
.Y(n_1714)
);

AND2x2_ASAP7_75t_L g1715 ( 
.A(n_1689),
.B(n_1639),
.Y(n_1715)
);

NAND2xp5_ASAP7_75t_L g1716 ( 
.A(n_1654),
.B(n_1613),
.Y(n_1716)
);

AND2x2_ASAP7_75t_L g1717 ( 
.A(n_1689),
.B(n_1641),
.Y(n_1717)
);

NAND2xp5_ASAP7_75t_L g1718 ( 
.A(n_1652),
.B(n_1614),
.Y(n_1718)
);

INVx1_ASAP7_75t_L g1719 ( 
.A(n_1662),
.Y(n_1719)
);

INVx1_ASAP7_75t_L g1720 ( 
.A(n_1662),
.Y(n_1720)
);

OR2x2_ASAP7_75t_L g1721 ( 
.A(n_1670),
.B(n_1671),
.Y(n_1721)
);

AND2x2_ASAP7_75t_L g1722 ( 
.A(n_1689),
.B(n_1641),
.Y(n_1722)
);

OR2x2_ASAP7_75t_L g1723 ( 
.A(n_1671),
.B(n_1626),
.Y(n_1723)
);

INVxp33_ASAP7_75t_SL g1724 ( 
.A(n_1673),
.Y(n_1724)
);

NAND3xp33_ASAP7_75t_L g1725 ( 
.A(n_1663),
.B(n_1618),
.C(n_1645),
.Y(n_1725)
);

OR2x2_ASAP7_75t_L g1726 ( 
.A(n_1660),
.B(n_1631),
.Y(n_1726)
);

NAND2xp5_ASAP7_75t_L g1727 ( 
.A(n_1660),
.B(n_1673),
.Y(n_1727)
);

INVx1_ASAP7_75t_L g1728 ( 
.A(n_1696),
.Y(n_1728)
);

OA222x2_ASAP7_75t_L g1729 ( 
.A1(n_1718),
.A2(n_1618),
.B1(n_1645),
.B2(n_1587),
.C1(n_1678),
.C2(n_1594),
.Y(n_1729)
);

NAND2xp5_ASAP7_75t_SL g1730 ( 
.A(n_1725),
.B(n_1669),
.Y(n_1730)
);

AOI21xp5_ASAP7_75t_L g1731 ( 
.A1(n_1713),
.A2(n_1618),
.B(n_1690),
.Y(n_1731)
);

INVx1_ASAP7_75t_SL g1732 ( 
.A(n_1697),
.Y(n_1732)
);

INVx1_ASAP7_75t_L g1733 ( 
.A(n_1691),
.Y(n_1733)
);

INVx1_ASAP7_75t_L g1734 ( 
.A(n_1691),
.Y(n_1734)
);

OAI221xp5_ASAP7_75t_SL g1735 ( 
.A1(n_1692),
.A2(n_1679),
.B1(n_1611),
.B2(n_1678),
.C(n_1642),
.Y(n_1735)
);

AND2x2_ASAP7_75t_L g1736 ( 
.A(n_1700),
.B(n_1688),
.Y(n_1736)
);

OAI22xp33_ASAP7_75t_L g1737 ( 
.A1(n_1713),
.A2(n_1587),
.B1(n_1679),
.B2(n_1604),
.Y(n_1737)
);

A2O1A1O1Ixp25_ASAP7_75t_L g1738 ( 
.A1(n_1693),
.A2(n_1663),
.B(n_1675),
.C(n_1677),
.D(n_1686),
.Y(n_1738)
);

OAI21xp5_ASAP7_75t_SL g1739 ( 
.A1(n_1711),
.A2(n_1688),
.B(n_1641),
.Y(n_1739)
);

AOI21xp5_ASAP7_75t_L g1740 ( 
.A1(n_1702),
.A2(n_1690),
.B(n_1684),
.Y(n_1740)
);

OAI22xp5_ASAP7_75t_L g1741 ( 
.A1(n_1702),
.A2(n_1631),
.B1(n_1611),
.B2(n_1674),
.Y(n_1741)
);

AOI21xp5_ASAP7_75t_L g1742 ( 
.A1(n_1724),
.A2(n_1684),
.B(n_1669),
.Y(n_1742)
);

INVx1_ASAP7_75t_L g1743 ( 
.A(n_1694),
.Y(n_1743)
);

OR2x2_ASAP7_75t_L g1744 ( 
.A(n_1721),
.B(n_1687),
.Y(n_1744)
);

AND2x2_ASAP7_75t_L g1745 ( 
.A(n_1700),
.B(n_1688),
.Y(n_1745)
);

OAI21xp33_ASAP7_75t_L g1746 ( 
.A1(n_1711),
.A2(n_1643),
.B(n_1687),
.Y(n_1746)
);

INVx1_ASAP7_75t_L g1747 ( 
.A(n_1694),
.Y(n_1747)
);

AND2x2_ASAP7_75t_L g1748 ( 
.A(n_1698),
.B(n_1674),
.Y(n_1748)
);

INVx1_ASAP7_75t_L g1749 ( 
.A(n_1708),
.Y(n_1749)
);

AOI21xp33_ASAP7_75t_L g1750 ( 
.A1(n_1695),
.A2(n_1677),
.B(n_1675),
.Y(n_1750)
);

INVx1_ASAP7_75t_L g1751 ( 
.A(n_1708),
.Y(n_1751)
);

INVx1_ASAP7_75t_L g1752 ( 
.A(n_1719),
.Y(n_1752)
);

NOR3xp33_ASAP7_75t_SL g1753 ( 
.A(n_1727),
.B(n_1681),
.C(n_1680),
.Y(n_1753)
);

INVxp33_ASAP7_75t_L g1754 ( 
.A(n_1730),
.Y(n_1754)
);

AND2x2_ASAP7_75t_L g1755 ( 
.A(n_1736),
.B(n_1709),
.Y(n_1755)
);

OR2x6_ASAP7_75t_L g1756 ( 
.A(n_1728),
.B(n_1666),
.Y(n_1756)
);

NAND4xp75_ASAP7_75t_L g1757 ( 
.A(n_1730),
.B(n_1715),
.C(n_1717),
.D(n_1722),
.Y(n_1757)
);

OAI22xp33_ASAP7_75t_L g1758 ( 
.A1(n_1738),
.A2(n_1714),
.B1(n_1716),
.B2(n_1704),
.Y(n_1758)
);

NAND2xp5_ASAP7_75t_L g1759 ( 
.A(n_1732),
.B(n_1724),
.Y(n_1759)
);

OAI22xp5_ASAP7_75t_L g1760 ( 
.A1(n_1731),
.A2(n_1722),
.B1(n_1715),
.B2(n_1717),
.Y(n_1760)
);

OAI31xp33_ASAP7_75t_L g1761 ( 
.A1(n_1737),
.A2(n_1643),
.A3(n_1604),
.B(n_1603),
.Y(n_1761)
);

INVx1_ASAP7_75t_L g1762 ( 
.A(n_1733),
.Y(n_1762)
);

INVx1_ASAP7_75t_L g1763 ( 
.A(n_1733),
.Y(n_1763)
);

AOI22xp33_ASAP7_75t_SL g1764 ( 
.A1(n_1741),
.A2(n_1643),
.B1(n_1701),
.B2(n_1698),
.Y(n_1764)
);

AOI22xp5_ASAP7_75t_L g1765 ( 
.A1(n_1753),
.A2(n_1604),
.B1(n_1603),
.B2(n_1709),
.Y(n_1765)
);

INVx2_ASAP7_75t_L g1766 ( 
.A(n_1744),
.Y(n_1766)
);

NAND2xp5_ASAP7_75t_L g1767 ( 
.A(n_1744),
.B(n_1701),
.Y(n_1767)
);

AND2x2_ASAP7_75t_L g1768 ( 
.A(n_1736),
.B(n_1710),
.Y(n_1768)
);

INVx1_ASAP7_75t_L g1769 ( 
.A(n_1734),
.Y(n_1769)
);

NAND2xp5_ASAP7_75t_L g1770 ( 
.A(n_1748),
.B(n_1721),
.Y(n_1770)
);

AND2x2_ASAP7_75t_L g1771 ( 
.A(n_1745),
.B(n_1683),
.Y(n_1771)
);

NAND2xp5_ASAP7_75t_L g1772 ( 
.A(n_1748),
.B(n_1705),
.Y(n_1772)
);

AOI22xp5_ASAP7_75t_L g1773 ( 
.A1(n_1746),
.A2(n_1603),
.B1(n_1581),
.B2(n_1599),
.Y(n_1773)
);

INVx2_ASAP7_75t_L g1774 ( 
.A(n_1745),
.Y(n_1774)
);

INVx2_ASAP7_75t_L g1775 ( 
.A(n_1755),
.Y(n_1775)
);

INVx1_ASAP7_75t_L g1776 ( 
.A(n_1766),
.Y(n_1776)
);

AOI32xp33_ASAP7_75t_L g1777 ( 
.A1(n_1754),
.A2(n_1729),
.A3(n_1735),
.B1(n_1752),
.B2(n_1749),
.Y(n_1777)
);

NOR2xp33_ASAP7_75t_L g1778 ( 
.A(n_1754),
.B(n_1739),
.Y(n_1778)
);

AND2x2_ASAP7_75t_L g1779 ( 
.A(n_1768),
.B(n_1683),
.Y(n_1779)
);

OR2x2_ASAP7_75t_L g1780 ( 
.A(n_1770),
.B(n_1712),
.Y(n_1780)
);

INVxp67_ASAP7_75t_L g1781 ( 
.A(n_1759),
.Y(n_1781)
);

OR2x2_ASAP7_75t_L g1782 ( 
.A(n_1767),
.B(n_1712),
.Y(n_1782)
);

AOI21xp33_ASAP7_75t_SL g1783 ( 
.A1(n_1758),
.A2(n_1750),
.B(n_1747),
.Y(n_1783)
);

AOI211xp5_ASAP7_75t_L g1784 ( 
.A1(n_1758),
.A2(n_1742),
.B(n_1743),
.C(n_1751),
.Y(n_1784)
);

INVx2_ASAP7_75t_L g1785 ( 
.A(n_1771),
.Y(n_1785)
);

INVx1_ASAP7_75t_L g1786 ( 
.A(n_1766),
.Y(n_1786)
);

NAND2xp5_ASAP7_75t_SL g1787 ( 
.A(n_1784),
.B(n_1774),
.Y(n_1787)
);

NAND2xp5_ASAP7_75t_L g1788 ( 
.A(n_1779),
.B(n_1774),
.Y(n_1788)
);

INVx1_ASAP7_75t_SL g1789 ( 
.A(n_1775),
.Y(n_1789)
);

AOI211x1_ASAP7_75t_L g1790 ( 
.A1(n_1776),
.A2(n_1760),
.B(n_1772),
.C(n_1740),
.Y(n_1790)
);

NAND2xp5_ASAP7_75t_L g1791 ( 
.A(n_1785),
.B(n_1757),
.Y(n_1791)
);

NAND2xp5_ASAP7_75t_SL g1792 ( 
.A(n_1784),
.B(n_1764),
.Y(n_1792)
);

NAND2xp5_ASAP7_75t_L g1793 ( 
.A(n_1781),
.B(n_1769),
.Y(n_1793)
);

INVx1_ASAP7_75t_L g1794 ( 
.A(n_1786),
.Y(n_1794)
);

AOI31xp33_ASAP7_75t_L g1795 ( 
.A1(n_1781),
.A2(n_1764),
.A3(n_1762),
.B(n_1763),
.Y(n_1795)
);

AOI22xp5_ASAP7_75t_L g1796 ( 
.A1(n_1792),
.A2(n_1778),
.B1(n_1765),
.B2(n_1780),
.Y(n_1796)
);

AOI221xp5_ASAP7_75t_L g1797 ( 
.A1(n_1795),
.A2(n_1783),
.B1(n_1777),
.B2(n_1761),
.C(n_1773),
.Y(n_1797)
);

NAND4xp25_ASAP7_75t_L g1798 ( 
.A(n_1790),
.B(n_1791),
.C(n_1788),
.D(n_1789),
.Y(n_1798)
);

NAND4xp25_ASAP7_75t_L g1799 ( 
.A(n_1787),
.B(n_1782),
.C(n_1719),
.D(n_1720),
.Y(n_1799)
);

AOI22xp5_ASAP7_75t_L g1800 ( 
.A1(n_1794),
.A2(n_1756),
.B1(n_1706),
.B2(n_1599),
.Y(n_1800)
);

INVx1_ASAP7_75t_L g1801 ( 
.A(n_1799),
.Y(n_1801)
);

NOR3xp33_ASAP7_75t_SL g1802 ( 
.A(n_1798),
.B(n_1793),
.C(n_1756),
.Y(n_1802)
);

NAND2xp5_ASAP7_75t_L g1803 ( 
.A(n_1796),
.B(n_1756),
.Y(n_1803)
);

AOI211xp5_ASAP7_75t_L g1804 ( 
.A1(n_1797),
.A2(n_1723),
.B(n_1726),
.C(n_1704),
.Y(n_1804)
);

NOR2xp33_ASAP7_75t_L g1805 ( 
.A(n_1800),
.B(n_1669),
.Y(n_1805)
);

O2A1O1Ixp33_ASAP7_75t_L g1806 ( 
.A1(n_1798),
.A2(n_1699),
.B(n_1706),
.C(n_1723),
.Y(n_1806)
);

XNOR2xp5_ASAP7_75t_L g1807 ( 
.A(n_1804),
.B(n_1567),
.Y(n_1807)
);

NAND4xp75_ASAP7_75t_L g1808 ( 
.A(n_1802),
.B(n_1474),
.C(n_1707),
.D(n_1703),
.Y(n_1808)
);

INVx1_ASAP7_75t_L g1809 ( 
.A(n_1806),
.Y(n_1809)
);

NAND4xp75_ASAP7_75t_L g1810 ( 
.A(n_1803),
.B(n_1685),
.C(n_1649),
.D(n_1657),
.Y(n_1810)
);

NAND4xp75_ASAP7_75t_L g1811 ( 
.A(n_1801),
.B(n_1685),
.C(n_1649),
.D(n_1657),
.Y(n_1811)
);

OA22x2_ASAP7_75t_L g1812 ( 
.A1(n_1807),
.A2(n_1666),
.B1(n_1805),
.B2(n_1682),
.Y(n_1812)
);

A2O1A1Ixp33_ASAP7_75t_SL g1813 ( 
.A1(n_1809),
.A2(n_1682),
.B(n_1686),
.C(n_1681),
.Y(n_1813)
);

INVx1_ASAP7_75t_L g1814 ( 
.A(n_1811),
.Y(n_1814)
);

HB1xp67_ASAP7_75t_L g1815 ( 
.A(n_1814),
.Y(n_1815)
);

INVx1_ASAP7_75t_L g1816 ( 
.A(n_1815),
.Y(n_1816)
);

OA21x2_ASAP7_75t_L g1817 ( 
.A1(n_1816),
.A2(n_1810),
.B(n_1808),
.Y(n_1817)
);

INVx2_ASAP7_75t_SL g1818 ( 
.A(n_1816),
.Y(n_1818)
);

XNOR2xp5_ASAP7_75t_L g1819 ( 
.A(n_1817),
.B(n_1812),
.Y(n_1819)
);

AOI22xp5_ASAP7_75t_L g1820 ( 
.A1(n_1818),
.A2(n_1813),
.B1(n_1657),
.B2(n_1650),
.Y(n_1820)
);

OAI22xp5_ASAP7_75t_SL g1821 ( 
.A1(n_1819),
.A2(n_1817),
.B1(n_1726),
.B2(n_1699),
.Y(n_1821)
);

NAND2xp5_ASAP7_75t_SL g1822 ( 
.A(n_1820),
.B(n_1649),
.Y(n_1822)
);

INVx2_ASAP7_75t_L g1823 ( 
.A(n_1821),
.Y(n_1823)
);

AOI22xp5_ASAP7_75t_L g1824 ( 
.A1(n_1823),
.A2(n_1822),
.B1(n_1650),
.B2(n_1667),
.Y(n_1824)
);

HB1xp67_ASAP7_75t_L g1825 ( 
.A(n_1824),
.Y(n_1825)
);

OAI221xp5_ASAP7_75t_R g1826 ( 
.A1(n_1825),
.A2(n_1682),
.B1(n_1680),
.B2(n_1650),
.C(n_1612),
.Y(n_1826)
);

AOI211xp5_ASAP7_75t_L g1827 ( 
.A1(n_1826),
.A2(n_1529),
.B(n_1536),
.C(n_1568),
.Y(n_1827)
);


endmodule