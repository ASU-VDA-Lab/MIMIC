module real_aes_505_n_99 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_43, n_96, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_817, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_816, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_99);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_817;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_816;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_99;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_800;
wire n_618;
wire n_778;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_357;
wire n_287;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_421;
wire n_364;
wire n_555;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_537;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_292;
wire n_539;
wire n_400;
wire n_626;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_781;
wire n_748;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_812;
wire n_565;
wire n_443;
wire n_782;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_808;
wire n_770;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_449;
wire n_417;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_783;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_807;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_790;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_735;
wire n_728;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_810;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_749;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_148;
wire n_498;
wire n_481;
wire n_765;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_789;
wire n_268;
wire n_544;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_809;
wire n_482;
wire n_520;
wire n_679;
wire n_633;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_753;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_771;
wire n_524;
wire n_219;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_740;
wire n_371;
wire n_698;
wire n_166;
wire n_103;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_804;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_802;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_554;
wire n_475;
wire n_264;
wire n_798;
wire n_797;
wire n_237;
wire n_668;
NAND2xp5_ASAP7_75t_L g531 ( .A(n_0), .B(n_217), .Y(n_531) );
NAND2xp5_ASAP7_75t_L g106 ( .A(n_1), .B(n_107), .Y(n_106) );
INVx1_ASAP7_75t_L g145 ( .A(n_2), .Y(n_145) );
NAND2xp5_ASAP7_75t_L g547 ( .A(n_3), .B(n_510), .Y(n_547) );
NAND2xp33_ASAP7_75t_SL g587 ( .A(n_4), .B(n_166), .Y(n_587) );
NAND2xp5_ASAP7_75t_SL g208 ( .A(n_5), .B(n_201), .Y(n_208) );
INVx1_ASAP7_75t_L g580 ( .A(n_6), .Y(n_580) );
INVx1_ASAP7_75t_L g188 ( .A(n_7), .Y(n_188) );
CKINVDCx16_ASAP7_75t_R g107 ( .A(n_8), .Y(n_107) );
CKINVDCx5p33_ASAP7_75t_R g276 ( .A(n_9), .Y(n_276) );
AND2x2_ASAP7_75t_L g545 ( .A(n_10), .B(n_169), .Y(n_545) );
INVx2_ASAP7_75t_L g137 ( .A(n_11), .Y(n_137) );
CKINVDCx16_ASAP7_75t_R g111 ( .A(n_12), .Y(n_111) );
INVx1_ASAP7_75t_L g218 ( .A(n_13), .Y(n_218) );
AOI221x1_ASAP7_75t_L g583 ( .A1(n_14), .A2(n_134), .B1(n_512), .B2(n_584), .C(n_586), .Y(n_583) );
NAND2xp5_ASAP7_75t_SL g509 ( .A(n_15), .B(n_510), .Y(n_509) );
INVx1_ASAP7_75t_L g115 ( .A(n_16), .Y(n_115) );
INVx1_ASAP7_75t_L g215 ( .A(n_17), .Y(n_215) );
INVx1_ASAP7_75t_SL g230 ( .A(n_18), .Y(n_230) );
NAND2xp5_ASAP7_75t_SL g204 ( .A(n_19), .B(n_160), .Y(n_204) );
AOI33xp33_ASAP7_75t_L g180 ( .A1(n_20), .A2(n_49), .A3(n_142), .B1(n_153), .B2(n_181), .B3(n_182), .Y(n_180) );
AOI221xp5_ASAP7_75t_SL g521 ( .A1(n_21), .A2(n_40), .B1(n_510), .B2(n_512), .C(n_522), .Y(n_521) );
AOI21xp5_ASAP7_75t_L g548 ( .A1(n_22), .A2(n_512), .B(n_549), .Y(n_548) );
NAND2xp5_ASAP7_75t_L g550 ( .A(n_23), .B(n_217), .Y(n_550) );
INVx1_ASAP7_75t_L g270 ( .A(n_24), .Y(n_270) );
OA21x2_ASAP7_75t_L g136 ( .A1(n_25), .A2(n_87), .B(n_137), .Y(n_136) );
OR2x2_ASAP7_75t_L g170 ( .A(n_25), .B(n_87), .Y(n_170) );
NAND2xp5_ASAP7_75t_L g515 ( .A(n_26), .B(n_220), .Y(n_515) );
INVxp67_ASAP7_75t_L g582 ( .A(n_27), .Y(n_582) );
AND2x2_ASAP7_75t_L g569 ( .A(n_28), .B(n_168), .Y(n_569) );
NAND2xp5_ASAP7_75t_L g227 ( .A(n_29), .B(n_140), .Y(n_227) );
AOI21xp5_ASAP7_75t_L g529 ( .A1(n_30), .A2(n_512), .B(n_530), .Y(n_529) );
NAND2xp5_ASAP7_75t_L g372 ( .A(n_31), .B(n_373), .Y(n_372) );
CKINVDCx16_ASAP7_75t_R g496 ( .A(n_31), .Y(n_496) );
OAI22x1_ASAP7_75t_R g796 ( .A1(n_31), .A2(n_35), .B1(n_496), .B2(n_797), .Y(n_796) );
NAND2xp5_ASAP7_75t_L g523 ( .A(n_32), .B(n_220), .Y(n_523) );
AND2x2_ASAP7_75t_L g147 ( .A(n_33), .B(n_148), .Y(n_147) );
INVx1_ASAP7_75t_L g152 ( .A(n_33), .Y(n_152) );
AND2x2_ASAP7_75t_L g166 ( .A(n_33), .B(n_145), .Y(n_166) );
OR2x6_ASAP7_75t_L g113 ( .A(n_34), .B(n_114), .Y(n_113) );
AOI222xp33_ASAP7_75t_L g99 ( .A1(n_35), .A2(n_100), .B1(n_117), .B2(n_789), .C1(n_804), .C2(n_808), .Y(n_99) );
CKINVDCx20_ASAP7_75t_R g797 ( .A(n_35), .Y(n_797) );
CKINVDCx20_ASAP7_75t_R g272 ( .A(n_36), .Y(n_272) );
NAND2xp5_ASAP7_75t_L g139 ( .A(n_37), .B(n_140), .Y(n_139) );
AOI22xp5_ASAP7_75t_L g196 ( .A1(n_38), .A2(n_135), .B1(n_197), .B2(n_201), .Y(n_196) );
NAND2xp5_ASAP7_75t_L g205 ( .A(n_39), .B(n_206), .Y(n_205) );
AOI22xp5_ASAP7_75t_L g541 ( .A1(n_41), .A2(n_79), .B1(n_150), .B2(n_512), .Y(n_541) );
NAND2xp5_ASAP7_75t_L g231 ( .A(n_42), .B(n_160), .Y(n_231) );
NAND2xp5_ASAP7_75t_L g567 ( .A(n_43), .B(n_217), .Y(n_567) );
NAND2xp5_ASAP7_75t_SL g190 ( .A(n_44), .B(n_175), .Y(n_190) );
NAND2xp5_ASAP7_75t_L g189 ( .A(n_45), .B(n_160), .Y(n_189) );
CKINVDCx5p33_ASAP7_75t_R g200 ( .A(n_46), .Y(n_200) );
AND2x2_ASAP7_75t_L g534 ( .A(n_47), .B(n_168), .Y(n_534) );
NAND2xp5_ASAP7_75t_L g525 ( .A(n_48), .B(n_168), .Y(n_525) );
NAND2xp5_ASAP7_75t_L g159 ( .A(n_50), .B(n_160), .Y(n_159) );
INVx1_ASAP7_75t_L g143 ( .A(n_51), .Y(n_143) );
INVx1_ASAP7_75t_L g162 ( .A(n_51), .Y(n_162) );
AND2x2_ASAP7_75t_L g167 ( .A(n_52), .B(n_168), .Y(n_167) );
AOI221xp5_ASAP7_75t_L g186 ( .A1(n_53), .A2(n_72), .B1(n_140), .B2(n_150), .C(n_187), .Y(n_186) );
NAND2xp5_ASAP7_75t_L g242 ( .A(n_54), .B(n_140), .Y(n_242) );
NAND2xp5_ASAP7_75t_SL g568 ( .A(n_55), .B(n_510), .Y(n_568) );
CKINVDCx20_ASAP7_75t_R g786 ( .A(n_56), .Y(n_786) );
NAND2xp5_ASAP7_75t_L g278 ( .A(n_57), .B(n_135), .Y(n_278) );
AOI21xp5_ASAP7_75t_SL g238 ( .A1(n_58), .A2(n_150), .B(n_239), .Y(n_238) );
AND2x2_ASAP7_75t_L g560 ( .A(n_59), .B(n_168), .Y(n_560) );
NAND2xp5_ASAP7_75t_L g532 ( .A(n_60), .B(n_220), .Y(n_532) );
CKINVDCx20_ASAP7_75t_R g803 ( .A(n_61), .Y(n_803) );
INVx1_ASAP7_75t_L g211 ( .A(n_62), .Y(n_211) );
AND2x2_ASAP7_75t_SL g516 ( .A(n_63), .B(n_169), .Y(n_516) );
NAND2xp5_ASAP7_75t_L g558 ( .A(n_64), .B(n_217), .Y(n_558) );
AOI21xp5_ASAP7_75t_L g564 ( .A1(n_65), .A2(n_512), .B(n_565), .Y(n_564) );
INVx1_ASAP7_75t_L g157 ( .A(n_66), .Y(n_157) );
NAND2xp5_ASAP7_75t_L g551 ( .A(n_67), .B(n_220), .Y(n_551) );
AND2x2_ASAP7_75t_SL g542 ( .A(n_68), .B(n_175), .Y(n_542) );
AOI21xp5_ASAP7_75t_L g149 ( .A1(n_69), .A2(n_150), .B(n_156), .Y(n_149) );
INVx1_ASAP7_75t_L g148 ( .A(n_70), .Y(n_148) );
INVx1_ASAP7_75t_L g164 ( .A(n_70), .Y(n_164) );
NAND2xp5_ASAP7_75t_L g183 ( .A(n_71), .B(n_140), .Y(n_183) );
AND2x2_ASAP7_75t_L g232 ( .A(n_73), .B(n_134), .Y(n_232) );
INVx1_ASAP7_75t_L g212 ( .A(n_74), .Y(n_212) );
AOI21xp5_ASAP7_75t_L g228 ( .A1(n_75), .A2(n_150), .B(n_229), .Y(n_228) );
A2O1A1Ixp33_ASAP7_75t_L g202 ( .A1(n_76), .A2(n_150), .B(n_174), .C(n_203), .Y(n_202) );
AOI22xp5_ASAP7_75t_L g540 ( .A1(n_77), .A2(n_82), .B1(n_140), .B2(n_510), .Y(n_540) );
NAND2xp5_ASAP7_75t_SL g559 ( .A(n_78), .B(n_510), .Y(n_559) );
INVx1_ASAP7_75t_L g116 ( .A(n_80), .Y(n_116) );
AND2x2_ASAP7_75t_SL g236 ( .A(n_81), .B(n_134), .Y(n_236) );
AOI22xp5_ASAP7_75t_L g177 ( .A1(n_83), .A2(n_150), .B1(n_178), .B2(n_179), .Y(n_177) );
NAND2xp5_ASAP7_75t_L g514 ( .A(n_84), .B(n_217), .Y(n_514) );
NAND2xp5_ASAP7_75t_L g524 ( .A(n_85), .B(n_217), .Y(n_524) );
AOI21xp5_ASAP7_75t_L g555 ( .A1(n_86), .A2(n_512), .B(n_556), .Y(n_555) );
INVx1_ASAP7_75t_L g240 ( .A(n_88), .Y(n_240) );
NAND2xp5_ASAP7_75t_L g557 ( .A(n_89), .B(n_220), .Y(n_557) );
AND2x2_ASAP7_75t_L g184 ( .A(n_90), .B(n_134), .Y(n_184) );
CKINVDCx20_ASAP7_75t_R g780 ( .A(n_91), .Y(n_780) );
A2O1A1Ixp33_ASAP7_75t_L g267 ( .A1(n_92), .A2(n_268), .B(n_269), .C(n_271), .Y(n_267) );
NAND2xp5_ASAP7_75t_L g533 ( .A(n_93), .B(n_510), .Y(n_533) );
INVxp67_ASAP7_75t_L g585 ( .A(n_94), .Y(n_585) );
NAND2xp5_ASAP7_75t_L g566 ( .A(n_95), .B(n_220), .Y(n_566) );
AOI21xp5_ASAP7_75t_L g511 ( .A1(n_96), .A2(n_512), .B(n_513), .Y(n_511) );
BUFx2_ASAP7_75t_L g108 ( .A(n_97), .Y(n_108) );
BUFx2_ASAP7_75t_SL g812 ( .A(n_97), .Y(n_812) );
NAND2xp5_ASAP7_75t_L g241 ( .A(n_98), .B(n_160), .Y(n_241) );
INVx1_ASAP7_75t_SL g100 ( .A(n_101), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_102), .Y(n_101) );
AND2x2_ASAP7_75t_L g102 ( .A(n_103), .B(n_109), .Y(n_102) );
INVxp67_ASAP7_75t_L g103 ( .A(n_104), .Y(n_103) );
NAND2xp5_ASAP7_75t_SL g104 ( .A(n_105), .B(n_108), .Y(n_104) );
INVx2_ASAP7_75t_L g105 ( .A(n_106), .Y(n_105) );
OR2x2_ASAP7_75t_SL g807 ( .A(n_106), .B(n_108), .Y(n_807) );
AOI21xp5_ASAP7_75t_L g809 ( .A1(n_106), .A2(n_810), .B(n_813), .Y(n_809) );
NOR2xp33_ASAP7_75t_SL g802 ( .A(n_109), .B(n_803), .Y(n_802) );
BUFx2_ASAP7_75t_L g109 ( .A(n_110), .Y(n_109) );
BUFx3_ASAP7_75t_L g793 ( .A(n_110), .Y(n_793) );
BUFx2_ASAP7_75t_L g814 ( .A(n_110), .Y(n_814) );
NAND2xp5_ASAP7_75t_L g110 ( .A(n_111), .B(n_112), .Y(n_110) );
AND2x6_ASAP7_75t_SL g122 ( .A(n_111), .B(n_113), .Y(n_122) );
OR2x6_ASAP7_75t_SL g500 ( .A(n_111), .B(n_112), .Y(n_500) );
OR2x2_ASAP7_75t_L g788 ( .A(n_111), .B(n_113), .Y(n_788) );
CKINVDCx5p33_ASAP7_75t_R g112 ( .A(n_113), .Y(n_112) );
NAND2xp5_ASAP7_75t_L g114 ( .A(n_115), .B(n_116), .Y(n_114) );
HB1xp67_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
OAI21xp5_ASAP7_75t_L g118 ( .A1(n_119), .A2(n_780), .B(n_781), .Y(n_118) );
INVxp33_ASAP7_75t_SL g119 ( .A(n_120), .Y(n_119) );
OAI22xp5_ASAP7_75t_L g120 ( .A1(n_121), .A2(n_123), .B1(n_498), .B2(n_501), .Y(n_120) );
OAI21x1_ASAP7_75t_L g782 ( .A1(n_121), .A2(n_783), .B(n_784), .Y(n_782) );
CKINVDCx11_ASAP7_75t_R g121 ( .A(n_122), .Y(n_121) );
INVx2_ASAP7_75t_L g783 ( .A(n_123), .Y(n_783) );
OR2x2_ASAP7_75t_L g123 ( .A(n_124), .B(n_493), .Y(n_123) );
NOR4xp25_ASAP7_75t_L g124 ( .A(n_125), .B(n_372), .C(n_396), .D(n_462), .Y(n_124) );
AOI22xp5_ASAP7_75t_L g497 ( .A1(n_125), .A2(n_396), .B1(n_496), .B2(n_816), .Y(n_497) );
INVx2_ASAP7_75t_L g801 ( .A(n_125), .Y(n_801) );
NAND3x1_ASAP7_75t_L g125 ( .A(n_126), .B(n_324), .C(n_358), .Y(n_125) );
NOR3x1_ASAP7_75t_L g126 ( .A(n_127), .B(n_283), .C(n_303), .Y(n_126) );
NAND2xp5_ASAP7_75t_L g127 ( .A(n_128), .B(n_258), .Y(n_127) );
AOI22xp5_ASAP7_75t_L g128 ( .A1(n_129), .A2(n_191), .B1(n_247), .B2(n_255), .Y(n_128) );
AND2x2_ASAP7_75t_L g129 ( .A(n_130), .B(n_171), .Y(n_129) );
AND2x2_ASAP7_75t_L g422 ( .A(n_130), .B(n_352), .Y(n_422) );
INVx1_ASAP7_75t_L g429 ( .A(n_130), .Y(n_429) );
NAND2xp5_ASAP7_75t_L g444 ( .A(n_130), .B(n_445), .Y(n_444) );
NAND2xp5_ASAP7_75t_L g481 ( .A(n_130), .B(n_292), .Y(n_481) );
OR2x2_ASAP7_75t_L g491 ( .A(n_130), .B(n_492), .Y(n_491) );
INVx3_ASAP7_75t_L g130 ( .A(n_131), .Y(n_130) );
NAND2x1p5_ASAP7_75t_L g312 ( .A(n_131), .B(n_249), .Y(n_312) );
AND2x4_ASAP7_75t_L g340 ( .A(n_131), .B(n_254), .Y(n_340) );
INVx3_ASAP7_75t_L g131 ( .A(n_132), .Y(n_131) );
AND2x2_ASAP7_75t_L g288 ( .A(n_132), .B(n_289), .Y(n_288) );
NAND2xp5_ASAP7_75t_L g378 ( .A(n_132), .B(n_173), .Y(n_378) );
HB1xp67_ASAP7_75t_L g392 ( .A(n_132), .Y(n_392) );
NAND2xp5_ASAP7_75t_L g415 ( .A(n_132), .B(n_265), .Y(n_415) );
AO21x2_ASAP7_75t_L g132 ( .A1(n_133), .A2(n_138), .B(n_167), .Y(n_132) );
AO21x2_ASAP7_75t_L g253 ( .A1(n_133), .A2(n_138), .B(n_167), .Y(n_253) );
OAI22xp5_ASAP7_75t_L g266 ( .A1(n_133), .A2(n_134), .B1(n_267), .B2(n_272), .Y(n_266) );
INVx3_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
INVx4_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
NAND2xp5_ASAP7_75t_L g274 ( .A(n_135), .B(n_275), .Y(n_274) );
AOI21x1_ASAP7_75t_L g527 ( .A1(n_135), .A2(n_528), .B(n_534), .Y(n_527) );
INVx3_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
BUFx4f_ASAP7_75t_L g175 ( .A(n_136), .Y(n_175) );
AND2x2_ASAP7_75t_SL g169 ( .A(n_137), .B(n_170), .Y(n_169) );
AND2x4_ASAP7_75t_L g201 ( .A(n_137), .B(n_170), .Y(n_201) );
NAND2xp5_ASAP7_75t_L g138 ( .A(n_139), .B(n_149), .Y(n_138) );
INVx1_ASAP7_75t_L g279 ( .A(n_140), .Y(n_279) );
AOI22xp5_ASAP7_75t_L g578 ( .A1(n_140), .A2(n_150), .B1(n_579), .B2(n_581), .Y(n_578) );
AND2x4_ASAP7_75t_L g140 ( .A(n_141), .B(n_146), .Y(n_140) );
INVx1_ASAP7_75t_L g198 ( .A(n_141), .Y(n_198) );
AND2x2_ASAP7_75t_L g141 ( .A(n_142), .B(n_144), .Y(n_141) );
OR2x6_ASAP7_75t_L g158 ( .A(n_142), .B(n_154), .Y(n_158) );
INVxp33_ASAP7_75t_L g181 ( .A(n_142), .Y(n_181) );
INVx2_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
AND2x2_ASAP7_75t_L g155 ( .A(n_143), .B(n_145), .Y(n_155) );
AND2x4_ASAP7_75t_L g220 ( .A(n_143), .B(n_163), .Y(n_220) );
HB1xp67_ASAP7_75t_L g144 ( .A(n_145), .Y(n_144) );
INVx1_ASAP7_75t_L g199 ( .A(n_146), .Y(n_199) );
BUFx3_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
AND2x6_ASAP7_75t_L g512 ( .A(n_147), .B(n_155), .Y(n_512) );
INVx2_ASAP7_75t_L g154 ( .A(n_148), .Y(n_154) );
AND2x6_ASAP7_75t_L g217 ( .A(n_148), .B(n_161), .Y(n_217) );
INVxp67_ASAP7_75t_L g277 ( .A(n_150), .Y(n_277) );
AND2x4_ASAP7_75t_L g150 ( .A(n_151), .B(n_155), .Y(n_150) );
NOR2x1p5_ASAP7_75t_L g151 ( .A(n_152), .B(n_153), .Y(n_151) );
INVx1_ASAP7_75t_L g182 ( .A(n_153), .Y(n_182) );
INVx3_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
O2A1O1Ixp33_ASAP7_75t_L g156 ( .A1(n_157), .A2(n_158), .B(n_159), .C(n_165), .Y(n_156) );
O2A1O1Ixp33_ASAP7_75t_SL g187 ( .A1(n_158), .A2(n_165), .B(n_188), .C(n_189), .Y(n_187) );
INVx2_ASAP7_75t_L g206 ( .A(n_158), .Y(n_206) );
OAI22xp5_ASAP7_75t_L g210 ( .A1(n_158), .A2(n_211), .B1(n_212), .B2(n_213), .Y(n_210) );
O2A1O1Ixp33_ASAP7_75t_SL g229 ( .A1(n_158), .A2(n_165), .B(n_230), .C(n_231), .Y(n_229) );
O2A1O1Ixp33_ASAP7_75t_L g239 ( .A1(n_158), .A2(n_165), .B(n_240), .C(n_241), .Y(n_239) );
INVxp67_ASAP7_75t_L g268 ( .A(n_158), .Y(n_268) );
INVx1_ASAP7_75t_L g213 ( .A(n_160), .Y(n_213) );
AND2x4_ASAP7_75t_L g510 ( .A(n_160), .B(n_166), .Y(n_510) );
AND2x4_ASAP7_75t_L g160 ( .A(n_161), .B(n_163), .Y(n_160) );
INVx2_ASAP7_75t_L g161 ( .A(n_162), .Y(n_161) );
INVx2_ASAP7_75t_L g163 ( .A(n_164), .Y(n_163) );
INVx1_ASAP7_75t_L g178 ( .A(n_165), .Y(n_178) );
AOI21xp5_ASAP7_75t_L g203 ( .A1(n_165), .A2(n_204), .B(n_205), .Y(n_203) );
NOR2xp33_ASAP7_75t_L g221 ( .A(n_165), .B(n_201), .Y(n_221) );
AOI21xp5_ASAP7_75t_L g513 ( .A1(n_165), .A2(n_514), .B(n_515), .Y(n_513) );
AOI21xp5_ASAP7_75t_L g522 ( .A1(n_165), .A2(n_523), .B(n_524), .Y(n_522) );
AOI21xp5_ASAP7_75t_L g530 ( .A1(n_165), .A2(n_531), .B(n_532), .Y(n_530) );
AOI21xp5_ASAP7_75t_L g549 ( .A1(n_165), .A2(n_550), .B(n_551), .Y(n_549) );
AOI21xp5_ASAP7_75t_L g556 ( .A1(n_165), .A2(n_557), .B(n_558), .Y(n_556) );
AOI21xp5_ASAP7_75t_L g565 ( .A1(n_165), .A2(n_566), .B(n_567), .Y(n_565) );
INVx5_ASAP7_75t_L g165 ( .A(n_166), .Y(n_165) );
HB1xp67_ASAP7_75t_L g271 ( .A(n_166), .Y(n_271) );
CKINVDCx5p33_ASAP7_75t_R g225 ( .A(n_168), .Y(n_225) );
OA21x2_ASAP7_75t_L g520 ( .A1(n_168), .A2(n_521), .B(n_525), .Y(n_520) );
BUFx6f_ASAP7_75t_L g168 ( .A(n_169), .Y(n_168) );
NAND2xp5_ASAP7_75t_L g428 ( .A(n_171), .B(n_429), .Y(n_428) );
AND2x2_ASAP7_75t_L g486 ( .A(n_171), .B(n_323), .Y(n_486) );
INVx2_ASAP7_75t_L g171 ( .A(n_172), .Y(n_171) );
OR2x2_ASAP7_75t_L g476 ( .A(n_172), .B(n_415), .Y(n_476) );
NAND2xp5_ASAP7_75t_L g172 ( .A(n_173), .B(n_185), .Y(n_172) );
INVx2_ASAP7_75t_L g254 ( .A(n_173), .Y(n_254) );
AO21x2_ASAP7_75t_L g173 ( .A1(n_174), .A2(n_176), .B(n_184), .Y(n_173) );
AO21x2_ASAP7_75t_L g282 ( .A1(n_174), .A2(n_176), .B(n_184), .Y(n_282) );
AOI21x1_ASAP7_75t_L g538 ( .A1(n_174), .A2(n_539), .B(n_542), .Y(n_538) );
INVx2_ASAP7_75t_SL g174 ( .A(n_175), .Y(n_174) );
OA21x2_ASAP7_75t_L g185 ( .A1(n_175), .A2(n_186), .B(n_190), .Y(n_185) );
AOI21xp5_ASAP7_75t_L g508 ( .A1(n_175), .A2(n_509), .B(n_511), .Y(n_508) );
NAND2xp5_ASAP7_75t_SL g176 ( .A(n_177), .B(n_183), .Y(n_176) );
INVx1_ASAP7_75t_L g179 ( .A(n_180), .Y(n_179) );
INVx1_ASAP7_75t_L g250 ( .A(n_185), .Y(n_250) );
INVx2_ASAP7_75t_L g264 ( .A(n_185), .Y(n_264) );
HB1xp67_ASAP7_75t_L g289 ( .A(n_185), .Y(n_289) );
INVx1_ASAP7_75t_L g302 ( .A(n_185), .Y(n_302) );
INVxp67_ASAP7_75t_L g321 ( .A(n_185), .Y(n_321) );
AND2x4_ASAP7_75t_L g352 ( .A(n_185), .B(n_353), .Y(n_352) );
NAND2xp5_ASAP7_75t_L g191 ( .A(n_192), .B(n_233), .Y(n_191) );
OR2x2_ASAP7_75t_L g192 ( .A(n_193), .B(n_222), .Y(n_192) );
INVx2_ASAP7_75t_L g193 ( .A(n_194), .Y(n_193) );
AND2x2_ASAP7_75t_L g394 ( .A(n_194), .B(n_381), .Y(n_394) );
AND2x2_ASAP7_75t_L g418 ( .A(n_194), .B(n_234), .Y(n_418) );
AND2x2_ASAP7_75t_L g194 ( .A(n_195), .B(n_207), .Y(n_194) );
INVx2_ASAP7_75t_L g246 ( .A(n_195), .Y(n_246) );
HB1xp67_ASAP7_75t_L g261 ( .A(n_195), .Y(n_261) );
INVx1_ASAP7_75t_L g318 ( .A(n_195), .Y(n_318) );
AND2x4_ASAP7_75t_L g327 ( .A(n_195), .B(n_245), .Y(n_327) );
AND2x2_ASAP7_75t_L g383 ( .A(n_195), .B(n_235), .Y(n_383) );
AND2x2_ASAP7_75t_L g195 ( .A(n_196), .B(n_202), .Y(n_195) );
NOR3xp33_ASAP7_75t_L g197 ( .A(n_198), .B(n_199), .C(n_200), .Y(n_197) );
AOI21xp5_ASAP7_75t_L g237 ( .A1(n_201), .A2(n_238), .B(n_242), .Y(n_237) );
AOI21xp5_ASAP7_75t_L g546 ( .A1(n_201), .A2(n_547), .B(n_548), .Y(n_546) );
NOR2xp33_ASAP7_75t_L g579 ( .A(n_201), .B(n_580), .Y(n_579) );
NOR2xp33_ASAP7_75t_L g581 ( .A(n_201), .B(n_582), .Y(n_581) );
NOR2xp33_ASAP7_75t_L g584 ( .A(n_201), .B(n_585), .Y(n_584) );
NOR3xp33_ASAP7_75t_L g586 ( .A(n_201), .B(n_213), .C(n_587), .Y(n_586) );
INVx3_ASAP7_75t_L g245 ( .A(n_207), .Y(n_245) );
AND2x2_ASAP7_75t_L g257 ( .A(n_207), .B(n_224), .Y(n_257) );
INVx2_ASAP7_75t_L g296 ( .A(n_207), .Y(n_296) );
NOR2x1_ASAP7_75t_SL g309 ( .A(n_207), .B(n_235), .Y(n_309) );
AND2x4_ASAP7_75t_L g207 ( .A(n_208), .B(n_209), .Y(n_207) );
OAI21xp5_ASAP7_75t_L g209 ( .A1(n_210), .A2(n_214), .B(n_221), .Y(n_209) );
NOR2xp33_ASAP7_75t_L g269 ( .A(n_213), .B(n_270), .Y(n_269) );
OAI22xp5_ASAP7_75t_L g214 ( .A1(n_215), .A2(n_216), .B1(n_218), .B2(n_219), .Y(n_214) );
INVxp67_ASAP7_75t_L g216 ( .A(n_217), .Y(n_216) );
INVxp67_ASAP7_75t_L g219 ( .A(n_220), .Y(n_219) );
INVx1_ASAP7_75t_L g411 ( .A(n_222), .Y(n_411) );
HB1xp67_ASAP7_75t_L g222 ( .A(n_223), .Y(n_222) );
INVx2_ASAP7_75t_L g334 ( .A(n_223), .Y(n_334) );
INVx2_ASAP7_75t_L g223 ( .A(n_224), .Y(n_223) );
HB1xp67_ASAP7_75t_L g292 ( .A(n_224), .Y(n_292) );
HB1xp67_ASAP7_75t_L g308 ( .A(n_224), .Y(n_308) );
AND2x2_ASAP7_75t_L g316 ( .A(n_224), .B(n_245), .Y(n_316) );
INVx1_ASAP7_75t_L g356 ( .A(n_224), .Y(n_356) );
INVx1_ASAP7_75t_L g381 ( .A(n_224), .Y(n_381) );
OR2x2_ASAP7_75t_L g442 ( .A(n_224), .B(n_235), .Y(n_442) );
AO21x2_ASAP7_75t_L g224 ( .A1(n_225), .A2(n_226), .B(n_232), .Y(n_224) );
AO21x2_ASAP7_75t_L g553 ( .A1(n_225), .A2(n_554), .B(n_560), .Y(n_553) );
AO21x2_ASAP7_75t_L g562 ( .A1(n_225), .A2(n_563), .B(n_569), .Y(n_562) );
AO21x2_ASAP7_75t_L g607 ( .A1(n_225), .A2(n_563), .B(n_569), .Y(n_607) );
NAND2xp5_ASAP7_75t_L g226 ( .A(n_227), .B(n_228), .Y(n_226) );
OA211x2_ASAP7_75t_L g463 ( .A1(n_233), .A2(n_464), .B(n_466), .C(n_473), .Y(n_463) );
OR2x6_ASAP7_75t_L g233 ( .A(n_234), .B(n_243), .Y(n_233) );
AND2x2_ASAP7_75t_L g384 ( .A(n_234), .B(n_257), .Y(n_384) );
AND2x2_ASAP7_75t_SL g402 ( .A(n_234), .B(n_244), .Y(n_402) );
BUFx6f_ASAP7_75t_L g234 ( .A(n_235), .Y(n_234) );
INVx4_ASAP7_75t_L g256 ( .A(n_235), .Y(n_256) );
INVx2_ASAP7_75t_L g298 ( .A(n_235), .Y(n_298) );
AND2x4_ASAP7_75t_L g361 ( .A(n_235), .B(n_318), .Y(n_361) );
NAND2xp5_ASAP7_75t_SL g412 ( .A(n_235), .B(n_357), .Y(n_412) );
AND2x2_ASAP7_75t_L g455 ( .A(n_235), .B(n_296), .Y(n_455) );
OR2x6_ASAP7_75t_L g235 ( .A(n_236), .B(n_237), .Y(n_235) );
INVx2_ASAP7_75t_L g243 ( .A(n_244), .Y(n_243) );
NAND2xp5_ASAP7_75t_L g449 ( .A(n_244), .B(n_356), .Y(n_449) );
AND2x2_ASAP7_75t_L g469 ( .A(n_244), .B(n_292), .Y(n_469) );
AND2x2_ASAP7_75t_L g244 ( .A(n_245), .B(n_246), .Y(n_244) );
INVx1_ASAP7_75t_L g357 ( .A(n_245), .Y(n_357) );
INVx1_ASAP7_75t_L g331 ( .A(n_246), .Y(n_331) );
NOR2xp67_ASAP7_75t_SL g247 ( .A(n_248), .B(n_251), .Y(n_247) );
INVx1_ASAP7_75t_L g425 ( .A(n_248), .Y(n_425) );
NOR2xp67_ASAP7_75t_L g472 ( .A(n_248), .B(n_426), .Y(n_472) );
INVx3_ASAP7_75t_L g248 ( .A(n_249), .Y(n_248) );
BUFx3_ASAP7_75t_L g249 ( .A(n_250), .Y(n_249) );
AND2x2_ASAP7_75t_L g445 ( .A(n_250), .B(n_287), .Y(n_445) );
OAI211xp5_ASAP7_75t_L g433 ( .A1(n_251), .A2(n_434), .B(n_437), .C(n_446), .Y(n_433) );
A2O1A1Ixp33_ASAP7_75t_L g477 ( .A1(n_251), .A2(n_471), .B(n_478), .C(n_482), .Y(n_477) );
INVx1_ASAP7_75t_L g251 ( .A(n_252), .Y(n_251) );
AND2x2_ASAP7_75t_L g362 ( .A(n_252), .B(n_363), .Y(n_362) );
AND2x2_ASAP7_75t_L g252 ( .A(n_253), .B(n_254), .Y(n_252) );
INVx2_ASAP7_75t_L g281 ( .A(n_253), .Y(n_281) );
NOR2x1_ASAP7_75t_L g301 ( .A(n_253), .B(n_302), .Y(n_301) );
AND2x2_ASAP7_75t_L g337 ( .A(n_253), .B(n_287), .Y(n_337) );
NOR2xp67_ASAP7_75t_L g447 ( .A(n_253), .B(n_287), .Y(n_447) );
AND2x2_ASAP7_75t_L g320 ( .A(n_254), .B(n_321), .Y(n_320) );
INVx1_ASAP7_75t_L g371 ( .A(n_254), .Y(n_371) );
AND2x2_ASAP7_75t_L g255 ( .A(n_256), .B(n_257), .Y(n_255) );
AND2x4_ASAP7_75t_SL g260 ( .A(n_256), .B(n_261), .Y(n_260) );
AND2x4_ASAP7_75t_L g317 ( .A(n_256), .B(n_318), .Y(n_317) );
NOR2x1_ASAP7_75t_L g346 ( .A(n_256), .B(n_347), .Y(n_346) );
OR2x2_ASAP7_75t_L g365 ( .A(n_256), .B(n_366), .Y(n_365) );
NOR2xp67_ASAP7_75t_SL g448 ( .A(n_256), .B(n_449), .Y(n_448) );
AND2x2_ASAP7_75t_SL g259 ( .A(n_257), .B(n_260), .Y(n_259) );
AND2x2_ASAP7_75t_SL g488 ( .A(n_257), .B(n_330), .Y(n_488) );
NAND2xp5_ASAP7_75t_L g258 ( .A(n_259), .B(n_262), .Y(n_258) );
INVx2_ASAP7_75t_SL g456 ( .A(n_262), .Y(n_456) );
AND2x2_ASAP7_75t_L g262 ( .A(n_263), .B(n_280), .Y(n_262) );
INVx3_ASAP7_75t_L g379 ( .A(n_263), .Y(n_379) );
AND2x2_ASAP7_75t_L g400 ( .A(n_263), .B(n_391), .Y(n_400) );
AND2x2_ASAP7_75t_L g458 ( .A(n_263), .B(n_340), .Y(n_458) );
AND2x4_ASAP7_75t_L g263 ( .A(n_264), .B(n_265), .Y(n_263) );
INVx2_ASAP7_75t_L g287 ( .A(n_265), .Y(n_287) );
INVx1_ASAP7_75t_L g323 ( .A(n_265), .Y(n_323) );
INVx1_ASAP7_75t_L g343 ( .A(n_265), .Y(n_343) );
OR2x2_ASAP7_75t_L g265 ( .A(n_266), .B(n_273), .Y(n_265) );
OAI22xp5_ASAP7_75t_L g273 ( .A1(n_274), .A2(n_277), .B1(n_278), .B2(n_279), .Y(n_273) );
INVx1_ASAP7_75t_L g275 ( .A(n_276), .Y(n_275) );
INVxp67_ASAP7_75t_L g426 ( .A(n_280), .Y(n_426) );
AND2x4_ASAP7_75t_L g280 ( .A(n_281), .B(n_282), .Y(n_280) );
AND2x2_ASAP7_75t_L g286 ( .A(n_282), .B(n_287), .Y(n_286) );
INVx2_ASAP7_75t_L g353 ( .A(n_282), .Y(n_353) );
OAI22xp5_ASAP7_75t_L g283 ( .A1(n_284), .A2(n_290), .B1(n_293), .B2(n_299), .Y(n_283) );
INVx1_ASAP7_75t_L g284 ( .A(n_285), .Y(n_284) );
AND2x4_ASAP7_75t_L g285 ( .A(n_286), .B(n_288), .Y(n_285) );
AND2x2_ASAP7_75t_L g300 ( .A(n_286), .B(n_301), .Y(n_300) );
INVx1_ASAP7_75t_L g311 ( .A(n_286), .Y(n_311) );
INVx1_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
AND2x2_ASAP7_75t_L g360 ( .A(n_291), .B(n_361), .Y(n_360) );
BUFx2_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
INVxp67_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
HB1xp67_ASAP7_75t_L g294 ( .A(n_295), .Y(n_294) );
AND2x2_ASAP7_75t_L g380 ( .A(n_295), .B(n_381), .Y(n_380) );
NOR2x1_ASAP7_75t_L g295 ( .A(n_296), .B(n_297), .Y(n_295) );
INVx1_ASAP7_75t_L g388 ( .A(n_296), .Y(n_388) );
INVx1_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
AND2x2_ASAP7_75t_L g436 ( .A(n_298), .B(n_327), .Y(n_436) );
INVx1_ASAP7_75t_SL g299 ( .A(n_300), .Y(n_299) );
OAI21xp5_ASAP7_75t_L g393 ( .A1(n_300), .A2(n_394), .B(n_395), .Y(n_393) );
OAI21xp5_ASAP7_75t_L g303 ( .A1(n_304), .A2(n_310), .B(n_313), .Y(n_303) );
INVx1_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
AND2x2_ASAP7_75t_L g305 ( .A(n_306), .B(n_309), .Y(n_305) );
INVx1_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
INVx1_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
AND2x2_ASAP7_75t_L g359 ( .A(n_309), .B(n_333), .Y(n_359) );
OAI22xp5_ASAP7_75t_L g416 ( .A1(n_310), .A2(n_417), .B1(n_419), .B2(n_421), .Y(n_416) );
OR2x2_ASAP7_75t_L g310 ( .A(n_311), .B(n_312), .Y(n_310) );
NAND2xp5_ASAP7_75t_L g313 ( .A(n_314), .B(n_319), .Y(n_313) );
INVxp67_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
NAND2xp5_ASAP7_75t_L g315 ( .A(n_316), .B(n_317), .Y(n_315) );
INVx1_ASAP7_75t_SL g366 ( .A(n_316), .Y(n_366) );
AND2x2_ASAP7_75t_L g395 ( .A(n_317), .B(n_333), .Y(n_395) );
NAND2xp5_ASAP7_75t_L g427 ( .A(n_317), .B(n_355), .Y(n_427) );
AND2x2_ASAP7_75t_L g431 ( .A(n_317), .B(n_388), .Y(n_431) );
OAI21xp5_ASAP7_75t_SL g375 ( .A1(n_319), .A2(n_376), .B(n_380), .Y(n_375) );
AND2x2_ASAP7_75t_L g319 ( .A(n_320), .B(n_322), .Y(n_319) );
AND2x2_ASAP7_75t_L g336 ( .A(n_320), .B(n_337), .Y(n_336) );
NAND2x1p5_ASAP7_75t_L g413 ( .A(n_320), .B(n_414), .Y(n_413) );
BUFx2_ASAP7_75t_L g322 ( .A(n_323), .Y(n_322) );
INVx1_ASAP7_75t_SL g405 ( .A(n_323), .Y(n_405) );
NOR2x1_ASAP7_75t_L g324 ( .A(n_325), .B(n_348), .Y(n_324) );
OAI22xp5_ASAP7_75t_L g325 ( .A1(n_326), .A2(n_335), .B1(n_338), .B2(n_344), .Y(n_325) );
NOR2xp33_ASAP7_75t_L g326 ( .A(n_327), .B(n_328), .Y(n_326) );
INVx4_ASAP7_75t_L g347 ( .A(n_327), .Y(n_347) );
NAND2xp5_ASAP7_75t_L g349 ( .A(n_327), .B(n_333), .Y(n_349) );
NAND2xp5_ASAP7_75t_L g479 ( .A(n_327), .B(n_480), .Y(n_479) );
INVxp67_ASAP7_75t_SL g328 ( .A(n_329), .Y(n_328) );
NAND2xp5_ASAP7_75t_L g329 ( .A(n_330), .B(n_332), .Y(n_329) );
AOI21xp5_ASAP7_75t_L g417 ( .A1(n_330), .A2(n_354), .B(n_418), .Y(n_417) );
AND2x4_ASAP7_75t_L g453 ( .A(n_330), .B(n_355), .Y(n_453) );
INVx2_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
AND2x2_ASAP7_75t_L g435 ( .A(n_332), .B(n_436), .Y(n_435) );
INVx1_ASAP7_75t_L g332 ( .A(n_333), .Y(n_332) );
AND2x2_ASAP7_75t_L g471 ( .A(n_333), .B(n_455), .Y(n_471) );
INVx3_ASAP7_75t_L g333 ( .A(n_334), .Y(n_333) );
INVx1_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
AND2x2_ASAP7_75t_L g351 ( .A(n_337), .B(n_352), .Y(n_351) );
NAND2x1p5_ASAP7_75t_L g370 ( .A(n_337), .B(n_371), .Y(n_370) );
OAI22xp5_ASAP7_75t_SL g348 ( .A1(n_338), .A2(n_349), .B1(n_350), .B2(n_354), .Y(n_348) );
INVx1_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
AND2x2_ASAP7_75t_L g339 ( .A(n_340), .B(n_341), .Y(n_339) );
INVx1_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
AND2x2_ASAP7_75t_L g465 ( .A(n_342), .B(n_352), .Y(n_465) );
INVx2_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
INVx1_ASAP7_75t_L g363 ( .A(n_343), .Y(n_363) );
AND2x2_ASAP7_75t_L g389 ( .A(n_343), .B(n_352), .Y(n_389) );
INVxp67_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
NAND2xp5_ASAP7_75t_L g485 ( .A(n_345), .B(n_486), .Y(n_485) );
BUFx2_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
NAND2xp5_ASAP7_75t_L g407 ( .A(n_346), .B(n_408), .Y(n_407) );
INVx2_ASAP7_75t_L g440 ( .A(n_347), .Y(n_440) );
INVx1_ASAP7_75t_L g452 ( .A(n_349), .Y(n_452) );
INVx1_ASAP7_75t_SL g350 ( .A(n_351), .Y(n_350) );
AOI22xp33_ASAP7_75t_L g473 ( .A1(n_351), .A2(n_395), .B1(n_474), .B2(n_475), .Y(n_473) );
AND2x2_ASAP7_75t_L g390 ( .A(n_352), .B(n_391), .Y(n_390) );
AND2x2_ASAP7_75t_L g461 ( .A(n_352), .B(n_414), .Y(n_461) );
INVx1_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
AOI211xp5_ASAP7_75t_SL g364 ( .A1(n_355), .A2(n_365), .B(n_367), .C(n_368), .Y(n_364) );
AND2x2_ASAP7_75t_SL g474 ( .A(n_355), .B(n_361), .Y(n_474) );
AND2x4_ASAP7_75t_SL g355 ( .A(n_356), .B(n_357), .Y(n_355) );
HB1xp67_ASAP7_75t_L g408 ( .A(n_356), .Y(n_408) );
O2A1O1Ixp5_ASAP7_75t_L g358 ( .A1(n_359), .A2(n_360), .B(n_362), .C(n_364), .Y(n_358) );
AOI22xp5_ASAP7_75t_L g386 ( .A1(n_359), .A2(n_387), .B1(n_389), .B2(n_390), .Y(n_386) );
INVx2_ASAP7_75t_L g367 ( .A(n_361), .Y(n_367) );
AND2x2_ASAP7_75t_L g387 ( .A(n_361), .B(n_388), .Y(n_387) );
HB1xp67_ASAP7_75t_L g454 ( .A(n_361), .Y(n_454) );
INVx1_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
INVx1_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
INVxp67_ASAP7_75t_L g495 ( .A(n_373), .Y(n_495) );
NAND4xp75_ASAP7_75t_L g798 ( .A(n_373), .B(n_799), .C(n_800), .D(n_801), .Y(n_798) );
NOR2x1_ASAP7_75t_SL g373 ( .A(n_374), .B(n_385), .Y(n_373) );
NAND2xp5_ASAP7_75t_L g374 ( .A(n_375), .B(n_382), .Y(n_374) );
OAI21xp5_ASAP7_75t_L g382 ( .A1(n_376), .A2(n_383), .B(n_384), .Y(n_382) );
INVx1_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
OR2x2_ASAP7_75t_L g377 ( .A(n_378), .B(n_379), .Y(n_377) );
INVx1_ASAP7_75t_L g406 ( .A(n_378), .Y(n_406) );
INVx1_ASAP7_75t_L g482 ( .A(n_379), .Y(n_482) );
AND2x2_ASAP7_75t_L g420 ( .A(n_383), .B(n_408), .Y(n_420) );
NAND2xp5_ASAP7_75t_L g489 ( .A(n_384), .B(n_490), .Y(n_489) );
NAND2xp5_ASAP7_75t_SL g385 ( .A(n_386), .B(n_393), .Y(n_385) );
AND2x2_ASAP7_75t_L g487 ( .A(n_389), .B(n_488), .Y(n_487) );
INVx1_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
INVx1_ASAP7_75t_L g799 ( .A(n_396), .Y(n_799) );
NAND2x1_ASAP7_75t_L g396 ( .A(n_397), .B(n_432), .Y(n_396) );
NOR3xp33_ASAP7_75t_L g397 ( .A(n_398), .B(n_416), .C(n_423), .Y(n_397) );
OAI222xp33_ASAP7_75t_L g398 ( .A1(n_399), .A2(n_401), .B1(n_403), .B2(n_407), .C1(n_409), .C2(n_413), .Y(n_398) );
INVxp67_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
INVx1_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
INVx1_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
AND2x2_ASAP7_75t_L g404 ( .A(n_405), .B(n_406), .Y(n_404) );
INVx1_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
NOR2x1_ASAP7_75t_L g410 ( .A(n_411), .B(n_412), .Y(n_410) );
INVx2_ASAP7_75t_SL g414 ( .A(n_415), .Y(n_414) );
INVx1_ASAP7_75t_L g459 ( .A(n_418), .Y(n_459) );
INVx1_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
INVx1_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
OAI22xp33_ASAP7_75t_L g423 ( .A1(n_424), .A2(n_427), .B1(n_428), .B2(n_430), .Y(n_423) );
NAND2xp5_ASAP7_75t_L g424 ( .A(n_425), .B(n_426), .Y(n_424) );
INVx1_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
NOR2xp67_ASAP7_75t_SL g432 ( .A(n_433), .B(n_450), .Y(n_432) );
INVx2_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
NAND2xp5_ASAP7_75t_L g437 ( .A(n_438), .B(n_443), .Y(n_437) );
INVx1_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
NAND2x1_ASAP7_75t_L g439 ( .A(n_440), .B(n_441), .Y(n_439) );
NAND2xp5_ASAP7_75t_L g460 ( .A(n_440), .B(n_461), .Y(n_460) );
INVx2_ASAP7_75t_SL g441 ( .A(n_442), .Y(n_441) );
INVx1_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
INVx2_ASAP7_75t_L g492 ( .A(n_445), .Y(n_492) );
NAND2xp33_ASAP7_75t_SL g446 ( .A(n_447), .B(n_448), .Y(n_446) );
OAI221xp5_ASAP7_75t_L g450 ( .A1(n_451), .A2(n_456), .B1(n_457), .B2(n_459), .C(n_460), .Y(n_450) );
NOR4xp25_ASAP7_75t_L g451 ( .A(n_452), .B(n_453), .C(n_454), .D(n_455), .Y(n_451) );
INVx2_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
OAI21xp5_ASAP7_75t_L g494 ( .A1(n_462), .A2(n_495), .B(n_496), .Y(n_494) );
INVx2_ASAP7_75t_L g800 ( .A(n_462), .Y(n_800) );
NAND4xp75_ASAP7_75t_L g462 ( .A(n_463), .B(n_477), .C(n_483), .D(n_489), .Y(n_462) );
INVx3_ASAP7_75t_L g464 ( .A(n_465), .Y(n_464) );
NAND2xp5_ASAP7_75t_SL g466 ( .A(n_467), .B(n_472), .Y(n_466) );
NAND2xp5_ASAP7_75t_L g467 ( .A(n_468), .B(n_470), .Y(n_467) );
INVx2_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
INVx1_ASAP7_75t_L g470 ( .A(n_471), .Y(n_470) );
INVx1_ASAP7_75t_SL g475 ( .A(n_476), .Y(n_475) );
INVxp67_ASAP7_75t_SL g478 ( .A(n_479), .Y(n_478) );
INVx1_ASAP7_75t_L g480 ( .A(n_481), .Y(n_480) );
NOR2x1_ASAP7_75t_L g483 ( .A(n_484), .B(n_487), .Y(n_483) );
INVx1_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
INVx1_ASAP7_75t_L g490 ( .A(n_491), .Y(n_490) );
NAND2xp5_ASAP7_75t_L g493 ( .A(n_494), .B(n_497), .Y(n_493) );
CKINVDCx20_ASAP7_75t_R g498 ( .A(n_499), .Y(n_498) );
NAND2x1_ASAP7_75t_SL g784 ( .A(n_499), .B(n_501), .Y(n_784) );
CKINVDCx11_ASAP7_75t_R g499 ( .A(n_500), .Y(n_499) );
INVx3_ASAP7_75t_SL g501 ( .A(n_502), .Y(n_501) );
AND2x4_ASAP7_75t_L g502 ( .A(n_503), .B(n_672), .Y(n_502) );
NOR3xp33_ASAP7_75t_L g503 ( .A(n_504), .B(n_600), .C(n_650), .Y(n_503) );
OAI211xp5_ASAP7_75t_SL g504 ( .A1(n_505), .A2(n_535), .B(n_570), .C(n_589), .Y(n_504) );
OR2x2_ASAP7_75t_L g505 ( .A(n_506), .B(n_517), .Y(n_505) );
AND2x2_ASAP7_75t_L g599 ( .A(n_506), .B(n_518), .Y(n_599) );
INVx1_ASAP7_75t_L g730 ( .A(n_506), .Y(n_730) );
NOR2x1p5_ASAP7_75t_L g762 ( .A(n_506), .B(n_763), .Y(n_762) );
INVx2_ASAP7_75t_L g506 ( .A(n_507), .Y(n_506) );
AND2x2_ASAP7_75t_L g575 ( .A(n_507), .B(n_576), .Y(n_575) );
INVx2_ASAP7_75t_L g621 ( .A(n_507), .Y(n_621) );
OR2x2_ASAP7_75t_L g625 ( .A(n_507), .B(n_626), .Y(n_625) );
NAND2xp5_ASAP7_75t_L g637 ( .A(n_507), .B(n_520), .Y(n_637) );
OR2x2_ASAP7_75t_L g659 ( .A(n_507), .B(n_520), .Y(n_659) );
AND2x4_ASAP7_75t_L g665 ( .A(n_507), .B(n_629), .Y(n_665) );
OR2x2_ASAP7_75t_L g682 ( .A(n_507), .B(n_577), .Y(n_682) );
INVx1_ASAP7_75t_L g717 ( .A(n_507), .Y(n_717) );
HB1xp67_ASAP7_75t_L g739 ( .A(n_507), .Y(n_739) );
OR2x2_ASAP7_75t_L g753 ( .A(n_507), .B(n_686), .Y(n_753) );
AND2x4_ASAP7_75t_SL g757 ( .A(n_507), .B(n_577), .Y(n_757) );
OR2x6_ASAP7_75t_L g507 ( .A(n_508), .B(n_516), .Y(n_507) );
INVx1_ASAP7_75t_L g517 ( .A(n_518), .Y(n_517) );
AND2x2_ASAP7_75t_L g709 ( .A(n_518), .B(n_665), .Y(n_709) );
AND2x2_ASAP7_75t_L g756 ( .A(n_518), .B(n_757), .Y(n_756) );
AND2x2_ASAP7_75t_L g518 ( .A(n_519), .B(n_526), .Y(n_518) );
INVx2_ASAP7_75t_L g519 ( .A(n_520), .Y(n_519) );
INVx1_ASAP7_75t_L g574 ( .A(n_520), .Y(n_574) );
AND2x2_ASAP7_75t_L g619 ( .A(n_520), .B(n_526), .Y(n_619) );
INVx2_ASAP7_75t_L g626 ( .A(n_520), .Y(n_626) );
HB1xp67_ASAP7_75t_L g747 ( .A(n_520), .Y(n_747) );
BUFx3_ASAP7_75t_L g763 ( .A(n_520), .Y(n_763) );
INVx2_ASAP7_75t_L g588 ( .A(n_526), .Y(n_588) );
NAND2xp5_ASAP7_75t_L g628 ( .A(n_526), .B(n_629), .Y(n_628) );
OR2x2_ASAP7_75t_L g686 ( .A(n_526), .B(n_626), .Y(n_686) );
INVx1_ASAP7_75t_L g704 ( .A(n_526), .Y(n_704) );
HB1xp67_ASAP7_75t_L g720 ( .A(n_526), .Y(n_720) );
INVx1_ASAP7_75t_L g742 ( .A(n_526), .Y(n_742) );
NAND2xp5_ASAP7_75t_L g769 ( .A(n_526), .B(n_621), .Y(n_769) );
NAND2xp5_ASAP7_75t_L g779 ( .A(n_526), .B(n_577), .Y(n_779) );
INVx3_ASAP7_75t_L g526 ( .A(n_527), .Y(n_526) );
NAND2xp5_ASAP7_75t_L g528 ( .A(n_529), .B(n_533), .Y(n_528) );
INVx1_ASAP7_75t_SL g535 ( .A(n_536), .Y(n_535) );
AND2x2_ASAP7_75t_L g536 ( .A(n_537), .B(n_543), .Y(n_536) );
AND2x4_ASAP7_75t_L g593 ( .A(n_537), .B(n_594), .Y(n_593) );
INVx2_ASAP7_75t_L g604 ( .A(n_537), .Y(n_604) );
AND2x2_ASAP7_75t_L g609 ( .A(n_537), .B(n_610), .Y(n_609) );
AND2x2_ASAP7_75t_L g644 ( .A(n_537), .B(n_552), .Y(n_644) );
AND2x2_ASAP7_75t_L g654 ( .A(n_537), .B(n_553), .Y(n_654) );
OR2x2_ASAP7_75t_L g734 ( .A(n_537), .B(n_649), .Y(n_734) );
OAI322xp33_ASAP7_75t_L g764 ( .A1(n_537), .A2(n_677), .A3(n_716), .B1(n_749), .B2(n_765), .C1(n_766), .C2(n_767), .Y(n_764) );
OR2x2_ASAP7_75t_L g765 ( .A(n_537), .B(n_747), .Y(n_765) );
BUFx6f_ASAP7_75t_L g537 ( .A(n_538), .Y(n_537) );
INVx2_ASAP7_75t_L g598 ( .A(n_538), .Y(n_598) );
NAND2xp5_ASAP7_75t_L g539 ( .A(n_540), .B(n_541), .Y(n_539) );
AOI22xp5_ASAP7_75t_L g710 ( .A1(n_543), .A2(n_711), .B1(n_715), .B2(n_718), .Y(n_710) );
AOI211xp5_ASAP7_75t_L g770 ( .A1(n_543), .A2(n_771), .B(n_772), .C(n_775), .Y(n_770) );
AND2x4_ASAP7_75t_SL g543 ( .A(n_544), .B(n_552), .Y(n_543) );
AND2x4_ASAP7_75t_L g592 ( .A(n_544), .B(n_562), .Y(n_592) );
HB1xp67_ASAP7_75t_L g596 ( .A(n_544), .Y(n_596) );
INVx5_ASAP7_75t_L g608 ( .A(n_544), .Y(n_608) );
INVx2_ASAP7_75t_L g617 ( .A(n_544), .Y(n_617) );
AND2x2_ASAP7_75t_L g640 ( .A(n_544), .B(n_553), .Y(n_640) );
AND2x2_ASAP7_75t_L g669 ( .A(n_544), .B(n_561), .Y(n_669) );
OR2x2_ASAP7_75t_L g678 ( .A(n_544), .B(n_598), .Y(n_678) );
OR2x2_ASAP7_75t_L g693 ( .A(n_544), .B(n_607), .Y(n_693) );
OR2x6_ASAP7_75t_L g544 ( .A(n_545), .B(n_546), .Y(n_544) );
NAND2xp5_ASAP7_75t_L g570 ( .A(n_552), .B(n_571), .Y(n_570) );
INVx3_ASAP7_75t_SL g677 ( .A(n_552), .Y(n_677) );
AND2x2_ASAP7_75t_L g700 ( .A(n_552), .B(n_608), .Y(n_700) );
AND2x4_ASAP7_75t_L g552 ( .A(n_553), .B(n_561), .Y(n_552) );
INVx2_ASAP7_75t_L g594 ( .A(n_553), .Y(n_594) );
AND2x2_ASAP7_75t_L g597 ( .A(n_553), .B(n_598), .Y(n_597) );
OR2x2_ASAP7_75t_L g611 ( .A(n_553), .B(n_562), .Y(n_611) );
INVx1_ASAP7_75t_L g615 ( .A(n_553), .Y(n_615) );
NAND2xp5_ASAP7_75t_L g649 ( .A(n_553), .B(n_562), .Y(n_649) );
HB1xp67_ASAP7_75t_L g713 ( .A(n_553), .Y(n_713) );
NAND2xp5_ASAP7_75t_L g724 ( .A(n_553), .B(n_608), .Y(n_724) );
NAND2xp5_ASAP7_75t_L g554 ( .A(n_555), .B(n_559), .Y(n_554) );
INVx2_ASAP7_75t_L g561 ( .A(n_562), .Y(n_561) );
HB1xp67_ASAP7_75t_L g630 ( .A(n_562), .Y(n_630) );
AND2x2_ASAP7_75t_L g714 ( .A(n_562), .B(n_598), .Y(n_714) );
NAND2xp5_ASAP7_75t_L g563 ( .A(n_564), .B(n_568), .Y(n_563) );
AND2x2_ASAP7_75t_L g571 ( .A(n_572), .B(n_575), .Y(n_571) );
NAND2xp5_ASAP7_75t_L g680 ( .A(n_572), .B(n_681), .Y(n_680) );
INVx1_ASAP7_75t_L g572 ( .A(n_573), .Y(n_572) );
OR2x6_ASAP7_75t_SL g778 ( .A(n_573), .B(n_779), .Y(n_778) );
INVxp67_ASAP7_75t_SL g573 ( .A(n_574), .Y(n_573) );
HB1xp67_ASAP7_75t_L g664 ( .A(n_574), .Y(n_664) );
NAND2xp5_ASAP7_75t_L g703 ( .A(n_574), .B(n_704), .Y(n_703) );
INVx1_ASAP7_75t_L g726 ( .A(n_574), .Y(n_726) );
AOI22xp5_ASAP7_75t_L g634 ( .A1(n_575), .A2(n_635), .B1(n_638), .B2(n_645), .Y(n_634) );
NAND2xp5_ASAP7_75t_L g657 ( .A(n_576), .B(n_658), .Y(n_657) );
AND2x2_ASAP7_75t_L g670 ( .A(n_576), .B(n_671), .Y(n_670) );
NAND2xp5_ASAP7_75t_L g716 ( .A(n_576), .B(n_717), .Y(n_716) );
AND2x2_ASAP7_75t_SL g725 ( .A(n_576), .B(n_726), .Y(n_725) );
AND2x4_ASAP7_75t_L g576 ( .A(n_577), .B(n_588), .Y(n_576) );
AND2x2_ASAP7_75t_L g620 ( .A(n_577), .B(n_621), .Y(n_620) );
INVx3_ASAP7_75t_L g629 ( .A(n_577), .Y(n_629) );
OAI22xp33_ASAP7_75t_L g687 ( .A1(n_577), .A2(n_636), .B1(n_688), .B2(n_690), .Y(n_687) );
INVx1_ASAP7_75t_L g695 ( .A(n_577), .Y(n_695) );
NOR2xp33_ASAP7_75t_L g735 ( .A(n_577), .B(n_689), .Y(n_735) );
NAND2xp5_ASAP7_75t_L g750 ( .A(n_577), .B(n_619), .Y(n_750) );
NAND2xp5_ASAP7_75t_L g768 ( .A(n_577), .B(n_626), .Y(n_768) );
AND2x4_ASAP7_75t_L g577 ( .A(n_578), .B(n_583), .Y(n_577) );
OAI21xp33_ASAP7_75t_L g589 ( .A1(n_590), .A2(n_595), .B(n_599), .Y(n_589) );
NOR2xp33_ASAP7_75t_L g590 ( .A(n_591), .B(n_593), .Y(n_590) );
NAND4xp25_ASAP7_75t_SL g638 ( .A(n_591), .B(n_639), .C(n_641), .D(n_643), .Y(n_638) );
INVx2_ASAP7_75t_SL g591 ( .A(n_592), .Y(n_591) );
NAND2xp5_ASAP7_75t_L g728 ( .A(n_592), .B(n_699), .Y(n_728) );
AND2x2_ASAP7_75t_L g755 ( .A(n_592), .B(n_593), .Y(n_755) );
NAND2xp5_ASAP7_75t_L g766 ( .A(n_592), .B(n_615), .Y(n_766) );
INVx1_ASAP7_75t_L g631 ( .A(n_593), .Y(n_631) );
AOI22xp5_ASAP7_75t_L g666 ( .A1(n_593), .A2(n_656), .B1(n_667), .B2(n_670), .Y(n_666) );
NAND3xp33_ASAP7_75t_L g688 ( .A(n_593), .B(n_606), .C(n_689), .Y(n_688) );
NAND2xp5_ASAP7_75t_L g707 ( .A(n_593), .B(n_608), .Y(n_707) );
NAND2xp5_ASAP7_75t_L g759 ( .A(n_593), .B(n_616), .Y(n_759) );
AND2x2_ASAP7_75t_L g691 ( .A(n_594), .B(n_598), .Y(n_691) );
HB1xp67_ASAP7_75t_L g752 ( .A(n_594), .Y(n_752) );
AND2x2_ASAP7_75t_L g595 ( .A(n_596), .B(n_597), .Y(n_595) );
INVx1_ASAP7_75t_L g647 ( .A(n_596), .Y(n_647) );
INVx1_ASAP7_75t_L g737 ( .A(n_597), .Y(n_737) );
AND2x2_ASAP7_75t_L g744 ( .A(n_597), .B(n_608), .Y(n_744) );
BUFx2_ASAP7_75t_L g699 ( .A(n_598), .Y(n_699) );
NAND3xp33_ASAP7_75t_SL g600 ( .A(n_601), .B(n_622), .C(n_634), .Y(n_600) );
OAI31xp33_ASAP7_75t_L g601 ( .A1(n_602), .A2(n_609), .A3(n_612), .B(n_618), .Y(n_601) );
AOI22xp5_ASAP7_75t_L g655 ( .A1(n_602), .A2(n_656), .B1(n_660), .B2(n_661), .Y(n_655) );
INVx1_ASAP7_75t_L g602 ( .A(n_603), .Y(n_602) );
OR2x2_ASAP7_75t_L g603 ( .A(n_604), .B(n_605), .Y(n_603) );
OR2x2_ASAP7_75t_L g641 ( .A(n_604), .B(n_642), .Y(n_641) );
NOR2x1_ASAP7_75t_L g667 ( .A(n_604), .B(n_668), .Y(n_667) );
O2A1O1Ixp33_ASAP7_75t_L g736 ( .A1(n_605), .A2(n_707), .B(n_737), .C(n_738), .Y(n_736) );
INVx2_ASAP7_75t_L g605 ( .A(n_606), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g751 ( .A(n_606), .B(n_752), .Y(n_751) );
AND2x4_ASAP7_75t_L g606 ( .A(n_607), .B(n_608), .Y(n_606) );
NAND2xp5_ASAP7_75t_L g642 ( .A(n_607), .B(n_615), .Y(n_642) );
AND2x2_ASAP7_75t_L g660 ( .A(n_607), .B(n_640), .Y(n_660) );
AND2x2_ASAP7_75t_L g777 ( .A(n_610), .B(n_699), .Y(n_777) );
INVx2_ASAP7_75t_L g610 ( .A(n_611), .Y(n_610) );
OR2x2_ASAP7_75t_L g633 ( .A(n_611), .B(n_617), .Y(n_633) );
NOR2xp33_ASAP7_75t_L g612 ( .A(n_613), .B(n_616), .Y(n_612) );
INVx1_ASAP7_75t_L g613 ( .A(n_614), .Y(n_613) );
HB1xp67_ASAP7_75t_L g614 ( .A(n_615), .Y(n_614) );
NAND2xp5_ASAP7_75t_L g653 ( .A(n_616), .B(n_654), .Y(n_653) );
AND2x2_ASAP7_75t_L g708 ( .A(n_616), .B(n_691), .Y(n_708) );
INVx2_ASAP7_75t_L g616 ( .A(n_617), .Y(n_616) );
NAND2xp5_ASAP7_75t_L g697 ( .A(n_617), .B(n_691), .Y(n_697) );
AND2x2_ASAP7_75t_L g618 ( .A(n_619), .B(n_620), .Y(n_618) );
INVx2_ASAP7_75t_L g689 ( .A(n_619), .Y(n_689) );
NAND2xp5_ASAP7_75t_L g719 ( .A(n_620), .B(n_720), .Y(n_719) );
AOI32xp33_ASAP7_75t_L g622 ( .A1(n_623), .A2(n_630), .A3(n_631), .B1(n_632), .B2(n_817), .Y(n_622) );
AOI221xp5_ASAP7_75t_L g743 ( .A1(n_623), .A2(n_708), .B1(n_744), .B2(n_745), .C(n_748), .Y(n_743) );
AND2x4_ASAP7_75t_L g623 ( .A(n_624), .B(n_627), .Y(n_623) );
INVx2_ASAP7_75t_L g624 ( .A(n_625), .Y(n_624) );
HB1xp67_ASAP7_75t_L g671 ( .A(n_626), .Y(n_671) );
INVx1_ASAP7_75t_L g627 ( .A(n_628), .Y(n_627) );
OR2x2_ASAP7_75t_L g636 ( .A(n_628), .B(n_637), .Y(n_636) );
AND2x2_ASAP7_75t_L g741 ( .A(n_629), .B(n_742), .Y(n_741) );
NAND2xp5_ASAP7_75t_SL g651 ( .A(n_630), .B(n_652), .Y(n_651) );
AOI221xp5_ASAP7_75t_L g674 ( .A1(n_632), .A2(n_675), .B1(n_679), .B2(n_683), .C(n_687), .Y(n_674) );
INVx1_ASAP7_75t_L g632 ( .A(n_633), .Y(n_632) );
INVx2_ASAP7_75t_L g635 ( .A(n_636), .Y(n_635) );
OAI211xp5_ASAP7_75t_L g650 ( .A1(n_637), .A2(n_651), .B(n_655), .C(n_666), .Y(n_650) );
INVx1_ASAP7_75t_L g639 ( .A(n_640), .Y(n_639) );
OAI322xp33_ASAP7_75t_L g748 ( .A1(n_643), .A2(n_653), .A3(n_702), .B1(n_749), .B2(n_750), .C1(n_751), .C2(n_753), .Y(n_748) );
INVx2_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
INVx2_ASAP7_75t_L g645 ( .A(n_646), .Y(n_645) );
AOI21xp33_ASAP7_75t_L g775 ( .A1(n_646), .A2(n_776), .B(n_778), .Y(n_775) );
NAND2xp5_ASAP7_75t_SL g646 ( .A(n_647), .B(n_648), .Y(n_646) );
INVx1_ASAP7_75t_L g648 ( .A(n_649), .Y(n_648) );
O2A1O1Ixp33_ASAP7_75t_L g732 ( .A1(n_652), .A2(n_733), .B(n_735), .C(n_736), .Y(n_732) );
INVx1_ASAP7_75t_L g652 ( .A(n_653), .Y(n_652) );
INVx1_ASAP7_75t_L g656 ( .A(n_657), .Y(n_656) );
INVx1_ASAP7_75t_SL g658 ( .A(n_659), .Y(n_658) );
OR2x2_ASAP7_75t_L g774 ( .A(n_659), .B(n_740), .Y(n_774) );
INVx1_ASAP7_75t_L g661 ( .A(n_662), .Y(n_661) );
NAND2xp5_ASAP7_75t_L g662 ( .A(n_663), .B(n_665), .Y(n_662) );
INVxp67_ASAP7_75t_L g663 ( .A(n_664), .Y(n_663) );
NAND2xp5_ASAP7_75t_L g684 ( .A(n_665), .B(n_685), .Y(n_684) );
INVx1_ASAP7_75t_L g749 ( .A(n_665), .Y(n_749) );
INVx2_ASAP7_75t_L g668 ( .A(n_669), .Y(n_668) );
OAI31xp33_ASAP7_75t_L g705 ( .A1(n_669), .A2(n_706), .A3(n_708), .B(n_709), .Y(n_705) );
NOR2x1_ASAP7_75t_L g672 ( .A(n_673), .B(n_731), .Y(n_672) );
NAND5xp2_ASAP7_75t_L g673 ( .A(n_674), .B(n_694), .C(n_705), .D(n_710), .E(n_721), .Y(n_673) );
INVx1_ASAP7_75t_L g675 ( .A(n_676), .Y(n_675) );
OR2x2_ASAP7_75t_L g676 ( .A(n_677), .B(n_678), .Y(n_676) );
AOI21xp33_ASAP7_75t_L g772 ( .A1(n_677), .A2(n_773), .B(n_774), .Y(n_772) );
INVx1_ASAP7_75t_SL g679 ( .A(n_680), .Y(n_679) );
AND2x2_ASAP7_75t_L g745 ( .A(n_681), .B(n_746), .Y(n_745) );
INVx1_ASAP7_75t_SL g681 ( .A(n_682), .Y(n_681) );
INVx1_ASAP7_75t_L g683 ( .A(n_684), .Y(n_683) );
INVx1_ASAP7_75t_L g685 ( .A(n_686), .Y(n_685) );
NAND2xp5_ASAP7_75t_L g690 ( .A(n_691), .B(n_692), .Y(n_690) );
INVx1_ASAP7_75t_SL g692 ( .A(n_693), .Y(n_692) );
A2O1A1Ixp33_ASAP7_75t_L g694 ( .A1(n_695), .A2(n_696), .B(n_698), .C(n_701), .Y(n_694) );
INVxp33_ASAP7_75t_L g696 ( .A(n_697), .Y(n_696) );
AND2x2_ASAP7_75t_L g698 ( .A(n_699), .B(n_700), .Y(n_698) );
OR2x2_ASAP7_75t_L g723 ( .A(n_699), .B(n_724), .Y(n_723) );
HB1xp67_ASAP7_75t_L g701 ( .A(n_702), .Y(n_701) );
NAND2xp5_ASAP7_75t_L g729 ( .A(n_702), .B(n_730), .Y(n_729) );
INVx1_ASAP7_75t_L g702 ( .A(n_703), .Y(n_702) );
INVx1_ASAP7_75t_L g706 ( .A(n_707), .Y(n_706) );
AND2x2_ASAP7_75t_SL g711 ( .A(n_712), .B(n_714), .Y(n_711) );
INVx1_ASAP7_75t_L g712 ( .A(n_713), .Y(n_712) );
INVx1_ASAP7_75t_L g773 ( .A(n_714), .Y(n_773) );
INVx1_ASAP7_75t_SL g715 ( .A(n_716), .Y(n_715) );
INVx1_ASAP7_75t_L g718 ( .A(n_719), .Y(n_718) );
AOI21xp5_ASAP7_75t_L g721 ( .A1(n_722), .A2(n_725), .B(n_727), .Y(n_721) );
INVx1_ASAP7_75t_L g722 ( .A(n_723), .Y(n_722) );
AOI21xp33_ASAP7_75t_L g727 ( .A1(n_723), .A2(n_728), .B(n_729), .Y(n_727) );
NAND4xp25_ASAP7_75t_L g731 ( .A(n_732), .B(n_743), .C(n_754), .D(n_770), .Y(n_731) );
INVx1_ASAP7_75t_SL g733 ( .A(n_734), .Y(n_733) );
OR2x2_ASAP7_75t_L g738 ( .A(n_739), .B(n_740), .Y(n_738) );
INVx1_ASAP7_75t_SL g740 ( .A(n_741), .Y(n_740) );
NAND2xp5_ASAP7_75t_L g761 ( .A(n_741), .B(n_762), .Y(n_761) );
HB1xp67_ASAP7_75t_L g746 ( .A(n_747), .Y(n_746) );
INVx1_ASAP7_75t_L g771 ( .A(n_753), .Y(n_771) );
AOI221xp5_ASAP7_75t_L g754 ( .A1(n_755), .A2(n_756), .B1(n_758), .B2(n_760), .C(n_764), .Y(n_754) );
INVx1_ASAP7_75t_L g758 ( .A(n_759), .Y(n_758) );
INVx1_ASAP7_75t_L g760 ( .A(n_761), .Y(n_760) );
OR2x2_ASAP7_75t_L g767 ( .A(n_768), .B(n_769), .Y(n_767) );
INVx2_ASAP7_75t_L g776 ( .A(n_777), .Y(n_776) );
AOI21xp33_ASAP7_75t_SL g781 ( .A1(n_780), .A2(n_782), .B(n_785), .Y(n_781) );
NOR2xp33_ASAP7_75t_L g785 ( .A(n_786), .B(n_787), .Y(n_785) );
BUFx2_ASAP7_75t_L g787 ( .A(n_788), .Y(n_787) );
INVxp67_ASAP7_75t_L g789 ( .A(n_790), .Y(n_789) );
AOI21xp5_ASAP7_75t_L g790 ( .A1(n_791), .A2(n_794), .B(n_802), .Y(n_790) );
CKINVDCx11_ASAP7_75t_R g791 ( .A(n_792), .Y(n_791) );
CKINVDCx20_ASAP7_75t_R g792 ( .A(n_793), .Y(n_792) );
INVx2_ASAP7_75t_L g794 ( .A(n_795), .Y(n_794) );
XNOR2x1_ASAP7_75t_L g795 ( .A(n_796), .B(n_798), .Y(n_795) );
CKINVDCx20_ASAP7_75t_R g804 ( .A(n_805), .Y(n_804) );
INVx2_ASAP7_75t_L g805 ( .A(n_806), .Y(n_805) );
INVx1_ASAP7_75t_L g806 ( .A(n_807), .Y(n_806) );
INVx1_ASAP7_75t_SL g808 ( .A(n_809), .Y(n_808) );
CKINVDCx11_ASAP7_75t_R g810 ( .A(n_811), .Y(n_810) );
CKINVDCx8_ASAP7_75t_R g811 ( .A(n_812), .Y(n_811) );
INVx2_ASAP7_75t_L g813 ( .A(n_814), .Y(n_813) );
endmodule