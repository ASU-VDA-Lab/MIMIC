module fake_jpeg_31290_n_521 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_521);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_521;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_518;
wire n_378;
wire n_132;
wire n_133;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx2_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_13),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

INVx8_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

BUFx16f_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

INVx13_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_3),
.Y(n_26)
);

BUFx8_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_11),
.Y(n_34)
);

BUFx10_ASAP7_75t_L g35 ( 
.A(n_0),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_3),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_0),
.Y(n_37)
);

INVx11_ASAP7_75t_L g38 ( 
.A(n_9),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_7),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_3),
.Y(n_40)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_5),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_13),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_1),
.Y(n_43)
);

BUFx16f_ASAP7_75t_L g44 ( 
.A(n_9),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_6),
.Y(n_45)
);

BUFx10_ASAP7_75t_L g46 ( 
.A(n_8),
.Y(n_46)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_7),
.Y(n_47)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_2),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_14),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_8),
.Y(n_50)
);

INVx8_ASAP7_75t_L g51 ( 
.A(n_13),
.Y(n_51)
);

BUFx10_ASAP7_75t_L g52 ( 
.A(n_11),
.Y(n_52)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_23),
.Y(n_53)
);

BUFx5_ASAP7_75t_L g129 ( 
.A(n_53),
.Y(n_129)
);

BUFx2_ASAP7_75t_L g54 ( 
.A(n_27),
.Y(n_54)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_54),
.Y(n_112)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_21),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g153 ( 
.A(n_55),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_17),
.B(n_7),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_56),
.B(n_57),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_17),
.B(n_7),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_21),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g159 ( 
.A(n_58),
.Y(n_159)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_16),
.Y(n_59)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_59),
.Y(n_110)
);

INVx5_ASAP7_75t_L g60 ( 
.A(n_22),
.Y(n_60)
);

INVx5_ASAP7_75t_L g144 ( 
.A(n_60),
.Y(n_144)
);

INVx2_ASAP7_75t_SL g61 ( 
.A(n_20),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_61),
.B(n_72),
.Y(n_148)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_47),
.Y(n_62)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_62),
.Y(n_113)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_29),
.Y(n_63)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_63),
.Y(n_130)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_25),
.Y(n_64)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_64),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_21),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g169 ( 
.A(n_65),
.Y(n_169)
);

INVx11_ASAP7_75t_L g66 ( 
.A(n_44),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g172 ( 
.A(n_66),
.Y(n_172)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_29),
.Y(n_67)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_67),
.Y(n_132)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_39),
.Y(n_68)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_68),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_21),
.Y(n_69)
);

INVx6_ASAP7_75t_L g119 ( 
.A(n_69),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_49),
.Y(n_70)
);

INVx6_ASAP7_75t_L g143 ( 
.A(n_70),
.Y(n_143)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_22),
.Y(n_71)
);

INVx4_ASAP7_75t_L g111 ( 
.A(n_71),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_34),
.B(n_9),
.Y(n_72)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_16),
.Y(n_73)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_73),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_49),
.Y(n_74)
);

INVx8_ASAP7_75t_L g149 ( 
.A(n_74),
.Y(n_149)
);

INVx2_ASAP7_75t_SL g75 ( 
.A(n_20),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_75),
.B(n_101),
.Y(n_158)
);

BUFx3_ASAP7_75t_L g76 ( 
.A(n_22),
.Y(n_76)
);

INVx4_ASAP7_75t_L g142 ( 
.A(n_76),
.Y(n_142)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_48),
.Y(n_77)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_77),
.Y(n_120)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_25),
.Y(n_78)
);

INVx3_ASAP7_75t_L g125 ( 
.A(n_78),
.Y(n_125)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_25),
.Y(n_79)
);

INVx3_ASAP7_75t_L g162 ( 
.A(n_79),
.Y(n_162)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_47),
.Y(n_80)
);

INVx3_ASAP7_75t_L g170 ( 
.A(n_80),
.Y(n_170)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_48),
.Y(n_81)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_81),
.Y(n_124)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_47),
.Y(n_82)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_82),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_49),
.Y(n_83)
);

INVx11_ASAP7_75t_L g141 ( 
.A(n_83),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_30),
.Y(n_84)
);

INVx5_ASAP7_75t_L g152 ( 
.A(n_84),
.Y(n_152)
);

BUFx2_ASAP7_75t_L g85 ( 
.A(n_27),
.Y(n_85)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_85),
.Y(n_131)
);

BUFx3_ASAP7_75t_L g86 ( 
.A(n_31),
.Y(n_86)
);

INVx4_ASAP7_75t_L g163 ( 
.A(n_86),
.Y(n_163)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_33),
.Y(n_87)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_87),
.Y(n_138)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_33),
.Y(n_88)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_88),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_30),
.Y(n_89)
);

INVx4_ASAP7_75t_L g109 ( 
.A(n_89),
.Y(n_109)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_31),
.Y(n_90)
);

INVx2_ASAP7_75t_SL g122 ( 
.A(n_90),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_30),
.Y(n_91)
);

INVx4_ASAP7_75t_L g121 ( 
.A(n_91),
.Y(n_121)
);

INVx8_ASAP7_75t_L g92 ( 
.A(n_27),
.Y(n_92)
);

BUFx5_ASAP7_75t_L g136 ( 
.A(n_92),
.Y(n_136)
);

INVx5_ASAP7_75t_L g93 ( 
.A(n_18),
.Y(n_93)
);

INVx4_ASAP7_75t_SL g128 ( 
.A(n_93),
.Y(n_128)
);

BUFx12_ASAP7_75t_L g94 ( 
.A(n_44),
.Y(n_94)
);

INVx1_ASAP7_75t_SL g117 ( 
.A(n_94),
.Y(n_117)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_33),
.Y(n_95)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_95),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_34),
.B(n_15),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_96),
.B(n_42),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_30),
.Y(n_97)
);

INVx4_ASAP7_75t_L g123 ( 
.A(n_97),
.Y(n_123)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_31),
.Y(n_98)
);

INVx4_ASAP7_75t_L g127 ( 
.A(n_98),
.Y(n_127)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_39),
.Y(n_99)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_99),
.Y(n_165)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_32),
.Y(n_100)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_100),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_42),
.B(n_14),
.Y(n_101)
);

BUFx12f_ASAP7_75t_L g102 ( 
.A(n_23),
.Y(n_102)
);

BUFx12f_ASAP7_75t_L g134 ( 
.A(n_102),
.Y(n_134)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_32),
.Y(n_103)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_103),
.Y(n_156)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_32),
.Y(n_104)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_104),
.Y(n_157)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_36),
.Y(n_105)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_105),
.Y(n_161)
);

BUFx12f_ASAP7_75t_L g106 ( 
.A(n_23),
.Y(n_106)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_106),
.Y(n_114)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_36),
.Y(n_107)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_107),
.Y(n_164)
);

BUFx3_ASAP7_75t_L g108 ( 
.A(n_18),
.Y(n_108)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_108),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_133),
.B(n_139),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_56),
.A2(n_41),
.B1(n_24),
.B2(n_26),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_135),
.A2(n_147),
.B1(n_151),
.B2(n_166),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_57),
.B(n_50),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_72),
.B(n_50),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_140),
.B(n_52),
.Y(n_209)
);

NOR2x1_ASAP7_75t_R g145 ( 
.A(n_101),
.B(n_44),
.Y(n_145)
);

AND2x2_ASAP7_75t_L g201 ( 
.A(n_145),
.B(n_27),
.Y(n_201)
);

AOI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_54),
.A2(n_36),
.B1(n_51),
.B2(n_24),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_SL g196 ( 
.A1(n_146),
.A2(n_160),
.B1(n_92),
.B2(n_102),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_70),
.A2(n_74),
.B1(n_83),
.B2(n_65),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_58),
.A2(n_41),
.B1(n_24),
.B2(n_45),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_SL g160 ( 
.A1(n_85),
.A2(n_51),
.B1(n_41),
.B2(n_19),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_L g166 ( 
.A1(n_55),
.A2(n_19),
.B1(n_51),
.B2(n_45),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_84),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_167),
.B(n_91),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_69),
.A2(n_26),
.B1(n_43),
.B2(n_40),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_171),
.A2(n_173),
.B1(n_37),
.B2(n_97),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_L g173 ( 
.A1(n_89),
.A2(n_43),
.B1(n_40),
.B2(n_28),
.Y(n_173)
);

INVx4_ASAP7_75t_SL g174 ( 
.A(n_129),
.Y(n_174)
);

INVx13_ASAP7_75t_L g239 ( 
.A(n_174),
.Y(n_239)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_130),
.Y(n_175)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_175),
.Y(n_229)
);

CKINVDCx14_ASAP7_75t_R g262 ( 
.A(n_176),
.Y(n_262)
);

CKINVDCx14_ASAP7_75t_R g178 ( 
.A(n_148),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_178),
.B(n_189),
.Y(n_230)
);

INVxp67_ASAP7_75t_SL g179 ( 
.A(n_114),
.Y(n_179)
);

INVx11_ASAP7_75t_L g269 ( 
.A(n_179),
.Y(n_269)
);

XOR2xp5_ASAP7_75t_L g180 ( 
.A(n_118),
.B(n_44),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_SL g235 ( 
.A(n_180),
.B(n_201),
.C(n_202),
.Y(n_235)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_132),
.Y(n_181)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_181),
.Y(n_243)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_137),
.Y(n_182)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_182),
.Y(n_258)
);

OAI21xp5_ASAP7_75t_L g183 ( 
.A1(n_148),
.A2(n_75),
.B(n_61),
.Y(n_183)
);

A2O1A1Ixp33_ASAP7_75t_L g240 ( 
.A1(n_183),
.A2(n_134),
.B(n_52),
.C(n_46),
.Y(n_240)
);

BUFx3_ASAP7_75t_L g184 ( 
.A(n_172),
.Y(n_184)
);

BUFx3_ASAP7_75t_L g231 ( 
.A(n_184),
.Y(n_231)
);

INVx4_ASAP7_75t_L g186 ( 
.A(n_172),
.Y(n_186)
);

HB1xp67_ASAP7_75t_L g264 ( 
.A(n_186),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_165),
.A2(n_37),
.B1(n_28),
.B2(n_20),
.Y(n_187)
);

AOI22xp33_ASAP7_75t_SL g256 ( 
.A1(n_187),
.A2(n_196),
.B1(n_218),
.B2(n_219),
.Y(n_256)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_110),
.Y(n_188)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_188),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_158),
.B(n_94),
.Y(n_189)
);

INVx4_ASAP7_75t_L g190 ( 
.A(n_112),
.Y(n_190)
);

INVx3_ASAP7_75t_L g270 ( 
.A(n_190),
.Y(n_270)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_116),
.Y(n_191)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_191),
.Y(n_265)
);

INVx1_ASAP7_75t_SL g192 ( 
.A(n_131),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_192),
.B(n_194),
.Y(n_233)
);

BUFx2_ASAP7_75t_L g193 ( 
.A(n_168),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_193),
.Y(n_238)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_126),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_158),
.B(n_106),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_195),
.B(n_197),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_118),
.B(n_53),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g250 ( 
.A1(n_198),
.A2(n_216),
.B1(n_169),
.B2(n_38),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_160),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_199),
.B(n_200),
.Y(n_257)
);

INVxp67_ASAP7_75t_L g200 ( 
.A(n_113),
.Y(n_200)
);

AOI21xp5_ASAP7_75t_L g202 ( 
.A1(n_122),
.A2(n_20),
.B(n_14),
.Y(n_202)
);

AO22x2_ASAP7_75t_L g203 ( 
.A1(n_146),
.A2(n_119),
.B1(n_123),
.B2(n_109),
.Y(n_203)
);

AO22x1_ASAP7_75t_L g236 ( 
.A1(n_203),
.A2(n_166),
.B1(n_117),
.B2(n_114),
.Y(n_236)
);

AOI21xp5_ASAP7_75t_SL g204 ( 
.A1(n_122),
.A2(n_27),
.B(n_46),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_204),
.B(n_206),
.Y(n_259)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_120),
.Y(n_205)
);

BUFx3_ASAP7_75t_L g232 ( 
.A(n_205),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_155),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_138),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_207),
.B(n_208),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_157),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_SL g252 ( 
.A(n_209),
.B(n_185),
.Y(n_252)
);

BUFx12f_ASAP7_75t_L g210 ( 
.A(n_144),
.Y(n_210)
);

BUFx12f_ASAP7_75t_L g242 ( 
.A(n_210),
.Y(n_242)
);

BUFx6f_ASAP7_75t_L g211 ( 
.A(n_159),
.Y(n_211)
);

INVx5_ASAP7_75t_L g245 ( 
.A(n_211),
.Y(n_245)
);

INVx6_ASAP7_75t_L g212 ( 
.A(n_141),
.Y(n_212)
);

BUFx3_ASAP7_75t_L g267 ( 
.A(n_212),
.Y(n_267)
);

BUFx3_ASAP7_75t_L g213 ( 
.A(n_136),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_213),
.Y(n_244)
);

OAI22xp33_ASAP7_75t_SL g214 ( 
.A1(n_143),
.A2(n_19),
.B1(n_38),
.B2(n_46),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_214),
.A2(n_123),
.B1(n_121),
.B2(n_143),
.Y(n_241)
);

HB1xp67_ASAP7_75t_L g215 ( 
.A(n_156),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_215),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_124),
.A2(n_38),
.B1(n_18),
.B2(n_11),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_150),
.B(n_52),
.C(n_46),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_217),
.B(n_220),
.Y(n_237)
);

INVx6_ASAP7_75t_L g218 ( 
.A(n_141),
.Y(n_218)
);

AOI22xp33_ASAP7_75t_SL g219 ( 
.A1(n_128),
.A2(n_111),
.B1(n_142),
.B2(n_149),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_154),
.B(n_52),
.Y(n_220)
);

INVx8_ASAP7_75t_L g221 ( 
.A(n_149),
.Y(n_221)
);

AOI22xp33_ASAP7_75t_SL g261 ( 
.A1(n_221),
.A2(n_222),
.B1(n_224),
.B2(n_225),
.Y(n_261)
);

AOI22xp33_ASAP7_75t_SL g222 ( 
.A1(n_128),
.A2(n_161),
.B1(n_127),
.B2(n_163),
.Y(n_222)
);

INVx11_ASAP7_75t_L g223 ( 
.A(n_152),
.Y(n_223)
);

CKINVDCx12_ASAP7_75t_R g246 ( 
.A(n_223),
.Y(n_246)
);

AOI22xp33_ASAP7_75t_SL g224 ( 
.A1(n_127),
.A2(n_52),
.B1(n_46),
.B2(n_35),
.Y(n_224)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_164),
.Y(n_225)
);

INVx3_ASAP7_75t_L g226 ( 
.A(n_134),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_226),
.B(n_228),
.Y(n_251)
);

BUFx6f_ASAP7_75t_L g227 ( 
.A(n_159),
.Y(n_227)
);

AOI22xp33_ASAP7_75t_L g247 ( 
.A1(n_227),
.A2(n_119),
.B1(n_169),
.B2(n_153),
.Y(n_247)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_109),
.Y(n_228)
);

AOI22x1_ASAP7_75t_L g284 ( 
.A1(n_236),
.A2(n_203),
.B1(n_225),
.B2(n_207),
.Y(n_284)
);

AND2x2_ASAP7_75t_L g274 ( 
.A(n_240),
.B(n_241),
.Y(n_274)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_247),
.Y(n_282)
);

OAI22xp33_ASAP7_75t_SL g248 ( 
.A1(n_177),
.A2(n_121),
.B1(n_153),
.B2(n_162),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_248),
.A2(n_250),
.B1(n_255),
.B2(n_200),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_252),
.B(n_194),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_220),
.B(n_35),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_253),
.B(n_203),
.Y(n_273)
);

AOI22xp33_ASAP7_75t_L g254 ( 
.A1(n_177),
.A2(n_125),
.B1(n_115),
.B2(n_170),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_254),
.A2(n_268),
.B1(n_216),
.B2(n_217),
.Y(n_272)
);

OAI22xp33_ASAP7_75t_SL g255 ( 
.A1(n_183),
.A2(n_52),
.B1(n_46),
.B2(n_35),
.Y(n_255)
);

A2O1A1Ixp33_ASAP7_75t_L g263 ( 
.A1(n_201),
.A2(n_134),
.B(n_35),
.C(n_15),
.Y(n_263)
);

AO22x1_ASAP7_75t_L g290 ( 
.A1(n_263),
.A2(n_240),
.B1(n_236),
.B2(n_235),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_201),
.A2(n_180),
.B1(n_202),
.B2(n_198),
.Y(n_268)
);

OR2x2_ASAP7_75t_L g271 ( 
.A(n_259),
.B(n_187),
.Y(n_271)
);

OR2x2_ASAP7_75t_L g324 ( 
.A(n_271),
.B(n_300),
.Y(n_324)
);

AOI22xp5_ASAP7_75t_L g311 ( 
.A1(n_272),
.A2(n_298),
.B1(n_279),
.B2(n_278),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_273),
.B(n_285),
.Y(n_308)
);

BUFx6f_ASAP7_75t_L g275 ( 
.A(n_239),
.Y(n_275)
);

HB1xp67_ASAP7_75t_L g328 ( 
.A(n_275),
.Y(n_328)
);

BUFx3_ASAP7_75t_L g276 ( 
.A(n_246),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g306 ( 
.A(n_276),
.Y(n_306)
);

BUFx2_ASAP7_75t_L g277 ( 
.A(n_245),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g317 ( 
.A(n_277),
.Y(n_317)
);

CKINVDCx16_ASAP7_75t_R g278 ( 
.A(n_257),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_278),
.B(n_279),
.Y(n_313)
);

CKINVDCx16_ASAP7_75t_R g279 ( 
.A(n_257),
.Y(n_279)
);

OAI21xp33_ASAP7_75t_SL g280 ( 
.A1(n_236),
.A2(n_203),
.B(n_204),
.Y(n_280)
);

INVxp67_ASAP7_75t_L g321 ( 
.A(n_280),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_SL g281 ( 
.A(n_230),
.B(n_175),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_281),
.B(n_286),
.Y(n_318)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_229),
.Y(n_283)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_283),
.Y(n_304)
);

OA22x2_ASAP7_75t_L g326 ( 
.A1(n_284),
.A2(n_289),
.B1(n_290),
.B2(n_270),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_237),
.B(n_181),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_232),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_229),
.Y(n_287)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_287),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_237),
.B(n_182),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_288),
.B(n_291),
.Y(n_310)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_243),
.Y(n_292)
);

CKINVDCx16_ASAP7_75t_R g309 ( 
.A(n_292),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_SL g293 ( 
.A(n_230),
.B(n_205),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_293),
.B(n_294),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_253),
.B(n_191),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_250),
.A2(n_188),
.B1(n_228),
.B2(n_193),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_SL g305 ( 
.A1(n_295),
.A2(n_296),
.B1(n_302),
.B2(n_241),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_259),
.A2(n_192),
.B1(n_221),
.B2(n_211),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_243),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_297),
.B(n_299),
.Y(n_332)
);

OAI22xp33_ASAP7_75t_SL g298 ( 
.A1(n_262),
.A2(n_212),
.B1(n_218),
.B2(n_186),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_258),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_262),
.B(n_190),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_L g301 ( 
.A(n_235),
.B(n_210),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_L g329 ( 
.A(n_301),
.B(n_303),
.Y(n_329)
);

AOI22xp5_ASAP7_75t_L g302 ( 
.A1(n_268),
.A2(n_227),
.B1(n_223),
.B2(n_184),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_252),
.B(n_35),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g359 ( 
.A1(n_305),
.A2(n_312),
.B1(n_319),
.B2(n_277),
.Y(n_359)
);

OAI22xp5_ASAP7_75t_SL g337 ( 
.A1(n_311),
.A2(n_322),
.B1(n_323),
.B2(n_327),
.Y(n_337)
);

OAI22xp5_ASAP7_75t_SL g312 ( 
.A1(n_273),
.A2(n_256),
.B1(n_261),
.B2(n_240),
.Y(n_312)
);

AOI21xp5_ASAP7_75t_SL g314 ( 
.A1(n_290),
.A2(n_263),
.B(n_266),
.Y(n_314)
);

CKINVDCx16_ASAP7_75t_R g356 ( 
.A(n_314),
.Y(n_356)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_285),
.B(n_234),
.C(n_251),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g351 ( 
.A(n_315),
.B(n_320),
.C(n_284),
.Y(n_351)
);

FAx1_ASAP7_75t_SL g316 ( 
.A(n_288),
.B(n_263),
.CI(n_251),
.CON(n_316),
.SN(n_316)
);

NAND2xp5_ASAP7_75t_SL g339 ( 
.A(n_316),
.B(n_271),
.Y(n_339)
);

OAI22xp5_ASAP7_75t_SL g319 ( 
.A1(n_290),
.A2(n_266),
.B1(n_258),
.B2(n_234),
.Y(n_319)
);

XOR2xp5_ASAP7_75t_L g320 ( 
.A(n_301),
.B(n_233),
.Y(n_320)
);

AOI22xp5_ASAP7_75t_L g322 ( 
.A1(n_272),
.A2(n_233),
.B1(n_249),
.B2(n_238),
.Y(n_322)
);

AOI22xp5_ASAP7_75t_L g323 ( 
.A1(n_274),
.A2(n_249),
.B1(n_238),
.B2(n_244),
.Y(n_323)
);

OAI21xp5_ASAP7_75t_SL g325 ( 
.A1(n_271),
.A2(n_246),
.B(n_270),
.Y(n_325)
);

AOI21xp5_ASAP7_75t_L g345 ( 
.A1(n_325),
.A2(n_276),
.B(n_289),
.Y(n_345)
);

AO21x1_ASAP7_75t_L g353 ( 
.A1(n_326),
.A2(n_282),
.B(n_295),
.Y(n_353)
);

AOI22xp5_ASAP7_75t_L g327 ( 
.A1(n_274),
.A2(n_244),
.B1(n_245),
.B2(n_265),
.Y(n_327)
);

AOI22xp5_ASAP7_75t_L g330 ( 
.A1(n_274),
.A2(n_265),
.B1(n_260),
.B2(n_264),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_330),
.B(n_296),
.Y(n_336)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_332),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g388 ( 
.A(n_333),
.Y(n_388)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_332),
.Y(n_334)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_334),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_SL g335 ( 
.A(n_310),
.B(n_281),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g370 ( 
.A(n_335),
.B(n_340),
.Y(n_370)
);

OAI21xp33_ASAP7_75t_SL g374 ( 
.A1(n_336),
.A2(n_352),
.B(n_311),
.Y(n_374)
);

XNOR2xp5_ASAP7_75t_L g338 ( 
.A(n_320),
.B(n_303),
.Y(n_338)
);

XNOR2xp5_ASAP7_75t_SL g366 ( 
.A(n_338),
.B(n_339),
.Y(n_366)
);

CKINVDCx20_ASAP7_75t_R g340 ( 
.A(n_318),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_SL g341 ( 
.A(n_313),
.B(n_293),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_L g377 ( 
.A(n_341),
.B(n_342),
.Y(n_377)
);

NOR2xp33_ASAP7_75t_SL g342 ( 
.A(n_313),
.B(n_283),
.Y(n_342)
);

XOR2xp5_ASAP7_75t_L g343 ( 
.A(n_320),
.B(n_294),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g361 ( 
.A(n_343),
.B(n_344),
.C(n_349),
.Y(n_361)
);

XNOR2xp5_ASAP7_75t_L g344 ( 
.A(n_329),
.B(n_302),
.Y(n_344)
);

OAI21xp5_ASAP7_75t_L g363 ( 
.A1(n_345),
.A2(n_347),
.B(n_323),
.Y(n_363)
);

BUFx6f_ASAP7_75t_L g346 ( 
.A(n_328),
.Y(n_346)
);

INVx2_ASAP7_75t_L g383 ( 
.A(n_346),
.Y(n_383)
);

AOI22xp5_ASAP7_75t_SL g347 ( 
.A1(n_321),
.A2(n_284),
.B1(n_282),
.B2(n_299),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_L g348 ( 
.A(n_306),
.B(n_269),
.Y(n_348)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_348),
.Y(n_367)
);

XOR2xp5_ASAP7_75t_L g349 ( 
.A(n_329),
.B(n_297),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_318),
.B(n_292),
.Y(n_350)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_350),
.Y(n_379)
);

XOR2xp5_ASAP7_75t_L g381 ( 
.A(n_351),
.B(n_325),
.Y(n_381)
);

OAI21xp33_ASAP7_75t_L g352 ( 
.A1(n_331),
.A2(n_287),
.B(n_286),
.Y(n_352)
);

OA22x2_ASAP7_75t_L g386 ( 
.A1(n_353),
.A2(n_326),
.B1(n_307),
.B2(n_309),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_SL g354 ( 
.A(n_310),
.B(n_275),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_354),
.B(n_360),
.Y(n_378)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_304),
.Y(n_355)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_355),
.Y(n_384)
);

CKINVDCx16_ASAP7_75t_R g357 ( 
.A(n_304),
.Y(n_357)
);

INVx1_ASAP7_75t_SL g382 ( 
.A(n_357),
.Y(n_382)
);

MAJIxp5_ASAP7_75t_L g358 ( 
.A(n_315),
.B(n_260),
.C(n_264),
.Y(n_358)
);

MAJIxp5_ASAP7_75t_L g364 ( 
.A(n_358),
.B(n_327),
.C(n_330),
.Y(n_364)
);

OAI22xp5_ASAP7_75t_SL g387 ( 
.A1(n_359),
.A2(n_309),
.B1(n_317),
.B2(n_306),
.Y(n_387)
);

NOR2xp33_ASAP7_75t_SL g360 ( 
.A(n_319),
.B(n_269),
.Y(n_360)
);

OAI21xp5_ASAP7_75t_SL g362 ( 
.A1(n_345),
.A2(n_314),
.B(n_324),
.Y(n_362)
);

AOI21xp5_ASAP7_75t_L g390 ( 
.A1(n_362),
.A2(n_363),
.B(n_369),
.Y(n_390)
);

MAJIxp5_ASAP7_75t_L g391 ( 
.A(n_364),
.B(n_365),
.C(n_368),
.Y(n_391)
);

MAJIxp5_ASAP7_75t_L g365 ( 
.A(n_351),
.B(n_308),
.C(n_331),
.Y(n_365)
);

MAJIxp5_ASAP7_75t_L g368 ( 
.A(n_343),
.B(n_308),
.C(n_316),
.Y(n_368)
);

OAI21xp5_ASAP7_75t_L g369 ( 
.A1(n_356),
.A2(n_314),
.B(n_324),
.Y(n_369)
);

AOI22xp5_ASAP7_75t_L g372 ( 
.A1(n_337),
.A2(n_312),
.B1(n_305),
.B2(n_326),
.Y(n_372)
);

AOI22xp5_ASAP7_75t_L g395 ( 
.A1(n_372),
.A2(n_374),
.B1(n_387),
.B2(n_337),
.Y(n_395)
);

XNOR2x1_ASAP7_75t_L g373 ( 
.A(n_349),
.B(n_316),
.Y(n_373)
);

XNOR2xp5_ASAP7_75t_SL g403 ( 
.A(n_373),
.B(n_381),
.Y(n_403)
);

MAJIxp5_ASAP7_75t_L g375 ( 
.A(n_358),
.B(n_316),
.C(n_322),
.Y(n_375)
);

MAJIxp5_ASAP7_75t_L g409 ( 
.A(n_375),
.B(n_341),
.C(n_342),
.Y(n_409)
);

OAI21xp5_ASAP7_75t_SL g376 ( 
.A1(n_360),
.A2(n_324),
.B(n_326),
.Y(n_376)
);

AOI21xp5_ASAP7_75t_L g413 ( 
.A1(n_376),
.A2(n_231),
.B(n_213),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_340),
.B(n_307),
.Y(n_380)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_380),
.Y(n_392)
);

XOR2x2_ASAP7_75t_L g385 ( 
.A(n_339),
.B(n_326),
.Y(n_385)
);

XNOR2xp5_ASAP7_75t_L g399 ( 
.A(n_385),
.B(n_344),
.Y(n_399)
);

CKINVDCx16_ASAP7_75t_R g394 ( 
.A(n_386),
.Y(n_394)
);

XOR2xp5_ASAP7_75t_L g389 ( 
.A(n_338),
.B(n_328),
.Y(n_389)
);

XOR2xp5_ASAP7_75t_L g405 ( 
.A(n_389),
.B(n_350),
.Y(n_405)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_380),
.Y(n_393)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_393),
.Y(n_418)
);

OAI22xp5_ASAP7_75t_SL g428 ( 
.A1(n_395),
.A2(n_407),
.B1(n_363),
.B2(n_364),
.Y(n_428)
);

CKINVDCx20_ASAP7_75t_R g396 ( 
.A(n_370),
.Y(n_396)
);

NOR2xp33_ASAP7_75t_L g420 ( 
.A(n_396),
.B(n_397),
.Y(n_420)
);

OAI21xp5_ASAP7_75t_SL g397 ( 
.A1(n_375),
.A2(n_367),
.B(n_377),
.Y(n_397)
);

BUFx12f_ASAP7_75t_L g398 ( 
.A(n_383),
.Y(n_398)
);

NOR2xp33_ASAP7_75t_L g421 ( 
.A(n_398),
.B(n_404),
.Y(n_421)
);

XNOR2xp5_ASAP7_75t_SL g433 ( 
.A(n_399),
.B(n_405),
.Y(n_433)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_382),
.Y(n_400)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_400),
.Y(n_425)
);

XNOR2xp5_ASAP7_75t_L g401 ( 
.A(n_361),
.B(n_359),
.Y(n_401)
);

MAJIxp5_ASAP7_75t_L g422 ( 
.A(n_401),
.B(n_406),
.C(n_408),
.Y(n_422)
);

CKINVDCx14_ASAP7_75t_R g402 ( 
.A(n_378),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_402),
.B(n_412),
.Y(n_435)
);

HB1xp67_ASAP7_75t_L g404 ( 
.A(n_367),
.Y(n_404)
);

XNOR2xp5_ASAP7_75t_L g406 ( 
.A(n_361),
.B(n_334),
.Y(n_406)
);

AOI22xp5_ASAP7_75t_L g407 ( 
.A1(n_387),
.A2(n_356),
.B1(n_333),
.B2(n_353),
.Y(n_407)
);

XNOR2xp5_ASAP7_75t_L g408 ( 
.A(n_381),
.B(n_347),
.Y(n_408)
);

XOR2xp5_ASAP7_75t_L g423 ( 
.A(n_409),
.B(n_415),
.Y(n_423)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_382),
.Y(n_410)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_410),
.Y(n_427)
);

XNOR2xp5_ASAP7_75t_L g411 ( 
.A(n_389),
.B(n_353),
.Y(n_411)
);

MAJIxp5_ASAP7_75t_L g438 ( 
.A(n_411),
.B(n_414),
.C(n_275),
.Y(n_438)
);

NAND5xp2_ASAP7_75t_L g412 ( 
.A(n_385),
.B(n_336),
.C(n_357),
.D(n_317),
.E(n_355),
.Y(n_412)
);

OAI21xp5_ASAP7_75t_SL g424 ( 
.A1(n_413),
.A2(n_384),
.B(n_383),
.Y(n_424)
);

MAJIxp5_ASAP7_75t_L g414 ( 
.A(n_365),
.B(n_267),
.C(n_232),
.Y(n_414)
);

XOR2xp5_ASAP7_75t_L g415 ( 
.A(n_373),
.B(n_239),
.Y(n_415)
);

NOR2xp33_ASAP7_75t_L g416 ( 
.A(n_388),
.B(n_368),
.Y(n_416)
);

CKINVDCx16_ASAP7_75t_R g417 ( 
.A(n_416),
.Y(n_417)
);

HB1xp67_ASAP7_75t_L g419 ( 
.A(n_392),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_419),
.B(n_432),
.Y(n_443)
);

XNOR2xp5_ASAP7_75t_L g440 ( 
.A(n_424),
.B(n_434),
.Y(n_440)
);

AOI22xp5_ASAP7_75t_L g426 ( 
.A1(n_394),
.A2(n_371),
.B1(n_379),
.B2(n_372),
.Y(n_426)
);

OAI22xp5_ASAP7_75t_SL g452 ( 
.A1(n_426),
.A2(n_429),
.B1(n_398),
.B2(n_269),
.Y(n_452)
);

AOI22xp5_ASAP7_75t_L g445 ( 
.A1(n_428),
.A2(n_437),
.B1(n_415),
.B2(n_405),
.Y(n_445)
);

AOI22xp5_ASAP7_75t_L g429 ( 
.A1(n_411),
.A2(n_379),
.B1(n_386),
.B2(n_376),
.Y(n_429)
);

XOR2xp5_ASAP7_75t_L g430 ( 
.A(n_408),
.B(n_366),
.Y(n_430)
);

XNOR2xp5_ASAP7_75t_SL g449 ( 
.A(n_430),
.B(n_438),
.Y(n_449)
);

OR2x2_ASAP7_75t_L g431 ( 
.A(n_407),
.B(n_378),
.Y(n_431)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_431),
.Y(n_446)
);

NOR3xp33_ASAP7_75t_SL g432 ( 
.A(n_390),
.B(n_369),
.C(n_362),
.Y(n_432)
);

FAx1_ASAP7_75t_SL g434 ( 
.A(n_399),
.B(n_366),
.CI(n_386),
.CON(n_434),
.SN(n_434)
);

INVx4_ASAP7_75t_L g436 ( 
.A(n_398),
.Y(n_436)
);

HB1xp67_ASAP7_75t_L g451 ( 
.A(n_436),
.Y(n_451)
);

OAI22xp5_ASAP7_75t_SL g437 ( 
.A1(n_395),
.A2(n_386),
.B1(n_384),
.B2(n_346),
.Y(n_437)
);

OAI21xp5_ASAP7_75t_L g439 ( 
.A1(n_435),
.A2(n_412),
.B(n_409),
.Y(n_439)
);

AOI21xp5_ASAP7_75t_L g470 ( 
.A1(n_439),
.A2(n_441),
.B(n_448),
.Y(n_470)
);

OAI21xp5_ASAP7_75t_L g441 ( 
.A1(n_435),
.A2(n_391),
.B(n_414),
.Y(n_441)
);

XNOR2xp5_ASAP7_75t_L g442 ( 
.A(n_438),
.B(n_401),
.Y(n_442)
);

MAJIxp5_ASAP7_75t_L g458 ( 
.A(n_442),
.B(n_444),
.C(n_453),
.Y(n_458)
);

MAJIxp5_ASAP7_75t_L g444 ( 
.A(n_422),
.B(n_391),
.C(n_406),
.Y(n_444)
);

OAI22xp5_ASAP7_75t_SL g462 ( 
.A1(n_445),
.A2(n_429),
.B1(n_426),
.B2(n_418),
.Y(n_462)
);

AOI22xp5_ASAP7_75t_L g447 ( 
.A1(n_428),
.A2(n_346),
.B1(n_403),
.B2(n_277),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_L g461 ( 
.A(n_447),
.B(n_456),
.Y(n_461)
);

OAI21xp5_ASAP7_75t_SL g448 ( 
.A1(n_420),
.A2(n_432),
.B(n_427),
.Y(n_448)
);

XOR2xp5_ASAP7_75t_L g450 ( 
.A(n_422),
.B(n_403),
.Y(n_450)
);

XOR2xp5_ASAP7_75t_L g469 ( 
.A(n_450),
.B(n_452),
.Y(n_469)
);

XOR2xp5_ASAP7_75t_L g453 ( 
.A(n_423),
.B(n_242),
.Y(n_453)
);

XOR2xp5_ASAP7_75t_L g454 ( 
.A(n_423),
.B(n_242),
.Y(n_454)
);

MAJIxp5_ASAP7_75t_L g459 ( 
.A(n_454),
.B(n_455),
.C(n_421),
.Y(n_459)
);

MAJIxp5_ASAP7_75t_L g455 ( 
.A(n_433),
.B(n_267),
.C(n_232),
.Y(n_455)
);

XNOR2xp5_ASAP7_75t_SL g456 ( 
.A(n_430),
.B(n_242),
.Y(n_456)
);

OAI22xp5_ASAP7_75t_L g457 ( 
.A1(n_431),
.A2(n_267),
.B1(n_231),
.B2(n_174),
.Y(n_457)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_457),
.Y(n_473)
);

XNOR2xp5_ASAP7_75t_L g487 ( 
.A(n_459),
.B(n_462),
.Y(n_487)
);

MAJIxp5_ASAP7_75t_L g460 ( 
.A(n_442),
.B(n_433),
.C(n_417),
.Y(n_460)
);

MAJIxp5_ASAP7_75t_L g474 ( 
.A(n_460),
.B(n_463),
.C(n_468),
.Y(n_474)
);

MAJIxp5_ASAP7_75t_L g463 ( 
.A(n_444),
.B(n_437),
.C(n_434),
.Y(n_463)
);

OAI22xp5_ASAP7_75t_SL g464 ( 
.A1(n_446),
.A2(n_427),
.B1(n_425),
.B2(n_424),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_464),
.B(n_465),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_L g465 ( 
.A(n_443),
.B(n_425),
.Y(n_465)
);

OAI321xp33_ASAP7_75t_L g466 ( 
.A1(n_439),
.A2(n_434),
.A3(n_436),
.B1(n_239),
.B2(n_242),
.C(n_231),
.Y(n_466)
);

OAI22xp5_ASAP7_75t_L g479 ( 
.A1(n_466),
.A2(n_450),
.B1(n_15),
.B2(n_12),
.Y(n_479)
);

OAI21xp5_ASAP7_75t_SL g467 ( 
.A1(n_451),
.A2(n_455),
.B(n_441),
.Y(n_467)
);

AOI21xp5_ASAP7_75t_L g484 ( 
.A1(n_467),
.A2(n_12),
.B(n_10),
.Y(n_484)
);

MAJIxp5_ASAP7_75t_L g468 ( 
.A(n_449),
.B(n_226),
.C(n_210),
.Y(n_468)
);

MAJIxp5_ASAP7_75t_L g471 ( 
.A(n_449),
.B(n_35),
.C(n_2),
.Y(n_471)
);

MAJIxp5_ASAP7_75t_L g478 ( 
.A(n_471),
.B(n_453),
.C(n_456),
.Y(n_478)
);

INVxp33_ASAP7_75t_L g472 ( 
.A(n_440),
.Y(n_472)
);

NOR2xp33_ASAP7_75t_L g480 ( 
.A(n_472),
.B(n_15),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_SL g476 ( 
.A(n_470),
.B(n_440),
.Y(n_476)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_476),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_L g477 ( 
.A(n_464),
.B(n_454),
.Y(n_477)
);

NOR2xp33_ASAP7_75t_L g496 ( 
.A(n_477),
.B(n_481),
.Y(n_496)
);

XNOR2xp5_ASAP7_75t_L g493 ( 
.A(n_478),
.B(n_1),
.Y(n_493)
);

AOI22xp5_ASAP7_75t_L g488 ( 
.A1(n_479),
.A2(n_462),
.B1(n_10),
.B2(n_3),
.Y(n_488)
);

XOR2xp5_ASAP7_75t_L g497 ( 
.A(n_480),
.B(n_1),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_L g481 ( 
.A(n_473),
.B(n_12),
.Y(n_481)
);

MAJIxp5_ASAP7_75t_L g482 ( 
.A(n_458),
.B(n_1),
.C(n_2),
.Y(n_482)
);

MAJIxp5_ASAP7_75t_L g489 ( 
.A(n_482),
.B(n_459),
.C(n_469),
.Y(n_489)
);

NOR2xp33_ASAP7_75t_L g483 ( 
.A(n_472),
.B(n_12),
.Y(n_483)
);

AOI21xp5_ASAP7_75t_L g490 ( 
.A1(n_483),
.A2(n_484),
.B(n_485),
.Y(n_490)
);

NOR2xp33_ASAP7_75t_SL g485 ( 
.A(n_460),
.B(n_10),
.Y(n_485)
);

NOR2xp67_ASAP7_75t_L g486 ( 
.A(n_463),
.B(n_10),
.Y(n_486)
);

NOR3xp33_ASAP7_75t_L g495 ( 
.A(n_486),
.B(n_6),
.C(n_2),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_SL g504 ( 
.A(n_488),
.B(n_492),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_489),
.Y(n_505)
);

OAI22xp5_ASAP7_75t_L g491 ( 
.A1(n_475),
.A2(n_461),
.B1(n_458),
.B2(n_468),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_L g499 ( 
.A(n_491),
.B(n_493),
.Y(n_499)
);

AOI21xp5_ASAP7_75t_L g492 ( 
.A1(n_474),
.A2(n_469),
.B(n_471),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_495),
.B(n_497),
.Y(n_500)
);

XNOR2xp5_ASAP7_75t_L g498 ( 
.A(n_474),
.B(n_6),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_L g503 ( 
.A(n_498),
.B(n_4),
.Y(n_503)
);

MAJIxp5_ASAP7_75t_L g501 ( 
.A(n_489),
.B(n_487),
.C(n_478),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_L g511 ( 
.A(n_501),
.B(n_502),
.Y(n_511)
);

OAI22xp5_ASAP7_75t_SL g502 ( 
.A1(n_494),
.A2(n_487),
.B1(n_482),
.B2(n_6),
.Y(n_502)
);

CKINVDCx16_ASAP7_75t_R g508 ( 
.A(n_503),
.Y(n_508)
);

INVxp67_ASAP7_75t_L g506 ( 
.A(n_498),
.Y(n_506)
);

NOR2xp33_ASAP7_75t_SL g509 ( 
.A(n_506),
.B(n_493),
.Y(n_509)
);

OAI21xp5_ASAP7_75t_SL g507 ( 
.A1(n_505),
.A2(n_496),
.B(n_490),
.Y(n_507)
);

NOR2xp33_ASAP7_75t_SL g512 ( 
.A(n_507),
.B(n_504),
.Y(n_512)
);

OAI21xp5_ASAP7_75t_L g514 ( 
.A1(n_509),
.A2(n_510),
.B(n_506),
.Y(n_514)
);

INVxp67_ASAP7_75t_L g510 ( 
.A(n_501),
.Y(n_510)
);

NOR3xp33_ASAP7_75t_L g515 ( 
.A(n_512),
.B(n_500),
.C(n_508),
.Y(n_515)
);

NAND2xp33_ASAP7_75t_SL g513 ( 
.A(n_511),
.B(n_499),
.Y(n_513)
);

A2O1A1Ixp33_ASAP7_75t_L g516 ( 
.A1(n_513),
.A2(n_514),
.B(n_497),
.C(n_4),
.Y(n_516)
);

INVxp67_ASAP7_75t_L g517 ( 
.A(n_515),
.Y(n_517)
);

HB1xp67_ASAP7_75t_L g518 ( 
.A(n_517),
.Y(n_518)
);

OAI21xp5_ASAP7_75t_SL g519 ( 
.A1(n_518),
.A2(n_516),
.B(n_4),
.Y(n_519)
);

AOI21xp5_ASAP7_75t_L g520 ( 
.A1(n_519),
.A2(n_5),
.B(n_443),
.Y(n_520)
);

XOR2x2_ASAP7_75t_SL g521 ( 
.A(n_520),
.B(n_5),
.Y(n_521)
);


endmodule