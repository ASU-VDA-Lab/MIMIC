module fake_jpeg_5452_n_251 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_251);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_251;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_212;
wire n_131;
wire n_56;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_4),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_4),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_12),
.Y(n_16)
);

INVx4_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

INVx11_ASAP7_75t_SL g18 ( 
.A(n_1),
.Y(n_18)
);

INVx8_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

INVx4_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_8),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

INVx11_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_1),
.Y(n_28)
);

BUFx10_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_18),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_30),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_23),
.Y(n_31)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_31),
.Y(n_54)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_18),
.Y(n_32)
);

INVx5_ASAP7_75t_L g44 ( 
.A(n_32),
.Y(n_44)
);

AND2x2_ASAP7_75t_SL g33 ( 
.A(n_29),
.B(n_0),
.Y(n_33)
);

AOI21xp33_ASAP7_75t_L g42 ( 
.A1(n_33),
.A2(n_29),
.B(n_23),
.Y(n_42)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_26),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_34),
.B(n_36),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_23),
.Y(n_35)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_35),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_27),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_15),
.B(n_6),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_SL g45 ( 
.A(n_37),
.B(n_15),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_27),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_38),
.B(n_39),
.Y(n_51)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_17),
.Y(n_39)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_33),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_40),
.B(n_43),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_SL g64 ( 
.A(n_42),
.B(n_49),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g43 ( 
.A(n_37),
.B(n_15),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_45),
.B(n_46),
.Y(n_71)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_33),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_L g47 ( 
.A1(n_33),
.A2(n_39),
.B1(n_19),
.B2(n_34),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_47),
.A2(n_57),
.B1(n_17),
.B2(n_20),
.Y(n_69)
);

OAI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_32),
.A2(n_19),
.B1(n_27),
.B2(n_25),
.Y(n_48)
);

OAI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_48),
.A2(n_14),
.B1(n_25),
.B2(n_28),
.Y(n_65)
);

AOI21xp33_ASAP7_75t_L g49 ( 
.A1(n_30),
.A2(n_29),
.B(n_23),
.Y(n_49)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_31),
.Y(n_52)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_52),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_35),
.B(n_21),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_SL g67 ( 
.A(n_55),
.B(n_22),
.Y(n_67)
);

INVx2_ASAP7_75t_SL g56 ( 
.A(n_36),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_56),
.B(n_58),
.Y(n_72)
);

OA22x2_ASAP7_75t_L g57 ( 
.A1(n_36),
.A2(n_29),
.B1(n_23),
.B2(n_19),
.Y(n_57)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_30),
.Y(n_58)
);

INVx13_ASAP7_75t_L g59 ( 
.A(n_44),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_59),
.B(n_70),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_40),
.A2(n_19),
.B1(n_20),
.B2(n_17),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_60),
.A2(n_74),
.B1(n_16),
.B2(n_54),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_55),
.B(n_29),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_62),
.B(n_65),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_47),
.B(n_29),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_66),
.B(n_67),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_41),
.B(n_52),
.Y(n_68)
);

XNOR2xp5_ASAP7_75t_L g97 ( 
.A(n_68),
.B(n_41),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_69),
.A2(n_56),
.B1(n_51),
.B2(n_58),
.Y(n_86)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_44),
.Y(n_70)
);

OR2x2_ASAP7_75t_L g73 ( 
.A(n_57),
.B(n_28),
.Y(n_73)
);

OAI21xp5_ASAP7_75t_SL g88 ( 
.A1(n_73),
.A2(n_51),
.B(n_16),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_46),
.A2(n_20),
.B1(n_24),
.B2(n_22),
.Y(n_74)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_57),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_75),
.B(n_78),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_57),
.A2(n_14),
.B1(n_21),
.B2(n_24),
.Y(n_76)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_76),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_45),
.B(n_24),
.Y(n_77)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_77),
.Y(n_89)
);

CKINVDCx9p33_ASAP7_75t_R g78 ( 
.A(n_53),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_43),
.B(n_22),
.Y(n_79)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_79),
.Y(n_101)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_50),
.Y(n_80)
);

INVx13_ASAP7_75t_L g84 ( 
.A(n_80),
.Y(n_84)
);

OR2x2_ASAP7_75t_L g81 ( 
.A(n_73),
.B(n_56),
.Y(n_81)
);

AND2x2_ASAP7_75t_L g122 ( 
.A(n_81),
.B(n_97),
.Y(n_122)
);

INVx1_ASAP7_75t_SL g82 ( 
.A(n_67),
.Y(n_82)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_82),
.Y(n_104)
);

INVx5_ASAP7_75t_L g83 ( 
.A(n_59),
.Y(n_83)
);

CKINVDCx16_ASAP7_75t_R g107 ( 
.A(n_83),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_86),
.A2(n_66),
.B1(n_74),
.B2(n_60),
.Y(n_105)
);

XNOR2xp5_ASAP7_75t_L g115 ( 
.A(n_88),
.B(n_95),
.Y(n_115)
);

BUFx2_ASAP7_75t_L g90 ( 
.A(n_78),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_90),
.Y(n_106)
);

CKINVDCx16_ASAP7_75t_R g91 ( 
.A(n_72),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_91),
.B(n_93),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_68),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_92),
.Y(n_113)
);

INVx13_ASAP7_75t_L g93 ( 
.A(n_61),
.Y(n_93)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_70),
.Y(n_94)
);

INVx4_ASAP7_75t_L g116 ( 
.A(n_94),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_L g95 ( 
.A1(n_64),
.A2(n_50),
.B(n_16),
.Y(n_95)
);

OR2x2_ASAP7_75t_SL g99 ( 
.A(n_71),
.B(n_10),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g124 ( 
.A(n_99),
.B(n_100),
.Y(n_124)
);

NAND3xp33_ASAP7_75t_L g103 ( 
.A(n_71),
.B(n_54),
.C(n_23),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_103),
.B(n_63),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_105),
.A2(n_112),
.B1(n_120),
.B2(n_63),
.Y(n_133)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_85),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_108),
.B(n_114),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_98),
.A2(n_66),
.B1(n_64),
.B2(n_69),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_109),
.A2(n_123),
.B1(n_121),
.B2(n_111),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_92),
.B(n_97),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_111),
.B(n_121),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_98),
.A2(n_75),
.B1(n_69),
.B2(n_76),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_101),
.B(n_89),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_117),
.B(n_119),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_102),
.B(n_62),
.C(n_68),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_118),
.B(n_125),
.C(n_91),
.Y(n_138)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_86),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_96),
.A2(n_75),
.B1(n_76),
.B2(n_73),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_102),
.Y(n_121)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_96),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_123),
.B(n_82),
.Y(n_142)
);

XNOR2x1_ASAP7_75t_L g125 ( 
.A(n_95),
.B(n_62),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_101),
.B(n_77),
.Y(n_126)
);

CKINVDCx14_ASAP7_75t_R g143 ( 
.A(n_126),
.Y(n_143)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_110),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_127),
.B(n_128),
.Y(n_162)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_118),
.Y(n_128)
);

AOI21xp5_ASAP7_75t_L g129 ( 
.A1(n_125),
.A2(n_88),
.B(n_81),
.Y(n_129)
);

INVxp67_ASAP7_75t_L g164 ( 
.A(n_129),
.Y(n_164)
);

HB1xp67_ASAP7_75t_L g130 ( 
.A(n_116),
.Y(n_130)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_130),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_119),
.A2(n_89),
.B1(n_81),
.B2(n_73),
.Y(n_131)
);

INVxp67_ASAP7_75t_L g168 ( 
.A(n_131),
.Y(n_168)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_109),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_132),
.B(n_135),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_133),
.B(n_144),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_134),
.A2(n_146),
.B1(n_124),
.B2(n_108),
.Y(n_152)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_122),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_122),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_136),
.B(n_142),
.Y(n_159)
);

BUFx5_ASAP7_75t_L g137 ( 
.A(n_116),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_137),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_138),
.B(n_141),
.C(n_148),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_122),
.B(n_61),
.C(n_80),
.Y(n_141)
);

AOI21xp5_ASAP7_75t_L g144 ( 
.A1(n_105),
.A2(n_87),
.B(n_79),
.Y(n_144)
);

OAI31xp33_ASAP7_75t_SL g145 ( 
.A1(n_120),
.A2(n_99),
.A3(n_65),
.B(n_84),
.Y(n_145)
);

A2O1A1O1Ixp25_ASAP7_75t_L g150 ( 
.A1(n_145),
.A2(n_115),
.B(n_124),
.C(n_112),
.D(n_104),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_113),
.A2(n_72),
.B1(n_70),
.B2(n_84),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_SL g148 ( 
.A1(n_104),
.A2(n_84),
.B(n_94),
.Y(n_148)
);

FAx1_ASAP7_75t_SL g177 ( 
.A(n_150),
.B(n_152),
.CI(n_144),
.CON(n_177),
.SN(n_177)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_146),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_151),
.B(n_153),
.Y(n_176)
);

NOR2x1_ASAP7_75t_L g153 ( 
.A(n_145),
.B(n_115),
.Y(n_153)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_140),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_156),
.B(n_158),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_SL g158 ( 
.A(n_143),
.B(n_124),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_SL g160 ( 
.A(n_139),
.B(n_107),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_160),
.B(n_161),
.Y(n_185)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_140),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_137),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_163),
.Y(n_183)
);

BUFx3_ASAP7_75t_L g165 ( 
.A(n_148),
.Y(n_165)
);

CKINVDCx16_ASAP7_75t_R g186 ( 
.A(n_165),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_128),
.B(n_83),
.C(n_93),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_166),
.B(n_138),
.C(n_141),
.Y(n_170)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_142),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_167),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_170),
.B(n_174),
.C(n_175),
.Y(n_192)
);

XNOR2x1_ASAP7_75t_SL g171 ( 
.A(n_153),
.B(n_136),
.Y(n_171)
);

XNOR2x1_ASAP7_75t_L g190 ( 
.A(n_171),
.B(n_168),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_151),
.A2(n_132),
.B1(n_135),
.B2(n_134),
.Y(n_172)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_172),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_164),
.A2(n_133),
.B1(n_131),
.B2(n_147),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_173),
.A2(n_180),
.B1(n_184),
.B2(n_162),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_L g174 ( 
.A(n_169),
.B(n_129),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_155),
.B(n_166),
.C(n_157),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_177),
.B(n_150),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_155),
.B(n_147),
.C(n_127),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_178),
.B(n_179),
.C(n_181),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_157),
.B(n_106),
.C(n_93),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_164),
.A2(n_38),
.B1(n_53),
.B2(n_26),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_159),
.B(n_38),
.C(n_53),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_168),
.A2(n_26),
.B1(n_59),
.B2(n_2),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_183),
.B(n_167),
.Y(n_188)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_188),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_L g207 ( 
.A(n_190),
.B(n_196),
.Y(n_207)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_185),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_191),
.B(n_195),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_183),
.B(n_156),
.Y(n_193)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_193),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_194),
.B(n_198),
.Y(n_208)
);

INVx1_ASAP7_75t_SL g195 ( 
.A(n_171),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g196 ( 
.A(n_170),
.B(n_169),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g197 ( 
.A(n_174),
.B(n_152),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_197),
.B(n_202),
.C(n_178),
.Y(n_210)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_181),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_186),
.A2(n_159),
.B1(n_161),
.B2(n_165),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_L g213 ( 
.A1(n_199),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_201),
.B(n_177),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_176),
.B(n_154),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_189),
.A2(n_172),
.B1(n_187),
.B2(n_177),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_204),
.A2(n_211),
.B1(n_213),
.B2(n_215),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_190),
.A2(n_173),
.B1(n_187),
.B2(n_175),
.Y(n_206)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_206),
.Y(n_220)
);

INVxp67_ASAP7_75t_L g221 ( 
.A(n_209),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_210),
.B(n_212),
.C(n_3),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_197),
.A2(n_179),
.B1(n_182),
.B2(n_180),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_192),
.B(n_149),
.C(n_184),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_195),
.A2(n_1),
.B1(n_2),
.B2(n_59),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_205),
.B(n_202),
.Y(n_216)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_216),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_214),
.B(n_200),
.Y(n_218)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_218),
.Y(n_232)
);

OAI321xp33_ASAP7_75t_L g219 ( 
.A1(n_203),
.A2(n_200),
.A3(n_192),
.B1(n_5),
.B2(n_6),
.C(n_7),
.Y(n_219)
);

OR2x2_ASAP7_75t_L g231 ( 
.A(n_219),
.B(n_222),
.Y(n_231)
);

OAI21x1_ASAP7_75t_L g222 ( 
.A1(n_211),
.A2(n_3),
.B(n_4),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_SL g233 ( 
.A(n_223),
.B(n_224),
.Y(n_233)
);

NOR2xp67_ASAP7_75t_L g224 ( 
.A(n_206),
.B(n_204),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_208),
.B(n_90),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_225),
.B(n_215),
.Y(n_226)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_226),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_220),
.A2(n_210),
.B1(n_212),
.B2(n_207),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_227),
.B(n_9),
.Y(n_239)
);

OAI21xp5_ASAP7_75t_SL g229 ( 
.A1(n_221),
.A2(n_207),
.B(n_5),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_229),
.B(n_13),
.C(n_10),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_217),
.B(n_90),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_SL g235 ( 
.A(n_230),
.B(n_223),
.Y(n_235)
);

CKINVDCx16_ASAP7_75t_R g241 ( 
.A(n_235),
.Y(n_241)
);

AOI21xp5_ASAP7_75t_SL g236 ( 
.A1(n_229),
.A2(n_221),
.B(n_7),
.Y(n_236)
);

CKINVDCx16_ASAP7_75t_R g244 ( 
.A(n_236),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_SL g237 ( 
.A(n_232),
.B(n_3),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_237),
.A2(n_238),
.B1(n_231),
.B2(n_11),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_239),
.B(n_234),
.C(n_228),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_240),
.B(n_243),
.C(n_231),
.Y(n_245)
);

AOI322xp5_ASAP7_75t_L g247 ( 
.A1(n_242),
.A2(n_244),
.A3(n_240),
.B1(n_12),
.B2(n_13),
.C1(n_11),
.C2(n_9),
.Y(n_247)
);

OAI21x1_ASAP7_75t_SL g243 ( 
.A1(n_239),
.A2(n_233),
.B(n_227),
.Y(n_243)
);

AND2x2_ASAP7_75t_L g248 ( 
.A(n_245),
.B(n_246),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_241),
.B(n_9),
.C(n_11),
.Y(n_246)
);

INVxp67_ASAP7_75t_L g249 ( 
.A(n_247),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_248),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_250),
.B(n_249),
.Y(n_251)
);


endmodule