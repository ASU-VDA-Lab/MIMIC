module fake_netlist_5_1795_n_83 (n_16, n_0, n_12, n_9, n_18, n_22, n_1, n_8, n_10, n_21, n_4, n_11, n_17, n_19, n_7, n_15, n_20, n_5, n_14, n_2, n_13, n_3, n_6, n_83);

input n_16;
input n_0;
input n_12;
input n_9;
input n_18;
input n_22;
input n_1;
input n_8;
input n_10;
input n_21;
input n_4;
input n_11;
input n_17;
input n_19;
input n_7;
input n_15;
input n_20;
input n_5;
input n_14;
input n_2;
input n_13;
input n_3;
input n_6;

output n_83;

wire n_82;
wire n_24;
wire n_61;
wire n_75;
wire n_65;
wire n_78;
wire n_74;
wire n_57;
wire n_37;
wire n_31;
wire n_66;
wire n_60;
wire n_43;
wire n_58;
wire n_69;
wire n_42;
wire n_45;
wire n_46;
wire n_38;
wire n_80;
wire n_35;
wire n_73;
wire n_30;
wire n_33;
wire n_23;
wire n_29;
wire n_79;
wire n_47;
wire n_25;
wire n_53;
wire n_44;
wire n_40;
wire n_34;
wire n_62;
wire n_71;
wire n_59;
wire n_26;
wire n_55;
wire n_49;
wire n_39;
wire n_54;
wire n_67;
wire n_36;
wire n_76;
wire n_27;
wire n_64;
wire n_77;
wire n_81;
wire n_28;
wire n_70;
wire n_68;
wire n_72;
wire n_32;
wire n_41;
wire n_56;
wire n_51;
wire n_63;
wire n_48;
wire n_50;
wire n_52;

BUFx2_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

AND2x2_ASAP7_75t_L g24 ( 
.A(n_21),
.B(n_16),
.Y(n_24)
);

AND2x2_ASAP7_75t_L g25 ( 
.A(n_22),
.B(n_10),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

BUFx8_ASAP7_75t_SL g27 ( 
.A(n_14),
.Y(n_27)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

AOI22xp5_ASAP7_75t_L g29 ( 
.A1(n_7),
.A2(n_15),
.B1(n_13),
.B2(n_20),
.Y(n_29)
);

INVx5_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

NAND2xp33_ASAP7_75t_L g32 ( 
.A(n_11),
.B(n_17),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_5),
.B(n_3),
.Y(n_33)
);

XNOR2x2_ASAP7_75t_L g34 ( 
.A(n_18),
.B(n_19),
.Y(n_34)
);

INVx5_ASAP7_75t_L g35 ( 
.A(n_4),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_1),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_4),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_8),
.Y(n_38)
);

AND2x2_ASAP7_75t_L g39 ( 
.A(n_9),
.B(n_2),
.Y(n_39)
);

INVx2_ASAP7_75t_SL g40 ( 
.A(n_30),
.Y(n_40)
);

INVxp67_ASAP7_75t_L g41 ( 
.A(n_23),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_26),
.B(n_0),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_26),
.B(n_2),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_L g44 ( 
.A1(n_39),
.A2(n_37),
.B1(n_28),
.B2(n_24),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_28),
.B(n_35),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_30),
.B(n_35),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_28),
.B(n_30),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_30),
.B(n_35),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_30),
.B(n_35),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_35),
.B(n_38),
.Y(n_50)
);

OAI21x1_ASAP7_75t_L g51 ( 
.A1(n_50),
.A2(n_25),
.B(n_24),
.Y(n_51)
);

OAI21x1_ASAP7_75t_L g52 ( 
.A1(n_46),
.A2(n_31),
.B(n_29),
.Y(n_52)
);

A2O1A1Ixp33_ASAP7_75t_L g53 ( 
.A1(n_45),
.A2(n_32),
.B(n_33),
.C(n_36),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_44),
.B(n_37),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_53),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_52),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_51),
.Y(n_57)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_54),
.Y(n_58)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_54),
.Y(n_59)
);

OR2x6_ASAP7_75t_L g60 ( 
.A(n_54),
.B(n_41),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_55),
.Y(n_61)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_56),
.Y(n_62)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_55),
.Y(n_63)
);

OR2x2_ASAP7_75t_L g64 ( 
.A(n_58),
.B(n_59),
.Y(n_64)
);

AND2x2_ASAP7_75t_L g65 ( 
.A(n_60),
.B(n_47),
.Y(n_65)
);

AND2x2_ASAP7_75t_L g66 ( 
.A(n_60),
.B(n_43),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_63),
.Y(n_67)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_63),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_61),
.B(n_57),
.Y(n_69)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_61),
.Y(n_70)
);

OR2x6_ASAP7_75t_L g71 ( 
.A(n_70),
.B(n_64),
.Y(n_71)
);

OAI21xp5_ASAP7_75t_L g72 ( 
.A1(n_69),
.A2(n_62),
.B(n_65),
.Y(n_72)
);

NAND3xp33_ASAP7_75t_L g73 ( 
.A(n_72),
.B(n_65),
.C(n_66),
.Y(n_73)
);

OAI211xp5_ASAP7_75t_SL g74 ( 
.A1(n_71),
.A2(n_42),
.B(n_32),
.C(n_67),
.Y(n_74)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_73),
.B(n_68),
.Y(n_75)
);

NOR2x1_ASAP7_75t_L g76 ( 
.A(n_74),
.B(n_69),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_75),
.Y(n_77)
);

OR2x2_ASAP7_75t_L g78 ( 
.A(n_76),
.B(n_34),
.Y(n_78)
);

AOI21xp5_ASAP7_75t_L g79 ( 
.A1(n_78),
.A2(n_62),
.B(n_34),
.Y(n_79)
);

OAI21x1_ASAP7_75t_L g80 ( 
.A1(n_77),
.A2(n_45),
.B(n_48),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_79),
.B(n_49),
.Y(n_81)
);

AOI21xp5_ASAP7_75t_L g82 ( 
.A1(n_80),
.A2(n_27),
.B(n_40),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_81),
.B(n_82),
.Y(n_83)
);


endmodule