module real_jpeg_21687_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_166;
wire n_176;
wire n_104;
wire n_194;
wire n_153;
wire n_161;
wire n_64;
wire n_177;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_200;
wire n_48;
wire n_164;
wire n_184;
wire n_140;
wire n_126;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_93;
wire n_141;
wire n_95;
wire n_65;
wire n_33;
wire n_188;
wire n_139;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_160;
wire n_172;
wire n_45;
wire n_112;
wire n_42;
wire n_145;
wire n_18;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_165;
wire n_134;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_198;
wire n_192;
wire n_100;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_117;
wire n_193;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_150;
wire n_30;
wire n_158;
wire n_149;
wire n_144;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_185;
wire n_55;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_167;
wire n_179;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;

AOI22xp5_ASAP7_75t_SL g39 ( 
.A1(n_0),
.A2(n_40),
.B1(n_41),
.B2(n_42),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_0),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_0),
.A2(n_27),
.B1(n_30),
.B2(n_42),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_1),
.A2(n_40),
.B1(n_41),
.B2(n_54),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_1),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_1),
.A2(n_54),
.B1(n_62),
.B2(n_63),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_1),
.A2(n_27),
.B1(n_30),
.B2(n_54),
.Y(n_162)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_2),
.A2(n_62),
.B1(n_63),
.B2(n_69),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_2),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_2),
.A2(n_27),
.B1(n_30),
.B2(n_69),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_SL g177 ( 
.A1(n_2),
.A2(n_40),
.B1(n_41),
.B2(n_69),
.Y(n_177)
);

BUFx16f_ASAP7_75t_L g72 ( 
.A(n_3),
.Y(n_72)
);

INVx13_ASAP7_75t_L g75 ( 
.A(n_4),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_4),
.A2(n_62),
.B1(n_63),
.B2(n_75),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_5),
.A2(n_62),
.B1(n_63),
.B2(n_67),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_5),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_5),
.A2(n_67),
.B1(n_72),
.B2(n_80),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_5),
.A2(n_27),
.B1(n_30),
.B2(n_67),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_SL g159 ( 
.A1(n_5),
.A2(n_40),
.B1(n_41),
.B2(n_67),
.Y(n_159)
);

AOI22xp33_ASAP7_75t_L g34 ( 
.A1(n_6),
.A2(n_27),
.B1(n_30),
.B2(n_35),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_6),
.Y(n_35)
);

OAI22xp33_ASAP7_75t_SL g44 ( 
.A1(n_6),
.A2(n_35),
.B1(n_40),
.B2(n_41),
.Y(n_44)
);

INVx6_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

INVx8_ASAP7_75t_L g88 ( 
.A(n_7),
.Y(n_88)
);

AOI21xp5_ASAP7_75t_L g113 ( 
.A1(n_7),
.A2(n_87),
.B(n_114),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g29 ( 
.A1(n_8),
.A2(n_27),
.B1(n_30),
.B2(n_31),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_8),
.Y(n_31)
);

BUFx8_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

BUFx12_ASAP7_75t_L g63 ( 
.A(n_10),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_11),
.A2(n_72),
.B1(n_79),
.B2(n_80),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_11),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_11),
.A2(n_62),
.B1(n_63),
.B2(n_79),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_11),
.A2(n_40),
.B1(n_41),
.B2(n_79),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_11),
.A2(n_27),
.B1(n_30),
.B2(n_79),
.Y(n_141)
);

INVx13_ASAP7_75t_L g61 ( 
.A(n_12),
.Y(n_61)
);

CKINVDCx14_ASAP7_75t_R g73 ( 
.A(n_13),
.Y(n_73)
);

AOI21xp33_ASAP7_75t_L g133 ( 
.A1(n_13),
.A2(n_14),
.B(n_27),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_SL g136 ( 
.A1(n_13),
.A2(n_40),
.B1(n_41),
.B2(n_73),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_13),
.A2(n_26),
.B1(n_141),
.B2(n_145),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_13),
.B(n_156),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_13),
.B(n_62),
.Y(n_170)
);

AOI21xp33_ASAP7_75t_L g174 ( 
.A1(n_13),
.A2(n_62),
.B(n_170),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_SL g37 ( 
.A1(n_14),
.A2(n_27),
.B1(n_30),
.B2(n_38),
.Y(n_37)
);

INVx11_ASAP7_75t_L g38 ( 
.A(n_14),
.Y(n_38)
);

A2O1A1Ixp33_ASAP7_75t_L g46 ( 
.A1(n_14),
.A2(n_37),
.B(n_40),
.C(n_47),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_14),
.B(n_40),
.Y(n_47)
);

INVx11_ASAP7_75t_SL g40 ( 
.A(n_15),
.Y(n_40)
);

XNOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_117),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_115),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_19),
.Y(n_18)
);

AND2x2_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_103),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_20),
.B(n_103),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g20 ( 
.A1(n_21),
.A2(n_22),
.B1(n_81),
.B2(n_102),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

XNOR2xp5_ASAP7_75t_SL g22 ( 
.A(n_23),
.B(n_49),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_25),
.B1(n_36),
.B2(n_48),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_25),
.Y(n_24)
);

OAI21xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_29),
.B(n_32),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_26),
.A2(n_29),
.B1(n_86),
.B2(n_88),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_26),
.B(n_34),
.Y(n_114)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_26),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_26),
.A2(n_88),
.B1(n_126),
.B2(n_141),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_L g160 ( 
.A1(n_26),
.A2(n_129),
.B(n_161),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_28),
.Y(n_26)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_27),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_28),
.B(n_34),
.Y(n_33)
);

INVx5_ASAP7_75t_L g127 ( 
.A(n_28),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_30),
.B(n_147),
.Y(n_146)
);

CKINVDCx14_ASAP7_75t_R g32 ( 
.A(n_33),
.Y(n_32)
);

AOI21xp5_ASAP7_75t_L g168 ( 
.A1(n_33),
.A2(n_124),
.B(n_162),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_36),
.Y(n_48)
);

OAI21xp5_ASAP7_75t_L g36 ( 
.A1(n_37),
.A2(n_39),
.B(n_43),
.Y(n_36)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_37),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_37),
.A2(n_46),
.B1(n_136),
.B2(n_137),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_37),
.B(n_73),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_37),
.A2(n_46),
.B1(n_137),
.B2(n_159),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_37),
.A2(n_46),
.B1(n_159),
.B2(n_177),
.Y(n_176)
);

A2O1A1Ixp33_ASAP7_75t_L g132 ( 
.A1(n_38),
.A2(n_41),
.B(n_73),
.C(n_133),
.Y(n_132)
);

INVx11_ASAP7_75t_L g41 ( 
.A(n_40),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_40),
.A2(n_41),
.B1(n_60),
.B2(n_61),
.Y(n_65)
);

AOI32xp33_ASAP7_75t_L g169 ( 
.A1(n_40),
.A2(n_61),
.A3(n_63),
.B1(n_170),
.B2(n_171),
.Y(n_169)
);

NAND2xp33_ASAP7_75t_SL g171 ( 
.A(n_41),
.B(n_60),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_44),
.B(n_45),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_SL g55 ( 
.A(n_44),
.B(n_56),
.Y(n_55)
);

INVxp67_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

OAI21xp5_ASAP7_75t_SL g51 ( 
.A1(n_46),
.A2(n_52),
.B(n_55),
.Y(n_51)
);

OAI21xp5_ASAP7_75t_SL g192 ( 
.A1(n_46),
.A2(n_177),
.B(n_193),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g49 ( 
.A(n_50),
.B(n_57),
.C(n_70),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_50),
.A2(n_51),
.B1(n_57),
.B2(n_58),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_51),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_53),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_53),
.B(n_56),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_58),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_59),
.A2(n_65),
.B1(n_66),
.B2(n_68),
.Y(n_58)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_59),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_59),
.A2(n_65),
.B1(n_66),
.B2(n_110),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_59),
.A2(n_65),
.B1(n_110),
.B2(n_174),
.Y(n_173)
);

A2O1A1Ixp33_ASAP7_75t_L g59 ( 
.A1(n_60),
.A2(n_62),
.B(n_64),
.C(n_65),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_60),
.B(n_62),
.Y(n_64)
);

INVx11_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_62),
.B(n_75),
.Y(n_84)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_63),
.A2(n_71),
.B1(n_76),
.B2(n_84),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_65),
.B(n_101),
.Y(n_100)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_65),
.Y(n_156)
);

CKINVDCx16_ASAP7_75t_R g99 ( 
.A(n_68),
.Y(n_99)
);

XNOR2xp5_ASAP7_75t_SL g104 ( 
.A(n_70),
.B(n_105),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_71),
.A2(n_74),
.B1(n_77),
.B2(n_78),
.Y(n_70)
);

HAxp5_ASAP7_75t_SL g71 ( 
.A(n_72),
.B(n_73),
.CON(n_71),
.SN(n_71)
);

O2A1O1Ixp33_ASAP7_75t_L g74 ( 
.A1(n_72),
.A2(n_75),
.B(n_76),
.C(n_77),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_72),
.B(n_75),
.Y(n_76)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_72),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_73),
.B(n_95),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_73),
.B(n_88),
.Y(n_147)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_74),
.Y(n_92)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_77),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_78),
.Y(n_93)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_81),
.Y(n_102)
);

XOR2xp5_ASAP7_75t_L g81 ( 
.A(n_82),
.B(n_89),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_83),
.B(n_85),
.Y(n_82)
);

XOR2xp5_ASAP7_75t_L g107 ( 
.A(n_83),
.B(n_85),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_87),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_90),
.A2(n_91),
.B1(n_96),
.B2(n_97),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_91),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_92),
.A2(n_93),
.B1(n_94),
.B2(n_95),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_97),
.Y(n_96)
);

AOI21xp5_ASAP7_75t_L g97 ( 
.A1(n_98),
.A2(n_99),
.B(n_100),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_104),
.B(n_106),
.C(n_108),
.Y(n_103)
);

XOR2xp5_ASAP7_75t_L g197 ( 
.A(n_104),
.B(n_198),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g198 ( 
.A1(n_106),
.A2(n_107),
.B1(n_108),
.B2(n_199),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_107),
.Y(n_106)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_108),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_109),
.B(n_111),
.C(n_112),
.Y(n_108)
);

XNOR2xp5_ASAP7_75t_SL g186 ( 
.A(n_109),
.B(n_187),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_111),
.A2(n_112),
.B1(n_113),
.B2(n_188),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_111),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_113),
.Y(n_112)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

AOI21xp5_ASAP7_75t_L g117 ( 
.A1(n_118),
.A2(n_195),
.B(n_200),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_SL g118 ( 
.A1(n_119),
.A2(n_182),
.B(n_194),
.Y(n_118)
);

AOI21xp5_ASAP7_75t_L g119 ( 
.A1(n_120),
.A2(n_164),
.B(n_181),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_SL g120 ( 
.A1(n_121),
.A2(n_150),
.B(n_163),
.Y(n_120)
);

AOI21xp5_ASAP7_75t_L g121 ( 
.A1(n_122),
.A2(n_138),
.B(n_149),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_123),
.B(n_130),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_123),
.B(n_130),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_124),
.A2(n_125),
.B1(n_127),
.B2(n_128),
.Y(n_123)
);

INVxp67_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVx4_ASAP7_75t_L g145 ( 
.A(n_127),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_127),
.B(n_162),
.Y(n_161)
);

INVxp67_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_131),
.A2(n_132),
.B1(n_134),
.B2(n_135),
.Y(n_130)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_SL g151 ( 
.A(n_132),
.B(n_134),
.Y(n_151)
);

CKINVDCx16_ASAP7_75t_R g134 ( 
.A(n_135),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_SL g138 ( 
.A1(n_139),
.A2(n_143),
.B(n_148),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_142),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_140),
.B(n_142),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_144),
.B(n_146),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_152),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_151),
.B(n_152),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_160),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_154),
.A2(n_155),
.B1(n_157),
.B2(n_158),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_154),
.B(n_158),
.C(n_160),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_155),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_158),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_165),
.B(n_166),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_165),
.B(n_166),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_167),
.A2(n_172),
.B1(n_179),
.B2(n_180),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_167),
.Y(n_179)
);

XOR2xp5_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_169),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_168),
.B(n_169),
.Y(n_191)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_172),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_173),
.A2(n_175),
.B1(n_176),
.B2(n_178),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_173),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_175),
.B(n_178),
.C(n_179),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_176),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_184),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_183),
.B(n_184),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_185),
.A2(n_186),
.B1(n_189),
.B2(n_190),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_185),
.B(n_191),
.C(n_192),
.Y(n_196)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

XOR2xp5_ASAP7_75t_L g190 ( 
.A(n_191),
.B(n_192),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_197),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_SL g200 ( 
.A(n_196),
.B(n_197),
.Y(n_200)
);


endmodule