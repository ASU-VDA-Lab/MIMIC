module fake_jpeg_28091_n_270 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_270);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_270;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_223;
wire n_187;
wire n_21;
wire n_57;
wire n_234;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_96;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_14),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_0),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_15),
.B(n_7),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_1),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

BUFx2_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

INVx6_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_0),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_3),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

BUFx16f_ASAP7_75t_L g35 ( 
.A(n_10),
.Y(n_35)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_21),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_36),
.Y(n_56)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_18),
.Y(n_37)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_37),
.Y(n_63)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_21),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_38),
.Y(n_51)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_26),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_39),
.Y(n_69)
);

INVx13_ASAP7_75t_L g40 ( 
.A(n_35),
.Y(n_40)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_40),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_23),
.B(n_9),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_SL g48 ( 
.A(n_41),
.B(n_23),
.Y(n_48)
);

INVx13_ASAP7_75t_L g42 ( 
.A(n_35),
.Y(n_42)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_42),
.Y(n_53)
);

HB1xp67_ASAP7_75t_L g43 ( 
.A(n_26),
.Y(n_43)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_43),
.Y(n_60)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_35),
.Y(n_44)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_44),
.Y(n_65)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_18),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_45),
.Y(n_70)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_21),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_46),
.B(n_21),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_18),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_47),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_SL g90 ( 
.A(n_48),
.B(n_62),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_L g49 ( 
.A1(n_36),
.A2(n_28),
.B1(n_27),
.B2(n_33),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_49),
.A2(n_76),
.B1(n_20),
.B2(n_19),
.Y(n_95)
);

OAI22xp33_ASAP7_75t_L g52 ( 
.A1(n_46),
.A2(n_28),
.B1(n_27),
.B2(n_31),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_52),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_SL g54 ( 
.A1(n_38),
.A2(n_28),
.B1(n_17),
.B2(n_33),
.Y(n_54)
);

OAI21xp5_ASAP7_75t_SL g89 ( 
.A1(n_54),
.A2(n_34),
.B(n_25),
.Y(n_89)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_57),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_41),
.B(n_17),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_58),
.B(n_67),
.Y(n_92)
);

AND2x2_ASAP7_75t_SL g59 ( 
.A(n_47),
.B(n_29),
.Y(n_59)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_59),
.B(n_31),
.C(n_29),
.Y(n_91)
);

AND2x2_ASAP7_75t_L g61 ( 
.A(n_37),
.B(n_31),
.Y(n_61)
);

A2O1A1Ixp33_ASAP7_75t_L g99 ( 
.A1(n_61),
.A2(n_0),
.B(n_1),
.C(n_2),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_43),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_45),
.B(n_30),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_64),
.B(n_72),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_SL g66 ( 
.A(n_40),
.B(n_17),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_66),
.B(n_71),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_40),
.B(n_24),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_42),
.B(n_24),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_68),
.B(n_73),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_42),
.B(n_25),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_47),
.B(n_30),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_44),
.B(n_32),
.Y(n_73)
);

BUFx12f_ASAP7_75t_L g74 ( 
.A(n_39),
.Y(n_74)
);

INVx5_ASAP7_75t_L g93 ( 
.A(n_74),
.Y(n_93)
);

BUFx12f_ASAP7_75t_L g75 ( 
.A(n_39),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_75),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_38),
.A2(n_28),
.B1(n_27),
.B2(n_32),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_L g78 ( 
.A1(n_72),
.A2(n_44),
.B1(n_26),
.B2(n_29),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_78),
.A2(n_97),
.B1(n_65),
.B2(n_56),
.Y(n_128)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_69),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_79),
.Y(n_115)
);

OA22x2_ASAP7_75t_L g80 ( 
.A1(n_59),
.A2(n_26),
.B1(n_35),
.B2(n_22),
.Y(n_80)
);

AO21x1_ASAP7_75t_L g129 ( 
.A1(n_80),
.A2(n_84),
.B(n_85),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_59),
.A2(n_30),
.B1(n_34),
.B2(n_20),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_81),
.A2(n_95),
.B1(n_96),
.B2(n_106),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_55),
.Y(n_82)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_82),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_62),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_83),
.B(n_86),
.Y(n_113)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_64),
.Y(n_84)
);

NOR2x1_ASAP7_75t_SL g85 ( 
.A(n_61),
.B(n_35),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_66),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_48),
.B(n_22),
.Y(n_88)
);

NOR3xp33_ASAP7_75t_SL g137 ( 
.A(n_88),
.B(n_6),
.C(n_8),
.Y(n_137)
);

CKINVDCx16_ASAP7_75t_R g132 ( 
.A(n_89),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_91),
.B(n_101),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_50),
.A2(n_25),
.B1(n_34),
.B2(n_20),
.Y(n_94)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_94),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_54),
.A2(n_19),
.B1(n_31),
.B2(n_29),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_L g97 ( 
.A1(n_63),
.A2(n_19),
.B1(n_9),
.B2(n_10),
.Y(n_97)
);

OAI32xp33_ASAP7_75t_L g98 ( 
.A1(n_61),
.A2(n_9),
.A3(n_15),
.B1(n_14),
.B2(n_3),
.Y(n_98)
);

NAND3xp33_ASAP7_75t_L g130 ( 
.A(n_98),
.B(n_6),
.C(n_7),
.Y(n_130)
);

NOR2x1_ASAP7_75t_L g119 ( 
.A(n_99),
.B(n_4),
.Y(n_119)
);

XNOR2xp5_ASAP7_75t_L g101 ( 
.A(n_60),
.B(n_10),
.Y(n_101)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_63),
.Y(n_102)
);

BUFx3_ASAP7_75t_L g134 ( 
.A(n_102),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_55),
.Y(n_104)
);

BUFx12f_ASAP7_75t_L g111 ( 
.A(n_104),
.Y(n_111)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_70),
.Y(n_105)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_105),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_55),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_107),
.Y(n_124)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_70),
.Y(n_108)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_108),
.Y(n_127)
);

AND2x2_ASAP7_75t_SL g109 ( 
.A(n_60),
.B(n_2),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_109),
.B(n_2),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_100),
.B(n_50),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_116),
.B(n_121),
.Y(n_160)
);

AND2x2_ASAP7_75t_L g150 ( 
.A(n_117),
.B(n_80),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_103),
.B(n_55),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_118),
.B(n_119),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_84),
.A2(n_52),
.B1(n_65),
.B2(n_56),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_120),
.A2(n_128),
.B1(n_81),
.B2(n_106),
.Y(n_141)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_89),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_92),
.B(n_53),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_122),
.B(n_123),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_90),
.B(n_53),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_130),
.B(n_8),
.Y(n_152)
);

NOR2x1_ASAP7_75t_L g131 ( 
.A(n_85),
.B(n_6),
.Y(n_131)
);

INVxp67_ASAP7_75t_L g164 ( 
.A(n_131),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_103),
.B(n_51),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_133),
.B(n_109),
.Y(n_151)
);

BUFx2_ASAP7_75t_L g136 ( 
.A(n_82),
.Y(n_136)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_136),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_SL g148 ( 
.A(n_137),
.B(n_101),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_124),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_138),
.Y(n_169)
);

CKINVDCx16_ASAP7_75t_R g140 ( 
.A(n_113),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_140),
.B(n_149),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_141),
.A2(n_134),
.B1(n_137),
.B2(n_75),
.Y(n_187)
);

AOI21xp5_ASAP7_75t_L g142 ( 
.A1(n_112),
.A2(n_99),
.B(n_86),
.Y(n_142)
);

AOI21xp5_ASAP7_75t_L g188 ( 
.A1(n_142),
.A2(n_156),
.B(n_150),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_112),
.A2(n_98),
.B1(n_77),
.B2(n_83),
.Y(n_143)
);

INVxp67_ASAP7_75t_L g173 ( 
.A(n_143),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_132),
.A2(n_77),
.B1(n_91),
.B2(n_90),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_144),
.A2(n_146),
.B1(n_165),
.B2(n_126),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_121),
.A2(n_109),
.B1(n_87),
.B2(n_80),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_148),
.B(n_152),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_124),
.B(n_108),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_150),
.B(n_151),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_135),
.A2(n_79),
.B1(n_102),
.B2(n_105),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_153),
.A2(n_154),
.B1(n_120),
.B2(n_156),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_135),
.A2(n_80),
.B1(n_93),
.B2(n_51),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_136),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_155),
.Y(n_180)
);

AND2x2_ASAP7_75t_L g156 ( 
.A(n_117),
.B(n_51),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_136),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_157),
.B(n_158),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_115),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_115),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_159),
.B(n_161),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_115),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_111),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_162),
.B(n_110),
.Y(n_190)
);

BUFx5_ASAP7_75t_L g163 ( 
.A(n_111),
.Y(n_163)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_163),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_128),
.A2(n_93),
.B1(n_69),
.B2(n_75),
.Y(n_165)
);

AOI322xp5_ASAP7_75t_L g168 ( 
.A1(n_154),
.A2(n_114),
.A3(n_129),
.B1(n_131),
.B2(n_133),
.C1(n_118),
.C2(n_119),
.Y(n_168)
);

AOI221xp5_ASAP7_75t_L g201 ( 
.A1(n_168),
.A2(n_164),
.B1(n_152),
.B2(n_161),
.C(n_159),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_170),
.A2(n_179),
.B1(n_187),
.B2(n_189),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g175 ( 
.A(n_144),
.B(n_114),
.Y(n_175)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_175),
.B(n_156),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_151),
.B(n_129),
.C(n_127),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_176),
.B(n_178),
.C(n_183),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_L g177 ( 
.A(n_146),
.B(n_129),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_177),
.B(n_188),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_160),
.B(n_127),
.C(n_125),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_153),
.A2(n_125),
.B1(n_126),
.B2(n_69),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_147),
.B(n_134),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_182),
.B(n_140),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_160),
.B(n_110),
.C(n_75),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_184),
.B(n_165),
.Y(n_197)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_138),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_185),
.B(n_186),
.Y(n_204)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_145),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_141),
.A2(n_74),
.B1(n_107),
.B2(n_104),
.Y(n_189)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_190),
.Y(n_206)
);

AOI22xp33_ASAP7_75t_SL g192 ( 
.A1(n_180),
.A2(n_157),
.B1(n_155),
.B2(n_158),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_192),
.A2(n_180),
.B1(n_183),
.B2(n_190),
.Y(n_213)
);

OAI32xp33_ASAP7_75t_L g194 ( 
.A1(n_174),
.A2(n_147),
.A3(n_150),
.B1(n_143),
.B2(n_142),
.Y(n_194)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_194),
.Y(n_215)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_196),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_197),
.B(n_198),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_SL g198 ( 
.A(n_166),
.B(n_148),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_SL g222 ( 
.A(n_199),
.B(n_172),
.Y(n_222)
);

INVx2_ASAP7_75t_SL g200 ( 
.A(n_169),
.Y(n_200)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_200),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_201),
.B(n_203),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_182),
.B(n_139),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_202),
.Y(n_212)
);

AOI21xp5_ASAP7_75t_L g203 ( 
.A1(n_169),
.A2(n_162),
.B(n_139),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_175),
.B(n_74),
.C(n_111),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_205),
.B(n_178),
.C(n_176),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_181),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_207),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_166),
.B(n_163),
.Y(n_208)
);

NAND3xp33_ASAP7_75t_L g214 ( 
.A(n_208),
.B(n_210),
.C(n_174),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_185),
.B(n_74),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_209),
.B(n_171),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_181),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_213),
.A2(n_219),
.B1(n_206),
.B2(n_200),
.Y(n_233)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_214),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_195),
.A2(n_184),
.B1(n_189),
.B2(n_173),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_216),
.A2(n_223),
.B1(n_202),
.B2(n_196),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_218),
.B(n_220),
.C(n_193),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_207),
.A2(n_170),
.B1(n_173),
.B2(n_179),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_191),
.B(n_188),
.C(n_177),
.Y(n_220)
);

MAJx2_ASAP7_75t_L g230 ( 
.A(n_222),
.B(n_205),
.C(n_199),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_195),
.A2(n_187),
.B1(n_186),
.B2(n_167),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_226),
.B(n_191),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_SL g245 ( 
.A(n_227),
.B(n_229),
.Y(n_245)
);

AOI31xp67_ASAP7_75t_L g228 ( 
.A1(n_225),
.A2(n_194),
.A3(n_210),
.B(n_206),
.Y(n_228)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_228),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_230),
.B(n_231),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_226),
.B(n_204),
.Y(n_232)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_232),
.Y(n_248)
);

AND2x2_ASAP7_75t_L g244 ( 
.A(n_233),
.B(n_236),
.Y(n_244)
);

AOI321xp33_ASAP7_75t_L g234 ( 
.A1(n_215),
.A2(n_193),
.A3(n_198),
.B1(n_204),
.B2(n_200),
.C(n_203),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_SL g242 ( 
.A(n_234),
.B(n_235),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_223),
.B(n_171),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_SL g236 ( 
.A(n_224),
.B(n_209),
.Y(n_236)
);

AOI21xp5_ASAP7_75t_L g237 ( 
.A1(n_213),
.A2(n_8),
.B(n_11),
.Y(n_237)
);

O2A1O1Ixp33_ASAP7_75t_L g240 ( 
.A1(n_237),
.A2(n_238),
.B(n_215),
.C(n_13),
.Y(n_240)
);

AOI31xp67_ASAP7_75t_L g238 ( 
.A1(n_212),
.A2(n_12),
.A3(n_13),
.B(n_15),
.Y(n_238)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_240),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_231),
.B(n_218),
.C(n_220),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_241),
.B(n_247),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_230),
.B(n_222),
.C(n_221),
.Y(n_247)
);

O2A1O1Ixp33_ASAP7_75t_L g249 ( 
.A1(n_228),
.A2(n_211),
.B(n_219),
.C(n_217),
.Y(n_249)
);

AOI21xp5_ASAP7_75t_L g252 ( 
.A1(n_249),
.A2(n_227),
.B(n_216),
.Y(n_252)
);

OAI221xp5_ASAP7_75t_L g250 ( 
.A1(n_245),
.A2(n_239),
.B1(n_234),
.B2(n_233),
.C(n_238),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_250),
.B(n_246),
.Y(n_260)
);

NOR2xp67_ASAP7_75t_SL g251 ( 
.A(n_243),
.B(n_221),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_SL g257 ( 
.A(n_251),
.B(n_256),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_252),
.B(n_253),
.Y(n_259)
);

CKINVDCx16_ASAP7_75t_R g253 ( 
.A(n_244),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_SL g256 ( 
.A(n_248),
.B(n_12),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_SL g258 ( 
.A(n_255),
.B(n_244),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_SL g262 ( 
.A(n_258),
.B(n_261),
.Y(n_262)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_260),
.Y(n_264)
);

AOI22xp33_ASAP7_75t_L g261 ( 
.A1(n_252),
.A2(n_249),
.B1(n_240),
.B2(n_242),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_257),
.B(n_254),
.C(n_241),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_SL g266 ( 
.A(n_263),
.B(n_265),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_259),
.B(n_247),
.C(n_111),
.Y(n_265)
);

OAI21x1_ASAP7_75t_L g267 ( 
.A1(n_262),
.A2(n_261),
.B(n_13),
.Y(n_267)
);

AOI21xp5_ASAP7_75t_SL g268 ( 
.A1(n_267),
.A2(n_264),
.B(n_16),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_268),
.B(n_266),
.C(n_16),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_269),
.B(n_16),
.Y(n_270)
);


endmodule