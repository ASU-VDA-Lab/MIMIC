module real_aes_7679_n_103 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_103);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_103;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_503;
wire n_357;
wire n_287;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_742;
wire n_112;
wire n_364;
wire n_319;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_537;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_693;
wire n_496;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_755;
wire n_153;
wire n_316;
wire n_532;
wire n_284;
wire n_656;
wire n_178;
wire n_409;
wire n_748;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_504;
wire n_310;
wire n_455;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_449;
wire n_363;
wire n_754;
wire n_417;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_505;
wire n_527;
wire n_434;
wire n_502;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_542;
wire n_163;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_756;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_749;
wire n_358;
wire n_275;
wire n_214;
wire n_385;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_679;
wire n_520;
wire n_633;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_753;
wire n_741;
wire n_283;
wire n_314;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_456;
wire n_359;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_524;
wire n_219;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_479;
wire n_338;
wire n_442;
wire n_740;
wire n_371;
wire n_698;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
NAND3xp33_ASAP7_75t_SL g111 ( .A(n_0), .B(n_112), .C(n_113), .Y(n_111) );
INVx1_ASAP7_75t_L g128 ( .A(n_0), .Y(n_128) );
INVx1_ASAP7_75t_L g496 ( .A(n_1), .Y(n_496) );
INVx1_ASAP7_75t_L g275 ( .A(n_2), .Y(n_275) );
AOI22xp33_ASAP7_75t_L g523 ( .A1(n_3), .A2(n_36), .B1(n_194), .B2(n_524), .Y(n_523) );
AOI21xp33_ASAP7_75t_L g182 ( .A1(n_4), .A2(n_183), .B(n_184), .Y(n_182) );
NAND2xp5_ASAP7_75t_L g473 ( .A(n_5), .B(n_181), .Y(n_473) );
AND2x6_ASAP7_75t_L g156 ( .A(n_6), .B(n_157), .Y(n_156) );
AOI21xp5_ASAP7_75t_L g250 ( .A1(n_7), .A2(n_251), .B(n_252), .Y(n_250) );
INVx1_ASAP7_75t_L g109 ( .A(n_8), .Y(n_109) );
NOR2xp33_ASAP7_75t_L g129 ( .A(n_8), .B(n_37), .Y(n_129) );
INVx1_ASAP7_75t_L g191 ( .A(n_9), .Y(n_191) );
NAND2xp5_ASAP7_75t_L g242 ( .A(n_10), .B(n_243), .Y(n_242) );
INVx1_ASAP7_75t_L g153 ( .A(n_11), .Y(n_153) );
INVx1_ASAP7_75t_L g492 ( .A(n_12), .Y(n_492) );
INVx1_ASAP7_75t_L g257 ( .A(n_13), .Y(n_257) );
NAND2xp5_ASAP7_75t_L g530 ( .A(n_14), .B(n_159), .Y(n_530) );
NAND2xp5_ASAP7_75t_L g501 ( .A(n_15), .B(n_149), .Y(n_501) );
AO32x2_ASAP7_75t_L g521 ( .A1(n_16), .A2(n_148), .A3(n_181), .B1(n_484), .B2(n_522), .Y(n_521) );
NAND2xp5_ASAP7_75t_SL g533 ( .A(n_17), .B(n_194), .Y(n_533) );
NAND2xp5_ASAP7_75t_L g229 ( .A(n_18), .B(n_202), .Y(n_229) );
NAND2xp5_ASAP7_75t_L g498 ( .A(n_19), .B(n_149), .Y(n_498) );
AOI22xp33_ASAP7_75t_L g525 ( .A1(n_20), .A2(n_50), .B1(n_194), .B2(n_524), .Y(n_525) );
NAND2xp5_ASAP7_75t_SL g211 ( .A(n_21), .B(n_183), .Y(n_211) );
AOI22xp33_ASAP7_75t_SL g544 ( .A1(n_22), .A2(n_76), .B1(n_159), .B2(n_194), .Y(n_544) );
NAND2xp5_ASAP7_75t_SL g516 ( .A(n_23), .B(n_194), .Y(n_516) );
NAND2xp5_ASAP7_75t_L g205 ( .A(n_24), .B(n_179), .Y(n_205) );
A2O1A1Ixp33_ASAP7_75t_L g254 ( .A1(n_25), .A2(n_255), .B(n_256), .C(n_258), .Y(n_254) );
BUFx6f_ASAP7_75t_L g164 ( .A(n_26), .Y(n_164) );
NAND2xp5_ASAP7_75t_L g485 ( .A(n_27), .B(n_196), .Y(n_485) );
NAND2xp5_ASAP7_75t_L g276 ( .A(n_28), .B(n_189), .Y(n_276) );
INVx1_ASAP7_75t_L g167 ( .A(n_29), .Y(n_167) );
NAND2xp5_ASAP7_75t_L g518 ( .A(n_30), .B(n_196), .Y(n_518) );
INVx2_ASAP7_75t_L g161 ( .A(n_31), .Y(n_161) );
NAND2xp5_ASAP7_75t_SL g478 ( .A(n_32), .B(n_194), .Y(n_478) );
NAND2xp5_ASAP7_75t_L g535 ( .A(n_33), .B(n_196), .Y(n_535) );
AOI22xp5_ASAP7_75t_L g751 ( .A1(n_34), .A2(n_42), .B1(n_752), .B2(n_753), .Y(n_751) );
CKINVDCx20_ASAP7_75t_R g753 ( .A(n_34), .Y(n_753) );
A2O1A1Ixp33_ASAP7_75t_L g212 ( .A1(n_35), .A2(n_156), .B(n_168), .C(n_213), .Y(n_212) );
NAND2xp5_ASAP7_75t_L g108 ( .A(n_37), .B(n_109), .Y(n_108) );
INVx1_ASAP7_75t_L g165 ( .A(n_38), .Y(n_165) );
CKINVDCx20_ASAP7_75t_R g130 ( .A(n_39), .Y(n_130) );
AOI22xp33_ASAP7_75t_L g103 ( .A1(n_40), .A2(n_104), .B1(n_116), .B2(n_756), .Y(n_103) );
NAND2xp5_ASAP7_75t_SL g228 ( .A(n_41), .B(n_189), .Y(n_228) );
CKINVDCx20_ASAP7_75t_R g752 ( .A(n_42), .Y(n_752) );
NAND2xp5_ASAP7_75t_SL g466 ( .A(n_43), .B(n_194), .Y(n_466) );
AOI22xp33_ASAP7_75t_L g543 ( .A1(n_44), .A2(n_87), .B1(n_219), .B2(n_524), .Y(n_543) );
NAND2xp5_ASAP7_75t_SL g469 ( .A(n_45), .B(n_194), .Y(n_469) );
NAND2xp5_ASAP7_75t_L g493 ( .A(n_46), .B(n_194), .Y(n_493) );
CKINVDCx16_ASAP7_75t_R g171 ( .A(n_47), .Y(n_171) );
NAND2xp5_ASAP7_75t_L g470 ( .A(n_48), .B(n_471), .Y(n_470) );
NAND2xp5_ASAP7_75t_L g245 ( .A(n_49), .B(n_183), .Y(n_245) );
AOI22xp33_ASAP7_75t_SL g505 ( .A1(n_51), .A2(n_60), .B1(n_159), .B2(n_194), .Y(n_505) );
AOI22xp5_ASAP7_75t_L g158 ( .A1(n_52), .A2(n_159), .B1(n_162), .B2(n_168), .Y(n_158) );
CKINVDCx20_ASAP7_75t_R g222 ( .A(n_53), .Y(n_222) );
NAND2xp5_ASAP7_75t_SL g483 ( .A(n_54), .B(n_194), .Y(n_483) );
CKINVDCx16_ASAP7_75t_R g272 ( .A(n_55), .Y(n_272) );
NAND2xp5_ASAP7_75t_SL g529 ( .A(n_56), .B(n_194), .Y(n_529) );
A2O1A1Ixp33_ASAP7_75t_L g187 ( .A1(n_57), .A2(n_188), .B(n_190), .C(n_193), .Y(n_187) );
CKINVDCx20_ASAP7_75t_R g232 ( .A(n_58), .Y(n_232) );
INVx1_ASAP7_75t_L g185 ( .A(n_59), .Y(n_185) );
INVx1_ASAP7_75t_L g157 ( .A(n_61), .Y(n_157) );
NAND2xp5_ASAP7_75t_L g497 ( .A(n_62), .B(n_194), .Y(n_497) );
INVx1_ASAP7_75t_L g152 ( .A(n_63), .Y(n_152) );
CKINVDCx20_ASAP7_75t_R g122 ( .A(n_64), .Y(n_122) );
AO32x2_ASAP7_75t_L g541 ( .A1(n_65), .A2(n_181), .A3(n_237), .B1(n_484), .B2(n_542), .Y(n_541) );
INVx1_ASAP7_75t_L g481 ( .A(n_66), .Y(n_481) );
INVx1_ASAP7_75t_L g513 ( .A(n_67), .Y(n_513) );
OAI22xp5_ASAP7_75t_SL g749 ( .A1(n_68), .A2(n_750), .B1(n_751), .B2(n_754), .Y(n_749) );
CKINVDCx20_ASAP7_75t_R g754 ( .A(n_68), .Y(n_754) );
A2O1A1Ixp33_ASAP7_75t_SL g201 ( .A1(n_69), .A2(n_193), .B(n_202), .C(n_203), .Y(n_201) );
INVxp67_ASAP7_75t_L g204 ( .A(n_70), .Y(n_204) );
NAND2xp5_ASAP7_75t_SL g514 ( .A(n_71), .B(n_159), .Y(n_514) );
INVx1_ASAP7_75t_L g115 ( .A(n_72), .Y(n_115) );
CKINVDCx20_ASAP7_75t_R g176 ( .A(n_73), .Y(n_176) );
INVx1_ASAP7_75t_L g225 ( .A(n_74), .Y(n_225) );
OAI22xp5_ASAP7_75t_L g136 ( .A1(n_75), .A2(n_101), .B1(n_137), .B2(n_138), .Y(n_136) );
CKINVDCx20_ASAP7_75t_R g137 ( .A(n_75), .Y(n_137) );
A2O1A1Ixp33_ASAP7_75t_L g226 ( .A1(n_77), .A2(n_156), .B(n_168), .C(n_227), .Y(n_226) );
NAND2xp5_ASAP7_75t_L g534 ( .A(n_78), .B(n_524), .Y(n_534) );
NAND2xp5_ASAP7_75t_SL g517 ( .A(n_79), .B(n_159), .Y(n_517) );
AOI222xp33_ASAP7_75t_SL g131 ( .A1(n_80), .A2(n_132), .B1(n_133), .B2(n_139), .C1(n_739), .C2(n_742), .Y(n_131) );
NAND2xp5_ASAP7_75t_SL g214 ( .A(n_81), .B(n_215), .Y(n_214) );
INVx2_ASAP7_75t_L g150 ( .A(n_82), .Y(n_150) );
NAND2xp5_ASAP7_75t_L g216 ( .A(n_83), .B(n_202), .Y(n_216) );
NAND2xp5_ASAP7_75t_L g467 ( .A(n_84), .B(n_159), .Y(n_467) );
A2O1A1Ixp33_ASAP7_75t_L g273 ( .A1(n_85), .A2(n_156), .B(n_168), .C(n_274), .Y(n_273) );
INVx2_ASAP7_75t_L g112 ( .A(n_86), .Y(n_112) );
OR2x2_ASAP7_75t_L g125 ( .A(n_86), .B(n_126), .Y(n_125) );
OR2x2_ASAP7_75t_L g455 ( .A(n_86), .B(n_127), .Y(n_455) );
AOI22xp33_ASAP7_75t_L g504 ( .A1(n_88), .A2(n_102), .B1(n_159), .B2(n_160), .Y(n_504) );
NAND2xp5_ASAP7_75t_L g195 ( .A(n_89), .B(n_196), .Y(n_195) );
CKINVDCx20_ASAP7_75t_R g279 ( .A(n_90), .Y(n_279) );
A2O1A1Ixp33_ASAP7_75t_L g239 ( .A1(n_91), .A2(n_156), .B(n_168), .C(n_240), .Y(n_239) );
CKINVDCx20_ASAP7_75t_R g247 ( .A(n_92), .Y(n_247) );
INVx1_ASAP7_75t_L g200 ( .A(n_93), .Y(n_200) );
CKINVDCx16_ASAP7_75t_R g253 ( .A(n_94), .Y(n_253) );
NAND2xp5_ASAP7_75t_SL g241 ( .A(n_95), .B(n_215), .Y(n_241) );
AOI22xp5_ASAP7_75t_L g133 ( .A1(n_96), .A2(n_134), .B1(n_135), .B2(n_136), .Y(n_133) );
CKINVDCx20_ASAP7_75t_R g134 ( .A(n_96), .Y(n_134) );
NAND2xp5_ASAP7_75t_L g479 ( .A(n_97), .B(n_159), .Y(n_479) );
NAND2xp5_ASAP7_75t_L g259 ( .A(n_98), .B(n_181), .Y(n_259) );
NAND2xp5_ASAP7_75t_L g114 ( .A(n_99), .B(n_115), .Y(n_114) );
AOI21xp5_ASAP7_75t_L g198 ( .A1(n_100), .A2(n_183), .B(n_199), .Y(n_198) );
CKINVDCx16_ASAP7_75t_R g138 ( .A(n_101), .Y(n_138) );
INVx1_ASAP7_75t_L g104 ( .A(n_105), .Y(n_104) );
INVx2_ASAP7_75t_L g105 ( .A(n_106), .Y(n_105) );
INVx2_ASAP7_75t_SL g756 ( .A(n_106), .Y(n_756) );
AND2x2_ASAP7_75t_L g106 ( .A(n_107), .B(n_110), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_108), .Y(n_107) );
INVx1_ASAP7_75t_L g110 ( .A(n_111), .Y(n_110) );
OR2x2_ASAP7_75t_L g738 ( .A(n_112), .B(n_127), .Y(n_738) );
NOR2x2_ASAP7_75t_L g744 ( .A(n_112), .B(n_126), .Y(n_744) );
INVx1_ASAP7_75t_SL g113 ( .A(n_114), .Y(n_113) );
BUFx2_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
AOI22xp5_ASAP7_75t_L g117 ( .A1(n_118), .A2(n_131), .B1(n_745), .B2(n_746), .Y(n_117) );
NOR2xp33_ASAP7_75t_L g118 ( .A(n_119), .B(n_123), .Y(n_118) );
INVx1_ASAP7_75t_SL g119 ( .A(n_120), .Y(n_119) );
INVx1_ASAP7_75t_SL g745 ( .A(n_120), .Y(n_745) );
BUFx2_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
INVx2_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
AOI21xp5_ASAP7_75t_L g746 ( .A1(n_123), .A2(n_747), .B(n_755), .Y(n_746) );
NOR2xp33_ASAP7_75t_SL g123 ( .A(n_124), .B(n_130), .Y(n_123) );
BUFx2_ASAP7_75t_L g124 ( .A(n_125), .Y(n_124) );
HB1xp67_ASAP7_75t_L g755 ( .A(n_125), .Y(n_755) );
INVx2_ASAP7_75t_L g126 ( .A(n_127), .Y(n_126) );
AND2x2_ASAP7_75t_L g127 ( .A(n_128), .B(n_129), .Y(n_127) );
INVx1_ASAP7_75t_L g132 ( .A(n_133), .Y(n_132) );
CKINVDCx14_ASAP7_75t_R g135 ( .A(n_136), .Y(n_135) );
OAI22xp5_ASAP7_75t_SL g139 ( .A1(n_140), .A2(n_453), .B1(n_456), .B2(n_736), .Y(n_139) );
OAI22xp5_ASAP7_75t_L g747 ( .A1(n_140), .A2(n_141), .B1(n_748), .B2(n_749), .Y(n_747) );
INVx1_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
OAI22xp5_ASAP7_75t_SL g739 ( .A1(n_141), .A2(n_453), .B1(n_740), .B2(n_741), .Y(n_739) );
AND3x1_ASAP7_75t_L g141 ( .A(n_142), .B(n_378), .C(n_427), .Y(n_141) );
NOR3xp33_ASAP7_75t_SL g142 ( .A(n_143), .B(n_285), .C(n_323), .Y(n_142) );
OAI222xp33_ASAP7_75t_L g143 ( .A1(n_144), .A2(n_206), .B1(n_260), .B2(n_266), .C1(n_280), .C2(n_283), .Y(n_143) );
NAND2xp5_ASAP7_75t_L g144 ( .A(n_145), .B(n_177), .Y(n_144) );
NAND2xp5_ASAP7_75t_L g352 ( .A(n_145), .B(n_353), .Y(n_352) );
NAND2xp5_ASAP7_75t_L g419 ( .A(n_145), .B(n_328), .Y(n_419) );
BUFx2_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
OR2x2_ASAP7_75t_L g296 ( .A(n_146), .B(n_197), .Y(n_296) );
NAND2xp5_ASAP7_75t_L g304 ( .A(n_146), .B(n_178), .Y(n_304) );
AND2x2_ASAP7_75t_L g339 ( .A(n_146), .B(n_316), .Y(n_339) );
OR2x2_ASAP7_75t_L g363 ( .A(n_146), .B(n_178), .Y(n_363) );
OR2x2_ASAP7_75t_L g371 ( .A(n_146), .B(n_270), .Y(n_371) );
AND2x2_ASAP7_75t_L g374 ( .A(n_146), .B(n_197), .Y(n_374) );
INVx3_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
OR2x2_ASAP7_75t_L g268 ( .A(n_147), .B(n_269), .Y(n_268) );
AND2x2_ASAP7_75t_L g282 ( .A(n_147), .B(n_197), .Y(n_282) );
AND2x2_ASAP7_75t_L g332 ( .A(n_147), .B(n_270), .Y(n_332) );
AND2x2_ASAP7_75t_L g345 ( .A(n_147), .B(n_178), .Y(n_345) );
NOR2xp33_ASAP7_75t_L g452 ( .A(n_147), .B(n_431), .Y(n_452) );
AO21x2_ASAP7_75t_L g147 ( .A1(n_148), .A2(n_154), .B(n_175), .Y(n_147) );
NOR2xp33_ASAP7_75t_L g175 ( .A(n_148), .B(n_176), .Y(n_175) );
INVx2_ASAP7_75t_L g220 ( .A(n_148), .Y(n_220) );
AO21x2_ASAP7_75t_L g270 ( .A1(n_148), .A2(n_271), .B(n_278), .Y(n_270) );
INVx1_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
BUFx6f_ASAP7_75t_L g181 ( .A(n_149), .Y(n_181) );
AND2x2_ASAP7_75t_L g149 ( .A(n_150), .B(n_151), .Y(n_149) );
AND2x2_ASAP7_75t_SL g196 ( .A(n_150), .B(n_151), .Y(n_196) );
NAND2xp5_ASAP7_75t_L g151 ( .A(n_152), .B(n_153), .Y(n_151) );
OAI22xp33_ASAP7_75t_L g154 ( .A1(n_155), .A2(n_158), .B1(n_171), .B2(n_172), .Y(n_154) );
O2A1O1Ixp33_ASAP7_75t_L g184 ( .A1(n_155), .A2(n_185), .B(n_186), .C(n_187), .Y(n_184) );
O2A1O1Ixp33_ASAP7_75t_L g199 ( .A1(n_155), .A2(n_186), .B(n_200), .C(n_201), .Y(n_199) );
O2A1O1Ixp33_ASAP7_75t_L g252 ( .A1(n_155), .A2(n_186), .B(n_253), .C(n_254), .Y(n_252) );
INVx4_ASAP7_75t_SL g155 ( .A(n_156), .Y(n_155) );
NAND2x1p5_ASAP7_75t_L g172 ( .A(n_156), .B(n_173), .Y(n_172) );
AND2x4_ASAP7_75t_L g183 ( .A(n_156), .B(n_173), .Y(n_183) );
OAI21xp5_ASAP7_75t_L g464 ( .A1(n_156), .A2(n_465), .B(n_468), .Y(n_464) );
BUFx3_ASAP7_75t_L g484 ( .A(n_156), .Y(n_484) );
OAI21xp5_ASAP7_75t_L g490 ( .A1(n_156), .A2(n_491), .B(n_495), .Y(n_490) );
OAI21xp5_ASAP7_75t_L g511 ( .A1(n_156), .A2(n_512), .B(n_515), .Y(n_511) );
OAI21xp5_ASAP7_75t_L g527 ( .A1(n_156), .A2(n_528), .B(n_532), .Y(n_527) );
INVx2_ASAP7_75t_L g277 ( .A(n_159), .Y(n_277) );
INVx3_ASAP7_75t_L g159 ( .A(n_160), .Y(n_159) );
INVx1_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
INVx2_ASAP7_75t_L g169 ( .A(n_161), .Y(n_169) );
INVx1_ASAP7_75t_L g174 ( .A(n_161), .Y(n_174) );
OAI22xp5_ASAP7_75t_SL g162 ( .A1(n_163), .A2(n_165), .B1(n_166), .B2(n_167), .Y(n_162) );
INVx2_ASAP7_75t_L g166 ( .A(n_163), .Y(n_166) );
INVx4_ASAP7_75t_L g255 ( .A(n_163), .Y(n_255) );
BUFx6f_ASAP7_75t_L g163 ( .A(n_164), .Y(n_163) );
INVx1_ASAP7_75t_L g170 ( .A(n_164), .Y(n_170) );
AND2x2_ASAP7_75t_L g173 ( .A(n_164), .B(n_174), .Y(n_173) );
BUFx6f_ASAP7_75t_L g189 ( .A(n_164), .Y(n_189) );
INVx3_ASAP7_75t_L g192 ( .A(n_164), .Y(n_192) );
INVx1_ASAP7_75t_L g202 ( .A(n_164), .Y(n_202) );
INVx5_ASAP7_75t_L g186 ( .A(n_168), .Y(n_186) );
AND2x6_ASAP7_75t_L g168 ( .A(n_169), .B(n_170), .Y(n_168) );
BUFx6f_ASAP7_75t_L g194 ( .A(n_169), .Y(n_194) );
BUFx3_ASAP7_75t_L g219 ( .A(n_169), .Y(n_219) );
INVx1_ASAP7_75t_L g524 ( .A(n_169), .Y(n_524) );
OAI21xp5_ASAP7_75t_L g224 ( .A1(n_172), .A2(n_225), .B(n_226), .Y(n_224) );
OAI21xp5_ASAP7_75t_L g271 ( .A1(n_172), .A2(n_272), .B(n_273), .Y(n_271) );
INVx1_ASAP7_75t_L g471 ( .A(n_174), .Y(n_471) );
O2A1O1Ixp33_ASAP7_75t_L g370 ( .A1(n_177), .A2(n_371), .B(n_372), .C(n_375), .Y(n_370) );
NAND2xp5_ASAP7_75t_L g399 ( .A(n_177), .B(n_400), .Y(n_399) );
NAND2xp5_ASAP7_75t_L g437 ( .A(n_177), .B(n_315), .Y(n_437) );
AND2x2_ASAP7_75t_L g177 ( .A(n_178), .B(n_197), .Y(n_177) );
AND2x2_ASAP7_75t_SL g281 ( .A(n_178), .B(n_282), .Y(n_281) );
INVx2_ASAP7_75t_L g295 ( .A(n_178), .Y(n_295) );
AND2x2_ASAP7_75t_L g322 ( .A(n_178), .B(n_316), .Y(n_322) );
INVx1_ASAP7_75t_SL g330 ( .A(n_178), .Y(n_330) );
AND2x2_ASAP7_75t_L g353 ( .A(n_178), .B(n_354), .Y(n_353) );
BUFx2_ASAP7_75t_L g431 ( .A(n_178), .Y(n_431) );
OA21x2_ASAP7_75t_L g178 ( .A1(n_179), .A2(n_182), .B(n_195), .Y(n_178) );
INVx3_ASAP7_75t_L g179 ( .A(n_180), .Y(n_179) );
NOR2xp33_ASAP7_75t_SL g221 ( .A(n_180), .B(n_222), .Y(n_221) );
NAND3xp33_ASAP7_75t_L g502 ( .A(n_180), .B(n_484), .C(n_503), .Y(n_502) );
AO21x1_ASAP7_75t_L g547 ( .A1(n_180), .A2(n_503), .B(n_548), .Y(n_547) );
INVx4_ASAP7_75t_L g180 ( .A(n_181), .Y(n_180) );
OA21x2_ASAP7_75t_L g197 ( .A1(n_181), .A2(n_198), .B(n_205), .Y(n_197) );
OA21x2_ASAP7_75t_L g463 ( .A1(n_181), .A2(n_464), .B(n_473), .Y(n_463) );
BUFx2_ASAP7_75t_L g251 ( .A(n_183), .Y(n_251) );
O2A1O1Ixp5_ASAP7_75t_L g480 ( .A1(n_188), .A2(n_481), .B(n_482), .C(n_483), .Y(n_480) );
AOI21xp5_ASAP7_75t_L g532 ( .A1(n_188), .A2(n_533), .B(n_534), .Y(n_532) );
INVx2_ASAP7_75t_L g188 ( .A(n_189), .Y(n_188) );
INVx4_ASAP7_75t_L g243 ( .A(n_189), .Y(n_243) );
OAI22xp5_ASAP7_75t_L g503 ( .A1(n_189), .A2(n_472), .B1(n_504), .B2(n_505), .Y(n_503) );
OAI22xp5_ASAP7_75t_L g522 ( .A1(n_189), .A2(n_472), .B1(n_523), .B2(n_525), .Y(n_522) );
OAI22xp5_ASAP7_75t_SL g542 ( .A1(n_189), .A2(n_192), .B1(n_543), .B2(n_544), .Y(n_542) );
NOR2xp33_ASAP7_75t_L g190 ( .A(n_191), .B(n_192), .Y(n_190) );
NOR2xp33_ASAP7_75t_L g203 ( .A(n_192), .B(n_204), .Y(n_203) );
INVx5_ASAP7_75t_L g215 ( .A(n_192), .Y(n_215) );
O2A1O1Ixp5_ASAP7_75t_SL g512 ( .A1(n_193), .A2(n_215), .B(n_513), .C(n_514), .Y(n_512) );
INVx3_ASAP7_75t_L g193 ( .A(n_194), .Y(n_193) );
HB1xp67_ASAP7_75t_L g244 ( .A(n_194), .Y(n_244) );
INVx1_ASAP7_75t_L g233 ( .A(n_196), .Y(n_233) );
INVx2_ASAP7_75t_L g237 ( .A(n_196), .Y(n_237) );
OA21x2_ASAP7_75t_L g249 ( .A1(n_196), .A2(n_250), .B(n_259), .Y(n_249) );
OA21x2_ASAP7_75t_L g510 ( .A1(n_196), .A2(n_511), .B(n_518), .Y(n_510) );
OA21x2_ASAP7_75t_L g526 ( .A1(n_196), .A2(n_527), .B(n_535), .Y(n_526) );
BUFx2_ASAP7_75t_L g267 ( .A(n_197), .Y(n_267) );
INVx1_ASAP7_75t_L g329 ( .A(n_197), .Y(n_329) );
INVx3_ASAP7_75t_L g354 ( .A(n_197), .Y(n_354) );
INVx1_ASAP7_75t_L g531 ( .A(n_202), .Y(n_531) );
NAND2xp5_ASAP7_75t_SL g287 ( .A(n_206), .B(n_288), .Y(n_287) );
OR2x2_ASAP7_75t_L g206 ( .A(n_207), .B(n_234), .Y(n_206) );
INVx1_ASAP7_75t_L g350 ( .A(n_207), .Y(n_350) );
OAI32xp33_ASAP7_75t_L g356 ( .A1(n_207), .A2(n_295), .A3(n_357), .B1(n_358), .B2(n_359), .Y(n_356) );
OAI22xp5_ASAP7_75t_L g360 ( .A1(n_207), .A2(n_361), .B1(n_364), .B2(n_369), .Y(n_360) );
INVx4_ASAP7_75t_L g207 ( .A(n_208), .Y(n_207) );
AND2x2_ASAP7_75t_L g298 ( .A(n_208), .B(n_299), .Y(n_298) );
AND2x2_ASAP7_75t_L g376 ( .A(n_208), .B(n_377), .Y(n_376) );
AND2x2_ASAP7_75t_L g446 ( .A(n_208), .B(n_392), .Y(n_446) );
AND2x2_ASAP7_75t_L g208 ( .A(n_209), .B(n_223), .Y(n_208) );
AND2x2_ASAP7_75t_L g261 ( .A(n_209), .B(n_262), .Y(n_261) );
INVx2_ASAP7_75t_L g291 ( .A(n_209), .Y(n_291) );
INVx1_ASAP7_75t_L g310 ( .A(n_209), .Y(n_310) );
OR2x2_ASAP7_75t_L g318 ( .A(n_209), .B(n_319), .Y(n_318) );
AND2x2_ASAP7_75t_L g325 ( .A(n_209), .B(n_299), .Y(n_325) );
NOR2xp33_ASAP7_75t_L g333 ( .A(n_209), .B(n_334), .Y(n_333) );
AND2x2_ASAP7_75t_L g346 ( .A(n_209), .B(n_264), .Y(n_346) );
INVx3_ASAP7_75t_L g368 ( .A(n_209), .Y(n_368) );
AND2x2_ASAP7_75t_L g393 ( .A(n_209), .B(n_265), .Y(n_393) );
NOR2xp33_ASAP7_75t_L g441 ( .A(n_209), .B(n_358), .Y(n_441) );
OR2x6_ASAP7_75t_L g209 ( .A(n_210), .B(n_221), .Y(n_209) );
AOI21xp5_ASAP7_75t_SL g210 ( .A1(n_211), .A2(n_212), .B(n_220), .Y(n_210) );
AOI21xp5_ASAP7_75t_L g213 ( .A1(n_214), .A2(n_216), .B(n_217), .Y(n_213) );
O2A1O1Ixp33_ASAP7_75t_L g274 ( .A1(n_215), .A2(n_275), .B(n_276), .C(n_277), .Y(n_274) );
AOI21xp5_ASAP7_75t_L g465 ( .A1(n_215), .A2(n_466), .B(n_467), .Y(n_465) );
INVx2_ASAP7_75t_L g472 ( .A(n_215), .Y(n_472) );
AOI21xp5_ASAP7_75t_L g477 ( .A1(n_215), .A2(n_478), .B(n_479), .Y(n_477) );
AOI21xp5_ASAP7_75t_L g227 ( .A1(n_217), .A2(n_228), .B(n_229), .Y(n_227) );
INVx2_ASAP7_75t_L g217 ( .A(n_218), .Y(n_217) );
INVx2_ASAP7_75t_L g218 ( .A(n_219), .Y(n_218) );
INVx1_ASAP7_75t_L g258 ( .A(n_219), .Y(n_258) );
INVx1_ASAP7_75t_L g230 ( .A(n_220), .Y(n_230) );
OA21x2_ASAP7_75t_L g475 ( .A1(n_220), .A2(n_476), .B(n_485), .Y(n_475) );
OA21x2_ASAP7_75t_L g489 ( .A1(n_220), .A2(n_490), .B(n_498), .Y(n_489) );
INVx2_ASAP7_75t_L g265 ( .A(n_223), .Y(n_265) );
AND2x2_ASAP7_75t_L g397 ( .A(n_223), .B(n_235), .Y(n_397) );
AO21x2_ASAP7_75t_L g223 ( .A1(n_224), .A2(n_230), .B(n_231), .Y(n_223) );
NOR2xp33_ASAP7_75t_L g231 ( .A(n_232), .B(n_233), .Y(n_231) );
NOR2xp33_ASAP7_75t_L g246 ( .A(n_233), .B(n_247), .Y(n_246) );
NOR2xp33_ASAP7_75t_L g278 ( .A(n_233), .B(n_279), .Y(n_278) );
INVx2_ASAP7_75t_L g439 ( .A(n_234), .Y(n_439) );
OR2x2_ASAP7_75t_L g234 ( .A(n_235), .B(n_248), .Y(n_234) );
INVx1_ASAP7_75t_L g284 ( .A(n_235), .Y(n_284) );
AND2x2_ASAP7_75t_L g311 ( .A(n_235), .B(n_312), .Y(n_311) );
NAND2xp5_ASAP7_75t_L g319 ( .A(n_235), .B(n_265), .Y(n_319) );
AND2x2_ASAP7_75t_L g377 ( .A(n_235), .B(n_300), .Y(n_377) );
INVx2_ASAP7_75t_L g235 ( .A(n_236), .Y(n_235) );
INVx1_ASAP7_75t_L g263 ( .A(n_236), .Y(n_263) );
AND2x2_ASAP7_75t_L g290 ( .A(n_236), .B(n_291), .Y(n_290) );
AND2x2_ASAP7_75t_L g299 ( .A(n_236), .B(n_300), .Y(n_299) );
NAND2xp5_ASAP7_75t_L g365 ( .A(n_236), .B(n_265), .Y(n_365) );
AO21x2_ASAP7_75t_L g236 ( .A1(n_237), .A2(n_238), .B(n_246), .Y(n_236) );
NAND2xp5_ASAP7_75t_L g238 ( .A(n_239), .B(n_245), .Y(n_238) );
AOI21xp5_ASAP7_75t_L g240 ( .A1(n_241), .A2(n_242), .B(n_244), .Y(n_240) );
NAND2xp5_ASAP7_75t_L g292 ( .A(n_248), .B(n_293), .Y(n_292) );
INVx2_ASAP7_75t_L g312 ( .A(n_248), .Y(n_312) );
NAND2xp5_ASAP7_75t_L g358 ( .A(n_248), .B(n_265), .Y(n_358) );
AND2x2_ASAP7_75t_L g367 ( .A(n_248), .B(n_368), .Y(n_367) );
INVx1_ASAP7_75t_L g392 ( .A(n_248), .Y(n_392) );
INVx2_ASAP7_75t_L g248 ( .A(n_249), .Y(n_248) );
AND2x2_ASAP7_75t_L g264 ( .A(n_249), .B(n_265), .Y(n_264) );
INVx1_ASAP7_75t_L g300 ( .A(n_249), .Y(n_300) );
NOR2xp33_ASAP7_75t_L g256 ( .A(n_255), .B(n_257), .Y(n_256) );
INVx1_ASAP7_75t_L g494 ( .A(n_255), .Y(n_494) );
AOI21xp5_ASAP7_75t_L g515 ( .A1(n_255), .A2(n_516), .B(n_517), .Y(n_515) );
OAI22xp5_ASAP7_75t_L g428 ( .A1(n_260), .A2(n_270), .B1(n_429), .B2(n_432), .Y(n_428) );
INVx1_ASAP7_75t_SL g260 ( .A(n_261), .Y(n_260) );
OAI21xp5_ASAP7_75t_SL g451 ( .A1(n_262), .A2(n_373), .B(n_452), .Y(n_451) );
AND2x2_ASAP7_75t_L g262 ( .A(n_263), .B(n_264), .Y(n_262) );
NOR2xp33_ASAP7_75t_L g385 ( .A(n_263), .B(n_368), .Y(n_385) );
INVx1_ASAP7_75t_L g410 ( .A(n_263), .Y(n_410) );
NAND2xp5_ASAP7_75t_L g283 ( .A(n_264), .B(n_284), .Y(n_283) );
AND2x2_ASAP7_75t_L g337 ( .A(n_264), .B(n_290), .Y(n_337) );
INVx2_ASAP7_75t_L g293 ( .A(n_265), .Y(n_293) );
INVx1_ASAP7_75t_L g343 ( .A(n_265), .Y(n_343) );
OAI221xp5_ASAP7_75t_L g434 ( .A1(n_266), .A2(n_418), .B1(n_435), .B2(n_438), .C(n_440), .Y(n_434) );
OR2x2_ASAP7_75t_L g266 ( .A(n_267), .B(n_268), .Y(n_266) );
INVx1_ASAP7_75t_L g305 ( .A(n_267), .Y(n_305) );
NAND2xp5_ASAP7_75t_L g357 ( .A(n_267), .B(n_316), .Y(n_357) );
NOR2xp33_ASAP7_75t_L g326 ( .A(n_268), .B(n_327), .Y(n_326) );
OR2x2_ASAP7_75t_L g359 ( .A(n_268), .B(n_305), .Y(n_359) );
INVx3_ASAP7_75t_SL g400 ( .A(n_268), .Y(n_400) );
AND2x2_ASAP7_75t_L g344 ( .A(n_269), .B(n_345), .Y(n_344) );
AND2x2_ASAP7_75t_L g373 ( .A(n_269), .B(n_374), .Y(n_373) );
NAND2xp5_ASAP7_75t_L g388 ( .A(n_269), .B(n_282), .Y(n_388) );
NAND2xp5_ASAP7_75t_L g414 ( .A(n_269), .B(n_328), .Y(n_414) );
INVx3_ASAP7_75t_L g269 ( .A(n_270), .Y(n_269) );
INVx3_ASAP7_75t_L g316 ( .A(n_270), .Y(n_316) );
OAI322xp33_ASAP7_75t_L g411 ( .A1(n_270), .A2(n_342), .A3(n_364), .B1(n_412), .B2(n_414), .C1(n_415), .C2(n_416), .Y(n_411) );
O2A1O1Ixp33_ASAP7_75t_L g491 ( .A1(n_277), .A2(n_492), .B(n_493), .C(n_494), .Y(n_491) );
INVx1_ASAP7_75t_L g280 ( .A(n_281), .Y(n_280) );
AOI21xp33_ASAP7_75t_L g435 ( .A1(n_281), .A2(n_284), .B(n_436), .Y(n_435) );
NOR2xp33_ASAP7_75t_SL g361 ( .A(n_282), .B(n_362), .Y(n_361) );
AND2x2_ASAP7_75t_L g383 ( .A(n_282), .B(n_295), .Y(n_383) );
NAND2xp5_ASAP7_75t_L g398 ( .A(n_282), .B(n_322), .Y(n_398) );
INVxp67_ASAP7_75t_L g349 ( .A(n_284), .Y(n_349) );
AOI211xp5_ASAP7_75t_L g355 ( .A1(n_284), .A2(n_356), .B(n_360), .C(n_370), .Y(n_355) );
OAI221xp5_ASAP7_75t_SL g285 ( .A1(n_286), .A2(n_294), .B1(n_297), .B2(n_301), .C(n_306), .Y(n_285) );
INVxp67_ASAP7_75t_L g286 ( .A(n_287), .Y(n_286) );
OR2x2_ASAP7_75t_L g288 ( .A(n_289), .B(n_292), .Y(n_288) );
INVx1_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
AND2x2_ASAP7_75t_L g309 ( .A(n_293), .B(n_310), .Y(n_309) );
INVx1_ASAP7_75t_L g426 ( .A(n_293), .Y(n_426) );
OAI221xp5_ASAP7_75t_L g442 ( .A1(n_294), .A2(n_443), .B1(n_448), .B2(n_449), .C(n_451), .Y(n_442) );
OR2x2_ASAP7_75t_L g294 ( .A(n_295), .B(n_296), .Y(n_294) );
NAND2xp5_ASAP7_75t_L g338 ( .A(n_295), .B(n_339), .Y(n_338) );
INVx1_ASAP7_75t_SL g342 ( .A(n_295), .Y(n_342) );
NAND2xp5_ASAP7_75t_L g380 ( .A(n_295), .B(n_373), .Y(n_380) );
AND2x2_ASAP7_75t_L g422 ( .A(n_295), .B(n_400), .Y(n_422) );
NOR2xp33_ASAP7_75t_L g320 ( .A(n_296), .B(n_321), .Y(n_320) );
OAI22xp33_ASAP7_75t_L g417 ( .A1(n_296), .A2(n_308), .B1(n_418), .B2(n_419), .Y(n_417) );
OR2x2_ASAP7_75t_L g448 ( .A(n_296), .B(n_316), .Y(n_448) );
CKINVDCx16_ASAP7_75t_R g297 ( .A(n_298), .Y(n_297) );
INVx1_ASAP7_75t_L g425 ( .A(n_299), .Y(n_425) );
AND2x2_ASAP7_75t_L g450 ( .A(n_299), .B(n_393), .Y(n_450) );
INVxp67_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
NOR2xp33_ASAP7_75t_SL g302 ( .A(n_303), .B(n_305), .Y(n_302) );
INVx1_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
OR2x2_ASAP7_75t_L g314 ( .A(n_304), .B(n_315), .Y(n_314) );
AOI22xp5_ASAP7_75t_L g306 ( .A1(n_307), .A2(n_313), .B1(n_317), .B2(n_320), .Y(n_306) );
INVx1_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
NAND2xp5_ASAP7_75t_L g308 ( .A(n_309), .B(n_311), .Y(n_308) );
INVx1_ASAP7_75t_L g381 ( .A(n_309), .Y(n_381) );
NAND2xp5_ASAP7_75t_L g416 ( .A(n_309), .B(n_349), .Y(n_416) );
AOI322xp5_ASAP7_75t_L g340 ( .A1(n_311), .A2(n_341), .A3(n_343), .B1(n_344), .B2(n_346), .C1(n_347), .C2(n_351), .Y(n_340) );
INVxp67_ASAP7_75t_L g334 ( .A(n_312), .Y(n_334) );
INVx1_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
OAI22xp5_ASAP7_75t_L g335 ( .A1(n_314), .A2(n_319), .B1(n_336), .B2(n_338), .Y(n_335) );
NAND2xp5_ASAP7_75t_L g415 ( .A(n_315), .B(n_328), .Y(n_415) );
INVx1_ASAP7_75t_SL g315 ( .A(n_316), .Y(n_315) );
NOR2xp33_ASAP7_75t_L g424 ( .A(n_316), .B(n_354), .Y(n_424) );
NOR2xp33_ASAP7_75t_L g430 ( .A(n_316), .B(n_431), .Y(n_430) );
INVx1_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
OR2x2_ASAP7_75t_L g412 ( .A(n_318), .B(n_413), .Y(n_412) );
INVx1_ASAP7_75t_SL g321 ( .A(n_322), .Y(n_321) );
NAND3xp33_ASAP7_75t_SL g323 ( .A(n_324), .B(n_340), .C(n_355), .Y(n_323) );
AOI221xp5_ASAP7_75t_L g324 ( .A1(n_325), .A2(n_326), .B1(n_331), .B2(n_333), .C(n_335), .Y(n_324) );
AND2x2_ASAP7_75t_L g331 ( .A(n_327), .B(n_332), .Y(n_331) );
INVx3_ASAP7_75t_SL g327 ( .A(n_328), .Y(n_327) );
AND2x4_ASAP7_75t_L g328 ( .A(n_329), .B(n_330), .Y(n_328) );
AND2x2_ASAP7_75t_L g341 ( .A(n_332), .B(n_342), .Y(n_341) );
HB1xp67_ASAP7_75t_L g413 ( .A(n_334), .Y(n_413) );
INVx1_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
NAND2xp5_ASAP7_75t_L g369 ( .A(n_339), .B(n_353), .Y(n_369) );
NAND2xp5_ASAP7_75t_L g406 ( .A(n_342), .B(n_400), .Y(n_406) );
NOR2xp33_ASAP7_75t_L g402 ( .A(n_343), .B(n_403), .Y(n_402) );
INVx1_ASAP7_75t_SL g418 ( .A(n_346), .Y(n_418) );
AND2x2_ASAP7_75t_L g433 ( .A(n_346), .B(n_410), .Y(n_433) );
INVx1_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
NAND2xp5_ASAP7_75t_L g348 ( .A(n_349), .B(n_350), .Y(n_348) );
INVx1_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
AOI211xp5_ASAP7_75t_L g427 ( .A1(n_357), .A2(n_428), .B(n_434), .C(n_442), .Y(n_427) );
INVx1_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
OR2x2_ASAP7_75t_L g364 ( .A(n_365), .B(n_366), .Y(n_364) );
INVx1_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
AND2x2_ASAP7_75t_L g396 ( .A(n_367), .B(n_397), .Y(n_396) );
NAND2x1_ASAP7_75t_SL g438 ( .A(n_368), .B(n_439), .Y(n_438) );
CKINVDCx16_ASAP7_75t_R g408 ( .A(n_371), .Y(n_408) );
INVx1_ASAP7_75t_SL g372 ( .A(n_373), .Y(n_372) );
INVx1_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
INVx1_ASAP7_75t_L g403 ( .A(n_377), .Y(n_403) );
AND2x2_ASAP7_75t_L g407 ( .A(n_377), .B(n_393), .Y(n_407) );
NOR5xp2_ASAP7_75t_L g378 ( .A(n_379), .B(n_394), .C(n_411), .D(n_417), .E(n_420), .Y(n_378) );
OAI221xp5_ASAP7_75t_L g379 ( .A1(n_380), .A2(n_381), .B1(n_382), .B2(n_384), .C(n_386), .Y(n_379) );
INVx2_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
NAND2xp5_ASAP7_75t_L g440 ( .A(n_383), .B(n_441), .Y(n_440) );
INVxp67_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
NAND2xp5_ASAP7_75t_L g386 ( .A(n_387), .B(n_389), .Y(n_386) );
INVx1_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
INVx1_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
NAND2xp5_ASAP7_75t_L g390 ( .A(n_391), .B(n_393), .Y(n_390) );
INVx1_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
AND2x2_ASAP7_75t_L g409 ( .A(n_393), .B(n_410), .Y(n_409) );
OAI221xp5_ASAP7_75t_SL g394 ( .A1(n_395), .A2(n_398), .B1(n_399), .B2(n_401), .C(n_404), .Y(n_394) );
INVx1_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
INVx1_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
AOI22xp33_ASAP7_75t_L g404 ( .A1(n_405), .A2(n_407), .B1(n_408), .B2(n_409), .Y(n_404) );
INVx1_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
INVx1_ASAP7_75t_L g447 ( .A(n_407), .Y(n_447) );
AOI211xp5_ASAP7_75t_SL g420 ( .A1(n_421), .A2(n_423), .B(n_425), .C(n_426), .Y(n_420) );
INVx1_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
INVx1_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
INVx1_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
INVx1_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
INVx1_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
INVxp67_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
NAND2xp5_ASAP7_75t_L g444 ( .A(n_445), .B(n_447), .Y(n_444) );
INVx1_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
CKINVDCx14_ASAP7_75t_R g449 ( .A(n_450), .Y(n_449) );
INVx2_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
INVx1_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
INVx2_ASAP7_75t_L g740 ( .A(n_456), .Y(n_740) );
NAND2x1p5_ASAP7_75t_L g456 ( .A(n_457), .B(n_660), .Y(n_456) );
AND2x2_ASAP7_75t_SL g457 ( .A(n_458), .B(n_618), .Y(n_457) );
NOR4xp25_ASAP7_75t_L g458 ( .A(n_459), .B(n_558), .C(n_594), .D(n_608), .Y(n_458) );
OAI221xp5_ASAP7_75t_SL g459 ( .A1(n_460), .A2(n_506), .B1(n_536), .B2(n_545), .C(n_549), .Y(n_459) );
NAND2xp5_ASAP7_75t_SL g692 ( .A(n_460), .B(n_693), .Y(n_692) );
OR2x2_ASAP7_75t_L g460 ( .A(n_461), .B(n_486), .Y(n_460) );
INVx1_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
AND2x2_ASAP7_75t_L g462 ( .A(n_463), .B(n_474), .Y(n_462) );
AND2x2_ASAP7_75t_L g555 ( .A(n_463), .B(n_475), .Y(n_555) );
INVx3_ASAP7_75t_L g563 ( .A(n_463), .Y(n_563) );
AND2x2_ASAP7_75t_L g617 ( .A(n_463), .B(n_489), .Y(n_617) );
NAND2xp5_ASAP7_75t_L g653 ( .A(n_463), .B(n_488), .Y(n_653) );
AND2x2_ASAP7_75t_L g711 ( .A(n_463), .B(n_573), .Y(n_711) );
AOI21xp5_ASAP7_75t_L g468 ( .A1(n_469), .A2(n_470), .B(n_472), .Y(n_468) );
INVx2_ASAP7_75t_L g482 ( .A(n_471), .Y(n_482) );
O2A1O1Ixp33_ASAP7_75t_L g495 ( .A1(n_472), .A2(n_482), .B(n_496), .C(n_497), .Y(n_495) );
AND2x2_ASAP7_75t_L g546 ( .A(n_474), .B(n_547), .Y(n_546) );
AND2x2_ASAP7_75t_L g560 ( .A(n_474), .B(n_489), .Y(n_560) );
INVx2_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
NAND2xp5_ASAP7_75t_L g575 ( .A(n_475), .B(n_489), .Y(n_575) );
AND2x2_ASAP7_75t_L g587 ( .A(n_475), .B(n_563), .Y(n_587) );
OR2x2_ASAP7_75t_L g589 ( .A(n_475), .B(n_547), .Y(n_589) );
AND2x2_ASAP7_75t_L g624 ( .A(n_475), .B(n_547), .Y(n_624) );
HB1xp67_ASAP7_75t_L g669 ( .A(n_475), .Y(n_669) );
INVx1_ASAP7_75t_L g677 ( .A(n_475), .Y(n_677) );
OAI21xp5_ASAP7_75t_L g476 ( .A1(n_477), .A2(n_480), .B(n_484), .Y(n_476) );
OAI221xp5_ASAP7_75t_L g594 ( .A1(n_486), .A2(n_595), .B1(n_599), .B2(n_603), .C(n_604), .Y(n_594) );
INVx1_ASAP7_75t_L g486 ( .A(n_487), .Y(n_486) );
AND2x2_ASAP7_75t_L g554 ( .A(n_487), .B(n_555), .Y(n_554) );
AND2x2_ASAP7_75t_L g487 ( .A(n_488), .B(n_499), .Y(n_487) );
INVx2_ASAP7_75t_L g553 ( .A(n_488), .Y(n_553) );
AND2x2_ASAP7_75t_L g606 ( .A(n_488), .B(n_607), .Y(n_606) );
AND2x2_ASAP7_75t_L g625 ( .A(n_488), .B(n_563), .Y(n_625) );
INVx2_ASAP7_75t_L g488 ( .A(n_489), .Y(n_488) );
AND2x2_ASAP7_75t_L g688 ( .A(n_489), .B(n_563), .Y(n_688) );
AND2x2_ASAP7_75t_L g610 ( .A(n_499), .B(n_555), .Y(n_610) );
OAI322xp33_ASAP7_75t_L g678 ( .A1(n_499), .A2(n_634), .A3(n_679), .B1(n_681), .B2(n_684), .C1(n_686), .C2(n_690), .Y(n_678) );
INVx3_ASAP7_75t_L g499 ( .A(n_500), .Y(n_499) );
NOR2x1_ASAP7_75t_L g561 ( .A(n_500), .B(n_562), .Y(n_561) );
INVx2_ASAP7_75t_L g574 ( .A(n_500), .Y(n_574) );
AND2x2_ASAP7_75t_L g683 ( .A(n_500), .B(n_563), .Y(n_683) );
AND2x2_ASAP7_75t_L g715 ( .A(n_500), .B(n_587), .Y(n_715) );
OR2x2_ASAP7_75t_L g718 ( .A(n_500), .B(n_719), .Y(n_718) );
AND2x4_ASAP7_75t_L g500 ( .A(n_501), .B(n_502), .Y(n_500) );
INVx1_ASAP7_75t_L g548 ( .A(n_501), .Y(n_548) );
INVx1_ASAP7_75t_L g506 ( .A(n_507), .Y(n_506) );
AND2x2_ASAP7_75t_L g507 ( .A(n_508), .B(n_519), .Y(n_507) );
INVx1_ASAP7_75t_L g731 ( .A(n_508), .Y(n_731) );
INVx1_ASAP7_75t_L g508 ( .A(n_509), .Y(n_508) );
OR2x2_ASAP7_75t_L g538 ( .A(n_509), .B(n_526), .Y(n_538) );
INVx2_ASAP7_75t_L g571 ( .A(n_509), .Y(n_571) );
INVx2_ASAP7_75t_L g509 ( .A(n_510), .Y(n_509) );
INVx2_ASAP7_75t_L g593 ( .A(n_510), .Y(n_593) );
HB1xp67_ASAP7_75t_L g601 ( .A(n_510), .Y(n_601) );
OR2x2_ASAP7_75t_L g725 ( .A(n_510), .B(n_726), .Y(n_725) );
AND2x2_ASAP7_75t_L g550 ( .A(n_519), .B(n_551), .Y(n_550) );
AND2x2_ASAP7_75t_L g590 ( .A(n_519), .B(n_591), .Y(n_590) );
AND2x2_ASAP7_75t_L g642 ( .A(n_519), .B(n_643), .Y(n_642) );
AND2x2_ASAP7_75t_L g519 ( .A(n_520), .B(n_526), .Y(n_519) );
AND2x2_ASAP7_75t_L g539 ( .A(n_520), .B(n_540), .Y(n_539) );
NOR2xp67_ASAP7_75t_L g597 ( .A(n_520), .B(n_598), .Y(n_597) );
AND2x2_ASAP7_75t_L g651 ( .A(n_520), .B(n_541), .Y(n_651) );
OR2x2_ASAP7_75t_L g659 ( .A(n_520), .B(n_593), .Y(n_659) );
INVx2_ASAP7_75t_L g520 ( .A(n_521), .Y(n_520) );
BUFx2_ASAP7_75t_L g568 ( .A(n_521), .Y(n_568) );
AND2x2_ASAP7_75t_L g578 ( .A(n_521), .B(n_579), .Y(n_578) );
AND2x2_ASAP7_75t_L g602 ( .A(n_521), .B(n_526), .Y(n_602) );
AND2x2_ASAP7_75t_L g666 ( .A(n_521), .B(n_541), .Y(n_666) );
NOR2xp33_ASAP7_75t_L g556 ( .A(n_526), .B(n_557), .Y(n_556) );
NAND2xp5_ASAP7_75t_L g570 ( .A(n_526), .B(n_571), .Y(n_570) );
INVx2_ASAP7_75t_L g579 ( .A(n_526), .Y(n_579) );
INVx1_ASAP7_75t_L g584 ( .A(n_526), .Y(n_584) );
AND2x2_ASAP7_75t_L g596 ( .A(n_526), .B(n_597), .Y(n_596) );
HB1xp67_ASAP7_75t_L g674 ( .A(n_526), .Y(n_674) );
INVx1_ASAP7_75t_L g726 ( .A(n_526), .Y(n_726) );
AOI21xp5_ASAP7_75t_L g528 ( .A1(n_529), .A2(n_530), .B(n_531), .Y(n_528) );
NAND2xp5_ASAP7_75t_L g536 ( .A(n_537), .B(n_539), .Y(n_536) );
AND2x2_ASAP7_75t_L g703 ( .A(n_537), .B(n_612), .Y(n_703) );
INVx2_ASAP7_75t_SL g537 ( .A(n_538), .Y(n_537) );
AND2x2_ASAP7_75t_L g630 ( .A(n_539), .B(n_631), .Y(n_630) );
AND2x2_ASAP7_75t_L g729 ( .A(n_539), .B(n_664), .Y(n_729) );
INVx1_ASAP7_75t_L g551 ( .A(n_540), .Y(n_551) );
AND2x2_ASAP7_75t_L g577 ( .A(n_540), .B(n_571), .Y(n_577) );
BUFx2_ASAP7_75t_L g636 ( .A(n_540), .Y(n_636) );
INVx1_ASAP7_75t_L g540 ( .A(n_541), .Y(n_540) );
BUFx6f_ASAP7_75t_L g557 ( .A(n_541), .Y(n_557) );
INVx1_ASAP7_75t_L g567 ( .A(n_541), .Y(n_567) );
NOR2xp67_ASAP7_75t_L g705 ( .A(n_545), .B(n_552), .Y(n_705) );
INVx2_ASAP7_75t_L g545 ( .A(n_546), .Y(n_545) );
AOI32xp33_ASAP7_75t_L g549 ( .A1(n_546), .A2(n_550), .A3(n_552), .B1(n_554), .B2(n_556), .Y(n_549) );
AND2x2_ASAP7_75t_L g689 ( .A(n_546), .B(n_562), .Y(n_689) );
AND2x2_ASAP7_75t_L g727 ( .A(n_546), .B(n_625), .Y(n_727) );
INVx1_ASAP7_75t_L g607 ( .A(n_547), .Y(n_607) );
NAND2xp5_ASAP7_75t_L g721 ( .A(n_551), .B(n_613), .Y(n_721) );
NAND2xp5_ASAP7_75t_L g586 ( .A(n_552), .B(n_587), .Y(n_586) );
NAND2xp5_ASAP7_75t_L g603 ( .A(n_552), .B(n_555), .Y(n_603) );
NAND2xp5_ASAP7_75t_SL g706 ( .A(n_552), .B(n_624), .Y(n_706) );
OR2x2_ASAP7_75t_L g720 ( .A(n_552), .B(n_589), .Y(n_720) );
INVx3_ASAP7_75t_L g552 ( .A(n_553), .Y(n_552) );
AND2x2_ASAP7_75t_L g647 ( .A(n_553), .B(n_555), .Y(n_647) );
OR2x2_ASAP7_75t_L g656 ( .A(n_553), .B(n_643), .Y(n_656) );
NAND2xp5_ASAP7_75t_L g628 ( .A(n_555), .B(n_606), .Y(n_628) );
INVx2_ASAP7_75t_L g643 ( .A(n_557), .Y(n_643) );
OR2x2_ASAP7_75t_L g658 ( .A(n_557), .B(n_659), .Y(n_658) );
AND2x2_ASAP7_75t_L g673 ( .A(n_557), .B(n_674), .Y(n_673) );
A2O1A1Ixp33_ASAP7_75t_L g730 ( .A1(n_557), .A2(n_650), .B(n_731), .C(n_732), .Y(n_730) );
OAI321xp33_ASAP7_75t_L g558 ( .A1(n_559), .A2(n_564), .A3(n_569), .B1(n_572), .B2(n_576), .C(n_580), .Y(n_558) );
INVx1_ASAP7_75t_L g671 ( .A(n_559), .Y(n_671) );
NAND2x1p5_ASAP7_75t_L g559 ( .A(n_560), .B(n_561), .Y(n_559) );
AND2x2_ASAP7_75t_L g682 ( .A(n_560), .B(n_683), .Y(n_682) );
INVx1_ASAP7_75t_L g634 ( .A(n_562), .Y(n_634) );
INVx2_ASAP7_75t_L g562 ( .A(n_563), .Y(n_562) );
NAND2xp5_ASAP7_75t_L g694 ( .A(n_563), .B(n_677), .Y(n_694) );
OAI221xp5_ASAP7_75t_L g701 ( .A1(n_564), .A2(n_702), .B1(n_704), .B2(n_706), .C(n_707), .Y(n_701) );
INVx1_ASAP7_75t_L g564 ( .A(n_565), .Y(n_564) );
AND2x2_ASAP7_75t_L g565 ( .A(n_566), .B(n_568), .Y(n_565) );
AND2x2_ASAP7_75t_L g639 ( .A(n_566), .B(n_613), .Y(n_639) );
HB1xp67_ASAP7_75t_L g566 ( .A(n_567), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g592 ( .A(n_567), .B(n_593), .Y(n_592) );
INVx2_ASAP7_75t_L g612 ( .A(n_568), .Y(n_612) );
A2O1A1Ixp33_ASAP7_75t_L g654 ( .A1(n_569), .A2(n_610), .B(n_655), .C(n_657), .Y(n_654) );
INVx1_ASAP7_75t_L g569 ( .A(n_570), .Y(n_569) );
AND2x2_ASAP7_75t_L g621 ( .A(n_571), .B(n_578), .Y(n_621) );
BUFx2_ASAP7_75t_L g631 ( .A(n_571), .Y(n_631) );
INVx1_ASAP7_75t_L g646 ( .A(n_571), .Y(n_646) );
INVx1_ASAP7_75t_L g572 ( .A(n_573), .Y(n_572) );
NOR2xp33_ASAP7_75t_L g573 ( .A(n_574), .B(n_575), .Y(n_573) );
OR2x2_ASAP7_75t_L g652 ( .A(n_574), .B(n_653), .Y(n_652) );
INVx1_ASAP7_75t_L g735 ( .A(n_574), .Y(n_735) );
INVx1_ASAP7_75t_L g728 ( .A(n_575), .Y(n_728) );
NAND2xp5_ASAP7_75t_L g576 ( .A(n_577), .B(n_578), .Y(n_576) );
AND2x2_ASAP7_75t_L g581 ( .A(n_577), .B(n_582), .Y(n_581) );
AND2x2_ASAP7_75t_L g685 ( .A(n_577), .B(n_602), .Y(n_685) );
INVx1_ASAP7_75t_L g614 ( .A(n_578), .Y(n_614) );
AOI22xp5_ASAP7_75t_L g580 ( .A1(n_581), .A2(n_585), .B1(n_588), .B2(n_590), .Y(n_580) );
NAND2xp5_ASAP7_75t_L g697 ( .A(n_582), .B(n_698), .Y(n_697) );
INVxp67_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
AND2x4_ASAP7_75t_L g650 ( .A(n_583), .B(n_651), .Y(n_650) );
BUFx3_ASAP7_75t_L g583 ( .A(n_584), .Y(n_583) );
AND2x2_ASAP7_75t_SL g613 ( .A(n_584), .B(n_593), .Y(n_613) );
INVx1_ASAP7_75t_L g585 ( .A(n_586), .Y(n_585) );
AND2x2_ASAP7_75t_L g605 ( .A(n_587), .B(n_606), .Y(n_605) );
INVx1_ASAP7_75t_SL g588 ( .A(n_589), .Y(n_588) );
OR2x2_ASAP7_75t_L g615 ( .A(n_589), .B(n_616), .Y(n_615) );
INVx1_ASAP7_75t_SL g591 ( .A(n_592), .Y(n_591) );
OAI221xp5_ASAP7_75t_L g709 ( .A1(n_592), .A2(n_710), .B1(n_712), .B2(n_713), .C(n_714), .Y(n_709) );
INVx1_ASAP7_75t_L g598 ( .A(n_593), .Y(n_598) );
HB1xp67_ASAP7_75t_L g664 ( .A(n_593), .Y(n_664) );
INVx1_ASAP7_75t_SL g595 ( .A(n_596), .Y(n_595) );
NAND2xp5_ASAP7_75t_L g714 ( .A(n_596), .B(n_715), .Y(n_714) );
OAI21xp5_ASAP7_75t_L g604 ( .A1(n_597), .A2(n_602), .B(n_605), .Y(n_604) );
INVx1_ASAP7_75t_L g599 ( .A(n_600), .Y(n_599) );
NAND2xp5_ASAP7_75t_L g707 ( .A(n_600), .B(n_610), .Y(n_707) );
AND2x2_ASAP7_75t_L g600 ( .A(n_601), .B(n_602), .Y(n_600) );
INVx1_ASAP7_75t_L g676 ( .A(n_601), .Y(n_676) );
AND2x2_ASAP7_75t_L g635 ( .A(n_602), .B(n_636), .Y(n_635) );
INVx2_ASAP7_75t_L g724 ( .A(n_602), .Y(n_724) );
INVx1_ASAP7_75t_L g640 ( .A(n_605), .Y(n_640) );
INVx1_ASAP7_75t_L g695 ( .A(n_606), .Y(n_695) );
OAI22xp5_ASAP7_75t_L g608 ( .A1(n_609), .A2(n_611), .B1(n_614), .B2(n_615), .Y(n_608) );
INVx1_ASAP7_75t_L g609 ( .A(n_610), .Y(n_609) );
NAND2xp5_ASAP7_75t_L g611 ( .A(n_612), .B(n_613), .Y(n_611) );
NAND2xp5_ASAP7_75t_L g645 ( .A(n_612), .B(n_646), .Y(n_645) );
INVx2_ASAP7_75t_L g680 ( .A(n_613), .Y(n_680) );
NAND2xp5_ASAP7_75t_SL g717 ( .A(n_613), .B(n_651), .Y(n_717) );
OR2x2_ASAP7_75t_L g690 ( .A(n_614), .B(n_643), .Y(n_690) );
INVx1_ASAP7_75t_L g629 ( .A(n_615), .Y(n_629) );
INVx1_ASAP7_75t_SL g616 ( .A(n_617), .Y(n_616) );
NAND2xp5_ASAP7_75t_L g667 ( .A(n_617), .B(n_668), .Y(n_667) );
NOR3xp33_ASAP7_75t_L g618 ( .A(n_619), .B(n_637), .C(n_648), .Y(n_618) );
OAI211xp5_ASAP7_75t_L g619 ( .A1(n_620), .A2(n_622), .B(n_626), .C(n_632), .Y(n_619) );
INVxp67_ASAP7_75t_L g620 ( .A(n_621), .Y(n_620) );
AOI221xp5_ASAP7_75t_L g691 ( .A1(n_621), .A2(n_692), .B1(n_696), .B2(n_699), .C(n_701), .Y(n_691) );
INVx1_ASAP7_75t_SL g622 ( .A(n_623), .Y(n_622) );
AND2x2_ASAP7_75t_L g623 ( .A(n_624), .B(n_625), .Y(n_623) );
AND2x2_ASAP7_75t_L g633 ( .A(n_624), .B(n_634), .Y(n_633) );
AND2x2_ASAP7_75t_L g687 ( .A(n_624), .B(n_688), .Y(n_687) );
OAI211xp5_ASAP7_75t_L g672 ( .A1(n_625), .A2(n_673), .B(n_675), .C(n_677), .Y(n_672) );
INVx2_ASAP7_75t_L g719 ( .A(n_625), .Y(n_719) );
OAI21xp5_ASAP7_75t_SL g626 ( .A1(n_627), .A2(n_629), .B(n_630), .Y(n_626) );
INVx1_ASAP7_75t_L g627 ( .A(n_628), .Y(n_627) );
AND2x2_ASAP7_75t_L g698 ( .A(n_631), .B(n_651), .Y(n_698) );
NAND2xp5_ASAP7_75t_L g632 ( .A(n_633), .B(n_635), .Y(n_632) );
OAI21xp5_ASAP7_75t_SL g637 ( .A1(n_638), .A2(n_640), .B(n_641), .Y(n_637) );
INVxp67_ASAP7_75t_L g638 ( .A(n_639), .Y(n_638) );
OAI21xp5_ASAP7_75t_SL g641 ( .A1(n_642), .A2(n_644), .B(n_647), .Y(n_641) );
NAND2xp5_ASAP7_75t_L g670 ( .A(n_642), .B(n_671), .Y(n_670) );
INVxp67_ASAP7_75t_L g644 ( .A(n_645), .Y(n_644) );
NAND2xp5_ASAP7_75t_L g733 ( .A(n_647), .B(n_734), .Y(n_733) );
OAI21xp33_ASAP7_75t_L g648 ( .A1(n_649), .A2(n_652), .B(n_654), .Y(n_648) );
INVx1_ASAP7_75t_SL g649 ( .A(n_650), .Y(n_649) );
AND2x2_ASAP7_75t_L g675 ( .A(n_651), .B(n_676), .Y(n_675) );
INVx1_ASAP7_75t_L g655 ( .A(n_656), .Y(n_655) );
INVx1_ASAP7_75t_L g657 ( .A(n_658), .Y(n_657) );
AND4x1_ASAP7_75t_L g660 ( .A(n_661), .B(n_691), .C(n_708), .D(n_730), .Y(n_660) );
NOR2xp33_ASAP7_75t_L g661 ( .A(n_662), .B(n_678), .Y(n_661) );
OAI211xp5_ASAP7_75t_SL g662 ( .A1(n_663), .A2(n_667), .B(n_670), .C(n_672), .Y(n_662) );
OR2x2_ASAP7_75t_L g663 ( .A(n_664), .B(n_665), .Y(n_663) );
INVx1_ASAP7_75t_SL g665 ( .A(n_666), .Y(n_665) );
NAND2xp5_ASAP7_75t_L g679 ( .A(n_666), .B(n_680), .Y(n_679) );
INVx1_ASAP7_75t_L g668 ( .A(n_669), .Y(n_668) );
NOR2xp33_ASAP7_75t_L g699 ( .A(n_677), .B(n_700), .Y(n_699) );
INVx1_ASAP7_75t_L g681 ( .A(n_682), .Y(n_681) );
INVx1_ASAP7_75t_L g684 ( .A(n_685), .Y(n_684) );
NOR2xp33_ASAP7_75t_L g686 ( .A(n_687), .B(n_689), .Y(n_686) );
INVx1_ASAP7_75t_L g712 ( .A(n_687), .Y(n_712) );
INVx2_ASAP7_75t_SL g700 ( .A(n_688), .Y(n_700) );
OR2x2_ASAP7_75t_L g693 ( .A(n_694), .B(n_695), .Y(n_693) );
INVx1_ASAP7_75t_L g696 ( .A(n_697), .Y(n_696) );
INVx1_ASAP7_75t_L g713 ( .A(n_698), .Y(n_713) );
INVx1_ASAP7_75t_L g702 ( .A(n_703), .Y(n_702) );
INVx1_ASAP7_75t_L g704 ( .A(n_705), .Y(n_704) );
NOR2xp33_ASAP7_75t_SL g708 ( .A(n_709), .B(n_716), .Y(n_708) );
INVx1_ASAP7_75t_SL g710 ( .A(n_711), .Y(n_710) );
OAI221xp5_ASAP7_75t_SL g716 ( .A1(n_717), .A2(n_718), .B1(n_720), .B2(n_721), .C(n_722), .Y(n_716) );
AOI22xp5_ASAP7_75t_L g722 ( .A1(n_723), .A2(n_727), .B1(n_728), .B2(n_729), .Y(n_722) );
NAND2xp5_ASAP7_75t_SL g723 ( .A(n_724), .B(n_725), .Y(n_723) );
INVx1_ASAP7_75t_L g732 ( .A(n_733), .Y(n_732) );
INVx1_ASAP7_75t_L g734 ( .A(n_735), .Y(n_734) );
INVx2_ASAP7_75t_L g736 ( .A(n_737), .Y(n_736) );
INVx2_ASAP7_75t_L g741 ( .A(n_737), .Y(n_741) );
INVx1_ASAP7_75t_L g737 ( .A(n_738), .Y(n_737) );
INVx1_ASAP7_75t_L g742 ( .A(n_743), .Y(n_742) );
INVx2_ASAP7_75t_L g743 ( .A(n_744), .Y(n_743) );
CKINVDCx20_ASAP7_75t_R g748 ( .A(n_749), .Y(n_748) );
CKINVDCx20_ASAP7_75t_R g750 ( .A(n_751), .Y(n_750) );
endmodule