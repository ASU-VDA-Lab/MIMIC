module real_jpeg_14170_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_80;
wire n_30;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_83;
wire n_288;
wire n_78;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_195;
wire n_110;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_312;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_299;
wire n_243;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx2_ASAP7_75t_L g116 ( 
.A(n_0),
.Y(n_116)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_1),
.Y(n_42)
);

BUFx4f_ASAP7_75t_L g71 ( 
.A(n_2),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_3),
.A2(n_39),
.B1(n_40),
.B2(n_103),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_3),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_3),
.A2(n_29),
.B1(n_30),
.B2(n_103),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_3),
.A2(n_25),
.B1(n_27),
.B2(n_103),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_3),
.A2(n_67),
.B1(n_72),
.B2(n_103),
.Y(n_209)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

INVx11_ASAP7_75t_L g69 ( 
.A(n_5),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_6),
.A2(n_29),
.B1(n_30),
.B2(n_109),
.Y(n_108)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_6),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g177 ( 
.A1(n_6),
.A2(n_25),
.B1(n_27),
.B2(n_109),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_6),
.A2(n_67),
.B1(n_72),
.B2(n_109),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_L g253 ( 
.A1(n_6),
.A2(n_39),
.B1(n_40),
.B2(n_109),
.Y(n_253)
);

OAI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_7),
.A2(n_39),
.B1(n_40),
.B2(n_51),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_7),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_L g58 ( 
.A1(n_7),
.A2(n_29),
.B1(n_30),
.B2(n_51),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_7),
.A2(n_25),
.B1(n_27),
.B2(n_51),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_7),
.A2(n_51),
.B1(n_67),
.B2(n_72),
.Y(n_129)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

AOI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_9),
.A2(n_39),
.B1(n_40),
.B2(n_62),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_9),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_9),
.A2(n_62),
.B1(n_67),
.B2(n_72),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_9),
.A2(n_25),
.B1(n_27),
.B2(n_62),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_9),
.A2(n_29),
.B1(n_30),
.B2(n_62),
.Y(n_272)
);

BUFx12_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_11),
.A2(n_39),
.B1(n_40),
.B2(n_101),
.Y(n_100)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_11),
.Y(n_101)
);

O2A1O1Ixp33_ASAP7_75t_L g120 ( 
.A1(n_11),
.A2(n_38),
.B(n_39),
.C(n_121),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_11),
.B(n_49),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_11),
.A2(n_25),
.B1(n_27),
.B2(n_101),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_L g208 ( 
.A1(n_11),
.A2(n_126),
.B1(n_151),
.B2(n_209),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_11),
.B(n_31),
.Y(n_222)
);

BUFx8_ASAP7_75t_L g38 ( 
.A(n_12),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_13),
.A2(n_29),
.B1(n_30),
.B2(n_107),
.Y(n_106)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_13),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_13),
.A2(n_39),
.B1(n_40),
.B2(n_107),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g186 ( 
.A1(n_13),
.A2(n_25),
.B1(n_27),
.B2(n_107),
.Y(n_186)
);

AOI22xp33_ASAP7_75t_L g201 ( 
.A1(n_13),
.A2(n_67),
.B1(n_72),
.B2(n_107),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_L g32 ( 
.A1(n_14),
.A2(n_29),
.B1(n_30),
.B2(n_33),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_14),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_14),
.A2(n_25),
.B1(n_27),
.B2(n_33),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_14),
.A2(n_33),
.B1(n_67),
.B2(n_72),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_14),
.A2(n_33),
.B1(n_39),
.B2(n_40),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_L g46 ( 
.A1(n_15),
.A2(n_39),
.B1(n_40),
.B2(n_47),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_15),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_15),
.A2(n_29),
.B1(n_30),
.B2(n_47),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_15),
.A2(n_47),
.B1(n_67),
.B2(n_72),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g246 ( 
.A1(n_15),
.A2(n_25),
.B1(n_27),
.B2(n_47),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_92),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_90),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_76),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_19),
.B(n_76),
.Y(n_91)
);

BUFx24_ASAP7_75t_SL g316 ( 
.A(n_19),
.Y(n_316)
);

FAx1_ASAP7_75t_SL g19 ( 
.A(n_20),
.B(n_34),
.CI(n_52),
.CON(n_19),
.SN(n_19)
);

OAI21xp5_ASAP7_75t_SL g20 ( 
.A1(n_21),
.A2(n_31),
.B(n_32),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_SL g56 ( 
.A(n_21),
.B(n_57),
.Y(n_56)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_21),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_21),
.A2(n_31),
.B1(n_106),
.B2(n_108),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_21),
.A2(n_31),
.B1(n_134),
.B2(n_170),
.Y(n_184)
);

AOI21xp5_ASAP7_75t_L g251 ( 
.A1(n_21),
.A2(n_32),
.B(n_89),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_21),
.A2(n_31),
.B1(n_86),
.B2(n_288),
.Y(n_287)
);

AND2x2_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_28),
.Y(n_21)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_22),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_22),
.B(n_58),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_22),
.A2(n_87),
.B1(n_133),
.B2(n_135),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_L g271 ( 
.A1(n_22),
.A2(n_56),
.B(n_272),
.Y(n_271)
);

OA22x2_ASAP7_75t_SL g22 ( 
.A1(n_23),
.A2(n_24),
.B1(n_25),
.B2(n_27),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_L g28 ( 
.A1(n_23),
.A2(n_24),
.B1(n_29),
.B2(n_30),
.Y(n_28)
);

O2A1O1Ixp33_ASAP7_75t_SL g168 ( 
.A1(n_23),
.A2(n_27),
.B(n_169),
.C(n_171),
.Y(n_168)
);

INVx8_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

NOR3xp33_ASAP7_75t_L g171 ( 
.A(n_24),
.B(n_25),
.C(n_29),
.Y(n_171)
);

INVx6_ASAP7_75t_SL g27 ( 
.A(n_25),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_25),
.A2(n_27),
.B1(n_70),
.B2(n_71),
.Y(n_74)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_SL g192 ( 
.A(n_27),
.B(n_193),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g44 ( 
.A1(n_29),
.A2(n_30),
.B1(n_38),
.B2(n_43),
.Y(n_44)
);

OAI21xp33_ASAP7_75t_L g121 ( 
.A1(n_29),
.A2(n_43),
.B(n_101),
.Y(n_121)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

HAxp5_ASAP7_75t_SL g170 ( 
.A(n_30),
.B(n_101),
.CON(n_170),
.SN(n_170)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_31),
.B(n_32),
.Y(n_55)
);

OAI21xp5_ASAP7_75t_SL g34 ( 
.A1(n_35),
.A2(n_45),
.B(n_48),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_35),
.A2(n_44),
.B1(n_142),
.B2(n_143),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_SL g273 ( 
.A1(n_35),
.A2(n_274),
.B(n_275),
.Y(n_273)
);

OAI21xp5_ASAP7_75t_SL g295 ( 
.A1(n_35),
.A2(n_48),
.B(n_296),
.Y(n_295)
);

CKINVDCx14_ASAP7_75t_R g35 ( 
.A(n_36),
.Y(n_35)
);

AOI22xp5_ASAP7_75t_L g59 ( 
.A1(n_36),
.A2(n_46),
.B1(n_49),
.B2(n_60),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_36),
.B(n_50),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_36),
.A2(n_49),
.B1(n_100),
.B2(n_102),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_36),
.A2(n_49),
.B1(n_144),
.B2(n_253),
.Y(n_252)
);

AND2x2_ASAP7_75t_L g36 ( 
.A(n_37),
.B(n_44),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_L g37 ( 
.A1(n_38),
.A2(n_39),
.B1(n_40),
.B2(n_43),
.Y(n_37)
);

INVx11_ASAP7_75t_L g43 ( 
.A(n_38),
.Y(n_43)
);

INVx5_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx13_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_44),
.Y(n_49)
);

OAI21xp5_ASAP7_75t_L g80 ( 
.A1(n_44),
.A2(n_61),
.B(n_81),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_46),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_49),
.B(n_50),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_49),
.B(n_276),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g52 ( 
.A(n_53),
.B(n_59),
.C(n_63),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_53),
.A2(n_54),
.B1(n_63),
.B2(n_64),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_54),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_55),
.B(n_56),
.Y(n_54)
);

OAI21xp5_ASAP7_75t_L g145 ( 
.A1(n_55),
.A2(n_87),
.B(n_146),
.Y(n_145)
);

INVxp67_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

XOR2xp5_ASAP7_75t_L g78 ( 
.A(n_59),
.B(n_79),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_61),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_63),
.A2(n_64),
.B1(n_83),
.B2(n_84),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_64),
.Y(n_63)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_64),
.B(n_80),
.C(n_83),
.Y(n_82)
);

OAI21xp5_ASAP7_75t_L g64 ( 
.A1(n_65),
.A2(n_73),
.B(n_75),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_65),
.B(n_75),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_65),
.A2(n_73),
.B1(n_177),
.B2(n_186),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_65),
.A2(n_73),
.B1(n_195),
.B2(n_196),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_65),
.A2(n_73),
.B1(n_186),
.B2(n_196),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_65),
.A2(n_73),
.B1(n_245),
.B2(n_246),
.Y(n_244)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

AND2x2_ASAP7_75t_L g73 ( 
.A(n_66),
.B(n_74),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_66),
.B(n_112),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_L g155 ( 
.A1(n_66),
.A2(n_156),
.B(n_157),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_66),
.B(n_101),
.Y(n_212)
);

OA22x2_ASAP7_75t_L g66 ( 
.A1(n_67),
.A2(n_70),
.B1(n_71),
.B2(n_72),
.Y(n_66)
);

CKINVDCx6p67_ASAP7_75t_R g72 ( 
.A(n_67),
.Y(n_72)
);

BUFx12f_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx5_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_70),
.B(n_72),
.C(n_101),
.Y(n_193)
);

INVx13_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_72),
.B(n_116),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_72),
.B(n_207),
.Y(n_206)
);

AOI21xp5_ASAP7_75t_L g110 ( 
.A1(n_73),
.A2(n_75),
.B(n_111),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_73),
.B(n_158),
.Y(n_157)
);

INVxp67_ASAP7_75t_L g175 ( 
.A(n_73),
.Y(n_175)
);

AOI21xp5_ASAP7_75t_L g265 ( 
.A1(n_73),
.A2(n_111),
.B(n_246),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g76 ( 
.A(n_77),
.B(n_80),
.C(n_82),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g309 ( 
.A1(n_77),
.A2(n_78),
.B1(n_80),
.B2(n_306),
.Y(n_309)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g303 ( 
.A1(n_80),
.A2(n_304),
.B1(n_305),
.B2(n_306),
.Y(n_303)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_80),
.Y(n_306)
);

XOR2xp5_ASAP7_75t_L g308 ( 
.A(n_82),
.B(n_309),
.Y(n_308)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

OAI21xp33_ASAP7_75t_L g84 ( 
.A1(n_85),
.A2(n_87),
.B(n_88),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_86),
.Y(n_85)
);

INVxp33_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVxp67_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

OAI21xp5_ASAP7_75t_SL g92 ( 
.A1(n_93),
.A2(n_300),
.B(n_313),
.Y(n_92)
);

AOI21xp5_ASAP7_75t_L g93 ( 
.A1(n_94),
.A2(n_281),
.B(n_299),
.Y(n_93)
);

OAI21xp5_ASAP7_75t_SL g94 ( 
.A1(n_95),
.A2(n_256),
.B(n_280),
.Y(n_94)
);

O2A1O1Ixp33_ASAP7_75t_L g95 ( 
.A1(n_96),
.A2(n_160),
.B(n_237),
.C(n_255),
.Y(n_95)
);

AND2x2_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_136),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_SL g161 ( 
.A(n_97),
.B(n_136),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_98),
.B(n_113),
.C(n_124),
.Y(n_97)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_98),
.B(n_234),
.Y(n_233)
);

XOR2xp5_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_104),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_99),
.B(n_105),
.C(n_110),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_SL g207 ( 
.A(n_101),
.B(n_126),
.Y(n_207)
);

INVxp67_ASAP7_75t_L g142 ( 
.A(n_102),
.Y(n_142)
);

XOR2xp5_ASAP7_75t_L g104 ( 
.A(n_105),
.B(n_110),
.Y(n_104)
);

CKINVDCx14_ASAP7_75t_R g135 ( 
.A(n_106),
.Y(n_135)
);

CKINVDCx14_ASAP7_75t_R g146 ( 
.A(n_108),
.Y(n_146)
);

INVxp67_ASAP7_75t_L g158 ( 
.A(n_112),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_113),
.B(n_124),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_114),
.A2(n_120),
.B1(n_122),
.B2(n_123),
.Y(n_113)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_114),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_115),
.A2(n_116),
.B1(n_117),
.B2(n_119),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_115),
.B(n_128),
.Y(n_127)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_115),
.Y(n_151)
);

AOI21xp5_ASAP7_75t_L g172 ( 
.A1(n_115),
.A2(n_154),
.B(n_173),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_115),
.A2(n_116),
.B1(n_200),
.B2(n_202),
.Y(n_199)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_116),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_116),
.B(n_173),
.Y(n_219)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_L g125 ( 
.A1(n_118),
.A2(n_126),
.B(n_127),
.Y(n_125)
);

CKINVDCx14_ASAP7_75t_R g152 ( 
.A(n_119),
.Y(n_152)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_120),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_120),
.B(n_122),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_125),
.B(n_130),
.C(n_132),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_125),
.A2(n_130),
.B1(n_131),
.B2(n_181),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_125),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_126),
.B(n_129),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g211 ( 
.A1(n_126),
.A2(n_151),
.B1(n_201),
.B2(n_209),
.Y(n_211)
);

AOI21xp5_ASAP7_75t_L g262 ( 
.A1(n_126),
.A2(n_151),
.B(n_263),
.Y(n_262)
);

AND2x2_ASAP7_75t_L g243 ( 
.A(n_127),
.B(n_219),
.Y(n_243)
);

INVxp67_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

XNOR2xp5_ASAP7_75t_SL g179 ( 
.A(n_132),
.B(n_180),
.Y(n_179)
);

INVxp67_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_148),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_137),
.B(n_149),
.C(n_159),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_138),
.A2(n_139),
.B1(n_140),
.B2(n_147),
.Y(n_137)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_138),
.Y(n_147)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_SL g140 ( 
.A(n_141),
.B(n_145),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_141),
.B(n_145),
.C(n_147),
.Y(n_239)
);

CKINVDCx14_ASAP7_75t_R g143 ( 
.A(n_144),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_159),
.Y(n_148)
);

XOR2xp5_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_155),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_150),
.B(n_155),
.Y(n_249)
);

OAI21xp5_ASAP7_75t_L g150 ( 
.A1(n_151),
.A2(n_152),
.B(n_153),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_L g218 ( 
.A1(n_151),
.A2(n_203),
.B(n_219),
.Y(n_218)
);

INVxp67_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

INVxp67_ASAP7_75t_L g245 ( 
.A(n_156),
.Y(n_245)
);

AND2x2_ASAP7_75t_L g289 ( 
.A(n_157),
.B(n_178),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_161),
.B(n_162),
.Y(n_160)
);

AOI21xp5_ASAP7_75t_SL g162 ( 
.A1(n_163),
.A2(n_232),
.B(n_236),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_L g163 ( 
.A1(n_164),
.A2(n_187),
.B(n_231),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_SL g164 ( 
.A(n_165),
.B(n_182),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_165),
.B(n_182),
.Y(n_231)
);

XOR2xp5_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_179),
.Y(n_165)
);

XOR2xp5_ASAP7_75t_L g166 ( 
.A(n_167),
.B(n_174),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_167),
.B(n_174),
.C(n_179),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_172),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_SL g183 ( 
.A(n_168),
.B(n_172),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_170),
.Y(n_169)
);

INVxp67_ASAP7_75t_L g263 ( 
.A(n_173),
.Y(n_263)
);

OAI21xp5_ASAP7_75t_SL g174 ( 
.A1(n_175),
.A2(n_176),
.B(n_178),
.Y(n_174)
);

INVxp67_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_184),
.C(n_185),
.Y(n_182)
);

XOR2xp5_ASAP7_75t_L g227 ( 
.A(n_183),
.B(n_228),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_184),
.B(n_185),
.Y(n_228)
);

AOI21xp5_ASAP7_75t_SL g187 ( 
.A1(n_188),
.A2(n_226),
.B(n_230),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_L g188 ( 
.A1(n_189),
.A2(n_215),
.B(n_225),
.Y(n_188)
);

AOI21xp5_ASAP7_75t_L g189 ( 
.A1(n_190),
.A2(n_204),
.B(n_214),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_191),
.B(n_199),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_191),
.B(n_199),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_192),
.A2(n_194),
.B1(n_197),
.B2(n_198),
.Y(n_191)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_192),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_194),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_194),
.B(n_197),
.Y(n_216)
);

INVxp67_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

CKINVDCx14_ASAP7_75t_R g202 ( 
.A(n_203),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_L g204 ( 
.A1(n_205),
.A2(n_210),
.B(n_213),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_206),
.B(n_208),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_SL g210 ( 
.A(n_211),
.B(n_212),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_211),
.B(n_212),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_216),
.B(n_217),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_216),
.B(n_217),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_220),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_218),
.B(n_221),
.C(n_224),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_221),
.A2(n_222),
.B1(n_223),
.B2(n_224),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_223),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_227),
.B(n_229),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_227),
.B(n_229),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_SL g232 ( 
.A(n_233),
.B(n_235),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_233),
.B(n_235),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_238),
.B(n_254),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_238),
.B(n_254),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_239),
.B(n_240),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_239),
.B(n_241),
.C(n_248),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_241),
.B(n_248),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_242),
.A2(n_243),
.B1(n_244),
.B2(n_247),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_242),
.B(n_247),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_243),
.Y(n_242)
);

CKINVDCx16_ASAP7_75t_R g247 ( 
.A(n_244),
.Y(n_247)
);

XOR2xp5_ASAP7_75t_L g248 ( 
.A(n_249),
.B(n_250),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_249),
.B(n_251),
.C(n_252),
.Y(n_279)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_251),
.B(n_252),
.Y(n_250)
);

CKINVDCx16_ASAP7_75t_R g274 ( 
.A(n_253),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_257),
.B(n_258),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_257),
.B(n_258),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g258 ( 
.A(n_259),
.B(n_279),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_260),
.A2(n_266),
.B1(n_277),
.B2(n_278),
.Y(n_259)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_260),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_260),
.B(n_278),
.C(n_279),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_L g260 ( 
.A1(n_261),
.A2(n_262),
.B1(n_264),
.B2(n_265),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_261),
.A2(n_262),
.B1(n_294),
.B2(n_295),
.Y(n_293)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_262),
.B(n_264),
.Y(n_292)
);

AOI21xp33_ASAP7_75t_L g307 ( 
.A1(n_262),
.A2(n_292),
.B(n_294),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_265),
.Y(n_264)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_266),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_267),
.A2(n_268),
.B1(n_269),
.B2(n_270),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_267),
.B(n_271),
.C(n_273),
.Y(n_284)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

XOR2xp5_ASAP7_75t_L g270 ( 
.A(n_271),
.B(n_273),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_272),
.Y(n_288)
);

CKINVDCx14_ASAP7_75t_R g296 ( 
.A(n_276),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_SL g281 ( 
.A(n_282),
.B(n_298),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_282),
.B(n_298),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g282 ( 
.A1(n_283),
.A2(n_284),
.B1(n_285),
.B2(n_297),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_283),
.B(n_286),
.C(n_291),
.Y(n_311)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_285),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_SL g285 ( 
.A(n_286),
.B(n_291),
.Y(n_285)
);

OAI21xp5_ASAP7_75t_L g286 ( 
.A1(n_287),
.A2(n_289),
.B(n_290),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_SL g290 ( 
.A(n_287),
.B(n_289),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_290),
.B(n_303),
.C(n_307),
.Y(n_302)
);

FAx1_ASAP7_75t_SL g312 ( 
.A(n_290),
.B(n_303),
.CI(n_307),
.CON(n_312),
.SN(n_312)
);

XOR2xp5_ASAP7_75t_L g291 ( 
.A(n_292),
.B(n_293),
.Y(n_291)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_SL g300 ( 
.A(n_301),
.B(n_310),
.Y(n_300)
);

AOI21xp33_ASAP7_75t_L g313 ( 
.A1(n_301),
.A2(n_314),
.B(n_315),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_302),
.B(n_308),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_302),
.B(n_308),
.Y(n_315)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_305),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_311),
.B(n_312),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_311),
.B(n_312),
.Y(n_314)
);

BUFx24_ASAP7_75t_SL g318 ( 
.A(n_312),
.Y(n_318)
);


endmodule