module fake_jpeg_12023_n_620 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_620);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_620;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_170;
wire n_602;
wire n_313;
wire n_574;
wire n_542;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_582;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_387;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_349;
wire n_21;
wire n_288;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_511;
wire n_486;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_615;
wire n_598;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_599;
wire n_239;
wire n_243;
wire n_481;
wire n_619;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_260;
wire n_199;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_613;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_616;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_17),
.Y(n_19)
);

INVx8_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_6),
.Y(n_22)
);

INVx11_ASAP7_75t_SL g23 ( 
.A(n_11),
.Y(n_23)
);

BUFx12_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

INVx6_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_15),
.Y(n_28)
);

INVx2_ASAP7_75t_R g29 ( 
.A(n_3),
.Y(n_29)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_4),
.Y(n_33)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_0),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_2),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_4),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_2),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_17),
.Y(n_38)
);

BUFx10_ASAP7_75t_L g39 ( 
.A(n_3),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_2),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_11),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_9),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_11),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_4),
.Y(n_44)
);

BUFx5_ASAP7_75t_L g45 ( 
.A(n_8),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_17),
.Y(n_46)
);

INVx2_ASAP7_75t_SL g47 ( 
.A(n_5),
.Y(n_47)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_0),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_2),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_8),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_5),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_6),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_10),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_13),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_4),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_15),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_12),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_10),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_11),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_28),
.B(n_8),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_60),
.B(n_76),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_35),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g138 ( 
.A(n_61),
.Y(n_138)
);

BUFx12f_ASAP7_75t_L g62 ( 
.A(n_27),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g149 ( 
.A(n_62),
.Y(n_149)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_27),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g183 ( 
.A(n_63),
.Y(n_183)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_27),
.Y(n_64)
);

BUFx2_ASAP7_75t_L g142 ( 
.A(n_64),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_35),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g154 ( 
.A(n_65),
.Y(n_154)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_36),
.Y(n_66)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_66),
.Y(n_140)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_36),
.Y(n_67)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_67),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_35),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g176 ( 
.A(n_68),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_35),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g180 ( 
.A(n_69),
.Y(n_180)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_59),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g185 ( 
.A(n_70),
.Y(n_185)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_59),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g204 ( 
.A(n_71),
.Y(n_204)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_59),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g207 ( 
.A(n_72),
.Y(n_207)
);

INVx2_ASAP7_75t_SL g73 ( 
.A(n_39),
.Y(n_73)
);

INVx13_ASAP7_75t_L g201 ( 
.A(n_73),
.Y(n_201)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_21),
.Y(n_74)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_74),
.Y(n_133)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_48),
.Y(n_75)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_75),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_28),
.B(n_9),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_21),
.Y(n_77)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_77),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_38),
.B(n_9),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_78),
.B(n_79),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_29),
.B(n_18),
.Y(n_79)
);

BUFx12f_ASAP7_75t_L g80 ( 
.A(n_45),
.Y(n_80)
);

INVx5_ASAP7_75t_L g144 ( 
.A(n_80),
.Y(n_144)
);

INVx8_ASAP7_75t_L g81 ( 
.A(n_45),
.Y(n_81)
);

BUFx2_ASAP7_75t_L g202 ( 
.A(n_81),
.Y(n_202)
);

OR2x2_ASAP7_75t_L g82 ( 
.A(n_31),
.B(n_18),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_82),
.B(n_105),
.Y(n_143)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_53),
.Y(n_83)
);

INVx3_ASAP7_75t_L g151 ( 
.A(n_83),
.Y(n_151)
);

BUFx12f_ASAP7_75t_L g84 ( 
.A(n_45),
.Y(n_84)
);

INVx5_ASAP7_75t_L g147 ( 
.A(n_84),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_29),
.B(n_18),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_85),
.B(n_92),
.Y(n_193)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_59),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g209 ( 
.A(n_86),
.Y(n_209)
);

INVx5_ASAP7_75t_L g87 ( 
.A(n_20),
.Y(n_87)
);

INVx5_ASAP7_75t_L g181 ( 
.A(n_87),
.Y(n_181)
);

INVx5_ASAP7_75t_L g88 ( 
.A(n_20),
.Y(n_88)
);

INVx3_ASAP7_75t_L g160 ( 
.A(n_88),
.Y(n_160)
);

INVx4_ASAP7_75t_SL g89 ( 
.A(n_39),
.Y(n_89)
);

INVx4_ASAP7_75t_L g161 ( 
.A(n_89),
.Y(n_161)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_48),
.Y(n_90)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_90),
.Y(n_156)
);

BUFx12f_ASAP7_75t_L g91 ( 
.A(n_53),
.Y(n_91)
);

INVx4_ASAP7_75t_L g162 ( 
.A(n_91),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_38),
.B(n_18),
.Y(n_92)
);

INVx6_ASAP7_75t_L g93 ( 
.A(n_32),
.Y(n_93)
);

INVx6_ASAP7_75t_L g157 ( 
.A(n_93),
.Y(n_157)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_25),
.Y(n_94)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_94),
.Y(n_172)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_25),
.Y(n_95)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_95),
.Y(n_174)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_26),
.Y(n_96)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_96),
.Y(n_191)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_53),
.Y(n_97)
);

INVx3_ASAP7_75t_L g167 ( 
.A(n_97),
.Y(n_167)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_26),
.Y(n_98)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_98),
.Y(n_194)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_33),
.Y(n_99)
);

INVx3_ASAP7_75t_SL g190 ( 
.A(n_99),
.Y(n_190)
);

INVx5_ASAP7_75t_L g100 ( 
.A(n_20),
.Y(n_100)
);

INVx3_ASAP7_75t_L g179 ( 
.A(n_100),
.Y(n_179)
);

BUFx12f_ASAP7_75t_L g101 ( 
.A(n_40),
.Y(n_101)
);

INVx4_ASAP7_75t_L g170 ( 
.A(n_101),
.Y(n_170)
);

INVx11_ASAP7_75t_L g102 ( 
.A(n_39),
.Y(n_102)
);

INVx11_ASAP7_75t_L g141 ( 
.A(n_102),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_33),
.Y(n_103)
);

INVx4_ASAP7_75t_L g152 ( 
.A(n_103),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_33),
.Y(n_104)
);

INVx4_ASAP7_75t_L g166 ( 
.A(n_104),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_SL g105 ( 
.A(n_29),
.B(n_17),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_37),
.Y(n_106)
);

INVx4_ASAP7_75t_L g169 ( 
.A(n_106),
.Y(n_169)
);

INVx6_ASAP7_75t_L g107 ( 
.A(n_32),
.Y(n_107)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_107),
.Y(n_200)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_26),
.Y(n_108)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_108),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_SL g109 ( 
.A(n_29),
.B(n_16),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_109),
.B(n_126),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_47),
.A2(n_16),
.B1(n_14),
.B2(n_13),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_110),
.A2(n_47),
.B1(n_22),
.B2(n_52),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_37),
.Y(n_111)
);

INVx4_ASAP7_75t_L g188 ( 
.A(n_111),
.Y(n_188)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_37),
.Y(n_112)
);

INVx4_ASAP7_75t_L g197 ( 
.A(n_112),
.Y(n_197)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_44),
.Y(n_113)
);

INVx4_ASAP7_75t_L g208 ( 
.A(n_113),
.Y(n_208)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_44),
.Y(n_114)
);

INVx4_ASAP7_75t_L g210 ( 
.A(n_114),
.Y(n_210)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_40),
.Y(n_115)
);

INVx3_ASAP7_75t_L g186 ( 
.A(n_115),
.Y(n_186)
);

BUFx5_ASAP7_75t_L g116 ( 
.A(n_39),
.Y(n_116)
);

INVx2_ASAP7_75t_SL g137 ( 
.A(n_116),
.Y(n_137)
);

BUFx3_ASAP7_75t_L g117 ( 
.A(n_19),
.Y(n_117)
);

INVx2_ASAP7_75t_SL g164 ( 
.A(n_117),
.Y(n_164)
);

BUFx3_ASAP7_75t_L g118 ( 
.A(n_19),
.Y(n_118)
);

INVx2_ASAP7_75t_SL g192 ( 
.A(n_118),
.Y(n_192)
);

INVx8_ASAP7_75t_L g119 ( 
.A(n_39),
.Y(n_119)
);

INVx3_ASAP7_75t_L g195 ( 
.A(n_119),
.Y(n_195)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_44),
.Y(n_120)
);

INVx3_ASAP7_75t_L g199 ( 
.A(n_120),
.Y(n_199)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_34),
.Y(n_121)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_121),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_49),
.Y(n_122)
);

INVx3_ASAP7_75t_L g206 ( 
.A(n_122),
.Y(n_206)
);

BUFx24_ASAP7_75t_L g123 ( 
.A(n_23),
.Y(n_123)
);

INVx6_ASAP7_75t_SL g173 ( 
.A(n_123),
.Y(n_173)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_49),
.Y(n_124)
);

INVx3_ASAP7_75t_L g211 ( 
.A(n_124),
.Y(n_211)
);

INVx11_ASAP7_75t_L g125 ( 
.A(n_23),
.Y(n_125)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_125),
.Y(n_168)
);

BUFx3_ASAP7_75t_L g126 ( 
.A(n_19),
.Y(n_126)
);

INVx6_ASAP7_75t_L g127 ( 
.A(n_32),
.Y(n_127)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_127),
.Y(n_177)
);

AOI22xp33_ASAP7_75t_L g128 ( 
.A1(n_93),
.A2(n_34),
.B1(n_47),
.B2(n_49),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g250 ( 
.A1(n_128),
.A2(n_131),
.B1(n_132),
.B2(n_134),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_129),
.A2(n_130),
.B1(n_158),
.B2(n_163),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_82),
.A2(n_30),
.B1(n_58),
.B2(n_42),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_64),
.A2(n_40),
.B1(n_51),
.B2(n_81),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_107),
.A2(n_30),
.B1(n_58),
.B2(n_43),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_127),
.A2(n_30),
.B1(n_58),
.B2(n_43),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_SL g135 ( 
.A1(n_63),
.A2(n_51),
.B1(n_34),
.B2(n_47),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_SL g215 ( 
.A1(n_135),
.A2(n_136),
.B1(n_145),
.B2(n_171),
.Y(n_215)
);

AOI22xp33_ASAP7_75t_SL g136 ( 
.A1(n_119),
.A2(n_51),
.B1(n_42),
.B2(n_43),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_SL g139 ( 
.A(n_62),
.B(n_41),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_SL g212 ( 
.A(n_139),
.B(n_153),
.Y(n_212)
);

AOI22xp33_ASAP7_75t_SL g145 ( 
.A1(n_73),
.A2(n_62),
.B1(n_80),
.B2(n_84),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_101),
.B(n_50),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g158 ( 
.A1(n_99),
.A2(n_57),
.B1(n_42),
.B2(n_50),
.Y(n_158)
);

OAI22xp33_ASAP7_75t_SL g163 ( 
.A1(n_103),
.A2(n_57),
.B1(n_55),
.B2(n_46),
.Y(n_163)
);

AOI22xp33_ASAP7_75t_SL g171 ( 
.A1(n_80),
.A2(n_57),
.B1(n_19),
.B2(n_46),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_123),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_SL g217 ( 
.A(n_175),
.B(n_178),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_101),
.B(n_56),
.Y(n_178)
);

AOI22xp33_ASAP7_75t_L g182 ( 
.A1(n_104),
.A2(n_22),
.B1(n_52),
.B2(n_55),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_182),
.A2(n_110),
.B1(n_61),
.B2(n_69),
.Y(n_233)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_117),
.Y(n_184)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_184),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_91),
.B(n_56),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_SL g264 ( 
.A(n_189),
.B(n_198),
.Y(n_264)
);

HAxp5_ASAP7_75t_SL g196 ( 
.A(n_102),
.B(n_123),
.CON(n_196),
.SN(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_196),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_91),
.B(n_41),
.Y(n_198)
);

AOI22xp33_ASAP7_75t_SL g203 ( 
.A1(n_84),
.A2(n_19),
.B1(n_31),
.B2(n_54),
.Y(n_203)
);

AOI22xp33_ASAP7_75t_SL g235 ( 
.A1(n_203),
.A2(n_125),
.B1(n_120),
.B2(n_114),
.Y(n_235)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_177),
.Y(n_213)
);

INVx2_ASAP7_75t_L g300 ( 
.A(n_213),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_159),
.B(n_54),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_SL g328 ( 
.A(n_214),
.B(n_219),
.Y(n_328)
);

INVxp67_ASAP7_75t_L g218 ( 
.A(n_145),
.Y(n_218)
);

HB1xp67_ASAP7_75t_L g337 ( 
.A(n_218),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_187),
.B(n_16),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_173),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_220),
.B(n_226),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_SL g221 ( 
.A(n_143),
.B(n_126),
.Y(n_221)
);

OAI21xp33_ASAP7_75t_L g333 ( 
.A1(n_221),
.A2(n_261),
.B(n_272),
.Y(n_333)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_200),
.Y(n_222)
);

INVx2_ASAP7_75t_L g306 ( 
.A(n_222),
.Y(n_306)
);

BUFx2_ASAP7_75t_L g223 ( 
.A(n_144),
.Y(n_223)
);

INVx1_ASAP7_75t_SL g302 ( 
.A(n_223),
.Y(n_302)
);

BUFx12f_ASAP7_75t_L g224 ( 
.A(n_149),
.Y(n_224)
);

BUFx3_ASAP7_75t_L g287 ( 
.A(n_224),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_133),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_163),
.A2(n_113),
.B1(n_124),
.B2(n_122),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_L g285 ( 
.A1(n_227),
.A2(n_239),
.B1(n_249),
.B2(n_262),
.Y(n_285)
);

BUFx3_ASAP7_75t_L g228 ( 
.A(n_149),
.Y(n_228)
);

BUFx12f_ASAP7_75t_L g315 ( 
.A(n_228),
.Y(n_315)
);

INVx4_ASAP7_75t_L g229 ( 
.A(n_162),
.Y(n_229)
);

INVx4_ASAP7_75t_L g289 ( 
.A(n_229),
.Y(n_289)
);

AND2x4_ASAP7_75t_L g230 ( 
.A(n_191),
.B(n_118),
.Y(n_230)
);

AND2x2_ASAP7_75t_L g317 ( 
.A(n_230),
.B(n_256),
.Y(n_317)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_194),
.Y(n_231)
);

INVx2_ASAP7_75t_L g332 ( 
.A(n_231),
.Y(n_332)
);

INVx3_ASAP7_75t_L g232 ( 
.A(n_181),
.Y(n_232)
);

INVx4_ASAP7_75t_L g298 ( 
.A(n_232),
.Y(n_298)
);

AOI22xp33_ASAP7_75t_L g294 ( 
.A1(n_233),
.A2(n_202),
.B1(n_210),
.B2(n_208),
.Y(n_294)
);

INVx2_ASAP7_75t_SL g234 ( 
.A(n_160),
.Y(n_234)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_234),
.Y(n_296)
);

AOI22xp33_ASAP7_75t_SL g297 ( 
.A1(n_235),
.A2(n_241),
.B1(n_245),
.B2(n_282),
.Y(n_297)
);

INVx4_ASAP7_75t_L g236 ( 
.A(n_147),
.Y(n_236)
);

INVx4_ASAP7_75t_L g304 ( 
.A(n_236),
.Y(n_304)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_150),
.Y(n_237)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_237),
.Y(n_310)
);

INVx4_ASAP7_75t_L g238 ( 
.A(n_179),
.Y(n_238)
);

INVx3_ASAP7_75t_L g301 ( 
.A(n_238),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_157),
.A2(n_112),
.B1(n_111),
.B2(n_106),
.Y(n_239)
);

INVx4_ASAP7_75t_L g240 ( 
.A(n_170),
.Y(n_240)
);

INVx5_ASAP7_75t_L g295 ( 
.A(n_240),
.Y(n_295)
);

AOI22xp33_ASAP7_75t_SL g241 ( 
.A1(n_196),
.A2(n_65),
.B1(n_68),
.B2(n_72),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_193),
.B(n_12),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_242),
.B(n_253),
.Y(n_307)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_205),
.Y(n_243)
);

INVx2_ASAP7_75t_L g341 ( 
.A(n_243),
.Y(n_341)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_165),
.Y(n_244)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_244),
.Y(n_321)
);

AOI22xp33_ASAP7_75t_SL g245 ( 
.A1(n_142),
.A2(n_86),
.B1(n_71),
.B2(n_70),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_151),
.Y(n_246)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_246),
.Y(n_322)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_167),
.Y(n_247)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_247),
.Y(n_339)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_140),
.Y(n_248)
);

BUFx6f_ASAP7_75t_L g290 ( 
.A(n_248),
.Y(n_290)
);

OAI22xp33_ASAP7_75t_SL g249 ( 
.A1(n_136),
.A2(n_89),
.B1(n_24),
.B2(n_16),
.Y(n_249)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_146),
.Y(n_251)
);

BUFx6f_ASAP7_75t_L g331 ( 
.A(n_251),
.Y(n_331)
);

INVxp33_ASAP7_75t_L g252 ( 
.A(n_201),
.Y(n_252)
);

INVx11_ASAP7_75t_L g327 ( 
.A(n_252),
.Y(n_327)
);

CKINVDCx16_ASAP7_75t_R g253 ( 
.A(n_141),
.Y(n_253)
);

INVx3_ASAP7_75t_L g254 ( 
.A(n_168),
.Y(n_254)
);

INVx6_ASAP7_75t_L g312 ( 
.A(n_254),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_182),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_255),
.B(n_258),
.Y(n_319)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_155),
.Y(n_256)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_156),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_148),
.B(n_0),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_259),
.B(n_266),
.Y(n_291)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_186),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_260),
.B(n_263),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_172),
.B(n_14),
.Y(n_261)
);

OAI22xp33_ASAP7_75t_SL g262 ( 
.A1(n_131),
.A2(n_24),
.B1(n_14),
.B2(n_13),
.Y(n_262)
);

INVxp67_ASAP7_75t_L g263 ( 
.A(n_203),
.Y(n_263)
);

AOI22xp33_ASAP7_75t_L g265 ( 
.A1(n_128),
.A2(n_24),
.B1(n_13),
.B2(n_12),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_L g308 ( 
.A1(n_265),
.A2(n_284),
.B1(n_227),
.B2(n_239),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_174),
.B(n_0),
.Y(n_266)
);

BUFx3_ASAP7_75t_L g267 ( 
.A(n_164),
.Y(n_267)
);

BUFx10_ASAP7_75t_L g305 ( 
.A(n_267),
.Y(n_305)
);

AO22x2_ASAP7_75t_L g268 ( 
.A1(n_135),
.A2(n_169),
.B1(n_210),
.B2(n_208),
.Y(n_268)
);

OR2x2_ASAP7_75t_L g340 ( 
.A(n_268),
.B(n_269),
.Y(n_340)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_161),
.Y(n_269)
);

INVx4_ASAP7_75t_L g270 ( 
.A(n_195),
.Y(n_270)
);

INVx6_ASAP7_75t_L g330 ( 
.A(n_270),
.Y(n_330)
);

INVx6_ASAP7_75t_L g271 ( 
.A(n_185),
.Y(n_271)
);

INVx8_ASAP7_75t_L g335 ( 
.A(n_271),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_164),
.B(n_10),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_141),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g293 ( 
.A(n_273),
.Y(n_293)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_157),
.Y(n_274)
);

AND2x2_ASAP7_75t_L g338 ( 
.A(n_274),
.B(n_275),
.Y(n_338)
);

INVx3_ASAP7_75t_L g275 ( 
.A(n_183),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_201),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g299 ( 
.A(n_276),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_152),
.B(n_0),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_277),
.B(n_283),
.Y(n_314)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_199),
.Y(n_278)
);

CKINVDCx16_ASAP7_75t_R g326 ( 
.A(n_278),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_192),
.B(n_1),
.Y(n_279)
);

CKINVDCx16_ASAP7_75t_R g329 ( 
.A(n_279),
.Y(n_329)
);

INVx4_ASAP7_75t_L g280 ( 
.A(n_183),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_280),
.Y(n_320)
);

INVx3_ASAP7_75t_L g281 ( 
.A(n_152),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g325 ( 
.A(n_281),
.Y(n_325)
);

INVx6_ASAP7_75t_L g282 ( 
.A(n_185),
.Y(n_282)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_192),
.Y(n_283)
);

AOI22xp33_ASAP7_75t_L g284 ( 
.A1(n_206),
.A2(n_24),
.B1(n_2),
.B2(n_3),
.Y(n_284)
);

A2O1A1Ixp33_ASAP7_75t_L g286 ( 
.A1(n_257),
.A2(n_171),
.B(n_137),
.C(n_142),
.Y(n_286)
);

A2O1A1Ixp33_ASAP7_75t_L g344 ( 
.A1(n_286),
.A2(n_303),
.B(n_230),
.C(n_268),
.Y(n_344)
);

XNOR2x1_ASAP7_75t_SL g292 ( 
.A(n_257),
.B(n_202),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g347 ( 
.A(n_292),
.B(n_317),
.Y(n_347)
);

OAI22xp5_ASAP7_75t_L g377 ( 
.A1(n_294),
.A2(n_324),
.B1(n_334),
.B2(n_282),
.Y(n_377)
);

A2O1A1Ixp33_ASAP7_75t_L g303 ( 
.A1(n_259),
.A2(n_137),
.B(n_190),
.C(n_197),
.Y(n_303)
);

AND2x2_ASAP7_75t_L g354 ( 
.A(n_308),
.B(n_268),
.Y(n_354)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_225),
.B(n_211),
.C(n_190),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g355 ( 
.A(n_309),
.B(n_230),
.C(n_234),
.Y(n_355)
);

OR2x2_ASAP7_75t_SL g311 ( 
.A(n_218),
.B(n_166),
.Y(n_311)
);

MAJx2_ASAP7_75t_L g361 ( 
.A(n_311),
.B(n_318),
.C(n_283),
.Y(n_361)
);

OAI22xp5_ASAP7_75t_L g313 ( 
.A1(n_216),
.A2(n_166),
.B1(n_197),
.B2(n_188),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_L g383 ( 
.A1(n_313),
.A2(n_222),
.B1(n_248),
.B2(n_267),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_266),
.B(n_188),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_316),
.B(n_336),
.Y(n_353)
);

OR2x2_ASAP7_75t_SL g318 ( 
.A(n_264),
.B(n_169),
.Y(n_318)
);

AOI22xp33_ASAP7_75t_L g324 ( 
.A1(n_233),
.A2(n_138),
.B1(n_180),
.B2(n_176),
.Y(n_324)
);

AOI22xp33_ASAP7_75t_L g334 ( 
.A1(n_263),
.A2(n_138),
.B1(n_180),
.B2(n_176),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_277),
.B(n_154),
.Y(n_336)
);

OAI22xp5_ASAP7_75t_SL g342 ( 
.A1(n_340),
.A2(n_216),
.B1(n_215),
.B2(n_250),
.Y(n_342)
);

AOI22xp5_ASAP7_75t_L g411 ( 
.A1(n_342),
.A2(n_359),
.B1(n_381),
.B2(n_301),
.Y(n_411)
);

OAI32xp33_ASAP7_75t_L g343 ( 
.A1(n_314),
.A2(n_212),
.A3(n_217),
.B1(n_231),
.B2(n_243),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_343),
.B(n_348),
.Y(n_388)
);

AOI21xp5_ASAP7_75t_L g394 ( 
.A1(n_344),
.A2(n_351),
.B(n_363),
.Y(n_394)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_296),
.Y(n_345)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_345),
.Y(n_397)
);

BUFx24_ASAP7_75t_SL g346 ( 
.A(n_328),
.Y(n_346)
);

NOR2xp33_ASAP7_75t_L g406 ( 
.A(n_346),
.B(n_349),
.Y(n_406)
);

XNOR2xp5_ASAP7_75t_SL g399 ( 
.A(n_347),
.B(n_355),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_SL g348 ( 
.A(n_291),
.B(n_254),
.Y(n_348)
);

INVxp67_ASAP7_75t_L g349 ( 
.A(n_327),
.Y(n_349)
);

OAI21xp5_ASAP7_75t_L g350 ( 
.A1(n_340),
.A2(n_230),
.B(n_252),
.Y(n_350)
);

OAI21xp5_ASAP7_75t_L g414 ( 
.A1(n_350),
.A2(n_301),
.B(n_339),
.Y(n_414)
);

AOI21xp5_ASAP7_75t_L g351 ( 
.A1(n_286),
.A2(n_268),
.B(n_234),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_296),
.Y(n_352)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_352),
.Y(n_400)
);

AOI22xp33_ASAP7_75t_L g390 ( 
.A1(n_354),
.A2(n_383),
.B1(n_338),
.B2(n_302),
.Y(n_390)
);

INVx1_ASAP7_75t_SL g356 ( 
.A(n_327),
.Y(n_356)
);

INVx2_ASAP7_75t_L g392 ( 
.A(n_356),
.Y(n_392)
);

AOI22xp33_ASAP7_75t_SL g357 ( 
.A1(n_337),
.A2(n_275),
.B1(n_280),
.B2(n_232),
.Y(n_357)
);

AOI22xp33_ASAP7_75t_SL g401 ( 
.A1(n_357),
.A2(n_358),
.B1(n_366),
.B2(n_367),
.Y(n_401)
);

AOI22xp33_ASAP7_75t_SL g358 ( 
.A1(n_311),
.A2(n_238),
.B1(n_270),
.B2(n_228),
.Y(n_358)
);

OAI22xp5_ASAP7_75t_SL g359 ( 
.A1(n_297),
.A2(n_274),
.B1(n_154),
.B2(n_207),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_310),
.Y(n_360)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_360),
.Y(n_404)
);

CKINVDCx14_ASAP7_75t_R g405 ( 
.A(n_361),
.Y(n_405)
);

AOI22xp33_ASAP7_75t_L g362 ( 
.A1(n_319),
.A2(n_209),
.B1(n_207),
.B2(n_204),
.Y(n_362)
);

OAI22xp5_ASAP7_75t_L g387 ( 
.A1(n_362),
.A2(n_302),
.B1(n_335),
.B2(n_299),
.Y(n_387)
);

AOI22xp5_ASAP7_75t_SL g363 ( 
.A1(n_329),
.A2(n_285),
.B1(n_317),
.B2(n_292),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_310),
.Y(n_364)
);

INVx2_ASAP7_75t_L g420 ( 
.A(n_364),
.Y(n_420)
);

INVx2_ASAP7_75t_L g365 ( 
.A(n_290),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_365),
.B(n_369),
.Y(n_389)
);

AOI22xp33_ASAP7_75t_SL g366 ( 
.A1(n_293),
.A2(n_330),
.B1(n_312),
.B2(n_298),
.Y(n_366)
);

INVx3_ASAP7_75t_L g367 ( 
.A(n_330),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_300),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_SL g417 ( 
.A(n_368),
.B(n_373),
.Y(n_417)
);

BUFx3_ASAP7_75t_L g369 ( 
.A(n_315),
.Y(n_369)
);

CKINVDCx20_ASAP7_75t_R g370 ( 
.A(n_288),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_370),
.B(n_374),
.Y(n_396)
);

MAJIxp5_ASAP7_75t_L g371 ( 
.A(n_314),
.B(n_256),
.C(n_251),
.Y(n_371)
);

XNOR2xp5_ASAP7_75t_SL g422 ( 
.A(n_371),
.B(n_372),
.Y(n_422)
);

AND2x2_ASAP7_75t_L g372 ( 
.A(n_317),
.B(n_323),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_300),
.Y(n_373)
);

CKINVDCx20_ASAP7_75t_R g374 ( 
.A(n_299),
.Y(n_374)
);

AOI21xp5_ASAP7_75t_L g375 ( 
.A1(n_293),
.A2(n_236),
.B(n_223),
.Y(n_375)
);

AOI21xp5_ASAP7_75t_L g395 ( 
.A1(n_375),
.A2(n_378),
.B(n_305),
.Y(n_395)
);

INVx2_ASAP7_75t_L g376 ( 
.A(n_290),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_376),
.B(n_380),
.Y(n_412)
);

CKINVDCx16_ASAP7_75t_R g391 ( 
.A(n_377),
.Y(n_391)
);

AOI22xp5_ASAP7_75t_SL g378 ( 
.A1(n_318),
.A2(n_281),
.B1(n_213),
.B2(n_229),
.Y(n_378)
);

BUFx2_ASAP7_75t_L g379 ( 
.A(n_335),
.Y(n_379)
);

CKINVDCx16_ASAP7_75t_R g402 ( 
.A(n_379),
.Y(n_402)
);

INVx2_ASAP7_75t_L g380 ( 
.A(n_331),
.Y(n_380)
);

OAI22xp5_ASAP7_75t_L g381 ( 
.A1(n_336),
.A2(n_204),
.B1(n_209),
.B2(n_271),
.Y(n_381)
);

INVxp67_ASAP7_75t_L g382 ( 
.A(n_307),
.Y(n_382)
);

NOR2xp33_ASAP7_75t_SL g398 ( 
.A(n_382),
.B(n_384),
.Y(n_398)
);

INVxp67_ASAP7_75t_L g384 ( 
.A(n_305),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_291),
.B(n_240),
.Y(n_385)
);

CKINVDCx20_ASAP7_75t_R g418 ( 
.A(n_385),
.Y(n_418)
);

OAI22xp5_ASAP7_75t_SL g386 ( 
.A1(n_363),
.A2(n_316),
.B1(n_309),
.B2(n_303),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_386),
.B(n_393),
.Y(n_443)
);

INVxp67_ASAP7_75t_SL g423 ( 
.A(n_387),
.Y(n_423)
);

OAI22xp5_ASAP7_75t_L g430 ( 
.A1(n_390),
.A2(n_403),
.B1(n_411),
.B2(n_419),
.Y(n_430)
);

OAI22xp5_ASAP7_75t_SL g393 ( 
.A1(n_351),
.A2(n_333),
.B1(n_321),
.B2(n_320),
.Y(n_393)
);

INVxp67_ASAP7_75t_L g425 ( 
.A(n_395),
.Y(n_425)
);

AOI22xp33_ASAP7_75t_L g403 ( 
.A1(n_354),
.A2(n_338),
.B1(n_320),
.B2(n_321),
.Y(n_403)
);

OAI22xp5_ASAP7_75t_L g407 ( 
.A1(n_342),
.A2(n_325),
.B1(n_312),
.B2(n_298),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g444 ( 
.A(n_407),
.B(n_413),
.Y(n_444)
);

AO22x1_ASAP7_75t_L g408 ( 
.A1(n_350),
.A2(n_339),
.B1(n_322),
.B2(n_332),
.Y(n_408)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_408),
.Y(n_456)
);

AOI21xp5_ASAP7_75t_L g409 ( 
.A1(n_347),
.A2(n_325),
.B(n_338),
.Y(n_409)
);

OAI21xp5_ASAP7_75t_L g447 ( 
.A1(n_409),
.A2(n_410),
.B(n_414),
.Y(n_447)
);

AOI21xp5_ASAP7_75t_L g410 ( 
.A1(n_344),
.A2(n_305),
.B(n_304),
.Y(n_410)
);

OAI22xp5_ASAP7_75t_SL g413 ( 
.A1(n_354),
.A2(n_344),
.B1(n_353),
.B2(n_385),
.Y(n_413)
);

AOI21xp5_ASAP7_75t_L g415 ( 
.A1(n_375),
.A2(n_305),
.B(n_304),
.Y(n_415)
);

INVxp67_ASAP7_75t_L g450 ( 
.A(n_415),
.Y(n_450)
);

OA21x2_ASAP7_75t_L g416 ( 
.A1(n_372),
.A2(n_322),
.B(n_332),
.Y(n_416)
);

NOR2xp33_ASAP7_75t_L g424 ( 
.A(n_416),
.B(n_374),
.Y(n_424)
);

AOI22xp5_ASAP7_75t_L g419 ( 
.A1(n_377),
.A2(n_331),
.B1(n_341),
.B2(n_306),
.Y(n_419)
);

AOI22xp5_ASAP7_75t_SL g421 ( 
.A1(n_372),
.A2(n_355),
.B1(n_359),
.B2(n_361),
.Y(n_421)
);

OAI22xp5_ASAP7_75t_SL g436 ( 
.A1(n_421),
.A2(n_356),
.B1(n_379),
.B2(n_373),
.Y(n_436)
);

OAI21xp5_ASAP7_75t_SL g478 ( 
.A1(n_424),
.A2(n_426),
.B(n_408),
.Y(n_478)
);

AOI32xp33_ASAP7_75t_L g426 ( 
.A1(n_388),
.A2(n_343),
.A3(n_361),
.B1(n_378),
.B2(n_348),
.Y(n_426)
);

CKINVDCx16_ASAP7_75t_R g427 ( 
.A(n_396),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_SL g462 ( 
.A(n_427),
.B(n_435),
.Y(n_462)
);

XNOR2xp5_ASAP7_75t_SL g428 ( 
.A(n_399),
.B(n_353),
.Y(n_428)
);

XOR2xp5_ASAP7_75t_L g469 ( 
.A(n_428),
.B(n_436),
.Y(n_469)
);

XNOR2xp5_ASAP7_75t_L g429 ( 
.A(n_399),
.B(n_422),
.Y(n_429)
);

MAJIxp5_ASAP7_75t_L g463 ( 
.A(n_429),
.B(n_431),
.C(n_422),
.Y(n_463)
);

MAJIxp5_ASAP7_75t_L g431 ( 
.A(n_399),
.B(n_371),
.C(n_370),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_SL g432 ( 
.A(n_396),
.B(n_345),
.Y(n_432)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_432),
.Y(n_458)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_420),
.Y(n_433)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_433),
.Y(n_468)
);

OAI22xp5_ASAP7_75t_L g434 ( 
.A1(n_391),
.A2(n_362),
.B1(n_383),
.B2(n_352),
.Y(n_434)
);

AOI22xp5_ASAP7_75t_L g460 ( 
.A1(n_434),
.A2(n_438),
.B1(n_387),
.B2(n_407),
.Y(n_460)
);

NAND3xp33_ASAP7_75t_L g435 ( 
.A(n_405),
.B(n_360),
.C(n_364),
.Y(n_435)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_420),
.Y(n_437)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_437),
.Y(n_486)
);

OAI22xp5_ASAP7_75t_SL g438 ( 
.A1(n_391),
.A2(n_381),
.B1(n_356),
.B2(n_379),
.Y(n_438)
);

NOR2xp33_ASAP7_75t_L g439 ( 
.A(n_398),
.B(n_368),
.Y(n_439)
);

INVxp33_ASAP7_75t_L g476 ( 
.A(n_439),
.Y(n_476)
);

CKINVDCx16_ASAP7_75t_R g440 ( 
.A(n_398),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_SL g466 ( 
.A(n_440),
.B(n_442),
.Y(n_466)
);

CKINVDCx20_ASAP7_75t_R g441 ( 
.A(n_417),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_L g464 ( 
.A(n_441),
.B(n_446),
.Y(n_464)
);

NOR2xp33_ASAP7_75t_L g442 ( 
.A(n_418),
.B(n_367),
.Y(n_442)
);

AOI22xp33_ASAP7_75t_SL g445 ( 
.A1(n_393),
.A2(n_369),
.B1(n_315),
.B2(n_287),
.Y(n_445)
);

A2O1A1Ixp33_ASAP7_75t_SL g461 ( 
.A1(n_445),
.A2(n_395),
.B(n_415),
.C(n_410),
.Y(n_461)
);

CKINVDCx20_ASAP7_75t_R g446 ( 
.A(n_417),
.Y(n_446)
);

NOR2xp33_ASAP7_75t_L g448 ( 
.A(n_418),
.B(n_380),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_L g465 ( 
.A(n_448),
.B(n_451),
.Y(n_465)
);

INVx2_ASAP7_75t_L g449 ( 
.A(n_397),
.Y(n_449)
);

INVx2_ASAP7_75t_L g459 ( 
.A(n_449),
.Y(n_459)
);

CKINVDCx20_ASAP7_75t_R g451 ( 
.A(n_412),
.Y(n_451)
);

CKINVDCx16_ASAP7_75t_R g452 ( 
.A(n_414),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_L g484 ( 
.A(n_452),
.B(n_454),
.Y(n_484)
);

AOI22xp33_ASAP7_75t_SL g453 ( 
.A1(n_401),
.A2(n_369),
.B1(n_315),
.B2(n_365),
.Y(n_453)
);

INVxp67_ASAP7_75t_L g457 ( 
.A(n_453),
.Y(n_457)
);

CKINVDCx20_ASAP7_75t_R g454 ( 
.A(n_412),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_397),
.Y(n_455)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_455),
.Y(n_482)
);

OAI22xp5_ASAP7_75t_L g512 ( 
.A1(n_460),
.A2(n_419),
.B1(n_455),
.B2(n_433),
.Y(n_512)
);

BUFx12f_ASAP7_75t_SL g492 ( 
.A(n_461),
.Y(n_492)
);

MAJIxp5_ASAP7_75t_L g493 ( 
.A(n_463),
.B(n_474),
.C(n_487),
.Y(n_493)
);

AOI22xp5_ASAP7_75t_L g467 ( 
.A1(n_430),
.A2(n_413),
.B1(n_386),
.B2(n_388),
.Y(n_467)
);

OAI22xp5_ASAP7_75t_SL g502 ( 
.A1(n_467),
.A2(n_472),
.B1(n_479),
.B2(n_485),
.Y(n_502)
);

CKINVDCx20_ASAP7_75t_R g470 ( 
.A(n_432),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_SL g495 ( 
.A(n_470),
.B(n_471),
.Y(n_495)
);

CKINVDCx20_ASAP7_75t_R g471 ( 
.A(n_439),
.Y(n_471)
);

AOI22xp5_ASAP7_75t_L g472 ( 
.A1(n_430),
.A2(n_413),
.B1(n_386),
.B2(n_416),
.Y(n_472)
);

AOI21xp5_ASAP7_75t_L g473 ( 
.A1(n_425),
.A2(n_394),
.B(n_414),
.Y(n_473)
);

AOI21xp5_ASAP7_75t_L g515 ( 
.A1(n_473),
.A2(n_434),
.B(n_389),
.Y(n_515)
);

MAJIxp5_ASAP7_75t_L g474 ( 
.A(n_429),
.B(n_422),
.C(n_421),
.Y(n_474)
);

XNOR2xp5_ASAP7_75t_L g475 ( 
.A(n_431),
.B(n_421),
.Y(n_475)
);

XOR2xp5_ASAP7_75t_L g505 ( 
.A(n_475),
.B(n_481),
.Y(n_505)
);

OAI22xp5_ASAP7_75t_SL g477 ( 
.A1(n_444),
.A2(n_394),
.B1(n_411),
.B2(n_403),
.Y(n_477)
);

AOI22xp5_ASAP7_75t_L g490 ( 
.A1(n_477),
.A2(n_456),
.B1(n_452),
.B2(n_447),
.Y(n_490)
);

INVxp67_ASAP7_75t_L g489 ( 
.A(n_478),
.Y(n_489)
);

AOI22xp5_ASAP7_75t_L g479 ( 
.A1(n_423),
.A2(n_444),
.B1(n_436),
.B2(n_427),
.Y(n_479)
);

INVxp67_ASAP7_75t_L g480 ( 
.A(n_445),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_L g499 ( 
.A(n_480),
.B(n_390),
.Y(n_499)
);

XOR2xp5_ASAP7_75t_L g481 ( 
.A(n_428),
.B(n_409),
.Y(n_481)
);

OAI21xp5_ASAP7_75t_L g483 ( 
.A1(n_447),
.A2(n_405),
.B(n_401),
.Y(n_483)
);

OAI21xp5_ASAP7_75t_L g497 ( 
.A1(n_483),
.A2(n_450),
.B(n_424),
.Y(n_497)
);

AOI22xp5_ASAP7_75t_L g485 ( 
.A1(n_423),
.A2(n_416),
.B1(n_411),
.B2(n_408),
.Y(n_485)
);

XNOR2xp5_ASAP7_75t_L g487 ( 
.A(n_428),
.B(n_408),
.Y(n_487)
);

AOI22xp5_ASAP7_75t_L g488 ( 
.A1(n_456),
.A2(n_416),
.B1(n_400),
.B2(n_404),
.Y(n_488)
);

OAI22xp5_ASAP7_75t_SL g503 ( 
.A1(n_488),
.A2(n_441),
.B1(n_446),
.B2(n_448),
.Y(n_503)
);

OAI22xp5_ASAP7_75t_SL g531 ( 
.A1(n_490),
.A2(n_516),
.B1(n_482),
.B2(n_461),
.Y(n_531)
);

NOR2xp33_ASAP7_75t_SL g491 ( 
.A(n_476),
.B(n_440),
.Y(n_491)
);

CKINVDCx14_ASAP7_75t_R g521 ( 
.A(n_491),
.Y(n_521)
);

XNOR2x1_ASAP7_75t_SL g494 ( 
.A(n_487),
.B(n_435),
.Y(n_494)
);

XOR2xp5_ASAP7_75t_L g520 ( 
.A(n_494),
.B(n_484),
.Y(n_520)
);

NOR2xp33_ASAP7_75t_L g496 ( 
.A(n_462),
.B(n_406),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_L g522 ( 
.A(n_496),
.B(n_499),
.Y(n_522)
);

XOR2x2_ASAP7_75t_L g525 ( 
.A(n_497),
.B(n_498),
.Y(n_525)
);

XNOR2xp5_ASAP7_75t_SL g498 ( 
.A(n_481),
.B(n_443),
.Y(n_498)
);

NOR2xp33_ASAP7_75t_L g500 ( 
.A(n_466),
.B(n_406),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_L g524 ( 
.A(n_500),
.B(n_508),
.Y(n_524)
);

MAJIxp5_ASAP7_75t_L g501 ( 
.A(n_463),
.B(n_475),
.C(n_474),
.Y(n_501)
);

MAJIxp5_ASAP7_75t_L g519 ( 
.A(n_501),
.B(n_483),
.C(n_467),
.Y(n_519)
);

AOI22xp5_ASAP7_75t_L g518 ( 
.A1(n_503),
.A2(n_504),
.B1(n_512),
.B2(n_517),
.Y(n_518)
);

NAND5xp2_ASAP7_75t_L g504 ( 
.A(n_484),
.B(n_443),
.C(n_454),
.D(n_451),
.E(n_426),
.Y(n_504)
);

XNOR2xp5_ASAP7_75t_L g506 ( 
.A(n_469),
.B(n_442),
.Y(n_506)
);

XNOR2xp5_ASAP7_75t_L g532 ( 
.A(n_506),
.B(n_511),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_L g507 ( 
.A(n_464),
.B(n_437),
.Y(n_507)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_507),
.Y(n_540)
);

CKINVDCx14_ASAP7_75t_R g508 ( 
.A(n_464),
.Y(n_508)
);

NOR2xp33_ASAP7_75t_L g509 ( 
.A(n_458),
.B(n_326),
.Y(n_509)
);

AOI21xp5_ASAP7_75t_L g537 ( 
.A1(n_509),
.A2(n_513),
.B(n_515),
.Y(n_537)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_465),
.Y(n_510)
);

INVx2_ASAP7_75t_L g523 ( 
.A(n_510),
.Y(n_523)
);

XNOR2xp5_ASAP7_75t_L g511 ( 
.A(n_469),
.B(n_416),
.Y(n_511)
);

NOR2xp33_ASAP7_75t_L g513 ( 
.A(n_478),
.B(n_289),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_L g514 ( 
.A(n_465),
.B(n_449),
.Y(n_514)
);

XNOR2xp5_ASAP7_75t_L g541 ( 
.A(n_514),
.B(n_295),
.Y(n_541)
);

AOI22xp5_ASAP7_75t_L g516 ( 
.A1(n_477),
.A2(n_438),
.B1(n_400),
.B2(n_404),
.Y(n_516)
);

OAI22xp5_ASAP7_75t_SL g517 ( 
.A1(n_479),
.A2(n_419),
.B1(n_402),
.B2(n_389),
.Y(n_517)
);

MAJIxp5_ASAP7_75t_L g544 ( 
.A(n_519),
.B(n_538),
.C(n_515),
.Y(n_544)
);

XNOR2xp5_ASAP7_75t_SL g543 ( 
.A(n_520),
.B(n_533),
.Y(n_543)
);

OAI22xp5_ASAP7_75t_SL g526 ( 
.A1(n_495),
.A2(n_460),
.B1(n_457),
.B2(n_480),
.Y(n_526)
);

INVxp67_ASAP7_75t_L g552 ( 
.A(n_526),
.Y(n_552)
);

MAJIxp5_ASAP7_75t_L g527 ( 
.A(n_493),
.B(n_473),
.C(n_472),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_L g549 ( 
.A(n_527),
.B(n_530),
.Y(n_549)
);

AOI22xp5_ASAP7_75t_L g528 ( 
.A1(n_502),
.A2(n_457),
.B1(n_461),
.B2(n_485),
.Y(n_528)
);

OAI22xp5_ASAP7_75t_SL g561 ( 
.A1(n_528),
.A2(n_529),
.B1(n_535),
.B2(n_504),
.Y(n_561)
);

AOI22xp5_ASAP7_75t_L g529 ( 
.A1(n_502),
.A2(n_461),
.B1(n_488),
.B2(n_482),
.Y(n_529)
);

MAJIxp5_ASAP7_75t_L g530 ( 
.A(n_493),
.B(n_461),
.C(n_486),
.Y(n_530)
);

XOR2xp5_ASAP7_75t_L g559 ( 
.A(n_531),
.B(n_512),
.Y(n_559)
);

XOR2xp5_ASAP7_75t_L g533 ( 
.A(n_505),
.B(n_468),
.Y(n_533)
);

OAI22xp5_ASAP7_75t_SL g534 ( 
.A1(n_489),
.A2(n_459),
.B1(n_402),
.B2(n_392),
.Y(n_534)
);

HB1xp67_ASAP7_75t_L g553 ( 
.A(n_534),
.Y(n_553)
);

AOI22xp5_ASAP7_75t_L g535 ( 
.A1(n_503),
.A2(n_459),
.B1(n_392),
.B2(n_376),
.Y(n_535)
);

XOR2xp5_ASAP7_75t_L g536 ( 
.A(n_505),
.B(n_287),
.Y(n_536)
);

XNOR2xp5_ASAP7_75t_SL g545 ( 
.A(n_536),
.B(n_539),
.Y(n_545)
);

MAJIxp5_ASAP7_75t_L g538 ( 
.A(n_501),
.B(n_341),
.C(n_306),
.Y(n_538)
);

XOR2xp5_ASAP7_75t_L g539 ( 
.A(n_506),
.B(n_289),
.Y(n_539)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_541),
.Y(n_542)
);

MAJIxp5_ASAP7_75t_L g570 ( 
.A(n_544),
.B(n_546),
.C(n_556),
.Y(n_570)
);

MAJIxp5_ASAP7_75t_L g546 ( 
.A(n_530),
.B(n_489),
.C(n_498),
.Y(n_546)
);

OAI21xp5_ASAP7_75t_SL g547 ( 
.A1(n_527),
.A2(n_492),
.B(n_507),
.Y(n_547)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_547),
.Y(n_564)
);

OAI22xp5_ASAP7_75t_SL g548 ( 
.A1(n_522),
.A2(n_491),
.B1(n_510),
.B2(n_516),
.Y(n_548)
);

NOR2xp33_ASAP7_75t_L g578 ( 
.A(n_548),
.B(n_558),
.Y(n_578)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_524),
.Y(n_550)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_550),
.Y(n_562)
);

NOR2xp33_ASAP7_75t_L g551 ( 
.A(n_521),
.B(n_490),
.Y(n_551)
);

NOR2xp33_ASAP7_75t_SL g573 ( 
.A(n_551),
.B(n_560),
.Y(n_573)
);

OR2x2_ASAP7_75t_L g554 ( 
.A(n_540),
.B(n_514),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_L g563 ( 
.A(n_554),
.B(n_518),
.Y(n_563)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_523),
.Y(n_555)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_555),
.Y(n_571)
);

MAJIxp5_ASAP7_75t_L g556 ( 
.A(n_538),
.B(n_511),
.C(n_497),
.Y(n_556)
);

MAJIxp5_ASAP7_75t_L g557 ( 
.A(n_519),
.B(n_494),
.C(n_499),
.Y(n_557)
);

MAJIxp5_ASAP7_75t_L g575 ( 
.A(n_557),
.B(n_545),
.C(n_544),
.Y(n_575)
);

XNOR2xp5_ASAP7_75t_L g558 ( 
.A(n_533),
.B(n_517),
.Y(n_558)
);

XOR2xp5_ASAP7_75t_L g567 ( 
.A(n_559),
.B(n_560),
.Y(n_567)
);

XNOR2xp5_ASAP7_75t_L g560 ( 
.A(n_532),
.B(n_504),
.Y(n_560)
);

AOI22xp5_ASAP7_75t_L g572 ( 
.A1(n_561),
.A2(n_520),
.B1(n_525),
.B2(n_534),
.Y(n_572)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_563),
.Y(n_583)
);

OAI21xp33_ASAP7_75t_L g565 ( 
.A1(n_549),
.A2(n_492),
.B(n_525),
.Y(n_565)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_565),
.Y(n_589)
);

OAI22xp5_ASAP7_75t_SL g566 ( 
.A1(n_552),
.A2(n_518),
.B1(n_528),
.B2(n_529),
.Y(n_566)
);

AOI22xp5_ASAP7_75t_L g579 ( 
.A1(n_566),
.A2(n_569),
.B1(n_559),
.B2(n_557),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_L g568 ( 
.A(n_554),
.B(n_541),
.Y(n_568)
);

AOI21xp33_ASAP7_75t_L g591 ( 
.A1(n_568),
.A2(n_577),
.B(n_1),
.Y(n_591)
);

OAI22xp5_ASAP7_75t_SL g569 ( 
.A1(n_552),
.A2(n_535),
.B1(n_537),
.B2(n_531),
.Y(n_569)
);

OAI22xp5_ASAP7_75t_SL g586 ( 
.A1(n_572),
.A2(n_574),
.B1(n_543),
.B2(n_545),
.Y(n_586)
);

AOI21xp5_ASAP7_75t_L g581 ( 
.A1(n_573),
.A2(n_546),
.B(n_558),
.Y(n_581)
);

AOI22xp5_ASAP7_75t_L g574 ( 
.A1(n_561),
.A2(n_539),
.B1(n_536),
.B2(n_532),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_SL g580 ( 
.A(n_575),
.B(n_576),
.Y(n_580)
);

MAJIxp5_ASAP7_75t_L g576 ( 
.A(n_556),
.B(n_295),
.C(n_224),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_L g577 ( 
.A(n_553),
.B(n_224),
.Y(n_577)
);

OAI22xp5_ASAP7_75t_SL g593 ( 
.A1(n_579),
.A2(n_588),
.B1(n_571),
.B2(n_574),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_581),
.Y(n_594)
);

NOR2xp67_ASAP7_75t_L g582 ( 
.A(n_564),
.B(n_542),
.Y(n_582)
);

AOI21xp5_ASAP7_75t_L g595 ( 
.A1(n_582),
.A2(n_562),
.B(n_563),
.Y(n_595)
);

XNOR2x1_ASAP7_75t_L g584 ( 
.A(n_572),
.B(n_543),
.Y(n_584)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_584),
.Y(n_597)
);

NOR2xp33_ASAP7_75t_SL g585 ( 
.A(n_562),
.B(n_570),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_SL g592 ( 
.A(n_585),
.B(n_578),
.Y(n_592)
);

NOR2xp33_ASAP7_75t_L g599 ( 
.A(n_586),
.B(n_567),
.Y(n_599)
);

XNOR2xp5_ASAP7_75t_L g587 ( 
.A(n_570),
.B(n_24),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_L g598 ( 
.A(n_587),
.B(n_590),
.Y(n_598)
);

AOI22xp5_ASAP7_75t_L g588 ( 
.A1(n_566),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_588)
);

MAJIxp5_ASAP7_75t_L g590 ( 
.A(n_575),
.B(n_1),
.C(n_5),
.Y(n_590)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_591),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_L g608 ( 
.A(n_592),
.B(n_593),
.Y(n_608)
);

AOI21xp5_ASAP7_75t_L g606 ( 
.A1(n_595),
.A2(n_600),
.B(n_590),
.Y(n_606)
);

CKINVDCx20_ASAP7_75t_R g596 ( 
.A(n_588),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_SL g602 ( 
.A(n_596),
.B(n_599),
.Y(n_602)
);

AOI21xp5_ASAP7_75t_L g600 ( 
.A1(n_589),
.A2(n_568),
.B(n_567),
.Y(n_600)
);

AND2x2_ASAP7_75t_L g603 ( 
.A(n_594),
.B(n_580),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_SL g610 ( 
.A(n_603),
.B(n_604),
.Y(n_610)
);

AND2x2_ASAP7_75t_L g604 ( 
.A(n_597),
.B(n_579),
.Y(n_604)
);

MAJIxp5_ASAP7_75t_L g605 ( 
.A(n_600),
.B(n_581),
.C(n_583),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_SL g611 ( 
.A(n_605),
.B(n_606),
.Y(n_611)
);

OR2x2_ASAP7_75t_L g607 ( 
.A(n_601),
.B(n_587),
.Y(n_607)
);

OAI21xp5_ASAP7_75t_SL g609 ( 
.A1(n_607),
.A2(n_576),
.B(n_571),
.Y(n_609)
);

MAJIxp5_ASAP7_75t_L g613 ( 
.A(n_609),
.B(n_612),
.C(n_602),
.Y(n_613)
);

MAJIxp5_ASAP7_75t_L g612 ( 
.A(n_608),
.B(n_593),
.C(n_584),
.Y(n_612)
);

OAI21xp5_ASAP7_75t_L g615 ( 
.A1(n_613),
.A2(n_614),
.B(n_610),
.Y(n_615)
);

MAJIxp5_ASAP7_75t_L g614 ( 
.A(n_611),
.B(n_569),
.C(n_577),
.Y(n_614)
);

AOI22xp5_ASAP7_75t_L g616 ( 
.A1(n_615),
.A2(n_586),
.B1(n_598),
.B2(n_6),
.Y(n_616)
);

MAJIxp5_ASAP7_75t_L g617 ( 
.A(n_616),
.B(n_1),
.C(n_5),
.Y(n_617)
);

A2O1A1Ixp33_ASAP7_75t_SL g618 ( 
.A1(n_617),
.A2(n_6),
.B(n_7),
.C(n_606),
.Y(n_618)
);

MAJIxp5_ASAP7_75t_L g619 ( 
.A(n_618),
.B(n_6),
.C(n_7),
.Y(n_619)
);

AO21x1_ASAP7_75t_L g620 ( 
.A1(n_619),
.A2(n_7),
.B(n_564),
.Y(n_620)
);


endmodule