module fake_jpeg_2472_n_557 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_557);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_557;

wire n_529;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_19;
wire n_182;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_547;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_541;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_11),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_16),
.Y(n_21)
);

INVxp67_ASAP7_75t_L g22 ( 
.A(n_14),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

BUFx10_ASAP7_75t_L g26 ( 
.A(n_16),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_10),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_4),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_9),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_15),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_9),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_11),
.Y(n_33)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_2),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_18),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_4),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_0),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_6),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_SL g39 ( 
.A(n_8),
.B(n_2),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_1),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_18),
.Y(n_41)
);

INVx11_ASAP7_75t_L g42 ( 
.A(n_11),
.Y(n_42)
);

INVx6_ASAP7_75t_SL g43 ( 
.A(n_3),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_1),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_7),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_11),
.Y(n_46)
);

BUFx16f_ASAP7_75t_L g47 ( 
.A(n_15),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_15),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_4),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_14),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_0),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_18),
.Y(n_52)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_4),
.Y(n_53)
);

INVx13_ASAP7_75t_L g54 ( 
.A(n_0),
.Y(n_54)
);

INVx13_ASAP7_75t_L g55 ( 
.A(n_8),
.Y(n_55)
);

INVx11_ASAP7_75t_L g56 ( 
.A(n_0),
.Y(n_56)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_52),
.Y(n_57)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_57),
.Y(n_131)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_47),
.Y(n_58)
);

INVx2_ASAP7_75t_SL g128 ( 
.A(n_58),
.Y(n_128)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_52),
.Y(n_59)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_59),
.Y(n_137)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_47),
.Y(n_60)
);

INVx2_ASAP7_75t_SL g198 ( 
.A(n_60),
.Y(n_198)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_43),
.Y(n_61)
);

INVx5_ASAP7_75t_L g133 ( 
.A(n_61),
.Y(n_133)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_43),
.Y(n_62)
);

BUFx2_ASAP7_75t_L g135 ( 
.A(n_62),
.Y(n_135)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_52),
.Y(n_63)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_63),
.Y(n_154)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_52),
.Y(n_64)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_64),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_39),
.B(n_1),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_65),
.B(n_106),
.Y(n_199)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_36),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_66),
.Y(n_134)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_43),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g190 ( 
.A(n_67),
.Y(n_190)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_52),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g160 ( 
.A(n_68),
.Y(n_160)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_36),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g197 ( 
.A(n_69),
.Y(n_197)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_23),
.Y(n_70)
);

INVx4_ASAP7_75t_L g129 ( 
.A(n_70),
.Y(n_129)
);

AND2x2_ASAP7_75t_L g71 ( 
.A(n_47),
.B(n_16),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_71),
.B(n_92),
.Y(n_127)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_47),
.Y(n_72)
);

INVx3_ASAP7_75t_L g130 ( 
.A(n_72),
.Y(n_130)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_32),
.Y(n_73)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_73),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_36),
.Y(n_74)
);

INVx6_ASAP7_75t_L g191 ( 
.A(n_74),
.Y(n_191)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_33),
.Y(n_75)
);

INVx3_ASAP7_75t_L g166 ( 
.A(n_75),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_36),
.Y(n_76)
);

INVx6_ASAP7_75t_L g193 ( 
.A(n_76),
.Y(n_193)
);

BUFx5_ASAP7_75t_L g77 ( 
.A(n_21),
.Y(n_77)
);

INVx4_ASAP7_75t_L g155 ( 
.A(n_77),
.Y(n_155)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_33),
.Y(n_78)
);

INVx3_ASAP7_75t_L g180 ( 
.A(n_78),
.Y(n_180)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_32),
.Y(n_79)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_79),
.Y(n_179)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_32),
.Y(n_80)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_80),
.Y(n_141)
);

INVx5_ASAP7_75t_L g81 ( 
.A(n_53),
.Y(n_81)
);

INVx4_ASAP7_75t_L g196 ( 
.A(n_81),
.Y(n_196)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_32),
.Y(n_82)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_82),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_38),
.Y(n_83)
);

INVx6_ASAP7_75t_L g211 ( 
.A(n_83),
.Y(n_211)
);

INVx6_ASAP7_75t_L g84 ( 
.A(n_31),
.Y(n_84)
);

INVx8_ASAP7_75t_L g136 ( 
.A(n_84),
.Y(n_136)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_32),
.Y(n_85)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_85),
.Y(n_174)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_45),
.Y(n_86)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_86),
.Y(n_178)
);

BUFx4f_ASAP7_75t_L g87 ( 
.A(n_54),
.Y(n_87)
);

BUFx4f_ASAP7_75t_SL g165 ( 
.A(n_87),
.Y(n_165)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_23),
.Y(n_88)
);

INVx4_ASAP7_75t_L g204 ( 
.A(n_88),
.Y(n_204)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_45),
.Y(n_89)
);

AND2x2_ASAP7_75t_L g161 ( 
.A(n_89),
.B(n_96),
.Y(n_161)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_23),
.Y(n_90)
);

INVx4_ASAP7_75t_L g213 ( 
.A(n_90),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_39),
.B(n_17),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g206 ( 
.A(n_91),
.B(n_98),
.Y(n_206)
);

AND2x2_ASAP7_75t_L g92 ( 
.A(n_45),
.B(n_17),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_38),
.Y(n_93)
);

INVx6_ASAP7_75t_L g215 ( 
.A(n_93),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_31),
.A2(n_17),
.B1(n_14),
.B2(n_13),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_94),
.A2(n_101),
.B1(n_28),
.B2(n_46),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_38),
.Y(n_95)
);

INVx8_ASAP7_75t_L g209 ( 
.A(n_95),
.Y(n_209)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_45),
.Y(n_96)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_33),
.Y(n_97)
);

INVx3_ASAP7_75t_L g182 ( 
.A(n_97),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_22),
.B(n_13),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_35),
.B(n_13),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_99),
.B(n_105),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_38),
.Y(n_100)
);

BUFx12f_ASAP7_75t_L g149 ( 
.A(n_100),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_31),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_101)
);

INVx6_ASAP7_75t_L g102 ( 
.A(n_44),
.Y(n_102)
);

INVx3_ASAP7_75t_L g183 ( 
.A(n_102),
.Y(n_183)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_34),
.Y(n_103)
);

INVx3_ASAP7_75t_L g203 ( 
.A(n_103),
.Y(n_203)
);

INVx5_ASAP7_75t_L g104 ( 
.A(n_53),
.Y(n_104)
);

INVx3_ASAP7_75t_L g210 ( 
.A(n_104),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_35),
.B(n_2),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_48),
.B(n_3),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_44),
.Y(n_107)
);

BUFx12f_ASAP7_75t_L g171 ( 
.A(n_107),
.Y(n_171)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_45),
.Y(n_108)
);

AND2x2_ASAP7_75t_L g181 ( 
.A(n_108),
.B(n_111),
.Y(n_181)
);

BUFx5_ASAP7_75t_L g109 ( 
.A(n_21),
.Y(n_109)
);

BUFx8_ASAP7_75t_L g167 ( 
.A(n_109),
.Y(n_167)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_37),
.Y(n_110)
);

INVx3_ASAP7_75t_L g214 ( 
.A(n_110),
.Y(n_214)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_24),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_41),
.B(n_3),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_112),
.B(n_115),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_SL g113 ( 
.A(n_41),
.B(n_5),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_113),
.B(n_114),
.Y(n_132)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_48),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_24),
.B(n_27),
.Y(n_115)
);

BUFx3_ASAP7_75t_L g116 ( 
.A(n_37),
.Y(n_116)
);

BUFx12f_ASAP7_75t_L g212 ( 
.A(n_116),
.Y(n_212)
);

BUFx12f_ASAP7_75t_L g117 ( 
.A(n_53),
.Y(n_117)
);

INVx11_ASAP7_75t_L g159 ( 
.A(n_117),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_50),
.B(n_5),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_118),
.B(n_29),
.Y(n_152)
);

INVx11_ASAP7_75t_L g119 ( 
.A(n_54),
.Y(n_119)
);

INVx11_ASAP7_75t_L g187 ( 
.A(n_119),
.Y(n_187)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_44),
.Y(n_120)
);

NAND2x1_ASAP7_75t_SL g201 ( 
.A(n_120),
.B(n_121),
.Y(n_201)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_44),
.Y(n_121)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_25),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_122),
.B(n_27),
.Y(n_139)
);

INVx5_ASAP7_75t_L g123 ( 
.A(n_37),
.Y(n_123)
);

CKINVDCx16_ASAP7_75t_R g156 ( 
.A(n_123),
.Y(n_156)
);

BUFx12_ASAP7_75t_L g124 ( 
.A(n_26),
.Y(n_124)
);

BUFx16f_ASAP7_75t_L g151 ( 
.A(n_124),
.Y(n_151)
);

BUFx5_ASAP7_75t_L g125 ( 
.A(n_21),
.Y(n_125)
);

CKINVDCx12_ASAP7_75t_R g169 ( 
.A(n_125),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_51),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_126),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_139),
.B(n_146),
.Y(n_225)
);

AOI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_87),
.A2(n_56),
.B1(n_42),
.B2(n_51),
.Y(n_140)
);

OA22x2_ASAP7_75t_L g237 ( 
.A1(n_140),
.A2(n_188),
.B1(n_192),
.B2(n_194),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_91),
.B(n_98),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_SL g246 ( 
.A(n_142),
.B(n_143),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_65),
.B(n_118),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_112),
.B(n_115),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_144),
.B(n_147),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_106),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_71),
.B(n_50),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_L g150 ( 
.A1(n_66),
.A2(n_95),
.B1(n_121),
.B2(n_120),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g255 ( 
.A1(n_150),
.A2(n_168),
.B1(n_207),
.B2(n_194),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_SL g257 ( 
.A(n_152),
.B(n_195),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_92),
.B(n_25),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_153),
.B(n_158),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_74),
.B(n_40),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_61),
.B(n_29),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_162),
.B(n_164),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_76),
.B(n_40),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_62),
.B(n_28),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_170),
.B(n_172),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_117),
.B(n_30),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_126),
.B(n_30),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_173),
.B(n_177),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_69),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_175),
.B(n_189),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_102),
.B(n_46),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_83),
.B(n_20),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_184),
.B(n_185),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_93),
.B(n_20),
.Y(n_185)
);

OAI22xp33_ASAP7_75t_SL g186 ( 
.A1(n_100),
.A2(n_51),
.B1(n_56),
.B2(n_42),
.Y(n_186)
);

AOI22xp33_ASAP7_75t_L g235 ( 
.A1(n_186),
.A2(n_26),
.B1(n_7),
.B2(n_12),
.Y(n_235)
);

AOI22xp33_ASAP7_75t_SL g188 ( 
.A1(n_107),
.A2(n_56),
.B1(n_42),
.B2(n_19),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_124),
.B(n_49),
.Y(n_189)
);

AOI22xp33_ASAP7_75t_SL g192 ( 
.A1(n_67),
.A2(n_19),
.B1(n_49),
.B2(n_55),
.Y(n_192)
);

AOI22xp33_ASAP7_75t_SL g194 ( 
.A1(n_67),
.A2(n_19),
.B1(n_54),
.B2(n_55),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_91),
.B(n_5),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_115),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_SL g265 ( 
.A(n_200),
.B(n_202),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_91),
.B(n_5),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_91),
.B(n_6),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g279 ( 
.A(n_205),
.B(n_208),
.Y(n_279)
);

AOI22xp33_ASAP7_75t_SL g207 ( 
.A1(n_67),
.A2(n_55),
.B1(n_34),
.B2(n_26),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_91),
.B(n_6),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_91),
.B(n_6),
.Y(n_216)
);

AOI21xp33_ASAP7_75t_L g251 ( 
.A1(n_216),
.A2(n_206),
.B(n_132),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_181),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_217),
.B(n_234),
.Y(n_309)
);

INVx3_ASAP7_75t_L g218 ( 
.A(n_133),
.Y(n_218)
);

BUFx2_ASAP7_75t_L g308 ( 
.A(n_218),
.Y(n_308)
);

FAx1_ASAP7_75t_SL g219 ( 
.A(n_148),
.B(n_26),
.CI(n_34),
.CON(n_219),
.SN(n_219)
);

FAx1_ASAP7_75t_SL g317 ( 
.A(n_219),
.B(n_261),
.CI(n_281),
.CON(n_317),
.SN(n_317)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_128),
.Y(n_220)
);

INVx1_ASAP7_75t_SL g310 ( 
.A(n_220),
.Y(n_310)
);

AOI22xp33_ASAP7_75t_SL g221 ( 
.A1(n_167),
.A2(n_26),
.B1(n_8),
.B2(n_10),
.Y(n_221)
);

INVxp67_ASAP7_75t_L g315 ( 
.A(n_221),
.Y(n_315)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_183),
.Y(n_222)
);

INVx4_ASAP7_75t_L g224 ( 
.A(n_159),
.Y(n_224)
);

INVx3_ASAP7_75t_L g297 ( 
.A(n_224),
.Y(n_297)
);

HB1xp67_ASAP7_75t_L g226 ( 
.A(n_166),
.Y(n_226)
);

INVxp67_ASAP7_75t_L g335 ( 
.A(n_226),
.Y(n_335)
);

INVx11_ASAP7_75t_L g227 ( 
.A(n_167),
.Y(n_227)
);

CKINVDCx16_ASAP7_75t_R g292 ( 
.A(n_227),
.Y(n_292)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_128),
.Y(n_228)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_228),
.Y(n_294)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_198),
.Y(n_229)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_229),
.Y(n_295)
);

INVx3_ASAP7_75t_L g230 ( 
.A(n_133),
.Y(n_230)
);

INVx3_ASAP7_75t_L g329 ( 
.A(n_230),
.Y(n_329)
);

INVx8_ASAP7_75t_L g231 ( 
.A(n_149),
.Y(n_231)
);

AOI22xp33_ASAP7_75t_SL g232 ( 
.A1(n_167),
.A2(n_26),
.B1(n_8),
.B2(n_10),
.Y(n_232)
);

AOI22xp33_ASAP7_75t_SL g299 ( 
.A1(n_232),
.A2(n_255),
.B1(n_261),
.B2(n_268),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_181),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_L g334 ( 
.A1(n_235),
.A2(n_239),
.B1(n_253),
.B2(n_259),
.Y(n_334)
);

OAI22xp33_ASAP7_75t_L g236 ( 
.A1(n_168),
.A2(n_7),
.B1(n_12),
.B2(n_188),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g302 ( 
.A1(n_236),
.A2(n_241),
.B1(n_250),
.B2(n_258),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_135),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_238),
.B(n_270),
.Y(n_318)
);

AOI22xp33_ASAP7_75t_L g239 ( 
.A1(n_186),
.A2(n_12),
.B1(n_145),
.B2(n_150),
.Y(n_239)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_183),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_199),
.A2(n_127),
.B1(n_207),
.B2(n_138),
.Y(n_241)
);

INVx4_ASAP7_75t_SL g242 ( 
.A(n_151),
.Y(n_242)
);

BUFx3_ASAP7_75t_L g336 ( 
.A(n_242),
.Y(n_336)
);

INVx8_ASAP7_75t_L g243 ( 
.A(n_149),
.Y(n_243)
);

INVx2_ASAP7_75t_L g325 ( 
.A(n_243),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_141),
.B(n_174),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_244),
.B(n_155),
.Y(n_301)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_166),
.Y(n_245)
);

INVx2_ASAP7_75t_L g339 ( 
.A(n_245),
.Y(n_339)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_198),
.Y(n_247)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_247),
.Y(n_296)
);

AND2x2_ASAP7_75t_L g249 ( 
.A(n_161),
.B(n_214),
.Y(n_249)
);

CKINVDCx16_ASAP7_75t_R g342 ( 
.A(n_249),
.Y(n_342)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_140),
.A2(n_197),
.B1(n_193),
.B2(n_211),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_SL g293 ( 
.A(n_251),
.B(n_190),
.Y(n_293)
);

INVx3_ASAP7_75t_L g252 ( 
.A(n_196),
.Y(n_252)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_252),
.Y(n_300)
);

AOI22xp33_ASAP7_75t_L g253 ( 
.A1(n_180),
.A2(n_214),
.B1(n_182),
.B2(n_134),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_157),
.Y(n_254)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_254),
.Y(n_306)
);

INVx8_ASAP7_75t_L g256 ( 
.A(n_149),
.Y(n_256)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_256),
.Y(n_311)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_197),
.A2(n_215),
.B1(n_211),
.B2(n_191),
.Y(n_258)
);

AOI22xp33_ASAP7_75t_L g259 ( 
.A1(n_180),
.A2(n_182),
.B1(n_134),
.B2(n_210),
.Y(n_259)
);

INVx5_ASAP7_75t_L g260 ( 
.A(n_212),
.Y(n_260)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_260),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_191),
.A2(n_215),
.B1(n_193),
.B2(n_192),
.Y(n_261)
);

BUFx6f_ASAP7_75t_L g262 ( 
.A(n_160),
.Y(n_262)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_262),
.Y(n_322)
);

AOI22xp33_ASAP7_75t_L g264 ( 
.A1(n_210),
.A2(n_201),
.B1(n_196),
.B2(n_178),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_SL g298 ( 
.A1(n_264),
.A2(n_155),
.B1(n_212),
.B2(n_190),
.Y(n_298)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_165),
.Y(n_266)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_266),
.Y(n_326)
);

INVx6_ASAP7_75t_L g267 ( 
.A(n_209),
.Y(n_267)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_267),
.Y(n_327)
);

OAI22xp5_ASAP7_75t_L g268 ( 
.A1(n_136),
.A2(n_209),
.B1(n_163),
.B2(n_131),
.Y(n_268)
);

BUFx6f_ASAP7_75t_L g269 ( 
.A(n_160),
.Y(n_269)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_269),
.Y(n_328)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_130),
.Y(n_270)
);

AND2x2_ASAP7_75t_L g271 ( 
.A(n_161),
.B(n_203),
.Y(n_271)
);

OAI21xp5_ASAP7_75t_SL g304 ( 
.A1(n_271),
.A2(n_272),
.B(n_282),
.Y(n_304)
);

OAI21xp33_ASAP7_75t_L g272 ( 
.A1(n_151),
.A2(n_203),
.B(n_130),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_151),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_273),
.B(n_275),
.Y(n_321)
);

INVx5_ASAP7_75t_L g274 ( 
.A(n_212),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g303 ( 
.A(n_274),
.Y(n_303)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_165),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_165),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_276),
.B(n_277),
.Y(n_324)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_176),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_201),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_280),
.B(n_283),
.Y(n_330)
);

OA22x2_ASAP7_75t_SL g281 ( 
.A1(n_169),
.A2(n_136),
.B1(n_159),
.B2(n_179),
.Y(n_281)
);

OA21x2_ASAP7_75t_L g305 ( 
.A1(n_281),
.A2(n_187),
.B(n_282),
.Y(n_305)
);

OAI21xp5_ASAP7_75t_L g282 ( 
.A1(n_129),
.A2(n_213),
.B(n_204),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_137),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_154),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g323 ( 
.A(n_284),
.Y(n_323)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_213),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g337 ( 
.A(n_287),
.Y(n_337)
);

INVxp67_ASAP7_75t_L g288 ( 
.A(n_187),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g340 ( 
.A(n_288),
.Y(n_340)
);

OAI22xp5_ASAP7_75t_L g289 ( 
.A1(n_129),
.A2(n_204),
.B1(n_156),
.B2(n_171),
.Y(n_289)
);

AOI22xp33_ASAP7_75t_SL g307 ( 
.A1(n_289),
.A2(n_290),
.B1(n_291),
.B2(n_227),
.Y(n_307)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_171),
.Y(n_290)
);

INVx2_ASAP7_75t_L g291 ( 
.A(n_171),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_SL g358 ( 
.A(n_293),
.B(n_274),
.Y(n_358)
);

AOI22xp33_ASAP7_75t_SL g374 ( 
.A1(n_298),
.A2(n_320),
.B1(n_308),
.B2(n_336),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_SL g346 ( 
.A(n_301),
.B(n_275),
.Y(n_346)
);

CKINVDCx9p33_ASAP7_75t_R g370 ( 
.A(n_305),
.Y(n_370)
);

INVxp33_ASAP7_75t_L g383 ( 
.A(n_307),
.Y(n_383)
);

AOI32xp33_ASAP7_75t_L g312 ( 
.A1(n_219),
.A2(n_278),
.A3(n_286),
.B1(n_248),
.B2(n_233),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g344 ( 
.A(n_312),
.B(n_218),
.Y(n_344)
);

OAI22xp5_ASAP7_75t_SL g314 ( 
.A1(n_219),
.A2(n_236),
.B1(n_241),
.B2(n_285),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_L g357 ( 
.A1(n_314),
.A2(n_331),
.B1(n_332),
.B2(n_260),
.Y(n_357)
);

OAI21xp5_ASAP7_75t_SL g316 ( 
.A1(n_271),
.A2(n_249),
.B(n_244),
.Y(n_316)
);

OAI21xp5_ASAP7_75t_SL g348 ( 
.A1(n_316),
.A2(n_317),
.B(n_252),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_279),
.B(n_225),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_319),
.B(n_333),
.Y(n_345)
);

AOI22xp33_ASAP7_75t_SL g320 ( 
.A1(n_250),
.A2(n_271),
.B1(n_237),
.B2(n_249),
.Y(n_320)
);

OAI22xp5_ASAP7_75t_SL g331 ( 
.A1(n_237),
.A2(n_265),
.B1(n_281),
.B2(n_263),
.Y(n_331)
);

OAI22xp5_ASAP7_75t_SL g332 ( 
.A1(n_237),
.A2(n_223),
.B1(n_257),
.B2(n_269),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_246),
.B(n_277),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_222),
.B(n_240),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_338),
.B(n_341),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_245),
.B(n_272),
.Y(n_341)
);

OAI22xp5_ASAP7_75t_SL g343 ( 
.A1(n_302),
.A2(n_237),
.B1(n_262),
.B2(n_230),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_343),
.B(n_346),
.Y(n_402)
);

XNOR2xp5_ASAP7_75t_SL g419 ( 
.A(n_344),
.B(n_365),
.Y(n_419)
);

OAI21xp5_ASAP7_75t_SL g401 ( 
.A1(n_348),
.A2(n_350),
.B(n_360),
.Y(n_401)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_338),
.Y(n_349)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_349),
.Y(n_389)
);

OAI21xp5_ASAP7_75t_L g350 ( 
.A1(n_330),
.A2(n_266),
.B(n_288),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_333),
.B(n_267),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_351),
.B(n_352),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_332),
.B(n_258),
.Y(n_352)
);

AOI22x1_ASAP7_75t_L g353 ( 
.A1(n_314),
.A2(n_291),
.B1(n_290),
.B2(n_242),
.Y(n_353)
);

OAI22xp5_ASAP7_75t_L g395 ( 
.A1(n_353),
.A2(n_368),
.B1(n_381),
.B2(n_292),
.Y(n_395)
);

AND2x2_ASAP7_75t_L g354 ( 
.A(n_342),
.B(n_301),
.Y(n_354)
);

INVxp67_ASAP7_75t_L g385 ( 
.A(n_354),
.Y(n_385)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_294),
.Y(n_355)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_355),
.Y(n_390)
);

CKINVDCx20_ASAP7_75t_R g356 ( 
.A(n_321),
.Y(n_356)
);

NOR2xp33_ASAP7_75t_L g396 ( 
.A(n_356),
.B(n_372),
.Y(n_396)
);

OAI22xp5_ASAP7_75t_SL g399 ( 
.A1(n_357),
.A2(n_308),
.B1(n_328),
.B2(n_322),
.Y(n_399)
);

INVxp67_ASAP7_75t_L g392 ( 
.A(n_358),
.Y(n_392)
);

NOR2xp33_ASAP7_75t_L g359 ( 
.A(n_319),
.B(n_224),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_SL g388 ( 
.A(n_359),
.B(n_363),
.Y(n_388)
);

AOI21xp5_ASAP7_75t_L g360 ( 
.A1(n_304),
.A2(n_231),
.B(n_243),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_331),
.B(n_256),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_361),
.B(n_364),
.Y(n_413)
);

AOI22xp5_ASAP7_75t_SL g362 ( 
.A1(n_315),
.A2(n_317),
.B1(n_293),
.B2(n_341),
.Y(n_362)
);

INVxp67_ASAP7_75t_L g397 ( 
.A(n_362),
.Y(n_397)
);

NOR2xp33_ASAP7_75t_L g363 ( 
.A(n_310),
.B(n_312),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_317),
.B(n_316),
.Y(n_364)
);

XNOR2xp5_ASAP7_75t_L g365 ( 
.A(n_309),
.B(n_306),
.Y(n_365)
);

MAJIxp5_ASAP7_75t_L g366 ( 
.A(n_306),
.B(n_304),
.C(n_294),
.Y(n_366)
);

XOR2xp5_ASAP7_75t_L g398 ( 
.A(n_366),
.B(n_376),
.Y(n_398)
);

NOR2xp33_ASAP7_75t_L g367 ( 
.A(n_310),
.B(n_337),
.Y(n_367)
);

NOR2xp33_ASAP7_75t_SL g409 ( 
.A(n_367),
.B(n_369),
.Y(n_409)
);

AOI22xp5_ASAP7_75t_L g368 ( 
.A1(n_302),
.A2(n_305),
.B1(n_334),
.B2(n_299),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_323),
.B(n_324),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_SL g371 ( 
.A(n_323),
.B(n_295),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_SL g411 ( 
.A(n_371),
.B(n_382),
.Y(n_411)
);

INVxp67_ASAP7_75t_L g372 ( 
.A(n_318),
.Y(n_372)
);

A2O1A1Ixp33_ASAP7_75t_L g373 ( 
.A1(n_305),
.A2(n_315),
.B(n_298),
.C(n_337),
.Y(n_373)
);

HB1xp67_ASAP7_75t_L g387 ( 
.A(n_373),
.Y(n_387)
);

AOI22xp33_ASAP7_75t_SL g406 ( 
.A1(n_374),
.A2(n_336),
.B1(n_308),
.B2(n_313),
.Y(n_406)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_295),
.Y(n_375)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_375),
.Y(n_405)
);

MAJIxp5_ASAP7_75t_L g376 ( 
.A(n_296),
.B(n_340),
.C(n_335),
.Y(n_376)
);

XOR2xp5_ASAP7_75t_L g377 ( 
.A(n_296),
.B(n_300),
.Y(n_377)
);

XOR2xp5_ASAP7_75t_L g403 ( 
.A(n_377),
.B(n_379),
.Y(n_403)
);

CKINVDCx20_ASAP7_75t_R g378 ( 
.A(n_335),
.Y(n_378)
);

NOR2xp33_ASAP7_75t_L g400 ( 
.A(n_378),
.B(n_384),
.Y(n_400)
);

MAJIxp5_ASAP7_75t_L g379 ( 
.A(n_340),
.B(n_326),
.C(n_300),
.Y(n_379)
);

AOI21xp5_ASAP7_75t_L g380 ( 
.A1(n_303),
.A2(n_326),
.B(n_297),
.Y(n_380)
);

BUFx12f_ASAP7_75t_L g418 ( 
.A(n_380),
.Y(n_418)
);

AOI22xp5_ASAP7_75t_L g381 ( 
.A1(n_327),
.A2(n_328),
.B1(n_322),
.B2(n_329),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_327),
.B(n_303),
.Y(n_382)
);

NOR2xp33_ASAP7_75t_L g384 ( 
.A(n_329),
.B(n_339),
.Y(n_384)
);

CKINVDCx20_ASAP7_75t_R g386 ( 
.A(n_371),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_386),
.B(n_391),
.Y(n_426)
);

CKINVDCx20_ASAP7_75t_R g391 ( 
.A(n_382),
.Y(n_391)
);

CKINVDCx20_ASAP7_75t_R g393 ( 
.A(n_384),
.Y(n_393)
);

NOR2xp33_ASAP7_75t_L g444 ( 
.A(n_393),
.B(n_394),
.Y(n_444)
);

CKINVDCx20_ASAP7_75t_R g394 ( 
.A(n_369),
.Y(n_394)
);

AOI22xp5_ASAP7_75t_L g420 ( 
.A1(n_395),
.A2(n_399),
.B1(n_373),
.B2(n_370),
.Y(n_420)
);

CKINVDCx20_ASAP7_75t_R g404 ( 
.A(n_367),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_SL g422 ( 
.A(n_404),
.B(n_408),
.Y(n_422)
);

OAI22xp5_ASAP7_75t_L g447 ( 
.A1(n_406),
.A2(n_378),
.B1(n_379),
.B2(n_350),
.Y(n_447)
);

INVx3_ASAP7_75t_L g407 ( 
.A(n_355),
.Y(n_407)
);

INVx2_ASAP7_75t_L g439 ( 
.A(n_407),
.Y(n_439)
);

CKINVDCx20_ASAP7_75t_R g408 ( 
.A(n_380),
.Y(n_408)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_375),
.Y(n_412)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_412),
.Y(n_429)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_349),
.Y(n_414)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_414),
.Y(n_433)
);

NOR2xp33_ASAP7_75t_L g415 ( 
.A(n_356),
.B(n_365),
.Y(n_415)
);

HB1xp67_ASAP7_75t_L g425 ( 
.A(n_415),
.Y(n_425)
);

INVx2_ASAP7_75t_L g416 ( 
.A(n_381),
.Y(n_416)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_416),
.Y(n_436)
);

CKINVDCx20_ASAP7_75t_R g417 ( 
.A(n_346),
.Y(n_417)
);

CKINVDCx20_ASAP7_75t_R g424 ( 
.A(n_417),
.Y(n_424)
);

OAI22xp5_ASAP7_75t_L g452 ( 
.A1(n_420),
.A2(n_432),
.B1(n_435),
.B2(n_447),
.Y(n_452)
);

OAI22xp5_ASAP7_75t_SL g421 ( 
.A1(n_387),
.A2(n_357),
.B1(n_368),
.B2(n_410),
.Y(n_421)
);

AOI22xp5_ASAP7_75t_L g465 ( 
.A1(n_421),
.A2(n_395),
.B1(n_410),
.B2(n_399),
.Y(n_465)
);

MAJIxp5_ASAP7_75t_L g423 ( 
.A(n_398),
.B(n_366),
.C(n_363),
.Y(n_423)
);

MAJIxp5_ASAP7_75t_L g458 ( 
.A(n_423),
.B(n_440),
.C(n_441),
.Y(n_458)
);

HB1xp67_ASAP7_75t_L g427 ( 
.A(n_396),
.Y(n_427)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_427),
.Y(n_461)
);

OAI21xp5_ASAP7_75t_SL g428 ( 
.A1(n_401),
.A2(n_362),
.B(n_348),
.Y(n_428)
);

OAI21xp5_ASAP7_75t_SL g451 ( 
.A1(n_428),
.A2(n_434),
.B(n_437),
.Y(n_451)
);

XNOR2xp5_ASAP7_75t_L g430 ( 
.A(n_398),
.B(n_364),
.Y(n_430)
);

XOR2xp5_ASAP7_75t_L g472 ( 
.A(n_430),
.B(n_431),
.Y(n_472)
);

XNOR2xp5_ASAP7_75t_L g431 ( 
.A(n_403),
.B(n_345),
.Y(n_431)
);

AOI22xp5_ASAP7_75t_L g432 ( 
.A1(n_402),
.A2(n_343),
.B1(n_361),
.B2(n_370),
.Y(n_432)
);

OAI21xp5_ASAP7_75t_L g434 ( 
.A1(n_401),
.A2(n_347),
.B(n_344),
.Y(n_434)
);

AOI22xp5_ASAP7_75t_L g435 ( 
.A1(n_402),
.A2(n_352),
.B1(n_373),
.B2(n_345),
.Y(n_435)
);

OAI21xp5_ASAP7_75t_L g437 ( 
.A1(n_397),
.A2(n_347),
.B(n_360),
.Y(n_437)
);

CKINVDCx16_ASAP7_75t_R g438 ( 
.A(n_400),
.Y(n_438)
);

NOR2xp33_ASAP7_75t_L g457 ( 
.A(n_438),
.B(n_445),
.Y(n_457)
);

XNOR2xp5_ASAP7_75t_L g440 ( 
.A(n_403),
.B(n_419),
.Y(n_440)
);

MAJIxp5_ASAP7_75t_L g441 ( 
.A(n_419),
.B(n_354),
.C(n_376),
.Y(n_441)
);

OAI21xp5_ASAP7_75t_L g442 ( 
.A1(n_413),
.A2(n_358),
.B(n_353),
.Y(n_442)
);

AOI21xp5_ASAP7_75t_L g454 ( 
.A1(n_442),
.A2(n_446),
.B(n_392),
.Y(n_454)
);

MAJIxp5_ASAP7_75t_L g443 ( 
.A(n_385),
.B(n_415),
.C(n_413),
.Y(n_443)
);

MAJIxp5_ASAP7_75t_L g460 ( 
.A(n_443),
.B(n_450),
.C(n_393),
.Y(n_460)
);

CKINVDCx20_ASAP7_75t_R g445 ( 
.A(n_400),
.Y(n_445)
);

OAI21xp5_ASAP7_75t_L g446 ( 
.A1(n_408),
.A2(n_353),
.B(n_351),
.Y(n_446)
);

A2O1A1O1Ixp25_ASAP7_75t_L g448 ( 
.A1(n_391),
.A2(n_354),
.B(n_359),
.C(n_377),
.D(n_383),
.Y(n_448)
);

XNOR2xp5_ASAP7_75t_SL g470 ( 
.A(n_448),
.B(n_389),
.Y(n_470)
);

CKINVDCx16_ASAP7_75t_R g449 ( 
.A(n_396),
.Y(n_449)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_449),
.Y(n_462)
);

XOR2xp5_ASAP7_75t_L g450 ( 
.A(n_388),
.B(n_354),
.Y(n_450)
);

CKINVDCx20_ASAP7_75t_R g453 ( 
.A(n_426),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g498 ( 
.A(n_453),
.B(n_455),
.Y(n_498)
);

INVxp67_ASAP7_75t_L g480 ( 
.A(n_454),
.Y(n_480)
);

INVx5_ASAP7_75t_L g455 ( 
.A(n_425),
.Y(n_455)
);

INVxp33_ASAP7_75t_L g456 ( 
.A(n_422),
.Y(n_456)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_456),
.Y(n_490)
);

CKINVDCx20_ASAP7_75t_R g459 ( 
.A(n_426),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_SL g484 ( 
.A(n_459),
.B(n_463),
.Y(n_484)
);

XNOR2xp5_ASAP7_75t_L g485 ( 
.A(n_460),
.B(n_467),
.Y(n_485)
);

NOR2xp33_ASAP7_75t_SL g463 ( 
.A(n_444),
.B(n_394),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_L g464 ( 
.A(n_424),
.B(n_386),
.Y(n_464)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_464),
.Y(n_491)
);

OAI22xp5_ASAP7_75t_L g481 ( 
.A1(n_465),
.A2(n_466),
.B1(n_468),
.B2(n_473),
.Y(n_481)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_433),
.Y(n_466)
);

MAJx2_ASAP7_75t_L g467 ( 
.A(n_440),
.B(n_388),
.C(n_409),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_433),
.Y(n_468)
);

CKINVDCx20_ASAP7_75t_R g469 ( 
.A(n_446),
.Y(n_469)
);

NOR2xp33_ASAP7_75t_L g478 ( 
.A(n_469),
.B(n_442),
.Y(n_478)
);

XOR2xp5_ASAP7_75t_L g479 ( 
.A(n_470),
.B(n_476),
.Y(n_479)
);

MAJIxp5_ASAP7_75t_L g471 ( 
.A(n_430),
.B(n_389),
.C(n_414),
.Y(n_471)
);

MAJIxp5_ASAP7_75t_L g486 ( 
.A(n_471),
.B(n_441),
.C(n_423),
.Y(n_486)
);

AOI22xp5_ASAP7_75t_L g473 ( 
.A1(n_421),
.A2(n_417),
.B1(n_404),
.B2(n_416),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_436),
.B(n_411),
.Y(n_474)
);

CKINVDCx20_ASAP7_75t_R g483 ( 
.A(n_474),
.Y(n_483)
);

AOI22xp5_ASAP7_75t_L g475 ( 
.A1(n_420),
.A2(n_411),
.B1(n_409),
.B2(n_418),
.Y(n_475)
);

OAI22xp5_ASAP7_75t_L g497 ( 
.A1(n_475),
.A2(n_477),
.B1(n_418),
.B2(n_412),
.Y(n_497)
);

XNOR2xp5_ASAP7_75t_L g476 ( 
.A(n_431),
.B(n_405),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_429),
.Y(n_477)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_478),
.Y(n_499)
);

AOI211xp5_ASAP7_75t_L g482 ( 
.A1(n_464),
.A2(n_434),
.B(n_448),
.C(n_443),
.Y(n_482)
);

OAI21xp33_ASAP7_75t_L g505 ( 
.A1(n_482),
.A2(n_451),
.B(n_457),
.Y(n_505)
);

XNOR2xp5_ASAP7_75t_L g503 ( 
.A(n_486),
.B(n_495),
.Y(n_503)
);

MAJIxp5_ASAP7_75t_L g487 ( 
.A(n_458),
.B(n_450),
.C(n_437),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_SL g506 ( 
.A(n_487),
.B(n_489),
.Y(n_506)
);

XOR2xp5_ASAP7_75t_L g488 ( 
.A(n_472),
.B(n_428),
.Y(n_488)
);

XOR2xp5_ASAP7_75t_L g510 ( 
.A(n_488),
.B(n_494),
.Y(n_510)
);

MAJIxp5_ASAP7_75t_L g489 ( 
.A(n_458),
.B(n_435),
.C(n_432),
.Y(n_489)
);

AOI22xp5_ASAP7_75t_L g492 ( 
.A1(n_452),
.A2(n_465),
.B1(n_473),
.B2(n_456),
.Y(n_492)
);

AOI22xp5_ASAP7_75t_L g500 ( 
.A1(n_492),
.A2(n_475),
.B1(n_454),
.B2(n_474),
.Y(n_500)
);

MAJIxp5_ASAP7_75t_L g493 ( 
.A(n_472),
.B(n_436),
.C(n_405),
.Y(n_493)
);

NOR2xp33_ASAP7_75t_L g501 ( 
.A(n_493),
.B(n_496),
.Y(n_501)
);

XOR2xp5_ASAP7_75t_L g494 ( 
.A(n_460),
.B(n_390),
.Y(n_494)
);

XNOR2xp5_ASAP7_75t_L g495 ( 
.A(n_471),
.B(n_390),
.Y(n_495)
);

MAJIxp5_ASAP7_75t_L g496 ( 
.A(n_476),
.B(n_467),
.C(n_451),
.Y(n_496)
);

AOI22xp33_ASAP7_75t_L g502 ( 
.A1(n_497),
.A2(n_461),
.B1(n_462),
.B2(n_455),
.Y(n_502)
);

OAI22xp5_ASAP7_75t_L g527 ( 
.A1(n_500),
.A2(n_502),
.B1(n_505),
.B2(n_509),
.Y(n_527)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_484),
.Y(n_504)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_504),
.Y(n_515)
);

XNOR2xp5_ASAP7_75t_L g507 ( 
.A(n_495),
.B(n_470),
.Y(n_507)
);

XNOR2xp5_ASAP7_75t_L g520 ( 
.A(n_507),
.B(n_514),
.Y(n_520)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_490),
.Y(n_508)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_508),
.Y(n_524)
);

AOI22xp33_ASAP7_75t_L g509 ( 
.A1(n_483),
.A2(n_462),
.B1(n_461),
.B2(n_477),
.Y(n_509)
);

NOR2x1_ASAP7_75t_L g511 ( 
.A(n_491),
.B(n_418),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_L g516 ( 
.A(n_511),
.B(n_513),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_L g512 ( 
.A(n_498),
.B(n_468),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_L g523 ( 
.A(n_512),
.B(n_493),
.Y(n_523)
);

NOR2xp33_ASAP7_75t_L g513 ( 
.A(n_494),
.B(n_466),
.Y(n_513)
);

XNOR2xp5_ASAP7_75t_SL g514 ( 
.A(n_488),
.B(n_418),
.Y(n_514)
);

AOI21xp5_ASAP7_75t_L g517 ( 
.A1(n_511),
.A2(n_480),
.B(n_492),
.Y(n_517)
);

NAND2xp33_ASAP7_75t_SL g528 ( 
.A(n_517),
.B(n_518),
.Y(n_528)
);

OAI21xp5_ASAP7_75t_L g518 ( 
.A1(n_500),
.A2(n_480),
.B(n_481),
.Y(n_518)
);

MAJIxp5_ASAP7_75t_L g519 ( 
.A(n_503),
.B(n_489),
.C(n_486),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_SL g529 ( 
.A(n_519),
.B(n_526),
.Y(n_529)
);

HB1xp67_ASAP7_75t_L g521 ( 
.A(n_499),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_L g537 ( 
.A(n_521),
.B(n_522),
.Y(n_537)
);

HB1xp67_ASAP7_75t_L g522 ( 
.A(n_503),
.Y(n_522)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_523),
.Y(n_533)
);

AOI22xp33_ASAP7_75t_SL g525 ( 
.A1(n_512),
.A2(n_439),
.B1(n_496),
.B2(n_505),
.Y(n_525)
);

OAI22xp5_ASAP7_75t_L g534 ( 
.A1(n_525),
.A2(n_507),
.B1(n_479),
.B2(n_510),
.Y(n_534)
);

NOR2xp33_ASAP7_75t_L g526 ( 
.A(n_501),
.B(n_485),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_SL g530 ( 
.A(n_515),
.B(n_506),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_L g539 ( 
.A(n_530),
.B(n_531),
.Y(n_539)
);

MAJIxp5_ASAP7_75t_L g531 ( 
.A(n_519),
.B(n_510),
.C(n_487),
.Y(n_531)
);

NOR2xp33_ASAP7_75t_L g532 ( 
.A(n_523),
.B(n_485),
.Y(n_532)
);

AOI21xp5_ASAP7_75t_L g542 ( 
.A1(n_532),
.A2(n_520),
.B(n_479),
.Y(n_542)
);

NAND2x1p5_ASAP7_75t_L g540 ( 
.A(n_534),
.B(n_527),
.Y(n_540)
);

CKINVDCx16_ASAP7_75t_R g535 ( 
.A(n_516),
.Y(n_535)
);

NOR2xp33_ASAP7_75t_L g538 ( 
.A(n_535),
.B(n_536),
.Y(n_538)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_524),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_L g547 ( 
.A(n_540),
.B(n_541),
.Y(n_547)
);

OA21x2_ASAP7_75t_SL g541 ( 
.A1(n_533),
.A2(n_517),
.B(n_537),
.Y(n_541)
);

AOI21xp33_ASAP7_75t_L g548 ( 
.A1(n_542),
.A2(n_531),
.B(n_514),
.Y(n_548)
);

AOI21xp5_ASAP7_75t_SL g543 ( 
.A1(n_533),
.A2(n_518),
.B(n_520),
.Y(n_543)
);

OAI21xp5_ASAP7_75t_SL g546 ( 
.A1(n_543),
.A2(n_528),
.B(n_536),
.Y(n_546)
);

NOR2xp33_ASAP7_75t_L g544 ( 
.A(n_529),
.B(n_439),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_SL g545 ( 
.A(n_544),
.B(n_537),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_L g550 ( 
.A(n_545),
.B(n_546),
.Y(n_550)
);

MAJIxp5_ASAP7_75t_L g551 ( 
.A(n_548),
.B(n_549),
.C(n_541),
.Y(n_551)
);

NOR2xp33_ASAP7_75t_L g549 ( 
.A(n_539),
.B(n_528),
.Y(n_549)
);

AOI31xp33_ASAP7_75t_L g553 ( 
.A1(n_551),
.A2(n_552),
.A3(n_311),
.B(n_313),
.Y(n_553)
);

OAI21xp5_ASAP7_75t_SL g552 ( 
.A1(n_547),
.A2(n_538),
.B(n_407),
.Y(n_552)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_553),
.Y(n_555)
);

OAI21x1_ASAP7_75t_SL g554 ( 
.A1(n_550),
.A2(n_311),
.B(n_325),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_SL g556 ( 
.A(n_555),
.B(n_554),
.Y(n_556)
);

AOI21xp5_ASAP7_75t_L g557 ( 
.A1(n_556),
.A2(n_325),
.B(n_297),
.Y(n_557)
);


endmodule