module fake_jpeg_29125_n_254 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_254);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_254;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_223;
wire n_187;
wire n_21;
wire n_57;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_155;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_4),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_11),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

BUFx2_ASAP7_75t_R g21 ( 
.A(n_5),
.Y(n_21)
);

INVx2_ASAP7_75t_R g22 ( 
.A(n_3),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_16),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_10),
.Y(n_25)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_10),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_1),
.Y(n_33)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_4),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_4),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_11),
.Y(n_36)
);

BUFx2_ASAP7_75t_L g37 ( 
.A(n_6),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_15),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_5),
.Y(n_39)
);

OR2x2_ASAP7_75t_L g40 ( 
.A(n_22),
.B(n_2),
.Y(n_40)
);

OR2x2_ASAP7_75t_L g86 ( 
.A(n_40),
.B(n_28),
.Y(n_86)
);

BUFx4f_ASAP7_75t_SL g41 ( 
.A(n_21),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g84 ( 
.A(n_41),
.Y(n_84)
);

BUFx5_ASAP7_75t_L g42 ( 
.A(n_21),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_42),
.Y(n_79)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_20),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_43),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_20),
.Y(n_44)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_44),
.Y(n_65)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_34),
.Y(n_45)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_45),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_SL g46 ( 
.A(n_22),
.B(n_15),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_46),
.B(n_52),
.Y(n_61)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_29),
.Y(n_47)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_47),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_20),
.Y(n_48)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_48),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g49 ( 
.A(n_22),
.B(n_2),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_49),
.B(n_19),
.Y(n_60)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_34),
.Y(n_50)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_50),
.Y(n_70)
);

INVx5_ASAP7_75t_L g51 ( 
.A(n_29),
.Y(n_51)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_51),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_24),
.B(n_14),
.Y(n_52)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_21),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_53),
.B(n_54),
.Y(n_62)
);

INVx13_ASAP7_75t_L g54 ( 
.A(n_34),
.Y(n_54)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_37),
.Y(n_55)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_55),
.Y(n_80)
);

INVx11_ASAP7_75t_L g56 ( 
.A(n_30),
.Y(n_56)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_56),
.Y(n_76)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_33),
.Y(n_57)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_57),
.Y(n_77)
);

BUFx5_ASAP7_75t_L g58 ( 
.A(n_30),
.Y(n_58)
);

AND2x2_ASAP7_75t_L g67 ( 
.A(n_58),
.B(n_39),
.Y(n_67)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_30),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_59),
.B(n_33),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_60),
.B(n_73),
.Y(n_104)
);

INVxp67_ASAP7_75t_L g111 ( 
.A(n_63),
.Y(n_111)
);

OAI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_43),
.A2(n_38),
.B1(n_37),
.B2(n_39),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_64),
.A2(n_71),
.B1(n_74),
.B2(n_58),
.Y(n_108)
);

AND2x2_ASAP7_75t_L g101 ( 
.A(n_67),
.B(n_81),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_53),
.A2(n_37),
.B1(n_26),
.B2(n_31),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_69),
.A2(n_51),
.B1(n_57),
.B2(n_31),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_56),
.A2(n_39),
.B1(n_36),
.B2(n_35),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_46),
.B(n_24),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_72),
.B(n_82),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_49),
.B(n_26),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_44),
.A2(n_36),
.B1(n_35),
.B2(n_38),
.Y(n_74)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_42),
.B(n_36),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_40),
.B(n_25),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_40),
.B(n_25),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_83),
.B(n_85),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_41),
.B(n_18),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_86),
.B(n_41),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_86),
.B(n_19),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_88),
.B(n_91),
.Y(n_141)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_87),
.Y(n_89)
);

INVx4_ASAP7_75t_L g128 ( 
.A(n_89),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_90),
.A2(n_96),
.B1(n_106),
.B2(n_112),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_60),
.B(n_28),
.Y(n_91)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_66),
.Y(n_92)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_92),
.Y(n_146)
);

BUFx8_ASAP7_75t_L g93 ( 
.A(n_84),
.Y(n_93)
);

BUFx2_ASAP7_75t_SL g138 ( 
.A(n_93),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_61),
.B(n_18),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_94),
.B(n_95),
.Y(n_152)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_66),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_73),
.A2(n_44),
.B1(n_48),
.B2(n_38),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_84),
.A2(n_53),
.B1(n_55),
.B2(n_31),
.Y(n_97)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_97),
.Y(n_129)
);

AO22x1_ASAP7_75t_L g98 ( 
.A1(n_85),
.A2(n_41),
.B1(n_53),
.B2(n_59),
.Y(n_98)
);

A2O1A1Ixp33_ASAP7_75t_L g145 ( 
.A1(n_98),
.A2(n_54),
.B(n_68),
.C(n_6),
.Y(n_145)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_70),
.Y(n_99)
);

INVxp67_ASAP7_75t_L g135 ( 
.A(n_99),
.Y(n_135)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_70),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g139 ( 
.A(n_100),
.Y(n_139)
);

BUFx2_ASAP7_75t_L g102 ( 
.A(n_75),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_102),
.B(n_116),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_62),
.B(n_23),
.Y(n_103)
);

OR2x2_ASAP7_75t_L g136 ( 
.A(n_103),
.B(n_107),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_84),
.A2(n_50),
.B1(n_45),
.B2(n_47),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_105),
.A2(n_68),
.B1(n_54),
.B2(n_6),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_81),
.A2(n_48),
.B1(n_35),
.B2(n_23),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_84),
.B(n_32),
.Y(n_107)
);

OA22x2_ASAP7_75t_L g143 ( 
.A1(n_108),
.A2(n_109),
.B1(n_115),
.B2(n_120),
.Y(n_143)
);

INVx8_ASAP7_75t_L g109 ( 
.A(n_87),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_81),
.B(n_77),
.C(n_67),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_110),
.B(n_80),
.C(n_76),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_74),
.A2(n_59),
.B1(n_47),
.B2(n_32),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_79),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_113),
.B(n_119),
.Y(n_127)
);

INVx6_ASAP7_75t_L g115 ( 
.A(n_65),
.Y(n_115)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_77),
.Y(n_116)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_76),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_117),
.B(n_121),
.Y(n_134)
);

OA22x2_ASAP7_75t_L g120 ( 
.A1(n_65),
.A2(n_59),
.B1(n_27),
.B2(n_17),
.Y(n_120)
);

INVx13_ASAP7_75t_L g121 ( 
.A(n_79),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_67),
.B(n_27),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_122),
.B(n_123),
.Y(n_137)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_78),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_75),
.B(n_17),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_124),
.B(n_125),
.Y(n_140)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_78),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_80),
.B(n_2),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_126),
.B(n_3),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_130),
.B(n_131),
.C(n_120),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_104),
.B(n_71),
.C(n_68),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_133),
.A2(n_148),
.B1(n_149),
.B2(n_12),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_142),
.B(n_150),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_SL g159 ( 
.A1(n_145),
.A2(n_101),
.B(n_111),
.Y(n_159)
);

AOI22xp33_ASAP7_75t_L g147 ( 
.A1(n_108),
.A2(n_3),
.B1(n_5),
.B2(n_7),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_147),
.A2(n_111),
.B1(n_120),
.B2(n_115),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_110),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_98),
.A2(n_7),
.B1(n_8),
.B2(n_11),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_126),
.B(n_8),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_101),
.B(n_12),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_151),
.B(n_93),
.Y(n_170)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_146),
.Y(n_153)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_153),
.Y(n_176)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_146),
.Y(n_154)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_154),
.Y(n_185)
);

XOR2xp5_ASAP7_75t_L g155 ( 
.A(n_130),
.B(n_118),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_L g181 ( 
.A(n_155),
.B(n_157),
.Y(n_181)
);

INVx6_ASAP7_75t_L g156 ( 
.A(n_128),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_156),
.B(n_165),
.Y(n_184)
);

XOR2x2_ASAP7_75t_L g157 ( 
.A(n_127),
.B(n_101),
.Y(n_157)
);

A2O1A1Ixp33_ASAP7_75t_L g158 ( 
.A1(n_151),
.A2(n_137),
.B(n_150),
.C(n_142),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_SL g175 ( 
.A1(n_158),
.A2(n_167),
.B(n_162),
.Y(n_175)
);

INVxp67_ASAP7_75t_L g183 ( 
.A(n_159),
.Y(n_183)
);

XOR2xp5_ASAP7_75t_L g174 ( 
.A(n_160),
.B(n_169),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_161),
.A2(n_163),
.B1(n_168),
.B2(n_144),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_144),
.A2(n_120),
.B1(n_112),
.B2(n_100),
.Y(n_163)
);

BUFx3_ASAP7_75t_L g164 ( 
.A(n_138),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_164),
.Y(n_177)
);

INVx3_ASAP7_75t_L g165 ( 
.A(n_138),
.Y(n_165)
);

OAI32xp33_ASAP7_75t_L g166 ( 
.A1(n_137),
.A2(n_114),
.A3(n_99),
.B1(n_95),
.B2(n_92),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_166),
.B(n_170),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_SL g167 ( 
.A1(n_145),
.A2(n_89),
.B(n_123),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_127),
.B(n_121),
.Y(n_169)
);

INVxp67_ASAP7_75t_L g171 ( 
.A(n_134),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_171),
.B(n_132),
.Y(n_187)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_128),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_172),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_136),
.B(n_152),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_SL g191 ( 
.A(n_173),
.B(n_141),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_175),
.B(n_186),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g178 ( 
.A(n_155),
.B(n_160),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_178),
.B(n_187),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_179),
.A2(n_180),
.B1(n_188),
.B2(n_143),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_168),
.A2(n_143),
.B1(n_131),
.B2(n_129),
.Y(n_180)
);

CKINVDCx16_ASAP7_75t_R g186 ( 
.A(n_172),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_L g188 ( 
.A1(n_161),
.A2(n_143),
.B1(n_140),
.B2(n_152),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_164),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_190),
.B(n_191),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_SL g192 ( 
.A1(n_183),
.A2(n_159),
.B(n_167),
.Y(n_192)
);

INVxp67_ASAP7_75t_L g218 ( 
.A(n_192),
.Y(n_218)
);

AOI21xp5_ASAP7_75t_SL g194 ( 
.A1(n_189),
.A2(n_157),
.B(n_169),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_194),
.B(n_201),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_183),
.A2(n_171),
.B1(n_133),
.B2(n_143),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g212 ( 
.A(n_196),
.B(n_156),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_SL g198 ( 
.A(n_175),
.B(n_166),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_198),
.B(n_200),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_187),
.B(n_136),
.Y(n_199)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_199),
.Y(n_216)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_176),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_176),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_SL g202 ( 
.A(n_181),
.B(n_141),
.Y(n_202)
);

NAND3xp33_ASAP7_75t_L g215 ( 
.A(n_202),
.B(n_203),
.C(n_205),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_SL g203 ( 
.A(n_181),
.B(n_140),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_185),
.B(n_136),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_204),
.Y(n_213)
);

NAND3xp33_ASAP7_75t_L g205 ( 
.A(n_185),
.B(n_134),
.C(n_158),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_206),
.A2(n_109),
.B1(n_102),
.B2(n_125),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_177),
.B(n_148),
.Y(n_207)
);

OAI322xp33_ASAP7_75t_L g210 ( 
.A1(n_207),
.A2(n_149),
.A3(n_190),
.B1(n_177),
.B2(n_143),
.C1(n_182),
.C2(n_184),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_195),
.B(n_178),
.C(n_174),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_208),
.B(n_209),
.C(n_199),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_195),
.B(n_174),
.C(n_132),
.Y(n_209)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_210),
.Y(n_222)
);

AOI321xp33_ASAP7_75t_L g211 ( 
.A1(n_194),
.A2(n_182),
.A3(n_93),
.B1(n_139),
.B2(n_135),
.C(n_165),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_211),
.B(n_193),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_212),
.A2(n_197),
.B1(n_198),
.B2(n_193),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_219),
.B(n_201),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_220),
.B(n_228),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_213),
.B(n_204),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_221),
.B(n_227),
.Y(n_230)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_208),
.B(n_209),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_223),
.B(n_224),
.Y(n_231)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_214),
.B(n_192),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_225),
.B(n_226),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_218),
.B(n_202),
.C(n_203),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_218),
.B(n_217),
.C(n_212),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_229),
.B(n_206),
.Y(n_237)
);

FAx1_ASAP7_75t_L g232 ( 
.A(n_224),
.B(n_215),
.CI(n_216),
.CON(n_232),
.SN(n_232)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_232),
.B(n_234),
.Y(n_238)
);

AOI22xp33_ASAP7_75t_SL g233 ( 
.A1(n_222),
.A2(n_196),
.B1(n_211),
.B2(n_219),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_233),
.A2(n_228),
.B1(n_200),
.B2(n_223),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_229),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_237),
.B(n_12),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_230),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_SL g244 ( 
.A(n_239),
.B(n_240),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_SL g246 ( 
.A(n_241),
.B(n_13),
.Y(n_246)
);

AOI21xp5_ASAP7_75t_L g242 ( 
.A1(n_232),
.A2(n_14),
.B(n_13),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_242),
.Y(n_243)
);

BUFx24_ASAP7_75t_SL g245 ( 
.A(n_238),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_245),
.B(n_246),
.Y(n_248)
);

AOI21xp5_ASAP7_75t_L g247 ( 
.A1(n_244),
.A2(n_235),
.B(n_236),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_SL g251 ( 
.A(n_247),
.B(n_231),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_243),
.B(n_240),
.C(n_241),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_249),
.B(n_242),
.Y(n_250)
);

AOI21xp5_ASAP7_75t_SL g252 ( 
.A1(n_250),
.A2(n_251),
.B(n_233),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_252),
.B(n_248),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_253),
.B(n_13),
.Y(n_254)
);


endmodule