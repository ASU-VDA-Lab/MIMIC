module real_jpeg_14913_n_14 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_2, n_13, n_6, n_7, n_3, n_10, n_9, n_14);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_2;
input n_13;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_14;

wire n_108;
wire n_54;
wire n_37;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_83;
wire n_78;
wire n_104;
wire n_64;
wire n_47;
wire n_131;
wire n_22;
wire n_87;
wire n_40;
wire n_105;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_126;
wire n_113;
wire n_120;
wire n_93;
wire n_95;
wire n_65;
wire n_33;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_66;
wire n_136;
wire n_44;
wire n_28;
wire n_62;
wire n_121;
wire n_106;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_69;
wire n_31;
wire n_129;
wire n_135;
wire n_134;
wire n_72;
wire n_100;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_117;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_30;
wire n_15;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_128;
wire n_133;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_101;
wire n_96;
wire n_89;
wire n_16;

BUFx2_ASAP7_75t_L g48 ( 
.A(n_0),
.Y(n_48)
);

BUFx4f_ASAP7_75t_L g73 ( 
.A(n_1),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g76 ( 
.A1(n_2),
.A2(n_23),
.B1(n_26),
.B2(n_77),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_2),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_2),
.A2(n_44),
.B1(n_47),
.B2(n_77),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_3),
.B(n_38),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_3),
.B(n_28),
.Y(n_59)
);

AOI21xp33_ASAP7_75t_SL g88 ( 
.A1(n_3),
.A2(n_28),
.B(n_59),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_3),
.B(n_44),
.C(n_71),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_3),
.A2(n_23),
.B1(n_26),
.B2(n_101),
.Y(n_100)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_3),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_3),
.A2(n_50),
.B1(n_51),
.B2(n_113),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_3),
.B(n_127),
.Y(n_126)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

BUFx12_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

AOI22xp33_ASAP7_75t_L g31 ( 
.A1(n_7),
.A2(n_28),
.B1(n_29),
.B2(n_32),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_7),
.A2(n_23),
.B1(n_26),
.B2(n_32),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_7),
.A2(n_32),
.B1(n_44),
.B2(n_47),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g43 ( 
.A1(n_8),
.A2(n_44),
.B1(n_46),
.B2(n_47),
.Y(n_43)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_8),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_L g52 ( 
.A1(n_9),
.A2(n_44),
.B1(n_47),
.B2(n_53),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_9),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_10),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_SL g33 ( 
.A1(n_11),
.A2(n_28),
.B1(n_29),
.B2(n_34),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_11),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_11),
.A2(n_23),
.B1(n_26),
.B2(n_34),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_L g105 ( 
.A1(n_11),
.A2(n_34),
.B1(n_44),
.B2(n_47),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_12),
.A2(n_44),
.B1(n_47),
.B2(n_64),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_12),
.Y(n_64)
);

OAI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_12),
.A2(n_23),
.B1(n_26),
.B2(n_64),
.Y(n_80)
);

INVx11_ASAP7_75t_L g45 ( 
.A(n_13),
.Y(n_45)
);

XNOR2xp5_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_92),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_91),
.Y(n_15)
);

INVxp67_ASAP7_75t_L g16 ( 
.A(n_17),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_SL g17 ( 
.A(n_18),
.B(n_83),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_18),
.B(n_83),
.Y(n_91)
);

XOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_55),
.Y(n_18)
);

XNOR2xp5_ASAP7_75t_SL g19 ( 
.A(n_20),
.B(n_35),
.Y(n_19)
);

OAI22xp5_ASAP7_75t_SL g20 ( 
.A1(n_21),
.A2(n_22),
.B1(n_31),
.B2(n_33),
.Y(n_20)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_21),
.A2(n_22),
.B1(n_31),
.B2(n_88),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g21 ( 
.A(n_22),
.B(n_27),
.Y(n_21)
);

CKINVDCx14_ASAP7_75t_R g127 ( 
.A(n_22),
.Y(n_127)
);

OA22x2_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_24),
.B1(n_25),
.B2(n_26),
.Y(n_22)
);

INVx4_ASAP7_75t_SL g26 ( 
.A(n_23),
.Y(n_26)
);

A2O1A1Ixp33_ASAP7_75t_L g57 ( 
.A1(n_23),
.A2(n_25),
.B(n_58),
.C(n_60),
.Y(n_57)
);

OAI22xp33_ASAP7_75t_L g70 ( 
.A1(n_23),
.A2(n_26),
.B1(n_71),
.B2(n_72),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_23),
.B(n_98),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g27 ( 
.A1(n_24),
.A2(n_25),
.B1(n_28),
.B2(n_29),
.Y(n_27)
);

NAND3xp33_ASAP7_75t_SL g60 ( 
.A(n_24),
.B(n_26),
.C(n_29),
.Y(n_60)
);

INVx8_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_L g39 ( 
.A1(n_28),
.A2(n_29),
.B1(n_40),
.B2(n_41),
.Y(n_39)
);

INVx5_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

AOI22xp5_ASAP7_75t_L g35 ( 
.A1(n_36),
.A2(n_37),
.B1(n_42),
.B2(n_54),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx1_ASAP7_75t_SL g41 ( 
.A(n_40),
.Y(n_41)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_42),
.Y(n_54)
);

AOI21xp5_ASAP7_75t_L g42 ( 
.A1(n_43),
.A2(n_48),
.B(n_49),
.Y(n_42)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_44),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_44),
.B(n_51),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_44),
.A2(n_47),
.B1(n_71),
.B2(n_72),
.Y(n_74)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_47),
.B(n_111),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_48),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_48),
.A2(n_65),
.B1(n_104),
.B2(n_106),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_48),
.B(n_63),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_50),
.B(n_52),
.Y(n_49)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_50),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_50),
.A2(n_51),
.B1(n_105),
.B2(n_113),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_L g122 ( 
.A1(n_50),
.A2(n_107),
.B(n_123),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_51),
.B(n_52),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_SL g111 ( 
.A(n_51),
.B(n_101),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_56),
.A2(n_67),
.B1(n_81),
.B2(n_82),
.Y(n_55)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_56),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_57),
.B(n_61),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_57),
.A2(n_61),
.B1(n_62),
.B2(n_85),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_57),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

AOI21xp5_ASAP7_75t_L g62 ( 
.A1(n_63),
.A2(n_65),
.B(n_66),
.Y(n_62)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_67),
.Y(n_82)
);

OAI21xp5_ASAP7_75t_SL g67 ( 
.A1(n_68),
.A2(n_75),
.B(n_78),
.Y(n_67)
);

CKINVDCx16_ASAP7_75t_R g68 ( 
.A(n_69),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_69),
.A2(n_76),
.B1(n_79),
.B2(n_90),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_69),
.A2(n_79),
.B1(n_100),
.B2(n_102),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_69),
.A2(n_79),
.B1(n_90),
.B2(n_102),
.Y(n_128)
);

AND2x2_ASAP7_75t_L g69 ( 
.A(n_70),
.B(n_74),
.Y(n_69)
);

CKINVDCx14_ASAP7_75t_SL g71 ( 
.A(n_72),
.Y(n_71)
);

INVx13_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_74),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_74),
.B(n_101),
.Y(n_116)
);

CKINVDCx16_ASAP7_75t_R g75 ( 
.A(n_76),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_79),
.B(n_80),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_84),
.B(n_86),
.C(n_89),
.Y(n_83)
);

XOR2xp5_ASAP7_75t_L g132 ( 
.A(n_84),
.B(n_133),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_86),
.A2(n_87),
.B1(n_89),
.B2(n_134),
.Y(n_133)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_89),
.Y(n_134)
);

AOI21xp5_ASAP7_75t_SL g92 ( 
.A1(n_93),
.A2(n_131),
.B(n_136),
.Y(n_92)
);

OAI21xp5_ASAP7_75t_L g93 ( 
.A1(n_94),
.A2(n_119),
.B(n_130),
.Y(n_93)
);

AOI21xp5_ASAP7_75t_L g94 ( 
.A1(n_95),
.A2(n_108),
.B(n_118),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_96),
.B(n_103),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_96),
.B(n_103),
.Y(n_118)
);

XNOR2xp5_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_99),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_97),
.B(n_99),
.Y(n_120)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_L g108 ( 
.A1(n_109),
.A2(n_114),
.B(n_117),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_110),
.B(n_112),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_115),
.B(n_116),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_115),
.B(n_116),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_120),
.B(n_121),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_120),
.B(n_121),
.Y(n_130)
);

XNOR2xp5_ASAP7_75t_L g121 ( 
.A(n_122),
.B(n_124),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_122),
.B(n_125),
.C(n_129),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_125),
.A2(n_126),
.B1(n_128),
.B2(n_129),
.Y(n_124)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_128),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_132),
.B(n_135),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_132),
.B(n_135),
.Y(n_136)
);


endmodule