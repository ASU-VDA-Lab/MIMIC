module real_jpeg_21967_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_233;
wire n_37;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_83;
wire n_78;
wire n_249;
wire n_166;
wire n_176;
wire n_215;
wire n_221;
wire n_104;
wire n_194;
wire n_153;
wire n_161;
wire n_207;
wire n_280;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_281;
wire n_271;
wire n_163;
wire n_276;
wire n_22;
wire n_237;
wire n_174;
wire n_87;
wire n_197;
wire n_105;
wire n_40;
wire n_173;
wire n_243;
wire n_255;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_200;
wire n_48;
wire n_184;
wire n_164;
wire n_275;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_120;
wire n_113;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_282;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_44;
wire n_28;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_262;
wire n_222;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_223;
wire n_159;
wire n_72;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_203;
wire n_192;
wire n_100;
wire n_198;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_195;
wire n_110;
wire n_205;
wire n_258;
wire n_117;
wire n_193;
wire n_99;
wire n_261;
wire n_86;
wire n_150;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_70;
wire n_228;
wire n_30;
wire n_204;
wire n_158;
wire n_149;
wire n_278;
wire n_130;
wire n_144;
wire n_241;
wire n_103;
wire n_225;
wire n_259;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_277;
wire n_226;
wire n_125;
wire n_240;
wire n_185;
wire n_209;
wire n_55;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_279;
wire n_167;
wire n_128;
wire n_213;
wire n_179;
wire n_244;
wire n_216;
wire n_133;
wire n_202;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_283;
wire n_101;
wire n_274;
wire n_256;
wire n_182;
wire n_273;
wire n_96;
wire n_253;
wire n_269;
wire n_89;

OAI22xp5_ASAP7_75t_SL g26 ( 
.A1(n_0),
.A2(n_27),
.B1(n_29),
.B2(n_30),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_0),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_0),
.A2(n_29),
.B1(n_33),
.B2(n_34),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_0),
.A2(n_29),
.B1(n_75),
.B2(n_80),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_0),
.A2(n_29),
.B1(n_46),
.B2(n_47),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_1),
.A2(n_75),
.B1(n_80),
.B2(n_97),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_1),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_1),
.A2(n_46),
.B1(n_47),
.B2(n_97),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_SL g196 ( 
.A1(n_1),
.A2(n_33),
.B1(n_34),
.B2(n_97),
.Y(n_196)
);

AOI22xp33_ASAP7_75t_SL g240 ( 
.A1(n_1),
.A2(n_27),
.B1(n_30),
.B2(n_97),
.Y(n_240)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_2),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_2),
.B(n_77),
.Y(n_178)
);

AOI21xp33_ASAP7_75t_L g200 ( 
.A1(n_2),
.A2(n_14),
.B(n_34),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_2),
.A2(n_27),
.B1(n_30),
.B2(n_150),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_L g211 ( 
.A1(n_2),
.A2(n_60),
.B1(n_122),
.B2(n_209),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_2),
.B(n_182),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_2),
.B(n_46),
.Y(n_233)
);

AOI21xp33_ASAP7_75t_L g237 ( 
.A1(n_2),
.A2(n_46),
.B(n_233),
.Y(n_237)
);

OAI22xp33_ASAP7_75t_SL g37 ( 
.A1(n_3),
.A2(n_27),
.B1(n_30),
.B2(n_38),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_3),
.Y(n_38)
);

OAI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_3),
.A2(n_38),
.B1(n_75),
.B2(n_80),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_L g90 ( 
.A1(n_3),
.A2(n_33),
.B1(n_34),
.B2(n_38),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_L g104 ( 
.A1(n_3),
.A2(n_38),
.B1(n_46),
.B2(n_47),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_4),
.A2(n_46),
.B1(n_47),
.B2(n_52),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_4),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_4),
.A2(n_27),
.B1(n_30),
.B2(n_52),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g158 ( 
.A1(n_4),
.A2(n_33),
.B1(n_34),
.B2(n_52),
.Y(n_158)
);

BUFx16f_ASAP7_75t_L g75 ( 
.A(n_5),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_6),
.A2(n_75),
.B1(n_80),
.B2(n_130),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_6),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_L g146 ( 
.A1(n_6),
.A2(n_46),
.B1(n_47),
.B2(n_130),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_SL g193 ( 
.A1(n_6),
.A2(n_33),
.B1(n_34),
.B2(n_130),
.Y(n_193)
);

AOI22xp33_ASAP7_75t_SL g224 ( 
.A1(n_6),
.A2(n_27),
.B1(n_30),
.B2(n_130),
.Y(n_224)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_7),
.Y(n_63)
);

INVx8_ASAP7_75t_L g122 ( 
.A(n_7),
.Y(n_122)
);

BUFx8_ASAP7_75t_L g34 ( 
.A(n_8),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_9),
.A2(n_75),
.B1(n_80),
.B2(n_152),
.Y(n_151)
);

CKINVDCx14_ASAP7_75t_R g152 ( 
.A(n_9),
.Y(n_152)
);

AOI22xp33_ASAP7_75t_SL g181 ( 
.A1(n_9),
.A2(n_46),
.B1(n_47),
.B2(n_152),
.Y(n_181)
);

AOI22xp33_ASAP7_75t_SL g204 ( 
.A1(n_9),
.A2(n_27),
.B1(n_30),
.B2(n_152),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_9),
.A2(n_33),
.B1(n_34),
.B2(n_152),
.Y(n_209)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_10),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_11),
.A2(n_46),
.B1(n_47),
.B2(n_54),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_11),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_11),
.A2(n_27),
.B1(n_30),
.B2(n_54),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_11),
.A2(n_33),
.B1(n_34),
.B2(n_54),
.Y(n_119)
);

INVx13_ASAP7_75t_L g45 ( 
.A(n_12),
.Y(n_45)
);

INVx13_ASAP7_75t_L g74 ( 
.A(n_13),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_13),
.A2(n_46),
.B1(n_47),
.B2(n_74),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_SL g32 ( 
.A1(n_14),
.A2(n_33),
.B1(n_34),
.B2(n_35),
.Y(n_32)
);

INVx11_ASAP7_75t_L g35 ( 
.A(n_14),
.Y(n_35)
);

A2O1A1Ixp33_ASAP7_75t_L g40 ( 
.A1(n_14),
.A2(n_30),
.B(n_32),
.C(n_41),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_14),
.B(n_30),
.Y(n_41)
);

INVx11_ASAP7_75t_SL g28 ( 
.A(n_15),
.Y(n_28)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_133),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_132),
.Y(n_17)
);

INVxp67_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_SL g19 ( 
.A(n_20),
.B(n_106),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_20),
.B(n_106),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_SL g20 ( 
.A1(n_21),
.A2(n_22),
.B1(n_85),
.B2(n_105),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

XOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_56),
.Y(n_22)
);

AOI21xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_42),
.B(n_55),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_24),
.B(n_42),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_36),
.Y(n_24)
);

OAI21xp5_ASAP7_75t_SL g255 ( 
.A1(n_25),
.A2(n_40),
.B(n_240),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_SL g25 ( 
.A(n_26),
.B(n_31),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_26),
.Y(n_143)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_27),
.Y(n_30)
);

AOI22xp5_ASAP7_75t_L g49 ( 
.A1(n_27),
.A2(n_30),
.B1(n_44),
.B2(n_50),
.Y(n_49)
);

A2O1A1Ixp33_ASAP7_75t_L g199 ( 
.A1(n_27),
.A2(n_35),
.B(n_150),
.C(n_200),
.Y(n_199)
);

NAND2xp33_ASAP7_75t_SL g234 ( 
.A(n_27),
.B(n_44),
.Y(n_234)
);

INVx11_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

AOI32xp33_ASAP7_75t_L g232 ( 
.A1(n_30),
.A2(n_47),
.A3(n_50),
.B1(n_233),
.B2(n_234),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_31),
.B(n_37),
.Y(n_68)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_32),
.A2(n_40),
.B1(n_67),
.B2(n_93),
.Y(n_92)
);

OAI21xp5_ASAP7_75t_L g116 ( 
.A1(n_32),
.A2(n_36),
.B(n_93),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_32),
.A2(n_40),
.B1(n_203),
.B2(n_204),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_32),
.B(n_150),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_32),
.A2(n_40),
.B1(n_204),
.B2(n_224),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_32),
.A2(n_40),
.B1(n_224),
.B2(n_240),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_33),
.B(n_62),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_33),
.B(n_213),
.Y(n_212)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_37),
.B(n_39),
.Y(n_36)
);

INVxp67_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

OAI21xp5_ASAP7_75t_SL g66 ( 
.A1(n_40),
.A2(n_67),
.B(n_68),
.Y(n_66)
);

OAI21xp5_ASAP7_75t_SL g142 ( 
.A1(n_40),
.A2(n_68),
.B(n_143),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g42 ( 
.A1(n_43),
.A2(n_49),
.B1(n_51),
.B2(n_53),
.Y(n_42)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_43),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_43),
.A2(n_49),
.B1(n_146),
.B2(n_147),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_43),
.A2(n_49),
.B1(n_181),
.B2(n_237),
.Y(n_236)
);

A2O1A1Ixp33_ASAP7_75t_L g43 ( 
.A1(n_44),
.A2(n_46),
.B(n_48),
.C(n_49),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_44),
.B(n_46),
.Y(n_48)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_44),
.Y(n_50)
);

INVx11_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_46),
.B(n_74),
.Y(n_156)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_47),
.A2(n_76),
.B1(n_149),
.B2(n_156),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_L g100 ( 
.A1(n_49),
.A2(n_51),
.B(n_101),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_49),
.B(n_104),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_49),
.B(n_125),
.Y(n_167)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_49),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g56 ( 
.A1(n_57),
.A2(n_58),
.B1(n_69),
.B2(n_70),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_58),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_59),
.B(n_66),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_59),
.A2(n_71),
.B1(n_83),
.B2(n_84),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_59),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_59),
.A2(n_66),
.B1(n_84),
.B2(n_111),
.Y(n_110)
);

AOI21xp5_ASAP7_75t_L g59 ( 
.A1(n_60),
.A2(n_63),
.B(n_64),
.Y(n_59)
);

OAI21xp5_ASAP7_75t_L g118 ( 
.A1(n_60),
.A2(n_119),
.B(n_120),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_60),
.A2(n_119),
.B1(n_158),
.B2(n_159),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_60),
.A2(n_63),
.B1(n_193),
.B2(n_209),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_L g225 ( 
.A1(n_60),
.A2(n_91),
.B(n_196),
.Y(n_225)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_61),
.B(n_89),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_61),
.A2(n_192),
.B1(n_194),
.B2(n_195),
.Y(n_191)
);

AOI21xp5_ASAP7_75t_L g231 ( 
.A1(n_61),
.A2(n_65),
.B(n_121),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_62),
.B(n_65),
.Y(n_91)
);

INVx4_ASAP7_75t_L g159 ( 
.A(n_62),
.Y(n_159)
);

INVx5_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_65),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_66),
.Y(n_111)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

CKINVDCx16_ASAP7_75t_R g83 ( 
.A(n_71),
.Y(n_83)
);

OAI21xp5_ASAP7_75t_SL g71 ( 
.A1(n_72),
.A2(n_78),
.B(n_81),
.Y(n_71)
);

OAI21xp5_ASAP7_75t_SL g95 ( 
.A1(n_72),
.A2(n_96),
.B(n_98),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_72),
.A2(n_96),
.B1(n_129),
.B2(n_131),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_72),
.A2(n_129),
.B1(n_131),
.B2(n_163),
.Y(n_162)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_73),
.A2(n_77),
.B1(n_149),
.B2(n_151),
.Y(n_148)
);

O2A1O1Ixp33_ASAP7_75t_L g73 ( 
.A1(n_74),
.A2(n_75),
.B(n_76),
.C(n_77),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_74),
.B(n_75),
.Y(n_76)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_75),
.Y(n_80)
);

HAxp5_ASAP7_75t_SL g149 ( 
.A(n_75),
.B(n_150),
.CON(n_149),
.SN(n_149)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_77),
.B(n_82),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_77),
.B(n_79),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_77),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_79),
.Y(n_78)
);

CKINVDCx16_ASAP7_75t_R g105 ( 
.A(n_85),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_86),
.B(n_94),
.C(n_99),
.Y(n_85)
);

XOR2xp5_ASAP7_75t_L g108 ( 
.A(n_86),
.B(n_109),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_92),
.Y(n_86)
);

XOR2xp5_ASAP7_75t_L g269 ( 
.A(n_87),
.B(n_92),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_88),
.B(n_91),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_L g177 ( 
.A1(n_88),
.A2(n_122),
.B(n_158),
.Y(n_177)
);

INVxp67_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_90),
.B(n_122),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_94),
.A2(n_95),
.B1(n_99),
.B2(n_100),
.Y(n_109)
);

CKINVDCx14_ASAP7_75t_R g94 ( 
.A(n_95),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_100),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_102),
.B(n_103),
.Y(n_101)
);

AOI21xp5_ASAP7_75t_L g123 ( 
.A1(n_102),
.A2(n_124),
.B(n_126),
.Y(n_123)
);

AOI21xp5_ASAP7_75t_L g165 ( 
.A1(n_102),
.A2(n_166),
.B(n_167),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_102),
.A2(n_180),
.B1(n_182),
.B2(n_183),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_104),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_107),
.B(n_110),
.C(n_112),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_107),
.A2(n_108),
.B1(n_110),
.B2(n_282),
.Y(n_281)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

CKINVDCx14_ASAP7_75t_R g282 ( 
.A(n_110),
.Y(n_282)
);

XOR2xp5_ASAP7_75t_L g280 ( 
.A(n_112),
.B(n_281),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_113),
.B(n_123),
.C(n_127),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_113),
.A2(n_114),
.B1(n_272),
.B2(n_273),
.Y(n_271)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_115),
.B(n_117),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_115),
.A2(n_116),
.B1(n_117),
.B2(n_118),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_116),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_118),
.Y(n_117)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_122),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_122),
.B(n_150),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_123),
.A2(n_127),
.B1(n_128),
.B2(n_274),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_123),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_125),
.Y(n_124)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_SL g133 ( 
.A1(n_134),
.A2(n_278),
.B(n_283),
.Y(n_133)
);

O2A1O1Ixp33_ASAP7_75t_SL g134 ( 
.A1(n_135),
.A2(n_184),
.B(n_263),
.C(n_277),
.Y(n_134)
);

AND2x2_ASAP7_75t_L g135 ( 
.A(n_136),
.B(n_169),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_136),
.B(n_169),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_137),
.A2(n_138),
.B1(n_153),
.B2(n_168),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_SL g138 ( 
.A(n_139),
.B(n_140),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_139),
.B(n_140),
.C(n_168),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_141),
.B(n_144),
.C(n_148),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_141),
.A2(n_142),
.B1(n_144),
.B2(n_145),
.Y(n_171)
);

CKINVDCx16_ASAP7_75t_R g141 ( 
.A(n_142),
.Y(n_141)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_146),
.Y(n_183)
);

CKINVDCx16_ASAP7_75t_R g166 ( 
.A(n_147),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_SL g170 ( 
.A(n_148),
.B(n_171),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_151),
.Y(n_163)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_153),
.Y(n_168)
);

XOR2xp5_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_160),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_154),
.B(n_161),
.C(n_165),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_157),
.Y(n_154)
);

XOR2xp5_ASAP7_75t_L g173 ( 
.A(n_155),
.B(n_157),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_161),
.A2(n_162),
.B1(n_164),
.B2(n_165),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

CKINVDCx16_ASAP7_75t_R g164 ( 
.A(n_165),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_172),
.C(n_174),
.Y(n_169)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_170),
.B(n_260),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_L g260 ( 
.A1(n_172),
.A2(n_173),
.B1(n_174),
.B2(n_175),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_173),
.Y(n_172)
);

CKINVDCx16_ASAP7_75t_R g174 ( 
.A(n_175),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_176),
.B(n_178),
.C(n_179),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_176),
.A2(n_177),
.B1(n_178),
.B2(n_251),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_177),
.Y(n_176)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_178),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_SL g249 ( 
.A(n_179),
.B(n_250),
.Y(n_249)
);

CKINVDCx14_ASAP7_75t_R g180 ( 
.A(n_181),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_SL g184 ( 
.A(n_185),
.B(n_262),
.Y(n_184)
);

AOI21xp5_ASAP7_75t_L g185 ( 
.A1(n_186),
.A2(n_257),
.B(n_261),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_SL g186 ( 
.A1(n_187),
.A2(n_245),
.B(n_256),
.Y(n_186)
);

AOI21xp5_ASAP7_75t_L g187 ( 
.A1(n_188),
.A2(n_227),
.B(n_244),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_SL g188 ( 
.A1(n_189),
.A2(n_216),
.B(n_226),
.Y(n_188)
);

AOI21xp5_ASAP7_75t_L g189 ( 
.A1(n_190),
.A2(n_205),
.B(n_215),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_191),
.B(n_197),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_191),
.B(n_197),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_193),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_196),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_198),
.A2(n_199),
.B1(n_201),
.B2(n_202),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_199),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_SL g217 ( 
.A(n_199),
.B(n_201),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_202),
.Y(n_201)
);

OAI21xp5_ASAP7_75t_SL g205 ( 
.A1(n_206),
.A2(n_210),
.B(n_214),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_207),
.B(n_208),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_207),
.B(n_208),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_211),
.B(n_212),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_217),
.B(n_218),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_217),
.B(n_218),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g218 ( 
.A(n_219),
.B(n_225),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_220),
.A2(n_221),
.B1(n_222),
.B2(n_223),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_220),
.B(n_223),
.C(n_225),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_221),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_223),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_228),
.B(n_229),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_228),
.B(n_229),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_230),
.A2(n_235),
.B1(n_242),
.B2(n_243),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_230),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_231),
.B(n_232),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_231),
.B(n_232),
.Y(n_254)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_235),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_236),
.A2(n_238),
.B1(n_239),
.B2(n_241),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_236),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_238),
.B(n_241),
.C(n_242),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_239),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_246),
.B(n_247),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_SL g256 ( 
.A(n_246),
.B(n_247),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_248),
.A2(n_249),
.B1(n_252),
.B2(n_253),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_248),
.B(n_254),
.C(n_255),
.Y(n_258)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_253),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_254),
.B(n_255),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_258),
.B(n_259),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_SL g261 ( 
.A(n_258),
.B(n_259),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_264),
.B(n_265),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_SL g277 ( 
.A(n_264),
.B(n_265),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_266),
.A2(n_267),
.B1(n_275),
.B2(n_276),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_L g267 ( 
.A1(n_268),
.A2(n_269),
.B1(n_270),
.B2(n_271),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_268),
.B(n_271),
.C(n_276),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_269),
.Y(n_268)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

CKINVDCx14_ASAP7_75t_R g276 ( 
.A(n_275),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_279),
.B(n_280),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_SL g283 ( 
.A(n_279),
.B(n_280),
.Y(n_283)
);


endmodule