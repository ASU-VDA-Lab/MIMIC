module fake_aes_181_n_853 (n_44, n_81, n_69, n_22, n_57, n_88, n_52, n_26, n_50, n_33, n_73, n_49, n_97, n_80, n_60, n_41, n_35, n_94, n_65, n_9, n_10, n_19, n_87, n_98, n_74, n_7, n_29, n_45, n_85, n_101, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_91, n_16, n_13, n_95, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_84, n_55, n_12, n_86, n_75, n_72, n_43, n_76, n_89, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_83, n_28, n_48, n_100, n_92, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_82, n_15, n_61, n_21, n_99, n_93, n_51, n_96, n_39, n_853);
input n_44;
input n_81;
input n_69;
input n_22;
input n_57;
input n_88;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_97;
input n_80;
input n_60;
input n_41;
input n_35;
input n_94;
input n_65;
input n_9;
input n_10;
input n_19;
input n_87;
input n_98;
input n_74;
input n_7;
input n_29;
input n_45;
input n_85;
input n_101;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_16;
input n_13;
input n_95;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_84;
input n_55;
input n_12;
input n_86;
input n_75;
input n_72;
input n_43;
input n_76;
input n_89;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_83;
input n_28;
input n_48;
input n_100;
input n_92;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_82;
input n_15;
input n_61;
input n_21;
input n_99;
input n_93;
input n_51;
input n_96;
input n_39;
output n_853;
wire n_117;
wire n_663;
wire n_707;
wire n_791;
wire n_361;
wire n_513;
wire n_838;
wire n_185;
wire n_705;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_755;
wire n_646;
wire n_792;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_848;
wire n_607;
wire n_808;
wire n_829;
wire n_125;
wire n_431;
wire n_484;
wire n_852;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_801;
wire n_292;
wire n_309;
wire n_160;
wire n_701;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_743;
wire n_523;
wire n_229;
wire n_757;
wire n_750;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_770;
wire n_252;
wire n_152;
wire n_113;
wire n_814;
wire n_637;
wire n_817;
wire n_802;
wire n_353;
wire n_564;
wire n_779;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_850;
wire n_762;
wire n_672;
wire n_532;
wire n_627;
wire n_758;
wire n_544;
wire n_400;
wire n_787;
wire n_296;
wire n_157;
wire n_765;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_807;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_783;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_715;
wire n_463;
wire n_131;
wire n_112;
wire n_789;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_476;
wire n_105;
wire n_227;
wire n_384;
wire n_434;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_812;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_777;
wire n_752;
wire n_732;
wire n_199;
wire n_351;
wire n_401;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_724;
wire n_786;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_796;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_702;
wire n_572;
wire n_324;
wire n_773;
wire n_847;
wire n_840;
wire n_392;
wire n_668;
wire n_846;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_830;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_623;
wire n_167;
wire n_593;
wire n_697;
wire n_554;
wire n_726;
wire n_780;
wire n_712;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_809;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_764;
wire n_314;
wire n_237;
wire n_181;
wire n_255;
wire n_426;
wire n_624;
wire n_725;
wire n_769;
wire n_818;
wire n_844;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_738;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_798;
wire n_241;
wire n_575;
wire n_711;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_767;
wire n_828;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_826;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_708;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_730;
wire n_771;
wire n_696;
wire n_735;
wire n_784;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_243;
wire n_235;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_813;
wire n_352;
wire n_746;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_803;
wire n_299;
wire n_338;
wire n_699;
wire n_519;
wire n_729;
wire n_805;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_849;
wire n_810;
wire n_172;
wire n_329;
wire n_251;
wire n_747;
wire n_635;
wire n_731;
wire n_689;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_719;
wire n_611;
wire n_704;
wire n_633;
wire n_271;
wire n_760;
wire n_751;
wire n_800;
wire n_626;
wire n_302;
wire n_466;
wire n_710;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_412;
wire n_664;
wire n_827;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_788;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_839;
wire n_450;
wire n_579;
wire n_107;
wire n_776;
wire n_403;
wire n_557;
wire n_516;
wire n_842;
wire n_254;
wire n_549;
wire n_622;
wire n_832;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_649;
wire n_526;
wire n_276;
wire n_320;
wire n_768;
wire n_797;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_621;
wire n_666;
wire n_799;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_706;
wire n_822;
wire n_823;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_720;
wire n_568;
wire n_245;
wire n_357;
wire n_716;
wire n_653;
wire n_260;
wire n_806;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_718;
wire n_111;
wire n_536;
wire n_816;
wire n_265;
wire n_264;
wire n_522;
wire n_208;
wire n_200;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_754;
wire n_775;
wire n_616;
wire n_118;
wire n_365;
wire n_717;
wire n_541;
wire n_179;
wire n_363;
wire n_315;
wire n_409;
wire n_733;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_794;
wire n_376;
wire n_639;
wire n_552;
wire n_744;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_756;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_790;
wire n_761;
wire n_615;
wire n_212;
wire n_472;
wire n_419;
wire n_851;
wire n_825;
wire n_396;
wire n_168;
wire n_804;
wire n_477;
wire n_815;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_721;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_821;
wire n_745;
wire n_684;
wire n_440;
wire n_106;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_597;
wire n_498;
wire n_723;
wire n_811;
wire n_749;
wire n_835;
wire n_225;
wire n_535;
wire n_530;
wire n_737;
wire n_778;
wire n_220;
wire n_358;
wire n_795;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_782;
wire n_102;
wire n_449;
wire n_115;
wire n_300;
wire n_158;
wire n_734;
wire n_524;
wire n_121;
wire n_584;
wire n_763;
wire n_497;
wire n_728;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_841;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_836;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_741;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_766;
wire n_602;
wire n_831;
wire n_198;
wire n_169;
wire n_424;
wire n_714;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_837;
wire n_128;
wire n_129;
wire n_410;
wire n_774;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_722;
wire n_618;
wire n_834;
wire n_727;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_785;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_748;
wire n_371;
wire n_688;
wire n_323;
wire n_473;
wire n_347;
wire n_820;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_843;
wire n_266;
wire n_683;
wire n_213;
wire n_824;
wire n_538;
wire n_793;
wire n_182;
wire n_492;
wire n_592;
wire n_753;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_695;
wire n_650;
wire n_469;
wire n_742;
wire n_585;
wire n_845;
wire n_713;
wire n_123;
wire n_457;
wire n_595;
wire n_759;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_453;
wire n_372;
wire n_631;
wire n_833;
wire n_736;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_781;
wire n_421;
wire n_175;
wire n_709;
wire n_739;
wire n_145;
wire n_740;
wire n_483;
wire n_408;
wire n_772;
wire n_290;
wire n_405;
wire n_819;
wire n_280;
wire n_132;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g102 ( .A(n_58), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_28), .Y(n_103) );
CKINVDCx5p33_ASAP7_75t_R g104 ( .A(n_62), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_2), .Y(n_105) );
CKINVDCx5p33_ASAP7_75t_R g106 ( .A(n_10), .Y(n_106) );
CKINVDCx5p33_ASAP7_75t_R g107 ( .A(n_63), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_101), .Y(n_108) );
CKINVDCx5p33_ASAP7_75t_R g109 ( .A(n_75), .Y(n_109) );
CKINVDCx5p33_ASAP7_75t_R g110 ( .A(n_20), .Y(n_110) );
INVx2_ASAP7_75t_SL g111 ( .A(n_39), .Y(n_111) );
INVx2_ASAP7_75t_L g112 ( .A(n_48), .Y(n_112) );
CKINVDCx5p33_ASAP7_75t_R g113 ( .A(n_1), .Y(n_113) );
CKINVDCx16_ASAP7_75t_R g114 ( .A(n_42), .Y(n_114) );
CKINVDCx20_ASAP7_75t_R g115 ( .A(n_7), .Y(n_115) );
HB1xp67_ASAP7_75t_L g116 ( .A(n_56), .Y(n_116) );
CKINVDCx5p33_ASAP7_75t_R g117 ( .A(n_86), .Y(n_117) );
CKINVDCx5p33_ASAP7_75t_R g118 ( .A(n_66), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_37), .Y(n_119) );
CKINVDCx5p33_ASAP7_75t_R g120 ( .A(n_43), .Y(n_120) );
CKINVDCx5p33_ASAP7_75t_R g121 ( .A(n_41), .Y(n_121) );
CKINVDCx5p33_ASAP7_75t_R g122 ( .A(n_69), .Y(n_122) );
INVx2_ASAP7_75t_L g123 ( .A(n_68), .Y(n_123) );
BUFx2_ASAP7_75t_L g124 ( .A(n_49), .Y(n_124) );
INVx1_ASAP7_75t_L g125 ( .A(n_92), .Y(n_125) );
CKINVDCx5p33_ASAP7_75t_R g126 ( .A(n_26), .Y(n_126) );
CKINVDCx5p33_ASAP7_75t_R g127 ( .A(n_78), .Y(n_127) );
INVx1_ASAP7_75t_L g128 ( .A(n_24), .Y(n_128) );
CKINVDCx20_ASAP7_75t_R g129 ( .A(n_93), .Y(n_129) );
INVx1_ASAP7_75t_L g130 ( .A(n_3), .Y(n_130) );
CKINVDCx20_ASAP7_75t_R g131 ( .A(n_30), .Y(n_131) );
INVx2_ASAP7_75t_L g132 ( .A(n_5), .Y(n_132) );
CKINVDCx5p33_ASAP7_75t_R g133 ( .A(n_80), .Y(n_133) );
INVx1_ASAP7_75t_L g134 ( .A(n_83), .Y(n_134) );
CKINVDCx5p33_ASAP7_75t_R g135 ( .A(n_45), .Y(n_135) );
CKINVDCx5p33_ASAP7_75t_R g136 ( .A(n_8), .Y(n_136) );
INVxp33_ASAP7_75t_L g137 ( .A(n_84), .Y(n_137) );
INVx1_ASAP7_75t_L g138 ( .A(n_60), .Y(n_138) );
NOR2xp67_ASAP7_75t_L g139 ( .A(n_90), .B(n_7), .Y(n_139) );
INVx2_ASAP7_75t_L g140 ( .A(n_112), .Y(n_140) );
NAND2xp5_ASAP7_75t_L g141 ( .A(n_124), .B(n_0), .Y(n_141) );
AND2x4_ASAP7_75t_L g142 ( .A(n_132), .B(n_0), .Y(n_142) );
INVx1_ASAP7_75t_L g143 ( .A(n_132), .Y(n_143) );
AND2x2_ASAP7_75t_L g144 ( .A(n_137), .B(n_1), .Y(n_144) );
INVx5_ASAP7_75t_L g145 ( .A(n_111), .Y(n_145) );
AND2x4_ASAP7_75t_L g146 ( .A(n_111), .B(n_2), .Y(n_146) );
INVx1_ASAP7_75t_L g147 ( .A(n_102), .Y(n_147) );
INVx3_ASAP7_75t_L g148 ( .A(n_112), .Y(n_148) );
OAI22xp5_ASAP7_75t_L g149 ( .A1(n_106), .A2(n_3), .B1(n_4), .B2(n_5), .Y(n_149) );
INVx3_ASAP7_75t_L g150 ( .A(n_123), .Y(n_150) );
INVx1_ASAP7_75t_L g151 ( .A(n_103), .Y(n_151) );
BUFx6f_ASAP7_75t_L g152 ( .A(n_123), .Y(n_152) );
BUFx6f_ASAP7_75t_L g153 ( .A(n_108), .Y(n_153) );
INVx1_ASAP7_75t_L g154 ( .A(n_119), .Y(n_154) );
AND2x4_ASAP7_75t_L g155 ( .A(n_116), .B(n_4), .Y(n_155) );
NAND2xp5_ASAP7_75t_L g156 ( .A(n_105), .B(n_6), .Y(n_156) );
BUFx3_ASAP7_75t_L g157 ( .A(n_125), .Y(n_157) );
BUFx6f_ASAP7_75t_L g158 ( .A(n_128), .Y(n_158) );
INVx1_ASAP7_75t_L g159 ( .A(n_134), .Y(n_159) );
NAND2xp5_ASAP7_75t_L g160 ( .A(n_130), .B(n_6), .Y(n_160) );
OAI22x1_ASAP7_75t_L g161 ( .A1(n_106), .A2(n_8), .B1(n_9), .B2(n_10), .Y(n_161) );
NAND2xp5_ASAP7_75t_L g162 ( .A(n_114), .B(n_9), .Y(n_162) );
INVx4_ASAP7_75t_L g163 ( .A(n_104), .Y(n_163) );
INVx2_ASAP7_75t_L g164 ( .A(n_152), .Y(n_164) );
NAND2xp5_ASAP7_75t_L g165 ( .A(n_163), .B(n_136), .Y(n_165) );
NAND2xp5_ASAP7_75t_L g166 ( .A(n_163), .B(n_136), .Y(n_166) );
INVx1_ASAP7_75t_L g167 ( .A(n_152), .Y(n_167) );
NOR2x1p5_ASAP7_75t_L g168 ( .A(n_141), .B(n_104), .Y(n_168) );
NOR2xp33_ASAP7_75t_L g169 ( .A(n_163), .B(n_138), .Y(n_169) );
INVx2_ASAP7_75t_L g170 ( .A(n_152), .Y(n_170) );
NAND2xp5_ASAP7_75t_L g171 ( .A(n_163), .B(n_107), .Y(n_171) );
BUFx4f_ASAP7_75t_L g172 ( .A(n_146), .Y(n_172) );
OR2x6_ASAP7_75t_L g173 ( .A(n_161), .B(n_139), .Y(n_173) );
INVx2_ASAP7_75t_L g174 ( .A(n_152), .Y(n_174) );
INVx1_ASAP7_75t_L g175 ( .A(n_152), .Y(n_175) );
NAND2xp5_ASAP7_75t_L g176 ( .A(n_147), .B(n_107), .Y(n_176) );
INVx2_ASAP7_75t_L g177 ( .A(n_152), .Y(n_177) );
INVx4_ASAP7_75t_L g178 ( .A(n_146), .Y(n_178) );
NAND2xp33_ASAP7_75t_SL g179 ( .A(n_144), .B(n_129), .Y(n_179) );
INVx2_ASAP7_75t_L g180 ( .A(n_152), .Y(n_180) );
AOI21x1_ASAP7_75t_L g181 ( .A1(n_140), .A2(n_135), .B(n_133), .Y(n_181) );
INVx1_ASAP7_75t_L g182 ( .A(n_153), .Y(n_182) );
AOI21x1_ASAP7_75t_L g183 ( .A1(n_140), .A2(n_135), .B(n_133), .Y(n_183) );
BUFx10_ASAP7_75t_L g184 ( .A(n_146), .Y(n_184) );
CKINVDCx6p67_ASAP7_75t_R g185 ( .A(n_162), .Y(n_185) );
INVx1_ASAP7_75t_L g186 ( .A(n_153), .Y(n_186) );
INVx2_ASAP7_75t_L g187 ( .A(n_153), .Y(n_187) );
INVx2_ASAP7_75t_L g188 ( .A(n_153), .Y(n_188) );
INVx2_ASAP7_75t_L g189 ( .A(n_153), .Y(n_189) );
INVx4_ASAP7_75t_L g190 ( .A(n_146), .Y(n_190) );
INVx2_ASAP7_75t_L g191 ( .A(n_153), .Y(n_191) );
OAI21xp33_ASAP7_75t_SL g192 ( .A1(n_147), .A2(n_11), .B(n_12), .Y(n_192) );
INVx1_ASAP7_75t_L g193 ( .A(n_153), .Y(n_193) );
INVx1_ASAP7_75t_L g194 ( .A(n_158), .Y(n_194) );
NAND2xp5_ASAP7_75t_SL g195 ( .A(n_155), .B(n_109), .Y(n_195) );
NAND2xp5_ASAP7_75t_SL g196 ( .A(n_155), .B(n_109), .Y(n_196) );
INVx3_ASAP7_75t_L g197 ( .A(n_142), .Y(n_197) );
INVx1_ASAP7_75t_L g198 ( .A(n_158), .Y(n_198) );
INVx2_ASAP7_75t_L g199 ( .A(n_158), .Y(n_199) );
INVx2_ASAP7_75t_L g200 ( .A(n_158), .Y(n_200) );
BUFx3_ASAP7_75t_L g201 ( .A(n_145), .Y(n_201) );
INVx2_ASAP7_75t_L g202 ( .A(n_158), .Y(n_202) );
INVx1_ASAP7_75t_L g203 ( .A(n_158), .Y(n_203) );
INVx3_ASAP7_75t_L g204 ( .A(n_142), .Y(n_204) );
AOI21x1_ASAP7_75t_L g205 ( .A1(n_140), .A2(n_110), .B(n_127), .Y(n_205) );
INVx1_ASAP7_75t_L g206 ( .A(n_158), .Y(n_206) );
INVx1_ASAP7_75t_L g207 ( .A(n_148), .Y(n_207) );
CKINVDCx5p33_ASAP7_75t_R g208 ( .A(n_144), .Y(n_208) );
INVx2_ASAP7_75t_L g209 ( .A(n_191), .Y(n_209) );
NOR2xp33_ASAP7_75t_L g210 ( .A(n_165), .B(n_151), .Y(n_210) );
NOR2xp33_ASAP7_75t_L g211 ( .A(n_166), .B(n_151), .Y(n_211) );
OAI22xp5_ASAP7_75t_L g212 ( .A1(n_172), .A2(n_162), .B1(n_131), .B2(n_155), .Y(n_212) );
NAND2xp5_ASAP7_75t_L g213 ( .A(n_176), .B(n_155), .Y(n_213) );
AOI22xp33_ASAP7_75t_L g214 ( .A1(n_172), .A2(n_142), .B1(n_157), .B2(n_159), .Y(n_214) );
NOR2xp33_ASAP7_75t_L g215 ( .A(n_171), .B(n_154), .Y(n_215) );
AOI22xp33_ASAP7_75t_L g216 ( .A1(n_172), .A2(n_142), .B1(n_157), .B2(n_159), .Y(n_216) );
NAND2xp5_ASAP7_75t_L g217 ( .A(n_168), .B(n_141), .Y(n_217) );
AND2x2_ASAP7_75t_L g218 ( .A(n_168), .B(n_154), .Y(n_218) );
OAI221xp5_ASAP7_75t_L g219 ( .A1(n_192), .A2(n_160), .B1(n_156), .B2(n_149), .C(n_157), .Y(n_219) );
O2A1O1Ixp33_ASAP7_75t_L g220 ( .A1(n_192), .A2(n_160), .B(n_156), .C(n_149), .Y(n_220) );
NAND2xp5_ASAP7_75t_L g221 ( .A(n_178), .B(n_110), .Y(n_221) );
AND2x6_ASAP7_75t_SL g222 ( .A(n_173), .B(n_143), .Y(n_222) );
NOR2xp67_ASAP7_75t_L g223 ( .A(n_178), .B(n_145), .Y(n_223) );
AND2x6_ASAP7_75t_SL g224 ( .A(n_173), .B(n_143), .Y(n_224) );
A2O1A1Ixp33_ASAP7_75t_L g225 ( .A1(n_172), .A2(n_150), .B(n_148), .C(n_145), .Y(n_225) );
O2A1O1Ixp5_ASAP7_75t_L g226 ( .A1(n_195), .A2(n_150), .B(n_148), .C(n_145), .Y(n_226) );
INVx1_ASAP7_75t_L g227 ( .A(n_197), .Y(n_227) );
NAND2xp5_ASAP7_75t_L g228 ( .A(n_178), .B(n_121), .Y(n_228) );
NAND2xp5_ASAP7_75t_L g229 ( .A(n_178), .B(n_121), .Y(n_229) );
INVx2_ASAP7_75t_L g230 ( .A(n_191), .Y(n_230) );
NAND2xp5_ASAP7_75t_L g231 ( .A(n_190), .B(n_127), .Y(n_231) );
AOI22xp33_ASAP7_75t_L g232 ( .A1(n_190), .A2(n_161), .B1(n_150), .B2(n_148), .Y(n_232) );
A2O1A1Ixp33_ASAP7_75t_L g233 ( .A1(n_197), .A2(n_150), .B(n_145), .C(n_113), .Y(n_233) );
NOR2xp33_ASAP7_75t_L g234 ( .A(n_196), .B(n_145), .Y(n_234) );
INVx2_ASAP7_75t_L g235 ( .A(n_199), .Y(n_235) );
BUFx3_ASAP7_75t_L g236 ( .A(n_184), .Y(n_236) );
INVx1_ASAP7_75t_L g237 ( .A(n_197), .Y(n_237) );
NOR3xp33_ASAP7_75t_L g238 ( .A(n_179), .B(n_126), .C(n_122), .Y(n_238) );
NOR2xp33_ASAP7_75t_L g239 ( .A(n_208), .B(n_145), .Y(n_239) );
INVx8_ASAP7_75t_L g240 ( .A(n_197), .Y(n_240) );
INVx2_ASAP7_75t_L g241 ( .A(n_199), .Y(n_241) );
INVx2_ASAP7_75t_SL g242 ( .A(n_184), .Y(n_242) );
AOI22xp5_ASAP7_75t_L g243 ( .A1(n_173), .A2(n_161), .B1(n_115), .B2(n_118), .Y(n_243) );
NAND2xp5_ASAP7_75t_SL g244 ( .A(n_184), .B(n_120), .Y(n_244) );
INVx2_ASAP7_75t_L g245 ( .A(n_200), .Y(n_245) );
NAND2xp5_ASAP7_75t_SL g246 ( .A(n_184), .B(n_117), .Y(n_246) );
INVx1_ASAP7_75t_L g247 ( .A(n_204), .Y(n_247) );
NOR2xp33_ASAP7_75t_L g248 ( .A(n_185), .B(n_54), .Y(n_248) );
INVx1_ASAP7_75t_L g249 ( .A(n_204), .Y(n_249) );
AOI22xp33_ASAP7_75t_L g250 ( .A1(n_190), .A2(n_11), .B1(n_12), .B2(n_13), .Y(n_250) );
NAND3xp33_ASAP7_75t_L g251 ( .A(n_169), .B(n_190), .C(n_204), .Y(n_251) );
INVx2_ASAP7_75t_SL g252 ( .A(n_204), .Y(n_252) );
O2A1O1Ixp5_ASAP7_75t_L g253 ( .A1(n_181), .A2(n_100), .B(n_55), .C(n_57), .Y(n_253) );
INVx1_ASAP7_75t_L g254 ( .A(n_207), .Y(n_254) );
NOR2xp33_ASAP7_75t_SL g255 ( .A(n_185), .B(n_13), .Y(n_255) );
INVx1_ASAP7_75t_L g256 ( .A(n_207), .Y(n_256) );
INVx2_ASAP7_75t_L g257 ( .A(n_200), .Y(n_257) );
NOR2xp33_ASAP7_75t_L g258 ( .A(n_181), .B(n_53), .Y(n_258) );
INVx3_ASAP7_75t_L g259 ( .A(n_183), .Y(n_259) );
AOI21xp5_ASAP7_75t_L g260 ( .A1(n_213), .A2(n_201), .B(n_186), .Y(n_260) );
NAND2xp5_ASAP7_75t_L g261 ( .A(n_210), .B(n_183), .Y(n_261) );
O2A1O1Ixp33_ASAP7_75t_L g262 ( .A1(n_219), .A2(n_173), .B(n_206), .C(n_203), .Y(n_262) );
BUFx2_ASAP7_75t_L g263 ( .A(n_240), .Y(n_263) );
NAND2xp5_ASAP7_75t_SL g264 ( .A(n_236), .B(n_205), .Y(n_264) );
O2A1O1Ixp5_ASAP7_75t_L g265 ( .A1(n_258), .A2(n_205), .B(n_182), .C(n_203), .Y(n_265) );
AOI22x1_ASAP7_75t_L g266 ( .A1(n_259), .A2(n_164), .B1(n_187), .B2(n_188), .Y(n_266) );
AOI21xp5_ASAP7_75t_L g267 ( .A1(n_259), .A2(n_201), .B(n_182), .Y(n_267) );
NOR2xp33_ASAP7_75t_L g268 ( .A(n_217), .B(n_173), .Y(n_268) );
AOI21xp5_ASAP7_75t_L g269 ( .A1(n_259), .A2(n_201), .B(n_186), .Y(n_269) );
O2A1O1Ixp33_ASAP7_75t_L g270 ( .A1(n_220), .A2(n_206), .B(n_198), .C(n_194), .Y(n_270) );
NAND2xp5_ASAP7_75t_L g271 ( .A(n_218), .B(n_14), .Y(n_271) );
NAND2xp5_ASAP7_75t_L g272 ( .A(n_211), .B(n_193), .Y(n_272) );
O2A1O1Ixp33_ASAP7_75t_L g273 ( .A1(n_212), .A2(n_198), .B(n_194), .C(n_193), .Y(n_273) );
AOI21x1_ASAP7_75t_L g274 ( .A1(n_223), .A2(n_167), .B(n_175), .Y(n_274) );
BUFx4f_ASAP7_75t_L g275 ( .A(n_218), .Y(n_275) );
AND2x2_ASAP7_75t_L g276 ( .A(n_243), .B(n_14), .Y(n_276) );
NOR2x1_ASAP7_75t_L g277 ( .A(n_248), .B(n_202), .Y(n_277) );
AND2x2_ASAP7_75t_L g278 ( .A(n_243), .B(n_15), .Y(n_278) );
NAND2xp5_ASAP7_75t_SL g279 ( .A(n_236), .B(n_189), .Y(n_279) );
AND2x2_ASAP7_75t_L g280 ( .A(n_215), .B(n_15), .Y(n_280) );
AOI21xp5_ASAP7_75t_L g281 ( .A1(n_227), .A2(n_167), .B(n_175), .Y(n_281) );
INVx5_ASAP7_75t_L g282 ( .A(n_240), .Y(n_282) );
AND2x2_ASAP7_75t_SL g283 ( .A(n_255), .B(n_16), .Y(n_283) );
NAND2xp5_ASAP7_75t_L g284 ( .A(n_227), .B(n_202), .Y(n_284) );
INVx1_ASAP7_75t_L g285 ( .A(n_237), .Y(n_285) );
OAI22xp5_ASAP7_75t_L g286 ( .A1(n_232), .A2(n_189), .B1(n_188), .B2(n_187), .Y(n_286) );
NAND3xp33_ASAP7_75t_L g287 ( .A(n_238), .B(n_189), .C(n_188), .Y(n_287) );
AOI21xp5_ASAP7_75t_L g288 ( .A1(n_237), .A2(n_187), .B(n_164), .Y(n_288) );
O2A1O1Ixp33_ASAP7_75t_L g289 ( .A1(n_233), .A2(n_180), .B(n_177), .C(n_174), .Y(n_289) );
BUFx6f_ASAP7_75t_L g290 ( .A(n_240), .Y(n_290) );
NAND2xp5_ASAP7_75t_SL g291 ( .A(n_242), .B(n_164), .Y(n_291) );
NOR2xp33_ASAP7_75t_L g292 ( .A(n_240), .B(n_16), .Y(n_292) );
NAND2xp5_ASAP7_75t_SL g293 ( .A(n_242), .B(n_180), .Y(n_293) );
NAND2xp5_ASAP7_75t_SL g294 ( .A(n_221), .B(n_177), .Y(n_294) );
HB1xp67_ASAP7_75t_L g295 ( .A(n_228), .Y(n_295) );
BUFx6f_ASAP7_75t_L g296 ( .A(n_252), .Y(n_296) );
BUFx8_ASAP7_75t_SL g297 ( .A(n_229), .Y(n_297) );
NAND2x1p5_ASAP7_75t_L g298 ( .A(n_252), .B(n_174), .Y(n_298) );
NOR2x1_ASAP7_75t_L g299 ( .A(n_244), .B(n_170), .Y(n_299) );
NAND2xp5_ASAP7_75t_SL g300 ( .A(n_282), .B(n_231), .Y(n_300) );
NAND2xp33_ASAP7_75t_SL g301 ( .A(n_290), .B(n_214), .Y(n_301) );
AOI221x1_ASAP7_75t_L g302 ( .A1(n_261), .A2(n_225), .B1(n_239), .B2(n_170), .C(n_251), .Y(n_302) );
NAND2xp5_ASAP7_75t_L g303 ( .A(n_268), .B(n_295), .Y(n_303) );
OAI21x1_ASAP7_75t_L g304 ( .A1(n_265), .A2(n_253), .B(n_226), .Y(n_304) );
INVx3_ASAP7_75t_L g305 ( .A(n_282), .Y(n_305) );
NAND3xp33_ASAP7_75t_L g306 ( .A(n_262), .B(n_250), .C(n_216), .Y(n_306) );
OAI21xp5_ASAP7_75t_L g307 ( .A1(n_261), .A2(n_249), .B(n_247), .Y(n_307) );
AO21x2_ASAP7_75t_L g308 ( .A1(n_264), .A2(n_256), .B(n_254), .Y(n_308) );
AO31x2_ASAP7_75t_L g309 ( .A1(n_286), .A2(n_256), .A3(n_254), .B(n_249), .Y(n_309) );
AO31x2_ASAP7_75t_L g310 ( .A1(n_286), .A2(n_247), .A3(n_234), .B(n_245), .Y(n_310) );
AOI221x1_ASAP7_75t_L g311 ( .A1(n_271), .A2(n_257), .B1(n_245), .B2(n_241), .C(n_235), .Y(n_311) );
OAI21x1_ASAP7_75t_L g312 ( .A1(n_266), .A2(n_223), .B(n_241), .Y(n_312) );
INVx2_ASAP7_75t_L g313 ( .A(n_285), .Y(n_313) );
AOI21xp5_ASAP7_75t_L g314 ( .A1(n_267), .A2(n_246), .B(n_257), .Y(n_314) );
NAND2x1p5_ASAP7_75t_L g315 ( .A(n_282), .B(n_235), .Y(n_315) );
AOI22xp33_ASAP7_75t_L g316 ( .A1(n_275), .A2(n_230), .B1(n_209), .B2(n_222), .Y(n_316) );
INVx1_ASAP7_75t_L g317 ( .A(n_270), .Y(n_317) );
NAND2xp5_ASAP7_75t_L g318 ( .A(n_282), .B(n_224), .Y(n_318) );
AND2x2_ASAP7_75t_L g319 ( .A(n_275), .B(n_230), .Y(n_319) );
AOI21xp5_ASAP7_75t_L g320 ( .A1(n_269), .A2(n_209), .B(n_64), .Y(n_320) );
AND2x2_ASAP7_75t_L g321 ( .A(n_280), .B(n_17), .Y(n_321) );
AO31x2_ASAP7_75t_L g322 ( .A1(n_272), .A2(n_17), .A3(n_18), .B(n_19), .Y(n_322) );
BUFx8_ASAP7_75t_L g323 ( .A(n_290), .Y(n_323) );
OAI21xp33_ASAP7_75t_L g324 ( .A1(n_272), .A2(n_18), .B(n_21), .Y(n_324) );
INVx1_ASAP7_75t_L g325 ( .A(n_284), .Y(n_325) );
AOI221x1_ASAP7_75t_L g326 ( .A1(n_260), .A2(n_22), .B1(n_23), .B2(n_25), .C(n_27), .Y(n_326) );
OAI21xp5_ASAP7_75t_L g327 ( .A1(n_317), .A2(n_273), .B(n_289), .Y(n_327) );
INVx1_ASAP7_75t_L g328 ( .A(n_325), .Y(n_328) );
OR2x2_ASAP7_75t_L g329 ( .A(n_325), .B(n_276), .Y(n_329) );
OAI21x1_ASAP7_75t_SL g330 ( .A1(n_307), .A2(n_277), .B(n_274), .Y(n_330) );
INVx1_ASAP7_75t_L g331 ( .A(n_313), .Y(n_331) );
AND2x4_ASAP7_75t_L g332 ( .A(n_305), .B(n_290), .Y(n_332) );
INVx1_ASAP7_75t_L g333 ( .A(n_313), .Y(n_333) );
OA21x2_ASAP7_75t_L g334 ( .A1(n_311), .A2(n_294), .B(n_288), .Y(n_334) );
INVx3_ASAP7_75t_L g335 ( .A(n_323), .Y(n_335) );
OAI21x1_ASAP7_75t_L g336 ( .A1(n_304), .A2(n_299), .B(n_281), .Y(n_336) );
INVx2_ASAP7_75t_L g337 ( .A(n_308), .Y(n_337) );
CKINVDCx5p33_ASAP7_75t_R g338 ( .A(n_323), .Y(n_338) );
OA21x2_ASAP7_75t_L g339 ( .A1(n_311), .A2(n_284), .B(n_287), .Y(n_339) );
INVx1_ASAP7_75t_L g340 ( .A(n_317), .Y(n_340) );
CKINVDCx11_ASAP7_75t_R g341 ( .A(n_323), .Y(n_341) );
OA21x2_ASAP7_75t_L g342 ( .A1(n_326), .A2(n_293), .B(n_291), .Y(n_342) );
INVx2_ASAP7_75t_L g343 ( .A(n_308), .Y(n_343) );
INVx1_ASAP7_75t_L g344 ( .A(n_309), .Y(n_344) );
AO31x2_ASAP7_75t_L g345 ( .A1(n_302), .A2(n_292), .A3(n_263), .B(n_283), .Y(n_345) );
AO31x2_ASAP7_75t_L g346 ( .A1(n_302), .A2(n_278), .A3(n_298), .B(n_296), .Y(n_346) );
OA21x2_ASAP7_75t_L g347 ( .A1(n_326), .A2(n_279), .B(n_298), .Y(n_347) );
OAI21x1_ASAP7_75t_L g348 ( .A1(n_304), .A2(n_296), .B(n_297), .Y(n_348) );
INVx1_ASAP7_75t_L g349 ( .A(n_309), .Y(n_349) );
INVx1_ASAP7_75t_L g350 ( .A(n_309), .Y(n_350) );
NAND3xp33_ASAP7_75t_L g351 ( .A(n_324), .B(n_296), .C(n_31), .Y(n_351) );
INVx1_ASAP7_75t_L g352 ( .A(n_309), .Y(n_352) );
OAI21x1_ASAP7_75t_SL g353 ( .A1(n_318), .A2(n_29), .B(n_32), .Y(n_353) );
INVxp67_ASAP7_75t_SL g354 ( .A(n_323), .Y(n_354) );
INVx1_ASAP7_75t_L g355 ( .A(n_331), .Y(n_355) );
AND2x2_ASAP7_75t_L g356 ( .A(n_331), .B(n_309), .Y(n_356) );
OAI21x1_ASAP7_75t_L g357 ( .A1(n_348), .A2(n_312), .B(n_320), .Y(n_357) );
AO21x2_ASAP7_75t_L g358 ( .A1(n_351), .A2(n_324), .B(n_308), .Y(n_358) );
BUFx4f_ASAP7_75t_L g359 ( .A(n_335), .Y(n_359) );
AND2x4_ASAP7_75t_L g360 ( .A(n_340), .B(n_310), .Y(n_360) );
AO21x1_ASAP7_75t_SL g361 ( .A1(n_344), .A2(n_310), .B(n_316), .Y(n_361) );
INVx1_ASAP7_75t_L g362 ( .A(n_333), .Y(n_362) );
OR2x2_ASAP7_75t_L g363 ( .A(n_333), .B(n_303), .Y(n_363) );
INVx1_ASAP7_75t_L g364 ( .A(n_328), .Y(n_364) );
INVx2_ASAP7_75t_L g365 ( .A(n_337), .Y(n_365) );
INVx3_ASAP7_75t_L g366 ( .A(n_335), .Y(n_366) );
INVx2_ASAP7_75t_L g367 ( .A(n_337), .Y(n_367) );
INVx1_ASAP7_75t_L g368 ( .A(n_328), .Y(n_368) );
INVx2_ASAP7_75t_L g369 ( .A(n_337), .Y(n_369) );
INVx1_ASAP7_75t_L g370 ( .A(n_340), .Y(n_370) );
INVx2_ASAP7_75t_L g371 ( .A(n_343), .Y(n_371) );
INVx2_ASAP7_75t_L g372 ( .A(n_343), .Y(n_372) );
OR2x2_ASAP7_75t_L g373 ( .A(n_329), .B(n_310), .Y(n_373) );
INVx2_ASAP7_75t_L g374 ( .A(n_343), .Y(n_374) );
INVx2_ASAP7_75t_L g375 ( .A(n_344), .Y(n_375) );
OAI21x1_ASAP7_75t_L g376 ( .A1(n_348), .A2(n_312), .B(n_314), .Y(n_376) );
INVx2_ASAP7_75t_L g377 ( .A(n_349), .Y(n_377) );
AND2x2_ASAP7_75t_L g378 ( .A(n_349), .B(n_322), .Y(n_378) );
INVx1_ASAP7_75t_L g379 ( .A(n_350), .Y(n_379) );
INVx1_ASAP7_75t_L g380 ( .A(n_350), .Y(n_380) );
AND2x2_ASAP7_75t_L g381 ( .A(n_352), .B(n_322), .Y(n_381) );
INVx1_ASAP7_75t_L g382 ( .A(n_352), .Y(n_382) );
HB1xp67_ASAP7_75t_L g383 ( .A(n_346), .Y(n_383) );
CKINVDCx5p33_ASAP7_75t_R g384 ( .A(n_341), .Y(n_384) );
OR2x2_ASAP7_75t_L g385 ( .A(n_329), .B(n_310), .Y(n_385) );
AOI22xp33_ASAP7_75t_L g386 ( .A1(n_335), .A2(n_321), .B1(n_306), .B2(n_301), .Y(n_386) );
INVx1_ASAP7_75t_L g387 ( .A(n_327), .Y(n_387) );
OAI21x1_ASAP7_75t_L g388 ( .A1(n_348), .A2(n_300), .B(n_321), .Y(n_388) );
AO21x2_ASAP7_75t_L g389 ( .A1(n_351), .A2(n_306), .B(n_310), .Y(n_389) );
INVx1_ASAP7_75t_L g390 ( .A(n_327), .Y(n_390) );
HB1xp67_ASAP7_75t_L g391 ( .A(n_346), .Y(n_391) );
BUFx3_ASAP7_75t_L g392 ( .A(n_335), .Y(n_392) );
INVx4_ASAP7_75t_L g393 ( .A(n_332), .Y(n_393) );
AND2x4_ASAP7_75t_L g394 ( .A(n_332), .B(n_305), .Y(n_394) );
AND2x2_ASAP7_75t_L g395 ( .A(n_346), .B(n_322), .Y(n_395) );
HB1xp67_ASAP7_75t_L g396 ( .A(n_346), .Y(n_396) );
INVx2_ASAP7_75t_L g397 ( .A(n_339), .Y(n_397) );
INVx1_ASAP7_75t_L g398 ( .A(n_346), .Y(n_398) );
INVx2_ASAP7_75t_L g399 ( .A(n_339), .Y(n_399) );
INVx2_ASAP7_75t_L g400 ( .A(n_339), .Y(n_400) );
BUFx2_ASAP7_75t_L g401 ( .A(n_392), .Y(n_401) );
INVx2_ASAP7_75t_L g402 ( .A(n_365), .Y(n_402) );
INVx1_ASAP7_75t_L g403 ( .A(n_364), .Y(n_403) );
AND2x4_ASAP7_75t_L g404 ( .A(n_379), .B(n_380), .Y(n_404) );
AND2x2_ASAP7_75t_L g405 ( .A(n_356), .B(n_346), .Y(n_405) );
INVx2_ASAP7_75t_L g406 ( .A(n_365), .Y(n_406) );
INVx1_ASAP7_75t_L g407 ( .A(n_364), .Y(n_407) );
INVx2_ASAP7_75t_L g408 ( .A(n_365), .Y(n_408) );
INVx1_ASAP7_75t_L g409 ( .A(n_368), .Y(n_409) );
INVx1_ASAP7_75t_L g410 ( .A(n_368), .Y(n_410) );
NAND2xp5_ASAP7_75t_L g411 ( .A(n_363), .B(n_354), .Y(n_411) );
NAND2xp5_ASAP7_75t_L g412 ( .A(n_363), .B(n_322), .Y(n_412) );
INVx1_ASAP7_75t_L g413 ( .A(n_355), .Y(n_413) );
AND2x2_ASAP7_75t_L g414 ( .A(n_356), .B(n_322), .Y(n_414) );
AND2x4_ASAP7_75t_L g415 ( .A(n_379), .B(n_345), .Y(n_415) );
BUFx3_ASAP7_75t_L g416 ( .A(n_359), .Y(n_416) );
AND2x2_ASAP7_75t_L g417 ( .A(n_356), .B(n_345), .Y(n_417) );
INVx2_ASAP7_75t_L g418 ( .A(n_367), .Y(n_418) );
INVx2_ASAP7_75t_L g419 ( .A(n_367), .Y(n_419) );
AND2x2_ASAP7_75t_L g420 ( .A(n_378), .B(n_345), .Y(n_420) );
INVxp67_ASAP7_75t_L g421 ( .A(n_363), .Y(n_421) );
INVx1_ASAP7_75t_L g422 ( .A(n_355), .Y(n_422) );
OR2x2_ASAP7_75t_L g423 ( .A(n_373), .B(n_345), .Y(n_423) );
INVx1_ASAP7_75t_L g424 ( .A(n_362), .Y(n_424) );
INVx2_ASAP7_75t_L g425 ( .A(n_367), .Y(n_425) );
OR2x2_ASAP7_75t_L g426 ( .A(n_373), .B(n_345), .Y(n_426) );
BUFx2_ASAP7_75t_L g427 ( .A(n_392), .Y(n_427) );
INVx2_ASAP7_75t_L g428 ( .A(n_369), .Y(n_428) );
INVx1_ASAP7_75t_L g429 ( .A(n_362), .Y(n_429) );
INVx1_ASAP7_75t_L g430 ( .A(n_370), .Y(n_430) );
INVx1_ASAP7_75t_L g431 ( .A(n_370), .Y(n_431) );
INVx4_ASAP7_75t_L g432 ( .A(n_359), .Y(n_432) );
INVx2_ASAP7_75t_L g433 ( .A(n_369), .Y(n_433) );
OR2x2_ASAP7_75t_L g434 ( .A(n_373), .B(n_345), .Y(n_434) );
OR2x2_ASAP7_75t_L g435 ( .A(n_385), .B(n_338), .Y(n_435) );
HB1xp67_ASAP7_75t_L g436 ( .A(n_392), .Y(n_436) );
INVx1_ASAP7_75t_L g437 ( .A(n_380), .Y(n_437) );
NOR4xp25_ASAP7_75t_SL g438 ( .A(n_384), .B(n_353), .C(n_347), .D(n_342), .Y(n_438) );
INVx1_ASAP7_75t_L g439 ( .A(n_382), .Y(n_439) );
AOI22xp5_ASAP7_75t_SL g440 ( .A1(n_384), .A2(n_332), .B1(n_305), .B2(n_347), .Y(n_440) );
INVx1_ASAP7_75t_L g441 ( .A(n_382), .Y(n_441) );
BUFx3_ASAP7_75t_L g442 ( .A(n_359), .Y(n_442) );
BUFx2_ASAP7_75t_L g443 ( .A(n_392), .Y(n_443) );
INVx1_ASAP7_75t_L g444 ( .A(n_375), .Y(n_444) );
BUFx3_ASAP7_75t_L g445 ( .A(n_359), .Y(n_445) );
AND2x2_ASAP7_75t_L g446 ( .A(n_378), .B(n_339), .Y(n_446) );
INVx3_ASAP7_75t_L g447 ( .A(n_366), .Y(n_447) );
INVx2_ASAP7_75t_L g448 ( .A(n_369), .Y(n_448) );
INVx1_ASAP7_75t_L g449 ( .A(n_375), .Y(n_449) );
BUFx6f_ASAP7_75t_L g450 ( .A(n_359), .Y(n_450) );
AND2x2_ASAP7_75t_L g451 ( .A(n_378), .B(n_332), .Y(n_451) );
OR2x2_ASAP7_75t_L g452 ( .A(n_385), .B(n_334), .Y(n_452) );
INVx1_ASAP7_75t_L g453 ( .A(n_375), .Y(n_453) );
CKINVDCx5p33_ASAP7_75t_R g454 ( .A(n_366), .Y(n_454) );
INVx1_ASAP7_75t_L g455 ( .A(n_377), .Y(n_455) );
INVx1_ASAP7_75t_L g456 ( .A(n_377), .Y(n_456) );
INVx3_ASAP7_75t_L g457 ( .A(n_366), .Y(n_457) );
AND2x4_ASAP7_75t_L g458 ( .A(n_377), .B(n_336), .Y(n_458) );
INVx1_ASAP7_75t_L g459 ( .A(n_385), .Y(n_459) );
NAND2xp5_ASAP7_75t_L g460 ( .A(n_387), .B(n_319), .Y(n_460) );
AND2x2_ASAP7_75t_L g461 ( .A(n_381), .B(n_347), .Y(n_461) );
OAI221xp5_ASAP7_75t_L g462 ( .A1(n_386), .A2(n_319), .B1(n_315), .B2(n_347), .C(n_342), .Y(n_462) );
AND2x4_ASAP7_75t_L g463 ( .A(n_360), .B(n_336), .Y(n_463) );
INVx2_ASAP7_75t_L g464 ( .A(n_371), .Y(n_464) );
INVx2_ASAP7_75t_L g465 ( .A(n_371), .Y(n_465) );
INVx1_ASAP7_75t_L g466 ( .A(n_381), .Y(n_466) );
OR2x2_ASAP7_75t_L g467 ( .A(n_387), .B(n_390), .Y(n_467) );
NAND2xp5_ASAP7_75t_L g468 ( .A(n_390), .B(n_353), .Y(n_468) );
INVx1_ASAP7_75t_L g469 ( .A(n_381), .Y(n_469) );
CKINVDCx20_ASAP7_75t_R g470 ( .A(n_393), .Y(n_470) );
AND2x2_ASAP7_75t_L g471 ( .A(n_395), .B(n_334), .Y(n_471) );
INVxp67_ASAP7_75t_L g472 ( .A(n_366), .Y(n_472) );
OR2x2_ASAP7_75t_L g473 ( .A(n_360), .B(n_334), .Y(n_473) );
INVx3_ASAP7_75t_L g474 ( .A(n_366), .Y(n_474) );
OR2x6_ASAP7_75t_L g475 ( .A(n_393), .B(n_315), .Y(n_475) );
AND2x2_ASAP7_75t_L g476 ( .A(n_395), .B(n_334), .Y(n_476) );
AND2x2_ASAP7_75t_L g477 ( .A(n_395), .B(n_342), .Y(n_477) );
AND2x2_ASAP7_75t_L g478 ( .A(n_360), .B(n_342), .Y(n_478) );
HB1xp67_ASAP7_75t_L g479 ( .A(n_402), .Y(n_479) );
INVx2_ASAP7_75t_L g480 ( .A(n_402), .Y(n_480) );
INVx3_ASAP7_75t_L g481 ( .A(n_458), .Y(n_481) );
AND2x2_ASAP7_75t_L g482 ( .A(n_451), .B(n_435), .Y(n_482) );
OR2x2_ASAP7_75t_L g483 ( .A(n_435), .B(n_374), .Y(n_483) );
INVx1_ASAP7_75t_L g484 ( .A(n_413), .Y(n_484) );
OR2x2_ASAP7_75t_L g485 ( .A(n_421), .B(n_459), .Y(n_485) );
NAND2xp5_ASAP7_75t_L g486 ( .A(n_466), .B(n_360), .Y(n_486) );
INVx1_ASAP7_75t_L g487 ( .A(n_422), .Y(n_487) );
AND2x2_ASAP7_75t_L g488 ( .A(n_451), .B(n_393), .Y(n_488) );
INVx1_ASAP7_75t_L g489 ( .A(n_424), .Y(n_489) );
BUFx8_ASAP7_75t_SL g490 ( .A(n_470), .Y(n_490) );
OR2x2_ASAP7_75t_L g491 ( .A(n_411), .B(n_374), .Y(n_491) );
INVx2_ASAP7_75t_L g492 ( .A(n_406), .Y(n_492) );
AND2x2_ASAP7_75t_L g493 ( .A(n_469), .B(n_393), .Y(n_493) );
HB1xp67_ASAP7_75t_L g494 ( .A(n_406), .Y(n_494) );
AND2x2_ASAP7_75t_L g495 ( .A(n_405), .B(n_360), .Y(n_495) );
INVx1_ASAP7_75t_L g496 ( .A(n_429), .Y(n_496) );
NAND2xp5_ASAP7_75t_L g497 ( .A(n_403), .B(n_407), .Y(n_497) );
INVx2_ASAP7_75t_L g498 ( .A(n_408), .Y(n_498) );
INVx1_ASAP7_75t_L g499 ( .A(n_409), .Y(n_499) );
INVx1_ASAP7_75t_L g500 ( .A(n_410), .Y(n_500) );
INVx2_ASAP7_75t_L g501 ( .A(n_408), .Y(n_501) );
OR2x2_ASAP7_75t_L g502 ( .A(n_405), .B(n_374), .Y(n_502) );
AND2x2_ASAP7_75t_L g503 ( .A(n_470), .B(n_393), .Y(n_503) );
AND2x2_ASAP7_75t_L g504 ( .A(n_417), .B(n_394), .Y(n_504) );
AND2x2_ASAP7_75t_L g505 ( .A(n_417), .B(n_394), .Y(n_505) );
INVx1_ASAP7_75t_L g506 ( .A(n_430), .Y(n_506) );
OR2x2_ASAP7_75t_L g507 ( .A(n_444), .B(n_449), .Y(n_507) );
AND2x2_ASAP7_75t_L g508 ( .A(n_404), .B(n_394), .Y(n_508) );
AND2x2_ASAP7_75t_L g509 ( .A(n_420), .B(n_398), .Y(n_509) );
CKINVDCx14_ASAP7_75t_R g510 ( .A(n_401), .Y(n_510) );
INVx1_ASAP7_75t_L g511 ( .A(n_431), .Y(n_511) );
OR2x2_ASAP7_75t_L g512 ( .A(n_453), .B(n_372), .Y(n_512) );
OR2x2_ASAP7_75t_L g513 ( .A(n_455), .B(n_372), .Y(n_513) );
AND2x4_ASAP7_75t_L g514 ( .A(n_463), .B(n_398), .Y(n_514) );
AND2x2_ASAP7_75t_L g515 ( .A(n_420), .B(n_383), .Y(n_515) );
INVx1_ASAP7_75t_L g516 ( .A(n_404), .Y(n_516) );
INVx1_ASAP7_75t_L g517 ( .A(n_404), .Y(n_517) );
BUFx3_ASAP7_75t_L g518 ( .A(n_401), .Y(n_518) );
AND2x2_ASAP7_75t_L g519 ( .A(n_427), .B(n_394), .Y(n_519) );
OR2x2_ASAP7_75t_L g520 ( .A(n_456), .B(n_371), .Y(n_520) );
INVx1_ASAP7_75t_L g521 ( .A(n_437), .Y(n_521) );
NAND2x1_ASAP7_75t_L g522 ( .A(n_432), .B(n_372), .Y(n_522) );
NAND2xp5_ASAP7_75t_L g523 ( .A(n_414), .B(n_386), .Y(n_523) );
HB1xp67_ASAP7_75t_L g524 ( .A(n_418), .Y(n_524) );
AND2x2_ASAP7_75t_L g525 ( .A(n_427), .B(n_394), .Y(n_525) );
BUFx3_ASAP7_75t_L g526 ( .A(n_443), .Y(n_526) );
AND2x2_ASAP7_75t_L g527 ( .A(n_414), .B(n_391), .Y(n_527) );
INVx2_ASAP7_75t_L g528 ( .A(n_418), .Y(n_528) );
INVx2_ASAP7_75t_L g529 ( .A(n_419), .Y(n_529) );
AND2x2_ASAP7_75t_L g530 ( .A(n_471), .B(n_391), .Y(n_530) );
INVx1_ASAP7_75t_L g531 ( .A(n_439), .Y(n_531) );
NAND2x1p5_ASAP7_75t_L g532 ( .A(n_432), .B(n_388), .Y(n_532) );
AND2x2_ASAP7_75t_L g533 ( .A(n_443), .B(n_361), .Y(n_533) );
NAND2xp5_ASAP7_75t_L g534 ( .A(n_441), .B(n_396), .Y(n_534) );
NAND2xp5_ASAP7_75t_L g535 ( .A(n_460), .B(n_396), .Y(n_535) );
INVx2_ASAP7_75t_L g536 ( .A(n_419), .Y(n_536) );
INVx1_ASAP7_75t_L g537 ( .A(n_467), .Y(n_537) );
INVx2_ASAP7_75t_L g538 ( .A(n_425), .Y(n_538) );
OR2x2_ASAP7_75t_L g539 ( .A(n_436), .B(n_383), .Y(n_539) );
INVx1_ASAP7_75t_L g540 ( .A(n_467), .Y(n_540) );
INVx1_ASAP7_75t_L g541 ( .A(n_425), .Y(n_541) );
INVx2_ASAP7_75t_L g542 ( .A(n_428), .Y(n_542) );
INVx2_ASAP7_75t_L g543 ( .A(n_428), .Y(n_543) );
INVx1_ASAP7_75t_L g544 ( .A(n_433), .Y(n_544) );
NAND2x1p5_ASAP7_75t_L g545 ( .A(n_432), .B(n_388), .Y(n_545) );
NAND2xp5_ASAP7_75t_L g546 ( .A(n_412), .B(n_400), .Y(n_546) );
INVx1_ASAP7_75t_L g547 ( .A(n_433), .Y(n_547) );
AND2x2_ASAP7_75t_L g548 ( .A(n_475), .B(n_361), .Y(n_548) );
AND2x4_ASAP7_75t_L g549 ( .A(n_463), .B(n_400), .Y(n_549) );
INVx1_ASAP7_75t_L g550 ( .A(n_448), .Y(n_550) );
INVx1_ASAP7_75t_L g551 ( .A(n_448), .Y(n_551) );
AND2x4_ASAP7_75t_L g552 ( .A(n_463), .B(n_400), .Y(n_552) );
HB1xp67_ASAP7_75t_L g553 ( .A(n_464), .Y(n_553) );
INVx1_ASAP7_75t_L g554 ( .A(n_464), .Y(n_554) );
AND2x2_ASAP7_75t_L g555 ( .A(n_475), .B(n_361), .Y(n_555) );
INVx1_ASAP7_75t_L g556 ( .A(n_465), .Y(n_556) );
INVx2_ASAP7_75t_SL g557 ( .A(n_475), .Y(n_557) );
INVxp67_ASAP7_75t_SL g558 ( .A(n_465), .Y(n_558) );
OR2x2_ASAP7_75t_L g559 ( .A(n_423), .B(n_399), .Y(n_559) );
INVx1_ASAP7_75t_L g560 ( .A(n_415), .Y(n_560) );
AND2x2_ASAP7_75t_L g561 ( .A(n_475), .B(n_388), .Y(n_561) );
HB1xp67_ASAP7_75t_L g562 ( .A(n_458), .Y(n_562) );
INVxp67_ASAP7_75t_L g563 ( .A(n_415), .Y(n_563) );
HB1xp67_ASAP7_75t_L g564 ( .A(n_458), .Y(n_564) );
AND2x2_ASAP7_75t_L g565 ( .A(n_471), .B(n_476), .Y(n_565) );
OR2x2_ASAP7_75t_L g566 ( .A(n_423), .B(n_399), .Y(n_566) );
INVx1_ASAP7_75t_L g567 ( .A(n_415), .Y(n_567) );
NAND2xp5_ASAP7_75t_L g568 ( .A(n_446), .B(n_399), .Y(n_568) );
INVx1_ASAP7_75t_L g569 ( .A(n_454), .Y(n_569) );
INVx3_ASAP7_75t_L g570 ( .A(n_447), .Y(n_570) );
INVx1_ASAP7_75t_L g571 ( .A(n_454), .Y(n_571) );
HB1xp67_ASAP7_75t_L g572 ( .A(n_473), .Y(n_572) );
INVxp67_ASAP7_75t_L g573 ( .A(n_440), .Y(n_573) );
AND2x4_ASAP7_75t_L g574 ( .A(n_478), .B(n_397), .Y(n_574) );
INVx1_ASAP7_75t_L g575 ( .A(n_472), .Y(n_575) );
INVx1_ASAP7_75t_L g576 ( .A(n_452), .Y(n_576) );
HB1xp67_ASAP7_75t_L g577 ( .A(n_473), .Y(n_577) );
NAND2xp5_ASAP7_75t_L g578 ( .A(n_446), .B(n_397), .Y(n_578) );
AND2x2_ASAP7_75t_L g579 ( .A(n_476), .B(n_397), .Y(n_579) );
AOI21xp5_ASAP7_75t_L g580 ( .A1(n_438), .A2(n_358), .B(n_330), .Y(n_580) );
INVx1_ASAP7_75t_L g581 ( .A(n_452), .Y(n_581) );
NAND2xp5_ASAP7_75t_SL g582 ( .A(n_573), .B(n_503), .Y(n_582) );
OR2x2_ASAP7_75t_L g583 ( .A(n_565), .B(n_426), .Y(n_583) );
AND2x2_ASAP7_75t_L g584 ( .A(n_504), .B(n_478), .Y(n_584) );
OR2x2_ASAP7_75t_L g585 ( .A(n_502), .B(n_434), .Y(n_585) );
NAND2xp5_ASAP7_75t_L g586 ( .A(n_537), .B(n_434), .Y(n_586) );
AND2x2_ASAP7_75t_L g587 ( .A(n_505), .B(n_477), .Y(n_587) );
NAND2x1p5_ASAP7_75t_L g588 ( .A(n_522), .B(n_445), .Y(n_588) );
NAND2xp5_ASAP7_75t_L g589 ( .A(n_540), .B(n_426), .Y(n_589) );
OAI21xp33_ASAP7_75t_L g590 ( .A1(n_573), .A2(n_442), .B(n_416), .Y(n_590) );
INVxp67_ASAP7_75t_L g591 ( .A(n_490), .Y(n_591) );
INVx1_ASAP7_75t_L g592 ( .A(n_484), .Y(n_592) );
NAND2xp5_ASAP7_75t_L g593 ( .A(n_576), .B(n_477), .Y(n_593) );
AND2x2_ASAP7_75t_L g594 ( .A(n_482), .B(n_461), .Y(n_594) );
HB1xp67_ASAP7_75t_L g595 ( .A(n_510), .Y(n_595) );
INVx1_ASAP7_75t_L g596 ( .A(n_487), .Y(n_596) );
NAND2xp5_ASAP7_75t_L g597 ( .A(n_581), .B(n_461), .Y(n_597) );
AND2x4_ASAP7_75t_L g598 ( .A(n_563), .B(n_474), .Y(n_598) );
INVx1_ASAP7_75t_L g599 ( .A(n_489), .Y(n_599) );
INVx1_ASAP7_75t_L g600 ( .A(n_496), .Y(n_600) );
INVx1_ASAP7_75t_L g601 ( .A(n_499), .Y(n_601) );
INVx2_ASAP7_75t_L g602 ( .A(n_479), .Y(n_602) );
AND2x2_ASAP7_75t_L g603 ( .A(n_510), .B(n_474), .Y(n_603) );
INVx2_ASAP7_75t_L g604 ( .A(n_479), .Y(n_604) );
HB1xp67_ASAP7_75t_L g605 ( .A(n_572), .Y(n_605) );
OR3x2_ASAP7_75t_L g606 ( .A(n_490), .B(n_445), .C(n_442), .Y(n_606) );
AND2x4_ASAP7_75t_L g607 ( .A(n_563), .B(n_474), .Y(n_607) );
OR2x2_ASAP7_75t_L g608 ( .A(n_515), .B(n_457), .Y(n_608) );
INVx1_ASAP7_75t_L g609 ( .A(n_500), .Y(n_609) );
AND2x2_ASAP7_75t_L g610 ( .A(n_495), .B(n_457), .Y(n_610) );
NAND2xp5_ASAP7_75t_L g611 ( .A(n_509), .B(n_468), .Y(n_611) );
AND2x2_ASAP7_75t_L g612 ( .A(n_495), .B(n_457), .Y(n_612) );
INVx1_ASAP7_75t_L g613 ( .A(n_506), .Y(n_613) );
AND2x4_ASAP7_75t_L g614 ( .A(n_514), .B(n_447), .Y(n_614) );
NAND2xp5_ASAP7_75t_L g615 ( .A(n_509), .B(n_389), .Y(n_615) );
OR2x2_ASAP7_75t_L g616 ( .A(n_515), .B(n_447), .Y(n_616) );
INVx1_ASAP7_75t_L g617 ( .A(n_511), .Y(n_617) );
INVxp67_ASAP7_75t_SL g618 ( .A(n_494), .Y(n_618) );
AND2x2_ASAP7_75t_L g619 ( .A(n_508), .B(n_416), .Y(n_619) );
INVx1_ASAP7_75t_L g620 ( .A(n_521), .Y(n_620) );
INVx1_ASAP7_75t_L g621 ( .A(n_531), .Y(n_621) );
NAND2xp5_ASAP7_75t_L g622 ( .A(n_527), .B(n_389), .Y(n_622) );
AND2x2_ASAP7_75t_L g623 ( .A(n_488), .B(n_450), .Y(n_623) );
INVx1_ASAP7_75t_L g624 ( .A(n_497), .Y(n_624) );
INVx1_ASAP7_75t_L g625 ( .A(n_485), .Y(n_625) );
CKINVDCx16_ASAP7_75t_R g626 ( .A(n_518), .Y(n_626) );
AND2x2_ASAP7_75t_L g627 ( .A(n_519), .B(n_450), .Y(n_627) );
INVx1_ASAP7_75t_L g628 ( .A(n_507), .Y(n_628) );
NAND2xp5_ASAP7_75t_L g629 ( .A(n_527), .B(n_389), .Y(n_629) );
AND2x2_ASAP7_75t_L g630 ( .A(n_525), .B(n_450), .Y(n_630) );
OR2x2_ASAP7_75t_L g631 ( .A(n_483), .B(n_491), .Y(n_631) );
INVx2_ASAP7_75t_L g632 ( .A(n_494), .Y(n_632) );
NOR2xp33_ASAP7_75t_L g633 ( .A(n_569), .B(n_450), .Y(n_633) );
INVx1_ASAP7_75t_L g634 ( .A(n_534), .Y(n_634) );
INVx1_ASAP7_75t_L g635 ( .A(n_516), .Y(n_635) );
INVx2_ASAP7_75t_L g636 ( .A(n_524), .Y(n_636) );
NAND2xp5_ASAP7_75t_L g637 ( .A(n_530), .B(n_389), .Y(n_637) );
AND2x4_ASAP7_75t_L g638 ( .A(n_514), .B(n_450), .Y(n_638) );
INVx1_ASAP7_75t_L g639 ( .A(n_517), .Y(n_639) );
INVx1_ASAP7_75t_L g640 ( .A(n_486), .Y(n_640) );
NAND2xp5_ASAP7_75t_L g641 ( .A(n_530), .B(n_389), .Y(n_641) );
OR2x2_ASAP7_75t_L g642 ( .A(n_559), .B(n_462), .Y(n_642) );
INVx2_ASAP7_75t_SL g643 ( .A(n_518), .Y(n_643) );
OAI21xp5_ASAP7_75t_SL g644 ( .A1(n_557), .A2(n_315), .B(n_358), .Y(n_644) );
INVx1_ASAP7_75t_L g645 ( .A(n_575), .Y(n_645) );
INVx1_ASAP7_75t_L g646 ( .A(n_524), .Y(n_646) );
INVx1_ASAP7_75t_L g647 ( .A(n_553), .Y(n_647) );
OR2x2_ASAP7_75t_L g648 ( .A(n_566), .B(n_358), .Y(n_648) );
AND2x2_ASAP7_75t_L g649 ( .A(n_579), .B(n_376), .Y(n_649) );
NOR2x1_ASAP7_75t_L g650 ( .A(n_526), .B(n_358), .Y(n_650) );
BUFx3_ASAP7_75t_L g651 ( .A(n_526), .Y(n_651) );
INVx2_ASAP7_75t_L g652 ( .A(n_553), .Y(n_652) );
OAI21xp33_ASAP7_75t_L g653 ( .A1(n_523), .A2(n_376), .B(n_357), .Y(n_653) );
INVx3_ASAP7_75t_L g654 ( .A(n_481), .Y(n_654) );
INVx2_ASAP7_75t_L g655 ( .A(n_512), .Y(n_655) );
OR2x2_ASAP7_75t_L g656 ( .A(n_568), .B(n_578), .Y(n_656) );
AND2x2_ASAP7_75t_L g657 ( .A(n_514), .B(n_376), .Y(n_657) );
OR2x2_ASAP7_75t_L g658 ( .A(n_572), .B(n_577), .Y(n_658) );
AND2x2_ASAP7_75t_L g659 ( .A(n_493), .B(n_358), .Y(n_659) );
INVx1_ASAP7_75t_SL g660 ( .A(n_577), .Y(n_660) );
INVx1_ASAP7_75t_L g661 ( .A(n_539), .Y(n_661) );
NAND2x1p5_ASAP7_75t_L g662 ( .A(n_557), .B(n_357), .Y(n_662) );
INVx2_ASAP7_75t_SL g663 ( .A(n_513), .Y(n_663) );
INVx1_ASAP7_75t_L g664 ( .A(n_558), .Y(n_664) );
INVx1_ASAP7_75t_L g665 ( .A(n_558), .Y(n_665) );
NAND2xp5_ASAP7_75t_L g666 ( .A(n_546), .B(n_357), .Y(n_666) );
AND2x2_ASAP7_75t_L g667 ( .A(n_560), .B(n_336), .Y(n_667) );
NAND2x1p5_ASAP7_75t_L g668 ( .A(n_571), .B(n_33), .Y(n_668) );
AND2x2_ASAP7_75t_L g669 ( .A(n_567), .B(n_34), .Y(n_669) );
INVx1_ASAP7_75t_L g670 ( .A(n_520), .Y(n_670) );
AND2x2_ASAP7_75t_L g671 ( .A(n_533), .B(n_35), .Y(n_671) );
INVx1_ASAP7_75t_L g672 ( .A(n_541), .Y(n_672) );
AOI21xp33_ASAP7_75t_L g673 ( .A1(n_535), .A2(n_561), .B(n_580), .Y(n_673) );
INVxp33_ASAP7_75t_L g674 ( .A(n_562), .Y(n_674) );
INVx2_ASAP7_75t_L g675 ( .A(n_480), .Y(n_675) );
OR2x2_ASAP7_75t_L g676 ( .A(n_574), .B(n_36), .Y(n_676) );
INVx1_ASAP7_75t_L g677 ( .A(n_544), .Y(n_677) );
OR2x2_ASAP7_75t_L g678 ( .A(n_574), .B(n_38), .Y(n_678) );
NAND2xp5_ASAP7_75t_L g679 ( .A(n_547), .B(n_330), .Y(n_679) );
NOR2xp67_ASAP7_75t_L g680 ( .A(n_562), .B(n_40), .Y(n_680) );
INVx2_ASAP7_75t_L g681 ( .A(n_480), .Y(n_681) );
AND2x2_ASAP7_75t_L g682 ( .A(n_548), .B(n_44), .Y(n_682) );
AND2x2_ASAP7_75t_L g683 ( .A(n_555), .B(n_46), .Y(n_683) );
INVx1_ASAP7_75t_L g684 ( .A(n_592), .Y(n_684) );
NAND2xp5_ASAP7_75t_L g685 ( .A(n_634), .B(n_574), .Y(n_685) );
NAND2xp5_ASAP7_75t_L g686 ( .A(n_640), .B(n_564), .Y(n_686) );
OR2x2_ASAP7_75t_L g687 ( .A(n_583), .B(n_564), .Y(n_687) );
OR2x2_ASAP7_75t_L g688 ( .A(n_656), .B(n_481), .Y(n_688) );
NOR4xp75_ASAP7_75t_L g689 ( .A(n_590), .B(n_570), .C(n_481), .D(n_545), .Y(n_689) );
AND2x2_ASAP7_75t_L g690 ( .A(n_587), .B(n_549), .Y(n_690) );
NAND2xp5_ASAP7_75t_L g691 ( .A(n_661), .B(n_556), .Y(n_691) );
NOR2xp33_ASAP7_75t_L g692 ( .A(n_591), .B(n_570), .Y(n_692) );
INVx2_ASAP7_75t_L g693 ( .A(n_660), .Y(n_693) );
AND2x2_ASAP7_75t_L g694 ( .A(n_594), .B(n_549), .Y(n_694) );
INVxp67_ASAP7_75t_L g695 ( .A(n_595), .Y(n_695) );
NAND2xp5_ASAP7_75t_SL g696 ( .A(n_626), .B(n_570), .Y(n_696) );
NAND2xp5_ASAP7_75t_L g697 ( .A(n_624), .B(n_554), .Y(n_697) );
INVx1_ASAP7_75t_L g698 ( .A(n_596), .Y(n_698) );
NAND2xp5_ASAP7_75t_L g699 ( .A(n_628), .B(n_551), .Y(n_699) );
OAI22xp5_ASAP7_75t_L g700 ( .A1(n_606), .A2(n_545), .B1(n_532), .B2(n_549), .Y(n_700) );
AND2x4_ASAP7_75t_L g701 ( .A(n_614), .B(n_552), .Y(n_701) );
OR2x2_ASAP7_75t_L g702 ( .A(n_631), .B(n_552), .Y(n_702) );
NAND2xp5_ASAP7_75t_L g703 ( .A(n_611), .B(n_550), .Y(n_703) );
OR2x2_ASAP7_75t_L g704 ( .A(n_658), .B(n_552), .Y(n_704) );
INVx1_ASAP7_75t_L g705 ( .A(n_599), .Y(n_705) );
NAND2xp5_ASAP7_75t_L g706 ( .A(n_611), .B(n_543), .Y(n_706) );
AND2x2_ASAP7_75t_L g707 ( .A(n_584), .B(n_532), .Y(n_707) );
NAND2xp5_ASAP7_75t_L g708 ( .A(n_625), .B(n_543), .Y(n_708) );
OR2x2_ASAP7_75t_L g709 ( .A(n_663), .B(n_542), .Y(n_709) );
INVx2_ASAP7_75t_SL g710 ( .A(n_651), .Y(n_710) );
OR2x2_ASAP7_75t_L g711 ( .A(n_585), .B(n_542), .Y(n_711) );
OR2x2_ASAP7_75t_L g712 ( .A(n_593), .B(n_538), .Y(n_712) );
OR2x2_ASAP7_75t_L g713 ( .A(n_593), .B(n_538), .Y(n_713) );
AND2x2_ASAP7_75t_L g714 ( .A(n_610), .B(n_536), .Y(n_714) );
NAND2xp5_ASAP7_75t_L g715 ( .A(n_605), .B(n_529), .Y(n_715) );
AOI21xp33_ASAP7_75t_SL g716 ( .A1(n_582), .A2(n_536), .B(n_529), .Y(n_716) );
INVx2_ASAP7_75t_L g717 ( .A(n_660), .Y(n_717) );
INVx2_ASAP7_75t_L g718 ( .A(n_602), .Y(n_718) );
NAND2xp5_ASAP7_75t_L g719 ( .A(n_670), .B(n_528), .Y(n_719) );
AND2x2_ASAP7_75t_L g720 ( .A(n_612), .B(n_528), .Y(n_720) );
INVx1_ASAP7_75t_L g721 ( .A(n_600), .Y(n_721) );
AND2x2_ASAP7_75t_L g722 ( .A(n_623), .B(n_501), .Y(n_722) );
OR2x2_ASAP7_75t_L g723 ( .A(n_597), .B(n_501), .Y(n_723) );
AOI211xp5_ASAP7_75t_L g724 ( .A1(n_590), .A2(n_498), .B(n_492), .C(n_51), .Y(n_724) );
INVx4_ASAP7_75t_L g725 ( .A(n_588), .Y(n_725) );
INVx1_ASAP7_75t_L g726 ( .A(n_601), .Y(n_726) );
NAND2xp5_ASAP7_75t_L g727 ( .A(n_645), .B(n_498), .Y(n_727) );
INVx1_ASAP7_75t_L g728 ( .A(n_609), .Y(n_728) );
INVx2_ASAP7_75t_L g729 ( .A(n_604), .Y(n_729) );
INVx1_ASAP7_75t_L g730 ( .A(n_613), .Y(n_730) );
OR2x2_ASAP7_75t_L g731 ( .A(n_597), .B(n_492), .Y(n_731) );
NAND2xp5_ASAP7_75t_L g732 ( .A(n_635), .B(n_47), .Y(n_732) );
NAND3x2_ASAP7_75t_L g733 ( .A(n_642), .B(n_50), .C(n_52), .Y(n_733) );
OR2x2_ASAP7_75t_L g734 ( .A(n_655), .B(n_59), .Y(n_734) );
OR2x2_ASAP7_75t_L g735 ( .A(n_586), .B(n_61), .Y(n_735) );
NAND2x1_ASAP7_75t_L g736 ( .A(n_643), .B(n_65), .Y(n_736) );
AND2x2_ASAP7_75t_L g737 ( .A(n_627), .B(n_67), .Y(n_737) );
INVx1_ASAP7_75t_L g738 ( .A(n_617), .Y(n_738) );
NOR2x1_ASAP7_75t_L g739 ( .A(n_644), .B(n_70), .Y(n_739) );
AOI22xp33_ASAP7_75t_L g740 ( .A1(n_657), .A2(n_71), .B1(n_72), .B2(n_73), .Y(n_740) );
INVx1_ASAP7_75t_L g741 ( .A(n_620), .Y(n_741) );
INVx1_ASAP7_75t_L g742 ( .A(n_621), .Y(n_742) );
INVx1_ASAP7_75t_L g743 ( .A(n_639), .Y(n_743) );
INVx1_ASAP7_75t_L g744 ( .A(n_672), .Y(n_744) );
OR2x2_ASAP7_75t_L g745 ( .A(n_586), .B(n_74), .Y(n_745) );
HB1xp67_ASAP7_75t_L g746 ( .A(n_618), .Y(n_746) );
AND2x2_ASAP7_75t_L g747 ( .A(n_630), .B(n_76), .Y(n_747) );
INVx4_ASAP7_75t_L g748 ( .A(n_668), .Y(n_748) );
OR2x2_ASAP7_75t_L g749 ( .A(n_589), .B(n_77), .Y(n_749) );
INVx1_ASAP7_75t_L g750 ( .A(n_677), .Y(n_750) );
NAND4xp25_ASAP7_75t_L g751 ( .A(n_673), .B(n_79), .C(n_81), .D(n_82), .Y(n_751) );
INVxp67_ASAP7_75t_L g752 ( .A(n_603), .Y(n_752) );
INVx3_ASAP7_75t_L g753 ( .A(n_654), .Y(n_753) );
BUFx2_ASAP7_75t_L g754 ( .A(n_614), .Y(n_754) );
INVxp67_ASAP7_75t_L g755 ( .A(n_633), .Y(n_755) );
AOI221xp5_ASAP7_75t_L g756 ( .A1(n_695), .A2(n_673), .B1(n_644), .B2(n_615), .C(n_674), .Y(n_756) );
INVx1_ASAP7_75t_L g757 ( .A(n_686), .Y(n_757) );
INVx1_ASAP7_75t_L g758 ( .A(n_697), .Y(n_758) );
INVx1_ASAP7_75t_L g759 ( .A(n_715), .Y(n_759) );
AND2x2_ASAP7_75t_L g760 ( .A(n_754), .B(n_619), .Y(n_760) );
HB1xp67_ASAP7_75t_L g761 ( .A(n_746), .Y(n_761) );
AOI22xp5_ASAP7_75t_L g762 ( .A1(n_755), .A2(n_659), .B1(n_589), .B2(n_649), .Y(n_762) );
INVx1_ASAP7_75t_L g763 ( .A(n_715), .Y(n_763) );
AOI22xp5_ASAP7_75t_L g764 ( .A1(n_725), .A2(n_629), .B1(n_622), .B2(n_641), .Y(n_764) );
INVx1_ASAP7_75t_L g765 ( .A(n_706), .Y(n_765) );
INVxp67_ASAP7_75t_L g766 ( .A(n_693), .Y(n_766) );
INVx1_ASAP7_75t_L g767 ( .A(n_684), .Y(n_767) );
NAND2xp5_ASAP7_75t_SL g768 ( .A(n_725), .B(n_680), .Y(n_768) );
INVxp67_ASAP7_75t_L g769 ( .A(n_717), .Y(n_769) );
OAI322xp33_ASAP7_75t_L g770 ( .A1(n_687), .A2(n_615), .A3(n_622), .B1(n_629), .B2(n_637), .C1(n_641), .C2(n_648), .Y(n_770) );
OAI21xp5_ASAP7_75t_SL g771 ( .A1(n_739), .A2(n_683), .B(n_682), .Y(n_771) );
AND2x2_ASAP7_75t_L g772 ( .A(n_694), .B(n_638), .Y(n_772) );
INVx1_ASAP7_75t_L g773 ( .A(n_698), .Y(n_773) );
OAI21xp33_ASAP7_75t_L g774 ( .A1(n_739), .A2(n_637), .B(n_650), .Y(n_774) );
INVx1_ASAP7_75t_L g775 ( .A(n_705), .Y(n_775) );
INVx2_ASAP7_75t_L g776 ( .A(n_709), .Y(n_776) );
AO22x1_ASAP7_75t_L g777 ( .A1(n_710), .A2(n_638), .B1(n_654), .B2(n_598), .Y(n_777) );
INVx2_ASAP7_75t_SL g778 ( .A(n_702), .Y(n_778) );
NOR2xp33_ASAP7_75t_L g779 ( .A(n_692), .B(n_616), .Y(n_779) );
INVx2_ASAP7_75t_L g780 ( .A(n_711), .Y(n_780) );
INVx1_ASAP7_75t_L g781 ( .A(n_721), .Y(n_781) );
NAND2xp5_ASAP7_75t_L g782 ( .A(n_726), .B(n_646), .Y(n_782) );
AND2x2_ASAP7_75t_SL g783 ( .A(n_748), .B(n_598), .Y(n_783) );
OR2x2_ASAP7_75t_L g784 ( .A(n_712), .B(n_647), .Y(n_784) );
INVx1_ASAP7_75t_L g785 ( .A(n_728), .Y(n_785) );
NOR2x1_ASAP7_75t_L g786 ( .A(n_748), .B(n_680), .Y(n_786) );
OAI22xp33_ASAP7_75t_L g787 ( .A1(n_751), .A2(n_608), .B1(n_676), .B2(n_678), .Y(n_787) );
INVx2_ASAP7_75t_SL g788 ( .A(n_690), .Y(n_788) );
INVx1_ASAP7_75t_L g789 ( .A(n_730), .Y(n_789) );
INVx1_ASAP7_75t_L g790 ( .A(n_738), .Y(n_790) );
NOR2x1_ASAP7_75t_L g791 ( .A(n_751), .B(n_671), .Y(n_791) );
INVxp67_ASAP7_75t_L g792 ( .A(n_741), .Y(n_792) );
INVx1_ASAP7_75t_SL g793 ( .A(n_701), .Y(n_793) );
AND2x2_ASAP7_75t_L g794 ( .A(n_701), .B(n_607), .Y(n_794) );
INVx2_ASAP7_75t_L g795 ( .A(n_722), .Y(n_795) );
INVx1_ASAP7_75t_L g796 ( .A(n_742), .Y(n_796) );
INVx1_ASAP7_75t_L g797 ( .A(n_761), .Y(n_797) );
OAI22xp5_ASAP7_75t_L g798 ( .A1(n_783), .A2(n_752), .B1(n_724), .B2(n_700), .Y(n_798) );
O2A1O1Ixp33_ASAP7_75t_L g799 ( .A1(n_761), .A2(n_716), .B(n_724), .C(n_736), .Y(n_799) );
AOI22xp33_ASAP7_75t_SL g800 ( .A1(n_793), .A2(n_700), .B1(n_733), .B2(n_707), .Y(n_800) );
OAI22xp33_ASAP7_75t_L g801 ( .A1(n_771), .A2(n_716), .B1(n_696), .B2(n_753), .Y(n_801) );
OAI22xp33_ASAP7_75t_L g802 ( .A1(n_793), .A2(n_753), .B1(n_688), .B2(n_704), .Y(n_802) );
OR2x2_ASAP7_75t_L g803 ( .A(n_759), .B(n_731), .Y(n_803) );
OAI22xp5_ASAP7_75t_L g804 ( .A1(n_791), .A2(n_685), .B1(n_703), .B2(n_723), .Y(n_804) );
NOR4xp25_ASAP7_75t_SL g805 ( .A(n_768), .B(n_689), .C(n_743), .D(n_750), .Y(n_805) );
INVxp67_ASAP7_75t_L g806 ( .A(n_782), .Y(n_806) );
NAND2xp5_ASAP7_75t_L g807 ( .A(n_763), .B(n_744), .Y(n_807) );
AOI22xp5_ASAP7_75t_L g808 ( .A1(n_787), .A2(n_699), .B1(n_691), .B2(n_720), .Y(n_808) );
OAI21xp5_ASAP7_75t_L g809 ( .A1(n_786), .A2(n_749), .B(n_735), .Y(n_809) );
AOI322xp5_ASAP7_75t_SL g810 ( .A1(n_760), .A2(n_714), .A3(n_689), .B1(n_747), .B2(n_737), .C1(n_669), .C2(n_667), .Y(n_810) );
OAI211xp5_ASAP7_75t_L g811 ( .A1(n_756), .A2(n_740), .B(n_653), .C(n_745), .Y(n_811) );
INVxp67_ASAP7_75t_L g812 ( .A(n_782), .Y(n_812) );
OR2x2_ASAP7_75t_L g813 ( .A(n_780), .B(n_713), .Y(n_813) );
NOR3xp33_ASAP7_75t_L g814 ( .A(n_756), .B(n_732), .C(n_708), .Y(n_814) );
AOI22xp5_ASAP7_75t_L g815 ( .A1(n_764), .A2(n_607), .B1(n_719), .B2(n_727), .Y(n_815) );
AOI21xp33_ASAP7_75t_L g816 ( .A1(n_774), .A2(n_734), .B(n_653), .Y(n_816) );
NAND2xp5_ASAP7_75t_L g817 ( .A(n_765), .B(n_729), .Y(n_817) );
AOI221xp5_ASAP7_75t_L g818 ( .A1(n_770), .A2(n_718), .B1(n_666), .B2(n_665), .C(n_664), .Y(n_818) );
OAI21xp5_ASAP7_75t_SL g819 ( .A1(n_800), .A2(n_762), .B(n_769), .Y(n_819) );
OAI21xp5_ASAP7_75t_SL g820 ( .A1(n_799), .A2(n_766), .B(n_769), .Y(n_820) );
OAI211xp5_ASAP7_75t_L g821 ( .A1(n_805), .A2(n_792), .B(n_766), .C(n_757), .Y(n_821) );
AOI22xp33_ASAP7_75t_L g822 ( .A1(n_814), .A2(n_758), .B1(n_792), .B2(n_796), .Y(n_822) );
OAI21xp33_ASAP7_75t_L g823 ( .A1(n_808), .A2(n_818), .B(n_804), .Y(n_823) );
AOI211xp5_ASAP7_75t_L g824 ( .A1(n_801), .A2(n_777), .B(n_779), .C(n_794), .Y(n_824) );
OAI221xp5_ASAP7_75t_SL g825 ( .A1(n_818), .A2(n_776), .B1(n_784), .B2(n_788), .C(n_778), .Y(n_825) );
NOR2xp33_ASAP7_75t_L g826 ( .A(n_806), .B(n_773), .Y(n_826) );
AOI221xp5_ASAP7_75t_SL g827 ( .A1(n_802), .A2(n_775), .B1(n_790), .B2(n_789), .C(n_785), .Y(n_827) );
NAND4xp25_ASAP7_75t_L g828 ( .A(n_798), .B(n_781), .C(n_767), .D(n_666), .Y(n_828) );
AND2x2_ASAP7_75t_L g829 ( .A(n_815), .B(n_772), .Y(n_829) );
NAND3xp33_ASAP7_75t_SL g830 ( .A(n_810), .B(n_662), .C(n_795), .Y(n_830) );
NAND2xp5_ASAP7_75t_L g831 ( .A(n_822), .B(n_812), .Y(n_831) );
OAI22xp5_ASAP7_75t_SL g832 ( .A1(n_824), .A2(n_809), .B1(n_797), .B2(n_811), .Y(n_832) );
INVxp67_ASAP7_75t_SL g833 ( .A(n_825), .Y(n_833) );
NAND4xp25_ASAP7_75t_L g834 ( .A(n_830), .B(n_816), .C(n_807), .D(n_817), .Y(n_834) );
NAND4xp25_ASAP7_75t_L g835 ( .A(n_823), .B(n_803), .C(n_813), .D(n_679), .Y(n_835) );
NOR3x1_ASAP7_75t_L g836 ( .A(n_828), .B(n_679), .C(n_87), .Y(n_836) );
OAI211xp5_ASAP7_75t_L g837 ( .A1(n_833), .A2(n_820), .B(n_821), .C(n_819), .Y(n_837) );
NAND2xp5_ASAP7_75t_L g838 ( .A(n_831), .B(n_822), .Y(n_838) );
NAND3xp33_ASAP7_75t_L g839 ( .A(n_834), .B(n_827), .C(n_826), .Y(n_839) );
NOR4xp25_ASAP7_75t_L g840 ( .A(n_835), .B(n_829), .C(n_652), .D(n_636), .Y(n_840) );
INVx2_ASAP7_75t_SL g841 ( .A(n_838), .Y(n_841) );
NAND4xp25_ASAP7_75t_L g842 ( .A(n_837), .B(n_836), .C(n_832), .D(n_632), .Y(n_842) );
OAI221xp5_ASAP7_75t_L g843 ( .A1(n_839), .A2(n_681), .B1(n_675), .B2(n_89), .C(n_91), .Y(n_843) );
INVx1_ASAP7_75t_L g844 ( .A(n_841), .Y(n_844) );
HB1xp67_ASAP7_75t_L g845 ( .A(n_842), .Y(n_845) );
AO21x2_ASAP7_75t_L g846 ( .A1(n_844), .A2(n_840), .B(n_843), .Y(n_846) );
XNOR2xp5_ASAP7_75t_L g847 ( .A(n_845), .B(n_85), .Y(n_847) );
AOI22x1_ASAP7_75t_L g848 ( .A1(n_847), .A2(n_844), .B1(n_94), .B2(n_95), .Y(n_848) );
INVx1_ASAP7_75t_L g849 ( .A(n_848), .Y(n_849) );
OA21x2_ASAP7_75t_L g850 ( .A1(n_849), .A2(n_846), .B(n_96), .Y(n_850) );
NAND2xp5_ASAP7_75t_L g851 ( .A(n_850), .B(n_846), .Y(n_851) );
OA21x2_ASAP7_75t_L g852 ( .A1(n_851), .A2(n_88), .B(n_97), .Y(n_852) );
AOI21xp33_ASAP7_75t_SL g853 ( .A1(n_852), .A2(n_98), .B(n_99), .Y(n_853) );
endmodule