module fake_jpeg_22792_n_335 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_335);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_335;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_6),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_9),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_10),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_10),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

BUFx10_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_10),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_1),
.Y(n_26)
);

CKINVDCx14_ASAP7_75t_R g27 ( 
.A(n_12),
.Y(n_27)
);

INVx13_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_2),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

INVx1_ASAP7_75t_SL g31 ( 
.A(n_3),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_5),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_15),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_32),
.Y(n_35)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_35),
.Y(n_62)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_32),
.Y(n_36)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_36),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_18),
.B(n_0),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_37),
.B(n_40),
.Y(n_59)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_30),
.Y(n_38)
);

INVx5_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_32),
.Y(n_39)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_39),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_31),
.B(n_15),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_32),
.Y(n_41)
);

INVx4_ASAP7_75t_SL g49 ( 
.A(n_41),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_32),
.Y(n_42)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_42),
.Y(n_47)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_30),
.Y(n_43)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_43),
.Y(n_46)
);

HB1xp67_ASAP7_75t_L g44 ( 
.A(n_19),
.Y(n_44)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_44),
.Y(n_56)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_19),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_45),
.B(n_22),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_39),
.Y(n_51)
);

INVx6_ASAP7_75t_L g89 ( 
.A(n_51),
.Y(n_89)
);

OAI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_38),
.A2(n_22),
.B1(n_28),
.B2(n_19),
.Y(n_52)
);

OAI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_52),
.A2(n_22),
.B1(n_28),
.B2(n_34),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_39),
.Y(n_53)
);

INVx11_ASAP7_75t_L g76 ( 
.A(n_53),
.Y(n_76)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_43),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_54),
.B(n_55),
.Y(n_92)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_43),
.Y(n_55)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_37),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_58),
.B(n_40),
.Y(n_82)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_60),
.Y(n_68)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_42),
.Y(n_61)
);

HB1xp67_ASAP7_75t_L g66 ( 
.A(n_61),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_L g63 ( 
.A1(n_58),
.A2(n_38),
.B1(n_19),
.B2(n_28),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_63),
.A2(n_80),
.B1(n_84),
.B2(n_86),
.Y(n_124)
);

AO22x2_ASAP7_75t_L g64 ( 
.A1(n_50),
.A2(n_42),
.B1(n_44),
.B2(n_35),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_64),
.A2(n_87),
.B1(n_91),
.B2(n_18),
.Y(n_106)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_62),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_65),
.B(n_69),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_50),
.A2(n_22),
.B1(n_36),
.B2(n_45),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_67),
.A2(n_83),
.B1(n_23),
.B2(n_30),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_59),
.Y(n_69)
);

BUFx12_ASAP7_75t_L g70 ( 
.A(n_47),
.Y(n_70)
);

INVx4_ASAP7_75t_L g122 ( 
.A(n_70),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_59),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_71),
.Y(n_95)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_48),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_72),
.B(n_79),
.Y(n_114)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_62),
.Y(n_73)
);

INVx4_ASAP7_75t_SL g115 ( 
.A(n_73),
.Y(n_115)
);

INVx5_ASAP7_75t_L g74 ( 
.A(n_57),
.Y(n_74)
);

BUFx10_ASAP7_75t_L g111 ( 
.A(n_74),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_L g116 ( 
.A1(n_75),
.A2(n_49),
.B1(n_27),
.B2(n_23),
.Y(n_116)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_62),
.Y(n_77)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_77),
.Y(n_120)
);

BUFx3_ASAP7_75t_L g78 ( 
.A(n_47),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_78),
.Y(n_98)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_48),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_56),
.A2(n_27),
.B1(n_34),
.B2(n_28),
.Y(n_80)
);

HB1xp67_ASAP7_75t_L g81 ( 
.A(n_49),
.Y(n_81)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_81),
.Y(n_96)
);

OAI21xp33_ASAP7_75t_L g101 ( 
.A1(n_82),
.A2(n_88),
.B(n_20),
.Y(n_101)
);

OA22x2_ASAP7_75t_L g83 ( 
.A1(n_46),
.A2(n_28),
.B1(n_35),
.B2(n_41),
.Y(n_83)
);

OAI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_46),
.A2(n_34),
.B1(n_25),
.B2(n_20),
.Y(n_84)
);

BUFx3_ASAP7_75t_L g85 ( 
.A(n_51),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_85),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_57),
.A2(n_31),
.B1(n_30),
.B2(n_41),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_54),
.A2(n_31),
.B1(n_30),
.B2(n_18),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_61),
.Y(n_88)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_51),
.Y(n_90)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_90),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_56),
.A2(n_27),
.B1(n_34),
.B2(n_18),
.Y(n_91)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_53),
.Y(n_93)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_93),
.Y(n_109)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_53),
.Y(n_94)
);

NAND2x1_ASAP7_75t_SL g103 ( 
.A(n_94),
.B(n_24),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_69),
.B(n_71),
.C(n_68),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_99),
.B(n_105),
.C(n_66),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_68),
.B(n_35),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_100),
.B(n_107),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_101),
.B(n_21),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_SL g102 ( 
.A1(n_64),
.A2(n_55),
.B(n_31),
.Y(n_102)
);

OAI21xp5_ASAP7_75t_SL g145 ( 
.A1(n_102),
.A2(n_113),
.B(n_33),
.Y(n_145)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_103),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_67),
.B(n_49),
.C(n_24),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_106),
.A2(n_121),
.B1(n_77),
.B2(n_76),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_88),
.B(n_24),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_92),
.B(n_24),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_108),
.B(n_110),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_72),
.B(n_24),
.Y(n_110)
);

AND2x4_ASAP7_75t_L g113 ( 
.A(n_64),
.B(n_24),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_L g133 ( 
.A1(n_116),
.A2(n_117),
.B1(n_74),
.B2(n_89),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_79),
.B(n_24),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_118),
.B(n_119),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_83),
.B(n_24),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_64),
.A2(n_86),
.B1(n_87),
.B2(n_83),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_83),
.B(n_70),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_123),
.B(n_0),
.Y(n_148)
);

XNOR2xp5_ASAP7_75t_L g125 ( 
.A(n_99),
.B(n_64),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_125),
.B(n_127),
.C(n_129),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_98),
.B(n_70),
.Y(n_126)
);

CKINVDCx14_ASAP7_75t_R g185 ( 
.A(n_126),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_105),
.B(n_78),
.C(n_85),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_112),
.B(n_93),
.Y(n_130)
);

CKINVDCx16_ASAP7_75t_R g183 ( 
.A(n_130),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_113),
.A2(n_89),
.B1(n_65),
.B2(n_73),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_SL g158 ( 
.A1(n_132),
.A2(n_145),
.B(n_147),
.Y(n_158)
);

AOI22xp33_ASAP7_75t_L g175 ( 
.A1(n_133),
.A2(n_143),
.B1(n_111),
.B2(n_109),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_134),
.B(n_123),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_135),
.A2(n_117),
.B1(n_102),
.B2(n_119),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_113),
.A2(n_94),
.B1(n_90),
.B2(n_76),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_136),
.A2(n_115),
.B1(n_103),
.B2(n_120),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_95),
.B(n_23),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_137),
.B(n_140),
.Y(n_154)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_112),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_139),
.B(n_142),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_L g140 ( 
.A(n_100),
.B(n_12),
.Y(n_140)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_114),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_L g143 ( 
.A1(n_113),
.A2(n_124),
.B1(n_106),
.B2(n_121),
.Y(n_143)
);

INVx3_ASAP7_75t_L g144 ( 
.A(n_111),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_144),
.B(n_153),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_98),
.B(n_21),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_146),
.B(n_150),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_L g147 ( 
.A1(n_113),
.A2(n_33),
.B(n_29),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_SL g169 ( 
.A1(n_148),
.A2(n_149),
.B(n_152),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_SL g149 ( 
.A(n_124),
.B(n_12),
.Y(n_149)
);

INVx1_ASAP7_75t_SL g150 ( 
.A(n_114),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_122),
.B(n_21),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_151),
.B(n_122),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_L g152 ( 
.A1(n_95),
.A2(n_33),
.B(n_29),
.Y(n_152)
);

INVx3_ASAP7_75t_L g153 ( 
.A(n_111),
.Y(n_153)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_130),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_155),
.B(n_157),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_156),
.A2(n_162),
.B1(n_164),
.B2(n_171),
.Y(n_187)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_128),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_159),
.B(n_163),
.Y(n_199)
);

AO22x1_ASAP7_75t_L g160 ( 
.A1(n_145),
.A2(n_116),
.B1(n_103),
.B2(n_107),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_SL g192 ( 
.A1(n_160),
.A2(n_167),
.B(n_178),
.Y(n_192)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_128),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_136),
.A2(n_96),
.B1(n_115),
.B2(n_118),
.Y(n_164)
);

AND2x2_ASAP7_75t_L g167 ( 
.A(n_125),
.B(n_110),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_138),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_168),
.Y(n_190)
);

AOI22xp33_ASAP7_75t_SL g171 ( 
.A1(n_144),
.A2(n_115),
.B1(n_120),
.B2(n_96),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_172),
.B(n_177),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_138),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_173),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_139),
.B(n_120),
.Y(n_174)
);

CKINVDCx16_ASAP7_75t_R g207 ( 
.A(n_174),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_L g217 ( 
.A1(n_175),
.A2(n_15),
.B1(n_14),
.B2(n_11),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_137),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_176),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_153),
.B(n_122),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_152),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_141),
.B(n_108),
.Y(n_179)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_179),
.Y(n_188)
);

BUFx2_ASAP7_75t_L g180 ( 
.A(n_150),
.Y(n_180)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_180),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_142),
.B(n_109),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_181),
.B(n_186),
.Y(n_195)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_129),
.Y(n_182)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_182),
.Y(n_191)
);

BUFx2_ASAP7_75t_L g184 ( 
.A(n_132),
.Y(n_184)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_184),
.Y(n_193)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_141),
.Y(n_186)
);

AOI21xp5_ASAP7_75t_L g194 ( 
.A1(n_158),
.A2(n_131),
.B(n_127),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_L g224 ( 
.A1(n_194),
.A2(n_206),
.B1(n_216),
.B2(n_178),
.Y(n_224)
);

OAI32xp33_ASAP7_75t_L g196 ( 
.A1(n_160),
.A2(n_148),
.A3(n_131),
.B1(n_149),
.B2(n_135),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_196),
.B(n_198),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_157),
.B(n_140),
.Y(n_197)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_197),
.Y(n_219)
);

OAI32xp33_ASAP7_75t_L g198 ( 
.A1(n_160),
.A2(n_147),
.A3(n_134),
.B1(n_97),
.B2(n_111),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g200 ( 
.A(n_161),
.B(n_111),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_200),
.B(n_211),
.C(n_169),
.Y(n_229)
);

NAND3xp33_ASAP7_75t_L g201 ( 
.A(n_154),
.B(n_163),
.C(n_155),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_201),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_161),
.B(n_97),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_202),
.B(n_169),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_186),
.A2(n_104),
.B1(n_29),
.B2(n_26),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_204),
.A2(n_213),
.B1(n_214),
.B2(n_217),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_SL g206 ( 
.A1(n_158),
.A2(n_104),
.B(n_26),
.Y(n_206)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_174),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_208),
.B(n_215),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_182),
.B(n_26),
.C(n_17),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_209),
.B(n_176),
.C(n_170),
.Y(n_244)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_166),
.Y(n_210)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_210),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_168),
.B(n_17),
.C(n_16),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_162),
.A2(n_17),
.B1(n_16),
.B2(n_25),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_173),
.A2(n_16),
.B1(n_25),
.B2(n_20),
.Y(n_214)
);

INVxp67_ASAP7_75t_L g215 ( 
.A(n_172),
.Y(n_215)
);

OAI32xp33_ASAP7_75t_L g216 ( 
.A1(n_156),
.A2(n_0),
.A3(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_216)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_195),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_220),
.B(n_226),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_193),
.A2(n_164),
.B1(n_184),
.B2(n_179),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_221),
.A2(n_224),
.B1(n_236),
.B2(n_213),
.Y(n_258)
);

INVxp67_ASAP7_75t_L g226 ( 
.A(n_205),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_190),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_SL g247 ( 
.A(n_228),
.B(n_231),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_229),
.B(n_234),
.C(n_243),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_230),
.B(n_206),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_203),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_195),
.Y(n_232)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_232),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_200),
.B(n_167),
.C(n_154),
.Y(n_234)
);

AO21x2_ASAP7_75t_SL g235 ( 
.A1(n_193),
.A2(n_184),
.B(n_180),
.Y(n_235)
);

AOI21xp5_ASAP7_75t_L g263 ( 
.A1(n_235),
.A2(n_189),
.B(n_210),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_192),
.A2(n_183),
.B1(n_167),
.B2(n_165),
.Y(n_236)
);

INVxp67_ASAP7_75t_L g237 ( 
.A(n_187),
.Y(n_237)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_237),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_194),
.B(n_159),
.Y(n_238)
);

XOR2xp5_ASAP7_75t_L g252 ( 
.A(n_238),
.B(n_198),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_212),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_L g260 ( 
.A1(n_239),
.A2(n_240),
.B1(n_241),
.B2(n_242),
.Y(n_260)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_199),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_218),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_204),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_202),
.B(n_185),
.C(n_165),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_244),
.B(n_183),
.C(n_170),
.Y(n_261)
);

OAI21xp5_ASAP7_75t_L g245 ( 
.A1(n_235),
.A2(n_225),
.B(n_237),
.Y(n_245)
);

OAI21xp5_ASAP7_75t_SL g269 ( 
.A1(n_245),
.A2(n_255),
.B(n_262),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_225),
.A2(n_192),
.B1(n_188),
.B2(n_191),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_246),
.A2(n_251),
.B1(n_264),
.B2(n_221),
.Y(n_268)
);

FAx1_ASAP7_75t_SL g248 ( 
.A(n_236),
.B(n_197),
.CI(n_196),
.CON(n_248),
.SN(n_248)
);

NAND2xp5_ASAP7_75t_SL g281 ( 
.A(n_248),
.B(n_223),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_222),
.A2(n_188),
.B1(n_191),
.B2(n_215),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g270 ( 
.A(n_252),
.B(n_254),
.Y(n_270)
);

OAI21xp5_ASAP7_75t_L g255 ( 
.A1(n_235),
.A2(n_207),
.B(n_208),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_234),
.B(n_209),
.Y(n_256)
);

XOR2xp5_ASAP7_75t_L g283 ( 
.A(n_256),
.B(n_214),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_SL g282 ( 
.A(n_258),
.B(n_181),
.Y(n_282)
);

HB1xp67_ASAP7_75t_L g259 ( 
.A(n_235),
.Y(n_259)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_259),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_261),
.B(n_219),
.C(n_244),
.Y(n_276)
);

INVxp67_ASAP7_75t_L g262 ( 
.A(n_233),
.Y(n_262)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_263),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_L g264 ( 
.A1(n_223),
.A2(n_220),
.B1(n_232),
.B2(n_233),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_230),
.B(n_216),
.Y(n_265)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_265),
.B(n_238),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_253),
.B(n_243),
.C(n_229),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_266),
.B(n_275),
.C(n_276),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_SL g298 ( 
.A1(n_268),
.A2(n_281),
.B1(n_248),
.B2(n_254),
.Y(n_298)
);

HB1xp67_ASAP7_75t_L g272 ( 
.A(n_262),
.Y(n_272)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_272),
.Y(n_285)
);

XOR2xp5_ASAP7_75t_L g290 ( 
.A(n_273),
.B(n_283),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_247),
.B(n_180),
.Y(n_274)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_274),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_253),
.B(n_219),
.C(n_189),
.Y(n_275)
);

CKINVDCx16_ASAP7_75t_R g277 ( 
.A(n_250),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_277),
.B(n_280),
.Y(n_286)
);

AND2x2_ASAP7_75t_L g278 ( 
.A(n_251),
.B(n_226),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_278),
.Y(n_287)
);

BUFx24_ASAP7_75t_SL g279 ( 
.A(n_260),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_279),
.B(n_258),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_256),
.B(n_227),
.C(n_211),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_282),
.B(n_265),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g304 ( 
.A(n_284),
.B(n_295),
.Y(n_304)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_288),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_SL g291 ( 
.A(n_275),
.B(n_261),
.Y(n_291)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_291),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_267),
.A2(n_257),
.B1(n_246),
.B2(n_249),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_SL g299 ( 
.A1(n_292),
.A2(n_248),
.B1(n_283),
.B2(n_270),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_271),
.A2(n_263),
.B1(n_269),
.B2(n_278),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_293),
.A2(n_270),
.B1(n_1),
.B2(n_2),
.Y(n_300)
);

INVxp67_ASAP7_75t_L g294 ( 
.A(n_282),
.Y(n_294)
);

AOI21xp5_ASAP7_75t_L g301 ( 
.A1(n_294),
.A2(n_296),
.B(n_14),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_L g295 ( 
.A(n_273),
.B(n_252),
.Y(n_295)
);

OAI21xp5_ASAP7_75t_L g296 ( 
.A1(n_266),
.A2(n_245),
.B(n_255),
.Y(n_296)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_298),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_299),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_SL g312 ( 
.A(n_300),
.B(n_306),
.Y(n_312)
);

AOI21xp5_ASAP7_75t_L g314 ( 
.A1(n_301),
.A2(n_309),
.B(n_285),
.Y(n_314)
);

AOI21xp5_ASAP7_75t_L g302 ( 
.A1(n_296),
.A2(n_11),
.B(n_1),
.Y(n_302)
);

OAI21xp5_ASAP7_75t_SL g313 ( 
.A1(n_302),
.A2(n_308),
.B(n_289),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_SL g306 ( 
.A1(n_293),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_SL g307 ( 
.A1(n_287),
.A2(n_11),
.B1(n_4),
.B2(n_5),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_L g317 ( 
.A(n_307),
.B(n_290),
.Y(n_317)
);

AOI21xp5_ASAP7_75t_L g308 ( 
.A1(n_294),
.A2(n_3),
.B(n_4),
.Y(n_308)
);

NOR2xp67_ASAP7_75t_SL g309 ( 
.A(n_297),
.B(n_4),
.Y(n_309)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_313),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_314),
.Y(n_324)
);

OR2x2_ASAP7_75t_L g315 ( 
.A(n_306),
.B(n_284),
.Y(n_315)
);

AOI21xp5_ASAP7_75t_SL g322 ( 
.A1(n_315),
.A2(n_319),
.B(n_6),
.Y(n_322)
);

OAI22xp5_ASAP7_75t_SL g316 ( 
.A1(n_310),
.A2(n_286),
.B1(n_297),
.B2(n_295),
.Y(n_316)
);

XOR2xp5_ASAP7_75t_L g321 ( 
.A(n_316),
.B(n_304),
.Y(n_321)
);

XNOR2xp5_ASAP7_75t_L g326 ( 
.A(n_317),
.B(n_7),
.Y(n_326)
);

OAI21x1_ASAP7_75t_L g318 ( 
.A1(n_304),
.A2(n_290),
.B(n_7),
.Y(n_318)
);

AOI21xp33_ASAP7_75t_L g325 ( 
.A1(n_318),
.A2(n_6),
.B(n_7),
.Y(n_325)
);

OAI21xp5_ASAP7_75t_L g319 ( 
.A1(n_305),
.A2(n_6),
.B(n_7),
.Y(n_319)
);

OAI21xp5_ASAP7_75t_SL g320 ( 
.A1(n_311),
.A2(n_300),
.B(n_303),
.Y(n_320)
);

AOI21xp5_ASAP7_75t_SL g329 ( 
.A1(n_320),
.A2(n_325),
.B(n_326),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_SL g327 ( 
.A(n_321),
.B(n_322),
.Y(n_327)
);

OAI21xp5_ASAP7_75t_L g328 ( 
.A1(n_323),
.A2(n_312),
.B(n_315),
.Y(n_328)
);

A2O1A1O1Ixp25_ASAP7_75t_L g330 ( 
.A1(n_328),
.A2(n_322),
.B(n_319),
.C(n_317),
.D(n_324),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_330),
.B(n_327),
.C(n_329),
.Y(n_331)
);

NAND2xp33_ASAP7_75t_L g332 ( 
.A(n_331),
.B(n_8),
.Y(n_332)
);

XOR2xp5_ASAP7_75t_L g333 ( 
.A(n_332),
.B(n_8),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_333),
.B(n_8),
.C(n_9),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_334),
.B(n_9),
.C(n_331),
.Y(n_335)
);


endmodule