module fake_jpeg_30299_n_160 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_160);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_160;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx2_ASAP7_75t_L g50 ( 
.A(n_26),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_16),
.Y(n_51)
);

BUFx10_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_34),
.Y(n_53)
);

BUFx5_ASAP7_75t_L g54 ( 
.A(n_47),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_41),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_14),
.B(n_13),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_20),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_22),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_4),
.Y(n_59)
);

BUFx12_ASAP7_75t_L g60 ( 
.A(n_3),
.Y(n_60)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_18),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_36),
.Y(n_62)
);

BUFx5_ASAP7_75t_L g63 ( 
.A(n_46),
.Y(n_63)
);

INVxp67_ASAP7_75t_L g64 ( 
.A(n_12),
.Y(n_64)
);

INVx2_ASAP7_75t_SL g65 ( 
.A(n_5),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_35),
.Y(n_66)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_32),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_17),
.Y(n_68)
);

HB1xp67_ASAP7_75t_L g69 ( 
.A(n_42),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_6),
.Y(n_70)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_9),
.Y(n_71)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_71),
.Y(n_72)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_72),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_55),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_73),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_59),
.B(n_0),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_74),
.Y(n_84)
);

INVx6_ASAP7_75t_L g75 ( 
.A(n_55),
.Y(n_75)
);

BUFx2_ASAP7_75t_L g93 ( 
.A(n_75),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_70),
.B(n_0),
.Y(n_76)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_76),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_58),
.Y(n_77)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_77),
.Y(n_91)
);

INVx5_ASAP7_75t_L g78 ( 
.A(n_54),
.Y(n_78)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_78),
.Y(n_92)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_63),
.Y(n_79)
);

HB1xp67_ASAP7_75t_L g88 ( 
.A(n_79),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_58),
.Y(n_80)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_80),
.Y(n_87)
);

AOI21xp5_ASAP7_75t_L g81 ( 
.A1(n_79),
.A2(n_65),
.B(n_64),
.Y(n_81)
);

OAI21xp5_ASAP7_75t_SL g106 ( 
.A1(n_81),
.A2(n_94),
.B(n_52),
.Y(n_106)
);

AOI222xp33_ASAP7_75t_L g83 ( 
.A1(n_77),
.A2(n_53),
.B1(n_51),
.B2(n_66),
.C1(n_57),
.C2(n_56),
.Y(n_83)
);

A2O1A1Ixp33_ASAP7_75t_L g104 ( 
.A1(n_83),
.A2(n_82),
.B(n_52),
.C(n_61),
.Y(n_104)
);

INVx1_ASAP7_75t_SL g86 ( 
.A(n_78),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_86),
.B(n_61),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_75),
.A2(n_50),
.B1(n_69),
.B2(n_67),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_90),
.A2(n_52),
.B1(n_61),
.B2(n_60),
.Y(n_102)
);

A2O1A1Ixp33_ASAP7_75t_L g94 ( 
.A1(n_72),
.A2(n_64),
.B(n_68),
.C(n_62),
.Y(n_94)
);

INVxp67_ASAP7_75t_L g95 ( 
.A(n_88),
.Y(n_95)
);

INVx13_ASAP7_75t_L g123 ( 
.A(n_95),
.Y(n_123)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_87),
.Y(n_96)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_96),
.Y(n_118)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_88),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_97),
.B(n_103),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_84),
.B(n_65),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_98),
.B(n_112),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_94),
.A2(n_80),
.B1(n_73),
.B2(n_69),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_99),
.A2(n_110),
.B1(n_15),
.B2(n_19),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_89),
.B(n_80),
.C(n_73),
.Y(n_100)
);

XOR2xp5_ASAP7_75t_L g116 ( 
.A(n_100),
.B(n_102),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_93),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_101),
.B(n_104),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_102),
.A2(n_108),
.B1(n_11),
.B2(n_12),
.Y(n_127)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_91),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_93),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_105),
.B(n_106),
.Y(n_117)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_107),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_L g108 ( 
.A1(n_85),
.A2(n_60),
.B1(n_2),
.B2(n_3),
.Y(n_108)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_92),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_109),
.B(n_7),
.Y(n_119)
);

AO21x1_ASAP7_75t_SL g110 ( 
.A1(n_92),
.A2(n_1),
.B(n_2),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_89),
.A2(n_1),
.B1(n_4),
.B2(n_5),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_111),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_84),
.B(n_6),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_84),
.B(n_7),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_113),
.B(n_11),
.Y(n_126)
);

XNOR2xp5_ASAP7_75t_L g138 ( 
.A(n_116),
.B(n_33),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_119),
.B(n_129),
.Y(n_136)
);

AOI21xp5_ASAP7_75t_L g120 ( 
.A1(n_95),
.A2(n_28),
.B(n_48),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_SL g137 ( 
.A1(n_120),
.A2(n_124),
.B(n_31),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_104),
.B(n_8),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_122),
.B(n_125),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_100),
.B(n_10),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_126),
.B(n_44),
.Y(n_144)
);

AND2x2_ASAP7_75t_L g143 ( 
.A(n_127),
.B(n_128),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_103),
.A2(n_21),
.B1(n_23),
.B2(n_24),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_129),
.B(n_132),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_111),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_131),
.B(n_39),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_110),
.B(n_49),
.Y(n_132)
);

OR2x2_ASAP7_75t_L g134 ( 
.A(n_117),
.B(n_25),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_134),
.B(n_136),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_SL g135 ( 
.A1(n_118),
.A2(n_27),
.B1(n_29),
.B2(n_30),
.Y(n_135)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_135),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_L g150 ( 
.A(n_137),
.B(n_138),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_L g139 ( 
.A(n_121),
.B(n_37),
.Y(n_139)
);

XOR2xp5_ASAP7_75t_L g148 ( 
.A(n_139),
.B(n_142),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_SL g140 ( 
.A(n_130),
.B(n_45),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_SL g151 ( 
.A(n_140),
.B(n_144),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_114),
.B(n_40),
.Y(n_145)
);

A2O1A1O1Ixp25_ASAP7_75t_L g147 ( 
.A1(n_145),
.A2(n_115),
.B(n_120),
.C(n_43),
.D(n_130),
.Y(n_147)
);

A2O1A1O1Ixp25_ASAP7_75t_L g154 ( 
.A1(n_147),
.A2(n_145),
.B(n_123),
.C(n_143),
.D(n_127),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_149),
.A2(n_143),
.B1(n_128),
.B2(n_136),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_SL g155 ( 
.A(n_152),
.B(n_153),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_L g153 ( 
.A1(n_146),
.A2(n_133),
.B(n_141),
.Y(n_153)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_155),
.Y(n_156)
);

OAI31xp33_ASAP7_75t_L g157 ( 
.A1(n_156),
.A2(n_147),
.A3(n_154),
.B(n_151),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_157),
.B(n_150),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_158),
.B(n_148),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_159),
.B(n_116),
.Y(n_160)
);


endmodule