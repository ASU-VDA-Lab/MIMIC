module fake_netlist_5_1564_n_2381 (n_137, n_210, n_168, n_164, n_191, n_91, n_208, n_82, n_122, n_194, n_142, n_176, n_10, n_214, n_140, n_24, n_124, n_86, n_136, n_146, n_182, n_143, n_83, n_132, n_61, n_237, n_90, n_127, n_75, n_101, n_180, n_184, n_226, n_235, n_65, n_78, n_74, n_144, n_207, n_114, n_57, n_96, n_37, n_189, n_220, n_165, n_111, n_229, n_108, n_231, n_213, n_129, n_31, n_13, n_66, n_98, n_177, n_60, n_155, n_152, n_197, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_236, n_18, n_116, n_195, n_42, n_22, n_227, n_1, n_45, n_117, n_46, n_233, n_21, n_94, n_203, n_205, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_179, n_125, n_35, n_167, n_128, n_73, n_234, n_17, n_92, n_19, n_149, n_120, n_232, n_135, n_30, n_156, n_5, n_33, n_126, n_14, n_225, n_84, n_23, n_202, n_130, n_219, n_157, n_29, n_79, n_193, n_131, n_151, n_47, n_173, n_192, n_25, n_53, n_160, n_198, n_223, n_188, n_190, n_8, n_201, n_158, n_44, n_224, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_228, n_109, n_112, n_212, n_85, n_159, n_163, n_95, n_119, n_183, n_185, n_175, n_169, n_59, n_26, n_133, n_215, n_55, n_196, n_99, n_2, n_211, n_218, n_181, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_178, n_221, n_12, n_67, n_121, n_36, n_76, n_200, n_87, n_150, n_162, n_27, n_170, n_64, n_77, n_102, n_106, n_161, n_209, n_222, n_230, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_174, n_186, n_199, n_134, n_187, n_32, n_41, n_104, n_172, n_103, n_56, n_51, n_63, n_97, n_141, n_166, n_11, n_206, n_217, n_171, n_153, n_7, n_15, n_145, n_48, n_204, n_50, n_52, n_88, n_110, n_216, n_2381);

input n_137;
input n_210;
input n_168;
input n_164;
input n_191;
input n_91;
input n_208;
input n_82;
input n_122;
input n_194;
input n_142;
input n_176;
input n_10;
input n_214;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_182;
input n_143;
input n_83;
input n_132;
input n_61;
input n_237;
input n_90;
input n_127;
input n_75;
input n_101;
input n_180;
input n_184;
input n_226;
input n_235;
input n_65;
input n_78;
input n_74;
input n_144;
input n_207;
input n_114;
input n_57;
input n_96;
input n_37;
input n_189;
input n_220;
input n_165;
input n_111;
input n_229;
input n_108;
input n_231;
input n_213;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_177;
input n_60;
input n_155;
input n_152;
input n_197;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_236;
input n_18;
input n_116;
input n_195;
input n_42;
input n_22;
input n_227;
input n_1;
input n_45;
input n_117;
input n_46;
input n_233;
input n_21;
input n_94;
input n_203;
input n_205;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_179;
input n_125;
input n_35;
input n_167;
input n_128;
input n_73;
input n_234;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_232;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_14;
input n_225;
input n_84;
input n_23;
input n_202;
input n_130;
input n_219;
input n_157;
input n_29;
input n_79;
input n_193;
input n_131;
input n_151;
input n_47;
input n_173;
input n_192;
input n_25;
input n_53;
input n_160;
input n_198;
input n_223;
input n_188;
input n_190;
input n_8;
input n_201;
input n_158;
input n_44;
input n_224;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_228;
input n_109;
input n_112;
input n_212;
input n_85;
input n_159;
input n_163;
input n_95;
input n_119;
input n_183;
input n_185;
input n_175;
input n_169;
input n_59;
input n_26;
input n_133;
input n_215;
input n_55;
input n_196;
input n_99;
input n_2;
input n_211;
input n_218;
input n_181;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_178;
input n_221;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_200;
input n_87;
input n_150;
input n_162;
input n_27;
input n_170;
input n_64;
input n_77;
input n_102;
input n_106;
input n_161;
input n_209;
input n_222;
input n_230;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_174;
input n_186;
input n_199;
input n_134;
input n_187;
input n_32;
input n_41;
input n_104;
input n_172;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_166;
input n_11;
input n_206;
input n_217;
input n_171;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_204;
input n_50;
input n_52;
input n_88;
input n_110;
input n_216;

output n_2381;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_2253;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1729;
wire n_1166;
wire n_2380;
wire n_1751;
wire n_469;
wire n_1508;
wire n_785;
wire n_549;
wire n_2200;
wire n_532;
wire n_1161;
wire n_1859;
wire n_1677;
wire n_1150;
wire n_2327;
wire n_1780;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_1501;
wire n_880;
wire n_544;
wire n_1007;
wire n_2369;
wire n_552;
wire n_1528;
wire n_1370;
wire n_1292;
wire n_2347;
wire n_1198;
wire n_1360;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1738;
wire n_2021;
wire n_2134;
wire n_1021;
wire n_1960;
wire n_2185;
wire n_551;
wire n_2143;
wire n_2059;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1695;
wire n_1353;
wire n_800;
wire n_1347;
wire n_1535;
wire n_1789;
wire n_1666;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_2302;
wire n_915;
wire n_1545;
wire n_2374;
wire n_864;
wire n_859;
wire n_951;
wire n_1947;
wire n_1264;
wire n_2114;
wire n_447;
wire n_247;
wire n_2001;
wire n_1494;
wire n_292;
wire n_625;
wire n_854;
wire n_1462;
wire n_1799;
wire n_2069;
wire n_1580;
wire n_674;
wire n_417;
wire n_1939;
wire n_1806;
wire n_516;
wire n_933;
wire n_2244;
wire n_2257;
wire n_1152;
wire n_497;
wire n_1869;
wire n_1607;
wire n_1563;
wire n_606;
wire n_275;
wire n_2011;
wire n_2096;
wire n_877;
wire n_2105;
wire n_2024;
wire n_1696;
wire n_755;
wire n_1118;
wire n_1686;
wire n_947;
wire n_1285;
wire n_373;
wire n_307;
wire n_1860;
wire n_1359;
wire n_530;
wire n_1107;
wire n_1728;
wire n_556;
wire n_2076;
wire n_2031;
wire n_1230;
wire n_668;
wire n_375;
wire n_301;
wire n_1896;
wire n_2165;
wire n_2147;
wire n_929;
wire n_1124;
wire n_1818;
wire n_2127;
wire n_902;
wire n_1576;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1705;
wire n_1257;
wire n_1182;
wire n_579;
wire n_1698;
wire n_1261;
wire n_2329;
wire n_938;
wire n_1098;
wire n_2142;
wire n_320;
wire n_1154;
wire n_2189;
wire n_1242;
wire n_1135;
wire n_406;
wire n_519;
wire n_2323;
wire n_2203;
wire n_1016;
wire n_1243;
wire n_546;
wire n_2047;
wire n_1280;
wire n_1845;
wire n_281;
wire n_240;
wire n_2052;
wire n_2193;
wire n_2058;
wire n_291;
wire n_257;
wire n_731;
wire n_371;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_317;
wire n_1236;
wire n_1633;
wire n_569;
wire n_2144;
wire n_1778;
wire n_2306;
wire n_920;
wire n_1289;
wire n_1517;
wire n_2091;
wire n_335;
wire n_2085;
wire n_1669;
wire n_370;
wire n_976;
wire n_1949;
wire n_343;
wire n_1449;
wire n_308;
wire n_1946;
wire n_1566;
wire n_2032;
wire n_297;
wire n_2149;
wire n_1078;
wire n_1670;
wire n_775;
wire n_600;
wire n_1484;
wire n_2071;
wire n_1374;
wire n_1328;
wire n_2141;
wire n_1948;
wire n_1984;
wire n_2099;
wire n_264;
wire n_1877;
wire n_1831;
wire n_1598;
wire n_1723;
wire n_955;
wire n_1850;
wire n_339;
wire n_1146;
wire n_882;
wire n_243;
wire n_1097;
wire n_1036;
wire n_1749;
wire n_347;
wire n_550;
wire n_696;
wire n_897;
wire n_798;
wire n_350;
wire n_646;
wire n_1428;
wire n_436;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_290;
wire n_580;
wire n_1040;
wire n_2202;
wire n_1872;
wire n_1852;
wire n_2159;
wire n_578;
wire n_926;
wire n_2180;
wire n_2249;
wire n_344;
wire n_2353;
wire n_1218;
wire n_1931;
wire n_2276;
wire n_475;
wire n_422;
wire n_777;
wire n_1070;
wire n_1547;
wire n_2089;
wire n_1030;
wire n_1755;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_1561;
wire n_496;
wire n_1801;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_1600;
wire n_521;
wire n_663;
wire n_845;
wire n_2235;
wire n_1862;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_2300;
wire n_1796;
wire n_680;
wire n_1473;
wire n_1587;
wire n_395;
wire n_901;
wire n_553;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_2174;
wire n_1748;
wire n_1672;
wire n_675;
wire n_888;
wire n_1880;
wire n_2337;
wire n_1167;
wire n_1626;
wire n_637;
wire n_1384;
wire n_1556;
wire n_446;
wire n_1863;
wire n_1064;
wire n_858;
wire n_2079;
wire n_2238;
wire n_923;
wire n_2118;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_1706;
wire n_468;
wire n_342;
wire n_464;
wire n_363;
wire n_1582;
wire n_1069;
wire n_1784;
wire n_1075;
wire n_1836;
wire n_1450;
wire n_1322;
wire n_2101;
wire n_1471;
wire n_1986;
wire n_2072;
wire n_1750;
wire n_1459;
wire n_460;
wire n_889;
wire n_2358;
wire n_973;
wire n_1700;
wire n_477;
wire n_571;
wire n_1585;
wire n_461;
wire n_1971;
wire n_1599;
wire n_2275;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_1950;
wire n_907;
wire n_1447;
wire n_2251;
wire n_1377;
wire n_2370;
wire n_989;
wire n_1039;
wire n_2214;
wire n_2055;
wire n_283;
wire n_1403;
wire n_2248;
wire n_2356;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_2062;
wire n_1002;
wire n_1463;
wire n_1581;
wire n_2100;
wire n_310;
wire n_593;
wire n_2258;
wire n_748;
wire n_586;
wire n_1058;
wire n_1667;
wire n_838;
wire n_332;
wire n_1053;
wire n_1224;
wire n_349;
wire n_1926;
wire n_1248;
wire n_1331;
wire n_953;
wire n_279;
wire n_1014;
wire n_1241;
wire n_2150;
wire n_2241;
wire n_2152;
wire n_289;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_440;
wire n_793;
wire n_478;
wire n_2140;
wire n_1819;
wire n_2330;
wire n_2139;
wire n_476;
wire n_1527;
wire n_2042;
wire n_534;
wire n_1882;
wire n_884;
wire n_345;
wire n_944;
wire n_1754;
wire n_1623;
wire n_2175;
wire n_2324;
wire n_1854;
wire n_1565;
wire n_1809;
wire n_1856;
wire n_647;
wire n_407;
wire n_1072;
wire n_2218;
wire n_2267;
wire n_832;
wire n_857;
wire n_2305;
wire n_561;
wire n_1319;
wire n_2379;
wire n_2154;
wire n_1825;
wire n_1951;
wire n_1883;
wire n_1906;
wire n_1712;
wire n_1387;
wire n_2262;
wire n_1532;
wire n_2322;
wire n_2271;
wire n_1027;
wire n_971;
wire n_1156;
wire n_326;
wire n_794;
wire n_404;
wire n_2331;
wire n_2293;
wire n_686;
wire n_847;
wire n_1393;
wire n_2319;
wire n_596;
wire n_1775;
wire n_2028;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_1709;
wire n_2108;
wire n_728;
wire n_266;
wire n_1162;
wire n_272;
wire n_1538;
wire n_1838;
wire n_1199;
wire n_1847;
wire n_1779;
wire n_352;
wire n_1884;
wire n_1038;
wire n_520;
wire n_1369;
wire n_409;
wire n_1841;
wire n_1660;
wire n_887;
wire n_1905;
wire n_2195;
wire n_300;
wire n_809;
wire n_931;
wire n_870;
wire n_599;
wire n_1711;
wire n_1662;
wire n_1891;
wire n_1481;
wire n_1942;
wire n_434;
wire n_1978;
wire n_1544;
wire n_868;
wire n_639;
wire n_914;
wire n_2120;
wire n_411;
wire n_414;
wire n_1629;
wire n_1293;
wire n_965;
wire n_1876;
wire n_1743;
wire n_935;
wire n_817;
wire n_1175;
wire n_360;
wire n_1479;
wire n_1810;
wire n_2350;
wire n_1888;
wire n_2009;
wire n_759;
wire n_2222;
wire n_1892;
wire n_806;
wire n_1997;
wire n_1766;
wire n_1477;
wire n_324;
wire n_1635;
wire n_1963;
wire n_2226;
wire n_1571;
wire n_1189;
wire n_2215;
wire n_1259;
wire n_1690;
wire n_706;
wire n_746;
wire n_1649;
wire n_747;
wire n_2064;
wire n_784;
wire n_1733;
wire n_1244;
wire n_431;
wire n_1194;
wire n_1925;
wire n_2297;
wire n_1815;
wire n_615;
wire n_851;
wire n_1759;
wire n_843;
wire n_1788;
wire n_2177;
wire n_523;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_2227;
wire n_678;
wire n_697;
wire n_1222;
wire n_1679;
wire n_2190;
wire n_776;
wire n_1798;
wire n_2022;
wire n_1790;
wire n_1415;
wire n_367;
wire n_452;
wire n_525;
wire n_1260;
wire n_1746;
wire n_1647;
wire n_2181;
wire n_1829;
wire n_1464;
wire n_649;
wire n_547;
wire n_1444;
wire n_1191;
wire n_1674;
wire n_1833;
wire n_1830;
wire n_2073;
wire n_1710;
wire n_284;
wire n_1128;
wire n_1734;
wire n_744;
wire n_629;
wire n_590;
wire n_1308;
wire n_2178;
wire n_1767;
wire n_2336;
wire n_254;
wire n_1680;
wire n_1233;
wire n_1615;
wire n_1529;
wire n_2005;
wire n_526;
wire n_1916;
wire n_372;
wire n_293;
wire n_677;
wire n_244;
wire n_1333;
wire n_1121;
wire n_433;
wire n_314;
wire n_368;
wire n_604;
wire n_2007;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_1001;
wire n_1503;
wire n_2054;
wire n_498;
wire n_1468;
wire n_1559;
wire n_1765;
wire n_1866;
wire n_689;
wire n_738;
wire n_1624;
wire n_640;
wire n_1510;
wire n_252;
wire n_624;
wire n_1380;
wire n_1744;
wire n_1617;
wire n_295;
wire n_1010;
wire n_1994;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_1195;
wire n_1839;
wire n_1837;
wire n_610;
wire n_1760;
wire n_936;
wire n_568;
wire n_1500;
wire n_1090;
wire n_757;
wire n_2342;
wire n_633;
wire n_439;
wire n_1832;
wire n_259;
wire n_448;
wire n_1851;
wire n_758;
wire n_999;
wire n_2046;
wire n_1933;
wire n_2290;
wire n_1656;
wire n_1158;
wire n_2045;
wire n_1509;
wire n_1874;
wire n_2040;
wire n_563;
wire n_2060;
wire n_1987;
wire n_1145;
wire n_878;
wire n_524;
wire n_394;
wire n_1678;
wire n_1049;
wire n_1153;
wire n_2145;
wire n_741;
wire n_1639;
wire n_1306;
wire n_1068;
wire n_1871;
wire n_1964;
wire n_331;
wire n_906;
wire n_1163;
wire n_2039;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_1781;
wire n_2084;
wire n_2035;
wire n_658;
wire n_2061;
wire n_2378;
wire n_1740;
wire n_1362;
wire n_1586;
wire n_456;
wire n_959;
wire n_535;
wire n_940;
wire n_1445;
wire n_1492;
wire n_2155;
wire n_1923;
wire n_1773;
wire n_592;
wire n_1169;
wire n_1596;
wire n_1692;
wire n_1017;
wire n_2171;
wire n_978;
wire n_2116;
wire n_2314;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_1095;
wire n_1828;
wire n_1614;
wire n_267;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_2093;
wire n_2038;
wire n_2320;
wire n_2339;
wire n_2137;
wire n_603;
wire n_1431;
wire n_484;
wire n_1593;
wire n_1033;
wire n_442;
wire n_2299;
wire n_636;
wire n_660;
wire n_2087;
wire n_1640;
wire n_2162;
wire n_1732;
wire n_1009;
wire n_1148;
wire n_2051;
wire n_742;
wire n_750;
wire n_2029;
wire n_995;
wire n_454;
wire n_2168;
wire n_1609;
wire n_374;
wire n_1989;
wire n_2359;
wire n_396;
wire n_1887;
wire n_1383;
wire n_1073;
wire n_255;
wire n_2346;
wire n_662;
wire n_459;
wire n_2312;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1920;
wire n_1065;
wire n_1592;
wire n_1336;
wire n_1721;
wire n_1959;
wire n_1758;
wire n_2338;
wire n_1574;
wire n_473;
wire n_2048;
wire n_2355;
wire n_2133;
wire n_1921;
wire n_1309;
wire n_1878;
wire n_1426;
wire n_1043;
wire n_355;
wire n_486;
wire n_1800;
wire n_1548;
wire n_614;
wire n_337;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_2124;
wire n_743;
wire n_2081;
wire n_299;
wire n_303;
wire n_296;
wire n_613;
wire n_1119;
wire n_2156;
wire n_1240;
wire n_2261;
wire n_1820;
wire n_829;
wire n_1612;
wire n_2179;
wire n_1416;
wire n_2077;
wire n_1724;
wire n_2111;
wire n_361;
wire n_700;
wire n_1237;
wire n_573;
wire n_1420;
wire n_1132;
wire n_388;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_2277;
wire n_761;
wire n_1785;
wire n_1568;
wire n_1006;
wire n_2110;
wire n_329;
wire n_274;
wire n_1270;
wire n_1664;
wire n_1486;
wire n_582;
wire n_1332;
wire n_2231;
wire n_1390;
wire n_2017;
wire n_2090;
wire n_1870;
wire n_309;
wire n_512;
wire n_2367;
wire n_1591;
wire n_2033;
wire n_322;
wire n_1682;
wire n_1980;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1927;
wire n_2132;
wire n_1349;
wire n_1093;
wire n_288;
wire n_1031;
wire n_263;
wire n_609;
wire n_1041;
wire n_1265;
wire n_1909;
wire n_1562;
wire n_383;
wire n_834;
wire n_765;
wire n_2255;
wire n_2272;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_1965;
wire n_239;
wire n_630;
wire n_1902;
wire n_2151;
wire n_1941;
wire n_2106;
wire n_1913;
wire n_504;
wire n_1823;
wire n_511;
wire n_874;
wire n_358;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_2230;
wire n_2015;
wire n_2365;
wire n_1875;
wire n_1982;
wire n_1304;
wire n_1324;
wire n_987;
wire n_1846;
wire n_261;
wire n_2066;
wire n_1885;
wire n_1455;
wire n_767;
wire n_993;
wire n_1903;
wire n_1407;
wire n_1551;
wire n_545;
wire n_860;
wire n_441;
wire n_450;
wire n_1805;
wire n_2176;
wire n_2204;
wire n_1816;
wire n_429;
wire n_948;
wire n_1217;
wire n_2220;
wire n_628;
wire n_365;
wire n_1849;
wire n_729;
wire n_1131;
wire n_1084;
wire n_1961;
wire n_970;
wire n_1935;
wire n_911;
wire n_1430;
wire n_513;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1534;
wire n_340;
wire n_2288;
wire n_1351;
wire n_2240;
wire n_1044;
wire n_1205;
wire n_346;
wire n_1209;
wire n_1552;
wire n_495;
wire n_602;
wire n_574;
wire n_1435;
wire n_879;
wire n_623;
wire n_2088;
wire n_405;
wire n_824;
wire n_359;
wire n_1645;
wire n_490;
wire n_1327;
wire n_2243;
wire n_996;
wire n_921;
wire n_1684;
wire n_1717;
wire n_572;
wire n_366;
wire n_815;
wire n_1795;
wire n_2128;
wire n_1821;
wire n_327;
wire n_1381;
wire n_1611;
wire n_1037;
wire n_2368;
wire n_1080;
wire n_2301;
wire n_1274;
wire n_1316;
wire n_1708;
wire n_426;
wire n_1438;
wire n_1082;
wire n_1840;
wire n_589;
wire n_716;
wire n_1630;
wire n_2122;
wire n_562;
wire n_1436;
wire n_1691;
wire n_952;
wire n_2092;
wire n_1229;
wire n_391;
wire n_701;
wire n_1437;
wire n_1023;
wire n_2075;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_238;
wire n_1776;
wire n_2198;
wire n_2281;
wire n_2131;
wire n_2216;
wire n_531;
wire n_1757;
wire n_890;
wire n_1897;
wire n_764;
wire n_1919;
wire n_1056;
wire n_1424;
wire n_960;
wire n_2308;
wire n_1893;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_2053;
wire n_2163;
wire n_634;
wire n_2328;
wire n_1958;
wire n_2254;
wire n_1252;
wire n_348;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_1311;
wire n_2191;
wire n_1519;
wire n_256;
wire n_950;
wire n_1553;
wire n_1811;
wire n_380;
wire n_419;
wire n_1346;
wire n_444;
wire n_1299;
wire n_2158;
wire n_1808;
wire n_1060;
wire n_1141;
wire n_316;
wire n_2266;
wire n_389;
wire n_418;
wire n_248;
wire n_912;
wire n_968;
wire n_315;
wire n_451;
wire n_619;
wire n_408;
wire n_1386;
wire n_1699;
wire n_376;
wire n_967;
wire n_1442;
wire n_1139;
wire n_515;
wire n_2333;
wire n_351;
wire n_885;
wire n_397;
wire n_1432;
wire n_1357;
wire n_483;
wire n_2125;
wire n_683;
wire n_1632;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_1954;
wire n_2265;
wire n_1608;
wire n_983;
wire n_1844;
wire n_280;
wire n_1305;
wire n_873;
wire n_1826;
wire n_378;
wire n_1112;
wire n_2304;
wire n_762;
wire n_1283;
wire n_1644;
wire n_2334;
wire n_690;
wire n_1974;
wire n_583;
wire n_2086;
wire n_2289;
wire n_302;
wire n_1343;
wire n_2263;
wire n_1203;
wire n_1631;
wire n_821;
wire n_1763;
wire n_2341;
wire n_1966;
wire n_1768;
wire n_321;
wire n_2294;
wire n_1179;
wire n_621;
wire n_753;
wire n_455;
wire n_1048;
wire n_1719;
wire n_1288;
wire n_385;
wire n_507;
wire n_2269;
wire n_2309;
wire n_1560;
wire n_1605;
wire n_2236;
wire n_330;
wire n_1228;
wire n_2123;
wire n_972;
wire n_692;
wire n_2037;
wire n_1953;
wire n_1938;
wire n_820;
wire n_1200;
wire n_1911;
wire n_1363;
wire n_1301;
wire n_1668;
wire n_1185;
wire n_991;
wire n_828;
wire n_1967;
wire n_779;
wire n_576;
wire n_1143;
wire n_1579;
wire n_2233;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_537;
wire n_1688;
wire n_945;
wire n_492;
wire n_1504;
wire n_943;
wire n_341;
wire n_250;
wire n_992;
wire n_1932;
wire n_543;
wire n_260;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_2082;
wire n_286;
wire n_1992;
wire n_1643;
wire n_883;
wire n_1983;
wire n_470;
wire n_449;
wire n_325;
wire n_1594;
wire n_1214;
wire n_1342;
wire n_1400;
wire n_900;
wire n_2362;
wire n_856;
wire n_1793;
wire n_1976;
wire n_2223;
wire n_918;
wire n_942;
wire n_2169;
wire n_1804;
wire n_1147;
wire n_1557;
wire n_1977;
wire n_2153;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_2364;
wire n_540;
wire n_618;
wire n_896;
wire n_2310;
wire n_323;
wire n_2287;
wire n_356;
wire n_2291;
wire n_894;
wire n_1636;
wire n_2056;
wire n_1730;
wire n_831;
wire n_2280;
wire n_2192;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1865;
wire n_1470;
wire n_1096;
wire n_2094;
wire n_1575;
wire n_1697;
wire n_1735;
wire n_833;
wire n_2318;
wire n_2020;
wire n_1646;
wire n_1307;
wire n_1881;
wire n_988;
wire n_2043;
wire n_1940;
wire n_814;
wire n_1549;
wire n_1934;
wire n_2311;
wire n_1201;
wire n_1114;
wire n_655;
wire n_2025;
wire n_1616;
wire n_1446;
wire n_2285;
wire n_669;
wire n_472;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_2298;
wire n_1807;
wire n_387;
wire n_1149;
wire n_398;
wire n_1671;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_2303;
wire n_1824;
wire n_1917;
wire n_2295;
wire n_1219;
wire n_1204;
wire n_2325;
wire n_1814;
wire n_1035;
wire n_287;
wire n_555;
wire n_783;
wire n_1848;
wire n_1928;
wire n_2126;
wire n_1188;
wire n_1722;
wire n_661;
wire n_1802;
wire n_849;
wire n_336;
wire n_681;
wire n_584;
wire n_1638;
wire n_1786;
wire n_430;
wire n_2002;
wire n_2282;
wire n_510;
wire n_2371;
wire n_311;
wire n_830;
wire n_2098;
wire n_1296;
wire n_2352;
wire n_1413;
wire n_801;
wire n_2207;
wire n_2080;
wire n_2377;
wire n_2340;
wire n_2068;
wire n_241;
wire n_875;
wire n_357;
wire n_1110;
wire n_1655;
wire n_445;
wire n_749;
wire n_1895;
wire n_1134;
wire n_1358;
wire n_717;
wire n_939;
wire n_482;
wire n_2361;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_249;
wire n_1998;
wire n_304;
wire n_1338;
wire n_577;
wire n_2016;
wire n_1522;
wire n_1687;
wire n_1637;
wire n_2034;
wire n_1419;
wire n_338;
wire n_1653;
wire n_693;
wire n_2270;
wire n_1506;
wire n_836;
wire n_990;
wire n_1886;
wire n_1389;
wire n_1894;
wire n_975;
wire n_1908;
wire n_1256;
wire n_1702;
wire n_2259;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_306;
wire n_770;
wire n_458;
wire n_1375;
wire n_1102;
wire n_1843;
wire n_711;
wire n_1499;
wire n_1187;
wire n_1441;
wire n_1392;
wire n_1597;
wire n_1929;
wire n_1164;
wire n_1659;
wire n_1834;
wire n_2097;
wire n_2313;
wire n_489;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_2206;
wire n_2063;
wire n_1572;
wire n_1968;
wire n_2252;
wire n_876;
wire n_1516;
wire n_1190;
wire n_1736;
wire n_1685;
wire n_601;
wire n_917;
wire n_1714;
wire n_966;
wire n_253;
wire n_1116;
wire n_2000;
wire n_1661;
wire n_1212;
wire n_2074;
wire n_1541;
wire n_726;
wire n_982;
wire n_1573;
wire n_1453;
wire n_1731;
wire n_2217;
wire n_818;
wire n_2373;
wire n_1970;
wire n_861;
wire n_1713;
wire n_1183;
wire n_2307;
wire n_1658;
wire n_899;
wire n_1253;
wire n_1737;
wire n_2201;
wire n_2117;
wire n_1904;
wire n_1993;
wire n_774;
wire n_1628;
wire n_2205;
wire n_1335;
wire n_1514;
wire n_1777;
wire n_1957;
wire n_1059;
wire n_1345;
wire n_1133;
wire n_1771;
wire n_1912;
wire n_1899;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_2067;
wire n_527;
wire n_707;
wire n_1168;
wire n_2219;
wire n_2148;
wire n_937;
wire n_1427;
wire n_393;
wire n_487;
wire n_1726;
wire n_665;
wire n_1584;
wire n_1835;
wire n_1440;
wire n_2164;
wire n_421;
wire n_1988;
wire n_2115;
wire n_1853;
wire n_1356;
wire n_1787;
wire n_910;
wire n_2232;
wire n_2212;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1302;
wire n_1774;
wire n_1725;
wire n_1136;
wire n_1313;
wire n_1491;
wire n_754;
wire n_1496;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_1812;
wire n_735;
wire n_1915;
wire n_1109;
wire n_895;
wire n_1310;
wire n_2121;
wire n_1803;
wire n_427;
wire n_1399;
wire n_1543;
wire n_1991;
wire n_1979;
wire n_791;
wire n_732;
wire n_1533;
wire n_2224;
wire n_808;
wire n_797;
wire n_1025;
wire n_1930;
wire n_1955;
wire n_500;
wire n_1067;
wire n_1720;
wire n_435;
wire n_2003;
wire n_766;
wire n_1457;
wire n_541;
wire n_538;
wire n_2354;
wire n_2246;
wire n_2008;
wire n_1117;
wire n_799;
wire n_2264;
wire n_687;
wire n_715;
wire n_1742;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_2012;
wire n_594;
wire n_1291;
wire n_1297;
wire n_1753;
wire n_2283;
wire n_1782;
wire n_2245;
wire n_1155;
wire n_1418;
wire n_1972;
wire n_1524;
wire n_1689;
wire n_1485;
wire n_1011;
wire n_1184;
wire n_2184;
wire n_985;
wire n_1855;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_1703;
wire n_1352;
wire n_626;
wire n_2197;
wire n_2199;
wire n_1650;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_1170;
wire n_305;
wire n_2023;
wire n_2213;
wire n_2351;
wire n_2211;
wire n_2095;
wire n_676;
wire n_294;
wire n_318;
wire n_2103;
wire n_653;
wire n_2160;
wire n_642;
wire n_2228;
wire n_1602;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_268;
wire n_2286;
wire n_664;
wire n_1999;
wire n_503;
wire n_2372;
wire n_2065;
wire n_2136;
wire n_1372;
wire n_605;
wire n_1273;
wire n_1822;
wire n_353;
wire n_620;
wire n_643;
wire n_2363;
wire n_916;
wire n_1081;
wire n_493;
wire n_2332;
wire n_1235;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_1282;
wire n_1318;
wire n_1783;
wire n_780;
wire n_998;
wire n_2375;
wire n_1454;
wire n_467;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_1907;
wire n_501;
wire n_823;
wire n_245;
wire n_725;
wire n_2344;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_2316;
wire n_672;
wire n_1985;
wire n_1898;
wire n_2107;
wire n_581;
wire n_382;
wire n_554;
wire n_1625;
wire n_2130;
wire n_2187;
wire n_2284;
wire n_898;
wire n_1762;
wire n_1013;
wire n_1452;
wire n_718;
wire n_265;
wire n_1120;
wire n_719;
wire n_443;
wire n_1791;
wire n_1890;
wire n_1747;
wire n_714;
wire n_1683;
wire n_1817;
wire n_909;
wire n_1944;
wire n_1497;
wire n_1530;
wire n_997;
wire n_932;
wire n_612;
wire n_2078;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_1981;
wire n_508;
wire n_2186;
wire n_506;
wire n_1320;
wire n_1663;
wire n_737;
wire n_1718;
wire n_986;
wire n_2315;
wire n_509;
wire n_1317;
wire n_1518;
wire n_1715;
wire n_2102;
wire n_1281;
wire n_1952;
wire n_1192;
wire n_2221;
wire n_1024;
wire n_1063;
wire n_1889;
wire n_1792;
wire n_1564;
wire n_1868;
wire n_1613;
wire n_733;
wire n_1489;
wire n_1922;
wire n_1376;
wire n_941;
wire n_2326;
wire n_981;
wire n_1569;
wire n_2188;
wire n_867;
wire n_2348;
wire n_2239;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_298;
wire n_2104;
wire n_518;
wire n_505;
wire n_2057;
wire n_1772;
wire n_282;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1861;
wire n_2129;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1901;
wire n_1900;
wire n_1620;
wire n_381;
wire n_390;
wire n_1330;
wire n_1867;
wire n_1945;
wire n_481;
wire n_1675;
wire n_1924;
wire n_1727;
wire n_1554;
wire n_1745;
wire n_769;
wire n_2006;
wire n_1995;
wire n_2138;
wire n_1046;
wire n_271;
wire n_934;
wire n_1618;
wire n_2260;
wire n_826;
wire n_2343;
wire n_1813;
wire n_886;
wire n_2014;
wire n_1221;
wire n_2345;
wire n_654;
wire n_1172;
wire n_428;
wire n_379;
wire n_1341;
wire n_570;
wire n_1641;
wire n_1361;
wire n_1707;
wire n_853;
wire n_377;
wire n_2317;
wire n_751;
wire n_2172;
wire n_1973;
wire n_786;
wire n_1083;
wire n_1142;
wire n_2376;
wire n_1129;
wire n_392;
wire n_704;
wire n_787;
wire n_1770;
wire n_961;
wire n_2250;
wire n_1756;
wire n_771;
wire n_276;
wire n_1716;
wire n_1225;
wire n_1520;
wire n_522;
wire n_1287;
wire n_1262;
wire n_400;
wire n_930;
wire n_1873;
wire n_1411;
wire n_622;
wire n_1962;
wire n_1577;
wire n_1087;
wire n_386;
wire n_994;
wire n_1701;
wire n_2194;
wire n_848;
wire n_1550;
wire n_1498;
wire n_2167;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1567;
wire n_1247;
wire n_922;
wire n_816;
wire n_1648;
wire n_591;
wire n_1536;
wire n_1857;
wire n_1344;
wire n_2041;
wire n_313;
wire n_631;
wire n_479;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_1797;
wire n_432;
wire n_1769;
wire n_839;
wire n_1210;
wire n_1364;
wire n_2357;
wire n_2183;
wire n_2360;
wire n_328;
wire n_2292;
wire n_1250;
wire n_2173;
wire n_369;
wire n_1842;
wire n_871;
wire n_685;
wire n_598;
wire n_608;
wire n_928;
wire n_1367;
wire n_1943;
wire n_1460;
wire n_772;
wire n_2018;
wire n_1555;
wire n_499;
wire n_1589;
wire n_517;
wire n_402;
wire n_413;
wire n_1086;
wire n_796;
wire n_1858;
wire n_1619;
wire n_2119;
wire n_1502;
wire n_2157;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_2030;
wire n_903;
wire n_1525;
wire n_1752;
wire n_740;
wire n_384;
wire n_2208;
wire n_1404;
wire n_1794;
wire n_2182;
wire n_1315;
wire n_2234;
wire n_277;
wire n_1061;
wire n_1910;
wire n_333;
wire n_1298;
wire n_1652;
wire n_2209;
wire n_462;
wire n_2050;
wire n_1193;
wire n_1676;
wire n_1255;
wire n_258;
wire n_1113;
wire n_2321;
wire n_1226;
wire n_722;
wire n_1277;
wire n_2146;
wire n_844;
wire n_471;
wire n_852;
wire n_1487;
wire n_1864;
wire n_1028;
wire n_1601;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_1546;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_1627;
wire n_1245;
wire n_846;
wire n_1673;
wire n_465;
wire n_1321;
wire n_362;
wire n_1975;
wire n_2296;
wire n_2070;
wire n_273;
wire n_1937;
wire n_585;
wire n_2112;
wire n_1739;
wire n_270;
wire n_616;
wire n_2278;
wire n_1914;
wire n_2135;
wire n_2335;
wire n_745;
wire n_1654;
wire n_2349;
wire n_1103;
wire n_648;
wire n_1379;
wire n_312;
wire n_2196;
wire n_2170;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_494;
wire n_1761;
wire n_641;
wire n_730;
wire n_2036;
wire n_1325;
wire n_1595;
wire n_2161;
wire n_354;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_2083;
wire n_695;
wire n_656;
wire n_1606;
wire n_1220;
wire n_1694;
wire n_1540;
wire n_1936;
wire n_1956;
wire n_437;
wire n_1642;
wire n_2279;
wire n_2027;
wire n_403;
wire n_453;
wire n_1130;
wire n_720;
wire n_2366;
wire n_1918;
wire n_1526;
wire n_863;
wire n_2210;
wire n_805;
wire n_1604;
wire n_1275;
wire n_1764;
wire n_712;
wire n_246;
wire n_1583;
wire n_1042;
wire n_1402;
wire n_269;
wire n_2049;
wire n_2273;
wire n_285;
wire n_412;
wire n_1493;
wire n_657;
wire n_644;
wire n_1741;
wire n_2229;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_2004;
wire n_1621;
wire n_2113;
wire n_251;
wire n_566;
wire n_565;
wire n_1448;
wire n_2225;
wire n_1507;
wire n_1398;
wire n_1879;
wire n_597;
wire n_1996;
wire n_1181;
wire n_1505;
wire n_1634;
wire n_1196;
wire n_2019;
wire n_651;
wire n_1340;
wire n_2274;
wire n_334;
wire n_811;
wire n_1558;
wire n_807;
wire n_2166;
wire n_835;
wire n_666;
wire n_262;
wire n_1433;
wire n_1704;
wire n_2256;
wire n_1254;
wire n_1026;
wire n_2026;
wire n_1969;
wire n_1234;
wire n_2109;
wire n_319;
wire n_364;
wire n_1138;
wire n_927;
wire n_1089;
wire n_2013;
wire n_1990;
wire n_2044;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_242;
wire n_1681;
wire n_2010;
wire n_1018;
wire n_2242;
wire n_2247;
wire n_1693;
wire n_438;
wire n_713;
wire n_904;
wire n_1588;
wire n_1622;
wire n_2237;
wire n_1180;
wire n_1827;
wire n_1271;
wire n_533;
wire n_1542;
wire n_1251;
wire n_278;
wire n_2268;

BUFx10_ASAP7_75t_L g238 ( 
.A(n_152),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_225),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_216),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_9),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_206),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_63),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_168),
.Y(n_244)
);

INVx1_ASAP7_75t_SL g245 ( 
.A(n_74),
.Y(n_245)
);

BUFx6f_ASAP7_75t_L g246 ( 
.A(n_31),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_229),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_176),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_19),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_17),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_150),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_43),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_14),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_196),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_66),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_156),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_209),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_203),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_89),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_113),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_39),
.Y(n_261)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_160),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_186),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_55),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_83),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_211),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_237),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_178),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_34),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_99),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_73),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_230),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_114),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_37),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_147),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_6),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_228),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_44),
.Y(n_278)
);

BUFx2_ASAP7_75t_SL g279 ( 
.A(n_67),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_70),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_173),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_195),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_1),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_183),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_32),
.Y(n_285)
);

CKINVDCx16_ASAP7_75t_R g286 ( 
.A(n_89),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_1),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_131),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_37),
.Y(n_289)
);

INVx1_ASAP7_75t_SL g290 ( 
.A(n_164),
.Y(n_290)
);

INVx1_ASAP7_75t_SL g291 ( 
.A(n_35),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_19),
.Y(n_292)
);

BUFx10_ASAP7_75t_L g293 ( 
.A(n_41),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_223),
.Y(n_294)
);

BUFx2_ASAP7_75t_L g295 ( 
.A(n_205),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_182),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g297 ( 
.A(n_97),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_214),
.Y(n_298)
);

BUFx6f_ASAP7_75t_L g299 ( 
.A(n_190),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_73),
.Y(n_300)
);

HB1xp67_ASAP7_75t_L g301 ( 
.A(n_204),
.Y(n_301)
);

INVx1_ASAP7_75t_SL g302 ( 
.A(n_79),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_148),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_47),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_149),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_38),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_187),
.Y(n_307)
);

BUFx10_ASAP7_75t_L g308 ( 
.A(n_227),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_226),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_107),
.Y(n_310)
);

BUFx2_ASAP7_75t_L g311 ( 
.A(n_232),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_191),
.Y(n_312)
);

INVx1_ASAP7_75t_SL g313 ( 
.A(n_133),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_224),
.Y(n_314)
);

HB1xp67_ASAP7_75t_L g315 ( 
.A(n_16),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_184),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_29),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_88),
.Y(n_318)
);

BUFx6f_ASAP7_75t_L g319 ( 
.A(n_33),
.Y(n_319)
);

INVx2_ASAP7_75t_L g320 ( 
.A(n_221),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_132),
.Y(n_321)
);

BUFx6f_ASAP7_75t_L g322 ( 
.A(n_91),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_82),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_188),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_81),
.Y(n_325)
);

INVx1_ASAP7_75t_SL g326 ( 
.A(n_20),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_14),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_87),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_122),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_24),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_134),
.Y(n_331)
);

CKINVDCx14_ASAP7_75t_R g332 ( 
.A(n_42),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_180),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_236),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_201),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_151),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_138),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_2),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_213),
.Y(n_339)
);

INVx2_ASAP7_75t_L g340 ( 
.A(n_219),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_175),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_39),
.Y(n_342)
);

BUFx6f_ASAP7_75t_L g343 ( 
.A(n_169),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_95),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_146),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_167),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_193),
.Y(n_347)
);

BUFx10_ASAP7_75t_L g348 ( 
.A(n_217),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_7),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_51),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_2),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_31),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_171),
.Y(n_353)
);

CKINVDCx20_ASAP7_75t_R g354 ( 
.A(n_30),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_102),
.Y(n_355)
);

INVx2_ASAP7_75t_L g356 ( 
.A(n_192),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_9),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_16),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_10),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_76),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_210),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_82),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_13),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_76),
.Y(n_364)
);

CKINVDCx16_ASAP7_75t_R g365 ( 
.A(n_108),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_212),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_105),
.Y(n_367)
);

INVx1_ASAP7_75t_SL g368 ( 
.A(n_11),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_218),
.Y(n_369)
);

CKINVDCx20_ASAP7_75t_R g370 ( 
.A(n_75),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_45),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_128),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_94),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_70),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_233),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_29),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_92),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_75),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_49),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_104),
.Y(n_380)
);

INVx2_ASAP7_75t_L g381 ( 
.A(n_142),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_10),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_159),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_126),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_21),
.Y(n_385)
);

CKINVDCx20_ASAP7_75t_R g386 ( 
.A(n_4),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_155),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_46),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_60),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_17),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_22),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_177),
.Y(n_392)
);

BUFx3_ASAP7_75t_L g393 ( 
.A(n_189),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_61),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_90),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_124),
.Y(n_396)
);

CKINVDCx20_ASAP7_75t_R g397 ( 
.A(n_137),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_52),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_57),
.Y(n_399)
);

BUFx3_ASAP7_75t_L g400 ( 
.A(n_207),
.Y(n_400)
);

CKINVDCx20_ASAP7_75t_R g401 ( 
.A(n_83),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_56),
.Y(n_402)
);

INVx1_ASAP7_75t_SL g403 ( 
.A(n_81),
.Y(n_403)
);

INVx2_ASAP7_75t_L g404 ( 
.A(n_43),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_3),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_121),
.Y(n_406)
);

CKINVDCx20_ASAP7_75t_R g407 ( 
.A(n_145),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_127),
.Y(n_408)
);

BUFx6f_ASAP7_75t_L g409 ( 
.A(n_78),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_49),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_88),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_129),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_110),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_40),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_79),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_22),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_60),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_179),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_64),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_24),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_91),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_0),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_112),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_111),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_116),
.Y(n_425)
);

CKINVDCx16_ASAP7_75t_R g426 ( 
.A(n_38),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_4),
.Y(n_427)
);

BUFx5_ASAP7_75t_L g428 ( 
.A(n_119),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_118),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_25),
.Y(n_430)
);

INVx2_ASAP7_75t_SL g431 ( 
.A(n_8),
.Y(n_431)
);

CKINVDCx5p33_ASAP7_75t_R g432 ( 
.A(n_67),
.Y(n_432)
);

BUFx3_ASAP7_75t_L g433 ( 
.A(n_66),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_20),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_40),
.Y(n_435)
);

CKINVDCx5p33_ASAP7_75t_R g436 ( 
.A(n_135),
.Y(n_436)
);

INVx2_ASAP7_75t_L g437 ( 
.A(n_50),
.Y(n_437)
);

BUFx3_ASAP7_75t_L g438 ( 
.A(n_21),
.Y(n_438)
);

BUFx10_ASAP7_75t_L g439 ( 
.A(n_68),
.Y(n_439)
);

CKINVDCx5p33_ASAP7_75t_R g440 ( 
.A(n_65),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_35),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_143),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_54),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_208),
.Y(n_444)
);

CKINVDCx5p33_ASAP7_75t_R g445 ( 
.A(n_144),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_235),
.Y(n_446)
);

CKINVDCx20_ASAP7_75t_R g447 ( 
.A(n_72),
.Y(n_447)
);

CKINVDCx20_ASAP7_75t_R g448 ( 
.A(n_69),
.Y(n_448)
);

BUFx3_ASAP7_75t_L g449 ( 
.A(n_158),
.Y(n_449)
);

CKINVDCx5p33_ASAP7_75t_R g450 ( 
.A(n_92),
.Y(n_450)
);

CKINVDCx5p33_ASAP7_75t_R g451 ( 
.A(n_7),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_117),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_231),
.Y(n_453)
);

CKINVDCx5p33_ASAP7_75t_R g454 ( 
.A(n_45),
.Y(n_454)
);

CKINVDCx5p33_ASAP7_75t_R g455 ( 
.A(n_93),
.Y(n_455)
);

CKINVDCx5p33_ASAP7_75t_R g456 ( 
.A(n_13),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_220),
.Y(n_457)
);

CKINVDCx5p33_ASAP7_75t_R g458 ( 
.A(n_15),
.Y(n_458)
);

CKINVDCx5p33_ASAP7_75t_R g459 ( 
.A(n_85),
.Y(n_459)
);

BUFx6f_ASAP7_75t_L g460 ( 
.A(n_5),
.Y(n_460)
);

INVx2_ASAP7_75t_L g461 ( 
.A(n_90),
.Y(n_461)
);

CKINVDCx5p33_ASAP7_75t_R g462 ( 
.A(n_200),
.Y(n_462)
);

CKINVDCx5p33_ASAP7_75t_R g463 ( 
.A(n_64),
.Y(n_463)
);

CKINVDCx5p33_ASAP7_75t_R g464 ( 
.A(n_62),
.Y(n_464)
);

CKINVDCx5p33_ASAP7_75t_R g465 ( 
.A(n_234),
.Y(n_465)
);

CKINVDCx5p33_ASAP7_75t_R g466 ( 
.A(n_239),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_246),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_246),
.Y(n_468)
);

CKINVDCx5p33_ASAP7_75t_R g469 ( 
.A(n_242),
.Y(n_469)
);

CKINVDCx5p33_ASAP7_75t_R g470 ( 
.A(n_244),
.Y(n_470)
);

CKINVDCx20_ASAP7_75t_R g471 ( 
.A(n_254),
.Y(n_471)
);

HB1xp67_ASAP7_75t_L g472 ( 
.A(n_286),
.Y(n_472)
);

NOR2xp33_ASAP7_75t_L g473 ( 
.A(n_295),
.B(n_0),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_246),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_246),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_246),
.Y(n_476)
);

CKINVDCx5p33_ASAP7_75t_R g477 ( 
.A(n_247),
.Y(n_477)
);

INVxp67_ASAP7_75t_L g478 ( 
.A(n_315),
.Y(n_478)
);

CKINVDCx5p33_ASAP7_75t_R g479 ( 
.A(n_248),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_319),
.Y(n_480)
);

CKINVDCx20_ASAP7_75t_R g481 ( 
.A(n_297),
.Y(n_481)
);

CKINVDCx16_ASAP7_75t_R g482 ( 
.A(n_426),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_319),
.Y(n_483)
);

BUFx2_ASAP7_75t_L g484 ( 
.A(n_433),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_319),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_319),
.Y(n_486)
);

CKINVDCx20_ASAP7_75t_R g487 ( 
.A(n_397),
.Y(n_487)
);

HB1xp67_ASAP7_75t_L g488 ( 
.A(n_286),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_319),
.Y(n_489)
);

INVxp33_ASAP7_75t_SL g490 ( 
.A(n_241),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_322),
.Y(n_491)
);

CKINVDCx20_ASAP7_75t_R g492 ( 
.A(n_407),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_322),
.Y(n_493)
);

INVxp33_ASAP7_75t_SL g494 ( 
.A(n_243),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_322),
.Y(n_495)
);

CKINVDCx5p33_ASAP7_75t_R g496 ( 
.A(n_251),
.Y(n_496)
);

INVxp33_ASAP7_75t_L g497 ( 
.A(n_249),
.Y(n_497)
);

NOR2xp67_ASAP7_75t_L g498 ( 
.A(n_431),
.B(n_3),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_322),
.Y(n_499)
);

CKINVDCx5p33_ASAP7_75t_R g500 ( 
.A(n_256),
.Y(n_500)
);

CKINVDCx5p33_ASAP7_75t_R g501 ( 
.A(n_257),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_322),
.Y(n_502)
);

CKINVDCx5p33_ASAP7_75t_R g503 ( 
.A(n_258),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_409),
.Y(n_504)
);

CKINVDCx16_ASAP7_75t_R g505 ( 
.A(n_365),
.Y(n_505)
);

NOR2xp33_ASAP7_75t_L g506 ( 
.A(n_295),
.B(n_5),
.Y(n_506)
);

CKINVDCx16_ASAP7_75t_R g507 ( 
.A(n_332),
.Y(n_507)
);

INVxp33_ASAP7_75t_L g508 ( 
.A(n_249),
.Y(n_508)
);

CKINVDCx20_ASAP7_75t_R g509 ( 
.A(n_260),
.Y(n_509)
);

CKINVDCx5p33_ASAP7_75t_R g510 ( 
.A(n_266),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_240),
.Y(n_511)
);

CKINVDCx5p33_ASAP7_75t_R g512 ( 
.A(n_267),
.Y(n_512)
);

CKINVDCx5p33_ASAP7_75t_R g513 ( 
.A(n_268),
.Y(n_513)
);

HB1xp67_ASAP7_75t_L g514 ( 
.A(n_250),
.Y(n_514)
);

CKINVDCx5p33_ASAP7_75t_R g515 ( 
.A(n_272),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_409),
.Y(n_516)
);

INVxp67_ASAP7_75t_SL g517 ( 
.A(n_301),
.Y(n_517)
);

BUFx6f_ASAP7_75t_L g518 ( 
.A(n_299),
.Y(n_518)
);

CKINVDCx5p33_ASAP7_75t_R g519 ( 
.A(n_277),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_409),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_L g521 ( 
.A(n_311),
.B(n_6),
.Y(n_521)
);

CKINVDCx5p33_ASAP7_75t_R g522 ( 
.A(n_281),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_409),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_409),
.Y(n_524)
);

CKINVDCx5p33_ASAP7_75t_R g525 ( 
.A(n_282),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_460),
.Y(n_526)
);

CKINVDCx5p33_ASAP7_75t_R g527 ( 
.A(n_288),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_460),
.Y(n_528)
);

INVxp67_ASAP7_75t_SL g529 ( 
.A(n_311),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_460),
.Y(n_530)
);

CKINVDCx5p33_ASAP7_75t_R g531 ( 
.A(n_296),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_460),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_240),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_460),
.Y(n_534)
);

INVxp67_ASAP7_75t_SL g535 ( 
.A(n_393),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_404),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_404),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_437),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_437),
.Y(n_539)
);

CKINVDCx20_ASAP7_75t_R g540 ( 
.A(n_303),
.Y(n_540)
);

HB1xp67_ASAP7_75t_L g541 ( 
.A(n_255),
.Y(n_541)
);

CKINVDCx20_ASAP7_75t_R g542 ( 
.A(n_309),
.Y(n_542)
);

CKINVDCx20_ASAP7_75t_R g543 ( 
.A(n_312),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_461),
.Y(n_544)
);

INVxp67_ASAP7_75t_L g545 ( 
.A(n_279),
.Y(n_545)
);

NOR2xp33_ASAP7_75t_L g546 ( 
.A(n_263),
.B(n_8),
.Y(n_546)
);

CKINVDCx5p33_ASAP7_75t_R g547 ( 
.A(n_314),
.Y(n_547)
);

HB1xp67_ASAP7_75t_L g548 ( 
.A(n_261),
.Y(n_548)
);

NOR2xp67_ASAP7_75t_L g549 ( 
.A(n_431),
.B(n_11),
.Y(n_549)
);

CKINVDCx20_ASAP7_75t_R g550 ( 
.A(n_321),
.Y(n_550)
);

CKINVDCx20_ASAP7_75t_R g551 ( 
.A(n_329),
.Y(n_551)
);

CKINVDCx20_ASAP7_75t_R g552 ( 
.A(n_331),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_461),
.Y(n_553)
);

INVxp67_ASAP7_75t_L g554 ( 
.A(n_279),
.Y(n_554)
);

CKINVDCx20_ASAP7_75t_R g555 ( 
.A(n_333),
.Y(n_555)
);

CKINVDCx16_ASAP7_75t_R g556 ( 
.A(n_293),
.Y(n_556)
);

CKINVDCx5p33_ASAP7_75t_R g557 ( 
.A(n_334),
.Y(n_557)
);

CKINVDCx20_ASAP7_75t_R g558 ( 
.A(n_335),
.Y(n_558)
);

INVx2_ASAP7_75t_L g559 ( 
.A(n_428),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_252),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_252),
.Y(n_561)
);

HB1xp67_ASAP7_75t_L g562 ( 
.A(n_264),
.Y(n_562)
);

CKINVDCx20_ASAP7_75t_R g563 ( 
.A(n_336),
.Y(n_563)
);

BUFx2_ASAP7_75t_L g564 ( 
.A(n_433),
.Y(n_564)
);

CKINVDCx5p33_ASAP7_75t_R g565 ( 
.A(n_337),
.Y(n_565)
);

CKINVDCx5p33_ASAP7_75t_R g566 ( 
.A(n_339),
.Y(n_566)
);

CKINVDCx20_ASAP7_75t_R g567 ( 
.A(n_341),
.Y(n_567)
);

INVxp33_ASAP7_75t_SL g568 ( 
.A(n_265),
.Y(n_568)
);

CKINVDCx5p33_ASAP7_75t_R g569 ( 
.A(n_344),
.Y(n_569)
);

CKINVDCx5p33_ASAP7_75t_R g570 ( 
.A(n_345),
.Y(n_570)
);

CKINVDCx20_ASAP7_75t_R g571 ( 
.A(n_346),
.Y(n_571)
);

CKINVDCx16_ASAP7_75t_R g572 ( 
.A(n_293),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_253),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_253),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_259),
.Y(n_575)
);

INVx2_ASAP7_75t_L g576 ( 
.A(n_428),
.Y(n_576)
);

INVxp67_ASAP7_75t_SL g577 ( 
.A(n_393),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_259),
.Y(n_578)
);

NOR2xp67_ASAP7_75t_L g579 ( 
.A(n_269),
.B(n_12),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_269),
.Y(n_580)
);

CKINVDCx20_ASAP7_75t_R g581 ( 
.A(n_355),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_271),
.Y(n_582)
);

NOR2xp33_ASAP7_75t_L g583 ( 
.A(n_263),
.B(n_12),
.Y(n_583)
);

CKINVDCx20_ASAP7_75t_R g584 ( 
.A(n_366),
.Y(n_584)
);

OR2x2_ASAP7_75t_L g585 ( 
.A(n_271),
.B(n_15),
.Y(n_585)
);

NOR2xp33_ASAP7_75t_L g586 ( 
.A(n_270),
.B(n_18),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_274),
.Y(n_587)
);

CKINVDCx5p33_ASAP7_75t_R g588 ( 
.A(n_367),
.Y(n_588)
);

OR2x2_ASAP7_75t_L g589 ( 
.A(n_274),
.B(n_18),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_278),
.Y(n_590)
);

NOR2xp33_ASAP7_75t_L g591 ( 
.A(n_270),
.B(n_23),
.Y(n_591)
);

INVxp67_ASAP7_75t_SL g592 ( 
.A(n_400),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_278),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_L g594 ( 
.A(n_535),
.B(n_372),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_L g595 ( 
.A(n_577),
.B(n_465),
.Y(n_595)
);

INVx3_ASAP7_75t_L g596 ( 
.A(n_518),
.Y(n_596)
);

HB1xp67_ASAP7_75t_L g597 ( 
.A(n_472),
.Y(n_597)
);

INVx2_ASAP7_75t_L g598 ( 
.A(n_518),
.Y(n_598)
);

BUFx6f_ASAP7_75t_L g599 ( 
.A(n_518),
.Y(n_599)
);

AND2x2_ASAP7_75t_L g600 ( 
.A(n_592),
.B(n_400),
.Y(n_600)
);

AND2x2_ASAP7_75t_L g601 ( 
.A(n_511),
.B(n_449),
.Y(n_601)
);

INVx2_ASAP7_75t_L g602 ( 
.A(n_518),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_467),
.Y(n_603)
);

INVx5_ASAP7_75t_L g604 ( 
.A(n_518),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_467),
.Y(n_605)
);

AND2x2_ASAP7_75t_L g606 ( 
.A(n_533),
.B(n_449),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_468),
.Y(n_607)
);

AND2x4_ASAP7_75t_L g608 ( 
.A(n_468),
.B(n_262),
.Y(n_608)
);

CKINVDCx5p33_ASAP7_75t_R g609 ( 
.A(n_509),
.Y(n_609)
);

BUFx6f_ASAP7_75t_L g610 ( 
.A(n_559),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_474),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_L g612 ( 
.A(n_474),
.B(n_373),
.Y(n_612)
);

INVx3_ASAP7_75t_L g613 ( 
.A(n_559),
.Y(n_613)
);

INVx2_ASAP7_75t_L g614 ( 
.A(n_576),
.Y(n_614)
);

INVx2_ASAP7_75t_L g615 ( 
.A(n_576),
.Y(n_615)
);

INVx3_ASAP7_75t_L g616 ( 
.A(n_475),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_475),
.Y(n_617)
);

BUFx2_ASAP7_75t_L g618 ( 
.A(n_488),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_476),
.Y(n_619)
);

INVx3_ASAP7_75t_L g620 ( 
.A(n_476),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_480),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_480),
.Y(n_622)
);

BUFx3_ASAP7_75t_L g623 ( 
.A(n_483),
.Y(n_623)
);

BUFx6f_ASAP7_75t_L g624 ( 
.A(n_483),
.Y(n_624)
);

INVx2_ASAP7_75t_L g625 ( 
.A(n_485),
.Y(n_625)
);

BUFx6f_ASAP7_75t_L g626 ( 
.A(n_485),
.Y(n_626)
);

INVx2_ASAP7_75t_L g627 ( 
.A(n_486),
.Y(n_627)
);

NOR2xp33_ASAP7_75t_L g628 ( 
.A(n_521),
.B(n_290),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_486),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_489),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_L g631 ( 
.A(n_489),
.B(n_380),
.Y(n_631)
);

INVx2_ASAP7_75t_L g632 ( 
.A(n_491),
.Y(n_632)
);

NAND2xp33_ASAP7_75t_L g633 ( 
.A(n_585),
.B(n_299),
.Y(n_633)
);

CKINVDCx5p33_ASAP7_75t_R g634 ( 
.A(n_540),
.Y(n_634)
);

OAI21x1_ASAP7_75t_L g635 ( 
.A1(n_491),
.A2(n_320),
.B(n_262),
.Y(n_635)
);

CKINVDCx20_ASAP7_75t_R g636 ( 
.A(n_471),
.Y(n_636)
);

BUFx6f_ASAP7_75t_L g637 ( 
.A(n_493),
.Y(n_637)
);

HB1xp67_ASAP7_75t_L g638 ( 
.A(n_484),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_493),
.Y(n_639)
);

INVx2_ASAP7_75t_L g640 ( 
.A(n_495),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_495),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_499),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_499),
.Y(n_643)
);

INVx3_ASAP7_75t_L g644 ( 
.A(n_502),
.Y(n_644)
);

HB1xp67_ASAP7_75t_L g645 ( 
.A(n_484),
.Y(n_645)
);

INVx3_ASAP7_75t_L g646 ( 
.A(n_502),
.Y(n_646)
);

BUFx2_ASAP7_75t_L g647 ( 
.A(n_564),
.Y(n_647)
);

AND2x4_ASAP7_75t_L g648 ( 
.A(n_504),
.B(n_320),
.Y(n_648)
);

INVx4_ASAP7_75t_L g649 ( 
.A(n_504),
.Y(n_649)
);

NAND3xp33_ASAP7_75t_L g650 ( 
.A(n_473),
.B(n_292),
.C(n_287),
.Y(n_650)
);

AND2x4_ASAP7_75t_L g651 ( 
.A(n_516),
.B(n_340),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_L g652 ( 
.A(n_516),
.B(n_384),
.Y(n_652)
);

BUFx2_ASAP7_75t_L g653 ( 
.A(n_564),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_520),
.Y(n_654)
);

CKINVDCx5p33_ASAP7_75t_R g655 ( 
.A(n_542),
.Y(n_655)
);

INVxp67_ASAP7_75t_L g656 ( 
.A(n_514),
.Y(n_656)
);

INVx2_ASAP7_75t_L g657 ( 
.A(n_520),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_L g658 ( 
.A(n_523),
.B(n_387),
.Y(n_658)
);

INVx3_ASAP7_75t_L g659 ( 
.A(n_523),
.Y(n_659)
);

HB1xp67_ASAP7_75t_L g660 ( 
.A(n_541),
.Y(n_660)
);

HB1xp67_ASAP7_75t_L g661 ( 
.A(n_548),
.Y(n_661)
);

BUFx6f_ASAP7_75t_L g662 ( 
.A(n_524),
.Y(n_662)
);

AND2x2_ASAP7_75t_L g663 ( 
.A(n_524),
.B(n_438),
.Y(n_663)
);

AND2x6_ASAP7_75t_L g664 ( 
.A(n_526),
.B(n_299),
.Y(n_664)
);

INVx2_ASAP7_75t_L g665 ( 
.A(n_526),
.Y(n_665)
);

BUFx6f_ASAP7_75t_L g666 ( 
.A(n_528),
.Y(n_666)
);

HB1xp67_ASAP7_75t_L g667 ( 
.A(n_562),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_L g668 ( 
.A(n_528),
.B(n_406),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_L g669 ( 
.A(n_530),
.B(n_408),
.Y(n_669)
);

OR2x6_ASAP7_75t_L g670 ( 
.A(n_585),
.B(n_340),
.Y(n_670)
);

INVx3_ASAP7_75t_L g671 ( 
.A(n_530),
.Y(n_671)
);

INVx1_ASAP7_75t_SL g672 ( 
.A(n_481),
.Y(n_672)
);

INVx2_ASAP7_75t_L g673 ( 
.A(n_532),
.Y(n_673)
);

CKINVDCx20_ASAP7_75t_R g674 ( 
.A(n_487),
.Y(n_674)
);

OA21x2_ASAP7_75t_L g675 ( 
.A1(n_532),
.A2(n_534),
.B(n_536),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_534),
.Y(n_676)
);

HB1xp67_ASAP7_75t_L g677 ( 
.A(n_498),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_560),
.Y(n_678)
);

INVx2_ASAP7_75t_L g679 ( 
.A(n_536),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_560),
.Y(n_680)
);

AND2x2_ASAP7_75t_L g681 ( 
.A(n_529),
.B(n_438),
.Y(n_681)
);

BUFx2_ASAP7_75t_L g682 ( 
.A(n_545),
.Y(n_682)
);

NOR2xp33_ASAP7_75t_SL g683 ( 
.A(n_506),
.B(n_293),
.Y(n_683)
);

BUFx6f_ASAP7_75t_L g684 ( 
.A(n_537),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_561),
.Y(n_685)
);

BUFx6f_ASAP7_75t_L g686 ( 
.A(n_537),
.Y(n_686)
);

BUFx6f_ASAP7_75t_L g687 ( 
.A(n_538),
.Y(n_687)
);

INVx3_ASAP7_75t_L g688 ( 
.A(n_538),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_561),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_573),
.Y(n_690)
);

INVx2_ASAP7_75t_L g691 ( 
.A(n_539),
.Y(n_691)
);

BUFx10_ASAP7_75t_L g692 ( 
.A(n_628),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_SL g693 ( 
.A(n_628),
.B(n_507),
.Y(n_693)
);

NOR2xp33_ASAP7_75t_L g694 ( 
.A(n_683),
.B(n_490),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_L g695 ( 
.A(n_594),
.B(n_466),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_675),
.Y(n_696)
);

INVx2_ASAP7_75t_L g697 ( 
.A(n_614),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_675),
.Y(n_698)
);

INVx3_ASAP7_75t_L g699 ( 
.A(n_610),
.Y(n_699)
);

INVx2_ASAP7_75t_L g700 ( 
.A(n_614),
.Y(n_700)
);

OAI21xp33_ASAP7_75t_SL g701 ( 
.A1(n_670),
.A2(n_583),
.B(n_546),
.Y(n_701)
);

INVx2_ASAP7_75t_L g702 ( 
.A(n_614),
.Y(n_702)
);

BUFx2_ASAP7_75t_L g703 ( 
.A(n_647),
.Y(n_703)
);

BUFx6f_ASAP7_75t_L g704 ( 
.A(n_599),
.Y(n_704)
);

INVx3_ASAP7_75t_L g705 ( 
.A(n_610),
.Y(n_705)
);

AND2x2_ASAP7_75t_L g706 ( 
.A(n_600),
.B(n_517),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_SL g707 ( 
.A(n_683),
.B(n_505),
.Y(n_707)
);

INVx2_ASAP7_75t_L g708 ( 
.A(n_614),
.Y(n_708)
);

INVx3_ASAP7_75t_L g709 ( 
.A(n_610),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_SL g710 ( 
.A(n_656),
.B(n_469),
.Y(n_710)
);

INVxp67_ASAP7_75t_SL g711 ( 
.A(n_610),
.Y(n_711)
);

INVx2_ASAP7_75t_L g712 ( 
.A(n_615),
.Y(n_712)
);

NOR2xp33_ASAP7_75t_L g713 ( 
.A(n_594),
.B(n_494),
.Y(n_713)
);

NAND2xp33_ASAP7_75t_L g714 ( 
.A(n_595),
.B(n_677),
.Y(n_714)
);

INVx2_ASAP7_75t_L g715 ( 
.A(n_615),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_L g716 ( 
.A(n_595),
.B(n_470),
.Y(n_716)
);

NOR2xp33_ASAP7_75t_L g717 ( 
.A(n_656),
.B(n_568),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_SL g718 ( 
.A(n_677),
.B(n_477),
.Y(n_718)
);

AND2x4_ASAP7_75t_L g719 ( 
.A(n_670),
.B(n_273),
.Y(n_719)
);

INVx2_ASAP7_75t_SL g720 ( 
.A(n_638),
.Y(n_720)
);

INVx2_ASAP7_75t_L g721 ( 
.A(n_615),
.Y(n_721)
);

NOR2xp33_ASAP7_75t_L g722 ( 
.A(n_682),
.B(n_479),
.Y(n_722)
);

INVx4_ASAP7_75t_L g723 ( 
.A(n_610),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_L g724 ( 
.A(n_612),
.B(n_496),
.Y(n_724)
);

NOR2xp33_ASAP7_75t_L g725 ( 
.A(n_682),
.B(n_500),
.Y(n_725)
);

NOR2xp33_ASAP7_75t_L g726 ( 
.A(n_682),
.B(n_501),
.Y(n_726)
);

INVx5_ASAP7_75t_L g727 ( 
.A(n_664),
.Y(n_727)
);

BUFx6f_ASAP7_75t_L g728 ( 
.A(n_599),
.Y(n_728)
);

NOR2xp33_ASAP7_75t_L g729 ( 
.A(n_600),
.B(n_503),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_SL g730 ( 
.A(n_681),
.B(n_510),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_675),
.Y(n_731)
);

INVx2_ASAP7_75t_SL g732 ( 
.A(n_638),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_675),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_L g734 ( 
.A(n_612),
.B(n_512),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_L g735 ( 
.A(n_631),
.B(n_513),
.Y(n_735)
);

INVx3_ASAP7_75t_L g736 ( 
.A(n_610),
.Y(n_736)
);

NOR2xp33_ASAP7_75t_L g737 ( 
.A(n_600),
.B(n_515),
.Y(n_737)
);

INVx2_ASAP7_75t_L g738 ( 
.A(n_615),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_675),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_L g740 ( 
.A(n_631),
.B(n_519),
.Y(n_740)
);

NAND2xp33_ASAP7_75t_L g741 ( 
.A(n_652),
.B(n_522),
.Y(n_741)
);

INVx8_ASAP7_75t_L g742 ( 
.A(n_670),
.Y(n_742)
);

NOR2xp33_ASAP7_75t_L g743 ( 
.A(n_647),
.B(n_525),
.Y(n_743)
);

AND2x2_ASAP7_75t_L g744 ( 
.A(n_663),
.B(n_554),
.Y(n_744)
);

INVx3_ASAP7_75t_L g745 ( 
.A(n_610),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_675),
.Y(n_746)
);

AND2x2_ASAP7_75t_L g747 ( 
.A(n_663),
.B(n_539),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_623),
.Y(n_748)
);

OAI22xp33_ASAP7_75t_L g749 ( 
.A1(n_670),
.A2(n_245),
.B1(n_302),
.B2(n_291),
.Y(n_749)
);

AND2x2_ASAP7_75t_L g750 ( 
.A(n_663),
.B(n_601),
.Y(n_750)
);

INVx2_ASAP7_75t_L g751 ( 
.A(n_625),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_L g752 ( 
.A(n_652),
.B(n_527),
.Y(n_752)
);

AND2x2_ASAP7_75t_L g753 ( 
.A(n_601),
.B(n_606),
.Y(n_753)
);

NOR2xp33_ASAP7_75t_L g754 ( 
.A(n_647),
.B(n_531),
.Y(n_754)
);

NAND3xp33_ASAP7_75t_L g755 ( 
.A(n_650),
.B(n_591),
.C(n_586),
.Y(n_755)
);

NOR2xp33_ASAP7_75t_L g756 ( 
.A(n_653),
.B(n_547),
.Y(n_756)
);

AOI22xp33_ASAP7_75t_L g757 ( 
.A1(n_670),
.A2(n_579),
.B1(n_589),
.B2(n_549),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_SL g758 ( 
.A(n_681),
.B(n_557),
.Y(n_758)
);

INVx2_ASAP7_75t_L g759 ( 
.A(n_625),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_SL g760 ( 
.A(n_681),
.B(n_565),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_623),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_SL g762 ( 
.A(n_653),
.B(n_566),
.Y(n_762)
);

INVx2_ASAP7_75t_L g763 ( 
.A(n_625),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_L g764 ( 
.A(n_658),
.B(n_569),
.Y(n_764)
);

INVx3_ASAP7_75t_L g765 ( 
.A(n_610),
.Y(n_765)
);

INVx2_ASAP7_75t_SL g766 ( 
.A(n_645),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_623),
.Y(n_767)
);

BUFx3_ASAP7_75t_L g768 ( 
.A(n_623),
.Y(n_768)
);

OAI22xp33_ASAP7_75t_L g769 ( 
.A1(n_670),
.A2(n_368),
.B1(n_403),
.B2(n_326),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_603),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_L g771 ( 
.A(n_658),
.B(n_570),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_603),
.Y(n_772)
);

AOI22xp33_ASAP7_75t_L g773 ( 
.A1(n_670),
.A2(n_589),
.B1(n_478),
.B2(n_292),
.Y(n_773)
);

INVx2_ASAP7_75t_L g774 ( 
.A(n_625),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_605),
.Y(n_775)
);

INVx3_ASAP7_75t_L g776 ( 
.A(n_599),
.Y(n_776)
);

INVxp33_ASAP7_75t_L g777 ( 
.A(n_597),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_605),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_L g779 ( 
.A(n_668),
.B(n_588),
.Y(n_779)
);

AND2x2_ASAP7_75t_L g780 ( 
.A(n_601),
.B(n_544),
.Y(n_780)
);

AND2x2_ASAP7_75t_L g781 ( 
.A(n_606),
.B(n_544),
.Y(n_781)
);

INVx1_ASAP7_75t_L g782 ( 
.A(n_607),
.Y(n_782)
);

INVx2_ASAP7_75t_L g783 ( 
.A(n_627),
.Y(n_783)
);

INVx2_ASAP7_75t_L g784 ( 
.A(n_627),
.Y(n_784)
);

AOI22xp33_ASAP7_75t_L g785 ( 
.A1(n_633),
.A2(n_650),
.B1(n_606),
.B2(n_648),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_L g786 ( 
.A(n_668),
.B(n_669),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_SL g787 ( 
.A(n_653),
.B(n_556),
.Y(n_787)
);

INVx3_ASAP7_75t_L g788 ( 
.A(n_599),
.Y(n_788)
);

INVx3_ASAP7_75t_L g789 ( 
.A(n_599),
.Y(n_789)
);

BUFx2_ASAP7_75t_L g790 ( 
.A(n_645),
.Y(n_790)
);

INVx3_ASAP7_75t_L g791 ( 
.A(n_599),
.Y(n_791)
);

INVx2_ASAP7_75t_L g792 ( 
.A(n_627),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_607),
.Y(n_793)
);

INVx3_ASAP7_75t_L g794 ( 
.A(n_599),
.Y(n_794)
);

INVx2_ASAP7_75t_SL g795 ( 
.A(n_660),
.Y(n_795)
);

INVx4_ASAP7_75t_L g796 ( 
.A(n_624),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_SL g797 ( 
.A(n_660),
.B(n_572),
.Y(n_797)
);

INVx2_ASAP7_75t_L g798 ( 
.A(n_627),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_611),
.Y(n_799)
);

OR2x2_ASAP7_75t_L g800 ( 
.A(n_597),
.B(n_482),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_L g801 ( 
.A(n_669),
.B(n_313),
.Y(n_801)
);

AND2x4_ASAP7_75t_L g802 ( 
.A(n_608),
.B(n_273),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_611),
.Y(n_803)
);

INVx2_ASAP7_75t_L g804 ( 
.A(n_632),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_617),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_617),
.Y(n_806)
);

NOR3xp33_ASAP7_75t_L g807 ( 
.A(n_618),
.B(n_280),
.C(n_276),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_619),
.Y(n_808)
);

INVxp67_ASAP7_75t_L g809 ( 
.A(n_661),
.Y(n_809)
);

OR2x2_ASAP7_75t_L g810 ( 
.A(n_618),
.B(n_497),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_619),
.Y(n_811)
);

NOR2xp33_ASAP7_75t_L g812 ( 
.A(n_661),
.B(n_543),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_SL g813 ( 
.A(n_667),
.B(n_550),
.Y(n_813)
);

AOI22xp33_ASAP7_75t_L g814 ( 
.A1(n_633),
.A2(n_300),
.B1(n_323),
.B2(n_287),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_SL g815 ( 
.A(n_667),
.B(n_551),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_621),
.Y(n_816)
);

INVx2_ASAP7_75t_L g817 ( 
.A(n_632),
.Y(n_817)
);

NAND3xp33_ASAP7_75t_L g818 ( 
.A(n_678),
.B(n_284),
.C(n_275),
.Y(n_818)
);

NOR2xp33_ASAP7_75t_L g819 ( 
.A(n_618),
.B(n_552),
.Y(n_819)
);

INVx2_ASAP7_75t_SL g820 ( 
.A(n_608),
.Y(n_820)
);

INVx2_ASAP7_75t_SL g821 ( 
.A(n_608),
.Y(n_821)
);

AOI22xp5_ASAP7_75t_L g822 ( 
.A1(n_608),
.A2(n_354),
.B1(n_370),
.B2(n_283),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_621),
.Y(n_823)
);

BUFx10_ASAP7_75t_L g824 ( 
.A(n_609),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_L g825 ( 
.A(n_649),
.B(n_418),
.Y(n_825)
);

INVx1_ASAP7_75t_SL g826 ( 
.A(n_672),
.Y(n_826)
);

INVx4_ASAP7_75t_L g827 ( 
.A(n_624),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_622),
.Y(n_828)
);

INVx2_ASAP7_75t_L g829 ( 
.A(n_632),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_622),
.Y(n_830)
);

OR2x6_ASAP7_75t_L g831 ( 
.A(n_608),
.B(n_275),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_629),
.Y(n_832)
);

AND2x2_ASAP7_75t_L g833 ( 
.A(n_678),
.B(n_680),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_SL g834 ( 
.A(n_609),
.B(n_555),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_629),
.Y(n_835)
);

NOR2xp33_ASAP7_75t_L g836 ( 
.A(n_649),
.B(n_558),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_SL g837 ( 
.A(n_634),
.B(n_563),
.Y(n_837)
);

INVx3_ASAP7_75t_L g838 ( 
.A(n_599),
.Y(n_838)
);

BUFx4f_ASAP7_75t_L g839 ( 
.A(n_648),
.Y(n_839)
);

OR2x6_ASAP7_75t_L g840 ( 
.A(n_648),
.B(n_284),
.Y(n_840)
);

INVx2_ASAP7_75t_L g841 ( 
.A(n_632),
.Y(n_841)
);

INVx2_ASAP7_75t_L g842 ( 
.A(n_640),
.Y(n_842)
);

NOR2xp33_ASAP7_75t_L g843 ( 
.A(n_649),
.B(n_567),
.Y(n_843)
);

INVx2_ASAP7_75t_L g844 ( 
.A(n_640),
.Y(n_844)
);

INVx1_ASAP7_75t_SL g845 ( 
.A(n_672),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_SL g846 ( 
.A(n_634),
.B(n_571),
.Y(n_846)
);

INVx2_ASAP7_75t_L g847 ( 
.A(n_640),
.Y(n_847)
);

AOI22xp33_ASAP7_75t_L g848 ( 
.A1(n_648),
.A2(n_323),
.B1(n_357),
.B2(n_300),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_630),
.Y(n_849)
);

AO22x2_ASAP7_75t_L g850 ( 
.A1(n_648),
.A2(n_363),
.B1(n_378),
.B2(n_357),
.Y(n_850)
);

INVx2_ASAP7_75t_L g851 ( 
.A(n_640),
.Y(n_851)
);

BUFx6f_ASAP7_75t_L g852 ( 
.A(n_635),
.Y(n_852)
);

NOR2xp33_ASAP7_75t_L g853 ( 
.A(n_649),
.B(n_581),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_L g854 ( 
.A(n_786),
.B(n_649),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_L g855 ( 
.A(n_713),
.B(n_613),
.Y(n_855)
);

AND2x2_ASAP7_75t_L g856 ( 
.A(n_753),
.B(n_508),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_L g857 ( 
.A(n_801),
.B(n_729),
.Y(n_857)
);

INVx2_ASAP7_75t_L g858 ( 
.A(n_770),
.Y(n_858)
);

AND2x2_ASAP7_75t_L g859 ( 
.A(n_753),
.B(n_492),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_L g860 ( 
.A(n_737),
.B(n_613),
.Y(n_860)
);

INVx2_ASAP7_75t_SL g861 ( 
.A(n_810),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_SL g862 ( 
.A(n_701),
.B(n_299),
.Y(n_862)
);

NOR2xp67_ASAP7_75t_L g863 ( 
.A(n_694),
.B(n_655),
.Y(n_863)
);

NAND2xp33_ASAP7_75t_L g864 ( 
.A(n_742),
.B(n_428),
.Y(n_864)
);

INVx1_ASAP7_75t_L g865 ( 
.A(n_833),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_L g866 ( 
.A(n_695),
.B(n_613),
.Y(n_866)
);

INVx2_ASAP7_75t_L g867 ( 
.A(n_770),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_833),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_748),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_748),
.Y(n_870)
);

NAND2x1p5_ASAP7_75t_L g871 ( 
.A(n_750),
.B(n_635),
.Y(n_871)
);

AOI22xp5_ASAP7_75t_L g872 ( 
.A1(n_714),
.A2(n_701),
.B1(n_706),
.B2(n_750),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_L g873 ( 
.A(n_716),
.B(n_613),
.Y(n_873)
);

INVx2_ASAP7_75t_L g874 ( 
.A(n_772),
.Y(n_874)
);

CKINVDCx5p33_ASAP7_75t_R g875 ( 
.A(n_824),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_L g876 ( 
.A(n_724),
.B(n_613),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_SL g877 ( 
.A(n_692),
.B(n_299),
.Y(n_877)
);

INVx2_ASAP7_75t_L g878 ( 
.A(n_772),
.Y(n_878)
);

NAND2x1_ASAP7_75t_L g879 ( 
.A(n_776),
.B(n_596),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_SL g880 ( 
.A(n_692),
.B(n_343),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_L g881 ( 
.A(n_734),
.B(n_651),
.Y(n_881)
);

AND2x2_ASAP7_75t_SL g882 ( 
.A(n_719),
.B(n_356),
.Y(n_882)
);

INVx2_ASAP7_75t_L g883 ( 
.A(n_775),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_SL g884 ( 
.A(n_692),
.B(n_785),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_761),
.Y(n_885)
);

AND2x6_ASAP7_75t_SL g886 ( 
.A(n_812),
.B(n_363),
.Y(n_886)
);

AO22x2_ASAP7_75t_L g887 ( 
.A1(n_755),
.A2(n_707),
.B1(n_719),
.B2(n_720),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_761),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_L g889 ( 
.A(n_735),
.B(n_651),
.Y(n_889)
);

AOI22xp5_ASAP7_75t_L g890 ( 
.A1(n_706),
.A2(n_755),
.B1(n_741),
.B2(n_719),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_L g891 ( 
.A(n_740),
.B(n_651),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_L g892 ( 
.A(n_752),
.B(n_651),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_SL g893 ( 
.A(n_692),
.B(n_343),
.Y(n_893)
);

INVxp67_ASAP7_75t_L g894 ( 
.A(n_810),
.Y(n_894)
);

INVx1_ASAP7_75t_L g895 ( 
.A(n_767),
.Y(n_895)
);

INVx2_ASAP7_75t_L g896 ( 
.A(n_775),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_SL g897 ( 
.A(n_839),
.B(n_343),
.Y(n_897)
);

BUFx2_ASAP7_75t_L g898 ( 
.A(n_703),
.Y(n_898)
);

NAND2xp5_ASAP7_75t_SL g899 ( 
.A(n_839),
.B(n_343),
.Y(n_899)
);

BUFx6f_ASAP7_75t_L g900 ( 
.A(n_742),
.Y(n_900)
);

NOR2xp33_ASAP7_75t_L g901 ( 
.A(n_722),
.B(n_584),
.Y(n_901)
);

INVx1_ASAP7_75t_L g902 ( 
.A(n_767),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_L g903 ( 
.A(n_764),
.B(n_651),
.Y(n_903)
);

INVx1_ASAP7_75t_L g904 ( 
.A(n_747),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_747),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_820),
.Y(n_906)
);

INVxp67_ASAP7_75t_L g907 ( 
.A(n_725),
.Y(n_907)
);

BUFx3_ASAP7_75t_L g908 ( 
.A(n_768),
.Y(n_908)
);

NOR2xp33_ASAP7_75t_L g909 ( 
.A(n_726),
.B(n_730),
.Y(n_909)
);

INVx2_ASAP7_75t_L g910 ( 
.A(n_778),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_820),
.Y(n_911)
);

BUFx8_ASAP7_75t_L g912 ( 
.A(n_790),
.Y(n_912)
);

INVx1_ASAP7_75t_L g913 ( 
.A(n_821),
.Y(n_913)
);

BUFx8_ASAP7_75t_L g914 ( 
.A(n_790),
.Y(n_914)
);

AO221x1_ASAP7_75t_L g915 ( 
.A1(n_749),
.A2(n_343),
.B1(n_382),
.B2(n_402),
.C(n_405),
.Y(n_915)
);

NAND2xp33_ASAP7_75t_SL g916 ( 
.A(n_795),
.B(n_386),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_821),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_SL g918 ( 
.A(n_839),
.B(n_428),
.Y(n_918)
);

BUFx6f_ASAP7_75t_L g919 ( 
.A(n_742),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_L g920 ( 
.A(n_771),
.B(n_630),
.Y(n_920)
);

BUFx6f_ASAP7_75t_L g921 ( 
.A(n_742),
.Y(n_921)
);

INVx1_ASAP7_75t_L g922 ( 
.A(n_780),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_780),
.Y(n_923)
);

AOI22xp5_ASAP7_75t_L g924 ( 
.A1(n_719),
.A2(n_424),
.B1(n_425),
.B2(n_423),
.Y(n_924)
);

INVx2_ASAP7_75t_L g925 ( 
.A(n_778),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_L g926 ( 
.A(n_779),
.B(n_639),
.Y(n_926)
);

INVx1_ASAP7_75t_L g927 ( 
.A(n_781),
.Y(n_927)
);

NAND2xp33_ASAP7_75t_L g928 ( 
.A(n_742),
.B(n_852),
.Y(n_928)
);

NAND2xp33_ASAP7_75t_L g929 ( 
.A(n_852),
.B(n_757),
.Y(n_929)
);

INVx2_ASAP7_75t_L g930 ( 
.A(n_782),
.Y(n_930)
);

OAI22xp33_ASAP7_75t_L g931 ( 
.A1(n_720),
.A2(n_298),
.B1(n_305),
.B2(n_294),
.Y(n_931)
);

NAND2xp5_ASAP7_75t_SL g932 ( 
.A(n_852),
.B(n_696),
.Y(n_932)
);

INVx2_ASAP7_75t_L g933 ( 
.A(n_782),
.Y(n_933)
);

CKINVDCx5p33_ASAP7_75t_R g934 ( 
.A(n_824),
.Y(n_934)
);

INVx2_ASAP7_75t_SL g935 ( 
.A(n_732),
.Y(n_935)
);

NAND2xp5_ASAP7_75t_SL g936 ( 
.A(n_852),
.B(n_428),
.Y(n_936)
);

NAND2xp5_ASAP7_75t_L g937 ( 
.A(n_696),
.B(n_639),
.Y(n_937)
);

O2A1O1Ixp33_ASAP7_75t_L g938 ( 
.A1(n_698),
.A2(n_685),
.B(n_689),
.C(n_680),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_L g939 ( 
.A(n_698),
.B(n_641),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_L g940 ( 
.A(n_731),
.B(n_641),
.Y(n_940)
);

INVx2_ASAP7_75t_L g941 ( 
.A(n_793),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_L g942 ( 
.A(n_731),
.B(n_642),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_L g943 ( 
.A(n_733),
.B(n_642),
.Y(n_943)
);

BUFx6f_ASAP7_75t_SL g944 ( 
.A(n_824),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_SL g945 ( 
.A(n_852),
.B(n_428),
.Y(n_945)
);

INVx1_ASAP7_75t_L g946 ( 
.A(n_781),
.Y(n_946)
);

INVx1_ASAP7_75t_L g947 ( 
.A(n_793),
.Y(n_947)
);

OAI22xp5_ASAP7_75t_L g948 ( 
.A1(n_758),
.A2(n_381),
.B1(n_356),
.B2(n_298),
.Y(n_948)
);

A2O1A1Ixp33_ASAP7_75t_L g949 ( 
.A1(n_733),
.A2(n_635),
.B(n_381),
.C(n_305),
.Y(n_949)
);

NOR2xp33_ASAP7_75t_L g950 ( 
.A(n_760),
.B(n_285),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_L g951 ( 
.A(n_739),
.B(n_643),
.Y(n_951)
);

AOI22xp5_ASAP7_75t_L g952 ( 
.A1(n_836),
.A2(n_444),
.B1(n_445),
.B2(n_436),
.Y(n_952)
);

INVx2_ASAP7_75t_L g953 ( 
.A(n_799),
.Y(n_953)
);

INVx1_ASAP7_75t_L g954 ( 
.A(n_799),
.Y(n_954)
);

INVx2_ASAP7_75t_L g955 ( 
.A(n_803),
.Y(n_955)
);

NAND2xp33_ASAP7_75t_L g956 ( 
.A(n_739),
.B(n_428),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_L g957 ( 
.A(n_746),
.B(n_643),
.Y(n_957)
);

INVxp67_ASAP7_75t_L g958 ( 
.A(n_743),
.Y(n_958)
);

NOR2xp33_ASAP7_75t_L g959 ( 
.A(n_717),
.B(n_289),
.Y(n_959)
);

INVx1_ASAP7_75t_L g960 ( 
.A(n_803),
.Y(n_960)
);

INVxp67_ASAP7_75t_L g961 ( 
.A(n_754),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_L g962 ( 
.A(n_746),
.B(n_654),
.Y(n_962)
);

NAND2xp5_ASAP7_75t_L g963 ( 
.A(n_805),
.B(n_654),
.Y(n_963)
);

NAND2xp5_ASAP7_75t_L g964 ( 
.A(n_805),
.B(n_676),
.Y(n_964)
);

NAND2xp5_ASAP7_75t_SL g965 ( 
.A(n_843),
.B(n_853),
.Y(n_965)
);

CKINVDCx5p33_ASAP7_75t_R g966 ( 
.A(n_824),
.Y(n_966)
);

NAND2xp5_ASAP7_75t_SL g967 ( 
.A(n_756),
.B(n_428),
.Y(n_967)
);

NAND2xp5_ASAP7_75t_L g968 ( 
.A(n_806),
.B(n_676),
.Y(n_968)
);

AND2x2_ASAP7_75t_L g969 ( 
.A(n_795),
.B(n_655),
.Y(n_969)
);

AOI22xp5_ASAP7_75t_L g970 ( 
.A1(n_744),
.A2(n_462),
.B1(n_294),
.B2(n_310),
.Y(n_970)
);

NOR2xp33_ASAP7_75t_L g971 ( 
.A(n_693),
.B(n_304),
.Y(n_971)
);

NAND2xp5_ASAP7_75t_L g972 ( 
.A(n_806),
.B(n_688),
.Y(n_972)
);

INVx2_ASAP7_75t_L g973 ( 
.A(n_808),
.Y(n_973)
);

AND2x2_ASAP7_75t_L g974 ( 
.A(n_732),
.B(n_685),
.Y(n_974)
);

NAND2xp5_ASAP7_75t_L g975 ( 
.A(n_808),
.B(n_688),
.Y(n_975)
);

INVx2_ASAP7_75t_SL g976 ( 
.A(n_766),
.Y(n_976)
);

INVx2_ASAP7_75t_L g977 ( 
.A(n_811),
.Y(n_977)
);

NAND2xp5_ASAP7_75t_L g978 ( 
.A(n_811),
.B(n_688),
.Y(n_978)
);

INVx3_ASAP7_75t_L g979 ( 
.A(n_768),
.Y(n_979)
);

NAND2xp5_ASAP7_75t_L g980 ( 
.A(n_816),
.B(n_688),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_SL g981 ( 
.A(n_802),
.B(n_428),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_L g982 ( 
.A(n_816),
.B(n_688),
.Y(n_982)
);

AOI22xp5_ASAP7_75t_L g983 ( 
.A1(n_744),
.A2(n_307),
.B1(n_316),
.B2(n_310),
.Y(n_983)
);

INVx1_ASAP7_75t_L g984 ( 
.A(n_823),
.Y(n_984)
);

NAND2xp5_ASAP7_75t_L g985 ( 
.A(n_823),
.B(n_616),
.Y(n_985)
);

NOR2xp67_ASAP7_75t_L g986 ( 
.A(n_809),
.B(n_689),
.Y(n_986)
);

NAND2xp5_ASAP7_75t_L g987 ( 
.A(n_828),
.B(n_616),
.Y(n_987)
);

INVx2_ASAP7_75t_L g988 ( 
.A(n_828),
.Y(n_988)
);

INVx1_ASAP7_75t_L g989 ( 
.A(n_830),
.Y(n_989)
);

NAND2xp5_ASAP7_75t_SL g990 ( 
.A(n_802),
.B(n_684),
.Y(n_990)
);

INVx2_ASAP7_75t_L g991 ( 
.A(n_830),
.Y(n_991)
);

INVx3_ASAP7_75t_L g992 ( 
.A(n_768),
.Y(n_992)
);

INVx2_ASAP7_75t_L g993 ( 
.A(n_832),
.Y(n_993)
);

INVxp67_ASAP7_75t_L g994 ( 
.A(n_819),
.Y(n_994)
);

INVx2_ASAP7_75t_L g995 ( 
.A(n_832),
.Y(n_995)
);

INVx2_ASAP7_75t_L g996 ( 
.A(n_835),
.Y(n_996)
);

NAND2xp5_ASAP7_75t_SL g997 ( 
.A(n_802),
.B(n_684),
.Y(n_997)
);

NAND2xp5_ASAP7_75t_L g998 ( 
.A(n_835),
.B(n_616),
.Y(n_998)
);

NOR2xp33_ASAP7_75t_L g999 ( 
.A(n_718),
.B(n_306),
.Y(n_999)
);

INVx1_ASAP7_75t_L g1000 ( 
.A(n_849),
.Y(n_1000)
);

INVx1_ASAP7_75t_L g1001 ( 
.A(n_849),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_L g1002 ( 
.A(n_711),
.B(n_616),
.Y(n_1002)
);

NOR2xp33_ASAP7_75t_L g1003 ( 
.A(n_710),
.B(n_317),
.Y(n_1003)
);

AND2x2_ASAP7_75t_SL g1004 ( 
.A(n_814),
.B(n_307),
.Y(n_1004)
);

A2O1A1Ixp33_ASAP7_75t_L g1005 ( 
.A1(n_802),
.A2(n_324),
.B(n_347),
.C(n_316),
.Y(n_1005)
);

NOR2xp33_ASAP7_75t_L g1006 ( 
.A(n_762),
.B(n_318),
.Y(n_1006)
);

AND2x4_ASAP7_75t_L g1007 ( 
.A(n_831),
.B(n_690),
.Y(n_1007)
);

INVx1_ASAP7_75t_L g1008 ( 
.A(n_831),
.Y(n_1008)
);

NOR2xp33_ASAP7_75t_SL g1009 ( 
.A(n_826),
.B(n_636),
.Y(n_1009)
);

AOI22xp33_ASAP7_75t_L g1010 ( 
.A1(n_850),
.A2(n_379),
.B1(n_382),
.B2(n_378),
.Y(n_1010)
);

NAND2xp5_ASAP7_75t_L g1011 ( 
.A(n_825),
.B(n_616),
.Y(n_1011)
);

NAND2xp5_ASAP7_75t_L g1012 ( 
.A(n_699),
.B(n_620),
.Y(n_1012)
);

INVx1_ASAP7_75t_L g1013 ( 
.A(n_831),
.Y(n_1013)
);

NOR2xp33_ASAP7_75t_L g1014 ( 
.A(n_766),
.B(n_325),
.Y(n_1014)
);

NAND2xp5_ASAP7_75t_L g1015 ( 
.A(n_699),
.B(n_620),
.Y(n_1015)
);

INVx1_ASAP7_75t_L g1016 ( 
.A(n_831),
.Y(n_1016)
);

NAND2xp5_ASAP7_75t_L g1017 ( 
.A(n_699),
.B(n_620),
.Y(n_1017)
);

INVx8_ASAP7_75t_L g1018 ( 
.A(n_831),
.Y(n_1018)
);

INVx2_ASAP7_75t_L g1019 ( 
.A(n_697),
.Y(n_1019)
);

INVx2_ASAP7_75t_L g1020 ( 
.A(n_697),
.Y(n_1020)
);

NOR2xp67_ASAP7_75t_L g1021 ( 
.A(n_800),
.B(n_690),
.Y(n_1021)
);

AOI22xp5_ASAP7_75t_L g1022 ( 
.A1(n_807),
.A2(n_347),
.B1(n_353),
.B2(n_324),
.Y(n_1022)
);

NOR3xp33_ASAP7_75t_L g1023 ( 
.A(n_787),
.B(n_328),
.C(n_327),
.Y(n_1023)
);

NOR2xp33_ASAP7_75t_L g1024 ( 
.A(n_769),
.B(n_330),
.Y(n_1024)
);

AOI22xp33_ASAP7_75t_L g1025 ( 
.A1(n_850),
.A2(n_416),
.B1(n_422),
.B2(n_410),
.Y(n_1025)
);

NAND2x1p5_ASAP7_75t_L g1026 ( 
.A(n_727),
.B(n_353),
.Y(n_1026)
);

NAND2xp5_ASAP7_75t_L g1027 ( 
.A(n_857),
.B(n_773),
.Y(n_1027)
);

INVx2_ASAP7_75t_L g1028 ( 
.A(n_858),
.Y(n_1028)
);

BUFx3_ASAP7_75t_L g1029 ( 
.A(n_898),
.Y(n_1029)
);

AOI21xp5_ASAP7_75t_L g1030 ( 
.A1(n_929),
.A2(n_723),
.B(n_796),
.Y(n_1030)
);

AOI21xp5_ASAP7_75t_L g1031 ( 
.A1(n_881),
.A2(n_723),
.B(n_796),
.Y(n_1031)
);

NOR2xp33_ASAP7_75t_L g1032 ( 
.A(n_907),
.B(n_703),
.Y(n_1032)
);

A2O1A1Ixp33_ASAP7_75t_L g1033 ( 
.A1(n_909),
.A2(n_818),
.B(n_822),
.C(n_848),
.Y(n_1033)
);

INVx4_ASAP7_75t_L g1034 ( 
.A(n_900),
.Y(n_1034)
);

NAND2xp5_ASAP7_75t_L g1035 ( 
.A(n_920),
.B(n_699),
.Y(n_1035)
);

INVx1_ASAP7_75t_L g1036 ( 
.A(n_858),
.Y(n_1036)
);

INVx1_ASAP7_75t_SL g1037 ( 
.A(n_969),
.Y(n_1037)
);

AO21x1_ASAP7_75t_L g1038 ( 
.A1(n_862),
.A2(n_884),
.B(n_965),
.Y(n_1038)
);

OAI21xp5_ASAP7_75t_L g1039 ( 
.A1(n_932),
.A2(n_709),
.B(n_705),
.Y(n_1039)
);

AOI33xp33_ASAP7_75t_L g1040 ( 
.A1(n_861),
.A2(n_575),
.A3(n_573),
.B1(n_574),
.B2(n_578),
.B3(n_580),
.Y(n_1040)
);

AOI22xp5_ASAP7_75t_L g1041 ( 
.A1(n_909),
.A2(n_813),
.B1(n_815),
.B2(n_840),
.Y(n_1041)
);

AND2x4_ASAP7_75t_L g1042 ( 
.A(n_865),
.B(n_826),
.Y(n_1042)
);

NOR2xp33_ASAP7_75t_L g1043 ( 
.A(n_958),
.B(n_822),
.Y(n_1043)
);

BUFx3_ASAP7_75t_L g1044 ( 
.A(n_912),
.Y(n_1044)
);

NAND2xp5_ASAP7_75t_L g1045 ( 
.A(n_926),
.B(n_705),
.Y(n_1045)
);

INVx1_ASAP7_75t_L g1046 ( 
.A(n_867),
.Y(n_1046)
);

NAND2xp5_ASAP7_75t_SL g1047 ( 
.A(n_872),
.B(n_845),
.Y(n_1047)
);

INVx2_ASAP7_75t_L g1048 ( 
.A(n_874),
.Y(n_1048)
);

O2A1O1Ixp33_ASAP7_75t_L g1049 ( 
.A1(n_884),
.A2(n_840),
.B(n_818),
.C(n_797),
.Y(n_1049)
);

OAI21xp5_ASAP7_75t_L g1050 ( 
.A1(n_932),
.A2(n_709),
.B(n_705),
.Y(n_1050)
);

AOI21xp5_ASAP7_75t_L g1051 ( 
.A1(n_889),
.A2(n_723),
.B(n_796),
.Y(n_1051)
);

INVx3_ASAP7_75t_L g1052 ( 
.A(n_908),
.Y(n_1052)
);

NAND2xp5_ASAP7_75t_L g1053 ( 
.A(n_855),
.B(n_705),
.Y(n_1053)
);

AOI21x1_ASAP7_75t_L g1054 ( 
.A1(n_936),
.A2(n_702),
.B(n_700),
.Y(n_1054)
);

OAI21xp5_ASAP7_75t_L g1055 ( 
.A1(n_862),
.A2(n_736),
.B(n_709),
.Y(n_1055)
);

NAND2xp5_ASAP7_75t_L g1056 ( 
.A(n_854),
.B(n_860),
.Y(n_1056)
);

NAND2xp5_ASAP7_75t_SL g1057 ( 
.A(n_890),
.B(n_845),
.Y(n_1057)
);

A2O1A1Ixp33_ASAP7_75t_L g1058 ( 
.A1(n_959),
.A2(n_388),
.B(n_402),
.C(n_379),
.Y(n_1058)
);

HB1xp67_ASAP7_75t_L g1059 ( 
.A(n_894),
.Y(n_1059)
);

AOI21xp5_ASAP7_75t_L g1060 ( 
.A1(n_891),
.A2(n_723),
.B(n_796),
.Y(n_1060)
);

AOI21xp5_ASAP7_75t_L g1061 ( 
.A1(n_892),
.A2(n_827),
.B(n_728),
.Y(n_1061)
);

BUFx2_ASAP7_75t_L g1062 ( 
.A(n_859),
.Y(n_1062)
);

NAND2xp5_ASAP7_75t_L g1063 ( 
.A(n_947),
.B(n_709),
.Y(n_1063)
);

NAND2xp5_ASAP7_75t_L g1064 ( 
.A(n_954),
.B(n_736),
.Y(n_1064)
);

NAND2xp5_ASAP7_75t_L g1065 ( 
.A(n_960),
.B(n_736),
.Y(n_1065)
);

NAND2xp5_ASAP7_75t_L g1066 ( 
.A(n_984),
.B(n_736),
.Y(n_1066)
);

AOI21xp5_ASAP7_75t_L g1067 ( 
.A1(n_903),
.A2(n_827),
.B(n_728),
.Y(n_1067)
);

NAND2xp5_ASAP7_75t_L g1068 ( 
.A(n_989),
.B(n_745),
.Y(n_1068)
);

INVx1_ASAP7_75t_SL g1069 ( 
.A(n_1009),
.Y(n_1069)
);

NOR2xp33_ASAP7_75t_SL g1070 ( 
.A(n_901),
.B(n_636),
.Y(n_1070)
);

NOR3xp33_ASAP7_75t_L g1071 ( 
.A(n_901),
.B(n_837),
.C(n_834),
.Y(n_1071)
);

INVxp67_ASAP7_75t_SL g1072 ( 
.A(n_979),
.Y(n_1072)
);

INVx11_ASAP7_75t_L g1073 ( 
.A(n_912),
.Y(n_1073)
);

NOR2xp33_ASAP7_75t_L g1074 ( 
.A(n_961),
.B(n_777),
.Y(n_1074)
);

AND2x2_ASAP7_75t_L g1075 ( 
.A(n_856),
.B(n_800),
.Y(n_1075)
);

NAND2xp5_ASAP7_75t_L g1076 ( 
.A(n_1000),
.B(n_745),
.Y(n_1076)
);

INVx1_ASAP7_75t_L g1077 ( 
.A(n_874),
.Y(n_1077)
);

INVx2_ASAP7_75t_L g1078 ( 
.A(n_878),
.Y(n_1078)
);

OAI22xp5_ASAP7_75t_L g1079 ( 
.A1(n_882),
.A2(n_840),
.B1(n_850),
.B2(n_369),
.Y(n_1079)
);

INVx3_ASAP7_75t_L g1080 ( 
.A(n_908),
.Y(n_1080)
);

AND2x4_ASAP7_75t_L g1081 ( 
.A(n_868),
.B(n_840),
.Y(n_1081)
);

NAND2xp5_ASAP7_75t_L g1082 ( 
.A(n_1001),
.B(n_959),
.Y(n_1082)
);

AOI21xp5_ASAP7_75t_L g1083 ( 
.A1(n_876),
.A2(n_827),
.B(n_728),
.Y(n_1083)
);

OAI21xp5_ASAP7_75t_L g1084 ( 
.A1(n_871),
.A2(n_765),
.B(n_745),
.Y(n_1084)
);

AOI21xp5_ASAP7_75t_L g1085 ( 
.A1(n_866),
.A2(n_827),
.B(n_728),
.Y(n_1085)
);

BUFx6f_ASAP7_75t_L g1086 ( 
.A(n_900),
.Y(n_1086)
);

O2A1O1Ixp5_ASAP7_75t_L g1087 ( 
.A1(n_877),
.A2(n_765),
.B(n_745),
.C(n_776),
.Y(n_1087)
);

AND2x4_ASAP7_75t_L g1088 ( 
.A(n_922),
.B(n_840),
.Y(n_1088)
);

NAND2xp33_ASAP7_75t_L g1089 ( 
.A(n_900),
.B(n_704),
.Y(n_1089)
);

NOR3xp33_ASAP7_75t_L g1090 ( 
.A(n_994),
.B(n_846),
.C(n_369),
.Y(n_1090)
);

NAND2xp5_ASAP7_75t_L g1091 ( 
.A(n_878),
.B(n_765),
.Y(n_1091)
);

A2O1A1Ixp33_ASAP7_75t_L g1092 ( 
.A1(n_1024),
.A2(n_405),
.B(n_410),
.C(n_388),
.Y(n_1092)
);

AOI22xp5_ASAP7_75t_L g1093 ( 
.A1(n_965),
.A2(n_850),
.B1(n_765),
.B2(n_674),
.Y(n_1093)
);

INVx1_ASAP7_75t_L g1094 ( 
.A(n_883),
.Y(n_1094)
);

AOI22xp33_ASAP7_75t_L g1095 ( 
.A1(n_1004),
.A2(n_422),
.B1(n_430),
.B2(n_416),
.Y(n_1095)
);

AOI21xp5_ASAP7_75t_L g1096 ( 
.A1(n_873),
.A2(n_728),
.B(n_704),
.Y(n_1096)
);

AOI22xp5_ASAP7_75t_L g1097 ( 
.A1(n_882),
.A2(n_674),
.B1(n_788),
.B2(n_776),
.Y(n_1097)
);

AOI21xp5_ASAP7_75t_L g1098 ( 
.A1(n_864),
.A2(n_704),
.B(n_727),
.Y(n_1098)
);

AOI21xp5_ASAP7_75t_L g1099 ( 
.A1(n_979),
.A2(n_704),
.B(n_727),
.Y(n_1099)
);

NAND2xp5_ASAP7_75t_SL g1100 ( 
.A(n_900),
.B(n_919),
.Y(n_1100)
);

NOR2xp33_ASAP7_75t_L g1101 ( 
.A(n_935),
.B(n_401),
.Y(n_1101)
);

NAND2xp5_ASAP7_75t_SL g1102 ( 
.A(n_919),
.B(n_727),
.Y(n_1102)
);

OAI321xp33_ASAP7_75t_L g1103 ( 
.A1(n_1024),
.A2(n_435),
.A3(n_430),
.B1(n_457),
.B2(n_383),
.C(n_429),
.Y(n_1103)
);

AOI21xp5_ASAP7_75t_L g1104 ( 
.A1(n_992),
.A2(n_704),
.B(n_727),
.Y(n_1104)
);

NOR2xp33_ASAP7_75t_SL g1105 ( 
.A(n_875),
.B(n_447),
.Y(n_1105)
);

NAND2xp5_ASAP7_75t_L g1106 ( 
.A(n_883),
.B(n_776),
.Y(n_1106)
);

NAND2xp5_ASAP7_75t_SL g1107 ( 
.A(n_919),
.B(n_727),
.Y(n_1107)
);

INVx1_ASAP7_75t_L g1108 ( 
.A(n_896),
.Y(n_1108)
);

AOI21xp5_ASAP7_75t_L g1109 ( 
.A1(n_992),
.A2(n_789),
.B(n_788),
.Y(n_1109)
);

INVx2_ASAP7_75t_L g1110 ( 
.A(n_896),
.Y(n_1110)
);

OAI21xp5_ASAP7_75t_L g1111 ( 
.A1(n_871),
.A2(n_702),
.B(n_700),
.Y(n_1111)
);

INVx2_ASAP7_75t_L g1112 ( 
.A(n_910),
.Y(n_1112)
);

AOI21xp5_ASAP7_75t_L g1113 ( 
.A1(n_1011),
.A2(n_928),
.B(n_956),
.Y(n_1113)
);

NAND2xp5_ASAP7_75t_L g1114 ( 
.A(n_910),
.B(n_788),
.Y(n_1114)
);

AOI21xp5_ASAP7_75t_L g1115 ( 
.A1(n_937),
.A2(n_940),
.B(n_939),
.Y(n_1115)
);

INVx1_ASAP7_75t_L g1116 ( 
.A(n_925),
.Y(n_1116)
);

OAI21xp5_ASAP7_75t_L g1117 ( 
.A1(n_936),
.A2(n_712),
.B(n_708),
.Y(n_1117)
);

BUFx3_ASAP7_75t_L g1118 ( 
.A(n_914),
.Y(n_1118)
);

INVx2_ASAP7_75t_L g1119 ( 
.A(n_925),
.Y(n_1119)
);

NAND2xp5_ASAP7_75t_L g1120 ( 
.A(n_930),
.B(n_788),
.Y(n_1120)
);

NAND2xp5_ASAP7_75t_L g1121 ( 
.A(n_930),
.B(n_789),
.Y(n_1121)
);

NAND2xp5_ASAP7_75t_L g1122 ( 
.A(n_933),
.B(n_941),
.Y(n_1122)
);

NAND2xp5_ASAP7_75t_L g1123 ( 
.A(n_933),
.B(n_789),
.Y(n_1123)
);

AND2x2_ASAP7_75t_L g1124 ( 
.A(n_974),
.B(n_293),
.Y(n_1124)
);

OAI21xp5_ASAP7_75t_L g1125 ( 
.A1(n_945),
.A2(n_712),
.B(n_708),
.Y(n_1125)
);

BUFx3_ASAP7_75t_L g1126 ( 
.A(n_914),
.Y(n_1126)
);

NAND2xp5_ASAP7_75t_L g1127 ( 
.A(n_941),
.B(n_789),
.Y(n_1127)
);

AND2x4_ASAP7_75t_L g1128 ( 
.A(n_923),
.B(n_574),
.Y(n_1128)
);

NOR2xp33_ASAP7_75t_L g1129 ( 
.A(n_976),
.B(n_448),
.Y(n_1129)
);

OAI22x1_ASAP7_75t_L g1130 ( 
.A1(n_1006),
.A2(n_342),
.B1(n_349),
.B2(n_338),
.Y(n_1130)
);

AOI21xp5_ASAP7_75t_L g1131 ( 
.A1(n_942),
.A2(n_794),
.B(n_791),
.Y(n_1131)
);

A2O1A1Ixp33_ASAP7_75t_L g1132 ( 
.A1(n_1010),
.A2(n_1025),
.B(n_938),
.C(n_971),
.Y(n_1132)
);

NOR2xp33_ASAP7_75t_L g1133 ( 
.A(n_1014),
.B(n_791),
.Y(n_1133)
);

BUFx6f_ASAP7_75t_L g1134 ( 
.A(n_919),
.Y(n_1134)
);

OAI21xp5_ASAP7_75t_L g1135 ( 
.A1(n_945),
.A2(n_721),
.B(n_715),
.Y(n_1135)
);

INVx1_ASAP7_75t_L g1136 ( 
.A(n_953),
.Y(n_1136)
);

INVx2_ASAP7_75t_SL g1137 ( 
.A(n_887),
.Y(n_1137)
);

AOI21xp5_ASAP7_75t_L g1138 ( 
.A1(n_943),
.A2(n_794),
.B(n_791),
.Y(n_1138)
);

AOI21xp5_ASAP7_75t_L g1139 ( 
.A1(n_951),
.A2(n_794),
.B(n_791),
.Y(n_1139)
);

INVx1_ASAP7_75t_L g1140 ( 
.A(n_953),
.Y(n_1140)
);

INVx2_ASAP7_75t_L g1141 ( 
.A(n_955),
.Y(n_1141)
);

BUFx8_ASAP7_75t_L g1142 ( 
.A(n_944),
.Y(n_1142)
);

NAND2xp5_ASAP7_75t_L g1143 ( 
.A(n_955),
.B(n_794),
.Y(n_1143)
);

AOI21xp5_ASAP7_75t_L g1144 ( 
.A1(n_957),
.A2(n_838),
.B(n_604),
.Y(n_1144)
);

AOI21xp5_ASAP7_75t_L g1145 ( 
.A1(n_962),
.A2(n_838),
.B(n_604),
.Y(n_1145)
);

OAI22xp5_ASAP7_75t_L g1146 ( 
.A1(n_906),
.A2(n_361),
.B1(n_375),
.B2(n_383),
.Y(n_1146)
);

OAI321xp33_ASAP7_75t_L g1147 ( 
.A1(n_931),
.A2(n_435),
.A3(n_442),
.B1(n_361),
.B2(n_453),
.C(n_412),
.Y(n_1147)
);

AOI21xp5_ASAP7_75t_L g1148 ( 
.A1(n_1002),
.A2(n_838),
.B(n_604),
.Y(n_1148)
);

AOI21xp5_ASAP7_75t_L g1149 ( 
.A1(n_990),
.A2(n_838),
.B(n_604),
.Y(n_1149)
);

NAND2xp5_ASAP7_75t_L g1150 ( 
.A(n_973),
.B(n_715),
.Y(n_1150)
);

OR2x2_ASAP7_75t_L g1151 ( 
.A(n_927),
.B(n_575),
.Y(n_1151)
);

AO21x1_ASAP7_75t_L g1152 ( 
.A1(n_967),
.A2(n_392),
.B(n_375),
.Y(n_1152)
);

INVx1_ASAP7_75t_SL g1153 ( 
.A(n_916),
.Y(n_1153)
);

NAND2xp5_ASAP7_75t_L g1154 ( 
.A(n_973),
.B(n_721),
.Y(n_1154)
);

AOI21xp5_ASAP7_75t_L g1155 ( 
.A1(n_990),
.A2(n_604),
.B(n_738),
.Y(n_1155)
);

NAND2xp5_ASAP7_75t_L g1156 ( 
.A(n_977),
.B(n_738),
.Y(n_1156)
);

NOR2xp33_ASAP7_75t_L g1157 ( 
.A(n_1014),
.B(n_350),
.Y(n_1157)
);

INVx3_ASAP7_75t_L g1158 ( 
.A(n_977),
.Y(n_1158)
);

OAI22xp5_ASAP7_75t_L g1159 ( 
.A1(n_911),
.A2(n_392),
.B1(n_396),
.B2(n_412),
.Y(n_1159)
);

OAI21xp5_ASAP7_75t_L g1160 ( 
.A1(n_949),
.A2(n_759),
.B(n_751),
.Y(n_1160)
);

OAI21xp33_ASAP7_75t_L g1161 ( 
.A1(n_1006),
.A2(n_352),
.B(n_351),
.Y(n_1161)
);

AOI21xp5_ASAP7_75t_L g1162 ( 
.A1(n_997),
.A2(n_899),
.B(n_897),
.Y(n_1162)
);

NOR2xp33_ASAP7_75t_SL g1163 ( 
.A(n_934),
.B(n_238),
.Y(n_1163)
);

OAI22xp5_ASAP7_75t_L g1164 ( 
.A1(n_913),
.A2(n_396),
.B1(n_413),
.B2(n_429),
.Y(n_1164)
);

AOI21xp5_ASAP7_75t_L g1165 ( 
.A1(n_997),
.A2(n_604),
.B(n_751),
.Y(n_1165)
);

NAND2xp5_ASAP7_75t_L g1166 ( 
.A(n_988),
.B(n_759),
.Y(n_1166)
);

INVx1_ASAP7_75t_L g1167 ( 
.A(n_988),
.Y(n_1167)
);

INVx2_ASAP7_75t_L g1168 ( 
.A(n_991),
.Y(n_1168)
);

NAND2xp5_ASAP7_75t_L g1169 ( 
.A(n_991),
.B(n_763),
.Y(n_1169)
);

AOI21xp5_ASAP7_75t_L g1170 ( 
.A1(n_897),
.A2(n_604),
.B(n_763),
.Y(n_1170)
);

OAI22xp5_ASAP7_75t_SL g1171 ( 
.A1(n_1003),
.A2(n_362),
.B1(n_358),
.B2(n_359),
.Y(n_1171)
);

BUFx6f_ASAP7_75t_L g1172 ( 
.A(n_921),
.Y(n_1172)
);

AOI21xp5_ASAP7_75t_L g1173 ( 
.A1(n_899),
.A2(n_604),
.B(n_774),
.Y(n_1173)
);

AND2x2_ASAP7_75t_L g1174 ( 
.A(n_1021),
.B(n_439),
.Y(n_1174)
);

OR2x2_ASAP7_75t_L g1175 ( 
.A(n_946),
.B(n_578),
.Y(n_1175)
);

OAI22xp5_ASAP7_75t_L g1176 ( 
.A1(n_917),
.A2(n_413),
.B1(n_442),
.B2(n_446),
.Y(n_1176)
);

INVx2_ASAP7_75t_L g1177 ( 
.A(n_993),
.Y(n_1177)
);

AOI21xp5_ASAP7_75t_L g1178 ( 
.A1(n_918),
.A2(n_604),
.B(n_774),
.Y(n_1178)
);

AOI21xp5_ASAP7_75t_L g1179 ( 
.A1(n_918),
.A2(n_784),
.B(n_783),
.Y(n_1179)
);

NAND2xp5_ASAP7_75t_SL g1180 ( 
.A(n_921),
.B(n_783),
.Y(n_1180)
);

AOI21xp5_ASAP7_75t_L g1181 ( 
.A1(n_1012),
.A2(n_792),
.B(n_784),
.Y(n_1181)
);

AOI21xp5_ASAP7_75t_L g1182 ( 
.A1(n_1015),
.A2(n_798),
.B(n_792),
.Y(n_1182)
);

BUFx2_ASAP7_75t_L g1183 ( 
.A(n_887),
.Y(n_1183)
);

INVx1_ASAP7_75t_L g1184 ( 
.A(n_993),
.Y(n_1184)
);

AOI21xp5_ASAP7_75t_L g1185 ( 
.A1(n_1017),
.A2(n_804),
.B(n_798),
.Y(n_1185)
);

AOI21xp5_ASAP7_75t_L g1186 ( 
.A1(n_972),
.A2(n_817),
.B(n_804),
.Y(n_1186)
);

AOI21xp5_ASAP7_75t_L g1187 ( 
.A1(n_975),
.A2(n_829),
.B(n_817),
.Y(n_1187)
);

INVxp67_ASAP7_75t_L g1188 ( 
.A(n_950),
.Y(n_1188)
);

AOI21xp5_ASAP7_75t_L g1189 ( 
.A1(n_978),
.A2(n_841),
.B(n_829),
.Y(n_1189)
);

NOR2xp67_ASAP7_75t_L g1190 ( 
.A(n_966),
.B(n_580),
.Y(n_1190)
);

OAI21xp33_ASAP7_75t_SL g1191 ( 
.A1(n_995),
.A2(n_452),
.B(n_446),
.Y(n_1191)
);

HB1xp67_ASAP7_75t_L g1192 ( 
.A(n_904),
.Y(n_1192)
);

INVx2_ASAP7_75t_SL g1193 ( 
.A(n_887),
.Y(n_1193)
);

AOI21xp5_ASAP7_75t_L g1194 ( 
.A1(n_980),
.A2(n_842),
.B(n_841),
.Y(n_1194)
);

AOI21xp5_ASAP7_75t_L g1195 ( 
.A1(n_982),
.A2(n_844),
.B(n_842),
.Y(n_1195)
);

NAND2xp5_ASAP7_75t_L g1196 ( 
.A(n_995),
.B(n_844),
.Y(n_1196)
);

NAND2xp5_ASAP7_75t_L g1197 ( 
.A(n_996),
.B(n_847),
.Y(n_1197)
);

NAND2xp5_ASAP7_75t_L g1198 ( 
.A(n_996),
.B(n_847),
.Y(n_1198)
);

NAND2xp5_ASAP7_75t_L g1199 ( 
.A(n_905),
.B(n_851),
.Y(n_1199)
);

NOR2xp33_ASAP7_75t_L g1200 ( 
.A(n_971),
.B(n_360),
.Y(n_1200)
);

NAND2xp5_ASAP7_75t_L g1201 ( 
.A(n_869),
.B(n_851),
.Y(n_1201)
);

NAND2xp5_ASAP7_75t_L g1202 ( 
.A(n_870),
.B(n_452),
.Y(n_1202)
);

NAND2xp5_ASAP7_75t_SL g1203 ( 
.A(n_921),
.B(n_1007),
.Y(n_1203)
);

NAND2xp5_ASAP7_75t_SL g1204 ( 
.A(n_921),
.B(n_684),
.Y(n_1204)
);

OAI21xp5_ASAP7_75t_L g1205 ( 
.A1(n_877),
.A2(n_457),
.B(n_453),
.Y(n_1205)
);

AOI21xp5_ASAP7_75t_L g1206 ( 
.A1(n_985),
.A2(n_596),
.B(n_598),
.Y(n_1206)
);

INVx3_ASAP7_75t_L g1207 ( 
.A(n_1007),
.Y(n_1207)
);

NAND2xp5_ASAP7_75t_SL g1208 ( 
.A(n_1010),
.B(n_684),
.Y(n_1208)
);

HB1xp67_ASAP7_75t_L g1209 ( 
.A(n_986),
.Y(n_1209)
);

NAND2xp5_ASAP7_75t_L g1210 ( 
.A(n_885),
.B(n_620),
.Y(n_1210)
);

NOR3xp33_ASAP7_75t_L g1211 ( 
.A(n_1003),
.B(n_371),
.C(n_364),
.Y(n_1211)
);

O2A1O1Ixp5_ASAP7_75t_L g1212 ( 
.A1(n_880),
.A2(n_620),
.B(n_644),
.C(n_646),
.Y(n_1212)
);

AND2x4_ASAP7_75t_L g1213 ( 
.A(n_1008),
.B(n_582),
.Y(n_1213)
);

INVx1_ASAP7_75t_SL g1214 ( 
.A(n_950),
.Y(n_1214)
);

NAND2xp5_ASAP7_75t_L g1215 ( 
.A(n_888),
.B(n_644),
.Y(n_1215)
);

NAND2xp5_ASAP7_75t_SL g1216 ( 
.A(n_1025),
.B(n_684),
.Y(n_1216)
);

OAI21x1_ASAP7_75t_L g1217 ( 
.A1(n_987),
.A2(n_646),
.B(n_644),
.Y(n_1217)
);

INVx2_ASAP7_75t_L g1218 ( 
.A(n_1019),
.Y(n_1218)
);

NAND2xp5_ASAP7_75t_L g1219 ( 
.A(n_895),
.B(n_644),
.Y(n_1219)
);

AOI21xp5_ASAP7_75t_L g1220 ( 
.A1(n_998),
.A2(n_596),
.B(n_598),
.Y(n_1220)
);

HB1xp67_ASAP7_75t_L g1221 ( 
.A(n_1029),
.Y(n_1221)
);

NOR2xp67_ASAP7_75t_L g1222 ( 
.A(n_1188),
.B(n_863),
.Y(n_1222)
);

INVx2_ASAP7_75t_L g1223 ( 
.A(n_1028),
.Y(n_1223)
);

OAI21x1_ASAP7_75t_L g1224 ( 
.A1(n_1054),
.A2(n_902),
.B(n_879),
.Y(n_1224)
);

O2A1O1Ixp33_ASAP7_75t_L g1225 ( 
.A1(n_1200),
.A2(n_948),
.B(n_967),
.C(n_999),
.Y(n_1225)
);

AND2x4_ASAP7_75t_L g1226 ( 
.A(n_1207),
.B(n_1013),
.Y(n_1226)
);

AOI21xp5_ASAP7_75t_L g1227 ( 
.A1(n_1115),
.A2(n_1018),
.B(n_893),
.Y(n_1227)
);

INVx1_ASAP7_75t_L g1228 ( 
.A(n_1078),
.Y(n_1228)
);

INVx2_ASAP7_75t_L g1229 ( 
.A(n_1078),
.Y(n_1229)
);

O2A1O1Ixp33_ASAP7_75t_L g1230 ( 
.A1(n_1200),
.A2(n_1047),
.B(n_1157),
.C(n_1057),
.Y(n_1230)
);

AOI21xp5_ASAP7_75t_L g1231 ( 
.A1(n_1113),
.A2(n_1018),
.B(n_893),
.Y(n_1231)
);

INVx1_ASAP7_75t_L g1232 ( 
.A(n_1110),
.Y(n_1232)
);

NOR2xp67_ASAP7_75t_SL g1233 ( 
.A(n_1086),
.B(n_1016),
.Y(n_1233)
);

AOI21xp5_ASAP7_75t_L g1234 ( 
.A1(n_1056),
.A2(n_1018),
.B(n_880),
.Y(n_1234)
);

INVx1_ASAP7_75t_L g1235 ( 
.A(n_1110),
.Y(n_1235)
);

INVx2_ASAP7_75t_L g1236 ( 
.A(n_1112),
.Y(n_1236)
);

AOI21xp5_ASAP7_75t_L g1237 ( 
.A1(n_1089),
.A2(n_981),
.B(n_1026),
.Y(n_1237)
);

NOR2xp33_ASAP7_75t_R g1238 ( 
.A(n_1070),
.B(n_944),
.Y(n_1238)
);

NAND2x1p5_ASAP7_75t_L g1239 ( 
.A(n_1034),
.B(n_981),
.Y(n_1239)
);

OR2x2_ASAP7_75t_L g1240 ( 
.A(n_1075),
.B(n_999),
.Y(n_1240)
);

AOI21xp5_ASAP7_75t_L g1241 ( 
.A1(n_1030),
.A2(n_1026),
.B(n_964),
.Y(n_1241)
);

A2O1A1Ixp33_ASAP7_75t_L g1242 ( 
.A1(n_1132),
.A2(n_1004),
.B(n_983),
.C(n_1022),
.Y(n_1242)
);

INVx2_ASAP7_75t_L g1243 ( 
.A(n_1141),
.Y(n_1243)
);

OAI22xp5_ASAP7_75t_L g1244 ( 
.A1(n_1082),
.A2(n_924),
.B1(n_952),
.B2(n_970),
.Y(n_1244)
);

AOI21x1_ASAP7_75t_L g1245 ( 
.A1(n_1180),
.A2(n_968),
.B(n_963),
.Y(n_1245)
);

AND2x4_ASAP7_75t_L g1246 ( 
.A(n_1207),
.B(n_1023),
.Y(n_1246)
);

NAND2x1p5_ASAP7_75t_L g1247 ( 
.A(n_1034),
.B(n_1020),
.Y(n_1247)
);

INVx2_ASAP7_75t_SL g1248 ( 
.A(n_1029),
.Y(n_1248)
);

BUFx2_ASAP7_75t_L g1249 ( 
.A(n_1062),
.Y(n_1249)
);

NAND2xp5_ASAP7_75t_L g1250 ( 
.A(n_1027),
.B(n_915),
.Y(n_1250)
);

INVx2_ASAP7_75t_L g1251 ( 
.A(n_1141),
.Y(n_1251)
);

BUFx2_ASAP7_75t_L g1252 ( 
.A(n_1042),
.Y(n_1252)
);

NAND3xp33_ASAP7_75t_L g1253 ( 
.A(n_1157),
.B(n_1005),
.C(n_376),
.Y(n_1253)
);

NAND2xp5_ASAP7_75t_L g1254 ( 
.A(n_1214),
.B(n_1047),
.Y(n_1254)
);

OAI22xp5_ASAP7_75t_L g1255 ( 
.A1(n_1132),
.A2(n_1020),
.B1(n_1019),
.B2(n_458),
.Y(n_1255)
);

INVx1_ASAP7_75t_L g1256 ( 
.A(n_1168),
.Y(n_1256)
);

AOI21xp5_ASAP7_75t_L g1257 ( 
.A1(n_1061),
.A2(n_1067),
.B(n_1051),
.Y(n_1257)
);

A2O1A1Ixp33_ASAP7_75t_L g1258 ( 
.A1(n_1033),
.A2(n_582),
.B(n_587),
.C(n_590),
.Y(n_1258)
);

AOI21xp5_ASAP7_75t_L g1259 ( 
.A1(n_1031),
.A2(n_596),
.B(n_598),
.Y(n_1259)
);

BUFx3_ASAP7_75t_L g1260 ( 
.A(n_1044),
.Y(n_1260)
);

INVx2_ASAP7_75t_SL g1261 ( 
.A(n_1042),
.Y(n_1261)
);

INVx2_ASAP7_75t_L g1262 ( 
.A(n_1168),
.Y(n_1262)
);

NOR2xp33_ASAP7_75t_SL g1263 ( 
.A(n_1105),
.B(n_238),
.Y(n_1263)
);

INVxp33_ASAP7_75t_SL g1264 ( 
.A(n_1074),
.Y(n_1264)
);

AOI21xp5_ASAP7_75t_L g1265 ( 
.A1(n_1060),
.A2(n_596),
.B(n_598),
.Y(n_1265)
);

OAI22xp5_ASAP7_75t_L g1266 ( 
.A1(n_1097),
.A2(n_1133),
.B1(n_1057),
.B2(n_1033),
.Y(n_1266)
);

BUFx3_ASAP7_75t_L g1267 ( 
.A(n_1044),
.Y(n_1267)
);

INVx2_ASAP7_75t_L g1268 ( 
.A(n_1177),
.Y(n_1268)
);

NAND2xp5_ASAP7_75t_L g1269 ( 
.A(n_1209),
.B(n_679),
.Y(n_1269)
);

BUFx2_ASAP7_75t_L g1270 ( 
.A(n_1059),
.Y(n_1270)
);

NOR2xp33_ASAP7_75t_L g1271 ( 
.A(n_1043),
.B(n_886),
.Y(n_1271)
);

NAND2xp5_ASAP7_75t_L g1272 ( 
.A(n_1209),
.B(n_679),
.Y(n_1272)
);

AOI22xp5_ASAP7_75t_L g1273 ( 
.A1(n_1071),
.A2(n_238),
.B1(n_308),
.B2(n_348),
.Y(n_1273)
);

AOI21xp5_ASAP7_75t_L g1274 ( 
.A1(n_1035),
.A2(n_1045),
.B(n_1083),
.Y(n_1274)
);

CKINVDCx16_ASAP7_75t_R g1275 ( 
.A(n_1118),
.Y(n_1275)
);

NOR2x1_ASAP7_75t_L g1276 ( 
.A(n_1052),
.B(n_587),
.Y(n_1276)
);

INVx1_ASAP7_75t_L g1277 ( 
.A(n_1177),
.Y(n_1277)
);

INVx3_ASAP7_75t_L g1278 ( 
.A(n_1086),
.Y(n_1278)
);

AOI21xp5_ASAP7_75t_L g1279 ( 
.A1(n_1085),
.A2(n_602),
.B(n_644),
.Y(n_1279)
);

AO22x1_ASAP7_75t_L g1280 ( 
.A1(n_1043),
.A2(n_421),
.B1(n_464),
.B2(n_463),
.Y(n_1280)
);

INVx1_ASAP7_75t_L g1281 ( 
.A(n_1036),
.Y(n_1281)
);

AOI21xp5_ASAP7_75t_L g1282 ( 
.A1(n_1162),
.A2(n_602),
.B(n_646),
.Y(n_1282)
);

AOI21x1_ASAP7_75t_L g1283 ( 
.A1(n_1180),
.A2(n_602),
.B(n_657),
.Y(n_1283)
);

AND2x2_ASAP7_75t_L g1284 ( 
.A(n_1124),
.B(n_439),
.Y(n_1284)
);

AND2x2_ASAP7_75t_L g1285 ( 
.A(n_1037),
.B(n_439),
.Y(n_1285)
);

INVx1_ASAP7_75t_SL g1286 ( 
.A(n_1069),
.Y(n_1286)
);

OAI22x1_ASAP7_75t_L g1287 ( 
.A1(n_1041),
.A2(n_374),
.B1(n_377),
.B2(n_385),
.Y(n_1287)
);

NAND2xp5_ASAP7_75t_L g1288 ( 
.A(n_1192),
.B(n_679),
.Y(n_1288)
);

NOR3xp33_ASAP7_75t_L g1289 ( 
.A(n_1171),
.B(n_593),
.C(n_590),
.Y(n_1289)
);

OAI22xp5_ASAP7_75t_L g1290 ( 
.A1(n_1133),
.A2(n_451),
.B1(n_389),
.B2(n_390),
.Y(n_1290)
);

BUFx6f_ASAP7_75t_L g1291 ( 
.A(n_1086),
.Y(n_1291)
);

NAND2xp5_ASAP7_75t_SL g1292 ( 
.A(n_1038),
.B(n_238),
.Y(n_1292)
);

OAI22xp5_ASAP7_75t_L g1293 ( 
.A1(n_1137),
.A2(n_455),
.B1(n_391),
.B2(n_394),
.Y(n_1293)
);

NAND2xp5_ASAP7_75t_L g1294 ( 
.A(n_1192),
.B(n_679),
.Y(n_1294)
);

NAND2xp5_ASAP7_75t_L g1295 ( 
.A(n_1174),
.B(n_691),
.Y(n_1295)
);

NAND3xp33_ASAP7_75t_SL g1296 ( 
.A(n_1163),
.B(n_443),
.C(n_415),
.Y(n_1296)
);

INVx5_ASAP7_75t_L g1297 ( 
.A(n_1086),
.Y(n_1297)
);

NOR3xp33_ASAP7_75t_SL g1298 ( 
.A(n_1032),
.B(n_432),
.C(n_459),
.Y(n_1298)
);

HB1xp67_ASAP7_75t_L g1299 ( 
.A(n_1059),
.Y(n_1299)
);

NAND2xp5_ASAP7_75t_L g1300 ( 
.A(n_1032),
.B(n_1128),
.Y(n_1300)
);

CKINVDCx16_ASAP7_75t_R g1301 ( 
.A(n_1118),
.Y(n_1301)
);

AOI21xp5_ASAP7_75t_L g1302 ( 
.A1(n_1084),
.A2(n_602),
.B(n_659),
.Y(n_1302)
);

INVxp67_ASAP7_75t_L g1303 ( 
.A(n_1074),
.Y(n_1303)
);

INVx2_ASAP7_75t_L g1304 ( 
.A(n_1158),
.Y(n_1304)
);

OAI22xp5_ASAP7_75t_L g1305 ( 
.A1(n_1193),
.A2(n_456),
.B1(n_395),
.B2(n_398),
.Y(n_1305)
);

BUFx6f_ASAP7_75t_L g1306 ( 
.A(n_1134),
.Y(n_1306)
);

OAI22xp5_ASAP7_75t_L g1307 ( 
.A1(n_1093),
.A2(n_1072),
.B1(n_1080),
.B2(n_1052),
.Y(n_1307)
);

A2O1A1Ixp33_ASAP7_75t_L g1308 ( 
.A1(n_1095),
.A2(n_593),
.B(n_399),
.C(n_411),
.Y(n_1308)
);

INVx3_ASAP7_75t_L g1309 ( 
.A(n_1134),
.Y(n_1309)
);

BUFx12f_ASAP7_75t_L g1310 ( 
.A(n_1142),
.Y(n_1310)
);

A2O1A1Ixp33_ASAP7_75t_L g1311 ( 
.A1(n_1095),
.A2(n_450),
.B(n_414),
.C(n_417),
.Y(n_1311)
);

NAND2xp5_ASAP7_75t_SL g1312 ( 
.A(n_1049),
.B(n_308),
.Y(n_1312)
);

NOR2xp33_ASAP7_75t_L g1313 ( 
.A(n_1101),
.B(n_419),
.Y(n_1313)
);

NAND2xp5_ASAP7_75t_L g1314 ( 
.A(n_1128),
.B(n_691),
.Y(n_1314)
);

AOI21xp5_ASAP7_75t_L g1315 ( 
.A1(n_1111),
.A2(n_646),
.B(n_659),
.Y(n_1315)
);

INVx1_ASAP7_75t_L g1316 ( 
.A(n_1046),
.Y(n_1316)
);

OAI22xp5_ASAP7_75t_L g1317 ( 
.A1(n_1080),
.A2(n_427),
.B1(n_441),
.B2(n_440),
.Y(n_1317)
);

INVx1_ASAP7_75t_L g1318 ( 
.A(n_1077),
.Y(n_1318)
);

AND2x2_ASAP7_75t_L g1319 ( 
.A(n_1101),
.B(n_439),
.Y(n_1319)
);

OAI21xp5_ASAP7_75t_L g1320 ( 
.A1(n_1087),
.A2(n_1212),
.B(n_1138),
.Y(n_1320)
);

AOI21xp5_ASAP7_75t_L g1321 ( 
.A1(n_1053),
.A2(n_646),
.B(n_659),
.Y(n_1321)
);

OAI21xp5_ASAP7_75t_L g1322 ( 
.A1(n_1131),
.A2(n_659),
.B(n_671),
.Y(n_1322)
);

OAI21x1_ASAP7_75t_L g1323 ( 
.A1(n_1217),
.A2(n_671),
.B(n_659),
.Y(n_1323)
);

OR2x6_ASAP7_75t_L g1324 ( 
.A(n_1126),
.B(n_553),
.Y(n_1324)
);

HAxp5_ASAP7_75t_L g1325 ( 
.A(n_1129),
.B(n_420),
.CON(n_1325),
.SN(n_1325)
);

OAI22xp5_ASAP7_75t_L g1326 ( 
.A1(n_1203),
.A2(n_434),
.B1(n_454),
.B2(n_671),
.Y(n_1326)
);

NAND2xp5_ASAP7_75t_L g1327 ( 
.A(n_1158),
.B(n_691),
.Y(n_1327)
);

INVx1_ASAP7_75t_L g1328 ( 
.A(n_1094),
.Y(n_1328)
);

INVx2_ASAP7_75t_L g1329 ( 
.A(n_1218),
.Y(n_1329)
);

AOI21xp5_ASAP7_75t_L g1330 ( 
.A1(n_1096),
.A2(n_671),
.B(n_657),
.Y(n_1330)
);

O2A1O1Ixp33_ASAP7_75t_L g1331 ( 
.A1(n_1092),
.A2(n_553),
.B(n_691),
.C(n_671),
.Y(n_1331)
);

NAND2xp5_ASAP7_75t_SL g1332 ( 
.A(n_1081),
.B(n_308),
.Y(n_1332)
);

NAND2xp5_ASAP7_75t_SL g1333 ( 
.A(n_1081),
.B(n_308),
.Y(n_1333)
);

NOR2xp33_ASAP7_75t_L g1334 ( 
.A(n_1129),
.B(n_23),
.Y(n_1334)
);

INVx1_ASAP7_75t_L g1335 ( 
.A(n_1108),
.Y(n_1335)
);

OAI22xp5_ASAP7_75t_L g1336 ( 
.A1(n_1203),
.A2(n_673),
.B1(n_657),
.B2(n_665),
.Y(n_1336)
);

AOI21xp5_ASAP7_75t_L g1337 ( 
.A1(n_1122),
.A2(n_665),
.B(n_657),
.Y(n_1337)
);

BUFx2_ASAP7_75t_L g1338 ( 
.A(n_1183),
.Y(n_1338)
);

AND2x2_ASAP7_75t_L g1339 ( 
.A(n_1153),
.B(n_348),
.Y(n_1339)
);

INVx2_ASAP7_75t_L g1340 ( 
.A(n_1218),
.Y(n_1340)
);

AOI22xp5_ASAP7_75t_L g1341 ( 
.A1(n_1211),
.A2(n_348),
.B1(n_686),
.B2(n_684),
.Y(n_1341)
);

NAND2xp5_ASAP7_75t_SL g1342 ( 
.A(n_1088),
.B(n_348),
.Y(n_1342)
);

NOR2xp33_ASAP7_75t_L g1343 ( 
.A(n_1161),
.B(n_25),
.Y(n_1343)
);

O2A1O1Ixp33_ASAP7_75t_L g1344 ( 
.A1(n_1092),
.A2(n_1058),
.B(n_1103),
.C(n_1090),
.Y(n_1344)
);

NOR2xp33_ASAP7_75t_L g1345 ( 
.A(n_1151),
.B(n_26),
.Y(n_1345)
);

INVx3_ASAP7_75t_L g1346 ( 
.A(n_1134),
.Y(n_1346)
);

AOI21xp5_ASAP7_75t_L g1347 ( 
.A1(n_1204),
.A2(n_665),
.B(n_673),
.Y(n_1347)
);

INVx3_ASAP7_75t_L g1348 ( 
.A(n_1134),
.Y(n_1348)
);

NAND2xp5_ASAP7_75t_L g1349 ( 
.A(n_1116),
.B(n_684),
.Y(n_1349)
);

OAI22xp5_ASAP7_75t_L g1350 ( 
.A1(n_1136),
.A2(n_665),
.B1(n_673),
.B2(n_684),
.Y(n_1350)
);

NAND2xp5_ASAP7_75t_L g1351 ( 
.A(n_1140),
.B(n_686),
.Y(n_1351)
);

INVx1_ASAP7_75t_L g1352 ( 
.A(n_1167),
.Y(n_1352)
);

AOI21xp5_ASAP7_75t_L g1353 ( 
.A1(n_1204),
.A2(n_673),
.B(n_626),
.Y(n_1353)
);

NAND2xp5_ASAP7_75t_L g1354 ( 
.A(n_1184),
.B(n_686),
.Y(n_1354)
);

AND2x4_ASAP7_75t_L g1355 ( 
.A(n_1088),
.B(n_96),
.Y(n_1355)
);

BUFx6f_ASAP7_75t_L g1356 ( 
.A(n_1172),
.Y(n_1356)
);

AO21x2_ASAP7_75t_L g1357 ( 
.A1(n_1160),
.A2(n_687),
.B(n_686),
.Y(n_1357)
);

AOI22xp33_ASAP7_75t_L g1358 ( 
.A1(n_1079),
.A2(n_687),
.B1(n_686),
.B2(n_664),
.Y(n_1358)
);

BUFx2_ASAP7_75t_L g1359 ( 
.A(n_1213),
.Y(n_1359)
);

NOR2xp33_ASAP7_75t_L g1360 ( 
.A(n_1175),
.B(n_26),
.Y(n_1360)
);

AOI21xp5_ASAP7_75t_L g1361 ( 
.A1(n_1099),
.A2(n_662),
.B(n_626),
.Y(n_1361)
);

NAND2xp5_ASAP7_75t_SL g1362 ( 
.A(n_1172),
.B(n_686),
.Y(n_1362)
);

NAND2xp5_ASAP7_75t_SL g1363 ( 
.A(n_1172),
.B(n_686),
.Y(n_1363)
);

INVx2_ASAP7_75t_L g1364 ( 
.A(n_1048),
.Y(n_1364)
);

AND2x2_ASAP7_75t_L g1365 ( 
.A(n_1190),
.B(n_1213),
.Y(n_1365)
);

CKINVDCx5p33_ASAP7_75t_R g1366 ( 
.A(n_1073),
.Y(n_1366)
);

INVxp67_ASAP7_75t_L g1367 ( 
.A(n_1202),
.Y(n_1367)
);

BUFx3_ASAP7_75t_L g1368 ( 
.A(n_1126),
.Y(n_1368)
);

OAI22xp5_ASAP7_75t_L g1369 ( 
.A1(n_1119),
.A2(n_1172),
.B1(n_1199),
.B2(n_1100),
.Y(n_1369)
);

NOR2xp33_ASAP7_75t_L g1370 ( 
.A(n_1063),
.B(n_27),
.Y(n_1370)
);

NOR3xp33_ASAP7_75t_SL g1371 ( 
.A(n_1147),
.B(n_27),
.C(n_28),
.Y(n_1371)
);

INVx6_ASAP7_75t_L g1372 ( 
.A(n_1142),
.Y(n_1372)
);

A2O1A1Ixp33_ASAP7_75t_L g1373 ( 
.A1(n_1058),
.A2(n_687),
.B(n_686),
.C(n_32),
.Y(n_1373)
);

INVxp67_ASAP7_75t_SL g1374 ( 
.A(n_1208),
.Y(n_1374)
);

INVxp67_ASAP7_75t_L g1375 ( 
.A(n_1146),
.Y(n_1375)
);

NAND2xp5_ASAP7_75t_L g1376 ( 
.A(n_1040),
.B(n_687),
.Y(n_1376)
);

AND2x2_ASAP7_75t_SL g1377 ( 
.A(n_1040),
.B(n_687),
.Y(n_1377)
);

INVx1_ASAP7_75t_L g1378 ( 
.A(n_1201),
.Y(n_1378)
);

OR2x2_ASAP7_75t_L g1379 ( 
.A(n_1130),
.B(n_687),
.Y(n_1379)
);

O2A1O1Ixp33_ASAP7_75t_L g1380 ( 
.A1(n_1159),
.A2(n_28),
.B(n_30),
.C(n_33),
.Y(n_1380)
);

NAND2xp5_ASAP7_75t_SL g1381 ( 
.A(n_1039),
.B(n_687),
.Y(n_1381)
);

NAND2xp5_ASAP7_75t_L g1382 ( 
.A(n_1166),
.B(n_687),
.Y(n_1382)
);

INVx1_ASAP7_75t_L g1383 ( 
.A(n_1169),
.Y(n_1383)
);

INVx1_ASAP7_75t_L g1384 ( 
.A(n_1196),
.Y(n_1384)
);

NAND2xp5_ASAP7_75t_SL g1385 ( 
.A(n_1050),
.B(n_624),
.Y(n_1385)
);

AO31x2_ASAP7_75t_L g1386 ( 
.A1(n_1266),
.A2(n_1152),
.A3(n_1164),
.B(n_1176),
.Y(n_1386)
);

AOI21xp5_ASAP7_75t_L g1387 ( 
.A1(n_1227),
.A2(n_1274),
.B(n_1241),
.Y(n_1387)
);

INVx1_ASAP7_75t_L g1388 ( 
.A(n_1281),
.Y(n_1388)
);

AOI21xp5_ASAP7_75t_L g1389 ( 
.A1(n_1257),
.A2(n_1100),
.B(n_1098),
.Y(n_1389)
);

INVx2_ASAP7_75t_L g1390 ( 
.A(n_1223),
.Y(n_1390)
);

CKINVDCx5p33_ASAP7_75t_R g1391 ( 
.A(n_1310),
.Y(n_1391)
);

OAI21x1_ASAP7_75t_L g1392 ( 
.A1(n_1323),
.A2(n_1179),
.B(n_1139),
.Y(n_1392)
);

OAI21x1_ASAP7_75t_L g1393 ( 
.A1(n_1283),
.A2(n_1187),
.B(n_1186),
.Y(n_1393)
);

AOI21xp5_ASAP7_75t_L g1394 ( 
.A1(n_1234),
.A2(n_1055),
.B(n_1107),
.Y(n_1394)
);

AOI21xp5_ASAP7_75t_L g1395 ( 
.A1(n_1231),
.A2(n_1107),
.B(n_1102),
.Y(n_1395)
);

AO31x2_ASAP7_75t_L g1396 ( 
.A1(n_1258),
.A2(n_1189),
.A3(n_1194),
.B(n_1195),
.Y(n_1396)
);

AOI21x1_ASAP7_75t_SL g1397 ( 
.A1(n_1250),
.A2(n_1064),
.B(n_1076),
.Y(n_1397)
);

HB1xp67_ASAP7_75t_L g1398 ( 
.A(n_1299),
.Y(n_1398)
);

AOI221xp5_ASAP7_75t_SL g1399 ( 
.A1(n_1242),
.A2(n_1205),
.B1(n_1191),
.B2(n_1216),
.C(n_1208),
.Y(n_1399)
);

HB1xp67_ASAP7_75t_L g1400 ( 
.A(n_1299),
.Y(n_1400)
);

O2A1O1Ixp5_ASAP7_75t_L g1401 ( 
.A1(n_1312),
.A2(n_1102),
.B(n_1216),
.C(n_1135),
.Y(n_1401)
);

NOR2xp33_ASAP7_75t_SL g1402 ( 
.A(n_1263),
.B(n_1065),
.Y(n_1402)
);

HB1xp67_ASAP7_75t_L g1403 ( 
.A(n_1270),
.Y(n_1403)
);

AOI21xp5_ASAP7_75t_L g1404 ( 
.A1(n_1230),
.A2(n_1091),
.B(n_1198),
.Y(n_1404)
);

INVx1_ASAP7_75t_SL g1405 ( 
.A(n_1286),
.Y(n_1405)
);

INVx1_ASAP7_75t_L g1406 ( 
.A(n_1316),
.Y(n_1406)
);

NAND2xp5_ASAP7_75t_SL g1407 ( 
.A(n_1264),
.B(n_1066),
.Y(n_1407)
);

INVx1_ASAP7_75t_L g1408 ( 
.A(n_1318),
.Y(n_1408)
);

O2A1O1Ixp33_ASAP7_75t_L g1409 ( 
.A1(n_1334),
.A2(n_1068),
.B(n_1219),
.C(n_1215),
.Y(n_1409)
);

NAND2xp5_ASAP7_75t_L g1410 ( 
.A(n_1254),
.B(n_1300),
.Y(n_1410)
);

O2A1O1Ixp5_ASAP7_75t_L g1411 ( 
.A1(n_1312),
.A2(n_1117),
.B(n_1125),
.C(n_1181),
.Y(n_1411)
);

NOR2xp33_ASAP7_75t_L g1412 ( 
.A(n_1303),
.B(n_1106),
.Y(n_1412)
);

OR2x2_ASAP7_75t_L g1413 ( 
.A(n_1240),
.B(n_1197),
.Y(n_1413)
);

OAI21xp5_ASAP7_75t_L g1414 ( 
.A1(n_1225),
.A2(n_1182),
.B(n_1185),
.Y(n_1414)
);

O2A1O1Ixp33_ASAP7_75t_L g1415 ( 
.A1(n_1334),
.A2(n_1271),
.B(n_1313),
.C(n_1325),
.Y(n_1415)
);

NAND2xp5_ASAP7_75t_L g1416 ( 
.A(n_1367),
.B(n_1150),
.Y(n_1416)
);

A2O1A1Ixp33_ASAP7_75t_L g1417 ( 
.A1(n_1313),
.A2(n_1220),
.B(n_1206),
.C(n_1144),
.Y(n_1417)
);

OAI21xp5_ASAP7_75t_L g1418 ( 
.A1(n_1242),
.A2(n_1127),
.B(n_1114),
.Y(n_1418)
);

AND2x2_ASAP7_75t_L g1419 ( 
.A(n_1284),
.B(n_1120),
.Y(n_1419)
);

NAND2xp5_ASAP7_75t_L g1420 ( 
.A(n_1367),
.B(n_1154),
.Y(n_1420)
);

O2A1O1Ixp33_ASAP7_75t_SL g1421 ( 
.A1(n_1308),
.A2(n_1210),
.B(n_1121),
.C(n_1123),
.Y(n_1421)
);

AND2x4_ASAP7_75t_L g1422 ( 
.A(n_1355),
.B(n_1143),
.Y(n_1422)
);

NOR2xp67_ASAP7_75t_L g1423 ( 
.A(n_1261),
.B(n_1149),
.Y(n_1423)
);

OAI21x1_ASAP7_75t_L g1424 ( 
.A1(n_1224),
.A2(n_1109),
.B(n_1148),
.Y(n_1424)
);

NOR2xp33_ASAP7_75t_L g1425 ( 
.A(n_1303),
.B(n_1156),
.Y(n_1425)
);

BUFx10_ASAP7_75t_L g1426 ( 
.A(n_1372),
.Y(n_1426)
);

O2A1O1Ixp5_ASAP7_75t_SL g1427 ( 
.A1(n_1292),
.A2(n_1173),
.B(n_1170),
.C(n_1178),
.Y(n_1427)
);

O2A1O1Ixp33_ASAP7_75t_L g1428 ( 
.A1(n_1271),
.A2(n_1145),
.B(n_1165),
.C(n_1155),
.Y(n_1428)
);

INVx1_ASAP7_75t_L g1429 ( 
.A(n_1328),
.Y(n_1429)
);

AND2x2_ASAP7_75t_L g1430 ( 
.A(n_1252),
.B(n_34),
.Y(n_1430)
);

AOI21xp5_ASAP7_75t_L g1431 ( 
.A1(n_1295),
.A2(n_1104),
.B(n_666),
.Y(n_1431)
);

NAND2xp5_ASAP7_75t_L g1432 ( 
.A(n_1378),
.B(n_36),
.Y(n_1432)
);

AOI22xp33_ASAP7_75t_L g1433 ( 
.A1(n_1343),
.A2(n_664),
.B1(n_662),
.B2(n_637),
.Y(n_1433)
);

AO31x2_ASAP7_75t_L g1434 ( 
.A1(n_1258),
.A2(n_664),
.A3(n_41),
.B(n_42),
.Y(n_1434)
);

OAI21xp5_ASAP7_75t_L g1435 ( 
.A1(n_1321),
.A2(n_664),
.B(n_666),
.Y(n_1435)
);

AOI221x1_ASAP7_75t_L g1436 ( 
.A1(n_1343),
.A2(n_666),
.B1(n_662),
.B2(n_637),
.C(n_626),
.Y(n_1436)
);

NOR2xp33_ASAP7_75t_L g1437 ( 
.A(n_1249),
.B(n_36),
.Y(n_1437)
);

OAI22xp5_ASAP7_75t_L g1438 ( 
.A1(n_1371),
.A2(n_44),
.B1(n_46),
.B2(n_47),
.Y(n_1438)
);

CKINVDCx5p33_ASAP7_75t_R g1439 ( 
.A(n_1366),
.Y(n_1439)
);

INVxp67_ASAP7_75t_SL g1440 ( 
.A(n_1221),
.Y(n_1440)
);

AO31x2_ASAP7_75t_L g1441 ( 
.A1(n_1373),
.A2(n_664),
.A3(n_50),
.B(n_51),
.Y(n_1441)
);

OAI21x1_ASAP7_75t_L g1442 ( 
.A1(n_1259),
.A2(n_666),
.B(n_662),
.Y(n_1442)
);

AND2x2_ASAP7_75t_L g1443 ( 
.A(n_1319),
.B(n_48),
.Y(n_1443)
);

BUFx6f_ASAP7_75t_L g1444 ( 
.A(n_1291),
.Y(n_1444)
);

NAND2xp5_ASAP7_75t_L g1445 ( 
.A(n_1383),
.B(n_48),
.Y(n_1445)
);

A2O1A1Ixp33_ASAP7_75t_L g1446 ( 
.A1(n_1344),
.A2(n_666),
.B(n_662),
.C(n_637),
.Y(n_1446)
);

AOI21xp5_ASAP7_75t_L g1447 ( 
.A1(n_1237),
.A2(n_666),
.B(n_662),
.Y(n_1447)
);

AO21x2_ASAP7_75t_L g1448 ( 
.A1(n_1292),
.A2(n_123),
.B(n_130),
.Y(n_1448)
);

INVx1_ASAP7_75t_L g1449 ( 
.A(n_1335),
.Y(n_1449)
);

CKINVDCx5p33_ASAP7_75t_R g1450 ( 
.A(n_1238),
.Y(n_1450)
);

O2A1O1Ixp33_ASAP7_75t_SL g1451 ( 
.A1(n_1308),
.A2(n_1311),
.B(n_1244),
.C(n_1373),
.Y(n_1451)
);

AND2x2_ASAP7_75t_L g1452 ( 
.A(n_1339),
.B(n_52),
.Y(n_1452)
);

AOI221xp5_ASAP7_75t_L g1453 ( 
.A1(n_1280),
.A2(n_666),
.B1(n_662),
.B2(n_637),
.C(n_626),
.Y(n_1453)
);

O2A1O1Ixp33_ASAP7_75t_L g1454 ( 
.A1(n_1325),
.A2(n_53),
.B(n_54),
.C(n_55),
.Y(n_1454)
);

O2A1O1Ixp33_ASAP7_75t_L g1455 ( 
.A1(n_1289),
.A2(n_53),
.B(n_56),
.C(n_57),
.Y(n_1455)
);

AOI221xp5_ASAP7_75t_SL g1456 ( 
.A1(n_1311),
.A2(n_666),
.B1(n_662),
.B2(n_637),
.C(n_626),
.Y(n_1456)
);

AO31x2_ASAP7_75t_L g1457 ( 
.A1(n_1255),
.A2(n_1307),
.A3(n_1369),
.B(n_1376),
.Y(n_1457)
);

NOR2xp33_ASAP7_75t_L g1458 ( 
.A(n_1221),
.B(n_58),
.Y(n_1458)
);

INVx1_ASAP7_75t_L g1459 ( 
.A(n_1352),
.Y(n_1459)
);

AOI21xp5_ASAP7_75t_L g1460 ( 
.A1(n_1320),
.A2(n_624),
.B(n_637),
.Y(n_1460)
);

OAI21x1_ASAP7_75t_L g1461 ( 
.A1(n_1265),
.A2(n_624),
.B(n_637),
.Y(n_1461)
);

NAND2xp5_ASAP7_75t_SL g1462 ( 
.A(n_1222),
.B(n_624),
.Y(n_1462)
);

OAI21xp5_ASAP7_75t_L g1463 ( 
.A1(n_1315),
.A2(n_664),
.B(n_637),
.Y(n_1463)
);

INVx1_ASAP7_75t_L g1464 ( 
.A(n_1228),
.Y(n_1464)
);

OAI22x1_ASAP7_75t_L g1465 ( 
.A1(n_1273),
.A2(n_58),
.B1(n_59),
.B2(n_61),
.Y(n_1465)
);

AO31x2_ASAP7_75t_L g1466 ( 
.A1(n_1302),
.A2(n_664),
.A3(n_62),
.B(n_63),
.Y(n_1466)
);

AOI21xp5_ASAP7_75t_L g1467 ( 
.A1(n_1374),
.A2(n_624),
.B(n_626),
.Y(n_1467)
);

AOI221x1_ASAP7_75t_L g1468 ( 
.A1(n_1287),
.A2(n_624),
.B1(n_626),
.B2(n_68),
.C(n_69),
.Y(n_1468)
);

NAND3x1_ASAP7_75t_L g1469 ( 
.A(n_1289),
.B(n_59),
.C(n_65),
.Y(n_1469)
);

NAND2xp5_ASAP7_75t_L g1470 ( 
.A(n_1384),
.B(n_71),
.Y(n_1470)
);

AND2x2_ASAP7_75t_L g1471 ( 
.A(n_1285),
.B(n_71),
.Y(n_1471)
);

INVxp67_ASAP7_75t_L g1472 ( 
.A(n_1248),
.Y(n_1472)
);

AO31x2_ASAP7_75t_L g1473 ( 
.A1(n_1370),
.A2(n_664),
.A3(n_74),
.B(n_77),
.Y(n_1473)
);

INVx3_ASAP7_75t_L g1474 ( 
.A(n_1291),
.Y(n_1474)
);

INVx1_ASAP7_75t_L g1475 ( 
.A(n_1232),
.Y(n_1475)
);

NOR2xp33_ASAP7_75t_L g1476 ( 
.A(n_1365),
.B(n_72),
.Y(n_1476)
);

NAND2xp5_ASAP7_75t_L g1477 ( 
.A(n_1374),
.B(n_626),
.Y(n_1477)
);

AO21x2_ASAP7_75t_L g1478 ( 
.A1(n_1357),
.A2(n_1381),
.B(n_1385),
.Y(n_1478)
);

A2O1A1Ixp33_ASAP7_75t_L g1479 ( 
.A1(n_1345),
.A2(n_77),
.B(n_78),
.C(n_80),
.Y(n_1479)
);

OAI21xp5_ASAP7_75t_L g1480 ( 
.A1(n_1381),
.A2(n_664),
.B(n_154),
.Y(n_1480)
);

INVx3_ASAP7_75t_L g1481 ( 
.A(n_1291),
.Y(n_1481)
);

INVx2_ASAP7_75t_L g1482 ( 
.A(n_1229),
.Y(n_1482)
);

BUFx6f_ASAP7_75t_L g1483 ( 
.A(n_1291),
.Y(n_1483)
);

OR2x6_ASAP7_75t_L g1484 ( 
.A(n_1355),
.B(n_153),
.Y(n_1484)
);

INVxp67_ASAP7_75t_L g1485 ( 
.A(n_1359),
.Y(n_1485)
);

INVx1_ASAP7_75t_L g1486 ( 
.A(n_1235),
.Y(n_1486)
);

AOI221xp5_ASAP7_75t_SL g1487 ( 
.A1(n_1380),
.A2(n_80),
.B1(n_84),
.B2(n_85),
.C(n_86),
.Y(n_1487)
);

AOI22xp5_ASAP7_75t_L g1488 ( 
.A1(n_1246),
.A2(n_84),
.B1(n_86),
.B2(n_87),
.Y(n_1488)
);

OAI21x1_ASAP7_75t_L g1489 ( 
.A1(n_1282),
.A2(n_1330),
.B(n_1279),
.Y(n_1489)
);

NAND2xp5_ASAP7_75t_L g1490 ( 
.A(n_1345),
.B(n_93),
.Y(n_1490)
);

BUFx2_ASAP7_75t_L g1491 ( 
.A(n_1338),
.Y(n_1491)
);

OA21x2_ASAP7_75t_L g1492 ( 
.A1(n_1322),
.A2(n_1385),
.B(n_1347),
.Y(n_1492)
);

INVx2_ASAP7_75t_L g1493 ( 
.A(n_1236),
.Y(n_1493)
);

AOI22xp5_ASAP7_75t_L g1494 ( 
.A1(n_1246),
.A2(n_98),
.B1(n_100),
.B2(n_101),
.Y(n_1494)
);

OAI21xp33_ASAP7_75t_L g1495 ( 
.A1(n_1360),
.A2(n_103),
.B(n_106),
.Y(n_1495)
);

AOI21xp5_ASAP7_75t_L g1496 ( 
.A1(n_1382),
.A2(n_109),
.B(n_115),
.Y(n_1496)
);

NOR2xp67_ASAP7_75t_L g1497 ( 
.A(n_1296),
.B(n_120),
.Y(n_1497)
);

INVx5_ASAP7_75t_L g1498 ( 
.A(n_1306),
.Y(n_1498)
);

CKINVDCx16_ASAP7_75t_R g1499 ( 
.A(n_1238),
.Y(n_1499)
);

INVx1_ASAP7_75t_L g1500 ( 
.A(n_1256),
.Y(n_1500)
);

AO31x2_ASAP7_75t_L g1501 ( 
.A1(n_1370),
.A2(n_125),
.A3(n_136),
.B(n_139),
.Y(n_1501)
);

BUFx2_ASAP7_75t_L g1502 ( 
.A(n_1260),
.Y(n_1502)
);

AOI21xp5_ASAP7_75t_L g1503 ( 
.A1(n_1357),
.A2(n_140),
.B(n_141),
.Y(n_1503)
);

AOI21xp5_ASAP7_75t_SL g1504 ( 
.A1(n_1306),
.A2(n_157),
.B(n_161),
.Y(n_1504)
);

O2A1O1Ixp5_ASAP7_75t_SL g1505 ( 
.A1(n_1332),
.A2(n_1333),
.B(n_1342),
.C(n_1293),
.Y(n_1505)
);

HB1xp67_ASAP7_75t_L g1506 ( 
.A(n_1226),
.Y(n_1506)
);

OAI21xp5_ASAP7_75t_L g1507 ( 
.A1(n_1337),
.A2(n_162),
.B(n_163),
.Y(n_1507)
);

OAI21x1_ASAP7_75t_L g1508 ( 
.A1(n_1361),
.A2(n_165),
.B(n_166),
.Y(n_1508)
);

OAI22x1_ASAP7_75t_L g1509 ( 
.A1(n_1360),
.A2(n_170),
.B1(n_172),
.B2(n_174),
.Y(n_1509)
);

NAND2xp5_ASAP7_75t_L g1510 ( 
.A(n_1375),
.B(n_181),
.Y(n_1510)
);

BUFx3_ASAP7_75t_L g1511 ( 
.A(n_1260),
.Y(n_1511)
);

OAI21x1_ASAP7_75t_L g1512 ( 
.A1(n_1245),
.A2(n_185),
.B(n_194),
.Y(n_1512)
);

OAI22xp5_ASAP7_75t_L g1513 ( 
.A1(n_1371),
.A2(n_197),
.B1(n_198),
.B2(n_199),
.Y(n_1513)
);

AOI21xp5_ASAP7_75t_L g1514 ( 
.A1(n_1297),
.A2(n_202),
.B(n_215),
.Y(n_1514)
);

AOI21xp5_ASAP7_75t_L g1515 ( 
.A1(n_1297),
.A2(n_1327),
.B(n_1314),
.Y(n_1515)
);

BUFx2_ASAP7_75t_L g1516 ( 
.A(n_1267),
.Y(n_1516)
);

AO31x2_ASAP7_75t_L g1517 ( 
.A1(n_1336),
.A2(n_222),
.A3(n_1350),
.B(n_1353),
.Y(n_1517)
);

INVx3_ASAP7_75t_SL g1518 ( 
.A(n_1372),
.Y(n_1518)
);

AOI211x1_ASAP7_75t_L g1519 ( 
.A1(n_1305),
.A2(n_1342),
.B(n_1332),
.C(n_1333),
.Y(n_1519)
);

NAND2xp5_ASAP7_75t_L g1520 ( 
.A(n_1375),
.B(n_1294),
.Y(n_1520)
);

AO31x2_ASAP7_75t_L g1521 ( 
.A1(n_1349),
.A2(n_1354),
.A3(n_1351),
.B(n_1277),
.Y(n_1521)
);

AND2x2_ASAP7_75t_L g1522 ( 
.A(n_1298),
.B(n_1226),
.Y(n_1522)
);

AOI21xp5_ASAP7_75t_L g1523 ( 
.A1(n_1297),
.A2(n_1253),
.B(n_1239),
.Y(n_1523)
);

INVx1_ASAP7_75t_L g1524 ( 
.A(n_1243),
.Y(n_1524)
);

INVx1_ASAP7_75t_L g1525 ( 
.A(n_1251),
.Y(n_1525)
);

AOI21xp5_ASAP7_75t_L g1526 ( 
.A1(n_1297),
.A2(n_1239),
.B(n_1362),
.Y(n_1526)
);

AOI21xp5_ASAP7_75t_L g1527 ( 
.A1(n_1362),
.A2(n_1363),
.B(n_1269),
.Y(n_1527)
);

AOI21xp5_ASAP7_75t_L g1528 ( 
.A1(n_1363),
.A2(n_1272),
.B(n_1247),
.Y(n_1528)
);

AOI22xp5_ASAP7_75t_L g1529 ( 
.A1(n_1298),
.A2(n_1290),
.B1(n_1276),
.B2(n_1324),
.Y(n_1529)
);

AOI21xp5_ASAP7_75t_L g1530 ( 
.A1(n_1247),
.A2(n_1288),
.B(n_1262),
.Y(n_1530)
);

NOR2xp67_ASAP7_75t_SL g1531 ( 
.A(n_1372),
.B(n_1267),
.Y(n_1531)
);

NOR2xp33_ASAP7_75t_L g1532 ( 
.A(n_1317),
.B(n_1304),
.Y(n_1532)
);

INVx1_ASAP7_75t_L g1533 ( 
.A(n_1268),
.Y(n_1533)
);

OAI22xp5_ASAP7_75t_SL g1534 ( 
.A1(n_1324),
.A2(n_1275),
.B1(n_1301),
.B2(n_1368),
.Y(n_1534)
);

O2A1O1Ixp33_ASAP7_75t_SL g1535 ( 
.A1(n_1379),
.A2(n_1341),
.B(n_1340),
.C(n_1329),
.Y(n_1535)
);

AOI21xp5_ASAP7_75t_L g1536 ( 
.A1(n_1377),
.A2(n_1358),
.B(n_1364),
.Y(n_1536)
);

O2A1O1Ixp33_ASAP7_75t_SL g1537 ( 
.A1(n_1331),
.A2(n_1326),
.B(n_1278),
.C(n_1348),
.Y(n_1537)
);

A2O1A1Ixp33_ASAP7_75t_L g1538 ( 
.A1(n_1377),
.A2(n_1233),
.B(n_1278),
.C(n_1348),
.Y(n_1538)
);

AOI221xp5_ASAP7_75t_L g1539 ( 
.A1(n_1368),
.A2(n_1358),
.B1(n_1309),
.B2(n_1346),
.C(n_1356),
.Y(n_1539)
);

INVx1_ASAP7_75t_L g1540 ( 
.A(n_1309),
.Y(n_1540)
);

NOR2xp33_ASAP7_75t_L g1541 ( 
.A(n_1324),
.B(n_1346),
.Y(n_1541)
);

AOI221xp5_ASAP7_75t_SL g1542 ( 
.A1(n_1306),
.A2(n_1095),
.B1(n_1242),
.B2(n_1344),
.C(n_1308),
.Y(n_1542)
);

OAI21x1_ASAP7_75t_L g1543 ( 
.A1(n_1356),
.A2(n_1323),
.B(n_1283),
.Y(n_1543)
);

AOI22xp5_ASAP7_75t_L g1544 ( 
.A1(n_1356),
.A2(n_901),
.B1(n_1070),
.B2(n_1200),
.Y(n_1544)
);

OR2x2_ASAP7_75t_L g1545 ( 
.A(n_1356),
.B(n_1240),
.Y(n_1545)
);

OAI21xp5_ASAP7_75t_L g1546 ( 
.A1(n_1230),
.A2(n_1266),
.B(n_1115),
.Y(n_1546)
);

BUFx6f_ASAP7_75t_L g1547 ( 
.A(n_1291),
.Y(n_1547)
);

NAND2x1p5_ASAP7_75t_L g1548 ( 
.A(n_1297),
.B(n_900),
.Y(n_1548)
);

NAND2xp5_ASAP7_75t_L g1549 ( 
.A(n_1254),
.B(n_857),
.Y(n_1549)
);

AOI22xp33_ASAP7_75t_L g1550 ( 
.A1(n_1271),
.A2(n_1200),
.B1(n_1043),
.B2(n_1157),
.Y(n_1550)
);

AOI21xp5_ASAP7_75t_L g1551 ( 
.A1(n_1227),
.A2(n_929),
.B(n_928),
.Y(n_1551)
);

OAI21xp5_ASAP7_75t_L g1552 ( 
.A1(n_1230),
.A2(n_1266),
.B(n_1115),
.Y(n_1552)
);

OAI22x1_ASAP7_75t_L g1553 ( 
.A1(n_1271),
.A2(n_1334),
.B1(n_1041),
.B2(n_1273),
.Y(n_1553)
);

AOI21xp5_ASAP7_75t_L g1554 ( 
.A1(n_1227),
.A2(n_929),
.B(n_928),
.Y(n_1554)
);

NOR2xp67_ASAP7_75t_L g1555 ( 
.A(n_1240),
.B(n_1188),
.Y(n_1555)
);

INVx1_ASAP7_75t_SL g1556 ( 
.A(n_1270),
.Y(n_1556)
);

NAND2xp5_ASAP7_75t_SL g1557 ( 
.A(n_1264),
.B(n_1214),
.Y(n_1557)
);

A2O1A1Ixp33_ASAP7_75t_L g1558 ( 
.A1(n_1230),
.A2(n_1200),
.B(n_1225),
.C(n_909),
.Y(n_1558)
);

AOI22xp5_ASAP7_75t_L g1559 ( 
.A1(n_1271),
.A2(n_901),
.B1(n_1070),
.B2(n_1200),
.Y(n_1559)
);

OAI21xp5_ASAP7_75t_L g1560 ( 
.A1(n_1230),
.A2(n_1266),
.B(n_1115),
.Y(n_1560)
);

BUFx8_ASAP7_75t_L g1561 ( 
.A(n_1310),
.Y(n_1561)
);

INVx1_ASAP7_75t_SL g1562 ( 
.A(n_1270),
.Y(n_1562)
);

OR2x6_ASAP7_75t_L g1563 ( 
.A(n_1355),
.B(n_900),
.Y(n_1563)
);

NAND2xp5_ASAP7_75t_L g1564 ( 
.A(n_1549),
.B(n_1410),
.Y(n_1564)
);

AOI22xp33_ASAP7_75t_L g1565 ( 
.A1(n_1550),
.A2(n_1553),
.B1(n_1559),
.B2(n_1490),
.Y(n_1565)
);

OAI22xp33_ASAP7_75t_L g1566 ( 
.A1(n_1438),
.A2(n_1488),
.B1(n_1544),
.B2(n_1513),
.Y(n_1566)
);

CKINVDCx11_ASAP7_75t_R g1567 ( 
.A(n_1518),
.Y(n_1567)
);

NAND2x1p5_ASAP7_75t_L g1568 ( 
.A(n_1498),
.B(n_1531),
.Y(n_1568)
);

CKINVDCx6p67_ASAP7_75t_R g1569 ( 
.A(n_1499),
.Y(n_1569)
);

NAND2xp5_ASAP7_75t_L g1570 ( 
.A(n_1413),
.B(n_1416),
.Y(n_1570)
);

INVx6_ASAP7_75t_L g1571 ( 
.A(n_1426),
.Y(n_1571)
);

AOI22xp33_ASAP7_75t_L g1572 ( 
.A1(n_1438),
.A2(n_1465),
.B1(n_1513),
.B2(n_1495),
.Y(n_1572)
);

BUFx6f_ASAP7_75t_L g1573 ( 
.A(n_1498),
.Y(n_1573)
);

CKINVDCx5p33_ASAP7_75t_R g1574 ( 
.A(n_1439),
.Y(n_1574)
);

OAI22xp5_ASAP7_75t_L g1575 ( 
.A1(n_1415),
.A2(n_1555),
.B1(n_1558),
.B2(n_1557),
.Y(n_1575)
);

INVx1_ASAP7_75t_L g1576 ( 
.A(n_1406),
.Y(n_1576)
);

AOI22xp33_ASAP7_75t_L g1577 ( 
.A1(n_1546),
.A2(n_1552),
.B1(n_1560),
.B2(n_1476),
.Y(n_1577)
);

BUFx2_ASAP7_75t_L g1578 ( 
.A(n_1491),
.Y(n_1578)
);

AOI22xp33_ASAP7_75t_L g1579 ( 
.A1(n_1546),
.A2(n_1552),
.B1(n_1560),
.B2(n_1443),
.Y(n_1579)
);

AND2x2_ASAP7_75t_L g1580 ( 
.A(n_1452),
.B(n_1471),
.Y(n_1580)
);

INVx2_ASAP7_75t_SL g1581 ( 
.A(n_1426),
.Y(n_1581)
);

BUFx12f_ASAP7_75t_L g1582 ( 
.A(n_1561),
.Y(n_1582)
);

OAI22xp33_ASAP7_75t_L g1583 ( 
.A1(n_1468),
.A2(n_1484),
.B1(n_1432),
.B2(n_1470),
.Y(n_1583)
);

NAND2xp5_ASAP7_75t_L g1584 ( 
.A(n_1420),
.B(n_1425),
.Y(n_1584)
);

HB1xp67_ASAP7_75t_SL g1585 ( 
.A(n_1561),
.Y(n_1585)
);

CKINVDCx20_ASAP7_75t_R g1586 ( 
.A(n_1450),
.Y(n_1586)
);

OAI22xp5_ASAP7_75t_L g1587 ( 
.A1(n_1563),
.A2(n_1407),
.B1(n_1556),
.B2(n_1562),
.Y(n_1587)
);

OAI22x1_ASAP7_75t_L g1588 ( 
.A1(n_1529),
.A2(n_1440),
.B1(n_1494),
.B2(n_1400),
.Y(n_1588)
);

INVx2_ASAP7_75t_SL g1589 ( 
.A(n_1511),
.Y(n_1589)
);

INVx1_ASAP7_75t_L g1590 ( 
.A(n_1408),
.Y(n_1590)
);

BUFx8_ASAP7_75t_L g1591 ( 
.A(n_1502),
.Y(n_1591)
);

OAI21xp5_ASAP7_75t_L g1592 ( 
.A1(n_1505),
.A2(n_1409),
.B(n_1428),
.Y(n_1592)
);

NAND2xp5_ASAP7_75t_L g1593 ( 
.A(n_1419),
.B(n_1412),
.Y(n_1593)
);

INVx2_ASAP7_75t_SL g1594 ( 
.A(n_1516),
.Y(n_1594)
);

INVx1_ASAP7_75t_L g1595 ( 
.A(n_1429),
.Y(n_1595)
);

INVx8_ASAP7_75t_L g1596 ( 
.A(n_1563),
.Y(n_1596)
);

OAI21xp5_ASAP7_75t_SL g1597 ( 
.A1(n_1454),
.A2(n_1455),
.B(n_1479),
.Y(n_1597)
);

INVx1_ASAP7_75t_L g1598 ( 
.A(n_1449),
.Y(n_1598)
);

INVx1_ASAP7_75t_L g1599 ( 
.A(n_1459),
.Y(n_1599)
);

AOI22xp5_ASAP7_75t_L g1600 ( 
.A1(n_1522),
.A2(n_1402),
.B1(n_1484),
.B2(n_1497),
.Y(n_1600)
);

BUFx2_ASAP7_75t_L g1601 ( 
.A(n_1403),
.Y(n_1601)
);

BUFx3_ASAP7_75t_L g1602 ( 
.A(n_1405),
.Y(n_1602)
);

BUFx2_ASAP7_75t_L g1603 ( 
.A(n_1398),
.Y(n_1603)
);

AOI22xp33_ASAP7_75t_SL g1604 ( 
.A1(n_1437),
.A2(n_1458),
.B1(n_1534),
.B2(n_1402),
.Y(n_1604)
);

BUFx6f_ASAP7_75t_SL g1605 ( 
.A(n_1484),
.Y(n_1605)
);

AOI22xp33_ASAP7_75t_L g1606 ( 
.A1(n_1509),
.A2(n_1445),
.B1(n_1520),
.B2(n_1507),
.Y(n_1606)
);

AOI22xp33_ASAP7_75t_L g1607 ( 
.A1(n_1507),
.A2(n_1532),
.B1(n_1510),
.B2(n_1422),
.Y(n_1607)
);

INVx6_ASAP7_75t_L g1608 ( 
.A(n_1444),
.Y(n_1608)
);

INVx2_ASAP7_75t_L g1609 ( 
.A(n_1482),
.Y(n_1609)
);

INVx1_ASAP7_75t_L g1610 ( 
.A(n_1524),
.Y(n_1610)
);

OAI22xp5_ASAP7_75t_L g1611 ( 
.A1(n_1563),
.A2(n_1562),
.B1(n_1556),
.B2(n_1545),
.Y(n_1611)
);

INVx6_ASAP7_75t_L g1612 ( 
.A(n_1483),
.Y(n_1612)
);

BUFx4f_ASAP7_75t_SL g1613 ( 
.A(n_1405),
.Y(n_1613)
);

INVx1_ASAP7_75t_L g1614 ( 
.A(n_1525),
.Y(n_1614)
);

CKINVDCx20_ASAP7_75t_R g1615 ( 
.A(n_1391),
.Y(n_1615)
);

INVx2_ASAP7_75t_L g1616 ( 
.A(n_1493),
.Y(n_1616)
);

INVx1_ASAP7_75t_L g1617 ( 
.A(n_1533),
.Y(n_1617)
);

AOI22xp33_ASAP7_75t_SL g1618 ( 
.A1(n_1469),
.A2(n_1480),
.B1(n_1430),
.B2(n_1487),
.Y(n_1618)
);

OAI22xp33_ASAP7_75t_L g1619 ( 
.A1(n_1436),
.A2(n_1480),
.B1(n_1464),
.B2(n_1475),
.Y(n_1619)
);

AOI22xp33_ASAP7_75t_L g1620 ( 
.A1(n_1422),
.A2(n_1418),
.B1(n_1500),
.B2(n_1486),
.Y(n_1620)
);

OAI22xp5_ASAP7_75t_L g1621 ( 
.A1(n_1485),
.A2(n_1538),
.B1(n_1446),
.B2(n_1519),
.Y(n_1621)
);

OAI22xp5_ASAP7_75t_L g1622 ( 
.A1(n_1472),
.A2(n_1506),
.B1(n_1539),
.B2(n_1541),
.Y(n_1622)
);

INVx1_ASAP7_75t_SL g1623 ( 
.A(n_1540),
.Y(n_1623)
);

CKINVDCx11_ASAP7_75t_R g1624 ( 
.A(n_1483),
.Y(n_1624)
);

AOI22xp33_ASAP7_75t_L g1625 ( 
.A1(n_1418),
.A2(n_1448),
.B1(n_1423),
.B2(n_1487),
.Y(n_1625)
);

CKINVDCx6p67_ASAP7_75t_R g1626 ( 
.A(n_1483),
.Y(n_1626)
);

AOI22xp33_ASAP7_75t_SL g1627 ( 
.A1(n_1542),
.A2(n_1536),
.B1(n_1451),
.B2(n_1448),
.Y(n_1627)
);

INVx1_ASAP7_75t_L g1628 ( 
.A(n_1474),
.Y(n_1628)
);

OAI22xp33_ASAP7_75t_L g1629 ( 
.A1(n_1542),
.A2(n_1477),
.B1(n_1404),
.B2(n_1514),
.Y(n_1629)
);

BUFx2_ASAP7_75t_L g1630 ( 
.A(n_1481),
.Y(n_1630)
);

OAI21xp5_ASAP7_75t_SL g1631 ( 
.A1(n_1496),
.A2(n_1554),
.B(n_1551),
.Y(n_1631)
);

BUFx6f_ASAP7_75t_L g1632 ( 
.A(n_1547),
.Y(n_1632)
);

AOI21xp5_ASAP7_75t_L g1633 ( 
.A1(n_1387),
.A2(n_1414),
.B(n_1389),
.Y(n_1633)
);

AOI22xp33_ASAP7_75t_L g1634 ( 
.A1(n_1414),
.A2(n_1478),
.B1(n_1503),
.B2(n_1523),
.Y(n_1634)
);

OAI22xp5_ASAP7_75t_L g1635 ( 
.A1(n_1548),
.A2(n_1515),
.B1(n_1528),
.B2(n_1462),
.Y(n_1635)
);

INVx2_ASAP7_75t_SL g1636 ( 
.A(n_1548),
.Y(n_1636)
);

INVx4_ASAP7_75t_L g1637 ( 
.A(n_1492),
.Y(n_1637)
);

AND2x2_ASAP7_75t_L g1638 ( 
.A(n_1501),
.B(n_1473),
.Y(n_1638)
);

AOI22xp33_ASAP7_75t_SL g1639 ( 
.A1(n_1399),
.A2(n_1508),
.B1(n_1394),
.B2(n_1441),
.Y(n_1639)
);

BUFx12f_ASAP7_75t_L g1640 ( 
.A(n_1504),
.Y(n_1640)
);

AOI22xp33_ASAP7_75t_SL g1641 ( 
.A1(n_1399),
.A2(n_1441),
.B1(n_1492),
.B2(n_1456),
.Y(n_1641)
);

OAI22xp5_ASAP7_75t_L g1642 ( 
.A1(n_1526),
.A2(n_1433),
.B1(n_1527),
.B2(n_1530),
.Y(n_1642)
);

BUFx2_ASAP7_75t_L g1643 ( 
.A(n_1501),
.Y(n_1643)
);

INVx2_ASAP7_75t_SL g1644 ( 
.A(n_1441),
.Y(n_1644)
);

OAI21xp33_ASAP7_75t_L g1645 ( 
.A1(n_1417),
.A2(n_1477),
.B(n_1453),
.Y(n_1645)
);

INVx1_ASAP7_75t_L g1646 ( 
.A(n_1473),
.Y(n_1646)
);

BUFx10_ASAP7_75t_L g1647 ( 
.A(n_1473),
.Y(n_1647)
);

AOI22xp33_ASAP7_75t_L g1648 ( 
.A1(n_1478),
.A2(n_1395),
.B1(n_1435),
.B2(n_1512),
.Y(n_1648)
);

INVx1_ASAP7_75t_L g1649 ( 
.A(n_1434),
.Y(n_1649)
);

CKINVDCx11_ASAP7_75t_R g1650 ( 
.A(n_1397),
.Y(n_1650)
);

AOI22xp33_ASAP7_75t_L g1651 ( 
.A1(n_1435),
.A2(n_1431),
.B1(n_1463),
.B2(n_1489),
.Y(n_1651)
);

CKINVDCx11_ASAP7_75t_R g1652 ( 
.A(n_1434),
.Y(n_1652)
);

AOI22xp33_ASAP7_75t_L g1653 ( 
.A1(n_1463),
.A2(n_1460),
.B1(n_1467),
.B2(n_1393),
.Y(n_1653)
);

NAND2xp5_ASAP7_75t_L g1654 ( 
.A(n_1457),
.B(n_1386),
.Y(n_1654)
);

BUFx12f_ASAP7_75t_L g1655 ( 
.A(n_1537),
.Y(n_1655)
);

INVx4_ASAP7_75t_L g1656 ( 
.A(n_1427),
.Y(n_1656)
);

AOI22xp33_ASAP7_75t_L g1657 ( 
.A1(n_1424),
.A2(n_1386),
.B1(n_1392),
.B2(n_1447),
.Y(n_1657)
);

BUFx3_ASAP7_75t_L g1658 ( 
.A(n_1457),
.Y(n_1658)
);

AOI22xp33_ASAP7_75t_L g1659 ( 
.A1(n_1386),
.A2(n_1461),
.B1(n_1442),
.B2(n_1543),
.Y(n_1659)
);

OAI22xp5_ASAP7_75t_L g1660 ( 
.A1(n_1535),
.A2(n_1421),
.B1(n_1401),
.B2(n_1456),
.Y(n_1660)
);

BUFx2_ASAP7_75t_L g1661 ( 
.A(n_1466),
.Y(n_1661)
);

AOI22xp33_ASAP7_75t_L g1662 ( 
.A1(n_1466),
.A2(n_1517),
.B1(n_1411),
.B2(n_1521),
.Y(n_1662)
);

AOI22xp33_ASAP7_75t_L g1663 ( 
.A1(n_1517),
.A2(n_1396),
.B1(n_1521),
.B2(n_1550),
.Y(n_1663)
);

INVx1_ASAP7_75t_SL g1664 ( 
.A(n_1517),
.Y(n_1664)
);

OAI22xp5_ASAP7_75t_L g1665 ( 
.A1(n_1396),
.A2(n_1550),
.B1(n_1559),
.B2(n_901),
.Y(n_1665)
);

BUFx12f_ASAP7_75t_L g1666 ( 
.A(n_1561),
.Y(n_1666)
);

INVx4_ASAP7_75t_L g1667 ( 
.A(n_1498),
.Y(n_1667)
);

NAND2x1p5_ASAP7_75t_L g1668 ( 
.A(n_1498),
.B(n_1297),
.Y(n_1668)
);

CKINVDCx6p67_ASAP7_75t_R g1669 ( 
.A(n_1518),
.Y(n_1669)
);

AOI22xp33_ASAP7_75t_SL g1670 ( 
.A1(n_1438),
.A2(n_1070),
.B1(n_1263),
.B2(n_1271),
.Y(n_1670)
);

HB1xp67_ASAP7_75t_SL g1671 ( 
.A(n_1561),
.Y(n_1671)
);

BUFx6f_ASAP7_75t_L g1672 ( 
.A(n_1498),
.Y(n_1672)
);

CKINVDCx20_ASAP7_75t_R g1673 ( 
.A(n_1561),
.Y(n_1673)
);

OAI21xp5_ASAP7_75t_SL g1674 ( 
.A1(n_1550),
.A2(n_1559),
.B(n_1415),
.Y(n_1674)
);

INVx3_ASAP7_75t_L g1675 ( 
.A(n_1444),
.Y(n_1675)
);

INVx8_ASAP7_75t_L g1676 ( 
.A(n_1498),
.Y(n_1676)
);

INVx1_ASAP7_75t_SL g1677 ( 
.A(n_1405),
.Y(n_1677)
);

OAI22xp5_ASAP7_75t_L g1678 ( 
.A1(n_1550),
.A2(n_1559),
.B1(n_901),
.B2(n_1544),
.Y(n_1678)
);

OAI22xp33_ASAP7_75t_L g1679 ( 
.A1(n_1559),
.A2(n_1263),
.B1(n_1438),
.B2(n_683),
.Y(n_1679)
);

AOI22xp33_ASAP7_75t_L g1680 ( 
.A1(n_1550),
.A2(n_1553),
.B1(n_1271),
.B2(n_1559),
.Y(n_1680)
);

INVx1_ASAP7_75t_L g1681 ( 
.A(n_1388),
.Y(n_1681)
);

OAI21xp5_ASAP7_75t_L g1682 ( 
.A1(n_1550),
.A2(n_1200),
.B(n_1415),
.Y(n_1682)
);

INVx6_ASAP7_75t_L g1683 ( 
.A(n_1426),
.Y(n_1683)
);

BUFx3_ASAP7_75t_L g1684 ( 
.A(n_1511),
.Y(n_1684)
);

INVx6_ASAP7_75t_L g1685 ( 
.A(n_1426),
.Y(n_1685)
);

CKINVDCx5p33_ASAP7_75t_R g1686 ( 
.A(n_1439),
.Y(n_1686)
);

AOI22xp33_ASAP7_75t_L g1687 ( 
.A1(n_1550),
.A2(n_1553),
.B1(n_1271),
.B2(n_1559),
.Y(n_1687)
);

CKINVDCx11_ASAP7_75t_R g1688 ( 
.A(n_1518),
.Y(n_1688)
);

BUFx8_ASAP7_75t_SL g1689 ( 
.A(n_1391),
.Y(n_1689)
);

INVx1_ASAP7_75t_L g1690 ( 
.A(n_1388),
.Y(n_1690)
);

AOI22xp33_ASAP7_75t_SL g1691 ( 
.A1(n_1438),
.A2(n_1070),
.B1(n_1263),
.B2(n_1271),
.Y(n_1691)
);

BUFx8_ASAP7_75t_SL g1692 ( 
.A(n_1391),
.Y(n_1692)
);

OAI22xp33_ASAP7_75t_L g1693 ( 
.A1(n_1559),
.A2(n_1263),
.B1(n_1438),
.B2(n_683),
.Y(n_1693)
);

AOI22xp33_ASAP7_75t_L g1694 ( 
.A1(n_1550),
.A2(n_1553),
.B1(n_1271),
.B2(n_1559),
.Y(n_1694)
);

NAND2xp5_ASAP7_75t_L g1695 ( 
.A(n_1549),
.B(n_1410),
.Y(n_1695)
);

AOI22xp33_ASAP7_75t_L g1696 ( 
.A1(n_1550),
.A2(n_1553),
.B1(n_1271),
.B2(n_1559),
.Y(n_1696)
);

OAI22x1_ASAP7_75t_L g1697 ( 
.A1(n_1559),
.A2(n_1544),
.B1(n_1334),
.B2(n_1488),
.Y(n_1697)
);

INVx2_ASAP7_75t_L g1698 ( 
.A(n_1390),
.Y(n_1698)
);

AOI22xp5_ASAP7_75t_L g1699 ( 
.A1(n_1550),
.A2(n_1559),
.B1(n_901),
.B2(n_1070),
.Y(n_1699)
);

INVx6_ASAP7_75t_L g1700 ( 
.A(n_1426),
.Y(n_1700)
);

NAND2xp5_ASAP7_75t_L g1701 ( 
.A(n_1549),
.B(n_1410),
.Y(n_1701)
);

BUFx6f_ASAP7_75t_L g1702 ( 
.A(n_1498),
.Y(n_1702)
);

INVx1_ASAP7_75t_L g1703 ( 
.A(n_1388),
.Y(n_1703)
);

BUFx3_ASAP7_75t_L g1704 ( 
.A(n_1511),
.Y(n_1704)
);

INVx1_ASAP7_75t_L g1705 ( 
.A(n_1388),
.Y(n_1705)
);

OAI22x1_ASAP7_75t_SL g1706 ( 
.A1(n_1391),
.A2(n_1366),
.B1(n_674),
.B2(n_636),
.Y(n_1706)
);

INVx1_ASAP7_75t_L g1707 ( 
.A(n_1388),
.Y(n_1707)
);

BUFx6f_ASAP7_75t_L g1708 ( 
.A(n_1498),
.Y(n_1708)
);

AOI22xp33_ASAP7_75t_L g1709 ( 
.A1(n_1550),
.A2(n_1553),
.B1(n_1271),
.B2(n_1559),
.Y(n_1709)
);

OAI22xp33_ASAP7_75t_L g1710 ( 
.A1(n_1559),
.A2(n_1263),
.B1(n_1438),
.B2(n_683),
.Y(n_1710)
);

AOI22xp33_ASAP7_75t_SL g1711 ( 
.A1(n_1438),
.A2(n_1070),
.B1(n_1263),
.B2(n_1271),
.Y(n_1711)
);

INVx1_ASAP7_75t_L g1712 ( 
.A(n_1388),
.Y(n_1712)
);

AOI22xp33_ASAP7_75t_SL g1713 ( 
.A1(n_1438),
.A2(n_1070),
.B1(n_1263),
.B2(n_1271),
.Y(n_1713)
);

OAI22xp5_ASAP7_75t_L g1714 ( 
.A1(n_1550),
.A2(n_1559),
.B1(n_901),
.B2(n_1544),
.Y(n_1714)
);

INVx1_ASAP7_75t_L g1715 ( 
.A(n_1388),
.Y(n_1715)
);

INVx1_ASAP7_75t_L g1716 ( 
.A(n_1388),
.Y(n_1716)
);

INVx6_ASAP7_75t_L g1717 ( 
.A(n_1426),
.Y(n_1717)
);

INVx1_ASAP7_75t_L g1718 ( 
.A(n_1388),
.Y(n_1718)
);

CKINVDCx20_ASAP7_75t_R g1719 ( 
.A(n_1561),
.Y(n_1719)
);

CKINVDCx6p67_ASAP7_75t_R g1720 ( 
.A(n_1518),
.Y(n_1720)
);

BUFx2_ASAP7_75t_SL g1721 ( 
.A(n_1511),
.Y(n_1721)
);

CKINVDCx11_ASAP7_75t_R g1722 ( 
.A(n_1518),
.Y(n_1722)
);

INVx6_ASAP7_75t_L g1723 ( 
.A(n_1426),
.Y(n_1723)
);

BUFx3_ASAP7_75t_L g1724 ( 
.A(n_1511),
.Y(n_1724)
);

INVx1_ASAP7_75t_L g1725 ( 
.A(n_1388),
.Y(n_1725)
);

AOI22xp5_ASAP7_75t_L g1726 ( 
.A1(n_1550),
.A2(n_1559),
.B1(n_901),
.B2(n_1070),
.Y(n_1726)
);

INVx1_ASAP7_75t_L g1727 ( 
.A(n_1388),
.Y(n_1727)
);

INVx1_ASAP7_75t_L g1728 ( 
.A(n_1388),
.Y(n_1728)
);

BUFx12f_ASAP7_75t_L g1729 ( 
.A(n_1561),
.Y(n_1729)
);

OAI22xp5_ASAP7_75t_L g1730 ( 
.A1(n_1550),
.A2(n_1559),
.B1(n_901),
.B2(n_1544),
.Y(n_1730)
);

AOI22xp33_ASAP7_75t_L g1731 ( 
.A1(n_1550),
.A2(n_1553),
.B1(n_1271),
.B2(n_1559),
.Y(n_1731)
);

INVx2_ASAP7_75t_SL g1732 ( 
.A(n_1426),
.Y(n_1732)
);

CKINVDCx8_ASAP7_75t_R g1733 ( 
.A(n_1721),
.Y(n_1733)
);

NAND2xp5_ASAP7_75t_L g1734 ( 
.A(n_1564),
.B(n_1695),
.Y(n_1734)
);

BUFx3_ASAP7_75t_L g1735 ( 
.A(n_1602),
.Y(n_1735)
);

BUFx6f_ASAP7_75t_L g1736 ( 
.A(n_1655),
.Y(n_1736)
);

AND2x4_ASAP7_75t_L g1737 ( 
.A(n_1658),
.B(n_1644),
.Y(n_1737)
);

HB1xp67_ASAP7_75t_L g1738 ( 
.A(n_1603),
.Y(n_1738)
);

OAI21x1_ASAP7_75t_L g1739 ( 
.A1(n_1633),
.A2(n_1657),
.B(n_1660),
.Y(n_1739)
);

AND2x2_ASAP7_75t_L g1740 ( 
.A(n_1577),
.B(n_1579),
.Y(n_1740)
);

OR2x2_ASAP7_75t_L g1741 ( 
.A(n_1654),
.B(n_1658),
.Y(n_1741)
);

NAND2x1_ASAP7_75t_L g1742 ( 
.A(n_1635),
.B(n_1577),
.Y(n_1742)
);

INVx2_ASAP7_75t_SL g1743 ( 
.A(n_1571),
.Y(n_1743)
);

HB1xp67_ASAP7_75t_L g1744 ( 
.A(n_1602),
.Y(n_1744)
);

CKINVDCx5p33_ASAP7_75t_R g1745 ( 
.A(n_1574),
.Y(n_1745)
);

OR2x6_ASAP7_75t_L g1746 ( 
.A(n_1631),
.B(n_1592),
.Y(n_1746)
);

INVx1_ASAP7_75t_L g1747 ( 
.A(n_1649),
.Y(n_1747)
);

INVx1_ASAP7_75t_L g1748 ( 
.A(n_1646),
.Y(n_1748)
);

OAI21x1_ASAP7_75t_L g1749 ( 
.A1(n_1657),
.A2(n_1648),
.B(n_1653),
.Y(n_1749)
);

BUFx6f_ASAP7_75t_L g1750 ( 
.A(n_1650),
.Y(n_1750)
);

INVx2_ASAP7_75t_L g1751 ( 
.A(n_1637),
.Y(n_1751)
);

BUFx6f_ASAP7_75t_L g1752 ( 
.A(n_1650),
.Y(n_1752)
);

BUFx3_ASAP7_75t_L g1753 ( 
.A(n_1591),
.Y(n_1753)
);

HB1xp67_ASAP7_75t_L g1754 ( 
.A(n_1601),
.Y(n_1754)
);

NAND2xp5_ASAP7_75t_L g1755 ( 
.A(n_1701),
.B(n_1593),
.Y(n_1755)
);

NOR2xp33_ASAP7_75t_L g1756 ( 
.A(n_1613),
.B(n_1674),
.Y(n_1756)
);

CKINVDCx20_ASAP7_75t_R g1757 ( 
.A(n_1586),
.Y(n_1757)
);

AND2x4_ASAP7_75t_L g1758 ( 
.A(n_1698),
.B(n_1638),
.Y(n_1758)
);

INVx1_ASAP7_75t_L g1759 ( 
.A(n_1661),
.Y(n_1759)
);

INVx1_ASAP7_75t_L g1760 ( 
.A(n_1643),
.Y(n_1760)
);

INVx1_ASAP7_75t_L g1761 ( 
.A(n_1647),
.Y(n_1761)
);

BUFx3_ASAP7_75t_L g1762 ( 
.A(n_1591),
.Y(n_1762)
);

AO21x1_ASAP7_75t_SL g1763 ( 
.A1(n_1572),
.A2(n_1625),
.B(n_1682),
.Y(n_1763)
);

INVx1_ASAP7_75t_L g1764 ( 
.A(n_1647),
.Y(n_1764)
);

BUFx2_ASAP7_75t_L g1765 ( 
.A(n_1637),
.Y(n_1765)
);

INVx2_ASAP7_75t_L g1766 ( 
.A(n_1576),
.Y(n_1766)
);

HB1xp67_ASAP7_75t_L g1767 ( 
.A(n_1611),
.Y(n_1767)
);

INVx2_ASAP7_75t_L g1768 ( 
.A(n_1590),
.Y(n_1768)
);

HB1xp67_ASAP7_75t_L g1769 ( 
.A(n_1677),
.Y(n_1769)
);

INVx1_ASAP7_75t_L g1770 ( 
.A(n_1595),
.Y(n_1770)
);

INVx1_ASAP7_75t_L g1771 ( 
.A(n_1598),
.Y(n_1771)
);

INVx1_ASAP7_75t_L g1772 ( 
.A(n_1599),
.Y(n_1772)
);

INVxp67_ASAP7_75t_L g1773 ( 
.A(n_1578),
.Y(n_1773)
);

NAND2xp5_ASAP7_75t_SL g1774 ( 
.A(n_1699),
.B(n_1726),
.Y(n_1774)
);

INVx2_ASAP7_75t_L g1775 ( 
.A(n_1656),
.Y(n_1775)
);

CKINVDCx5p33_ASAP7_75t_R g1776 ( 
.A(n_1686),
.Y(n_1776)
);

AOI221x1_ASAP7_75t_L g1777 ( 
.A1(n_1678),
.A2(n_1714),
.B1(n_1730),
.B2(n_1665),
.C(n_1697),
.Y(n_1777)
);

INVx1_ASAP7_75t_L g1778 ( 
.A(n_1681),
.Y(n_1778)
);

AOI22xp33_ASAP7_75t_L g1779 ( 
.A1(n_1670),
.A2(n_1711),
.B1(n_1691),
.B2(n_1713),
.Y(n_1779)
);

INVx1_ASAP7_75t_L g1780 ( 
.A(n_1690),
.Y(n_1780)
);

INVxp67_ASAP7_75t_SL g1781 ( 
.A(n_1570),
.Y(n_1781)
);

INVx2_ASAP7_75t_L g1782 ( 
.A(n_1703),
.Y(n_1782)
);

OAI21x1_ASAP7_75t_L g1783 ( 
.A1(n_1648),
.A2(n_1653),
.B(n_1659),
.Y(n_1783)
);

HB1xp67_ASAP7_75t_L g1784 ( 
.A(n_1623),
.Y(n_1784)
);

AND2x2_ASAP7_75t_L g1785 ( 
.A(n_1579),
.B(n_1663),
.Y(n_1785)
);

INVx1_ASAP7_75t_L g1786 ( 
.A(n_1705),
.Y(n_1786)
);

INVx1_ASAP7_75t_L g1787 ( 
.A(n_1707),
.Y(n_1787)
);

INVx3_ASAP7_75t_L g1788 ( 
.A(n_1656),
.Y(n_1788)
);

INVx2_ASAP7_75t_SL g1789 ( 
.A(n_1571),
.Y(n_1789)
);

OAI21x1_ASAP7_75t_SL g1790 ( 
.A1(n_1621),
.A2(n_1600),
.B(n_1620),
.Y(n_1790)
);

NOR2xp33_ASAP7_75t_L g1791 ( 
.A(n_1613),
.B(n_1584),
.Y(n_1791)
);

HB1xp67_ASAP7_75t_L g1792 ( 
.A(n_1587),
.Y(n_1792)
);

INVx2_ASAP7_75t_SL g1793 ( 
.A(n_1571),
.Y(n_1793)
);

AOI21x1_ASAP7_75t_L g1794 ( 
.A1(n_1642),
.A2(n_1575),
.B(n_1588),
.Y(n_1794)
);

AO21x2_ASAP7_75t_L g1795 ( 
.A1(n_1619),
.A2(n_1629),
.B(n_1645),
.Y(n_1795)
);

INVx1_ASAP7_75t_L g1796 ( 
.A(n_1712),
.Y(n_1796)
);

INVx1_ASAP7_75t_L g1797 ( 
.A(n_1715),
.Y(n_1797)
);

INVx2_ASAP7_75t_L g1798 ( 
.A(n_1716),
.Y(n_1798)
);

INVx3_ASAP7_75t_L g1799 ( 
.A(n_1664),
.Y(n_1799)
);

A2O1A1Ixp33_ASAP7_75t_L g1800 ( 
.A1(n_1680),
.A2(n_1687),
.B(n_1709),
.C(n_1731),
.Y(n_1800)
);

INVx2_ASAP7_75t_L g1801 ( 
.A(n_1718),
.Y(n_1801)
);

AOI21xp5_ASAP7_75t_L g1802 ( 
.A1(n_1629),
.A2(n_1607),
.B(n_1619),
.Y(n_1802)
);

INVx1_ASAP7_75t_L g1803 ( 
.A(n_1725),
.Y(n_1803)
);

INVx1_ASAP7_75t_SL g1804 ( 
.A(n_1580),
.Y(n_1804)
);

OAI21xp5_ASAP7_75t_L g1805 ( 
.A1(n_1680),
.A2(n_1687),
.B(n_1694),
.Y(n_1805)
);

NAND2xp5_ASAP7_75t_L g1806 ( 
.A(n_1694),
.B(n_1696),
.Y(n_1806)
);

NAND2xp33_ASAP7_75t_L g1807 ( 
.A(n_1696),
.B(n_1709),
.Y(n_1807)
);

INVx1_ASAP7_75t_L g1808 ( 
.A(n_1727),
.Y(n_1808)
);

OAI21x1_ASAP7_75t_L g1809 ( 
.A1(n_1659),
.A2(n_1634),
.B(n_1651),
.Y(n_1809)
);

INVx1_ASAP7_75t_L g1810 ( 
.A(n_1728),
.Y(n_1810)
);

INVx1_ASAP7_75t_L g1811 ( 
.A(n_1610),
.Y(n_1811)
);

CKINVDCx5p33_ASAP7_75t_R g1812 ( 
.A(n_1689),
.Y(n_1812)
);

INVx1_ASAP7_75t_L g1813 ( 
.A(n_1614),
.Y(n_1813)
);

INVx4_ASAP7_75t_SL g1814 ( 
.A(n_1605),
.Y(n_1814)
);

INVx2_ASAP7_75t_L g1815 ( 
.A(n_1617),
.Y(n_1815)
);

INVx1_ASAP7_75t_L g1816 ( 
.A(n_1641),
.Y(n_1816)
);

AND2x2_ASAP7_75t_L g1817 ( 
.A(n_1663),
.B(n_1620),
.Y(n_1817)
);

HB1xp67_ASAP7_75t_L g1818 ( 
.A(n_1630),
.Y(n_1818)
);

HB1xp67_ASAP7_75t_L g1819 ( 
.A(n_1622),
.Y(n_1819)
);

HB1xp67_ASAP7_75t_L g1820 ( 
.A(n_1594),
.Y(n_1820)
);

INVx1_ASAP7_75t_L g1821 ( 
.A(n_1641),
.Y(n_1821)
);

AO21x2_ASAP7_75t_L g1822 ( 
.A1(n_1566),
.A2(n_1693),
.B(n_1679),
.Y(n_1822)
);

AND2x2_ASAP7_75t_L g1823 ( 
.A(n_1652),
.B(n_1565),
.Y(n_1823)
);

INVx1_ASAP7_75t_L g1824 ( 
.A(n_1662),
.Y(n_1824)
);

AOI221xp5_ASAP7_75t_L g1825 ( 
.A1(n_1679),
.A2(n_1693),
.B1(n_1710),
.B2(n_1566),
.C(n_1731),
.Y(n_1825)
);

BUFx6f_ASAP7_75t_L g1826 ( 
.A(n_1652),
.Y(n_1826)
);

INVx3_ASAP7_75t_L g1827 ( 
.A(n_1596),
.Y(n_1827)
);

INVx1_ASAP7_75t_L g1828 ( 
.A(n_1662),
.Y(n_1828)
);

HB1xp67_ASAP7_75t_L g1829 ( 
.A(n_1628),
.Y(n_1829)
);

INVx1_ASAP7_75t_L g1830 ( 
.A(n_1609),
.Y(n_1830)
);

INVx1_ASAP7_75t_L g1831 ( 
.A(n_1616),
.Y(n_1831)
);

AO32x2_ASAP7_75t_L g1832 ( 
.A1(n_1636),
.A2(n_1639),
.A3(n_1627),
.B1(n_1711),
.B2(n_1713),
.Y(n_1832)
);

INVx1_ASAP7_75t_L g1833 ( 
.A(n_1639),
.Y(n_1833)
);

BUFx2_ASAP7_75t_L g1834 ( 
.A(n_1568),
.Y(n_1834)
);

AO21x2_ASAP7_75t_L g1835 ( 
.A1(n_1710),
.A2(n_1583),
.B(n_1597),
.Y(n_1835)
);

INVx2_ASAP7_75t_L g1836 ( 
.A(n_1573),
.Y(n_1836)
);

INVx2_ASAP7_75t_L g1837 ( 
.A(n_1573),
.Y(n_1837)
);

OR2x2_ASAP7_75t_L g1838 ( 
.A(n_1565),
.B(n_1625),
.Y(n_1838)
);

INVx2_ASAP7_75t_SL g1839 ( 
.A(n_1683),
.Y(n_1839)
);

INVx1_ASAP7_75t_L g1840 ( 
.A(n_1627),
.Y(n_1840)
);

INVx1_ASAP7_75t_L g1841 ( 
.A(n_1634),
.Y(n_1841)
);

INVx1_ASAP7_75t_L g1842 ( 
.A(n_1651),
.Y(n_1842)
);

INVx1_ASAP7_75t_L g1843 ( 
.A(n_1607),
.Y(n_1843)
);

OAI21x1_ASAP7_75t_L g1844 ( 
.A1(n_1606),
.A2(n_1572),
.B(n_1668),
.Y(n_1844)
);

INVx1_ASAP7_75t_L g1845 ( 
.A(n_1583),
.Y(n_1845)
);

INVx2_ASAP7_75t_SL g1846 ( 
.A(n_1683),
.Y(n_1846)
);

BUFx4f_ASAP7_75t_SL g1847 ( 
.A(n_1582),
.Y(n_1847)
);

AOI22xp33_ASAP7_75t_L g1848 ( 
.A1(n_1670),
.A2(n_1691),
.B1(n_1604),
.B2(n_1618),
.Y(n_1848)
);

INVx1_ASAP7_75t_L g1849 ( 
.A(n_1606),
.Y(n_1849)
);

OA21x2_ASAP7_75t_L g1850 ( 
.A1(n_1618),
.A2(n_1604),
.B(n_1732),
.Y(n_1850)
);

BUFx6f_ASAP7_75t_L g1851 ( 
.A(n_1596),
.Y(n_1851)
);

INVx2_ASAP7_75t_L g1852 ( 
.A(n_1672),
.Y(n_1852)
);

INVx1_ASAP7_75t_L g1853 ( 
.A(n_1702),
.Y(n_1853)
);

INVx3_ASAP7_75t_L g1854 ( 
.A(n_1596),
.Y(n_1854)
);

BUFx3_ASAP7_75t_L g1855 ( 
.A(n_1676),
.Y(n_1855)
);

NAND2xp5_ASAP7_75t_L g1856 ( 
.A(n_1589),
.B(n_1704),
.Y(n_1856)
);

INVx1_ASAP7_75t_L g1857 ( 
.A(n_1708),
.Y(n_1857)
);

INVx3_ASAP7_75t_L g1858 ( 
.A(n_1640),
.Y(n_1858)
);

BUFx2_ASAP7_75t_L g1859 ( 
.A(n_1632),
.Y(n_1859)
);

INVx1_ASAP7_75t_L g1860 ( 
.A(n_1708),
.Y(n_1860)
);

NAND2xp5_ASAP7_75t_L g1861 ( 
.A(n_1684),
.B(n_1704),
.Y(n_1861)
);

INVx3_ASAP7_75t_L g1862 ( 
.A(n_1667),
.Y(n_1862)
);

INVx3_ASAP7_75t_L g1863 ( 
.A(n_1676),
.Y(n_1863)
);

INVx1_ASAP7_75t_L g1864 ( 
.A(n_1675),
.Y(n_1864)
);

AND2x2_ASAP7_75t_L g1865 ( 
.A(n_1626),
.B(n_1608),
.Y(n_1865)
);

AOI221xp5_ASAP7_75t_L g1866 ( 
.A1(n_1825),
.A2(n_1706),
.B1(n_1684),
.B2(n_1724),
.C(n_1581),
.Y(n_1866)
);

AND2x4_ASAP7_75t_L g1867 ( 
.A(n_1758),
.B(n_1724),
.Y(n_1867)
);

AND2x2_ASAP7_75t_L g1868 ( 
.A(n_1735),
.B(n_1569),
.Y(n_1868)
);

OR2x2_ASAP7_75t_L g1869 ( 
.A(n_1767),
.B(n_1669),
.Y(n_1869)
);

BUFx8_ASAP7_75t_L g1870 ( 
.A(n_1753),
.Y(n_1870)
);

AND2x2_ASAP7_75t_L g1871 ( 
.A(n_1735),
.B(n_1624),
.Y(n_1871)
);

AOI221xp5_ASAP7_75t_L g1872 ( 
.A1(n_1807),
.A2(n_1673),
.B1(n_1719),
.B2(n_1676),
.C(n_1615),
.Y(n_1872)
);

BUFx3_ASAP7_75t_L g1873 ( 
.A(n_1861),
.Y(n_1873)
);

NAND2xp5_ASAP7_75t_L g1874 ( 
.A(n_1781),
.B(n_1700),
.Y(n_1874)
);

AND2x2_ASAP7_75t_L g1875 ( 
.A(n_1735),
.B(n_1744),
.Y(n_1875)
);

NOR2xp33_ASAP7_75t_L g1876 ( 
.A(n_1791),
.B(n_1567),
.Y(n_1876)
);

AND2x2_ASAP7_75t_L g1877 ( 
.A(n_1792),
.B(n_1624),
.Y(n_1877)
);

INVx4_ASAP7_75t_L g1878 ( 
.A(n_1858),
.Y(n_1878)
);

AND2x2_ASAP7_75t_L g1879 ( 
.A(n_1823),
.B(n_1612),
.Y(n_1879)
);

BUFx2_ASAP7_75t_L g1880 ( 
.A(n_1859),
.Y(n_1880)
);

OAI22xp5_ASAP7_75t_L g1881 ( 
.A1(n_1848),
.A2(n_1671),
.B1(n_1585),
.B2(n_1700),
.Y(n_1881)
);

AND2x4_ASAP7_75t_L g1882 ( 
.A(n_1758),
.B(n_1720),
.Y(n_1882)
);

INVxp33_ASAP7_75t_L g1883 ( 
.A(n_1769),
.Y(n_1883)
);

AND2x2_ASAP7_75t_L g1884 ( 
.A(n_1823),
.B(n_1612),
.Y(n_1884)
);

AND2x2_ASAP7_75t_L g1885 ( 
.A(n_1804),
.B(n_1612),
.Y(n_1885)
);

CKINVDCx20_ASAP7_75t_R g1886 ( 
.A(n_1757),
.Y(n_1886)
);

A2O1A1Ixp33_ASAP7_75t_L g1887 ( 
.A1(n_1800),
.A2(n_1685),
.B(n_1717),
.C(n_1723),
.Y(n_1887)
);

NOR2xp33_ASAP7_75t_L g1888 ( 
.A(n_1734),
.B(n_1567),
.Y(n_1888)
);

INVx1_ASAP7_75t_SL g1889 ( 
.A(n_1784),
.Y(n_1889)
);

AND2x4_ASAP7_75t_L g1890 ( 
.A(n_1758),
.B(n_1688),
.Y(n_1890)
);

BUFx3_ASAP7_75t_L g1891 ( 
.A(n_1753),
.Y(n_1891)
);

OR2x2_ASAP7_75t_L g1892 ( 
.A(n_1741),
.B(n_1722),
.Y(n_1892)
);

INVx1_ASAP7_75t_L g1893 ( 
.A(n_1770),
.Y(n_1893)
);

NAND2xp5_ASAP7_75t_L g1894 ( 
.A(n_1740),
.B(n_1723),
.Y(n_1894)
);

INVxp67_ASAP7_75t_L g1895 ( 
.A(n_1754),
.Y(n_1895)
);

AOI221xp5_ASAP7_75t_L g1896 ( 
.A1(n_1805),
.A2(n_1688),
.B1(n_1722),
.B2(n_1685),
.C(n_1723),
.Y(n_1896)
);

NOR2x1_ASAP7_75t_SL g1897 ( 
.A(n_1826),
.B(n_1666),
.Y(n_1897)
);

O2A1O1Ixp33_ASAP7_75t_L g1898 ( 
.A1(n_1774),
.A2(n_1683),
.B(n_1685),
.C(n_1700),
.Y(n_1898)
);

OAI21x1_ASAP7_75t_L g1899 ( 
.A1(n_1739),
.A2(n_1717),
.B(n_1729),
.Y(n_1899)
);

CKINVDCx5p33_ASAP7_75t_R g1900 ( 
.A(n_1745),
.Y(n_1900)
);

OR2x2_ASAP7_75t_L g1901 ( 
.A(n_1741),
.B(n_1798),
.Y(n_1901)
);

BUFx12f_ASAP7_75t_L g1902 ( 
.A(n_1812),
.Y(n_1902)
);

OR2x2_ASAP7_75t_L g1903 ( 
.A(n_1798),
.B(n_1717),
.Y(n_1903)
);

INVx1_ASAP7_75t_L g1904 ( 
.A(n_1770),
.Y(n_1904)
);

A2O1A1Ixp33_ASAP7_75t_L g1905 ( 
.A1(n_1802),
.A2(n_1689),
.B(n_1692),
.C(n_1779),
.Y(n_1905)
);

AND2x2_ASAP7_75t_L g1906 ( 
.A(n_1826),
.B(n_1692),
.Y(n_1906)
);

INVx1_ASAP7_75t_L g1907 ( 
.A(n_1771),
.Y(n_1907)
);

NOR2xp33_ASAP7_75t_L g1908 ( 
.A(n_1755),
.B(n_1756),
.Y(n_1908)
);

OAI211xp5_ASAP7_75t_L g1909 ( 
.A1(n_1777),
.A2(n_1806),
.B(n_1845),
.C(n_1819),
.Y(n_1909)
);

A2O1A1Ixp33_ASAP7_75t_L g1910 ( 
.A1(n_1742),
.A2(n_1844),
.B(n_1845),
.C(n_1849),
.Y(n_1910)
);

AOI21xp5_ASAP7_75t_L g1911 ( 
.A1(n_1742),
.A2(n_1746),
.B(n_1795),
.Y(n_1911)
);

NAND2xp5_ASAP7_75t_L g1912 ( 
.A(n_1740),
.B(n_1849),
.Y(n_1912)
);

OR2x2_ASAP7_75t_L g1913 ( 
.A(n_1798),
.B(n_1801),
.Y(n_1913)
);

A2O1A1Ixp33_ASAP7_75t_L g1914 ( 
.A1(n_1844),
.A2(n_1838),
.B(n_1843),
.C(n_1785),
.Y(n_1914)
);

AND2x4_ASAP7_75t_L g1915 ( 
.A(n_1758),
.B(n_1814),
.Y(n_1915)
);

AND2x2_ASAP7_75t_L g1916 ( 
.A(n_1826),
.B(n_1738),
.Y(n_1916)
);

AOI22xp33_ASAP7_75t_L g1917 ( 
.A1(n_1822),
.A2(n_1835),
.B1(n_1763),
.B2(n_1790),
.Y(n_1917)
);

NAND2xp5_ASAP7_75t_L g1918 ( 
.A(n_1843),
.B(n_1801),
.Y(n_1918)
);

INVxp67_ASAP7_75t_L g1919 ( 
.A(n_1820),
.Y(n_1919)
);

OR2x6_ASAP7_75t_L g1920 ( 
.A(n_1746),
.B(n_1794),
.Y(n_1920)
);

INVx1_ASAP7_75t_L g1921 ( 
.A(n_1772),
.Y(n_1921)
);

OR2x2_ASAP7_75t_L g1922 ( 
.A(n_1766),
.B(n_1768),
.Y(n_1922)
);

AO21x2_ASAP7_75t_L g1923 ( 
.A1(n_1795),
.A2(n_1790),
.B(n_1775),
.Y(n_1923)
);

HB1xp67_ASAP7_75t_L g1924 ( 
.A(n_1818),
.Y(n_1924)
);

OAI21xp5_ASAP7_75t_L g1925 ( 
.A1(n_1777),
.A2(n_1794),
.B(n_1838),
.Y(n_1925)
);

INVx4_ASAP7_75t_L g1926 ( 
.A(n_1858),
.Y(n_1926)
);

A2O1A1Ixp33_ASAP7_75t_L g1927 ( 
.A1(n_1785),
.A2(n_1809),
.B(n_1817),
.C(n_1840),
.Y(n_1927)
);

AND2x2_ASAP7_75t_L g1928 ( 
.A(n_1782),
.B(n_1822),
.Y(n_1928)
);

A2O1A1Ixp33_ASAP7_75t_L g1929 ( 
.A1(n_1809),
.A2(n_1817),
.B(n_1840),
.C(n_1841),
.Y(n_1929)
);

AND4x1_ASAP7_75t_L g1930 ( 
.A(n_1814),
.B(n_1833),
.C(n_1835),
.D(n_1733),
.Y(n_1930)
);

OAI21xp5_ASAP7_75t_L g1931 ( 
.A1(n_1746),
.A2(n_1841),
.B(n_1850),
.Y(n_1931)
);

O2A1O1Ixp33_ASAP7_75t_SL g1932 ( 
.A1(n_1743),
.A2(n_1793),
.B(n_1846),
.C(n_1839),
.Y(n_1932)
);

AOI22xp5_ASAP7_75t_L g1933 ( 
.A1(n_1835),
.A2(n_1822),
.B1(n_1850),
.B2(n_1795),
.Y(n_1933)
);

AO32x2_ASAP7_75t_L g1934 ( 
.A1(n_1832),
.A2(n_1743),
.A3(n_1846),
.B1(n_1839),
.B2(n_1793),
.Y(n_1934)
);

AND2x2_ASAP7_75t_L g1935 ( 
.A(n_1815),
.B(n_1746),
.Y(n_1935)
);

AND2x2_ASAP7_75t_L g1936 ( 
.A(n_1815),
.B(n_1746),
.Y(n_1936)
);

AOI21xp5_ASAP7_75t_L g1937 ( 
.A1(n_1749),
.A2(n_1783),
.B(n_1833),
.Y(n_1937)
);

AO32x2_ASAP7_75t_L g1938 ( 
.A1(n_1832),
.A2(n_1789),
.A3(n_1816),
.B1(n_1821),
.B2(n_1759),
.Y(n_1938)
);

INVx1_ASAP7_75t_L g1939 ( 
.A(n_1778),
.Y(n_1939)
);

AOI221xp5_ASAP7_75t_L g1940 ( 
.A1(n_1816),
.A2(n_1821),
.B1(n_1842),
.B2(n_1824),
.C(n_1828),
.Y(n_1940)
);

A2O1A1Ixp33_ASAP7_75t_L g1941 ( 
.A1(n_1858),
.A2(n_1783),
.B(n_1752),
.C(n_1750),
.Y(n_1941)
);

INVx1_ASAP7_75t_L g1942 ( 
.A(n_1778),
.Y(n_1942)
);

OR2x6_ASAP7_75t_L g1943 ( 
.A(n_1750),
.B(n_1752),
.Y(n_1943)
);

NAND4xp25_ASAP7_75t_L g1944 ( 
.A(n_1773),
.B(n_1856),
.C(n_1842),
.D(n_1753),
.Y(n_1944)
);

AND2x4_ASAP7_75t_L g1945 ( 
.A(n_1834),
.B(n_1836),
.Y(n_1945)
);

NOR2x1_ASAP7_75t_L g1946 ( 
.A(n_1858),
.B(n_1855),
.Y(n_1946)
);

INVx3_ASAP7_75t_L g1947 ( 
.A(n_1836),
.Y(n_1947)
);

CKINVDCx5p33_ASAP7_75t_R g1948 ( 
.A(n_1776),
.Y(n_1948)
);

A2O1A1Ixp33_ASAP7_75t_L g1949 ( 
.A1(n_1750),
.A2(n_1752),
.B(n_1749),
.C(n_1828),
.Y(n_1949)
);

AND2x4_ASAP7_75t_L g1950 ( 
.A(n_1834),
.B(n_1836),
.Y(n_1950)
);

INVx1_ASAP7_75t_L g1951 ( 
.A(n_1780),
.Y(n_1951)
);

AND2x4_ASAP7_75t_L g1952 ( 
.A(n_1837),
.B(n_1852),
.Y(n_1952)
);

CKINVDCx8_ASAP7_75t_R g1953 ( 
.A(n_1750),
.Y(n_1953)
);

INVx1_ASAP7_75t_L g1954 ( 
.A(n_1786),
.Y(n_1954)
);

AND2x4_ASAP7_75t_L g1955 ( 
.A(n_1837),
.B(n_1852),
.Y(n_1955)
);

BUFx3_ASAP7_75t_L g1956 ( 
.A(n_1762),
.Y(n_1956)
);

NAND2xp5_ASAP7_75t_L g1957 ( 
.A(n_1811),
.B(n_1813),
.Y(n_1957)
);

BUFx6f_ASAP7_75t_L g1958 ( 
.A(n_1733),
.Y(n_1958)
);

AND2x2_ASAP7_75t_L g1959 ( 
.A(n_1787),
.B(n_1796),
.Y(n_1959)
);

OR2x2_ASAP7_75t_L g1960 ( 
.A(n_1797),
.B(n_1803),
.Y(n_1960)
);

NAND2xp5_ASAP7_75t_L g1961 ( 
.A(n_1811),
.B(n_1813),
.Y(n_1961)
);

INVx1_ASAP7_75t_L g1962 ( 
.A(n_1803),
.Y(n_1962)
);

AO21x2_ASAP7_75t_L g1963 ( 
.A1(n_1775),
.A2(n_1764),
.B(n_1761),
.Y(n_1963)
);

A2O1A1Ixp33_ASAP7_75t_L g1964 ( 
.A1(n_1750),
.A2(n_1752),
.B(n_1824),
.C(n_1762),
.Y(n_1964)
);

AND2x2_ASAP7_75t_L g1965 ( 
.A(n_1808),
.B(n_1810),
.Y(n_1965)
);

AO32x2_ASAP7_75t_L g1966 ( 
.A1(n_1832),
.A2(n_1789),
.A3(n_1759),
.B1(n_1775),
.B2(n_1788),
.Y(n_1966)
);

AND2x2_ASAP7_75t_L g1967 ( 
.A(n_1808),
.B(n_1810),
.Y(n_1967)
);

OR2x2_ASAP7_75t_L g1968 ( 
.A(n_1760),
.B(n_1799),
.Y(n_1968)
);

INVx1_ASAP7_75t_L g1969 ( 
.A(n_1893),
.Y(n_1969)
);

INVx1_ASAP7_75t_L g1970 ( 
.A(n_1904),
.Y(n_1970)
);

OR2x2_ASAP7_75t_L g1971 ( 
.A(n_1901),
.B(n_1760),
.Y(n_1971)
);

AND2x2_ASAP7_75t_L g1972 ( 
.A(n_1935),
.B(n_1765),
.Y(n_1972)
);

INVx1_ASAP7_75t_L g1973 ( 
.A(n_1907),
.Y(n_1973)
);

AND2x2_ASAP7_75t_L g1974 ( 
.A(n_1936),
.B(n_1928),
.Y(n_1974)
);

OR2x2_ASAP7_75t_L g1975 ( 
.A(n_1968),
.B(n_1937),
.Y(n_1975)
);

BUFx2_ASAP7_75t_L g1976 ( 
.A(n_1934),
.Y(n_1976)
);

INVx2_ASAP7_75t_L g1977 ( 
.A(n_1913),
.Y(n_1977)
);

AND2x4_ASAP7_75t_L g1978 ( 
.A(n_1945),
.B(n_1737),
.Y(n_1978)
);

INVx1_ASAP7_75t_L g1979 ( 
.A(n_1921),
.Y(n_1979)
);

INVx1_ASAP7_75t_L g1980 ( 
.A(n_1939),
.Y(n_1980)
);

BUFx3_ASAP7_75t_L g1981 ( 
.A(n_1870),
.Y(n_1981)
);

AND2x2_ASAP7_75t_L g1982 ( 
.A(n_1931),
.B(n_1765),
.Y(n_1982)
);

AND2x2_ASAP7_75t_L g1983 ( 
.A(n_1931),
.B(n_1751),
.Y(n_1983)
);

AND2x2_ASAP7_75t_L g1984 ( 
.A(n_1927),
.B(n_1799),
.Y(n_1984)
);

HB1xp67_ASAP7_75t_L g1985 ( 
.A(n_1889),
.Y(n_1985)
);

INVx1_ASAP7_75t_L g1986 ( 
.A(n_1942),
.Y(n_1986)
);

AOI21xp33_ASAP7_75t_L g1987 ( 
.A1(n_1909),
.A2(n_1925),
.B(n_1908),
.Y(n_1987)
);

NAND2xp5_ASAP7_75t_L g1988 ( 
.A(n_1889),
.B(n_1895),
.Y(n_1988)
);

AOI22xp5_ASAP7_75t_L g1989 ( 
.A1(n_1881),
.A2(n_1850),
.B1(n_1752),
.B2(n_1736),
.Y(n_1989)
);

OR2x2_ASAP7_75t_L g1990 ( 
.A(n_1937),
.B(n_1748),
.Y(n_1990)
);

AND2x2_ASAP7_75t_L g1991 ( 
.A(n_1934),
.B(n_1799),
.Y(n_1991)
);

INVxp67_ASAP7_75t_SL g1992 ( 
.A(n_1924),
.Y(n_1992)
);

AND2x2_ASAP7_75t_L g1993 ( 
.A(n_1934),
.B(n_1799),
.Y(n_1993)
);

AND2x4_ASAP7_75t_L g1994 ( 
.A(n_1945),
.B(n_1950),
.Y(n_1994)
);

NOR2xp33_ASAP7_75t_SL g1995 ( 
.A(n_1902),
.B(n_1847),
.Y(n_1995)
);

HB1xp67_ASAP7_75t_L g1996 ( 
.A(n_1880),
.Y(n_1996)
);

AND2x2_ASAP7_75t_L g1997 ( 
.A(n_1966),
.B(n_1788),
.Y(n_1997)
);

AOI22xp33_ASAP7_75t_L g1998 ( 
.A1(n_1866),
.A2(n_1850),
.B1(n_1762),
.B2(n_1851),
.Y(n_1998)
);

HB1xp67_ASAP7_75t_L g1999 ( 
.A(n_1947),
.Y(n_1999)
);

AOI22xp33_ASAP7_75t_L g2000 ( 
.A1(n_1866),
.A2(n_1851),
.B1(n_1854),
.B2(n_1827),
.Y(n_2000)
);

OR2x2_ASAP7_75t_L g2001 ( 
.A(n_1929),
.B(n_1748),
.Y(n_2001)
);

INVx2_ASAP7_75t_SL g2002 ( 
.A(n_1950),
.Y(n_2002)
);

HB1xp67_ASAP7_75t_L g2003 ( 
.A(n_1918),
.Y(n_2003)
);

AND2x2_ASAP7_75t_L g2004 ( 
.A(n_1966),
.B(n_1788),
.Y(n_2004)
);

INVx1_ASAP7_75t_L g2005 ( 
.A(n_1951),
.Y(n_2005)
);

HB1xp67_ASAP7_75t_L g2006 ( 
.A(n_1918),
.Y(n_2006)
);

AOI22xp33_ASAP7_75t_SL g2007 ( 
.A1(n_1881),
.A2(n_1832),
.B1(n_1736),
.B2(n_1851),
.Y(n_2007)
);

INVx1_ASAP7_75t_L g2008 ( 
.A(n_1954),
.Y(n_2008)
);

AND2x4_ASAP7_75t_L g2009 ( 
.A(n_1915),
.B(n_1737),
.Y(n_2009)
);

INVx1_ASAP7_75t_L g2010 ( 
.A(n_1962),
.Y(n_2010)
);

CKINVDCx5p33_ASAP7_75t_R g2011 ( 
.A(n_1886),
.Y(n_2011)
);

AOI22xp33_ASAP7_75t_L g2012 ( 
.A1(n_1896),
.A2(n_1851),
.B1(n_1827),
.B2(n_1854),
.Y(n_2012)
);

NOR2x1_ASAP7_75t_L g2013 ( 
.A(n_1963),
.B(n_1761),
.Y(n_2013)
);

INVx2_ASAP7_75t_SL g2014 ( 
.A(n_1890),
.Y(n_2014)
);

NOR2xp67_ASAP7_75t_L g2015 ( 
.A(n_1911),
.B(n_1764),
.Y(n_2015)
);

INVx2_ASAP7_75t_SL g2016 ( 
.A(n_1890),
.Y(n_2016)
);

AND2x4_ASAP7_75t_SL g2017 ( 
.A(n_1943),
.B(n_1958),
.Y(n_2017)
);

INVx3_ASAP7_75t_L g2018 ( 
.A(n_1952),
.Y(n_2018)
);

INVx1_ASAP7_75t_SL g2019 ( 
.A(n_1873),
.Y(n_2019)
);

INVx1_ASAP7_75t_L g2020 ( 
.A(n_1957),
.Y(n_2020)
);

INVx1_ASAP7_75t_L g2021 ( 
.A(n_1957),
.Y(n_2021)
);

AND2x2_ASAP7_75t_L g2022 ( 
.A(n_1959),
.B(n_1965),
.Y(n_2022)
);

AND2x2_ASAP7_75t_L g2023 ( 
.A(n_1967),
.B(n_1832),
.Y(n_2023)
);

OR2x2_ASAP7_75t_L g2024 ( 
.A(n_1960),
.B(n_1961),
.Y(n_2024)
);

INVx1_ASAP7_75t_L g2025 ( 
.A(n_1961),
.Y(n_2025)
);

NOR2x1_ASAP7_75t_SL g2026 ( 
.A(n_1920),
.B(n_1747),
.Y(n_2026)
);

INVx3_ASAP7_75t_L g2027 ( 
.A(n_1955),
.Y(n_2027)
);

NAND3xp33_ASAP7_75t_L g2028 ( 
.A(n_1911),
.B(n_1830),
.C(n_1831),
.Y(n_2028)
);

INVx2_ASAP7_75t_SL g2029 ( 
.A(n_1875),
.Y(n_2029)
);

NAND2xp5_ASAP7_75t_L g2030 ( 
.A(n_1874),
.B(n_1829),
.Y(n_2030)
);

NOR2xp33_ASAP7_75t_L g2031 ( 
.A(n_1888),
.B(n_1736),
.Y(n_2031)
);

AOI22xp5_ASAP7_75t_L g2032 ( 
.A1(n_1896),
.A2(n_1736),
.B1(n_1827),
.B2(n_1854),
.Y(n_2032)
);

BUFx3_ASAP7_75t_L g2033 ( 
.A(n_1870),
.Y(n_2033)
);

BUFx12f_ASAP7_75t_L g2034 ( 
.A(n_1900),
.Y(n_2034)
);

NAND2xp5_ASAP7_75t_L g2035 ( 
.A(n_1874),
.B(n_1830),
.Y(n_2035)
);

NAND2xp5_ASAP7_75t_L g2036 ( 
.A(n_1912),
.B(n_1831),
.Y(n_2036)
);

OR2x2_ASAP7_75t_L g2037 ( 
.A(n_1922),
.B(n_1914),
.Y(n_2037)
);

INVxp67_ASAP7_75t_SL g2038 ( 
.A(n_1894),
.Y(n_2038)
);

AND2x2_ASAP7_75t_L g2039 ( 
.A(n_1938),
.B(n_1832),
.Y(n_2039)
);

OR2x6_ASAP7_75t_L g2040 ( 
.A(n_2015),
.B(n_1920),
.Y(n_2040)
);

INVx1_ASAP7_75t_L g2041 ( 
.A(n_1969),
.Y(n_2041)
);

AND2x2_ASAP7_75t_L g2042 ( 
.A(n_1974),
.B(n_1916),
.Y(n_2042)
);

HB1xp67_ASAP7_75t_L g2043 ( 
.A(n_1985),
.Y(n_2043)
);

INVx1_ASAP7_75t_L g2044 ( 
.A(n_1969),
.Y(n_2044)
);

AND2x2_ASAP7_75t_L g2045 ( 
.A(n_2029),
.B(n_1920),
.Y(n_2045)
);

AOI22xp5_ASAP7_75t_L g2046 ( 
.A1(n_2007),
.A2(n_1905),
.B1(n_1909),
.B2(n_1917),
.Y(n_2046)
);

INVx2_ASAP7_75t_SL g2047 ( 
.A(n_1994),
.Y(n_2047)
);

INVx1_ASAP7_75t_L g2048 ( 
.A(n_1970),
.Y(n_2048)
);

INVx1_ASAP7_75t_L g2049 ( 
.A(n_1970),
.Y(n_2049)
);

NAND2xp5_ASAP7_75t_L g2050 ( 
.A(n_2038),
.B(n_1910),
.Y(n_2050)
);

AND2x2_ASAP7_75t_L g2051 ( 
.A(n_2018),
.B(n_1949),
.Y(n_2051)
);

AND2x2_ASAP7_75t_L g2052 ( 
.A(n_2018),
.B(n_1963),
.Y(n_2052)
);

INVx1_ASAP7_75t_L g2053 ( 
.A(n_1973),
.Y(n_2053)
);

NAND3xp33_ASAP7_75t_L g2054 ( 
.A(n_1987),
.B(n_1925),
.C(n_1933),
.Y(n_2054)
);

AND2x2_ASAP7_75t_L g2055 ( 
.A(n_2018),
.B(n_2027),
.Y(n_2055)
);

CKINVDCx16_ASAP7_75t_R g2056 ( 
.A(n_1981),
.Y(n_2056)
);

INVx2_ASAP7_75t_L g2057 ( 
.A(n_1990),
.Y(n_2057)
);

INVx2_ASAP7_75t_L g2058 ( 
.A(n_1990),
.Y(n_2058)
);

AO21x2_ASAP7_75t_L g2059 ( 
.A1(n_2015),
.A2(n_1941),
.B(n_1933),
.Y(n_2059)
);

AND2x2_ASAP7_75t_L g2060 ( 
.A(n_2027),
.B(n_1994),
.Y(n_2060)
);

AOI221xp5_ASAP7_75t_L g2061 ( 
.A1(n_2039),
.A2(n_1998),
.B1(n_1976),
.B2(n_1992),
.C(n_1940),
.Y(n_2061)
);

BUFx2_ASAP7_75t_L g2062 ( 
.A(n_2027),
.Y(n_2062)
);

NOR2x1_ASAP7_75t_SL g2063 ( 
.A(n_2001),
.B(n_1943),
.Y(n_2063)
);

AND2x2_ASAP7_75t_L g2064 ( 
.A(n_1994),
.B(n_1892),
.Y(n_2064)
);

OR2x2_ASAP7_75t_L g2065 ( 
.A(n_1975),
.B(n_1977),
.Y(n_2065)
);

OR2x2_ASAP7_75t_L g2066 ( 
.A(n_1975),
.B(n_1977),
.Y(n_2066)
);

AOI22xp33_ASAP7_75t_L g2067 ( 
.A1(n_2012),
.A2(n_1872),
.B1(n_1944),
.B2(n_1882),
.Y(n_2067)
);

NAND2xp5_ASAP7_75t_L g2068 ( 
.A(n_2030),
.B(n_1912),
.Y(n_2068)
);

INVx2_ASAP7_75t_L g2069 ( 
.A(n_1979),
.Y(n_2069)
);

HB1xp67_ASAP7_75t_L g2070 ( 
.A(n_2003),
.Y(n_2070)
);

BUFx2_ASAP7_75t_L g2071 ( 
.A(n_1978),
.Y(n_2071)
);

OAI33xp33_ASAP7_75t_L g2072 ( 
.A1(n_2001),
.A2(n_1988),
.A3(n_2035),
.B1(n_2021),
.B2(n_2025),
.B3(n_2020),
.Y(n_2072)
);

INVx2_ASAP7_75t_L g2073 ( 
.A(n_1980),
.Y(n_2073)
);

NOR2xp33_ASAP7_75t_L g2074 ( 
.A(n_2011),
.B(n_1883),
.Y(n_2074)
);

AND2x2_ASAP7_75t_L g2075 ( 
.A(n_2022),
.B(n_1938),
.Y(n_2075)
);

INVx2_ASAP7_75t_L g2076 ( 
.A(n_1986),
.Y(n_2076)
);

INVx1_ASAP7_75t_SL g2077 ( 
.A(n_2011),
.Y(n_2077)
);

AND2x4_ASAP7_75t_L g2078 ( 
.A(n_2026),
.B(n_1943),
.Y(n_2078)
);

OR2x6_ASAP7_75t_L g2079 ( 
.A(n_2028),
.B(n_1899),
.Y(n_2079)
);

NAND3xp33_ASAP7_75t_L g2080 ( 
.A(n_1989),
.B(n_1930),
.C(n_1940),
.Y(n_2080)
);

INVx2_ASAP7_75t_L g2081 ( 
.A(n_2005),
.Y(n_2081)
);

OAI221xp5_ASAP7_75t_L g2082 ( 
.A1(n_2032),
.A2(n_1887),
.B1(n_1872),
.B2(n_1930),
.C(n_1964),
.Y(n_2082)
);

AND2x2_ASAP7_75t_L g2083 ( 
.A(n_2022),
.B(n_1938),
.Y(n_2083)
);

BUFx6f_ASAP7_75t_L g2084 ( 
.A(n_1981),
.Y(n_2084)
);

INVx5_ASAP7_75t_SL g2085 ( 
.A(n_2009),
.Y(n_2085)
);

AND4x1_ASAP7_75t_L g2086 ( 
.A(n_1995),
.B(n_1898),
.C(n_1946),
.D(n_1906),
.Y(n_2086)
);

AOI22xp33_ASAP7_75t_L g2087 ( 
.A1(n_1984),
.A2(n_1944),
.B1(n_1882),
.B2(n_1869),
.Y(n_2087)
);

AOI22xp33_ASAP7_75t_L g2088 ( 
.A1(n_1984),
.A2(n_1867),
.B1(n_1879),
.B2(n_1884),
.Y(n_2088)
);

OAI33xp33_ASAP7_75t_L g2089 ( 
.A1(n_2020),
.A2(n_1919),
.A3(n_1894),
.B1(n_1903),
.B2(n_1898),
.B3(n_1864),
.Y(n_2089)
);

AOI22xp33_ASAP7_75t_L g2090 ( 
.A1(n_2000),
.A2(n_1877),
.B1(n_1923),
.B2(n_1876),
.Y(n_2090)
);

NOR2x1_ASAP7_75t_L g2091 ( 
.A(n_2013),
.B(n_2037),
.Y(n_2091)
);

HB1xp67_ASAP7_75t_L g2092 ( 
.A(n_2006),
.Y(n_2092)
);

BUFx2_ASAP7_75t_L g2093 ( 
.A(n_1978),
.Y(n_2093)
);

HB1xp67_ASAP7_75t_L g2094 ( 
.A(n_1999),
.Y(n_2094)
);

AND2x2_ASAP7_75t_L g2095 ( 
.A(n_1972),
.B(n_1923),
.Y(n_2095)
);

AND2x2_ASAP7_75t_L g2096 ( 
.A(n_2002),
.B(n_1982),
.Y(n_2096)
);

INVx3_ASAP7_75t_L g2097 ( 
.A(n_2078),
.Y(n_2097)
);

INVx1_ASAP7_75t_L g2098 ( 
.A(n_2069),
.Y(n_2098)
);

INVx1_ASAP7_75t_L g2099 ( 
.A(n_2069),
.Y(n_2099)
);

INVx2_ASAP7_75t_L g2100 ( 
.A(n_2069),
.Y(n_2100)
);

AND2x2_ASAP7_75t_L g2101 ( 
.A(n_2071),
.B(n_1976),
.Y(n_2101)
);

OR2x2_ASAP7_75t_L g2102 ( 
.A(n_2065),
.B(n_2037),
.Y(n_2102)
);

AND2x2_ASAP7_75t_L g2103 ( 
.A(n_2071),
.B(n_2093),
.Y(n_2103)
);

AND2x2_ASAP7_75t_L g2104 ( 
.A(n_2093),
.B(n_1982),
.Y(n_2104)
);

INVx1_ASAP7_75t_L g2105 ( 
.A(n_2076),
.Y(n_2105)
);

NAND2xp5_ASAP7_75t_L g2106 ( 
.A(n_2057),
.B(n_2021),
.Y(n_2106)
);

INVx1_ASAP7_75t_L g2107 ( 
.A(n_2076),
.Y(n_2107)
);

INVx1_ASAP7_75t_L g2108 ( 
.A(n_2076),
.Y(n_2108)
);

NAND2xp5_ASAP7_75t_L g2109 ( 
.A(n_2057),
.B(n_2025),
.Y(n_2109)
);

AND2x2_ASAP7_75t_L g2110 ( 
.A(n_2075),
.B(n_2039),
.Y(n_2110)
);

BUFx2_ASAP7_75t_L g2111 ( 
.A(n_2078),
.Y(n_2111)
);

OR2x2_ASAP7_75t_L g2112 ( 
.A(n_2065),
.B(n_2024),
.Y(n_2112)
);

OR2x2_ASAP7_75t_L g2113 ( 
.A(n_2066),
.B(n_2024),
.Y(n_2113)
);

NAND2xp5_ASAP7_75t_L g2114 ( 
.A(n_2057),
.B(n_2023),
.Y(n_2114)
);

AND2x4_ASAP7_75t_L g2115 ( 
.A(n_2078),
.B(n_2026),
.Y(n_2115)
);

NAND2xp5_ASAP7_75t_L g2116 ( 
.A(n_2058),
.B(n_2023),
.Y(n_2116)
);

AND2x2_ASAP7_75t_L g2117 ( 
.A(n_2075),
.B(n_1983),
.Y(n_2117)
);

AND2x2_ASAP7_75t_L g2118 ( 
.A(n_2083),
.B(n_1983),
.Y(n_2118)
);

NAND3xp33_ASAP7_75t_SL g2119 ( 
.A(n_2086),
.B(n_2019),
.C(n_2031),
.Y(n_2119)
);

INVx1_ASAP7_75t_L g2120 ( 
.A(n_2081),
.Y(n_2120)
);

OAI221xp5_ASAP7_75t_L g2121 ( 
.A1(n_2080),
.A2(n_2033),
.B1(n_1958),
.B2(n_1891),
.C(n_1956),
.Y(n_2121)
);

INVx1_ASAP7_75t_L g2122 ( 
.A(n_2081),
.Y(n_2122)
);

INVx2_ASAP7_75t_L g2123 ( 
.A(n_2081),
.Y(n_2123)
);

INVx1_ASAP7_75t_L g2124 ( 
.A(n_2073),
.Y(n_2124)
);

AND2x2_ASAP7_75t_L g2125 ( 
.A(n_2083),
.B(n_1991),
.Y(n_2125)
);

INVx2_ASAP7_75t_L g2126 ( 
.A(n_2058),
.Y(n_2126)
);

AND2x4_ASAP7_75t_L g2127 ( 
.A(n_2078),
.B(n_2013),
.Y(n_2127)
);

AND2x4_ASAP7_75t_L g2128 ( 
.A(n_2063),
.B(n_2009),
.Y(n_2128)
);

AND2x2_ASAP7_75t_L g2129 ( 
.A(n_2060),
.B(n_1991),
.Y(n_2129)
);

AND2x2_ASAP7_75t_L g2130 ( 
.A(n_2051),
.B(n_1993),
.Y(n_2130)
);

OR2x2_ASAP7_75t_L g2131 ( 
.A(n_2066),
.B(n_2058),
.Y(n_2131)
);

AND2x2_ASAP7_75t_L g2132 ( 
.A(n_2051),
.B(n_2002),
.Y(n_2132)
);

INVx1_ASAP7_75t_L g2133 ( 
.A(n_2073),
.Y(n_2133)
);

INVx2_ASAP7_75t_L g2134 ( 
.A(n_2052),
.Y(n_2134)
);

INVx4_ASAP7_75t_L g2135 ( 
.A(n_2084),
.Y(n_2135)
);

INVx2_ASAP7_75t_SL g2136 ( 
.A(n_2084),
.Y(n_2136)
);

NOR2xp33_ASAP7_75t_L g2137 ( 
.A(n_2056),
.B(n_2033),
.Y(n_2137)
);

INVxp67_ASAP7_75t_SL g2138 ( 
.A(n_2091),
.Y(n_2138)
);

AND2x2_ASAP7_75t_L g2139 ( 
.A(n_2096),
.B(n_1996),
.Y(n_2139)
);

OR2x2_ASAP7_75t_L g2140 ( 
.A(n_2050),
.B(n_1971),
.Y(n_2140)
);

NAND2xp5_ASAP7_75t_L g2141 ( 
.A(n_2070),
.B(n_2008),
.Y(n_2141)
);

OR2x6_ASAP7_75t_L g2142 ( 
.A(n_2040),
.B(n_2079),
.Y(n_2142)
);

INVx1_ASAP7_75t_L g2143 ( 
.A(n_2041),
.Y(n_2143)
);

INVx1_ASAP7_75t_L g2144 ( 
.A(n_2041),
.Y(n_2144)
);

INVx2_ASAP7_75t_L g2145 ( 
.A(n_2052),
.Y(n_2145)
);

INVx1_ASAP7_75t_L g2146 ( 
.A(n_2044),
.Y(n_2146)
);

OR2x2_ASAP7_75t_L g2147 ( 
.A(n_2092),
.B(n_1971),
.Y(n_2147)
);

NAND2xp5_ASAP7_75t_L g2148 ( 
.A(n_2044),
.B(n_2010),
.Y(n_2148)
);

AND2x2_ASAP7_75t_L g2149 ( 
.A(n_2055),
.B(n_1997),
.Y(n_2149)
);

AND2x2_ASAP7_75t_L g2150 ( 
.A(n_2055),
.B(n_2004),
.Y(n_2150)
);

AND2x2_ASAP7_75t_L g2151 ( 
.A(n_2085),
.B(n_2004),
.Y(n_2151)
);

INVx1_ASAP7_75t_L g2152 ( 
.A(n_2048),
.Y(n_2152)
);

NAND2xp5_ASAP7_75t_L g2153 ( 
.A(n_2048),
.B(n_2010),
.Y(n_2153)
);

OR2x2_ASAP7_75t_L g2154 ( 
.A(n_2102),
.B(n_2054),
.Y(n_2154)
);

OAI211xp5_ASAP7_75t_SL g2155 ( 
.A1(n_2121),
.A2(n_2061),
.B(n_2046),
.C(n_2091),
.Y(n_2155)
);

AOI32xp33_ASAP7_75t_L g2156 ( 
.A1(n_2121),
.A2(n_2082),
.A3(n_2090),
.B1(n_2087),
.B2(n_2067),
.Y(n_2156)
);

INVx1_ASAP7_75t_L g2157 ( 
.A(n_2143),
.Y(n_2157)
);

INVx1_ASAP7_75t_L g2158 ( 
.A(n_2143),
.Y(n_2158)
);

INVx1_ASAP7_75t_L g2159 ( 
.A(n_2144),
.Y(n_2159)
);

INVx1_ASAP7_75t_L g2160 ( 
.A(n_2144),
.Y(n_2160)
);

INVx3_ASAP7_75t_L g2161 ( 
.A(n_2128),
.Y(n_2161)
);

INVx1_ASAP7_75t_L g2162 ( 
.A(n_2146),
.Y(n_2162)
);

AND2x4_ASAP7_75t_L g2163 ( 
.A(n_2136),
.B(n_2063),
.Y(n_2163)
);

NAND3xp33_ASAP7_75t_L g2164 ( 
.A(n_2138),
.B(n_2046),
.C(n_2086),
.Y(n_2164)
);

AND2x2_ASAP7_75t_L g2165 ( 
.A(n_2132),
.B(n_2085),
.Y(n_2165)
);

INVx1_ASAP7_75t_L g2166 ( 
.A(n_2146),
.Y(n_2166)
);

INVx1_ASAP7_75t_L g2167 ( 
.A(n_2152),
.Y(n_2167)
);

AND2x2_ASAP7_75t_L g2168 ( 
.A(n_2132),
.B(n_2085),
.Y(n_2168)
);

INVxp67_ASAP7_75t_L g2169 ( 
.A(n_2140),
.Y(n_2169)
);

INVx1_ASAP7_75t_L g2170 ( 
.A(n_2152),
.Y(n_2170)
);

NAND2xp5_ASAP7_75t_L g2171 ( 
.A(n_2140),
.B(n_2043),
.Y(n_2171)
);

AND2x2_ASAP7_75t_L g2172 ( 
.A(n_2128),
.B(n_2130),
.Y(n_2172)
);

INVx2_ASAP7_75t_SL g2173 ( 
.A(n_2136),
.Y(n_2173)
);

OR2x6_ASAP7_75t_L g2174 ( 
.A(n_2135),
.B(n_2084),
.Y(n_2174)
);

INVx2_ASAP7_75t_L g2175 ( 
.A(n_2111),
.Y(n_2175)
);

OR2x2_ASAP7_75t_L g2176 ( 
.A(n_2102),
.B(n_2112),
.Y(n_2176)
);

INVx1_ASAP7_75t_L g2177 ( 
.A(n_2148),
.Y(n_2177)
);

NAND2xp5_ASAP7_75t_L g2178 ( 
.A(n_2130),
.B(n_2068),
.Y(n_2178)
);

AOI22xp5_ASAP7_75t_L g2179 ( 
.A1(n_2119),
.A2(n_2089),
.B1(n_2056),
.B2(n_2084),
.Y(n_2179)
);

INVx1_ASAP7_75t_L g2180 ( 
.A(n_2148),
.Y(n_2180)
);

INVx1_ASAP7_75t_L g2181 ( 
.A(n_2153),
.Y(n_2181)
);

INVx1_ASAP7_75t_L g2182 ( 
.A(n_2153),
.Y(n_2182)
);

NAND2xp5_ASAP7_75t_L g2183 ( 
.A(n_2106),
.B(n_2049),
.Y(n_2183)
);

NAND2xp5_ASAP7_75t_L g2184 ( 
.A(n_2106),
.B(n_2109),
.Y(n_2184)
);

INVx1_ASAP7_75t_L g2185 ( 
.A(n_2141),
.Y(n_2185)
);

OR2x2_ASAP7_75t_L g2186 ( 
.A(n_2112),
.B(n_2113),
.Y(n_2186)
);

AND2x4_ASAP7_75t_SL g2187 ( 
.A(n_2137),
.B(n_1958),
.Y(n_2187)
);

NAND2xp5_ASAP7_75t_L g2188 ( 
.A(n_2109),
.B(n_2049),
.Y(n_2188)
);

INVx1_ASAP7_75t_L g2189 ( 
.A(n_2141),
.Y(n_2189)
);

INVx1_ASAP7_75t_L g2190 ( 
.A(n_2147),
.Y(n_2190)
);

INVx1_ASAP7_75t_L g2191 ( 
.A(n_2147),
.Y(n_2191)
);

INVx1_ASAP7_75t_L g2192 ( 
.A(n_2124),
.Y(n_2192)
);

NAND2xp5_ASAP7_75t_L g2193 ( 
.A(n_2139),
.B(n_2095),
.Y(n_2193)
);

INVx1_ASAP7_75t_L g2194 ( 
.A(n_2124),
.Y(n_2194)
);

INVx1_ASAP7_75t_L g2195 ( 
.A(n_2133),
.Y(n_2195)
);

AND2x2_ASAP7_75t_L g2196 ( 
.A(n_2128),
.B(n_2085),
.Y(n_2196)
);

OR2x6_ASAP7_75t_L g2197 ( 
.A(n_2135),
.B(n_2084),
.Y(n_2197)
);

NAND2xp5_ASAP7_75t_L g2198 ( 
.A(n_2139),
.B(n_2095),
.Y(n_2198)
);

NOR2xp33_ASAP7_75t_L g2199 ( 
.A(n_2119),
.B(n_2084),
.Y(n_2199)
);

OR2x2_ASAP7_75t_L g2200 ( 
.A(n_2113),
.B(n_2094),
.Y(n_2200)
);

INVx1_ASAP7_75t_L g2201 ( 
.A(n_2133),
.Y(n_2201)
);

INVx2_ASAP7_75t_L g2202 ( 
.A(n_2111),
.Y(n_2202)
);

OR2x2_ASAP7_75t_L g2203 ( 
.A(n_2114),
.B(n_2036),
.Y(n_2203)
);

OR2x2_ASAP7_75t_L g2204 ( 
.A(n_2114),
.B(n_2042),
.Y(n_2204)
);

INVx1_ASAP7_75t_L g2205 ( 
.A(n_2098),
.Y(n_2205)
);

OR2x2_ASAP7_75t_L g2206 ( 
.A(n_2116),
.B(n_2042),
.Y(n_2206)
);

NAND2xp5_ASAP7_75t_L g2207 ( 
.A(n_2117),
.B(n_2053),
.Y(n_2207)
);

INVx1_ASAP7_75t_L g2208 ( 
.A(n_2098),
.Y(n_2208)
);

INVx1_ASAP7_75t_L g2209 ( 
.A(n_2099),
.Y(n_2209)
);

INVx1_ASAP7_75t_L g2210 ( 
.A(n_2099),
.Y(n_2210)
);

INVx1_ASAP7_75t_L g2211 ( 
.A(n_2157),
.Y(n_2211)
);

OR2x2_ASAP7_75t_L g2212 ( 
.A(n_2176),
.B(n_2186),
.Y(n_2212)
);

AND2x4_ASAP7_75t_L g2213 ( 
.A(n_2172),
.B(n_2128),
.Y(n_2213)
);

INVx2_ASAP7_75t_L g2214 ( 
.A(n_2173),
.Y(n_2214)
);

INVxp67_ASAP7_75t_SL g2215 ( 
.A(n_2199),
.Y(n_2215)
);

INVx1_ASAP7_75t_L g2216 ( 
.A(n_2158),
.Y(n_2216)
);

OR2x2_ASAP7_75t_L g2217 ( 
.A(n_2154),
.B(n_2131),
.Y(n_2217)
);

INVxp67_ASAP7_75t_L g2218 ( 
.A(n_2164),
.Y(n_2218)
);

NOR2xp33_ASAP7_75t_L g2219 ( 
.A(n_2187),
.B(n_2077),
.Y(n_2219)
);

NAND2xp5_ASAP7_75t_L g2220 ( 
.A(n_2156),
.B(n_2136),
.Y(n_2220)
);

OR2x2_ASAP7_75t_L g2221 ( 
.A(n_2178),
.B(n_2207),
.Y(n_2221)
);

NAND2xp5_ASAP7_75t_L g2222 ( 
.A(n_2179),
.B(n_2117),
.Y(n_2222)
);

NAND2xp5_ASAP7_75t_L g2223 ( 
.A(n_2179),
.B(n_2118),
.Y(n_2223)
);

INVx1_ASAP7_75t_SL g2224 ( 
.A(n_2165),
.Y(n_2224)
);

INVx1_ASAP7_75t_L g2225 ( 
.A(n_2159),
.Y(n_2225)
);

HB1xp67_ASAP7_75t_L g2226 ( 
.A(n_2175),
.Y(n_2226)
);

NOR2x1_ASAP7_75t_R g2227 ( 
.A(n_2163),
.B(n_2034),
.Y(n_2227)
);

INVx1_ASAP7_75t_L g2228 ( 
.A(n_2160),
.Y(n_2228)
);

NAND2xp5_ASAP7_75t_L g2229 ( 
.A(n_2169),
.B(n_2118),
.Y(n_2229)
);

AND2x2_ASAP7_75t_L g2230 ( 
.A(n_2196),
.B(n_2115),
.Y(n_2230)
);

INVx2_ASAP7_75t_L g2231 ( 
.A(n_2202),
.Y(n_2231)
);

INVx1_ASAP7_75t_L g2232 ( 
.A(n_2162),
.Y(n_2232)
);

OAI21xp5_ASAP7_75t_L g2233 ( 
.A1(n_2164),
.A2(n_2138),
.B(n_2142),
.Y(n_2233)
);

INVx1_ASAP7_75t_L g2234 ( 
.A(n_2166),
.Y(n_2234)
);

NAND2xp5_ASAP7_75t_L g2235 ( 
.A(n_2190),
.B(n_2135),
.Y(n_2235)
);

INVx2_ASAP7_75t_L g2236 ( 
.A(n_2161),
.Y(n_2236)
);

OR2x2_ASAP7_75t_L g2237 ( 
.A(n_2178),
.B(n_2131),
.Y(n_2237)
);

CKINVDCx16_ASAP7_75t_R g2238 ( 
.A(n_2174),
.Y(n_2238)
);

INVx1_ASAP7_75t_L g2239 ( 
.A(n_2167),
.Y(n_2239)
);

AOI22xp33_ASAP7_75t_L g2240 ( 
.A1(n_2155),
.A2(n_2142),
.B1(n_2059),
.B2(n_2072),
.Y(n_2240)
);

INVx1_ASAP7_75t_L g2241 ( 
.A(n_2170),
.Y(n_2241)
);

INVx1_ASAP7_75t_L g2242 ( 
.A(n_2192),
.Y(n_2242)
);

OR2x2_ASAP7_75t_L g2243 ( 
.A(n_2207),
.B(n_2116),
.Y(n_2243)
);

OR2x2_ASAP7_75t_L g2244 ( 
.A(n_2191),
.B(n_2126),
.Y(n_2244)
);

INVx2_ASAP7_75t_L g2245 ( 
.A(n_2161),
.Y(n_2245)
);

AND2x2_ASAP7_75t_L g2246 ( 
.A(n_2168),
.B(n_2115),
.Y(n_2246)
);

INVx1_ASAP7_75t_L g2247 ( 
.A(n_2194),
.Y(n_2247)
);

AND2x4_ASAP7_75t_L g2248 ( 
.A(n_2174),
.B(n_2115),
.Y(n_2248)
);

HB1xp67_ASAP7_75t_L g2249 ( 
.A(n_2174),
.Y(n_2249)
);

INVx1_ASAP7_75t_L g2250 ( 
.A(n_2195),
.Y(n_2250)
);

OR2x6_ASAP7_75t_L g2251 ( 
.A(n_2197),
.B(n_2135),
.Y(n_2251)
);

NAND2xp5_ASAP7_75t_L g2252 ( 
.A(n_2185),
.B(n_2104),
.Y(n_2252)
);

INVx2_ASAP7_75t_L g2253 ( 
.A(n_2197),
.Y(n_2253)
);

NAND2xp33_ASAP7_75t_SL g2254 ( 
.A(n_2240),
.B(n_2163),
.Y(n_2254)
);

AOI211xp5_ASAP7_75t_L g2255 ( 
.A1(n_2218),
.A2(n_2189),
.B(n_2171),
.C(n_2115),
.Y(n_2255)
);

OAI322xp33_ASAP7_75t_L g2256 ( 
.A1(n_2220),
.A2(n_2182),
.A3(n_2181),
.B1(n_2177),
.B2(n_2180),
.C1(n_2184),
.C2(n_2200),
.Y(n_2256)
);

INVx1_ASAP7_75t_L g2257 ( 
.A(n_2232),
.Y(n_2257)
);

OAI21xp5_ASAP7_75t_L g2258 ( 
.A1(n_2233),
.A2(n_2197),
.B(n_2142),
.Y(n_2258)
);

INVx1_ASAP7_75t_L g2259 ( 
.A(n_2232),
.Y(n_2259)
);

INVx1_ASAP7_75t_L g2260 ( 
.A(n_2241),
.Y(n_2260)
);

AOI222xp33_ASAP7_75t_L g2261 ( 
.A1(n_2222),
.A2(n_2101),
.B1(n_2127),
.B2(n_2184),
.C1(n_2074),
.C2(n_2198),
.Y(n_2261)
);

INVx2_ASAP7_75t_L g2262 ( 
.A(n_2236),
.Y(n_2262)
);

AOI322xp5_ASAP7_75t_L g2263 ( 
.A1(n_2223),
.A2(n_2101),
.A3(n_2125),
.B1(n_2110),
.B2(n_2193),
.C1(n_2104),
.C2(n_2127),
.Y(n_2263)
);

NAND2xp5_ASAP7_75t_L g2264 ( 
.A(n_2215),
.B(n_2204),
.Y(n_2264)
);

NOR2xp33_ASAP7_75t_L g2265 ( 
.A(n_2227),
.B(n_2034),
.Y(n_2265)
);

OAI211xp5_ASAP7_75t_SL g2266 ( 
.A1(n_2224),
.A2(n_2201),
.B(n_2097),
.C(n_2208),
.Y(n_2266)
);

OR2x2_ASAP7_75t_L g2267 ( 
.A(n_2212),
.B(n_2206),
.Y(n_2267)
);

INVx2_ASAP7_75t_L g2268 ( 
.A(n_2236),
.Y(n_2268)
);

NAND4xp25_ASAP7_75t_SL g2269 ( 
.A(n_2230),
.B(n_2088),
.C(n_2151),
.D(n_2103),
.Y(n_2269)
);

NAND2xp5_ASAP7_75t_L g2270 ( 
.A(n_2226),
.B(n_2203),
.Y(n_2270)
);

AOI21xp33_ASAP7_75t_L g2271 ( 
.A1(n_2235),
.A2(n_2142),
.B(n_2059),
.Y(n_2271)
);

AOI22xp33_ASAP7_75t_SL g2272 ( 
.A1(n_2238),
.A2(n_2059),
.B1(n_2142),
.B2(n_2097),
.Y(n_2272)
);

NAND2xp5_ASAP7_75t_L g2273 ( 
.A(n_2231),
.B(n_2103),
.Y(n_2273)
);

NOR2xp33_ASAP7_75t_L g2274 ( 
.A(n_2219),
.B(n_1948),
.Y(n_2274)
);

NOR2xp33_ASAP7_75t_L g2275 ( 
.A(n_2212),
.B(n_2064),
.Y(n_2275)
);

INVx1_ASAP7_75t_SL g2276 ( 
.A(n_2217),
.Y(n_2276)
);

NAND2xp5_ASAP7_75t_SL g2277 ( 
.A(n_2248),
.B(n_2217),
.Y(n_2277)
);

OAI311xp33_ASAP7_75t_L g2278 ( 
.A1(n_2229),
.A2(n_2097),
.A3(n_2188),
.B1(n_2183),
.C1(n_2205),
.Y(n_2278)
);

OAI21xp33_ASAP7_75t_L g2279 ( 
.A1(n_2252),
.A2(n_2079),
.B(n_2097),
.Y(n_2279)
);

AND2x2_ASAP7_75t_L g2280 ( 
.A(n_2230),
.B(n_2246),
.Y(n_2280)
);

INVx2_ASAP7_75t_L g2281 ( 
.A(n_2245),
.Y(n_2281)
);

INVx1_ASAP7_75t_SL g2282 ( 
.A(n_2249),
.Y(n_2282)
);

AOI22xp5_ASAP7_75t_L g2283 ( 
.A1(n_2246),
.A2(n_2040),
.B1(n_2079),
.B2(n_2127),
.Y(n_2283)
);

NAND2xp5_ASAP7_75t_L g2284 ( 
.A(n_2282),
.B(n_2231),
.Y(n_2284)
);

AND2x2_ASAP7_75t_L g2285 ( 
.A(n_2280),
.B(n_2213),
.Y(n_2285)
);

NAND2xp5_ASAP7_75t_L g2286 ( 
.A(n_2276),
.B(n_2253),
.Y(n_2286)
);

NAND2xp5_ASAP7_75t_L g2287 ( 
.A(n_2277),
.B(n_2253),
.Y(n_2287)
);

NOR3xp33_ASAP7_75t_SL g2288 ( 
.A(n_2254),
.B(n_2269),
.C(n_2258),
.Y(n_2288)
);

INVx1_ASAP7_75t_L g2289 ( 
.A(n_2257),
.Y(n_2289)
);

OAI21xp5_ASAP7_75t_L g2290 ( 
.A1(n_2278),
.A2(n_2251),
.B(n_2248),
.Y(n_2290)
);

NAND2xp5_ASAP7_75t_L g2291 ( 
.A(n_2277),
.B(n_2214),
.Y(n_2291)
);

INVx2_ASAP7_75t_L g2292 ( 
.A(n_2262),
.Y(n_2292)
);

INVx1_ASAP7_75t_SL g2293 ( 
.A(n_2273),
.Y(n_2293)
);

INVx1_ASAP7_75t_L g2294 ( 
.A(n_2259),
.Y(n_2294)
);

OAI21xp5_ASAP7_75t_L g2295 ( 
.A1(n_2272),
.A2(n_2251),
.B(n_2248),
.Y(n_2295)
);

AOI221xp5_ASAP7_75t_L g2296 ( 
.A1(n_2256),
.A2(n_2241),
.B1(n_2216),
.B2(n_2234),
.C(n_2225),
.Y(n_2296)
);

AOI21xp33_ASAP7_75t_SL g2297 ( 
.A1(n_2265),
.A2(n_2251),
.B(n_2214),
.Y(n_2297)
);

INVx1_ASAP7_75t_L g2298 ( 
.A(n_2260),
.Y(n_2298)
);

OAI211xp5_ASAP7_75t_L g2299 ( 
.A1(n_2261),
.A2(n_2245),
.B(n_2239),
.C(n_2211),
.Y(n_2299)
);

NOR2xp33_ASAP7_75t_L g2300 ( 
.A(n_2274),
.B(n_2265),
.Y(n_2300)
);

OAI21xp5_ASAP7_75t_SL g2301 ( 
.A1(n_2263),
.A2(n_2213),
.B(n_2221),
.Y(n_2301)
);

AND2x2_ASAP7_75t_L g2302 ( 
.A(n_2275),
.B(n_2213),
.Y(n_2302)
);

INVx1_ASAP7_75t_L g2303 ( 
.A(n_2262),
.Y(n_2303)
);

INVx1_ASAP7_75t_L g2304 ( 
.A(n_2268),
.Y(n_2304)
);

INVx1_ASAP7_75t_L g2305 ( 
.A(n_2268),
.Y(n_2305)
);

INVx1_ASAP7_75t_L g2306 ( 
.A(n_2281),
.Y(n_2306)
);

XNOR2x1_ASAP7_75t_L g2307 ( 
.A(n_2293),
.B(n_2264),
.Y(n_2307)
);

INVx1_ASAP7_75t_L g2308 ( 
.A(n_2292),
.Y(n_2308)
);

AOI221xp5_ASAP7_75t_L g2309 ( 
.A1(n_2288),
.A2(n_2255),
.B1(n_2271),
.B2(n_2266),
.C(n_2279),
.Y(n_2309)
);

AOI221xp5_ASAP7_75t_L g2310 ( 
.A1(n_2301),
.A2(n_2270),
.B1(n_2281),
.B2(n_2275),
.C(n_2267),
.Y(n_2310)
);

AOI22xp5_ASAP7_75t_L g2311 ( 
.A1(n_2285),
.A2(n_2302),
.B1(n_2300),
.B2(n_2287),
.Y(n_2311)
);

A2O1A1Ixp33_ASAP7_75t_L g2312 ( 
.A1(n_2290),
.A2(n_2283),
.B(n_2274),
.C(n_2127),
.Y(n_2312)
);

AND2x2_ASAP7_75t_L g2313 ( 
.A(n_2285),
.B(n_2251),
.Y(n_2313)
);

NAND2xp5_ASAP7_75t_L g2314 ( 
.A(n_2291),
.B(n_2228),
.Y(n_2314)
);

AOI21xp33_ASAP7_75t_L g2315 ( 
.A1(n_2284),
.A2(n_2247),
.B(n_2242),
.Y(n_2315)
);

INVx1_ASAP7_75t_L g2316 ( 
.A(n_2292),
.Y(n_2316)
);

OAI322xp33_ASAP7_75t_L g2317 ( 
.A1(n_2286),
.A2(n_2221),
.A3(n_2247),
.B1(n_2250),
.B2(n_2244),
.C1(n_2243),
.C2(n_2237),
.Y(n_2317)
);

OAI22xp33_ASAP7_75t_SL g2318 ( 
.A1(n_2295),
.A2(n_2244),
.B1(n_2237),
.B2(n_2243),
.Y(n_2318)
);

NAND2xp33_ASAP7_75t_L g2319 ( 
.A(n_2302),
.B(n_1736),
.Y(n_2319)
);

OAI21xp33_ASAP7_75t_L g2320 ( 
.A1(n_2297),
.A2(n_2079),
.B(n_2209),
.Y(n_2320)
);

INVx1_ASAP7_75t_L g2321 ( 
.A(n_2303),
.Y(n_2321)
);

INVx1_ASAP7_75t_L g2322 ( 
.A(n_2308),
.Y(n_2322)
);

INVx1_ASAP7_75t_L g2323 ( 
.A(n_2316),
.Y(n_2323)
);

NAND4xp25_ASAP7_75t_L g2324 ( 
.A(n_2311),
.B(n_2296),
.C(n_2299),
.D(n_2298),
.Y(n_2324)
);

NAND2xp5_ASAP7_75t_L g2325 ( 
.A(n_2310),
.B(n_2306),
.Y(n_2325)
);

OAI211xp5_ASAP7_75t_L g2326 ( 
.A1(n_2309),
.A2(n_2289),
.B(n_2294),
.C(n_2303),
.Y(n_2326)
);

NAND2xp5_ASAP7_75t_L g2327 ( 
.A(n_2307),
.B(n_2304),
.Y(n_2327)
);

INVx1_ASAP7_75t_L g2328 ( 
.A(n_2321),
.Y(n_2328)
);

NOR3xp33_ASAP7_75t_L g2329 ( 
.A(n_2318),
.B(n_2305),
.C(n_2304),
.Y(n_2329)
);

NOR3xp33_ASAP7_75t_L g2330 ( 
.A(n_2312),
.B(n_2305),
.C(n_2289),
.Y(n_2330)
);

NAND4xp25_ASAP7_75t_L g2331 ( 
.A(n_2313),
.B(n_1868),
.C(n_1871),
.D(n_1926),
.Y(n_2331)
);

INVx1_ASAP7_75t_L g2332 ( 
.A(n_2314),
.Y(n_2332)
);

O2A1O1Ixp33_ASAP7_75t_L g2333 ( 
.A1(n_2315),
.A2(n_2079),
.B(n_2210),
.C(n_2183),
.Y(n_2333)
);

NAND2xp5_ASAP7_75t_L g2334 ( 
.A(n_2315),
.B(n_2188),
.Y(n_2334)
);

XNOR2xp5_ASAP7_75t_L g2335 ( 
.A(n_2320),
.B(n_2064),
.Y(n_2335)
);

NAND4xp25_ASAP7_75t_SL g2336 ( 
.A(n_2327),
.B(n_2319),
.C(n_2317),
.D(n_2151),
.Y(n_2336)
);

NOR2xp33_ASAP7_75t_L g2337 ( 
.A(n_2324),
.B(n_2126),
.Y(n_2337)
);

AOI221xp5_ASAP7_75t_L g2338 ( 
.A1(n_2325),
.A2(n_2126),
.B1(n_2134),
.B2(n_2145),
.C(n_1932),
.Y(n_2338)
);

OAI221xp5_ASAP7_75t_L g2339 ( 
.A1(n_2330),
.A2(n_2040),
.B1(n_1878),
.B2(n_1926),
.C(n_2014),
.Y(n_2339)
);

NAND2xp5_ASAP7_75t_L g2340 ( 
.A(n_2329),
.B(n_2110),
.Y(n_2340)
);

NAND2xp5_ASAP7_75t_L g2341 ( 
.A(n_2332),
.B(n_2326),
.Y(n_2341)
);

NAND4xp25_ASAP7_75t_L g2342 ( 
.A(n_2326),
.B(n_1878),
.C(n_1885),
.D(n_1855),
.Y(n_2342)
);

INVx1_ASAP7_75t_L g2343 ( 
.A(n_2322),
.Y(n_2343)
);

AOI211xp5_ASAP7_75t_L g2344 ( 
.A1(n_2334),
.A2(n_1736),
.B(n_2045),
.C(n_2145),
.Y(n_2344)
);

NAND2xp5_ASAP7_75t_L g2345 ( 
.A(n_2323),
.B(n_2125),
.Y(n_2345)
);

OAI21xp5_ASAP7_75t_L g2346 ( 
.A1(n_2333),
.A2(n_2145),
.B(n_2134),
.Y(n_2346)
);

AOI22xp5_ASAP7_75t_L g2347 ( 
.A1(n_2331),
.A2(n_2040),
.B1(n_2017),
.B2(n_2014),
.Y(n_2347)
);

INVx1_ASAP7_75t_L g2348 ( 
.A(n_2345),
.Y(n_2348)
);

AOI21xp5_ASAP7_75t_L g2349 ( 
.A1(n_2341),
.A2(n_2328),
.B(n_2335),
.Y(n_2349)
);

OAI211xp5_ASAP7_75t_SL g2350 ( 
.A1(n_2337),
.A2(n_2016),
.B(n_1953),
.C(n_2134),
.Y(n_2350)
);

NAND2xp5_ASAP7_75t_L g2351 ( 
.A(n_2340),
.B(n_2129),
.Y(n_2351)
);

INVx1_ASAP7_75t_L g2352 ( 
.A(n_2343),
.Y(n_2352)
);

AOI211xp5_ASAP7_75t_L g2353 ( 
.A1(n_2336),
.A2(n_2045),
.B(n_1855),
.C(n_2016),
.Y(n_2353)
);

OAI211xp5_ASAP7_75t_L g2354 ( 
.A1(n_2342),
.A2(n_2062),
.B(n_1863),
.C(n_1865),
.Y(n_2354)
);

INVx1_ASAP7_75t_L g2355 ( 
.A(n_2344),
.Y(n_2355)
);

OAI211xp5_ASAP7_75t_SL g2356 ( 
.A1(n_2338),
.A2(n_2120),
.B(n_2108),
.C(n_2107),
.Y(n_2356)
);

NOR2xp33_ASAP7_75t_L g2357 ( 
.A(n_2351),
.B(n_2339),
.Y(n_2357)
);

INVxp67_ASAP7_75t_SL g2358 ( 
.A(n_2349),
.Y(n_2358)
);

NOR2x1_ASAP7_75t_L g2359 ( 
.A(n_2352),
.B(n_2346),
.Y(n_2359)
);

OR2x2_ASAP7_75t_L g2360 ( 
.A(n_2355),
.B(n_2347),
.Y(n_2360)
);

NOR2xp33_ASAP7_75t_L g2361 ( 
.A(n_2348),
.B(n_1897),
.Y(n_2361)
);

AND2x2_ASAP7_75t_L g2362 ( 
.A(n_2353),
.B(n_2129),
.Y(n_2362)
);

HB1xp67_ASAP7_75t_L g2363 ( 
.A(n_2354),
.Y(n_2363)
);

OAI22xp5_ASAP7_75t_L g2364 ( 
.A1(n_2358),
.A2(n_2350),
.B1(n_2356),
.B2(n_2100),
.Y(n_2364)
);

NAND3xp33_ASAP7_75t_SL g2365 ( 
.A(n_2360),
.B(n_1865),
.C(n_2062),
.Y(n_2365)
);

INVx1_ASAP7_75t_SL g2366 ( 
.A(n_2359),
.Y(n_2366)
);

INVx2_ASAP7_75t_L g2367 ( 
.A(n_2362),
.Y(n_2367)
);

INVx1_ASAP7_75t_L g2368 ( 
.A(n_2366),
.Y(n_2368)
);

AO22x2_ASAP7_75t_L g2369 ( 
.A1(n_2367),
.A2(n_2363),
.B1(n_2361),
.B2(n_2357),
.Y(n_2369)
);

AO22x2_ASAP7_75t_L g2370 ( 
.A1(n_2368),
.A2(n_2364),
.B1(n_2365),
.B2(n_2100),
.Y(n_2370)
);

INVx1_ASAP7_75t_L g2371 ( 
.A(n_2370),
.Y(n_2371)
);

AOI22xp5_ASAP7_75t_L g2372 ( 
.A1(n_2370),
.A2(n_2369),
.B1(n_2150),
.B2(n_2149),
.Y(n_2372)
);

OAI22xp5_ASAP7_75t_L g2373 ( 
.A1(n_2372),
.A2(n_2100),
.B1(n_2123),
.B2(n_2105),
.Y(n_2373)
);

OAI22xp5_ASAP7_75t_L g2374 ( 
.A1(n_2371),
.A2(n_2123),
.B1(n_2105),
.B2(n_2107),
.Y(n_2374)
);

OAI21xp5_ASAP7_75t_SL g2375 ( 
.A1(n_2373),
.A2(n_2017),
.B(n_1863),
.Y(n_2375)
);

AOI221xp5_ASAP7_75t_L g2376 ( 
.A1(n_2374),
.A2(n_2120),
.B1(n_2108),
.B2(n_2122),
.C(n_2123),
.Y(n_2376)
);

INVxp67_ASAP7_75t_L g2377 ( 
.A(n_2375),
.Y(n_2377)
);

AO21x2_ASAP7_75t_L g2378 ( 
.A1(n_2377),
.A2(n_2376),
.B(n_2122),
.Y(n_2378)
);

OAI22xp33_ASAP7_75t_L g2379 ( 
.A1(n_2378),
.A2(n_2040),
.B1(n_2047),
.B2(n_1863),
.Y(n_2379)
);

AOI32xp33_ASAP7_75t_L g2380 ( 
.A1(n_2379),
.A2(n_1863),
.A3(n_1862),
.B1(n_2150),
.B2(n_2149),
.Y(n_2380)
);

AOI211xp5_ASAP7_75t_L g2381 ( 
.A1(n_2380),
.A2(n_1857),
.B(n_1860),
.C(n_1853),
.Y(n_2381)
);


endmodule