module real_aes_58_n_104 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_103, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_104);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_103;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_104;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_185;
wire n_285;
wire n_624;
wire n_800;
wire n_618;
wire n_778;
wire n_522;
wire n_485;
wire n_822;
wire n_222;
wire n_750;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_421;
wire n_364;
wire n_555;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_551;
wire n_320;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_824;
wire n_467;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_535;
wire n_732;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_748;
wire n_781;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_504;
wire n_310;
wire n_455;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_454;
wire n_122;
wire n_812;
wire n_817;
wire n_565;
wire n_443;
wire n_782;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_449;
wire n_363;
wire n_417;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_527;
wire n_434;
wire n_502;
wire n_505;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_552;
wire n_402;
wire n_617;
wire n_733;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_807;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_288;
wire n_147;
wire n_150;
wire n_404;
wire n_598;
wire n_756;
wire n_735;
wire n_728;
wire n_713;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_810;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_765;
wire n_826;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_829;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_241;
wire n_175;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_802;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_798;
wire n_797;
wire n_237;
wire n_668;
NAND2xp5_ASAP7_75t_L g527 ( .A(n_0), .B(n_224), .Y(n_527) );
NAND2xp5_ASAP7_75t_L g113 ( .A(n_1), .B(n_114), .Y(n_113) );
INVx1_ASAP7_75t_L g158 ( .A(n_2), .Y(n_158) );
NAND2xp5_ASAP7_75t_L g549 ( .A(n_3), .B(n_530), .Y(n_549) );
NAND2xp33_ASAP7_75t_SL g520 ( .A(n_4), .B(n_179), .Y(n_520) );
NAND2xp5_ASAP7_75t_SL g215 ( .A(n_5), .B(n_192), .Y(n_215) );
INVx1_ASAP7_75t_L g512 ( .A(n_6), .Y(n_512) );
INVx1_ASAP7_75t_L g249 ( .A(n_7), .Y(n_249) );
CKINVDCx16_ASAP7_75t_R g114 ( .A(n_8), .Y(n_114) );
CKINVDCx5p33_ASAP7_75t_R g266 ( .A(n_9), .Y(n_266) );
AND2x2_ASAP7_75t_L g547 ( .A(n_10), .B(n_148), .Y(n_547) );
AOI22xp33_ASAP7_75t_SL g800 ( .A1(n_11), .A2(n_794), .B1(n_801), .B2(n_803), .Y(n_800) );
INVx2_ASAP7_75t_L g149 ( .A(n_12), .Y(n_149) );
CKINVDCx16_ASAP7_75t_R g115 ( .A(n_13), .Y(n_115) );
INVx1_ASAP7_75t_L g225 ( .A(n_14), .Y(n_225) );
AOI221x1_ASAP7_75t_L g515 ( .A1(n_15), .A2(n_181), .B1(n_516), .B2(n_518), .C(n_519), .Y(n_515) );
NAND2xp5_ASAP7_75t_SL g583 ( .A(n_16), .B(n_530), .Y(n_583) );
NOR2xp33_ASAP7_75t_SL g110 ( .A(n_17), .B(n_111), .Y(n_110) );
INVx1_ASAP7_75t_L g131 ( .A(n_17), .Y(n_131) );
INVx1_ASAP7_75t_L g222 ( .A(n_18), .Y(n_222) );
INVx1_ASAP7_75t_SL g170 ( .A(n_19), .Y(n_170) );
NAND2xp5_ASAP7_75t_SL g195 ( .A(n_20), .B(n_173), .Y(n_195) );
AOI33xp33_ASAP7_75t_L g240 ( .A1(n_21), .A2(n_48), .A3(n_155), .B1(n_166), .B2(n_241), .B3(n_242), .Y(n_240) );
AOI21xp5_ASAP7_75t_L g550 ( .A1(n_22), .A2(n_518), .B(n_551), .Y(n_550) );
NAND2xp5_ASAP7_75t_L g552 ( .A(n_23), .B(n_224), .Y(n_552) );
AOI221xp5_ASAP7_75t_SL g592 ( .A1(n_24), .A2(n_39), .B1(n_518), .B2(n_530), .C(n_593), .Y(n_592) );
INVx1_ASAP7_75t_L g259 ( .A(n_25), .Y(n_259) );
OR2x2_ASAP7_75t_L g150 ( .A(n_26), .B(n_91), .Y(n_150) );
OA21x2_ASAP7_75t_L g183 ( .A1(n_26), .A2(n_91), .B(n_149), .Y(n_183) );
INVxp67_ASAP7_75t_L g514 ( .A(n_27), .Y(n_514) );
NAND2xp5_ASAP7_75t_L g587 ( .A(n_28), .B(n_227), .Y(n_587) );
AND2x2_ASAP7_75t_L g541 ( .A(n_29), .B(n_147), .Y(n_541) );
NAND2xp5_ASAP7_75t_L g152 ( .A(n_30), .B(n_153), .Y(n_152) );
AOI21xp5_ASAP7_75t_L g525 ( .A1(n_31), .A2(n_518), .B(n_526), .Y(n_525) );
NAND2xp5_ASAP7_75t_L g594 ( .A(n_32), .B(n_227), .Y(n_594) );
AND2x2_ASAP7_75t_L g160 ( .A(n_33), .B(n_161), .Y(n_160) );
INVx1_ASAP7_75t_L g165 ( .A(n_33), .Y(n_165) );
AND2x2_ASAP7_75t_L g179 ( .A(n_33), .B(n_158), .Y(n_179) );
NOR3xp33_ASAP7_75t_L g112 ( .A(n_34), .B(n_113), .C(n_115), .Y(n_112) );
OR2x6_ASAP7_75t_L g129 ( .A(n_34), .B(n_130), .Y(n_129) );
CKINVDCx20_ASAP7_75t_R g261 ( .A(n_35), .Y(n_261) );
NAND2xp5_ASAP7_75t_L g286 ( .A(n_36), .B(n_153), .Y(n_286) );
AOI22xp5_ASAP7_75t_L g187 ( .A1(n_37), .A2(n_182), .B1(n_188), .B2(n_192), .Y(n_187) );
NAND2xp5_ASAP7_75t_L g196 ( .A(n_38), .B(n_197), .Y(n_196) );
AOI22xp5_ASAP7_75t_L g559 ( .A1(n_40), .A2(n_82), .B1(n_163), .B2(n_518), .Y(n_559) );
NAND2xp5_ASAP7_75t_L g172 ( .A(n_41), .B(n_173), .Y(n_172) );
NAND2xp5_ASAP7_75t_L g539 ( .A(n_42), .B(n_224), .Y(n_539) );
NAND2xp5_ASAP7_75t_SL g251 ( .A(n_43), .B(n_199), .Y(n_251) );
NAND2xp5_ASAP7_75t_L g250 ( .A(n_44), .B(n_173), .Y(n_250) );
CKINVDCx5p33_ASAP7_75t_R g191 ( .A(n_45), .Y(n_191) );
AND2x2_ASAP7_75t_L g531 ( .A(n_46), .B(n_147), .Y(n_531) );
NAND2xp5_ASAP7_75t_L g596 ( .A(n_47), .B(n_147), .Y(n_596) );
NAND2xp5_ASAP7_75t_L g290 ( .A(n_49), .B(n_173), .Y(n_290) );
CKINVDCx20_ASAP7_75t_R g438 ( .A(n_50), .Y(n_438) );
OAI22xp5_ASAP7_75t_L g818 ( .A1(n_50), .A2(n_62), .B1(n_438), .B2(n_819), .Y(n_818) );
INVx1_ASAP7_75t_L g156 ( .A(n_51), .Y(n_156) );
INVx1_ASAP7_75t_L g175 ( .A(n_51), .Y(n_175) );
AOI22x1_ASAP7_75t_L g794 ( .A1(n_52), .A2(n_795), .B1(n_796), .B2(n_797), .Y(n_794) );
CKINVDCx20_ASAP7_75t_R g795 ( .A(n_52), .Y(n_795) );
AND2x2_ASAP7_75t_L g291 ( .A(n_53), .B(n_147), .Y(n_291) );
AOI221xp5_ASAP7_75t_L g247 ( .A1(n_54), .A2(n_75), .B1(n_153), .B2(n_163), .C(n_248), .Y(n_247) );
NAND2xp5_ASAP7_75t_L g208 ( .A(n_55), .B(n_153), .Y(n_208) );
NAND2xp5_ASAP7_75t_SL g540 ( .A(n_56), .B(n_530), .Y(n_540) );
OAI21xp5_ASAP7_75t_L g805 ( .A1(n_57), .A2(n_806), .B(n_821), .Y(n_805) );
INVx1_ASAP7_75t_L g824 ( .A(n_57), .Y(n_824) );
NAND2xp5_ASAP7_75t_L g268 ( .A(n_58), .B(n_182), .Y(n_268) );
AOI21xp5_ASAP7_75t_SL g204 ( .A1(n_59), .A2(n_163), .B(n_205), .Y(n_204) );
AND2x2_ASAP7_75t_L g568 ( .A(n_60), .B(n_147), .Y(n_568) );
NAND2xp5_ASAP7_75t_L g528 ( .A(n_61), .B(n_227), .Y(n_528) );
CKINVDCx20_ASAP7_75t_R g819 ( .A(n_62), .Y(n_819) );
INVx1_ASAP7_75t_L g218 ( .A(n_63), .Y(n_218) );
NAND2xp5_ASAP7_75t_L g566 ( .A(n_64), .B(n_224), .Y(n_566) );
AND2x2_ASAP7_75t_SL g588 ( .A(n_65), .B(n_148), .Y(n_588) );
AOI21xp5_ASAP7_75t_L g536 ( .A1(n_66), .A2(n_518), .B(n_537), .Y(n_536) );
INVx1_ASAP7_75t_L g289 ( .A(n_67), .Y(n_289) );
NAND2xp5_ASAP7_75t_L g553 ( .A(n_68), .B(n_227), .Y(n_553) );
AND2x2_ASAP7_75t_SL g560 ( .A(n_69), .B(n_199), .Y(n_560) );
OAI22xp5_ASAP7_75t_L g797 ( .A1(n_70), .A2(n_103), .B1(n_798), .B2(n_799), .Y(n_797) );
CKINVDCx20_ASAP7_75t_R g798 ( .A(n_70), .Y(n_798) );
AOI21xp5_ASAP7_75t_L g287 ( .A1(n_71), .A2(n_163), .B(n_288), .Y(n_287) );
OAI22xp5_ASAP7_75t_L g816 ( .A1(n_72), .A2(n_817), .B1(n_818), .B2(n_820), .Y(n_816) );
CKINVDCx20_ASAP7_75t_R g817 ( .A(n_72), .Y(n_817) );
INVx1_ASAP7_75t_L g161 ( .A(n_73), .Y(n_161) );
INVx1_ASAP7_75t_L g177 ( .A(n_73), .Y(n_177) );
NAND2xp5_ASAP7_75t_L g243 ( .A(n_74), .B(n_153), .Y(n_243) );
AND2x2_ASAP7_75t_L g180 ( .A(n_76), .B(n_181), .Y(n_180) );
INVx1_ASAP7_75t_L g219 ( .A(n_77), .Y(n_219) );
AOI21xp5_ASAP7_75t_L g162 ( .A1(n_78), .A2(n_163), .B(n_169), .Y(n_162) );
A2O1A1Ixp33_ASAP7_75t_L g193 ( .A1(n_79), .A2(n_163), .B(n_194), .C(n_198), .Y(n_193) );
AOI22xp5_ASAP7_75t_L g558 ( .A1(n_80), .A2(n_85), .B1(n_153), .B2(n_530), .Y(n_558) );
NAND2xp5_ASAP7_75t_SL g567 ( .A(n_81), .B(n_530), .Y(n_567) );
INVx1_ASAP7_75t_L g111 ( .A(n_83), .Y(n_111) );
AND2x2_ASAP7_75t_SL g202 ( .A(n_84), .B(n_181), .Y(n_202) );
AOI22xp5_ASAP7_75t_L g237 ( .A1(n_86), .A2(n_163), .B1(n_238), .B2(n_239), .Y(n_237) );
NAND2xp5_ASAP7_75t_L g586 ( .A(n_87), .B(n_224), .Y(n_586) );
NAND2xp5_ASAP7_75t_L g595 ( .A(n_88), .B(n_224), .Y(n_595) );
CKINVDCx20_ASAP7_75t_R g829 ( .A(n_89), .Y(n_829) );
AOI21xp5_ASAP7_75t_L g563 ( .A1(n_90), .A2(n_518), .B(n_564), .Y(n_563) );
INVx1_ASAP7_75t_L g206 ( .A(n_92), .Y(n_206) );
NAND2xp5_ASAP7_75t_L g565 ( .A(n_93), .B(n_227), .Y(n_565) );
AND2x2_ASAP7_75t_L g244 ( .A(n_94), .B(n_181), .Y(n_244) );
A2O1A1Ixp33_ASAP7_75t_L g256 ( .A1(n_95), .A2(n_257), .B(n_258), .C(n_260), .Y(n_256) );
INVxp67_ASAP7_75t_L g517 ( .A(n_96), .Y(n_517) );
NAND2xp5_ASAP7_75t_L g529 ( .A(n_97), .B(n_530), .Y(n_529) );
NAND2xp5_ASAP7_75t_L g538 ( .A(n_98), .B(n_227), .Y(n_538) );
AOI21xp5_ASAP7_75t_L g584 ( .A1(n_99), .A2(n_518), .B(n_585), .Y(n_584) );
CKINVDCx20_ASAP7_75t_R g125 ( .A(n_100), .Y(n_125) );
BUFx2_ASAP7_75t_L g121 ( .A(n_101), .Y(n_121) );
NAND2xp5_ASAP7_75t_L g207 ( .A(n_102), .B(n_173), .Y(n_207) );
CKINVDCx20_ASAP7_75t_R g799 ( .A(n_103), .Y(n_799) );
AOI21xp33_ASAP7_75t_L g104 ( .A1(n_105), .A2(n_116), .B(n_828), .Y(n_104) );
CKINVDCx5p33_ASAP7_75t_R g105 ( .A(n_106), .Y(n_105) );
CKINVDCx20_ASAP7_75t_R g106 ( .A(n_107), .Y(n_106) );
NOR2xp67_ASAP7_75t_R g828 ( .A(n_107), .B(n_829), .Y(n_828) );
INVx2_ASAP7_75t_L g107 ( .A(n_108), .Y(n_107) );
INVx2_ASAP7_75t_L g108 ( .A(n_109), .Y(n_108) );
AND2x2_ASAP7_75t_SL g109 ( .A(n_110), .B(n_112), .Y(n_109) );
NAND2xp5_ASAP7_75t_L g130 ( .A(n_111), .B(n_131), .Y(n_130) );
NAND2xp5_ASAP7_75t_L g127 ( .A(n_115), .B(n_128), .Y(n_127) );
AND2x6_ASAP7_75t_SL g502 ( .A(n_115), .B(n_129), .Y(n_502) );
OR2x6_ASAP7_75t_SL g793 ( .A(n_115), .B(n_128), .Y(n_793) );
OR2x2_ASAP7_75t_L g804 ( .A(n_115), .B(n_129), .Y(n_804) );
OA22x2_ASAP7_75t_L g116 ( .A1(n_117), .A2(n_132), .B1(n_805), .B2(n_826), .Y(n_116) );
NAND2xp5_ASAP7_75t_L g117 ( .A(n_118), .B(n_122), .Y(n_117) );
CKINVDCx11_ASAP7_75t_R g118 ( .A(n_119), .Y(n_118) );
BUFx3_ASAP7_75t_L g827 ( .A(n_119), .Y(n_827) );
CKINVDCx20_ASAP7_75t_R g119 ( .A(n_120), .Y(n_119) );
HB1xp67_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
CKINVDCx16_ASAP7_75t_R g122 ( .A(n_123), .Y(n_122) );
HB1xp67_ASAP7_75t_L g123 ( .A(n_124), .Y(n_123) );
AOI21xp5_ASAP7_75t_L g821 ( .A1(n_124), .A2(n_822), .B(n_823), .Y(n_821) );
NOR2xp33_ASAP7_75t_L g124 ( .A(n_125), .B(n_126), .Y(n_124) );
INVx1_ASAP7_75t_L g825 ( .A(n_126), .Y(n_825) );
BUFx2_ASAP7_75t_L g126 ( .A(n_127), .Y(n_126) );
BUFx3_ASAP7_75t_L g809 ( .A(n_127), .Y(n_809) );
CKINVDCx5p33_ASAP7_75t_R g128 ( .A(n_129), .Y(n_128) );
OAI21xp5_ASAP7_75t_L g132 ( .A1(n_133), .A2(n_794), .B(n_800), .Y(n_132) );
INVxp67_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
OAI22x1_ASAP7_75t_L g134 ( .A1(n_135), .A2(n_501), .B1(n_503), .B2(n_791), .Y(n_134) );
INVx1_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
OAI22xp5_ASAP7_75t_L g801 ( .A1(n_136), .A2(n_501), .B1(n_504), .B2(n_802), .Y(n_801) );
AND3x1_ASAP7_75t_L g136 ( .A(n_137), .B(n_495), .C(n_498), .Y(n_136) );
NAND5xp2_ASAP7_75t_L g137 ( .A(n_138), .B(n_395), .C(n_425), .D(n_439), .E(n_465), .Y(n_137) );
INVx1_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
OAI21xp33_ASAP7_75t_L g495 ( .A1(n_139), .A2(n_438), .B(n_496), .Y(n_495) );
INVx1_ASAP7_75t_L g813 ( .A(n_139), .Y(n_813) );
NAND2xp5_ASAP7_75t_L g139 ( .A(n_140), .B(n_344), .Y(n_139) );
NOR3xp33_ASAP7_75t_SL g140 ( .A(n_141), .B(n_292), .C(n_326), .Y(n_140) );
A2O1A1Ixp33_ASAP7_75t_L g141 ( .A1(n_142), .A2(n_209), .B(n_231), .C(n_270), .Y(n_141) );
NAND2xp5_ASAP7_75t_L g142 ( .A(n_143), .B(n_184), .Y(n_142) );
BUFx2_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
NAND2xp5_ASAP7_75t_L g347 ( .A(n_144), .B(n_282), .Y(n_347) );
AND2x2_ASAP7_75t_L g434 ( .A(n_144), .B(n_212), .Y(n_434) );
HB1xp67_ASAP7_75t_L g144 ( .A(n_145), .Y(n_144) );
OR2x2_ASAP7_75t_L g230 ( .A(n_145), .B(n_201), .Y(n_230) );
INVx1_ASAP7_75t_L g272 ( .A(n_145), .Y(n_272) );
INVx2_ASAP7_75t_L g277 ( .A(n_145), .Y(n_277) );
HB1xp67_ASAP7_75t_L g305 ( .A(n_145), .Y(n_305) );
INVx1_ASAP7_75t_L g319 ( .A(n_145), .Y(n_319) );
AND2x2_ASAP7_75t_L g323 ( .A(n_145), .B(n_214), .Y(n_323) );
AND2x2_ASAP7_75t_L g404 ( .A(n_145), .B(n_213), .Y(n_404) );
AO21x2_ASAP7_75t_L g145 ( .A1(n_146), .A2(n_151), .B(n_180), .Y(n_145) );
AO21x2_ASAP7_75t_L g534 ( .A1(n_146), .A2(n_535), .B(n_541), .Y(n_534) );
AO21x2_ASAP7_75t_L g561 ( .A1(n_146), .A2(n_562), .B(n_568), .Y(n_561) );
AO21x2_ASAP7_75t_L g599 ( .A1(n_146), .A2(n_535), .B(n_541), .Y(n_599) );
CKINVDCx5p33_ASAP7_75t_R g146 ( .A(n_147), .Y(n_146) );
OA21x2_ASAP7_75t_L g591 ( .A1(n_147), .A2(n_592), .B(n_596), .Y(n_591) );
BUFx6f_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
AND2x2_ASAP7_75t_SL g148 ( .A(n_149), .B(n_150), .Y(n_148) );
AND2x4_ASAP7_75t_L g192 ( .A(n_149), .B(n_150), .Y(n_192) );
NAND2xp5_ASAP7_75t_L g151 ( .A(n_152), .B(n_162), .Y(n_151) );
INVx1_ASAP7_75t_L g269 ( .A(n_153), .Y(n_269) );
AOI22xp5_ASAP7_75t_L g510 ( .A1(n_153), .A2(n_163), .B1(n_511), .B2(n_513), .Y(n_510) );
AND2x4_ASAP7_75t_L g153 ( .A(n_154), .B(n_159), .Y(n_153) );
INVx1_ASAP7_75t_L g189 ( .A(n_154), .Y(n_189) );
AND2x2_ASAP7_75t_L g154 ( .A(n_155), .B(n_157), .Y(n_154) );
OR2x6_ASAP7_75t_L g171 ( .A(n_155), .B(n_167), .Y(n_171) );
INVxp33_ASAP7_75t_L g241 ( .A(n_155), .Y(n_241) );
INVx2_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
AND2x2_ASAP7_75t_L g168 ( .A(n_156), .B(n_158), .Y(n_168) );
AND2x4_ASAP7_75t_L g227 ( .A(n_156), .B(n_176), .Y(n_227) );
HB1xp67_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
INVx1_ASAP7_75t_L g190 ( .A(n_159), .Y(n_190) );
BUFx3_ASAP7_75t_L g159 ( .A(n_160), .Y(n_159) );
AND2x6_ASAP7_75t_L g518 ( .A(n_160), .B(n_168), .Y(n_518) );
INVx2_ASAP7_75t_L g167 ( .A(n_161), .Y(n_167) );
AND2x6_ASAP7_75t_L g224 ( .A(n_161), .B(n_174), .Y(n_224) );
INVxp67_ASAP7_75t_L g267 ( .A(n_163), .Y(n_267) );
AND2x4_ASAP7_75t_L g163 ( .A(n_164), .B(n_168), .Y(n_163) );
NOR2x1p5_ASAP7_75t_L g164 ( .A(n_165), .B(n_166), .Y(n_164) );
INVx1_ASAP7_75t_L g242 ( .A(n_166), .Y(n_242) );
INVx3_ASAP7_75t_L g166 ( .A(n_167), .Y(n_166) );
O2A1O1Ixp33_ASAP7_75t_SL g169 ( .A1(n_170), .A2(n_171), .B(n_172), .C(n_178), .Y(n_169) );
INVx2_ASAP7_75t_L g197 ( .A(n_171), .Y(n_197) );
O2A1O1Ixp33_ASAP7_75t_L g205 ( .A1(n_171), .A2(n_178), .B(n_206), .C(n_207), .Y(n_205) );
OAI22xp5_ASAP7_75t_L g217 ( .A1(n_171), .A2(n_218), .B1(n_219), .B2(n_220), .Y(n_217) );
O2A1O1Ixp33_ASAP7_75t_SL g248 ( .A1(n_171), .A2(n_178), .B(n_249), .C(n_250), .Y(n_248) );
INVxp67_ASAP7_75t_L g257 ( .A(n_171), .Y(n_257) );
O2A1O1Ixp33_ASAP7_75t_L g288 ( .A1(n_171), .A2(n_178), .B(n_289), .C(n_290), .Y(n_288) );
INVx1_ASAP7_75t_L g220 ( .A(n_173), .Y(n_220) );
AND2x4_ASAP7_75t_L g530 ( .A(n_173), .B(n_179), .Y(n_530) );
AND2x4_ASAP7_75t_L g173 ( .A(n_174), .B(n_176), .Y(n_173) );
INVx2_ASAP7_75t_L g174 ( .A(n_175), .Y(n_174) );
INVx2_ASAP7_75t_L g176 ( .A(n_177), .Y(n_176) );
AOI21xp5_ASAP7_75t_L g194 ( .A1(n_178), .A2(n_195), .B(n_196), .Y(n_194) );
NOR2xp33_ASAP7_75t_L g228 ( .A(n_178), .B(n_192), .Y(n_228) );
INVx1_ASAP7_75t_L g238 ( .A(n_178), .Y(n_238) );
AOI21xp5_ASAP7_75t_L g526 ( .A1(n_178), .A2(n_527), .B(n_528), .Y(n_526) );
AOI21xp5_ASAP7_75t_L g537 ( .A1(n_178), .A2(n_538), .B(n_539), .Y(n_537) );
AOI21xp5_ASAP7_75t_L g551 ( .A1(n_178), .A2(n_552), .B(n_553), .Y(n_551) );
AOI21xp5_ASAP7_75t_L g564 ( .A1(n_178), .A2(n_565), .B(n_566), .Y(n_564) );
AOI21xp5_ASAP7_75t_L g585 ( .A1(n_178), .A2(n_586), .B(n_587), .Y(n_585) );
AOI21xp5_ASAP7_75t_L g593 ( .A1(n_178), .A2(n_594), .B(n_595), .Y(n_593) );
INVx5_ASAP7_75t_L g178 ( .A(n_179), .Y(n_178) );
HB1xp67_ASAP7_75t_L g260 ( .A(n_179), .Y(n_260) );
OAI22xp5_ASAP7_75t_L g255 ( .A1(n_181), .A2(n_256), .B1(n_261), .B2(n_262), .Y(n_255) );
INVx3_ASAP7_75t_L g262 ( .A(n_181), .Y(n_262) );
INVx4_ASAP7_75t_L g181 ( .A(n_182), .Y(n_181) );
NAND2xp5_ASAP7_75t_L g264 ( .A(n_182), .B(n_265), .Y(n_264) );
AOI21x1_ASAP7_75t_L g523 ( .A1(n_182), .A2(n_524), .B(n_531), .Y(n_523) );
INVx3_ASAP7_75t_L g182 ( .A(n_183), .Y(n_182) );
BUFx4f_ASAP7_75t_L g199 ( .A(n_183), .Y(n_199) );
AND2x4_ASAP7_75t_SL g184 ( .A(n_185), .B(n_200), .Y(n_184) );
HB1xp67_ASAP7_75t_L g185 ( .A(n_186), .Y(n_185) );
INVx2_ASAP7_75t_L g229 ( .A(n_186), .Y(n_229) );
AND2x2_ASAP7_75t_L g273 ( .A(n_186), .B(n_214), .Y(n_273) );
AND2x2_ASAP7_75t_L g294 ( .A(n_186), .B(n_201), .Y(n_294) );
INVx1_ASAP7_75t_L g317 ( .A(n_186), .Y(n_317) );
AND2x4_ASAP7_75t_L g384 ( .A(n_186), .B(n_213), .Y(n_384) );
AND2x2_ASAP7_75t_L g186 ( .A(n_187), .B(n_193), .Y(n_186) );
NOR3xp33_ASAP7_75t_L g188 ( .A(n_189), .B(n_190), .C(n_191), .Y(n_188) );
AOI21xp5_ASAP7_75t_L g203 ( .A1(n_192), .A2(n_204), .B(n_208), .Y(n_203) );
NOR2xp33_ASAP7_75t_L g511 ( .A(n_192), .B(n_512), .Y(n_511) );
NOR2xp33_ASAP7_75t_L g513 ( .A(n_192), .B(n_514), .Y(n_513) );
NOR2xp33_ASAP7_75t_L g516 ( .A(n_192), .B(n_517), .Y(n_516) );
NOR3xp33_ASAP7_75t_L g519 ( .A(n_192), .B(n_220), .C(n_520), .Y(n_519) );
AOI21xp5_ASAP7_75t_L g548 ( .A1(n_192), .A2(n_549), .B(n_550), .Y(n_548) );
AO21x2_ASAP7_75t_L g235 ( .A1(n_198), .A2(n_236), .B(n_244), .Y(n_235) );
AO21x2_ASAP7_75t_L g299 ( .A1(n_198), .A2(n_236), .B(n_244), .Y(n_299) );
AOI21x1_ASAP7_75t_L g556 ( .A1(n_198), .A2(n_557), .B(n_560), .Y(n_556) );
INVx2_ASAP7_75t_SL g198 ( .A(n_199), .Y(n_198) );
OA21x2_ASAP7_75t_L g246 ( .A1(n_199), .A2(n_247), .B(n_251), .Y(n_246) );
AOI21xp5_ASAP7_75t_L g582 ( .A1(n_199), .A2(n_583), .B(n_584), .Y(n_582) );
AND2x4_ASAP7_75t_L g400 ( .A(n_200), .B(n_317), .Y(n_400) );
OR2x2_ASAP7_75t_L g441 ( .A(n_200), .B(n_442), .Y(n_441) );
NOR2xp67_ASAP7_75t_SL g460 ( .A(n_200), .B(n_333), .Y(n_460) );
NOR2x1_ASAP7_75t_L g478 ( .A(n_200), .B(n_392), .Y(n_478) );
INVx4_ASAP7_75t_L g200 ( .A(n_201), .Y(n_200) );
NOR2x1_ASAP7_75t_SL g278 ( .A(n_201), .B(n_214), .Y(n_278) );
AND2x4_ASAP7_75t_L g316 ( .A(n_201), .B(n_317), .Y(n_316) );
BUFx6f_ASAP7_75t_L g322 ( .A(n_201), .Y(n_322) );
NAND2xp5_ASAP7_75t_L g354 ( .A(n_201), .B(n_276), .Y(n_354) );
INVx2_ASAP7_75t_L g368 ( .A(n_201), .Y(n_368) );
NAND2xp5_ASAP7_75t_SL g390 ( .A(n_201), .B(n_320), .Y(n_390) );
AND2x2_ASAP7_75t_L g482 ( .A(n_201), .B(n_340), .Y(n_482) );
OR2x6_ASAP7_75t_L g201 ( .A(n_202), .B(n_203), .Y(n_201) );
INVx1_ASAP7_75t_L g209 ( .A(n_210), .Y(n_209) );
NOR2x1_ASAP7_75t_L g210 ( .A(n_211), .B(n_230), .Y(n_210) );
INVx2_ASAP7_75t_L g211 ( .A(n_212), .Y(n_211) );
NAND2xp5_ASAP7_75t_L g333 ( .A(n_212), .B(n_319), .Y(n_333) );
AND2x2_ASAP7_75t_SL g342 ( .A(n_212), .B(n_322), .Y(n_342) );
AND2x2_ASAP7_75t_L g212 ( .A(n_213), .B(n_229), .Y(n_212) );
INVx1_ASAP7_75t_L g320 ( .A(n_213), .Y(n_320) );
INVx3_ASAP7_75t_L g213 ( .A(n_214), .Y(n_213) );
INVx2_ASAP7_75t_L g340 ( .A(n_214), .Y(n_340) );
AND2x4_ASAP7_75t_L g214 ( .A(n_215), .B(n_216), .Y(n_214) );
OAI21xp5_ASAP7_75t_L g216 ( .A1(n_217), .A2(n_221), .B(n_228), .Y(n_216) );
NOR2xp33_ASAP7_75t_L g258 ( .A(n_220), .B(n_259), .Y(n_258) );
OAI22xp5_ASAP7_75t_L g221 ( .A1(n_222), .A2(n_223), .B1(n_225), .B2(n_226), .Y(n_221) );
INVxp67_ASAP7_75t_L g223 ( .A(n_224), .Y(n_223) );
INVxp67_ASAP7_75t_L g226 ( .A(n_227), .Y(n_226) );
INVx1_ASAP7_75t_L g373 ( .A(n_229), .Y(n_373) );
INVx2_ASAP7_75t_SL g418 ( .A(n_230), .Y(n_418) );
INVx1_ASAP7_75t_L g231 ( .A(n_232), .Y(n_231) );
AND2x2_ASAP7_75t_L g232 ( .A(n_233), .B(n_252), .Y(n_232) );
NAND2x1p5_ASAP7_75t_L g327 ( .A(n_233), .B(n_328), .Y(n_327) );
BUFx2_ASAP7_75t_L g364 ( .A(n_233), .Y(n_364) );
AND2x2_ASAP7_75t_L g488 ( .A(n_233), .B(n_313), .Y(n_488) );
AND2x2_ASAP7_75t_L g233 ( .A(n_234), .B(n_245), .Y(n_233) );
AND2x4_ASAP7_75t_L g301 ( .A(n_234), .B(n_283), .Y(n_301) );
INVx1_ASAP7_75t_L g312 ( .A(n_234), .Y(n_312) );
AND2x2_ASAP7_75t_L g343 ( .A(n_234), .B(n_298), .Y(n_343) );
INVx2_ASAP7_75t_L g234 ( .A(n_235), .Y(n_234) );
NAND2xp5_ASAP7_75t_L g337 ( .A(n_235), .B(n_246), .Y(n_337) );
NAND2xp5_ASAP7_75t_L g375 ( .A(n_235), .B(n_284), .Y(n_375) );
NAND2xp5_ASAP7_75t_SL g236 ( .A(n_237), .B(n_243), .Y(n_236) );
INVx1_ASAP7_75t_L g239 ( .A(n_240), .Y(n_239) );
INVxp67_ASAP7_75t_L g245 ( .A(n_246), .Y(n_245) );
INVx2_ASAP7_75t_L g281 ( .A(n_246), .Y(n_281) );
AND2x4_ASAP7_75t_L g349 ( .A(n_246), .B(n_350), .Y(n_349) );
INVx1_ASAP7_75t_L g361 ( .A(n_246), .Y(n_361) );
INVx1_ASAP7_75t_L g403 ( .A(n_246), .Y(n_403) );
HB1xp67_ASAP7_75t_L g415 ( .A(n_246), .Y(n_415) );
AND2x2_ASAP7_75t_L g431 ( .A(n_246), .B(n_254), .Y(n_431) );
BUFx2_ASAP7_75t_L g252 ( .A(n_253), .Y(n_252) );
AND2x2_ASAP7_75t_L g378 ( .A(n_253), .B(n_336), .Y(n_378) );
INVx1_ASAP7_75t_SL g380 ( .A(n_253), .Y(n_380) );
AND2x2_ASAP7_75t_L g401 ( .A(n_253), .B(n_402), .Y(n_401) );
INVx1_ASAP7_75t_L g253 ( .A(n_254), .Y(n_253) );
AND2x4_ASAP7_75t_L g280 ( .A(n_254), .B(n_281), .Y(n_280) );
INVx1_ASAP7_75t_L g308 ( .A(n_254), .Y(n_308) );
INVx2_ASAP7_75t_L g314 ( .A(n_254), .Y(n_314) );
NAND2xp5_ASAP7_75t_L g329 ( .A(n_254), .B(n_284), .Y(n_329) );
OR2x2_ASAP7_75t_L g254 ( .A(n_255), .B(n_263), .Y(n_254) );
AO21x2_ASAP7_75t_L g284 ( .A1(n_262), .A2(n_285), .B(n_291), .Y(n_284) );
AO21x2_ASAP7_75t_L g298 ( .A1(n_262), .A2(n_285), .B(n_291), .Y(n_298) );
OAI22xp5_ASAP7_75t_L g263 ( .A1(n_264), .A2(n_267), .B1(n_268), .B2(n_269), .Y(n_263) );
INVx1_ASAP7_75t_L g265 ( .A(n_266), .Y(n_265) );
OAI21xp5_ASAP7_75t_L g270 ( .A1(n_271), .A2(n_274), .B(n_279), .Y(n_270) );
INVx1_ASAP7_75t_L g410 ( .A(n_271), .Y(n_410) );
AND2x2_ASAP7_75t_L g271 ( .A(n_272), .B(n_273), .Y(n_271) );
INVx2_ASAP7_75t_L g330 ( .A(n_273), .Y(n_330) );
AND2x2_ASAP7_75t_L g386 ( .A(n_273), .B(n_322), .Y(n_386) );
AND2x2_ASAP7_75t_L g274 ( .A(n_275), .B(n_278), .Y(n_274) );
INVx1_ASAP7_75t_L g300 ( .A(n_275), .Y(n_300) );
NAND2xp5_ASAP7_75t_L g362 ( .A(n_275), .B(n_316), .Y(n_362) );
NOR2xp33_ASAP7_75t_L g391 ( .A(n_275), .B(n_392), .Y(n_391) );
AND2x2_ASAP7_75t_L g407 ( .A(n_275), .B(n_400), .Y(n_407) );
AND2x2_ASAP7_75t_L g481 ( .A(n_275), .B(n_482), .Y(n_481) );
INVx3_ASAP7_75t_L g275 ( .A(n_276), .Y(n_275) );
HB1xp67_ASAP7_75t_L g469 ( .A(n_276), .Y(n_469) );
INVx2_ASAP7_75t_L g276 ( .A(n_277), .Y(n_276) );
HB1xp67_ASAP7_75t_L g389 ( .A(n_277), .Y(n_389) );
AND2x2_ASAP7_75t_L g302 ( .A(n_278), .B(n_303), .Y(n_302) );
OAI21xp33_ASAP7_75t_L g490 ( .A1(n_278), .A2(n_491), .B(n_493), .Y(n_490) );
AND2x2_ASAP7_75t_L g279 ( .A(n_280), .B(n_282), .Y(n_279) );
INVx3_ASAP7_75t_L g376 ( .A(n_280), .Y(n_376) );
NAND2x1_ASAP7_75t_SL g420 ( .A(n_280), .B(n_421), .Y(n_420) );
AND2x2_ASAP7_75t_L g423 ( .A(n_280), .B(n_301), .Y(n_423) );
AND2x2_ASAP7_75t_L g335 ( .A(n_282), .B(n_336), .Y(n_335) );
OR2x2_ASAP7_75t_L g472 ( .A(n_282), .B(n_473), .Y(n_472) );
AND2x2_ASAP7_75t_L g483 ( .A(n_282), .B(n_431), .Y(n_483) );
INVx3_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
NAND2x1p5_ASAP7_75t_L g359 ( .A(n_283), .B(n_360), .Y(n_359) );
INVx3_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
AND2x2_ASAP7_75t_L g414 ( .A(n_284), .B(n_415), .Y(n_414) );
NAND2xp5_ASAP7_75t_L g285 ( .A(n_286), .B(n_287), .Y(n_285) );
OAI21xp5_ASAP7_75t_SL g292 ( .A1(n_293), .A2(n_306), .B(n_309), .Y(n_292) );
AOI22xp5_ASAP7_75t_L g293 ( .A1(n_294), .A2(n_295), .B1(n_301), .B2(n_302), .Y(n_293) );
HB1xp67_ASAP7_75t_L g351 ( .A(n_294), .Y(n_351) );
AND2x2_ASAP7_75t_L g295 ( .A(n_296), .B(n_300), .Y(n_295) );
AND2x2_ASAP7_75t_L g324 ( .A(n_296), .B(n_325), .Y(n_324) );
AND2x2_ASAP7_75t_L g430 ( .A(n_296), .B(n_431), .Y(n_430) );
AOI22xp5_ASAP7_75t_L g448 ( .A1(n_296), .A2(n_449), .B1(n_450), .B2(n_451), .Y(n_448) );
NAND2xp5_ASAP7_75t_L g456 ( .A(n_296), .B(n_457), .Y(n_456) );
AND2x4_ASAP7_75t_L g296 ( .A(n_297), .B(n_299), .Y(n_296) );
INVx2_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
AND2x2_ASAP7_75t_L g313 ( .A(n_298), .B(n_314), .Y(n_313) );
NOR2xp67_ASAP7_75t_L g394 ( .A(n_298), .B(n_314), .Y(n_394) );
NOR2x1_ASAP7_75t_L g402 ( .A(n_298), .B(n_403), .Y(n_402) );
INVx2_ASAP7_75t_L g350 ( .A(n_299), .Y(n_350) );
AND2x2_ASAP7_75t_L g358 ( .A(n_299), .B(n_314), .Y(n_358) );
INVx1_ASAP7_75t_L g421 ( .A(n_299), .Y(n_421) );
INVx1_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
NAND2x1_ASAP7_75t_L g339 ( .A(n_304), .B(n_340), .Y(n_339) );
INVx1_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
INVx1_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
AND2x2_ASAP7_75t_L g451 ( .A(n_307), .B(n_336), .Y(n_451) );
INVx1_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
INVx2_ASAP7_75t_L g325 ( .A(n_308), .Y(n_325) );
AND2x2_ASAP7_75t_L g348 ( .A(n_308), .B(n_349), .Y(n_348) );
AND2x2_ASAP7_75t_L g436 ( .A(n_308), .B(n_343), .Y(n_436) );
AOI22xp5_ASAP7_75t_L g309 ( .A1(n_310), .A2(n_315), .B1(n_321), .B2(n_324), .Y(n_309) );
INVx1_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
OR2x2_ASAP7_75t_L g444 ( .A(n_311), .B(n_445), .Y(n_444) );
NAND2x1p5_ASAP7_75t_L g311 ( .A(n_312), .B(n_313), .Y(n_311) );
AND2x2_ASAP7_75t_L g474 ( .A(n_314), .B(n_361), .Y(n_474) );
AND2x2_ASAP7_75t_SL g315 ( .A(n_316), .B(n_318), .Y(n_315) );
INVx2_ASAP7_75t_L g341 ( .A(n_316), .Y(n_341) );
OAI21xp33_ASAP7_75t_SL g487 ( .A1(n_316), .A2(n_488), .B(n_489), .Y(n_487) );
AND2x4_ASAP7_75t_SL g318 ( .A(n_319), .B(n_320), .Y(n_318) );
HB1xp67_ASAP7_75t_L g477 ( .A(n_319), .Y(n_477) );
AND2x2_ASAP7_75t_L g321 ( .A(n_322), .B(n_323), .Y(n_321) );
O2A1O1Ixp33_ASAP7_75t_SL g419 ( .A1(n_322), .A2(n_420), .B(n_422), .C(n_424), .Y(n_419) );
AND2x2_ASAP7_75t_SL g371 ( .A(n_323), .B(n_372), .Y(n_371) );
INVx1_ASAP7_75t_L g424 ( .A(n_323), .Y(n_424) );
NAND2xp5_ASAP7_75t_L g464 ( .A(n_323), .B(n_400), .Y(n_464) );
INVx1_ASAP7_75t_SL g331 ( .A(n_324), .Y(n_331) );
AND2x2_ASAP7_75t_L g412 ( .A(n_325), .B(n_349), .Y(n_412) );
INVx1_ASAP7_75t_L g457 ( .A(n_325), .Y(n_457) );
OAI221xp5_ASAP7_75t_L g326 ( .A1(n_327), .A2(n_330), .B1(n_331), .B2(n_332), .C(n_334), .Y(n_326) );
HB1xp67_ASAP7_75t_L g446 ( .A(n_327), .Y(n_446) );
INVx2_ASAP7_75t_SL g328 ( .A(n_329), .Y(n_328) );
OR2x2_ASAP7_75t_L g494 ( .A(n_329), .B(n_337), .Y(n_494) );
OR2x2_ASAP7_75t_L g353 ( .A(n_330), .B(n_354), .Y(n_353) );
NOR2x1_ASAP7_75t_L g366 ( .A(n_330), .B(n_367), .Y(n_366) );
NOR2xp33_ASAP7_75t_L g453 ( .A(n_330), .B(n_454), .Y(n_453) );
OR2x2_ASAP7_75t_L g492 ( .A(n_330), .B(n_389), .Y(n_492) );
BUFx2_ASAP7_75t_L g332 ( .A(n_333), .Y(n_332) );
AOI32xp33_ASAP7_75t_L g334 ( .A1(n_335), .A2(n_338), .A3(n_341), .B1(n_342), .B2(n_343), .Y(n_334) );
INVx1_ASAP7_75t_L g355 ( .A(n_336), .Y(n_355) );
INVx2_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
NOR2xp33_ASAP7_75t_L g398 ( .A(n_338), .B(n_399), .Y(n_398) );
INVx2_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
INVx1_ASAP7_75t_L g450 ( .A(n_339), .Y(n_450) );
OAI22xp33_ASAP7_75t_SL g432 ( .A1(n_341), .A2(n_433), .B1(n_435), .B2(n_437), .Y(n_432) );
INVx1_ASAP7_75t_L g463 ( .A(n_342), .Y(n_463) );
AOI211x1_ASAP7_75t_L g344 ( .A1(n_345), .A2(n_351), .B(n_352), .C(n_369), .Y(n_344) );
AND2x2_ASAP7_75t_L g345 ( .A(n_346), .B(n_348), .Y(n_345) );
NAND2xp5_ASAP7_75t_L g437 ( .A(n_346), .B(n_431), .Y(n_437) );
INVx1_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
AND2x4_ASAP7_75t_L g393 ( .A(n_349), .B(n_394), .Y(n_393) );
INVx1_ASAP7_75t_L g459 ( .A(n_349), .Y(n_459) );
OAI222xp33_ASAP7_75t_L g352 ( .A1(n_353), .A2(n_355), .B1(n_356), .B2(n_362), .C1(n_363), .C2(n_365), .Y(n_352) );
INVxp67_ASAP7_75t_L g449 ( .A(n_353), .Y(n_449) );
OR2x2_ASAP7_75t_L g356 ( .A(n_357), .B(n_359), .Y(n_356) );
NOR2xp33_ASAP7_75t_L g489 ( .A(n_357), .B(n_442), .Y(n_489) );
INVx1_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
AND2x2_ASAP7_75t_L g405 ( .A(n_358), .B(n_402), .Y(n_405) );
INVx3_ASAP7_75t_L g445 ( .A(n_360), .Y(n_445) );
BUFx3_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
INVx1_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
INVx1_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
INVx1_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
AND2x2_ASAP7_75t_L g383 ( .A(n_368), .B(n_384), .Y(n_383) );
OAI221xp5_ASAP7_75t_L g369 ( .A1(n_370), .A2(n_374), .B1(n_377), .B2(n_382), .C(n_385), .Y(n_369) );
INVx1_ASAP7_75t_SL g370 ( .A(n_371), .Y(n_370) );
OAI21xp5_ASAP7_75t_L g427 ( .A1(n_371), .A2(n_428), .B(n_430), .Y(n_427) );
INVx2_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
OR2x2_ASAP7_75t_L g374 ( .A(n_375), .B(n_376), .Y(n_374) );
INVx1_ASAP7_75t_L g381 ( .A(n_375), .Y(n_381) );
OR2x2_ASAP7_75t_L g485 ( .A(n_376), .B(n_421), .Y(n_485) );
NOR2xp67_ASAP7_75t_L g377 ( .A(n_378), .B(n_379), .Y(n_377) );
NAND2xp5_ASAP7_75t_L g406 ( .A(n_379), .B(n_407), .Y(n_406) );
AND2x2_ASAP7_75t_L g379 ( .A(n_380), .B(n_381), .Y(n_379) );
OAI21xp5_ASAP7_75t_L g479 ( .A1(n_382), .A2(n_411), .B(n_480), .Y(n_479) );
INVx1_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
OAI21xp5_ASAP7_75t_L g461 ( .A1(n_383), .A2(n_455), .B(n_462), .Y(n_461) );
INVx4_ASAP7_75t_L g392 ( .A(n_384), .Y(n_392) );
OAI31xp33_ASAP7_75t_SL g385 ( .A1(n_386), .A2(n_387), .A3(n_391), .B(n_393), .Y(n_385) );
INVx1_ASAP7_75t_L g443 ( .A(n_387), .Y(n_443) );
NOR2x1_ASAP7_75t_L g387 ( .A(n_388), .B(n_390), .Y(n_387) );
INVx1_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
INVx2_ASAP7_75t_L g417 ( .A(n_392), .Y(n_417) );
AND2x2_ASAP7_75t_L g395 ( .A(n_396), .B(n_408), .Y(n_395) );
NAND4xp25_ASAP7_75t_L g496 ( .A(n_396), .B(n_408), .C(n_427), .D(n_497), .Y(n_496) );
AND2x2_ASAP7_75t_L g396 ( .A(n_397), .B(n_406), .Y(n_396) );
AOI22xp5_ASAP7_75t_L g397 ( .A1(n_398), .A2(n_401), .B1(n_404), .B2(n_405), .Y(n_397) );
INVx1_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
AND2x2_ASAP7_75t_L g468 ( .A(n_400), .B(n_469), .Y(n_468) );
NAND2xp5_ASAP7_75t_L g429 ( .A(n_401), .B(n_421), .Y(n_429) );
INVx1_ASAP7_75t_SL g442 ( .A(n_404), .Y(n_442) );
NOR2xp33_ASAP7_75t_L g408 ( .A(n_409), .B(n_419), .Y(n_408) );
OAI22xp5_ASAP7_75t_L g409 ( .A1(n_410), .A2(n_411), .B1(n_413), .B2(n_416), .Y(n_409) );
INVx3_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
INVxp67_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
NAND2x1_ASAP7_75t_L g416 ( .A(n_417), .B(n_418), .Y(n_416) );
AOI22xp5_ASAP7_75t_L g480 ( .A1(n_418), .A2(n_481), .B1(n_483), .B2(n_484), .Y(n_480) );
INVx2_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
NOR3xp33_ASAP7_75t_L g425 ( .A(n_426), .B(n_432), .C(n_438), .Y(n_425) );
INVxp67_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
INVx1_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
INVx1_ASAP7_75t_L g497 ( .A(n_432), .Y(n_497) );
INVx2_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
INVx1_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
OAI21xp33_ASAP7_75t_L g498 ( .A1(n_438), .A2(n_499), .B(n_500), .Y(n_498) );
INVxp33_ASAP7_75t_L g499 ( .A(n_439), .Y(n_499) );
AND2x2_ASAP7_75t_L g812 ( .A(n_439), .B(n_465), .Y(n_812) );
NOR2xp67_ASAP7_75t_L g439 ( .A(n_440), .B(n_447), .Y(n_439) );
AOI22xp33_ASAP7_75t_L g440 ( .A1(n_441), .A2(n_443), .B1(n_444), .B2(n_446), .Y(n_440) );
OAI21xp5_ASAP7_75t_L g466 ( .A1(n_444), .A2(n_467), .B(n_470), .Y(n_466) );
INVx2_ASAP7_75t_L g454 ( .A(n_445), .Y(n_454) );
NAND3xp33_ASAP7_75t_SL g447 ( .A(n_448), .B(n_452), .C(n_461), .Y(n_447) );
AOI22xp5_ASAP7_75t_L g452 ( .A1(n_453), .A2(n_455), .B1(n_458), .B2(n_460), .Y(n_452) );
INVx1_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
INVx1_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
NAND2xp5_ASAP7_75t_L g462 ( .A(n_463), .B(n_464), .Y(n_462) );
INVxp33_ASAP7_75t_SL g500 ( .A(n_465), .Y(n_500) );
NOR3x1_ASAP7_75t_L g465 ( .A(n_466), .B(n_479), .C(n_486), .Y(n_465) );
INVx1_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
NAND2xp5_ASAP7_75t_L g470 ( .A(n_471), .B(n_475), .Y(n_470) );
INVx1_ASAP7_75t_L g471 ( .A(n_472), .Y(n_471) );
INVx2_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
INVx1_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
NAND2xp5_ASAP7_75t_L g476 ( .A(n_477), .B(n_478), .Y(n_476) );
INVx1_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
NAND2xp5_ASAP7_75t_SL g486 ( .A(n_487), .B(n_490), .Y(n_486) );
INVx1_ASAP7_75t_L g491 ( .A(n_492), .Y(n_491) );
INVx1_ASAP7_75t_SL g493 ( .A(n_494), .Y(n_493) );
INVx1_ASAP7_75t_L g814 ( .A(n_496), .Y(n_814) );
CKINVDCx11_ASAP7_75t_R g501 ( .A(n_502), .Y(n_501) );
INVx3_ASAP7_75t_L g503 ( .A(n_504), .Y(n_503) );
AND2x4_ASAP7_75t_L g504 ( .A(n_505), .B(n_668), .Y(n_504) );
NOR4xp25_ASAP7_75t_L g505 ( .A(n_506), .B(n_611), .C(n_650), .D(n_657), .Y(n_505) );
OAI221xp5_ASAP7_75t_L g506 ( .A1(n_507), .A2(n_532), .B1(n_569), .B2(n_578), .C(n_597), .Y(n_506) );
OR2x2_ASAP7_75t_L g741 ( .A(n_507), .B(n_603), .Y(n_741) );
INVx1_ASAP7_75t_L g507 ( .A(n_508), .Y(n_507) );
AND2x2_ASAP7_75t_L g656 ( .A(n_508), .B(n_581), .Y(n_656) );
NAND2xp5_ASAP7_75t_L g675 ( .A(n_508), .B(n_676), .Y(n_675) );
AND2x2_ASAP7_75t_SL g721 ( .A(n_508), .B(n_722), .Y(n_721) );
AND2x4_ASAP7_75t_L g508 ( .A(n_509), .B(n_521), .Y(n_508) );
AND2x4_ASAP7_75t_SL g580 ( .A(n_509), .B(n_581), .Y(n_580) );
INVx3_ASAP7_75t_L g602 ( .A(n_509), .Y(n_602) );
AND2x2_ASAP7_75t_L g637 ( .A(n_509), .B(n_610), .Y(n_637) );
NAND2xp5_ASAP7_75t_L g651 ( .A(n_509), .B(n_522), .Y(n_651) );
NAND2xp5_ASAP7_75t_L g689 ( .A(n_509), .B(n_604), .Y(n_689) );
OR2x2_ASAP7_75t_L g767 ( .A(n_509), .B(n_581), .Y(n_767) );
AND2x4_ASAP7_75t_L g509 ( .A(n_510), .B(n_515), .Y(n_509) );
INVx2_ASAP7_75t_L g521 ( .A(n_522), .Y(n_521) );
AND2x2_ASAP7_75t_L g589 ( .A(n_522), .B(n_590), .Y(n_589) );
NAND2xp5_ASAP7_75t_L g609 ( .A(n_522), .B(n_610), .Y(n_609) );
INVx1_ASAP7_75t_L g615 ( .A(n_522), .Y(n_615) );
OR2x2_ASAP7_75t_L g620 ( .A(n_522), .B(n_604), .Y(n_620) );
AND2x2_ASAP7_75t_L g633 ( .A(n_522), .B(n_591), .Y(n_633) );
HB1xp67_ASAP7_75t_L g636 ( .A(n_522), .Y(n_636) );
INVx1_ASAP7_75t_L g648 ( .A(n_522), .Y(n_648) );
NAND2xp5_ASAP7_75t_L g713 ( .A(n_522), .B(n_602), .Y(n_713) );
INVx3_ASAP7_75t_L g522 ( .A(n_523), .Y(n_522) );
NAND2xp5_ASAP7_75t_L g524 ( .A(n_525), .B(n_529), .Y(n_524) );
NAND2xp5_ASAP7_75t_SL g532 ( .A(n_533), .B(n_542), .Y(n_532) );
HB1xp67_ASAP7_75t_L g533 ( .A(n_534), .Y(n_533) );
OR2x2_ASAP7_75t_L g577 ( .A(n_534), .B(n_561), .Y(n_577) );
AND2x4_ASAP7_75t_L g607 ( .A(n_534), .B(n_546), .Y(n_607) );
INVx2_ASAP7_75t_L g641 ( .A(n_534), .Y(n_641) );
NAND2xp5_ASAP7_75t_L g699 ( .A(n_534), .B(n_561), .Y(n_699) );
AND2x2_ASAP7_75t_L g746 ( .A(n_534), .B(n_575), .Y(n_746) );
NAND2xp5_ASAP7_75t_L g535 ( .A(n_536), .B(n_540), .Y(n_535) );
AOI222xp33_ASAP7_75t_L g734 ( .A1(n_542), .A2(n_606), .B1(n_649), .B2(n_709), .C1(n_735), .C2(n_737), .Y(n_734) );
INVx1_ASAP7_75t_L g542 ( .A(n_543), .Y(n_542) );
NAND2xp5_ASAP7_75t_L g543 ( .A(n_544), .B(n_554), .Y(n_543) );
AND2x2_ASAP7_75t_L g653 ( .A(n_544), .B(n_573), .Y(n_653) );
NAND2xp5_ASAP7_75t_L g703 ( .A(n_544), .B(n_704), .Y(n_703) );
AND2x2_ASAP7_75t_L g782 ( .A(n_544), .B(n_622), .Y(n_782) );
INVx2_ASAP7_75t_L g544 ( .A(n_545), .Y(n_544) );
AOI21xp5_ASAP7_75t_L g612 ( .A1(n_545), .A2(n_613), .B(n_617), .Y(n_612) );
AND2x2_ASAP7_75t_L g693 ( .A(n_545), .B(n_576), .Y(n_693) );
OR2x2_ASAP7_75t_L g718 ( .A(n_545), .B(n_577), .Y(n_718) );
INVx2_ASAP7_75t_L g545 ( .A(n_546), .Y(n_545) );
INVx5_ASAP7_75t_L g572 ( .A(n_546), .Y(n_572) );
AND2x2_ASAP7_75t_L g659 ( .A(n_546), .B(n_641), .Y(n_659) );
AND2x2_ASAP7_75t_L g685 ( .A(n_546), .B(n_561), .Y(n_685) );
OR2x2_ASAP7_75t_L g688 ( .A(n_546), .B(n_575), .Y(n_688) );
HB1xp67_ASAP7_75t_L g706 ( .A(n_546), .Y(n_706) );
AND2x4_ASAP7_75t_SL g763 ( .A(n_546), .B(n_640), .Y(n_763) );
OR2x2_ASAP7_75t_L g772 ( .A(n_546), .B(n_599), .Y(n_772) );
OR2x6_ASAP7_75t_L g546 ( .A(n_547), .B(n_548), .Y(n_546) );
INVx1_ASAP7_75t_L g605 ( .A(n_554), .Y(n_605) );
AOI221xp5_ASAP7_75t_SL g723 ( .A1(n_554), .A2(n_607), .B1(n_724), .B2(n_726), .C(n_727), .Y(n_723) );
AND2x2_ASAP7_75t_L g554 ( .A(n_555), .B(n_561), .Y(n_554) );
OR2x2_ASAP7_75t_L g662 ( .A(n_555), .B(n_632), .Y(n_662) );
OR2x2_ASAP7_75t_L g672 ( .A(n_555), .B(n_673), .Y(n_672) );
OR2x2_ASAP7_75t_L g698 ( .A(n_555), .B(n_699), .Y(n_698) );
AND2x4_ASAP7_75t_L g704 ( .A(n_555), .B(n_623), .Y(n_704) );
NOR2xp33_ASAP7_75t_L g716 ( .A(n_555), .B(n_687), .Y(n_716) );
INVx2_ASAP7_75t_L g729 ( .A(n_555), .Y(n_729) );
NAND2xp5_ASAP7_75t_SL g750 ( .A(n_555), .B(n_607), .Y(n_750) );
AND2x2_ASAP7_75t_L g754 ( .A(n_555), .B(n_576), .Y(n_754) );
AND2x2_ASAP7_75t_L g762 ( .A(n_555), .B(n_763), .Y(n_762) );
BUFx6f_ASAP7_75t_L g555 ( .A(n_556), .Y(n_555) );
INVx2_ASAP7_75t_L g575 ( .A(n_556), .Y(n_575) );
NAND2xp5_ASAP7_75t_L g557 ( .A(n_558), .B(n_559), .Y(n_557) );
NAND2xp5_ASAP7_75t_L g571 ( .A(n_561), .B(n_572), .Y(n_571) );
AND2x2_ASAP7_75t_L g606 ( .A(n_561), .B(n_575), .Y(n_606) );
INVx2_ASAP7_75t_L g623 ( .A(n_561), .Y(n_623) );
AND2x4_ASAP7_75t_L g640 ( .A(n_561), .B(n_641), .Y(n_640) );
HB1xp67_ASAP7_75t_L g745 ( .A(n_561), .Y(n_745) );
NAND2xp5_ASAP7_75t_L g562 ( .A(n_563), .B(n_567), .Y(n_562) );
NOR2xp33_ASAP7_75t_L g569 ( .A(n_570), .B(n_573), .Y(n_569) );
INVx1_ASAP7_75t_L g570 ( .A(n_571), .Y(n_570) );
OR2x2_ASAP7_75t_L g752 ( .A(n_571), .B(n_574), .Y(n_752) );
AND2x4_ASAP7_75t_L g598 ( .A(n_572), .B(n_599), .Y(n_598) );
AND2x2_ASAP7_75t_L g639 ( .A(n_572), .B(n_640), .Y(n_639) );
AND2x2_ASAP7_75t_L g666 ( .A(n_572), .B(n_606), .Y(n_666) );
AND2x2_ASAP7_75t_L g573 ( .A(n_574), .B(n_576), .Y(n_573) );
AND2x2_ASAP7_75t_L g770 ( .A(n_574), .B(n_771), .Y(n_770) );
BUFx2_ASAP7_75t_L g574 ( .A(n_575), .Y(n_574) );
AND2x2_ASAP7_75t_L g622 ( .A(n_575), .B(n_623), .Y(n_622) );
OAI21xp5_ASAP7_75t_SL g642 ( .A1(n_576), .A2(n_643), .B(n_649), .Y(n_642) );
INVx2_ASAP7_75t_L g576 ( .A(n_577), .Y(n_576) );
INVx1_ASAP7_75t_SL g578 ( .A(n_579), .Y(n_578) );
AND2x2_ASAP7_75t_L g579 ( .A(n_580), .B(n_589), .Y(n_579) );
INVx1_ASAP7_75t_SL g696 ( .A(n_580), .Y(n_696) );
AND2x2_ASAP7_75t_L g726 ( .A(n_580), .B(n_636), .Y(n_726) );
AND2x4_ASAP7_75t_L g737 ( .A(n_580), .B(n_738), .Y(n_737) );
OR2x2_ASAP7_75t_L g603 ( .A(n_581), .B(n_604), .Y(n_603) );
INVx2_ASAP7_75t_L g610 ( .A(n_581), .Y(n_610) );
AND2x4_ASAP7_75t_L g616 ( .A(n_581), .B(n_602), .Y(n_616) );
INVx2_ASAP7_75t_L g627 ( .A(n_581), .Y(n_627) );
INVx1_ASAP7_75t_L g676 ( .A(n_581), .Y(n_676) );
OR2x2_ASAP7_75t_L g697 ( .A(n_581), .B(n_681), .Y(n_697) );
OR2x2_ASAP7_75t_L g711 ( .A(n_581), .B(n_591), .Y(n_711) );
HB1xp67_ASAP7_75t_L g777 ( .A(n_581), .Y(n_777) );
NAND2xp5_ASAP7_75t_L g783 ( .A(n_581), .B(n_633), .Y(n_783) );
OR2x6_ASAP7_75t_L g581 ( .A(n_582), .B(n_588), .Y(n_581) );
INVx1_ASAP7_75t_L g628 ( .A(n_589), .Y(n_628) );
AND2x2_ASAP7_75t_L g761 ( .A(n_589), .B(n_627), .Y(n_761) );
AND2x2_ASAP7_75t_L g786 ( .A(n_589), .B(n_616), .Y(n_786) );
INVx2_ASAP7_75t_L g590 ( .A(n_591), .Y(n_590) );
INVx2_ASAP7_75t_L g604 ( .A(n_591), .Y(n_604) );
BUFx3_ASAP7_75t_L g646 ( .A(n_591), .Y(n_646) );
HB1xp67_ASAP7_75t_L g673 ( .A(n_591), .Y(n_673) );
INVx1_ASAP7_75t_L g682 ( .A(n_591), .Y(n_682) );
AOI33xp33_ASAP7_75t_L g597 ( .A1(n_598), .A2(n_600), .A3(n_605), .B1(n_606), .B2(n_607), .B3(n_608), .Y(n_597) );
AOI21x1_ASAP7_75t_SL g700 ( .A1(n_598), .A2(n_622), .B(n_684), .Y(n_700) );
INVx2_ASAP7_75t_L g730 ( .A(n_598), .Y(n_730) );
NAND2xp5_ASAP7_75t_L g736 ( .A(n_598), .B(n_729), .Y(n_736) );
AND2x2_ASAP7_75t_L g684 ( .A(n_599), .B(n_685), .Y(n_684) );
INVx1_ASAP7_75t_SL g600 ( .A(n_601), .Y(n_600) );
OR2x2_ASAP7_75t_L g601 ( .A(n_602), .B(n_603), .Y(n_601) );
AND2x2_ASAP7_75t_L g647 ( .A(n_602), .B(n_648), .Y(n_647) );
INVx2_ASAP7_75t_L g748 ( .A(n_603), .Y(n_748) );
HB1xp67_ASAP7_75t_L g738 ( .A(n_604), .Y(n_738) );
OAI32xp33_ASAP7_75t_L g787 ( .A1(n_605), .A2(n_607), .A3(n_783), .B1(n_788), .B2(n_790), .Y(n_787) );
AND2x2_ASAP7_75t_L g705 ( .A(n_606), .B(n_706), .Y(n_705) );
INVx2_ASAP7_75t_SL g695 ( .A(n_607), .Y(n_695) );
AND2x2_ASAP7_75t_L g760 ( .A(n_607), .B(n_704), .Y(n_760) );
INVx1_ASAP7_75t_L g608 ( .A(n_609), .Y(n_608) );
OAI221xp5_ASAP7_75t_L g611 ( .A1(n_612), .A2(n_621), .B1(n_624), .B2(n_638), .C(n_642), .Y(n_611) );
INVx1_ASAP7_75t_L g613 ( .A(n_614), .Y(n_613) );
NAND2xp5_ASAP7_75t_L g614 ( .A(n_615), .B(n_616), .Y(n_614) );
NAND2xp5_ASAP7_75t_L g681 ( .A(n_615), .B(n_682), .Y(n_681) );
NAND2xp5_ASAP7_75t_L g618 ( .A(n_616), .B(n_619), .Y(n_618) );
NAND2xp5_ASAP7_75t_L g731 ( .A(n_616), .B(n_732), .Y(n_731) );
NAND2xp5_ASAP7_75t_L g755 ( .A(n_616), .B(n_756), .Y(n_755) );
INVx1_ASAP7_75t_L g617 ( .A(n_618), .Y(n_617) );
INVx1_ASAP7_75t_L g619 ( .A(n_620), .Y(n_619) );
INVx1_ASAP7_75t_L g665 ( .A(n_620), .Y(n_665) );
INVx1_ASAP7_75t_L g621 ( .A(n_622), .Y(n_621) );
NOR3xp33_ASAP7_75t_L g624 ( .A(n_625), .B(n_629), .C(n_634), .Y(n_624) );
INVx1_ASAP7_75t_SL g625 ( .A(n_626), .Y(n_625) );
OAI22xp33_ASAP7_75t_L g727 ( .A1(n_626), .A2(n_688), .B1(n_728), .B2(n_731), .Y(n_727) );
OR2x2_ASAP7_75t_L g626 ( .A(n_627), .B(n_628), .Y(n_626) );
INVx1_ASAP7_75t_L g631 ( .A(n_627), .Y(n_631) );
NOR2x1p5_ASAP7_75t_L g645 ( .A(n_627), .B(n_646), .Y(n_645) );
HB1xp67_ASAP7_75t_L g667 ( .A(n_627), .Y(n_667) );
INVx1_ASAP7_75t_L g629 ( .A(n_630), .Y(n_629) );
OAI322xp33_ASAP7_75t_L g694 ( .A1(n_630), .A2(n_672), .A3(n_695), .B1(n_696), .B2(n_697), .C1(n_698), .C2(n_700), .Y(n_694) );
OR2x2_ASAP7_75t_L g630 ( .A(n_631), .B(n_632), .Y(n_630) );
A2O1A1Ixp33_ASAP7_75t_L g650 ( .A1(n_632), .A2(n_651), .B(n_652), .C(n_654), .Y(n_650) );
OR2x2_ASAP7_75t_L g742 ( .A(n_632), .B(n_696), .Y(n_742) );
INVx2_ASAP7_75t_L g632 ( .A(n_633), .Y(n_632) );
AND2x2_ASAP7_75t_L g649 ( .A(n_633), .B(n_637), .Y(n_649) );
INVx1_ASAP7_75t_L g634 ( .A(n_635), .Y(n_634) );
NAND2xp5_ASAP7_75t_L g635 ( .A(n_636), .B(n_637), .Y(n_635) );
INVx2_ASAP7_75t_L g638 ( .A(n_639), .Y(n_638) );
AND2x2_ASAP7_75t_L g655 ( .A(n_639), .B(n_656), .Y(n_655) );
INVx3_ASAP7_75t_SL g687 ( .A(n_640), .Y(n_687) );
INVx1_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
NAND2xp5_ASAP7_75t_L g707 ( .A(n_644), .B(n_708), .Y(n_707) );
NAND2xp5_ASAP7_75t_L g644 ( .A(n_645), .B(n_647), .Y(n_644) );
INVx1_ASAP7_75t_SL g691 ( .A(n_647), .Y(n_691) );
HB1xp67_ASAP7_75t_L g733 ( .A(n_648), .Y(n_733) );
OR2x6_ASAP7_75t_SL g788 ( .A(n_651), .B(n_789), .Y(n_788) );
INVx1_ASAP7_75t_L g652 ( .A(n_653), .Y(n_652) );
INVxp67_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
AOI211xp5_ASAP7_75t_L g778 ( .A1(n_656), .A2(n_779), .B(n_780), .C(n_787), .Y(n_778) );
O2A1O1Ixp33_ASAP7_75t_SL g657 ( .A1(n_658), .A2(n_660), .B(n_663), .C(n_667), .Y(n_657) );
OAI211xp5_ASAP7_75t_SL g669 ( .A1(n_658), .A2(n_670), .B(n_677), .C(n_701), .Y(n_669) );
INVx2_ASAP7_75t_L g658 ( .A(n_659), .Y(n_658) );
INVx1_ASAP7_75t_L g660 ( .A(n_661), .Y(n_660) );
INVx3_ASAP7_75t_L g661 ( .A(n_662), .Y(n_661) );
INVxp67_ASAP7_75t_L g663 ( .A(n_664), .Y(n_663) );
AND2x2_ASAP7_75t_L g664 ( .A(n_665), .B(n_666), .Y(n_664) );
NOR3xp33_ASAP7_75t_L g668 ( .A(n_669), .B(n_714), .C(n_758), .Y(n_668) );
NAND2xp5_ASAP7_75t_L g670 ( .A(n_671), .B(n_674), .Y(n_670) );
INVx1_ASAP7_75t_SL g671 ( .A(n_672), .Y(n_671) );
HB1xp67_ASAP7_75t_L g765 ( .A(n_673), .Y(n_765) );
INVx1_ASAP7_75t_SL g674 ( .A(n_675), .Y(n_674) );
INVx1_ASAP7_75t_L g720 ( .A(n_676), .Y(n_720) );
NOR3xp33_ASAP7_75t_SL g677 ( .A(n_678), .B(n_690), .C(n_694), .Y(n_677) );
OAI22xp5_ASAP7_75t_L g678 ( .A1(n_679), .A2(n_683), .B1(n_686), .B2(n_689), .Y(n_678) );
INVx1_ASAP7_75t_L g679 ( .A(n_680), .Y(n_679) );
INVx1_ASAP7_75t_L g680 ( .A(n_681), .Y(n_680) );
INVx1_ASAP7_75t_L g722 ( .A(n_682), .Y(n_722) );
INVxp67_ASAP7_75t_SL g789 ( .A(n_682), .Y(n_789) );
INVx1_ASAP7_75t_L g683 ( .A(n_684), .Y(n_683) );
OR2x2_ASAP7_75t_L g686 ( .A(n_687), .B(n_688), .Y(n_686) );
INVx1_ASAP7_75t_SL g775 ( .A(n_688), .Y(n_775) );
NOR2xp33_ASAP7_75t_L g690 ( .A(n_691), .B(n_692), .Y(n_690) );
OR2x2_ASAP7_75t_L g725 ( .A(n_691), .B(n_711), .Y(n_725) );
OR2x2_ASAP7_75t_L g776 ( .A(n_691), .B(n_777), .Y(n_776) );
INVx2_ASAP7_75t_L g692 ( .A(n_693), .Y(n_692) );
INVx1_ASAP7_75t_L g774 ( .A(n_699), .Y(n_774) );
OR2x2_ASAP7_75t_L g790 ( .A(n_699), .B(n_729), .Y(n_790) );
OAI21xp33_ASAP7_75t_L g701 ( .A1(n_702), .A2(n_705), .B(n_707), .Y(n_701) );
OAI31xp33_ASAP7_75t_L g715 ( .A1(n_702), .A2(n_716), .A3(n_717), .B(n_719), .Y(n_715) );
INVx1_ASAP7_75t_L g702 ( .A(n_703), .Y(n_702) );
INVx1_ASAP7_75t_L g708 ( .A(n_709), .Y(n_708) );
AND2x2_ASAP7_75t_L g709 ( .A(n_710), .B(n_712), .Y(n_709) );
INVx1_ASAP7_75t_SL g710 ( .A(n_711), .Y(n_710) );
AND2x4_ASAP7_75t_L g747 ( .A(n_712), .B(n_748), .Y(n_747) );
INVx1_ASAP7_75t_L g712 ( .A(n_713), .Y(n_712) );
NAND4xp25_ASAP7_75t_SL g714 ( .A(n_715), .B(n_723), .C(n_734), .D(n_739), .Y(n_714) );
INVx1_ASAP7_75t_L g717 ( .A(n_718), .Y(n_717) );
AND2x2_ASAP7_75t_L g719 ( .A(n_720), .B(n_721), .Y(n_719) );
HB1xp67_ASAP7_75t_L g757 ( .A(n_722), .Y(n_757) );
INVx1_ASAP7_75t_SL g724 ( .A(n_725), .Y(n_724) );
OR2x2_ASAP7_75t_L g728 ( .A(n_729), .B(n_730), .Y(n_728) );
INVxp67_ASAP7_75t_L g732 ( .A(n_733), .Y(n_732) );
INVx1_ASAP7_75t_L g735 ( .A(n_736), .Y(n_735) );
AOI221xp5_ASAP7_75t_L g739 ( .A1(n_740), .A2(n_743), .B1(n_747), .B2(n_749), .C(n_751), .Y(n_739) );
NAND2xp33_ASAP7_75t_SL g740 ( .A(n_741), .B(n_742), .Y(n_740) );
INVx1_ASAP7_75t_L g784 ( .A(n_743), .Y(n_784) );
AND2x2_ASAP7_75t_SL g743 ( .A(n_744), .B(n_746), .Y(n_743) );
INVx1_ASAP7_75t_L g744 ( .A(n_745), .Y(n_744) );
INVx1_ASAP7_75t_L g749 ( .A(n_750), .Y(n_749) );
AOI21xp33_ASAP7_75t_L g751 ( .A1(n_752), .A2(n_753), .B(n_755), .Y(n_751) );
INVx1_ASAP7_75t_L g779 ( .A(n_753), .Y(n_779) );
INVx2_ASAP7_75t_L g753 ( .A(n_754), .Y(n_753) );
INVx1_ASAP7_75t_L g756 ( .A(n_757), .Y(n_756) );
NAND2xp5_ASAP7_75t_SL g758 ( .A(n_759), .B(n_778), .Y(n_758) );
AOI221xp5_ASAP7_75t_L g759 ( .A1(n_760), .A2(n_761), .B1(n_762), .B2(n_764), .C(n_768), .Y(n_759) );
AND2x2_ASAP7_75t_L g764 ( .A(n_765), .B(n_766), .Y(n_764) );
INVx1_ASAP7_75t_SL g766 ( .A(n_767), .Y(n_766) );
AOI21xp33_ASAP7_75t_L g768 ( .A1(n_769), .A2(n_773), .B(n_776), .Y(n_768) );
INVxp33_ASAP7_75t_L g769 ( .A(n_770), .Y(n_769) );
INVx1_ASAP7_75t_SL g771 ( .A(n_772), .Y(n_771) );
NAND2xp5_ASAP7_75t_L g773 ( .A(n_774), .B(n_775), .Y(n_773) );
OAI22xp5_ASAP7_75t_L g780 ( .A1(n_781), .A2(n_783), .B1(n_784), .B2(n_785), .Y(n_780) );
INVx1_ASAP7_75t_L g781 ( .A(n_782), .Y(n_781) );
INVx1_ASAP7_75t_L g785 ( .A(n_786), .Y(n_785) );
CKINVDCx5p33_ASAP7_75t_R g791 ( .A(n_792), .Y(n_791) );
CKINVDCx20_ASAP7_75t_R g802 ( .A(n_792), .Y(n_802) );
CKINVDCx11_ASAP7_75t_R g792 ( .A(n_793), .Y(n_792) );
INVx1_ASAP7_75t_L g796 ( .A(n_797), .Y(n_796) );
INVx2_ASAP7_75t_L g803 ( .A(n_804), .Y(n_803) );
NAND2xp5_ASAP7_75t_L g806 ( .A(n_807), .B(n_810), .Y(n_806) );
CKINVDCx11_ASAP7_75t_R g807 ( .A(n_808), .Y(n_807) );
CKINVDCx20_ASAP7_75t_R g808 ( .A(n_809), .Y(n_808) );
INVxp67_ASAP7_75t_SL g822 ( .A(n_810), .Y(n_822) );
XNOR2xp5_ASAP7_75t_L g810 ( .A(n_811), .B(n_815), .Y(n_810) );
NAND3x1_ASAP7_75t_L g811 ( .A(n_812), .B(n_813), .C(n_814), .Y(n_811) );
CKINVDCx5p33_ASAP7_75t_R g815 ( .A(n_816), .Y(n_815) );
INVx1_ASAP7_75t_L g820 ( .A(n_818), .Y(n_820) );
NOR2xp33_ASAP7_75t_L g823 ( .A(n_824), .B(n_825), .Y(n_823) );
CKINVDCx5p33_ASAP7_75t_R g826 ( .A(n_827), .Y(n_826) );
endmodule