module real_aes_8363_n_101 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_101);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_101;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_357;
wire n_287;
wire n_635;
wire n_503;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_744;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_178;
wire n_409;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_725;
wire n_455;
wire n_310;
wire n_504;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_527;
wire n_434;
wire n_502;
wire n_505;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_733;
wire n_402;
wire n_552;
wire n_602;
wire n_617;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_713;
wire n_288;
wire n_404;
wire n_598;
wire n_728;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_720;
wire n_354;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_233;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_679;
wire n_633;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_456;
wire n_359;
wire n_717;
wire n_712;
wire n_266;
wire n_183;
wire n_312;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_479;
wire n_338;
wire n_442;
wire n_740;
wire n_371;
wire n_698;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_639;
wire n_546;
wire n_587;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_719;
wire n_473;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_424;
wire n_225;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
A2O1A1Ixp33_ASAP7_75t_SL g261 ( .A1(n_0), .A2(n_262), .B(n_263), .C(n_266), .Y(n_261) );
NAND2xp5_ASAP7_75t_L g267 ( .A(n_1), .B(n_203), .Y(n_267) );
NAND3xp33_ASAP7_75t_SL g109 ( .A(n_2), .B(n_110), .C(n_111), .Y(n_109) );
INVx1_ASAP7_75t_L g441 ( .A(n_2), .Y(n_441) );
NAND2xp5_ASAP7_75t_SL g239 ( .A(n_3), .B(n_173), .Y(n_239) );
A2O1A1Ixp33_ASAP7_75t_L g453 ( .A1(n_4), .A2(n_143), .B(n_146), .C(n_454), .Y(n_453) );
AOI21xp5_ASAP7_75t_L g493 ( .A1(n_5), .A2(n_163), .B(n_494), .Y(n_493) );
AOI21xp5_ASAP7_75t_L g193 ( .A1(n_6), .A2(n_163), .B(n_194), .Y(n_193) );
NAND2xp5_ASAP7_75t_L g500 ( .A(n_7), .B(n_203), .Y(n_500) );
AO21x2_ASAP7_75t_L g182 ( .A1(n_8), .A2(n_130), .B(n_183), .Y(n_182) );
AND2x6_ASAP7_75t_L g143 ( .A(n_9), .B(n_144), .Y(n_143) );
A2O1A1Ixp33_ASAP7_75t_L g145 ( .A1(n_10), .A2(n_143), .B(n_146), .C(n_149), .Y(n_145) );
OAI22xp5_ASAP7_75t_L g116 ( .A1(n_11), .A2(n_45), .B1(n_117), .B2(n_118), .Y(n_116) );
CKINVDCx20_ASAP7_75t_R g117 ( .A(n_11), .Y(n_117) );
INVx1_ASAP7_75t_L g107 ( .A(n_12), .Y(n_107) );
NOR2xp33_ASAP7_75t_L g442 ( .A(n_12), .B(n_41), .Y(n_442) );
INVx1_ASAP7_75t_L g470 ( .A(n_13), .Y(n_470) );
NAND2xp5_ASAP7_75t_SL g456 ( .A(n_14), .B(n_153), .Y(n_456) );
INVx1_ASAP7_75t_L g135 ( .A(n_15), .Y(n_135) );
NAND2xp5_ASAP7_75t_SL g189 ( .A(n_16), .B(n_173), .Y(n_189) );
AOI22xp33_ASAP7_75t_L g101 ( .A1(n_17), .A2(n_102), .B1(n_114), .B2(n_744), .Y(n_101) );
A2O1A1Ixp33_ASAP7_75t_L g477 ( .A1(n_18), .A2(n_151), .B(n_478), .C(n_480), .Y(n_477) );
NAND2xp5_ASAP7_75t_L g481 ( .A(n_19), .B(n_203), .Y(n_481) );
NAND2xp5_ASAP7_75t_L g513 ( .A(n_20), .B(n_227), .Y(n_513) );
A2O1A1Ixp33_ASAP7_75t_L g222 ( .A1(n_21), .A2(n_146), .B(n_190), .C(n_223), .Y(n_222) );
A2O1A1Ixp33_ASAP7_75t_L g486 ( .A1(n_22), .A2(n_155), .B(n_265), .C(n_487), .Y(n_486) );
NAND2xp5_ASAP7_75t_SL g532 ( .A(n_23), .B(n_153), .Y(n_532) );
CKINVDCx20_ASAP7_75t_R g741 ( .A(n_24), .Y(n_741) );
NAND2xp5_ASAP7_75t_SL g521 ( .A(n_25), .B(n_153), .Y(n_521) );
CKINVDCx16_ASAP7_75t_R g528 ( .A(n_26), .Y(n_528) );
INVx1_ASAP7_75t_L g520 ( .A(n_27), .Y(n_520) );
A2O1A1Ixp33_ASAP7_75t_L g185 ( .A1(n_28), .A2(n_146), .B(n_186), .C(n_190), .Y(n_185) );
BUFx6f_ASAP7_75t_L g142 ( .A(n_29), .Y(n_142) );
CKINVDCx20_ASAP7_75t_R g452 ( .A(n_30), .Y(n_452) );
INVx1_ASAP7_75t_L g511 ( .A(n_31), .Y(n_511) );
AOI21xp5_ASAP7_75t_L g258 ( .A1(n_32), .A2(n_163), .B(n_259), .Y(n_258) );
INVx2_ASAP7_75t_L g141 ( .A(n_33), .Y(n_141) );
A2O1A1Ixp33_ASAP7_75t_L g210 ( .A1(n_34), .A2(n_165), .B(n_176), .C(n_211), .Y(n_210) );
CKINVDCx20_ASAP7_75t_R g459 ( .A(n_35), .Y(n_459) );
A2O1A1Ixp33_ASAP7_75t_L g496 ( .A1(n_36), .A2(n_265), .B(n_497), .C(n_499), .Y(n_496) );
INVxp67_ASAP7_75t_L g512 ( .A(n_37), .Y(n_512) );
NAND2xp5_ASAP7_75t_L g187 ( .A(n_38), .B(n_188), .Y(n_187) );
CKINVDCx14_ASAP7_75t_R g495 ( .A(n_39), .Y(n_495) );
A2O1A1Ixp33_ASAP7_75t_L g518 ( .A1(n_40), .A2(n_146), .B(n_190), .C(n_519), .Y(n_518) );
NAND2xp5_ASAP7_75t_L g106 ( .A(n_41), .B(n_107), .Y(n_106) );
A2O1A1Ixp33_ASAP7_75t_L g467 ( .A1(n_42), .A2(n_266), .B(n_468), .C(n_469), .Y(n_467) );
NAND2xp5_ASAP7_75t_L g220 ( .A(n_43), .B(n_221), .Y(n_220) );
CKINVDCx20_ASAP7_75t_R g158 ( .A(n_44), .Y(n_158) );
INVx1_ASAP7_75t_L g118 ( .A(n_45), .Y(n_118) );
NAND2xp5_ASAP7_75t_L g172 ( .A(n_46), .B(n_173), .Y(n_172) );
NAND2xp5_ASAP7_75t_L g184 ( .A(n_47), .B(n_163), .Y(n_184) );
CKINVDCx20_ASAP7_75t_R g523 ( .A(n_48), .Y(n_523) );
CKINVDCx20_ASAP7_75t_R g508 ( .A(n_49), .Y(n_508) );
A2O1A1Ixp33_ASAP7_75t_L g164 ( .A1(n_50), .A2(n_165), .B(n_167), .C(n_176), .Y(n_164) );
INVx1_ASAP7_75t_L g264 ( .A(n_51), .Y(n_264) );
INVx1_ASAP7_75t_L g168 ( .A(n_52), .Y(n_168) );
INVx1_ASAP7_75t_L g485 ( .A(n_53), .Y(n_485) );
NAND2xp5_ASAP7_75t_L g162 ( .A(n_54), .B(n_163), .Y(n_162) );
OAI22xp5_ASAP7_75t_SL g732 ( .A1(n_55), .A2(n_59), .B1(n_733), .B2(n_734), .Y(n_732) );
CKINVDCx20_ASAP7_75t_R g734 ( .A(n_55), .Y(n_734) );
CKINVDCx20_ASAP7_75t_R g719 ( .A(n_56), .Y(n_719) );
CKINVDCx20_ASAP7_75t_R g230 ( .A(n_57), .Y(n_230) );
CKINVDCx14_ASAP7_75t_R g466 ( .A(n_58), .Y(n_466) );
CKINVDCx20_ASAP7_75t_R g733 ( .A(n_59), .Y(n_733) );
INVx1_ASAP7_75t_L g144 ( .A(n_60), .Y(n_144) );
NAND2xp5_ASAP7_75t_L g242 ( .A(n_61), .B(n_163), .Y(n_242) );
NAND2xp5_ASAP7_75t_L g202 ( .A(n_62), .B(n_203), .Y(n_202) );
A2O1A1Ixp33_ASAP7_75t_L g196 ( .A1(n_63), .A2(n_197), .B(n_199), .C(n_201), .Y(n_196) );
INVx1_ASAP7_75t_L g134 ( .A(n_64), .Y(n_134) );
INVx1_ASAP7_75t_SL g498 ( .A(n_65), .Y(n_498) );
CKINVDCx20_ASAP7_75t_R g727 ( .A(n_66), .Y(n_727) );
NAND2xp5_ASAP7_75t_SL g213 ( .A(n_67), .B(n_173), .Y(n_213) );
NAND2xp5_ASAP7_75t_L g489 ( .A(n_68), .B(n_203), .Y(n_489) );
NAND2xp5_ASAP7_75t_L g150 ( .A(n_69), .B(n_151), .Y(n_150) );
INVx1_ASAP7_75t_L g531 ( .A(n_70), .Y(n_531) );
CKINVDCx16_ASAP7_75t_R g260 ( .A(n_71), .Y(n_260) );
NAND2xp5_ASAP7_75t_L g224 ( .A(n_72), .B(n_170), .Y(n_224) );
A2O1A1Ixp33_ASAP7_75t_L g236 ( .A1(n_73), .A2(n_146), .B(n_176), .C(n_237), .Y(n_236) );
CKINVDCx16_ASAP7_75t_R g195 ( .A(n_74), .Y(n_195) );
INVx1_ASAP7_75t_L g113 ( .A(n_75), .Y(n_113) );
AOI21xp5_ASAP7_75t_L g464 ( .A1(n_76), .A2(n_163), .B(n_465), .Y(n_464) );
CKINVDCx20_ASAP7_75t_R g534 ( .A(n_77), .Y(n_534) );
AOI21xp5_ASAP7_75t_L g474 ( .A1(n_78), .A2(n_163), .B(n_475), .Y(n_474) );
AOI21xp5_ASAP7_75t_L g506 ( .A1(n_79), .A2(n_221), .B(n_507), .Y(n_506) );
INVx1_ASAP7_75t_L g476 ( .A(n_80), .Y(n_476) );
CKINVDCx16_ASAP7_75t_R g517 ( .A(n_81), .Y(n_517) );
NAND2xp5_ASAP7_75t_SL g225 ( .A(n_82), .B(n_169), .Y(n_225) );
CKINVDCx20_ASAP7_75t_R g215 ( .A(n_83), .Y(n_215) );
AOI21xp5_ASAP7_75t_L g483 ( .A1(n_84), .A2(n_163), .B(n_484), .Y(n_483) );
INVx1_ASAP7_75t_L g479 ( .A(n_85), .Y(n_479) );
INVx2_ASAP7_75t_L g132 ( .A(n_86), .Y(n_132) );
INVx1_ASAP7_75t_L g455 ( .A(n_87), .Y(n_455) );
CKINVDCx20_ASAP7_75t_R g244 ( .A(n_88), .Y(n_244) );
NAND2xp5_ASAP7_75t_SL g152 ( .A(n_89), .B(n_153), .Y(n_152) );
INVx2_ASAP7_75t_L g110 ( .A(n_90), .Y(n_110) );
OR2x2_ASAP7_75t_L g439 ( .A(n_90), .B(n_440), .Y(n_439) );
OR2x2_ASAP7_75t_L g737 ( .A(n_90), .B(n_724), .Y(n_737) );
A2O1A1Ixp33_ASAP7_75t_L g529 ( .A1(n_91), .A2(n_146), .B(n_176), .C(n_530), .Y(n_529) );
NAND2xp5_ASAP7_75t_L g209 ( .A(n_92), .B(n_163), .Y(n_209) );
INVx1_ASAP7_75t_L g212 ( .A(n_93), .Y(n_212) );
INVxp67_ASAP7_75t_L g200 ( .A(n_94), .Y(n_200) );
NAND2xp5_ASAP7_75t_L g471 ( .A(n_95), .B(n_130), .Y(n_471) );
INVx2_ASAP7_75t_L g488 ( .A(n_96), .Y(n_488) );
NAND2xp5_ASAP7_75t_L g112 ( .A(n_97), .B(n_113), .Y(n_112) );
INVx1_ASAP7_75t_L g137 ( .A(n_98), .Y(n_137) );
INVx1_ASAP7_75t_L g238 ( .A(n_99), .Y(n_238) );
AND2x2_ASAP7_75t_L g179 ( .A(n_100), .B(n_178), .Y(n_179) );
INVx1_ASAP7_75t_SL g102 ( .A(n_103), .Y(n_102) );
INVx2_ASAP7_75t_SL g103 ( .A(n_104), .Y(n_103) );
INVx2_ASAP7_75t_SL g744 ( .A(n_104), .Y(n_744) );
AND2x2_ASAP7_75t_L g104 ( .A(n_105), .B(n_108), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_106), .Y(n_105) );
INVx1_ASAP7_75t_L g108 ( .A(n_109), .Y(n_108) );
OR2x2_ASAP7_75t_L g711 ( .A(n_110), .B(n_440), .Y(n_711) );
NOR2x2_ASAP7_75t_L g723 ( .A(n_110), .B(n_724), .Y(n_723) );
INVx1_ASAP7_75t_SL g111 ( .A(n_112), .Y(n_111) );
AO221x1_ASAP7_75t_L g114 ( .A1(n_115), .A2(n_725), .B1(n_728), .B2(n_738), .C(n_740), .Y(n_114) );
OAI222xp33_ASAP7_75t_SL g115 ( .A1(n_116), .A2(n_119), .B1(n_712), .B2(n_713), .C1(n_719), .C2(n_720), .Y(n_115) );
INVx1_ASAP7_75t_L g712 ( .A(n_116), .Y(n_712) );
INVxp67_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
OAI22xp5_ASAP7_75t_SL g120 ( .A1(n_121), .A2(n_437), .B1(n_443), .B2(n_709), .Y(n_120) );
INVx2_ASAP7_75t_L g716 ( .A(n_121), .Y(n_716) );
AOI22xp5_ASAP7_75t_L g730 ( .A1(n_121), .A2(n_716), .B1(n_731), .B2(n_732), .Y(n_730) );
OR3x1_ASAP7_75t_L g121 ( .A(n_122), .B(n_335), .C(n_400), .Y(n_121) );
NAND4xp25_ASAP7_75t_SL g122 ( .A(n_123), .B(n_276), .C(n_302), .D(n_325), .Y(n_122) );
AOI221xp5_ASAP7_75t_L g123 ( .A1(n_124), .A2(n_204), .B1(n_245), .B2(n_252), .C(n_268), .Y(n_123) );
CKINVDCx14_ASAP7_75t_R g124 ( .A(n_125), .Y(n_124) );
OAI22xp5_ASAP7_75t_L g423 ( .A1(n_125), .A2(n_269), .B1(n_293), .B2(n_424), .Y(n_423) );
OR2x2_ASAP7_75t_L g125 ( .A(n_126), .B(n_180), .Y(n_125) );
INVx1_ASAP7_75t_SL g329 ( .A(n_126), .Y(n_329) );
OR2x2_ASAP7_75t_L g126 ( .A(n_127), .B(n_160), .Y(n_126) );
OR2x2_ASAP7_75t_L g250 ( .A(n_127), .B(n_251), .Y(n_250) );
AND2x2_ASAP7_75t_L g271 ( .A(n_127), .B(n_181), .Y(n_271) );
NAND2xp5_ASAP7_75t_L g284 ( .A(n_127), .B(n_191), .Y(n_284) );
AND2x2_ASAP7_75t_L g301 ( .A(n_127), .B(n_160), .Y(n_301) );
NAND2xp5_ASAP7_75t_L g323 ( .A(n_127), .B(n_248), .Y(n_323) );
NAND2xp5_ASAP7_75t_L g412 ( .A(n_127), .B(n_300), .Y(n_412) );
NOR2xp33_ASAP7_75t_L g422 ( .A(n_127), .B(n_180), .Y(n_422) );
AOI211xp5_ASAP7_75t_SL g433 ( .A1(n_127), .A2(n_339), .B(n_434), .C(n_435), .Y(n_433) );
INVx5_ASAP7_75t_SL g127 ( .A(n_128), .Y(n_127) );
NAND2xp5_ASAP7_75t_SL g305 ( .A(n_128), .B(n_181), .Y(n_305) );
AND2x2_ASAP7_75t_L g308 ( .A(n_128), .B(n_182), .Y(n_308) );
OR2x2_ASAP7_75t_L g353 ( .A(n_128), .B(n_181), .Y(n_353) );
NAND2xp5_ASAP7_75t_L g362 ( .A(n_128), .B(n_191), .Y(n_362) );
AO21x2_ASAP7_75t_L g128 ( .A1(n_129), .A2(n_136), .B(n_157), .Y(n_128) );
INVx3_ASAP7_75t_L g203 ( .A(n_129), .Y(n_203) );
NOR2xp33_ASAP7_75t_L g214 ( .A(n_129), .B(n_215), .Y(n_214) );
AO21x2_ASAP7_75t_L g234 ( .A1(n_129), .A2(n_235), .B(n_243), .Y(n_234) );
NOR2xp33_ASAP7_75t_L g243 ( .A(n_129), .B(n_244), .Y(n_243) );
NOR2xp33_ASAP7_75t_L g458 ( .A(n_129), .B(n_459), .Y(n_458) );
NOR2xp33_ASAP7_75t_L g522 ( .A(n_129), .B(n_523), .Y(n_522) );
AO21x2_ASAP7_75t_L g526 ( .A1(n_129), .A2(n_527), .B(n_533), .Y(n_526) );
INVx4_ASAP7_75t_L g129 ( .A(n_130), .Y(n_129) );
AOI21xp5_ASAP7_75t_L g183 ( .A1(n_130), .A2(n_184), .B(n_185), .Y(n_183) );
HB1xp67_ASAP7_75t_L g192 ( .A(n_130), .Y(n_192) );
BUFx6f_ASAP7_75t_L g130 ( .A(n_131), .Y(n_130) );
INVx1_ASAP7_75t_L g159 ( .A(n_131), .Y(n_159) );
AND2x2_ASAP7_75t_L g131 ( .A(n_132), .B(n_133), .Y(n_131) );
AND2x2_ASAP7_75t_SL g178 ( .A(n_132), .B(n_133), .Y(n_178) );
NAND2xp5_ASAP7_75t_L g133 ( .A(n_134), .B(n_135), .Y(n_133) );
OAI21xp5_ASAP7_75t_L g136 ( .A1(n_137), .A2(n_138), .B(n_145), .Y(n_136) );
OAI21xp5_ASAP7_75t_L g451 ( .A1(n_138), .A2(n_452), .B(n_453), .Y(n_451) );
O2A1O1Ixp33_ASAP7_75t_L g516 ( .A1(n_138), .A2(n_178), .B(n_517), .C(n_518), .Y(n_516) );
OAI21xp5_ASAP7_75t_L g527 ( .A1(n_138), .A2(n_528), .B(n_529), .Y(n_527) );
NAND2x1p5_ASAP7_75t_L g138 ( .A(n_139), .B(n_143), .Y(n_138) );
AND2x4_ASAP7_75t_L g163 ( .A(n_139), .B(n_143), .Y(n_163) );
AND2x2_ASAP7_75t_L g139 ( .A(n_140), .B(n_142), .Y(n_139) );
INVx1_ASAP7_75t_L g201 ( .A(n_140), .Y(n_201) );
INVx1_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
INVx2_ASAP7_75t_L g147 ( .A(n_141), .Y(n_147) );
INVx1_ASAP7_75t_L g156 ( .A(n_141), .Y(n_156) );
INVx1_ASAP7_75t_L g148 ( .A(n_142), .Y(n_148) );
INVx3_ASAP7_75t_L g151 ( .A(n_142), .Y(n_151) );
BUFx6f_ASAP7_75t_L g153 ( .A(n_142), .Y(n_153) );
BUFx6f_ASAP7_75t_L g171 ( .A(n_142), .Y(n_171) );
INVx1_ASAP7_75t_L g188 ( .A(n_142), .Y(n_188) );
INVx4_ASAP7_75t_SL g177 ( .A(n_143), .Y(n_177) );
BUFx3_ASAP7_75t_L g190 ( .A(n_143), .Y(n_190) );
INVx5_ASAP7_75t_L g166 ( .A(n_146), .Y(n_166) );
AND2x6_ASAP7_75t_L g146 ( .A(n_147), .B(n_148), .Y(n_146) );
BUFx3_ASAP7_75t_L g175 ( .A(n_147), .Y(n_175) );
BUFx6f_ASAP7_75t_L g241 ( .A(n_147), .Y(n_241) );
AOI21xp5_ASAP7_75t_L g149 ( .A1(n_150), .A2(n_152), .B(n_154), .Y(n_149) );
INVx5_ASAP7_75t_L g173 ( .A(n_151), .Y(n_173) );
NOR2xp33_ASAP7_75t_L g469 ( .A(n_151), .B(n_470), .Y(n_469) );
INVx4_ASAP7_75t_L g265 ( .A(n_153), .Y(n_265) );
INVx2_ASAP7_75t_L g468 ( .A(n_153), .Y(n_468) );
AOI21xp5_ASAP7_75t_L g186 ( .A1(n_154), .A2(n_187), .B(n_189), .Y(n_186) );
INVx2_ASAP7_75t_L g154 ( .A(n_155), .Y(n_154) );
INVx3_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
NOR2xp33_ASAP7_75t_L g157 ( .A(n_158), .B(n_159), .Y(n_157) );
INVx2_ASAP7_75t_L g505 ( .A(n_159), .Y(n_505) );
INVx5_ASAP7_75t_SL g251 ( .A(n_160), .Y(n_251) );
AND2x2_ASAP7_75t_L g270 ( .A(n_160), .B(n_271), .Y(n_270) );
NOR2xp33_ASAP7_75t_L g352 ( .A(n_160), .B(n_353), .Y(n_352) );
AND2x2_ASAP7_75t_L g356 ( .A(n_160), .B(n_357), .Y(n_356) );
AND2x2_ASAP7_75t_L g388 ( .A(n_160), .B(n_191), .Y(n_388) );
OR2x2_ASAP7_75t_L g394 ( .A(n_160), .B(n_284), .Y(n_394) );
NAND2xp5_ASAP7_75t_L g403 ( .A(n_160), .B(n_344), .Y(n_403) );
OR2x6_ASAP7_75t_L g160 ( .A(n_161), .B(n_179), .Y(n_160) );
AOI21xp5_ASAP7_75t_L g161 ( .A1(n_162), .A2(n_164), .B(n_178), .Y(n_161) );
BUFx2_ASAP7_75t_L g221 ( .A(n_163), .Y(n_221) );
INVx2_ASAP7_75t_L g165 ( .A(n_166), .Y(n_165) );
O2A1O1Ixp33_ASAP7_75t_L g194 ( .A1(n_166), .A2(n_177), .B(n_195), .C(n_196), .Y(n_194) );
O2A1O1Ixp33_ASAP7_75t_SL g259 ( .A1(n_166), .A2(n_177), .B(n_260), .C(n_261), .Y(n_259) );
O2A1O1Ixp33_ASAP7_75t_SL g465 ( .A1(n_166), .A2(n_177), .B(n_466), .C(n_467), .Y(n_465) );
O2A1O1Ixp33_ASAP7_75t_SL g475 ( .A1(n_166), .A2(n_177), .B(n_476), .C(n_477), .Y(n_475) );
O2A1O1Ixp33_ASAP7_75t_SL g484 ( .A1(n_166), .A2(n_177), .B(n_485), .C(n_486), .Y(n_484) );
O2A1O1Ixp33_ASAP7_75t_L g494 ( .A1(n_166), .A2(n_177), .B(n_495), .C(n_496), .Y(n_494) );
O2A1O1Ixp33_ASAP7_75t_SL g507 ( .A1(n_166), .A2(n_177), .B(n_508), .C(n_509), .Y(n_507) );
O2A1O1Ixp33_ASAP7_75t_L g167 ( .A1(n_168), .A2(n_169), .B(n_172), .C(n_174), .Y(n_167) );
O2A1O1Ixp33_ASAP7_75t_L g211 ( .A1(n_169), .A2(n_174), .B(n_212), .C(n_213), .Y(n_211) );
O2A1O1Ixp5_ASAP7_75t_L g454 ( .A1(n_169), .A2(n_455), .B(n_456), .C(n_457), .Y(n_454) );
O2A1O1Ixp33_ASAP7_75t_L g530 ( .A1(n_169), .A2(n_457), .B(n_531), .C(n_532), .Y(n_530) );
INVx2_ASAP7_75t_L g169 ( .A(n_170), .Y(n_169) );
INVx2_ASAP7_75t_L g170 ( .A(n_171), .Y(n_170) );
INVx4_ASAP7_75t_L g198 ( .A(n_171), .Y(n_198) );
NOR2xp33_ASAP7_75t_L g199 ( .A(n_173), .B(n_200), .Y(n_199) );
INVx2_ASAP7_75t_L g262 ( .A(n_173), .Y(n_262) );
OAI22xp33_ASAP7_75t_L g510 ( .A1(n_173), .A2(n_198), .B1(n_511), .B2(n_512), .Y(n_510) );
O2A1O1Ixp33_ASAP7_75t_L g519 ( .A1(n_173), .A2(n_226), .B(n_520), .C(n_521), .Y(n_519) );
HB1xp67_ASAP7_75t_L g174 ( .A(n_175), .Y(n_174) );
INVx2_ASAP7_75t_L g266 ( .A(n_175), .Y(n_266) );
INVx1_ASAP7_75t_L g480 ( .A(n_175), .Y(n_480) );
INVx1_ASAP7_75t_L g176 ( .A(n_177), .Y(n_176) );
AOI21xp5_ASAP7_75t_L g208 ( .A1(n_178), .A2(n_209), .B(n_210), .Y(n_208) );
INVx2_ASAP7_75t_L g228 ( .A(n_178), .Y(n_228) );
INVx1_ASAP7_75t_L g231 ( .A(n_178), .Y(n_231) );
OA21x2_ASAP7_75t_L g463 ( .A1(n_178), .A2(n_464), .B(n_471), .Y(n_463) );
NAND2xp5_ASAP7_75t_L g180 ( .A(n_181), .B(n_191), .Y(n_180) );
AND2x2_ASAP7_75t_L g285 ( .A(n_181), .B(n_251), .Y(n_285) );
INVx1_ASAP7_75t_SL g298 ( .A(n_181), .Y(n_298) );
OR2x2_ASAP7_75t_L g333 ( .A(n_181), .B(n_334), .Y(n_333) );
OR2x2_ASAP7_75t_L g339 ( .A(n_181), .B(n_191), .Y(n_339) );
AND2x2_ASAP7_75t_L g397 ( .A(n_181), .B(n_248), .Y(n_397) );
INVx2_ASAP7_75t_L g181 ( .A(n_182), .Y(n_181) );
NAND2xp5_ASAP7_75t_L g324 ( .A(n_182), .B(n_251), .Y(n_324) );
INVx3_ASAP7_75t_L g248 ( .A(n_191), .Y(n_248) );
OR2x2_ASAP7_75t_L g290 ( .A(n_191), .B(n_251), .Y(n_290) );
AND2x2_ASAP7_75t_L g300 ( .A(n_191), .B(n_298), .Y(n_300) );
HB1xp67_ASAP7_75t_L g348 ( .A(n_191), .Y(n_348) );
AND2x2_ASAP7_75t_L g357 ( .A(n_191), .B(n_271), .Y(n_357) );
OA21x2_ASAP7_75t_L g191 ( .A1(n_192), .A2(n_193), .B(n_202), .Y(n_191) );
OA21x2_ASAP7_75t_L g473 ( .A1(n_192), .A2(n_474), .B(n_481), .Y(n_473) );
OA21x2_ASAP7_75t_L g482 ( .A1(n_192), .A2(n_483), .B(n_489), .Y(n_482) );
OA21x2_ASAP7_75t_L g492 ( .A1(n_192), .A2(n_493), .B(n_500), .Y(n_492) );
O2A1O1Ixp33_ASAP7_75t_L g237 ( .A1(n_197), .A2(n_238), .B(n_239), .C(n_240), .Y(n_237) );
INVx1_ASAP7_75t_L g197 ( .A(n_198), .Y(n_197) );
NOR2xp33_ASAP7_75t_L g478 ( .A(n_198), .B(n_479), .Y(n_478) );
NOR2xp33_ASAP7_75t_L g487 ( .A(n_198), .B(n_488), .Y(n_487) );
INVx2_ASAP7_75t_L g226 ( .A(n_201), .Y(n_226) );
NAND2xp5_ASAP7_75t_SL g509 ( .A(n_201), .B(n_510), .Y(n_509) );
OA21x2_ASAP7_75t_L g257 ( .A1(n_203), .A2(n_258), .B(n_267), .Y(n_257) );
AOI221xp5_ASAP7_75t_L g373 ( .A1(n_204), .A2(n_374), .B1(n_376), .B2(n_378), .C(n_381), .Y(n_373) );
INVx2_ASAP7_75t_L g204 ( .A(n_205), .Y(n_204) );
OR2x2_ASAP7_75t_L g205 ( .A(n_206), .B(n_216), .Y(n_205) );
AND2x2_ASAP7_75t_L g347 ( .A(n_206), .B(n_328), .Y(n_347) );
NAND2xp5_ASAP7_75t_L g410 ( .A(n_206), .B(n_406), .Y(n_410) );
OR2x2_ASAP7_75t_L g431 ( .A(n_206), .B(n_432), .Y(n_431) );
NAND2xp5_ASAP7_75t_L g435 ( .A(n_206), .B(n_436), .Y(n_435) );
BUFx2_ASAP7_75t_L g206 ( .A(n_207), .Y(n_206) );
INVx5_ASAP7_75t_L g278 ( .A(n_207), .Y(n_278) );
AND2x2_ASAP7_75t_L g355 ( .A(n_207), .B(n_218), .Y(n_355) );
AND2x2_ASAP7_75t_L g416 ( .A(n_207), .B(n_295), .Y(n_416) );
AND2x2_ASAP7_75t_L g429 ( .A(n_207), .B(n_248), .Y(n_429) );
OR2x6_ASAP7_75t_L g207 ( .A(n_208), .B(n_214), .Y(n_207) );
NAND2xp5_ASAP7_75t_L g216 ( .A(n_217), .B(n_232), .Y(n_216) );
AND2x4_ASAP7_75t_L g255 ( .A(n_217), .B(n_256), .Y(n_255) );
AND2x2_ASAP7_75t_L g274 ( .A(n_217), .B(n_275), .Y(n_274) );
INVx2_ASAP7_75t_L g281 ( .A(n_217), .Y(n_281) );
AND2x2_ASAP7_75t_L g350 ( .A(n_217), .B(n_328), .Y(n_350) );
AND2x2_ASAP7_75t_L g360 ( .A(n_217), .B(n_278), .Y(n_360) );
HB1xp67_ASAP7_75t_L g368 ( .A(n_217), .Y(n_368) );
AND2x2_ASAP7_75t_L g380 ( .A(n_217), .B(n_257), .Y(n_380) );
NOR2xp33_ASAP7_75t_L g384 ( .A(n_217), .B(n_312), .Y(n_384) );
AND2x2_ASAP7_75t_L g421 ( .A(n_217), .B(n_416), .Y(n_421) );
NAND2xp5_ASAP7_75t_L g432 ( .A(n_217), .B(n_295), .Y(n_432) );
OR2x2_ASAP7_75t_L g434 ( .A(n_217), .B(n_370), .Y(n_434) );
INVx5_ASAP7_75t_L g217 ( .A(n_218), .Y(n_217) );
AND2x2_ASAP7_75t_L g320 ( .A(n_218), .B(n_321), .Y(n_320) );
AND2x2_ASAP7_75t_L g330 ( .A(n_218), .B(n_275), .Y(n_330) );
AND2x2_ASAP7_75t_L g342 ( .A(n_218), .B(n_257), .Y(n_342) );
HB1xp67_ASAP7_75t_L g372 ( .A(n_218), .Y(n_372) );
AND2x4_ASAP7_75t_L g406 ( .A(n_218), .B(n_256), .Y(n_406) );
OR2x6_ASAP7_75t_L g218 ( .A(n_219), .B(n_229), .Y(n_218) );
AOI21xp5_ASAP7_75t_SL g219 ( .A1(n_220), .A2(n_222), .B(n_227), .Y(n_219) );
AOI21xp5_ASAP7_75t_L g223 ( .A1(n_224), .A2(n_225), .B(n_226), .Y(n_223) );
INVx1_ASAP7_75t_L g227 ( .A(n_228), .Y(n_227) );
NOR2xp33_ASAP7_75t_L g533 ( .A(n_228), .B(n_534), .Y(n_533) );
NOR2xp33_ASAP7_75t_L g229 ( .A(n_230), .B(n_231), .Y(n_229) );
AO21x2_ASAP7_75t_L g450 ( .A1(n_231), .A2(n_451), .B(n_458), .Y(n_450) );
BUFx2_ASAP7_75t_L g254 ( .A(n_232), .Y(n_254) );
HB1xp67_ASAP7_75t_L g232 ( .A(n_233), .Y(n_232) );
INVx2_ASAP7_75t_L g295 ( .A(n_233), .Y(n_295) );
AND2x2_ASAP7_75t_L g328 ( .A(n_233), .B(n_257), .Y(n_328) );
INVx2_ASAP7_75t_L g233 ( .A(n_234), .Y(n_233) );
AND2x2_ASAP7_75t_L g275 ( .A(n_234), .B(n_257), .Y(n_275) );
BUFx2_ASAP7_75t_L g321 ( .A(n_234), .Y(n_321) );
NAND2xp5_ASAP7_75t_L g235 ( .A(n_236), .B(n_242), .Y(n_235) );
HB1xp67_ASAP7_75t_L g240 ( .A(n_241), .Y(n_240) );
INVx3_ASAP7_75t_L g499 ( .A(n_241), .Y(n_499) );
INVx1_ASAP7_75t_L g245 ( .A(n_246), .Y(n_245) );
NAND2xp5_ASAP7_75t_L g246 ( .A(n_247), .B(n_249), .Y(n_246) );
NAND2xp5_ASAP7_75t_L g408 ( .A(n_247), .B(n_329), .Y(n_408) );
INVx1_ASAP7_75t_L g247 ( .A(n_248), .Y(n_247) );
NAND2xp5_ASAP7_75t_L g272 ( .A(n_248), .B(n_271), .Y(n_272) );
NAND2xp5_ASAP7_75t_L g310 ( .A(n_248), .B(n_251), .Y(n_310) );
AND2x2_ASAP7_75t_L g365 ( .A(n_248), .B(n_301), .Y(n_365) );
AOI221xp5_ASAP7_75t_SL g302 ( .A1(n_249), .A2(n_303), .B1(n_311), .B2(n_313), .C(n_317), .Y(n_302) );
INVx2_ASAP7_75t_L g249 ( .A(n_250), .Y(n_249) );
OR2x2_ASAP7_75t_L g297 ( .A(n_250), .B(n_298), .Y(n_297) );
OR2x2_ASAP7_75t_L g338 ( .A(n_250), .B(n_339), .Y(n_338) );
OAI321xp33_ASAP7_75t_L g345 ( .A1(n_250), .A2(n_304), .A3(n_346), .B1(n_348), .B2(n_349), .C(n_351), .Y(n_345) );
NAND2xp5_ASAP7_75t_L g396 ( .A(n_251), .B(n_397), .Y(n_396) );
INVx1_ASAP7_75t_L g252 ( .A(n_253), .Y(n_252) );
NAND2xp5_ASAP7_75t_L g253 ( .A(n_254), .B(n_255), .Y(n_253) );
NAND2xp5_ASAP7_75t_L g424 ( .A(n_254), .B(n_406), .Y(n_424) );
AND2x2_ASAP7_75t_L g311 ( .A(n_255), .B(n_312), .Y(n_311) );
NAND2xp5_ASAP7_75t_L g314 ( .A(n_255), .B(n_315), .Y(n_314) );
HB1xp67_ASAP7_75t_L g287 ( .A(n_256), .Y(n_287) );
AND2x2_ASAP7_75t_L g294 ( .A(n_256), .B(n_295), .Y(n_294) );
NAND2xp5_ASAP7_75t_L g399 ( .A(n_256), .B(n_369), .Y(n_399) );
INVx1_ASAP7_75t_L g436 ( .A(n_256), .Y(n_436) );
INVx2_ASAP7_75t_L g256 ( .A(n_257), .Y(n_256) );
NOR2xp33_ASAP7_75t_L g263 ( .A(n_264), .B(n_265), .Y(n_263) );
NOR2xp33_ASAP7_75t_L g497 ( .A(n_265), .B(n_498), .Y(n_497) );
INVx2_ASAP7_75t_L g457 ( .A(n_266), .Y(n_457) );
AOI21xp5_ASAP7_75t_L g268 ( .A1(n_269), .A2(n_272), .B(n_273), .Y(n_268) );
INVx1_ASAP7_75t_SL g269 ( .A(n_270), .Y(n_269) );
A2O1A1Ixp33_ASAP7_75t_L g428 ( .A1(n_270), .A2(n_380), .B(n_429), .C(n_430), .Y(n_428) );
NAND2xp5_ASAP7_75t_L g288 ( .A(n_271), .B(n_289), .Y(n_288) );
NAND2xp5_ASAP7_75t_L g375 ( .A(n_271), .B(n_309), .Y(n_375) );
INVx1_ASAP7_75t_SL g273 ( .A(n_274), .Y(n_273) );
INVx1_ASAP7_75t_L g318 ( .A(n_275), .Y(n_318) );
NAND2xp5_ASAP7_75t_L g332 ( .A(n_275), .B(n_278), .Y(n_332) );
NOR2xp33_ASAP7_75t_L g341 ( .A(n_275), .B(n_342), .Y(n_341) );
NAND2xp5_ASAP7_75t_L g359 ( .A(n_275), .B(n_360), .Y(n_359) );
AOI22xp33_ASAP7_75t_L g276 ( .A1(n_277), .A2(n_279), .B1(n_291), .B2(n_296), .Y(n_276) );
HB1xp67_ASAP7_75t_L g277 ( .A(n_278), .Y(n_277) );
OR2x2_ASAP7_75t_L g292 ( .A(n_278), .B(n_293), .Y(n_292) );
AND2x2_ASAP7_75t_L g315 ( .A(n_278), .B(n_316), .Y(n_315) );
AND2x2_ASAP7_75t_L g327 ( .A(n_278), .B(n_328), .Y(n_327) );
NAND2xp5_ASAP7_75t_L g363 ( .A(n_278), .B(n_321), .Y(n_363) );
OR2x2_ASAP7_75t_L g370 ( .A(n_278), .B(n_295), .Y(n_370) );
NAND2xp5_ASAP7_75t_L g379 ( .A(n_278), .B(n_380), .Y(n_379) );
AND2x2_ASAP7_75t_L g420 ( .A(n_278), .B(n_406), .Y(n_420) );
OAI22xp33_ASAP7_75t_L g279 ( .A1(n_280), .A2(n_282), .B1(n_286), .B2(n_288), .Y(n_279) );
INVx1_ASAP7_75t_L g280 ( .A(n_281), .Y(n_280) );
AND2x2_ASAP7_75t_L g326 ( .A(n_281), .B(n_327), .Y(n_326) );
NAND2xp5_ASAP7_75t_L g282 ( .A(n_283), .B(n_285), .Y(n_282) );
INVx1_ASAP7_75t_SL g283 ( .A(n_284), .Y(n_283) );
OAI22xp33_ASAP7_75t_L g366 ( .A1(n_284), .A2(n_299), .B1(n_367), .B2(n_371), .Y(n_366) );
INVx1_ASAP7_75t_L g414 ( .A(n_285), .Y(n_414) );
INVx1_ASAP7_75t_L g286 ( .A(n_287), .Y(n_286) );
AOI221xp5_ASAP7_75t_L g325 ( .A1(n_289), .A2(n_326), .B1(n_329), .B2(n_330), .C(n_331), .Y(n_325) );
INVx1_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
OR2x2_ASAP7_75t_L g304 ( .A(n_290), .B(n_305), .Y(n_304) );
INVx1_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
INVx1_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
NAND2xp5_ASAP7_75t_L g392 ( .A(n_294), .B(n_360), .Y(n_392) );
HB1xp67_ASAP7_75t_L g312 ( .A(n_295), .Y(n_312) );
INVx1_ASAP7_75t_L g316 ( .A(n_295), .Y(n_316) );
NAND2xp33_ASAP7_75t_L g296 ( .A(n_297), .B(n_299), .Y(n_296) );
NAND2xp5_ASAP7_75t_L g299 ( .A(n_300), .B(n_301), .Y(n_299) );
INVx1_ASAP7_75t_L g334 ( .A(n_301), .Y(n_334) );
AND2x2_ASAP7_75t_L g343 ( .A(n_301), .B(n_344), .Y(n_343) );
NAND2xp33_ASAP7_75t_L g303 ( .A(n_304), .B(n_306), .Y(n_303) );
INVx2_ASAP7_75t_SL g306 ( .A(n_307), .Y(n_306) );
AND2x4_ASAP7_75t_L g307 ( .A(n_308), .B(n_309), .Y(n_307) );
AND2x2_ASAP7_75t_L g387 ( .A(n_308), .B(n_388), .Y(n_387) );
INVx2_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
AOI221xp5_ASAP7_75t_L g336 ( .A1(n_311), .A2(n_337), .B1(n_340), .B2(n_343), .C(n_345), .Y(n_336) );
INVx1_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
NAND2xp5_ASAP7_75t_L g371 ( .A(n_315), .B(n_372), .Y(n_371) );
AOI21xp33_ASAP7_75t_SL g317 ( .A1(n_318), .A2(n_319), .B(n_322), .Y(n_317) );
INVx2_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
CKINVDCx16_ASAP7_75t_R g419 ( .A(n_322), .Y(n_419) );
OR2x2_ASAP7_75t_L g322 ( .A(n_323), .B(n_324), .Y(n_322) );
OR2x2_ASAP7_75t_L g361 ( .A(n_324), .B(n_362), .Y(n_361) );
INVx1_ASAP7_75t_SL g382 ( .A(n_327), .Y(n_382) );
NAND2xp5_ASAP7_75t_L g427 ( .A(n_327), .B(n_387), .Y(n_427) );
NAND2xp5_ASAP7_75t_L g351 ( .A(n_330), .B(n_352), .Y(n_351) );
NOR2xp33_ASAP7_75t_L g331 ( .A(n_332), .B(n_333), .Y(n_331) );
NAND4xp25_ASAP7_75t_L g335 ( .A(n_336), .B(n_354), .C(n_373), .D(n_386), .Y(n_335) );
INVx1_ASAP7_75t_SL g337 ( .A(n_338), .Y(n_337) );
INVx1_ASAP7_75t_SL g344 ( .A(n_339), .Y(n_344) );
INVxp67_ASAP7_75t_L g340 ( .A(n_341), .Y(n_340) );
INVx1_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
OR2x2_ASAP7_75t_L g377 ( .A(n_348), .B(n_353), .Y(n_377) );
INVxp67_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
AOI211xp5_ASAP7_75t_L g354 ( .A1(n_355), .A2(n_356), .B(n_358), .C(n_366), .Y(n_354) );
AOI211xp5_ASAP7_75t_L g425 ( .A1(n_356), .A2(n_398), .B(n_426), .C(n_433), .Y(n_425) );
INVx1_ASAP7_75t_SL g385 ( .A(n_357), .Y(n_385) );
OAI22xp5_ASAP7_75t_L g358 ( .A1(n_359), .A2(n_361), .B1(n_363), .B2(n_364), .Y(n_358) );
INVx1_ASAP7_75t_L g389 ( .A(n_363), .Y(n_389) );
INVx1_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
NAND2xp5_ASAP7_75t_L g367 ( .A(n_368), .B(n_369), .Y(n_367) );
NAND2xp5_ASAP7_75t_L g405 ( .A(n_369), .B(n_406), .Y(n_405) );
NAND2xp5_ASAP7_75t_L g413 ( .A(n_369), .B(n_380), .Y(n_413) );
INVx2_ASAP7_75t_SL g369 ( .A(n_370), .Y(n_369) );
INVx1_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
INVx1_ASAP7_75t_SL g376 ( .A(n_377), .Y(n_376) );
INVx1_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
INVx1_ASAP7_75t_L g390 ( .A(n_380), .Y(n_390) );
AOI21xp33_ASAP7_75t_L g381 ( .A1(n_382), .A2(n_383), .B(n_385), .Y(n_381) );
INVxp33_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
AOI322xp5_ASAP7_75t_L g386 ( .A1(n_387), .A2(n_389), .A3(n_390), .B1(n_391), .B2(n_393), .C1(n_395), .C2(n_398), .Y(n_386) );
INVxp67_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
INVx1_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
INVx1_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
INVx1_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
NAND3xp33_ASAP7_75t_SL g400 ( .A(n_401), .B(n_418), .C(n_425), .Y(n_400) );
AOI221xp5_ASAP7_75t_L g401 ( .A1(n_402), .A2(n_404), .B1(n_407), .B2(n_409), .C(n_411), .Y(n_401) );
INVx1_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
INVx1_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
INVx1_ASAP7_75t_SL g417 ( .A(n_406), .Y(n_417) );
INVx1_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
INVxp67_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
OAI22xp33_ASAP7_75t_L g411 ( .A1(n_412), .A2(n_413), .B1(n_414), .B2(n_415), .Y(n_411) );
NAND2xp5_ASAP7_75t_L g415 ( .A(n_416), .B(n_417), .Y(n_415) );
AOI221xp5_ASAP7_75t_L g418 ( .A1(n_419), .A2(n_420), .B1(n_421), .B2(n_422), .C(n_423), .Y(n_418) );
NAND2xp33_ASAP7_75t_L g426 ( .A(n_427), .B(n_428), .Y(n_426) );
INVxp67_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
INVx2_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
INVx2_ASAP7_75t_L g715 ( .A(n_438), .Y(n_715) );
INVx1_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
INVx2_ASAP7_75t_L g724 ( .A(n_440), .Y(n_724) );
AND2x2_ASAP7_75t_L g440 ( .A(n_441), .B(n_442), .Y(n_440) );
INVx2_ASAP7_75t_L g717 ( .A(n_443), .Y(n_717) );
OR2x2_ASAP7_75t_SL g443 ( .A(n_444), .B(n_664), .Y(n_443) );
NAND5xp2_ASAP7_75t_L g444 ( .A(n_445), .B(n_576), .C(n_614), .D(n_635), .E(n_652), .Y(n_444) );
NOR3xp33_ASAP7_75t_L g445 ( .A(n_446), .B(n_548), .C(n_569), .Y(n_445) );
OAI221xp5_ASAP7_75t_SL g446 ( .A1(n_447), .A2(n_490), .B1(n_514), .B2(n_535), .C(n_539), .Y(n_446) );
NAND2xp5_ASAP7_75t_L g447 ( .A(n_448), .B(n_460), .Y(n_447) );
INVx1_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
NAND2xp5_ASAP7_75t_L g556 ( .A(n_449), .B(n_537), .Y(n_556) );
OR2x2_ASAP7_75t_L g583 ( .A(n_449), .B(n_473), .Y(n_583) );
AND2x2_ASAP7_75t_L g597 ( .A(n_449), .B(n_473), .Y(n_597) );
NOR2xp33_ASAP7_75t_L g611 ( .A(n_449), .B(n_463), .Y(n_611) );
AND2x2_ASAP7_75t_L g649 ( .A(n_449), .B(n_613), .Y(n_649) );
AND2x2_ASAP7_75t_L g678 ( .A(n_449), .B(n_588), .Y(n_678) );
NAND2xp5_ASAP7_75t_L g695 ( .A(n_449), .B(n_560), .Y(n_695) );
INVx4_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
AND2x2_ASAP7_75t_L g575 ( .A(n_450), .B(n_472), .Y(n_575) );
BUFx3_ASAP7_75t_L g600 ( .A(n_450), .Y(n_600) );
AND2x2_ASAP7_75t_L g629 ( .A(n_450), .B(n_473), .Y(n_629) );
AND3x2_ASAP7_75t_L g642 ( .A(n_450), .B(n_643), .C(n_644), .Y(n_642) );
INVx1_ASAP7_75t_L g565 ( .A(n_460), .Y(n_565) );
AND2x2_ASAP7_75t_L g460 ( .A(n_461), .B(n_472), .Y(n_460) );
AOI32xp33_ASAP7_75t_L g620 ( .A1(n_461), .A2(n_572), .A3(n_621), .B1(n_624), .B2(n_625), .Y(n_620) );
INVx1_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
AND2x2_ASAP7_75t_L g547 ( .A(n_462), .B(n_472), .Y(n_547) );
NAND2xp5_ASAP7_75t_SL g618 ( .A(n_462), .B(n_575), .Y(n_618) );
AND2x2_ASAP7_75t_L g625 ( .A(n_462), .B(n_597), .Y(n_625) );
OR2x2_ASAP7_75t_L g631 ( .A(n_462), .B(n_632), .Y(n_631) );
NAND2xp5_ASAP7_75t_L g656 ( .A(n_462), .B(n_586), .Y(n_656) );
OR2x2_ASAP7_75t_L g674 ( .A(n_462), .B(n_502), .Y(n_674) );
BUFx3_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
AND2x2_ASAP7_75t_L g538 ( .A(n_463), .B(n_482), .Y(n_538) );
INVx2_ASAP7_75t_L g560 ( .A(n_463), .Y(n_560) );
OR2x2_ASAP7_75t_L g582 ( .A(n_463), .B(n_482), .Y(n_582) );
AND2x2_ASAP7_75t_L g587 ( .A(n_463), .B(n_588), .Y(n_587) );
NAND2xp5_ASAP7_75t_L g638 ( .A(n_463), .B(n_639), .Y(n_638) );
AND2x2_ASAP7_75t_L g643 ( .A(n_463), .B(n_537), .Y(n_643) );
INVx1_ASAP7_75t_SL g694 ( .A(n_472), .Y(n_694) );
AND2x2_ASAP7_75t_L g472 ( .A(n_473), .B(n_482), .Y(n_472) );
INVx1_ASAP7_75t_SL g537 ( .A(n_473), .Y(n_537) );
HB1xp67_ASAP7_75t_L g586 ( .A(n_473), .Y(n_586) );
NAND2xp5_ASAP7_75t_L g622 ( .A(n_473), .B(n_623), .Y(n_622) );
NAND3xp33_ASAP7_75t_L g689 ( .A(n_473), .B(n_560), .C(n_678), .Y(n_689) );
INVx2_ASAP7_75t_L g588 ( .A(n_482), .Y(n_588) );
HB1xp67_ASAP7_75t_L g602 ( .A(n_482), .Y(n_602) );
NAND2xp5_ASAP7_75t_L g490 ( .A(n_491), .B(n_501), .Y(n_490) );
INVx1_ASAP7_75t_L g624 ( .A(n_491), .Y(n_624) );
INVx1_ASAP7_75t_L g491 ( .A(n_492), .Y(n_491) );
AND2x2_ASAP7_75t_L g542 ( .A(n_492), .B(n_525), .Y(n_542) );
INVx2_ASAP7_75t_L g559 ( .A(n_492), .Y(n_559) );
AND2x2_ASAP7_75t_L g564 ( .A(n_492), .B(n_526), .Y(n_564) );
AND2x2_ASAP7_75t_L g579 ( .A(n_492), .B(n_515), .Y(n_579) );
AND2x2_ASAP7_75t_L g591 ( .A(n_492), .B(n_563), .Y(n_591) );
NAND2xp5_ASAP7_75t_L g606 ( .A(n_501), .B(n_607), .Y(n_606) );
NAND2x1p5_ASAP7_75t_L g663 ( .A(n_501), .B(n_564), .Y(n_663) );
NAND2xp5_ASAP7_75t_L g682 ( .A(n_501), .B(n_683), .Y(n_682) );
NAND2xp5_ASAP7_75t_L g686 ( .A(n_501), .B(n_558), .Y(n_686) );
BUFx3_ASAP7_75t_L g501 ( .A(n_502), .Y(n_501) );
OR2x2_ASAP7_75t_L g524 ( .A(n_502), .B(n_525), .Y(n_524) );
NAND2xp5_ASAP7_75t_L g541 ( .A(n_502), .B(n_542), .Y(n_541) );
AND2x2_ASAP7_75t_L g568 ( .A(n_502), .B(n_515), .Y(n_568) );
AND2x2_ASAP7_75t_L g594 ( .A(n_502), .B(n_525), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g633 ( .A(n_502), .B(n_634), .Y(n_633) );
OA21x2_ASAP7_75t_L g502 ( .A1(n_503), .A2(n_506), .B(n_513), .Y(n_502) );
INVx1_ASAP7_75t_L g503 ( .A(n_504), .Y(n_503) );
AO21x2_ASAP7_75t_L g552 ( .A1(n_504), .A2(n_553), .B(n_554), .Y(n_552) );
INVx1_ASAP7_75t_L g504 ( .A(n_505), .Y(n_504) );
INVx1_ASAP7_75t_L g553 ( .A(n_506), .Y(n_553) );
INVx1_ASAP7_75t_L g554 ( .A(n_513), .Y(n_554) );
OR2x2_ASAP7_75t_L g514 ( .A(n_515), .B(n_524), .Y(n_514) );
NAND2xp5_ASAP7_75t_L g544 ( .A(n_515), .B(n_545), .Y(n_544) );
AND2x4_ASAP7_75t_L g558 ( .A(n_515), .B(n_559), .Y(n_558) );
INVx3_ASAP7_75t_SL g563 ( .A(n_515), .Y(n_563) );
NAND2xp5_ASAP7_75t_L g616 ( .A(n_515), .B(n_550), .Y(n_616) );
OR2x2_ASAP7_75t_L g626 ( .A(n_515), .B(n_552), .Y(n_626) );
NAND2xp5_ASAP7_75t_L g654 ( .A(n_515), .B(n_594), .Y(n_654) );
OR2x2_ASAP7_75t_L g684 ( .A(n_515), .B(n_525), .Y(n_684) );
AND2x2_ASAP7_75t_L g688 ( .A(n_515), .B(n_526), .Y(n_688) );
NAND2xp5_ASAP7_75t_SL g701 ( .A(n_515), .B(n_564), .Y(n_701) );
AND2x2_ASAP7_75t_L g708 ( .A(n_515), .B(n_590), .Y(n_708) );
OR2x6_ASAP7_75t_L g515 ( .A(n_516), .B(n_522), .Y(n_515) );
INVx1_ASAP7_75t_SL g651 ( .A(n_524), .Y(n_651) );
AND2x2_ASAP7_75t_L g590 ( .A(n_525), .B(n_552), .Y(n_590) );
AND2x2_ASAP7_75t_L g604 ( .A(n_525), .B(n_559), .Y(n_604) );
AND2x2_ASAP7_75t_L g607 ( .A(n_525), .B(n_563), .Y(n_607) );
INVx1_ASAP7_75t_L g634 ( .A(n_525), .Y(n_634) );
INVx2_ASAP7_75t_SL g525 ( .A(n_526), .Y(n_525) );
BUFx2_ASAP7_75t_L g546 ( .A(n_526), .Y(n_546) );
NAND2xp5_ASAP7_75t_L g535 ( .A(n_536), .B(n_538), .Y(n_535) );
A2O1A1Ixp33_ASAP7_75t_L g705 ( .A1(n_536), .A2(n_582), .B(n_706), .C(n_707), .Y(n_705) );
HB1xp67_ASAP7_75t_L g536 ( .A(n_537), .Y(n_536) );
AND2x2_ASAP7_75t_L g612 ( .A(n_537), .B(n_613), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g570 ( .A(n_538), .B(n_555), .Y(n_570) );
AND2x2_ASAP7_75t_L g596 ( .A(n_538), .B(n_597), .Y(n_596) );
OAI21xp5_ASAP7_75t_SL g539 ( .A1(n_540), .A2(n_543), .B(n_547), .Y(n_539) );
INVx1_ASAP7_75t_L g540 ( .A(n_541), .Y(n_540) );
NOR2xp33_ASAP7_75t_L g640 ( .A(n_541), .B(n_641), .Y(n_640) );
AND2x2_ASAP7_75t_L g567 ( .A(n_542), .B(n_568), .Y(n_567) );
NAND2xp5_ASAP7_75t_L g608 ( .A(n_542), .B(n_563), .Y(n_608) );
AND2x2_ASAP7_75t_L g699 ( .A(n_542), .B(n_550), .Y(n_699) );
INVxp67_ASAP7_75t_L g543 ( .A(n_544), .Y(n_543) );
INVx1_ASAP7_75t_L g545 ( .A(n_546), .Y(n_545) );
AND2x2_ASAP7_75t_L g572 ( .A(n_546), .B(n_559), .Y(n_572) );
OR2x2_ASAP7_75t_L g573 ( .A(n_546), .B(n_557), .Y(n_573) );
OAI322xp33_ASAP7_75t_L g548 ( .A1(n_549), .A2(n_556), .A3(n_557), .B1(n_560), .B2(n_561), .C1(n_565), .C2(n_566), .Y(n_548) );
NAND2xp5_ASAP7_75t_L g549 ( .A(n_550), .B(n_555), .Y(n_549) );
AND2x2_ASAP7_75t_L g660 ( .A(n_550), .B(n_572), .Y(n_660) );
NAND2xp5_ASAP7_75t_L g706 ( .A(n_550), .B(n_624), .Y(n_706) );
INVx2_ASAP7_75t_L g550 ( .A(n_551), .Y(n_550) );
INVx1_ASAP7_75t_SL g551 ( .A(n_552), .Y(n_551) );
AND2x2_ASAP7_75t_L g603 ( .A(n_552), .B(n_604), .Y(n_603) );
INVx1_ASAP7_75t_L g555 ( .A(n_556), .Y(n_555) );
OR2x2_ASAP7_75t_L g669 ( .A(n_556), .B(n_582), .Y(n_669) );
NAND2xp5_ASAP7_75t_L g650 ( .A(n_557), .B(n_651), .Y(n_650) );
INVx3_ASAP7_75t_L g557 ( .A(n_558), .Y(n_557) );
NAND2xp5_ASAP7_75t_L g647 ( .A(n_558), .B(n_590), .Y(n_647) );
AND2x2_ASAP7_75t_L g593 ( .A(n_559), .B(n_563), .Y(n_593) );
AND2x2_ASAP7_75t_L g601 ( .A(n_560), .B(n_602), .Y(n_601) );
A2O1A1Ixp33_ASAP7_75t_L g698 ( .A1(n_560), .A2(n_639), .B(n_699), .C(n_700), .Y(n_698) );
AOI21xp33_ASAP7_75t_L g671 ( .A1(n_561), .A2(n_574), .B(n_672), .Y(n_671) );
INVx1_ASAP7_75t_SL g561 ( .A(n_562), .Y(n_561) );
AND2x2_ASAP7_75t_L g562 ( .A(n_563), .B(n_564), .Y(n_562) );
NAND2xp5_ASAP7_75t_L g630 ( .A(n_563), .B(n_590), .Y(n_630) );
AND2x2_ASAP7_75t_L g636 ( .A(n_563), .B(n_604), .Y(n_636) );
AND2x2_ASAP7_75t_L g670 ( .A(n_563), .B(n_572), .Y(n_670) );
NOR2xp33_ASAP7_75t_L g578 ( .A(n_564), .B(n_579), .Y(n_578) );
INVx2_ASAP7_75t_SL g680 ( .A(n_564), .Y(n_680) );
INVx1_ASAP7_75t_L g566 ( .A(n_567), .Y(n_566) );
AOI22xp5_ASAP7_75t_L g595 ( .A1(n_568), .A2(n_596), .B1(n_598), .B2(n_603), .Y(n_595) );
OAI22xp5_ASAP7_75t_SL g569 ( .A1(n_570), .A2(n_571), .B1(n_573), .B2(n_574), .Y(n_569) );
OAI22xp33_ASAP7_75t_L g605 ( .A1(n_570), .A2(n_606), .B1(n_608), .B2(n_609), .Y(n_605) );
INVxp67_ASAP7_75t_L g571 ( .A(n_572), .Y(n_571) );
INVx1_ASAP7_75t_SL g574 ( .A(n_575), .Y(n_574) );
AOI221xp5_ASAP7_75t_L g676 ( .A1(n_575), .A2(n_677), .B1(n_679), .B2(n_681), .C(n_685), .Y(n_676) );
AOI211xp5_ASAP7_75t_L g576 ( .A1(n_577), .A2(n_580), .B(n_584), .C(n_605), .Y(n_576) );
INVxp67_ASAP7_75t_L g577 ( .A(n_578), .Y(n_577) );
INVx1_ASAP7_75t_L g580 ( .A(n_581), .Y(n_580) );
OR2x2_ASAP7_75t_L g581 ( .A(n_582), .B(n_583), .Y(n_581) );
OR2x2_ASAP7_75t_L g646 ( .A(n_582), .B(n_599), .Y(n_646) );
INVx1_ASAP7_75t_L g697 ( .A(n_582), .Y(n_697) );
OAI221xp5_ASAP7_75t_L g584 ( .A1(n_583), .A2(n_585), .B1(n_589), .B2(n_592), .C(n_595), .Y(n_584) );
INVx2_ASAP7_75t_SL g639 ( .A(n_583), .Y(n_639) );
NAND2xp5_ASAP7_75t_L g585 ( .A(n_586), .B(n_587), .Y(n_585) );
INVx1_ASAP7_75t_L g704 ( .A(n_586), .Y(n_704) );
AND2x2_ASAP7_75t_L g628 ( .A(n_587), .B(n_629), .Y(n_628) );
INVx2_ASAP7_75t_L g613 ( .A(n_588), .Y(n_613) );
NAND2xp5_ASAP7_75t_L g589 ( .A(n_590), .B(n_591), .Y(n_589) );
INVx1_ASAP7_75t_L g675 ( .A(n_591), .Y(n_675) );
NAND2xp5_ASAP7_75t_L g592 ( .A(n_593), .B(n_594), .Y(n_592) );
AND2x2_ASAP7_75t_L g598 ( .A(n_599), .B(n_601), .Y(n_598) );
NOR2xp33_ASAP7_75t_L g700 ( .A(n_599), .B(n_701), .Y(n_700) );
CKINVDCx16_ASAP7_75t_R g599 ( .A(n_600), .Y(n_599) );
INVxp67_ASAP7_75t_L g644 ( .A(n_602), .Y(n_644) );
O2A1O1Ixp33_ASAP7_75t_L g614 ( .A1(n_603), .A2(n_615), .B(n_617), .C(n_619), .Y(n_614) );
INVx1_ASAP7_75t_L g692 ( .A(n_606), .Y(n_692) );
INVx1_ASAP7_75t_L g609 ( .A(n_610), .Y(n_609) );
NOR2xp33_ASAP7_75t_L g667 ( .A(n_610), .B(n_668), .Y(n_667) );
AND2x2_ASAP7_75t_L g610 ( .A(n_611), .B(n_612), .Y(n_610) );
INVx2_ASAP7_75t_L g623 ( .A(n_613), .Y(n_623) );
INVx1_ASAP7_75t_L g615 ( .A(n_616), .Y(n_615) );
INVx1_ASAP7_75t_L g617 ( .A(n_618), .Y(n_617) );
OAI222xp33_ASAP7_75t_L g619 ( .A1(n_620), .A2(n_626), .B1(n_627), .B2(n_630), .C1(n_631), .C2(n_633), .Y(n_619) );
INVx1_ASAP7_75t_L g621 ( .A(n_622), .Y(n_621) );
INVx1_ASAP7_75t_SL g659 ( .A(n_623), .Y(n_659) );
NOR2xp33_ASAP7_75t_L g679 ( .A(n_626), .B(n_680), .Y(n_679) );
NAND2xp33_ASAP7_75t_SL g657 ( .A(n_627), .B(n_658), .Y(n_657) );
INVx1_ASAP7_75t_SL g627 ( .A(n_628), .Y(n_627) );
INVx1_ASAP7_75t_SL g632 ( .A(n_629), .Y(n_632) );
AND2x2_ASAP7_75t_L g696 ( .A(n_629), .B(n_697), .Y(n_696) );
OR2x2_ASAP7_75t_L g662 ( .A(n_632), .B(n_659), .Y(n_662) );
INVx1_ASAP7_75t_L g691 ( .A(n_633), .Y(n_691) );
AOI211xp5_ASAP7_75t_L g635 ( .A1(n_636), .A2(n_637), .B(n_640), .C(n_645), .Y(n_635) );
INVx1_ASAP7_75t_L g637 ( .A(n_638), .Y(n_637) );
NAND2xp5_ASAP7_75t_L g658 ( .A(n_639), .B(n_659), .Y(n_658) );
INVx2_ASAP7_75t_SL g641 ( .A(n_642), .Y(n_641) );
AOI322xp5_ASAP7_75t_L g690 ( .A1(n_642), .A2(n_670), .A3(n_675), .B1(n_691), .B2(n_692), .C1(n_693), .C2(n_696), .Y(n_690) );
AND2x2_ASAP7_75t_L g677 ( .A(n_643), .B(n_678), .Y(n_677) );
OAI22xp33_ASAP7_75t_L g645 ( .A1(n_646), .A2(n_647), .B1(n_648), .B2(n_650), .Y(n_645) );
INVxp33_ASAP7_75t_L g648 ( .A(n_649), .Y(n_648) );
AOI221xp5_ASAP7_75t_L g652 ( .A1(n_653), .A2(n_655), .B1(n_657), .B2(n_660), .C(n_661), .Y(n_652) );
INVx1_ASAP7_75t_L g653 ( .A(n_654), .Y(n_653) );
INVx1_ASAP7_75t_L g655 ( .A(n_656), .Y(n_655) );
NOR2xp33_ASAP7_75t_L g661 ( .A(n_662), .B(n_663), .Y(n_661) );
NAND5xp2_ASAP7_75t_L g664 ( .A(n_665), .B(n_676), .C(n_690), .D(n_698), .E(n_702), .Y(n_664) );
AOI21xp5_ASAP7_75t_L g665 ( .A1(n_666), .A2(n_670), .B(n_671), .Y(n_665) );
INVxp67_ASAP7_75t_L g666 ( .A(n_667), .Y(n_666) );
INVx2_ASAP7_75t_L g668 ( .A(n_669), .Y(n_668) );
INVxp33_ASAP7_75t_L g672 ( .A(n_673), .Y(n_672) );
NOR2xp33_ASAP7_75t_L g673 ( .A(n_674), .B(n_675), .Y(n_673) );
A2O1A1Ixp33_ASAP7_75t_L g702 ( .A1(n_678), .A2(n_703), .B(n_704), .C(n_705), .Y(n_702) );
AOI31xp33_ASAP7_75t_L g685 ( .A1(n_680), .A2(n_686), .A3(n_687), .B(n_689), .Y(n_685) );
INVx1_ASAP7_75t_L g681 ( .A(n_682), .Y(n_681) );
INVx1_ASAP7_75t_L g683 ( .A(n_684), .Y(n_683) );
INVx1_ASAP7_75t_L g687 ( .A(n_688), .Y(n_687) );
NOR2xp33_ASAP7_75t_L g693 ( .A(n_694), .B(n_695), .Y(n_693) );
INVx1_ASAP7_75t_L g703 ( .A(n_701), .Y(n_703) );
INVx1_ASAP7_75t_L g707 ( .A(n_708), .Y(n_707) );
INVx2_ASAP7_75t_L g709 ( .A(n_710), .Y(n_709) );
INVx2_ASAP7_75t_L g718 ( .A(n_710), .Y(n_718) );
INVx1_ASAP7_75t_L g710 ( .A(n_711), .Y(n_710) );
INVxp67_ASAP7_75t_L g713 ( .A(n_714), .Y(n_713) );
OAI22x1_ASAP7_75t_SL g714 ( .A1(n_715), .A2(n_716), .B1(n_717), .B2(n_718), .Y(n_714) );
INVx1_ASAP7_75t_SL g720 ( .A(n_721), .Y(n_720) );
INVx1_ASAP7_75t_L g721 ( .A(n_722), .Y(n_721) );
INVx2_ASAP7_75t_L g722 ( .A(n_723), .Y(n_722) );
BUFx2_ASAP7_75t_L g725 ( .A(n_726), .Y(n_725) );
INVx2_ASAP7_75t_L g726 ( .A(n_727), .Y(n_726) );
INVx1_ASAP7_75t_L g739 ( .A(n_727), .Y(n_739) );
INVxp67_ASAP7_75t_L g728 ( .A(n_729), .Y(n_728) );
NAND2xp5_ASAP7_75t_SL g729 ( .A(n_730), .B(n_735), .Y(n_729) );
INVx1_ASAP7_75t_L g731 ( .A(n_732), .Y(n_731) );
INVx1_ASAP7_75t_SL g735 ( .A(n_736), .Y(n_735) );
INVx1_ASAP7_75t_SL g736 ( .A(n_737), .Y(n_736) );
INVx1_ASAP7_75t_SL g743 ( .A(n_737), .Y(n_743) );
INVx1_ASAP7_75t_L g738 ( .A(n_739), .Y(n_738) );
NOR2xp33_ASAP7_75t_L g740 ( .A(n_741), .B(n_742), .Y(n_740) );
INVx1_ASAP7_75t_SL g742 ( .A(n_743), .Y(n_742) );
endmodule