module fake_jpeg_22229_n_339 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_339);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_339;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_256;
wire n_221;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVxp67_ASAP7_75t_L g17 ( 
.A(n_16),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

INVx6_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

INVx6_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

BUFx2_ASAP7_75t_L g22 ( 
.A(n_16),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_11),
.Y(n_24)
);

BUFx12_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_12),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_15),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_0),
.B(n_8),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_1),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_9),
.Y(n_34)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_9),
.Y(n_35)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_4),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_24),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_37),
.B(n_39),
.Y(n_50)
);

INVx11_ASAP7_75t_L g38 ( 
.A(n_25),
.Y(n_38)
);

INVx8_ASAP7_75t_L g55 ( 
.A(n_38),
.Y(n_55)
);

INVxp67_ASAP7_75t_L g39 ( 
.A(n_35),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_22),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_40),
.B(n_44),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_19),
.Y(n_41)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_41),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_19),
.Y(n_42)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_42),
.Y(n_60)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_23),
.Y(n_43)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_43),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_24),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_19),
.Y(n_45)
);

INVx5_ASAP7_75t_L g52 ( 
.A(n_45),
.Y(n_52)
);

INVx5_ASAP7_75t_L g46 ( 
.A(n_20),
.Y(n_46)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_46),
.Y(n_58)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_36),
.Y(n_47)
);

INVx11_ASAP7_75t_L g57 ( 
.A(n_47),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_19),
.Y(n_48)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_48),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g49 ( 
.A1(n_46),
.A2(n_21),
.B1(n_20),
.B2(n_29),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_49),
.A2(n_34),
.B1(n_29),
.B2(n_21),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_37),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_SL g70 ( 
.A(n_51),
.B(n_59),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_43),
.B(n_40),
.Y(n_53)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_53),
.B(n_30),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_46),
.A2(n_21),
.B1(n_20),
.B2(n_36),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_54),
.A2(n_49),
.B1(n_34),
.B2(n_43),
.Y(n_95)
);

OR2x2_ASAP7_75t_L g59 ( 
.A(n_45),
.B(n_19),
.Y(n_59)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_45),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_62),
.B(n_48),
.Y(n_76)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_45),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_64),
.B(n_40),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_37),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_65),
.B(n_44),
.Y(n_75)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_57),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_67),
.B(n_69),
.Y(n_101)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_53),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_68),
.B(n_73),
.Y(n_99)
);

BUFx12_ASAP7_75t_L g69 ( 
.A(n_52),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_71),
.A2(n_95),
.B1(n_47),
.B2(n_55),
.Y(n_122)
);

INVx1_ASAP7_75t_SL g104 ( 
.A(n_72),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_51),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_56),
.Y(n_74)
);

INVx6_ASAP7_75t_L g121 ( 
.A(n_74),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_SL g119 ( 
.A(n_75),
.B(n_94),
.Y(n_119)
);

AND2x2_ASAP7_75t_L g117 ( 
.A(n_76),
.B(n_81),
.Y(n_117)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_57),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_77),
.B(n_80),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_53),
.B(n_48),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_78),
.B(n_87),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_65),
.B(n_44),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_79),
.B(n_83),
.Y(n_112)
);

BUFx8_ASAP7_75t_L g80 ( 
.A(n_57),
.Y(n_80)
);

BUFx12f_ASAP7_75t_L g82 ( 
.A(n_62),
.Y(n_82)
);

CKINVDCx14_ASAP7_75t_R g113 ( 
.A(n_82),
.Y(n_113)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_61),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_58),
.A2(n_29),
.B1(n_34),
.B2(n_36),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_84),
.A2(n_89),
.B1(n_91),
.B2(n_55),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_61),
.B(n_25),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_SL g120 ( 
.A(n_85),
.B(n_92),
.Y(n_120)
);

BUFx10_ASAP7_75t_L g86 ( 
.A(n_55),
.Y(n_86)
);

BUFx3_ASAP7_75t_L g106 ( 
.A(n_86),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_59),
.B(n_48),
.Y(n_87)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_58),
.Y(n_88)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_88),
.Y(n_103)
);

INVx8_ASAP7_75t_L g89 ( 
.A(n_66),
.Y(n_89)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_58),
.Y(n_90)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_90),
.Y(n_124)
);

INVx6_ASAP7_75t_L g91 ( 
.A(n_66),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_50),
.B(n_25),
.Y(n_92)
);

BUFx2_ASAP7_75t_L g93 ( 
.A(n_63),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_93),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_50),
.B(n_25),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_59),
.B(n_42),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_96),
.B(n_62),
.C(n_64),
.Y(n_116)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_49),
.Y(n_97)
);

OAI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_97),
.A2(n_66),
.B1(n_47),
.B2(n_63),
.Y(n_111)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_89),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_98),
.B(n_100),
.Y(n_132)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_69),
.Y(n_100)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_69),
.Y(n_102)
);

INVx13_ASAP7_75t_L g155 ( 
.A(n_102),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_74),
.Y(n_105)
);

BUFx3_ASAP7_75t_L g149 ( 
.A(n_105),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_82),
.Y(n_108)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_108),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_97),
.A2(n_55),
.B1(n_35),
.B2(n_43),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_109),
.A2(n_122),
.B1(n_54),
.B2(n_88),
.Y(n_129)
);

A2O1A1Ixp33_ASAP7_75t_L g110 ( 
.A1(n_87),
.A2(n_59),
.B(n_28),
.C(n_45),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_SL g131 ( 
.A(n_110),
.B(n_75),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_111),
.B(n_90),
.Y(n_133)
);

AO22x2_ASAP7_75t_L g114 ( 
.A1(n_81),
.A2(n_96),
.B1(n_71),
.B2(n_45),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_114),
.A2(n_38),
.B1(n_52),
.B2(n_60),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_116),
.B(n_128),
.C(n_33),
.Y(n_145)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_82),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_118),
.Y(n_135)
);

A2O1A1Ixp33_ASAP7_75t_SL g125 ( 
.A1(n_70),
.A2(n_18),
.B(n_33),
.C(n_30),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_125),
.A2(n_126),
.B1(n_127),
.B2(n_91),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_SL g127 ( 
.A1(n_83),
.A2(n_52),
.B1(n_56),
.B2(n_60),
.Y(n_127)
);

MAJx2_ASAP7_75t_L g128 ( 
.A(n_81),
.B(n_68),
.C(n_70),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_129),
.A2(n_138),
.B1(n_120),
.B2(n_104),
.Y(n_162)
);

AND2x6_ASAP7_75t_L g130 ( 
.A(n_114),
.B(n_73),
.Y(n_130)
);

NOR3xp33_ASAP7_75t_L g166 ( 
.A(n_130),
.B(n_142),
.C(n_144),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_131),
.B(n_150),
.Y(n_165)
);

O2A1O1Ixp33_ASAP7_75t_L g181 ( 
.A1(n_133),
.A2(n_106),
.B(n_80),
.C(n_30),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_136),
.A2(n_121),
.B1(n_38),
.B2(n_109),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_123),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_137),
.Y(n_179)
);

O2A1O1Ixp33_ASAP7_75t_L g138 ( 
.A1(n_125),
.A2(n_76),
.B(n_82),
.C(n_78),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_139),
.A2(n_152),
.B1(n_101),
.B2(n_100),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_L g140 ( 
.A1(n_115),
.A2(n_32),
.B(n_18),
.Y(n_140)
);

AOI21xp5_ASAP7_75t_SL g160 ( 
.A1(n_140),
.A2(n_125),
.B(n_18),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_114),
.A2(n_35),
.B1(n_17),
.B2(n_33),
.Y(n_141)
);

INVxp67_ASAP7_75t_L g164 ( 
.A(n_141),
.Y(n_164)
);

AND2x6_ASAP7_75t_L g142 ( 
.A(n_114),
.B(n_15),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_115),
.B(n_86),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_143),
.B(n_146),
.Y(n_167)
);

AND2x6_ASAP7_75t_L g144 ( 
.A(n_117),
.B(n_15),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_145),
.B(n_125),
.C(n_113),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_117),
.B(n_86),
.Y(n_146)
);

AND2x2_ASAP7_75t_L g147 ( 
.A(n_117),
.B(n_116),
.Y(n_147)
);

AOI21xp5_ASAP7_75t_L g178 ( 
.A1(n_147),
.A2(n_124),
.B(n_103),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_99),
.B(n_86),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_148),
.B(n_151),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_123),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_119),
.B(n_67),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_122),
.A2(n_56),
.B1(n_60),
.B2(n_77),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_107),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_153),
.B(n_154),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_119),
.B(n_38),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_128),
.B(n_80),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_156),
.B(n_108),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_139),
.A2(n_136),
.B1(n_152),
.B2(n_146),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_157),
.A2(n_176),
.B1(n_181),
.B2(n_182),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_158),
.B(n_185),
.C(n_150),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_SL g159 ( 
.A(n_131),
.B(n_110),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_159),
.B(n_170),
.Y(n_190)
);

OAI21xp5_ASAP7_75t_L g199 ( 
.A1(n_160),
.A2(n_183),
.B(n_135),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_161),
.A2(n_162),
.B1(n_173),
.B2(n_177),
.Y(n_189)
);

CKINVDCx14_ASAP7_75t_R g163 ( 
.A(n_132),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_163),
.B(n_171),
.Y(n_212)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_143),
.Y(n_170)
);

FAx1_ASAP7_75t_SL g171 ( 
.A(n_156),
.B(n_104),
.CI(n_112),
.CON(n_171),
.SN(n_171)
);

AND2x2_ASAP7_75t_L g172 ( 
.A(n_145),
.B(n_106),
.Y(n_172)
);

AOI21xp5_ASAP7_75t_L g202 ( 
.A1(n_172),
.A2(n_135),
.B(n_153),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_129),
.A2(n_138),
.B1(n_130),
.B2(n_142),
.Y(n_173)
);

INVx1_ASAP7_75t_SL g174 ( 
.A(n_149),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_174),
.B(n_155),
.Y(n_191)
);

INVxp67_ASAP7_75t_L g175 ( 
.A(n_132),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_175),
.B(n_180),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_141),
.A2(n_121),
.B1(n_63),
.B2(n_98),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_138),
.A2(n_124),
.B1(n_103),
.B2(n_118),
.Y(n_177)
);

XOR2xp5_ASAP7_75t_L g215 ( 
.A(n_178),
.B(n_22),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_SL g180 ( 
.A(n_151),
.B(n_27),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_140),
.B(n_154),
.Y(n_184)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_184),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_147),
.B(n_42),
.C(n_41),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_148),
.B(n_80),
.Y(n_186)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_186),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_133),
.A2(n_102),
.B1(n_93),
.B2(n_32),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_L g203 ( 
.A1(n_187),
.A2(n_155),
.B1(n_134),
.B2(n_149),
.Y(n_203)
);

AOI21xp5_ASAP7_75t_SL g188 ( 
.A1(n_160),
.A2(n_144),
.B(n_147),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_L g227 ( 
.A1(n_188),
.A2(n_199),
.B(n_202),
.Y(n_227)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_191),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_179),
.B(n_137),
.Y(n_192)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_192),
.Y(n_228)
);

INVx3_ASAP7_75t_L g194 ( 
.A(n_174),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_194),
.B(n_203),
.Y(n_245)
);

BUFx12f_ASAP7_75t_L g195 ( 
.A(n_179),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_195),
.Y(n_225)
);

CKINVDCx14_ASAP7_75t_R g196 ( 
.A(n_186),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g221 ( 
.A(n_196),
.B(n_200),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_197),
.B(n_205),
.Y(n_226)
);

INVxp67_ASAP7_75t_L g200 ( 
.A(n_183),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_173),
.A2(n_134),
.B1(n_155),
.B2(n_105),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_204),
.A2(n_208),
.B1(n_216),
.B2(n_187),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_167),
.B(n_41),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_185),
.B(n_41),
.C(n_42),
.Y(n_206)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_206),
.B(n_211),
.Y(n_238)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_168),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_207),
.B(n_209),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_157),
.A2(n_182),
.B1(n_176),
.B2(n_164),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_168),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_177),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_210),
.B(n_218),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_167),
.B(n_28),
.C(n_31),
.Y(n_211)
);

AO22x1_ASAP7_75t_L g214 ( 
.A1(n_162),
.A2(n_22),
.B1(n_23),
.B2(n_2),
.Y(n_214)
);

OAI21xp5_ASAP7_75t_L g233 ( 
.A1(n_214),
.A2(n_164),
.B(n_180),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_215),
.B(n_158),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_161),
.A2(n_32),
.B1(n_31),
.B2(n_27),
.Y(n_216)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_175),
.Y(n_217)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_217),
.Y(n_232)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_169),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_169),
.Y(n_219)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_219),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_220),
.B(n_231),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_197),
.B(n_184),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_222),
.B(n_230),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_229),
.A2(n_240),
.B1(n_242),
.B2(n_214),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_199),
.B(n_178),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_212),
.B(n_205),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_SL g251 ( 
.A(n_233),
.B(n_216),
.Y(n_251)
);

OAI21xp5_ASAP7_75t_L g234 ( 
.A1(n_188),
.A2(n_193),
.B(n_200),
.Y(n_234)
);

OAI21xp5_ASAP7_75t_SL g264 ( 
.A1(n_234),
.A2(n_229),
.B(n_227),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_189),
.B(n_172),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_236),
.B(n_237),
.C(n_215),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g237 ( 
.A(n_202),
.B(n_172),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_195),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_239),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_208),
.A2(n_166),
.B1(n_170),
.B2(n_165),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_195),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_241),
.B(n_244),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_198),
.A2(n_171),
.B1(n_159),
.B2(n_181),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_213),
.Y(n_244)
);

XOR2xp5_ASAP7_75t_L g268 ( 
.A(n_246),
.B(n_255),
.Y(n_268)
);

CKINVDCx16_ASAP7_75t_R g247 ( 
.A(n_245),
.Y(n_247)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_247),
.Y(n_270)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_251),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_SL g273 ( 
.A(n_252),
.B(n_236),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_228),
.B(n_190),
.Y(n_253)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_253),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_226),
.B(n_201),
.C(n_206),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_254),
.B(n_226),
.C(n_238),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_SL g255 ( 
.A(n_242),
.B(n_204),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_243),
.A2(n_198),
.B1(n_217),
.B2(n_194),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_256),
.A2(n_223),
.B1(n_222),
.B2(n_225),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_240),
.A2(n_171),
.B1(n_211),
.B2(n_26),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_257),
.A2(n_261),
.B1(n_266),
.B2(n_13),
.Y(n_283)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_221),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_258),
.B(n_260),
.Y(n_269)
);

OR2x2_ASAP7_75t_L g260 ( 
.A(n_243),
.B(n_26),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_235),
.A2(n_23),
.B1(n_10),
.B2(n_16),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_224),
.Y(n_262)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_262),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_SL g263 ( 
.A(n_238),
.B(n_10),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_263),
.Y(n_282)
);

AOI21xp5_ASAP7_75t_L g274 ( 
.A1(n_264),
.A2(n_233),
.B(n_232),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_SL g265 ( 
.A(n_227),
.B(n_22),
.Y(n_265)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_265),
.B(n_25),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_234),
.A2(n_23),
.B1(n_8),
.B2(n_14),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_L g267 ( 
.A1(n_264),
.A2(n_252),
.B1(n_266),
.B2(n_249),
.Y(n_267)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_267),
.Y(n_285)
);

AOI21x1_ASAP7_75t_SL g272 ( 
.A1(n_256),
.A2(n_230),
.B(n_237),
.Y(n_272)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_272),
.Y(n_294)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_273),
.Y(n_296)
);

AOI21xp5_ASAP7_75t_L g291 ( 
.A1(n_274),
.A2(n_246),
.B(n_261),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_275),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_276),
.B(n_277),
.C(n_250),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_254),
.B(n_220),
.C(n_231),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_L g278 ( 
.A1(n_257),
.A2(n_13),
.B1(n_12),
.B2(n_11),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_278),
.A2(n_11),
.B1(n_10),
.B2(n_3),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_SL g299 ( 
.A(n_279),
.B(n_0),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_259),
.B(n_13),
.Y(n_280)
);

XOR2xp5_ASAP7_75t_L g289 ( 
.A(n_280),
.B(n_259),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_SL g297 ( 
.A(n_283),
.B(n_12),
.Y(n_297)
);

A2O1A1Ixp33_ASAP7_75t_SL g286 ( 
.A1(n_272),
.A2(n_255),
.B(n_265),
.C(n_248),
.Y(n_286)
);

AOI22xp33_ASAP7_75t_SL g300 ( 
.A1(n_286),
.A2(n_288),
.B1(n_284),
.B2(n_281),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_270),
.B(n_269),
.Y(n_287)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_287),
.Y(n_303)
);

INVx3_ASAP7_75t_L g288 ( 
.A(n_271),
.Y(n_288)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_289),
.Y(n_306)
);

OA21x2_ASAP7_75t_SL g290 ( 
.A1(n_280),
.A2(n_250),
.B(n_260),
.Y(n_290)
);

NOR2xp67_ASAP7_75t_L g311 ( 
.A(n_290),
.B(n_268),
.Y(n_311)
);

AOI21xp5_ASAP7_75t_L g305 ( 
.A1(n_291),
.A2(n_269),
.B(n_273),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_292),
.B(n_276),
.C(n_277),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_SL g308 ( 
.A(n_293),
.B(n_298),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_SL g295 ( 
.A1(n_274),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_SL g307 ( 
.A1(n_295),
.A2(n_275),
.B1(n_282),
.B2(n_5),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_297),
.B(n_283),
.Y(n_304)
);

XOR2xp5_ASAP7_75t_L g301 ( 
.A(n_299),
.B(n_279),
.Y(n_301)
);

AOI21xp5_ASAP7_75t_L g316 ( 
.A1(n_300),
.A2(n_305),
.B(n_311),
.Y(n_316)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_301),
.Y(n_312)
);

HB1xp67_ASAP7_75t_L g302 ( 
.A(n_286),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_302),
.B(n_304),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_307),
.B(n_309),
.Y(n_314)
);

OAI22xp5_ASAP7_75t_SL g309 ( 
.A1(n_294),
.A2(n_285),
.B1(n_296),
.B2(n_286),
.Y(n_309)
);

OAI21xp5_ASAP7_75t_L g318 ( 
.A1(n_310),
.A2(n_292),
.B(n_286),
.Y(n_318)
);

XNOR2xp5_ASAP7_75t_L g315 ( 
.A(n_310),
.B(n_289),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_315),
.B(n_319),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_307),
.B(n_298),
.Y(n_317)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_317),
.Y(n_324)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_318),
.Y(n_327)
);

XNOR2xp5_ASAP7_75t_L g319 ( 
.A(n_305),
.B(n_268),
.Y(n_319)
);

AOI22xp5_ASAP7_75t_SL g320 ( 
.A1(n_303),
.A2(n_288),
.B1(n_295),
.B2(n_299),
.Y(n_320)
);

A2O1A1Ixp33_ASAP7_75t_SL g326 ( 
.A1(n_320),
.A2(n_301),
.B(n_4),
.C(n_5),
.Y(n_326)
);

OAI21x1_ASAP7_75t_L g322 ( 
.A1(n_319),
.A2(n_309),
.B(n_306),
.Y(n_322)
);

OAI21x1_ASAP7_75t_L g328 ( 
.A1(n_322),
.A2(n_325),
.B(n_316),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_320),
.B(n_308),
.Y(n_323)
);

OAI22xp5_ASAP7_75t_L g331 ( 
.A1(n_323),
.A2(n_326),
.B1(n_4),
.B2(n_5),
.Y(n_331)
);

INVxp33_ASAP7_75t_L g325 ( 
.A(n_313),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_328),
.B(n_330),
.Y(n_332)
);

NOR3xp33_ASAP7_75t_L g329 ( 
.A(n_327),
.B(n_312),
.C(n_314),
.Y(n_329)
);

AOI21xp33_ASAP7_75t_L g333 ( 
.A1(n_329),
.A2(n_331),
.B(n_324),
.Y(n_333)
);

OAI21xp5_ASAP7_75t_L g330 ( 
.A1(n_321),
.A2(n_1),
.B(n_4),
.Y(n_330)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_333),
.Y(n_334)
);

NAND2xp33_ASAP7_75t_SL g335 ( 
.A(n_334),
.B(n_332),
.Y(n_335)
);

AOI22xp33_ASAP7_75t_L g336 ( 
.A1(n_335),
.A2(n_326),
.B1(n_6),
.B2(n_7),
.Y(n_336)
);

OAI21xp5_ASAP7_75t_L g337 ( 
.A1(n_336),
.A2(n_6),
.B(n_7),
.Y(n_337)
);

OAI21xp5_ASAP7_75t_SL g338 ( 
.A1(n_337),
.A2(n_6),
.B(n_7),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_338),
.B(n_6),
.Y(n_339)
);


endmodule