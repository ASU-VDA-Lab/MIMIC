module fake_jpeg_1297_n_206 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_206);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_206;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_143;
wire n_202;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_0),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_9),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_29),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_13),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_27),
.Y(n_52)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_21),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_34),
.B(n_14),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_20),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_26),
.Y(n_56)
);

BUFx16f_ASAP7_75t_L g57 ( 
.A(n_3),
.Y(n_57)
);

INVx5_ASAP7_75t_L g58 ( 
.A(n_5),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_38),
.Y(n_59)
);

BUFx5_ASAP7_75t_L g60 ( 
.A(n_14),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_35),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_2),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_45),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_46),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_10),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_43),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_13),
.Y(n_67)
);

INVx1_ASAP7_75t_SL g68 ( 
.A(n_23),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_19),
.Y(n_69)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_1),
.Y(n_70)
);

INVx5_ASAP7_75t_L g71 ( 
.A(n_57),
.Y(n_71)
);

INVx1_ASAP7_75t_SL g91 ( 
.A(n_71),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_47),
.B(n_48),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_72),
.B(n_59),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_63),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_73),
.Y(n_84)
);

BUFx3_ASAP7_75t_L g74 ( 
.A(n_57),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_74),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_63),
.Y(n_75)
);

INVx6_ASAP7_75t_L g81 ( 
.A(n_75),
.Y(n_81)
);

INVx5_ASAP7_75t_L g76 ( 
.A(n_53),
.Y(n_76)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_76),
.Y(n_79)
);

BUFx5_ASAP7_75t_L g77 ( 
.A(n_57),
.Y(n_77)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_77),
.Y(n_83)
);

INVx6_ASAP7_75t_L g78 ( 
.A(n_67),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_78),
.Y(n_82)
);

O2A1O1Ixp33_ASAP7_75t_SL g80 ( 
.A1(n_76),
.A2(n_78),
.B(n_74),
.C(n_53),
.Y(n_80)
);

AOI21xp5_ASAP7_75t_L g102 ( 
.A1(n_80),
.A2(n_86),
.B(n_91),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_73),
.B(n_54),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_85),
.B(n_89),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_75),
.A2(n_67),
.B1(n_49),
.B2(n_58),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_L g87 ( 
.A1(n_73),
.A2(n_58),
.B1(n_69),
.B2(n_51),
.Y(n_87)
);

OAI22xp33_ASAP7_75t_L g111 ( 
.A1(n_87),
.A2(n_56),
.B1(n_68),
.B2(n_66),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_78),
.B(n_55),
.Y(n_88)
);

NOR2x1_ASAP7_75t_L g109 ( 
.A(n_88),
.B(n_70),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_72),
.B(n_62),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_92),
.B(n_61),
.Y(n_95)
);

INVx8_ASAP7_75t_L g94 ( 
.A(n_90),
.Y(n_94)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_94),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_95),
.B(n_109),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_90),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_96),
.B(n_100),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_84),
.Y(n_97)
);

CKINVDCx14_ASAP7_75t_R g116 ( 
.A(n_97),
.Y(n_116)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_79),
.Y(n_98)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_98),
.Y(n_112)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_81),
.Y(n_99)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_99),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_88),
.B(n_64),
.Y(n_100)
);

OR2x4_ASAP7_75t_L g101 ( 
.A(n_80),
.B(n_53),
.Y(n_101)
);

AO21x1_ASAP7_75t_L g119 ( 
.A1(n_101),
.A2(n_110),
.B(n_83),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_102),
.A2(n_24),
.B1(n_42),
.B2(n_41),
.Y(n_129)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_79),
.Y(n_103)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_103),
.Y(n_128)
);

INVx6_ASAP7_75t_L g104 ( 
.A(n_84),
.Y(n_104)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_104),
.Y(n_130)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_91),
.Y(n_105)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_105),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_83),
.B(n_64),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_106),
.B(n_107),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_81),
.Y(n_107)
);

INVx5_ASAP7_75t_L g108 ( 
.A(n_80),
.Y(n_108)
);

AND2x2_ASAP7_75t_L g118 ( 
.A(n_108),
.B(n_111),
.Y(n_118)
);

AOI21xp5_ASAP7_75t_L g110 ( 
.A1(n_86),
.A2(n_68),
.B(n_65),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_109),
.B(n_82),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_114),
.B(n_115),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_93),
.B(n_108),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_101),
.A2(n_82),
.B1(n_49),
.B2(n_70),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_117),
.A2(n_120),
.B1(n_129),
.B2(n_44),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_SL g143 ( 
.A1(n_119),
.A2(n_127),
.B(n_118),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_111),
.A2(n_66),
.B1(n_55),
.B2(n_52),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_99),
.B(n_50),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_122),
.B(n_123),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_107),
.B(n_50),
.Y(n_123)
);

OAI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_97),
.A2(n_52),
.B1(n_60),
.B2(n_22),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_L g153 ( 
.A1(n_124),
.A2(n_36),
.B1(n_33),
.B2(n_32),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_SL g127 ( 
.A1(n_94),
.A2(n_60),
.B1(n_1),
.B2(n_2),
.Y(n_127)
);

XOR2xp5_ASAP7_75t_L g133 ( 
.A(n_115),
.B(n_104),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_133),
.B(n_28),
.C(n_30),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_121),
.B(n_0),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_135),
.B(n_136),
.Y(n_158)
);

INVx4_ASAP7_75t_L g137 ( 
.A(n_125),
.Y(n_137)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_137),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g138 ( 
.A(n_130),
.Y(n_138)
);

INVxp67_ASAP7_75t_L g172 ( 
.A(n_138),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_114),
.A2(n_118),
.B1(n_119),
.B2(n_132),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_140),
.B(n_156),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_126),
.B(n_40),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_141),
.B(n_144),
.Y(n_167)
);

INVx13_ASAP7_75t_L g142 ( 
.A(n_116),
.Y(n_142)
);

INVx1_ASAP7_75t_SL g157 ( 
.A(n_142),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_SL g169 ( 
.A1(n_143),
.A2(n_149),
.B(n_150),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_122),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_123),
.B(n_39),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_145),
.B(n_146),
.Y(n_170)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_112),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_120),
.B(n_3),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_147),
.B(n_148),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_128),
.B(n_4),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_L g149 ( 
.A1(n_118),
.A2(n_4),
.B(n_5),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_L g150 ( 
.A1(n_117),
.A2(n_6),
.B(n_7),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_113),
.Y(n_151)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_151),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_131),
.B(n_6),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_152),
.B(n_153),
.Y(n_168)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_125),
.Y(n_154)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_154),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_SL g155 ( 
.A(n_132),
.B(n_7),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_155),
.B(n_17),
.Y(n_174)
);

OAI32xp33_ASAP7_75t_L g156 ( 
.A1(n_115),
.A2(n_8),
.A3(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_134),
.A2(n_8),
.B1(n_11),
.B2(n_12),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_160),
.B(n_161),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_140),
.A2(n_12),
.B1(n_15),
.B2(n_16),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_138),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_162),
.B(n_175),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g180 ( 
.A(n_163),
.B(n_156),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_133),
.A2(n_15),
.B1(n_16),
.B2(n_17),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_173),
.B(n_160),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_174),
.B(n_31),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_141),
.B(n_18),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_167),
.B(n_139),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_176),
.B(n_178),
.C(n_180),
.Y(n_189)
);

AOI21xp5_ASAP7_75t_L g177 ( 
.A1(n_169),
.A2(n_143),
.B(n_149),
.Y(n_177)
);

AOI21xp5_ASAP7_75t_L g192 ( 
.A1(n_177),
.A2(n_173),
.B(n_150),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_L g178 ( 
.A(n_170),
.B(n_145),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_179),
.B(n_182),
.Y(n_188)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_164),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_165),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_183),
.A2(n_185),
.B1(n_168),
.B2(n_171),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_L g186 ( 
.A1(n_176),
.A2(n_166),
.B1(n_158),
.B2(n_136),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_186),
.B(n_187),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_180),
.B(n_163),
.C(n_166),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_190),
.B(n_191),
.C(n_181),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_184),
.B(n_169),
.C(n_161),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_192),
.B(n_157),
.C(n_172),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_193),
.B(n_189),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_188),
.B(n_172),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_194),
.B(n_196),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_195),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_197),
.B(n_198),
.C(n_157),
.Y(n_201)
);

XOR2xp5_ASAP7_75t_L g200 ( 
.A(n_199),
.B(n_186),
.Y(n_200)
);

OAI21xp33_ASAP7_75t_L g202 ( 
.A1(n_200),
.A2(n_201),
.B(n_159),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_202),
.B(n_159),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_203),
.B(n_142),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_204),
.B(n_137),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_205),
.B(n_25),
.Y(n_206)
);


endmodule