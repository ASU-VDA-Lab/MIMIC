module fake_jpeg_4534_n_333 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_333);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_333;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_3),
.Y(n_16)
);

INVx6_ASAP7_75t_SL g17 ( 
.A(n_7),
.Y(n_17)
);

BUFx16f_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_3),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_15),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

BUFx4f_ASAP7_75t_L g25 ( 
.A(n_15),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

BUFx2_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_0),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_9),
.Y(n_33)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_25),
.Y(n_34)
);

INVx8_ASAP7_75t_L g65 ( 
.A(n_34),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_20),
.B(n_0),
.Y(n_35)
);

AND2x2_ASAP7_75t_L g49 ( 
.A(n_35),
.B(n_36),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_20),
.B(n_0),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_27),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_37),
.B(n_38),
.Y(n_53)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_27),
.Y(n_38)
);

INVx11_ASAP7_75t_L g39 ( 
.A(n_19),
.Y(n_39)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_39),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_18),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_40),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_27),
.B(n_15),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_SL g58 ( 
.A(n_41),
.B(n_42),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_27),
.B(n_14),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_18),
.Y(n_43)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_43),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_18),
.Y(n_44)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_44),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_34),
.A2(n_30),
.B1(n_17),
.B2(n_33),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_45),
.A2(n_68),
.B1(n_60),
.B2(n_26),
.Y(n_86)
);

BUFx16f_ASAP7_75t_L g46 ( 
.A(n_40),
.Y(n_46)
);

CKINVDCx16_ASAP7_75t_R g97 ( 
.A(n_46),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_35),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_47),
.B(n_54),
.Y(n_77)
);

NAND2x1_ASAP7_75t_SL g48 ( 
.A(n_41),
.B(n_17),
.Y(n_48)
);

NAND2xp33_ASAP7_75t_SL g95 ( 
.A(n_48),
.B(n_18),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_39),
.Y(n_50)
);

INVx8_ASAP7_75t_L g73 ( 
.A(n_50),
.Y(n_73)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_40),
.Y(n_52)
);

INVxp67_ASAP7_75t_L g83 ( 
.A(n_52),
.Y(n_83)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_37),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_35),
.B(n_22),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_55),
.B(n_57),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_36),
.B(n_22),
.Y(n_57)
);

CKINVDCx16_ASAP7_75t_R g59 ( 
.A(n_41),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_59),
.B(n_62),
.Y(n_81)
);

AO22x1_ASAP7_75t_SL g60 ( 
.A1(n_34),
.A2(n_17),
.B1(n_26),
.B2(n_18),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_60),
.A2(n_70),
.B1(n_22),
.B2(n_32),
.Y(n_88)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_37),
.Y(n_61)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_61),
.Y(n_78)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_37),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_40),
.B(n_33),
.Y(n_63)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_63),
.Y(n_89)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_36),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_64),
.B(n_71),
.Y(n_91)
);

INVx5_ASAP7_75t_L g66 ( 
.A(n_38),
.Y(n_66)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_66),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_34),
.A2(n_30),
.B1(n_23),
.B2(n_33),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_39),
.A2(n_30),
.B1(n_31),
.B2(n_16),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_SL g71 ( 
.A(n_42),
.B(n_23),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_42),
.B(n_32),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_72),
.B(n_49),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_75),
.B(n_79),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g76 ( 
.A(n_64),
.B(n_34),
.C(n_38),
.Y(n_76)
);

OAI21xp5_ASAP7_75t_SL g105 ( 
.A1(n_76),
.A2(n_95),
.B(n_53),
.Y(n_105)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_66),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_L g82 ( 
.A1(n_47),
.A2(n_30),
.B1(n_39),
.B2(n_38),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_82),
.A2(n_96),
.B1(n_51),
.B2(n_56),
.Y(n_109)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_46),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_84),
.B(n_85),
.Y(n_118)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_46),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_86),
.A2(n_48),
.B1(n_65),
.B2(n_28),
.Y(n_99)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_60),
.Y(n_87)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_87),
.Y(n_103)
);

CKINVDCx16_ASAP7_75t_R g98 ( 
.A(n_88),
.Y(n_98)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_67),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_90),
.Y(n_108)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_55),
.Y(n_92)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_92),
.Y(n_101)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_67),
.Y(n_93)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_93),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_49),
.B(n_20),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_94),
.B(n_57),
.Y(n_100)
);

AO22x1_ASAP7_75t_SL g96 ( 
.A1(n_49),
.A2(n_39),
.B1(n_25),
.B2(n_26),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_99),
.A2(n_107),
.B1(n_113),
.B2(n_56),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_SL g126 ( 
.A(n_100),
.B(n_89),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_74),
.B(n_72),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_102),
.B(n_110),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_L g104 ( 
.A1(n_94),
.A2(n_48),
.B(n_58),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_104),
.B(n_28),
.C(n_29),
.Y(n_136)
);

AND2x2_ASAP7_75t_L g141 ( 
.A(n_105),
.B(n_122),
.Y(n_141)
);

CKINVDCx16_ASAP7_75t_R g106 ( 
.A(n_81),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_106),
.B(n_112),
.Y(n_127)
);

OAI22x1_ASAP7_75t_SL g107 ( 
.A1(n_96),
.A2(n_65),
.B1(n_54),
.B2(n_62),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_109),
.A2(n_114),
.B1(n_124),
.B2(n_69),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_74),
.B(n_58),
.Y(n_110)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_77),
.Y(n_112)
);

OA22x2_ASAP7_75t_L g113 ( 
.A1(n_96),
.A2(n_61),
.B1(n_70),
.B2(n_51),
.Y(n_113)
);

O2A1O1Ixp33_ASAP7_75t_SL g114 ( 
.A1(n_88),
.A2(n_71),
.B(n_25),
.C(n_21),
.Y(n_114)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_81),
.Y(n_116)
);

CKINVDCx14_ASAP7_75t_R g143 ( 
.A(n_116),
.Y(n_143)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_77),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_117),
.B(n_120),
.Y(n_130)
);

AOI32xp33_ASAP7_75t_L g119 ( 
.A1(n_96),
.A2(n_44),
.A3(n_40),
.B1(n_43),
.B2(n_25),
.Y(n_119)
);

A2O1A1Ixp33_ASAP7_75t_L g128 ( 
.A1(n_119),
.A2(n_93),
.B(n_25),
.C(n_83),
.Y(n_128)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_91),
.Y(n_120)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_79),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_121),
.B(n_123),
.Y(n_145)
);

OR2x2_ASAP7_75t_L g122 ( 
.A(n_95),
.B(n_16),
.Y(n_122)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_91),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_87),
.A2(n_92),
.B1(n_75),
.B2(n_76),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_126),
.B(n_147),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_128),
.A2(n_134),
.B1(n_142),
.B2(n_113),
.Y(n_161)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_114),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_129),
.B(n_133),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_110),
.B(n_89),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_131),
.B(n_137),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_132),
.A2(n_146),
.B1(n_109),
.B2(n_107),
.Y(n_154)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_114),
.Y(n_133)
);

INVx4_ASAP7_75t_L g135 ( 
.A(n_107),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_135),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_L g164 ( 
.A(n_136),
.B(n_104),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_102),
.B(n_78),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_100),
.B(n_78),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_L g158 ( 
.A1(n_138),
.A2(n_139),
.B(n_144),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_101),
.B(n_29),
.Y(n_139)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_121),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_140),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_98),
.A2(n_69),
.B1(n_73),
.B2(n_25),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_101),
.B(n_32),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_98),
.A2(n_80),
.B1(n_90),
.B2(n_73),
.Y(n_146)
);

CKINVDCx14_ASAP7_75t_R g147 ( 
.A(n_118),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_120),
.B(n_80),
.Y(n_148)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_148),
.Y(n_157)
);

BUFx12_ASAP7_75t_L g149 ( 
.A(n_118),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_149),
.Y(n_177)
);

CKINVDCx14_ASAP7_75t_R g150 ( 
.A(n_111),
.Y(n_150)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_150),
.Y(n_160)
);

CKINVDCx16_ASAP7_75t_R g151 ( 
.A(n_111),
.Y(n_151)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_151),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_123),
.B(n_16),
.Y(n_152)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_152),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g207 ( 
.A1(n_154),
.A2(n_179),
.B1(n_149),
.B2(n_115),
.Y(n_207)
);

OR2x2_ASAP7_75t_L g155 ( 
.A(n_151),
.B(n_113),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_155),
.B(n_162),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_132),
.A2(n_129),
.B1(n_133),
.B2(n_103),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_156),
.A2(n_165),
.B1(n_169),
.B2(n_173),
.Y(n_201)
);

AND2x6_ASAP7_75t_L g159 ( 
.A(n_141),
.B(n_113),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_159),
.B(n_142),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_161),
.A2(n_152),
.B1(n_149),
.B2(n_73),
.Y(n_206)
);

BUFx6f_ASAP7_75t_L g162 ( 
.A(n_140),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_164),
.B(n_166),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_134),
.A2(n_103),
.B1(n_113),
.B2(n_114),
.Y(n_165)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_149),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g167 ( 
.A(n_125),
.B(n_124),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_167),
.B(n_174),
.C(n_126),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_141),
.A2(n_103),
.B1(n_146),
.B2(n_135),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_137),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_170),
.B(n_171),
.Y(n_200)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_145),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_L g172 ( 
.A1(n_141),
.A2(n_125),
.B(n_105),
.Y(n_172)
);

AOI21xp5_ASAP7_75t_L g188 ( 
.A1(n_172),
.A2(n_128),
.B(n_136),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_135),
.A2(n_119),
.B1(n_104),
.B2(n_117),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_138),
.B(n_112),
.C(n_106),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_128),
.A2(n_99),
.B1(n_122),
.B2(n_108),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_SL g181 ( 
.A1(n_168),
.A2(n_127),
.B(n_131),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_L g227 ( 
.A1(n_181),
.A2(n_188),
.B(n_190),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_176),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_182),
.B(n_191),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_183),
.B(n_185),
.Y(n_208)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_175),
.Y(n_185)
);

BUFx6f_ASAP7_75t_L g186 ( 
.A(n_162),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_186),
.B(n_189),
.Y(n_211)
);

BUFx5_ASAP7_75t_L g187 ( 
.A(n_159),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_187),
.Y(n_216)
);

AOI21xp5_ASAP7_75t_L g190 ( 
.A1(n_172),
.A2(n_127),
.B(n_130),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_175),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_L g192 ( 
.A(n_167),
.B(n_130),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_SL g213 ( 
.A(n_192),
.B(n_205),
.Y(n_213)
);

INVxp67_ASAP7_75t_L g193 ( 
.A(n_169),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_193),
.B(n_196),
.Y(n_209)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_178),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_194),
.B(n_195),
.Y(n_215)
);

OAI21xp5_ASAP7_75t_SL g195 ( 
.A1(n_153),
.A2(n_145),
.B(n_122),
.Y(n_195)
);

INVxp67_ASAP7_75t_L g196 ( 
.A(n_156),
.Y(n_196)
);

NOR2xp67_ASAP7_75t_L g197 ( 
.A(n_173),
.B(n_143),
.Y(n_197)
);

NOR4xp25_ASAP7_75t_L g221 ( 
.A(n_197),
.B(n_158),
.C(n_160),
.D(n_180),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_177),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_198),
.Y(n_220)
);

INVx2_ASAP7_75t_SL g202 ( 
.A(n_166),
.Y(n_202)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_202),
.Y(n_210)
);

INVxp67_ASAP7_75t_L g203 ( 
.A(n_165),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_203),
.B(n_163),
.Y(n_233)
);

OAI21xp5_ASAP7_75t_L g204 ( 
.A1(n_179),
.A2(n_139),
.B(n_144),
.Y(n_204)
);

AO21x1_ASAP7_75t_L g231 ( 
.A1(n_204),
.A2(n_163),
.B(n_23),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_164),
.B(n_148),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_L g212 ( 
.A1(n_206),
.A2(n_193),
.B1(n_203),
.B2(n_196),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_207),
.A2(n_161),
.B1(n_174),
.B2(n_158),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_212),
.A2(n_214),
.B1(n_97),
.B2(n_21),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_L g214 ( 
.A1(n_187),
.A2(n_155),
.B1(n_154),
.B2(n_170),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_202),
.B(n_171),
.Y(n_217)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_217),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_218),
.A2(n_219),
.B1(n_221),
.B2(n_226),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_201),
.A2(n_184),
.B1(n_183),
.B2(n_204),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_200),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_222),
.B(n_223),
.Y(n_234)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_206),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_199),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_224),
.B(n_228),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_202),
.B(n_186),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_225),
.B(n_232),
.Y(n_235)
);

OA22x2_ASAP7_75t_L g226 ( 
.A1(n_201),
.A2(n_180),
.B1(n_160),
.B2(n_157),
.Y(n_226)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_190),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_189),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_229),
.B(n_228),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_231),
.A2(n_28),
.B1(n_29),
.B2(n_31),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_194),
.B(n_108),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_L g250 ( 
.A1(n_233),
.A2(n_21),
.B1(n_31),
.B2(n_84),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_213),
.B(n_192),
.Y(n_236)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_236),
.B(n_239),
.Y(n_273)
);

HB1xp67_ASAP7_75t_L g237 ( 
.A(n_226),
.Y(n_237)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_237),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_229),
.B(n_188),
.C(n_185),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_238),
.B(n_241),
.C(n_243),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_SL g239 ( 
.A(n_219),
.B(n_205),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_213),
.B(n_224),
.C(n_211),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_208),
.B(n_195),
.Y(n_243)
);

OAI21xp5_ASAP7_75t_SL g259 ( 
.A1(n_245),
.A2(n_255),
.B(n_230),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_214),
.B(n_181),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_246),
.B(n_253),
.Y(n_262)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_227),
.B(n_52),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_247),
.B(n_251),
.C(n_252),
.Y(n_258)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_248),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_SL g249 ( 
.A(n_220),
.B(n_85),
.Y(n_249)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_249),
.Y(n_261)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_250),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_216),
.B(n_97),
.C(n_44),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g252 ( 
.A(n_227),
.B(n_52),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_216),
.B(n_44),
.C(n_43),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_254),
.B(n_209),
.C(n_210),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_SL g255 ( 
.A(n_220),
.B(n_11),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_259),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_263),
.B(n_265),
.C(n_268),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_244),
.A2(n_212),
.B1(n_223),
.B2(n_209),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_L g277 ( 
.A1(n_264),
.A2(n_266),
.B1(n_234),
.B2(n_240),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_241),
.B(n_218),
.C(n_215),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_254),
.A2(n_226),
.B1(n_233),
.B2(n_222),
.Y(n_266)
);

OAI21xp5_ASAP7_75t_SL g267 ( 
.A1(n_251),
.A2(n_226),
.B(n_210),
.Y(n_267)
);

OAI21xp5_ASAP7_75t_SL g280 ( 
.A1(n_267),
.A2(n_247),
.B(n_19),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_238),
.B(n_221),
.C(n_231),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_235),
.B(n_231),
.Y(n_270)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_270),
.Y(n_276)
);

XNOR2x1_ASAP7_75t_L g271 ( 
.A(n_239),
.B(n_246),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g287 ( 
.A(n_271),
.B(n_274),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_242),
.B(n_67),
.C(n_52),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_272),
.B(n_24),
.C(n_19),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_236),
.B(n_252),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_263),
.Y(n_275)
);

OAI21xp5_ASAP7_75t_SL g302 ( 
.A1(n_275),
.A2(n_280),
.B(n_281),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_277),
.B(n_279),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_271),
.B(n_243),
.Y(n_279)
);

OR2x2_ASAP7_75t_L g281 ( 
.A(n_256),
.B(n_0),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_261),
.B(n_24),
.Y(n_282)
);

AOI21xp5_ASAP7_75t_L g292 ( 
.A1(n_282),
.A2(n_288),
.B(n_257),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_272),
.B(n_50),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_SL g293 ( 
.A(n_283),
.B(n_284),
.Y(n_293)
);

NOR5xp2_ASAP7_75t_L g284 ( 
.A(n_262),
.B(n_10),
.C(n_14),
.D(n_13),
.E(n_12),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_SL g294 ( 
.A(n_285),
.B(n_257),
.Y(n_294)
);

OAI21xp5_ASAP7_75t_L g288 ( 
.A1(n_268),
.A2(n_265),
.B(n_258),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_260),
.B(n_19),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_SL g295 ( 
.A(n_289),
.B(n_290),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_258),
.A2(n_24),
.B1(n_2),
.B2(n_3),
.Y(n_290)
);

OAI21xp5_ASAP7_75t_L g311 ( 
.A1(n_292),
.A2(n_298),
.B(n_299),
.Y(n_311)
);

AOI21xp5_ASAP7_75t_L g310 ( 
.A1(n_294),
.A2(n_296),
.B(n_297),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_282),
.B(n_269),
.Y(n_296)
);

AO221x1_ASAP7_75t_L g297 ( 
.A1(n_275),
.A2(n_273),
.B1(n_44),
.B2(n_43),
.C(n_24),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_276),
.B(n_273),
.Y(n_298)
);

OAI21xp5_ASAP7_75t_L g299 ( 
.A1(n_280),
.A2(n_1),
.B(n_2),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_290),
.B(n_24),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_300),
.B(n_301),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_286),
.B(n_24),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_285),
.B(n_24),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_303),
.B(n_288),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_L g304 ( 
.A1(n_278),
.A2(n_14),
.B1(n_13),
.B2(n_12),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_L g313 ( 
.A1(n_304),
.A2(n_2),
.B1(n_4),
.B2(n_5),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_SL g319 ( 
.A(n_306),
.B(n_308),
.Y(n_319)
);

AOI322xp5_ASAP7_75t_L g307 ( 
.A1(n_293),
.A2(n_278),
.A3(n_279),
.B1(n_281),
.B2(n_287),
.C1(n_9),
.C2(n_13),
.Y(n_307)
);

OAI21x1_ASAP7_75t_L g321 ( 
.A1(n_307),
.A2(n_314),
.B(n_5),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_300),
.B(n_287),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_291),
.B(n_11),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_309),
.B(n_302),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_295),
.B(n_1),
.Y(n_312)
);

OAI21xp5_ASAP7_75t_L g317 ( 
.A1(n_312),
.A2(n_313),
.B(n_298),
.Y(n_317)
);

AOI322xp5_ASAP7_75t_L g314 ( 
.A1(n_299),
.A2(n_2),
.A3(n_4),
.B1(n_5),
.B2(n_6),
.C1(n_7),
.C2(n_8),
.Y(n_314)
);

AO21x1_ASAP7_75t_L g315 ( 
.A1(n_311),
.A2(n_292),
.B(n_302),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_315),
.B(n_317),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_SL g323 ( 
.A(n_316),
.B(n_318),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_313),
.B(n_43),
.Y(n_318)
);

XNOR2xp5_ASAP7_75t_L g320 ( 
.A(n_310),
.B(n_4),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_320),
.B(n_322),
.Y(n_327)
);

AO21x1_ASAP7_75t_L g324 ( 
.A1(n_321),
.A2(n_305),
.B(n_7),
.Y(n_324)
);

XNOR2xp5_ASAP7_75t_L g322 ( 
.A(n_311),
.B(n_8),
.Y(n_322)
);

OAI21xp5_ASAP7_75t_L g330 ( 
.A1(n_324),
.A2(n_326),
.B(n_6),
.Y(n_330)
);

AOI21xp5_ASAP7_75t_SL g325 ( 
.A1(n_319),
.A2(n_6),
.B(n_7),
.Y(n_325)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_325),
.Y(n_329)
);

INVxp67_ASAP7_75t_L g326 ( 
.A(n_319),
.Y(n_326)
);

O2A1O1Ixp33_ASAP7_75t_SL g331 ( 
.A1(n_330),
.A2(n_323),
.B(n_328),
.C(n_327),
.Y(n_331)
);

OAI21xp5_ASAP7_75t_SL g332 ( 
.A1(n_331),
.A2(n_329),
.B(n_8),
.Y(n_332)
);

XOR2xp5_ASAP7_75t_L g333 ( 
.A(n_332),
.B(n_8),
.Y(n_333)
);


endmodule