module fake_jpeg_21911_n_41 (n_3, n_2, n_1, n_0, n_4, n_5, n_41);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_41;

wire n_13;
wire n_21;
wire n_33;
wire n_10;
wire n_23;
wire n_27;
wire n_6;
wire n_22;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_34;
wire n_30;
wire n_39;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

INVx2_ASAP7_75t_L g6 ( 
.A(n_3),
.Y(n_6)
);

INVx2_ASAP7_75t_L g7 ( 
.A(n_2),
.Y(n_7)
);

BUFx6f_ASAP7_75t_L g8 ( 
.A(n_0),
.Y(n_8)
);

BUFx6f_ASAP7_75t_L g9 ( 
.A(n_5),
.Y(n_9)
);

NAND2xp5_ASAP7_75t_L g10 ( 
.A(n_5),
.B(n_1),
.Y(n_10)
);

INVx1_ASAP7_75t_L g11 ( 
.A(n_2),
.Y(n_11)
);

BUFx12f_ASAP7_75t_L g12 ( 
.A(n_0),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_3),
.Y(n_13)
);

MAJIxp5_ASAP7_75t_L g14 ( 
.A(n_10),
.B(n_0),
.C(n_1),
.Y(n_14)
);

OAI21xp5_ASAP7_75t_SL g27 ( 
.A1(n_14),
.A2(n_18),
.B(n_20),
.Y(n_27)
);

OAI22xp33_ASAP7_75t_SL g15 ( 
.A1(n_6),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_15)
);

AOI22xp5_ASAP7_75t_L g21 ( 
.A1(n_15),
.A2(n_20),
.B1(n_7),
.B2(n_12),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g16 ( 
.A(n_11),
.B(n_2),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_16),
.B(n_4),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_SL g17 ( 
.A(n_13),
.B(n_3),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_SL g26 ( 
.A(n_17),
.B(n_19),
.Y(n_26)
);

AOI21xp5_ASAP7_75t_L g18 ( 
.A1(n_6),
.A2(n_3),
.B(n_4),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_SL g19 ( 
.A(n_11),
.B(n_4),
.Y(n_19)
);

OAI22xp5_ASAP7_75t_SL g20 ( 
.A1(n_7),
.A2(n_4),
.B1(n_5),
.B2(n_12),
.Y(n_20)
);

OAI21xp5_ASAP7_75t_L g29 ( 
.A1(n_21),
.A2(n_22),
.B(n_25),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_SL g23 ( 
.A1(n_18),
.A2(n_12),
.B1(n_8),
.B2(n_9),
.Y(n_23)
);

MAJIxp5_ASAP7_75t_L g28 ( 
.A(n_23),
.B(n_27),
.C(n_19),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_16),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_24),
.Y(n_32)
);

A2O1A1Ixp33_ASAP7_75t_L g25 ( 
.A1(n_14),
.A2(n_12),
.B(n_8),
.C(n_9),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_L g35 ( 
.A1(n_28),
.A2(n_23),
.B1(n_26),
.B2(n_31),
.Y(n_35)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_25),
.Y(n_30)
);

MAJx2_ASAP7_75t_L g31 ( 
.A(n_27),
.B(n_17),
.C(n_24),
.Y(n_31)
);

OAI21xp5_ASAP7_75t_L g34 ( 
.A1(n_31),
.A2(n_26),
.B(n_21),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_32),
.B(n_22),
.Y(n_33)
);

MAJIxp5_ASAP7_75t_L g38 ( 
.A(n_33),
.B(n_34),
.C(n_35),
.Y(n_38)
);

O2A1O1Ixp33_ASAP7_75t_SL g36 ( 
.A1(n_29),
.A2(n_30),
.B(n_31),
.C(n_27),
.Y(n_36)
);

OAI21xp5_ASAP7_75t_SL g37 ( 
.A1(n_36),
.A2(n_28),
.B(n_29),
.Y(n_37)
);

OR2x2_ASAP7_75t_L g40 ( 
.A(n_37),
.B(n_39),
.Y(n_40)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_36),
.Y(n_39)
);

MAJx2_ASAP7_75t_L g41 ( 
.A(n_40),
.B(n_38),
.C(n_34),
.Y(n_41)
);


endmodule