module fake_jpeg_29435_n_313 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_313);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_313;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_256;
wire n_221;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

INVx11_ASAP7_75t_SL g19 ( 
.A(n_5),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_1),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_11),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_3),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_8),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_7),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

BUFx10_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_9),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_1),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_1),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_4),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_16),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_7),
.Y(n_39)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_9),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_13),
.Y(n_41)
);

BUFx5_ASAP7_75t_L g42 ( 
.A(n_12),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_17),
.Y(n_43)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_43),
.Y(n_79)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_40),
.Y(n_44)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_44),
.Y(n_70)
);

INVx4_ASAP7_75t_SL g45 ( 
.A(n_42),
.Y(n_45)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_45),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g46 ( 
.A1(n_18),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_46),
.A2(n_26),
.B1(n_39),
.B2(n_34),
.Y(n_68)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_42),
.Y(n_47)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_47),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_33),
.B(n_16),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_48),
.B(n_51),
.Y(n_73)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_19),
.Y(n_49)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_49),
.Y(n_89)
);

INVx11_ASAP7_75t_L g50 ( 
.A(n_18),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_50),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_32),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_17),
.Y(n_52)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_52),
.Y(n_102)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_21),
.Y(n_53)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_53),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_18),
.Y(n_54)
);

BUFx2_ASAP7_75t_L g88 ( 
.A(n_54),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g55 ( 
.A(n_40),
.B(n_0),
.C(n_2),
.Y(n_55)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_55),
.B(n_35),
.C(n_29),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_33),
.B(n_15),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_56),
.B(n_57),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_41),
.B(n_14),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_32),
.B(n_0),
.Y(n_58)
);

AND2x2_ASAP7_75t_L g108 ( 
.A(n_58),
.B(n_67),
.Y(n_108)
);

INVx2_ASAP7_75t_R g59 ( 
.A(n_20),
.Y(n_59)
);

CKINVDCx14_ASAP7_75t_R g87 ( 
.A(n_59),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_32),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_60),
.B(n_25),
.Y(n_81)
);

INVx13_ASAP7_75t_L g61 ( 
.A(n_40),
.Y(n_61)
);

CKINVDCx5p33_ASAP7_75t_R g71 ( 
.A(n_61),
.Y(n_71)
);

HB1xp67_ASAP7_75t_L g62 ( 
.A(n_28),
.Y(n_62)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_62),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_28),
.Y(n_63)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_63),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_28),
.Y(n_64)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_64),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_31),
.Y(n_65)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_65),
.Y(n_98)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_31),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_66),
.Y(n_69)
);

BUFx5_ASAP7_75t_L g67 ( 
.A(n_31),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_68),
.B(n_78),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_59),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_72),
.B(n_76),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_SL g74 ( 
.A(n_59),
.B(n_26),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g113 ( 
.A(n_74),
.B(n_91),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_66),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_45),
.A2(n_30),
.B1(n_27),
.B2(n_38),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_77),
.A2(n_97),
.B1(n_99),
.B2(n_110),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_58),
.B(n_32),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_55),
.B(n_32),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_80),
.B(n_103),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_81),
.B(n_82),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_47),
.Y(n_82)
);

OR2x2_ASAP7_75t_L g84 ( 
.A(n_43),
.B(n_25),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_84),
.B(n_86),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_52),
.B(n_41),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_53),
.B(n_39),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_90),
.B(n_100),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_SL g91 ( 
.A(n_51),
.B(n_23),
.Y(n_91)
);

AOI21xp33_ASAP7_75t_L g92 ( 
.A1(n_46),
.A2(n_24),
.B(n_37),
.Y(n_92)
);

AOI21xp33_ASAP7_75t_L g137 ( 
.A1(n_92),
.A2(n_6),
.B(n_10),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_60),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_SL g132 ( 
.A(n_93),
.B(n_67),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_45),
.A2(n_30),
.B1(n_38),
.B2(n_27),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_44),
.A2(n_30),
.B1(n_38),
.B2(n_27),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_61),
.B(n_36),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_49),
.B(n_36),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_101),
.B(n_106),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_50),
.A2(n_35),
.B1(n_34),
.B2(n_29),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_105),
.B(n_4),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_49),
.B(n_20),
.Y(n_106)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_49),
.Y(n_107)
);

INVxp67_ASAP7_75t_SL g143 ( 
.A(n_107),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_64),
.A2(n_37),
.B1(n_24),
.B2(n_22),
.Y(n_110)
);

INVx8_ASAP7_75t_L g112 ( 
.A(n_94),
.Y(n_112)
);

INVx4_ASAP7_75t_L g164 ( 
.A(n_112),
.Y(n_164)
);

INVx5_ASAP7_75t_L g116 ( 
.A(n_89),
.Y(n_116)
);

INVx1_ASAP7_75t_SL g158 ( 
.A(n_116),
.Y(n_158)
);

OR2x2_ASAP7_75t_L g117 ( 
.A(n_72),
.B(n_23),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_L g163 ( 
.A1(n_117),
.A2(n_146),
.B(n_71),
.Y(n_163)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_98),
.Y(n_118)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_118),
.Y(n_174)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_79),
.Y(n_119)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_119),
.Y(n_171)
);

AOI21xp5_ASAP7_75t_L g123 ( 
.A1(n_80),
.A2(n_21),
.B(n_22),
.Y(n_123)
);

AOI21xp5_ASAP7_75t_L g149 ( 
.A1(n_123),
.A2(n_135),
.B(n_107),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_78),
.B(n_65),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_124),
.B(n_127),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_73),
.B(n_4),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_SL g180 ( 
.A(n_125),
.B(n_129),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_126),
.B(n_105),
.C(n_87),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_108),
.B(n_65),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_75),
.B(n_5),
.Y(n_129)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_98),
.Y(n_130)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_130),
.Y(n_154)
);

INVx3_ASAP7_75t_L g131 ( 
.A(n_89),
.Y(n_131)
);

INVx2_ASAP7_75t_SL g170 ( 
.A(n_131),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_132),
.B(n_138),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_108),
.B(n_54),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_133),
.B(n_134),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_108),
.B(n_54),
.Y(n_134)
);

NAND2x1_ASAP7_75t_SL g135 ( 
.A(n_71),
.B(n_83),
.Y(n_135)
);

INVx4_ASAP7_75t_L g136 ( 
.A(n_83),
.Y(n_136)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_136),
.Y(n_155)
);

FAx1_ASAP7_75t_SL g177 ( 
.A(n_137),
.B(n_11),
.CI(n_12),
.CON(n_177),
.SN(n_177)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_74),
.B(n_6),
.Y(n_138)
);

INVx1_ASAP7_75t_SL g139 ( 
.A(n_95),
.Y(n_139)
);

AND2x2_ASAP7_75t_L g157 ( 
.A(n_139),
.B(n_109),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g141 ( 
.A(n_94),
.Y(n_141)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_141),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_91),
.B(n_10),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_142),
.B(n_145),
.Y(n_162)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_79),
.Y(n_144)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_144),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_84),
.B(n_10),
.Y(n_145)
);

OR2x2_ASAP7_75t_L g146 ( 
.A(n_93),
.B(n_11),
.Y(n_146)
);

CKINVDCx16_ASAP7_75t_R g147 ( 
.A(n_95),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_147),
.B(n_82),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_148),
.B(n_159),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_SL g189 ( 
.A1(n_149),
.A2(n_146),
.B(n_117),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_115),
.A2(n_68),
.B1(n_104),
.B2(n_102),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_150),
.A2(n_160),
.B1(n_165),
.B2(n_173),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_124),
.B(n_104),
.C(n_102),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_152),
.B(n_131),
.C(n_112),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_115),
.A2(n_103),
.B1(n_109),
.B2(n_63),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_153),
.A2(n_172),
.B1(n_148),
.B2(n_181),
.Y(n_196)
);

INVxp67_ASAP7_75t_L g203 ( 
.A(n_157),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_128),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_114),
.A2(n_63),
.B1(n_96),
.B2(n_85),
.Y(n_160)
);

NAND2xp67_ASAP7_75t_SL g205 ( 
.A(n_163),
.B(n_177),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_114),
.A2(n_96),
.B1(n_85),
.B2(n_88),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_123),
.B(n_76),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_166),
.B(n_111),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_168),
.B(n_179),
.Y(n_195)
);

INVxp67_ASAP7_75t_L g169 ( 
.A(n_135),
.Y(n_169)
);

INVx13_ASAP7_75t_L g209 ( 
.A(n_169),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_133),
.A2(n_126),
.B1(n_122),
.B2(n_127),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_134),
.A2(n_144),
.B1(n_119),
.B2(n_111),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_120),
.B(n_70),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_SL g198 ( 
.A(n_176),
.B(n_178),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_128),
.B(n_70),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_140),
.B(n_69),
.Y(n_179)
);

INVxp67_ASAP7_75t_L g181 ( 
.A(n_135),
.Y(n_181)
);

INVxp33_ASAP7_75t_L g183 ( 
.A(n_181),
.Y(n_183)
);

AO22x1_ASAP7_75t_L g182 ( 
.A1(n_147),
.A2(n_69),
.B1(n_88),
.B2(n_94),
.Y(n_182)
);

AOI21xp5_ASAP7_75t_SL g186 ( 
.A1(n_182),
.A2(n_139),
.B(n_116),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_L g184 ( 
.A1(n_149),
.A2(n_146),
.B(n_132),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_L g226 ( 
.A1(n_184),
.A2(n_194),
.B(n_170),
.Y(n_226)
);

OAI21xp33_ASAP7_75t_L g216 ( 
.A1(n_185),
.A2(n_177),
.B(n_180),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_SL g234 ( 
.A1(n_186),
.A2(n_213),
.B(n_203),
.Y(n_234)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_171),
.Y(n_187)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_187),
.Y(n_220)
);

AOI21xp5_ASAP7_75t_L g232 ( 
.A1(n_189),
.A2(n_164),
.B(n_167),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_157),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_190),
.B(n_192),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_150),
.A2(n_88),
.B1(n_121),
.B2(n_118),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_191),
.A2(n_200),
.B1(n_188),
.B2(n_203),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_157),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_L g194 ( 
.A1(n_166),
.A2(n_117),
.B(n_140),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_196),
.A2(n_207),
.B1(n_208),
.B2(n_170),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_182),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_197),
.B(n_204),
.Y(n_221)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_171),
.Y(n_199)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_199),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_173),
.A2(n_130),
.B1(n_113),
.B2(n_136),
.Y(n_200)
);

MAJx2_ASAP7_75t_L g201 ( 
.A(n_152),
.B(n_113),
.C(n_143),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_SL g230 ( 
.A(n_201),
.B(n_202),
.Y(n_230)
);

AND2x6_ASAP7_75t_L g204 ( 
.A(n_172),
.B(n_112),
.Y(n_204)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_175),
.Y(n_206)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_206),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_153),
.A2(n_12),
.B1(n_141),
.B2(n_151),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_L g208 ( 
.A1(n_151),
.A2(n_141),
.B1(n_169),
.B2(n_156),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_156),
.B(n_163),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_210),
.B(n_212),
.Y(n_235)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_154),
.Y(n_211)
);

CKINVDCx16_ASAP7_75t_R g225 ( 
.A(n_211),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_161),
.B(n_160),
.Y(n_212)
);

AOI21xp5_ASAP7_75t_SL g213 ( 
.A1(n_182),
.A2(n_177),
.B(n_162),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_193),
.B(n_165),
.C(n_155),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_214),
.B(n_219),
.Y(n_248)
);

A2O1A1O1Ixp25_ASAP7_75t_L g241 ( 
.A1(n_216),
.A2(n_226),
.B(n_205),
.C(n_183),
.D(n_209),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_185),
.B(n_210),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_217),
.B(n_224),
.Y(n_244)
);

CKINVDCx14_ASAP7_75t_R g218 ( 
.A(n_198),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_218),
.B(n_223),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_196),
.B(n_158),
.C(n_174),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_195),
.B(n_200),
.Y(n_222)
);

INVxp67_ASAP7_75t_L g239 ( 
.A(n_222),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_186),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_202),
.B(n_158),
.C(n_174),
.Y(n_224)
);

CKINVDCx14_ASAP7_75t_R g228 ( 
.A(n_213),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_228),
.B(n_229),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_201),
.B(n_170),
.C(n_164),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_231),
.B(n_237),
.Y(n_251)
);

OAI21xp5_ASAP7_75t_SL g247 ( 
.A1(n_232),
.A2(n_183),
.B(n_209),
.Y(n_247)
);

INVxp67_ASAP7_75t_L g243 ( 
.A(n_233),
.Y(n_243)
);

INVxp67_ASAP7_75t_L g257 ( 
.A(n_234),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_191),
.B(n_212),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_236),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_194),
.B(n_184),
.C(n_189),
.Y(n_237)
);

XOR2xp5_ASAP7_75t_L g261 ( 
.A(n_241),
.B(n_226),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_215),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_242),
.B(n_245),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_225),
.Y(n_245)
);

AOI21xp5_ASAP7_75t_L g260 ( 
.A1(n_247),
.A2(n_255),
.B(n_258),
.Y(n_260)
);

INVx6_ASAP7_75t_L g250 ( 
.A(n_225),
.Y(n_250)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_250),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_217),
.B(n_207),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_252),
.Y(n_264)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_227),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_253),
.Y(n_266)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_227),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_SL g262 ( 
.A(n_254),
.B(n_256),
.Y(n_262)
);

BUFx12f_ASAP7_75t_SL g255 ( 
.A(n_234),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_238),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_238),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_243),
.A2(n_221),
.B1(n_223),
.B2(n_231),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_L g274 ( 
.A1(n_259),
.A2(n_263),
.B1(n_272),
.B2(n_252),
.Y(n_274)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_261),
.B(n_268),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_251),
.A2(n_219),
.B1(n_204),
.B2(n_235),
.Y(n_263)
);

BUFx12_ASAP7_75t_L g267 ( 
.A(n_255),
.Y(n_267)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_267),
.Y(n_277)
);

XOR2xp5_ASAP7_75t_L g268 ( 
.A(n_248),
.B(n_230),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_L g269 ( 
.A(n_248),
.B(n_230),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_269),
.B(n_270),
.Y(n_282)
);

XOR2xp5_ASAP7_75t_L g270 ( 
.A(n_249),
.B(n_237),
.Y(n_270)
);

AND2x2_ASAP7_75t_L g271 ( 
.A(n_246),
.B(n_205),
.Y(n_271)
);

AOI21xp5_ASAP7_75t_L g284 ( 
.A1(n_271),
.A2(n_247),
.B(n_240),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_251),
.A2(n_246),
.B1(n_239),
.B2(n_257),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_SL g286 ( 
.A1(n_274),
.A2(n_275),
.B1(n_263),
.B2(n_272),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_264),
.A2(n_249),
.B1(n_240),
.B2(n_244),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_SL g276 ( 
.A(n_265),
.B(n_242),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_276),
.B(n_280),
.Y(n_287)
);

AOI21xp5_ASAP7_75t_SL g278 ( 
.A1(n_260),
.A2(n_232),
.B(n_235),
.Y(n_278)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_278),
.Y(n_292)
);

FAx1_ASAP7_75t_SL g280 ( 
.A(n_271),
.B(n_244),
.CI(n_229),
.CON(n_280),
.SN(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_262),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_281),
.B(n_245),
.Y(n_288)
);

OAI21xp5_ASAP7_75t_SL g283 ( 
.A1(n_267),
.A2(n_214),
.B(n_224),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_SL g289 ( 
.A(n_283),
.B(n_285),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g290 ( 
.A(n_284),
.B(n_261),
.Y(n_290)
);

AOI21xp5_ASAP7_75t_L g285 ( 
.A1(n_267),
.A2(n_233),
.B(n_258),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_286),
.B(n_290),
.Y(n_297)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_288),
.Y(n_295)
);

OR2x2_ASAP7_75t_L g291 ( 
.A(n_277),
.B(n_259),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_291),
.B(n_293),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_282),
.B(n_270),
.C(n_269),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_282),
.B(n_268),
.C(n_273),
.Y(n_294)
);

OAI21xp5_ASAP7_75t_L g301 ( 
.A1(n_294),
.A2(n_280),
.B(n_279),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_292),
.A2(n_275),
.B1(n_285),
.B2(n_284),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_296),
.B(n_298),
.Y(n_302)
);

NOR3xp33_ASAP7_75t_SL g298 ( 
.A(n_287),
.B(n_241),
.C(n_278),
.Y(n_298)
);

NOR2xp67_ASAP7_75t_L g299 ( 
.A(n_289),
.B(n_280),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_299),
.B(n_266),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_L g304 ( 
.A(n_301),
.B(n_294),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_300),
.B(n_291),
.Y(n_303)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_303),
.Y(n_308)
);

OAI21xp5_ASAP7_75t_SL g309 ( 
.A1(n_304),
.A2(n_305),
.B(n_306),
.Y(n_309)
);

AOI21xp5_ASAP7_75t_L g305 ( 
.A1(n_295),
.A2(n_293),
.B(n_279),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_L g307 ( 
.A1(n_302),
.A2(n_298),
.B1(n_254),
.B2(n_256),
.Y(n_307)
);

AOI322xp5_ASAP7_75t_L g311 ( 
.A1(n_307),
.A2(n_250),
.A3(n_220),
.B1(n_199),
.B2(n_206),
.C1(n_297),
.C2(n_188),
.Y(n_311)
);

NOR5xp2_ASAP7_75t_L g310 ( 
.A(n_309),
.B(n_304),
.C(n_297),
.D(n_250),
.E(n_253),
.Y(n_310)
);

NAND4xp25_ASAP7_75t_L g312 ( 
.A(n_310),
.B(n_311),
.C(n_308),
.D(n_220),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_L g313 ( 
.A(n_312),
.B(n_211),
.Y(n_313)
);


endmodule