module fake_ibex_80_n_3731 (n_151, n_85, n_599, n_507, n_540, n_395, n_84, n_64, n_171, n_103, n_529, n_389, n_204, n_274, n_387, n_130, n_177, n_76, n_273, n_309, n_330, n_9, n_328, n_293, n_341, n_372, n_124, n_37, n_256, n_418, n_193, n_510, n_446, n_108, n_350, n_601, n_621, n_610, n_165, n_452, n_86, n_70, n_255, n_175, n_586, n_398, n_59, n_28, n_125, n_304, n_191, n_593, n_5, n_62, n_71, n_153, n_545, n_583, n_194, n_249, n_334, n_312, n_578, n_478, n_239, n_94, n_134, n_432, n_371, n_403, n_423, n_608, n_357, n_88, n_412, n_457, n_494, n_142, n_226, n_336, n_258, n_40, n_90, n_17, n_74, n_449, n_547, n_176, n_58, n_43, n_216, n_33, n_421, n_475, n_166, n_163, n_500, n_542, n_114, n_236, n_34, n_376, n_377, n_584, n_531, n_15, n_556, n_24, n_189, n_498, n_280, n_317, n_340, n_375, n_105, n_187, n_1, n_154, n_182, n_196, n_326, n_327, n_89, n_50, n_144, n_170, n_270, n_346, n_383, n_113, n_561, n_117, n_417, n_471, n_265, n_504, n_158, n_259, n_276, n_339, n_470, n_210, n_348, n_220, n_91, n_481, n_287, n_54, n_243, n_19, n_497, n_228, n_147, n_552, n_251, n_384, n_373, n_458, n_244, n_73, n_343, n_310, n_426, n_323, n_469, n_598, n_143, n_106, n_386, n_549, n_8, n_224, n_183, n_533, n_508, n_67, n_453, n_591, n_333, n_110, n_306, n_400, n_47, n_550, n_169, n_10, n_21, n_242, n_278, n_316, n_16, n_404, n_60, n_557, n_7, n_109, n_127, n_121, n_527, n_590, n_465, n_48, n_325, n_57, n_301, n_496, n_617, n_434, n_296, n_120, n_168, n_526, n_155, n_315, n_441, n_604, n_13, n_122, n_523, n_116, n_614, n_370, n_431, n_574, n_0, n_289, n_12, n_515, n_150, n_286, n_321, n_133, n_569, n_600, n_51, n_215, n_279, n_49, n_374, n_235, n_464, n_538, n_22, n_136, n_261, n_521, n_459, n_30, n_518, n_367, n_221, n_437, n_602, n_355, n_474, n_594, n_407, n_102, n_490, n_568, n_52, n_448, n_595, n_99, n_466, n_269, n_156, n_570, n_126, n_585, n_530, n_356, n_25, n_104, n_45, n_420, n_483, n_543, n_580, n_141, n_487, n_222, n_186, n_524, n_349, n_454, n_295, n_331, n_576, n_230, n_96, n_185, n_388, n_619, n_536, n_611, n_352, n_290, n_558, n_174, n_467, n_427, n_607, n_157, n_219, n_246, n_31, n_442, n_146, n_207, n_438, n_167, n_128, n_253, n_208, n_234, n_3, n_152, n_300, n_145, n_65, n_358, n_205, n_618, n_488, n_139, n_514, n_429, n_560, n_275, n_541, n_98, n_129, n_613, n_267, n_245, n_589, n_571, n_229, n_209, n_472, n_347, n_473, n_445, n_335, n_413, n_82, n_263, n_27, n_573, n_353, n_359, n_299, n_87, n_262, n_433, n_75, n_439, n_137, n_338, n_173, n_477, n_363, n_402, n_180, n_369, n_596, n_201, n_14, n_351, n_368, n_456, n_257, n_77, n_44, n_401, n_553, n_554, n_66, n_305, n_307, n_192, n_140, n_484, n_566, n_480, n_416, n_581, n_365, n_4, n_6, n_605, n_539, n_100, n_179, n_354, n_206, n_392, n_516, n_548, n_567, n_329, n_447, n_26, n_188, n_200, n_444, n_506, n_562, n_564, n_546, n_199, n_592, n_495, n_410, n_308, n_463, n_411, n_135, n_520, n_512, n_615, n_283, n_366, n_397, n_111, n_36, n_18, n_322, n_53, n_227, n_499, n_115, n_11, n_248, n_92, n_451, n_101, n_190, n_138, n_409, n_582, n_214, n_238, n_579, n_332, n_517, n_211, n_218, n_314, n_563, n_132, n_277, n_555, n_337, n_522, n_479, n_534, n_225, n_360, n_272, n_511, n_23, n_468, n_223, n_381, n_525, n_535, n_382, n_502, n_532, n_95, n_405, n_415, n_597, n_285, n_288, n_247, n_320, n_379, n_551, n_55, n_612, n_291, n_318, n_63, n_161, n_237, n_29, n_203, n_268, n_440, n_148, n_2, n_342, n_233, n_385, n_414, n_430, n_118, n_603, n_378, n_486, n_422, n_164, n_38, n_198, n_264, n_616, n_217, n_324, n_391, n_537, n_78, n_20, n_69, n_390, n_544, n_39, n_178, n_509, n_303, n_362, n_93, n_505, n_162, n_482, n_240, n_282, n_61, n_501, n_266, n_42, n_294, n_112, n_485, n_46, n_284, n_80, n_172, n_250, n_493, n_460, n_609, n_476, n_461, n_575, n_313, n_519, n_345, n_408, n_119, n_361, n_455, n_419, n_72, n_319, n_195, n_513, n_212, n_588, n_311, n_406, n_606, n_97, n_197, n_528, n_181, n_131, n_123, n_260, n_620, n_462, n_302, n_450, n_443, n_572, n_577, n_344, n_393, n_436, n_428, n_491, n_297, n_435, n_41, n_252, n_396, n_83, n_32, n_107, n_149, n_489, n_399, n_254, n_213, n_424, n_565, n_271, n_241, n_68, n_503, n_292, n_394, n_79, n_81, n_35, n_364, n_159, n_202, n_231, n_298, n_587, n_160, n_184, n_56, n_492, n_232, n_380, n_281, n_559, n_425, n_3731);

input n_151;
input n_85;
input n_599;
input n_507;
input n_540;
input n_395;
input n_84;
input n_64;
input n_171;
input n_103;
input n_529;
input n_389;
input n_204;
input n_274;
input n_387;
input n_130;
input n_177;
input n_76;
input n_273;
input n_309;
input n_330;
input n_9;
input n_328;
input n_293;
input n_341;
input n_372;
input n_124;
input n_37;
input n_256;
input n_418;
input n_193;
input n_510;
input n_446;
input n_108;
input n_350;
input n_601;
input n_621;
input n_610;
input n_165;
input n_452;
input n_86;
input n_70;
input n_255;
input n_175;
input n_586;
input n_398;
input n_59;
input n_28;
input n_125;
input n_304;
input n_191;
input n_593;
input n_5;
input n_62;
input n_71;
input n_153;
input n_545;
input n_583;
input n_194;
input n_249;
input n_334;
input n_312;
input n_578;
input n_478;
input n_239;
input n_94;
input n_134;
input n_432;
input n_371;
input n_403;
input n_423;
input n_608;
input n_357;
input n_88;
input n_412;
input n_457;
input n_494;
input n_142;
input n_226;
input n_336;
input n_258;
input n_40;
input n_90;
input n_17;
input n_74;
input n_449;
input n_547;
input n_176;
input n_58;
input n_43;
input n_216;
input n_33;
input n_421;
input n_475;
input n_166;
input n_163;
input n_500;
input n_542;
input n_114;
input n_236;
input n_34;
input n_376;
input n_377;
input n_584;
input n_531;
input n_15;
input n_556;
input n_24;
input n_189;
input n_498;
input n_280;
input n_317;
input n_340;
input n_375;
input n_105;
input n_187;
input n_1;
input n_154;
input n_182;
input n_196;
input n_326;
input n_327;
input n_89;
input n_50;
input n_144;
input n_170;
input n_270;
input n_346;
input n_383;
input n_113;
input n_561;
input n_117;
input n_417;
input n_471;
input n_265;
input n_504;
input n_158;
input n_259;
input n_276;
input n_339;
input n_470;
input n_210;
input n_348;
input n_220;
input n_91;
input n_481;
input n_287;
input n_54;
input n_243;
input n_19;
input n_497;
input n_228;
input n_147;
input n_552;
input n_251;
input n_384;
input n_373;
input n_458;
input n_244;
input n_73;
input n_343;
input n_310;
input n_426;
input n_323;
input n_469;
input n_598;
input n_143;
input n_106;
input n_386;
input n_549;
input n_8;
input n_224;
input n_183;
input n_533;
input n_508;
input n_67;
input n_453;
input n_591;
input n_333;
input n_110;
input n_306;
input n_400;
input n_47;
input n_550;
input n_169;
input n_10;
input n_21;
input n_242;
input n_278;
input n_316;
input n_16;
input n_404;
input n_60;
input n_557;
input n_7;
input n_109;
input n_127;
input n_121;
input n_527;
input n_590;
input n_465;
input n_48;
input n_325;
input n_57;
input n_301;
input n_496;
input n_617;
input n_434;
input n_296;
input n_120;
input n_168;
input n_526;
input n_155;
input n_315;
input n_441;
input n_604;
input n_13;
input n_122;
input n_523;
input n_116;
input n_614;
input n_370;
input n_431;
input n_574;
input n_0;
input n_289;
input n_12;
input n_515;
input n_150;
input n_286;
input n_321;
input n_133;
input n_569;
input n_600;
input n_51;
input n_215;
input n_279;
input n_49;
input n_374;
input n_235;
input n_464;
input n_538;
input n_22;
input n_136;
input n_261;
input n_521;
input n_459;
input n_30;
input n_518;
input n_367;
input n_221;
input n_437;
input n_602;
input n_355;
input n_474;
input n_594;
input n_407;
input n_102;
input n_490;
input n_568;
input n_52;
input n_448;
input n_595;
input n_99;
input n_466;
input n_269;
input n_156;
input n_570;
input n_126;
input n_585;
input n_530;
input n_356;
input n_25;
input n_104;
input n_45;
input n_420;
input n_483;
input n_543;
input n_580;
input n_141;
input n_487;
input n_222;
input n_186;
input n_524;
input n_349;
input n_454;
input n_295;
input n_331;
input n_576;
input n_230;
input n_96;
input n_185;
input n_388;
input n_619;
input n_536;
input n_611;
input n_352;
input n_290;
input n_558;
input n_174;
input n_467;
input n_427;
input n_607;
input n_157;
input n_219;
input n_246;
input n_31;
input n_442;
input n_146;
input n_207;
input n_438;
input n_167;
input n_128;
input n_253;
input n_208;
input n_234;
input n_3;
input n_152;
input n_300;
input n_145;
input n_65;
input n_358;
input n_205;
input n_618;
input n_488;
input n_139;
input n_514;
input n_429;
input n_560;
input n_275;
input n_541;
input n_98;
input n_129;
input n_613;
input n_267;
input n_245;
input n_589;
input n_571;
input n_229;
input n_209;
input n_472;
input n_347;
input n_473;
input n_445;
input n_335;
input n_413;
input n_82;
input n_263;
input n_27;
input n_573;
input n_353;
input n_359;
input n_299;
input n_87;
input n_262;
input n_433;
input n_75;
input n_439;
input n_137;
input n_338;
input n_173;
input n_477;
input n_363;
input n_402;
input n_180;
input n_369;
input n_596;
input n_201;
input n_14;
input n_351;
input n_368;
input n_456;
input n_257;
input n_77;
input n_44;
input n_401;
input n_553;
input n_554;
input n_66;
input n_305;
input n_307;
input n_192;
input n_140;
input n_484;
input n_566;
input n_480;
input n_416;
input n_581;
input n_365;
input n_4;
input n_6;
input n_605;
input n_539;
input n_100;
input n_179;
input n_354;
input n_206;
input n_392;
input n_516;
input n_548;
input n_567;
input n_329;
input n_447;
input n_26;
input n_188;
input n_200;
input n_444;
input n_506;
input n_562;
input n_564;
input n_546;
input n_199;
input n_592;
input n_495;
input n_410;
input n_308;
input n_463;
input n_411;
input n_135;
input n_520;
input n_512;
input n_615;
input n_283;
input n_366;
input n_397;
input n_111;
input n_36;
input n_18;
input n_322;
input n_53;
input n_227;
input n_499;
input n_115;
input n_11;
input n_248;
input n_92;
input n_451;
input n_101;
input n_190;
input n_138;
input n_409;
input n_582;
input n_214;
input n_238;
input n_579;
input n_332;
input n_517;
input n_211;
input n_218;
input n_314;
input n_563;
input n_132;
input n_277;
input n_555;
input n_337;
input n_522;
input n_479;
input n_534;
input n_225;
input n_360;
input n_272;
input n_511;
input n_23;
input n_468;
input n_223;
input n_381;
input n_525;
input n_535;
input n_382;
input n_502;
input n_532;
input n_95;
input n_405;
input n_415;
input n_597;
input n_285;
input n_288;
input n_247;
input n_320;
input n_379;
input n_551;
input n_55;
input n_612;
input n_291;
input n_318;
input n_63;
input n_161;
input n_237;
input n_29;
input n_203;
input n_268;
input n_440;
input n_148;
input n_2;
input n_342;
input n_233;
input n_385;
input n_414;
input n_430;
input n_118;
input n_603;
input n_378;
input n_486;
input n_422;
input n_164;
input n_38;
input n_198;
input n_264;
input n_616;
input n_217;
input n_324;
input n_391;
input n_537;
input n_78;
input n_20;
input n_69;
input n_390;
input n_544;
input n_39;
input n_178;
input n_509;
input n_303;
input n_362;
input n_93;
input n_505;
input n_162;
input n_482;
input n_240;
input n_282;
input n_61;
input n_501;
input n_266;
input n_42;
input n_294;
input n_112;
input n_485;
input n_46;
input n_284;
input n_80;
input n_172;
input n_250;
input n_493;
input n_460;
input n_609;
input n_476;
input n_461;
input n_575;
input n_313;
input n_519;
input n_345;
input n_408;
input n_119;
input n_361;
input n_455;
input n_419;
input n_72;
input n_319;
input n_195;
input n_513;
input n_212;
input n_588;
input n_311;
input n_406;
input n_606;
input n_97;
input n_197;
input n_528;
input n_181;
input n_131;
input n_123;
input n_260;
input n_620;
input n_462;
input n_302;
input n_450;
input n_443;
input n_572;
input n_577;
input n_344;
input n_393;
input n_436;
input n_428;
input n_491;
input n_297;
input n_435;
input n_41;
input n_252;
input n_396;
input n_83;
input n_32;
input n_107;
input n_149;
input n_489;
input n_399;
input n_254;
input n_213;
input n_424;
input n_565;
input n_271;
input n_241;
input n_68;
input n_503;
input n_292;
input n_394;
input n_79;
input n_81;
input n_35;
input n_364;
input n_159;
input n_202;
input n_231;
input n_298;
input n_587;
input n_160;
input n_184;
input n_56;
input n_492;
input n_232;
input n_380;
input n_281;
input n_559;
input n_425;

output n_3731;

wire n_1084;
wire n_2594;
wire n_1474;
wire n_1295;
wire n_1983;
wire n_2804;
wire n_3150;
wire n_992;
wire n_1582;
wire n_2201;
wire n_2512;
wire n_766;
wire n_3590;
wire n_2960;
wire n_2175;
wire n_2071;
wire n_2796;
wire n_1110;
wire n_3548;
wire n_2607;
wire n_1382;
wire n_3610;
wire n_3144;
wire n_2569;
wire n_2949;
wire n_1998;
wire n_2840;
wire n_1596;
wire n_926;
wire n_3319;
wire n_1079;
wire n_3077;
wire n_2835;
wire n_1100;
wire n_3559;
wire n_845;
wire n_2177;
wire n_1930;
wire n_2123;
wire n_1234;
wire n_3019;
wire n_2047;
wire n_1594;
wire n_1944;
wire n_2235;
wire n_1802;
wire n_2498;
wire n_773;
wire n_2038;
wire n_2504;
wire n_1469;
wire n_821;
wire n_2017;
wire n_873;
wire n_1227;
wire n_962;
wire n_1080;
wire n_862;
wire n_909;
wire n_2290;
wire n_957;
wire n_3255;
wire n_3272;
wire n_3674;
wire n_1652;
wire n_678;
wire n_969;
wire n_1859;
wire n_1954;
wire n_2183;
wire n_2074;
wire n_2897;
wire n_1883;
wire n_1125;
wire n_733;
wire n_2687;
wire n_3456;
wire n_2037;
wire n_622;
wire n_1226;
wire n_1034;
wire n_2383;
wire n_3132;
wire n_1765;
wire n_872;
wire n_2392;
wire n_1873;
wire n_1619;
wire n_1666;
wire n_2682;
wire n_2640;
wire n_3605;
wire n_930;
wire n_1044;
wire n_3280;
wire n_3105;
wire n_3146;
wire n_1492;
wire n_1134;
wire n_1478;
wire n_1684;
wire n_1796;
wire n_3569;
wire n_1614;
wire n_2374;
wire n_3334;
wire n_2598;
wire n_1722;
wire n_911;
wire n_2023;
wire n_652;
wire n_781;
wire n_2720;
wire n_802;
wire n_3340;
wire n_2322;
wire n_1233;
wire n_2335;
wire n_3025;
wire n_3411;
wire n_2955;
wire n_3458;
wire n_3653;
wire n_3519;
wire n_2276;
wire n_1045;
wire n_3235;
wire n_2989;
wire n_1856;
wire n_963;
wire n_1782;
wire n_2230;
wire n_2889;
wire n_2139;
wire n_2847;
wire n_3693;
wire n_3033;
wire n_1308;
wire n_1138;
wire n_2943;
wire n_708;
wire n_1096;
wire n_2151;
wire n_2391;
wire n_1391;
wire n_3338;
wire n_3168;
wire n_667;
wire n_884;
wire n_2396;
wire n_3135;
wire n_3440;
wire n_850;
wire n_3175;
wire n_3729;
wire n_3484;
wire n_1971;
wire n_2485;
wire n_2479;
wire n_3570;
wire n_879;
wire n_2179;
wire n_1957;
wire n_2188;
wire n_723;
wire n_1144;
wire n_2359;
wire n_2360;
wire n_2506;
wire n_1392;
wire n_2158;
wire n_1268;
wire n_2571;
wire n_3187;
wire n_739;
wire n_3598;
wire n_2724;
wire n_3086;
wire n_2475;
wire n_853;
wire n_3721;
wire n_948;
wire n_2799;
wire n_1752;
wire n_1829;
wire n_1338;
wire n_3726;
wire n_1730;
wire n_875;
wire n_1307;
wire n_1327;
wire n_2644;
wire n_876;
wire n_3211;
wire n_3479;
wire n_711;
wire n_1840;
wire n_2837;
wire n_671;
wire n_989;
wire n_3262;
wire n_3407;
wire n_1908;
wire n_3315;
wire n_3537;
wire n_1668;
wire n_2343;
wire n_2605;
wire n_2887;
wire n_1641;
wire n_829;
wire n_2565;
wire n_825;
wire n_1480;
wire n_1463;
wire n_1823;
wire n_3251;
wire n_1681;
wire n_2921;
wire n_3724;
wire n_939;
wire n_1636;
wire n_1687;
wire n_655;
wire n_3192;
wire n_3533;
wire n_2192;
wire n_1766;
wire n_3184;
wire n_3566;
wire n_3469;
wire n_3170;
wire n_1922;
wire n_2032;
wire n_2820;
wire n_3323;
wire n_641;
wire n_1937;
wire n_2311;
wire n_3392;
wire n_3347;
wire n_893;
wire n_3242;
wire n_3395;
wire n_1654;
wire n_3577;
wire n_2995;
wire n_3330;
wire n_1258;
wire n_1344;
wire n_2208;
wire n_2198;
wire n_1929;
wire n_2707;
wire n_3472;
wire n_3509;
wire n_1749;
wire n_1680;
wire n_835;
wire n_1981;
wire n_1195;
wire n_2918;
wire n_3353;
wire n_824;
wire n_1945;
wire n_2638;
wire n_694;
wire n_787;
wire n_2860;
wire n_2448;
wire n_3631;
wire n_2015;
wire n_2537;
wire n_1130;
wire n_2643;
wire n_1228;
wire n_2998;
wire n_2336;
wire n_3641;
wire n_2163;
wire n_1081;
wire n_2354;
wire n_3639;
wire n_1155;
wire n_1292;
wire n_2432;
wire n_3043;
wire n_2873;
wire n_1576;
wire n_1664;
wire n_2273;
wire n_3298;
wire n_852;
wire n_1427;
wire n_1133;
wire n_3049;
wire n_2421;
wire n_1926;
wire n_3208;
wire n_904;
wire n_2363;
wire n_2814;
wire n_3237;
wire n_3264;
wire n_3204;
wire n_2003;
wire n_1970;
wire n_3671;
wire n_3727;
wire n_2621;
wire n_3620;
wire n_1778;
wire n_646;
wire n_2558;
wire n_2953;
wire n_2922;
wire n_2347;
wire n_3507;
wire n_3103;
wire n_2839;
wire n_1030;
wire n_1698;
wire n_3688;
wire n_1094;
wire n_2462;
wire n_1496;
wire n_1910;
wire n_715;
wire n_2436;
wire n_1663;
wire n_2705;
wire n_1214;
wire n_1274;
wire n_2333;
wire n_2527;
wire n_1606;
wire n_769;
wire n_1595;
wire n_2164;
wire n_3711;
wire n_1509;
wire n_1648;
wire n_1618;
wire n_2944;
wire n_1886;
wire n_2269;
wire n_857;
wire n_765;
wire n_1070;
wire n_2472;
wire n_1841;
wire n_777;
wire n_2846;
wire n_3197;
wire n_2685;
wire n_3668;
wire n_1955;
wire n_3699;
wire n_917;
wire n_2413;
wire n_3022;
wire n_2362;
wire n_968;
wire n_2249;
wire n_3148;
wire n_2822;
wire n_1253;
wire n_3707;
wire n_1306;
wire n_1484;
wire n_2686;
wire n_1493;
wire n_2597;
wire n_1313;
wire n_2774;
wire n_3151;
wire n_2090;
wire n_666;
wire n_2260;
wire n_3722;
wire n_3125;
wire n_2812;
wire n_3681;
wire n_2753;
wire n_3603;
wire n_1638;
wire n_2215;
wire n_1071;
wire n_1449;
wire n_1960;
wire n_2663;
wire n_1723;
wire n_793;
wire n_3129;
wire n_937;
wire n_2595;
wire n_2116;
wire n_3714;
wire n_3592;
wire n_1645;
wire n_3186;
wire n_973;
wire n_1038;
wire n_2280;
wire n_1943;
wire n_3541;
wire n_1863;
wire n_2844;
wire n_1269;
wire n_2393;
wire n_2773;
wire n_3565;
wire n_662;
wire n_2906;
wire n_3030;
wire n_3097;
wire n_979;
wire n_1309;
wire n_1999;
wire n_3718;
wire n_1316;
wire n_1562;
wire n_1215;
wire n_629;
wire n_3679;
wire n_3579;
wire n_2777;
wire n_2480;
wire n_1445;
wire n_2806;
wire n_2283;
wire n_2813;
wire n_2147;
wire n_1716;
wire n_1466;
wire n_1412;
wire n_3210;
wire n_3221;
wire n_3667;
wire n_1672;
wire n_1007;
wire n_2253;
wire n_643;
wire n_1276;
wire n_1637;
wire n_3310;
wire n_841;
wire n_2900;
wire n_772;
wire n_810;
wire n_1401;
wire n_1817;
wire n_2951;
wire n_2145;
wire n_2122;
wire n_1588;
wire n_2216;
wire n_1301;
wire n_2579;
wire n_2876;
wire n_2242;
wire n_869;
wire n_1620;
wire n_1561;
wire n_718;
wire n_3301;
wire n_2370;
wire n_2025;
wire n_1078;
wire n_2247;
wire n_3451;
wire n_1219;
wire n_713;
wire n_1865;
wire n_3177;
wire n_3518;
wire n_3399;
wire n_1252;
wire n_2022;
wire n_2730;
wire n_1170;
wire n_1927;
wire n_2373;
wire n_630;
wire n_1869;
wire n_1853;
wire n_2275;
wire n_2980;
wire n_2189;
wire n_2482;
wire n_745;
wire n_2767;
wire n_3676;
wire n_2826;
wire n_2899;
wire n_2112;
wire n_1753;
wire n_3351;
wire n_1322;
wire n_2008;
wire n_1305;
wire n_2088;
wire n_795;
wire n_1248;
wire n_2762;
wire n_2171;
wire n_3307;
wire n_762;
wire n_1388;
wire n_2859;
wire n_800;
wire n_2564;
wire n_706;
wire n_3023;
wire n_784;
wire n_684;
wire n_1653;
wire n_1375;
wire n_3224;
wire n_1356;
wire n_894;
wire n_1118;
wire n_692;
wire n_2591;
wire n_1881;
wire n_1969;
wire n_709;
wire n_1296;
wire n_3060;
wire n_702;
wire n_1326;
wire n_971;
wire n_1350;
wire n_3627;
wire n_906;
wire n_2957;
wire n_2586;
wire n_1093;
wire n_1764;
wire n_2412;
wire n_2783;
wire n_978;
wire n_899;
wire n_3293;
wire n_1799;
wire n_1019;
wire n_902;
wire n_1689;
wire n_1250;
wire n_2550;
wire n_1190;
wire n_1304;
wire n_744;
wire n_2541;
wire n_2987;
wire n_881;
wire n_3259;
wire n_1702;
wire n_3381;
wire n_3630;
wire n_734;
wire n_1558;
wire n_2750;
wire n_1650;
wire n_1520;
wire n_1073;
wire n_1453;
wire n_1108;
wire n_2722;
wire n_2509;
wire n_2727;
wire n_3618;
wire n_1794;
wire n_1423;
wire n_1239;
wire n_2399;
wire n_1370;
wire n_2719;
wire n_1209;
wire n_1708;
wire n_2213;
wire n_3038;
wire n_3521;
wire n_3203;
wire n_3295;
wire n_2723;
wire n_1616;
wire n_3199;
wire n_3093;
wire n_729;
wire n_1569;
wire n_2664;
wire n_1434;
wire n_3716;
wire n_1649;
wire n_2389;
wire n_3450;
wire n_1936;
wire n_2114;
wire n_1717;
wire n_3567;
wire n_2107;
wire n_1609;
wire n_2257;
wire n_3435;
wire n_3530;
wire n_1613;
wire n_820;
wire n_805;
wire n_1988;
wire n_670;
wire n_1132;
wire n_892;
wire n_1467;
wire n_1803;
wire n_2401;
wire n_1787;
wire n_2782;
wire n_2511;
wire n_3217;
wire n_1281;
wire n_3094;
wire n_1447;
wire n_2166;
wire n_2451;
wire n_2150;
wire n_695;
wire n_1549;
wire n_639;
wire n_2631;
wire n_1867;
wire n_1531;
wire n_2919;
wire n_1332;
wire n_2660;
wire n_2661;
wire n_2292;
wire n_3573;
wire n_3563;
wire n_3510;
wire n_3560;
wire n_2334;
wire n_1424;
wire n_3467;
wire n_2444;
wire n_2625;
wire n_1742;
wire n_2350;
wire n_3652;
wire n_1818;
wire n_870;
wire n_2199;
wire n_1709;
wire n_1610;
wire n_2219;
wire n_1298;
wire n_1844;
wire n_1387;
wire n_2649;
wire n_1040;
wire n_2203;
wire n_2693;
wire n_3194;
wire n_3607;
wire n_3371;
wire n_1159;
wire n_1368;
wire n_2281;
wire n_1154;
wire n_3202;
wire n_2539;
wire n_2431;
wire n_1701;
wire n_2084;
wire n_1243;
wire n_3572;
wire n_2387;
wire n_2646;
wire n_3375;
wire n_2397;
wire n_1121;
wire n_693;
wire n_2746;
wire n_3241;
wire n_2256;
wire n_3317;
wire n_737;
wire n_2445;
wire n_3461;
wire n_2729;
wire n_1571;
wire n_1980;
wire n_3355;
wire n_2529;
wire n_3583;
wire n_2019;
wire n_1407;
wire n_3282;
wire n_1235;
wire n_1821;
wire n_3508;
wire n_1003;
wire n_889;
wire n_2708;
wire n_3156;
wire n_3457;
wire n_2748;
wire n_816;
wire n_1058;
wire n_1835;
wire n_2224;
wire n_1862;
wire n_2697;
wire n_3531;
wire n_3415;
wire n_2470;
wire n_2355;
wire n_2890;
wire n_3698;
wire n_2731;
wire n_1543;
wire n_3466;
wire n_3386;
wire n_823;
wire n_2233;
wire n_2499;
wire n_3370;
wire n_1504;
wire n_1519;
wire n_1425;
wire n_1781;
wire n_2069;
wire n_2602;
wire n_1441;
wire n_2028;
wire n_3309;
wire n_3678;
wire n_1924;
wire n_2856;
wire n_1921;
wire n_3024;
wire n_657;
wire n_1156;
wire n_2857;
wire n_1293;
wire n_1360;
wire n_749;
wire n_1555;
wire n_1394;
wire n_1347;
wire n_819;
wire n_2070;
wire n_822;
wire n_1042;
wire n_1888;
wire n_3471;
wire n_743;
wire n_3117;
wire n_3320;
wire n_754;
wire n_1786;
wire n_2033;
wire n_3039;
wire n_1319;
wire n_1553;
wire n_3478;
wire n_3701;
wire n_3542;
wire n_1041;
wire n_2766;
wire n_2828;
wire n_1964;
wire n_1090;
wire n_3720;
wire n_3374;
wire n_1196;
wire n_3704;
wire n_1182;
wire n_1271;
wire n_2416;
wire n_3633;
wire n_2786;
wire n_1731;
wire n_1905;
wire n_2962;
wire n_1031;
wire n_3416;
wire n_2879;
wire n_2958;
wire n_3147;
wire n_3694;
wire n_2052;
wire n_3690;
wire n_981;
wire n_3628;
wire n_2425;
wire n_2800;
wire n_3514;
wire n_3091;
wire n_3006;
wire n_3348;
wire n_2118;
wire n_2259;
wire n_2162;
wire n_2236;
wire n_3455;
wire n_3660;
wire n_2377;
wire n_2718;
wire n_2577;
wire n_1591;
wire n_3426;
wire n_3165;
wire n_2289;
wire n_2288;
wire n_2841;
wire n_3075;
wire n_1671;
wire n_1795;
wire n_1409;
wire n_1015;
wire n_663;
wire n_3448;
wire n_3634;
wire n_2744;
wire n_2101;
wire n_2795;
wire n_3524;
wire n_1377;
wire n_2473;
wire n_1583;
wire n_3520;
wire n_1521;
wire n_2632;
wire n_1152;
wire n_2456;
wire n_2924;
wire n_3054;
wire n_2264;
wire n_2076;
wire n_2599;
wire n_974;
wire n_1036;
wire n_1831;
wire n_3626;
wire n_864;
wire n_1987;
wire n_959;
wire n_1106;
wire n_1312;
wire n_1129;
wire n_1244;
wire n_3171;
wire n_1733;
wire n_3365;
wire n_3684;
wire n_1634;
wire n_2853;
wire n_1932;
wire n_1452;
wire n_1552;
wire n_1318;
wire n_1508;
wire n_2217;
wire n_738;
wire n_1217;
wire n_3594;
wire n_2866;
wire n_3153;
wire n_3291;
wire n_2655;
wire n_3487;
wire n_2454;
wire n_1715;
wire n_1189;
wire n_3300;
wire n_761;
wire n_748;
wire n_1713;
wire n_3621;
wire n_901;
wire n_1577;
wire n_2036;
wire n_1255;
wire n_2829;
wire n_2968;
wire n_2740;
wire n_3473;
wire n_1700;
wire n_2623;
wire n_2622;
wire n_3232;
wire n_2819;
wire n_1218;
wire n_2178;
wire n_1181;
wire n_3263;
wire n_1140;
wire n_1985;
wire n_1772;
wire n_2858;
wire n_3708;
wire n_1056;
wire n_2626;
wire n_1283;
wire n_3007;
wire n_1446;
wire n_2404;
wire n_1487;
wire n_3078;
wire n_2789;
wire n_2603;
wire n_840;
wire n_1203;
wire n_1421;
wire n_3640;
wire n_3218;
wire n_2821;
wire n_2573;
wire n_846;
wire n_1793;
wire n_1237;
wire n_2424;
wire n_2880;
wire n_2390;
wire n_2423;
wire n_859;
wire n_1109;
wire n_965;
wire n_2741;
wire n_2793;
wire n_3098;
wire n_3490;
wire n_3055;
wire n_1633;
wire n_3299;
wire n_2580;
wire n_3222;
wire n_1711;
wire n_3529;
wire n_3069;
wire n_3107;
wire n_3352;
wire n_3436;
wire n_1051;
wire n_1008;
wire n_3065;
wire n_2964;
wire n_2375;
wire n_1498;
wire n_2312;
wire n_2572;
wire n_2946;
wire n_1053;
wire n_1656;
wire n_1207;
wire n_1076;
wire n_1735;
wire n_2063;
wire n_1032;
wire n_936;
wire n_3082;
wire n_1884;
wire n_2176;
wire n_1825;
wire n_2805;
wire n_1589;
wire n_2717;
wire n_2204;
wire n_2863;
wire n_2575;
wire n_1210;
wire n_2319;
wire n_2877;
wire n_1933;
wire n_2522;
wire n_3357;
wire n_1996;
wire n_1510;
wire n_1201;
wire n_1842;
wire n_2852;
wire n_2132;
wire n_3110;
wire n_1246;
wire n_1677;
wire n_732;
wire n_1236;
wire n_3364;
wire n_832;
wire n_2297;
wire n_3429;
wire n_3306;
wire n_3412;
wire n_3037;
wire n_3188;
wire n_2780;
wire n_1792;
wire n_1712;
wire n_3250;
wire n_1984;
wire n_1568;
wire n_2885;
wire n_1877;
wire n_3445;
wire n_1184;
wire n_1477;
wire n_2080;
wire n_2220;
wire n_2585;
wire n_1724;
wire n_2554;
wire n_3155;
wire n_2838;
wire n_1364;
wire n_3183;
wire n_1540;
wire n_1676;
wire n_1013;
wire n_3243;
wire n_2468;
wire n_929;
wire n_3248;
wire n_3214;
wire n_637;
wire n_1136;
wire n_1890;
wire n_1075;
wire n_1249;
wire n_3128;
wire n_1918;
wire n_2606;
wire n_3642;
wire n_2549;
wire n_2461;
wire n_3468;
wire n_2006;
wire n_2440;
wire n_1229;
wire n_1440;
wire n_1490;
wire n_2152;
wire n_907;
wire n_1179;
wire n_1990;
wire n_3680;
wire n_1153;
wire n_3624;
wire n_1751;
wire n_669;
wire n_2787;
wire n_2467;
wire n_2146;
wire n_2341;
wire n_3525;
wire n_1737;
wire n_3145;
wire n_2779;
wire n_1117;
wire n_1273;
wire n_2547;
wire n_2930;
wire n_2616;
wire n_1748;
wire n_2662;
wire n_1083;
wire n_3205;
wire n_1014;
wire n_724;
wire n_2883;
wire n_938;
wire n_1178;
wire n_2935;
wire n_878;
wire n_2441;
wire n_3503;
wire n_2358;
wire n_2490;
wire n_3127;
wire n_3496;
wire n_2361;
wire n_1464;
wire n_1566;
wire n_3568;
wire n_944;
wire n_3312;
wire n_3003;
wire n_1848;
wire n_623;
wire n_2062;
wire n_2277;
wire n_2650;
wire n_1982;
wire n_2252;
wire n_2888;
wire n_2339;
wire n_3614;
wire n_1334;
wire n_1963;
wire n_3394;
wire n_1695;
wire n_1418;
wire n_2999;
wire n_2402;
wire n_1137;
wire n_2552;
wire n_2910;
wire n_3331;
wire n_660;
wire n_2590;
wire n_3119;
wire n_1977;
wire n_2294;
wire n_1200;
wire n_2295;
wire n_2530;
wire n_3345;
wire n_2379;
wire n_1120;
wire n_2300;
wire n_2792;
wire n_1602;
wire n_2965;
wire n_1776;
wire n_2372;
wire n_3341;
wire n_2382;
wire n_1852;
wire n_1522;
wire n_2523;
wire n_2557;
wire n_3544;
wire n_1279;
wire n_2505;
wire n_931;
wire n_3488;
wire n_827;
wire n_3554;
wire n_2481;
wire n_3692;
wire n_1064;
wire n_1408;
wire n_2832;
wire n_1028;
wire n_1264;
wire n_3535;
wire n_3730;
wire n_2808;
wire n_2287;
wire n_3597;
wire n_3396;
wire n_2954;
wire n_3526;
wire n_2102;
wire n_1935;
wire n_2046;
wire n_3367;
wire n_3492;
wire n_1146;
wire n_2785;
wire n_2751;
wire n_3558;
wire n_705;
wire n_2142;
wire n_1548;
wire n_3703;
wire n_2977;
wire n_1682;
wire n_1608;
wire n_3599;
wire n_1009;
wire n_1260;
wire n_1896;
wire n_1704;
wire n_2160;
wire n_2699;
wire n_2234;
wire n_2991;
wire n_847;
wire n_1436;
wire n_3239;
wire n_2303;
wire n_2600;
wire n_1069;
wire n_1485;
wire n_2239;
wire n_1465;
wire n_1352;
wire n_1171;
wire n_1126;
wire n_1232;
wire n_1979;
wire n_2328;
wire n_2715;
wire n_679;
wire n_1345;
wire n_2434;
wire n_696;
wire n_837;
wire n_1590;
wire n_2332;
wire n_640;
wire n_2971;
wire n_954;
wire n_3578;
wire n_1628;
wire n_725;
wire n_1773;
wire n_2133;
wire n_3553;
wire n_3072;
wire n_1545;
wire n_3249;
wire n_3580;
wire n_2369;
wire n_3470;
wire n_3584;
wire n_1471;
wire n_1738;
wire n_3441;
wire n_1115;
wire n_998;
wire n_1395;
wire n_1729;
wire n_2551;
wire n_3281;
wire n_801;
wire n_2823;
wire n_3274;
wire n_2613;
wire n_2094;
wire n_1479;
wire n_3505;
wire n_2306;
wire n_1046;
wire n_2419;
wire n_3397;
wire n_2934;
wire n_2807;
wire n_882;
wire n_942;
wire n_1627;
wire n_1431;
wire n_651;
wire n_721;
wire n_2525;
wire n_814;
wire n_1864;
wire n_943;
wire n_2568;
wire n_3087;
wire n_2629;
wire n_3587;
wire n_1086;
wire n_1523;
wire n_2197;
wire n_2010;
wire n_1756;
wire n_2097;
wire n_2733;
wire n_2241;
wire n_1470;
wire n_2109;
wire n_2098;
wire n_1761;
wire n_2648;
wire n_2458;
wire n_1836;
wire n_2398;
wire n_3032;
wire n_3401;
wire n_1593;
wire n_986;
wire n_1420;
wire n_2651;
wire n_1750;
wire n_1775;
wire n_2833;
wire n_1699;
wire n_3179;
wire n_927;
wire n_1563;
wire n_2905;
wire n_3460;
wire n_803;
wire n_2570;
wire n_3123;
wire n_1875;
wire n_3379;
wire n_1615;
wire n_2418;
wire n_2184;
wire n_1087;
wire n_3390;
wire n_3719;
wire n_757;
wire n_1400;
wire n_712;
wire n_1539;
wire n_1599;
wire n_1806;
wire n_2711;
wire n_3070;
wire n_2842;
wire n_3477;
wire n_650;
wire n_2635;
wire n_3646;
wire n_2469;
wire n_1575;
wire n_2209;
wire n_3074;
wire n_3020;
wire n_3142;
wire n_3164;
wire n_3475;
wire n_1448;
wire n_2077;
wire n_3136;
wire n_2520;
wire n_817;
wire n_2612;
wire n_2193;
wire n_3034;
wire n_2095;
wire n_3108;
wire n_2486;
wire n_2628;
wire n_2395;
wire n_951;
wire n_2521;
wire n_2908;
wire n_2053;
wire n_2752;
wire n_1580;
wire n_2124;
wire n_1574;
wire n_780;
wire n_2200;
wire n_1705;
wire n_3625;
wire n_633;
wire n_2304;
wire n_1746;
wire n_726;
wire n_1439;
wire n_2352;
wire n_2212;
wire n_2263;
wire n_2716;
wire n_3495;
wire n_863;
wire n_2185;
wire n_3169;
wire n_1832;
wire n_1128;
wire n_2476;
wire n_2376;
wire n_2979;
wire n_3398;
wire n_1266;
wire n_1300;
wire n_2781;
wire n_3419;
wire n_3629;
wire n_807;
wire n_741;
wire n_2460;
wire n_2170;
wire n_3600;
wire n_1785;
wire n_1870;
wire n_2484;
wire n_2721;
wire n_1405;
wire n_2884;
wire n_3383;
wire n_3167;
wire n_3687;
wire n_997;
wire n_2308;
wire n_3459;
wire n_3238;
wire n_2986;
wire n_3498;
wire n_1428;
wire n_2691;
wire n_2243;
wire n_2400;
wire n_3092;
wire n_3555;
wire n_2903;
wire n_891;
wire n_3659;
wire n_3254;
wire n_2507;
wire n_2759;
wire n_3434;
wire n_1528;
wire n_1495;
wire n_3131;
wire n_3682;
wire n_2463;
wire n_2654;
wire n_717;
wire n_2975;
wire n_1357;
wire n_2503;
wire n_2478;
wire n_3178;
wire n_2794;
wire n_1512;
wire n_3672;
wire n_2496;
wire n_3378;
wire n_3481;
wire n_668;
wire n_2974;
wire n_871;
wire n_2990;
wire n_2923;
wire n_1339;
wire n_1544;
wire n_1426;
wire n_2365;
wire n_3449;
wire n_3517;
wire n_3350;
wire n_2245;
wire n_1315;
wire n_1413;
wire n_2464;
wire n_811;
wire n_808;
wire n_945;
wire n_2925;
wire n_2270;
wire n_3260;
wire n_1706;
wire n_1560;
wire n_1592;
wire n_2776;
wire n_1461;
wire n_3166;
wire n_2695;
wire n_2630;
wire n_903;
wire n_1967;
wire n_2340;
wire n_3385;
wire n_2117;
wire n_1095;
wire n_1328;
wire n_1265;
wire n_2488;
wire n_1378;
wire n_2042;
wire n_3656;
wire n_3257;
wire n_1048;
wire n_774;
wire n_2459;
wire n_3137;
wire n_3116;
wire n_1925;
wire n_2439;
wire n_3638;
wire n_2106;
wire n_1430;
wire n_2414;
wire n_1251;
wire n_3090;
wire n_1247;
wire n_2450;
wire n_836;
wire n_1475;
wire n_3316;
wire n_2465;
wire n_1263;
wire n_3337;
wire n_1683;
wire n_1185;
wire n_3575;
wire n_1122;
wire n_2765;
wire n_3387;
wire n_890;
wire n_628;
wire n_874;
wire n_1505;
wire n_3010;
wire n_2941;
wire n_1163;
wire n_677;
wire n_1514;
wire n_964;
wire n_2728;
wire n_2948;
wire n_916;
wire n_3428;
wire n_2298;
wire n_2771;
wire n_3219;
wire n_2936;
wire n_895;
wire n_687;
wire n_1035;
wire n_2427;
wire n_2045;
wire n_2985;
wire n_1535;
wire n_3158;
wire n_3106;
wire n_751;
wire n_2190;
wire n_1127;
wire n_932;
wire n_3657;
wire n_1972;
wire n_3080;
wire n_2772;
wire n_2778;
wire n_947;
wire n_1004;
wire n_831;
wire n_778;
wire n_1898;
wire n_1254;
wire n_1148;
wire n_1667;
wire n_1104;
wire n_1845;
wire n_1011;
wire n_2205;
wire n_2684;
wire n_2875;
wire n_2524;
wire n_3284;
wire n_1437;
wire n_3723;
wire n_2747;
wire n_3389;
wire n_626;
wire n_1707;
wire n_1941;
wire n_2422;
wire n_2064;
wire n_3088;
wire n_1679;
wire n_2342;
wire n_2755;
wire n_2301;
wire n_1497;
wire n_2002;
wire n_2055;
wire n_3564;
wire n_2385;
wire n_3095;
wire n_3026;
wire n_2545;
wire n_1578;
wire n_3294;
wire n_2050;
wire n_1143;
wire n_1783;
wire n_2712;
wire n_3695;
wire n_3279;
wire n_2584;
wire n_972;
wire n_1815;
wire n_2500;
wire n_3344;
wire n_1917;
wire n_1444;
wire n_920;
wire n_664;
wire n_2442;
wire n_1067;
wire n_3328;
wire n_2763;
wire n_2788;
wire n_994;
wire n_2000;
wire n_2089;
wire n_1857;
wire n_2761;
wire n_1920;
wire n_2696;
wire n_3252;
wire n_887;
wire n_1162;
wire n_1997;
wire n_2578;
wire n_2745;
wire n_1894;
wire n_2110;
wire n_2904;
wire n_2896;
wire n_3064;
wire n_2997;
wire n_3314;
wire n_634;
wire n_961;
wire n_991;
wire n_1223;
wire n_1349;
wire n_1331;
wire n_2127;
wire n_1323;
wire n_1739;
wire n_3130;
wire n_1777;
wire n_3028;
wire n_3228;
wire n_3710;
wire n_1353;
wire n_3409;
wire n_2386;
wire n_3706;
wire n_3324;
wire n_1429;
wire n_3073;
wire n_2029;
wire n_3209;
wire n_2026;
wire n_1546;
wire n_3588;
wire n_3420;
wire n_1432;
wire n_2103;
wire n_3322;
wire n_1950;
wire n_1320;
wire n_996;
wire n_3632;
wire n_915;
wire n_2238;
wire n_3289;
wire n_1174;
wire n_1834;
wire n_1874;
wire n_3372;
wire n_3499;
wire n_3552;
wire n_2862;
wire n_3100;
wire n_3405;
wire n_1727;
wire n_3377;
wire n_1286;
wire n_1657;
wire n_1741;
wire n_1294;
wire n_1601;
wire n_900;
wire n_3414;
wire n_1351;
wire n_2933;
wire n_2138;
wire n_647;
wire n_1380;
wire n_1367;
wire n_3336;
wire n_3240;
wire n_1291;
wire n_2895;
wire n_1914;
wire n_1458;
wire n_1694;
wire n_1460;
wire n_2041;
wire n_3201;
wire n_2271;
wire n_2356;
wire n_3339;
wire n_1830;
wire n_2261;
wire n_3016;
wire n_1629;
wire n_3476;
wire n_3673;
wire n_2994;
wire n_2011;
wire n_2620;
wire n_1826;
wire n_1855;
wire n_1662;
wire n_2105;
wire n_2187;
wire n_3556;
wire n_1340;
wire n_2694;
wire n_3443;
wire n_2562;
wire n_2642;
wire n_3029;
wire n_3269;
wire n_3609;
wire n_3447;
wire n_2647;
wire n_1626;
wire n_674;
wire n_2223;
wire n_1660;
wire n_1850;
wire n_1643;
wire n_1670;
wire n_1789;
wire n_2415;
wire n_3152;
wire n_3154;
wire n_2344;
wire n_3589;
wire n_2317;
wire n_2556;
wire n_1112;
wire n_1267;
wire n_2384;
wire n_2683;
wire n_1384;
wire n_1376;
wire n_1537;
wire n_1858;
wire n_3432;
wire n_3523;
wire n_2815;
wire n_1816;
wire n_2446;
wire n_3388;
wire n_1612;
wire n_703;
wire n_2318;
wire n_1172;
wire n_2659;
wire n_3616;
wire n_1099;
wire n_2141;
wire n_3113;
wire n_3696;
wire n_2902;
wire n_2909;
wire n_1422;
wire n_1527;
wire n_3174;
wire n_3608;
wire n_3190;
wire n_1055;
wire n_1524;
wire n_673;
wire n_798;
wire n_2849;
wire n_2947;
wire n_1754;
wire n_3048;
wire n_3686;
wire n_1177;
wire n_1025;
wire n_1991;
wire n_2566;
wire n_2679;
wire n_3292;
wire n_2210;
wire n_1517;
wire n_690;
wire n_2502;
wire n_1225;
wire n_1962;
wire n_2346;
wire n_982;
wire n_3670;
wire n_1624;
wire n_785;
wire n_1952;
wire n_2180;
wire n_3002;
wire n_3376;
wire n_2087;
wire n_2920;
wire n_3290;
wire n_1598;
wire n_2952;
wire n_2617;
wire n_3585;
wire n_977;
wire n_2878;
wire n_1895;
wire n_2250;
wire n_719;
wire n_1491;
wire n_1860;
wire n_2831;
wire n_716;
wire n_1810;
wire n_1763;
wire n_923;
wire n_642;
wire n_1607;
wire n_2865;
wire n_2075;
wire n_3047;
wire n_1625;
wire n_2959;
wire n_2610;
wire n_2420;
wire n_2380;
wire n_3335;
wire n_3265;
wire n_2240;
wire n_933;
wire n_2221;
wire n_1774;
wire n_1797;
wire n_2516;
wire n_2120;
wire n_1037;
wire n_1899;
wire n_2031;
wire n_3669;
wire n_3427;
wire n_1289;
wire n_838;
wire n_1348;
wire n_2892;
wire n_1021;
wire n_746;
wire n_1557;
wire n_1188;
wire n_1567;
wire n_2007;
wire n_742;
wire n_1191;
wire n_2004;
wire n_3356;
wire n_3431;
wire n_3220;
wire n_2024;
wire n_2086;
wire n_1503;
wire n_3422;
wire n_1052;
wire n_789;
wire n_1942;
wire n_656;
wire n_3666;
wire n_3141;
wire n_2309;
wire n_842;
wire n_2274;
wire n_2698;
wire n_767;
wire n_1617;
wire n_1839;
wire n_1587;
wire n_2330;
wire n_2555;
wire n_2639;
wire n_636;
wire n_1259;
wire n_2108;
wire n_3099;
wire n_3712;
wire n_2535;
wire n_1001;
wire n_2945;
wire n_3057;
wire n_2143;
wire n_2410;
wire n_1396;
wire n_2916;
wire n_1224;
wire n_1923;
wire n_3206;
wire n_2196;
wire n_2739;
wire n_2611;
wire n_1538;
wire n_2528;
wire n_2548;
wire n_3216;
wire n_2709;
wire n_3061;
wire n_3717;
wire n_2633;
wire n_1017;
wire n_2244;
wire n_730;
wire n_2604;
wire n_3462;
wire n_3424;
wire n_2351;
wire n_2437;
wire n_3664;
wire n_2049;
wire n_1456;
wire n_3245;
wire n_1889;
wire n_625;
wire n_2113;
wire n_2665;
wire n_1124;
wire n_1690;
wire n_3063;
wire n_2688;
wire n_2881;
wire n_3302;
wire n_1673;
wire n_3361;
wire n_2018;
wire n_3134;
wire n_922;
wire n_2817;
wire n_1790;
wire n_851;
wire n_993;
wire n_3196;
wire n_2085;
wire n_3304;
wire n_2581;
wire n_1725;
wire n_2809;
wire n_2149;
wire n_2237;
wire n_2320;
wire n_2268;
wire n_1135;
wire n_2255;
wire n_2001;
wire n_1820;
wire n_1800;
wire n_3277;
wire n_3480;
wire n_2758;
wire n_659;
wire n_1494;
wire n_1550;
wire n_2060;
wire n_1066;
wire n_2214;
wire n_3474;
wire n_648;
wire n_1169;
wire n_1726;
wire n_1946;
wire n_3111;
wire n_1938;
wire n_830;
wire n_3452;
wire n_1241;
wire n_3645;
wire n_2589;
wire n_1072;
wire n_2194;
wire n_1231;
wire n_1173;
wire n_2736;
wire n_1208;
wire n_1639;
wire n_1604;
wire n_2735;
wire n_2845;
wire n_3506;
wire n_826;
wire n_2154;
wire n_1976;
wire n_2035;
wire n_1337;
wire n_2984;
wire n_3162;
wire n_2732;
wire n_1906;
wire n_3004;
wire n_1647;
wire n_1901;
wire n_3096;
wire n_3333;
wire n_768;
wire n_839;
wire n_3705;
wire n_3031;
wire n_1278;
wire n_2059;
wire n_796;
wire n_797;
wire n_3276;
wire n_1006;
wire n_2956;
wire n_1238;
wire n_1415;
wire n_976;
wire n_1710;
wire n_3021;
wire n_1063;
wire n_2153;
wire n_2452;
wire n_1270;
wire n_2891;
wire n_834;
wire n_2457;
wire n_2144;
wire n_1476;
wire n_935;
wire n_1603;
wire n_925;
wire n_2592;
wire n_1054;
wire n_2027;
wire n_3404;
wire n_2072;
wire n_2737;
wire n_2012;
wire n_722;
wire n_2251;
wire n_2963;
wire n_3512;
wire n_1644;
wire n_1406;
wire n_1489;
wire n_3591;
wire n_1880;
wire n_1993;
wire n_2137;
wire n_804;
wire n_1642;
wire n_1455;
wire n_1871;
wire n_2182;
wire n_3044;
wire n_2868;
wire n_2447;
wire n_3493;
wire n_2818;
wire n_3358;
wire n_3115;
wire n_1057;
wire n_1473;
wire n_3140;
wire n_3486;
wire n_2125;
wire n_2426;
wire n_2894;
wire n_1403;
wire n_3253;
wire n_2181;
wire n_2587;
wire n_1149;
wire n_1176;
wire n_1502;
wire n_1605;
wire n_868;
wire n_2099;
wire n_1202;
wire n_1065;
wire n_1897;
wire n_2477;
wire n_1457;
wire n_3172;
wire n_905;
wire n_2159;
wire n_3410;
wire n_975;
wire n_675;
wire n_624;
wire n_934;
wire n_775;
wire n_3273;
wire n_950;
wire n_2700;
wire n_685;
wire n_1222;
wire n_3139;
wire n_1630;
wire n_3408;
wire n_2286;
wire n_3182;
wire n_1879;
wire n_1959;
wire n_2563;
wire n_1198;
wire n_2206;
wire n_3637;
wire n_1311;
wire n_3393;
wire n_1261;
wire n_2299;
wire n_3538;
wire n_2078;
wire n_3650;
wire n_3327;
wire n_2265;
wire n_776;
wire n_1114;
wire n_3513;
wire n_3709;
wire n_3011;
wire n_1167;
wire n_818;
wire n_3231;
wire n_2677;
wire n_2531;
wire n_2315;
wire n_3623;
wire n_3647;
wire n_3138;
wire n_2157;
wire n_3212;
wire n_1282;
wire n_2067;
wire n_2517;
wire n_1321;
wire n_700;
wire n_1779;
wire n_3446;
wire n_3349;
wire n_3619;
wire n_2489;
wire n_1770;
wire n_1107;
wire n_3058;
wire n_3454;
wire n_1846;
wire n_2211;
wire n_1573;
wire n_2950;
wire n_815;
wire n_919;
wire n_2272;
wire n_1956;
wire n_3574;
wire n_681;
wire n_2608;
wire n_3384;
wire n_2983;
wire n_1718;
wire n_2225;
wire n_3229;
wire n_2546;
wire n_1411;
wire n_2825;
wire n_1139;
wire n_1018;
wire n_858;
wire n_2345;
wire n_1324;
wire n_1669;
wire n_1501;
wire n_2742;
wire n_782;
wire n_1885;
wire n_1740;
wire n_1989;
wire n_3540;
wire n_1838;
wire n_3604;
wire n_833;
wire n_3649;
wire n_2680;
wire n_1343;
wire n_1801;
wire n_3439;
wire n_1371;
wire n_1513;
wire n_728;
wire n_3001;
wire n_2861;
wire n_2976;
wire n_2161;
wire n_2191;
wire n_3611;
wire n_2329;
wire n_1788;
wire n_2348;
wire n_2093;
wire n_786;
wire n_2576;
wire n_2417;
wire n_2675;
wire n_2043;
wire n_3601;
wire n_2366;
wire n_1621;
wire n_2338;
wire n_3571;
wire n_1919;
wire n_1342;
wire n_752;
wire n_2756;
wire n_2893;
wire n_2009;
wire n_2248;
wire n_958;
wire n_1175;
wire n_3500;
wire n_1416;
wire n_1659;
wire n_2850;
wire n_3465;
wire n_1221;
wire n_1047;
wire n_1878;
wire n_1515;
wire n_1374;
wire n_2851;
wire n_2438;
wire n_1435;
wire n_1688;
wire n_792;
wire n_2973;
wire n_3651;
wire n_1314;
wire n_1433;
wire n_2567;
wire n_3059;
wire n_3085;
wire n_1242;
wire n_1119;
wire n_2229;
wire n_2810;
wire n_2867;
wire n_1085;
wire n_3027;
wire n_2388;
wire n_2981;
wire n_3438;
wire n_2222;
wire n_3112;
wire n_1907;
wire n_3464;
wire n_885;
wire n_1530;
wire n_3215;
wire n_3413;
wire n_877;
wire n_2871;
wire n_2135;
wire n_1088;
wire n_896;
wire n_2764;
wire n_2624;
wire n_1813;
wire n_1451;
wire n_1005;
wire n_1102;
wire n_3234;
wire n_631;
wire n_794;
wire n_3648;
wire n_2471;
wire n_1288;
wire n_1275;
wire n_985;
wire n_1165;
wire n_897;
wire n_1622;
wire n_2757;
wire n_2714;
wire n_3066;
wire n_2669;
wire n_697;
wire n_2869;
wire n_1105;
wire n_1459;
wire n_912;
wire n_2898;
wire n_2232;
wire n_3121;
wire n_2455;
wire n_2121;
wire n_1893;
wire n_2519;
wire n_1570;
wire n_2231;
wire n_2874;
wire n_701;
wire n_995;
wire n_2278;
wire n_1000;
wire n_2284;
wire n_2433;
wire n_2816;
wire n_2803;
wire n_1931;
wire n_3402;
wire n_1256;
wire n_2798;
wire n_3425;
wire n_1303;
wire n_1994;
wire n_1771;
wire n_3308;
wire n_1526;
wire n_764;
wire n_1507;
wire n_1206;
wire n_1809;
wire n_855;
wire n_2367;
wire n_812;
wire n_2658;
wire n_3236;
wire n_3491;
wire n_3109;
wire n_1961;
wire n_3576;
wire n_3271;
wire n_3013;
wire n_2553;
wire n_1050;
wire n_2218;
wire n_2667;
wire n_3062;
wire n_1769;
wire n_2130;
wire n_3256;
wire n_1060;
wire n_3126;
wire n_1372;
wire n_1847;
wire n_756;
wire n_1565;
wire n_1257;
wire n_2325;
wire n_2406;
wire n_1632;
wire n_2864;
wire n_3346;
wire n_688;
wire n_3104;
wire n_3391;
wire n_1542;
wire n_946;
wire n_1586;
wire n_707;
wire n_1362;
wire n_1547;
wire n_3497;
wire n_1097;
wire n_3354;
wire n_3288;
wire n_3373;
wire n_3382;
wire n_3122;
wire n_2518;
wire n_2784;
wire n_3012;
wire n_3045;
wire n_1909;
wire n_2543;
wire n_3368;
wire n_2381;
wire n_2313;
wire n_3561;
wire n_956;
wire n_3586;
wire n_790;
wire n_2495;
wire n_2992;
wire n_1541;
wire n_2703;
wire n_1812;
wire n_3014;
wire n_1951;
wire n_1330;
wire n_638;
wire n_2574;
wire n_1697;
wire n_2128;
wire n_1872;
wire n_1940;
wire n_2690;
wire n_1747;
wire n_1212;
wire n_1887;
wire n_1199;
wire n_3400;
wire n_2020;
wire n_3504;
wire n_1978;
wire n_2508;
wire n_3511;
wire n_2540;
wire n_1767;
wire n_1939;
wire n_2428;
wire n_3159;
wire n_1768;
wire n_1443;
wire n_3697;
wire n_2068;
wire n_2636;
wire n_2672;
wire n_3360;
wire n_1585;
wire n_1861;
wire n_2316;
wire n_3101;
wire n_1564;
wire n_1995;
wire n_1631;
wire n_2593;
wire n_2911;
wire n_1623;
wire n_861;
wire n_1828;
wire n_2364;
wire n_1389;
wire n_3303;
wire n_1131;
wire n_2641;
wire n_1798;
wire n_727;
wire n_1077;
wire n_3120;
wire n_1554;
wire n_3549;
wire n_1584;
wire n_1481;
wire n_2021;
wire n_1928;
wire n_2713;
wire n_828;
wire n_2938;
wire n_3227;
wire n_1438;
wire n_3342;
wire n_1973;
wire n_2314;
wire n_2939;
wire n_2156;
wire n_2494;
wire n_753;
wire n_2126;
wire n_645;
wire n_1147;
wire n_747;
wire n_3403;
wire n_1363;
wire n_2228;
wire n_1691;
wire n_1098;
wire n_1366;
wire n_1518;
wire n_1187;
wire n_1361;
wire n_2034;
wire n_1693;
wire n_698;
wire n_2790;
wire n_3173;
wire n_2872;
wire n_3102;
wire n_2411;
wire n_2081;
wire n_1892;
wire n_1061;
wire n_3539;
wire n_2266;
wire n_2993;
wire n_682;
wire n_3433;
wire n_2061;
wire n_3018;
wire n_1373;
wire n_2449;
wire n_1686;
wire n_2131;
wire n_2526;
wire n_2830;
wire n_1302;
wire n_3017;
wire n_3083;
wire n_2083;
wire n_886;
wire n_2119;
wire n_1010;
wire n_883;
wire n_2207;
wire n_2044;
wire n_2542;
wire n_755;
wire n_2091;
wire n_2843;
wire n_3362;
wire n_3035;
wire n_3191;
wire n_1029;
wire n_3485;
wire n_2394;
wire n_3051;
wire n_770;
wire n_1572;
wire n_1635;
wire n_3305;
wire n_3149;
wire n_2827;
wire n_941;
wire n_1245;
wire n_1317;
wire n_3643;
wire n_2615;
wire n_3278;
wire n_2487;
wire n_2701;
wire n_2929;
wire n_3163;
wire n_3343;
wire n_632;
wire n_1329;
wire n_2409;
wire n_2637;
wire n_2337;
wire n_854;
wire n_2405;
wire n_2601;
wire n_2513;
wire n_3118;
wire n_1369;
wire n_714;
wire n_1297;
wire n_1912;
wire n_3143;
wire n_1734;
wire n_3543;
wire n_3655;
wire n_1876;
wire n_2666;
wire n_3050;
wire n_2323;
wire n_3532;
wire n_740;
wire n_1811;
wire n_898;
wire n_928;
wire n_1285;
wire n_3042;
wire n_967;
wire n_2561;
wire n_736;
wire n_3725;
wire n_2913;
wire n_2491;
wire n_1529;
wire n_1381;
wire n_1824;
wire n_2254;
wire n_1597;
wire n_1161;
wire n_1103;
wire n_3522;
wire n_1486;
wire n_1068;
wire n_1833;
wire n_2914;
wire n_3551;
wire n_2371;
wire n_914;
wire n_3444;
wire n_1986;
wire n_3366;
wire n_2882;
wire n_1024;
wire n_3009;
wire n_1141;
wire n_3453;
wire n_3297;
wire n_3176;
wire n_1949;
wire n_1197;
wire n_2493;
wire n_2408;
wire n_2429;
wire n_3326;
wire n_1168;
wire n_865;
wire n_3581;
wire n_3000;
wire n_2115;
wire n_2013;
wire n_2140;
wire n_2134;
wire n_2483;
wire n_2305;
wire n_1556;
wire n_3423;
wire n_3547;
wire n_1192;
wire n_1646;
wire n_1290;
wire n_3700;
wire n_2514;
wire n_2466;
wire n_3661;
wire n_1759;
wire n_2048;
wire n_2760;
wire n_987;
wire n_750;
wire n_1299;
wire n_2942;
wire n_2096;
wire n_3663;
wire n_2129;
wire n_3230;
wire n_665;
wire n_3545;
wire n_1101;
wire n_2532;
wire n_3665;
wire n_2079;
wire n_2296;
wire n_1720;
wire n_880;
wire n_654;
wire n_2671;
wire n_1911;
wire n_2293;
wire n_3296;
wire n_731;
wire n_1336;
wire n_3068;
wire n_3071;
wire n_3683;
wire n_2734;
wire n_2870;
wire n_1166;
wire n_758;
wire n_710;
wire n_720;
wire n_1390;
wire n_2775;
wire n_1023;
wire n_1358;
wire n_813;
wire n_2310;
wire n_3318;
wire n_3223;
wire n_1397;
wire n_1211;
wire n_2674;
wire n_1284;
wire n_2005;
wire n_1359;
wire n_1116;
wire n_2811;
wire n_1758;
wire n_3226;
wire n_3702;
wire n_791;
wire n_1532;
wire n_2848;
wire n_1419;
wire n_2689;
wire n_1784;
wire n_1685;
wire n_1992;
wire n_1082;
wire n_3200;
wire n_3430;
wire n_1213;
wire n_2596;
wire n_2801;
wire n_980;
wire n_1193;
wire n_849;
wire n_1488;
wire n_2928;
wire n_3067;
wire n_2227;
wire n_2652;
wire n_3225;
wire n_1074;
wire n_3380;
wire n_3557;
wire n_3207;
wire n_3596;
wire n_759;
wire n_1379;
wire n_1721;
wire n_2972;
wire n_2627;
wire n_1827;
wire n_953;
wire n_1180;
wire n_1462;
wire n_3606;
wire n_3369;
wire n_3185;
wire n_2326;
wire n_1866;
wire n_1220;
wire n_1398;
wire n_2111;
wire n_2169;
wire n_1262;
wire n_1904;
wire n_2966;
wire n_3084;
wire n_3036;
wire n_1692;
wire n_2501;
wire n_2051;
wire n_1012;
wire n_1805;
wire n_960;
wire n_689;
wire n_1022;
wire n_1760;
wire n_676;
wire n_1240;
wire n_2173;
wire n_1183;
wire n_3285;
wire n_3160;
wire n_3483;
wire n_1204;
wire n_1151;
wire n_2824;
wire n_1814;
wire n_771;
wire n_2982;
wire n_999;
wire n_2634;
wire n_3124;
wire n_3286;
wire n_1092;
wire n_1808;
wire n_2768;
wire n_2668;
wire n_1658;
wire n_1386;
wire n_3015;
wire n_2588;
wire n_2931;
wire n_3321;
wire n_2492;
wire n_3081;
wire n_3636;
wire n_910;
wire n_2291;
wire n_635;
wire n_3612;
wire n_3046;
wire n_844;
wire n_2172;
wire n_1728;
wire n_1020;
wire n_3076;
wire n_783;
wire n_1385;
wire n_1142;
wire n_2927;
wire n_1062;
wire n_1230;
wire n_1027;
wire n_1516;
wire n_3622;
wire n_2533;
wire n_1499;
wire n_1500;
wire n_2155;
wire n_2706;
wire n_1868;
wire n_966;
wire n_2148;
wire n_2104;
wire n_949;
wire n_704;
wire n_2653;
wire n_2618;
wire n_2357;
wire n_2855;
wire n_924;
wire n_2937;
wire n_3728;
wire n_3359;
wire n_3114;
wire n_2331;
wire n_3332;
wire n_1600;
wire n_1661;
wire n_2967;
wire n_1965;
wire n_3005;
wire n_1757;
wire n_699;
wire n_2136;
wire n_3617;
wire n_3602;
wire n_2403;
wire n_918;
wire n_3053;
wire n_2056;
wire n_1913;
wire n_672;
wire n_2702;
wire n_2054;
wire n_1039;
wire n_2226;
wire n_2407;
wire n_2791;
wire n_1043;
wire n_1402;
wire n_2267;
wire n_735;
wire n_1450;
wire n_2082;
wire n_2302;
wire n_2453;
wire n_3056;
wire n_2560;
wire n_3267;
wire n_2092;
wire n_3008;
wire n_1365;
wire n_1472;
wire n_2443;
wire n_2802;
wire n_3052;
wire n_3189;
wire n_2797;
wire n_2279;
wire n_1089;
wire n_1536;
wire n_1049;
wire n_1719;
wire n_1974;
wire n_1158;
wire n_2066;
wire n_2988;
wire n_763;
wire n_1882;
wire n_2770;
wire n_2961;
wire n_2704;
wire n_2996;
wire n_1915;
wire n_2836;
wire n_940;
wire n_1762;
wire n_2534;
wire n_1404;
wire n_3582;
wire n_3689;
wire n_788;
wire n_3283;
wire n_1736;
wire n_3421;
wire n_2907;
wire n_3311;
wire n_1160;
wire n_1442;
wire n_658;
wire n_1948;
wire n_2168;
wire n_1216;
wire n_2681;
wire n_1891;
wire n_1026;
wire n_3247;
wire n_2886;
wire n_1454;
wire n_1033;
wire n_3613;
wire n_627;
wire n_990;
wire n_1383;
wire n_3675;
wire n_1968;
wire n_2057;
wire n_2609;
wire n_2378;
wire n_888;
wire n_2749;
wire n_3658;
wire n_1325;
wire n_3133;
wire n_2754;
wire n_3527;
wire n_2014;
wire n_3041;
wire n_1483;
wire n_1703;
wire n_653;
wire n_1205;
wire n_1822;
wire n_843;
wire n_1953;
wire n_3715;
wire n_1059;
wire n_2969;
wire n_799;
wire n_3713;
wire n_2692;
wire n_3261;
wire n_3550;
wire n_691;
wire n_1804;
wire n_1581;
wire n_3287;
wire n_3534;
wire n_1837;
wire n_3325;
wire n_1744;
wire n_1975;
wire n_3437;
wire n_1414;
wire n_2246;
wire n_2738;
wire n_2324;
wire n_3161;
wire n_1002;
wire n_1851;
wire n_1755;
wire n_2195;
wire n_2940;
wire n_1111;
wire n_1819;
wire n_3313;
wire n_1341;
wire n_1807;
wire n_2670;
wire n_2645;
wire n_2202;
wire n_1310;
wire n_3275;
wire n_1745;
wire n_1714;
wire n_3198;
wire n_3463;
wire n_1958;
wire n_1611;
wire n_2559;
wire n_3516;
wire n_2262;
wire n_3562;
wire n_955;
wire n_1333;
wire n_1916;
wire n_2619;
wire n_2917;
wire n_2726;
wire n_2073;
wire n_952;
wire n_1675;
wire n_1947;
wire n_2165;
wire n_1640;
wire n_2016;
wire n_3157;
wire n_1551;
wire n_1145;
wire n_1533;
wire n_2307;
wire n_2515;
wire n_3546;
wire n_1511;
wire n_1791;
wire n_1113;
wire n_3089;
wire n_1651;
wire n_1966;
wire n_2058;
wire n_2678;
wire n_3406;
wire n_1468;
wire n_3442;
wire n_2327;
wire n_2656;
wire n_913;
wire n_2353;
wire n_1164;
wire n_2258;
wire n_3662;
wire n_3595;
wire n_1732;
wire n_2167;
wire n_3079;
wire n_1354;
wire n_3329;
wire n_2039;
wire n_1277;
wire n_1696;
wire n_1016;
wire n_3233;
wire n_680;
wire n_1355;
wire n_809;
wire n_3691;
wire n_2544;
wire n_856;
wire n_779;
wire n_3193;
wire n_3501;
wire n_3635;
wire n_866;
wire n_2538;
wire n_3270;
wire n_2582;
wire n_1559;
wire n_2321;
wire n_2915;
wire n_1579;
wire n_1280;
wire n_2854;
wire n_2932;
wire n_3258;
wire n_1335;
wire n_3266;
wire n_2285;
wire n_3213;
wire n_1934;
wire n_1900;
wire n_2040;
wire n_2174;
wire n_3246;
wire n_1843;
wire n_2186;
wire n_2510;
wire n_2030;
wire n_2614;
wire n_3418;
wire n_2435;
wire n_1665;
wire n_2583;
wire n_3417;
wire n_1091;
wire n_1678;
wire n_1780;
wire n_2725;
wire n_1287;
wire n_2769;
wire n_1482;
wire n_860;
wire n_1525;
wire n_661;
wire n_848;
wire n_3244;
wire n_3195;
wire n_3593;
wire n_2100;
wire n_2349;
wire n_1902;
wire n_2536;
wire n_2474;
wire n_683;
wire n_1150;
wire n_1194;
wire n_1399;
wire n_3685;
wire n_1903;
wire n_1674;
wire n_1849;
wire n_686;
wire n_867;
wire n_983;
wire n_1417;
wire n_644;
wire n_3482;
wire n_2282;
wire n_970;
wire n_3654;
wire n_2430;
wire n_2673;
wire n_921;
wire n_2676;
wire n_3515;
wire n_3489;
wire n_2926;
wire n_1534;
wire n_2912;
wire n_3181;
wire n_908;
wire n_3536;
wire n_1346;
wire n_2834;
wire n_3644;
wire n_3268;
wire n_1123;
wire n_2710;
wire n_1272;
wire n_2497;
wire n_1393;
wire n_2970;
wire n_984;
wire n_1655;
wire n_3040;
wire n_3494;
wire n_2978;
wire n_3615;
wire n_1410;
wire n_988;
wire n_2368;
wire n_3363;
wire n_760;
wire n_3528;
wire n_1157;
wire n_3502;
wire n_806;
wire n_3677;
wire n_2657;
wire n_1186;
wire n_2065;
wire n_2901;
wire n_3180;
wire n_1743;
wire n_2743;
wire n_649;
wire n_1854;
wire n_1506;

CKINVDCx5p33_ASAP7_75t_R g622 ( 
.A(n_580),
.Y(n_622)
);

CKINVDCx5p33_ASAP7_75t_R g623 ( 
.A(n_202),
.Y(n_623)
);

CKINVDCx5p33_ASAP7_75t_R g624 ( 
.A(n_280),
.Y(n_624)
);

BUFx6f_ASAP7_75t_L g625 ( 
.A(n_379),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_564),
.Y(n_626)
);

BUFx2_ASAP7_75t_L g627 ( 
.A(n_527),
.Y(n_627)
);

CKINVDCx5p33_ASAP7_75t_R g628 ( 
.A(n_63),
.Y(n_628)
);

CKINVDCx5p33_ASAP7_75t_R g629 ( 
.A(n_410),
.Y(n_629)
);

CKINVDCx14_ASAP7_75t_R g630 ( 
.A(n_539),
.Y(n_630)
);

CKINVDCx20_ASAP7_75t_R g631 ( 
.A(n_430),
.Y(n_631)
);

CKINVDCx5p33_ASAP7_75t_R g632 ( 
.A(n_535),
.Y(n_632)
);

CKINVDCx5p33_ASAP7_75t_R g633 ( 
.A(n_281),
.Y(n_633)
);

CKINVDCx5p33_ASAP7_75t_R g634 ( 
.A(n_181),
.Y(n_634)
);

CKINVDCx5p33_ASAP7_75t_R g635 ( 
.A(n_415),
.Y(n_635)
);

BUFx10_ASAP7_75t_L g636 ( 
.A(n_416),
.Y(n_636)
);

INVx1_ASAP7_75t_SL g637 ( 
.A(n_96),
.Y(n_637)
);

INVx1_ASAP7_75t_SL g638 ( 
.A(n_101),
.Y(n_638)
);

CKINVDCx5p33_ASAP7_75t_R g639 ( 
.A(n_614),
.Y(n_639)
);

CKINVDCx20_ASAP7_75t_R g640 ( 
.A(n_524),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_69),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_588),
.Y(n_642)
);

CKINVDCx5p33_ASAP7_75t_R g643 ( 
.A(n_226),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_142),
.Y(n_644)
);

INVxp67_ASAP7_75t_L g645 ( 
.A(n_5),
.Y(n_645)
);

BUFx10_ASAP7_75t_L g646 ( 
.A(n_258),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_593),
.Y(n_647)
);

CKINVDCx20_ASAP7_75t_R g648 ( 
.A(n_102),
.Y(n_648)
);

CKINVDCx5p33_ASAP7_75t_R g649 ( 
.A(n_401),
.Y(n_649)
);

CKINVDCx5p33_ASAP7_75t_R g650 ( 
.A(n_442),
.Y(n_650)
);

CKINVDCx5p33_ASAP7_75t_R g651 ( 
.A(n_382),
.Y(n_651)
);

CKINVDCx5p33_ASAP7_75t_R g652 ( 
.A(n_452),
.Y(n_652)
);

CKINVDCx5p33_ASAP7_75t_R g653 ( 
.A(n_230),
.Y(n_653)
);

BUFx2_ASAP7_75t_L g654 ( 
.A(n_380),
.Y(n_654)
);

CKINVDCx5p33_ASAP7_75t_R g655 ( 
.A(n_506),
.Y(n_655)
);

INVx2_ASAP7_75t_L g656 ( 
.A(n_165),
.Y(n_656)
);

CKINVDCx5p33_ASAP7_75t_R g657 ( 
.A(n_522),
.Y(n_657)
);

INVx2_ASAP7_75t_L g658 ( 
.A(n_81),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_152),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_204),
.Y(n_660)
);

HB1xp67_ASAP7_75t_L g661 ( 
.A(n_328),
.Y(n_661)
);

CKINVDCx5p33_ASAP7_75t_R g662 ( 
.A(n_202),
.Y(n_662)
);

CKINVDCx20_ASAP7_75t_R g663 ( 
.A(n_384),
.Y(n_663)
);

CKINVDCx5p33_ASAP7_75t_R g664 ( 
.A(n_545),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_99),
.Y(n_665)
);

INVx3_ASAP7_75t_L g666 ( 
.A(n_107),
.Y(n_666)
);

CKINVDCx5p33_ASAP7_75t_R g667 ( 
.A(n_237),
.Y(n_667)
);

CKINVDCx5p33_ASAP7_75t_R g668 ( 
.A(n_548),
.Y(n_668)
);

CKINVDCx16_ASAP7_75t_R g669 ( 
.A(n_150),
.Y(n_669)
);

CKINVDCx5p33_ASAP7_75t_R g670 ( 
.A(n_298),
.Y(n_670)
);

CKINVDCx5p33_ASAP7_75t_R g671 ( 
.A(n_245),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_467),
.Y(n_672)
);

CKINVDCx20_ASAP7_75t_R g673 ( 
.A(n_592),
.Y(n_673)
);

CKINVDCx5p33_ASAP7_75t_R g674 ( 
.A(n_397),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_576),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_620),
.Y(n_676)
);

CKINVDCx5p33_ASAP7_75t_R g677 ( 
.A(n_568),
.Y(n_677)
);

CKINVDCx5p33_ASAP7_75t_R g678 ( 
.A(n_16),
.Y(n_678)
);

HB1xp67_ASAP7_75t_L g679 ( 
.A(n_372),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_384),
.Y(n_680)
);

CKINVDCx5p33_ASAP7_75t_R g681 ( 
.A(n_387),
.Y(n_681)
);

INVx2_ASAP7_75t_L g682 ( 
.A(n_268),
.Y(n_682)
);

CKINVDCx5p33_ASAP7_75t_R g683 ( 
.A(n_604),
.Y(n_683)
);

CKINVDCx5p33_ASAP7_75t_R g684 ( 
.A(n_248),
.Y(n_684)
);

CKINVDCx5p33_ASAP7_75t_R g685 ( 
.A(n_547),
.Y(n_685)
);

CKINVDCx14_ASAP7_75t_R g686 ( 
.A(n_135),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_303),
.Y(n_687)
);

CKINVDCx5p33_ASAP7_75t_R g688 ( 
.A(n_244),
.Y(n_688)
);

CKINVDCx5p33_ASAP7_75t_R g689 ( 
.A(n_450),
.Y(n_689)
);

BUFx10_ASAP7_75t_L g690 ( 
.A(n_273),
.Y(n_690)
);

CKINVDCx14_ASAP7_75t_R g691 ( 
.A(n_595),
.Y(n_691)
);

CKINVDCx5p33_ASAP7_75t_R g692 ( 
.A(n_383),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_407),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_601),
.Y(n_694)
);

CKINVDCx5p33_ASAP7_75t_R g695 ( 
.A(n_514),
.Y(n_695)
);

CKINVDCx5p33_ASAP7_75t_R g696 ( 
.A(n_382),
.Y(n_696)
);

INVx2_ASAP7_75t_L g697 ( 
.A(n_443),
.Y(n_697)
);

CKINVDCx5p33_ASAP7_75t_R g698 ( 
.A(n_480),
.Y(n_698)
);

CKINVDCx5p33_ASAP7_75t_R g699 ( 
.A(n_578),
.Y(n_699)
);

BUFx10_ASAP7_75t_L g700 ( 
.A(n_48),
.Y(n_700)
);

CKINVDCx5p33_ASAP7_75t_R g701 ( 
.A(n_355),
.Y(n_701)
);

CKINVDCx5p33_ASAP7_75t_R g702 ( 
.A(n_281),
.Y(n_702)
);

BUFx6f_ASAP7_75t_L g703 ( 
.A(n_262),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_164),
.Y(n_704)
);

CKINVDCx5p33_ASAP7_75t_R g705 ( 
.A(n_586),
.Y(n_705)
);

CKINVDCx5p33_ASAP7_75t_R g706 ( 
.A(n_79),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_6),
.Y(n_707)
);

CKINVDCx5p33_ASAP7_75t_R g708 ( 
.A(n_46),
.Y(n_708)
);

CKINVDCx5p33_ASAP7_75t_R g709 ( 
.A(n_326),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_569),
.Y(n_710)
);

BUFx5_ASAP7_75t_L g711 ( 
.A(n_590),
.Y(n_711)
);

CKINVDCx5p33_ASAP7_75t_R g712 ( 
.A(n_460),
.Y(n_712)
);

INVx1_ASAP7_75t_SL g713 ( 
.A(n_500),
.Y(n_713)
);

BUFx6f_ASAP7_75t_L g714 ( 
.A(n_558),
.Y(n_714)
);

CKINVDCx5p33_ASAP7_75t_R g715 ( 
.A(n_541),
.Y(n_715)
);

BUFx6f_ASAP7_75t_L g716 ( 
.A(n_273),
.Y(n_716)
);

INVx1_ASAP7_75t_SL g717 ( 
.A(n_389),
.Y(n_717)
);

CKINVDCx5p33_ASAP7_75t_R g718 ( 
.A(n_315),
.Y(n_718)
);

CKINVDCx5p33_ASAP7_75t_R g719 ( 
.A(n_62),
.Y(n_719)
);

CKINVDCx5p33_ASAP7_75t_R g720 ( 
.A(n_512),
.Y(n_720)
);

CKINVDCx5p33_ASAP7_75t_R g721 ( 
.A(n_549),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_232),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_104),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_574),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_310),
.Y(n_725)
);

CKINVDCx5p33_ASAP7_75t_R g726 ( 
.A(n_257),
.Y(n_726)
);

CKINVDCx5p33_ASAP7_75t_R g727 ( 
.A(n_38),
.Y(n_727)
);

CKINVDCx20_ASAP7_75t_R g728 ( 
.A(n_209),
.Y(n_728)
);

CKINVDCx5p33_ASAP7_75t_R g729 ( 
.A(n_247),
.Y(n_729)
);

CKINVDCx5p33_ASAP7_75t_R g730 ( 
.A(n_429),
.Y(n_730)
);

INVx1_ASAP7_75t_SL g731 ( 
.A(n_1),
.Y(n_731)
);

BUFx6f_ASAP7_75t_L g732 ( 
.A(n_199),
.Y(n_732)
);

CKINVDCx5p33_ASAP7_75t_R g733 ( 
.A(n_37),
.Y(n_733)
);

CKINVDCx5p33_ASAP7_75t_R g734 ( 
.A(n_528),
.Y(n_734)
);

CKINVDCx5p33_ASAP7_75t_R g735 ( 
.A(n_613),
.Y(n_735)
);

CKINVDCx5p33_ASAP7_75t_R g736 ( 
.A(n_226),
.Y(n_736)
);

BUFx3_ASAP7_75t_L g737 ( 
.A(n_422),
.Y(n_737)
);

BUFx6f_ASAP7_75t_L g738 ( 
.A(n_432),
.Y(n_738)
);

CKINVDCx5p33_ASAP7_75t_R g739 ( 
.A(n_20),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_611),
.Y(n_740)
);

CKINVDCx5p33_ASAP7_75t_R g741 ( 
.A(n_465),
.Y(n_741)
);

CKINVDCx20_ASAP7_75t_R g742 ( 
.A(n_478),
.Y(n_742)
);

CKINVDCx5p33_ASAP7_75t_R g743 ( 
.A(n_144),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_46),
.Y(n_744)
);

CKINVDCx5p33_ASAP7_75t_R g745 ( 
.A(n_561),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_223),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_209),
.Y(n_747)
);

CKINVDCx16_ASAP7_75t_R g748 ( 
.A(n_159),
.Y(n_748)
);

CKINVDCx5p33_ASAP7_75t_R g749 ( 
.A(n_175),
.Y(n_749)
);

CKINVDCx5p33_ASAP7_75t_R g750 ( 
.A(n_520),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_117),
.Y(n_751)
);

INVxp67_ASAP7_75t_L g752 ( 
.A(n_552),
.Y(n_752)
);

INVx1_ASAP7_75t_SL g753 ( 
.A(n_505),
.Y(n_753)
);

CKINVDCx5p33_ASAP7_75t_R g754 ( 
.A(n_200),
.Y(n_754)
);

CKINVDCx5p33_ASAP7_75t_R g755 ( 
.A(n_308),
.Y(n_755)
);

CKINVDCx5p33_ASAP7_75t_R g756 ( 
.A(n_366),
.Y(n_756)
);

CKINVDCx20_ASAP7_75t_R g757 ( 
.A(n_567),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_546),
.Y(n_758)
);

CKINVDCx5p33_ASAP7_75t_R g759 ( 
.A(n_60),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_272),
.Y(n_760)
);

BUFx6f_ASAP7_75t_L g761 ( 
.A(n_553),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_110),
.Y(n_762)
);

CKINVDCx5p33_ASAP7_75t_R g763 ( 
.A(n_27),
.Y(n_763)
);

CKINVDCx5p33_ASAP7_75t_R g764 ( 
.A(n_591),
.Y(n_764)
);

CKINVDCx5p33_ASAP7_75t_R g765 ( 
.A(n_612),
.Y(n_765)
);

CKINVDCx5p33_ASAP7_75t_R g766 ( 
.A(n_361),
.Y(n_766)
);

CKINVDCx5p33_ASAP7_75t_R g767 ( 
.A(n_147),
.Y(n_767)
);

CKINVDCx20_ASAP7_75t_R g768 ( 
.A(n_200),
.Y(n_768)
);

CKINVDCx20_ASAP7_75t_R g769 ( 
.A(n_184),
.Y(n_769)
);

CKINVDCx5p33_ASAP7_75t_R g770 ( 
.A(n_204),
.Y(n_770)
);

CKINVDCx20_ASAP7_75t_R g771 ( 
.A(n_299),
.Y(n_771)
);

BUFx6f_ASAP7_75t_L g772 ( 
.A(n_518),
.Y(n_772)
);

INVx3_ASAP7_75t_L g773 ( 
.A(n_606),
.Y(n_773)
);

CKINVDCx5p33_ASAP7_75t_R g774 ( 
.A(n_257),
.Y(n_774)
);

CKINVDCx5p33_ASAP7_75t_R g775 ( 
.A(n_411),
.Y(n_775)
);

CKINVDCx5p33_ASAP7_75t_R g776 ( 
.A(n_92),
.Y(n_776)
);

INVx2_ASAP7_75t_L g777 ( 
.A(n_599),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_618),
.Y(n_778)
);

CKINVDCx5p33_ASAP7_75t_R g779 ( 
.A(n_602),
.Y(n_779)
);

CKINVDCx5p33_ASAP7_75t_R g780 ( 
.A(n_275),
.Y(n_780)
);

CKINVDCx5p33_ASAP7_75t_R g781 ( 
.A(n_59),
.Y(n_781)
);

CKINVDCx5p33_ASAP7_75t_R g782 ( 
.A(n_92),
.Y(n_782)
);

INVx2_ASAP7_75t_L g783 ( 
.A(n_83),
.Y(n_783)
);

CKINVDCx5p33_ASAP7_75t_R g784 ( 
.A(n_538),
.Y(n_784)
);

INVx1_ASAP7_75t_SL g785 ( 
.A(n_43),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_85),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_534),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_551),
.Y(n_788)
);

INVx1_ASAP7_75t_L g789 ( 
.A(n_48),
.Y(n_789)
);

CKINVDCx5p33_ASAP7_75t_R g790 ( 
.A(n_100),
.Y(n_790)
);

CKINVDCx20_ASAP7_75t_R g791 ( 
.A(n_562),
.Y(n_791)
);

CKINVDCx5p33_ASAP7_75t_R g792 ( 
.A(n_598),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_502),
.Y(n_793)
);

CKINVDCx5p33_ASAP7_75t_R g794 ( 
.A(n_608),
.Y(n_794)
);

CKINVDCx5p33_ASAP7_75t_R g795 ( 
.A(n_584),
.Y(n_795)
);

BUFx6f_ASAP7_75t_L g796 ( 
.A(n_73),
.Y(n_796)
);

CKINVDCx5p33_ASAP7_75t_R g797 ( 
.A(n_283),
.Y(n_797)
);

CKINVDCx5p33_ASAP7_75t_R g798 ( 
.A(n_27),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_168),
.Y(n_799)
);

CKINVDCx5p33_ASAP7_75t_R g800 ( 
.A(n_507),
.Y(n_800)
);

BUFx10_ASAP7_75t_L g801 ( 
.A(n_555),
.Y(n_801)
);

CKINVDCx5p33_ASAP7_75t_R g802 ( 
.A(n_573),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_181),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_581),
.Y(n_804)
);

CKINVDCx5p33_ASAP7_75t_R g805 ( 
.A(n_471),
.Y(n_805)
);

CKINVDCx5p33_ASAP7_75t_R g806 ( 
.A(n_363),
.Y(n_806)
);

CKINVDCx5p33_ASAP7_75t_R g807 ( 
.A(n_536),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_374),
.Y(n_808)
);

CKINVDCx5p33_ASAP7_75t_R g809 ( 
.A(n_78),
.Y(n_809)
);

INVx1_ASAP7_75t_SL g810 ( 
.A(n_560),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_453),
.Y(n_811)
);

CKINVDCx5p33_ASAP7_75t_R g812 ( 
.A(n_201),
.Y(n_812)
);

BUFx6f_ASAP7_75t_L g813 ( 
.A(n_424),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_302),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_212),
.Y(n_815)
);

CKINVDCx5p33_ASAP7_75t_R g816 ( 
.A(n_377),
.Y(n_816)
);

CKINVDCx20_ASAP7_75t_R g817 ( 
.A(n_222),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_582),
.Y(n_818)
);

CKINVDCx5p33_ASAP7_75t_R g819 ( 
.A(n_302),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_417),
.Y(n_820)
);

CKINVDCx20_ASAP7_75t_R g821 ( 
.A(n_494),
.Y(n_821)
);

CKINVDCx5p33_ASAP7_75t_R g822 ( 
.A(n_354),
.Y(n_822)
);

BUFx6f_ASAP7_75t_L g823 ( 
.A(n_155),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_308),
.Y(n_824)
);

CKINVDCx5p33_ASAP7_75t_R g825 ( 
.A(n_14),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_472),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_331),
.Y(n_827)
);

BUFx6f_ASAP7_75t_L g828 ( 
.A(n_504),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_339),
.Y(n_829)
);

CKINVDCx5p33_ASAP7_75t_R g830 ( 
.A(n_10),
.Y(n_830)
);

CKINVDCx20_ASAP7_75t_R g831 ( 
.A(n_247),
.Y(n_831)
);

CKINVDCx5p33_ASAP7_75t_R g832 ( 
.A(n_120),
.Y(n_832)
);

CKINVDCx5p33_ASAP7_75t_R g833 ( 
.A(n_515),
.Y(n_833)
);

CKINVDCx20_ASAP7_75t_R g834 ( 
.A(n_407),
.Y(n_834)
);

CKINVDCx5p33_ASAP7_75t_R g835 ( 
.A(n_570),
.Y(n_835)
);

CKINVDCx5p33_ASAP7_75t_R g836 ( 
.A(n_385),
.Y(n_836)
);

CKINVDCx14_ASAP7_75t_R g837 ( 
.A(n_24),
.Y(n_837)
);

CKINVDCx5p33_ASAP7_75t_R g838 ( 
.A(n_381),
.Y(n_838)
);

CKINVDCx5p33_ASAP7_75t_R g839 ( 
.A(n_433),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_275),
.Y(n_840)
);

CKINVDCx20_ASAP7_75t_R g841 ( 
.A(n_221),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_78),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_557),
.Y(n_843)
);

CKINVDCx5p33_ASAP7_75t_R g844 ( 
.A(n_340),
.Y(n_844)
);

INVx2_ASAP7_75t_SL g845 ( 
.A(n_262),
.Y(n_845)
);

CKINVDCx20_ASAP7_75t_R g846 ( 
.A(n_87),
.Y(n_846)
);

CKINVDCx5p33_ASAP7_75t_R g847 ( 
.A(n_544),
.Y(n_847)
);

CKINVDCx20_ASAP7_75t_R g848 ( 
.A(n_532),
.Y(n_848)
);

INVx2_ASAP7_75t_L g849 ( 
.A(n_531),
.Y(n_849)
);

CKINVDCx5p33_ASAP7_75t_R g850 ( 
.A(n_26),
.Y(n_850)
);

BUFx5_ASAP7_75t_L g851 ( 
.A(n_187),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_339),
.Y(n_852)
);

CKINVDCx5p33_ASAP7_75t_R g853 ( 
.A(n_24),
.Y(n_853)
);

CKINVDCx5p33_ASAP7_75t_R g854 ( 
.A(n_105),
.Y(n_854)
);

BUFx6f_ASAP7_75t_L g855 ( 
.A(n_583),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_84),
.Y(n_856)
);

CKINVDCx20_ASAP7_75t_R g857 ( 
.A(n_132),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_360),
.Y(n_858)
);

CKINVDCx5p33_ASAP7_75t_R g859 ( 
.A(n_30),
.Y(n_859)
);

CKINVDCx5p33_ASAP7_75t_R g860 ( 
.A(n_158),
.Y(n_860)
);

CKINVDCx5p33_ASAP7_75t_R g861 ( 
.A(n_530),
.Y(n_861)
);

INVx1_ASAP7_75t_SL g862 ( 
.A(n_176),
.Y(n_862)
);

INVx2_ASAP7_75t_L g863 ( 
.A(n_123),
.Y(n_863)
);

CKINVDCx5p33_ASAP7_75t_R g864 ( 
.A(n_597),
.Y(n_864)
);

CKINVDCx5p33_ASAP7_75t_R g865 ( 
.A(n_23),
.Y(n_865)
);

CKINVDCx5p33_ASAP7_75t_R g866 ( 
.A(n_196),
.Y(n_866)
);

CKINVDCx20_ASAP7_75t_R g867 ( 
.A(n_73),
.Y(n_867)
);

CKINVDCx5p33_ASAP7_75t_R g868 ( 
.A(n_346),
.Y(n_868)
);

CKINVDCx5p33_ASAP7_75t_R g869 ( 
.A(n_463),
.Y(n_869)
);

BUFx3_ASAP7_75t_L g870 ( 
.A(n_213),
.Y(n_870)
);

CKINVDCx5p33_ASAP7_75t_R g871 ( 
.A(n_498),
.Y(n_871)
);

CKINVDCx5p33_ASAP7_75t_R g872 ( 
.A(n_317),
.Y(n_872)
);

BUFx6f_ASAP7_75t_L g873 ( 
.A(n_563),
.Y(n_873)
);

CKINVDCx5p33_ASAP7_75t_R g874 ( 
.A(n_64),
.Y(n_874)
);

CKINVDCx5p33_ASAP7_75t_R g875 ( 
.A(n_43),
.Y(n_875)
);

INVx2_ASAP7_75t_L g876 ( 
.A(n_431),
.Y(n_876)
);

CKINVDCx5p33_ASAP7_75t_R g877 ( 
.A(n_318),
.Y(n_877)
);

CKINVDCx5p33_ASAP7_75t_R g878 ( 
.A(n_71),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_55),
.Y(n_879)
);

CKINVDCx5p33_ASAP7_75t_R g880 ( 
.A(n_188),
.Y(n_880)
);

INVx1_ASAP7_75t_L g881 ( 
.A(n_289),
.Y(n_881)
);

INVx2_ASAP7_75t_L g882 ( 
.A(n_533),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_222),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_83),
.Y(n_884)
);

CKINVDCx5p33_ASAP7_75t_R g885 ( 
.A(n_525),
.Y(n_885)
);

CKINVDCx20_ASAP7_75t_R g886 ( 
.A(n_425),
.Y(n_886)
);

CKINVDCx20_ASAP7_75t_R g887 ( 
.A(n_13),
.Y(n_887)
);

CKINVDCx5p33_ASAP7_75t_R g888 ( 
.A(n_206),
.Y(n_888)
);

BUFx10_ASAP7_75t_L g889 ( 
.A(n_30),
.Y(n_889)
);

CKINVDCx20_ASAP7_75t_R g890 ( 
.A(n_215),
.Y(n_890)
);

CKINVDCx5p33_ASAP7_75t_R g891 ( 
.A(n_366),
.Y(n_891)
);

CKINVDCx5p33_ASAP7_75t_R g892 ( 
.A(n_15),
.Y(n_892)
);

CKINVDCx5p33_ASAP7_75t_R g893 ( 
.A(n_251),
.Y(n_893)
);

BUFx2_ASAP7_75t_L g894 ( 
.A(n_11),
.Y(n_894)
);

INVx1_ASAP7_75t_L g895 ( 
.A(n_162),
.Y(n_895)
);

BUFx10_ASAP7_75t_L g896 ( 
.A(n_333),
.Y(n_896)
);

CKINVDCx5p33_ASAP7_75t_R g897 ( 
.A(n_249),
.Y(n_897)
);

CKINVDCx20_ASAP7_75t_R g898 ( 
.A(n_401),
.Y(n_898)
);

CKINVDCx5p33_ASAP7_75t_R g899 ( 
.A(n_390),
.Y(n_899)
);

CKINVDCx14_ASAP7_75t_R g900 ( 
.A(n_359),
.Y(n_900)
);

INVx2_ASAP7_75t_SL g901 ( 
.A(n_41),
.Y(n_901)
);

CKINVDCx20_ASAP7_75t_R g902 ( 
.A(n_235),
.Y(n_902)
);

CKINVDCx5p33_ASAP7_75t_R g903 ( 
.A(n_240),
.Y(n_903)
);

BUFx6f_ASAP7_75t_L g904 ( 
.A(n_521),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_15),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_100),
.Y(n_906)
);

CKINVDCx5p33_ASAP7_75t_R g907 ( 
.A(n_94),
.Y(n_907)
);

CKINVDCx5p33_ASAP7_75t_R g908 ( 
.A(n_529),
.Y(n_908)
);

CKINVDCx5p33_ASAP7_75t_R g909 ( 
.A(n_149),
.Y(n_909)
);

CKINVDCx5p33_ASAP7_75t_R g910 ( 
.A(n_458),
.Y(n_910)
);

CKINVDCx20_ASAP7_75t_R g911 ( 
.A(n_313),
.Y(n_911)
);

CKINVDCx5p33_ASAP7_75t_R g912 ( 
.A(n_457),
.Y(n_912)
);

INVx1_ASAP7_75t_L g913 ( 
.A(n_351),
.Y(n_913)
);

CKINVDCx5p33_ASAP7_75t_R g914 ( 
.A(n_37),
.Y(n_914)
);

CKINVDCx5p33_ASAP7_75t_R g915 ( 
.A(n_135),
.Y(n_915)
);

INVx2_ASAP7_75t_L g916 ( 
.A(n_16),
.Y(n_916)
);

CKINVDCx5p33_ASAP7_75t_R g917 ( 
.A(n_128),
.Y(n_917)
);

INVx1_ASAP7_75t_L g918 ( 
.A(n_134),
.Y(n_918)
);

INVx1_ASAP7_75t_SL g919 ( 
.A(n_84),
.Y(n_919)
);

INVx1_ASAP7_75t_L g920 ( 
.A(n_155),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_596),
.Y(n_921)
);

HB1xp67_ASAP7_75t_L g922 ( 
.A(n_331),
.Y(n_922)
);

CKINVDCx5p33_ASAP7_75t_R g923 ( 
.A(n_440),
.Y(n_923)
);

INVx1_ASAP7_75t_L g924 ( 
.A(n_368),
.Y(n_924)
);

CKINVDCx5p33_ASAP7_75t_R g925 ( 
.A(n_232),
.Y(n_925)
);

CKINVDCx20_ASAP7_75t_R g926 ( 
.A(n_484),
.Y(n_926)
);

INVx1_ASAP7_75t_L g927 ( 
.A(n_287),
.Y(n_927)
);

CKINVDCx20_ASAP7_75t_R g928 ( 
.A(n_29),
.Y(n_928)
);

CKINVDCx5p33_ASAP7_75t_R g929 ( 
.A(n_328),
.Y(n_929)
);

INVx1_ASAP7_75t_L g930 ( 
.A(n_540),
.Y(n_930)
);

CKINVDCx5p33_ASAP7_75t_R g931 ( 
.A(n_607),
.Y(n_931)
);

CKINVDCx5p33_ASAP7_75t_R g932 ( 
.A(n_221),
.Y(n_932)
);

CKINVDCx5p33_ASAP7_75t_R g933 ( 
.A(n_523),
.Y(n_933)
);

CKINVDCx5p33_ASAP7_75t_R g934 ( 
.A(n_167),
.Y(n_934)
);

INVx1_ASAP7_75t_L g935 ( 
.A(n_437),
.Y(n_935)
);

CKINVDCx16_ASAP7_75t_R g936 ( 
.A(n_372),
.Y(n_936)
);

CKINVDCx5p33_ASAP7_75t_R g937 ( 
.A(n_177),
.Y(n_937)
);

INVx2_ASAP7_75t_L g938 ( 
.A(n_47),
.Y(n_938)
);

CKINVDCx5p33_ASAP7_75t_R g939 ( 
.A(n_438),
.Y(n_939)
);

CKINVDCx5p33_ASAP7_75t_R g940 ( 
.A(n_157),
.Y(n_940)
);

CKINVDCx16_ASAP7_75t_R g941 ( 
.A(n_332),
.Y(n_941)
);

CKINVDCx5p33_ASAP7_75t_R g942 ( 
.A(n_579),
.Y(n_942)
);

CKINVDCx5p33_ASAP7_75t_R g943 ( 
.A(n_298),
.Y(n_943)
);

CKINVDCx5p33_ASAP7_75t_R g944 ( 
.A(n_35),
.Y(n_944)
);

INVx2_ASAP7_75t_SL g945 ( 
.A(n_301),
.Y(n_945)
);

CKINVDCx20_ASAP7_75t_R g946 ( 
.A(n_473),
.Y(n_946)
);

CKINVDCx5p33_ASAP7_75t_R g947 ( 
.A(n_251),
.Y(n_947)
);

CKINVDCx5p33_ASAP7_75t_R g948 ( 
.A(n_250),
.Y(n_948)
);

CKINVDCx5p33_ASAP7_75t_R g949 ( 
.A(n_603),
.Y(n_949)
);

INVx1_ASAP7_75t_L g950 ( 
.A(n_609),
.Y(n_950)
);

BUFx3_ASAP7_75t_L g951 ( 
.A(n_587),
.Y(n_951)
);

INVx2_ASAP7_75t_L g952 ( 
.A(n_217),
.Y(n_952)
);

HB1xp67_ASAP7_75t_L g953 ( 
.A(n_235),
.Y(n_953)
);

CKINVDCx5p33_ASAP7_75t_R g954 ( 
.A(n_338),
.Y(n_954)
);

CKINVDCx5p33_ASAP7_75t_R g955 ( 
.A(n_594),
.Y(n_955)
);

INVx1_ASAP7_75t_L g956 ( 
.A(n_427),
.Y(n_956)
);

INVx1_ASAP7_75t_L g957 ( 
.A(n_185),
.Y(n_957)
);

BUFx5_ASAP7_75t_L g958 ( 
.A(n_537),
.Y(n_958)
);

INVx1_ASAP7_75t_L g959 ( 
.A(n_26),
.Y(n_959)
);

CKINVDCx5p33_ASAP7_75t_R g960 ( 
.A(n_58),
.Y(n_960)
);

CKINVDCx5p33_ASAP7_75t_R g961 ( 
.A(n_368),
.Y(n_961)
);

CKINVDCx5p33_ASAP7_75t_R g962 ( 
.A(n_71),
.Y(n_962)
);

INVx1_ASAP7_75t_L g963 ( 
.A(n_411),
.Y(n_963)
);

CKINVDCx20_ASAP7_75t_R g964 ( 
.A(n_170),
.Y(n_964)
);

CKINVDCx5p33_ASAP7_75t_R g965 ( 
.A(n_88),
.Y(n_965)
);

INVx1_ASAP7_75t_L g966 ( 
.A(n_225),
.Y(n_966)
);

INVx1_ASAP7_75t_L g967 ( 
.A(n_543),
.Y(n_967)
);

CKINVDCx5p33_ASAP7_75t_R g968 ( 
.A(n_334),
.Y(n_968)
);

INVx1_ASAP7_75t_L g969 ( 
.A(n_0),
.Y(n_969)
);

BUFx6f_ASAP7_75t_L g970 ( 
.A(n_332),
.Y(n_970)
);

CKINVDCx5p33_ASAP7_75t_R g971 ( 
.A(n_8),
.Y(n_971)
);

CKINVDCx5p33_ASAP7_75t_R g972 ( 
.A(n_455),
.Y(n_972)
);

CKINVDCx5p33_ASAP7_75t_R g973 ( 
.A(n_35),
.Y(n_973)
);

CKINVDCx5p33_ASAP7_75t_R g974 ( 
.A(n_322),
.Y(n_974)
);

CKINVDCx5p33_ASAP7_75t_R g975 ( 
.A(n_447),
.Y(n_975)
);

CKINVDCx5p33_ASAP7_75t_R g976 ( 
.A(n_190),
.Y(n_976)
);

CKINVDCx20_ASAP7_75t_R g977 ( 
.A(n_404),
.Y(n_977)
);

CKINVDCx5p33_ASAP7_75t_R g978 ( 
.A(n_163),
.Y(n_978)
);

CKINVDCx5p33_ASAP7_75t_R g979 ( 
.A(n_94),
.Y(n_979)
);

INVx1_ASAP7_75t_L g980 ( 
.A(n_231),
.Y(n_980)
);

CKINVDCx5p33_ASAP7_75t_R g981 ( 
.A(n_550),
.Y(n_981)
);

INVx1_ASAP7_75t_L g982 ( 
.A(n_605),
.Y(n_982)
);

CKINVDCx5p33_ASAP7_75t_R g983 ( 
.A(n_559),
.Y(n_983)
);

INVx1_ASAP7_75t_L g984 ( 
.A(n_102),
.Y(n_984)
);

CKINVDCx5p33_ASAP7_75t_R g985 ( 
.A(n_565),
.Y(n_985)
);

CKINVDCx5p33_ASAP7_75t_R g986 ( 
.A(n_370),
.Y(n_986)
);

INVx1_ASAP7_75t_L g987 ( 
.A(n_354),
.Y(n_987)
);

BUFx3_ASAP7_75t_L g988 ( 
.A(n_56),
.Y(n_988)
);

INVx1_ASAP7_75t_SL g989 ( 
.A(n_571),
.Y(n_989)
);

INVx1_ASAP7_75t_L g990 ( 
.A(n_406),
.Y(n_990)
);

CKINVDCx5p33_ASAP7_75t_R g991 ( 
.A(n_294),
.Y(n_991)
);

BUFx3_ASAP7_75t_L g992 ( 
.A(n_158),
.Y(n_992)
);

INVx1_ASAP7_75t_L g993 ( 
.A(n_333),
.Y(n_993)
);

CKINVDCx5p33_ASAP7_75t_R g994 ( 
.A(n_324),
.Y(n_994)
);

CKINVDCx5p33_ASAP7_75t_R g995 ( 
.A(n_616),
.Y(n_995)
);

INVx1_ASAP7_75t_L g996 ( 
.A(n_163),
.Y(n_996)
);

CKINVDCx5p33_ASAP7_75t_R g997 ( 
.A(n_542),
.Y(n_997)
);

CKINVDCx5p33_ASAP7_75t_R g998 ( 
.A(n_324),
.Y(n_998)
);

CKINVDCx5p33_ASAP7_75t_R g999 ( 
.A(n_406),
.Y(n_999)
);

BUFx2_ASAP7_75t_L g1000 ( 
.A(n_495),
.Y(n_1000)
);

CKINVDCx16_ASAP7_75t_R g1001 ( 
.A(n_93),
.Y(n_1001)
);

CKINVDCx5p33_ASAP7_75t_R g1002 ( 
.A(n_34),
.Y(n_1002)
);

CKINVDCx5p33_ASAP7_75t_R g1003 ( 
.A(n_230),
.Y(n_1003)
);

INVx1_ASAP7_75t_L g1004 ( 
.A(n_51),
.Y(n_1004)
);

CKINVDCx20_ASAP7_75t_R g1005 ( 
.A(n_554),
.Y(n_1005)
);

CKINVDCx20_ASAP7_75t_R g1006 ( 
.A(n_310),
.Y(n_1006)
);

INVx1_ASAP7_75t_SL g1007 ( 
.A(n_481),
.Y(n_1007)
);

CKINVDCx5p33_ASAP7_75t_R g1008 ( 
.A(n_575),
.Y(n_1008)
);

BUFx6f_ASAP7_75t_L g1009 ( 
.A(n_526),
.Y(n_1009)
);

CKINVDCx5p33_ASAP7_75t_R g1010 ( 
.A(n_389),
.Y(n_1010)
);

CKINVDCx5p33_ASAP7_75t_R g1011 ( 
.A(n_413),
.Y(n_1011)
);

INVx1_ASAP7_75t_L g1012 ( 
.A(n_149),
.Y(n_1012)
);

CKINVDCx5p33_ASAP7_75t_R g1013 ( 
.A(n_577),
.Y(n_1013)
);

CKINVDCx20_ASAP7_75t_R g1014 ( 
.A(n_299),
.Y(n_1014)
);

INVx2_ASAP7_75t_L g1015 ( 
.A(n_385),
.Y(n_1015)
);

INVx1_ASAP7_75t_L g1016 ( 
.A(n_315),
.Y(n_1016)
);

INVx1_ASAP7_75t_SL g1017 ( 
.A(n_585),
.Y(n_1017)
);

INVx2_ASAP7_75t_SL g1018 ( 
.A(n_287),
.Y(n_1018)
);

CKINVDCx5p33_ASAP7_75t_R g1019 ( 
.A(n_503),
.Y(n_1019)
);

CKINVDCx5p33_ASAP7_75t_R g1020 ( 
.A(n_174),
.Y(n_1020)
);

INVx2_ASAP7_75t_L g1021 ( 
.A(n_208),
.Y(n_1021)
);

CKINVDCx5p33_ASAP7_75t_R g1022 ( 
.A(n_619),
.Y(n_1022)
);

CKINVDCx5p33_ASAP7_75t_R g1023 ( 
.A(n_556),
.Y(n_1023)
);

CKINVDCx5p33_ASAP7_75t_R g1024 ( 
.A(n_572),
.Y(n_1024)
);

CKINVDCx5p33_ASAP7_75t_R g1025 ( 
.A(n_22),
.Y(n_1025)
);

INVx1_ASAP7_75t_SL g1026 ( 
.A(n_127),
.Y(n_1026)
);

INVx1_ASAP7_75t_L g1027 ( 
.A(n_234),
.Y(n_1027)
);

INVx1_ASAP7_75t_L g1028 ( 
.A(n_89),
.Y(n_1028)
);

CKINVDCx5p33_ASAP7_75t_R g1029 ( 
.A(n_268),
.Y(n_1029)
);

BUFx10_ASAP7_75t_L g1030 ( 
.A(n_334),
.Y(n_1030)
);

CKINVDCx20_ASAP7_75t_R g1031 ( 
.A(n_237),
.Y(n_1031)
);

BUFx10_ASAP7_75t_L g1032 ( 
.A(n_123),
.Y(n_1032)
);

INVx1_ASAP7_75t_L g1033 ( 
.A(n_276),
.Y(n_1033)
);

CKINVDCx5p33_ASAP7_75t_R g1034 ( 
.A(n_589),
.Y(n_1034)
);

CKINVDCx5p33_ASAP7_75t_R g1035 ( 
.A(n_141),
.Y(n_1035)
);

CKINVDCx5p33_ASAP7_75t_R g1036 ( 
.A(n_566),
.Y(n_1036)
);

CKINVDCx5p33_ASAP7_75t_R g1037 ( 
.A(n_31),
.Y(n_1037)
);

CKINVDCx5p33_ASAP7_75t_R g1038 ( 
.A(n_203),
.Y(n_1038)
);

CKINVDCx5p33_ASAP7_75t_R g1039 ( 
.A(n_117),
.Y(n_1039)
);

CKINVDCx5p33_ASAP7_75t_R g1040 ( 
.A(n_25),
.Y(n_1040)
);

CKINVDCx5p33_ASAP7_75t_R g1041 ( 
.A(n_174),
.Y(n_1041)
);

CKINVDCx5p33_ASAP7_75t_R g1042 ( 
.A(n_600),
.Y(n_1042)
);

INVx1_ASAP7_75t_L g1043 ( 
.A(n_375),
.Y(n_1043)
);

INVx1_ASAP7_75t_L g1044 ( 
.A(n_150),
.Y(n_1044)
);

CKINVDCx5p33_ASAP7_75t_R g1045 ( 
.A(n_370),
.Y(n_1045)
);

CKINVDCx5p33_ASAP7_75t_R g1046 ( 
.A(n_161),
.Y(n_1046)
);

CKINVDCx5p33_ASAP7_75t_R g1047 ( 
.A(n_290),
.Y(n_1047)
);

INVx1_ASAP7_75t_L g1048 ( 
.A(n_166),
.Y(n_1048)
);

INVx1_ASAP7_75t_L g1049 ( 
.A(n_125),
.Y(n_1049)
);

INVx1_ASAP7_75t_L g1050 ( 
.A(n_85),
.Y(n_1050)
);

INVx1_ASAP7_75t_SL g1051 ( 
.A(n_116),
.Y(n_1051)
);

BUFx2_ASAP7_75t_L g1052 ( 
.A(n_686),
.Y(n_1052)
);

AND2x2_ASAP7_75t_L g1053 ( 
.A(n_686),
.B(n_0),
.Y(n_1053)
);

BUFx6f_ASAP7_75t_L g1054 ( 
.A(n_714),
.Y(n_1054)
);

NAND2xp5_ASAP7_75t_SL g1055 ( 
.A(n_773),
.B(n_1),
.Y(n_1055)
);

INVx1_ASAP7_75t_SL g1056 ( 
.A(n_654),
.Y(n_1056)
);

BUFx6f_ASAP7_75t_L g1057 ( 
.A(n_714),
.Y(n_1057)
);

CKINVDCx5p33_ASAP7_75t_R g1058 ( 
.A(n_673),
.Y(n_1058)
);

NOR2xp33_ASAP7_75t_L g1059 ( 
.A(n_773),
.B(n_2),
.Y(n_1059)
);

NOR2xp33_ASAP7_75t_L g1060 ( 
.A(n_627),
.B(n_2),
.Y(n_1060)
);

INVx2_ASAP7_75t_L g1061 ( 
.A(n_851),
.Y(n_1061)
);

NOR2xp33_ASAP7_75t_L g1062 ( 
.A(n_1000),
.B(n_3),
.Y(n_1062)
);

INVx1_ASAP7_75t_SL g1063 ( 
.A(n_894),
.Y(n_1063)
);

INVx5_ASAP7_75t_L g1064 ( 
.A(n_714),
.Y(n_1064)
);

INVx5_ASAP7_75t_L g1065 ( 
.A(n_714),
.Y(n_1065)
);

AND2x4_ASAP7_75t_L g1066 ( 
.A(n_666),
.B(n_3),
.Y(n_1066)
);

INVx2_ASAP7_75t_SL g1067 ( 
.A(n_646),
.Y(n_1067)
);

NOR2xp33_ASAP7_75t_L g1068 ( 
.A(n_626),
.B(n_4),
.Y(n_1068)
);

INVx5_ASAP7_75t_L g1069 ( 
.A(n_738),
.Y(n_1069)
);

INVx5_ASAP7_75t_L g1070 ( 
.A(n_738),
.Y(n_1070)
);

BUFx2_ASAP7_75t_L g1071 ( 
.A(n_837),
.Y(n_1071)
);

AND2x2_ASAP7_75t_L g1072 ( 
.A(n_837),
.B(n_4),
.Y(n_1072)
);

NOR2xp33_ASAP7_75t_L g1073 ( 
.A(n_642),
.B(n_5),
.Y(n_1073)
);

AND2x6_ASAP7_75t_L g1074 ( 
.A(n_737),
.B(n_621),
.Y(n_1074)
);

AND2x4_ASAP7_75t_L g1075 ( 
.A(n_666),
.B(n_6),
.Y(n_1075)
);

BUFx3_ASAP7_75t_L g1076 ( 
.A(n_636),
.Y(n_1076)
);

NOR2xp33_ASAP7_75t_SL g1077 ( 
.A(n_622),
.B(n_617),
.Y(n_1077)
);

AND2x2_ASAP7_75t_L g1078 ( 
.A(n_900),
.B(n_7),
.Y(n_1078)
);

NOR2xp33_ASAP7_75t_L g1079 ( 
.A(n_647),
.B(n_7),
.Y(n_1079)
);

INVx5_ASAP7_75t_L g1080 ( 
.A(n_738),
.Y(n_1080)
);

BUFx6f_ASAP7_75t_L g1081 ( 
.A(n_738),
.Y(n_1081)
);

INVx3_ASAP7_75t_L g1082 ( 
.A(n_646),
.Y(n_1082)
);

INVx1_ASAP7_75t_L g1083 ( 
.A(n_851),
.Y(n_1083)
);

INVx2_ASAP7_75t_L g1084 ( 
.A(n_851),
.Y(n_1084)
);

NOR2xp33_ASAP7_75t_L g1085 ( 
.A(n_672),
.B(n_8),
.Y(n_1085)
);

AND2x2_ASAP7_75t_L g1086 ( 
.A(n_900),
.B(n_669),
.Y(n_1086)
);

BUFx8_ASAP7_75t_L g1087 ( 
.A(n_851),
.Y(n_1087)
);

INVx2_ASAP7_75t_L g1088 ( 
.A(n_851),
.Y(n_1088)
);

AND2x4_ASAP7_75t_L g1089 ( 
.A(n_870),
.B(n_9),
.Y(n_1089)
);

CKINVDCx6p67_ASAP7_75t_R g1090 ( 
.A(n_636),
.Y(n_1090)
);

HB1xp67_ASAP7_75t_L g1091 ( 
.A(n_661),
.Y(n_1091)
);

BUFx6f_ASAP7_75t_L g1092 ( 
.A(n_761),
.Y(n_1092)
);

NOR2xp33_ASAP7_75t_L g1093 ( 
.A(n_675),
.B(n_9),
.Y(n_1093)
);

NOR2x1_ASAP7_75t_L g1094 ( 
.A(n_870),
.B(n_10),
.Y(n_1094)
);

NAND2xp5_ASAP7_75t_L g1095 ( 
.A(n_679),
.B(n_11),
.Y(n_1095)
);

BUFx6f_ASAP7_75t_L g1096 ( 
.A(n_761),
.Y(n_1096)
);

BUFx6f_ASAP7_75t_L g1097 ( 
.A(n_761),
.Y(n_1097)
);

BUFx8_ASAP7_75t_SL g1098 ( 
.A(n_887),
.Y(n_1098)
);

AND2x4_ASAP7_75t_L g1099 ( 
.A(n_988),
.B(n_12),
.Y(n_1099)
);

BUFx8_ASAP7_75t_L g1100 ( 
.A(n_851),
.Y(n_1100)
);

BUFx2_ASAP7_75t_L g1101 ( 
.A(n_922),
.Y(n_1101)
);

NOR2xp33_ASAP7_75t_L g1102 ( 
.A(n_676),
.B(n_12),
.Y(n_1102)
);

BUFx6f_ASAP7_75t_L g1103 ( 
.A(n_761),
.Y(n_1103)
);

INVx5_ASAP7_75t_L g1104 ( 
.A(n_772),
.Y(n_1104)
);

AND2x4_ASAP7_75t_L g1105 ( 
.A(n_988),
.B(n_13),
.Y(n_1105)
);

NAND2xp5_ASAP7_75t_L g1106 ( 
.A(n_953),
.B(n_14),
.Y(n_1106)
);

INVx1_ASAP7_75t_L g1107 ( 
.A(n_851),
.Y(n_1107)
);

INVx3_ASAP7_75t_L g1108 ( 
.A(n_646),
.Y(n_1108)
);

AND2x4_ASAP7_75t_L g1109 ( 
.A(n_992),
.B(n_17),
.Y(n_1109)
);

AND2x2_ASAP7_75t_L g1110 ( 
.A(n_748),
.B(n_17),
.Y(n_1110)
);

NAND2xp5_ASAP7_75t_L g1111 ( 
.A(n_845),
.B(n_18),
.Y(n_1111)
);

INVx2_ASAP7_75t_L g1112 ( 
.A(n_992),
.Y(n_1112)
);

INVx2_ASAP7_75t_L g1113 ( 
.A(n_901),
.Y(n_1113)
);

CKINVDCx6p67_ASAP7_75t_R g1114 ( 
.A(n_636),
.Y(n_1114)
);

NOR2xp33_ASAP7_75t_L g1115 ( 
.A(n_694),
.B(n_18),
.Y(n_1115)
);

AND2x4_ASAP7_75t_L g1116 ( 
.A(n_656),
.B(n_19),
.Y(n_1116)
);

NAND2xp5_ASAP7_75t_L g1117 ( 
.A(n_945),
.B(n_19),
.Y(n_1117)
);

HB1xp67_ASAP7_75t_L g1118 ( 
.A(n_645),
.Y(n_1118)
);

AND2x2_ASAP7_75t_L g1119 ( 
.A(n_936),
.B(n_20),
.Y(n_1119)
);

BUFx12f_ASAP7_75t_L g1120 ( 
.A(n_690),
.Y(n_1120)
);

INVx5_ASAP7_75t_L g1121 ( 
.A(n_772),
.Y(n_1121)
);

BUFx12f_ASAP7_75t_L g1122 ( 
.A(n_690),
.Y(n_1122)
);

BUFx6f_ASAP7_75t_L g1123 ( 
.A(n_772),
.Y(n_1123)
);

BUFx2_ASAP7_75t_L g1124 ( 
.A(n_941),
.Y(n_1124)
);

BUFx3_ASAP7_75t_L g1125 ( 
.A(n_801),
.Y(n_1125)
);

INVx3_ASAP7_75t_L g1126 ( 
.A(n_690),
.Y(n_1126)
);

NAND2xp5_ASAP7_75t_L g1127 ( 
.A(n_1018),
.B(n_21),
.Y(n_1127)
);

INVx1_ASAP7_75t_L g1128 ( 
.A(n_656),
.Y(n_1128)
);

BUFx12f_ASAP7_75t_L g1129 ( 
.A(n_700),
.Y(n_1129)
);

INVx1_ASAP7_75t_L g1130 ( 
.A(n_658),
.Y(n_1130)
);

INVx5_ASAP7_75t_L g1131 ( 
.A(n_772),
.Y(n_1131)
);

AND2x4_ASAP7_75t_L g1132 ( 
.A(n_658),
.B(n_21),
.Y(n_1132)
);

INVx2_ASAP7_75t_L g1133 ( 
.A(n_711),
.Y(n_1133)
);

BUFx8_ASAP7_75t_SL g1134 ( 
.A(n_887),
.Y(n_1134)
);

BUFx8_ASAP7_75t_SL g1135 ( 
.A(n_890),
.Y(n_1135)
);

XOR2xp5_ASAP7_75t_L g1136 ( 
.A(n_890),
.B(n_22),
.Y(n_1136)
);

INVx3_ASAP7_75t_L g1137 ( 
.A(n_700),
.Y(n_1137)
);

NAND2xp5_ASAP7_75t_L g1138 ( 
.A(n_1001),
.B(n_23),
.Y(n_1138)
);

NAND2xp5_ASAP7_75t_L g1139 ( 
.A(n_641),
.B(n_25),
.Y(n_1139)
);

INVx3_ASAP7_75t_L g1140 ( 
.A(n_700),
.Y(n_1140)
);

BUFx2_ASAP7_75t_L g1141 ( 
.A(n_623),
.Y(n_1141)
);

BUFx6f_ASAP7_75t_L g1142 ( 
.A(n_813),
.Y(n_1142)
);

BUFx2_ASAP7_75t_L g1143 ( 
.A(n_624),
.Y(n_1143)
);

HB1xp67_ASAP7_75t_L g1144 ( 
.A(n_628),
.Y(n_1144)
);

NOR2xp33_ASAP7_75t_R g1145 ( 
.A(n_630),
.B(n_412),
.Y(n_1145)
);

BUFx3_ASAP7_75t_L g1146 ( 
.A(n_801),
.Y(n_1146)
);

BUFx2_ASAP7_75t_L g1147 ( 
.A(n_629),
.Y(n_1147)
);

NAND2xp5_ASAP7_75t_L g1148 ( 
.A(n_644),
.B(n_28),
.Y(n_1148)
);

INVx2_ASAP7_75t_L g1149 ( 
.A(n_711),
.Y(n_1149)
);

INVx1_ASAP7_75t_L g1150 ( 
.A(n_682),
.Y(n_1150)
);

BUFx6f_ASAP7_75t_L g1151 ( 
.A(n_813),
.Y(n_1151)
);

INVx4_ASAP7_75t_L g1152 ( 
.A(n_801),
.Y(n_1152)
);

AND2x2_ASAP7_75t_L g1153 ( 
.A(n_889),
.B(n_28),
.Y(n_1153)
);

NAND2xp5_ASAP7_75t_L g1154 ( 
.A(n_659),
.B(n_29),
.Y(n_1154)
);

AND2x4_ASAP7_75t_L g1155 ( 
.A(n_682),
.B(n_31),
.Y(n_1155)
);

INVx5_ASAP7_75t_L g1156 ( 
.A(n_813),
.Y(n_1156)
);

NAND2xp5_ASAP7_75t_L g1157 ( 
.A(n_660),
.B(n_32),
.Y(n_1157)
);

NAND2xp5_ASAP7_75t_L g1158 ( 
.A(n_665),
.B(n_32),
.Y(n_1158)
);

INVx5_ASAP7_75t_L g1159 ( 
.A(n_813),
.Y(n_1159)
);

INVx2_ASAP7_75t_L g1160 ( 
.A(n_711),
.Y(n_1160)
);

NAND2xp5_ASAP7_75t_L g1161 ( 
.A(n_680),
.B(n_33),
.Y(n_1161)
);

HB1xp67_ASAP7_75t_L g1162 ( 
.A(n_633),
.Y(n_1162)
);

NAND2xp5_ASAP7_75t_L g1163 ( 
.A(n_687),
.B(n_33),
.Y(n_1163)
);

BUFx12f_ASAP7_75t_L g1164 ( 
.A(n_889),
.Y(n_1164)
);

INVx5_ASAP7_75t_L g1165 ( 
.A(n_828),
.Y(n_1165)
);

INVx1_ASAP7_75t_L g1166 ( 
.A(n_783),
.Y(n_1166)
);

AND2x6_ASAP7_75t_L g1167 ( 
.A(n_737),
.B(n_951),
.Y(n_1167)
);

BUFx6f_ASAP7_75t_L g1168 ( 
.A(n_828),
.Y(n_1168)
);

NAND2xp5_ASAP7_75t_L g1169 ( 
.A(n_693),
.B(n_34),
.Y(n_1169)
);

CKINVDCx11_ASAP7_75t_R g1170 ( 
.A(n_898),
.Y(n_1170)
);

BUFx6f_ASAP7_75t_L g1171 ( 
.A(n_828),
.Y(n_1171)
);

INVx5_ASAP7_75t_L g1172 ( 
.A(n_828),
.Y(n_1172)
);

AND2x4_ASAP7_75t_L g1173 ( 
.A(n_783),
.B(n_36),
.Y(n_1173)
);

INVx5_ASAP7_75t_L g1174 ( 
.A(n_855),
.Y(n_1174)
);

INVx2_ASAP7_75t_L g1175 ( 
.A(n_711),
.Y(n_1175)
);

BUFx2_ASAP7_75t_L g1176 ( 
.A(n_634),
.Y(n_1176)
);

AND2x4_ASAP7_75t_L g1177 ( 
.A(n_863),
.B(n_36),
.Y(n_1177)
);

BUFx6f_ASAP7_75t_L g1178 ( 
.A(n_855),
.Y(n_1178)
);

NAND2xp5_ASAP7_75t_L g1179 ( 
.A(n_704),
.B(n_38),
.Y(n_1179)
);

HB1xp67_ASAP7_75t_L g1180 ( 
.A(n_643),
.Y(n_1180)
);

AOI22xp5_ASAP7_75t_L g1181 ( 
.A1(n_1056),
.A2(n_640),
.B1(n_926),
.B2(n_631),
.Y(n_1181)
);

AOI22xp5_ASAP7_75t_L g1182 ( 
.A1(n_1063),
.A2(n_640),
.B1(n_926),
.B2(n_631),
.Y(n_1182)
);

BUFx6f_ASAP7_75t_SL g1183 ( 
.A(n_1116),
.Y(n_1183)
);

AO22x2_ASAP7_75t_L g1184 ( 
.A1(n_1136),
.A2(n_638),
.B1(n_717),
.B2(n_637),
.Y(n_1184)
);

OAI22xp33_ASAP7_75t_L g1185 ( 
.A1(n_1124),
.A2(n_902),
.B1(n_911),
.B2(n_898),
.Y(n_1185)
);

INVx2_ASAP7_75t_L g1186 ( 
.A(n_1112),
.Y(n_1186)
);

OAI22xp5_ASAP7_75t_SL g1187 ( 
.A1(n_1058),
.A2(n_911),
.B1(n_928),
.B2(n_902),
.Y(n_1187)
);

AND2x2_ASAP7_75t_L g1188 ( 
.A(n_1052),
.B(n_630),
.Y(n_1188)
);

AOI22xp5_ASAP7_75t_L g1189 ( 
.A1(n_1086),
.A2(n_946),
.B1(n_651),
.B2(n_653),
.Y(n_1189)
);

AO22x2_ASAP7_75t_L g1190 ( 
.A1(n_1110),
.A2(n_785),
.B1(n_862),
.B2(n_731),
.Y(n_1190)
);

AND2x2_ASAP7_75t_L g1191 ( 
.A(n_1071),
.B(n_691),
.Y(n_1191)
);

AND2x2_ASAP7_75t_L g1192 ( 
.A(n_1101),
.B(n_691),
.Y(n_1192)
);

AND2x2_ASAP7_75t_L g1193 ( 
.A(n_1091),
.B(n_889),
.Y(n_1193)
);

OAI22xp33_ASAP7_75t_SL g1194 ( 
.A1(n_1138),
.A2(n_649),
.B1(n_667),
.B2(n_662),
.Y(n_1194)
);

OR2x6_ASAP7_75t_L g1195 ( 
.A(n_1120),
.B(n_863),
.Y(n_1195)
);

INVx2_ASAP7_75t_L g1196 ( 
.A(n_1061),
.Y(n_1196)
);

AND2x2_ASAP7_75t_L g1197 ( 
.A(n_1152),
.B(n_896),
.Y(n_1197)
);

AO22x2_ASAP7_75t_L g1198 ( 
.A1(n_1119),
.A2(n_1066),
.B1(n_1075),
.B2(n_1089),
.Y(n_1198)
);

OAI22xp5_ASAP7_75t_L g1199 ( 
.A1(n_1090),
.A2(n_946),
.B1(n_757),
.B2(n_791),
.Y(n_1199)
);

INVx1_ASAP7_75t_L g1200 ( 
.A(n_1066),
.Y(n_1200)
);

INVx2_ASAP7_75t_SL g1201 ( 
.A(n_1152),
.Y(n_1201)
);

AO22x2_ASAP7_75t_L g1202 ( 
.A1(n_1075),
.A2(n_1026),
.B1(n_1051),
.B2(n_919),
.Y(n_1202)
);

AND2x2_ASAP7_75t_L g1203 ( 
.A(n_1118),
.B(n_896),
.Y(n_1203)
);

INVx1_ASAP7_75t_L g1204 ( 
.A(n_1116),
.Y(n_1204)
);

OAI22xp33_ASAP7_75t_SL g1205 ( 
.A1(n_1095),
.A2(n_671),
.B1(n_674),
.B2(n_670),
.Y(n_1205)
);

INVx2_ASAP7_75t_L g1206 ( 
.A(n_1084),
.Y(n_1206)
);

OAI22xp33_ASAP7_75t_L g1207 ( 
.A1(n_1106),
.A2(n_1114),
.B1(n_1129),
.B2(n_1122),
.Y(n_1207)
);

AND2x2_ASAP7_75t_L g1208 ( 
.A(n_1141),
.B(n_896),
.Y(n_1208)
);

BUFx3_ASAP7_75t_L g1209 ( 
.A(n_1164),
.Y(n_1209)
);

AOI22xp5_ASAP7_75t_L g1210 ( 
.A1(n_1089),
.A2(n_681),
.B1(n_684),
.B2(n_678),
.Y(n_1210)
);

OAI22xp33_ASAP7_75t_L g1211 ( 
.A1(n_1139),
.A2(n_964),
.B1(n_928),
.B2(n_648),
.Y(n_1211)
);

INVx2_ASAP7_75t_L g1212 ( 
.A(n_1088),
.Y(n_1212)
);

NOR2xp33_ASAP7_75t_L g1213 ( 
.A(n_1076),
.B(n_752),
.Y(n_1213)
);

OAI22xp33_ASAP7_75t_L g1214 ( 
.A1(n_1148),
.A2(n_964),
.B1(n_663),
.B2(n_768),
.Y(n_1214)
);

INVx1_ASAP7_75t_SL g1215 ( 
.A(n_1143),
.Y(n_1215)
);

OAI22xp33_ASAP7_75t_L g1216 ( 
.A1(n_1154),
.A2(n_769),
.B1(n_771),
.B2(n_728),
.Y(n_1216)
);

INVx1_ASAP7_75t_L g1217 ( 
.A(n_1132),
.Y(n_1217)
);

OAI22xp5_ASAP7_75t_SL g1218 ( 
.A1(n_1170),
.A2(n_817),
.B1(n_834),
.B2(n_831),
.Y(n_1218)
);

OAI22xp5_ASAP7_75t_SL g1219 ( 
.A1(n_1098),
.A2(n_846),
.B1(n_857),
.B2(n_841),
.Y(n_1219)
);

CKINVDCx11_ASAP7_75t_R g1220 ( 
.A(n_1134),
.Y(n_1220)
);

AOI22xp5_ASAP7_75t_L g1221 ( 
.A1(n_1099),
.A2(n_688),
.B1(n_696),
.B2(n_692),
.Y(n_1221)
);

AOI22xp5_ASAP7_75t_L g1222 ( 
.A1(n_1099),
.A2(n_701),
.B1(n_706),
.B2(n_702),
.Y(n_1222)
);

INVx2_ASAP7_75t_L g1223 ( 
.A(n_1083),
.Y(n_1223)
);

INVx1_ASAP7_75t_L g1224 ( 
.A(n_1132),
.Y(n_1224)
);

INVx1_ASAP7_75t_L g1225 ( 
.A(n_1155),
.Y(n_1225)
);

BUFx6f_ASAP7_75t_L g1226 ( 
.A(n_1054),
.Y(n_1226)
);

AO22x2_ASAP7_75t_L g1227 ( 
.A1(n_1105),
.A2(n_707),
.B1(n_723),
.B2(n_722),
.Y(n_1227)
);

INVx1_ASAP7_75t_L g1228 ( 
.A(n_1155),
.Y(n_1228)
);

AOI22x1_ASAP7_75t_SL g1229 ( 
.A1(n_1135),
.A2(n_977),
.B1(n_1006),
.B2(n_867),
.Y(n_1229)
);

INVx1_ASAP7_75t_L g1230 ( 
.A(n_1173),
.Y(n_1230)
);

INVx2_ASAP7_75t_SL g1231 ( 
.A(n_1125),
.Y(n_1231)
);

BUFx6f_ASAP7_75t_L g1232 ( 
.A(n_1054),
.Y(n_1232)
);

NAND2xp33_ASAP7_75t_SL g1233 ( 
.A(n_1145),
.B(n_742),
.Y(n_1233)
);

AND2x2_ASAP7_75t_L g1234 ( 
.A(n_1147),
.B(n_1176),
.Y(n_1234)
);

AO22x2_ASAP7_75t_L g1235 ( 
.A1(n_1105),
.A2(n_1044),
.B1(n_1048),
.B2(n_1043),
.Y(n_1235)
);

AO22x2_ASAP7_75t_L g1236 ( 
.A1(n_1109),
.A2(n_1050),
.B1(n_1049),
.B2(n_744),
.Y(n_1236)
);

INVx2_ASAP7_75t_L g1237 ( 
.A(n_1083),
.Y(n_1237)
);

OAI22xp5_ASAP7_75t_L g1238 ( 
.A1(n_1180),
.A2(n_848),
.B1(n_886),
.B2(n_821),
.Y(n_1238)
);

AO22x2_ASAP7_75t_L g1239 ( 
.A1(n_1109),
.A2(n_746),
.B1(n_747),
.B2(n_725),
.Y(n_1239)
);

INVx2_ASAP7_75t_SL g1240 ( 
.A(n_1146),
.Y(n_1240)
);

OAI22xp33_ASAP7_75t_SL g1241 ( 
.A1(n_1055),
.A2(n_709),
.B1(n_718),
.B2(n_708),
.Y(n_1241)
);

NOR2xp33_ASAP7_75t_L g1242 ( 
.A(n_1082),
.B(n_1108),
.Y(n_1242)
);

AO22x2_ASAP7_75t_L g1243 ( 
.A1(n_1173),
.A2(n_760),
.B1(n_762),
.B2(n_751),
.Y(n_1243)
);

INVx2_ASAP7_75t_SL g1244 ( 
.A(n_1087),
.Y(n_1244)
);

INVx2_ASAP7_75t_L g1245 ( 
.A(n_1107),
.Y(n_1245)
);

AO22x2_ASAP7_75t_L g1246 ( 
.A1(n_1177),
.A2(n_789),
.B1(n_799),
.B2(n_786),
.Y(n_1246)
);

OAI22xp33_ASAP7_75t_SL g1247 ( 
.A1(n_1111),
.A2(n_719),
.B1(n_727),
.B2(n_726),
.Y(n_1247)
);

BUFx6f_ASAP7_75t_L g1248 ( 
.A(n_1054),
.Y(n_1248)
);

AND2x2_ASAP7_75t_L g1249 ( 
.A(n_1082),
.B(n_1030),
.Y(n_1249)
);

INVx2_ASAP7_75t_L g1250 ( 
.A(n_1107),
.Y(n_1250)
);

INVx1_ASAP7_75t_L g1251 ( 
.A(n_1177),
.Y(n_1251)
);

INVx1_ASAP7_75t_L g1252 ( 
.A(n_1113),
.Y(n_1252)
);

AND2x2_ASAP7_75t_L g1253 ( 
.A(n_1108),
.B(n_1126),
.Y(n_1253)
);

OAI22xp33_ASAP7_75t_L g1254 ( 
.A1(n_1157),
.A2(n_1031),
.B1(n_1014),
.B2(n_808),
.Y(n_1254)
);

AO22x2_ASAP7_75t_L g1255 ( 
.A1(n_1153),
.A2(n_1033),
.B1(n_814),
.B2(n_815),
.Y(n_1255)
);

OAI22xp33_ASAP7_75t_SL g1256 ( 
.A1(n_1117),
.A2(n_733),
.B1(n_736),
.B2(n_729),
.Y(n_1256)
);

AOI22xp5_ASAP7_75t_L g1257 ( 
.A1(n_1144),
.A2(n_743),
.B1(n_749),
.B2(n_739),
.Y(n_1257)
);

INVx1_ASAP7_75t_L g1258 ( 
.A(n_1127),
.Y(n_1258)
);

INVx2_ASAP7_75t_L g1259 ( 
.A(n_1133),
.Y(n_1259)
);

CKINVDCx6p67_ASAP7_75t_R g1260 ( 
.A(n_1053),
.Y(n_1260)
);

OAI22xp33_ASAP7_75t_SL g1261 ( 
.A1(n_1126),
.A2(n_755),
.B1(n_756),
.B2(n_754),
.Y(n_1261)
);

AOI22xp5_ASAP7_75t_L g1262 ( 
.A1(n_1162),
.A2(n_763),
.B1(n_766),
.B2(n_759),
.Y(n_1262)
);

INVx1_ASAP7_75t_L g1263 ( 
.A(n_1059),
.Y(n_1263)
);

AND2x2_ASAP7_75t_L g1264 ( 
.A(n_1137),
.B(n_1030),
.Y(n_1264)
);

AOI22xp5_ASAP7_75t_L g1265 ( 
.A1(n_1072),
.A2(n_770),
.B1(n_774),
.B2(n_767),
.Y(n_1265)
);

AOI22xp5_ASAP7_75t_L g1266 ( 
.A1(n_1078),
.A2(n_776),
.B1(n_780),
.B2(n_775),
.Y(n_1266)
);

CKINVDCx5p33_ASAP7_75t_R g1267 ( 
.A(n_1087),
.Y(n_1267)
);

AOI22xp5_ASAP7_75t_L g1268 ( 
.A1(n_1067),
.A2(n_782),
.B1(n_790),
.B2(n_781),
.Y(n_1268)
);

OA22x2_ASAP7_75t_L g1269 ( 
.A1(n_1137),
.A2(n_838),
.B1(n_850),
.B2(n_816),
.Y(n_1269)
);

AND2x2_ASAP7_75t_L g1270 ( 
.A(n_1140),
.B(n_1030),
.Y(n_1270)
);

AOI22xp5_ASAP7_75t_L g1271 ( 
.A1(n_1140),
.A2(n_798),
.B1(n_806),
.B2(n_797),
.Y(n_1271)
);

OAI22xp33_ASAP7_75t_SL g1272 ( 
.A1(n_1158),
.A2(n_809),
.B1(n_819),
.B2(n_812),
.Y(n_1272)
);

AND2x2_ASAP7_75t_L g1273 ( 
.A(n_1060),
.B(n_1032),
.Y(n_1273)
);

OAI22xp33_ASAP7_75t_SL g1274 ( 
.A1(n_1161),
.A2(n_822),
.B1(n_830),
.B2(n_825),
.Y(n_1274)
);

OAI22xp33_ASAP7_75t_SL g1275 ( 
.A1(n_1163),
.A2(n_836),
.B1(n_844),
.B2(n_832),
.Y(n_1275)
);

AOI22xp5_ASAP7_75t_L g1276 ( 
.A1(n_1062),
.A2(n_854),
.B1(n_859),
.B2(n_853),
.Y(n_1276)
);

OAI22xp33_ASAP7_75t_L g1277 ( 
.A1(n_1169),
.A2(n_824),
.B1(n_827),
.B2(n_803),
.Y(n_1277)
);

AND2x2_ASAP7_75t_SL g1278 ( 
.A(n_1077),
.B(n_916),
.Y(n_1278)
);

CKINVDCx6p67_ASAP7_75t_R g1279 ( 
.A(n_1179),
.Y(n_1279)
);

INVx2_ASAP7_75t_L g1280 ( 
.A(n_1149),
.Y(n_1280)
);

INVx1_ASAP7_75t_L g1281 ( 
.A(n_1128),
.Y(n_1281)
);

OAI22xp5_ASAP7_75t_L g1282 ( 
.A1(n_1068),
.A2(n_1005),
.B1(n_865),
.B2(n_866),
.Y(n_1282)
);

OAI22xp33_ASAP7_75t_L g1283 ( 
.A1(n_1077),
.A2(n_840),
.B1(n_842),
.B2(n_829),
.Y(n_1283)
);

AO22x2_ASAP7_75t_L g1284 ( 
.A1(n_1128),
.A2(n_856),
.B1(n_858),
.B2(n_852),
.Y(n_1284)
);

INVx2_ASAP7_75t_L g1285 ( 
.A(n_1160),
.Y(n_1285)
);

NAND2xp5_ASAP7_75t_L g1286 ( 
.A(n_1100),
.B(n_1039),
.Y(n_1286)
);

AOI22xp5_ASAP7_75t_L g1287 ( 
.A1(n_1100),
.A2(n_868),
.B1(n_872),
.B2(n_860),
.Y(n_1287)
);

NAND2xp5_ASAP7_75t_SL g1288 ( 
.A(n_1175),
.B(n_632),
.Y(n_1288)
);

AO22x2_ASAP7_75t_L g1289 ( 
.A1(n_1130),
.A2(n_881),
.B1(n_883),
.B2(n_879),
.Y(n_1289)
);

OAI22xp33_ASAP7_75t_SL g1290 ( 
.A1(n_1094),
.A2(n_875),
.B1(n_877),
.B2(n_874),
.Y(n_1290)
);

INVx1_ASAP7_75t_L g1291 ( 
.A(n_1130),
.Y(n_1291)
);

NOR2x1p5_ASAP7_75t_L g1292 ( 
.A(n_1150),
.B(n_905),
.Y(n_1292)
);

AND2x2_ASAP7_75t_L g1293 ( 
.A(n_1150),
.B(n_1032),
.Y(n_1293)
);

AOI22xp5_ASAP7_75t_L g1294 ( 
.A1(n_1073),
.A2(n_880),
.B1(n_888),
.B2(n_878),
.Y(n_1294)
);

AND2x2_ASAP7_75t_L g1295 ( 
.A(n_1166),
.B(n_1032),
.Y(n_1295)
);

BUFx10_ASAP7_75t_L g1296 ( 
.A(n_1079),
.Y(n_1296)
);

INVx2_ASAP7_75t_SL g1297 ( 
.A(n_1167),
.Y(n_1297)
);

CKINVDCx6p67_ASAP7_75t_R g1298 ( 
.A(n_1074),
.Y(n_1298)
);

AO22x2_ASAP7_75t_L g1299 ( 
.A1(n_1166),
.A2(n_895),
.B1(n_906),
.B2(n_884),
.Y(n_1299)
);

BUFx10_ASAP7_75t_L g1300 ( 
.A(n_1085),
.Y(n_1300)
);

AOI22xp5_ASAP7_75t_L g1301 ( 
.A1(n_1093),
.A2(n_892),
.B1(n_893),
.B2(n_891),
.Y(n_1301)
);

OAI22xp33_ASAP7_75t_L g1302 ( 
.A1(n_1094),
.A2(n_918),
.B1(n_920),
.B2(n_913),
.Y(n_1302)
);

AND2x2_ASAP7_75t_L g1303 ( 
.A(n_1102),
.B(n_916),
.Y(n_1303)
);

INVx2_ASAP7_75t_L g1304 ( 
.A(n_1064),
.Y(n_1304)
);

AND2x2_ASAP7_75t_L g1305 ( 
.A(n_1115),
.B(n_938),
.Y(n_1305)
);

OR2x6_ASAP7_75t_L g1306 ( 
.A(n_1057),
.B(n_952),
.Y(n_1306)
);

AO22x2_ASAP7_75t_L g1307 ( 
.A1(n_1074),
.A2(n_1028),
.B1(n_927),
.B2(n_957),
.Y(n_1307)
);

OAI22xp33_ASAP7_75t_SL g1308 ( 
.A1(n_1064),
.A2(n_899),
.B1(n_903),
.B2(n_897),
.Y(n_1308)
);

OAI22xp33_ASAP7_75t_SL g1309 ( 
.A1(n_1064),
.A2(n_909),
.B1(n_914),
.B2(n_907),
.Y(n_1309)
);

AO22x2_ASAP7_75t_L g1310 ( 
.A1(n_1074),
.A2(n_959),
.B1(n_963),
.B2(n_924),
.Y(n_1310)
);

AOI22xp5_ASAP7_75t_L g1311 ( 
.A1(n_1074),
.A2(n_917),
.B1(n_925),
.B2(n_915),
.Y(n_1311)
);

AND2x2_ASAP7_75t_L g1312 ( 
.A(n_1167),
.B(n_938),
.Y(n_1312)
);

AOI22xp5_ASAP7_75t_L g1313 ( 
.A1(n_1167),
.A2(n_932),
.B1(n_934),
.B2(n_929),
.Y(n_1313)
);

AOI22xp5_ASAP7_75t_L g1314 ( 
.A1(n_1167),
.A2(n_940),
.B1(n_943),
.B2(n_937),
.Y(n_1314)
);

AND2x2_ASAP7_75t_L g1315 ( 
.A(n_1065),
.B(n_952),
.Y(n_1315)
);

OAI22xp33_ASAP7_75t_L g1316 ( 
.A1(n_1065),
.A2(n_969),
.B1(n_980),
.B2(n_966),
.Y(n_1316)
);

INVx1_ASAP7_75t_L g1317 ( 
.A(n_1065),
.Y(n_1317)
);

INVx1_ASAP7_75t_L g1318 ( 
.A(n_1069),
.Y(n_1318)
);

AO22x2_ASAP7_75t_L g1319 ( 
.A1(n_1069),
.A2(n_987),
.B1(n_990),
.B2(n_984),
.Y(n_1319)
);

OAI22xp5_ASAP7_75t_SL g1320 ( 
.A1(n_1069),
.A2(n_947),
.B1(n_948),
.B2(n_944),
.Y(n_1320)
);

HB1xp67_ASAP7_75t_L g1321 ( 
.A(n_1070),
.Y(n_1321)
);

AO22x2_ASAP7_75t_L g1322 ( 
.A1(n_1070),
.A2(n_1027),
.B1(n_996),
.B2(n_1004),
.Y(n_1322)
);

OAI22xp33_ASAP7_75t_L g1323 ( 
.A1(n_1070),
.A2(n_1012),
.B1(n_1016),
.B2(n_993),
.Y(n_1323)
);

OAI22xp33_ASAP7_75t_SL g1324 ( 
.A1(n_1080),
.A2(n_960),
.B1(n_961),
.B2(n_954),
.Y(n_1324)
);

OAI22xp33_ASAP7_75t_L g1325 ( 
.A1(n_1080),
.A2(n_1046),
.B1(n_1047),
.B2(n_1045),
.Y(n_1325)
);

OAI22xp33_ASAP7_75t_SL g1326 ( 
.A1(n_1080),
.A2(n_965),
.B1(n_968),
.B2(n_962),
.Y(n_1326)
);

AOI22xp5_ASAP7_75t_L g1327 ( 
.A1(n_1104),
.A2(n_973),
.B1(n_974),
.B2(n_971),
.Y(n_1327)
);

OAI22xp33_ASAP7_75t_SL g1328 ( 
.A1(n_1104),
.A2(n_978),
.B1(n_979),
.B2(n_976),
.Y(n_1328)
);

OAI22xp33_ASAP7_75t_L g1329 ( 
.A1(n_1104),
.A2(n_1037),
.B1(n_1038),
.B2(n_1035),
.Y(n_1329)
);

AO22x2_ASAP7_75t_L g1330 ( 
.A1(n_1121),
.A2(n_1021),
.B1(n_1015),
.B2(n_710),
.Y(n_1330)
);

OAI22xp33_ASAP7_75t_L g1331 ( 
.A1(n_1121),
.A2(n_991),
.B1(n_994),
.B2(n_986),
.Y(n_1331)
);

NAND2xp5_ASAP7_75t_L g1332 ( 
.A(n_1121),
.B(n_998),
.Y(n_1332)
);

AOI22xp5_ASAP7_75t_L g1333 ( 
.A1(n_1131),
.A2(n_1002),
.B1(n_1003),
.B2(n_999),
.Y(n_1333)
);

OAI22xp5_ASAP7_75t_L g1334 ( 
.A1(n_1131),
.A2(n_1020),
.B1(n_1025),
.B2(n_1010),
.Y(n_1334)
);

INVx1_ASAP7_75t_L g1335 ( 
.A(n_1131),
.Y(n_1335)
);

CKINVDCx6p67_ASAP7_75t_R g1336 ( 
.A(n_1156),
.Y(n_1336)
);

AO22x2_ASAP7_75t_L g1337 ( 
.A1(n_1156),
.A2(n_1021),
.B1(n_1015),
.B2(n_724),
.Y(n_1337)
);

AO22x2_ASAP7_75t_L g1338 ( 
.A1(n_1156),
.A2(n_740),
.B1(n_778),
.B2(n_758),
.Y(n_1338)
);

BUFx6f_ASAP7_75t_SL g1339 ( 
.A(n_1057),
.Y(n_1339)
);

OAI22xp33_ASAP7_75t_SL g1340 ( 
.A1(n_1159),
.A2(n_1040),
.B1(n_1041),
.B2(n_1029),
.Y(n_1340)
);

INVx2_ASAP7_75t_SL g1341 ( 
.A(n_1159),
.Y(n_1341)
);

AOI22xp5_ASAP7_75t_L g1342 ( 
.A1(n_1159),
.A2(n_703),
.B1(n_716),
.B2(n_625),
.Y(n_1342)
);

AND2x2_ASAP7_75t_L g1343 ( 
.A(n_1165),
.B(n_951),
.Y(n_1343)
);

INVx3_ASAP7_75t_L g1344 ( 
.A(n_1165),
.Y(n_1344)
);

AND2x2_ASAP7_75t_L g1345 ( 
.A(n_1165),
.B(n_625),
.Y(n_1345)
);

NAND2xp5_ASAP7_75t_SL g1346 ( 
.A(n_1172),
.B(n_635),
.Y(n_1346)
);

INVx2_ASAP7_75t_L g1347 ( 
.A(n_1172),
.Y(n_1347)
);

INVx2_ASAP7_75t_L g1348 ( 
.A(n_1172),
.Y(n_1348)
);

INVx2_ASAP7_75t_L g1349 ( 
.A(n_1174),
.Y(n_1349)
);

AND2x2_ASAP7_75t_L g1350 ( 
.A(n_1174),
.B(n_625),
.Y(n_1350)
);

AOI22xp5_ASAP7_75t_L g1351 ( 
.A1(n_1174),
.A2(n_703),
.B1(n_716),
.B2(n_625),
.Y(n_1351)
);

NOR2xp33_ASAP7_75t_L g1352 ( 
.A(n_1057),
.B(n_787),
.Y(n_1352)
);

AOI22xp5_ASAP7_75t_L g1353 ( 
.A1(n_1081),
.A2(n_716),
.B1(n_732),
.B2(n_703),
.Y(n_1353)
);

AND2x2_ASAP7_75t_L g1354 ( 
.A(n_1178),
.B(n_703),
.Y(n_1354)
);

AOI22xp5_ASAP7_75t_L g1355 ( 
.A1(n_1081),
.A2(n_732),
.B1(n_796),
.B2(n_716),
.Y(n_1355)
);

INVx8_ASAP7_75t_L g1356 ( 
.A(n_1081),
.Y(n_1356)
);

AOI22xp5_ASAP7_75t_L g1357 ( 
.A1(n_1092),
.A2(n_796),
.B1(n_823),
.B2(n_732),
.Y(n_1357)
);

INVx1_ASAP7_75t_L g1358 ( 
.A(n_1092),
.Y(n_1358)
);

AND2x2_ASAP7_75t_L g1359 ( 
.A(n_1092),
.B(n_732),
.Y(n_1359)
);

AOI22xp5_ASAP7_75t_SL g1360 ( 
.A1(n_1096),
.A2(n_650),
.B1(n_652),
.B2(n_639),
.Y(n_1360)
);

NOR2xp33_ASAP7_75t_L g1361 ( 
.A(n_1096),
.B(n_788),
.Y(n_1361)
);

AND2x2_ASAP7_75t_L g1362 ( 
.A(n_1178),
.B(n_796),
.Y(n_1362)
);

AND2x2_ASAP7_75t_L g1363 ( 
.A(n_1178),
.B(n_796),
.Y(n_1363)
);

INVx3_ASAP7_75t_L g1364 ( 
.A(n_1096),
.Y(n_1364)
);

INVx1_ASAP7_75t_L g1365 ( 
.A(n_1097),
.Y(n_1365)
);

INVx2_ASAP7_75t_SL g1366 ( 
.A(n_1171),
.Y(n_1366)
);

OAI22xp33_ASAP7_75t_L g1367 ( 
.A1(n_1097),
.A2(n_970),
.B1(n_823),
.B2(n_804),
.Y(n_1367)
);

INVx2_ASAP7_75t_SL g1368 ( 
.A(n_1171),
.Y(n_1368)
);

AOI22xp5_ASAP7_75t_L g1369 ( 
.A1(n_1097),
.A2(n_970),
.B1(n_823),
.B2(n_811),
.Y(n_1369)
);

INVx1_ASAP7_75t_L g1370 ( 
.A(n_1103),
.Y(n_1370)
);

INVx2_ASAP7_75t_L g1371 ( 
.A(n_1103),
.Y(n_1371)
);

AND2x2_ASAP7_75t_L g1372 ( 
.A(n_1103),
.B(n_823),
.Y(n_1372)
);

OAI22xp33_ASAP7_75t_SL g1373 ( 
.A1(n_1171),
.A2(n_818),
.B1(n_820),
.B2(n_793),
.Y(n_1373)
);

AND2x2_ASAP7_75t_L g1374 ( 
.A(n_1123),
.B(n_970),
.Y(n_1374)
);

INVx2_ASAP7_75t_L g1375 ( 
.A(n_1123),
.Y(n_1375)
);

NAND2xp33_ASAP7_75t_SL g1376 ( 
.A(n_1123),
.B(n_970),
.Y(n_1376)
);

OAI22xp33_ASAP7_75t_L g1377 ( 
.A1(n_1142),
.A2(n_843),
.B1(n_921),
.B2(n_826),
.Y(n_1377)
);

OR2x6_ASAP7_75t_L g1378 ( 
.A(n_1142),
.B(n_930),
.Y(n_1378)
);

AOI22xp5_ASAP7_75t_L g1379 ( 
.A1(n_1142),
.A2(n_950),
.B1(n_956),
.B2(n_935),
.Y(n_1379)
);

AOI22xp5_ASAP7_75t_L g1380 ( 
.A1(n_1151),
.A2(n_982),
.B1(n_967),
.B2(n_657),
.Y(n_1380)
);

AOI22xp5_ASAP7_75t_L g1381 ( 
.A1(n_1151),
.A2(n_664),
.B1(n_668),
.B2(n_655),
.Y(n_1381)
);

OA22x2_ASAP7_75t_L g1382 ( 
.A1(n_1151),
.A2(n_713),
.B1(n_810),
.B2(n_753),
.Y(n_1382)
);

AND2x2_ASAP7_75t_L g1383 ( 
.A(n_1168),
.B(n_677),
.Y(n_1383)
);

INVx2_ASAP7_75t_L g1384 ( 
.A(n_1168),
.Y(n_1384)
);

OAI22xp33_ASAP7_75t_L g1385 ( 
.A1(n_1168),
.A2(n_777),
.B1(n_849),
.B2(n_697),
.Y(n_1385)
);

OAI22xp33_ASAP7_75t_R g1386 ( 
.A1(n_1056),
.A2(n_777),
.B1(n_849),
.B2(n_697),
.Y(n_1386)
);

AO22x2_ASAP7_75t_L g1387 ( 
.A1(n_1136),
.A2(n_882),
.B1(n_876),
.B2(n_989),
.Y(n_1387)
);

AOI22xp5_ASAP7_75t_L g1388 ( 
.A1(n_1056),
.A2(n_685),
.B1(n_689),
.B2(n_683),
.Y(n_1388)
);

AOI22xp5_ASAP7_75t_L g1389 ( 
.A1(n_1056),
.A2(n_698),
.B1(n_699),
.B2(n_695),
.Y(n_1389)
);

OR2x6_ASAP7_75t_L g1390 ( 
.A(n_1120),
.B(n_876),
.Y(n_1390)
);

AND2x2_ASAP7_75t_L g1391 ( 
.A(n_1052),
.B(n_705),
.Y(n_1391)
);

INVx2_ASAP7_75t_L g1392 ( 
.A(n_1112),
.Y(n_1392)
);

AND2x2_ASAP7_75t_L g1393 ( 
.A(n_1052),
.B(n_712),
.Y(n_1393)
);

AOI22xp5_ASAP7_75t_L g1394 ( 
.A1(n_1056),
.A2(n_715),
.B1(n_721),
.B2(n_720),
.Y(n_1394)
);

INVx1_ASAP7_75t_L g1395 ( 
.A(n_1066),
.Y(n_1395)
);

OR2x6_ASAP7_75t_L g1396 ( 
.A(n_1120),
.B(n_882),
.Y(n_1396)
);

AO22x2_ASAP7_75t_L g1397 ( 
.A1(n_1136),
.A2(n_1017),
.B1(n_1007),
.B2(n_41),
.Y(n_1397)
);

NOR2xp33_ASAP7_75t_L g1398 ( 
.A(n_1258),
.B(n_1042),
.Y(n_1398)
);

INVx1_ASAP7_75t_L g1399 ( 
.A(n_1252),
.Y(n_1399)
);

AND2x2_ASAP7_75t_L g1400 ( 
.A(n_1215),
.B(n_1192),
.Y(n_1400)
);

INVx1_ASAP7_75t_L g1401 ( 
.A(n_1253),
.Y(n_1401)
);

INVx1_ASAP7_75t_L g1402 ( 
.A(n_1315),
.Y(n_1402)
);

NOR2xp33_ASAP7_75t_L g1403 ( 
.A(n_1201),
.B(n_730),
.Y(n_1403)
);

BUFx3_ASAP7_75t_L g1404 ( 
.A(n_1209),
.Y(n_1404)
);

XNOR2xp5_ASAP7_75t_L g1405 ( 
.A(n_1199),
.B(n_39),
.Y(n_1405)
);

INVxp33_ASAP7_75t_L g1406 ( 
.A(n_1234),
.Y(n_1406)
);

INVx1_ASAP7_75t_L g1407 ( 
.A(n_1281),
.Y(n_1407)
);

AND2x2_ASAP7_75t_L g1408 ( 
.A(n_1193),
.B(n_1036),
.Y(n_1408)
);

XNOR2xp5_ASAP7_75t_L g1409 ( 
.A(n_1238),
.B(n_39),
.Y(n_1409)
);

NOR2xp33_ASAP7_75t_L g1410 ( 
.A(n_1231),
.B(n_734),
.Y(n_1410)
);

HB1xp67_ASAP7_75t_L g1411 ( 
.A(n_1330),
.Y(n_1411)
);

INVx1_ASAP7_75t_L g1412 ( 
.A(n_1291),
.Y(n_1412)
);

INVx2_ASAP7_75t_L g1413 ( 
.A(n_1345),
.Y(n_1413)
);

INVx1_ASAP7_75t_L g1414 ( 
.A(n_1293),
.Y(n_1414)
);

INVx1_ASAP7_75t_L g1415 ( 
.A(n_1295),
.Y(n_1415)
);

INVx1_ASAP7_75t_L g1416 ( 
.A(n_1186),
.Y(n_1416)
);

AND2x2_ASAP7_75t_L g1417 ( 
.A(n_1203),
.B(n_735),
.Y(n_1417)
);

NOR2xp33_ASAP7_75t_L g1418 ( 
.A(n_1263),
.B(n_1034),
.Y(n_1418)
);

INVxp67_ASAP7_75t_L g1419 ( 
.A(n_1188),
.Y(n_1419)
);

INVx2_ASAP7_75t_L g1420 ( 
.A(n_1350),
.Y(n_1420)
);

INVx2_ASAP7_75t_L g1421 ( 
.A(n_1354),
.Y(n_1421)
);

OR2x2_ASAP7_75t_L g1422 ( 
.A(n_1185),
.B(n_40),
.Y(n_1422)
);

NAND2xp5_ASAP7_75t_L g1423 ( 
.A(n_1200),
.B(n_741),
.Y(n_1423)
);

XOR2x2_ASAP7_75t_L g1424 ( 
.A(n_1187),
.B(n_40),
.Y(n_1424)
);

BUFx6f_ASAP7_75t_L g1425 ( 
.A(n_1298),
.Y(n_1425)
);

INVx2_ASAP7_75t_SL g1426 ( 
.A(n_1197),
.Y(n_1426)
);

OR2x2_ASAP7_75t_L g1427 ( 
.A(n_1181),
.B(n_42),
.Y(n_1427)
);

INVx1_ASAP7_75t_L g1428 ( 
.A(n_1392),
.Y(n_1428)
);

CKINVDCx20_ASAP7_75t_R g1429 ( 
.A(n_1182),
.Y(n_1429)
);

AND2x2_ASAP7_75t_L g1430 ( 
.A(n_1191),
.B(n_745),
.Y(n_1430)
);

CKINVDCx20_ASAP7_75t_R g1431 ( 
.A(n_1219),
.Y(n_1431)
);

NAND2xp33_ASAP7_75t_R g1432 ( 
.A(n_1267),
.B(n_750),
.Y(n_1432)
);

INVx1_ASAP7_75t_L g1433 ( 
.A(n_1284),
.Y(n_1433)
);

INVx1_ASAP7_75t_L g1434 ( 
.A(n_1284),
.Y(n_1434)
);

INVx1_ASAP7_75t_L g1435 ( 
.A(n_1289),
.Y(n_1435)
);

AND2x6_ASAP7_75t_L g1436 ( 
.A(n_1312),
.B(n_855),
.Y(n_1436)
);

INVx1_ASAP7_75t_L g1437 ( 
.A(n_1289),
.Y(n_1437)
);

INVx2_ASAP7_75t_SL g1438 ( 
.A(n_1208),
.Y(n_1438)
);

AND2x2_ASAP7_75t_L g1439 ( 
.A(n_1279),
.B(n_1391),
.Y(n_1439)
);

NAND2xp5_ASAP7_75t_L g1440 ( 
.A(n_1395),
.B(n_764),
.Y(n_1440)
);

XNOR2xp5_ASAP7_75t_L g1441 ( 
.A(n_1189),
.B(n_42),
.Y(n_1441)
);

INVx1_ASAP7_75t_L g1442 ( 
.A(n_1299),
.Y(n_1442)
);

NAND2xp5_ASAP7_75t_SL g1443 ( 
.A(n_1311),
.B(n_765),
.Y(n_1443)
);

INVx2_ASAP7_75t_L g1444 ( 
.A(n_1359),
.Y(n_1444)
);

AND2x2_ASAP7_75t_L g1445 ( 
.A(n_1393),
.B(n_1024),
.Y(n_1445)
);

AND2x2_ASAP7_75t_L g1446 ( 
.A(n_1255),
.B(n_779),
.Y(n_1446)
);

INVx1_ASAP7_75t_L g1447 ( 
.A(n_1299),
.Y(n_1447)
);

INVx1_ASAP7_75t_L g1448 ( 
.A(n_1243),
.Y(n_1448)
);

NOR2xp33_ASAP7_75t_SL g1449 ( 
.A(n_1278),
.B(n_1023),
.Y(n_1449)
);

INVx1_ASAP7_75t_L g1450 ( 
.A(n_1243),
.Y(n_1450)
);

INVx1_ASAP7_75t_L g1451 ( 
.A(n_1246),
.Y(n_1451)
);

NOR2xp67_ASAP7_75t_L g1452 ( 
.A(n_1257),
.B(n_44),
.Y(n_1452)
);

INVxp67_ASAP7_75t_SL g1453 ( 
.A(n_1204),
.Y(n_1453)
);

NAND2xp5_ASAP7_75t_L g1454 ( 
.A(n_1217),
.B(n_784),
.Y(n_1454)
);

INVx1_ASAP7_75t_L g1455 ( 
.A(n_1246),
.Y(n_1455)
);

BUFx6f_ASAP7_75t_SL g1456 ( 
.A(n_1195),
.Y(n_1456)
);

INVx1_ASAP7_75t_L g1457 ( 
.A(n_1224),
.Y(n_1457)
);

NAND2xp5_ASAP7_75t_L g1458 ( 
.A(n_1225),
.B(n_792),
.Y(n_1458)
);

XNOR2x2_ASAP7_75t_L g1459 ( 
.A(n_1190),
.B(n_44),
.Y(n_1459)
);

INVx1_ASAP7_75t_L g1460 ( 
.A(n_1228),
.Y(n_1460)
);

INVx1_ASAP7_75t_L g1461 ( 
.A(n_1230),
.Y(n_1461)
);

INVx1_ASAP7_75t_L g1462 ( 
.A(n_1251),
.Y(n_1462)
);

AND2x2_ASAP7_75t_SL g1463 ( 
.A(n_1286),
.B(n_855),
.Y(n_1463)
);

BUFx8_ASAP7_75t_L g1464 ( 
.A(n_1183),
.Y(n_1464)
);

INVx1_ASAP7_75t_L g1465 ( 
.A(n_1330),
.Y(n_1465)
);

AND2x2_ASAP7_75t_SL g1466 ( 
.A(n_1287),
.B(n_873),
.Y(n_1466)
);

XOR2xp5_ASAP7_75t_L g1467 ( 
.A(n_1229),
.B(n_45),
.Y(n_1467)
);

INVx1_ASAP7_75t_L g1468 ( 
.A(n_1337),
.Y(n_1468)
);

INVx1_ASAP7_75t_L g1469 ( 
.A(n_1337),
.Y(n_1469)
);

INVx1_ASAP7_75t_L g1470 ( 
.A(n_1198),
.Y(n_1470)
);

INVx1_ASAP7_75t_L g1471 ( 
.A(n_1198),
.Y(n_1471)
);

BUFx2_ASAP7_75t_L g1472 ( 
.A(n_1260),
.Y(n_1472)
);

NAND2xp5_ASAP7_75t_L g1473 ( 
.A(n_1292),
.B(n_794),
.Y(n_1473)
);

INVxp33_ASAP7_75t_L g1474 ( 
.A(n_1218),
.Y(n_1474)
);

XOR2xp5_ASAP7_75t_L g1475 ( 
.A(n_1387),
.B(n_45),
.Y(n_1475)
);

NAND2xp5_ASAP7_75t_L g1476 ( 
.A(n_1302),
.B(n_795),
.Y(n_1476)
);

INVx1_ASAP7_75t_L g1477 ( 
.A(n_1227),
.Y(n_1477)
);

NAND2xp5_ASAP7_75t_L g1478 ( 
.A(n_1223),
.B(n_1237),
.Y(n_1478)
);

INVx2_ASAP7_75t_L g1479 ( 
.A(n_1362),
.Y(n_1479)
);

INVx3_ASAP7_75t_L g1480 ( 
.A(n_1306),
.Y(n_1480)
);

INVx1_ASAP7_75t_L g1481 ( 
.A(n_1227),
.Y(n_1481)
);

INVx1_ASAP7_75t_L g1482 ( 
.A(n_1235),
.Y(n_1482)
);

AND2x2_ASAP7_75t_L g1483 ( 
.A(n_1255),
.B(n_1022),
.Y(n_1483)
);

CKINVDCx5p33_ASAP7_75t_R g1484 ( 
.A(n_1220),
.Y(n_1484)
);

CKINVDCx20_ASAP7_75t_R g1485 ( 
.A(n_1233),
.Y(n_1485)
);

AND2x2_ASAP7_75t_L g1486 ( 
.A(n_1195),
.B(n_800),
.Y(n_1486)
);

INVx1_ASAP7_75t_L g1487 ( 
.A(n_1235),
.Y(n_1487)
);

AND2x2_ASAP7_75t_L g1488 ( 
.A(n_1273),
.B(n_1019),
.Y(n_1488)
);

XNOR2x2_ASAP7_75t_L g1489 ( 
.A(n_1190),
.B(n_1397),
.Y(n_1489)
);

NOR2xp67_ASAP7_75t_L g1490 ( 
.A(n_1262),
.B(n_47),
.Y(n_1490)
);

INVx1_ASAP7_75t_L g1491 ( 
.A(n_1236),
.Y(n_1491)
);

INVx1_ASAP7_75t_L g1492 ( 
.A(n_1236),
.Y(n_1492)
);

INVx1_ASAP7_75t_L g1493 ( 
.A(n_1239),
.Y(n_1493)
);

INVx1_ASAP7_75t_L g1494 ( 
.A(n_1239),
.Y(n_1494)
);

INVxp33_ASAP7_75t_L g1495 ( 
.A(n_1249),
.Y(n_1495)
);

INVx3_ASAP7_75t_L g1496 ( 
.A(n_1306),
.Y(n_1496)
);

INVx1_ASAP7_75t_L g1497 ( 
.A(n_1264),
.Y(n_1497)
);

INVxp33_ASAP7_75t_L g1498 ( 
.A(n_1270),
.Y(n_1498)
);

INVx1_ASAP7_75t_L g1499 ( 
.A(n_1242),
.Y(n_1499)
);

INVx1_ASAP7_75t_L g1500 ( 
.A(n_1336),
.Y(n_1500)
);

AND2x2_ASAP7_75t_L g1501 ( 
.A(n_1390),
.B(n_1013),
.Y(n_1501)
);

CKINVDCx20_ASAP7_75t_R g1502 ( 
.A(n_1282),
.Y(n_1502)
);

INVx1_ASAP7_75t_L g1503 ( 
.A(n_1303),
.Y(n_1503)
);

INVx1_ASAP7_75t_SL g1504 ( 
.A(n_1307),
.Y(n_1504)
);

AND2x2_ASAP7_75t_L g1505 ( 
.A(n_1390),
.B(n_1396),
.Y(n_1505)
);

AND2x6_ASAP7_75t_L g1506 ( 
.A(n_1307),
.B(n_873),
.Y(n_1506)
);

INVx1_ASAP7_75t_L g1507 ( 
.A(n_1305),
.Y(n_1507)
);

NOR2xp33_ASAP7_75t_L g1508 ( 
.A(n_1213),
.B(n_802),
.Y(n_1508)
);

INVx1_ASAP7_75t_L g1509 ( 
.A(n_1319),
.Y(n_1509)
);

INVx1_ASAP7_75t_L g1510 ( 
.A(n_1319),
.Y(n_1510)
);

OAI21xp5_ASAP7_75t_L g1511 ( 
.A1(n_1245),
.A2(n_807),
.B(n_805),
.Y(n_1511)
);

INVx1_ASAP7_75t_L g1512 ( 
.A(n_1322),
.Y(n_1512)
);

BUFx3_ASAP7_75t_L g1513 ( 
.A(n_1396),
.Y(n_1513)
);

INVx1_ASAP7_75t_L g1514 ( 
.A(n_1322),
.Y(n_1514)
);

INVx1_ASAP7_75t_L g1515 ( 
.A(n_1343),
.Y(n_1515)
);

XOR2xp5_ASAP7_75t_L g1516 ( 
.A(n_1387),
.B(n_49),
.Y(n_1516)
);

CKINVDCx20_ASAP7_75t_R g1517 ( 
.A(n_1244),
.Y(n_1517)
);

NOR2xp33_ASAP7_75t_L g1518 ( 
.A(n_1240),
.B(n_1296),
.Y(n_1518)
);

INVx1_ASAP7_75t_L g1519 ( 
.A(n_1382),
.Y(n_1519)
);

CKINVDCx20_ASAP7_75t_R g1520 ( 
.A(n_1320),
.Y(n_1520)
);

XOR2xp5_ASAP7_75t_L g1521 ( 
.A(n_1184),
.B(n_49),
.Y(n_1521)
);

NOR2xp33_ASAP7_75t_L g1522 ( 
.A(n_1300),
.B(n_833),
.Y(n_1522)
);

INVx2_ASAP7_75t_L g1523 ( 
.A(n_1363),
.Y(n_1523)
);

AND2x2_ASAP7_75t_L g1524 ( 
.A(n_1265),
.B(n_1011),
.Y(n_1524)
);

INVx1_ASAP7_75t_L g1525 ( 
.A(n_1269),
.Y(n_1525)
);

AND2x4_ASAP7_75t_L g1526 ( 
.A(n_1210),
.B(n_835),
.Y(n_1526)
);

INVx1_ASAP7_75t_L g1527 ( 
.A(n_1383),
.Y(n_1527)
);

NOR2xp33_ASAP7_75t_L g1528 ( 
.A(n_1221),
.B(n_839),
.Y(n_1528)
);

INVx1_ASAP7_75t_L g1529 ( 
.A(n_1310),
.Y(n_1529)
);

INVx1_ASAP7_75t_L g1530 ( 
.A(n_1310),
.Y(n_1530)
);

INVx1_ASAP7_75t_L g1531 ( 
.A(n_1321),
.Y(n_1531)
);

INVx1_ASAP7_75t_L g1532 ( 
.A(n_1372),
.Y(n_1532)
);

INVxp33_ASAP7_75t_L g1533 ( 
.A(n_1202),
.Y(n_1533)
);

HB1xp67_ASAP7_75t_L g1534 ( 
.A(n_1202),
.Y(n_1534)
);

INVx1_ASAP7_75t_L g1535 ( 
.A(n_1374),
.Y(n_1535)
);

CKINVDCx5p33_ASAP7_75t_R g1536 ( 
.A(n_1388),
.Y(n_1536)
);

INVx1_ASAP7_75t_L g1537 ( 
.A(n_1332),
.Y(n_1537)
);

NOR2xp33_ASAP7_75t_L g1538 ( 
.A(n_1222),
.B(n_847),
.Y(n_1538)
);

INVx1_ASAP7_75t_L g1539 ( 
.A(n_1342),
.Y(n_1539)
);

INVx1_ASAP7_75t_L g1540 ( 
.A(n_1351),
.Y(n_1540)
);

NAND2x1p5_ASAP7_75t_L g1541 ( 
.A(n_1360),
.B(n_1313),
.Y(n_1541)
);

INVx1_ASAP7_75t_L g1542 ( 
.A(n_1316),
.Y(n_1542)
);

NAND2xp5_ASAP7_75t_SL g1543 ( 
.A(n_1314),
.B(n_1283),
.Y(n_1543)
);

NOR2xp33_ASAP7_75t_SL g1544 ( 
.A(n_1297),
.B(n_861),
.Y(n_1544)
);

NAND2xp5_ASAP7_75t_SL g1545 ( 
.A(n_1389),
.B(n_864),
.Y(n_1545)
);

INVx1_ASAP7_75t_L g1546 ( 
.A(n_1323),
.Y(n_1546)
);

INVx1_ASAP7_75t_L g1547 ( 
.A(n_1352),
.Y(n_1547)
);

INVx1_ASAP7_75t_L g1548 ( 
.A(n_1361),
.Y(n_1548)
);

INVx1_ASAP7_75t_L g1549 ( 
.A(n_1379),
.Y(n_1549)
);

INVx1_ASAP7_75t_L g1550 ( 
.A(n_1338),
.Y(n_1550)
);

INVx1_ASAP7_75t_L g1551 ( 
.A(n_1338),
.Y(n_1551)
);

XOR2xp5_ASAP7_75t_SL g1552 ( 
.A(n_1386),
.B(n_50),
.Y(n_1552)
);

INVx1_ASAP7_75t_L g1553 ( 
.A(n_1317),
.Y(n_1553)
);

INVx1_ASAP7_75t_L g1554 ( 
.A(n_1318),
.Y(n_1554)
);

OR2x2_ASAP7_75t_L g1555 ( 
.A(n_1211),
.B(n_50),
.Y(n_1555)
);

NAND2xp33_ASAP7_75t_R g1556 ( 
.A(n_1378),
.B(n_869),
.Y(n_1556)
);

INVx1_ASAP7_75t_L g1557 ( 
.A(n_1335),
.Y(n_1557)
);

AND2x2_ASAP7_75t_L g1558 ( 
.A(n_1266),
.B(n_871),
.Y(n_1558)
);

AND2x2_ASAP7_75t_L g1559 ( 
.A(n_1271),
.B(n_885),
.Y(n_1559)
);

INVx1_ASAP7_75t_L g1560 ( 
.A(n_1385),
.Y(n_1560)
);

INVx2_ASAP7_75t_L g1561 ( 
.A(n_1304),
.Y(n_1561)
);

AND2x4_ASAP7_75t_L g1562 ( 
.A(n_1327),
.B(n_908),
.Y(n_1562)
);

AND2x2_ASAP7_75t_L g1563 ( 
.A(n_1276),
.B(n_910),
.Y(n_1563)
);

INVx1_ASAP7_75t_L g1564 ( 
.A(n_1277),
.Y(n_1564)
);

INVx1_ASAP7_75t_L g1565 ( 
.A(n_1290),
.Y(n_1565)
);

INVx1_ASAP7_75t_L g1566 ( 
.A(n_1377),
.Y(n_1566)
);

CKINVDCx16_ASAP7_75t_R g1567 ( 
.A(n_1394),
.Y(n_1567)
);

INVx1_ASAP7_75t_L g1568 ( 
.A(n_1373),
.Y(n_1568)
);

INVx1_ASAP7_75t_L g1569 ( 
.A(n_1380),
.Y(n_1569)
);

INVx1_ASAP7_75t_L g1570 ( 
.A(n_1241),
.Y(n_1570)
);

INVx1_ASAP7_75t_L g1571 ( 
.A(n_1344),
.Y(n_1571)
);

AND2x4_ASAP7_75t_L g1572 ( 
.A(n_1333),
.B(n_1268),
.Y(n_1572)
);

NOR2xp33_ASAP7_75t_L g1573 ( 
.A(n_1294),
.B(n_912),
.Y(n_1573)
);

BUFx6f_ASAP7_75t_L g1574 ( 
.A(n_1378),
.Y(n_1574)
);

INVx2_ASAP7_75t_L g1575 ( 
.A(n_1347),
.Y(n_1575)
);

INVx1_ASAP7_75t_L g1576 ( 
.A(n_1259),
.Y(n_1576)
);

OR2x2_ASAP7_75t_L g1577 ( 
.A(n_1214),
.B(n_51),
.Y(n_1577)
);

INVx1_ASAP7_75t_L g1578 ( 
.A(n_1280),
.Y(n_1578)
);

NOR2xp67_ASAP7_75t_L g1579 ( 
.A(n_1301),
.B(n_52),
.Y(n_1579)
);

INVx2_ASAP7_75t_L g1580 ( 
.A(n_1348),
.Y(n_1580)
);

BUFx3_ASAP7_75t_L g1581 ( 
.A(n_1341),
.Y(n_1581)
);

NOR2xp33_ASAP7_75t_SL g1582 ( 
.A(n_1207),
.B(n_923),
.Y(n_1582)
);

AND2x4_ASAP7_75t_L g1583 ( 
.A(n_1346),
.B(n_931),
.Y(n_1583)
);

INVx1_ASAP7_75t_L g1584 ( 
.A(n_1285),
.Y(n_1584)
);

NAND2xp5_ASAP7_75t_L g1585 ( 
.A(n_1250),
.B(n_933),
.Y(n_1585)
);

XNOR2xp5_ASAP7_75t_L g1586 ( 
.A(n_1216),
.B(n_52),
.Y(n_1586)
);

CKINVDCx20_ASAP7_75t_R g1587 ( 
.A(n_1334),
.Y(n_1587)
);

AND2x2_ASAP7_75t_L g1588 ( 
.A(n_1184),
.B(n_939),
.Y(n_1588)
);

CKINVDCx20_ASAP7_75t_R g1589 ( 
.A(n_1381),
.Y(n_1589)
);

INVx3_ASAP7_75t_L g1590 ( 
.A(n_1349),
.Y(n_1590)
);

NOR2xp33_ASAP7_75t_L g1591 ( 
.A(n_1288),
.B(n_1325),
.Y(n_1591)
);

INVx1_ASAP7_75t_L g1592 ( 
.A(n_1308),
.Y(n_1592)
);

NAND2x1p5_ASAP7_75t_L g1593 ( 
.A(n_1369),
.B(n_873),
.Y(n_1593)
);

INVx1_ASAP7_75t_L g1594 ( 
.A(n_1309),
.Y(n_1594)
);

NOR2xp67_ASAP7_75t_L g1595 ( 
.A(n_1353),
.B(n_53),
.Y(n_1595)
);

CKINVDCx20_ASAP7_75t_R g1596 ( 
.A(n_1254),
.Y(n_1596)
);

HB1xp67_ASAP7_75t_L g1597 ( 
.A(n_1397),
.Y(n_1597)
);

CKINVDCx20_ASAP7_75t_R g1598 ( 
.A(n_1329),
.Y(n_1598)
);

INVxp33_ASAP7_75t_SL g1599 ( 
.A(n_1194),
.Y(n_1599)
);

INVx1_ASAP7_75t_L g1600 ( 
.A(n_1324),
.Y(n_1600)
);

INVx1_ASAP7_75t_L g1601 ( 
.A(n_1326),
.Y(n_1601)
);

CKINVDCx20_ASAP7_75t_R g1602 ( 
.A(n_1331),
.Y(n_1602)
);

AND2x2_ASAP7_75t_L g1603 ( 
.A(n_1196),
.B(n_942),
.Y(n_1603)
);

INVx1_ASAP7_75t_L g1604 ( 
.A(n_1328),
.Y(n_1604)
);

AND2x2_ASAP7_75t_L g1605 ( 
.A(n_1206),
.B(n_949),
.Y(n_1605)
);

XOR2xp5_ASAP7_75t_L g1606 ( 
.A(n_1205),
.B(n_53),
.Y(n_1606)
);

INVx1_ASAP7_75t_L g1607 ( 
.A(n_1340),
.Y(n_1607)
);

INVx1_ASAP7_75t_L g1608 ( 
.A(n_1261),
.Y(n_1608)
);

INVx1_ASAP7_75t_L g1609 ( 
.A(n_1272),
.Y(n_1609)
);

AND2x2_ASAP7_75t_L g1610 ( 
.A(n_1212),
.B(n_955),
.Y(n_1610)
);

INVx1_ASAP7_75t_L g1611 ( 
.A(n_1274),
.Y(n_1611)
);

INVx1_ASAP7_75t_L g1612 ( 
.A(n_1275),
.Y(n_1612)
);

INVx1_ASAP7_75t_L g1613 ( 
.A(n_1247),
.Y(n_1613)
);

INVx1_ASAP7_75t_L g1614 ( 
.A(n_1256),
.Y(n_1614)
);

INVx1_ASAP7_75t_L g1615 ( 
.A(n_1339),
.Y(n_1615)
);

OAI21xp5_ASAP7_75t_L g1616 ( 
.A1(n_1355),
.A2(n_975),
.B(n_972),
.Y(n_1616)
);

NOR2xp67_ASAP7_75t_L g1617 ( 
.A(n_1357),
.B(n_54),
.Y(n_1617)
);

NOR2xp33_ASAP7_75t_L g1618 ( 
.A(n_1367),
.B(n_981),
.Y(n_1618)
);

INVx1_ASAP7_75t_L g1619 ( 
.A(n_1356),
.Y(n_1619)
);

INVx2_ASAP7_75t_SL g1620 ( 
.A(n_1356),
.Y(n_1620)
);

INVx1_ASAP7_75t_L g1621 ( 
.A(n_1366),
.Y(n_1621)
);

INVxp67_ASAP7_75t_SL g1622 ( 
.A(n_1364),
.Y(n_1622)
);

INVx1_ASAP7_75t_L g1623 ( 
.A(n_1368),
.Y(n_1623)
);

CKINVDCx20_ASAP7_75t_R g1624 ( 
.A(n_1376),
.Y(n_1624)
);

INVx1_ASAP7_75t_L g1625 ( 
.A(n_1358),
.Y(n_1625)
);

CKINVDCx5p33_ASAP7_75t_R g1626 ( 
.A(n_1226),
.Y(n_1626)
);

AND2x2_ASAP7_75t_L g1627 ( 
.A(n_1365),
.B(n_983),
.Y(n_1627)
);

INVx1_ASAP7_75t_L g1628 ( 
.A(n_1370),
.Y(n_1628)
);

NOR2xp33_ASAP7_75t_L g1629 ( 
.A(n_1371),
.B(n_985),
.Y(n_1629)
);

INVx1_ASAP7_75t_L g1630 ( 
.A(n_1384),
.Y(n_1630)
);

INVx1_ASAP7_75t_L g1631 ( 
.A(n_1375),
.Y(n_1631)
);

INVx1_ASAP7_75t_L g1632 ( 
.A(n_1226),
.Y(n_1632)
);

NOR2xp33_ASAP7_75t_L g1633 ( 
.A(n_1232),
.B(n_995),
.Y(n_1633)
);

AOI21x1_ASAP7_75t_L g1634 ( 
.A1(n_1232),
.A2(n_958),
.B(n_711),
.Y(n_1634)
);

INVxp33_ASAP7_75t_L g1635 ( 
.A(n_1248),
.Y(n_1635)
);

AND2x2_ASAP7_75t_L g1636 ( 
.A(n_1248),
.B(n_997),
.Y(n_1636)
);

INVx1_ASAP7_75t_L g1637 ( 
.A(n_1252),
.Y(n_1637)
);

AOI21xp5_ASAP7_75t_L g1638 ( 
.A1(n_1258),
.A2(n_1008),
.B(n_904),
.Y(n_1638)
);

AND2x2_ASAP7_75t_L g1639 ( 
.A(n_1215),
.B(n_711),
.Y(n_1639)
);

NOR2xp33_ASAP7_75t_L g1640 ( 
.A(n_1258),
.B(n_873),
.Y(n_1640)
);

CKINVDCx16_ASAP7_75t_R g1641 ( 
.A(n_1199),
.Y(n_1641)
);

INVx1_ASAP7_75t_L g1642 ( 
.A(n_1252),
.Y(n_1642)
);

INVx1_ASAP7_75t_L g1643 ( 
.A(n_1252),
.Y(n_1643)
);

NOR2xp33_ASAP7_75t_L g1644 ( 
.A(n_1258),
.B(n_904),
.Y(n_1644)
);

NAND2x1p5_ASAP7_75t_L g1645 ( 
.A(n_1244),
.B(n_904),
.Y(n_1645)
);

NAND2xp5_ASAP7_75t_L g1646 ( 
.A(n_1258),
.B(n_711),
.Y(n_1646)
);

INVx1_ASAP7_75t_L g1647 ( 
.A(n_1252),
.Y(n_1647)
);

NAND2xp5_ASAP7_75t_L g1648 ( 
.A(n_1258),
.B(n_958),
.Y(n_1648)
);

BUFx6f_ASAP7_75t_L g1649 ( 
.A(n_1298),
.Y(n_1649)
);

OR2x6_ASAP7_75t_L g1650 ( 
.A(n_1195),
.B(n_904),
.Y(n_1650)
);

NOR2xp33_ASAP7_75t_L g1651 ( 
.A(n_1258),
.B(n_1009),
.Y(n_1651)
);

XOR2xp5_ASAP7_75t_L g1652 ( 
.A(n_1199),
.B(n_54),
.Y(n_1652)
);

INVx1_ASAP7_75t_L g1653 ( 
.A(n_1252),
.Y(n_1653)
);

XNOR2xp5_ASAP7_75t_L g1654 ( 
.A(n_1199),
.B(n_55),
.Y(n_1654)
);

INVx1_ASAP7_75t_L g1655 ( 
.A(n_1252),
.Y(n_1655)
);

INVx2_ASAP7_75t_L g1656 ( 
.A(n_1345),
.Y(n_1656)
);

INVx1_ASAP7_75t_L g1657 ( 
.A(n_1252),
.Y(n_1657)
);

AND2x2_ASAP7_75t_L g1658 ( 
.A(n_1215),
.B(n_958),
.Y(n_1658)
);

XOR2xp5_ASAP7_75t_L g1659 ( 
.A(n_1199),
.B(n_56),
.Y(n_1659)
);

NOR2xp33_ASAP7_75t_L g1660 ( 
.A(n_1258),
.B(n_1009),
.Y(n_1660)
);

AND2x2_ASAP7_75t_L g1661 ( 
.A(n_1215),
.B(n_958),
.Y(n_1661)
);

INVx2_ASAP7_75t_L g1662 ( 
.A(n_1345),
.Y(n_1662)
);

INVx1_ASAP7_75t_L g1663 ( 
.A(n_1252),
.Y(n_1663)
);

XOR2xp5_ASAP7_75t_L g1664 ( 
.A(n_1199),
.B(n_57),
.Y(n_1664)
);

INVx1_ASAP7_75t_L g1665 ( 
.A(n_1252),
.Y(n_1665)
);

INVx2_ASAP7_75t_SL g1666 ( 
.A(n_1215),
.Y(n_1666)
);

NOR2xp33_ASAP7_75t_L g1667 ( 
.A(n_1258),
.B(n_1009),
.Y(n_1667)
);

AND2x2_ASAP7_75t_L g1668 ( 
.A(n_1215),
.B(n_958),
.Y(n_1668)
);

INVx1_ASAP7_75t_L g1669 ( 
.A(n_1252),
.Y(n_1669)
);

NAND2xp5_ASAP7_75t_L g1670 ( 
.A(n_1258),
.B(n_958),
.Y(n_1670)
);

CKINVDCx20_ASAP7_75t_R g1671 ( 
.A(n_1238),
.Y(n_1671)
);

INVx1_ASAP7_75t_L g1672 ( 
.A(n_1252),
.Y(n_1672)
);

NOR2xp33_ASAP7_75t_L g1673 ( 
.A(n_1258),
.B(n_1009),
.Y(n_1673)
);

INVx1_ASAP7_75t_L g1674 ( 
.A(n_1252),
.Y(n_1674)
);

INVx1_ASAP7_75t_L g1675 ( 
.A(n_1252),
.Y(n_1675)
);

INVx2_ASAP7_75t_L g1676 ( 
.A(n_1345),
.Y(n_1676)
);

XOR2xp5_ASAP7_75t_L g1677 ( 
.A(n_1199),
.B(n_57),
.Y(n_1677)
);

NOR2xp33_ASAP7_75t_L g1678 ( 
.A(n_1258),
.B(n_958),
.Y(n_1678)
);

INVx2_ASAP7_75t_SL g1679 ( 
.A(n_1215),
.Y(n_1679)
);

AND2x2_ASAP7_75t_L g1680 ( 
.A(n_1215),
.B(n_58),
.Y(n_1680)
);

NOR2xp33_ASAP7_75t_L g1681 ( 
.A(n_1258),
.B(n_414),
.Y(n_1681)
);

INVx2_ASAP7_75t_L g1682 ( 
.A(n_1345),
.Y(n_1682)
);

INVx3_ASAP7_75t_L g1683 ( 
.A(n_1306),
.Y(n_1683)
);

INVx1_ASAP7_75t_L g1684 ( 
.A(n_1252),
.Y(n_1684)
);

INVx1_ASAP7_75t_L g1685 ( 
.A(n_1252),
.Y(n_1685)
);

INVx2_ASAP7_75t_L g1686 ( 
.A(n_1345),
.Y(n_1686)
);

XOR2x2_ASAP7_75t_L g1687 ( 
.A(n_1187),
.B(n_59),
.Y(n_1687)
);

INVx1_ASAP7_75t_L g1688 ( 
.A(n_1252),
.Y(n_1688)
);

AND2x2_ASAP7_75t_L g1689 ( 
.A(n_1215),
.B(n_60),
.Y(n_1689)
);

INVx2_ASAP7_75t_L g1690 ( 
.A(n_1345),
.Y(n_1690)
);

INVx3_ASAP7_75t_L g1691 ( 
.A(n_1574),
.Y(n_1691)
);

AOI22xp5_ASAP7_75t_L g1692 ( 
.A1(n_1666),
.A2(n_63),
.B1(n_61),
.B2(n_62),
.Y(n_1692)
);

INVx1_ASAP7_75t_L g1693 ( 
.A(n_1401),
.Y(n_1693)
);

OAI21xp5_ASAP7_75t_L g1694 ( 
.A1(n_1478),
.A2(n_419),
.B(n_418),
.Y(n_1694)
);

AND2x6_ASAP7_75t_L g1695 ( 
.A(n_1504),
.B(n_1574),
.Y(n_1695)
);

AND2x2_ASAP7_75t_L g1696 ( 
.A(n_1679),
.B(n_61),
.Y(n_1696)
);

NAND2xp5_ASAP7_75t_L g1697 ( 
.A(n_1453),
.B(n_64),
.Y(n_1697)
);

INVx2_ASAP7_75t_SL g1698 ( 
.A(n_1574),
.Y(n_1698)
);

INVx2_ASAP7_75t_L g1699 ( 
.A(n_1576),
.Y(n_1699)
);

INVx1_ASAP7_75t_L g1700 ( 
.A(n_1497),
.Y(n_1700)
);

AND2x2_ASAP7_75t_L g1701 ( 
.A(n_1400),
.B(n_65),
.Y(n_1701)
);

AND2x2_ASAP7_75t_L g1702 ( 
.A(n_1453),
.B(n_65),
.Y(n_1702)
);

INVx2_ASAP7_75t_L g1703 ( 
.A(n_1578),
.Y(n_1703)
);

NAND2xp5_ASAP7_75t_SL g1704 ( 
.A(n_1509),
.B(n_420),
.Y(n_1704)
);

NAND2xp5_ASAP7_75t_L g1705 ( 
.A(n_1414),
.B(n_66),
.Y(n_1705)
);

NOR2xp33_ASAP7_75t_L g1706 ( 
.A(n_1415),
.B(n_66),
.Y(n_1706)
);

AND2x2_ASAP7_75t_SL g1707 ( 
.A(n_1449),
.B(n_67),
.Y(n_1707)
);

HB1xp67_ASAP7_75t_L g1708 ( 
.A(n_1411),
.Y(n_1708)
);

BUFx3_ASAP7_75t_L g1709 ( 
.A(n_1425),
.Y(n_1709)
);

INVx4_ASAP7_75t_L g1710 ( 
.A(n_1506),
.Y(n_1710)
);

AND2x2_ASAP7_75t_L g1711 ( 
.A(n_1439),
.B(n_67),
.Y(n_1711)
);

AND2x2_ASAP7_75t_L g1712 ( 
.A(n_1406),
.B(n_1446),
.Y(n_1712)
);

AND2x2_ASAP7_75t_SL g1713 ( 
.A(n_1449),
.B(n_68),
.Y(n_1713)
);

INVx1_ASAP7_75t_L g1714 ( 
.A(n_1407),
.Y(n_1714)
);

AND2x2_ASAP7_75t_SL g1715 ( 
.A(n_1411),
.B(n_68),
.Y(n_1715)
);

INVx3_ASAP7_75t_L g1716 ( 
.A(n_1506),
.Y(n_1716)
);

HB1xp67_ASAP7_75t_L g1717 ( 
.A(n_1650),
.Y(n_1717)
);

NAND2xp5_ASAP7_75t_L g1718 ( 
.A(n_1398),
.B(n_69),
.Y(n_1718)
);

AND2x2_ASAP7_75t_SL g1719 ( 
.A(n_1466),
.B(n_70),
.Y(n_1719)
);

AND2x2_ASAP7_75t_L g1720 ( 
.A(n_1483),
.B(n_70),
.Y(n_1720)
);

INVx1_ASAP7_75t_L g1721 ( 
.A(n_1412),
.Y(n_1721)
);

AND2x2_ASAP7_75t_L g1722 ( 
.A(n_1680),
.B(n_72),
.Y(n_1722)
);

NAND2xp5_ASAP7_75t_SL g1723 ( 
.A(n_1510),
.B(n_421),
.Y(n_1723)
);

AND2x2_ASAP7_75t_L g1724 ( 
.A(n_1689),
.B(n_72),
.Y(n_1724)
);

INVx4_ASAP7_75t_L g1725 ( 
.A(n_1506),
.Y(n_1725)
);

AND2x2_ASAP7_75t_L g1726 ( 
.A(n_1419),
.B(n_74),
.Y(n_1726)
);

HB1xp67_ASAP7_75t_L g1727 ( 
.A(n_1650),
.Y(n_1727)
);

INVx3_ASAP7_75t_L g1728 ( 
.A(n_1506),
.Y(n_1728)
);

NAND2xp5_ASAP7_75t_L g1729 ( 
.A(n_1398),
.B(n_74),
.Y(n_1729)
);

AND2x2_ASAP7_75t_L g1730 ( 
.A(n_1419),
.B(n_75),
.Y(n_1730)
);

HB1xp67_ASAP7_75t_L g1731 ( 
.A(n_1650),
.Y(n_1731)
);

BUFx3_ASAP7_75t_L g1732 ( 
.A(n_1425),
.Y(n_1732)
);

NOR2xp33_ASAP7_75t_L g1733 ( 
.A(n_1495),
.B(n_75),
.Y(n_1733)
);

AND2x2_ASAP7_75t_L g1734 ( 
.A(n_1408),
.B(n_1417),
.Y(n_1734)
);

INVx2_ASAP7_75t_SL g1735 ( 
.A(n_1480),
.Y(n_1735)
);

BUFx6f_ASAP7_75t_L g1736 ( 
.A(n_1425),
.Y(n_1736)
);

INVx2_ASAP7_75t_L g1737 ( 
.A(n_1584),
.Y(n_1737)
);

INVx4_ASAP7_75t_L g1738 ( 
.A(n_1649),
.Y(n_1738)
);

OR2x6_ASAP7_75t_L g1739 ( 
.A(n_1513),
.B(n_76),
.Y(n_1739)
);

INVx3_ASAP7_75t_L g1740 ( 
.A(n_1421),
.Y(n_1740)
);

AND2x2_ASAP7_75t_L g1741 ( 
.A(n_1526),
.B(n_76),
.Y(n_1741)
);

BUFx3_ASAP7_75t_L g1742 ( 
.A(n_1649),
.Y(n_1742)
);

INVxp67_ASAP7_75t_L g1743 ( 
.A(n_1456),
.Y(n_1743)
);

INVx1_ASAP7_75t_L g1744 ( 
.A(n_1527),
.Y(n_1744)
);

AND2x2_ASAP7_75t_L g1745 ( 
.A(n_1526),
.B(n_77),
.Y(n_1745)
);

INVx2_ASAP7_75t_L g1746 ( 
.A(n_1478),
.Y(n_1746)
);

AND2x2_ASAP7_75t_L g1747 ( 
.A(n_1438),
.B(n_77),
.Y(n_1747)
);

BUFx6f_ASAP7_75t_L g1748 ( 
.A(n_1649),
.Y(n_1748)
);

AND2x2_ASAP7_75t_L g1749 ( 
.A(n_1488),
.B(n_1498),
.Y(n_1749)
);

HB1xp67_ASAP7_75t_L g1750 ( 
.A(n_1504),
.Y(n_1750)
);

INVx2_ASAP7_75t_L g1751 ( 
.A(n_1416),
.Y(n_1751)
);

INVx1_ASAP7_75t_L g1752 ( 
.A(n_1457),
.Y(n_1752)
);

OAI21xp33_ASAP7_75t_L g1753 ( 
.A1(n_1582),
.A2(n_79),
.B(n_80),
.Y(n_1753)
);

NAND2xp5_ASAP7_75t_L g1754 ( 
.A(n_1564),
.B(n_80),
.Y(n_1754)
);

AND2x2_ASAP7_75t_SL g1755 ( 
.A(n_1463),
.B(n_81),
.Y(n_1755)
);

AND3x1_ASAP7_75t_SL g1756 ( 
.A(n_1609),
.B(n_82),
.C(n_86),
.Y(n_1756)
);

NAND2x1p5_ASAP7_75t_L g1757 ( 
.A(n_1480),
.B(n_1683),
.Y(n_1757)
);

HB1xp67_ASAP7_75t_L g1758 ( 
.A(n_1404),
.Y(n_1758)
);

INVx1_ASAP7_75t_L g1759 ( 
.A(n_1460),
.Y(n_1759)
);

NAND2xp5_ASAP7_75t_L g1760 ( 
.A(n_1461),
.B(n_82),
.Y(n_1760)
);

BUFx3_ASAP7_75t_L g1761 ( 
.A(n_1619),
.Y(n_1761)
);

AND2x2_ASAP7_75t_L g1762 ( 
.A(n_1588),
.B(n_86),
.Y(n_1762)
);

NAND2xp5_ASAP7_75t_SL g1763 ( 
.A(n_1512),
.B(n_615),
.Y(n_1763)
);

AND2x2_ASAP7_75t_L g1764 ( 
.A(n_1524),
.B(n_87),
.Y(n_1764)
);

OAI21xp5_ASAP7_75t_L g1765 ( 
.A1(n_1638),
.A2(n_426),
.B(n_423),
.Y(n_1765)
);

INVx2_ASAP7_75t_SL g1766 ( 
.A(n_1496),
.Y(n_1766)
);

NAND2xp5_ASAP7_75t_L g1767 ( 
.A(n_1462),
.B(n_88),
.Y(n_1767)
);

NOR2xp33_ASAP7_75t_R g1768 ( 
.A(n_1556),
.B(n_1517),
.Y(n_1768)
);

INVx1_ASAP7_75t_L g1769 ( 
.A(n_1399),
.Y(n_1769)
);

INVx3_ASAP7_75t_L g1770 ( 
.A(n_1444),
.Y(n_1770)
);

AND2x2_ASAP7_75t_L g1771 ( 
.A(n_1558),
.B(n_89),
.Y(n_1771)
);

OR2x2_ASAP7_75t_L g1772 ( 
.A(n_1641),
.B(n_90),
.Y(n_1772)
);

INVx2_ASAP7_75t_L g1773 ( 
.A(n_1428),
.Y(n_1773)
);

INVx1_ASAP7_75t_L g1774 ( 
.A(n_1637),
.Y(n_1774)
);

AND2x4_ASAP7_75t_L g1775 ( 
.A(n_1470),
.B(n_90),
.Y(n_1775)
);

AND2x2_ASAP7_75t_L g1776 ( 
.A(n_1445),
.B(n_91),
.Y(n_1776)
);

INVx4_ASAP7_75t_L g1777 ( 
.A(n_1645),
.Y(n_1777)
);

AND2x2_ASAP7_75t_L g1778 ( 
.A(n_1503),
.B(n_91),
.Y(n_1778)
);

INVxp67_ASAP7_75t_L g1779 ( 
.A(n_1456),
.Y(n_1779)
);

INVx1_ASAP7_75t_L g1780 ( 
.A(n_1642),
.Y(n_1780)
);

NAND2xp5_ASAP7_75t_L g1781 ( 
.A(n_1499),
.B(n_93),
.Y(n_1781)
);

NAND2xp5_ASAP7_75t_L g1782 ( 
.A(n_1507),
.B(n_95),
.Y(n_1782)
);

NAND2xp5_ASAP7_75t_L g1783 ( 
.A(n_1569),
.B(n_95),
.Y(n_1783)
);

AND2x4_ASAP7_75t_L g1784 ( 
.A(n_1471),
.B(n_96),
.Y(n_1784)
);

INVx4_ASAP7_75t_L g1785 ( 
.A(n_1645),
.Y(n_1785)
);

INVx2_ASAP7_75t_SL g1786 ( 
.A(n_1496),
.Y(n_1786)
);

INVx2_ASAP7_75t_L g1787 ( 
.A(n_1479),
.Y(n_1787)
);

BUFx3_ASAP7_75t_L g1788 ( 
.A(n_1620),
.Y(n_1788)
);

INVx2_ASAP7_75t_SL g1789 ( 
.A(n_1683),
.Y(n_1789)
);

AND2x4_ASAP7_75t_L g1790 ( 
.A(n_1448),
.B(n_97),
.Y(n_1790)
);

INVx1_ASAP7_75t_SL g1791 ( 
.A(n_1472),
.Y(n_1791)
);

INVx3_ASAP7_75t_L g1792 ( 
.A(n_1523),
.Y(n_1792)
);

AND2x2_ASAP7_75t_L g1793 ( 
.A(n_1563),
.B(n_97),
.Y(n_1793)
);

INVx1_ASAP7_75t_L g1794 ( 
.A(n_1643),
.Y(n_1794)
);

AND2x2_ASAP7_75t_L g1795 ( 
.A(n_1596),
.B(n_98),
.Y(n_1795)
);

AOI22xp5_ASAP7_75t_L g1796 ( 
.A1(n_1572),
.A2(n_101),
.B1(n_98),
.B2(n_99),
.Y(n_1796)
);

INVx2_ASAP7_75t_L g1797 ( 
.A(n_1553),
.Y(n_1797)
);

INVx2_ASAP7_75t_L g1798 ( 
.A(n_1554),
.Y(n_1798)
);

BUFx6f_ASAP7_75t_L g1799 ( 
.A(n_1634),
.Y(n_1799)
);

AND2x2_ASAP7_75t_L g1800 ( 
.A(n_1433),
.B(n_103),
.Y(n_1800)
);

NAND2xp5_ASAP7_75t_L g1801 ( 
.A(n_1542),
.B(n_103),
.Y(n_1801)
);

INVx1_ASAP7_75t_L g1802 ( 
.A(n_1647),
.Y(n_1802)
);

BUFx3_ASAP7_75t_L g1803 ( 
.A(n_1464),
.Y(n_1803)
);

AND2x2_ASAP7_75t_L g1804 ( 
.A(n_1430),
.B(n_104),
.Y(n_1804)
);

AND2x2_ASAP7_75t_L g1805 ( 
.A(n_1559),
.B(n_105),
.Y(n_1805)
);

AND2x2_ASAP7_75t_SL g1806 ( 
.A(n_1597),
.B(n_106),
.Y(n_1806)
);

INVx1_ASAP7_75t_L g1807 ( 
.A(n_1653),
.Y(n_1807)
);

NAND2xp5_ASAP7_75t_SL g1808 ( 
.A(n_1514),
.B(n_610),
.Y(n_1808)
);

AND2x2_ASAP7_75t_L g1809 ( 
.A(n_1597),
.B(n_106),
.Y(n_1809)
);

INVxp67_ASAP7_75t_L g1810 ( 
.A(n_1464),
.Y(n_1810)
);

AND2x2_ASAP7_75t_L g1811 ( 
.A(n_1562),
.B(n_107),
.Y(n_1811)
);

INVx1_ASAP7_75t_L g1812 ( 
.A(n_1655),
.Y(n_1812)
);

AND2x2_ASAP7_75t_SL g1813 ( 
.A(n_1534),
.B(n_108),
.Y(n_1813)
);

INVx1_ASAP7_75t_L g1814 ( 
.A(n_1657),
.Y(n_1814)
);

AND2x4_ASAP7_75t_L g1815 ( 
.A(n_1450),
.B(n_108),
.Y(n_1815)
);

NAND2xp5_ASAP7_75t_L g1816 ( 
.A(n_1546),
.B(n_1663),
.Y(n_1816)
);

AND2x4_ASAP7_75t_L g1817 ( 
.A(n_1451),
.B(n_109),
.Y(n_1817)
);

NAND2xp5_ASAP7_75t_L g1818 ( 
.A(n_1665),
.B(n_109),
.Y(n_1818)
);

INVx2_ASAP7_75t_L g1819 ( 
.A(n_1557),
.Y(n_1819)
);

AND2x2_ASAP7_75t_L g1820 ( 
.A(n_1434),
.B(n_110),
.Y(n_1820)
);

AND2x2_ASAP7_75t_SL g1821 ( 
.A(n_1534),
.B(n_111),
.Y(n_1821)
);

AND2x2_ASAP7_75t_L g1822 ( 
.A(n_1435),
.B(n_111),
.Y(n_1822)
);

AND2x2_ASAP7_75t_L g1823 ( 
.A(n_1437),
.B(n_112),
.Y(n_1823)
);

NOR2xp33_ASAP7_75t_L g1824 ( 
.A(n_1591),
.B(n_112),
.Y(n_1824)
);

INVx1_ASAP7_75t_L g1825 ( 
.A(n_1669),
.Y(n_1825)
);

INVx2_ASAP7_75t_L g1826 ( 
.A(n_1532),
.Y(n_1826)
);

INVx1_ASAP7_75t_SL g1827 ( 
.A(n_1671),
.Y(n_1827)
);

INVxp33_ASAP7_75t_L g1828 ( 
.A(n_1505),
.Y(n_1828)
);

AND2x2_ASAP7_75t_L g1829 ( 
.A(n_1442),
.B(n_113),
.Y(n_1829)
);

AND2x2_ASAP7_75t_L g1830 ( 
.A(n_1562),
.B(n_113),
.Y(n_1830)
);

AND2x2_ASAP7_75t_SL g1831 ( 
.A(n_1529),
.B(n_114),
.Y(n_1831)
);

NAND2xp5_ASAP7_75t_L g1832 ( 
.A(n_1672),
.B(n_1674),
.Y(n_1832)
);

NOR2xp33_ASAP7_75t_R g1833 ( 
.A(n_1484),
.B(n_114),
.Y(n_1833)
);

INVx2_ASAP7_75t_L g1834 ( 
.A(n_1535),
.Y(n_1834)
);

BUFx6f_ASAP7_75t_L g1835 ( 
.A(n_1561),
.Y(n_1835)
);

AND2x4_ASAP7_75t_L g1836 ( 
.A(n_1455),
.B(n_115),
.Y(n_1836)
);

AND2x2_ASAP7_75t_L g1837 ( 
.A(n_1422),
.B(n_115),
.Y(n_1837)
);

OAI21xp5_ASAP7_75t_L g1838 ( 
.A1(n_1638),
.A2(n_434),
.B(n_428),
.Y(n_1838)
);

OAI21xp5_ASAP7_75t_L g1839 ( 
.A1(n_1646),
.A2(n_436),
.B(n_435),
.Y(n_1839)
);

INVx2_ASAP7_75t_SL g1840 ( 
.A(n_1426),
.Y(n_1840)
);

OAI21xp5_ASAP7_75t_L g1841 ( 
.A1(n_1646),
.A2(n_441),
.B(n_439),
.Y(n_1841)
);

AND2x2_ASAP7_75t_L g1842 ( 
.A(n_1533),
.B(n_116),
.Y(n_1842)
);

INVx1_ASAP7_75t_L g1843 ( 
.A(n_1675),
.Y(n_1843)
);

NAND2xp5_ASAP7_75t_L g1844 ( 
.A(n_1684),
.B(n_118),
.Y(n_1844)
);

INVx4_ASAP7_75t_L g1845 ( 
.A(n_1626),
.Y(n_1845)
);

INVx1_ASAP7_75t_L g1846 ( 
.A(n_1685),
.Y(n_1846)
);

AND2x2_ASAP7_75t_L g1847 ( 
.A(n_1486),
.B(n_118),
.Y(n_1847)
);

AND2x2_ASAP7_75t_L g1848 ( 
.A(n_1572),
.B(n_119),
.Y(n_1848)
);

HB1xp67_ASAP7_75t_L g1849 ( 
.A(n_1465),
.Y(n_1849)
);

INVx2_ASAP7_75t_L g1850 ( 
.A(n_1575),
.Y(n_1850)
);

INVx2_ASAP7_75t_L g1851 ( 
.A(n_1580),
.Y(n_1851)
);

AND2x2_ASAP7_75t_L g1852 ( 
.A(n_1502),
.B(n_119),
.Y(n_1852)
);

OR2x2_ASAP7_75t_L g1853 ( 
.A(n_1611),
.B(n_120),
.Y(n_1853)
);

INVx1_ASAP7_75t_L g1854 ( 
.A(n_1688),
.Y(n_1854)
);

AND2x2_ASAP7_75t_L g1855 ( 
.A(n_1501),
.B(n_121),
.Y(n_1855)
);

HB1xp67_ASAP7_75t_L g1856 ( 
.A(n_1468),
.Y(n_1856)
);

INVx1_ASAP7_75t_L g1857 ( 
.A(n_1648),
.Y(n_1857)
);

INVx2_ASAP7_75t_L g1858 ( 
.A(n_1625),
.Y(n_1858)
);

BUFx3_ASAP7_75t_L g1859 ( 
.A(n_1581),
.Y(n_1859)
);

AND2x2_ASAP7_75t_SL g1860 ( 
.A(n_1530),
.B(n_121),
.Y(n_1860)
);

AND2x2_ASAP7_75t_L g1861 ( 
.A(n_1447),
.B(n_1477),
.Y(n_1861)
);

NAND2xp5_ASAP7_75t_L g1862 ( 
.A(n_1639),
.B(n_122),
.Y(n_1862)
);

NAND2x1p5_ASAP7_75t_L g1863 ( 
.A(n_1481),
.B(n_122),
.Y(n_1863)
);

AND2x2_ASAP7_75t_L g1864 ( 
.A(n_1567),
.B(n_124),
.Y(n_1864)
);

AND2x2_ASAP7_75t_L g1865 ( 
.A(n_1612),
.B(n_124),
.Y(n_1865)
);

NAND2xp5_ASAP7_75t_L g1866 ( 
.A(n_1658),
.B(n_125),
.Y(n_1866)
);

INVx1_ASAP7_75t_L g1867 ( 
.A(n_1648),
.Y(n_1867)
);

INVx2_ASAP7_75t_L g1868 ( 
.A(n_1628),
.Y(n_1868)
);

OAI21xp5_ASAP7_75t_L g1869 ( 
.A1(n_1670),
.A2(n_445),
.B(n_444),
.Y(n_1869)
);

NAND2xp5_ASAP7_75t_L g1870 ( 
.A(n_1661),
.B(n_1668),
.Y(n_1870)
);

OR2x2_ASAP7_75t_L g1871 ( 
.A(n_1613),
.B(n_126),
.Y(n_1871)
);

HB1xp67_ASAP7_75t_L g1872 ( 
.A(n_1469),
.Y(n_1872)
);

AND2x2_ASAP7_75t_L g1873 ( 
.A(n_1614),
.B(n_126),
.Y(n_1873)
);

INVx2_ASAP7_75t_L g1874 ( 
.A(n_1413),
.Y(n_1874)
);

INVx1_ASAP7_75t_L g1875 ( 
.A(n_1670),
.Y(n_1875)
);

NAND2xp5_ASAP7_75t_L g1876 ( 
.A(n_1418),
.B(n_127),
.Y(n_1876)
);

HB1xp67_ASAP7_75t_L g1877 ( 
.A(n_1577),
.Y(n_1877)
);

NAND2xp5_ASAP7_75t_L g1878 ( 
.A(n_1418),
.B(n_128),
.Y(n_1878)
);

INVx2_ASAP7_75t_L g1879 ( 
.A(n_1420),
.Y(n_1879)
);

INVx1_ASAP7_75t_SL g1880 ( 
.A(n_1603),
.Y(n_1880)
);

NOR2xp33_ASAP7_75t_L g1881 ( 
.A(n_1592),
.B(n_129),
.Y(n_1881)
);

NAND2xp5_ASAP7_75t_L g1882 ( 
.A(n_1537),
.B(n_129),
.Y(n_1882)
);

NOR2xp33_ASAP7_75t_L g1883 ( 
.A(n_1594),
.B(n_1600),
.Y(n_1883)
);

NAND2xp5_ASAP7_75t_L g1884 ( 
.A(n_1605),
.B(n_130),
.Y(n_1884)
);

INVx2_ASAP7_75t_L g1885 ( 
.A(n_1690),
.Y(n_1885)
);

AND2x2_ASAP7_75t_L g1886 ( 
.A(n_1555),
.B(n_130),
.Y(n_1886)
);

INVx1_ASAP7_75t_L g1887 ( 
.A(n_1515),
.Y(n_1887)
);

AND2x2_ASAP7_75t_L g1888 ( 
.A(n_1608),
.B(n_131),
.Y(n_1888)
);

INVx3_ASAP7_75t_L g1889 ( 
.A(n_1590),
.Y(n_1889)
);

INVx2_ASAP7_75t_L g1890 ( 
.A(n_1656),
.Y(n_1890)
);

OAI21xp5_ASAP7_75t_L g1891 ( 
.A1(n_1678),
.A2(n_448),
.B(n_446),
.Y(n_1891)
);

INVx2_ASAP7_75t_L g1892 ( 
.A(n_1662),
.Y(n_1892)
);

BUFx6f_ASAP7_75t_L g1893 ( 
.A(n_1590),
.Y(n_1893)
);

AND2x4_ASAP7_75t_L g1894 ( 
.A(n_1482),
.B(n_1487),
.Y(n_1894)
);

AND2x2_ASAP7_75t_L g1895 ( 
.A(n_1427),
.B(n_131),
.Y(n_1895)
);

INVx4_ASAP7_75t_L g1896 ( 
.A(n_1436),
.Y(n_1896)
);

AND2x2_ASAP7_75t_L g1897 ( 
.A(n_1522),
.B(n_1409),
.Y(n_1897)
);

INVx2_ASAP7_75t_L g1898 ( 
.A(n_1676),
.Y(n_1898)
);

INVx1_ASAP7_75t_L g1899 ( 
.A(n_1402),
.Y(n_1899)
);

OAI21xp5_ASAP7_75t_L g1900 ( 
.A1(n_1539),
.A2(n_451),
.B(n_449),
.Y(n_1900)
);

AND2x2_ASAP7_75t_L g1901 ( 
.A(n_1565),
.B(n_132),
.Y(n_1901)
);

AND2x2_ASAP7_75t_L g1902 ( 
.A(n_1491),
.B(n_133),
.Y(n_1902)
);

BUFx6f_ASAP7_75t_L g1903 ( 
.A(n_1436),
.Y(n_1903)
);

AND2x2_ASAP7_75t_L g1904 ( 
.A(n_1492),
.B(n_133),
.Y(n_1904)
);

INVx2_ASAP7_75t_L g1905 ( 
.A(n_1682),
.Y(n_1905)
);

NOR2xp33_ASAP7_75t_L g1906 ( 
.A(n_1601),
.B(n_134),
.Y(n_1906)
);

AND2x4_ASAP7_75t_L g1907 ( 
.A(n_1493),
.B(n_136),
.Y(n_1907)
);

OR2x2_ASAP7_75t_SL g1908 ( 
.A(n_1431),
.B(n_136),
.Y(n_1908)
);

NAND2xp5_ASAP7_75t_L g1909 ( 
.A(n_1610),
.B(n_1549),
.Y(n_1909)
);

AND2x2_ASAP7_75t_L g1910 ( 
.A(n_1494),
.B(n_137),
.Y(n_1910)
);

INVxp67_ASAP7_75t_L g1911 ( 
.A(n_1432),
.Y(n_1911)
);

INVx2_ASAP7_75t_L g1912 ( 
.A(n_1686),
.Y(n_1912)
);

INVx3_ASAP7_75t_L g1913 ( 
.A(n_1436),
.Y(n_1913)
);

AND2x2_ASAP7_75t_L g1914 ( 
.A(n_1528),
.B(n_137),
.Y(n_1914)
);

NAND2xp5_ASAP7_75t_L g1915 ( 
.A(n_1454),
.B(n_138),
.Y(n_1915)
);

NAND2x1p5_ASAP7_75t_L g1916 ( 
.A(n_1500),
.B(n_138),
.Y(n_1916)
);

NAND2xp5_ASAP7_75t_L g1917 ( 
.A(n_1454),
.B(n_139),
.Y(n_1917)
);

AND2x2_ASAP7_75t_L g1918 ( 
.A(n_1538),
.B(n_139),
.Y(n_1918)
);

AND2x2_ASAP7_75t_L g1919 ( 
.A(n_1570),
.B(n_140),
.Y(n_1919)
);

BUFx3_ASAP7_75t_L g1920 ( 
.A(n_1436),
.Y(n_1920)
);

INVx2_ASAP7_75t_L g1921 ( 
.A(n_1630),
.Y(n_1921)
);

INVx1_ASAP7_75t_L g1922 ( 
.A(n_1531),
.Y(n_1922)
);

BUFx6f_ASAP7_75t_L g1923 ( 
.A(n_1550),
.Y(n_1923)
);

INVx2_ASAP7_75t_L g1924 ( 
.A(n_1631),
.Y(n_1924)
);

INVx3_ASAP7_75t_L g1925 ( 
.A(n_1551),
.Y(n_1925)
);

INVx2_ASAP7_75t_L g1926 ( 
.A(n_1540),
.Y(n_1926)
);

AND2x2_ASAP7_75t_L g1927 ( 
.A(n_1518),
.B(n_140),
.Y(n_1927)
);

AND2x2_ASAP7_75t_L g1928 ( 
.A(n_1582),
.B(n_141),
.Y(n_1928)
);

INVx3_ASAP7_75t_L g1929 ( 
.A(n_1571),
.Y(n_1929)
);

INVx1_ASAP7_75t_L g1930 ( 
.A(n_1525),
.Y(n_1930)
);

INVx2_ASAP7_75t_L g1931 ( 
.A(n_1632),
.Y(n_1931)
);

BUFx3_ASAP7_75t_L g1932 ( 
.A(n_1624),
.Y(n_1932)
);

NAND2xp5_ASAP7_75t_L g1933 ( 
.A(n_1458),
.B(n_142),
.Y(n_1933)
);

AND2x2_ASAP7_75t_L g1934 ( 
.A(n_1441),
.B(n_143),
.Y(n_1934)
);

INVxp67_ASAP7_75t_L g1935 ( 
.A(n_1652),
.Y(n_1935)
);

INVx2_ASAP7_75t_L g1936 ( 
.A(n_1560),
.Y(n_1936)
);

BUFx6f_ASAP7_75t_L g1937 ( 
.A(n_1593),
.Y(n_1937)
);

BUFx6f_ASAP7_75t_L g1938 ( 
.A(n_1593),
.Y(n_1938)
);

AND2x2_ASAP7_75t_L g1939 ( 
.A(n_1536),
.B(n_143),
.Y(n_1939)
);

INVx1_ASAP7_75t_L g1940 ( 
.A(n_1458),
.Y(n_1940)
);

INVx2_ASAP7_75t_SL g1941 ( 
.A(n_1636),
.Y(n_1941)
);

AND2x2_ASAP7_75t_L g1942 ( 
.A(n_1586),
.B(n_1573),
.Y(n_1942)
);

INVx1_ASAP7_75t_L g1943 ( 
.A(n_1519),
.Y(n_1943)
);

INVx2_ASAP7_75t_L g1944 ( 
.A(n_1621),
.Y(n_1944)
);

AND2x2_ASAP7_75t_SL g1945 ( 
.A(n_1544),
.B(n_144),
.Y(n_1945)
);

AND2x2_ASAP7_75t_L g1946 ( 
.A(n_1604),
.B(n_145),
.Y(n_1946)
);

HB1xp67_ASAP7_75t_L g1947 ( 
.A(n_1489),
.Y(n_1947)
);

INVxp67_ASAP7_75t_SL g1948 ( 
.A(n_1544),
.Y(n_1948)
);

INVx1_ASAP7_75t_L g1949 ( 
.A(n_1423),
.Y(n_1949)
);

INVx1_ASAP7_75t_L g1950 ( 
.A(n_1423),
.Y(n_1950)
);

AND2x2_ASAP7_75t_L g1951 ( 
.A(n_1607),
.B(n_145),
.Y(n_1951)
);

INVxp67_ASAP7_75t_L g1952 ( 
.A(n_1659),
.Y(n_1952)
);

AND2x2_ASAP7_75t_L g1953 ( 
.A(n_1429),
.B(n_146),
.Y(n_1953)
);

INVx2_ASAP7_75t_L g1954 ( 
.A(n_1623),
.Y(n_1954)
);

INVx1_ASAP7_75t_L g1955 ( 
.A(n_1440),
.Y(n_1955)
);

BUFx3_ASAP7_75t_L g1956 ( 
.A(n_1615),
.Y(n_1956)
);

INVx3_ASAP7_75t_L g1957 ( 
.A(n_1583),
.Y(n_1957)
);

NAND2x1p5_ASAP7_75t_L g1958 ( 
.A(n_1579),
.B(n_146),
.Y(n_1958)
);

NOR2xp33_ASAP7_75t_R g1959 ( 
.A(n_1485),
.B(n_147),
.Y(n_1959)
);

AND2x4_ASAP7_75t_L g1960 ( 
.A(n_1583),
.B(n_148),
.Y(n_1960)
);

INVx1_ASAP7_75t_L g1961 ( 
.A(n_1440),
.Y(n_1961)
);

NAND2xp5_ASAP7_75t_L g1962 ( 
.A(n_1566),
.B(n_1476),
.Y(n_1962)
);

INVx2_ASAP7_75t_L g1963 ( 
.A(n_1547),
.Y(n_1963)
);

BUFx3_ASAP7_75t_L g1964 ( 
.A(n_1541),
.Y(n_1964)
);

AND2x2_ASAP7_75t_L g1965 ( 
.A(n_1405),
.B(n_148),
.Y(n_1965)
);

AND2x2_ASAP7_75t_L g1966 ( 
.A(n_1654),
.B(n_151),
.Y(n_1966)
);

NOR2xp33_ASAP7_75t_L g1967 ( 
.A(n_1443),
.B(n_151),
.Y(n_1967)
);

OAI21xp5_ASAP7_75t_L g1968 ( 
.A1(n_1681),
.A2(n_456),
.B(n_454),
.Y(n_1968)
);

BUFx6f_ASAP7_75t_L g1969 ( 
.A(n_1541),
.Y(n_1969)
);

INVx3_ASAP7_75t_L g1970 ( 
.A(n_1568),
.Y(n_1970)
);

INVx1_ASAP7_75t_L g1971 ( 
.A(n_1585),
.Y(n_1971)
);

INVx1_ASAP7_75t_L g1972 ( 
.A(n_1585),
.Y(n_1972)
);

INVx1_ASAP7_75t_L g1973 ( 
.A(n_1627),
.Y(n_1973)
);

INVx4_ASAP7_75t_L g1974 ( 
.A(n_1548),
.Y(n_1974)
);

NAND2xp5_ASAP7_75t_L g1975 ( 
.A(n_1476),
.B(n_152),
.Y(n_1975)
);

NAND2xp5_ASAP7_75t_L g1976 ( 
.A(n_1508),
.B(n_153),
.Y(n_1976)
);

AND2x4_ASAP7_75t_L g1977 ( 
.A(n_1452),
.B(n_153),
.Y(n_1977)
);

CKINVDCx5p33_ASAP7_75t_R g1978 ( 
.A(n_1520),
.Y(n_1978)
);

AND2x2_ASAP7_75t_L g1979 ( 
.A(n_1475),
.B(n_154),
.Y(n_1979)
);

INVx1_ASAP7_75t_L g1980 ( 
.A(n_1640),
.Y(n_1980)
);

NAND2xp5_ASAP7_75t_L g1981 ( 
.A(n_1508),
.B(n_154),
.Y(n_1981)
);

AND2x2_ASAP7_75t_L g1982 ( 
.A(n_1516),
.B(n_156),
.Y(n_1982)
);

HB1xp67_ASAP7_75t_L g1983 ( 
.A(n_1552),
.Y(n_1983)
);

BUFx2_ASAP7_75t_L g1984 ( 
.A(n_1664),
.Y(n_1984)
);

AND2x2_ASAP7_75t_L g1985 ( 
.A(n_1490),
.B(n_156),
.Y(n_1985)
);

INVx2_ASAP7_75t_SL g1986 ( 
.A(n_1473),
.Y(n_1986)
);

AND2x2_ASAP7_75t_L g1987 ( 
.A(n_1511),
.B(n_157),
.Y(n_1987)
);

AND2x2_ASAP7_75t_SL g1988 ( 
.A(n_1618),
.B(n_159),
.Y(n_1988)
);

INVx1_ASAP7_75t_L g1989 ( 
.A(n_1644),
.Y(n_1989)
);

BUFx3_ASAP7_75t_L g1990 ( 
.A(n_1599),
.Y(n_1990)
);

AND2x2_ASAP7_75t_L g1991 ( 
.A(n_1511),
.B(n_160),
.Y(n_1991)
);

AND2x2_ASAP7_75t_L g1992 ( 
.A(n_1677),
.B(n_160),
.Y(n_1992)
);

NAND2xp5_ASAP7_75t_L g1993 ( 
.A(n_1543),
.B(n_1473),
.Y(n_1993)
);

AND2x2_ASAP7_75t_SL g1994 ( 
.A(n_1459),
.B(n_161),
.Y(n_1994)
);

NOR2xp33_ASAP7_75t_L g1995 ( 
.A(n_1545),
.B(n_162),
.Y(n_1995)
);

BUFx6f_ASAP7_75t_L g1996 ( 
.A(n_1651),
.Y(n_1996)
);

INVx4_ASAP7_75t_L g1997 ( 
.A(n_1635),
.Y(n_1997)
);

NAND2xp5_ASAP7_75t_L g1998 ( 
.A(n_1410),
.B(n_164),
.Y(n_1998)
);

AND2x2_ASAP7_75t_L g1999 ( 
.A(n_1598),
.B(n_165),
.Y(n_1999)
);

INVx2_ASAP7_75t_SL g2000 ( 
.A(n_1660),
.Y(n_2000)
);

INVx2_ASAP7_75t_L g2001 ( 
.A(n_1622),
.Y(n_2001)
);

BUFx3_ASAP7_75t_L g2002 ( 
.A(n_1589),
.Y(n_2002)
);

NOR2xp67_ASAP7_75t_SL g2003 ( 
.A(n_1616),
.B(n_166),
.Y(n_2003)
);

AND2x2_ASAP7_75t_L g2004 ( 
.A(n_1667),
.B(n_167),
.Y(n_2004)
);

INVx2_ASAP7_75t_L g2005 ( 
.A(n_1622),
.Y(n_2005)
);

BUFx5_ASAP7_75t_L g2006 ( 
.A(n_1595),
.Y(n_2006)
);

BUFx5_ASAP7_75t_L g2007 ( 
.A(n_1617),
.Y(n_2007)
);

INVx2_ASAP7_75t_L g2008 ( 
.A(n_1673),
.Y(n_2008)
);

INVx2_ASAP7_75t_L g2009 ( 
.A(n_1629),
.Y(n_2009)
);

AND2x4_ASAP7_75t_L g2010 ( 
.A(n_1587),
.B(n_168),
.Y(n_2010)
);

OAI21x1_ASAP7_75t_L g2011 ( 
.A1(n_1616),
.A2(n_461),
.B(n_459),
.Y(n_2011)
);

AND2x2_ASAP7_75t_L g2012 ( 
.A(n_1606),
.B(n_169),
.Y(n_2012)
);

INVx2_ASAP7_75t_L g2013 ( 
.A(n_1629),
.Y(n_2013)
);

AND2x2_ASAP7_75t_L g2014 ( 
.A(n_1602),
.B(n_169),
.Y(n_2014)
);

NAND2xp5_ASAP7_75t_L g2015 ( 
.A(n_1403),
.B(n_170),
.Y(n_2015)
);

INVx1_ASAP7_75t_SL g2016 ( 
.A(n_1424),
.Y(n_2016)
);

BUFx3_ASAP7_75t_L g2017 ( 
.A(n_1633),
.Y(n_2017)
);

INVx1_ASAP7_75t_L g2018 ( 
.A(n_1521),
.Y(n_2018)
);

HB1xp67_ASAP7_75t_L g2019 ( 
.A(n_1687),
.Y(n_2019)
);

NAND2xp5_ASAP7_75t_L g2020 ( 
.A(n_1474),
.B(n_171),
.Y(n_2020)
);

BUFx3_ASAP7_75t_L g2021 ( 
.A(n_1467),
.Y(n_2021)
);

NAND2xp5_ASAP7_75t_L g2022 ( 
.A(n_1453),
.B(n_171),
.Y(n_2022)
);

NOR2xp33_ASAP7_75t_SL g2023 ( 
.A(n_1666),
.B(n_172),
.Y(n_2023)
);

BUFx3_ASAP7_75t_L g2024 ( 
.A(n_1574),
.Y(n_2024)
);

AND2x2_ASAP7_75t_L g2025 ( 
.A(n_1666),
.B(n_172),
.Y(n_2025)
);

INVx1_ASAP7_75t_L g2026 ( 
.A(n_1401),
.Y(n_2026)
);

AND2x2_ASAP7_75t_L g2027 ( 
.A(n_1666),
.B(n_173),
.Y(n_2027)
);

INVx2_ASAP7_75t_L g2028 ( 
.A(n_1576),
.Y(n_2028)
);

AND2x2_ASAP7_75t_L g2029 ( 
.A(n_1666),
.B(n_173),
.Y(n_2029)
);

OAI21xp5_ASAP7_75t_L g2030 ( 
.A1(n_1478),
.A2(n_464),
.B(n_462),
.Y(n_2030)
);

NOR2xp33_ASAP7_75t_L g2031 ( 
.A(n_1414),
.B(n_175),
.Y(n_2031)
);

BUFx2_ASAP7_75t_L g2032 ( 
.A(n_1739),
.Y(n_2032)
);

AND2x4_ASAP7_75t_L g2033 ( 
.A(n_1964),
.B(n_1940),
.Y(n_2033)
);

NAND2xp5_ASAP7_75t_SL g2034 ( 
.A(n_1945),
.B(n_176),
.Y(n_2034)
);

BUFx2_ASAP7_75t_L g2035 ( 
.A(n_1739),
.Y(n_2035)
);

NOR2xp33_ASAP7_75t_L g2036 ( 
.A(n_1877),
.B(n_177),
.Y(n_2036)
);

BUFx6f_ASAP7_75t_L g2037 ( 
.A(n_1736),
.Y(n_2037)
);

OR2x6_ASAP7_75t_L g2038 ( 
.A(n_1739),
.B(n_178),
.Y(n_2038)
);

OR2x6_ASAP7_75t_L g2039 ( 
.A(n_1803),
.B(n_178),
.Y(n_2039)
);

INVx2_ASAP7_75t_L g2040 ( 
.A(n_1746),
.Y(n_2040)
);

AND2x2_ASAP7_75t_L g2041 ( 
.A(n_1877),
.B(n_179),
.Y(n_2041)
);

INVx1_ASAP7_75t_L g2042 ( 
.A(n_1963),
.Y(n_2042)
);

OR2x2_ASAP7_75t_L g2043 ( 
.A(n_1827),
.B(n_179),
.Y(n_2043)
);

BUFx2_ASAP7_75t_L g2044 ( 
.A(n_1768),
.Y(n_2044)
);

OR2x2_ASAP7_75t_L g2045 ( 
.A(n_1791),
.B(n_180),
.Y(n_2045)
);

BUFx3_ASAP7_75t_L g2046 ( 
.A(n_1803),
.Y(n_2046)
);

INVx2_ASAP7_75t_L g2047 ( 
.A(n_1746),
.Y(n_2047)
);

NAND2xp5_ASAP7_75t_L g2048 ( 
.A(n_1926),
.B(n_180),
.Y(n_2048)
);

INVx1_ASAP7_75t_L g2049 ( 
.A(n_1963),
.Y(n_2049)
);

INVx2_ASAP7_75t_L g2050 ( 
.A(n_1974),
.Y(n_2050)
);

AOI21x1_ASAP7_75t_L g2051 ( 
.A1(n_2003),
.A2(n_468),
.B(n_466),
.Y(n_2051)
);

BUFx2_ASAP7_75t_L g2052 ( 
.A(n_1768),
.Y(n_2052)
);

BUFx2_ASAP7_75t_L g2053 ( 
.A(n_1717),
.Y(n_2053)
);

INVx4_ASAP7_75t_L g2054 ( 
.A(n_1736),
.Y(n_2054)
);

INVx1_ASAP7_75t_SL g2055 ( 
.A(n_1708),
.Y(n_2055)
);

NAND2x1_ASAP7_75t_L g2056 ( 
.A(n_1777),
.B(n_469),
.Y(n_2056)
);

AND2x2_ASAP7_75t_L g2057 ( 
.A(n_2010),
.B(n_182),
.Y(n_2057)
);

AND2x4_ASAP7_75t_L g2058 ( 
.A(n_1964),
.B(n_182),
.Y(n_2058)
);

NOR2xp33_ASAP7_75t_L g2059 ( 
.A(n_1828),
.B(n_183),
.Y(n_2059)
);

NAND2xp5_ASAP7_75t_L g2060 ( 
.A(n_1926),
.B(n_183),
.Y(n_2060)
);

AND2x4_ASAP7_75t_L g2061 ( 
.A(n_1949),
.B(n_184),
.Y(n_2061)
);

INVx6_ASAP7_75t_L g2062 ( 
.A(n_1845),
.Y(n_2062)
);

INVxp67_ASAP7_75t_SL g2063 ( 
.A(n_1708),
.Y(n_2063)
);

NAND2x1p5_ASAP7_75t_L g2064 ( 
.A(n_2024),
.B(n_185),
.Y(n_2064)
);

NAND2xp5_ASAP7_75t_L g2065 ( 
.A(n_1970),
.B(n_186),
.Y(n_2065)
);

BUFx6f_ASAP7_75t_L g2066 ( 
.A(n_1736),
.Y(n_2066)
);

INVx1_ASAP7_75t_L g2067 ( 
.A(n_1922),
.Y(n_2067)
);

AND2x2_ASAP7_75t_SL g2068 ( 
.A(n_1719),
.B(n_1945),
.Y(n_2068)
);

INVxp67_ASAP7_75t_L g2069 ( 
.A(n_1960),
.Y(n_2069)
);

INVx3_ASAP7_75t_L g2070 ( 
.A(n_1777),
.Y(n_2070)
);

INVx2_ASAP7_75t_L g2071 ( 
.A(n_1974),
.Y(n_2071)
);

INVx3_ASAP7_75t_L g2072 ( 
.A(n_1777),
.Y(n_2072)
);

AND2x2_ASAP7_75t_L g2073 ( 
.A(n_2010),
.B(n_186),
.Y(n_2073)
);

BUFx2_ASAP7_75t_L g2074 ( 
.A(n_1717),
.Y(n_2074)
);

INVx2_ASAP7_75t_L g2075 ( 
.A(n_1974),
.Y(n_2075)
);

NAND2xp5_ASAP7_75t_L g2076 ( 
.A(n_1970),
.B(n_187),
.Y(n_2076)
);

INVx1_ASAP7_75t_L g2077 ( 
.A(n_1714),
.Y(n_2077)
);

OR2x6_ASAP7_75t_L g2078 ( 
.A(n_1710),
.B(n_188),
.Y(n_2078)
);

CKINVDCx5p33_ASAP7_75t_R g2079 ( 
.A(n_1810),
.Y(n_2079)
);

NAND2xp5_ASAP7_75t_L g2080 ( 
.A(n_1970),
.B(n_189),
.Y(n_2080)
);

AND2x2_ASAP7_75t_L g2081 ( 
.A(n_2010),
.B(n_189),
.Y(n_2081)
);

BUFx3_ASAP7_75t_L g2082 ( 
.A(n_1845),
.Y(n_2082)
);

AND2x2_ASAP7_75t_L g2083 ( 
.A(n_1852),
.B(n_190),
.Y(n_2083)
);

NAND2x1p5_ASAP7_75t_L g2084 ( 
.A(n_2024),
.B(n_191),
.Y(n_2084)
);

NOR2xp33_ASAP7_75t_SL g2085 ( 
.A(n_1710),
.B(n_470),
.Y(n_2085)
);

BUFx2_ASAP7_75t_L g2086 ( 
.A(n_1727),
.Y(n_2086)
);

INVx3_ASAP7_75t_L g2087 ( 
.A(n_1785),
.Y(n_2087)
);

AND2x2_ASAP7_75t_SL g2088 ( 
.A(n_1719),
.B(n_191),
.Y(n_2088)
);

AND2x2_ASAP7_75t_L g2089 ( 
.A(n_1999),
.B(n_192),
.Y(n_2089)
);

BUFx4f_ASAP7_75t_L g2090 ( 
.A(n_1695),
.Y(n_2090)
);

AND2x4_ASAP7_75t_L g2091 ( 
.A(n_1950),
.B(n_192),
.Y(n_2091)
);

AND2x6_ASAP7_75t_L g2092 ( 
.A(n_1790),
.B(n_193),
.Y(n_2092)
);

NOR2xp33_ASAP7_75t_SL g2093 ( 
.A(n_1710),
.B(n_474),
.Y(n_2093)
);

NAND2xp5_ASAP7_75t_L g2094 ( 
.A(n_1861),
.B(n_193),
.Y(n_2094)
);

NAND2xp5_ASAP7_75t_L g2095 ( 
.A(n_1861),
.B(n_194),
.Y(n_2095)
);

INVxp67_ASAP7_75t_SL g2096 ( 
.A(n_1727),
.Y(n_2096)
);

BUFx3_ASAP7_75t_L g2097 ( 
.A(n_1845),
.Y(n_2097)
);

INVxp67_ASAP7_75t_L g2098 ( 
.A(n_1960),
.Y(n_2098)
);

OR2x6_ASAP7_75t_L g2099 ( 
.A(n_1725),
.B(n_194),
.Y(n_2099)
);

INVx2_ASAP7_75t_L g2100 ( 
.A(n_1797),
.Y(n_2100)
);

NOR2xp33_ASAP7_75t_SL g2101 ( 
.A(n_1725),
.B(n_475),
.Y(n_2101)
);

AND2x6_ASAP7_75t_L g2102 ( 
.A(n_1790),
.B(n_195),
.Y(n_2102)
);

NAND2xp5_ASAP7_75t_L g2103 ( 
.A(n_1955),
.B(n_1961),
.Y(n_2103)
);

INVx2_ASAP7_75t_L g2104 ( 
.A(n_1797),
.Y(n_2104)
);

NAND2xp5_ASAP7_75t_L g2105 ( 
.A(n_1721),
.B(n_195),
.Y(n_2105)
);

OR2x2_ASAP7_75t_L g2106 ( 
.A(n_2002),
.B(n_196),
.Y(n_2106)
);

HB1xp67_ASAP7_75t_L g2107 ( 
.A(n_1731),
.Y(n_2107)
);

AND2x2_ASAP7_75t_L g2108 ( 
.A(n_2014),
.B(n_197),
.Y(n_2108)
);

INVx1_ASAP7_75t_L g2109 ( 
.A(n_1769),
.Y(n_2109)
);

INVx2_ASAP7_75t_SL g2110 ( 
.A(n_1859),
.Y(n_2110)
);

INVxp67_ASAP7_75t_L g2111 ( 
.A(n_1960),
.Y(n_2111)
);

BUFx12f_ASAP7_75t_L g2112 ( 
.A(n_1908),
.Y(n_2112)
);

BUFx2_ASAP7_75t_L g2113 ( 
.A(n_1731),
.Y(n_2113)
);

INVx1_ASAP7_75t_L g2114 ( 
.A(n_1774),
.Y(n_2114)
);

NAND2xp5_ASAP7_75t_L g2115 ( 
.A(n_1883),
.B(n_197),
.Y(n_2115)
);

OR2x6_ASAP7_75t_L g2116 ( 
.A(n_1725),
.B(n_198),
.Y(n_2116)
);

OR2x6_ASAP7_75t_L g2117 ( 
.A(n_1790),
.B(n_198),
.Y(n_2117)
);

NAND2xp5_ASAP7_75t_L g2118 ( 
.A(n_1883),
.B(n_199),
.Y(n_2118)
);

INVx2_ASAP7_75t_L g2119 ( 
.A(n_1798),
.Y(n_2119)
);

AND2x2_ASAP7_75t_L g2120 ( 
.A(n_1795),
.B(n_201),
.Y(n_2120)
);

NAND2xp5_ASAP7_75t_L g2121 ( 
.A(n_1993),
.B(n_203),
.Y(n_2121)
);

INVx1_ASAP7_75t_L g2122 ( 
.A(n_1780),
.Y(n_2122)
);

OR2x6_ASAP7_75t_SL g2123 ( 
.A(n_1978),
.B(n_205),
.Y(n_2123)
);

INVx2_ASAP7_75t_SL g2124 ( 
.A(n_1859),
.Y(n_2124)
);

OR2x2_ASAP7_75t_L g2125 ( 
.A(n_2002),
.B(n_205),
.Y(n_2125)
);

INVx2_ASAP7_75t_L g2126 ( 
.A(n_1798),
.Y(n_2126)
);

BUFx4_ASAP7_75t_SL g2127 ( 
.A(n_1956),
.Y(n_2127)
);

BUFx2_ASAP7_75t_L g2128 ( 
.A(n_1695),
.Y(n_2128)
);

INVxp67_ASAP7_75t_L g2129 ( 
.A(n_2023),
.Y(n_2129)
);

CKINVDCx11_ASAP7_75t_R g2130 ( 
.A(n_1932),
.Y(n_2130)
);

INVx1_ASAP7_75t_L g2131 ( 
.A(n_1794),
.Y(n_2131)
);

HB1xp67_ASAP7_75t_L g2132 ( 
.A(n_1758),
.Y(n_2132)
);

NAND2xp5_ASAP7_75t_L g2133 ( 
.A(n_1971),
.B(n_206),
.Y(n_2133)
);

BUFx12f_ASAP7_75t_L g2134 ( 
.A(n_1916),
.Y(n_2134)
);

NAND2xp5_ASAP7_75t_L g2135 ( 
.A(n_1972),
.B(n_207),
.Y(n_2135)
);

INVx4_ASAP7_75t_L g2136 ( 
.A(n_1736),
.Y(n_2136)
);

INVx2_ASAP7_75t_L g2137 ( 
.A(n_1819),
.Y(n_2137)
);

NAND2xp5_ASAP7_75t_L g2138 ( 
.A(n_1962),
.B(n_207),
.Y(n_2138)
);

NOR2xp33_ASAP7_75t_L g2139 ( 
.A(n_1828),
.B(n_208),
.Y(n_2139)
);

BUFx6f_ASAP7_75t_L g2140 ( 
.A(n_1748),
.Y(n_2140)
);

INVx1_ASAP7_75t_L g2141 ( 
.A(n_1802),
.Y(n_2141)
);

NOR2xp33_ASAP7_75t_SL g2142 ( 
.A(n_1707),
.B(n_476),
.Y(n_2142)
);

NOR2xp33_ASAP7_75t_SL g2143 ( 
.A(n_1707),
.B(n_477),
.Y(n_2143)
);

AO21x2_ASAP7_75t_L g2144 ( 
.A1(n_1900),
.A2(n_482),
.B(n_479),
.Y(n_2144)
);

BUFx3_ASAP7_75t_L g2145 ( 
.A(n_1748),
.Y(n_2145)
);

BUFx3_ASAP7_75t_L g2146 ( 
.A(n_1748),
.Y(n_2146)
);

BUFx6f_ASAP7_75t_L g2147 ( 
.A(n_1748),
.Y(n_2147)
);

NAND2xp5_ASAP7_75t_L g2148 ( 
.A(n_1701),
.B(n_1909),
.Y(n_2148)
);

AND2x4_ASAP7_75t_L g2149 ( 
.A(n_1957),
.B(n_210),
.Y(n_2149)
);

INVx1_ASAP7_75t_L g2150 ( 
.A(n_1807),
.Y(n_2150)
);

OR2x2_ASAP7_75t_L g2151 ( 
.A(n_1984),
.B(n_210),
.Y(n_2151)
);

BUFx3_ASAP7_75t_L g2152 ( 
.A(n_1758),
.Y(n_2152)
);

INVx4_ASAP7_75t_L g2153 ( 
.A(n_1695),
.Y(n_2153)
);

INVx3_ASAP7_75t_L g2154 ( 
.A(n_1785),
.Y(n_2154)
);

NAND2xp5_ASAP7_75t_SL g2155 ( 
.A(n_1713),
.B(n_211),
.Y(n_2155)
);

BUFx6f_ASAP7_75t_L g2156 ( 
.A(n_1903),
.Y(n_2156)
);

INVxp67_ASAP7_75t_L g2157 ( 
.A(n_1701),
.Y(n_2157)
);

INVx5_ASAP7_75t_L g2158 ( 
.A(n_1695),
.Y(n_2158)
);

INVx3_ASAP7_75t_L g2159 ( 
.A(n_1785),
.Y(n_2159)
);

AND2x4_ASAP7_75t_L g2160 ( 
.A(n_1957),
.B(n_211),
.Y(n_2160)
);

INVx6_ASAP7_75t_L g2161 ( 
.A(n_1738),
.Y(n_2161)
);

INVx2_ASAP7_75t_SL g2162 ( 
.A(n_1788),
.Y(n_2162)
);

NAND2xp5_ASAP7_75t_L g2163 ( 
.A(n_1702),
.B(n_1700),
.Y(n_2163)
);

OR2x2_ASAP7_75t_L g2164 ( 
.A(n_1880),
.B(n_212),
.Y(n_2164)
);

INVx4_ASAP7_75t_L g2165 ( 
.A(n_1695),
.Y(n_2165)
);

BUFx4f_ASAP7_75t_L g2166 ( 
.A(n_1715),
.Y(n_2166)
);

BUFx2_ASAP7_75t_L g2167 ( 
.A(n_1713),
.Y(n_2167)
);

INVx2_ASAP7_75t_L g2168 ( 
.A(n_1819),
.Y(n_2168)
);

OR2x2_ASAP7_75t_L g2169 ( 
.A(n_1935),
.B(n_1952),
.Y(n_2169)
);

NAND2x1p5_ASAP7_75t_L g2170 ( 
.A(n_1738),
.B(n_213),
.Y(n_2170)
);

INVx1_ASAP7_75t_L g2171 ( 
.A(n_1812),
.Y(n_2171)
);

OR2x2_ASAP7_75t_L g2172 ( 
.A(n_1712),
.B(n_214),
.Y(n_2172)
);

INVx2_ASAP7_75t_SL g2173 ( 
.A(n_1788),
.Y(n_2173)
);

AND2x4_ASAP7_75t_L g2174 ( 
.A(n_1957),
.B(n_214),
.Y(n_2174)
);

NAND2xp5_ASAP7_75t_L g2175 ( 
.A(n_1702),
.B(n_1734),
.Y(n_2175)
);

INVxp67_ASAP7_75t_L g2176 ( 
.A(n_1711),
.Y(n_2176)
);

OR2x6_ASAP7_75t_L g2177 ( 
.A(n_1815),
.B(n_215),
.Y(n_2177)
);

AND2x2_ASAP7_75t_L g2178 ( 
.A(n_1965),
.B(n_216),
.Y(n_2178)
);

AND2x4_ASAP7_75t_L g2179 ( 
.A(n_1894),
.B(n_216),
.Y(n_2179)
);

AND2x2_ASAP7_75t_L g2180 ( 
.A(n_1966),
.B(n_217),
.Y(n_2180)
);

BUFx6f_ASAP7_75t_L g2181 ( 
.A(n_1903),
.Y(n_2181)
);

CKINVDCx5p33_ASAP7_75t_R g2182 ( 
.A(n_1833),
.Y(n_2182)
);

INVx2_ASAP7_75t_L g2183 ( 
.A(n_1826),
.Y(n_2183)
);

INVx2_ASAP7_75t_L g2184 ( 
.A(n_1826),
.Y(n_2184)
);

INVx3_ASAP7_75t_L g2185 ( 
.A(n_1691),
.Y(n_2185)
);

INVx1_ASAP7_75t_L g2186 ( 
.A(n_1814),
.Y(n_2186)
);

NAND2xp5_ASAP7_75t_L g2187 ( 
.A(n_1894),
.B(n_218),
.Y(n_2187)
);

NAND2xp5_ASAP7_75t_L g2188 ( 
.A(n_1894),
.B(n_218),
.Y(n_2188)
);

INVx1_ASAP7_75t_SL g2189 ( 
.A(n_2001),
.Y(n_2189)
);

NOR2xp33_ASAP7_75t_SL g2190 ( 
.A(n_1896),
.B(n_483),
.Y(n_2190)
);

INVx3_ASAP7_75t_L g2191 ( 
.A(n_1691),
.Y(n_2191)
);

CKINVDCx10_ASAP7_75t_R g2192 ( 
.A(n_1833),
.Y(n_2192)
);

INVx2_ASAP7_75t_L g2193 ( 
.A(n_1834),
.Y(n_2193)
);

INVx1_ASAP7_75t_L g2194 ( 
.A(n_1825),
.Y(n_2194)
);

AND2x2_ASAP7_75t_L g2195 ( 
.A(n_1953),
.B(n_219),
.Y(n_2195)
);

INVx2_ASAP7_75t_L g2196 ( 
.A(n_1834),
.Y(n_2196)
);

OR2x6_ASAP7_75t_L g2197 ( 
.A(n_1815),
.B(n_219),
.Y(n_2197)
);

NAND2xp5_ASAP7_75t_L g2198 ( 
.A(n_1752),
.B(n_220),
.Y(n_2198)
);

AND2x2_ASAP7_75t_L g2199 ( 
.A(n_1934),
.B(n_220),
.Y(n_2199)
);

NAND2x1p5_ASAP7_75t_L g2200 ( 
.A(n_1738),
.B(n_223),
.Y(n_2200)
);

AND2x2_ASAP7_75t_L g2201 ( 
.A(n_1749),
.B(n_224),
.Y(n_2201)
);

AND2x4_ASAP7_75t_L g2202 ( 
.A(n_1986),
.B(n_1735),
.Y(n_2202)
);

NAND2xp5_ASAP7_75t_L g2203 ( 
.A(n_1759),
.B(n_224),
.Y(n_2203)
);

INVx1_ASAP7_75t_L g2204 ( 
.A(n_1843),
.Y(n_2204)
);

NAND2x1p5_ASAP7_75t_L g2205 ( 
.A(n_1709),
.B(n_225),
.Y(n_2205)
);

OR2x2_ASAP7_75t_L g2206 ( 
.A(n_1897),
.B(n_227),
.Y(n_2206)
);

INVxp67_ASAP7_75t_SL g2207 ( 
.A(n_2001),
.Y(n_2207)
);

NAND2xp5_ASAP7_75t_L g2208 ( 
.A(n_1857),
.B(n_227),
.Y(n_2208)
);

INVx1_ASAP7_75t_L g2209 ( 
.A(n_1846),
.Y(n_2209)
);

INVx1_ASAP7_75t_L g2210 ( 
.A(n_1854),
.Y(n_2210)
);

BUFx2_ASAP7_75t_L g2211 ( 
.A(n_1750),
.Y(n_2211)
);

HB1xp67_ASAP7_75t_L g2212 ( 
.A(n_1750),
.Y(n_2212)
);

NAND2xp5_ASAP7_75t_L g2213 ( 
.A(n_1867),
.B(n_228),
.Y(n_2213)
);

AND2x4_ASAP7_75t_L g2214 ( 
.A(n_1986),
.B(n_228),
.Y(n_2214)
);

INVx2_ASAP7_75t_L g2215 ( 
.A(n_1699),
.Y(n_2215)
);

INVx2_ASAP7_75t_L g2216 ( 
.A(n_1699),
.Y(n_2216)
);

INVx4_ASAP7_75t_L g2217 ( 
.A(n_1691),
.Y(n_2217)
);

BUFx4f_ASAP7_75t_L g2218 ( 
.A(n_1715),
.Y(n_2218)
);

NAND2xp5_ASAP7_75t_L g2219 ( 
.A(n_1875),
.B(n_229),
.Y(n_2219)
);

INVx2_ASAP7_75t_L g2220 ( 
.A(n_1703),
.Y(n_2220)
);

NOR2xp67_ASAP7_75t_L g2221 ( 
.A(n_1896),
.B(n_485),
.Y(n_2221)
);

OR2x2_ASAP7_75t_L g2222 ( 
.A(n_1942),
.B(n_229),
.Y(n_2222)
);

OR2x6_ASAP7_75t_L g2223 ( 
.A(n_1815),
.B(n_1817),
.Y(n_2223)
);

CKINVDCx6p67_ASAP7_75t_R g2224 ( 
.A(n_1932),
.Y(n_2224)
);

INVx1_ASAP7_75t_L g2225 ( 
.A(n_1778),
.Y(n_2225)
);

AND2x2_ASAP7_75t_L g2226 ( 
.A(n_1864),
.B(n_231),
.Y(n_2226)
);

NOR2xp33_ASAP7_75t_SL g2227 ( 
.A(n_1896),
.B(n_486),
.Y(n_2227)
);

INVx1_ASAP7_75t_L g2228 ( 
.A(n_1787),
.Y(n_2228)
);

INVxp67_ASAP7_75t_L g2229 ( 
.A(n_1733),
.Y(n_2229)
);

OR2x2_ASAP7_75t_L g2230 ( 
.A(n_1772),
.B(n_233),
.Y(n_2230)
);

NAND2xp5_ASAP7_75t_L g2231 ( 
.A(n_1936),
.B(n_233),
.Y(n_2231)
);

INVx1_ASAP7_75t_L g2232 ( 
.A(n_1787),
.Y(n_2232)
);

AND2x4_ASAP7_75t_L g2233 ( 
.A(n_1735),
.B(n_234),
.Y(n_2233)
);

NAND2xp5_ASAP7_75t_L g2234 ( 
.A(n_1936),
.B(n_236),
.Y(n_2234)
);

NOR2xp33_ASAP7_75t_SL g2235 ( 
.A(n_1755),
.B(n_487),
.Y(n_2235)
);

BUFx2_ASAP7_75t_L g2236 ( 
.A(n_1959),
.Y(n_2236)
);

BUFx12f_ASAP7_75t_L g2237 ( 
.A(n_1916),
.Y(n_2237)
);

INVx1_ASAP7_75t_L g2238 ( 
.A(n_1744),
.Y(n_2238)
);

BUFx2_ASAP7_75t_L g2239 ( 
.A(n_1959),
.Y(n_2239)
);

AND2x4_ASAP7_75t_L g2240 ( 
.A(n_1766),
.B(n_236),
.Y(n_2240)
);

NAND2xp5_ASAP7_75t_L g2241 ( 
.A(n_1816),
.B(n_238),
.Y(n_2241)
);

AND2x4_ASAP7_75t_L g2242 ( 
.A(n_1766),
.B(n_238),
.Y(n_2242)
);

INVx1_ASAP7_75t_L g2243 ( 
.A(n_1832),
.Y(n_2243)
);

INVx1_ASAP7_75t_L g2244 ( 
.A(n_1874),
.Y(n_2244)
);

INVx1_ASAP7_75t_L g2245 ( 
.A(n_1874),
.Y(n_2245)
);

NAND2xp5_ASAP7_75t_L g2246 ( 
.A(n_1848),
.B(n_239),
.Y(n_2246)
);

INVx3_ASAP7_75t_L g2247 ( 
.A(n_1709),
.Y(n_2247)
);

BUFx12f_ASAP7_75t_L g2248 ( 
.A(n_1978),
.Y(n_2248)
);

INVx1_ASAP7_75t_L g2249 ( 
.A(n_1879),
.Y(n_2249)
);

INVx2_ASAP7_75t_L g2250 ( 
.A(n_1703),
.Y(n_2250)
);

INVx1_ASAP7_75t_L g2251 ( 
.A(n_1879),
.Y(n_2251)
);

BUFx6f_ASAP7_75t_L g2252 ( 
.A(n_1903),
.Y(n_2252)
);

INVx4_ASAP7_75t_L g2253 ( 
.A(n_1732),
.Y(n_2253)
);

AND2x2_ASAP7_75t_L g2254 ( 
.A(n_1741),
.B(n_239),
.Y(n_2254)
);

INVx3_ASAP7_75t_L g2255 ( 
.A(n_1732),
.Y(n_2255)
);

INVx1_ASAP7_75t_L g2256 ( 
.A(n_1885),
.Y(n_2256)
);

INVx3_ASAP7_75t_L g2257 ( 
.A(n_1742),
.Y(n_2257)
);

INVx1_ASAP7_75t_L g2258 ( 
.A(n_1885),
.Y(n_2258)
);

INVx1_ASAP7_75t_SL g2259 ( 
.A(n_2005),
.Y(n_2259)
);

BUFx6f_ASAP7_75t_L g2260 ( 
.A(n_1903),
.Y(n_2260)
);

INVxp67_ASAP7_75t_L g2261 ( 
.A(n_1733),
.Y(n_2261)
);

AND2x2_ASAP7_75t_L g2262 ( 
.A(n_1745),
.B(n_240),
.Y(n_2262)
);

NAND2xp5_ASAP7_75t_L g2263 ( 
.A(n_1824),
.B(n_241),
.Y(n_2263)
);

INVx1_ASAP7_75t_L g2264 ( 
.A(n_1890),
.Y(n_2264)
);

BUFx6f_ASAP7_75t_L g2265 ( 
.A(n_1920),
.Y(n_2265)
);

INVx5_ASAP7_75t_L g2266 ( 
.A(n_1698),
.Y(n_2266)
);

AND2x2_ASAP7_75t_L g2267 ( 
.A(n_1939),
.B(n_241),
.Y(n_2267)
);

INVx1_ASAP7_75t_L g2268 ( 
.A(n_1890),
.Y(n_2268)
);

AND2x4_ASAP7_75t_L g2269 ( 
.A(n_1786),
.B(n_242),
.Y(n_2269)
);

CKINVDCx11_ASAP7_75t_R g2270 ( 
.A(n_2021),
.Y(n_2270)
);

AND2x2_ASAP7_75t_L g2271 ( 
.A(n_1813),
.B(n_242),
.Y(n_2271)
);

BUFx2_ASAP7_75t_L g2272 ( 
.A(n_1817),
.Y(n_2272)
);

AND2x4_ASAP7_75t_L g2273 ( 
.A(n_1786),
.B(n_243),
.Y(n_2273)
);

AND2x4_ASAP7_75t_L g2274 ( 
.A(n_1789),
.B(n_243),
.Y(n_2274)
);

INVx2_ASAP7_75t_L g2275 ( 
.A(n_1737),
.Y(n_2275)
);

BUFx2_ASAP7_75t_L g2276 ( 
.A(n_1817),
.Y(n_2276)
);

NAND2x1_ASAP7_75t_SL g2277 ( 
.A(n_1983),
.B(n_244),
.Y(n_2277)
);

INVx1_ASAP7_75t_L g2278 ( 
.A(n_1892),
.Y(n_2278)
);

BUFx4_ASAP7_75t_SL g2279 ( 
.A(n_1956),
.Y(n_2279)
);

INVx1_ASAP7_75t_L g2280 ( 
.A(n_1892),
.Y(n_2280)
);

AND2x4_ASAP7_75t_L g2281 ( 
.A(n_1789),
.B(n_245),
.Y(n_2281)
);

OR2x6_ASAP7_75t_L g2282 ( 
.A(n_1836),
.B(n_246),
.Y(n_2282)
);

NOR2xp67_ASAP7_75t_L g2283 ( 
.A(n_1716),
.B(n_488),
.Y(n_2283)
);

BUFx12f_ASAP7_75t_L g2284 ( 
.A(n_1977),
.Y(n_2284)
);

CKINVDCx5p33_ASAP7_75t_R g2285 ( 
.A(n_1743),
.Y(n_2285)
);

INVx3_ASAP7_75t_L g2286 ( 
.A(n_1742),
.Y(n_2286)
);

AND2x4_ASAP7_75t_L g2287 ( 
.A(n_1973),
.B(n_246),
.Y(n_2287)
);

CKINVDCx5p33_ASAP7_75t_R g2288 ( 
.A(n_1779),
.Y(n_2288)
);

NAND2xp5_ASAP7_75t_L g2289 ( 
.A(n_1824),
.B(n_248),
.Y(n_2289)
);

INVx1_ASAP7_75t_L g2290 ( 
.A(n_1898),
.Y(n_2290)
);

BUFx6f_ASAP7_75t_L g2291 ( 
.A(n_1920),
.Y(n_2291)
);

OR2x6_ASAP7_75t_L g2292 ( 
.A(n_1836),
.B(n_249),
.Y(n_2292)
);

AND2x4_ASAP7_75t_L g2293 ( 
.A(n_1693),
.B(n_250),
.Y(n_2293)
);

INVx3_ASAP7_75t_L g2294 ( 
.A(n_2005),
.Y(n_2294)
);

BUFx6f_ASAP7_75t_L g2295 ( 
.A(n_1698),
.Y(n_2295)
);

INVx5_ASAP7_75t_L g2296 ( 
.A(n_1913),
.Y(n_2296)
);

OR2x6_ASAP7_75t_L g2297 ( 
.A(n_1836),
.B(n_1907),
.Y(n_2297)
);

NAND2xp5_ASAP7_75t_L g2298 ( 
.A(n_1849),
.B(n_252),
.Y(n_2298)
);

INVxp67_ASAP7_75t_L g2299 ( 
.A(n_1806),
.Y(n_2299)
);

NOR2x1_ASAP7_75t_L g2300 ( 
.A(n_1716),
.B(n_252),
.Y(n_2300)
);

BUFx3_ASAP7_75t_L g2301 ( 
.A(n_1761),
.Y(n_2301)
);

AND2x2_ASAP7_75t_L g2302 ( 
.A(n_1813),
.B(n_253),
.Y(n_2302)
);

INVx5_ASAP7_75t_L g2303 ( 
.A(n_1913),
.Y(n_2303)
);

CKINVDCx16_ASAP7_75t_R g2304 ( 
.A(n_1983),
.Y(n_2304)
);

AND2x4_ASAP7_75t_L g2305 ( 
.A(n_2026),
.B(n_253),
.Y(n_2305)
);

AND2x2_ASAP7_75t_L g2306 ( 
.A(n_1821),
.B(n_254),
.Y(n_2306)
);

BUFx12f_ASAP7_75t_L g2307 ( 
.A(n_1977),
.Y(n_2307)
);

INVx2_ASAP7_75t_L g2308 ( 
.A(n_1737),
.Y(n_2308)
);

BUFx3_ASAP7_75t_L g2309 ( 
.A(n_1761),
.Y(n_2309)
);

AND2x2_ASAP7_75t_L g2310 ( 
.A(n_1821),
.B(n_254),
.Y(n_2310)
);

NOR2xp67_ASAP7_75t_SL g2311 ( 
.A(n_1716),
.B(n_255),
.Y(n_2311)
);

BUFx2_ASAP7_75t_L g2312 ( 
.A(n_1907),
.Y(n_2312)
);

OR2x6_ASAP7_75t_L g2313 ( 
.A(n_1907),
.B(n_255),
.Y(n_2313)
);

BUFx3_ASAP7_75t_L g2314 ( 
.A(n_1757),
.Y(n_2314)
);

NOR2xp67_ASAP7_75t_L g2315 ( 
.A(n_1728),
.B(n_1913),
.Y(n_2315)
);

AND2x4_ASAP7_75t_L g2316 ( 
.A(n_1941),
.B(n_256),
.Y(n_2316)
);

INVx1_ASAP7_75t_L g2317 ( 
.A(n_1898),
.Y(n_2317)
);

INVx1_ASAP7_75t_L g2318 ( 
.A(n_1905),
.Y(n_2318)
);

NOR2x1_ASAP7_75t_L g2319 ( 
.A(n_1728),
.B(n_256),
.Y(n_2319)
);

BUFx2_ASAP7_75t_L g2320 ( 
.A(n_1775),
.Y(n_2320)
);

OR2x6_ASAP7_75t_L g2321 ( 
.A(n_1775),
.B(n_258),
.Y(n_2321)
);

OR2x2_ASAP7_75t_L g2322 ( 
.A(n_2016),
.B(n_2019),
.Y(n_2322)
);

INVxp67_ASAP7_75t_L g2323 ( 
.A(n_1806),
.Y(n_2323)
);

INVx1_ASAP7_75t_L g2324 ( 
.A(n_1905),
.Y(n_2324)
);

INVx1_ASAP7_75t_L g2325 ( 
.A(n_1912),
.Y(n_2325)
);

AND2x6_ASAP7_75t_L g2326 ( 
.A(n_1775),
.B(n_259),
.Y(n_2326)
);

INVx1_ASAP7_75t_L g2327 ( 
.A(n_1912),
.Y(n_2327)
);

AND2x2_ASAP7_75t_L g2328 ( 
.A(n_2012),
.B(n_259),
.Y(n_2328)
);

NAND2xp5_ASAP7_75t_SL g2329 ( 
.A(n_1755),
.B(n_260),
.Y(n_2329)
);

HB1xp67_ASAP7_75t_L g2330 ( 
.A(n_1784),
.Y(n_2330)
);

INVx2_ASAP7_75t_L g2331 ( 
.A(n_1751),
.Y(n_2331)
);

INVx1_ASAP7_75t_SL g2332 ( 
.A(n_1784),
.Y(n_2332)
);

NAND2xp5_ASAP7_75t_L g2333 ( 
.A(n_1849),
.B(n_260),
.Y(n_2333)
);

BUFx2_ASAP7_75t_L g2334 ( 
.A(n_1784),
.Y(n_2334)
);

NAND2xp5_ASAP7_75t_L g2335 ( 
.A(n_1856),
.B(n_261),
.Y(n_2335)
);

INVx2_ASAP7_75t_L g2336 ( 
.A(n_1751),
.Y(n_2336)
);

AND2x4_ASAP7_75t_L g2337 ( 
.A(n_1941),
.B(n_261),
.Y(n_2337)
);

NAND2xp5_ASAP7_75t_L g2338 ( 
.A(n_1856),
.B(n_263),
.Y(n_2338)
);

NAND2x1p5_ASAP7_75t_L g2339 ( 
.A(n_1997),
.B(n_263),
.Y(n_2339)
);

INVx1_ASAP7_75t_L g2340 ( 
.A(n_1899),
.Y(n_2340)
);

INVx2_ASAP7_75t_L g2341 ( 
.A(n_1773),
.Y(n_2341)
);

NAND2x1p5_ASAP7_75t_L g2342 ( 
.A(n_1997),
.B(n_264),
.Y(n_2342)
);

BUFx4f_ASAP7_75t_L g2343 ( 
.A(n_1831),
.Y(n_2343)
);

BUFx6f_ASAP7_75t_L g2344 ( 
.A(n_1937),
.Y(n_2344)
);

BUFx2_ASAP7_75t_SL g2345 ( 
.A(n_1997),
.Y(n_2345)
);

HB1xp67_ASAP7_75t_L g2346 ( 
.A(n_1840),
.Y(n_2346)
);

NAND2xp5_ASAP7_75t_L g2347 ( 
.A(n_1872),
.B(n_264),
.Y(n_2347)
);

BUFx3_ASAP7_75t_L g2348 ( 
.A(n_1757),
.Y(n_2348)
);

OR2x2_ASAP7_75t_L g2349 ( 
.A(n_2019),
.B(n_265),
.Y(n_2349)
);

NAND2xp5_ASAP7_75t_L g2350 ( 
.A(n_1872),
.B(n_265),
.Y(n_2350)
);

OR2x6_ASAP7_75t_SL g2351 ( 
.A(n_2018),
.B(n_266),
.Y(n_2351)
);

BUFx2_ASAP7_75t_L g2352 ( 
.A(n_1840),
.Y(n_2352)
);

INVx2_ASAP7_75t_L g2353 ( 
.A(n_1773),
.Y(n_2353)
);

AND2x2_ASAP7_75t_L g2354 ( 
.A(n_2012),
.B(n_266),
.Y(n_2354)
);

INVxp67_ASAP7_75t_L g2355 ( 
.A(n_1696),
.Y(n_2355)
);

INVx3_ASAP7_75t_L g2356 ( 
.A(n_1893),
.Y(n_2356)
);

AND2x2_ASAP7_75t_L g2357 ( 
.A(n_1811),
.B(n_267),
.Y(n_2357)
);

AND2x6_ASAP7_75t_L g2358 ( 
.A(n_1728),
.B(n_267),
.Y(n_2358)
);

NAND2x1p5_ASAP7_75t_L g2359 ( 
.A(n_1988),
.B(n_269),
.Y(n_2359)
);

INVx1_ASAP7_75t_L g2360 ( 
.A(n_1782),
.Y(n_2360)
);

INVx2_ASAP7_75t_L g2361 ( 
.A(n_2028),
.Y(n_2361)
);

INVx2_ASAP7_75t_L g2362 ( 
.A(n_2028),
.Y(n_2362)
);

INVx1_ASAP7_75t_L g2363 ( 
.A(n_1705),
.Y(n_2363)
);

BUFx8_ASAP7_75t_L g2364 ( 
.A(n_1977),
.Y(n_2364)
);

AND2x4_ASAP7_75t_L g2365 ( 
.A(n_1887),
.B(n_269),
.Y(n_2365)
);

AND2x2_ASAP7_75t_L g2366 ( 
.A(n_1830),
.B(n_270),
.Y(n_2366)
);

AND2x2_ASAP7_75t_L g2367 ( 
.A(n_1837),
.B(n_270),
.Y(n_2367)
);

INVx6_ASAP7_75t_L g2368 ( 
.A(n_1990),
.Y(n_2368)
);

NOR2x1_ASAP7_75t_L g2369 ( 
.A(n_1925),
.B(n_271),
.Y(n_2369)
);

AND2x6_ASAP7_75t_L g2370 ( 
.A(n_1969),
.B(n_1925),
.Y(n_2370)
);

INVx3_ASAP7_75t_L g2371 ( 
.A(n_1893),
.Y(n_2371)
);

BUFx8_ASAP7_75t_L g2372 ( 
.A(n_1979),
.Y(n_2372)
);

AND2x4_ASAP7_75t_L g2373 ( 
.A(n_1969),
.B(n_271),
.Y(n_2373)
);

BUFx5_ASAP7_75t_L g2374 ( 
.A(n_1800),
.Y(n_2374)
);

INVx2_ASAP7_75t_L g2375 ( 
.A(n_1740),
.Y(n_2375)
);

NAND2xp5_ASAP7_75t_L g2376 ( 
.A(n_1706),
.B(n_272),
.Y(n_2376)
);

INVx1_ASAP7_75t_SL g2377 ( 
.A(n_2025),
.Y(n_2377)
);

OR2x2_ASAP7_75t_L g2378 ( 
.A(n_1990),
.B(n_274),
.Y(n_2378)
);

AND2x4_ASAP7_75t_L g2379 ( 
.A(n_1969),
.B(n_1726),
.Y(n_2379)
);

INVx2_ASAP7_75t_L g2380 ( 
.A(n_1740),
.Y(n_2380)
);

AND2x4_ASAP7_75t_L g2381 ( 
.A(n_1969),
.B(n_274),
.Y(n_2381)
);

NAND2xp5_ASAP7_75t_L g2382 ( 
.A(n_1895),
.B(n_276),
.Y(n_2382)
);

AND2x4_ASAP7_75t_L g2383 ( 
.A(n_1730),
.B(n_277),
.Y(n_2383)
);

AND2x4_ASAP7_75t_L g2384 ( 
.A(n_1776),
.B(n_277),
.Y(n_2384)
);

NOR2xp33_ASAP7_75t_L g2385 ( 
.A(n_1847),
.B(n_278),
.Y(n_2385)
);

INVx3_ASAP7_75t_L g2386 ( 
.A(n_1893),
.Y(n_2386)
);

AND2x2_ASAP7_75t_L g2387 ( 
.A(n_1988),
.B(n_278),
.Y(n_2387)
);

AND2x4_ASAP7_75t_L g2388 ( 
.A(n_1855),
.B(n_279),
.Y(n_2388)
);

BUFx2_ASAP7_75t_L g2389 ( 
.A(n_2027),
.Y(n_2389)
);

INVx3_ASAP7_75t_L g2390 ( 
.A(n_1893),
.Y(n_2390)
);

AND2x2_ASAP7_75t_L g2391 ( 
.A(n_1992),
.B(n_279),
.Y(n_2391)
);

HB1xp67_ASAP7_75t_L g2392 ( 
.A(n_2029),
.Y(n_2392)
);

CKINVDCx5p33_ASAP7_75t_R g2393 ( 
.A(n_1911),
.Y(n_2393)
);

AND2x2_ASAP7_75t_L g2394 ( 
.A(n_1886),
.B(n_280),
.Y(n_2394)
);

BUFx2_ASAP7_75t_L g2395 ( 
.A(n_1863),
.Y(n_2395)
);

AND2x4_ASAP7_75t_L g2396 ( 
.A(n_1804),
.B(n_282),
.Y(n_2396)
);

OR2x2_ASAP7_75t_L g2397 ( 
.A(n_1764),
.B(n_282),
.Y(n_2397)
);

NAND2xp5_ASAP7_75t_L g2398 ( 
.A(n_1706),
.B(n_283),
.Y(n_2398)
);

BUFx8_ASAP7_75t_SL g2399 ( 
.A(n_2021),
.Y(n_2399)
);

AND2x4_ASAP7_75t_L g2400 ( 
.A(n_1747),
.B(n_1930),
.Y(n_2400)
);

INVx2_ASAP7_75t_L g2401 ( 
.A(n_1740),
.Y(n_2401)
);

CKINVDCx6p67_ASAP7_75t_R g2402 ( 
.A(n_1994),
.Y(n_2402)
);

AND2x2_ASAP7_75t_L g2403 ( 
.A(n_1982),
.B(n_284),
.Y(n_2403)
);

INVx6_ASAP7_75t_L g2404 ( 
.A(n_1985),
.Y(n_2404)
);

INVx4_ASAP7_75t_L g2405 ( 
.A(n_1831),
.Y(n_2405)
);

NAND2x1p5_ASAP7_75t_L g2406 ( 
.A(n_1860),
.B(n_284),
.Y(n_2406)
);

INVx3_ASAP7_75t_L g2407 ( 
.A(n_1770),
.Y(n_2407)
);

BUFx3_ASAP7_75t_L g2408 ( 
.A(n_1958),
.Y(n_2408)
);

HB1xp67_ASAP7_75t_L g2409 ( 
.A(n_1863),
.Y(n_2409)
);

AND2x2_ASAP7_75t_L g2410 ( 
.A(n_1771),
.B(n_285),
.Y(n_2410)
);

NOR2xp33_ASAP7_75t_SL g2411 ( 
.A(n_1948),
.B(n_489),
.Y(n_2411)
);

NOR2xp33_ASAP7_75t_L g2412 ( 
.A(n_1793),
.B(n_285),
.Y(n_2412)
);

OR2x2_ASAP7_75t_L g2413 ( 
.A(n_1947),
.B(n_1805),
.Y(n_2413)
);

INVx1_ASAP7_75t_SL g2414 ( 
.A(n_1910),
.Y(n_2414)
);

BUFx6f_ASAP7_75t_L g2415 ( 
.A(n_1937),
.Y(n_2415)
);

HB1xp67_ASAP7_75t_L g2416 ( 
.A(n_1928),
.Y(n_2416)
);

AND2x4_ASAP7_75t_L g2417 ( 
.A(n_1943),
.B(n_286),
.Y(n_2417)
);

BUFx2_ASAP7_75t_L g2418 ( 
.A(n_1987),
.Y(n_2418)
);

NAND2xp5_ASAP7_75t_L g2419 ( 
.A(n_1925),
.B(n_286),
.Y(n_2419)
);

CKINVDCx5p33_ASAP7_75t_R g2420 ( 
.A(n_1994),
.Y(n_2420)
);

INVx1_ASAP7_75t_L g2421 ( 
.A(n_1910),
.Y(n_2421)
);

AND2x2_ASAP7_75t_L g2422 ( 
.A(n_1860),
.B(n_1720),
.Y(n_2422)
);

AND2x4_ASAP7_75t_L g2423 ( 
.A(n_1800),
.B(n_288),
.Y(n_2423)
);

INVx3_ASAP7_75t_L g2424 ( 
.A(n_1770),
.Y(n_2424)
);

AND2x2_ASAP7_75t_L g2425 ( 
.A(n_1762),
.B(n_288),
.Y(n_2425)
);

AND2x4_ASAP7_75t_L g2426 ( 
.A(n_1820),
.B(n_1822),
.Y(n_2426)
);

BUFx6f_ASAP7_75t_L g2427 ( 
.A(n_1937),
.Y(n_2427)
);

AND2x2_ASAP7_75t_L g2428 ( 
.A(n_1947),
.B(n_1914),
.Y(n_2428)
);

NOR2xp33_ASAP7_75t_L g2429 ( 
.A(n_1918),
.B(n_289),
.Y(n_2429)
);

HB1xp67_ASAP7_75t_L g2430 ( 
.A(n_1991),
.Y(n_2430)
);

NOR2x1_ASAP7_75t_L g2431 ( 
.A(n_1915),
.B(n_290),
.Y(n_2431)
);

INVx3_ASAP7_75t_L g2432 ( 
.A(n_1770),
.Y(n_2432)
);

NOR2xp33_ASAP7_75t_L g2433 ( 
.A(n_1927),
.B(n_291),
.Y(n_2433)
);

AND2x2_ASAP7_75t_L g2434 ( 
.A(n_1958),
.B(n_291),
.Y(n_2434)
);

NAND2xp5_ASAP7_75t_L g2435 ( 
.A(n_2031),
.B(n_292),
.Y(n_2435)
);

BUFx4f_ASAP7_75t_L g2436 ( 
.A(n_1809),
.Y(n_2436)
);

INVx2_ASAP7_75t_L g2437 ( 
.A(n_1792),
.Y(n_2437)
);

HB1xp67_ASAP7_75t_L g2438 ( 
.A(n_1850),
.Y(n_2438)
);

NOR2xp33_ASAP7_75t_SL g2439 ( 
.A(n_1753),
.B(n_490),
.Y(n_2439)
);

INVx1_ASAP7_75t_L g2440 ( 
.A(n_1820),
.Y(n_2440)
);

NAND2xp5_ASAP7_75t_L g2441 ( 
.A(n_2031),
.B(n_292),
.Y(n_2441)
);

NAND2xp5_ASAP7_75t_L g2442 ( 
.A(n_1881),
.B(n_1906),
.Y(n_2442)
);

INVx6_ASAP7_75t_L g2443 ( 
.A(n_1946),
.Y(n_2443)
);

BUFx6f_ASAP7_75t_L g2444 ( 
.A(n_1937),
.Y(n_2444)
);

BUFx2_ASAP7_75t_L g2445 ( 
.A(n_1842),
.Y(n_2445)
);

OR2x2_ASAP7_75t_L g2446 ( 
.A(n_1853),
.B(n_293),
.Y(n_2446)
);

AND2x2_ASAP7_75t_L g2447 ( 
.A(n_1888),
.B(n_293),
.Y(n_2447)
);

NAND2xp5_ASAP7_75t_L g2448 ( 
.A(n_1881),
.B(n_294),
.Y(n_2448)
);

AND2x4_ASAP7_75t_L g2449 ( 
.A(n_1822),
.B(n_295),
.Y(n_2449)
);

NAND2xp5_ASAP7_75t_L g2450 ( 
.A(n_1801),
.B(n_295),
.Y(n_2450)
);

INVx4_ASAP7_75t_L g2451 ( 
.A(n_1792),
.Y(n_2451)
);

NOR2xp33_ASAP7_75t_L g2452 ( 
.A(n_2020),
.B(n_1884),
.Y(n_2452)
);

AND2x2_ASAP7_75t_L g2453 ( 
.A(n_1865),
.B(n_296),
.Y(n_2453)
);

INVx3_ASAP7_75t_L g2454 ( 
.A(n_1792),
.Y(n_2454)
);

BUFx3_ASAP7_75t_L g2455 ( 
.A(n_1951),
.Y(n_2455)
);

INVx1_ASAP7_75t_L g2456 ( 
.A(n_1823),
.Y(n_2456)
);

NAND2xp5_ASAP7_75t_L g2457 ( 
.A(n_1754),
.B(n_296),
.Y(n_2457)
);

BUFx3_ASAP7_75t_L g2458 ( 
.A(n_1873),
.Y(n_2458)
);

INVx2_ASAP7_75t_L g2459 ( 
.A(n_1858),
.Y(n_2459)
);

NOR2xp33_ASAP7_75t_L g2460 ( 
.A(n_1929),
.B(n_297),
.Y(n_2460)
);

NAND2xp5_ASAP7_75t_SL g2461 ( 
.A(n_1923),
.B(n_297),
.Y(n_2461)
);

INVx2_ASAP7_75t_L g2462 ( 
.A(n_1858),
.Y(n_2462)
);

BUFx6f_ASAP7_75t_L g2463 ( 
.A(n_1938),
.Y(n_2463)
);

AND2x4_ASAP7_75t_L g2464 ( 
.A(n_1823),
.B(n_300),
.Y(n_2464)
);

AND2x4_ASAP7_75t_L g2465 ( 
.A(n_1829),
.B(n_300),
.Y(n_2465)
);

OR2x2_ASAP7_75t_L g2466 ( 
.A(n_1871),
.B(n_301),
.Y(n_2466)
);

INVx2_ASAP7_75t_L g2467 ( 
.A(n_1868),
.Y(n_2467)
);

INVx2_ASAP7_75t_L g2468 ( 
.A(n_1868),
.Y(n_2468)
);

AND2x2_ASAP7_75t_L g2469 ( 
.A(n_1901),
.B(n_303),
.Y(n_2469)
);

INVxp67_ASAP7_75t_L g2470 ( 
.A(n_1722),
.Y(n_2470)
);

NAND2x1p5_ASAP7_75t_L g2471 ( 
.A(n_2090),
.B(n_1889),
.Y(n_2471)
);

BUFx12f_ASAP7_75t_L g2472 ( 
.A(n_2130),
.Y(n_2472)
);

INVx2_ASAP7_75t_L g2473 ( 
.A(n_2040),
.Y(n_2473)
);

BUFx6f_ASAP7_75t_L g2474 ( 
.A(n_2037),
.Y(n_2474)
);

INVxp67_ASAP7_75t_SL g2475 ( 
.A(n_2189),
.Y(n_2475)
);

INVx1_ASAP7_75t_L g2476 ( 
.A(n_2067),
.Y(n_2476)
);

INVx1_ASAP7_75t_L g2477 ( 
.A(n_2048),
.Y(n_2477)
);

BUFx2_ASAP7_75t_L g2478 ( 
.A(n_2038),
.Y(n_2478)
);

AND2x4_ASAP7_75t_L g2479 ( 
.A(n_2223),
.B(n_1829),
.Y(n_2479)
);

INVx1_ASAP7_75t_L g2480 ( 
.A(n_2048),
.Y(n_2480)
);

BUFx3_ASAP7_75t_L g2481 ( 
.A(n_2046),
.Y(n_2481)
);

NAND2xp5_ASAP7_75t_L g2482 ( 
.A(n_2243),
.B(n_2009),
.Y(n_2482)
);

AOI22xp33_ASAP7_75t_L g2483 ( 
.A1(n_2166),
.A2(n_1906),
.B1(n_1796),
.B2(n_1919),
.Y(n_2483)
);

INVx1_ASAP7_75t_SL g2484 ( 
.A(n_2223),
.Y(n_2484)
);

INVx3_ASAP7_75t_SL g2485 ( 
.A(n_2079),
.Y(n_2485)
);

INVx5_ASAP7_75t_L g2486 ( 
.A(n_2223),
.Y(n_2486)
);

BUFx6f_ASAP7_75t_L g2487 ( 
.A(n_2037),
.Y(n_2487)
);

INVx1_ASAP7_75t_SL g2488 ( 
.A(n_2297),
.Y(n_2488)
);

AND2x2_ASAP7_75t_L g2489 ( 
.A(n_2166),
.B(n_1724),
.Y(n_2489)
);

NAND2x1p5_ASAP7_75t_L g2490 ( 
.A(n_2090),
.B(n_2158),
.Y(n_2490)
);

INVx1_ASAP7_75t_SL g2491 ( 
.A(n_2297),
.Y(n_2491)
);

INVx5_ASAP7_75t_L g2492 ( 
.A(n_2297),
.Y(n_2492)
);

AND2x2_ASAP7_75t_L g2493 ( 
.A(n_2218),
.B(n_2328),
.Y(n_2493)
);

BUFx2_ASAP7_75t_L g2494 ( 
.A(n_2038),
.Y(n_2494)
);

BUFx3_ASAP7_75t_L g2495 ( 
.A(n_2152),
.Y(n_2495)
);

AO22x1_ASAP7_75t_L g2496 ( 
.A1(n_2364),
.A2(n_1995),
.B1(n_1967),
.B2(n_1756),
.Y(n_2496)
);

INVx2_ASAP7_75t_L g2497 ( 
.A(n_2047),
.Y(n_2497)
);

NAND2xp5_ASAP7_75t_SL g2498 ( 
.A(n_2142),
.B(n_2143),
.Y(n_2498)
);

INVx1_ASAP7_75t_L g2499 ( 
.A(n_2060),
.Y(n_2499)
);

INVx1_ASAP7_75t_L g2500 ( 
.A(n_2060),
.Y(n_2500)
);

INVx2_ASAP7_75t_L g2501 ( 
.A(n_2100),
.Y(n_2501)
);

NAND2xp5_ASAP7_75t_L g2502 ( 
.A(n_2103),
.B(n_2009),
.Y(n_2502)
);

INVx1_ASAP7_75t_L g2503 ( 
.A(n_2103),
.Y(n_2503)
);

INVx1_ASAP7_75t_L g2504 ( 
.A(n_2077),
.Y(n_2504)
);

HB1xp67_ASAP7_75t_L g2505 ( 
.A(n_2189),
.Y(n_2505)
);

INVx5_ASAP7_75t_L g2506 ( 
.A(n_2078),
.Y(n_2506)
);

INVx3_ASAP7_75t_L g2507 ( 
.A(n_2070),
.Y(n_2507)
);

BUFx3_ASAP7_75t_L g2508 ( 
.A(n_2082),
.Y(n_2508)
);

NAND2xp5_ASAP7_75t_L g2509 ( 
.A(n_2148),
.B(n_2013),
.Y(n_2509)
);

BUFx3_ASAP7_75t_L g2510 ( 
.A(n_2097),
.Y(n_2510)
);

BUFx12f_ASAP7_75t_L g2511 ( 
.A(n_2270),
.Y(n_2511)
);

INVx2_ASAP7_75t_SL g2512 ( 
.A(n_2127),
.Y(n_2512)
);

INVx5_ASAP7_75t_L g2513 ( 
.A(n_2078),
.Y(n_2513)
);

BUFx6f_ASAP7_75t_L g2514 ( 
.A(n_2037),
.Y(n_2514)
);

NOR2xp33_ASAP7_75t_L g2515 ( 
.A(n_2422),
.B(n_1718),
.Y(n_2515)
);

INVx1_ASAP7_75t_L g2516 ( 
.A(n_2109),
.Y(n_2516)
);

BUFx6f_ASAP7_75t_L g2517 ( 
.A(n_2066),
.Y(n_2517)
);

INVx8_ASAP7_75t_L g2518 ( 
.A(n_2038),
.Y(n_2518)
);

INVx1_ASAP7_75t_L g2519 ( 
.A(n_2114),
.Y(n_2519)
);

INVx3_ASAP7_75t_SL g2520 ( 
.A(n_2039),
.Y(n_2520)
);

BUFx12f_ASAP7_75t_L g2521 ( 
.A(n_2039),
.Y(n_2521)
);

BUFx6f_ASAP7_75t_L g2522 ( 
.A(n_2066),
.Y(n_2522)
);

BUFx2_ASAP7_75t_SL g2523 ( 
.A(n_2158),
.Y(n_2523)
);

INVx3_ASAP7_75t_L g2524 ( 
.A(n_2070),
.Y(n_2524)
);

BUFx2_ASAP7_75t_SL g2525 ( 
.A(n_2158),
.Y(n_2525)
);

BUFx6f_ASAP7_75t_L g2526 ( 
.A(n_2066),
.Y(n_2526)
);

AO21x2_ASAP7_75t_L g2527 ( 
.A1(n_2065),
.A2(n_1968),
.B(n_1838),
.Y(n_2527)
);

INVx2_ASAP7_75t_L g2528 ( 
.A(n_2104),
.Y(n_2528)
);

NAND2x1p5_ASAP7_75t_L g2529 ( 
.A(n_2153),
.B(n_1889),
.Y(n_2529)
);

AOI22xp5_ASAP7_75t_L g2530 ( 
.A1(n_2068),
.A2(n_1756),
.B1(n_1995),
.B2(n_1967),
.Y(n_2530)
);

INVx2_ASAP7_75t_L g2531 ( 
.A(n_2119),
.Y(n_2531)
);

INVx1_ASAP7_75t_L g2532 ( 
.A(n_2122),
.Y(n_2532)
);

INVx2_ASAP7_75t_L g2533 ( 
.A(n_2126),
.Y(n_2533)
);

BUFx3_ASAP7_75t_L g2534 ( 
.A(n_2134),
.Y(n_2534)
);

INVx1_ASAP7_75t_SL g2535 ( 
.A(n_2055),
.Y(n_2535)
);

AND2x2_ASAP7_75t_L g2536 ( 
.A(n_2218),
.B(n_1902),
.Y(n_2536)
);

INVx2_ASAP7_75t_SL g2537 ( 
.A(n_2279),
.Y(n_2537)
);

INVx2_ASAP7_75t_L g2538 ( 
.A(n_2137),
.Y(n_2538)
);

INVx3_ASAP7_75t_L g2539 ( 
.A(n_2072),
.Y(n_2539)
);

BUFx2_ASAP7_75t_L g2540 ( 
.A(n_2364),
.Y(n_2540)
);

BUFx6f_ASAP7_75t_L g2541 ( 
.A(n_2140),
.Y(n_2541)
);

BUFx4_ASAP7_75t_SL g2542 ( 
.A(n_2039),
.Y(n_2542)
);

BUFx2_ASAP7_75t_SL g2543 ( 
.A(n_2058),
.Y(n_2543)
);

BUFx2_ASAP7_75t_L g2544 ( 
.A(n_2078),
.Y(n_2544)
);

BUFx12f_ASAP7_75t_L g2545 ( 
.A(n_2248),
.Y(n_2545)
);

INVx6_ASAP7_75t_SL g2546 ( 
.A(n_2099),
.Y(n_2546)
);

AOI22xp33_ASAP7_75t_L g2547 ( 
.A1(n_2343),
.A2(n_2013),
.B1(n_1975),
.B2(n_1783),
.Y(n_2547)
);

INVx6_ASAP7_75t_L g2548 ( 
.A(n_2062),
.Y(n_2548)
);

INVx1_ASAP7_75t_L g2549 ( 
.A(n_2131),
.Y(n_2549)
);

INVx3_ASAP7_75t_L g2550 ( 
.A(n_2072),
.Y(n_2550)
);

BUFx12f_ASAP7_75t_L g2551 ( 
.A(n_2285),
.Y(n_2551)
);

INVx1_ASAP7_75t_L g2552 ( 
.A(n_2141),
.Y(n_2552)
);

INVx1_ASAP7_75t_L g2553 ( 
.A(n_2150),
.Y(n_2553)
);

BUFx3_ASAP7_75t_L g2554 ( 
.A(n_2237),
.Y(n_2554)
);

AND2x2_ASAP7_75t_L g2555 ( 
.A(n_2354),
.B(n_1904),
.Y(n_2555)
);

INVx5_ASAP7_75t_L g2556 ( 
.A(n_2099),
.Y(n_2556)
);

CKINVDCx5p33_ASAP7_75t_R g2557 ( 
.A(n_2192),
.Y(n_2557)
);

INVx1_ASAP7_75t_L g2558 ( 
.A(n_2171),
.Y(n_2558)
);

INVx1_ASAP7_75t_L g2559 ( 
.A(n_2186),
.Y(n_2559)
);

BUFx6f_ASAP7_75t_L g2560 ( 
.A(n_2140),
.Y(n_2560)
);

INVx2_ASAP7_75t_L g2561 ( 
.A(n_2168),
.Y(n_2561)
);

INVx1_ASAP7_75t_L g2562 ( 
.A(n_2194),
.Y(n_2562)
);

BUFx3_ASAP7_75t_L g2563 ( 
.A(n_2314),
.Y(n_2563)
);

INVx1_ASAP7_75t_SL g2564 ( 
.A(n_2055),
.Y(n_2564)
);

BUFx2_ASAP7_75t_SL g2565 ( 
.A(n_2058),
.Y(n_2565)
);

INVx2_ASAP7_75t_SL g2566 ( 
.A(n_2062),
.Y(n_2566)
);

INVx1_ASAP7_75t_SL g2567 ( 
.A(n_2259),
.Y(n_2567)
);

BUFx12f_ASAP7_75t_L g2568 ( 
.A(n_2288),
.Y(n_2568)
);

INVx3_ASAP7_75t_L g2569 ( 
.A(n_2087),
.Y(n_2569)
);

INVx2_ASAP7_75t_SL g2570 ( 
.A(n_2192),
.Y(n_2570)
);

AND2x2_ASAP7_75t_L g2571 ( 
.A(n_2343),
.B(n_1692),
.Y(n_2571)
);

INVx3_ASAP7_75t_SL g2572 ( 
.A(n_2182),
.Y(n_2572)
);

BUFx3_ASAP7_75t_L g2573 ( 
.A(n_2348),
.Y(n_2573)
);

INVx1_ASAP7_75t_SL g2574 ( 
.A(n_2259),
.Y(n_2574)
);

BUFx2_ASAP7_75t_L g2575 ( 
.A(n_2099),
.Y(n_2575)
);

INVx1_ASAP7_75t_L g2576 ( 
.A(n_2204),
.Y(n_2576)
);

INVx1_ASAP7_75t_L g2577 ( 
.A(n_2209),
.Y(n_2577)
);

BUFx6f_ASAP7_75t_L g2578 ( 
.A(n_2140),
.Y(n_2578)
);

INVx1_ASAP7_75t_SL g2579 ( 
.A(n_2332),
.Y(n_2579)
);

INVx3_ASAP7_75t_L g2580 ( 
.A(n_2087),
.Y(n_2580)
);

INVx8_ASAP7_75t_L g2581 ( 
.A(n_2117),
.Y(n_2581)
);

BUFx8_ASAP7_75t_SL g2582 ( 
.A(n_2399),
.Y(n_2582)
);

INVx1_ASAP7_75t_L g2583 ( 
.A(n_2210),
.Y(n_2583)
);

INVx4_ASAP7_75t_L g2584 ( 
.A(n_2117),
.Y(n_2584)
);

BUFx10_ASAP7_75t_L g2585 ( 
.A(n_2061),
.Y(n_2585)
);

BUFx12f_ASAP7_75t_L g2586 ( 
.A(n_2112),
.Y(n_2586)
);

BUFx12f_ASAP7_75t_L g2587 ( 
.A(n_2044),
.Y(n_2587)
);

INVx3_ASAP7_75t_L g2588 ( 
.A(n_2154),
.Y(n_2588)
);

BUFx3_ASAP7_75t_L g2589 ( 
.A(n_2224),
.Y(n_2589)
);

INVx3_ASAP7_75t_L g2590 ( 
.A(n_2154),
.Y(n_2590)
);

NAND2xp5_ASAP7_75t_L g2591 ( 
.A(n_2442),
.B(n_1923),
.Y(n_2591)
);

INVx3_ASAP7_75t_L g2592 ( 
.A(n_2159),
.Y(n_2592)
);

AND2x4_ASAP7_75t_L g2593 ( 
.A(n_2033),
.B(n_1929),
.Y(n_2593)
);

INVx4_ASAP7_75t_L g2594 ( 
.A(n_2117),
.Y(n_2594)
);

INVx1_ASAP7_75t_L g2595 ( 
.A(n_2238),
.Y(n_2595)
);

INVx1_ASAP7_75t_SL g2596 ( 
.A(n_2332),
.Y(n_2596)
);

INVx5_ASAP7_75t_L g2597 ( 
.A(n_2116),
.Y(n_2597)
);

INVx1_ASAP7_75t_L g2598 ( 
.A(n_2340),
.Y(n_2598)
);

INVx4_ASAP7_75t_L g2599 ( 
.A(n_2177),
.Y(n_2599)
);

HB1xp67_ASAP7_75t_L g2600 ( 
.A(n_2177),
.Y(n_2600)
);

INVx1_ASAP7_75t_L g2601 ( 
.A(n_2105),
.Y(n_2601)
);

BUFx4f_ASAP7_75t_L g2602 ( 
.A(n_2177),
.Y(n_2602)
);

INVx3_ASAP7_75t_L g2603 ( 
.A(n_2159),
.Y(n_2603)
);

INVx1_ASAP7_75t_SL g2604 ( 
.A(n_2211),
.Y(n_2604)
);

BUFx12f_ASAP7_75t_L g2605 ( 
.A(n_2052),
.Y(n_2605)
);

INVx2_ASAP7_75t_L g2606 ( 
.A(n_2459),
.Y(n_2606)
);

INVx1_ASAP7_75t_SL g2607 ( 
.A(n_2352),
.Y(n_2607)
);

INVx2_ASAP7_75t_SL g2608 ( 
.A(n_2301),
.Y(n_2608)
);

AND2x2_ASAP7_75t_L g2609 ( 
.A(n_2402),
.B(n_2033),
.Y(n_2609)
);

NOR2xp33_ASAP7_75t_L g2610 ( 
.A(n_2069),
.B(n_1729),
.Y(n_2610)
);

INVx2_ASAP7_75t_L g2611 ( 
.A(n_2462),
.Y(n_2611)
);

AOI22xp33_ASAP7_75t_L g2612 ( 
.A1(n_2088),
.A2(n_1781),
.B1(n_1878),
.B2(n_1876),
.Y(n_2612)
);

BUFx3_ASAP7_75t_L g2613 ( 
.A(n_2368),
.Y(n_2613)
);

BUFx3_ASAP7_75t_L g2614 ( 
.A(n_2368),
.Y(n_2614)
);

CKINVDCx8_ASAP7_75t_R g2615 ( 
.A(n_2304),
.Y(n_2615)
);

INVx3_ASAP7_75t_L g2616 ( 
.A(n_2153),
.Y(n_2616)
);

BUFx12f_ASAP7_75t_L g2617 ( 
.A(n_2284),
.Y(n_2617)
);

BUFx12f_ASAP7_75t_L g2618 ( 
.A(n_2307),
.Y(n_2618)
);

BUFx3_ASAP7_75t_L g2619 ( 
.A(n_2309),
.Y(n_2619)
);

INVx1_ASAP7_75t_SL g2620 ( 
.A(n_2197),
.Y(n_2620)
);

INVx3_ASAP7_75t_L g2621 ( 
.A(n_2165),
.Y(n_2621)
);

INVx5_ASAP7_75t_SL g2622 ( 
.A(n_2116),
.Y(n_2622)
);

NOR2xp33_ASAP7_75t_L g2623 ( 
.A(n_2098),
.B(n_1882),
.Y(n_2623)
);

BUFx12f_ASAP7_75t_L g2624 ( 
.A(n_2372),
.Y(n_2624)
);

INVx1_ASAP7_75t_SL g2625 ( 
.A(n_2197),
.Y(n_2625)
);

INVx4_ASAP7_75t_L g2626 ( 
.A(n_2197),
.Y(n_2626)
);

NAND2xp5_ASAP7_75t_L g2627 ( 
.A(n_2175),
.B(n_1923),
.Y(n_2627)
);

NAND2xp5_ASAP7_75t_L g2628 ( 
.A(n_2421),
.B(n_1923),
.Y(n_2628)
);

INVx1_ASAP7_75t_L g2629 ( 
.A(n_2105),
.Y(n_2629)
);

CKINVDCx5p33_ASAP7_75t_R g2630 ( 
.A(n_2123),
.Y(n_2630)
);

BUFx12f_ASAP7_75t_L g2631 ( 
.A(n_2372),
.Y(n_2631)
);

BUFx12f_ASAP7_75t_L g2632 ( 
.A(n_2032),
.Y(n_2632)
);

INVx2_ASAP7_75t_SL g2633 ( 
.A(n_2161),
.Y(n_2633)
);

INVx3_ASAP7_75t_L g2634 ( 
.A(n_2165),
.Y(n_2634)
);

BUFx3_ASAP7_75t_L g2635 ( 
.A(n_2110),
.Y(n_2635)
);

BUFx3_ASAP7_75t_L g2636 ( 
.A(n_2124),
.Y(n_2636)
);

OR2x6_ASAP7_75t_L g2637 ( 
.A(n_2282),
.B(n_1944),
.Y(n_2637)
);

BUFx6f_ASAP7_75t_L g2638 ( 
.A(n_2147),
.Y(n_2638)
);

BUFx6f_ASAP7_75t_L g2639 ( 
.A(n_2147),
.Y(n_2639)
);

INVx1_ASAP7_75t_L g2640 ( 
.A(n_2198),
.Y(n_2640)
);

BUFx12f_ASAP7_75t_L g2641 ( 
.A(n_2035),
.Y(n_2641)
);

INVx1_ASAP7_75t_L g2642 ( 
.A(n_2198),
.Y(n_2642)
);

NAND2x1p5_ASAP7_75t_L g2643 ( 
.A(n_2272),
.B(n_1889),
.Y(n_2643)
);

BUFx3_ASAP7_75t_L g2644 ( 
.A(n_2161),
.Y(n_2644)
);

INVxp67_ASAP7_75t_SL g2645 ( 
.A(n_2207),
.Y(n_2645)
);

BUFx3_ASAP7_75t_L g2646 ( 
.A(n_2132),
.Y(n_2646)
);

BUFx3_ASAP7_75t_L g2647 ( 
.A(n_2236),
.Y(n_2647)
);

INVx4_ASAP7_75t_L g2648 ( 
.A(n_2282),
.Y(n_2648)
);

INVx1_ASAP7_75t_L g2649 ( 
.A(n_2203),
.Y(n_2649)
);

CKINVDCx11_ASAP7_75t_R g2650 ( 
.A(n_2351),
.Y(n_2650)
);

INVx2_ASAP7_75t_L g2651 ( 
.A(n_2467),
.Y(n_2651)
);

HB1xp67_ASAP7_75t_L g2652 ( 
.A(n_2282),
.Y(n_2652)
);

INVx2_ASAP7_75t_L g2653 ( 
.A(n_2468),
.Y(n_2653)
);

BUFx4_ASAP7_75t_SL g2654 ( 
.A(n_2116),
.Y(n_2654)
);

NAND2x1p5_ASAP7_75t_L g2655 ( 
.A(n_2276),
.B(n_1929),
.Y(n_2655)
);

BUFx6f_ASAP7_75t_L g2656 ( 
.A(n_2147),
.Y(n_2656)
);

INVx1_ASAP7_75t_L g2657 ( 
.A(n_2203),
.Y(n_2657)
);

AND2x2_ASAP7_75t_L g2658 ( 
.A(n_2428),
.B(n_1944),
.Y(n_2658)
);

INVx6_ASAP7_75t_SL g2659 ( 
.A(n_2292),
.Y(n_2659)
);

NAND2x1p5_ASAP7_75t_L g2660 ( 
.A(n_2312),
.B(n_1954),
.Y(n_2660)
);

NAND2x1p5_ASAP7_75t_L g2661 ( 
.A(n_2320),
.B(n_1954),
.Y(n_2661)
);

BUFx3_ASAP7_75t_L g2662 ( 
.A(n_2239),
.Y(n_2662)
);

BUFx4_ASAP7_75t_SL g2663 ( 
.A(n_2292),
.Y(n_2663)
);

INVx2_ASAP7_75t_L g2664 ( 
.A(n_2215),
.Y(n_2664)
);

INVx2_ASAP7_75t_L g2665 ( 
.A(n_2216),
.Y(n_2665)
);

BUFx5_ASAP7_75t_L g2666 ( 
.A(n_2370),
.Y(n_2666)
);

NAND2xp5_ASAP7_75t_L g2667 ( 
.A(n_2440),
.B(n_1697),
.Y(n_2667)
);

OR2x6_ASAP7_75t_L g2668 ( 
.A(n_2292),
.B(n_1760),
.Y(n_2668)
);

BUFx3_ASAP7_75t_L g2669 ( 
.A(n_2162),
.Y(n_2669)
);

INVx1_ASAP7_75t_L g2670 ( 
.A(n_2042),
.Y(n_2670)
);

BUFx2_ASAP7_75t_SL g2671 ( 
.A(n_2092),
.Y(n_2671)
);

NAND2x1p5_ASAP7_75t_L g2672 ( 
.A(n_2334),
.B(n_1850),
.Y(n_2672)
);

INVx6_ASAP7_75t_L g2673 ( 
.A(n_2266),
.Y(n_2673)
);

INVx2_ASAP7_75t_SL g2674 ( 
.A(n_2408),
.Y(n_2674)
);

BUFx3_ASAP7_75t_L g2675 ( 
.A(n_2173),
.Y(n_2675)
);

BUFx3_ASAP7_75t_L g2676 ( 
.A(n_2266),
.Y(n_2676)
);

INVx2_ASAP7_75t_L g2677 ( 
.A(n_2220),
.Y(n_2677)
);

CKINVDCx12_ASAP7_75t_R g2678 ( 
.A(n_2313),
.Y(n_2678)
);

INVx3_ASAP7_75t_L g2679 ( 
.A(n_2370),
.Y(n_2679)
);

BUFx8_ASAP7_75t_SL g2680 ( 
.A(n_2313),
.Y(n_2680)
);

INVx1_ASAP7_75t_L g2681 ( 
.A(n_2049),
.Y(n_2681)
);

INVx2_ASAP7_75t_SL g2682 ( 
.A(n_2061),
.Y(n_2682)
);

BUFx12f_ASAP7_75t_L g2683 ( 
.A(n_2393),
.Y(n_2683)
);

INVx2_ASAP7_75t_L g2684 ( 
.A(n_2250),
.Y(n_2684)
);

BUFx6f_ASAP7_75t_L g2685 ( 
.A(n_2344),
.Y(n_2685)
);

CKINVDCx16_ASAP7_75t_R g2686 ( 
.A(n_2304),
.Y(n_2686)
);

INVx2_ASAP7_75t_L g2687 ( 
.A(n_2275),
.Y(n_2687)
);

INVx5_ASAP7_75t_L g2688 ( 
.A(n_2313),
.Y(n_2688)
);

INVx2_ASAP7_75t_SL g2689 ( 
.A(n_2091),
.Y(n_2689)
);

BUFx6f_ASAP7_75t_L g2690 ( 
.A(n_2344),
.Y(n_2690)
);

BUFx8_ASAP7_75t_L g2691 ( 
.A(n_2057),
.Y(n_2691)
);

CKINVDCx6p67_ASAP7_75t_R g2692 ( 
.A(n_2321),
.Y(n_2692)
);

INVx2_ASAP7_75t_L g2693 ( 
.A(n_2308),
.Y(n_2693)
);

INVxp67_ASAP7_75t_SL g2694 ( 
.A(n_2330),
.Y(n_2694)
);

NAND2xp5_ASAP7_75t_L g2695 ( 
.A(n_2456),
.B(n_2430),
.Y(n_2695)
);

HB1xp67_ASAP7_75t_L g2696 ( 
.A(n_2321),
.Y(n_2696)
);

INVx1_ASAP7_75t_L g2697 ( 
.A(n_2316),
.Y(n_2697)
);

CKINVDCx5p33_ASAP7_75t_R g2698 ( 
.A(n_2420),
.Y(n_2698)
);

INVx4_ASAP7_75t_L g2699 ( 
.A(n_2321),
.Y(n_2699)
);

INVx2_ASAP7_75t_SL g2700 ( 
.A(n_2091),
.Y(n_2700)
);

BUFx3_ASAP7_75t_L g2701 ( 
.A(n_2266),
.Y(n_2701)
);

NAND2x1p5_ASAP7_75t_L g2702 ( 
.A(n_2179),
.B(n_1851),
.Y(n_2702)
);

INVx4_ASAP7_75t_L g2703 ( 
.A(n_2092),
.Y(n_2703)
);

NOR2xp33_ASAP7_75t_L g2704 ( 
.A(n_2111),
.B(n_1917),
.Y(n_2704)
);

BUFx4f_ASAP7_75t_SL g2705 ( 
.A(n_2092),
.Y(n_2705)
);

INVx1_ASAP7_75t_L g2706 ( 
.A(n_2316),
.Y(n_2706)
);

BUFx12f_ASAP7_75t_L g2707 ( 
.A(n_2151),
.Y(n_2707)
);

BUFx3_ASAP7_75t_L g2708 ( 
.A(n_2346),
.Y(n_2708)
);

BUFx2_ASAP7_75t_SL g2709 ( 
.A(n_2092),
.Y(n_2709)
);

INVx1_ASAP7_75t_SL g2710 ( 
.A(n_2053),
.Y(n_2710)
);

INVx2_ASAP7_75t_SL g2711 ( 
.A(n_2179),
.Y(n_2711)
);

BUFx6f_ASAP7_75t_L g2712 ( 
.A(n_2344),
.Y(n_2712)
);

INVx2_ASAP7_75t_L g2713 ( 
.A(n_2331),
.Y(n_2713)
);

INVx2_ASAP7_75t_SL g2714 ( 
.A(n_2287),
.Y(n_2714)
);

INVx3_ASAP7_75t_L g2715 ( 
.A(n_2370),
.Y(n_2715)
);

INVx1_ASAP7_75t_L g2716 ( 
.A(n_2337),
.Y(n_2716)
);

CKINVDCx5p33_ASAP7_75t_R g2717 ( 
.A(n_2322),
.Y(n_2717)
);

BUFx3_ASAP7_75t_L g2718 ( 
.A(n_2287),
.Y(n_2718)
);

INVx1_ASAP7_75t_L g2719 ( 
.A(n_2337),
.Y(n_2719)
);

INVx3_ASAP7_75t_L g2720 ( 
.A(n_2370),
.Y(n_2720)
);

INVx8_ASAP7_75t_L g2721 ( 
.A(n_2102),
.Y(n_2721)
);

CKINVDCx16_ASAP7_75t_R g2722 ( 
.A(n_2235),
.Y(n_2722)
);

AOI22xp33_ASAP7_75t_L g2723 ( 
.A1(n_2405),
.A2(n_1933),
.B1(n_2022),
.B2(n_1981),
.Y(n_2723)
);

INVx2_ASAP7_75t_L g2724 ( 
.A(n_2336),
.Y(n_2724)
);

HB1xp67_ASAP7_75t_L g2725 ( 
.A(n_2438),
.Y(n_2725)
);

BUFx6f_ASAP7_75t_L g2726 ( 
.A(n_2415),
.Y(n_2726)
);

OR2x2_ASAP7_75t_L g2727 ( 
.A(n_2222),
.B(n_1818),
.Y(n_2727)
);

BUFx6f_ASAP7_75t_L g2728 ( 
.A(n_2415),
.Y(n_2728)
);

INVx3_ASAP7_75t_L g2729 ( 
.A(n_2054),
.Y(n_2729)
);

INVx1_ASAP7_75t_L g2730 ( 
.A(n_2133),
.Y(n_2730)
);

AO21x2_ASAP7_75t_L g2731 ( 
.A1(n_2065),
.A2(n_2080),
.B(n_2076),
.Y(n_2731)
);

BUFx6f_ASAP7_75t_L g2732 ( 
.A(n_2415),
.Y(n_2732)
);

NAND2xp5_ASAP7_75t_SL g2733 ( 
.A(n_2142),
.B(n_1694),
.Y(n_2733)
);

CKINVDCx5p33_ASAP7_75t_R g2734 ( 
.A(n_2345),
.Y(n_2734)
);

BUFx3_ASAP7_75t_L g2735 ( 
.A(n_2169),
.Y(n_2735)
);

CKINVDCx11_ASAP7_75t_R g2736 ( 
.A(n_2395),
.Y(n_2736)
);

BUFx2_ASAP7_75t_SL g2737 ( 
.A(n_2102),
.Y(n_2737)
);

INVx3_ASAP7_75t_SL g2738 ( 
.A(n_2106),
.Y(n_2738)
);

INVx5_ASAP7_75t_L g2739 ( 
.A(n_2102),
.Y(n_2739)
);

AOI22xp33_ASAP7_75t_L g2740 ( 
.A1(n_2405),
.A2(n_1976),
.B1(n_1767),
.B2(n_1844),
.Y(n_2740)
);

NAND2xp5_ASAP7_75t_L g2741 ( 
.A(n_2426),
.B(n_1870),
.Y(n_2741)
);

BUFx2_ASAP7_75t_L g2742 ( 
.A(n_2102),
.Y(n_2742)
);

CKINVDCx20_ASAP7_75t_R g2743 ( 
.A(n_2045),
.Y(n_2743)
);

BUFx4f_ASAP7_75t_SL g2744 ( 
.A(n_2326),
.Y(n_2744)
);

INVx1_ASAP7_75t_SL g2745 ( 
.A(n_2074),
.Y(n_2745)
);

INVx1_ASAP7_75t_SL g2746 ( 
.A(n_2086),
.Y(n_2746)
);

INVx1_ASAP7_75t_L g2747 ( 
.A(n_2133),
.Y(n_2747)
);

INVx3_ASAP7_75t_L g2748 ( 
.A(n_2054),
.Y(n_2748)
);

BUFx3_ASAP7_75t_L g2749 ( 
.A(n_2113),
.Y(n_2749)
);

BUFx3_ASAP7_75t_L g2750 ( 
.A(n_2265),
.Y(n_2750)
);

INVx8_ASAP7_75t_L g2751 ( 
.A(n_2326),
.Y(n_2751)
);

BUFx6f_ASAP7_75t_SL g2752 ( 
.A(n_2326),
.Y(n_2752)
);

BUFx6f_ASAP7_75t_L g2753 ( 
.A(n_2427),
.Y(n_2753)
);

AOI22xp33_ASAP7_75t_L g2754 ( 
.A1(n_2359),
.A2(n_2015),
.B1(n_1998),
.B2(n_2004),
.Y(n_2754)
);

AND2x2_ASAP7_75t_L g2755 ( 
.A(n_2073),
.B(n_1851),
.Y(n_2755)
);

INVx3_ASAP7_75t_L g2756 ( 
.A(n_2136),
.Y(n_2756)
);

NOR2xp33_ASAP7_75t_SL g2757 ( 
.A(n_2143),
.B(n_2030),
.Y(n_2757)
);

BUFx6f_ASAP7_75t_L g2758 ( 
.A(n_2427),
.Y(n_2758)
);

AOI22xp5_ASAP7_75t_L g2759 ( 
.A1(n_2326),
.A2(n_1866),
.B1(n_1862),
.B2(n_2004),
.Y(n_2759)
);

BUFx6f_ASAP7_75t_L g2760 ( 
.A(n_2427),
.Y(n_2760)
);

INVx1_ASAP7_75t_L g2761 ( 
.A(n_2135),
.Y(n_2761)
);

BUFx3_ASAP7_75t_L g2762 ( 
.A(n_2265),
.Y(n_2762)
);

BUFx6f_ASAP7_75t_L g2763 ( 
.A(n_2444),
.Y(n_2763)
);

BUFx6f_ASAP7_75t_L g2764 ( 
.A(n_2444),
.Y(n_2764)
);

BUFx6f_ASAP7_75t_L g2765 ( 
.A(n_2444),
.Y(n_2765)
);

BUFx3_ASAP7_75t_L g2766 ( 
.A(n_2265),
.Y(n_2766)
);

INVx3_ASAP7_75t_SL g2767 ( 
.A(n_2293),
.Y(n_2767)
);

CKINVDCx20_ASAP7_75t_R g2768 ( 
.A(n_2043),
.Y(n_2768)
);

BUFx12f_ASAP7_75t_L g2769 ( 
.A(n_2125),
.Y(n_2769)
);

INVx1_ASAP7_75t_L g2770 ( 
.A(n_2135),
.Y(n_2770)
);

BUFx2_ASAP7_75t_L g2771 ( 
.A(n_2063),
.Y(n_2771)
);

BUFx2_ASAP7_75t_L g2772 ( 
.A(n_2409),
.Y(n_2772)
);

BUFx2_ASAP7_75t_L g2773 ( 
.A(n_2214),
.Y(n_2773)
);

CKINVDCx20_ASAP7_75t_R g2774 ( 
.A(n_2349),
.Y(n_2774)
);

INVx2_ASAP7_75t_L g2775 ( 
.A(n_2341),
.Y(n_2775)
);

INVx1_ASAP7_75t_SL g2776 ( 
.A(n_2214),
.Y(n_2776)
);

BUFx3_ASAP7_75t_L g2777 ( 
.A(n_2291),
.Y(n_2777)
);

NAND2xp5_ASAP7_75t_SL g2778 ( 
.A(n_2235),
.B(n_1839),
.Y(n_2778)
);

INVx3_ASAP7_75t_SL g2779 ( 
.A(n_2293),
.Y(n_2779)
);

INVx3_ASAP7_75t_L g2780 ( 
.A(n_2136),
.Y(n_2780)
);

INVx2_ASAP7_75t_L g2781 ( 
.A(n_2353),
.Y(n_2781)
);

NAND2xp5_ASAP7_75t_L g2782 ( 
.A(n_2426),
.B(n_1921),
.Y(n_2782)
);

BUFx3_ASAP7_75t_L g2783 ( 
.A(n_2291),
.Y(n_2783)
);

INVx5_ASAP7_75t_L g2784 ( 
.A(n_2156),
.Y(n_2784)
);

INVx2_ASAP7_75t_L g2785 ( 
.A(n_2361),
.Y(n_2785)
);

CKINVDCx5p33_ASAP7_75t_R g2786 ( 
.A(n_2081),
.Y(n_2786)
);

INVx2_ASAP7_75t_SL g2787 ( 
.A(n_2202),
.Y(n_2787)
);

BUFx3_ASAP7_75t_L g2788 ( 
.A(n_2291),
.Y(n_2788)
);

CKINVDCx5p33_ASAP7_75t_R g2789 ( 
.A(n_2403),
.Y(n_2789)
);

INVx1_ASAP7_75t_L g2790 ( 
.A(n_2233),
.Y(n_2790)
);

BUFx3_ASAP7_75t_L g2791 ( 
.A(n_2305),
.Y(n_2791)
);

BUFx6f_ASAP7_75t_L g2792 ( 
.A(n_2463),
.Y(n_2792)
);

INVx1_ASAP7_75t_L g2793 ( 
.A(n_2233),
.Y(n_2793)
);

INVx1_ASAP7_75t_L g2794 ( 
.A(n_2240),
.Y(n_2794)
);

INVx4_ASAP7_75t_L g2795 ( 
.A(n_2253),
.Y(n_2795)
);

BUFx5_ASAP7_75t_L g2796 ( 
.A(n_2145),
.Y(n_2796)
);

NAND2xp5_ASAP7_75t_L g2797 ( 
.A(n_2163),
.B(n_2414),
.Y(n_2797)
);

BUFx4f_ASAP7_75t_SL g2798 ( 
.A(n_2253),
.Y(n_2798)
);

BUFx6f_ASAP7_75t_L g2799 ( 
.A(n_2463),
.Y(n_2799)
);

INVx1_ASAP7_75t_L g2800 ( 
.A(n_2240),
.Y(n_2800)
);

BUFx6f_ASAP7_75t_L g2801 ( 
.A(n_2463),
.Y(n_2801)
);

CKINVDCx16_ASAP7_75t_R g2802 ( 
.A(n_2271),
.Y(n_2802)
);

INVx2_ASAP7_75t_L g2803 ( 
.A(n_2362),
.Y(n_2803)
);

BUFx6f_ASAP7_75t_L g2804 ( 
.A(n_2146),
.Y(n_2804)
);

INVx2_ASAP7_75t_SL g2805 ( 
.A(n_2202),
.Y(n_2805)
);

CKINVDCx5p33_ASAP7_75t_R g2806 ( 
.A(n_2391),
.Y(n_2806)
);

INVx1_ASAP7_75t_SL g2807 ( 
.A(n_2212),
.Y(n_2807)
);

INVx8_ASAP7_75t_L g2808 ( 
.A(n_2305),
.Y(n_2808)
);

INVx3_ASAP7_75t_L g2809 ( 
.A(n_2217),
.Y(n_2809)
);

INVx3_ASAP7_75t_L g2810 ( 
.A(n_2217),
.Y(n_2810)
);

BUFx4f_ASAP7_75t_SL g2811 ( 
.A(n_2358),
.Y(n_2811)
);

INVx5_ASAP7_75t_L g2812 ( 
.A(n_2156),
.Y(n_2812)
);

BUFx6f_ASAP7_75t_L g2813 ( 
.A(n_2156),
.Y(n_2813)
);

INVx3_ASAP7_75t_L g2814 ( 
.A(n_2451),
.Y(n_2814)
);

INVx3_ASAP7_75t_L g2815 ( 
.A(n_2451),
.Y(n_2815)
);

INVx8_ASAP7_75t_L g2816 ( 
.A(n_2365),
.Y(n_2816)
);

INVx3_ASAP7_75t_SL g2817 ( 
.A(n_2365),
.Y(n_2817)
);

BUFx3_ASAP7_75t_L g2818 ( 
.A(n_2170),
.Y(n_2818)
);

INVx1_ASAP7_75t_SL g2819 ( 
.A(n_2149),
.Y(n_2819)
);

INVx3_ASAP7_75t_L g2820 ( 
.A(n_2294),
.Y(n_2820)
);

INVx2_ASAP7_75t_SL g2821 ( 
.A(n_2149),
.Y(n_2821)
);

INVx2_ASAP7_75t_SL g2822 ( 
.A(n_2160),
.Y(n_2822)
);

NAND2x1p5_ASAP7_75t_L g2823 ( 
.A(n_2128),
.B(n_1835),
.Y(n_2823)
);

BUFx2_ASAP7_75t_L g2824 ( 
.A(n_2358),
.Y(n_2824)
);

INVx2_ASAP7_75t_L g2825 ( 
.A(n_2183),
.Y(n_2825)
);

BUFx3_ASAP7_75t_L g2826 ( 
.A(n_2200),
.Y(n_2826)
);

CKINVDCx5p33_ASAP7_75t_R g2827 ( 
.A(n_2434),
.Y(n_2827)
);

INVx1_ASAP7_75t_SL g2828 ( 
.A(n_2736),
.Y(n_2828)
);

AOI22xp33_ASAP7_75t_SL g2829 ( 
.A1(n_2602),
.A2(n_2406),
.B1(n_2167),
.B2(n_2387),
.Y(n_2829)
);

BUFx6f_ASAP7_75t_L g2830 ( 
.A(n_2474),
.Y(n_2830)
);

NAND2xp5_ASAP7_75t_L g2831 ( 
.A(n_2503),
.B(n_2658),
.Y(n_2831)
);

INVx1_ASAP7_75t_L g2832 ( 
.A(n_2476),
.Y(n_2832)
);

INVx6_ASAP7_75t_L g2833 ( 
.A(n_2624),
.Y(n_2833)
);

OAI22xp33_ASAP7_75t_L g2834 ( 
.A1(n_2602),
.A2(n_2323),
.B1(n_2299),
.B2(n_2418),
.Y(n_2834)
);

AOI22xp33_ASAP7_75t_SL g2835 ( 
.A1(n_2581),
.A2(n_2306),
.B1(n_2310),
.B2(n_2302),
.Y(n_2835)
);

CKINVDCx20_ASAP7_75t_R g2836 ( 
.A(n_2582),
.Y(n_2836)
);

AOI22xp33_ASAP7_75t_L g2837 ( 
.A1(n_2518),
.A2(n_2329),
.B1(n_2452),
.B2(n_2155),
.Y(n_2837)
);

INVx1_ASAP7_75t_L g2838 ( 
.A(n_2504),
.Y(n_2838)
);

INVx6_ASAP7_75t_L g2839 ( 
.A(n_2631),
.Y(n_2839)
);

AOI21xp5_ASAP7_75t_L g2840 ( 
.A1(n_2733),
.A2(n_2093),
.B(n_2085),
.Y(n_2840)
);

OAI22xp5_ASAP7_75t_L g2841 ( 
.A1(n_2637),
.A2(n_2436),
.B1(n_2157),
.B2(n_2414),
.Y(n_2841)
);

CKINVDCx11_ASAP7_75t_R g2842 ( 
.A(n_2511),
.Y(n_2842)
);

INVx6_ASAP7_75t_L g2843 ( 
.A(n_2534),
.Y(n_2843)
);

INVx1_ASAP7_75t_L g2844 ( 
.A(n_2516),
.Y(n_2844)
);

AND2x2_ASAP7_75t_L g2845 ( 
.A(n_2771),
.B(n_2041),
.Y(n_2845)
);

OAI22xp5_ASAP7_75t_L g2846 ( 
.A1(n_2637),
.A2(n_2436),
.B1(n_2396),
.B2(n_2384),
.Y(n_2846)
);

AOI22xp33_ASAP7_75t_L g2847 ( 
.A1(n_2518),
.A2(n_2034),
.B1(n_2458),
.B2(n_2455),
.Y(n_2847)
);

AOI22xp33_ASAP7_75t_SL g2848 ( 
.A1(n_2581),
.A2(n_2417),
.B1(n_2342),
.B2(n_2339),
.Y(n_2848)
);

AOI22xp33_ASAP7_75t_L g2849 ( 
.A1(n_2518),
.A2(n_2388),
.B1(n_2443),
.B2(n_2429),
.Y(n_2849)
);

AOI22xp33_ASAP7_75t_L g2850 ( 
.A1(n_2581),
.A2(n_2388),
.B1(n_2443),
.B2(n_2396),
.Y(n_2850)
);

INVx4_ASAP7_75t_L g2851 ( 
.A(n_2705),
.Y(n_2851)
);

INVx1_ASAP7_75t_L g2852 ( 
.A(n_2519),
.Y(n_2852)
);

INVx1_ASAP7_75t_L g2853 ( 
.A(n_2532),
.Y(n_2853)
);

AOI21xp5_ASAP7_75t_L g2854 ( 
.A1(n_2733),
.A2(n_2093),
.B(n_2085),
.Y(n_2854)
);

OAI22xp33_ASAP7_75t_L g2855 ( 
.A1(n_2637),
.A2(n_2378),
.B1(n_2129),
.B2(n_2206),
.Y(n_2855)
);

INVx1_ASAP7_75t_SL g2856 ( 
.A(n_2554),
.Y(n_2856)
);

INVx1_ASAP7_75t_L g2857 ( 
.A(n_2549),
.Y(n_2857)
);

AOI22xp33_ASAP7_75t_L g2858 ( 
.A1(n_2584),
.A2(n_2384),
.B1(n_2036),
.B2(n_2423),
.Y(n_2858)
);

INVx1_ASAP7_75t_L g2859 ( 
.A(n_2552),
.Y(n_2859)
);

AOI22xp33_ASAP7_75t_L g2860 ( 
.A1(n_2584),
.A2(n_2423),
.B1(n_2464),
.B2(n_2449),
.Y(n_2860)
);

INVx1_ASAP7_75t_L g2861 ( 
.A(n_2553),
.Y(n_2861)
);

NAND2xp5_ASAP7_75t_L g2862 ( 
.A(n_2482),
.B(n_2413),
.Y(n_2862)
);

AOI22xp33_ASAP7_75t_L g2863 ( 
.A1(n_2594),
.A2(n_2464),
.B1(n_2465),
.B2(n_2449),
.Y(n_2863)
);

BUFx4f_ASAP7_75t_SL g2864 ( 
.A(n_2472),
.Y(n_2864)
);

NAND2xp5_ASAP7_75t_L g2865 ( 
.A(n_2482),
.B(n_2178),
.Y(n_2865)
);

NAND2xp5_ASAP7_75t_L g2866 ( 
.A(n_2509),
.B(n_2797),
.Y(n_2866)
);

INVx6_ASAP7_75t_L g2867 ( 
.A(n_2545),
.Y(n_2867)
);

INVx6_ASAP7_75t_L g2868 ( 
.A(n_2617),
.Y(n_2868)
);

INVx2_ASAP7_75t_L g2869 ( 
.A(n_2473),
.Y(n_2869)
);

OAI22xp5_ASAP7_75t_L g2870 ( 
.A1(n_2705),
.A2(n_2465),
.B1(n_2269),
.B2(n_2273),
.Y(n_2870)
);

BUFx6f_ASAP7_75t_SL g2871 ( 
.A(n_2570),
.Y(n_2871)
);

CKINVDCx5p33_ASAP7_75t_R g2872 ( 
.A(n_2557),
.Y(n_2872)
);

CKINVDCx11_ASAP7_75t_R g2873 ( 
.A(n_2485),
.Y(n_2873)
);

BUFx12f_ASAP7_75t_L g2874 ( 
.A(n_2618),
.Y(n_2874)
);

AOI22xp5_ASAP7_75t_SL g2875 ( 
.A1(n_2630),
.A2(n_2417),
.B1(n_2269),
.B2(n_2273),
.Y(n_2875)
);

INVx6_ASAP7_75t_L g2876 ( 
.A(n_2481),
.Y(n_2876)
);

OAI22xp5_ASAP7_75t_L g2877 ( 
.A1(n_2744),
.A2(n_2274),
.B1(n_2281),
.B2(n_2242),
.Y(n_2877)
);

AOI22xp33_ASAP7_75t_L g2878 ( 
.A1(n_2594),
.A2(n_2445),
.B1(n_2404),
.B2(n_2412),
.Y(n_2878)
);

CKINVDCx6p67_ASAP7_75t_R g2879 ( 
.A(n_2520),
.Y(n_2879)
);

CKINVDCx11_ASAP7_75t_R g2880 ( 
.A(n_2551),
.Y(n_2880)
);

INVx6_ASAP7_75t_L g2881 ( 
.A(n_2568),
.Y(n_2881)
);

INVx4_ASAP7_75t_L g2882 ( 
.A(n_2744),
.Y(n_2882)
);

INVx1_ASAP7_75t_L g2883 ( 
.A(n_2558),
.Y(n_2883)
);

INVxp67_ASAP7_75t_SL g2884 ( 
.A(n_2702),
.Y(n_2884)
);

CKINVDCx14_ASAP7_75t_R g2885 ( 
.A(n_2540),
.Y(n_2885)
);

INVx1_ASAP7_75t_L g2886 ( 
.A(n_2559),
.Y(n_2886)
);

INVx1_ASAP7_75t_L g2887 ( 
.A(n_2562),
.Y(n_2887)
);

BUFx6f_ASAP7_75t_L g2888 ( 
.A(n_2474),
.Y(n_2888)
);

AOI22xp33_ASAP7_75t_L g2889 ( 
.A1(n_2599),
.A2(n_2404),
.B1(n_2108),
.B2(n_2120),
.Y(n_2889)
);

OAI22xp33_ASAP7_75t_L g2890 ( 
.A1(n_2692),
.A2(n_2230),
.B1(n_2397),
.B2(n_2446),
.Y(n_2890)
);

CKINVDCx20_ASAP7_75t_R g2891 ( 
.A(n_2680),
.Y(n_2891)
);

AOI22xp33_ASAP7_75t_L g2892 ( 
.A1(n_2599),
.A2(n_2089),
.B1(n_2195),
.B2(n_2229),
.Y(n_2892)
);

AND2x2_ASAP7_75t_L g2893 ( 
.A(n_2767),
.B(n_2083),
.Y(n_2893)
);

OR2x6_ASAP7_75t_L g2894 ( 
.A(n_2808),
.B(n_2205),
.Y(n_2894)
);

INVx5_ASAP7_75t_L g2895 ( 
.A(n_2721),
.Y(n_2895)
);

AOI22xp33_ASAP7_75t_SL g2896 ( 
.A1(n_2808),
.A2(n_2274),
.B1(n_2281),
.B2(n_2242),
.Y(n_2896)
);

INVx2_ASAP7_75t_SL g2897 ( 
.A(n_2734),
.Y(n_2897)
);

INVx4_ASAP7_75t_L g2898 ( 
.A(n_2721),
.Y(n_2898)
);

INVx1_ASAP7_75t_SL g2899 ( 
.A(n_2495),
.Y(n_2899)
);

INVx2_ASAP7_75t_SL g2900 ( 
.A(n_2542),
.Y(n_2900)
);

INVx6_ASAP7_75t_L g2901 ( 
.A(n_2589),
.Y(n_2901)
);

INVx1_ASAP7_75t_L g2902 ( 
.A(n_2576),
.Y(n_2902)
);

BUFx12f_ASAP7_75t_L g2903 ( 
.A(n_2512),
.Y(n_2903)
);

AOI22xp33_ASAP7_75t_L g2904 ( 
.A1(n_2626),
.A2(n_2261),
.B1(n_2416),
.B2(n_2433),
.Y(n_2904)
);

AOI22xp33_ASAP7_75t_SL g2905 ( 
.A1(n_2808),
.A2(n_2190),
.B1(n_2227),
.B2(n_2101),
.Y(n_2905)
);

OAI22xp5_ASAP7_75t_L g2906 ( 
.A1(n_2622),
.A2(n_2174),
.B1(n_2160),
.B2(n_2383),
.Y(n_2906)
);

BUFx3_ASAP7_75t_L g2907 ( 
.A(n_2537),
.Y(n_2907)
);

INVx2_ASAP7_75t_L g2908 ( 
.A(n_2497),
.Y(n_2908)
);

CKINVDCx11_ASAP7_75t_R g2909 ( 
.A(n_2586),
.Y(n_2909)
);

AOI22xp5_ASAP7_75t_L g2910 ( 
.A1(n_2515),
.A2(n_2226),
.B1(n_2267),
.B2(n_2180),
.Y(n_2910)
);

AOI21xp5_ASAP7_75t_L g2911 ( 
.A1(n_2778),
.A2(n_2101),
.B(n_2411),
.Y(n_2911)
);

AOI22xp33_ASAP7_75t_L g2912 ( 
.A1(n_2626),
.A2(n_2174),
.B1(n_2385),
.B2(n_2199),
.Y(n_2912)
);

INVx2_ASAP7_75t_L g2913 ( 
.A(n_2501),
.Y(n_2913)
);

AOI22xp5_ASAP7_75t_SL g2914 ( 
.A1(n_2542),
.A2(n_2663),
.B1(n_2478),
.B2(n_2494),
.Y(n_2914)
);

INVx3_ASAP7_75t_L g2915 ( 
.A(n_2721),
.Y(n_2915)
);

INVx1_ASAP7_75t_L g2916 ( 
.A(n_2577),
.Y(n_2916)
);

BUFx2_ASAP7_75t_L g2917 ( 
.A(n_2546),
.Y(n_2917)
);

BUFx4f_ASAP7_75t_L g2918 ( 
.A(n_2751),
.Y(n_2918)
);

BUFx8_ASAP7_75t_L g2919 ( 
.A(n_2521),
.Y(n_2919)
);

OAI22x1_ASAP7_75t_L g2920 ( 
.A1(n_2520),
.A2(n_2084),
.B1(n_2064),
.B2(n_2373),
.Y(n_2920)
);

INVx2_ASAP7_75t_SL g2921 ( 
.A(n_2798),
.Y(n_2921)
);

OAI22xp5_ASAP7_75t_L g2922 ( 
.A1(n_2622),
.A2(n_2383),
.B1(n_2289),
.B2(n_2263),
.Y(n_2922)
);

CKINVDCx5p33_ASAP7_75t_R g2923 ( 
.A(n_2663),
.Y(n_2923)
);

AOI22xp33_ASAP7_75t_L g2924 ( 
.A1(n_2648),
.A2(n_2139),
.B1(n_2059),
.B2(n_2360),
.Y(n_2924)
);

INVx1_ASAP7_75t_L g2925 ( 
.A(n_2583),
.Y(n_2925)
);

INVx2_ASAP7_75t_L g2926 ( 
.A(n_2528),
.Y(n_2926)
);

BUFx6f_ASAP7_75t_L g2927 ( 
.A(n_2474),
.Y(n_2927)
);

HB1xp67_ASAP7_75t_L g2928 ( 
.A(n_2535),
.Y(n_2928)
);

INVx2_ASAP7_75t_L g2929 ( 
.A(n_2531),
.Y(n_2929)
);

AOI22xp33_ASAP7_75t_SL g2930 ( 
.A1(n_2816),
.A2(n_2190),
.B1(n_2227),
.B2(n_2439),
.Y(n_2930)
);

INVx2_ASAP7_75t_SL g2931 ( 
.A(n_2798),
.Y(n_2931)
);

BUFx3_ASAP7_75t_L g2932 ( 
.A(n_2563),
.Y(n_2932)
);

INVx2_ASAP7_75t_L g2933 ( 
.A(n_2533),
.Y(n_2933)
);

OR2x2_ASAP7_75t_L g2934 ( 
.A(n_2802),
.B(n_2164),
.Y(n_2934)
);

INVxp67_ASAP7_75t_SL g2935 ( 
.A(n_2702),
.Y(n_2935)
);

CKINVDCx11_ASAP7_75t_R g2936 ( 
.A(n_2572),
.Y(n_2936)
);

OAI21xp5_ASAP7_75t_SL g2937 ( 
.A1(n_2620),
.A2(n_2369),
.B(n_2367),
.Y(n_2937)
);

NAND2x1p5_ASAP7_75t_L g2938 ( 
.A(n_2688),
.B(n_2373),
.Y(n_2938)
);

INVx2_ASAP7_75t_L g2939 ( 
.A(n_2538),
.Y(n_2939)
);

INVx1_ASAP7_75t_L g2940 ( 
.A(n_2595),
.Y(n_2940)
);

NAND2x1p5_ASAP7_75t_L g2941 ( 
.A(n_2688),
.B(n_2381),
.Y(n_2941)
);

INVx2_ASAP7_75t_L g2942 ( 
.A(n_2561),
.Y(n_2942)
);

INVx1_ASAP7_75t_SL g2943 ( 
.A(n_2619),
.Y(n_2943)
);

INVxp67_ASAP7_75t_SL g2944 ( 
.A(n_2645),
.Y(n_2944)
);

CKINVDCx11_ASAP7_75t_R g2945 ( 
.A(n_2572),
.Y(n_2945)
);

INVx2_ASAP7_75t_L g2946 ( 
.A(n_2606),
.Y(n_2946)
);

AOI22xp33_ASAP7_75t_L g2947 ( 
.A1(n_2648),
.A2(n_2363),
.B1(n_2431),
.B2(n_2374),
.Y(n_2947)
);

BUFx12f_ASAP7_75t_L g2948 ( 
.A(n_2650),
.Y(n_2948)
);

AOI22xp33_ASAP7_75t_SL g2949 ( 
.A1(n_2816),
.A2(n_2439),
.B1(n_2411),
.B2(n_2381),
.Y(n_2949)
);

INVx1_ASAP7_75t_L g2950 ( 
.A(n_2598),
.Y(n_2950)
);

OAI22xp5_ASAP7_75t_L g2951 ( 
.A1(n_2622),
.A2(n_2289),
.B1(n_2263),
.B2(n_2176),
.Y(n_2951)
);

CKINVDCx6p67_ASAP7_75t_R g2952 ( 
.A(n_2678),
.Y(n_2952)
);

AOI22xp33_ASAP7_75t_L g2953 ( 
.A1(n_2699),
.A2(n_2431),
.B1(n_2374),
.B2(n_2448),
.Y(n_2953)
);

AOI22xp33_ASAP7_75t_SL g2954 ( 
.A1(n_2816),
.A2(n_2358),
.B1(n_2374),
.B2(n_2394),
.Y(n_2954)
);

INVx2_ASAP7_75t_L g2955 ( 
.A(n_2611),
.Y(n_2955)
);

INVx1_ASAP7_75t_L g2956 ( 
.A(n_2695),
.Y(n_2956)
);

INVx3_ASAP7_75t_L g2957 ( 
.A(n_2751),
.Y(n_2957)
);

INVx2_ASAP7_75t_L g2958 ( 
.A(n_2651),
.Y(n_2958)
);

BUFx3_ASAP7_75t_L g2959 ( 
.A(n_2573),
.Y(n_2959)
);

CKINVDCx11_ASAP7_75t_R g2960 ( 
.A(n_2615),
.Y(n_2960)
);

INVx3_ASAP7_75t_L g2961 ( 
.A(n_2751),
.Y(n_2961)
);

BUFx12f_ASAP7_75t_L g2962 ( 
.A(n_2683),
.Y(n_2962)
);

CKINVDCx14_ASAP7_75t_R g2963 ( 
.A(n_2827),
.Y(n_2963)
);

BUFx8_ASAP7_75t_SL g2964 ( 
.A(n_2632),
.Y(n_2964)
);

AOI22xp5_ASAP7_75t_L g2965 ( 
.A1(n_2515),
.A2(n_2377),
.B1(n_2470),
.B2(n_2254),
.Y(n_2965)
);

INVx6_ASAP7_75t_L g2966 ( 
.A(n_2795),
.Y(n_2966)
);

INVx1_ASAP7_75t_L g2967 ( 
.A(n_2695),
.Y(n_2967)
);

AOI22xp33_ASAP7_75t_L g2968 ( 
.A1(n_2699),
.A2(n_2374),
.B1(n_2201),
.B2(n_2389),
.Y(n_2968)
);

INVx2_ASAP7_75t_L g2969 ( 
.A(n_2653),
.Y(n_2969)
);

CKINVDCx20_ASAP7_75t_R g2970 ( 
.A(n_2686),
.Y(n_2970)
);

OAI22xp33_ASAP7_75t_L g2971 ( 
.A1(n_2767),
.A2(n_2466),
.B1(n_2172),
.B2(n_2377),
.Y(n_2971)
);

BUFx5_ASAP7_75t_L g2972 ( 
.A(n_2750),
.Y(n_2972)
);

BUFx8_ASAP7_75t_SL g2973 ( 
.A(n_2641),
.Y(n_2973)
);

INVx6_ASAP7_75t_L g2974 ( 
.A(n_2795),
.Y(n_2974)
);

OAI22xp5_ASAP7_75t_L g2975 ( 
.A1(n_2722),
.A2(n_2435),
.B1(n_2441),
.B2(n_2382),
.Y(n_2975)
);

INVx2_ASAP7_75t_L g2976 ( 
.A(n_2664),
.Y(n_2976)
);

INVx2_ASAP7_75t_L g2977 ( 
.A(n_2665),
.Y(n_2977)
);

AOI22xp33_ASAP7_75t_SL g2978 ( 
.A1(n_2543),
.A2(n_2358),
.B1(n_2374),
.B2(n_2410),
.Y(n_2978)
);

AOI22xp33_ASAP7_75t_L g2979 ( 
.A1(n_2546),
.A2(n_2262),
.B1(n_2366),
.B2(n_2357),
.Y(n_2979)
);

INVx1_ASAP7_75t_L g2980 ( 
.A(n_2670),
.Y(n_2980)
);

BUFx3_ASAP7_75t_L g2981 ( 
.A(n_2613),
.Y(n_2981)
);

INVx4_ASAP7_75t_L g2982 ( 
.A(n_2811),
.Y(n_2982)
);

BUFx12f_ASAP7_75t_L g2983 ( 
.A(n_2587),
.Y(n_2983)
);

NAND2xp5_ASAP7_75t_L g2984 ( 
.A(n_2509),
.B(n_2225),
.Y(n_2984)
);

NAND2x1p5_ASAP7_75t_L g2985 ( 
.A(n_2688),
.B(n_2247),
.Y(n_2985)
);

INVx2_ASAP7_75t_SL g2986 ( 
.A(n_2654),
.Y(n_2986)
);

INVx1_ASAP7_75t_L g2987 ( 
.A(n_2681),
.Y(n_2987)
);

INVx2_ASAP7_75t_L g2988 ( 
.A(n_2677),
.Y(n_2988)
);

OAI22xp5_ASAP7_75t_L g2989 ( 
.A1(n_2688),
.A2(n_2435),
.B1(n_2441),
.B2(n_2382),
.Y(n_2989)
);

AOI22xp33_ASAP7_75t_SL g2990 ( 
.A1(n_2565),
.A2(n_2425),
.B1(n_2460),
.B2(n_2096),
.Y(n_2990)
);

INVx4_ASAP7_75t_L g2991 ( 
.A(n_2811),
.Y(n_2991)
);

INVx4_ASAP7_75t_L g2992 ( 
.A(n_2506),
.Y(n_2992)
);

INVx2_ASAP7_75t_L g2993 ( 
.A(n_2684),
.Y(n_2993)
);

OAI21xp5_ASAP7_75t_L g2994 ( 
.A1(n_2483),
.A2(n_2118),
.B(n_2115),
.Y(n_2994)
);

BUFx2_ASAP7_75t_R g2995 ( 
.A(n_2698),
.Y(n_2995)
);

CKINVDCx11_ASAP7_75t_R g2996 ( 
.A(n_2605),
.Y(n_2996)
);

AOI22xp33_ASAP7_75t_L g2997 ( 
.A1(n_2659),
.A2(n_2453),
.B1(n_2469),
.B2(n_2447),
.Y(n_2997)
);

NAND2xp5_ASAP7_75t_L g2998 ( 
.A(n_2797),
.B(n_2246),
.Y(n_2998)
);

INVx1_ASAP7_75t_L g2999 ( 
.A(n_2725),
.Y(n_2999)
);

AOI22xp5_ASAP7_75t_L g3000 ( 
.A1(n_2774),
.A2(n_2355),
.B1(n_2246),
.B2(n_2400),
.Y(n_3000)
);

INVx8_ASAP7_75t_L g3001 ( 
.A(n_2752),
.Y(n_3001)
);

CKINVDCx11_ASAP7_75t_R g3002 ( 
.A(n_2779),
.Y(n_3002)
);

INVx1_ASAP7_75t_L g3003 ( 
.A(n_2725),
.Y(n_3003)
);

INVx8_ASAP7_75t_L g3004 ( 
.A(n_2752),
.Y(n_3004)
);

AOI22xp33_ASAP7_75t_L g3005 ( 
.A1(n_2659),
.A2(n_2376),
.B1(n_2398),
.B2(n_2379),
.Y(n_3005)
);

AOI22xp33_ASAP7_75t_L g3006 ( 
.A1(n_2483),
.A2(n_2379),
.B1(n_2392),
.B2(n_2400),
.Y(n_3006)
);

INVx2_ASAP7_75t_L g3007 ( 
.A(n_2687),
.Y(n_3007)
);

INVx1_ASAP7_75t_L g3008 ( 
.A(n_2505),
.Y(n_3008)
);

AOI22xp33_ASAP7_75t_L g3009 ( 
.A1(n_2612),
.A2(n_2138),
.B1(n_2241),
.B2(n_2050),
.Y(n_3009)
);

AOI22xp33_ASAP7_75t_L g3010 ( 
.A1(n_2612),
.A2(n_2571),
.B1(n_2652),
.B2(n_2600),
.Y(n_3010)
);

INVx1_ASAP7_75t_L g3011 ( 
.A(n_2693),
.Y(n_3011)
);

INVx2_ASAP7_75t_L g3012 ( 
.A(n_2713),
.Y(n_3012)
);

INVx2_ASAP7_75t_L g3013 ( 
.A(n_2724),
.Y(n_3013)
);

BUFx2_ASAP7_75t_L g3014 ( 
.A(n_2817),
.Y(n_3014)
);

AOI22xp33_ASAP7_75t_L g3015 ( 
.A1(n_2600),
.A2(n_2138),
.B1(n_2241),
.B2(n_2071),
.Y(n_3015)
);

INVx2_ASAP7_75t_SL g3016 ( 
.A(n_2654),
.Y(n_3016)
);

INVx2_ASAP7_75t_L g3017 ( 
.A(n_2775),
.Y(n_3017)
);

INVx2_ASAP7_75t_SL g3018 ( 
.A(n_2508),
.Y(n_3018)
);

BUFx2_ASAP7_75t_R g3019 ( 
.A(n_2671),
.Y(n_3019)
);

AOI21xp33_ASAP7_75t_L g3020 ( 
.A1(n_2723),
.A2(n_2457),
.B(n_2450),
.Y(n_3020)
);

AOI22xp33_ASAP7_75t_L g3021 ( 
.A1(n_2652),
.A2(n_2075),
.B1(n_2369),
.B2(n_2017),
.Y(n_3021)
);

INVx1_ASAP7_75t_L g3022 ( 
.A(n_2781),
.Y(n_3022)
);

AOI22xp33_ASAP7_75t_L g3023 ( 
.A1(n_2696),
.A2(n_2017),
.B1(n_2457),
.B2(n_2450),
.Y(n_3023)
);

BUFx8_ASAP7_75t_SL g3024 ( 
.A(n_2735),
.Y(n_3024)
);

NAND2x1p5_ASAP7_75t_L g3025 ( 
.A(n_2506),
.B(n_2247),
.Y(n_3025)
);

INVx2_ASAP7_75t_SL g3026 ( 
.A(n_2510),
.Y(n_3026)
);

OAI22x1_ASAP7_75t_L g3027 ( 
.A1(n_2620),
.A2(n_2625),
.B1(n_2696),
.B2(n_2575),
.Y(n_3027)
);

BUFx3_ASAP7_75t_L g3028 ( 
.A(n_2614),
.Y(n_3028)
);

BUFx6f_ASAP7_75t_L g3029 ( 
.A(n_2487),
.Y(n_3029)
);

AOI22xp33_ASAP7_75t_L g3030 ( 
.A1(n_2544),
.A2(n_2095),
.B1(n_2094),
.B2(n_2107),
.Y(n_3030)
);

INVx1_ASAP7_75t_L g3031 ( 
.A(n_2785),
.Y(n_3031)
);

AOI22xp33_ASAP7_75t_SL g3032 ( 
.A1(n_2625),
.A2(n_2144),
.B1(n_2188),
.B2(n_2187),
.Y(n_3032)
);

INVx2_ASAP7_75t_L g3033 ( 
.A(n_2803),
.Y(n_3033)
);

INVx1_ASAP7_75t_L g3034 ( 
.A(n_2825),
.Y(n_3034)
);

CKINVDCx20_ASAP7_75t_R g3035 ( 
.A(n_2691),
.Y(n_3035)
);

CKINVDCx5p33_ASAP7_75t_R g3036 ( 
.A(n_2717),
.Y(n_3036)
);

INVx1_ASAP7_75t_L g3037 ( 
.A(n_2535),
.Y(n_3037)
);

CKINVDCx20_ASAP7_75t_R g3038 ( 
.A(n_2691),
.Y(n_3038)
);

AOI22xp33_ASAP7_75t_L g3039 ( 
.A1(n_2668),
.A2(n_2095),
.B1(n_2094),
.B2(n_2298),
.Y(n_3039)
);

INVx1_ASAP7_75t_L g3040 ( 
.A(n_2564),
.Y(n_3040)
);

AOI22xp33_ASAP7_75t_L g3041 ( 
.A1(n_2668),
.A2(n_2333),
.B1(n_2335),
.B2(n_2298),
.Y(n_3041)
);

INVx2_ASAP7_75t_L g3042 ( 
.A(n_2505),
.Y(n_3042)
);

AOI22xp5_ASAP7_75t_SL g3043 ( 
.A1(n_2709),
.A2(n_2335),
.B1(n_2338),
.B2(n_2333),
.Y(n_3043)
);

INVx1_ASAP7_75t_L g3044 ( 
.A(n_2564),
.Y(n_3044)
);

INVx1_ASAP7_75t_L g3045 ( 
.A(n_2502),
.Y(n_3045)
);

AOI22xp33_ASAP7_75t_L g3046 ( 
.A1(n_2668),
.A2(n_2347),
.B1(n_2350),
.B2(n_2338),
.Y(n_3046)
);

INVxp67_ASAP7_75t_SL g3047 ( 
.A(n_2645),
.Y(n_3047)
);

CKINVDCx20_ASAP7_75t_R g3048 ( 
.A(n_2743),
.Y(n_3048)
);

OAI22xp5_ASAP7_75t_L g3049 ( 
.A1(n_2506),
.A2(n_2556),
.B1(n_2597),
.B2(n_2513),
.Y(n_3049)
);

INVx2_ASAP7_75t_L g3050 ( 
.A(n_2567),
.Y(n_3050)
);

AOI22xp33_ASAP7_75t_L g3051 ( 
.A1(n_2530),
.A2(n_2350),
.B1(n_2347),
.B2(n_2187),
.Y(n_3051)
);

INVx5_ASAP7_75t_L g3052 ( 
.A(n_2506),
.Y(n_3052)
);

INVx3_ASAP7_75t_L g3053 ( 
.A(n_2703),
.Y(n_3053)
);

CKINVDCx20_ASAP7_75t_R g3054 ( 
.A(n_2768),
.Y(n_3054)
);

INVx1_ASAP7_75t_L g3055 ( 
.A(n_2502),
.Y(n_3055)
);

INVx6_ASAP7_75t_L g3056 ( 
.A(n_2673),
.Y(n_3056)
);

AOI22xp33_ASAP7_75t_SL g3057 ( 
.A1(n_2737),
.A2(n_2144),
.B1(n_2188),
.B2(n_2080),
.Y(n_3057)
);

INVx2_ASAP7_75t_L g3058 ( 
.A(n_2567),
.Y(n_3058)
);

INVx1_ASAP7_75t_L g3059 ( 
.A(n_2477),
.Y(n_3059)
);

AOI22xp5_ASAP7_75t_L g3060 ( 
.A1(n_2789),
.A2(n_2806),
.B1(n_2530),
.B2(n_2479),
.Y(n_3060)
);

OAI22xp5_ASAP7_75t_L g3061 ( 
.A1(n_2513),
.A2(n_2213),
.B1(n_2219),
.B2(n_2208),
.Y(n_3061)
);

INVx1_ASAP7_75t_L g3062 ( 
.A(n_2807),
.Y(n_3062)
);

BUFx8_ASAP7_75t_L g3063 ( 
.A(n_2609),
.Y(n_3063)
);

OAI22x1_ASAP7_75t_L g3064 ( 
.A1(n_2513),
.A2(n_2319),
.B1(n_2300),
.B2(n_2277),
.Y(n_3064)
);

AOI22xp33_ASAP7_75t_L g3065 ( 
.A1(n_2703),
.A2(n_2213),
.B1(n_2219),
.B2(n_2208),
.Y(n_3065)
);

AOI22xp33_ASAP7_75t_L g3066 ( 
.A1(n_2773),
.A2(n_2121),
.B1(n_2193),
.B2(n_2184),
.Y(n_3066)
);

BUFx2_ASAP7_75t_L g3067 ( 
.A(n_2676),
.Y(n_3067)
);

BUFx2_ASAP7_75t_SL g3068 ( 
.A(n_2513),
.Y(n_3068)
);

OAI22x1_ASAP7_75t_L g3069 ( 
.A1(n_2556),
.A2(n_2597),
.B1(n_2738),
.B2(n_2742),
.Y(n_3069)
);

BUFx12f_ASAP7_75t_L g3070 ( 
.A(n_2585),
.Y(n_3070)
);

INVx1_ASAP7_75t_L g3071 ( 
.A(n_2807),
.Y(n_3071)
);

INVxp67_ASAP7_75t_SL g3072 ( 
.A(n_2475),
.Y(n_3072)
);

BUFx2_ASAP7_75t_L g3073 ( 
.A(n_2701),
.Y(n_3073)
);

INVxp67_ASAP7_75t_SL g3074 ( 
.A(n_2475),
.Y(n_3074)
);

OAI22xp33_ASAP7_75t_L g3075 ( 
.A1(n_2556),
.A2(n_2076),
.B1(n_2419),
.B2(n_2234),
.Y(n_3075)
);

BUFx4f_ASAP7_75t_SL g3076 ( 
.A(n_2647),
.Y(n_3076)
);

OAI22xp5_ASAP7_75t_L g3077 ( 
.A1(n_2556),
.A2(n_2231),
.B1(n_2234),
.B2(n_2419),
.Y(n_3077)
);

CKINVDCx11_ASAP7_75t_R g3078 ( 
.A(n_2707),
.Y(n_3078)
);

INVx2_ASAP7_75t_L g3079 ( 
.A(n_2574),
.Y(n_3079)
);

NAND2xp5_ASAP7_75t_L g3080 ( 
.A(n_2555),
.B(n_2196),
.Y(n_3080)
);

INVx6_ASAP7_75t_L g3081 ( 
.A(n_2673),
.Y(n_3081)
);

INVx1_ASAP7_75t_L g3082 ( 
.A(n_2782),
.Y(n_3082)
);

NAND2xp5_ASAP7_75t_L g3083 ( 
.A(n_2741),
.B(n_2755),
.Y(n_3083)
);

OAI22xp5_ASAP7_75t_L g3084 ( 
.A1(n_2597),
.A2(n_2231),
.B1(n_2121),
.B2(n_2294),
.Y(n_3084)
);

INVx2_ASAP7_75t_L g3085 ( 
.A(n_2574),
.Y(n_3085)
);

INVx1_ASAP7_75t_L g3086 ( 
.A(n_2782),
.Y(n_3086)
);

BUFx6f_ASAP7_75t_L g3087 ( 
.A(n_2487),
.Y(n_3087)
);

BUFx6f_ASAP7_75t_L g3088 ( 
.A(n_2487),
.Y(n_3088)
);

AND2x2_ASAP7_75t_L g3089 ( 
.A(n_2604),
.B(n_2228),
.Y(n_3089)
);

AOI22xp33_ASAP7_75t_SL g3090 ( 
.A1(n_2597),
.A2(n_2791),
.B1(n_2718),
.B2(n_2739),
.Y(n_3090)
);

AOI22xp33_ASAP7_75t_SL g3091 ( 
.A1(n_2739),
.A2(n_2006),
.B1(n_2007),
.B2(n_2011),
.Y(n_3091)
);

INVx1_ASAP7_75t_L g3092 ( 
.A(n_2480),
.Y(n_3092)
);

BUFx3_ASAP7_75t_L g3093 ( 
.A(n_2646),
.Y(n_3093)
);

INVx1_ASAP7_75t_L g3094 ( 
.A(n_2832),
.Y(n_3094)
);

NAND2xp33_ASAP7_75t_SL g3095 ( 
.A(n_2920),
.B(n_2824),
.Y(n_3095)
);

AND2x2_ASAP7_75t_L g3096 ( 
.A(n_3089),
.B(n_2604),
.Y(n_3096)
);

OAI22xp5_ASAP7_75t_L g3097 ( 
.A1(n_2905),
.A2(n_2739),
.B1(n_2819),
.B2(n_2759),
.Y(n_3097)
);

AOI22xp33_ASAP7_75t_SL g3098 ( 
.A1(n_2875),
.A2(n_2906),
.B1(n_2870),
.B2(n_2914),
.Y(n_3098)
);

NAND2xp5_ASAP7_75t_L g3099 ( 
.A(n_2956),
.B(n_2710),
.Y(n_3099)
);

NAND2xp5_ASAP7_75t_L g3100 ( 
.A(n_2967),
.B(n_2831),
.Y(n_3100)
);

AOI22xp5_ASAP7_75t_L g3101 ( 
.A1(n_2877),
.A2(n_2479),
.B1(n_2496),
.B2(n_2610),
.Y(n_3101)
);

AOI22xp33_ASAP7_75t_SL g3102 ( 
.A1(n_2922),
.A2(n_2739),
.B1(n_2585),
.B2(n_2492),
.Y(n_3102)
);

OAI22xp5_ASAP7_75t_L g3103 ( 
.A1(n_2896),
.A2(n_2819),
.B1(n_2759),
.B2(n_2776),
.Y(n_3103)
);

NAND2xp5_ASAP7_75t_L g3104 ( 
.A(n_2862),
.B(n_2710),
.Y(n_3104)
);

AND2x2_ASAP7_75t_L g3105 ( 
.A(n_2845),
.B(n_2607),
.Y(n_3105)
);

AOI22xp33_ASAP7_75t_L g3106 ( 
.A1(n_3010),
.A2(n_2547),
.B1(n_2754),
.B2(n_2769),
.Y(n_3106)
);

AND2x2_ASAP7_75t_L g3107 ( 
.A(n_2893),
.B(n_2607),
.Y(n_3107)
);

OAI21xp33_ASAP7_75t_L g3108 ( 
.A1(n_2937),
.A2(n_3060),
.B(n_3000),
.Y(n_3108)
);

NAND2xp5_ASAP7_75t_L g3109 ( 
.A(n_3083),
.B(n_2745),
.Y(n_3109)
);

NAND2xp5_ASAP7_75t_L g3110 ( 
.A(n_3059),
.B(n_2745),
.Y(n_3110)
);

AOI22xp33_ASAP7_75t_L g3111 ( 
.A1(n_2975),
.A2(n_2547),
.B1(n_2754),
.B2(n_2723),
.Y(n_3111)
);

HB1xp67_ASAP7_75t_L g3112 ( 
.A(n_2928),
.Y(n_3112)
);

AOI22xp33_ASAP7_75t_L g3113 ( 
.A1(n_2951),
.A2(n_2740),
.B1(n_2689),
.B2(n_2700),
.Y(n_3113)
);

AOI22xp33_ASAP7_75t_L g3114 ( 
.A1(n_3006),
.A2(n_2740),
.B1(n_2682),
.B2(n_2493),
.Y(n_3114)
);

INVx1_ASAP7_75t_L g3115 ( 
.A(n_2838),
.Y(n_3115)
);

OAI21xp5_ASAP7_75t_SL g3116 ( 
.A1(n_2848),
.A2(n_2490),
.B(n_2489),
.Y(n_3116)
);

OAI22xp5_ASAP7_75t_L g3117 ( 
.A1(n_2860),
.A2(n_2711),
.B1(n_2776),
.B2(n_2486),
.Y(n_3117)
);

AOI22xp33_ASAP7_75t_SL g3118 ( 
.A1(n_2846),
.A2(n_2492),
.B1(n_2486),
.B2(n_2818),
.Y(n_3118)
);

OAI22xp5_ASAP7_75t_L g3119 ( 
.A1(n_2863),
.A2(n_2486),
.B1(n_2492),
.B2(n_2821),
.Y(n_3119)
);

AND2x2_ASAP7_75t_L g3120 ( 
.A(n_3093),
.B(n_2708),
.Y(n_3120)
);

INVx2_ASAP7_75t_L g3121 ( 
.A(n_2869),
.Y(n_3121)
);

AND2x2_ASAP7_75t_L g3122 ( 
.A(n_3062),
.B(n_3071),
.Y(n_3122)
);

NAND2xp5_ASAP7_75t_L g3123 ( 
.A(n_3059),
.B(n_2746),
.Y(n_3123)
);

AND2x2_ASAP7_75t_L g3124 ( 
.A(n_3080),
.B(n_2749),
.Y(n_3124)
);

BUFx12f_ASAP7_75t_L g3125 ( 
.A(n_2909),
.Y(n_3125)
);

OAI22xp5_ASAP7_75t_L g3126 ( 
.A1(n_2930),
.A2(n_2498),
.B1(n_2486),
.B2(n_2492),
.Y(n_3126)
);

BUFx6f_ASAP7_75t_L g3127 ( 
.A(n_2966),
.Y(n_3127)
);

AOI22xp33_ASAP7_75t_SL g3128 ( 
.A1(n_3043),
.A2(n_2841),
.B1(n_3004),
.B2(n_3001),
.Y(n_3128)
);

OAI22xp5_ASAP7_75t_L g3129 ( 
.A1(n_2850),
.A2(n_2822),
.B1(n_2498),
.B2(n_2714),
.Y(n_3129)
);

AOI222xp33_ASAP7_75t_L g3130 ( 
.A1(n_2948),
.A2(n_2601),
.B1(n_2629),
.B2(n_2649),
.C1(n_2642),
.C2(n_2640),
.Y(n_3130)
);

AOI22xp5_ASAP7_75t_SL g3131 ( 
.A1(n_2891),
.A2(n_2786),
.B1(n_2826),
.B2(n_2525),
.Y(n_3131)
);

CKINVDCx11_ASAP7_75t_R g3132 ( 
.A(n_2874),
.Y(n_3132)
);

AOI22xp33_ASAP7_75t_SL g3133 ( 
.A1(n_3001),
.A2(n_3004),
.B1(n_3068),
.B2(n_2966),
.Y(n_3133)
);

OAI21xp33_ASAP7_75t_L g3134 ( 
.A1(n_2910),
.A2(n_2727),
.B(n_2610),
.Y(n_3134)
);

AOI22xp33_ASAP7_75t_SL g3135 ( 
.A1(n_2974),
.A2(n_2484),
.B1(n_2491),
.B2(n_2488),
.Y(n_3135)
);

INVx1_ASAP7_75t_L g3136 ( 
.A(n_2844),
.Y(n_3136)
);

BUFx6f_ASAP7_75t_L g3137 ( 
.A(n_2974),
.Y(n_3137)
);

INVx1_ASAP7_75t_SL g3138 ( 
.A(n_3067),
.Y(n_3138)
);

AND2x2_ASAP7_75t_L g3139 ( 
.A(n_2835),
.B(n_2772),
.Y(n_3139)
);

BUFx2_ASAP7_75t_L g3140 ( 
.A(n_3024),
.Y(n_3140)
);

OAI21xp5_ASAP7_75t_SL g3141 ( 
.A1(n_2829),
.A2(n_2490),
.B(n_2488),
.Y(n_3141)
);

OAI22xp5_ASAP7_75t_L g3142 ( 
.A1(n_2944),
.A2(n_2491),
.B1(n_2484),
.B2(n_2694),
.Y(n_3142)
);

INVx1_ASAP7_75t_L g3143 ( 
.A(n_2852),
.Y(n_3143)
);

INVx1_ASAP7_75t_L g3144 ( 
.A(n_2853),
.Y(n_3144)
);

NOR2xp33_ASAP7_75t_L g3145 ( 
.A(n_2856),
.B(n_2662),
.Y(n_3145)
);

AOI22xp33_ASAP7_75t_L g3146 ( 
.A1(n_3020),
.A2(n_2730),
.B1(n_2761),
.B2(n_2747),
.Y(n_3146)
);

INVx1_ASAP7_75t_L g3147 ( 
.A(n_2857),
.Y(n_3147)
);

OAI22xp5_ASAP7_75t_L g3148 ( 
.A1(n_3047),
.A2(n_2694),
.B1(n_2770),
.B2(n_2500),
.Y(n_3148)
);

INVx4_ASAP7_75t_L g3149 ( 
.A(n_2895),
.Y(n_3149)
);

INVx1_ASAP7_75t_L g3150 ( 
.A(n_2859),
.Y(n_3150)
);

INVx3_ASAP7_75t_L g3151 ( 
.A(n_2898),
.Y(n_3151)
);

OAI21xp5_ASAP7_75t_L g3152 ( 
.A1(n_2994),
.A2(n_2704),
.B(n_2778),
.Y(n_3152)
);

CKINVDCx5p33_ASAP7_75t_R g3153 ( 
.A(n_2885),
.Y(n_3153)
);

INVx1_ASAP7_75t_L g3154 ( 
.A(n_2861),
.Y(n_3154)
);

INVx2_ASAP7_75t_L g3155 ( 
.A(n_2908),
.Y(n_3155)
);

INVx3_ASAP7_75t_L g3156 ( 
.A(n_2898),
.Y(n_3156)
);

AOI22xp33_ASAP7_75t_L g3157 ( 
.A1(n_3039),
.A2(n_2536),
.B1(n_2657),
.B2(n_2499),
.Y(n_3157)
);

INVx2_ASAP7_75t_L g3158 ( 
.A(n_2913),
.Y(n_3158)
);

INVx1_ASAP7_75t_L g3159 ( 
.A(n_2883),
.Y(n_3159)
);

INVx2_ASAP7_75t_L g3160 ( 
.A(n_2926),
.Y(n_3160)
);

AOI22xp33_ASAP7_75t_SL g3161 ( 
.A1(n_2918),
.A2(n_2757),
.B1(n_2523),
.B2(n_2746),
.Y(n_3161)
);

HB1xp67_ASAP7_75t_L g3162 ( 
.A(n_3042),
.Y(n_3162)
);

OAI21xp5_ASAP7_75t_SL g3163 ( 
.A1(n_2963),
.A2(n_2471),
.B(n_2660),
.Y(n_3163)
);

AOI22xp33_ASAP7_75t_SL g3164 ( 
.A1(n_2918),
.A2(n_2757),
.B1(n_2679),
.B2(n_2720),
.Y(n_3164)
);

AOI22xp33_ASAP7_75t_L g3165 ( 
.A1(n_3041),
.A2(n_2704),
.B1(n_2623),
.B2(n_2741),
.Y(n_3165)
);

AND2x2_ASAP7_75t_L g3166 ( 
.A(n_2899),
.B(n_2608),
.Y(n_3166)
);

INVx3_ASAP7_75t_L g3167 ( 
.A(n_2895),
.Y(n_3167)
);

BUFx3_ASAP7_75t_L g3168 ( 
.A(n_2843),
.Y(n_3168)
);

HB1xp67_ASAP7_75t_L g3169 ( 
.A(n_2999),
.Y(n_3169)
);

AOI22xp33_ASAP7_75t_L g3170 ( 
.A1(n_3046),
.A2(n_2623),
.B1(n_2793),
.B2(n_2790),
.Y(n_3170)
);

AOI22xp33_ASAP7_75t_L g3171 ( 
.A1(n_3009),
.A2(n_2800),
.B1(n_2794),
.B2(n_2706),
.Y(n_3171)
);

AOI22xp33_ASAP7_75t_L g3172 ( 
.A1(n_3051),
.A2(n_2716),
.B1(n_2719),
.B2(n_2697),
.Y(n_3172)
);

AOI22xp33_ASAP7_75t_L g3173 ( 
.A1(n_3023),
.A2(n_2971),
.B1(n_2890),
.B2(n_2924),
.Y(n_3173)
);

OAI222xp33_ASAP7_75t_L g3174 ( 
.A1(n_2990),
.A2(n_2661),
.B1(n_2660),
.B2(n_2319),
.C1(n_2300),
.C2(n_2672),
.Y(n_3174)
);

AND2x2_ASAP7_75t_L g3175 ( 
.A(n_3073),
.B(n_2635),
.Y(n_3175)
);

INVx5_ASAP7_75t_SL g3176 ( 
.A(n_2894),
.Y(n_3176)
);

OAI21xp33_ASAP7_75t_L g3177 ( 
.A1(n_2997),
.A2(n_2675),
.B(n_2669),
.Y(n_3177)
);

AOI22xp33_ASAP7_75t_L g3178 ( 
.A1(n_2837),
.A2(n_2805),
.B1(n_2787),
.B2(n_2667),
.Y(n_3178)
);

AOI22xp33_ASAP7_75t_SL g3179 ( 
.A1(n_2986),
.A2(n_2715),
.B1(n_2720),
.B2(n_2679),
.Y(n_3179)
);

OAI22xp5_ASAP7_75t_L g3180 ( 
.A1(n_2858),
.A2(n_2661),
.B1(n_2672),
.B2(n_2655),
.Y(n_3180)
);

OAI22xp5_ASAP7_75t_L g3181 ( 
.A1(n_2949),
.A2(n_2655),
.B1(n_2627),
.B2(n_2643),
.Y(n_3181)
);

HB1xp67_ASAP7_75t_L g3182 ( 
.A(n_3003),
.Y(n_3182)
);

OAI21xp5_ASAP7_75t_SL g3183 ( 
.A1(n_3016),
.A2(n_2471),
.B(n_2715),
.Y(n_3183)
);

AOI22xp33_ASAP7_75t_L g3184 ( 
.A1(n_3015),
.A2(n_2667),
.B1(n_2593),
.B2(n_2627),
.Y(n_3184)
);

INVx2_ASAP7_75t_L g3185 ( 
.A(n_2929),
.Y(n_3185)
);

BUFx2_ASAP7_75t_L g3186 ( 
.A(n_3076),
.Y(n_3186)
);

INVx1_ASAP7_75t_L g3187 ( 
.A(n_2886),
.Y(n_3187)
);

OAI22xp5_ASAP7_75t_L g3188 ( 
.A1(n_2954),
.A2(n_2643),
.B1(n_2591),
.B2(n_2814),
.Y(n_3188)
);

INVx1_ASAP7_75t_L g3189 ( 
.A(n_2887),
.Y(n_3189)
);

BUFx8_ASAP7_75t_SL g3190 ( 
.A(n_2836),
.Y(n_3190)
);

OAI22xp5_ASAP7_75t_SL g3191 ( 
.A1(n_2923),
.A2(n_2674),
.B1(n_2636),
.B2(n_2548),
.Y(n_3191)
);

AND2x2_ASAP7_75t_L g3192 ( 
.A(n_3018),
.B(n_3026),
.Y(n_3192)
);

OAI21xp5_ASAP7_75t_SL g3193 ( 
.A1(n_2900),
.A2(n_2621),
.B(n_2616),
.Y(n_3193)
);

AND2x2_ASAP7_75t_L g3194 ( 
.A(n_2902),
.B(n_2916),
.Y(n_3194)
);

OAI22xp5_ASAP7_75t_L g3195 ( 
.A1(n_2978),
.A2(n_2591),
.B1(n_2596),
.B2(n_2579),
.Y(n_3195)
);

AND2x2_ASAP7_75t_L g3196 ( 
.A(n_2925),
.B(n_2593),
.Y(n_3196)
);

BUFx4f_ASAP7_75t_SL g3197 ( 
.A(n_2962),
.Y(n_3197)
);

INVx2_ASAP7_75t_L g3198 ( 
.A(n_2933),
.Y(n_3198)
);

INVx1_ASAP7_75t_L g3199 ( 
.A(n_2940),
.Y(n_3199)
);

INVx2_ASAP7_75t_L g3200 ( 
.A(n_2939),
.Y(n_3200)
);

INVx1_ASAP7_75t_L g3201 ( 
.A(n_2950),
.Y(n_3201)
);

NAND2xp5_ASAP7_75t_L g3202 ( 
.A(n_3092),
.B(n_2628),
.Y(n_3202)
);

INVx1_ASAP7_75t_L g3203 ( 
.A(n_2980),
.Y(n_3203)
);

OAI21xp33_ASAP7_75t_L g3204 ( 
.A1(n_2965),
.A2(n_2566),
.B(n_1765),
.Y(n_3204)
);

OAI22xp5_ASAP7_75t_L g3205 ( 
.A1(n_3045),
.A2(n_2596),
.B1(n_2579),
.B2(n_2628),
.Y(n_3205)
);

CKINVDCx5p33_ASAP7_75t_R g3206 ( 
.A(n_2873),
.Y(n_3206)
);

AOI22xp33_ASAP7_75t_L g3207 ( 
.A1(n_2855),
.A2(n_2892),
.B1(n_2912),
.B2(n_2934),
.Y(n_3207)
);

OAI22xp5_ASAP7_75t_L g3208 ( 
.A1(n_2849),
.A2(n_2815),
.B1(n_2814),
.B2(n_2810),
.Y(n_3208)
);

INVxp67_ASAP7_75t_L g3209 ( 
.A(n_3014),
.Y(n_3209)
);

AND2x2_ASAP7_75t_L g3210 ( 
.A(n_2943),
.B(n_3037),
.Y(n_3210)
);

INVx1_ASAP7_75t_L g3211 ( 
.A(n_2987),
.Y(n_3211)
);

AOI22xp33_ASAP7_75t_SL g3212 ( 
.A1(n_2895),
.A2(n_2815),
.B1(n_2666),
.B2(n_2524),
.Y(n_3212)
);

INVx1_ASAP7_75t_L g3213 ( 
.A(n_3092),
.Y(n_3213)
);

INVx1_ASAP7_75t_L g3214 ( 
.A(n_3011),
.Y(n_3214)
);

BUFx4f_ASAP7_75t_SL g3215 ( 
.A(n_3035),
.Y(n_3215)
);

OAI22xp5_ASAP7_75t_L g3216 ( 
.A1(n_3055),
.A2(n_2866),
.B1(n_3030),
.B2(n_2865),
.Y(n_3216)
);

AOI22xp33_ASAP7_75t_L g3217 ( 
.A1(n_2904),
.A2(n_2424),
.B1(n_2432),
.B2(n_2407),
.Y(n_3217)
);

AOI22xp33_ASAP7_75t_L g3218 ( 
.A1(n_3065),
.A2(n_2424),
.B1(n_2432),
.B2(n_2407),
.Y(n_3218)
);

AOI222xp33_ASAP7_75t_L g3219 ( 
.A1(n_2871),
.A2(n_2461),
.B1(n_2325),
.B2(n_2264),
.C1(n_2327),
.C2(n_2324),
.Y(n_3219)
);

NAND2xp5_ASAP7_75t_SL g3220 ( 
.A(n_3052),
.B(n_2666),
.Y(n_3220)
);

AOI22xp33_ASAP7_75t_SL g3221 ( 
.A1(n_3053),
.A2(n_2666),
.B1(n_2524),
.B2(n_2539),
.Y(n_3221)
);

BUFx2_ASAP7_75t_L g3222 ( 
.A(n_3063),
.Y(n_3222)
);

CKINVDCx5p33_ASAP7_75t_R g3223 ( 
.A(n_3038),
.Y(n_3223)
);

INVx1_ASAP7_75t_L g3224 ( 
.A(n_3022),
.Y(n_3224)
);

AOI22xp33_ASAP7_75t_L g3225 ( 
.A1(n_3005),
.A2(n_2454),
.B1(n_2007),
.B2(n_2006),
.Y(n_3225)
);

AOI222xp33_ASAP7_75t_L g3226 ( 
.A1(n_2871),
.A2(n_2318),
.B1(n_2317),
.B2(n_2290),
.C1(n_2280),
.C2(n_2278),
.Y(n_3226)
);

AND2x2_ASAP7_75t_L g3227 ( 
.A(n_3040),
.B(n_2633),
.Y(n_3227)
);

NAND2xp5_ASAP7_75t_L g3228 ( 
.A(n_3082),
.B(n_2232),
.Y(n_3228)
);

AOI22xp33_ASAP7_75t_L g3229 ( 
.A1(n_2952),
.A2(n_2454),
.B1(n_2007),
.B2(n_2006),
.Y(n_3229)
);

INVx1_ASAP7_75t_L g3230 ( 
.A(n_3031),
.Y(n_3230)
);

BUFx4f_ASAP7_75t_SL g3231 ( 
.A(n_2903),
.Y(n_3231)
);

AOI22xp33_ASAP7_75t_L g3232 ( 
.A1(n_2989),
.A2(n_2007),
.B1(n_2006),
.B2(n_2820),
.Y(n_3232)
);

AOI22xp33_ASAP7_75t_SL g3233 ( 
.A1(n_3053),
.A2(n_2666),
.B1(n_2539),
.B2(n_2550),
.Y(n_3233)
);

INVx1_ASAP7_75t_L g3234 ( 
.A(n_3034),
.Y(n_3234)
);

NAND3xp33_ASAP7_75t_L g3235 ( 
.A(n_2979),
.B(n_2311),
.C(n_1891),
.Y(n_3235)
);

AOI22xp33_ASAP7_75t_L g3236 ( 
.A1(n_2894),
.A2(n_2007),
.B1(n_2006),
.B2(n_2820),
.Y(n_3236)
);

OAI22xp33_ASAP7_75t_L g3237 ( 
.A1(n_2879),
.A2(n_2810),
.B1(n_2809),
.B2(n_2621),
.Y(n_3237)
);

INVx2_ASAP7_75t_L g3238 ( 
.A(n_2942),
.Y(n_3238)
);

INVx2_ASAP7_75t_SL g3239 ( 
.A(n_2843),
.Y(n_3239)
);

AOI22xp33_ASAP7_75t_L g3240 ( 
.A1(n_3066),
.A2(n_2007),
.B1(n_2006),
.B2(n_2731),
.Y(n_3240)
);

NAND2xp5_ASAP7_75t_L g3241 ( 
.A(n_3086),
.B(n_2244),
.Y(n_3241)
);

AOI22xp33_ASAP7_75t_SL g3242 ( 
.A1(n_3052),
.A2(n_2666),
.B1(n_2507),
.B2(n_2569),
.Y(n_3242)
);

AOI222xp33_ASAP7_75t_L g3243 ( 
.A1(n_2919),
.A2(n_2245),
.B1(n_2249),
.B2(n_2251),
.C1(n_2256),
.C2(n_2268),
.Y(n_3243)
);

OAI22xp33_ASAP7_75t_L g3244 ( 
.A1(n_2851),
.A2(n_2809),
.B1(n_2634),
.B2(n_2616),
.Y(n_3244)
);

INVx1_ASAP7_75t_SL g3245 ( 
.A(n_3069),
.Y(n_3245)
);

AOI21xp33_ASAP7_75t_L g3246 ( 
.A1(n_3064),
.A2(n_2748),
.B(n_2729),
.Y(n_3246)
);

AOI22xp33_ASAP7_75t_SL g3247 ( 
.A1(n_3052),
.A2(n_2507),
.B1(n_2569),
.B2(n_2550),
.Y(n_3247)
);

AOI22xp33_ASAP7_75t_SL g3248 ( 
.A1(n_2915),
.A2(n_2580),
.B1(n_2590),
.B2(n_2588),
.Y(n_3248)
);

OAI21xp5_ASAP7_75t_SL g3249 ( 
.A1(n_3090),
.A2(n_2634),
.B(n_2529),
.Y(n_3249)
);

INVx1_ASAP7_75t_L g3250 ( 
.A(n_3008),
.Y(n_3250)
);

AOI22xp33_ASAP7_75t_L g3251 ( 
.A1(n_2889),
.A2(n_2731),
.B1(n_2580),
.B2(n_2590),
.Y(n_3251)
);

NAND2xp5_ASAP7_75t_L g3252 ( 
.A(n_2984),
.B(n_2258),
.Y(n_3252)
);

OAI22xp5_ASAP7_75t_L g3253 ( 
.A1(n_2878),
.A2(n_2588),
.B1(n_2603),
.B2(n_2592),
.Y(n_3253)
);

INVx2_ASAP7_75t_L g3254 ( 
.A(n_2946),
.Y(n_3254)
);

AOI22xp5_ASAP7_75t_L g3255 ( 
.A1(n_2834),
.A2(n_2548),
.B1(n_2603),
.B2(n_2592),
.Y(n_3255)
);

AOI21x1_ASAP7_75t_L g3256 ( 
.A1(n_2840),
.A2(n_2051),
.B(n_2011),
.Y(n_3256)
);

INVx2_ASAP7_75t_L g3257 ( 
.A(n_2955),
.Y(n_3257)
);

AOI22xp33_ASAP7_75t_L g3258 ( 
.A1(n_2953),
.A2(n_2644),
.B1(n_2000),
.B2(n_2380),
.Y(n_3258)
);

INVx1_ASAP7_75t_L g3259 ( 
.A(n_3008),
.Y(n_3259)
);

OAI22xp5_ASAP7_75t_L g3260 ( 
.A1(n_2847),
.A2(n_2529),
.B1(n_2748),
.B2(n_2729),
.Y(n_3260)
);

INVx1_ASAP7_75t_L g3261 ( 
.A(n_2958),
.Y(n_3261)
);

HB1xp67_ASAP7_75t_L g3262 ( 
.A(n_3050),
.Y(n_3262)
);

INVx1_ASAP7_75t_L g3263 ( 
.A(n_2969),
.Y(n_3263)
);

OAI21xp33_ASAP7_75t_L g3264 ( 
.A1(n_3044),
.A2(n_1869),
.B(n_1841),
.Y(n_3264)
);

OAI222xp33_ASAP7_75t_L g3265 ( 
.A1(n_2992),
.A2(n_2756),
.B1(n_2780),
.B2(n_2823),
.C1(n_2056),
.C2(n_2784),
.Y(n_3265)
);

AOI22xp33_ASAP7_75t_L g3266 ( 
.A1(n_3027),
.A2(n_2000),
.B1(n_2401),
.B2(n_2375),
.Y(n_3266)
);

BUFx4f_ASAP7_75t_SL g3267 ( 
.A(n_2983),
.Y(n_3267)
);

AOI22xp33_ASAP7_75t_L g3268 ( 
.A1(n_3061),
.A2(n_2437),
.B1(n_1996),
.B2(n_2756),
.Y(n_3268)
);

AOI22xp33_ASAP7_75t_L g3269 ( 
.A1(n_2947),
.A2(n_1996),
.B1(n_2780),
.B2(n_1989),
.Y(n_3269)
);

OAI22xp5_ASAP7_75t_L g3270 ( 
.A1(n_2938),
.A2(n_2941),
.B1(n_2998),
.B2(n_3021),
.Y(n_3270)
);

BUFx3_ASAP7_75t_L g3271 ( 
.A(n_2932),
.Y(n_3271)
);

INVx1_ASAP7_75t_L g3272 ( 
.A(n_2976),
.Y(n_3272)
);

INVx2_ASAP7_75t_L g3273 ( 
.A(n_2977),
.Y(n_3273)
);

NAND2xp5_ASAP7_75t_L g3274 ( 
.A(n_2988),
.B(n_2993),
.Y(n_3274)
);

OAI222xp33_ASAP7_75t_L g3275 ( 
.A1(n_2992),
.A2(n_2823),
.B1(n_2812),
.B2(n_2784),
.C1(n_1704),
.C2(n_1723),
.Y(n_3275)
);

AOI22xp33_ASAP7_75t_L g3276 ( 
.A1(n_2851),
.A2(n_1996),
.B1(n_1980),
.B2(n_2527),
.Y(n_3276)
);

INVx1_ASAP7_75t_L g3277 ( 
.A(n_3007),
.Y(n_3277)
);

AOI22xp33_ASAP7_75t_SL g3278 ( 
.A1(n_2915),
.A2(n_2812),
.B1(n_2784),
.B2(n_2796),
.Y(n_3278)
);

OAI21xp33_ASAP7_75t_L g3279 ( 
.A1(n_3032),
.A2(n_2766),
.B(n_2762),
.Y(n_3279)
);

INVx2_ASAP7_75t_L g3280 ( 
.A(n_3012),
.Y(n_3280)
);

AOI22xp33_ASAP7_75t_L g3281 ( 
.A1(n_2882),
.A2(n_1996),
.B1(n_2527),
.B2(n_2008),
.Y(n_3281)
);

INVx3_ASAP7_75t_L g3282 ( 
.A(n_2982),
.Y(n_3282)
);

OAI21xp5_ASAP7_75t_SL g3283 ( 
.A1(n_2957),
.A2(n_2257),
.B(n_2255),
.Y(n_3283)
);

OAI22xp5_ASAP7_75t_SL g3284 ( 
.A1(n_2970),
.A2(n_2812),
.B1(n_2784),
.B2(n_2783),
.Y(n_3284)
);

INVx4_ASAP7_75t_L g3285 ( 
.A(n_2982),
.Y(n_3285)
);

AOI22xp33_ASAP7_75t_L g3286 ( 
.A1(n_2882),
.A2(n_2991),
.B1(n_2968),
.B2(n_2960),
.Y(n_3286)
);

AND2x2_ASAP7_75t_L g3287 ( 
.A(n_3013),
.B(n_304),
.Y(n_3287)
);

INVx1_ASAP7_75t_L g3288 ( 
.A(n_3169),
.Y(n_3288)
);

AOI22xp33_ASAP7_75t_L g3289 ( 
.A1(n_3098),
.A2(n_2991),
.B1(n_3077),
.B2(n_3084),
.Y(n_3289)
);

AOI22xp33_ASAP7_75t_L g3290 ( 
.A1(n_3130),
.A2(n_3075),
.B1(n_2917),
.B2(n_2961),
.Y(n_3290)
);

OAI21xp33_ASAP7_75t_L g3291 ( 
.A1(n_3108),
.A2(n_3057),
.B(n_2828),
.Y(n_3291)
);

AOI22xp33_ASAP7_75t_SL g3292 ( 
.A1(n_3103),
.A2(n_2961),
.B1(n_2957),
.B2(n_3049),
.Y(n_3292)
);

AOI22xp33_ASAP7_75t_SL g3293 ( 
.A1(n_3103),
.A2(n_3097),
.B1(n_3216),
.B2(n_3138),
.Y(n_3293)
);

AOI22xp33_ASAP7_75t_L g3294 ( 
.A1(n_3130),
.A2(n_2935),
.B1(n_2884),
.B2(n_2907),
.Y(n_3294)
);

INVx1_ASAP7_75t_L g3295 ( 
.A(n_3182),
.Y(n_3295)
);

NAND2xp5_ASAP7_75t_L g3296 ( 
.A(n_3194),
.B(n_3058),
.Y(n_3296)
);

INVx1_ASAP7_75t_L g3297 ( 
.A(n_3094),
.Y(n_3297)
);

AOI22xp33_ASAP7_75t_L g3298 ( 
.A1(n_3111),
.A2(n_3070),
.B1(n_2876),
.B2(n_3056),
.Y(n_3298)
);

AOI22xp33_ASAP7_75t_SL g3299 ( 
.A1(n_3097),
.A2(n_3048),
.B1(n_3054),
.B2(n_2919),
.Y(n_3299)
);

INVx1_ASAP7_75t_L g3300 ( 
.A(n_3115),
.Y(n_3300)
);

OAI22xp33_ASAP7_75t_L g3301 ( 
.A1(n_3101),
.A2(n_2931),
.B1(n_2921),
.B2(n_2833),
.Y(n_3301)
);

OAI222xp33_ASAP7_75t_L g3302 ( 
.A1(n_3128),
.A2(n_3072),
.B1(n_3074),
.B2(n_2854),
.C1(n_2911),
.C2(n_3091),
.Y(n_3302)
);

OA21x2_ASAP7_75t_L g3303 ( 
.A1(n_3276),
.A2(n_3085),
.B(n_3079),
.Y(n_3303)
);

AOI22xp33_ASAP7_75t_L g3304 ( 
.A1(n_3173),
.A2(n_2876),
.B1(n_3081),
.B2(n_3056),
.Y(n_3304)
);

OAI22xp5_ASAP7_75t_L g3305 ( 
.A1(n_3106),
.A2(n_3019),
.B1(n_3036),
.B2(n_3025),
.Y(n_3305)
);

AOI21xp5_ASAP7_75t_L g3306 ( 
.A1(n_3126),
.A2(n_1723),
.B(n_1704),
.Y(n_3306)
);

AOI22xp33_ASAP7_75t_L g3307 ( 
.A1(n_3243),
.A2(n_3081),
.B1(n_3002),
.B2(n_3063),
.Y(n_3307)
);

OAI22xp5_ASAP7_75t_L g3308 ( 
.A1(n_3165),
.A2(n_2985),
.B1(n_2833),
.B2(n_2839),
.Y(n_3308)
);

AOI22xp33_ASAP7_75t_L g3309 ( 
.A1(n_3243),
.A2(n_3134),
.B1(n_3207),
.B2(n_3216),
.Y(n_3309)
);

OAI22xp5_ASAP7_75t_L g3310 ( 
.A1(n_3118),
.A2(n_3116),
.B1(n_3178),
.B2(n_3113),
.Y(n_3310)
);

AND2x2_ASAP7_75t_L g3311 ( 
.A(n_3105),
.B(n_3017),
.Y(n_3311)
);

OAI22xp5_ASAP7_75t_L g3312 ( 
.A1(n_3157),
.A2(n_2839),
.B1(n_2868),
.B2(n_2897),
.Y(n_3312)
);

AOI22xp5_ASAP7_75t_L g3313 ( 
.A1(n_3226),
.A2(n_2868),
.B1(n_2867),
.B2(n_2901),
.Y(n_3313)
);

AOI221xp5_ASAP7_75t_L g3314 ( 
.A1(n_3146),
.A2(n_2981),
.B1(n_3028),
.B2(n_2959),
.C(n_3033),
.Y(n_3314)
);

AOI22xp33_ASAP7_75t_SL g3315 ( 
.A1(n_3148),
.A2(n_2867),
.B1(n_2864),
.B2(n_2881),
.Y(n_3315)
);

NAND2xp5_ASAP7_75t_L g3316 ( 
.A(n_3096),
.B(n_3100),
.Y(n_3316)
);

NAND3xp33_ASAP7_75t_L g3317 ( 
.A(n_3226),
.B(n_2945),
.C(n_2936),
.Y(n_3317)
);

NAND2xp5_ASAP7_75t_L g3318 ( 
.A(n_3104),
.B(n_2972),
.Y(n_3318)
);

OAI222xp33_ASAP7_75t_L g3319 ( 
.A1(n_3148),
.A2(n_2872),
.B1(n_2812),
.B2(n_1763),
.C1(n_1808),
.C2(n_2777),
.Y(n_3319)
);

AOI22xp33_ASAP7_75t_L g3320 ( 
.A1(n_3219),
.A2(n_2972),
.B1(n_2257),
.B2(n_2286),
.Y(n_3320)
);

OAI22xp5_ASAP7_75t_L g3321 ( 
.A1(n_3102),
.A2(n_2901),
.B1(n_2995),
.B2(n_2881),
.Y(n_3321)
);

AOI22xp33_ASAP7_75t_L g3322 ( 
.A1(n_3219),
.A2(n_2972),
.B1(n_2286),
.B2(n_2255),
.Y(n_3322)
);

AOI221xp5_ASAP7_75t_L g3323 ( 
.A1(n_3170),
.A2(n_1921),
.B1(n_1924),
.B2(n_2788),
.C(n_2008),
.Y(n_3323)
);

AOI22xp5_ASAP7_75t_L g3324 ( 
.A1(n_3114),
.A2(n_3078),
.B1(n_2996),
.B2(n_1808),
.Y(n_3324)
);

AND4x1_ASAP7_75t_L g3325 ( 
.A(n_3132),
.B(n_3197),
.C(n_3267),
.D(n_3231),
.Y(n_3325)
);

AOI222xp33_ASAP7_75t_L g3326 ( 
.A1(n_3222),
.A2(n_3139),
.B1(n_3177),
.B2(n_3152),
.C1(n_3109),
.C2(n_3176),
.Y(n_3326)
);

AOI22xp33_ASAP7_75t_L g3327 ( 
.A1(n_3129),
.A2(n_2972),
.B1(n_1763),
.B2(n_2191),
.Y(n_3327)
);

AOI22xp33_ASAP7_75t_L g3328 ( 
.A1(n_3152),
.A2(n_2972),
.B1(n_2185),
.B2(n_2191),
.Y(n_3328)
);

AND2x2_ASAP7_75t_L g3329 ( 
.A(n_3107),
.B(n_2830),
.Y(n_3329)
);

OAI22xp5_ASAP7_75t_L g3330 ( 
.A1(n_3184),
.A2(n_2804),
.B1(n_2221),
.B2(n_3088),
.Y(n_3330)
);

AOI22xp33_ASAP7_75t_L g3331 ( 
.A1(n_3270),
.A2(n_2185),
.B1(n_2804),
.B2(n_2796),
.Y(n_3331)
);

OAI221xp5_ASAP7_75t_SL g3332 ( 
.A1(n_3163),
.A2(n_1924),
.B1(n_2842),
.B2(n_1931),
.C(n_2973),
.Y(n_3332)
);

NAND2xp5_ASAP7_75t_L g3333 ( 
.A(n_3214),
.B(n_3088),
.Y(n_3333)
);

AOI22xp5_ASAP7_75t_L g3334 ( 
.A1(n_3270),
.A2(n_2221),
.B1(n_2796),
.B2(n_2880),
.Y(n_3334)
);

AOI22xp33_ASAP7_75t_L g3335 ( 
.A1(n_3235),
.A2(n_2804),
.B1(n_2796),
.B2(n_2296),
.Y(n_3335)
);

NAND2xp5_ASAP7_75t_SL g3336 ( 
.A(n_3127),
.B(n_2830),
.Y(n_3336)
);

AOI22xp33_ASAP7_75t_L g3337 ( 
.A1(n_3124),
.A2(n_3204),
.B1(n_3251),
.B2(n_3095),
.Y(n_3337)
);

OAI21xp33_ASAP7_75t_L g3338 ( 
.A1(n_3112),
.A2(n_1931),
.B(n_2830),
.Y(n_3338)
);

OAI222xp33_ASAP7_75t_L g3339 ( 
.A1(n_3195),
.A2(n_2296),
.B1(n_2303),
.B2(n_2964),
.C1(n_2371),
.C2(n_2386),
.Y(n_3339)
);

AOI22xp33_ASAP7_75t_L g3340 ( 
.A1(n_3126),
.A2(n_2796),
.B1(n_2296),
.B2(n_2303),
.Y(n_3340)
);

INVx2_ASAP7_75t_L g3341 ( 
.A(n_3121),
.Y(n_3341)
);

INVx1_ASAP7_75t_L g3342 ( 
.A(n_3136),
.Y(n_3342)
);

NAND2xp5_ASAP7_75t_SL g3343 ( 
.A(n_3127),
.B(n_2888),
.Y(n_3343)
);

NOR2xp33_ASAP7_75t_L g3344 ( 
.A(n_3271),
.B(n_304),
.Y(n_3344)
);

AOI22xp33_ASAP7_75t_L g3345 ( 
.A1(n_3195),
.A2(n_2303),
.B1(n_1938),
.B2(n_2295),
.Y(n_3345)
);

AOI22xp33_ASAP7_75t_L g3346 ( 
.A1(n_3188),
.A2(n_1938),
.B1(n_2295),
.B2(n_2356),
.Y(n_3346)
);

INVx4_ASAP7_75t_SL g3347 ( 
.A(n_3127),
.Y(n_3347)
);

AOI22xp33_ASAP7_75t_L g3348 ( 
.A1(n_3210),
.A2(n_3117),
.B1(n_3161),
.B2(n_3171),
.Y(n_3348)
);

AOI22xp5_ASAP7_75t_L g3349 ( 
.A1(n_3141),
.A2(n_2315),
.B1(n_2283),
.B2(n_2295),
.Y(n_3349)
);

OAI22xp5_ASAP7_75t_L g3350 ( 
.A1(n_3176),
.A2(n_2927),
.B1(n_3029),
.B2(n_2888),
.Y(n_3350)
);

AOI22xp33_ASAP7_75t_L g3351 ( 
.A1(n_3196),
.A2(n_3172),
.B1(n_3181),
.B2(n_3227),
.Y(n_3351)
);

NAND2xp5_ASAP7_75t_L g3352 ( 
.A(n_3224),
.B(n_2888),
.Y(n_3352)
);

AOI22xp33_ASAP7_75t_L g3353 ( 
.A1(n_3138),
.A2(n_3180),
.B1(n_3285),
.B2(n_3218),
.Y(n_3353)
);

AOI22xp33_ASAP7_75t_L g3354 ( 
.A1(n_3285),
.A2(n_1938),
.B1(n_2371),
.B2(n_2356),
.Y(n_3354)
);

AOI22xp33_ASAP7_75t_L g3355 ( 
.A1(n_3176),
.A2(n_2386),
.B1(n_2390),
.B2(n_2927),
.Y(n_3355)
);

AOI22xp33_ASAP7_75t_L g3356 ( 
.A1(n_3122),
.A2(n_2390),
.B1(n_3029),
.B2(n_2927),
.Y(n_3356)
);

AOI22xp33_ASAP7_75t_L g3357 ( 
.A1(n_3119),
.A2(n_3029),
.B1(n_3087),
.B2(n_3088),
.Y(n_3357)
);

NOR3xp33_ASAP7_75t_L g3358 ( 
.A(n_3209),
.B(n_2315),
.C(n_2283),
.Y(n_3358)
);

AOI22xp33_ASAP7_75t_L g3359 ( 
.A1(n_3217),
.A2(n_3087),
.B1(n_2690),
.B2(n_2712),
.Y(n_3359)
);

OAI221xp5_ASAP7_75t_SL g3360 ( 
.A1(n_3286),
.A2(n_305),
.B1(n_306),
.B2(n_307),
.C(n_309),
.Y(n_3360)
);

AOI22xp33_ASAP7_75t_L g3361 ( 
.A1(n_3287),
.A2(n_3087),
.B1(n_2690),
.B2(n_2712),
.Y(n_3361)
);

AOI22xp33_ASAP7_75t_L g3362 ( 
.A1(n_3258),
.A2(n_2690),
.B1(n_2712),
.B2(n_2685),
.Y(n_3362)
);

AND2x2_ASAP7_75t_L g3363 ( 
.A(n_3162),
.B(n_305),
.Y(n_3363)
);

AOI222xp33_ASAP7_75t_L g3364 ( 
.A1(n_3215),
.A2(n_306),
.B1(n_307),
.B2(n_309),
.C1(n_311),
.C2(n_312),
.Y(n_3364)
);

AOI22xp33_ASAP7_75t_L g3365 ( 
.A1(n_3279),
.A2(n_2726),
.B1(n_2728),
.B2(n_2685),
.Y(n_3365)
);

NAND2xp5_ASAP7_75t_L g3366 ( 
.A(n_3230),
.B(n_311),
.Y(n_3366)
);

AND2x2_ASAP7_75t_L g3367 ( 
.A(n_3120),
.B(n_312),
.Y(n_3367)
);

AOI22xp33_ASAP7_75t_SL g3368 ( 
.A1(n_3131),
.A2(n_2726),
.B1(n_2728),
.B2(n_2685),
.Y(n_3368)
);

OAI22xp5_ASAP7_75t_L g3369 ( 
.A1(n_3133),
.A2(n_2728),
.B1(n_2732),
.B2(n_2726),
.Y(n_3369)
);

OAI22xp33_ASAP7_75t_L g3370 ( 
.A1(n_3151),
.A2(n_2753),
.B1(n_2758),
.B2(n_2732),
.Y(n_3370)
);

NAND2xp33_ASAP7_75t_SL g3371 ( 
.A(n_3153),
.B(n_2732),
.Y(n_3371)
);

OR2x2_ASAP7_75t_L g3372 ( 
.A(n_3110),
.B(n_313),
.Y(n_3372)
);

OAI222xp33_ASAP7_75t_L g3373 ( 
.A1(n_3142),
.A2(n_314),
.B1(n_316),
.B2(n_317),
.C1(n_318),
.C2(n_319),
.Y(n_3373)
);

AOI22xp33_ASAP7_75t_L g3374 ( 
.A1(n_3282),
.A2(n_3164),
.B1(n_3213),
.B2(n_3250),
.Y(n_3374)
);

AOI22xp33_ASAP7_75t_L g3375 ( 
.A1(n_3282),
.A2(n_2758),
.B1(n_2760),
.B2(n_2753),
.Y(n_3375)
);

BUFx6f_ASAP7_75t_L g3376 ( 
.A(n_3137),
.Y(n_3376)
);

AOI22xp33_ASAP7_75t_L g3377 ( 
.A1(n_3259),
.A2(n_2758),
.B1(n_2760),
.B2(n_2753),
.Y(n_3377)
);

OAI21xp33_ASAP7_75t_L g3378 ( 
.A1(n_3245),
.A2(n_3123),
.B(n_3281),
.Y(n_3378)
);

AOI22xp33_ASAP7_75t_L g3379 ( 
.A1(n_3208),
.A2(n_2763),
.B1(n_2764),
.B2(n_2760),
.Y(n_3379)
);

OAI22xp5_ASAP7_75t_L g3380 ( 
.A1(n_3151),
.A2(n_2764),
.B1(n_2765),
.B2(n_2763),
.Y(n_3380)
);

AND2x2_ASAP7_75t_L g3381 ( 
.A(n_3143),
.B(n_314),
.Y(n_3381)
);

AOI22xp33_ASAP7_75t_L g3382 ( 
.A1(n_3142),
.A2(n_2764),
.B1(n_2765),
.B2(n_2763),
.Y(n_3382)
);

OAI22xp5_ASAP7_75t_L g3383 ( 
.A1(n_3156),
.A2(n_2792),
.B1(n_2799),
.B2(n_2765),
.Y(n_3383)
);

AOI22xp33_ASAP7_75t_L g3384 ( 
.A1(n_3166),
.A2(n_2799),
.B1(n_2801),
.B2(n_2792),
.Y(n_3384)
);

AND2x2_ASAP7_75t_L g3385 ( 
.A(n_3144),
.B(n_316),
.Y(n_3385)
);

AOI22xp5_ASAP7_75t_L g3386 ( 
.A1(n_3253),
.A2(n_1835),
.B1(n_2801),
.B2(n_2799),
.Y(n_3386)
);

AOI22xp33_ASAP7_75t_L g3387 ( 
.A1(n_3240),
.A2(n_2801),
.B1(n_2792),
.B2(n_1835),
.Y(n_3387)
);

AND2x2_ASAP7_75t_L g3388 ( 
.A(n_3147),
.B(n_319),
.Y(n_3388)
);

NAND2xp5_ASAP7_75t_L g3389 ( 
.A(n_3234),
.B(n_320),
.Y(n_3389)
);

AOI22xp33_ASAP7_75t_L g3390 ( 
.A1(n_3225),
.A2(n_1835),
.B1(n_2813),
.B2(n_2639),
.Y(n_3390)
);

NAND2xp5_ASAP7_75t_SL g3391 ( 
.A(n_3137),
.B(n_2514),
.Y(n_3391)
);

OAI22xp5_ASAP7_75t_L g3392 ( 
.A1(n_3156),
.A2(n_2526),
.B1(n_2656),
.B2(n_2639),
.Y(n_3392)
);

OAI222xp33_ASAP7_75t_L g3393 ( 
.A1(n_3205),
.A2(n_320),
.B1(n_321),
.B2(n_322),
.C1(n_323),
.C2(n_325),
.Y(n_3393)
);

AOI22xp33_ASAP7_75t_L g3394 ( 
.A1(n_3192),
.A2(n_2813),
.B1(n_2656),
.B2(n_2639),
.Y(n_3394)
);

NAND3xp33_ASAP7_75t_L g3395 ( 
.A(n_3266),
.B(n_2813),
.C(n_2517),
.Y(n_3395)
);

NAND3xp33_ASAP7_75t_L g3396 ( 
.A(n_3099),
.B(n_2517),
.C(n_2514),
.Y(n_3396)
);

AOI22xp33_ASAP7_75t_SL g3397 ( 
.A1(n_3149),
.A2(n_2656),
.B1(n_2638),
.B2(n_2578),
.Y(n_3397)
);

AOI22xp33_ASAP7_75t_L g3398 ( 
.A1(n_3205),
.A2(n_2638),
.B1(n_2578),
.B2(n_2560),
.Y(n_3398)
);

AND2x2_ASAP7_75t_L g3399 ( 
.A(n_3150),
.B(n_321),
.Y(n_3399)
);

AOI22xp33_ASAP7_75t_L g3400 ( 
.A1(n_3269),
.A2(n_2638),
.B1(n_2578),
.B2(n_2560),
.Y(n_3400)
);

OAI222xp33_ASAP7_75t_L g3401 ( 
.A1(n_3245),
.A2(n_323),
.B1(n_325),
.B2(n_326),
.C1(n_327),
.C2(n_329),
.Y(n_3401)
);

OAI221xp5_ASAP7_75t_L g3402 ( 
.A1(n_3193),
.A2(n_2560),
.B1(n_2541),
.B2(n_2526),
.C(n_2522),
.Y(n_3402)
);

AND2x2_ASAP7_75t_L g3403 ( 
.A(n_3154),
.B(n_327),
.Y(n_3403)
);

INVx2_ASAP7_75t_L g3404 ( 
.A(n_3155),
.Y(n_3404)
);

OAI22xp5_ASAP7_75t_L g3405 ( 
.A1(n_3248),
.A2(n_2514),
.B1(n_2526),
.B2(n_2522),
.Y(n_3405)
);

AOI22xp5_ASAP7_75t_L g3406 ( 
.A1(n_3183),
.A2(n_2541),
.B1(n_2522),
.B2(n_2517),
.Y(n_3406)
);

OAI222xp33_ASAP7_75t_L g3407 ( 
.A1(n_3135),
.A2(n_329),
.B1(n_330),
.B2(n_335),
.C1(n_336),
.C2(n_337),
.Y(n_3407)
);

AOI22xp33_ASAP7_75t_SL g3408 ( 
.A1(n_3149),
.A2(n_2541),
.B1(n_2260),
.B2(n_2252),
.Y(n_3408)
);

NAND4xp25_ASAP7_75t_L g3409 ( 
.A(n_3309),
.B(n_3145),
.C(n_3232),
.D(n_3140),
.Y(n_3409)
);

NAND2xp5_ASAP7_75t_SL g3410 ( 
.A(n_3315),
.B(n_3237),
.Y(n_3410)
);

OAI221xp5_ASAP7_75t_SL g3411 ( 
.A1(n_3307),
.A2(n_3249),
.B1(n_3186),
.B2(n_3236),
.C(n_3175),
.Y(n_3411)
);

NAND2xp5_ASAP7_75t_L g3412 ( 
.A(n_3288),
.B(n_3159),
.Y(n_3412)
);

AND2x2_ASAP7_75t_L g3413 ( 
.A(n_3329),
.B(n_3262),
.Y(n_3413)
);

NAND2xp5_ASAP7_75t_L g3414 ( 
.A(n_3295),
.B(n_3187),
.Y(n_3414)
);

NAND2xp5_ASAP7_75t_L g3415 ( 
.A(n_3316),
.B(n_3189),
.Y(n_3415)
);

NAND2xp5_ASAP7_75t_L g3416 ( 
.A(n_3311),
.B(n_3199),
.Y(n_3416)
);

AOI21xp5_ASAP7_75t_SL g3417 ( 
.A1(n_3321),
.A2(n_3220),
.B(n_3260),
.Y(n_3417)
);

OAI21xp33_ASAP7_75t_L g3418 ( 
.A1(n_3293),
.A2(n_3291),
.B(n_3292),
.Y(n_3418)
);

AND2x2_ASAP7_75t_L g3419 ( 
.A(n_3296),
.B(n_3201),
.Y(n_3419)
);

NAND2xp5_ASAP7_75t_L g3420 ( 
.A(n_3297),
.B(n_3203),
.Y(n_3420)
);

AND2x2_ASAP7_75t_L g3421 ( 
.A(n_3300),
.B(n_3211),
.Y(n_3421)
);

NAND3xp33_ASAP7_75t_L g3422 ( 
.A(n_3299),
.B(n_3246),
.C(n_3137),
.Y(n_3422)
);

AND2x2_ASAP7_75t_L g3423 ( 
.A(n_3342),
.B(n_3158),
.Y(n_3423)
);

NAND3xp33_ASAP7_75t_L g3424 ( 
.A(n_3315),
.B(n_3268),
.C(n_3263),
.Y(n_3424)
);

NAND4xp25_ASAP7_75t_L g3425 ( 
.A(n_3326),
.B(n_3255),
.C(n_3179),
.D(n_3229),
.Y(n_3425)
);

NAND2xp5_ASAP7_75t_SL g3426 ( 
.A(n_3368),
.B(n_3167),
.Y(n_3426)
);

AOI221xp5_ASAP7_75t_L g3427 ( 
.A1(n_3310),
.A2(n_3401),
.B1(n_3373),
.B2(n_3393),
.C(n_3301),
.Y(n_3427)
);

NAND3xp33_ASAP7_75t_L g3428 ( 
.A(n_3337),
.B(n_3272),
.C(n_3261),
.Y(n_3428)
);

AND2x2_ASAP7_75t_L g3429 ( 
.A(n_3341),
.B(n_3160),
.Y(n_3429)
);

OA21x2_ASAP7_75t_L g3430 ( 
.A1(n_3302),
.A2(n_3256),
.B(n_3274),
.Y(n_3430)
);

NAND3xp33_ASAP7_75t_L g3431 ( 
.A(n_3364),
.B(n_3277),
.C(n_3239),
.Y(n_3431)
);

AND2x2_ASAP7_75t_L g3432 ( 
.A(n_3404),
.B(n_3185),
.Y(n_3432)
);

NAND2xp5_ASAP7_75t_L g3433 ( 
.A(n_3318),
.B(n_3198),
.Y(n_3433)
);

NAND3xp33_ASAP7_75t_L g3434 ( 
.A(n_3317),
.B(n_3233),
.C(n_3221),
.Y(n_3434)
);

NAND2xp5_ASAP7_75t_L g3435 ( 
.A(n_3351),
.B(n_3200),
.Y(n_3435)
);

NAND3xp33_ASAP7_75t_L g3436 ( 
.A(n_3378),
.B(n_3254),
.C(n_3238),
.Y(n_3436)
);

NAND2xp5_ASAP7_75t_L g3437 ( 
.A(n_3363),
.B(n_3257),
.Y(n_3437)
);

OAI221xp5_ASAP7_75t_SL g3438 ( 
.A1(n_3294),
.A2(n_3167),
.B1(n_3283),
.B2(n_3252),
.C(n_3244),
.Y(n_3438)
);

NAND2xp5_ASAP7_75t_SL g3439 ( 
.A(n_3338),
.B(n_3242),
.Y(n_3439)
);

AND2x2_ASAP7_75t_L g3440 ( 
.A(n_3367),
.B(n_3273),
.Y(n_3440)
);

AND2x2_ASAP7_75t_L g3441 ( 
.A(n_3353),
.B(n_3280),
.Y(n_3441)
);

NOR2xp33_ASAP7_75t_R g3442 ( 
.A(n_3371),
.B(n_3125),
.Y(n_3442)
);

AND2x2_ASAP7_75t_L g3443 ( 
.A(n_3333),
.B(n_3168),
.Y(n_3443)
);

OAI21xp5_ASAP7_75t_SL g3444 ( 
.A1(n_3313),
.A2(n_3174),
.B(n_3212),
.Y(n_3444)
);

AND2x2_ASAP7_75t_L g3445 ( 
.A(n_3352),
.B(n_3202),
.Y(n_3445)
);

NAND2xp5_ASAP7_75t_SL g3446 ( 
.A(n_3334),
.B(n_3247),
.Y(n_3446)
);

NAND3xp33_ASAP7_75t_L g3447 ( 
.A(n_3314),
.B(n_3278),
.C(n_3241),
.Y(n_3447)
);

OAI22xp5_ASAP7_75t_L g3448 ( 
.A1(n_3332),
.A2(n_3284),
.B1(n_3228),
.B2(n_3223),
.Y(n_3448)
);

NAND2xp5_ASAP7_75t_L g3449 ( 
.A(n_3381),
.B(n_3264),
.Y(n_3449)
);

NAND2xp5_ASAP7_75t_L g3450 ( 
.A(n_3385),
.B(n_330),
.Y(n_3450)
);

NAND2xp5_ASAP7_75t_L g3451 ( 
.A(n_3388),
.B(n_335),
.Y(n_3451)
);

OAI21xp5_ASAP7_75t_SL g3452 ( 
.A1(n_3401),
.A2(n_3265),
.B(n_3275),
.Y(n_3452)
);

NAND4xp25_ASAP7_75t_L g3453 ( 
.A(n_3290),
.B(n_336),
.C(n_337),
.D(n_338),
.Y(n_3453)
);

NAND2xp5_ASAP7_75t_L g3454 ( 
.A(n_3399),
.B(n_340),
.Y(n_3454)
);

AOI22xp33_ASAP7_75t_L g3455 ( 
.A1(n_3305),
.A2(n_3191),
.B1(n_3190),
.B2(n_3206),
.Y(n_3455)
);

AND2x2_ASAP7_75t_L g3456 ( 
.A(n_3348),
.B(n_341),
.Y(n_3456)
);

NAND2xp5_ASAP7_75t_L g3457 ( 
.A(n_3403),
.B(n_341),
.Y(n_3457)
);

AND2x2_ASAP7_75t_L g3458 ( 
.A(n_3376),
.B(n_342),
.Y(n_3458)
);

NOR2xp67_ASAP7_75t_L g3459 ( 
.A(n_3369),
.B(n_342),
.Y(n_3459)
);

NAND4xp25_ASAP7_75t_L g3460 ( 
.A(n_3289),
.B(n_343),
.C(n_344),
.D(n_345),
.Y(n_3460)
);

OAI22xp5_ASAP7_75t_L g3461 ( 
.A1(n_3320),
.A2(n_2260),
.B1(n_2252),
.B2(n_2181),
.Y(n_3461)
);

AND2x2_ASAP7_75t_L g3462 ( 
.A(n_3376),
.B(n_343),
.Y(n_3462)
);

NOR2xp67_ASAP7_75t_L g3463 ( 
.A(n_3312),
.B(n_344),
.Y(n_3463)
);

AND2x2_ASAP7_75t_L g3464 ( 
.A(n_3376),
.B(n_345),
.Y(n_3464)
);

NAND3xp33_ASAP7_75t_L g3465 ( 
.A(n_3344),
.B(n_2252),
.C(n_2181),
.Y(n_3465)
);

NAND4xp25_ASAP7_75t_L g3466 ( 
.A(n_3298),
.B(n_346),
.C(n_347),
.D(n_348),
.Y(n_3466)
);

NOR3xp33_ASAP7_75t_L g3467 ( 
.A(n_3407),
.B(n_347),
.C(n_348),
.Y(n_3467)
);

OAI221xp5_ASAP7_75t_L g3468 ( 
.A1(n_3304),
.A2(n_349),
.B1(n_350),
.B2(n_351),
.C(n_352),
.Y(n_3468)
);

NOR3xp33_ASAP7_75t_L g3469 ( 
.A(n_3407),
.B(n_349),
.C(n_350),
.Y(n_3469)
);

AND2x2_ASAP7_75t_L g3470 ( 
.A(n_3356),
.B(n_352),
.Y(n_3470)
);

AND2x2_ASAP7_75t_L g3471 ( 
.A(n_3413),
.B(n_3382),
.Y(n_3471)
);

AOI22xp5_ASAP7_75t_L g3472 ( 
.A1(n_3418),
.A2(n_3308),
.B1(n_3324),
.B2(n_3374),
.Y(n_3472)
);

NAND2xp5_ASAP7_75t_L g3473 ( 
.A(n_3441),
.B(n_3372),
.Y(n_3473)
);

NAND2xp5_ASAP7_75t_L g3474 ( 
.A(n_3419),
.B(n_3331),
.Y(n_3474)
);

NAND2xp5_ASAP7_75t_L g3475 ( 
.A(n_3421),
.B(n_3303),
.Y(n_3475)
);

NOR2x1_ASAP7_75t_L g3476 ( 
.A(n_3417),
.B(n_3339),
.Y(n_3476)
);

AND2x2_ASAP7_75t_L g3477 ( 
.A(n_3443),
.B(n_3398),
.Y(n_3477)
);

NAND3xp33_ASAP7_75t_L g3478 ( 
.A(n_3427),
.B(n_3360),
.C(n_3366),
.Y(n_3478)
);

AND2x2_ASAP7_75t_SL g3479 ( 
.A(n_3455),
.B(n_3325),
.Y(n_3479)
);

OAI21xp5_ASAP7_75t_L g3480 ( 
.A1(n_3467),
.A2(n_3469),
.B(n_3452),
.Y(n_3480)
);

NAND2xp5_ASAP7_75t_L g3481 ( 
.A(n_3445),
.B(n_3389),
.Y(n_3481)
);

AND2x2_ASAP7_75t_L g3482 ( 
.A(n_3440),
.B(n_3303),
.Y(n_3482)
);

BUFx3_ASAP7_75t_L g3483 ( 
.A(n_3429),
.Y(n_3483)
);

OR2x2_ASAP7_75t_L g3484 ( 
.A(n_3416),
.B(n_3396),
.Y(n_3484)
);

OAI21xp5_ASAP7_75t_L g3485 ( 
.A1(n_3467),
.A2(n_3393),
.B(n_3373),
.Y(n_3485)
);

INVx1_ASAP7_75t_L g3486 ( 
.A(n_3420),
.Y(n_3486)
);

NAND2xp5_ASAP7_75t_L g3487 ( 
.A(n_3449),
.B(n_3345),
.Y(n_3487)
);

AO21x2_ASAP7_75t_L g3488 ( 
.A1(n_3428),
.A2(n_3302),
.B(n_3306),
.Y(n_3488)
);

OR2x2_ASAP7_75t_L g3489 ( 
.A(n_3412),
.B(n_3395),
.Y(n_3489)
);

NAND4xp75_ASAP7_75t_L g3490 ( 
.A(n_3410),
.B(n_3406),
.C(n_3336),
.D(n_3343),
.Y(n_3490)
);

AND2x2_ASAP7_75t_L g3491 ( 
.A(n_3423),
.B(n_3379),
.Y(n_3491)
);

AND2x2_ASAP7_75t_L g3492 ( 
.A(n_3432),
.B(n_3357),
.Y(n_3492)
);

NOR3xp33_ASAP7_75t_L g3493 ( 
.A(n_3411),
.B(n_3339),
.C(n_3319),
.Y(n_3493)
);

NOR3xp33_ASAP7_75t_L g3494 ( 
.A(n_3411),
.B(n_3319),
.C(n_3330),
.Y(n_3494)
);

AND2x2_ASAP7_75t_L g3495 ( 
.A(n_3415),
.B(n_3365),
.Y(n_3495)
);

NAND2xp5_ASAP7_75t_L g3496 ( 
.A(n_3435),
.B(n_3346),
.Y(n_3496)
);

NAND2xp5_ASAP7_75t_L g3497 ( 
.A(n_3414),
.B(n_3384),
.Y(n_3497)
);

OR2x2_ASAP7_75t_L g3498 ( 
.A(n_3433),
.B(n_3405),
.Y(n_3498)
);

OAI221xp5_ASAP7_75t_L g3499 ( 
.A1(n_3444),
.A2(n_3322),
.B1(n_3340),
.B2(n_3335),
.C(n_3394),
.Y(n_3499)
);

NOR2xp33_ASAP7_75t_L g3500 ( 
.A(n_3409),
.B(n_3347),
.Y(n_3500)
);

AND2x2_ASAP7_75t_L g3501 ( 
.A(n_3437),
.B(n_3386),
.Y(n_3501)
);

OAI21xp5_ASAP7_75t_L g3502 ( 
.A1(n_3469),
.A2(n_3402),
.B(n_3350),
.Y(n_3502)
);

NAND2xp5_ASAP7_75t_L g3503 ( 
.A(n_3436),
.B(n_3377),
.Y(n_3503)
);

OAI211xp5_ASAP7_75t_L g3504 ( 
.A1(n_3410),
.A2(n_3397),
.B(n_3362),
.C(n_3361),
.Y(n_3504)
);

NOR3xp33_ASAP7_75t_L g3505 ( 
.A(n_3438),
.B(n_3358),
.C(n_3323),
.Y(n_3505)
);

NOR3xp33_ASAP7_75t_SL g3506 ( 
.A(n_3438),
.B(n_3370),
.C(n_3380),
.Y(n_3506)
);

AOI22xp33_ASAP7_75t_L g3507 ( 
.A1(n_3425),
.A2(n_3328),
.B1(n_3400),
.B2(n_3359),
.Y(n_3507)
);

OR2x2_ASAP7_75t_L g3508 ( 
.A(n_3426),
.B(n_3383),
.Y(n_3508)
);

AOI22xp5_ASAP7_75t_L g3509 ( 
.A1(n_3448),
.A2(n_3327),
.B1(n_3347),
.B2(n_3349),
.Y(n_3509)
);

AND2x2_ASAP7_75t_L g3510 ( 
.A(n_3455),
.B(n_3458),
.Y(n_3510)
);

OAI211xp5_ASAP7_75t_L g3511 ( 
.A1(n_3442),
.A2(n_3375),
.B(n_3355),
.C(n_3408),
.Y(n_3511)
);

AND2x2_ASAP7_75t_L g3512 ( 
.A(n_3462),
.B(n_3347),
.Y(n_3512)
);

NAND3xp33_ASAP7_75t_L g3513 ( 
.A(n_3431),
.B(n_3354),
.C(n_3392),
.Y(n_3513)
);

BUFx2_ASAP7_75t_L g3514 ( 
.A(n_3442),
.Y(n_3514)
);

AOI22xp5_ASAP7_75t_L g3515 ( 
.A1(n_3460),
.A2(n_3391),
.B1(n_3387),
.B2(n_3390),
.Y(n_3515)
);

AOI22xp33_ASAP7_75t_SL g3516 ( 
.A1(n_3434),
.A2(n_2260),
.B1(n_2181),
.B2(n_356),
.Y(n_3516)
);

AO21x2_ASAP7_75t_L g3517 ( 
.A1(n_3446),
.A2(n_353),
.B(n_355),
.Y(n_3517)
);

OR2x6_ASAP7_75t_L g3518 ( 
.A(n_3459),
.B(n_353),
.Y(n_3518)
);

INVx1_ASAP7_75t_SL g3519 ( 
.A(n_3514),
.Y(n_3519)
);

XNOR2xp5_ASAP7_75t_L g3520 ( 
.A(n_3479),
.B(n_3422),
.Y(n_3520)
);

INVx1_ASAP7_75t_L g3521 ( 
.A(n_3486),
.Y(n_3521)
);

NAND4xp75_ASAP7_75t_SL g3522 ( 
.A(n_3500),
.B(n_3463),
.C(n_3430),
.D(n_3456),
.Y(n_3522)
);

HB1xp67_ASAP7_75t_L g3523 ( 
.A(n_3483),
.Y(n_3523)
);

XNOR2xp5_ASAP7_75t_L g3524 ( 
.A(n_3510),
.B(n_3466),
.Y(n_3524)
);

XNOR2xp5_ASAP7_75t_L g3525 ( 
.A(n_3476),
.B(n_3447),
.Y(n_3525)
);

INVx1_ASAP7_75t_L g3526 ( 
.A(n_3484),
.Y(n_3526)
);

NOR4xp25_ASAP7_75t_L g3527 ( 
.A(n_3480),
.B(n_3453),
.C(n_3468),
.D(n_3450),
.Y(n_3527)
);

XOR2x2_ASAP7_75t_L g3528 ( 
.A(n_3472),
.B(n_3480),
.Y(n_3528)
);

INVx1_ASAP7_75t_L g3529 ( 
.A(n_3489),
.Y(n_3529)
);

NAND4xp75_ASAP7_75t_L g3530 ( 
.A(n_3506),
.B(n_3446),
.C(n_3439),
.D(n_3464),
.Y(n_3530)
);

AND2x2_ASAP7_75t_L g3531 ( 
.A(n_3482),
.B(n_3430),
.Y(n_3531)
);

NAND2xp5_ASAP7_75t_L g3532 ( 
.A(n_3495),
.B(n_3439),
.Y(n_3532)
);

INVx2_ASAP7_75t_SL g3533 ( 
.A(n_3512),
.Y(n_3533)
);

INVx2_ASAP7_75t_SL g3534 ( 
.A(n_3492),
.Y(n_3534)
);

INVx1_ASAP7_75t_L g3535 ( 
.A(n_3475),
.Y(n_3535)
);

NAND2xp5_ASAP7_75t_L g3536 ( 
.A(n_3487),
.B(n_3424),
.Y(n_3536)
);

INVx1_ASAP7_75t_L g3537 ( 
.A(n_3475),
.Y(n_3537)
);

INVx1_ASAP7_75t_L g3538 ( 
.A(n_3497),
.Y(n_3538)
);

NOR2x1_ASAP7_75t_L g3539 ( 
.A(n_3490),
.B(n_3513),
.Y(n_3539)
);

INVx2_ASAP7_75t_SL g3540 ( 
.A(n_3508),
.Y(n_3540)
);

AOI22xp5_ASAP7_75t_L g3541 ( 
.A1(n_3478),
.A2(n_3457),
.B1(n_3454),
.B2(n_3451),
.Y(n_3541)
);

INVx1_ASAP7_75t_L g3542 ( 
.A(n_3498),
.Y(n_3542)
);

HB1xp67_ASAP7_75t_L g3543 ( 
.A(n_3491),
.Y(n_3543)
);

INVx1_ASAP7_75t_L g3544 ( 
.A(n_3481),
.Y(n_3544)
);

XOR2x2_ASAP7_75t_L g3545 ( 
.A(n_3478),
.B(n_3465),
.Y(n_3545)
);

OAI31xp33_ASAP7_75t_L g3546 ( 
.A1(n_3493),
.A2(n_3470),
.A3(n_3461),
.B(n_358),
.Y(n_3546)
);

AND2x2_ASAP7_75t_L g3547 ( 
.A(n_3471),
.B(n_356),
.Y(n_3547)
);

INVx1_ASAP7_75t_L g3548 ( 
.A(n_3474),
.Y(n_3548)
);

AND2x2_ASAP7_75t_L g3549 ( 
.A(n_3477),
.B(n_357),
.Y(n_3549)
);

AOI22xp5_ASAP7_75t_L g3550 ( 
.A1(n_3505),
.A2(n_3485),
.B1(n_3494),
.B2(n_3518),
.Y(n_3550)
);

XNOR2x2_ASAP7_75t_L g3551 ( 
.A(n_3513),
.B(n_357),
.Y(n_3551)
);

AND2x4_ASAP7_75t_L g3552 ( 
.A(n_3501),
.B(n_358),
.Y(n_3552)
);

INVx1_ASAP7_75t_L g3553 ( 
.A(n_3473),
.Y(n_3553)
);

XOR2xp5_ASAP7_75t_L g3554 ( 
.A(n_3509),
.B(n_3496),
.Y(n_3554)
);

OR2x2_ASAP7_75t_L g3555 ( 
.A(n_3503),
.B(n_359),
.Y(n_3555)
);

INVx2_ASAP7_75t_L g3556 ( 
.A(n_3488),
.Y(n_3556)
);

AND2x4_ASAP7_75t_L g3557 ( 
.A(n_3488),
.B(n_360),
.Y(n_3557)
);

XNOR2xp5_ASAP7_75t_L g3558 ( 
.A(n_3507),
.B(n_361),
.Y(n_3558)
);

NAND4xp75_ASAP7_75t_L g3559 ( 
.A(n_3485),
.B(n_362),
.C(n_363),
.D(n_364),
.Y(n_3559)
);

AND2x2_ASAP7_75t_L g3560 ( 
.A(n_3502),
.B(n_362),
.Y(n_3560)
);

NAND2xp5_ASAP7_75t_L g3561 ( 
.A(n_3517),
.B(n_364),
.Y(n_3561)
);

XOR2x2_ASAP7_75t_L g3562 ( 
.A(n_3528),
.B(n_3520),
.Y(n_3562)
);

INVx2_ASAP7_75t_SL g3563 ( 
.A(n_3523),
.Y(n_3563)
);

XNOR2xp5_ASAP7_75t_L g3564 ( 
.A(n_3530),
.B(n_3504),
.Y(n_3564)
);

INVx1_ASAP7_75t_L g3565 ( 
.A(n_3526),
.Y(n_3565)
);

INVx1_ASAP7_75t_L g3566 ( 
.A(n_3542),
.Y(n_3566)
);

XOR2x2_ASAP7_75t_L g3567 ( 
.A(n_3550),
.B(n_3499),
.Y(n_3567)
);

INVx1_ASAP7_75t_L g3568 ( 
.A(n_3529),
.Y(n_3568)
);

XOR2x2_ASAP7_75t_L g3569 ( 
.A(n_3550),
.B(n_3502),
.Y(n_3569)
);

INVx1_ASAP7_75t_L g3570 ( 
.A(n_3521),
.Y(n_3570)
);

INVxp67_ASAP7_75t_L g3571 ( 
.A(n_3519),
.Y(n_3571)
);

HB1xp67_ASAP7_75t_L g3572 ( 
.A(n_3519),
.Y(n_3572)
);

INVxp67_ASAP7_75t_L g3573 ( 
.A(n_3560),
.Y(n_3573)
);

INVx2_ASAP7_75t_L g3574 ( 
.A(n_3540),
.Y(n_3574)
);

INVx1_ASAP7_75t_SL g3575 ( 
.A(n_3552),
.Y(n_3575)
);

INVxp67_ASAP7_75t_L g3576 ( 
.A(n_3556),
.Y(n_3576)
);

INVx1_ASAP7_75t_L g3577 ( 
.A(n_3538),
.Y(n_3577)
);

INVx1_ASAP7_75t_L g3578 ( 
.A(n_3535),
.Y(n_3578)
);

OAI22x1_ASAP7_75t_L g3579 ( 
.A1(n_3525),
.A2(n_3515),
.B1(n_3518),
.B2(n_3511),
.Y(n_3579)
);

INVx1_ASAP7_75t_L g3580 ( 
.A(n_3537),
.Y(n_3580)
);

INVx1_ASAP7_75t_L g3581 ( 
.A(n_3548),
.Y(n_3581)
);

NAND2xp5_ASAP7_75t_L g3582 ( 
.A(n_3543),
.B(n_3517),
.Y(n_3582)
);

INVx1_ASAP7_75t_L g3583 ( 
.A(n_3544),
.Y(n_3583)
);

INVx2_ASAP7_75t_L g3584 ( 
.A(n_3534),
.Y(n_3584)
);

XNOR2xp5_ASAP7_75t_L g3585 ( 
.A(n_3558),
.B(n_3554),
.Y(n_3585)
);

XNOR2xp5_ASAP7_75t_L g3586 ( 
.A(n_3524),
.B(n_3516),
.Y(n_3586)
);

NOR2xp33_ASAP7_75t_L g3587 ( 
.A(n_3536),
.B(n_3518),
.Y(n_3587)
);

INVxp67_ASAP7_75t_L g3588 ( 
.A(n_3539),
.Y(n_3588)
);

INVx1_ASAP7_75t_SL g3589 ( 
.A(n_3552),
.Y(n_3589)
);

AOI22xp5_ASAP7_75t_L g3590 ( 
.A1(n_3579),
.A2(n_3545),
.B1(n_3557),
.B2(n_3532),
.Y(n_3590)
);

OA22x2_ASAP7_75t_L g3591 ( 
.A1(n_3588),
.A2(n_3557),
.B1(n_3541),
.B2(n_3531),
.Y(n_3591)
);

INVx1_ASAP7_75t_L g3592 ( 
.A(n_3572),
.Y(n_3592)
);

INVx1_ASAP7_75t_L g3593 ( 
.A(n_3578),
.Y(n_3593)
);

INVx2_ASAP7_75t_L g3594 ( 
.A(n_3563),
.Y(n_3594)
);

INVx1_ASAP7_75t_L g3595 ( 
.A(n_3571),
.Y(n_3595)
);

INVx1_ASAP7_75t_L g3596 ( 
.A(n_3583),
.Y(n_3596)
);

XOR2x2_ASAP7_75t_L g3597 ( 
.A(n_3562),
.B(n_3569),
.Y(n_3597)
);

OAI22xp5_ASAP7_75t_L g3598 ( 
.A1(n_3575),
.A2(n_3533),
.B1(n_3553),
.B2(n_3541),
.Y(n_3598)
);

INVx2_ASAP7_75t_L g3599 ( 
.A(n_3574),
.Y(n_3599)
);

INVx1_ASAP7_75t_L g3600 ( 
.A(n_3577),
.Y(n_3600)
);

INVx2_ASAP7_75t_L g3601 ( 
.A(n_3584),
.Y(n_3601)
);

INVx1_ASAP7_75t_L g3602 ( 
.A(n_3580),
.Y(n_3602)
);

XOR2x2_ASAP7_75t_L g3603 ( 
.A(n_3567),
.B(n_3551),
.Y(n_3603)
);

OA22x2_ASAP7_75t_L g3604 ( 
.A1(n_3564),
.A2(n_3549),
.B1(n_3547),
.B2(n_3561),
.Y(n_3604)
);

INVxp33_ASAP7_75t_SL g3605 ( 
.A(n_3585),
.Y(n_3605)
);

INVx2_ASAP7_75t_SL g3606 ( 
.A(n_3575),
.Y(n_3606)
);

INVx1_ASAP7_75t_L g3607 ( 
.A(n_3570),
.Y(n_3607)
);

INVx2_ASAP7_75t_SL g3608 ( 
.A(n_3589),
.Y(n_3608)
);

BUFx3_ASAP7_75t_L g3609 ( 
.A(n_3589),
.Y(n_3609)
);

INVx1_ASAP7_75t_L g3610 ( 
.A(n_3566),
.Y(n_3610)
);

OA22x2_ASAP7_75t_L g3611 ( 
.A1(n_3586),
.A2(n_3561),
.B1(n_3522),
.B2(n_3546),
.Y(n_3611)
);

XNOR2x1_ASAP7_75t_L g3612 ( 
.A(n_3565),
.B(n_3559),
.Y(n_3612)
);

OAI22xp5_ASAP7_75t_L g3613 ( 
.A1(n_3573),
.A2(n_3555),
.B1(n_3546),
.B2(n_3527),
.Y(n_3613)
);

INVx1_ASAP7_75t_SL g3614 ( 
.A(n_3582),
.Y(n_3614)
);

OAI22xp5_ASAP7_75t_L g3615 ( 
.A1(n_3573),
.A2(n_3527),
.B1(n_1799),
.B2(n_369),
.Y(n_3615)
);

OAI22xp5_ASAP7_75t_L g3616 ( 
.A1(n_3587),
.A2(n_1799),
.B1(n_367),
.B2(n_369),
.Y(n_3616)
);

OA22x2_ASAP7_75t_L g3617 ( 
.A1(n_3582),
.A2(n_365),
.B1(n_367),
.B2(n_371),
.Y(n_3617)
);

OA22x2_ASAP7_75t_L g3618 ( 
.A1(n_3568),
.A2(n_365),
.B1(n_371),
.B2(n_373),
.Y(n_3618)
);

INVx1_ASAP7_75t_L g3619 ( 
.A(n_3592),
.Y(n_3619)
);

INVxp67_ASAP7_75t_L g3620 ( 
.A(n_3609),
.Y(n_3620)
);

INVx3_ASAP7_75t_L g3621 ( 
.A(n_3594),
.Y(n_3621)
);

INVx1_ASAP7_75t_L g3622 ( 
.A(n_3592),
.Y(n_3622)
);

INVx2_ASAP7_75t_L g3623 ( 
.A(n_3606),
.Y(n_3623)
);

INVx2_ASAP7_75t_L g3624 ( 
.A(n_3608),
.Y(n_3624)
);

INVx1_ASAP7_75t_L g3625 ( 
.A(n_3595),
.Y(n_3625)
);

INVx1_ASAP7_75t_L g3626 ( 
.A(n_3593),
.Y(n_3626)
);

INVx1_ASAP7_75t_L g3627 ( 
.A(n_3593),
.Y(n_3627)
);

INVx2_ASAP7_75t_L g3628 ( 
.A(n_3599),
.Y(n_3628)
);

INVx1_ASAP7_75t_L g3629 ( 
.A(n_3602),
.Y(n_3629)
);

HB1xp67_ASAP7_75t_L g3630 ( 
.A(n_3614),
.Y(n_3630)
);

INVx2_ASAP7_75t_L g3631 ( 
.A(n_3601),
.Y(n_3631)
);

INVx1_ASAP7_75t_L g3632 ( 
.A(n_3602),
.Y(n_3632)
);

INVx1_ASAP7_75t_L g3633 ( 
.A(n_3596),
.Y(n_3633)
);

INVx1_ASAP7_75t_L g3634 ( 
.A(n_3600),
.Y(n_3634)
);

INVx1_ASAP7_75t_L g3635 ( 
.A(n_3607),
.Y(n_3635)
);

OAI322xp33_ASAP7_75t_L g3636 ( 
.A1(n_3590),
.A2(n_3613),
.A3(n_3591),
.B1(n_3611),
.B2(n_3604),
.C1(n_3598),
.C2(n_3615),
.Y(n_3636)
);

INVx1_ASAP7_75t_L g3637 ( 
.A(n_3607),
.Y(n_3637)
);

INVx2_ASAP7_75t_L g3638 ( 
.A(n_3610),
.Y(n_3638)
);

INVx1_ASAP7_75t_L g3639 ( 
.A(n_3617),
.Y(n_3639)
);

INVx1_ASAP7_75t_L g3640 ( 
.A(n_3618),
.Y(n_3640)
);

INVx1_ASAP7_75t_L g3641 ( 
.A(n_3612),
.Y(n_3641)
);

INVx1_ASAP7_75t_L g3642 ( 
.A(n_3620),
.Y(n_3642)
);

INVx1_ASAP7_75t_L g3643 ( 
.A(n_3620),
.Y(n_3643)
);

OAI22xp5_ASAP7_75t_L g3644 ( 
.A1(n_3641),
.A2(n_3605),
.B1(n_3581),
.B2(n_3576),
.Y(n_3644)
);

INVxp67_ASAP7_75t_L g3645 ( 
.A(n_3630),
.Y(n_3645)
);

OA22x2_ASAP7_75t_L g3646 ( 
.A1(n_3639),
.A2(n_3597),
.B1(n_3603),
.B2(n_3616),
.Y(n_3646)
);

AOI221xp5_ASAP7_75t_L g3647 ( 
.A1(n_3636),
.A2(n_3630),
.B1(n_3625),
.B2(n_3640),
.C(n_3623),
.Y(n_3647)
);

INVx1_ASAP7_75t_L g3648 ( 
.A(n_3623),
.Y(n_3648)
);

AO22x2_ASAP7_75t_L g3649 ( 
.A1(n_3624),
.A2(n_3576),
.B1(n_374),
.B2(n_375),
.Y(n_3649)
);

INVx1_ASAP7_75t_SL g3650 ( 
.A(n_3624),
.Y(n_3650)
);

OA22x2_ASAP7_75t_L g3651 ( 
.A1(n_3621),
.A2(n_373),
.B1(n_376),
.B2(n_377),
.Y(n_3651)
);

OAI31xp33_ASAP7_75t_L g3652 ( 
.A1(n_3621),
.A2(n_376),
.A3(n_378),
.B(n_379),
.Y(n_3652)
);

OAI22xp5_ASAP7_75t_L g3653 ( 
.A1(n_3628),
.A2(n_1799),
.B1(n_380),
.B2(n_381),
.Y(n_3653)
);

AND4x1_ASAP7_75t_L g3654 ( 
.A(n_3619),
.B(n_3622),
.C(n_3633),
.D(n_3634),
.Y(n_3654)
);

AOI22xp5_ASAP7_75t_L g3655 ( 
.A1(n_3631),
.A2(n_1799),
.B1(n_383),
.B2(n_386),
.Y(n_3655)
);

HB1xp67_ASAP7_75t_L g3656 ( 
.A(n_3638),
.Y(n_3656)
);

INVx1_ASAP7_75t_L g3657 ( 
.A(n_3638),
.Y(n_3657)
);

AOI22xp5_ASAP7_75t_L g3658 ( 
.A1(n_3626),
.A2(n_378),
.B1(n_386),
.B2(n_387),
.Y(n_3658)
);

INVx2_ASAP7_75t_L g3659 ( 
.A(n_3627),
.Y(n_3659)
);

HB1xp67_ASAP7_75t_L g3660 ( 
.A(n_3629),
.Y(n_3660)
);

NOR2xp67_ASAP7_75t_L g3661 ( 
.A(n_3645),
.B(n_3642),
.Y(n_3661)
);

OAI22xp5_ASAP7_75t_L g3662 ( 
.A1(n_3647),
.A2(n_3637),
.B1(n_3635),
.B2(n_3632),
.Y(n_3662)
);

BUFx2_ASAP7_75t_L g3663 ( 
.A(n_3643),
.Y(n_3663)
);

INVx1_ASAP7_75t_L g3664 ( 
.A(n_3656),
.Y(n_3664)
);

INVx1_ASAP7_75t_L g3665 ( 
.A(n_3648),
.Y(n_3665)
);

INVx1_ASAP7_75t_L g3666 ( 
.A(n_3649),
.Y(n_3666)
);

BUFx2_ASAP7_75t_L g3667 ( 
.A(n_3649),
.Y(n_3667)
);

INVx1_ASAP7_75t_L g3668 ( 
.A(n_3650),
.Y(n_3668)
);

INVx1_ASAP7_75t_L g3669 ( 
.A(n_3657),
.Y(n_3669)
);

INVx1_ASAP7_75t_L g3670 ( 
.A(n_3651),
.Y(n_3670)
);

INVx1_ASAP7_75t_L g3671 ( 
.A(n_3660),
.Y(n_3671)
);

AOI22xp5_ASAP7_75t_L g3672 ( 
.A1(n_3646),
.A2(n_388),
.B1(n_390),
.B2(n_391),
.Y(n_3672)
);

INVx1_ASAP7_75t_L g3673 ( 
.A(n_3659),
.Y(n_3673)
);

INVxp67_ASAP7_75t_L g3674 ( 
.A(n_3644),
.Y(n_3674)
);

AND4x1_ASAP7_75t_L g3675 ( 
.A(n_3652),
.B(n_388),
.C(n_391),
.D(n_392),
.Y(n_3675)
);

OAI22x1_ASAP7_75t_L g3676 ( 
.A1(n_3654),
.A2(n_3658),
.B1(n_3655),
.B2(n_3653),
.Y(n_3676)
);

INVx1_ASAP7_75t_L g3677 ( 
.A(n_3642),
.Y(n_3677)
);

OAI22xp5_ASAP7_75t_SL g3678 ( 
.A1(n_3672),
.A2(n_392),
.B1(n_393),
.B2(n_394),
.Y(n_3678)
);

INVx1_ASAP7_75t_L g3679 ( 
.A(n_3668),
.Y(n_3679)
);

INVx1_ASAP7_75t_L g3680 ( 
.A(n_3663),
.Y(n_3680)
);

AOI22xp5_ASAP7_75t_L g3681 ( 
.A1(n_3670),
.A2(n_393),
.B1(n_394),
.B2(n_395),
.Y(n_3681)
);

NOR2xp67_ASAP7_75t_L g3682 ( 
.A(n_3664),
.B(n_395),
.Y(n_3682)
);

NAND2xp5_ASAP7_75t_L g3683 ( 
.A(n_3674),
.B(n_396),
.Y(n_3683)
);

NAND2xp5_ASAP7_75t_SL g3684 ( 
.A(n_3662),
.B(n_396),
.Y(n_3684)
);

INVx2_ASAP7_75t_L g3685 ( 
.A(n_3665),
.Y(n_3685)
);

AOI22xp5_ASAP7_75t_L g3686 ( 
.A1(n_3661),
.A2(n_397),
.B1(n_398),
.B2(n_399),
.Y(n_3686)
);

AOI22xp5_ASAP7_75t_L g3687 ( 
.A1(n_3676),
.A2(n_398),
.B1(n_399),
.B2(n_400),
.Y(n_3687)
);

NAND2xp5_ASAP7_75t_L g3688 ( 
.A(n_3667),
.B(n_400),
.Y(n_3688)
);

INVx1_ASAP7_75t_L g3689 ( 
.A(n_3671),
.Y(n_3689)
);

AOI22xp5_ASAP7_75t_L g3690 ( 
.A1(n_3666),
.A2(n_402),
.B1(n_403),
.B2(n_404),
.Y(n_3690)
);

INVx1_ASAP7_75t_L g3691 ( 
.A(n_3677),
.Y(n_3691)
);

INVx1_ASAP7_75t_L g3692 ( 
.A(n_3680),
.Y(n_3692)
);

INVx1_ASAP7_75t_L g3693 ( 
.A(n_3681),
.Y(n_3693)
);

INVx1_ASAP7_75t_L g3694 ( 
.A(n_3683),
.Y(n_3694)
);

AOI22xp5_ASAP7_75t_L g3695 ( 
.A1(n_3687),
.A2(n_3673),
.B1(n_3669),
.B2(n_3675),
.Y(n_3695)
);

AOI22xp5_ASAP7_75t_L g3696 ( 
.A1(n_3678),
.A2(n_3679),
.B1(n_3684),
.B2(n_3682),
.Y(n_3696)
);

INVx1_ASAP7_75t_L g3697 ( 
.A(n_3688),
.Y(n_3697)
);

AO22x2_ASAP7_75t_L g3698 ( 
.A1(n_3689),
.A2(n_3675),
.B1(n_403),
.B2(n_405),
.Y(n_3698)
);

NAND2xp5_ASAP7_75t_L g3699 ( 
.A(n_3686),
.B(n_402),
.Y(n_3699)
);

INVx1_ASAP7_75t_L g3700 ( 
.A(n_3685),
.Y(n_3700)
);

NAND2xp5_ASAP7_75t_L g3701 ( 
.A(n_3690),
.B(n_405),
.Y(n_3701)
);

NAND2xp5_ASAP7_75t_SL g3702 ( 
.A(n_3691),
.B(n_408),
.Y(n_3702)
);

NAND2xp5_ASAP7_75t_L g3703 ( 
.A(n_3687),
.B(n_408),
.Y(n_3703)
);

INVx1_ASAP7_75t_L g3704 ( 
.A(n_3680),
.Y(n_3704)
);

INVx1_ASAP7_75t_SL g3705 ( 
.A(n_3679),
.Y(n_3705)
);

NAND5xp2_ASAP7_75t_L g3706 ( 
.A(n_3696),
.B(n_409),
.C(n_410),
.D(n_491),
.E(n_492),
.Y(n_3706)
);

INVx2_ASAP7_75t_L g3707 ( 
.A(n_3700),
.Y(n_3707)
);

AND2x2_ASAP7_75t_L g3708 ( 
.A(n_3698),
.B(n_409),
.Y(n_3708)
);

NOR2x1_ASAP7_75t_L g3709 ( 
.A(n_3692),
.B(n_493),
.Y(n_3709)
);

INVx1_ASAP7_75t_L g3710 ( 
.A(n_3703),
.Y(n_3710)
);

INVx1_ASAP7_75t_L g3711 ( 
.A(n_3699),
.Y(n_3711)
);

BUFx2_ASAP7_75t_L g3712 ( 
.A(n_3704),
.Y(n_3712)
);

OAI22xp5_ASAP7_75t_L g3713 ( 
.A1(n_3707),
.A2(n_3695),
.B1(n_3693),
.B2(n_3705),
.Y(n_3713)
);

INVx2_ASAP7_75t_L g3714 ( 
.A(n_3708),
.Y(n_3714)
);

AND2x4_ASAP7_75t_L g3715 ( 
.A(n_3711),
.B(n_3694),
.Y(n_3715)
);

INVx2_ASAP7_75t_L g3716 ( 
.A(n_3712),
.Y(n_3716)
);

INVx1_ASAP7_75t_L g3717 ( 
.A(n_3710),
.Y(n_3717)
);

INVx1_ASAP7_75t_L g3718 ( 
.A(n_3714),
.Y(n_3718)
);

OAI22x1_ASAP7_75t_L g3719 ( 
.A1(n_3716),
.A2(n_3697),
.B1(n_3702),
.B2(n_3709),
.Y(n_3719)
);

OAI22xp5_ASAP7_75t_L g3720 ( 
.A1(n_3713),
.A2(n_3701),
.B1(n_3706),
.B2(n_499),
.Y(n_3720)
);

INVx1_ASAP7_75t_L g3721 ( 
.A(n_3717),
.Y(n_3721)
);

AOI22xp5_ASAP7_75t_L g3722 ( 
.A1(n_3715),
.A2(n_3706),
.B1(n_497),
.B2(n_501),
.Y(n_3722)
);

INVx2_ASAP7_75t_L g3723 ( 
.A(n_3718),
.Y(n_3723)
);

INVx1_ASAP7_75t_L g3724 ( 
.A(n_3721),
.Y(n_3724)
);

INVx1_ASAP7_75t_L g3725 ( 
.A(n_3719),
.Y(n_3725)
);

AOI22xp5_ASAP7_75t_L g3726 ( 
.A1(n_3723),
.A2(n_3720),
.B1(n_3722),
.B2(n_509),
.Y(n_3726)
);

INVx1_ASAP7_75t_SL g3727 ( 
.A(n_3726),
.Y(n_3727)
);

AO22x2_ASAP7_75t_L g3728 ( 
.A1(n_3727),
.A2(n_3725),
.B1(n_3724),
.B2(n_510),
.Y(n_3728)
);

INVx2_ASAP7_75t_L g3729 ( 
.A(n_3728),
.Y(n_3729)
);

AOI221xp5_ASAP7_75t_L g3730 ( 
.A1(n_3729),
.A2(n_496),
.B1(n_508),
.B2(n_511),
.C(n_513),
.Y(n_3730)
);

AOI211xp5_ASAP7_75t_L g3731 ( 
.A1(n_3730),
.A2(n_516),
.B(n_517),
.C(n_519),
.Y(n_3731)
);


endmodule