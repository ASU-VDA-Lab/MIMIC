module fake_jpeg_13716_n_307 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_307);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_307;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_208;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_4),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_1),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_12),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

BUFx12_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_14),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_7),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_12),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_2),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_6),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_6),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_4),
.Y(n_35)
);

INVx13_ASAP7_75t_L g36 ( 
.A(n_0),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_8),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_2),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_3),
.Y(n_39)
);

BUFx10_ASAP7_75t_L g40 ( 
.A(n_9),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_16),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_1),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_13),
.Y(n_43)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_0),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_14),
.Y(n_45)
);

CKINVDCx14_ASAP7_75t_R g46 ( 
.A(n_16),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_14),
.Y(n_47)
);

BUFx12_ASAP7_75t_L g48 ( 
.A(n_13),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_46),
.B(n_0),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_SL g108 ( 
.A(n_49),
.B(n_68),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_20),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_50),
.Y(n_97)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_22),
.Y(n_51)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_51),
.Y(n_114)
);

INVx5_ASAP7_75t_L g52 ( 
.A(n_18),
.Y(n_52)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_52),
.Y(n_116)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_18),
.Y(n_53)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_53),
.Y(n_96)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_18),
.Y(n_54)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_54),
.Y(n_102)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_22),
.Y(n_55)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_55),
.Y(n_127)
);

INVx4_ASAP7_75t_SL g56 ( 
.A(n_40),
.Y(n_56)
);

INVx13_ASAP7_75t_L g119 ( 
.A(n_56),
.Y(n_119)
);

INVx5_ASAP7_75t_L g57 ( 
.A(n_18),
.Y(n_57)
);

INVx3_ASAP7_75t_L g131 ( 
.A(n_57),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_20),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_58),
.Y(n_103)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_26),
.Y(n_59)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_59),
.Y(n_135)
);

INVx11_ASAP7_75t_L g60 ( 
.A(n_40),
.Y(n_60)
);

BUFx5_ASAP7_75t_L g99 ( 
.A(n_60),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_41),
.B(n_1),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_61),
.B(n_81),
.Y(n_106)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_24),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g144 ( 
.A(n_62),
.Y(n_144)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_26),
.Y(n_63)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_63),
.Y(n_138)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_20),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_64),
.Y(n_104)
);

BUFx12f_ASAP7_75t_L g65 ( 
.A(n_24),
.Y(n_65)
);

INVx5_ASAP7_75t_L g124 ( 
.A(n_65),
.Y(n_124)
);

BUFx12f_ASAP7_75t_L g66 ( 
.A(n_47),
.Y(n_66)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_66),
.Y(n_101)
);

HB1xp67_ASAP7_75t_L g67 ( 
.A(n_40),
.Y(n_67)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_67),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_17),
.B(n_2),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_17),
.B(n_3),
.Y(n_69)
);

AND2x2_ASAP7_75t_L g105 ( 
.A(n_69),
.B(n_73),
.Y(n_105)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_40),
.Y(n_70)
);

INVx4_ASAP7_75t_L g111 ( 
.A(n_70),
.Y(n_111)
);

BUFx4f_ASAP7_75t_SL g71 ( 
.A(n_40),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_71),
.Y(n_118)
);

BUFx5_ASAP7_75t_L g72 ( 
.A(n_27),
.Y(n_72)
);

INVx4_ASAP7_75t_L g120 ( 
.A(n_72),
.Y(n_120)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_44),
.Y(n_73)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_27),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_74),
.Y(n_129)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_47),
.Y(n_75)
);

INVx3_ASAP7_75t_L g134 ( 
.A(n_75),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_SL g76 ( 
.A(n_41),
.B(n_15),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_76),
.B(n_80),
.Y(n_98)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_44),
.Y(n_77)
);

INVx6_ASAP7_75t_L g94 ( 
.A(n_77),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_27),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g141 ( 
.A(n_78),
.Y(n_141)
);

INVx8_ASAP7_75t_L g79 ( 
.A(n_29),
.Y(n_79)
);

BUFx10_ASAP7_75t_L g143 ( 
.A(n_79),
.Y(n_143)
);

BUFx12f_ASAP7_75t_L g80 ( 
.A(n_29),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_19),
.B(n_4),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_SL g82 ( 
.A(n_19),
.B(n_30),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_82),
.B(n_89),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_35),
.B(n_5),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_83),
.B(n_85),
.Y(n_107)
);

INVx5_ASAP7_75t_L g84 ( 
.A(n_29),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g117 ( 
.A(n_84),
.B(n_86),
.Y(n_117)
);

CKINVDCx16_ASAP7_75t_R g85 ( 
.A(n_36),
.Y(n_85)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_31),
.Y(n_86)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_31),
.Y(n_87)
);

AND2x2_ASAP7_75t_L g126 ( 
.A(n_87),
.B(n_88),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_31),
.Y(n_88)
);

INVx5_ASAP7_75t_L g89 ( 
.A(n_33),
.Y(n_89)
);

INVx5_ASAP7_75t_L g90 ( 
.A(n_33),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_90),
.B(n_91),
.Y(n_113)
);

INVx5_ASAP7_75t_L g91 ( 
.A(n_33),
.Y(n_91)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_34),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_92),
.B(n_93),
.Y(n_130)
);

BUFx5_ASAP7_75t_L g93 ( 
.A(n_34),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_64),
.A2(n_88),
.B1(n_78),
.B2(n_58),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_95),
.A2(n_110),
.B1(n_115),
.B2(n_122),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_83),
.B(n_35),
.C(n_45),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_100),
.B(n_11),
.C(n_13),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_67),
.A2(n_37),
.B1(n_45),
.B2(n_43),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_68),
.B(n_28),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_112),
.B(n_121),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_65),
.A2(n_34),
.B1(n_43),
.B2(n_42),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_69),
.B(n_25),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_79),
.A2(n_37),
.B1(n_42),
.B2(n_39),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_50),
.A2(n_49),
.B1(n_38),
.B2(n_32),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_125),
.A2(n_128),
.B1(n_120),
.B2(n_99),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_80),
.A2(n_28),
.B1(n_21),
.B2(n_25),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_85),
.B(n_21),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_132),
.B(n_136),
.Y(n_174)
);

AOI22xp33_ASAP7_75t_L g133 ( 
.A1(n_56),
.A2(n_39),
.B1(n_38),
.B2(n_32),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_133),
.A2(n_140),
.B1(n_142),
.B2(n_115),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_66),
.B(n_30),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_71),
.B(n_15),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_SL g179 ( 
.A(n_137),
.B(n_139),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_83),
.B(n_7),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_73),
.A2(n_48),
.B1(n_23),
.B2(n_10),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_L g142 ( 
.A1(n_74),
.A2(n_36),
.B1(n_48),
.B2(n_23),
.Y(n_142)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_123),
.Y(n_145)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_145),
.Y(n_190)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_135),
.Y(n_146)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_146),
.Y(n_192)
);

AND2x2_ASAP7_75t_L g147 ( 
.A(n_105),
.B(n_107),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_147),
.B(n_172),
.C(n_185),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_108),
.B(n_7),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_SL g191 ( 
.A(n_148),
.B(n_151),
.Y(n_191)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_104),
.Y(n_150)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_150),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_98),
.B(n_8),
.Y(n_151)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_104),
.Y(n_152)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_152),
.Y(n_199)
);

INVx4_ASAP7_75t_L g153 ( 
.A(n_118),
.Y(n_153)
);

INVx4_ASAP7_75t_L g214 ( 
.A(n_153),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_133),
.A2(n_36),
.B1(n_48),
.B2(n_23),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_154),
.A2(n_176),
.B1(n_178),
.B2(n_185),
.Y(n_197)
);

A2O1A1Ixp33_ASAP7_75t_L g155 ( 
.A1(n_105),
.A2(n_8),
.B(n_11),
.C(n_12),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_155),
.B(n_167),
.Y(n_193)
);

BUFx8_ASAP7_75t_L g156 ( 
.A(n_119),
.Y(n_156)
);

INVxp67_ASAP7_75t_L g216 ( 
.A(n_156),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_157),
.B(n_169),
.Y(n_189)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_138),
.Y(n_158)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_158),
.Y(n_213)
);

BUFx6f_ASAP7_75t_L g159 ( 
.A(n_97),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g206 ( 
.A(n_159),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_109),
.B(n_106),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_SL g200 ( 
.A(n_160),
.B(n_162),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_114),
.B(n_23),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_127),
.B(n_48),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_SL g207 ( 
.A(n_163),
.B(n_166),
.Y(n_207)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_96),
.Y(n_164)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_164),
.Y(n_218)
);

BUFx3_ASAP7_75t_L g165 ( 
.A(n_118),
.Y(n_165)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_165),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_134),
.B(n_102),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_122),
.B(n_126),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_130),
.B(n_131),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_SL g208 ( 
.A(n_168),
.B(n_170),
.Y(n_208)
);

INVx3_ASAP7_75t_L g169 ( 
.A(n_101),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_116),
.B(n_113),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_94),
.B(n_101),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_171),
.B(n_180),
.Y(n_222)
);

MAJx2_ASAP7_75t_L g172 ( 
.A(n_117),
.B(n_126),
.C(n_143),
.Y(n_172)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_111),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_173),
.B(n_175),
.Y(n_201)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_94),
.Y(n_175)
);

INVx13_ASAP7_75t_L g177 ( 
.A(n_119),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_177),
.B(n_183),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_142),
.A2(n_129),
.B1(n_103),
.B2(n_141),
.Y(n_178)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_117),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_111),
.B(n_97),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_181),
.B(n_182),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_103),
.B(n_141),
.Y(n_182)
);

INVx3_ASAP7_75t_SL g183 ( 
.A(n_143),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_129),
.B(n_143),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_184),
.B(n_187),
.Y(n_211)
);

AND2x2_ASAP7_75t_L g185 ( 
.A(n_124),
.B(n_144),
.Y(n_185)
);

OAI32xp33_ASAP7_75t_L g186 ( 
.A1(n_120),
.A2(n_107),
.A3(n_106),
.B1(n_139),
.B2(n_108),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g195 ( 
.A(n_186),
.B(n_147),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_144),
.B(n_124),
.Y(n_187)
);

OA22x2_ASAP7_75t_L g204 ( 
.A1(n_188),
.A2(n_150),
.B1(n_152),
.B2(n_155),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_167),
.A2(n_188),
.B1(n_180),
.B2(n_149),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_194),
.A2(n_196),
.B1(n_198),
.B2(n_204),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_195),
.B(n_202),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_184),
.A2(n_182),
.B1(n_181),
.B2(n_147),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_L g240 ( 
.A1(n_197),
.A2(n_211),
.B1(n_202),
.B2(n_194),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_172),
.A2(n_174),
.B1(n_186),
.B2(n_154),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_161),
.B(n_157),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_205),
.B(n_212),
.C(n_211),
.Y(n_247)
);

AOI22x1_ASAP7_75t_SL g209 ( 
.A1(n_146),
.A2(n_153),
.B1(n_173),
.B2(n_158),
.Y(n_209)
);

AOI21xp5_ASAP7_75t_L g231 ( 
.A1(n_209),
.A2(n_210),
.B(n_165),
.Y(n_231)
);

AOI21xp5_ASAP7_75t_L g210 ( 
.A1(n_185),
.A2(n_169),
.B(n_177),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_L g212 ( 
.A(n_145),
.B(n_164),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_156),
.B(n_159),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_215),
.B(n_217),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_156),
.B(n_183),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_200),
.B(n_208),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_SL g263 ( 
.A(n_223),
.B(n_232),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_201),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_224),
.B(n_227),
.Y(n_250)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_192),
.Y(n_226)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_226),
.Y(n_253)
);

BUFx4f_ASAP7_75t_SL g227 ( 
.A(n_216),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_190),
.Y(n_228)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_228),
.Y(n_262)
);

HAxp5_ASAP7_75t_SL g229 ( 
.A(n_193),
.B(n_179),
.CON(n_229),
.SN(n_229)
);

BUFx24_ASAP7_75t_SL g255 ( 
.A(n_229),
.Y(n_255)
);

CKINVDCx14_ASAP7_75t_R g230 ( 
.A(n_217),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_230),
.B(n_233),
.Y(n_258)
);

OAI21xp5_ASAP7_75t_L g257 ( 
.A1(n_231),
.A2(n_236),
.B(n_239),
.Y(n_257)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_199),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_207),
.B(n_222),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_SL g234 ( 
.A(n_205),
.B(n_189),
.Y(n_234)
);

AOI221xp5_ASAP7_75t_L g251 ( 
.A1(n_234),
.A2(n_244),
.B1(n_245),
.B2(n_246),
.C(n_203),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_215),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_235),
.Y(n_249)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_213),
.Y(n_236)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_220),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_237),
.A2(n_240),
.B1(n_241),
.B2(n_243),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_238),
.B(n_247),
.C(n_196),
.Y(n_248)
);

INVxp33_ASAP7_75t_L g239 ( 
.A(n_219),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_197),
.A2(n_203),
.B1(n_193),
.B2(n_198),
.Y(n_241)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_220),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_191),
.B(n_195),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_218),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_209),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_248),
.B(n_260),
.C(n_264),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_SL g265 ( 
.A(n_251),
.B(n_254),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_242),
.A2(n_204),
.B1(n_210),
.B2(n_212),
.Y(n_252)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_252),
.Y(n_267)
);

AOI322xp5_ASAP7_75t_L g254 ( 
.A1(n_240),
.A2(n_204),
.A3(n_206),
.B1(n_214),
.B2(n_216),
.C1(n_221),
.C2(n_241),
.Y(n_254)
);

OAI32xp33_ASAP7_75t_L g259 ( 
.A1(n_242),
.A2(n_204),
.A3(n_206),
.B1(n_214),
.B2(n_238),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_259),
.B(n_227),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_247),
.B(n_234),
.C(n_235),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_246),
.A2(n_225),
.B1(n_224),
.B2(n_231),
.Y(n_261)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_261),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_225),
.B(n_223),
.C(n_228),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_264),
.B(n_226),
.Y(n_266)
);

AOI21xp33_ASAP7_75t_L g280 ( 
.A1(n_266),
.A2(n_268),
.B(n_263),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_263),
.B(n_250),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_248),
.B(n_236),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_269),
.B(n_274),
.C(n_270),
.Y(n_282)
);

OAI21xp5_ASAP7_75t_SL g271 ( 
.A1(n_261),
.A2(n_227),
.B(n_232),
.Y(n_271)
);

OAI21xp5_ASAP7_75t_SL g278 ( 
.A1(n_271),
.A2(n_277),
.B(n_249),
.Y(n_278)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_253),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_260),
.B(n_245),
.C(n_237),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_253),
.Y(n_275)
);

NAND2xp33_ASAP7_75t_SL g283 ( 
.A(n_275),
.B(n_276),
.Y(n_283)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_262),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_278),
.B(n_271),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_L g279 ( 
.A1(n_272),
.A2(n_256),
.B1(n_249),
.B2(n_257),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_SL g291 ( 
.A1(n_279),
.A2(n_284),
.B1(n_267),
.B2(n_276),
.Y(n_291)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_280),
.Y(n_288)
);

XOR2xp5_ASAP7_75t_L g281 ( 
.A(n_269),
.B(n_259),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_281),
.B(n_282),
.C(n_285),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_267),
.A2(n_256),
.B1(n_257),
.B2(n_252),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_270),
.B(n_258),
.C(n_262),
.Y(n_285)
);

OR2x2_ASAP7_75t_L g296 ( 
.A(n_286),
.B(n_279),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_282),
.B(n_274),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_287),
.B(n_290),
.C(n_284),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_285),
.B(n_265),
.C(n_272),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_291),
.B(n_292),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_281),
.B(n_273),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_294),
.B(n_289),
.C(n_290),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_288),
.B(n_278),
.Y(n_295)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_295),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_296),
.B(n_297),
.Y(n_298)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_292),
.Y(n_297)
);

INVxp67_ASAP7_75t_L g302 ( 
.A(n_299),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_293),
.B(n_289),
.C(n_255),
.Y(n_300)
);

INVxp67_ASAP7_75t_L g303 ( 
.A(n_300),
.Y(n_303)
);

AOI21xp5_ASAP7_75t_SL g304 ( 
.A1(n_302),
.A2(n_301),
.B(n_298),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_304),
.B(n_305),
.Y(n_306)
);

INVxp67_ASAP7_75t_L g305 ( 
.A(n_303),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_L g307 ( 
.A(n_306),
.B(n_283),
.Y(n_307)
);


endmodule