module fake_jpeg_7572_n_202 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_202);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_202;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_154;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g15 ( 
.A(n_0),
.Y(n_15)
);

BUFx12_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_3),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

INVx5_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_1),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_10),
.Y(n_22)
);

BUFx10_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

CKINVDCx14_ASAP7_75t_R g26 ( 
.A(n_11),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_5),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_20),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_32),
.B(n_40),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_29),
.Y(n_33)
);

INVx4_ASAP7_75t_SL g62 ( 
.A(n_33),
.Y(n_62)
);

INVx4_ASAP7_75t_SL g34 ( 
.A(n_25),
.Y(n_34)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_34),
.A2(n_20),
.B1(n_30),
.B2(n_17),
.Y(n_54)
);

BUFx16f_ASAP7_75t_L g35 ( 
.A(n_23),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_27),
.B(n_1),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_36),
.B(n_38),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_27),
.B(n_31),
.Y(n_37)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_37),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_18),
.B(n_1),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_18),
.B(n_2),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_39),
.B(n_19),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_29),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_29),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_41),
.Y(n_48)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_25),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_42),
.B(n_24),
.Y(n_44)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_44),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_47),
.B(n_49),
.Y(n_75)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_L g50 ( 
.A1(n_36),
.A2(n_24),
.B1(n_20),
.B2(n_21),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_50),
.A2(n_23),
.B1(n_16),
.B2(n_5),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_38),
.B(n_15),
.Y(n_51)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_51),
.Y(n_72)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_35),
.Y(n_52)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_52),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_35),
.Y(n_53)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_53),
.Y(n_77)
);

OAI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_54),
.A2(n_23),
.B1(n_16),
.B2(n_5),
.Y(n_80)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_35),
.Y(n_56)
);

BUFx2_ASAP7_75t_L g65 ( 
.A(n_56),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g57 ( 
.A1(n_32),
.A2(n_26),
.B1(n_30),
.B2(n_28),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_57),
.A2(n_26),
.B1(n_17),
.B2(n_28),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_42),
.Y(n_58)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_58),
.Y(n_67)
);

BUFx4f_ASAP7_75t_SL g59 ( 
.A(n_33),
.Y(n_59)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_59),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_37),
.B(n_29),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_60),
.B(n_22),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_39),
.B(n_40),
.Y(n_61)
);

OR2x2_ASAP7_75t_L g71 ( 
.A(n_61),
.B(n_16),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_63),
.B(n_71),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_45),
.A2(n_42),
.B1(n_34),
.B2(n_32),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_64),
.A2(n_69),
.B1(n_81),
.B2(n_62),
.Y(n_83)
);

O2A1O1Ixp33_ASAP7_75t_L g66 ( 
.A1(n_57),
.A2(n_15),
.B(n_19),
.C(n_34),
.Y(n_66)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_66),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_45),
.A2(n_34),
.B1(n_21),
.B2(n_31),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_L g70 ( 
.A1(n_55),
.A2(n_22),
.B1(n_25),
.B2(n_23),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_70),
.A2(n_80),
.B1(n_62),
.B2(n_47),
.Y(n_82)
);

XNOR2xp5_ASAP7_75t_L g96 ( 
.A(n_73),
.B(n_52),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_55),
.B(n_60),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_76),
.B(n_52),
.C(n_46),
.Y(n_95)
);

OR2x2_ASAP7_75t_L g79 ( 
.A(n_43),
.B(n_16),
.Y(n_79)
);

OAI21xp5_ASAP7_75t_L g88 ( 
.A1(n_79),
.A2(n_23),
.B(n_59),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_82),
.A2(n_83),
.B1(n_85),
.B2(n_91),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_81),
.A2(n_62),
.B1(n_58),
.B2(n_41),
.Y(n_85)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_64),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_86),
.B(n_87),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_78),
.B(n_56),
.Y(n_87)
);

XNOR2x1_ASAP7_75t_SL g113 ( 
.A(n_88),
.B(n_102),
.Y(n_113)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_75),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_90),
.B(n_98),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_76),
.A2(n_33),
.B1(n_41),
.B2(n_48),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_76),
.A2(n_68),
.B1(n_73),
.B2(n_72),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_92),
.A2(n_93),
.B1(n_94),
.B2(n_97),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_68),
.A2(n_33),
.B1(n_41),
.B2(n_48),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_72),
.A2(n_59),
.B1(n_49),
.B2(n_53),
.Y(n_94)
);

XOR2xp5_ASAP7_75t_L g107 ( 
.A(n_95),
.B(n_69),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_SL g106 ( 
.A(n_96),
.B(n_71),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_75),
.A2(n_52),
.B1(n_46),
.B2(n_14),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_78),
.B(n_46),
.Y(n_98)
);

INVxp67_ASAP7_75t_L g99 ( 
.A(n_66),
.Y(n_99)
);

INVxp67_ASAP7_75t_SL g109 ( 
.A(n_99),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_74),
.B(n_79),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_100),
.B(n_101),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_74),
.B(n_46),
.Y(n_101)
);

NAND2x1_ASAP7_75t_SL g102 ( 
.A(n_79),
.B(n_2),
.Y(n_102)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_94),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_104),
.B(n_111),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_106),
.B(n_107),
.C(n_112),
.Y(n_127)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_93),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_108),
.B(n_115),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_97),
.Y(n_111)
);

XOR2xp5_ASAP7_75t_L g112 ( 
.A(n_96),
.B(n_71),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_86),
.A2(n_63),
.B1(n_77),
.B2(n_7),
.Y(n_114)
);

INVxp67_ASAP7_75t_L g135 ( 
.A(n_114),
.Y(n_135)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_91),
.Y(n_115)
);

AND2x4_ASAP7_75t_L g117 ( 
.A(n_88),
.B(n_67),
.Y(n_117)
);

AND2x2_ASAP7_75t_L g131 ( 
.A(n_117),
.B(n_102),
.Y(n_131)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_85),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_118),
.B(n_120),
.Y(n_126)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_95),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_90),
.B(n_65),
.Y(n_121)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_121),
.Y(n_128)
);

OAI22xp33_ASAP7_75t_L g123 ( 
.A1(n_118),
.A2(n_99),
.B1(n_84),
.B2(n_89),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_123),
.A2(n_104),
.B1(n_108),
.B2(n_115),
.Y(n_141)
);

XOR2xp5_ASAP7_75t_L g124 ( 
.A(n_112),
.B(n_107),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_124),
.B(n_133),
.C(n_137),
.Y(n_146)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_121),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_125),
.B(n_130),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_111),
.A2(n_89),
.B1(n_84),
.B2(n_83),
.Y(n_129)
);

CKINVDCx14_ASAP7_75t_R g142 ( 
.A(n_129),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_109),
.B(n_77),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_L g140 ( 
.A1(n_131),
.A2(n_132),
.B(n_117),
.Y(n_140)
);

AOI21xp5_ASAP7_75t_L g132 ( 
.A1(n_117),
.A2(n_113),
.B(n_103),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_120),
.B(n_92),
.C(n_82),
.Y(n_133)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_105),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_134),
.B(n_136),
.Y(n_150)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_119),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_106),
.B(n_102),
.C(n_65),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_113),
.B(n_65),
.C(n_67),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_138),
.B(n_6),
.Y(n_154)
);

XOR2xp5_ASAP7_75t_L g155 ( 
.A(n_140),
.B(n_154),
.Y(n_155)
);

CKINVDCx14_ASAP7_75t_R g163 ( 
.A(n_141),
.Y(n_163)
);

INVx1_ASAP7_75t_SL g143 ( 
.A(n_122),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_143),
.B(n_151),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_SL g144 ( 
.A(n_126),
.B(n_114),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_SL g158 ( 
.A(n_144),
.B(n_137),
.Y(n_158)
);

AND2x2_ASAP7_75t_L g147 ( 
.A(n_138),
.B(n_117),
.Y(n_147)
);

AOI21xp5_ASAP7_75t_SL g162 ( 
.A1(n_147),
.A2(n_152),
.B(n_127),
.Y(n_162)
);

HB1xp67_ASAP7_75t_L g148 ( 
.A(n_128),
.Y(n_148)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_148),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_139),
.A2(n_110),
.B1(n_116),
.B2(n_7),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_149),
.A2(n_153),
.B1(n_8),
.B2(n_9),
.Y(n_167)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_128),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_L g152 ( 
.A1(n_132),
.A2(n_4),
.B(n_6),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_135),
.A2(n_4),
.B1(n_6),
.B2(n_8),
.Y(n_153)
);

A2O1A1Ixp33_ASAP7_75t_L g157 ( 
.A1(n_142),
.A2(n_135),
.B(n_131),
.C(n_123),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_157),
.B(n_158),
.Y(n_177)
);

OAI211xp5_ASAP7_75t_SL g160 ( 
.A1(n_140),
.A2(n_131),
.B(n_133),
.C(n_124),
.Y(n_160)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_160),
.Y(n_168)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_145),
.Y(n_161)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_161),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_L g173 ( 
.A1(n_162),
.A2(n_165),
.B(n_166),
.Y(n_173)
);

INVx13_ASAP7_75t_L g164 ( 
.A(n_143),
.Y(n_164)
);

CKINVDCx16_ASAP7_75t_R g170 ( 
.A(n_164),
.Y(n_170)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_150),
.Y(n_165)
);

INVx13_ASAP7_75t_L g166 ( 
.A(n_151),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_L g174 ( 
.A(n_167),
.B(n_153),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g169 ( 
.A(n_160),
.B(n_146),
.Y(n_169)
);

XOR2xp5_ASAP7_75t_L g183 ( 
.A(n_169),
.B(n_156),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_155),
.B(n_146),
.C(n_127),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_172),
.B(n_175),
.C(n_176),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_174),
.B(n_167),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_155),
.B(n_147),
.C(n_149),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_158),
.B(n_147),
.C(n_144),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_178),
.B(n_179),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_170),
.B(n_156),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_172),
.B(n_165),
.C(n_161),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_180),
.B(n_183),
.Y(n_190)
);

NOR2xp67_ASAP7_75t_SL g181 ( 
.A(n_173),
.B(n_162),
.Y(n_181)
);

INVxp67_ASAP7_75t_SL g188 ( 
.A(n_181),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_168),
.A2(n_171),
.B1(n_163),
.B2(n_157),
.Y(n_182)
);

AOI322xp5_ASAP7_75t_L g189 ( 
.A1(n_182),
.A2(n_184),
.A3(n_166),
.B1(n_152),
.B2(n_174),
.C1(n_141),
.C2(n_175),
.Y(n_189)
);

OAI22xp33_ASAP7_75t_SL g184 ( 
.A1(n_177),
.A2(n_166),
.B1(n_159),
.B2(n_164),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_SL g187 ( 
.A(n_183),
.B(n_159),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_187),
.B(n_184),
.Y(n_192)
);

INVxp67_ASAP7_75t_SL g195 ( 
.A(n_189),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_185),
.B(n_176),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_191),
.B(n_185),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_192),
.B(n_193),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_187),
.B(n_169),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_194),
.B(n_9),
.C(n_10),
.Y(n_197)
);

AOI22xp33_ASAP7_75t_L g196 ( 
.A1(n_195),
.A2(n_186),
.B1(n_188),
.B2(n_190),
.Y(n_196)
);

AOI21x1_ASAP7_75t_L g199 ( 
.A1(n_196),
.A2(n_11),
.B(n_12),
.Y(n_199)
);

MAJx2_ASAP7_75t_L g200 ( 
.A(n_197),
.B(n_11),
.C(n_12),
.Y(n_200)
);

O2A1O1Ixp33_ASAP7_75t_SL g201 ( 
.A1(n_199),
.A2(n_200),
.B(n_12),
.C(n_13),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_201),
.A2(n_13),
.B1(n_198),
.B2(n_167),
.Y(n_202)
);


endmodule