module fake_netlist_6_3957_n_1113 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_193, n_147, n_154, n_191, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_199, n_138, n_22, n_161, n_68, n_166, n_28, n_184, n_50, n_158, n_49, n_7, n_83, n_206, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_178, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_188, n_102, n_186, n_204, n_0, n_87, n_195, n_189, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_197, n_11, n_137, n_17, n_23, n_203, n_142, n_20, n_143, n_207, n_2, n_180, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_205, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_181, n_76, n_36, n_182, n_26, n_124, n_55, n_126, n_202, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_175, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_196, n_200, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_198, n_104, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_6, n_190, n_14, n_123, n_136, n_72, n_187, n_89, n_173, n_201, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_185, n_35, n_183, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_194, n_171, n_31, n_192, n_57, n_169, n_53, n_51, n_44, n_56, n_1113);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_193;
input n_147;
input n_154;
input n_191;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_199;
input n_138;
input n_22;
input n_161;
input n_68;
input n_166;
input n_28;
input n_184;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_206;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_178;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_188;
input n_102;
input n_186;
input n_204;
input n_0;
input n_87;
input n_195;
input n_189;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_197;
input n_11;
input n_137;
input n_17;
input n_23;
input n_203;
input n_142;
input n_20;
input n_143;
input n_207;
input n_2;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_205;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_55;
input n_126;
input n_202;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_175;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_196;
input n_200;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_190;
input n_14;
input n_123;
input n_136;
input n_72;
input n_187;
input n_89;
input n_173;
input n_201;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_185;
input n_35;
input n_183;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_194;
input n_171;
input n_31;
input n_192;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1113;

wire n_992;
wire n_591;
wire n_435;
wire n_793;
wire n_326;
wire n_801;
wire n_256;
wire n_853;
wire n_440;
wire n_587;
wire n_695;
wire n_507;
wire n_968;
wire n_909;
wire n_580;
wire n_762;
wire n_1030;
wire n_881;
wire n_875;
wire n_209;
wire n_367;
wire n_465;
wire n_680;
wire n_741;
wire n_760;
wire n_1008;
wire n_1027;
wire n_590;
wire n_625;
wire n_661;
wire n_223;
wire n_278;
wire n_1079;
wire n_341;
wire n_362;
wire n_226;
wire n_828;
wire n_208;
wire n_462;
wire n_607;
wire n_671;
wire n_726;
wire n_1033;
wire n_316;
wire n_419;
wire n_304;
wire n_212;
wire n_700;
wire n_694;
wire n_1103;
wire n_933;
wire n_740;
wire n_1038;
wire n_578;
wire n_703;
wire n_1003;
wire n_365;
wire n_978;
wire n_1061;
wire n_384;
wire n_297;
wire n_595;
wire n_627;
wire n_524;
wire n_342;
wire n_820;
wire n_1044;
wire n_951;
wire n_783;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_751;
wire n_449;
wire n_749;
wire n_798;
wire n_310;
wire n_509;
wire n_245;
wire n_368;
wire n_575;
wire n_994;
wire n_1072;
wire n_677;
wire n_969;
wire n_988;
wire n_805;
wire n_396;
wire n_495;
wire n_1065;
wire n_815;
wire n_350;
wire n_1100;
wire n_585;
wire n_732;
wire n_974;
wire n_568;
wire n_392;
wire n_840;
wire n_442;
wire n_480;
wire n_874;
wire n_724;
wire n_382;
wire n_673;
wire n_1020;
wire n_1009;
wire n_1042;
wire n_1071;
wire n_628;
wire n_1067;
wire n_883;
wire n_557;
wire n_823;
wire n_349;
wire n_643;
wire n_233;
wire n_617;
wire n_698;
wire n_898;
wire n_1074;
wire n_1032;
wire n_845;
wire n_255;
wire n_807;
wire n_1036;
wire n_739;
wire n_284;
wire n_400;
wire n_337;
wire n_955;
wire n_865;
wire n_893;
wire n_214;
wire n_925;
wire n_485;
wire n_1101;
wire n_1026;
wire n_443;
wire n_1099;
wire n_246;
wire n_892;
wire n_768;
wire n_1097;
wire n_471;
wire n_289;
wire n_935;
wire n_421;
wire n_781;
wire n_424;
wire n_789;
wire n_615;
wire n_238;
wire n_1095;
wire n_573;
wire n_769;
wire n_320;
wire n_639;
wire n_676;
wire n_327;
wire n_794;
wire n_963;
wire n_727;
wire n_894;
wire n_369;
wire n_597;
wire n_685;
wire n_280;
wire n_287;
wire n_832;
wire n_353;
wire n_610;
wire n_555;
wire n_389;
wire n_814;
wire n_415;
wire n_830;
wire n_230;
wire n_605;
wire n_461;
wire n_873;
wire n_383;
wire n_826;
wire n_1024;
wire n_669;
wire n_447;
wire n_872;
wire n_300;
wire n_222;
wire n_248;
wire n_718;
wire n_517;
wire n_1018;
wire n_747;
wire n_852;
wire n_667;
wire n_229;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_1105;
wire n_621;
wire n_305;
wire n_1037;
wire n_721;
wire n_996;
wire n_750;
wire n_532;
wire n_742;
wire n_535;
wire n_691;
wire n_250;
wire n_372;
wire n_468;
wire n_544;
wire n_901;
wire n_504;
wire n_923;
wire n_314;
wire n_378;
wire n_413;
wire n_377;
wire n_791;
wire n_510;
wire n_837;
wire n_836;
wire n_1015;
wire n_863;
wire n_375;
wire n_601;
wire n_338;
wire n_522;
wire n_948;
wire n_466;
wire n_704;
wire n_918;
wire n_748;
wire n_506;
wire n_763;
wire n_1057;
wire n_360;
wire n_977;
wire n_945;
wire n_603;
wire n_1005;
wire n_991;
wire n_957;
wire n_235;
wire n_536;
wire n_895;
wire n_866;
wire n_622;
wire n_340;
wire n_710;
wire n_1108;
wire n_387;
wire n_452;
wire n_616;
wire n_658;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_581;
wire n_428;
wire n_761;
wire n_785;
wire n_746;
wire n_609;
wire n_765;
wire n_432;
wire n_987;
wire n_641;
wire n_822;
wire n_693;
wire n_1056;
wire n_631;
wire n_516;
wire n_720;
wire n_758;
wire n_525;
wire n_842;
wire n_611;
wire n_943;
wire n_491;
wire n_878;
wire n_656;
wire n_772;
wire n_843;
wire n_989;
wire n_797;
wire n_666;
wire n_1016;
wire n_371;
wire n_795;
wire n_770;
wire n_940;
wire n_567;
wire n_899;
wire n_738;
wire n_405;
wire n_213;
wire n_538;
wire n_1035;
wire n_294;
wire n_302;
wire n_499;
wire n_380;
wire n_838;
wire n_705;
wire n_647;
wire n_343;
wire n_844;
wire n_448;
wire n_886;
wire n_1017;
wire n_1004;
wire n_953;
wire n_1094;
wire n_494;
wire n_539;
wire n_493;
wire n_397;
wire n_1022;
wire n_1083;
wire n_614;
wire n_529;
wire n_445;
wire n_425;
wire n_684;
wire n_930;
wire n_888;
wire n_1112;
wire n_454;
wire n_218;
wire n_638;
wire n_234;
wire n_910;
wire n_486;
wire n_911;
wire n_381;
wire n_947;
wire n_236;
wire n_653;
wire n_887;
wire n_1087;
wire n_752;
wire n_908;
wire n_944;
wire n_713;
wire n_648;
wire n_657;
wire n_1049;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_239;
wire n_414;
wire n_563;
wire n_782;
wire n_976;
wire n_490;
wire n_803;
wire n_290;
wire n_220;
wire n_809;
wire n_1043;
wire n_1011;
wire n_224;
wire n_926;
wire n_927;
wire n_839;
wire n_986;
wire n_734;
wire n_1088;
wire n_708;
wire n_919;
wire n_1081;
wire n_402;
wire n_352;
wire n_917;
wire n_668;
wire n_478;
wire n_626;
wire n_990;
wire n_574;
wire n_779;
wire n_800;
wire n_929;
wire n_460;
wire n_1084;
wire n_1104;
wire n_907;
wire n_854;
wire n_1058;
wire n_417;
wire n_446;
wire n_498;
wire n_662;
wire n_374;
wire n_659;
wire n_709;
wire n_870;
wire n_366;
wire n_904;
wire n_777;
wire n_407;
wire n_913;
wire n_450;
wire n_808;
wire n_867;
wire n_272;
wire n_526;
wire n_1109;
wire n_921;
wire n_712;
wire n_348;
wire n_711;
wire n_579;
wire n_376;
wire n_937;
wire n_390;
wire n_473;
wire n_293;
wire n_1054;
wire n_334;
wire n_559;
wire n_370;
wire n_458;
wire n_1070;
wire n_1085;
wire n_232;
wire n_650;
wire n_998;
wire n_1046;
wire n_717;
wire n_330;
wire n_771;
wire n_470;
wire n_475;
wire n_924;
wire n_1102;
wire n_298;
wire n_492;
wire n_972;
wire n_281;
wire n_258;
wire n_551;
wire n_699;
wire n_456;
wire n_564;
wire n_260;
wire n_265;
wire n_313;
wire n_451;
wire n_624;
wire n_824;
wire n_962;
wire n_1073;
wire n_1000;
wire n_279;
wire n_686;
wire n_796;
wire n_1041;
wire n_252;
wire n_757;
wire n_228;
wire n_594;
wire n_565;
wire n_719;
wire n_356;
wire n_577;
wire n_936;
wire n_552;
wire n_1062;
wire n_619;
wire n_885;
wire n_216;
wire n_455;
wire n_896;
wire n_521;
wire n_363;
wire n_572;
wire n_912;
wire n_395;
wire n_813;
wire n_592;
wire n_1090;
wire n_745;
wire n_654;
wire n_323;
wire n_829;
wire n_606;
wire n_393;
wire n_818;
wire n_984;
wire n_411;
wire n_503;
wire n_716;
wire n_623;
wire n_1048;
wire n_884;
wire n_599;
wire n_513;
wire n_855;
wire n_776;
wire n_321;
wire n_645;
wire n_331;
wire n_916;
wire n_227;
wire n_1078;
wire n_868;
wire n_570;
wire n_731;
wire n_859;
wire n_406;
wire n_483;
wire n_735;
wire n_482;
wire n_934;
wire n_755;
wire n_1021;
wire n_931;
wire n_474;
wire n_527;
wire n_261;
wire n_608;
wire n_620;
wire n_420;
wire n_683;
wire n_630;
wire n_312;
wire n_394;
wire n_519;
wire n_541;
wire n_512;
wire n_958;
wire n_292;
wire n_307;
wire n_469;
wire n_433;
wire n_500;
wire n_942;
wire n_792;
wire n_880;
wire n_476;
wire n_981;
wire n_714;
wire n_291;
wire n_219;
wire n_543;
wire n_889;
wire n_357;
wire n_264;
wire n_263;
wire n_985;
wire n_589;
wire n_860;
wire n_481;
wire n_788;
wire n_819;
wire n_939;
wire n_997;
wire n_821;
wire n_325;
wire n_938;
wire n_1068;
wire n_767;
wire n_804;
wire n_329;
wire n_464;
wire n_600;
wire n_831;
wire n_802;
wire n_964;
wire n_982;
wire n_561;
wire n_477;
wire n_549;
wire n_980;
wire n_533;
wire n_954;
wire n_1075;
wire n_408;
wire n_932;
wire n_806;
wire n_864;
wire n_879;
wire n_959;
wire n_237;
wire n_584;
wire n_1110;
wire n_244;
wire n_399;
wire n_243;
wire n_979;
wire n_548;
wire n_905;
wire n_282;
wire n_436;
wire n_833;
wire n_211;
wire n_523;
wire n_707;
wire n_322;
wire n_993;
wire n_345;
wire n_409;
wire n_231;
wire n_354;
wire n_689;
wire n_799;
wire n_505;
wire n_240;
wire n_756;
wire n_319;
wire n_547;
wire n_537;
wire n_273;
wire n_558;
wire n_810;
wire n_635;
wire n_787;
wire n_311;
wire n_1064;
wire n_403;
wire n_1080;
wire n_723;
wire n_253;
wire n_634;
wire n_1051;
wire n_583;
wire n_596;
wire n_966;
wire n_546;
wire n_562;
wire n_249;
wire n_386;
wire n_764;
wire n_1039;
wire n_556;
wire n_1034;
wire n_1086;
wire n_1066;
wire n_692;
wire n_733;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_487;
wire n_550;
wire n_241;
wire n_275;
wire n_553;
wire n_652;
wire n_849;
wire n_970;
wire n_1107;
wire n_560;
wire n_1014;
wire n_753;
wire n_642;
wire n_995;
wire n_276;
wire n_569;
wire n_1092;
wire n_441;
wire n_221;
wire n_811;
wire n_1060;
wire n_882;
wire n_444;
wire n_586;
wire n_423;
wire n_737;
wire n_318;
wire n_1111;
wire n_303;
wire n_511;
wire n_715;
wire n_467;
wire n_306;
wire n_269;
wire n_359;
wire n_973;
wire n_346;
wire n_416;
wire n_1053;
wire n_530;
wire n_277;
wire n_520;
wire n_1029;
wire n_418;
wire n_1093;
wire n_618;
wire n_1055;
wire n_790;
wire n_1106;
wire n_582;
wire n_266;
wire n_296;
wire n_861;
wire n_674;
wire n_857;
wire n_871;
wire n_967;
wire n_775;
wire n_922;
wire n_571;
wire n_268;
wire n_271;
wire n_404;
wire n_651;
wire n_439;
wire n_217;
wire n_210;
wire n_299;
wire n_518;
wire n_679;
wire n_1069;
wire n_453;
wire n_612;
wire n_633;
wire n_665;
wire n_902;
wire n_333;
wire n_588;
wire n_215;
wire n_247;
wire n_225;
wire n_308;
wire n_309;
wire n_914;
wire n_759;
wire n_1047;
wire n_1010;
wire n_355;
wire n_426;
wire n_317;
wire n_1040;
wire n_915;
wire n_632;
wire n_702;
wire n_431;
wire n_347;
wire n_812;
wire n_459;
wire n_1052;
wire n_502;
wire n_328;
wire n_672;
wire n_534;
wire n_488;
wire n_429;
wire n_1006;
wire n_373;
wire n_1012;
wire n_497;
wire n_285;
wire n_780;
wire n_773;
wire n_675;
wire n_920;
wire n_257;
wire n_903;
wire n_730;
wire n_655;
wire n_706;
wire n_1045;
wire n_786;
wire n_670;
wire n_286;
wire n_254;
wire n_834;
wire n_242;
wire n_835;
wire n_928;
wire n_690;
wire n_850;
wire n_1089;
wire n_401;
wire n_324;
wire n_743;
wire n_766;
wire n_816;
wire n_335;
wire n_430;
wire n_1002;
wire n_463;
wire n_545;
wire n_489;
wire n_877;
wire n_604;
wire n_848;
wire n_251;
wire n_1019;
wire n_301;
wire n_274;
wire n_636;
wire n_825;
wire n_728;
wire n_681;
wire n_1096;
wire n_1063;
wire n_729;
wire n_1091;
wire n_876;
wire n_774;
wire n_412;
wire n_640;
wire n_660;
wire n_965;
wire n_267;
wire n_438;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_515;
wire n_983;
wire n_288;
wire n_427;
wire n_1059;
wire n_479;
wire n_496;
wire n_598;
wire n_422;
wire n_696;
wire n_906;
wire n_722;
wire n_688;
wire n_1077;
wire n_961;
wire n_862;
wire n_351;
wire n_869;
wire n_437;
wire n_1082;
wire n_259;
wire n_540;
wire n_593;
wire n_514;
wire n_646;
wire n_528;
wire n_457;
wire n_391;
wire n_1098;
wire n_687;
wire n_697;
wire n_364;
wire n_890;
wire n_637;
wire n_295;
wire n_385;
wire n_701;
wire n_817;
wire n_950;
wire n_629;
wire n_388;
wire n_858;
wire n_262;
wire n_484;
wire n_613;
wire n_736;
wire n_897;
wire n_900;
wire n_846;
wire n_501;
wire n_841;
wire n_960;
wire n_956;
wire n_531;
wire n_827;
wire n_1001;
wire n_361;
wire n_508;
wire n_663;
wire n_856;
wire n_1050;
wire n_379;
wire n_778;
wire n_1025;
wire n_332;
wire n_891;
wire n_336;
wire n_398;
wire n_410;
wire n_566;
wire n_554;
wire n_602;
wire n_1013;
wire n_1023;
wire n_1076;
wire n_664;
wire n_949;
wire n_678;
wire n_1007;
wire n_649;
wire n_283;

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_191),
.Y(n_208)
);

INVx1_ASAP7_75t_SL g209 ( 
.A(n_50),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_154),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_183),
.Y(n_211)
);

BUFx6f_ASAP7_75t_L g212 ( 
.A(n_179),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_11),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_145),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_45),
.Y(n_215)
);

INVx1_ASAP7_75t_SL g216 ( 
.A(n_105),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_75),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_35),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_17),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_40),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_119),
.Y(n_221)
);

INVx2_ASAP7_75t_SL g222 ( 
.A(n_100),
.Y(n_222)
);

BUFx6f_ASAP7_75t_L g223 ( 
.A(n_199),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_160),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_60),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_126),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_114),
.Y(n_227)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_120),
.Y(n_228)
);

CKINVDCx14_ASAP7_75t_R g229 ( 
.A(n_167),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_121),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_162),
.Y(n_231)
);

INVx1_ASAP7_75t_SL g232 ( 
.A(n_113),
.Y(n_232)
);

BUFx6f_ASAP7_75t_L g233 ( 
.A(n_152),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_187),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_161),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_9),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_13),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_83),
.Y(n_238)
);

BUFx6f_ASAP7_75t_L g239 ( 
.A(n_200),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_102),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_125),
.Y(n_241)
);

BUFx10_ASAP7_75t_L g242 ( 
.A(n_182),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_22),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_73),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_33),
.Y(n_245)
);

BUFx3_ASAP7_75t_L g246 ( 
.A(n_197),
.Y(n_246)
);

BUFx6f_ASAP7_75t_L g247 ( 
.A(n_131),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_72),
.Y(n_248)
);

INVxp67_ASAP7_75t_L g249 ( 
.A(n_112),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_98),
.Y(n_250)
);

INVx2_ASAP7_75t_SL g251 ( 
.A(n_86),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_173),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_70),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_71),
.Y(n_254)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_30),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_95),
.Y(n_256)
);

INVx1_ASAP7_75t_SL g257 ( 
.A(n_1),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_108),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_2),
.Y(n_259)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_93),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_194),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_118),
.Y(n_262)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_7),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_3),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_156),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_165),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_198),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_27),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_42),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_81),
.Y(n_270)
);

BUFx10_ASAP7_75t_L g271 ( 
.A(n_37),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_205),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_52),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_149),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_157),
.Y(n_275)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_136),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_29),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_243),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_215),
.Y(n_279)
);

INVxp67_ASAP7_75t_SL g280 ( 
.A(n_246),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_214),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_231),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_234),
.Y(n_283)
);

BUFx3_ASAP7_75t_L g284 ( 
.A(n_242),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g285 ( 
.A(n_220),
.Y(n_285)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_255),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_235),
.Y(n_287)
);

BUFx2_ASAP7_75t_SL g288 ( 
.A(n_238),
.Y(n_288)
);

BUFx2_ASAP7_75t_L g289 ( 
.A(n_213),
.Y(n_289)
);

INVxp33_ASAP7_75t_L g290 ( 
.A(n_263),
.Y(n_290)
);

INVxp67_ASAP7_75t_SL g291 ( 
.A(n_249),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_219),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_244),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_270),
.Y(n_294)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_212),
.Y(n_295)
);

INVxp67_ASAP7_75t_SL g296 ( 
.A(n_249),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_236),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g298 ( 
.A(n_273),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_248),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_253),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_258),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_237),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_262),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_259),
.Y(n_304)
);

INVxp67_ASAP7_75t_SL g305 ( 
.A(n_228),
.Y(n_305)
);

INVx2_ASAP7_75t_L g306 ( 
.A(n_212),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_268),
.Y(n_307)
);

INVxp33_ASAP7_75t_SL g308 ( 
.A(n_257),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_260),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_208),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_276),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_210),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_212),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_212),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_223),
.Y(n_315)
);

INVx2_ASAP7_75t_L g316 ( 
.A(n_223),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_223),
.Y(n_317)
);

INVxp67_ASAP7_75t_L g318 ( 
.A(n_242),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_223),
.Y(n_319)
);

INVx1_ASAP7_75t_SL g320 ( 
.A(n_264),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_233),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_211),
.Y(n_322)
);

INVx2_ASAP7_75t_L g323 ( 
.A(n_233),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_217),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_218),
.Y(n_325)
);

BUFx2_ASAP7_75t_SL g326 ( 
.A(n_274),
.Y(n_326)
);

HB1xp67_ASAP7_75t_L g327 ( 
.A(n_277),
.Y(n_327)
);

CKINVDCx16_ASAP7_75t_R g328 ( 
.A(n_229),
.Y(n_328)
);

BUFx6f_ASAP7_75t_L g329 ( 
.A(n_295),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_291),
.B(n_209),
.Y(n_330)
);

AND2x4_ASAP7_75t_L g331 ( 
.A(n_280),
.B(n_222),
.Y(n_331)
);

AOI22xp5_ASAP7_75t_L g332 ( 
.A1(n_308),
.A2(n_292),
.B1(n_302),
.B2(n_297),
.Y(n_332)
);

OA21x2_ASAP7_75t_L g333 ( 
.A1(n_295),
.A2(n_251),
.B(n_224),
.Y(n_333)
);

OAI22xp5_ASAP7_75t_L g334 ( 
.A1(n_308),
.A2(n_216),
.B1(n_232),
.B2(n_275),
.Y(n_334)
);

INVx2_ASAP7_75t_L g335 ( 
.A(n_306),
.Y(n_335)
);

BUFx6f_ASAP7_75t_L g336 ( 
.A(n_306),
.Y(n_336)
);

NOR2x1_ASAP7_75t_L g337 ( 
.A(n_284),
.B(n_233),
.Y(n_337)
);

AND2x4_ASAP7_75t_L g338 ( 
.A(n_284),
.B(n_233),
.Y(n_338)
);

NOR2x1_ASAP7_75t_L g339 ( 
.A(n_313),
.B(n_314),
.Y(n_339)
);

BUFx6f_ASAP7_75t_L g340 ( 
.A(n_316),
.Y(n_340)
);

BUFx6f_ASAP7_75t_L g341 ( 
.A(n_316),
.Y(n_341)
);

INVx2_ASAP7_75t_L g342 ( 
.A(n_323),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_279),
.Y(n_343)
);

OAI22xp5_ASAP7_75t_L g344 ( 
.A1(n_296),
.A2(n_272),
.B1(n_221),
.B2(n_269),
.Y(n_344)
);

BUFx6f_ASAP7_75t_L g345 ( 
.A(n_323),
.Y(n_345)
);

INVx2_ASAP7_75t_L g346 ( 
.A(n_315),
.Y(n_346)
);

NOR2x1_ASAP7_75t_L g347 ( 
.A(n_317),
.B(n_239),
.Y(n_347)
);

INVx6_ASAP7_75t_L g348 ( 
.A(n_328),
.Y(n_348)
);

INVx2_ASAP7_75t_L g349 ( 
.A(n_319),
.Y(n_349)
);

BUFx3_ASAP7_75t_L g350 ( 
.A(n_282),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_283),
.Y(n_351)
);

INVx2_ASAP7_75t_SL g352 ( 
.A(n_292),
.Y(n_352)
);

BUFx6f_ASAP7_75t_L g353 ( 
.A(n_286),
.Y(n_353)
);

AND2x2_ASAP7_75t_L g354 ( 
.A(n_289),
.B(n_271),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_SL g355 ( 
.A(n_318),
.B(n_271),
.Y(n_355)
);

BUFx6f_ASAP7_75t_L g356 ( 
.A(n_286),
.Y(n_356)
);

BUFx6f_ASAP7_75t_L g357 ( 
.A(n_321),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_287),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_305),
.B(n_225),
.Y(n_359)
);

OA21x2_ASAP7_75t_L g360 ( 
.A1(n_293),
.A2(n_227),
.B(n_226),
.Y(n_360)
);

BUFx3_ASAP7_75t_L g361 ( 
.A(n_310),
.Y(n_361)
);

BUFx6f_ASAP7_75t_L g362 ( 
.A(n_278),
.Y(n_362)
);

AND2x4_ASAP7_75t_L g363 ( 
.A(n_289),
.B(n_239),
.Y(n_363)
);

INVxp33_ASAP7_75t_SL g364 ( 
.A(n_310),
.Y(n_364)
);

BUFx6f_ASAP7_75t_L g365 ( 
.A(n_293),
.Y(n_365)
);

NAND2xp33_ASAP7_75t_L g366 ( 
.A(n_303),
.B(n_239),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_299),
.B(n_267),
.Y(n_367)
);

OAI22xp5_ASAP7_75t_SL g368 ( 
.A1(n_320),
.A2(n_266),
.B1(n_265),
.B2(n_261),
.Y(n_368)
);

BUFx2_ASAP7_75t_L g369 ( 
.A(n_297),
.Y(n_369)
);

INVx2_ASAP7_75t_L g370 ( 
.A(n_309),
.Y(n_370)
);

NOR2x1_ASAP7_75t_L g371 ( 
.A(n_303),
.B(n_239),
.Y(n_371)
);

BUFx6f_ASAP7_75t_L g372 ( 
.A(n_311),
.Y(n_372)
);

INVx5_ASAP7_75t_L g373 ( 
.A(n_300),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_301),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_290),
.Y(n_375)
);

OA21x2_ASAP7_75t_L g376 ( 
.A1(n_302),
.A2(n_240),
.B(n_230),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_304),
.Y(n_377)
);

NAND2xp33_ASAP7_75t_L g378 ( 
.A(n_304),
.B(n_247),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_307),
.Y(n_379)
);

AND2x4_ASAP7_75t_L g380 ( 
.A(n_312),
.B(n_247),
.Y(n_380)
);

INVx2_ASAP7_75t_L g381 ( 
.A(n_312),
.Y(n_381)
);

INVx3_ASAP7_75t_L g382 ( 
.A(n_322),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_322),
.B(n_241),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_365),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_365),
.Y(n_385)
);

INVx5_ASAP7_75t_L g386 ( 
.A(n_329),
.Y(n_386)
);

INVxp67_ASAP7_75t_SL g387 ( 
.A(n_329),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_365),
.Y(n_388)
);

INVx2_ASAP7_75t_L g389 ( 
.A(n_335),
.Y(n_389)
);

INVx5_ASAP7_75t_L g390 ( 
.A(n_329),
.Y(n_390)
);

INVx2_ASAP7_75t_L g391 ( 
.A(n_342),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_365),
.Y(n_392)
);

INVx2_ASAP7_75t_L g393 ( 
.A(n_353),
.Y(n_393)
);

INVx2_ASAP7_75t_L g394 ( 
.A(n_353),
.Y(n_394)
);

AND3x2_ASAP7_75t_L g395 ( 
.A(n_369),
.B(n_327),
.C(n_326),
.Y(n_395)
);

INVx2_ASAP7_75t_L g396 ( 
.A(n_353),
.Y(n_396)
);

INVx2_ASAP7_75t_SL g397 ( 
.A(n_375),
.Y(n_397)
);

INVx2_ASAP7_75t_L g398 ( 
.A(n_353),
.Y(n_398)
);

INVx2_ASAP7_75t_L g399 ( 
.A(n_356),
.Y(n_399)
);

INVx2_ASAP7_75t_L g400 ( 
.A(n_356),
.Y(n_400)
);

AND2x2_ASAP7_75t_L g401 ( 
.A(n_363),
.B(n_307),
.Y(n_401)
);

INVx2_ASAP7_75t_L g402 ( 
.A(n_356),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_356),
.Y(n_403)
);

INVx2_ASAP7_75t_L g404 ( 
.A(n_329),
.Y(n_404)
);

NAND2xp33_ASAP7_75t_SL g405 ( 
.A(n_354),
.B(n_324),
.Y(n_405)
);

AND2x2_ASAP7_75t_L g406 ( 
.A(n_363),
.B(n_324),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_346),
.Y(n_407)
);

INVx2_ASAP7_75t_L g408 ( 
.A(n_336),
.Y(n_408)
);

OR2x6_ASAP7_75t_L g409 ( 
.A(n_381),
.B(n_288),
.Y(n_409)
);

INVx2_ASAP7_75t_L g410 ( 
.A(n_336),
.Y(n_410)
);

INVx2_ASAP7_75t_L g411 ( 
.A(n_336),
.Y(n_411)
);

INVx2_ASAP7_75t_L g412 ( 
.A(n_336),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_349),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_SL g414 ( 
.A(n_330),
.B(n_325),
.Y(n_414)
);

AND3x2_ASAP7_75t_L g415 ( 
.A(n_330),
.B(n_326),
.C(n_288),
.Y(n_415)
);

INVx2_ASAP7_75t_L g416 ( 
.A(n_340),
.Y(n_416)
);

INVx2_ASAP7_75t_L g417 ( 
.A(n_340),
.Y(n_417)
);

NOR2xp33_ASAP7_75t_L g418 ( 
.A(n_383),
.B(n_325),
.Y(n_418)
);

INVx2_ASAP7_75t_L g419 ( 
.A(n_340),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_380),
.B(n_245),
.Y(n_420)
);

CKINVDCx6p67_ASAP7_75t_R g421 ( 
.A(n_361),
.Y(n_421)
);

AOI22xp5_ASAP7_75t_L g422 ( 
.A1(n_334),
.A2(n_298),
.B1(n_294),
.B2(n_285),
.Y(n_422)
);

INVx3_ASAP7_75t_L g423 ( 
.A(n_340),
.Y(n_423)
);

INVx2_ASAP7_75t_L g424 ( 
.A(n_341),
.Y(n_424)
);

INVx2_ASAP7_75t_L g425 ( 
.A(n_341),
.Y(n_425)
);

INVx2_ASAP7_75t_L g426 ( 
.A(n_341),
.Y(n_426)
);

NOR2xp33_ASAP7_75t_L g427 ( 
.A(n_383),
.B(n_281),
.Y(n_427)
);

BUFx6f_ASAP7_75t_L g428 ( 
.A(n_341),
.Y(n_428)
);

AND3x2_ASAP7_75t_L g429 ( 
.A(n_377),
.B(n_0),
.C(n_1),
.Y(n_429)
);

INVx2_ASAP7_75t_L g430 ( 
.A(n_345),
.Y(n_430)
);

INVx2_ASAP7_75t_L g431 ( 
.A(n_345),
.Y(n_431)
);

NOR2xp33_ASAP7_75t_L g432 ( 
.A(n_379),
.B(n_256),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_SL g433 ( 
.A(n_380),
.B(n_332),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_362),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_362),
.Y(n_435)
);

BUFx3_ASAP7_75t_L g436 ( 
.A(n_350),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_362),
.Y(n_437)
);

INVx1_ASAP7_75t_SL g438 ( 
.A(n_348),
.Y(n_438)
);

INVx2_ASAP7_75t_SL g439 ( 
.A(n_338),
.Y(n_439)
);

INVx2_ASAP7_75t_L g440 ( 
.A(n_345),
.Y(n_440)
);

INVx2_ASAP7_75t_L g441 ( 
.A(n_345),
.Y(n_441)
);

BUFx2_ASAP7_75t_L g442 ( 
.A(n_338),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_362),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g444 ( 
.A(n_359),
.B(n_250),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_SL g445 ( 
.A(n_382),
.B(n_254),
.Y(n_445)
);

INVx3_ASAP7_75t_L g446 ( 
.A(n_357),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_343),
.Y(n_447)
);

INVx2_ASAP7_75t_L g448 ( 
.A(n_357),
.Y(n_448)
);

INVx4_ASAP7_75t_L g449 ( 
.A(n_357),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_351),
.Y(n_450)
);

INVx2_ASAP7_75t_L g451 ( 
.A(n_357),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_358),
.Y(n_452)
);

CKINVDCx6p67_ASAP7_75t_R g453 ( 
.A(n_355),
.Y(n_453)
);

INVx2_ASAP7_75t_L g454 ( 
.A(n_370),
.Y(n_454)
);

INVx2_ASAP7_75t_SL g455 ( 
.A(n_331),
.Y(n_455)
);

BUFx6f_ASAP7_75t_L g456 ( 
.A(n_372),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_374),
.Y(n_457)
);

NOR2xp33_ASAP7_75t_L g458 ( 
.A(n_359),
.B(n_252),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_447),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_447),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_450),
.Y(n_461)
);

AND2x4_ASAP7_75t_L g462 ( 
.A(n_439),
.B(n_350),
.Y(n_462)
);

CKINVDCx20_ASAP7_75t_R g463 ( 
.A(n_421),
.Y(n_463)
);

AND2x2_ASAP7_75t_L g464 ( 
.A(n_397),
.B(n_382),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_450),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_452),
.Y(n_466)
);

BUFx6f_ASAP7_75t_L g467 ( 
.A(n_436),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_452),
.Y(n_468)
);

BUFx6f_ASAP7_75t_L g469 ( 
.A(n_436),
.Y(n_469)
);

CKINVDCx5p33_ASAP7_75t_R g470 ( 
.A(n_421),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_457),
.Y(n_471)
);

BUFx6f_ASAP7_75t_L g472 ( 
.A(n_442),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_457),
.Y(n_473)
);

CKINVDCx20_ASAP7_75t_R g474 ( 
.A(n_422),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_454),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_407),
.Y(n_476)
);

AND2x4_ASAP7_75t_L g477 ( 
.A(n_439),
.B(n_337),
.Y(n_477)
);

HB1xp67_ASAP7_75t_L g478 ( 
.A(n_401),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_413),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_413),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_L g481 ( 
.A(n_458),
.B(n_331),
.Y(n_481)
);

CKINVDCx20_ASAP7_75t_R g482 ( 
.A(n_422),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_389),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_391),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_391),
.Y(n_485)
);

BUFx6f_ASAP7_75t_L g486 ( 
.A(n_442),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_397),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_455),
.Y(n_488)
);

BUFx6f_ASAP7_75t_L g489 ( 
.A(n_456),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_455),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_434),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_434),
.Y(n_492)
);

NOR2xp33_ASAP7_75t_L g493 ( 
.A(n_418),
.B(n_364),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_435),
.Y(n_494)
);

XNOR2x2_ASAP7_75t_L g495 ( 
.A(n_414),
.B(n_334),
.Y(n_495)
);

CKINVDCx20_ASAP7_75t_R g496 ( 
.A(n_405),
.Y(n_496)
);

AND2x2_ASAP7_75t_L g497 ( 
.A(n_401),
.B(n_406),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_435),
.Y(n_498)
);

NAND2x1p5_ASAP7_75t_L g499 ( 
.A(n_438),
.B(n_333),
.Y(n_499)
);

NOR2xp33_ASAP7_75t_L g500 ( 
.A(n_432),
.B(n_352),
.Y(n_500)
);

AND2x2_ASAP7_75t_L g501 ( 
.A(n_406),
.B(n_427),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_437),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_437),
.Y(n_503)
);

AND2x2_ASAP7_75t_L g504 ( 
.A(n_409),
.B(n_348),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_443),
.Y(n_505)
);

CKINVDCx5p33_ASAP7_75t_R g506 ( 
.A(n_453),
.Y(n_506)
);

AND2x2_ASAP7_75t_L g507 ( 
.A(n_409),
.B(n_348),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_443),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_384),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_385),
.Y(n_510)
);

BUFx6f_ASAP7_75t_L g511 ( 
.A(n_456),
.Y(n_511)
);

INVx2_ASAP7_75t_L g512 ( 
.A(n_428),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_385),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_388),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_388),
.Y(n_515)
);

OR2x6_ASAP7_75t_L g516 ( 
.A(n_409),
.B(n_368),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_392),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_392),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_393),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_393),
.Y(n_520)
);

OAI21xp5_ASAP7_75t_L g521 ( 
.A1(n_444),
.A2(n_360),
.B(n_333),
.Y(n_521)
);

CKINVDCx20_ASAP7_75t_R g522 ( 
.A(n_453),
.Y(n_522)
);

INVxp67_ASAP7_75t_SL g523 ( 
.A(n_428),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_394),
.Y(n_524)
);

AND2x2_ASAP7_75t_L g525 ( 
.A(n_409),
.B(n_355),
.Y(n_525)
);

CKINVDCx20_ASAP7_75t_R g526 ( 
.A(n_433),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_394),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_396),
.Y(n_528)
);

NOR2xp33_ASAP7_75t_L g529 ( 
.A(n_445),
.B(n_344),
.Y(n_529)
);

INVx4_ASAP7_75t_L g530 ( 
.A(n_456),
.Y(n_530)
);

BUFx6f_ASAP7_75t_SL g531 ( 
.A(n_395),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_396),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_398),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_398),
.Y(n_534)
);

CKINVDCx5p33_ASAP7_75t_R g535 ( 
.A(n_420),
.Y(n_535)
);

XNOR2xp5_ASAP7_75t_L g536 ( 
.A(n_415),
.B(n_376),
.Y(n_536)
);

XOR2xp5_ASAP7_75t_L g537 ( 
.A(n_403),
.B(n_376),
.Y(n_537)
);

AND2x2_ASAP7_75t_L g538 ( 
.A(n_399),
.B(n_344),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_399),
.Y(n_539)
);

NOR2xp33_ASAP7_75t_L g540 ( 
.A(n_493),
.B(n_367),
.Y(n_540)
);

NOR2xp33_ASAP7_75t_L g541 ( 
.A(n_501),
.B(n_481),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_L g542 ( 
.A(n_481),
.B(n_500),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_L g543 ( 
.A(n_464),
.B(n_459),
.Y(n_543)
);

CKINVDCx5p33_ASAP7_75t_R g544 ( 
.A(n_470),
.Y(n_544)
);

NOR2xp33_ASAP7_75t_L g545 ( 
.A(n_478),
.B(n_367),
.Y(n_545)
);

INVxp33_ASAP7_75t_L g546 ( 
.A(n_497),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_SL g547 ( 
.A(n_535),
.B(n_456),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_L g548 ( 
.A(n_460),
.B(n_360),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_483),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_SL g550 ( 
.A(n_472),
.B(n_456),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_484),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_L g552 ( 
.A(n_461),
.B(n_403),
.Y(n_552)
);

OAI22xp5_ASAP7_75t_L g553 ( 
.A1(n_529),
.A2(n_402),
.B1(n_400),
.B2(n_404),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_L g554 ( 
.A(n_465),
.B(n_400),
.Y(n_554)
);

BUFx3_ASAP7_75t_L g555 ( 
.A(n_467),
.Y(n_555)
);

AND2x2_ASAP7_75t_SL g556 ( 
.A(n_525),
.B(n_378),
.Y(n_556)
);

AND2x6_ASAP7_75t_SL g557 ( 
.A(n_516),
.B(n_429),
.Y(n_557)
);

NOR3xp33_ASAP7_75t_L g558 ( 
.A(n_538),
.B(n_378),
.C(n_366),
.Y(n_558)
);

INVx2_ASAP7_75t_SL g559 ( 
.A(n_487),
.Y(n_559)
);

NOR2xp33_ASAP7_75t_L g560 ( 
.A(n_495),
.B(n_402),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_L g561 ( 
.A(n_466),
.B(n_446),
.Y(n_561)
);

NOR2xp33_ASAP7_75t_L g562 ( 
.A(n_488),
.B(n_423),
.Y(n_562)
);

NOR2xp33_ASAP7_75t_L g563 ( 
.A(n_490),
.B(n_423),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_L g564 ( 
.A(n_468),
.B(n_446),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_L g565 ( 
.A(n_471),
.B(n_446),
.Y(n_565)
);

AOI22xp33_ASAP7_75t_L g566 ( 
.A1(n_473),
.A2(n_247),
.B1(n_408),
.B2(n_404),
.Y(n_566)
);

NOR2xp33_ASAP7_75t_L g567 ( 
.A(n_472),
.B(n_423),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_SL g568 ( 
.A(n_472),
.B(n_448),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_L g569 ( 
.A(n_462),
.B(n_408),
.Y(n_569)
);

INVxp67_ASAP7_75t_SL g570 ( 
.A(n_489),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_485),
.Y(n_571)
);

AND2x2_ASAP7_75t_L g572 ( 
.A(n_486),
.B(n_372),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_SL g573 ( 
.A(n_486),
.B(n_462),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_L g574 ( 
.A(n_477),
.B(n_410),
.Y(n_574)
);

BUFx6f_ASAP7_75t_L g575 ( 
.A(n_489),
.Y(n_575)
);

INVx3_ASAP7_75t_L g576 ( 
.A(n_512),
.Y(n_576)
);

NOR2xp33_ASAP7_75t_L g577 ( 
.A(n_486),
.B(n_526),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_SL g578 ( 
.A(n_477),
.B(n_448),
.Y(n_578)
);

INVx2_ASAP7_75t_L g579 ( 
.A(n_475),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_L g580 ( 
.A(n_476),
.B(n_410),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_479),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_480),
.Y(n_582)
);

AOI22xp5_ASAP7_75t_L g583 ( 
.A1(n_537),
.A2(n_387),
.B1(n_451),
.B2(n_441),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_509),
.Y(n_584)
);

NAND2xp5_ASAP7_75t_SL g585 ( 
.A(n_467),
.B(n_451),
.Y(n_585)
);

INVx5_ASAP7_75t_L g586 ( 
.A(n_489),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_510),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_513),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_514),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_SL g590 ( 
.A(n_467),
.B(n_372),
.Y(n_590)
);

INVx3_ASAP7_75t_L g591 ( 
.A(n_511),
.Y(n_591)
);

INVx3_ASAP7_75t_L g592 ( 
.A(n_511),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_515),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_L g594 ( 
.A(n_517),
.B(n_411),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_L g595 ( 
.A(n_518),
.B(n_412),
.Y(n_595)
);

OAI21xp5_ASAP7_75t_L g596 ( 
.A1(n_521),
.A2(n_416),
.B(n_412),
.Y(n_596)
);

AND2x2_ASAP7_75t_L g597 ( 
.A(n_504),
.B(n_372),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_L g598 ( 
.A(n_491),
.B(n_416),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_SL g599 ( 
.A(n_469),
.B(n_428),
.Y(n_599)
);

AND2x2_ASAP7_75t_L g600 ( 
.A(n_507),
.B(n_371),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_492),
.Y(n_601)
);

AND2x2_ASAP7_75t_L g602 ( 
.A(n_469),
.B(n_339),
.Y(n_602)
);

AND2x4_ASAP7_75t_SL g603 ( 
.A(n_463),
.B(n_417),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_L g604 ( 
.A(n_494),
.B(n_417),
.Y(n_604)
);

AND2x4_ASAP7_75t_L g605 ( 
.A(n_555),
.B(n_516),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_L g606 ( 
.A(n_542),
.B(n_499),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_554),
.Y(n_607)
);

BUFx8_ASAP7_75t_L g608 ( 
.A(n_602),
.Y(n_608)
);

BUFx4f_ASAP7_75t_SL g609 ( 
.A(n_573),
.Y(n_609)
);

NOR2xp33_ASAP7_75t_R g610 ( 
.A(n_544),
.B(n_506),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_SL g611 ( 
.A(n_541),
.B(n_536),
.Y(n_611)
);

INVx3_ASAP7_75t_L g612 ( 
.A(n_575),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_594),
.Y(n_613)
);

A2O1A1Ixp33_ASAP7_75t_L g614 ( 
.A1(n_540),
.A2(n_521),
.B(n_498),
.C(n_503),
.Y(n_614)
);

INVx2_ASAP7_75t_SL g615 ( 
.A(n_603),
.Y(n_615)
);

AOI22xp33_ASAP7_75t_L g616 ( 
.A1(n_540),
.A2(n_474),
.B1(n_482),
.B2(n_516),
.Y(n_616)
);

NOR2xp67_ASAP7_75t_L g617 ( 
.A(n_577),
.B(n_545),
.Y(n_617)
);

INVx3_ASAP7_75t_SL g618 ( 
.A(n_556),
.Y(n_618)
);

INVx2_ASAP7_75t_L g619 ( 
.A(n_579),
.Y(n_619)
);

NOR2xp33_ASAP7_75t_L g620 ( 
.A(n_546),
.B(n_522),
.Y(n_620)
);

NOR2xp33_ASAP7_75t_R g621 ( 
.A(n_556),
.B(n_496),
.Y(n_621)
);

NOR2xp33_ASAP7_75t_L g622 ( 
.A(n_541),
.B(n_499),
.Y(n_622)
);

NAND3xp33_ASAP7_75t_SL g623 ( 
.A(n_545),
.B(n_505),
.C(n_502),
.Y(n_623)
);

BUFx3_ASAP7_75t_L g624 ( 
.A(n_577),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_581),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_582),
.Y(n_626)
);

NOR2xp33_ASAP7_75t_R g627 ( 
.A(n_560),
.B(n_531),
.Y(n_627)
);

BUFx6f_ASAP7_75t_L g628 ( 
.A(n_575),
.Y(n_628)
);

BUFx10_ASAP7_75t_L g629 ( 
.A(n_557),
.Y(n_629)
);

BUFx12f_ASAP7_75t_L g630 ( 
.A(n_559),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_SL g631 ( 
.A(n_543),
.B(n_511),
.Y(n_631)
);

BUFx2_ASAP7_75t_L g632 ( 
.A(n_572),
.Y(n_632)
);

OR2x6_ASAP7_75t_L g633 ( 
.A(n_600),
.B(n_508),
.Y(n_633)
);

BUFx6f_ASAP7_75t_L g634 ( 
.A(n_575),
.Y(n_634)
);

BUFx6f_ASAP7_75t_L g635 ( 
.A(n_575),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_595),
.Y(n_636)
);

INVx3_ASAP7_75t_L g637 ( 
.A(n_591),
.Y(n_637)
);

INVx2_ASAP7_75t_L g638 ( 
.A(n_584),
.Y(n_638)
);

OR2x6_ASAP7_75t_L g639 ( 
.A(n_597),
.B(n_519),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_L g640 ( 
.A(n_560),
.B(n_523),
.Y(n_640)
);

AOI211xp5_ASAP7_75t_L g641 ( 
.A1(n_558),
.A2(n_366),
.B(n_247),
.C(n_533),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_598),
.Y(n_642)
);

NAND2xp33_ASAP7_75t_SL g643 ( 
.A(n_547),
.B(n_531),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_604),
.Y(n_644)
);

INVx4_ASAP7_75t_L g645 ( 
.A(n_586),
.Y(n_645)
);

BUFx2_ASAP7_75t_L g646 ( 
.A(n_587),
.Y(n_646)
);

INVx2_ASAP7_75t_L g647 ( 
.A(n_588),
.Y(n_647)
);

AND2x2_ASAP7_75t_L g648 ( 
.A(n_589),
.B(n_539),
.Y(n_648)
);

CKINVDCx20_ASAP7_75t_R g649 ( 
.A(n_583),
.Y(n_649)
);

HB1xp67_ASAP7_75t_L g650 ( 
.A(n_567),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_L g651 ( 
.A(n_593),
.B(n_601),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_L g652 ( 
.A(n_574),
.B(n_520),
.Y(n_652)
);

INVx5_ASAP7_75t_L g653 ( 
.A(n_586),
.Y(n_653)
);

NOR2xp67_ASAP7_75t_L g654 ( 
.A(n_549),
.B(n_551),
.Y(n_654)
);

INVx2_ASAP7_75t_L g655 ( 
.A(n_571),
.Y(n_655)
);

NOR2xp33_ASAP7_75t_R g656 ( 
.A(n_591),
.B(n_534),
.Y(n_656)
);

NOR2xp33_ASAP7_75t_L g657 ( 
.A(n_569),
.B(n_524),
.Y(n_657)
);

NOR3xp33_ASAP7_75t_SL g658 ( 
.A(n_550),
.B(n_528),
.C(n_527),
.Y(n_658)
);

NOR3xp33_ASAP7_75t_SL g659 ( 
.A(n_567),
.B(n_532),
.C(n_0),
.Y(n_659)
);

CKINVDCx6p67_ASAP7_75t_R g660 ( 
.A(n_586),
.Y(n_660)
);

INVx5_ASAP7_75t_L g661 ( 
.A(n_586),
.Y(n_661)
);

BUFx6f_ASAP7_75t_L g662 ( 
.A(n_592),
.Y(n_662)
);

INVx2_ASAP7_75t_L g663 ( 
.A(n_576),
.Y(n_663)
);

AOI22xp5_ASAP7_75t_L g664 ( 
.A1(n_558),
.A2(n_530),
.B1(n_425),
.B2(n_441),
.Y(n_664)
);

BUFx6f_ASAP7_75t_L g665 ( 
.A(n_592),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_L g666 ( 
.A(n_552),
.B(n_530),
.Y(n_666)
);

NOR2xp33_ASAP7_75t_R g667 ( 
.A(n_576),
.B(n_31),
.Y(n_667)
);

AND2x2_ASAP7_75t_L g668 ( 
.A(n_578),
.B(n_373),
.Y(n_668)
);

OAI21xp5_ASAP7_75t_L g669 ( 
.A1(n_614),
.A2(n_548),
.B(n_596),
.Y(n_669)
);

AOI21xp33_ASAP7_75t_L g670 ( 
.A1(n_616),
.A2(n_564),
.B(n_561),
.Y(n_670)
);

AOI21xp5_ASAP7_75t_SL g671 ( 
.A1(n_640),
.A2(n_570),
.B(n_553),
.Y(n_671)
);

O2A1O1Ixp5_ASAP7_75t_L g672 ( 
.A1(n_611),
.A2(n_568),
.B(n_563),
.C(n_562),
.Y(n_672)
);

NAND2x1p5_ASAP7_75t_L g673 ( 
.A(n_653),
.B(n_599),
.Y(n_673)
);

AO31x2_ASAP7_75t_L g674 ( 
.A1(n_622),
.A2(n_562),
.A3(n_563),
.B(n_565),
.Y(n_674)
);

CKINVDCx20_ASAP7_75t_R g675 ( 
.A(n_610),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_625),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_L g677 ( 
.A(n_617),
.B(n_607),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_L g678 ( 
.A(n_607),
.B(n_570),
.Y(n_678)
);

AND2x4_ASAP7_75t_L g679 ( 
.A(n_633),
.B(n_585),
.Y(n_679)
);

OAI21x1_ASAP7_75t_L g680 ( 
.A1(n_664),
.A2(n_580),
.B(n_590),
.Y(n_680)
);

OAI22x1_ASAP7_75t_L g681 ( 
.A1(n_618),
.A2(n_419),
.B1(n_424),
.B2(n_425),
.Y(n_681)
);

INVx2_ASAP7_75t_L g682 ( 
.A(n_638),
.Y(n_682)
);

AOI21x1_ASAP7_75t_L g683 ( 
.A1(n_606),
.A2(n_424),
.B(n_419),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_613),
.B(n_566),
.Y(n_684)
);

AOI21xp5_ASAP7_75t_L g685 ( 
.A1(n_653),
.A2(n_566),
.B(n_449),
.Y(n_685)
);

OAI21x1_ASAP7_75t_L g686 ( 
.A1(n_631),
.A2(n_430),
.B(n_426),
.Y(n_686)
);

BUFx3_ASAP7_75t_L g687 ( 
.A(n_630),
.Y(n_687)
);

AND2x2_ASAP7_75t_L g688 ( 
.A(n_624),
.B(n_373),
.Y(n_688)
);

AOI21x1_ASAP7_75t_SL g689 ( 
.A1(n_666),
.A2(n_652),
.B(n_650),
.Y(n_689)
);

OAI21xp5_ASAP7_75t_L g690 ( 
.A1(n_641),
.A2(n_657),
.B(n_636),
.Y(n_690)
);

INVx2_ASAP7_75t_L g691 ( 
.A(n_647),
.Y(n_691)
);

AOI21xp5_ASAP7_75t_L g692 ( 
.A1(n_661),
.A2(n_449),
.B(n_390),
.Y(n_692)
);

OAI21xp5_ASAP7_75t_L g693 ( 
.A1(n_636),
.A2(n_440),
.B(n_431),
.Y(n_693)
);

INVx5_ASAP7_75t_L g694 ( 
.A(n_661),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_L g695 ( 
.A(n_642),
.B(n_431),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_L g696 ( 
.A(n_642),
.B(n_644),
.Y(n_696)
);

OAI21xp33_ASAP7_75t_L g697 ( 
.A1(n_627),
.A2(n_347),
.B(n_440),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_L g698 ( 
.A(n_644),
.B(n_632),
.Y(n_698)
);

OAI21xp5_ASAP7_75t_L g699 ( 
.A1(n_623),
.A2(n_449),
.B(n_390),
.Y(n_699)
);

INVx3_ASAP7_75t_L g700 ( 
.A(n_645),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_L g701 ( 
.A(n_651),
.B(n_373),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_626),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_L g703 ( 
.A(n_646),
.B(n_373),
.Y(n_703)
);

NOR2xp33_ASAP7_75t_L g704 ( 
.A(n_649),
.B(n_2),
.Y(n_704)
);

AOI21xp5_ASAP7_75t_L g705 ( 
.A1(n_661),
.A2(n_390),
.B(n_386),
.Y(n_705)
);

CKINVDCx5p33_ASAP7_75t_R g706 ( 
.A(n_608),
.Y(n_706)
);

OAI21x1_ASAP7_75t_L g707 ( 
.A1(n_637),
.A2(n_386),
.B(n_390),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_L g708 ( 
.A(n_655),
.B(n_3),
.Y(n_708)
);

HB1xp67_ASAP7_75t_L g709 ( 
.A(n_633),
.Y(n_709)
);

A2O1A1Ixp33_ASAP7_75t_L g710 ( 
.A1(n_654),
.A2(n_390),
.B(n_386),
.C(n_6),
.Y(n_710)
);

OAI21x1_ASAP7_75t_L g711 ( 
.A1(n_637),
.A2(n_386),
.B(n_34),
.Y(n_711)
);

OAI21xp5_ASAP7_75t_L g712 ( 
.A1(n_658),
.A2(n_386),
.B(n_36),
.Y(n_712)
);

AOI21xp5_ASAP7_75t_L g713 ( 
.A1(n_645),
.A2(n_38),
.B(n_32),
.Y(n_713)
);

BUFx3_ASAP7_75t_L g714 ( 
.A(n_608),
.Y(n_714)
);

INVx2_ASAP7_75t_L g715 ( 
.A(n_648),
.Y(n_715)
);

AOI21xp5_ASAP7_75t_L g716 ( 
.A1(n_639),
.A2(n_41),
.B(n_39),
.Y(n_716)
);

NOR2xp33_ASAP7_75t_R g717 ( 
.A(n_643),
.B(n_43),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_619),
.Y(n_718)
);

BUFx6f_ASAP7_75t_L g719 ( 
.A(n_628),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_663),
.Y(n_720)
);

NOR2xp33_ASAP7_75t_R g721 ( 
.A(n_615),
.B(n_44),
.Y(n_721)
);

OAI22xp5_ASAP7_75t_L g722 ( 
.A1(n_609),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_722)
);

AND2x2_ASAP7_75t_L g723 ( 
.A(n_605),
.B(n_4),
.Y(n_723)
);

OAI21x1_ASAP7_75t_L g724 ( 
.A1(n_612),
.A2(n_47),
.B(n_46),
.Y(n_724)
);

OAI21x1_ASAP7_75t_L g725 ( 
.A1(n_612),
.A2(n_49),
.B(n_48),
.Y(n_725)
);

OAI21x1_ASAP7_75t_L g726 ( 
.A1(n_668),
.A2(n_53),
.B(n_51),
.Y(n_726)
);

INVx5_ASAP7_75t_L g727 ( 
.A(n_628),
.Y(n_727)
);

OAI22xp5_ASAP7_75t_L g728 ( 
.A1(n_605),
.A2(n_5),
.B1(n_7),
.B2(n_8),
.Y(n_728)
);

AO31x2_ASAP7_75t_L g729 ( 
.A1(n_681),
.A2(n_659),
.A3(n_620),
.B(n_667),
.Y(n_729)
);

AOI21xp5_ASAP7_75t_L g730 ( 
.A1(n_671),
.A2(n_634),
.B(n_628),
.Y(n_730)
);

AO32x2_ASAP7_75t_L g731 ( 
.A1(n_728),
.A2(n_621),
.A3(n_629),
.B1(n_656),
.B2(n_11),
.Y(n_731)
);

AOI21xp33_ASAP7_75t_L g732 ( 
.A1(n_690),
.A2(n_665),
.B(n_662),
.Y(n_732)
);

BUFx10_ASAP7_75t_L g733 ( 
.A(n_706),
.Y(n_733)
);

O2A1O1Ixp33_ASAP7_75t_L g734 ( 
.A1(n_722),
.A2(n_629),
.B(n_9),
.C(n_10),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_676),
.Y(n_735)
);

INVx3_ASAP7_75t_L g736 ( 
.A(n_719),
.Y(n_736)
);

NAND2x1p5_ASAP7_75t_L g737 ( 
.A(n_694),
.B(n_727),
.Y(n_737)
);

NOR2xp67_ASAP7_75t_L g738 ( 
.A(n_694),
.B(n_662),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_L g739 ( 
.A(n_696),
.B(n_662),
.Y(n_739)
);

AOI21xp5_ASAP7_75t_L g740 ( 
.A1(n_669),
.A2(n_635),
.B(n_634),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_L g741 ( 
.A(n_715),
.B(n_665),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_L g742 ( 
.A(n_677),
.B(n_665),
.Y(n_742)
);

INVx2_ASAP7_75t_L g743 ( 
.A(n_682),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_702),
.Y(n_744)
);

NOR2xp33_ASAP7_75t_L g745 ( 
.A(n_704),
.B(n_634),
.Y(n_745)
);

AOI21xp5_ASAP7_75t_L g746 ( 
.A1(n_669),
.A2(n_635),
.B(n_660),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_691),
.Y(n_747)
);

AND2x2_ASAP7_75t_L g748 ( 
.A(n_723),
.B(n_635),
.Y(n_748)
);

AO31x2_ASAP7_75t_L g749 ( 
.A1(n_710),
.A2(n_115),
.A3(n_206),
.B(n_204),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_718),
.Y(n_750)
);

NAND3xp33_ASAP7_75t_SL g751 ( 
.A(n_717),
.B(n_8),
.C(n_10),
.Y(n_751)
);

AOI21xp5_ASAP7_75t_L g752 ( 
.A1(n_690),
.A2(n_207),
.B(n_55),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_L g753 ( 
.A(n_698),
.B(n_12),
.Y(n_753)
);

BUFx3_ASAP7_75t_L g754 ( 
.A(n_675),
.Y(n_754)
);

AND2x2_ASAP7_75t_L g755 ( 
.A(n_688),
.B(n_12),
.Y(n_755)
);

OAI22xp5_ASAP7_75t_L g756 ( 
.A1(n_678),
.A2(n_13),
.B1(n_14),
.B2(n_15),
.Y(n_756)
);

A2O1A1Ixp33_ASAP7_75t_L g757 ( 
.A1(n_670),
.A2(n_14),
.B(n_15),
.C(n_16),
.Y(n_757)
);

INVxp67_ASAP7_75t_L g758 ( 
.A(n_709),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_720),
.Y(n_759)
);

AND2x2_ASAP7_75t_L g760 ( 
.A(n_679),
.B(n_16),
.Y(n_760)
);

AOI221xp5_ASAP7_75t_L g761 ( 
.A1(n_728),
.A2(n_17),
.B1(n_18),
.B2(n_19),
.C(n_20),
.Y(n_761)
);

OR2x6_ASAP7_75t_L g762 ( 
.A(n_714),
.B(n_54),
.Y(n_762)
);

BUFx6f_ASAP7_75t_L g763 ( 
.A(n_719),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_708),
.Y(n_764)
);

AOI21xp5_ASAP7_75t_L g765 ( 
.A1(n_685),
.A2(n_117),
.B(n_202),
.Y(n_765)
);

AOI21xp5_ASAP7_75t_L g766 ( 
.A1(n_684),
.A2(n_116),
.B(n_201),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_695),
.Y(n_767)
);

AOI21xp5_ASAP7_75t_L g768 ( 
.A1(n_699),
.A2(n_693),
.B(n_712),
.Y(n_768)
);

O2A1O1Ixp33_ASAP7_75t_SL g769 ( 
.A1(n_712),
.A2(n_18),
.B(n_19),
.C(n_20),
.Y(n_769)
);

INVx3_ASAP7_75t_SL g770 ( 
.A(n_687),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_SL g771 ( 
.A(n_694),
.B(n_21),
.Y(n_771)
);

AOI21xp5_ASAP7_75t_L g772 ( 
.A1(n_672),
.A2(n_203),
.B(n_122),
.Y(n_772)
);

AO31x2_ASAP7_75t_L g773 ( 
.A1(n_692),
.A2(n_713),
.A3(n_716),
.B(n_705),
.Y(n_773)
);

AO31x2_ASAP7_75t_L g774 ( 
.A1(n_701),
.A2(n_111),
.A3(n_195),
.B(n_193),
.Y(n_774)
);

BUFx10_ASAP7_75t_L g775 ( 
.A(n_719),
.Y(n_775)
);

AOI21xp5_ASAP7_75t_L g776 ( 
.A1(n_680),
.A2(n_110),
.B(n_192),
.Y(n_776)
);

O2A1O1Ixp33_ASAP7_75t_L g777 ( 
.A1(n_703),
.A2(n_21),
.B(n_22),
.C(n_23),
.Y(n_777)
);

AO32x2_ASAP7_75t_L g778 ( 
.A1(n_689),
.A2(n_23),
.A3(n_24),
.B1(n_25),
.B2(n_26),
.Y(n_778)
);

AOI21xp5_ASAP7_75t_L g779 ( 
.A1(n_711),
.A2(n_196),
.B(n_123),
.Y(n_779)
);

AOI21xp5_ASAP7_75t_L g780 ( 
.A1(n_726),
.A2(n_697),
.B(n_707),
.Y(n_780)
);

BUFx4f_ASAP7_75t_L g781 ( 
.A(n_673),
.Y(n_781)
);

INVx3_ASAP7_75t_L g782 ( 
.A(n_727),
.Y(n_782)
);

AND2x2_ASAP7_75t_L g783 ( 
.A(n_721),
.B(n_24),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_L g784 ( 
.A(n_697),
.B(n_25),
.Y(n_784)
);

AO32x2_ASAP7_75t_L g785 ( 
.A1(n_674),
.A2(n_26),
.A3(n_27),
.B1(n_28),
.B2(n_29),
.Y(n_785)
);

AOI21x1_ASAP7_75t_SL g786 ( 
.A1(n_674),
.A2(n_28),
.B(n_30),
.Y(n_786)
);

CKINVDCx5p33_ASAP7_75t_R g787 ( 
.A(n_727),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_686),
.Y(n_788)
);

NOR2xp33_ASAP7_75t_R g789 ( 
.A(n_700),
.B(n_683),
.Y(n_789)
);

OA21x2_ASAP7_75t_L g790 ( 
.A1(n_724),
.A2(n_725),
.B(n_674),
.Y(n_790)
);

INVx2_ASAP7_75t_SL g791 ( 
.A(n_700),
.Y(n_791)
);

A2O1A1Ixp33_ASAP7_75t_L g792 ( 
.A1(n_690),
.A2(n_56),
.B(n_57),
.C(n_58),
.Y(n_792)
);

O2A1O1Ixp33_ASAP7_75t_L g793 ( 
.A1(n_722),
.A2(n_59),
.B(n_61),
.C(n_62),
.Y(n_793)
);

OR2x2_ASAP7_75t_L g794 ( 
.A(n_698),
.B(n_63),
.Y(n_794)
);

A2O1A1Ixp33_ASAP7_75t_L g795 ( 
.A1(n_690),
.A2(n_64),
.B(n_65),
.C(n_66),
.Y(n_795)
);

BUFx3_ASAP7_75t_L g796 ( 
.A(n_754),
.Y(n_796)
);

AOI22xp33_ASAP7_75t_L g797 ( 
.A1(n_751),
.A2(n_67),
.B1(n_68),
.B2(n_69),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_735),
.Y(n_798)
);

AOI22xp5_ASAP7_75t_L g799 ( 
.A1(n_761),
.A2(n_74),
.B1(n_76),
.B2(n_77),
.Y(n_799)
);

OR2x2_ASAP7_75t_L g800 ( 
.A(n_744),
.B(n_78),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_750),
.Y(n_801)
);

CKINVDCx6p67_ASAP7_75t_R g802 ( 
.A(n_770),
.Y(n_802)
);

BUFx6f_ASAP7_75t_L g803 ( 
.A(n_763),
.Y(n_803)
);

BUFx2_ASAP7_75t_SL g804 ( 
.A(n_738),
.Y(n_804)
);

OAI22xp5_ASAP7_75t_L g805 ( 
.A1(n_764),
.A2(n_79),
.B1(n_80),
.B2(n_82),
.Y(n_805)
);

BUFx4_ASAP7_75t_R g806 ( 
.A(n_733),
.Y(n_806)
);

OAI22xp5_ASAP7_75t_SL g807 ( 
.A1(n_784),
.A2(n_84),
.B1(n_85),
.B2(n_87),
.Y(n_807)
);

INVx2_ASAP7_75t_L g808 ( 
.A(n_743),
.Y(n_808)
);

AO22x1_ASAP7_75t_L g809 ( 
.A1(n_783),
.A2(n_88),
.B1(n_89),
.B2(n_90),
.Y(n_809)
);

INVx2_ASAP7_75t_SL g810 ( 
.A(n_787),
.Y(n_810)
);

AOI21xp5_ASAP7_75t_L g811 ( 
.A1(n_768),
.A2(n_91),
.B(n_92),
.Y(n_811)
);

NAND2x1p5_ASAP7_75t_L g812 ( 
.A(n_781),
.B(n_94),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_759),
.Y(n_813)
);

AOI22xp33_ASAP7_75t_L g814 ( 
.A1(n_756),
.A2(n_96),
.B1(n_97),
.B2(n_99),
.Y(n_814)
);

INVx1_ASAP7_75t_SL g815 ( 
.A(n_742),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_747),
.Y(n_816)
);

BUFx12f_ASAP7_75t_L g817 ( 
.A(n_775),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_778),
.Y(n_818)
);

AOI22xp33_ASAP7_75t_SL g819 ( 
.A1(n_752),
.A2(n_101),
.B1(n_103),
.B2(n_104),
.Y(n_819)
);

INVx2_ASAP7_75t_L g820 ( 
.A(n_739),
.Y(n_820)
);

BUFx6f_ASAP7_75t_L g821 ( 
.A(n_763),
.Y(n_821)
);

BUFx12f_ASAP7_75t_L g822 ( 
.A(n_762),
.Y(n_822)
);

BUFx12f_ASAP7_75t_L g823 ( 
.A(n_762),
.Y(n_823)
);

AOI21xp33_ASAP7_75t_L g824 ( 
.A1(n_734),
.A2(n_106),
.B(n_107),
.Y(n_824)
);

AOI22xp33_ASAP7_75t_L g825 ( 
.A1(n_771),
.A2(n_109),
.B1(n_124),
.B2(n_127),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_L g826 ( 
.A(n_767),
.B(n_128),
.Y(n_826)
);

INVx2_ASAP7_75t_SL g827 ( 
.A(n_748),
.Y(n_827)
);

OAI22xp5_ASAP7_75t_L g828 ( 
.A1(n_757),
.A2(n_129),
.B1(n_130),
.B2(n_132),
.Y(n_828)
);

AOI21xp33_ASAP7_75t_L g829 ( 
.A1(n_793),
.A2(n_133),
.B(n_134),
.Y(n_829)
);

AOI21xp33_ASAP7_75t_L g830 ( 
.A1(n_777),
.A2(n_758),
.B(n_732),
.Y(n_830)
);

INVx2_ASAP7_75t_L g831 ( 
.A(n_741),
.Y(n_831)
);

INVx6_ASAP7_75t_L g832 ( 
.A(n_760),
.Y(n_832)
);

AOI22xp33_ASAP7_75t_L g833 ( 
.A1(n_755),
.A2(n_135),
.B1(n_137),
.B2(n_138),
.Y(n_833)
);

INVx2_ASAP7_75t_L g834 ( 
.A(n_791),
.Y(n_834)
);

BUFx6f_ASAP7_75t_L g835 ( 
.A(n_737),
.Y(n_835)
);

CKINVDCx11_ASAP7_75t_R g836 ( 
.A(n_745),
.Y(n_836)
);

AOI22xp33_ASAP7_75t_SL g837 ( 
.A1(n_731),
.A2(n_139),
.B1(n_140),
.B2(n_141),
.Y(n_837)
);

AOI22xp33_ASAP7_75t_L g838 ( 
.A1(n_794),
.A2(n_142),
.B1(n_143),
.B2(n_144),
.Y(n_838)
);

OAI22xp5_ASAP7_75t_SL g839 ( 
.A1(n_731),
.A2(n_146),
.B1(n_147),
.B2(n_148),
.Y(n_839)
);

AOI22xp33_ASAP7_75t_L g840 ( 
.A1(n_753),
.A2(n_150),
.B1(n_151),
.B2(n_153),
.Y(n_840)
);

AOI22xp33_ASAP7_75t_L g841 ( 
.A1(n_766),
.A2(n_155),
.B1(n_158),
.B2(n_159),
.Y(n_841)
);

BUFx3_ASAP7_75t_L g842 ( 
.A(n_736),
.Y(n_842)
);

OAI22xp33_ASAP7_75t_L g843 ( 
.A1(n_765),
.A2(n_163),
.B1(n_164),
.B2(n_166),
.Y(n_843)
);

INVx3_ASAP7_75t_L g844 ( 
.A(n_782),
.Y(n_844)
);

NAND2xp33_ASAP7_75t_R g845 ( 
.A(n_789),
.B(n_168),
.Y(n_845)
);

CKINVDCx20_ASAP7_75t_R g846 ( 
.A(n_746),
.Y(n_846)
);

CKINVDCx6p67_ASAP7_75t_R g847 ( 
.A(n_786),
.Y(n_847)
);

AOI22xp33_ASAP7_75t_L g848 ( 
.A1(n_772),
.A2(n_169),
.B1(n_170),
.B2(n_171),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_785),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_740),
.Y(n_850)
);

BUFx4f_ASAP7_75t_SL g851 ( 
.A(n_788),
.Y(n_851)
);

OAI22xp5_ASAP7_75t_L g852 ( 
.A1(n_792),
.A2(n_172),
.B1(n_174),
.B2(n_175),
.Y(n_852)
);

OAI22xp33_ASAP7_75t_L g853 ( 
.A1(n_730),
.A2(n_176),
.B1(n_177),
.B2(n_178),
.Y(n_853)
);

AOI22xp33_ASAP7_75t_L g854 ( 
.A1(n_776),
.A2(n_180),
.B1(n_181),
.B2(n_184),
.Y(n_854)
);

AOI22xp33_ASAP7_75t_SL g855 ( 
.A1(n_839),
.A2(n_769),
.B1(n_779),
.B2(n_780),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_798),
.Y(n_856)
);

AOI221xp5_ASAP7_75t_L g857 ( 
.A1(n_839),
.A2(n_824),
.B1(n_830),
.B2(n_828),
.C(n_837),
.Y(n_857)
);

INVx2_ASAP7_75t_L g858 ( 
.A(n_801),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_813),
.Y(n_859)
);

AOI21x1_ASAP7_75t_L g860 ( 
.A1(n_811),
.A2(n_790),
.B(n_749),
.Y(n_860)
);

OA21x2_ASAP7_75t_L g861 ( 
.A1(n_850),
.A2(n_795),
.B(n_790),
.Y(n_861)
);

BUFx2_ASAP7_75t_L g862 ( 
.A(n_851),
.Y(n_862)
);

HB1xp67_ASAP7_75t_L g863 ( 
.A(n_815),
.Y(n_863)
);

CKINVDCx11_ASAP7_75t_R g864 ( 
.A(n_802),
.Y(n_864)
);

INVx2_ASAP7_75t_L g865 ( 
.A(n_816),
.Y(n_865)
);

A2O1A1Ixp33_ASAP7_75t_L g866 ( 
.A1(n_799),
.A2(n_729),
.B(n_749),
.C(n_774),
.Y(n_866)
);

INVx2_ASAP7_75t_L g867 ( 
.A(n_808),
.Y(n_867)
);

HB1xp67_ASAP7_75t_L g868 ( 
.A(n_815),
.Y(n_868)
);

INVx2_ASAP7_75t_L g869 ( 
.A(n_820),
.Y(n_869)
);

NAND2xp5_ASAP7_75t_L g870 ( 
.A(n_831),
.B(n_729),
.Y(n_870)
);

BUFx2_ASAP7_75t_L g871 ( 
.A(n_849),
.Y(n_871)
);

CKINVDCx11_ASAP7_75t_R g872 ( 
.A(n_836),
.Y(n_872)
);

BUFx2_ASAP7_75t_L g873 ( 
.A(n_846),
.Y(n_873)
);

INVx2_ASAP7_75t_L g874 ( 
.A(n_818),
.Y(n_874)
);

AND2x2_ASAP7_75t_L g875 ( 
.A(n_827),
.B(n_773),
.Y(n_875)
);

INVx1_ASAP7_75t_L g876 ( 
.A(n_847),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_800),
.Y(n_877)
);

HB1xp67_ASAP7_75t_L g878 ( 
.A(n_834),
.Y(n_878)
);

CKINVDCx8_ASAP7_75t_R g879 ( 
.A(n_804),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_826),
.Y(n_880)
);

INVx1_ASAP7_75t_L g881 ( 
.A(n_844),
.Y(n_881)
);

INVx3_ASAP7_75t_L g882 ( 
.A(n_835),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_844),
.Y(n_883)
);

INVx2_ASAP7_75t_L g884 ( 
.A(n_835),
.Y(n_884)
);

INVx4_ASAP7_75t_L g885 ( 
.A(n_835),
.Y(n_885)
);

BUFx3_ASAP7_75t_L g886 ( 
.A(n_817),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_807),
.Y(n_887)
);

INVx3_ASAP7_75t_L g888 ( 
.A(n_803),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_807),
.Y(n_889)
);

AO21x2_ASAP7_75t_L g890 ( 
.A1(n_829),
.A2(n_773),
.B(n_186),
.Y(n_890)
);

INVx2_ASAP7_75t_L g891 ( 
.A(n_803),
.Y(n_891)
);

INVx3_ASAP7_75t_L g892 ( 
.A(n_803),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_828),
.Y(n_893)
);

INVx1_ASAP7_75t_L g894 ( 
.A(n_852),
.Y(n_894)
);

OAI22xp5_ASAP7_75t_L g895 ( 
.A1(n_799),
.A2(n_185),
.B1(n_188),
.B2(n_189),
.Y(n_895)
);

BUFx2_ASAP7_75t_L g896 ( 
.A(n_842),
.Y(n_896)
);

INVx1_ASAP7_75t_L g897 ( 
.A(n_852),
.Y(n_897)
);

OAI22xp33_ASAP7_75t_SL g898 ( 
.A1(n_832),
.A2(n_805),
.B1(n_812),
.B2(n_845),
.Y(n_898)
);

INVx3_ASAP7_75t_L g899 ( 
.A(n_821),
.Y(n_899)
);

INVx1_ASAP7_75t_L g900 ( 
.A(n_821),
.Y(n_900)
);

INVx1_ASAP7_75t_L g901 ( 
.A(n_821),
.Y(n_901)
);

INVx2_ASAP7_75t_L g902 ( 
.A(n_832),
.Y(n_902)
);

INVx2_ASAP7_75t_L g903 ( 
.A(n_809),
.Y(n_903)
);

AO21x2_ASAP7_75t_L g904 ( 
.A1(n_860),
.A2(n_843),
.B(n_853),
.Y(n_904)
);

AND2x2_ASAP7_75t_L g905 ( 
.A(n_874),
.B(n_796),
.Y(n_905)
);

BUFx6f_ASAP7_75t_L g906 ( 
.A(n_885),
.Y(n_906)
);

OR2x2_ASAP7_75t_L g907 ( 
.A(n_871),
.B(n_810),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_856),
.Y(n_908)
);

AND2x2_ASAP7_75t_L g909 ( 
.A(n_874),
.B(n_819),
.Y(n_909)
);

AOI22xp33_ASAP7_75t_L g910 ( 
.A1(n_857),
.A2(n_797),
.B1(n_814),
.B2(n_823),
.Y(n_910)
);

INVxp67_ASAP7_75t_SL g911 ( 
.A(n_863),
.Y(n_911)
);

OR2x2_ASAP7_75t_L g912 ( 
.A(n_871),
.B(n_848),
.Y(n_912)
);

INVx2_ASAP7_75t_L g913 ( 
.A(n_858),
.Y(n_913)
);

INVx3_ASAP7_75t_L g914 ( 
.A(n_858),
.Y(n_914)
);

OR2x2_ASAP7_75t_L g915 ( 
.A(n_868),
.B(n_854),
.Y(n_915)
);

AND2x2_ASAP7_75t_L g916 ( 
.A(n_856),
.B(n_841),
.Y(n_916)
);

BUFx4f_ASAP7_75t_SL g917 ( 
.A(n_886),
.Y(n_917)
);

INVx1_ASAP7_75t_L g918 ( 
.A(n_859),
.Y(n_918)
);

INVx2_ASAP7_75t_SL g919 ( 
.A(n_884),
.Y(n_919)
);

INVx1_ASAP7_75t_L g920 ( 
.A(n_859),
.Y(n_920)
);

NAND2xp5_ASAP7_75t_L g921 ( 
.A(n_877),
.B(n_822),
.Y(n_921)
);

INVx2_ASAP7_75t_L g922 ( 
.A(n_865),
.Y(n_922)
);

OR2x6_ASAP7_75t_L g923 ( 
.A(n_875),
.B(n_806),
.Y(n_923)
);

BUFx2_ASAP7_75t_L g924 ( 
.A(n_875),
.Y(n_924)
);

OAI21x1_ASAP7_75t_L g925 ( 
.A1(n_861),
.A2(n_838),
.B(n_840),
.Y(n_925)
);

AND2x2_ASAP7_75t_L g926 ( 
.A(n_883),
.B(n_833),
.Y(n_926)
);

BUFx4f_ASAP7_75t_SL g927 ( 
.A(n_886),
.Y(n_927)
);

INVx1_ASAP7_75t_L g928 ( 
.A(n_867),
.Y(n_928)
);

INVx3_ASAP7_75t_L g929 ( 
.A(n_884),
.Y(n_929)
);

INVx1_ASAP7_75t_L g930 ( 
.A(n_869),
.Y(n_930)
);

BUFx6f_ASAP7_75t_L g931 ( 
.A(n_885),
.Y(n_931)
);

HB1xp67_ASAP7_75t_L g932 ( 
.A(n_878),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_L g933 ( 
.A(n_877),
.B(n_825),
.Y(n_933)
);

OR2x2_ASAP7_75t_L g934 ( 
.A(n_870),
.B(n_190),
.Y(n_934)
);

CKINVDCx5p33_ASAP7_75t_R g935 ( 
.A(n_872),
.Y(n_935)
);

INVx1_ASAP7_75t_L g936 ( 
.A(n_908),
.Y(n_936)
);

AND2x2_ASAP7_75t_L g937 ( 
.A(n_924),
.B(n_902),
.Y(n_937)
);

HB1xp67_ASAP7_75t_L g938 ( 
.A(n_924),
.Y(n_938)
);

INVx2_ASAP7_75t_L g939 ( 
.A(n_914),
.Y(n_939)
);

AND2x2_ASAP7_75t_L g940 ( 
.A(n_932),
.B(n_902),
.Y(n_940)
);

INVx1_ASAP7_75t_L g941 ( 
.A(n_908),
.Y(n_941)
);

INVx1_ASAP7_75t_L g942 ( 
.A(n_918),
.Y(n_942)
);

INVx1_ASAP7_75t_L g943 ( 
.A(n_918),
.Y(n_943)
);

INVx1_ASAP7_75t_L g944 ( 
.A(n_920),
.Y(n_944)
);

INVxp67_ASAP7_75t_SL g945 ( 
.A(n_914),
.Y(n_945)
);

AND2x2_ASAP7_75t_L g946 ( 
.A(n_923),
.B(n_873),
.Y(n_946)
);

AND2x2_ASAP7_75t_L g947 ( 
.A(n_923),
.B(n_873),
.Y(n_947)
);

INVx5_ASAP7_75t_L g948 ( 
.A(n_923),
.Y(n_948)
);

INVx1_ASAP7_75t_L g949 ( 
.A(n_920),
.Y(n_949)
);

INVx4_ASAP7_75t_L g950 ( 
.A(n_935),
.Y(n_950)
);

NOR2xp33_ASAP7_75t_SL g951 ( 
.A(n_935),
.B(n_879),
.Y(n_951)
);

NAND2xp5_ASAP7_75t_L g952 ( 
.A(n_911),
.B(n_880),
.Y(n_952)
);

INVx2_ASAP7_75t_L g953 ( 
.A(n_914),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_L g954 ( 
.A(n_905),
.B(n_880),
.Y(n_954)
);

BUFx2_ASAP7_75t_L g955 ( 
.A(n_923),
.Y(n_955)
);

INVx1_ASAP7_75t_L g956 ( 
.A(n_913),
.Y(n_956)
);

INVx2_ASAP7_75t_L g957 ( 
.A(n_913),
.Y(n_957)
);

OR2x2_ASAP7_75t_L g958 ( 
.A(n_922),
.B(n_883),
.Y(n_958)
);

AND2x2_ASAP7_75t_L g959 ( 
.A(n_923),
.B(n_896),
.Y(n_959)
);

AND2x2_ASAP7_75t_L g960 ( 
.A(n_905),
.B(n_896),
.Y(n_960)
);

INVx4_ASAP7_75t_L g961 ( 
.A(n_950),
.Y(n_961)
);

OR2x2_ASAP7_75t_L g962 ( 
.A(n_938),
.B(n_907),
.Y(n_962)
);

INVx2_ASAP7_75t_L g963 ( 
.A(n_939),
.Y(n_963)
);

BUFx3_ASAP7_75t_L g964 ( 
.A(n_950),
.Y(n_964)
);

BUFx6f_ASAP7_75t_L g965 ( 
.A(n_950),
.Y(n_965)
);

AND2x2_ASAP7_75t_L g966 ( 
.A(n_955),
.B(n_929),
.Y(n_966)
);

INVx1_ASAP7_75t_L g967 ( 
.A(n_942),
.Y(n_967)
);

OR2x2_ASAP7_75t_L g968 ( 
.A(n_954),
.B(n_907),
.Y(n_968)
);

INVx1_ASAP7_75t_L g969 ( 
.A(n_942),
.Y(n_969)
);

OR2x2_ASAP7_75t_L g970 ( 
.A(n_955),
.B(n_928),
.Y(n_970)
);

INVx1_ASAP7_75t_L g971 ( 
.A(n_943),
.Y(n_971)
);

NAND2xp5_ASAP7_75t_L g972 ( 
.A(n_940),
.B(n_930),
.Y(n_972)
);

HB1xp67_ASAP7_75t_L g973 ( 
.A(n_943),
.Y(n_973)
);

INVx2_ASAP7_75t_L g974 ( 
.A(n_939),
.Y(n_974)
);

AND2x2_ASAP7_75t_L g975 ( 
.A(n_948),
.B(n_929),
.Y(n_975)
);

INVx1_ASAP7_75t_L g976 ( 
.A(n_944),
.Y(n_976)
);

AND2x2_ASAP7_75t_L g977 ( 
.A(n_948),
.B(n_959),
.Y(n_977)
);

INVx2_ASAP7_75t_L g978 ( 
.A(n_963),
.Y(n_978)
);

AND2x4_ASAP7_75t_L g979 ( 
.A(n_977),
.B(n_948),
.Y(n_979)
);

AND2x4_ASAP7_75t_L g980 ( 
.A(n_977),
.B(n_948),
.Y(n_980)
);

OR2x2_ASAP7_75t_L g981 ( 
.A(n_970),
.B(n_952),
.Y(n_981)
);

AND2x2_ASAP7_75t_L g982 ( 
.A(n_966),
.B(n_948),
.Y(n_982)
);

AND2x2_ASAP7_75t_L g983 ( 
.A(n_966),
.B(n_975),
.Y(n_983)
);

INVx1_ASAP7_75t_L g984 ( 
.A(n_973),
.Y(n_984)
);

INVx1_ASAP7_75t_L g985 ( 
.A(n_967),
.Y(n_985)
);

OR2x2_ASAP7_75t_L g986 ( 
.A(n_968),
.B(n_940),
.Y(n_986)
);

INVx1_ASAP7_75t_L g987 ( 
.A(n_969),
.Y(n_987)
);

INVx3_ASAP7_75t_L g988 ( 
.A(n_961),
.Y(n_988)
);

AND2x2_ASAP7_75t_L g989 ( 
.A(n_975),
.B(n_959),
.Y(n_989)
);

INVx2_ASAP7_75t_L g990 ( 
.A(n_963),
.Y(n_990)
);

AND2x2_ASAP7_75t_L g991 ( 
.A(n_962),
.B(n_946),
.Y(n_991)
);

INVxp67_ASAP7_75t_L g992 ( 
.A(n_988),
.Y(n_992)
);

INVx2_ASAP7_75t_L g993 ( 
.A(n_979),
.Y(n_993)
);

OR2x2_ASAP7_75t_L g994 ( 
.A(n_986),
.B(n_968),
.Y(n_994)
);

INVx1_ASAP7_75t_L g995 ( 
.A(n_985),
.Y(n_995)
);

AND2x4_ASAP7_75t_L g996 ( 
.A(n_988),
.B(n_964),
.Y(n_996)
);

AND2x2_ASAP7_75t_L g997 ( 
.A(n_989),
.B(n_964),
.Y(n_997)
);

INVx1_ASAP7_75t_L g998 ( 
.A(n_987),
.Y(n_998)
);

AND2x2_ASAP7_75t_L g999 ( 
.A(n_989),
.B(n_961),
.Y(n_999)
);

INVxp67_ASAP7_75t_L g1000 ( 
.A(n_988),
.Y(n_1000)
);

OAI22xp33_ASAP7_75t_L g1001 ( 
.A1(n_993),
.A2(n_887),
.B1(n_889),
.B2(n_951),
.Y(n_1001)
);

AO221x2_ASAP7_75t_L g1002 ( 
.A1(n_995),
.A2(n_984),
.B1(n_876),
.B2(n_887),
.C(n_889),
.Y(n_1002)
);

NOR2xp33_ASAP7_75t_L g1003 ( 
.A(n_997),
.B(n_961),
.Y(n_1003)
);

INVx4_ASAP7_75t_L g1004 ( 
.A(n_996),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_L g1005 ( 
.A(n_996),
.B(n_991),
.Y(n_1005)
);

OAI22xp33_ASAP7_75t_L g1006 ( 
.A1(n_994),
.A2(n_903),
.B1(n_965),
.B2(n_981),
.Y(n_1006)
);

INVx1_ASAP7_75t_L g1007 ( 
.A(n_1005),
.Y(n_1007)
);

INVx2_ASAP7_75t_L g1008 ( 
.A(n_1004),
.Y(n_1008)
);

OR2x2_ASAP7_75t_L g1009 ( 
.A(n_1002),
.B(n_998),
.Y(n_1009)
);

INVx1_ASAP7_75t_L g1010 ( 
.A(n_1003),
.Y(n_1010)
);

INVx2_ASAP7_75t_SL g1011 ( 
.A(n_1001),
.Y(n_1011)
);

INVx2_ASAP7_75t_L g1012 ( 
.A(n_1006),
.Y(n_1012)
);

AND2x2_ASAP7_75t_L g1013 ( 
.A(n_1004),
.B(n_999),
.Y(n_1013)
);

INVx1_ASAP7_75t_L g1014 ( 
.A(n_1005),
.Y(n_1014)
);

AND2x2_ASAP7_75t_SL g1015 ( 
.A(n_1004),
.B(n_965),
.Y(n_1015)
);

OR2x2_ASAP7_75t_L g1016 ( 
.A(n_1005),
.B(n_992),
.Y(n_1016)
);

AND2x2_ASAP7_75t_L g1017 ( 
.A(n_1013),
.B(n_979),
.Y(n_1017)
);

AOI211xp5_ASAP7_75t_L g1018 ( 
.A1(n_1008),
.A2(n_1000),
.B(n_992),
.C(n_965),
.Y(n_1018)
);

NAND3xp33_ASAP7_75t_L g1019 ( 
.A(n_1008),
.B(n_1007),
.C(n_1014),
.Y(n_1019)
);

INVxp67_ASAP7_75t_L g1020 ( 
.A(n_1015),
.Y(n_1020)
);

NAND3xp33_ASAP7_75t_L g1021 ( 
.A(n_1016),
.B(n_1000),
.C(n_965),
.Y(n_1021)
);

INVx1_ASAP7_75t_L g1022 ( 
.A(n_1009),
.Y(n_1022)
);

INVx1_ASAP7_75t_L g1023 ( 
.A(n_1015),
.Y(n_1023)
);

AOI22xp5_ASAP7_75t_L g1024 ( 
.A1(n_1011),
.A2(n_979),
.B1(n_980),
.B2(n_982),
.Y(n_1024)
);

OAI22xp33_ASAP7_75t_SL g1025 ( 
.A1(n_1022),
.A2(n_1012),
.B1(n_1010),
.B2(n_980),
.Y(n_1025)
);

OAI21xp33_ASAP7_75t_L g1026 ( 
.A1(n_1024),
.A2(n_1012),
.B(n_980),
.Y(n_1026)
);

XOR2x2_ASAP7_75t_L g1027 ( 
.A(n_1019),
.B(n_864),
.Y(n_1027)
);

INVx1_ASAP7_75t_L g1028 ( 
.A(n_1023),
.Y(n_1028)
);

INVx2_ASAP7_75t_L g1029 ( 
.A(n_1017),
.Y(n_1029)
);

O2A1O1Ixp5_ASAP7_75t_L g1030 ( 
.A1(n_1021),
.A2(n_982),
.B(n_990),
.C(n_978),
.Y(n_1030)
);

OAI22xp33_ASAP7_75t_L g1031 ( 
.A1(n_1020),
.A2(n_879),
.B1(n_927),
.B2(n_917),
.Y(n_1031)
);

OAI322xp33_ASAP7_75t_SL g1032 ( 
.A1(n_1028),
.A2(n_1029),
.A3(n_1025),
.B1(n_1026),
.B2(n_1027),
.C1(n_1018),
.C2(n_1030),
.Y(n_1032)
);

INVx1_ASAP7_75t_L g1033 ( 
.A(n_1031),
.Y(n_1033)
);

AOI21xp33_ASAP7_75t_L g1034 ( 
.A1(n_1025),
.A2(n_876),
.B(n_934),
.Y(n_1034)
);

AO22x2_ASAP7_75t_L g1035 ( 
.A1(n_1029),
.A2(n_990),
.B1(n_978),
.B2(n_983),
.Y(n_1035)
);

INVx2_ASAP7_75t_L g1036 ( 
.A(n_1029),
.Y(n_1036)
);

INVx1_ASAP7_75t_L g1037 ( 
.A(n_1036),
.Y(n_1037)
);

INVx2_ASAP7_75t_L g1038 ( 
.A(n_1035),
.Y(n_1038)
);

INVx1_ASAP7_75t_L g1039 ( 
.A(n_1033),
.Y(n_1039)
);

INVx1_ASAP7_75t_SL g1040 ( 
.A(n_1034),
.Y(n_1040)
);

INVxp67_ASAP7_75t_L g1041 ( 
.A(n_1032),
.Y(n_1041)
);

INVx3_ASAP7_75t_L g1042 ( 
.A(n_1035),
.Y(n_1042)
);

AOI211xp5_ASAP7_75t_L g1043 ( 
.A1(n_1041),
.A2(n_895),
.B(n_898),
.C(n_862),
.Y(n_1043)
);

AOI21xp5_ASAP7_75t_L g1044 ( 
.A1(n_1040),
.A2(n_983),
.B(n_921),
.Y(n_1044)
);

NOR2xp33_ASAP7_75t_L g1045 ( 
.A(n_1037),
.B(n_991),
.Y(n_1045)
);

INVx1_ASAP7_75t_L g1046 ( 
.A(n_1042),
.Y(n_1046)
);

AOI211x1_ASAP7_75t_L g1047 ( 
.A1(n_1039),
.A2(n_946),
.B(n_947),
.C(n_971),
.Y(n_1047)
);

HB1xp67_ASAP7_75t_L g1048 ( 
.A(n_1042),
.Y(n_1048)
);

NAND3xp33_ASAP7_75t_SL g1049 ( 
.A(n_1046),
.B(n_1038),
.C(n_862),
.Y(n_1049)
);

NOR2xp33_ASAP7_75t_L g1050 ( 
.A(n_1045),
.B(n_981),
.Y(n_1050)
);

AOI222xp33_ASAP7_75t_L g1051 ( 
.A1(n_1048),
.A2(n_910),
.B1(n_947),
.B2(n_903),
.C1(n_893),
.C2(n_897),
.Y(n_1051)
);

NAND3xp33_ASAP7_75t_L g1052 ( 
.A(n_1043),
.B(n_934),
.C(n_962),
.Y(n_1052)
);

NAND4xp25_ASAP7_75t_L g1053 ( 
.A(n_1044),
.B(n_933),
.C(n_885),
.D(n_915),
.Y(n_1053)
);

AOI221xp5_ASAP7_75t_L g1054 ( 
.A1(n_1049),
.A2(n_1047),
.B1(n_976),
.B2(n_866),
.C(n_974),
.Y(n_1054)
);

OAI221xp5_ASAP7_75t_SL g1055 ( 
.A1(n_1053),
.A2(n_1050),
.B1(n_1052),
.B2(n_1051),
.C(n_855),
.Y(n_1055)
);

AND2x2_ASAP7_75t_L g1056 ( 
.A(n_1050),
.B(n_960),
.Y(n_1056)
);

OAI211xp5_ASAP7_75t_SL g1057 ( 
.A1(n_1050),
.A2(n_972),
.B(n_915),
.C(n_901),
.Y(n_1057)
);

NAND5xp2_ASAP7_75t_L g1058 ( 
.A(n_1050),
.B(n_909),
.C(n_926),
.D(n_893),
.E(n_894),
.Y(n_1058)
);

OAI22xp5_ASAP7_75t_L g1059 ( 
.A1(n_1052),
.A2(n_974),
.B1(n_906),
.B2(n_931),
.Y(n_1059)
);

OR2x2_ASAP7_75t_L g1060 ( 
.A(n_1049),
.B(n_960),
.Y(n_1060)
);

OAI211xp5_ASAP7_75t_L g1061 ( 
.A1(n_1049),
.A2(n_945),
.B(n_901),
.C(n_900),
.Y(n_1061)
);

NAND2xp5_ASAP7_75t_SL g1062 ( 
.A(n_1060),
.B(n_931),
.Y(n_1062)
);

NOR2x1_ASAP7_75t_L g1063 ( 
.A(n_1061),
.B(n_892),
.Y(n_1063)
);

A2O1A1Ixp33_ASAP7_75t_L g1064 ( 
.A1(n_1055),
.A2(n_900),
.B(n_882),
.C(n_919),
.Y(n_1064)
);

AND2x4_ASAP7_75t_L g1065 ( 
.A(n_1056),
.B(n_882),
.Y(n_1065)
);

NOR2x1_ASAP7_75t_L g1066 ( 
.A(n_1058),
.B(n_899),
.Y(n_1066)
);

NOR3xp33_ASAP7_75t_L g1067 ( 
.A(n_1057),
.B(n_882),
.C(n_899),
.Y(n_1067)
);

INVx1_ASAP7_75t_SL g1068 ( 
.A(n_1059),
.Y(n_1068)
);

NAND4xp25_ASAP7_75t_SL g1069 ( 
.A(n_1054),
.B(n_891),
.C(n_937),
.D(n_912),
.Y(n_1069)
);

NAND3x2_ASAP7_75t_L g1070 ( 
.A(n_1060),
.B(n_958),
.C(n_937),
.Y(n_1070)
);

NAND2x1p5_ASAP7_75t_L g1071 ( 
.A(n_1068),
.B(n_899),
.Y(n_1071)
);

INVxp67_ASAP7_75t_SL g1072 ( 
.A(n_1062),
.Y(n_1072)
);

NAND2xp5_ASAP7_75t_L g1073 ( 
.A(n_1066),
.B(n_881),
.Y(n_1073)
);

INVx1_ASAP7_75t_L g1074 ( 
.A(n_1065),
.Y(n_1074)
);

INVxp67_ASAP7_75t_L g1075 ( 
.A(n_1063),
.Y(n_1075)
);

NOR3xp33_ASAP7_75t_L g1076 ( 
.A(n_1064),
.B(n_888),
.C(n_892),
.Y(n_1076)
);

XNOR2xp5_ASAP7_75t_L g1077 ( 
.A(n_1070),
.B(n_926),
.Y(n_1077)
);

AND2x2_ASAP7_75t_SL g1078 ( 
.A(n_1065),
.B(n_931),
.Y(n_1078)
);

NAND2xp5_ASAP7_75t_SL g1079 ( 
.A(n_1067),
.B(n_906),
.Y(n_1079)
);

NOR2xp33_ASAP7_75t_L g1080 ( 
.A(n_1069),
.B(n_906),
.Y(n_1080)
);

NOR2xp67_ASAP7_75t_L g1081 ( 
.A(n_1069),
.B(n_888),
.Y(n_1081)
);

AND2x4_ASAP7_75t_L g1082 ( 
.A(n_1066),
.B(n_906),
.Y(n_1082)
);

INVx2_ASAP7_75t_L g1083 ( 
.A(n_1071),
.Y(n_1083)
);

AND3x4_ASAP7_75t_L g1084 ( 
.A(n_1082),
.B(n_891),
.C(n_953),
.Y(n_1084)
);

AOI211xp5_ASAP7_75t_SL g1085 ( 
.A1(n_1075),
.A2(n_888),
.B(n_892),
.C(n_909),
.Y(n_1085)
);

AOI21xp5_ASAP7_75t_L g1086 ( 
.A1(n_1072),
.A2(n_890),
.B(n_904),
.Y(n_1086)
);

INVx1_ASAP7_75t_SL g1087 ( 
.A(n_1074),
.Y(n_1087)
);

AND2x2_ASAP7_75t_L g1088 ( 
.A(n_1077),
.B(n_931),
.Y(n_1088)
);

NAND2x1_ASAP7_75t_SL g1089 ( 
.A(n_1081),
.B(n_1080),
.Y(n_1089)
);

AOI22xp5_ASAP7_75t_L g1090 ( 
.A1(n_1079),
.A2(n_931),
.B1(n_906),
.B2(n_919),
.Y(n_1090)
);

NOR2x1_ASAP7_75t_L g1091 ( 
.A(n_1083),
.B(n_1073),
.Y(n_1091)
);

OAI22x1_ASAP7_75t_L g1092 ( 
.A1(n_1087),
.A2(n_1078),
.B1(n_1076),
.B2(n_953),
.Y(n_1092)
);

INVx1_ASAP7_75t_L g1093 ( 
.A(n_1088),
.Y(n_1093)
);

INVx1_ASAP7_75t_L g1094 ( 
.A(n_1089),
.Y(n_1094)
);

HB1xp67_ASAP7_75t_L g1095 ( 
.A(n_1084),
.Y(n_1095)
);

HB1xp67_ASAP7_75t_L g1096 ( 
.A(n_1085),
.Y(n_1096)
);

INVx1_ASAP7_75t_L g1097 ( 
.A(n_1096),
.Y(n_1097)
);

OR2x2_ASAP7_75t_L g1098 ( 
.A(n_1094),
.B(n_1090),
.Y(n_1098)
);

INVx1_ASAP7_75t_L g1099 ( 
.A(n_1095),
.Y(n_1099)
);

OR2x2_ASAP7_75t_L g1100 ( 
.A(n_1097),
.B(n_1093),
.Y(n_1100)
);

INVx1_ASAP7_75t_L g1101 ( 
.A(n_1100),
.Y(n_1101)
);

NAND2xp5_ASAP7_75t_L g1102 ( 
.A(n_1101),
.B(n_1091),
.Y(n_1102)
);

NAND2xp33_ASAP7_75t_L g1103 ( 
.A(n_1101),
.B(n_1099),
.Y(n_1103)
);

AOI22xp33_ASAP7_75t_L g1104 ( 
.A1(n_1103),
.A2(n_1102),
.B1(n_1092),
.B2(n_1098),
.Y(n_1104)
);

AOI22xp5_ASAP7_75t_L g1105 ( 
.A1(n_1103),
.A2(n_1086),
.B1(n_929),
.B2(n_941),
.Y(n_1105)
);

OAI22xp5_ASAP7_75t_SL g1106 ( 
.A1(n_1102),
.A2(n_912),
.B1(n_936),
.B2(n_949),
.Y(n_1106)
);

OAI21xp5_ASAP7_75t_L g1107 ( 
.A1(n_1104),
.A2(n_916),
.B(n_925),
.Y(n_1107)
);

NAND2xp5_ASAP7_75t_L g1108 ( 
.A(n_1105),
.B(n_890),
.Y(n_1108)
);

NAND2xp5_ASAP7_75t_SL g1109 ( 
.A(n_1106),
.B(n_957),
.Y(n_1109)
);

OAI21xp5_ASAP7_75t_L g1110 ( 
.A1(n_1108),
.A2(n_925),
.B(n_916),
.Y(n_1110)
);

OA22x2_ASAP7_75t_L g1111 ( 
.A1(n_1109),
.A2(n_944),
.B1(n_956),
.B2(n_957),
.Y(n_1111)
);

AO22x2_ASAP7_75t_L g1112 ( 
.A1(n_1110),
.A2(n_1107),
.B1(n_956),
.B2(n_958),
.Y(n_1112)
);

AOI211xp5_ASAP7_75t_L g1113 ( 
.A1(n_1112),
.A2(n_1111),
.B(n_897),
.C(n_894),
.Y(n_1113)
);


endmodule