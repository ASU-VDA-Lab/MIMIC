module real_jpeg_23444_n_14 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_2, n_13, n_6, n_7, n_3, n_10, n_9, n_14);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_2;
input n_13;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_14;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_80;
wire n_30;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_216;
wire n_202;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_323;
wire n_166;
wire n_176;
wire n_215;
wire n_286;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_16;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_299;
wire n_243;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_32;
wire n_228;
wire n_15;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

INVx3_ASAP7_75t_L g99 ( 
.A(n_0),
.Y(n_99)
);

INVx6_ASAP7_75t_L g100 ( 
.A(n_0),
.Y(n_100)
);

INVx6_ASAP7_75t_L g203 ( 
.A(n_0),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_0),
.B(n_2),
.Y(n_265)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_SL g37 ( 
.A1(n_2),
.A2(n_23),
.B1(n_38),
.B2(n_39),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_2),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_2),
.A2(n_38),
.B1(n_58),
.B2(n_59),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_2),
.A2(n_38),
.B1(n_74),
.B2(n_75),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_2),
.A2(n_28),
.B1(n_29),
.B2(n_38),
.Y(n_125)
);

O2A1O1Ixp33_ASAP7_75t_L g197 ( 
.A1(n_2),
.A2(n_26),
.B(n_198),
.C(n_199),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_2),
.B(n_27),
.Y(n_214)
);

O2A1O1Ixp33_ASAP7_75t_L g224 ( 
.A1(n_2),
.A2(n_29),
.B(n_56),
.C(n_225),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_2),
.B(n_72),
.C(n_74),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_SL g246 ( 
.A(n_2),
.B(n_54),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_SL g269 ( 
.A(n_2),
.B(n_70),
.Y(n_269)
);

BUFx12f_ASAP7_75t_L g73 ( 
.A(n_3),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g14 ( 
.A1(n_4),
.A2(n_5),
.B1(n_15),
.B2(n_16),
.Y(n_14)
);

INVx13_ASAP7_75t_L g15 ( 
.A(n_5),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_6),
.Y(n_76)
);

BUFx10_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_SL g31 ( 
.A1(n_8),
.A2(n_32),
.B1(n_33),
.B2(n_34),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_8),
.Y(n_33)
);

AOI22xp33_ASAP7_75t_L g64 ( 
.A1(n_8),
.A2(n_28),
.B1(n_29),
.B2(n_33),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_8),
.A2(n_33),
.B1(n_58),
.B2(n_59),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_8),
.A2(n_33),
.B1(n_74),
.B2(n_75),
.Y(n_120)
);

OAI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_9),
.A2(n_23),
.B1(n_24),
.B2(n_130),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_9),
.Y(n_130)
);

OAI22xp33_ASAP7_75t_SL g185 ( 
.A1(n_9),
.A2(n_28),
.B1(n_29),
.B2(n_130),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_L g229 ( 
.A1(n_9),
.A2(n_58),
.B1(n_59),
.B2(n_130),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_9),
.A2(n_74),
.B1(n_75),
.B2(n_130),
.Y(n_254)
);

BUFx5_ASAP7_75t_L g57 ( 
.A(n_10),
.Y(n_57)
);

INVx13_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_12),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_SL g52 ( 
.A1(n_13),
.A2(n_28),
.B1(n_29),
.B2(n_53),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_13),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_13),
.A2(n_53),
.B1(n_58),
.B2(n_59),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_13),
.A2(n_23),
.B1(n_39),
.B2(n_53),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_13),
.A2(n_53),
.B1(n_74),
.B2(n_75),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g16 ( 
.A(n_17),
.B(n_325),
.Y(n_16)
);

OAI221xp5_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_41),
.B1(n_45),
.B2(n_322),
.C(n_324),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_18),
.B(n_323),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_SL g324 ( 
.A(n_18),
.B(n_323),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_18),
.B(n_41),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_SL g18 ( 
.A(n_19),
.B(n_35),
.Y(n_18)
);

AOI21xp5_ASAP7_75t_L g142 ( 
.A1(n_19),
.A2(n_27),
.B(n_143),
.Y(n_142)
);

CKINVDCx14_ASAP7_75t_R g19 ( 
.A(n_20),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_20),
.B(n_168),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g20 ( 
.A(n_21),
.B(n_31),
.Y(n_20)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_21),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_21),
.B(n_37),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_21),
.B(n_129),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_27),
.Y(n_21)
);

AOI22xp33_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_24),
.B1(n_25),
.B2(n_26),
.Y(n_22)
);

INVx8_ASAP7_75t_L g199 ( 
.A(n_23),
.Y(n_199)
);

INVx11_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_24),
.Y(n_32)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_24),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_L g27 ( 
.A1(n_25),
.A2(n_26),
.B1(n_28),
.B2(n_29),
.Y(n_27)
);

OAI21xp33_ASAP7_75t_L g198 ( 
.A1(n_25),
.A2(n_29),
.B(n_38),
.Y(n_198)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_SL g36 ( 
.A(n_27),
.B(n_37),
.Y(n_36)
);

INVxp67_ASAP7_75t_L g43 ( 
.A(n_27),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_27),
.B(n_31),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_27),
.B(n_129),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_L g63 ( 
.A1(n_28),
.A2(n_29),
.B1(n_56),
.B2(n_60),
.Y(n_63)
);

INVx3_ASAP7_75t_SL g28 ( 
.A(n_29),
.Y(n_28)
);

CKINVDCx6p67_ASAP7_75t_R g29 ( 
.A(n_30),
.Y(n_29)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_32),
.Y(n_34)
);

INVxp33_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_36),
.B(n_128),
.Y(n_127)
);

INVxp67_ASAP7_75t_L g44 ( 
.A(n_37),
.Y(n_44)
);

OAI21xp33_ASAP7_75t_L g225 ( 
.A1(n_38),
.A2(n_58),
.B(n_60),
.Y(n_225)
);

INVx11_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_41),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_41),
.A2(n_97),
.B1(n_106),
.B2(n_111),
.Y(n_110)
);

AOI21xp5_ASAP7_75t_SL g41 ( 
.A1(n_42),
.A2(n_43),
.B(n_44),
.Y(n_41)
);

OAI21xp5_ASAP7_75t_SL g316 ( 
.A1(n_42),
.A2(n_85),
.B(n_317),
.Y(n_316)
);

AOI21xp5_ASAP7_75t_L g45 ( 
.A1(n_46),
.A2(n_311),
.B(n_321),
.Y(n_45)
);

OAI211xp5_ASAP7_75t_L g46 ( 
.A1(n_47),
.A2(n_131),
.B(n_146),
.C(n_310),
.Y(n_46)
);

OR2x2_ASAP7_75t_L g47 ( 
.A(n_48),
.B(n_107),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_48),
.B(n_107),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_L g48 ( 
.A(n_49),
.B(n_96),
.Y(n_48)
);

XOR2xp5_ASAP7_75t_L g49 ( 
.A(n_50),
.B(n_82),
.Y(n_49)
);

OAI21xp5_ASAP7_75t_SL g112 ( 
.A1(n_50),
.A2(n_51),
.B(n_65),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_50),
.B(n_82),
.C(n_96),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_51),
.B(n_65),
.Y(n_50)
);

AOI21xp5_ASAP7_75t_L g51 ( 
.A1(n_52),
.A2(n_54),
.B(n_61),
.Y(n_51)
);

AOI21xp5_ASAP7_75t_L g88 ( 
.A1(n_52),
.A2(n_89),
.B(n_90),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_54),
.B(n_185),
.Y(n_184)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_55),
.B(n_63),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_SL g90 ( 
.A(n_55),
.B(n_64),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_55),
.B(n_141),
.Y(n_140)
);

AOI21xp5_ASAP7_75t_L g166 ( 
.A1(n_55),
.A2(n_62),
.B(n_141),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g55 ( 
.A1(n_56),
.A2(n_58),
.B1(n_59),
.B2(n_60),
.Y(n_55)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_56),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_L g80 ( 
.A1(n_58),
.A2(n_59),
.B1(n_71),
.B2(n_72),
.Y(n_80)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_59),
.B(n_242),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_61),
.B(n_140),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_SL g182 ( 
.A(n_61),
.B(n_183),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_SL g61 ( 
.A(n_62),
.B(n_64),
.Y(n_61)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_62),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_SL g191 ( 
.A(n_62),
.B(n_192),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_66),
.B(n_77),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_66),
.B(n_227),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_SL g66 ( 
.A(n_67),
.B(n_69),
.Y(n_66)
);

AOI21xp5_ASAP7_75t_SL g92 ( 
.A1(n_67),
.A2(n_69),
.B(n_93),
.Y(n_92)
);

CKINVDCx16_ASAP7_75t_R g67 ( 
.A(n_68),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_68),
.B(n_79),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_L g121 ( 
.A1(n_69),
.A2(n_78),
.B(n_104),
.Y(n_121)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_70),
.B(n_80),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_70),
.B(n_81),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_70),
.B(n_229),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_71),
.A2(n_72),
.B1(n_74),
.B2(n_75),
.Y(n_70)
);

INVx13_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

BUFx24_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_74),
.B(n_99),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g264 ( 
.A(n_74),
.B(n_265),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g74 ( 
.A(n_75),
.Y(n_74)
);

INVx6_ASAP7_75t_SL g75 ( 
.A(n_76),
.Y(n_75)
);

INVxp33_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_78),
.B(n_239),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_79),
.B(n_81),
.Y(n_78)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_79),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_79),
.B(n_229),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_83),
.A2(n_86),
.B1(n_94),
.B2(n_95),
.Y(n_82)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_83),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_83),
.A2(n_94),
.B1(n_136),
.B2(n_144),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_83),
.B(n_88),
.C(n_91),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_83),
.B(n_136),
.C(n_145),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_84),
.B(n_85),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_84),
.B(n_168),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_85),
.B(n_128),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_86),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_87),
.A2(n_88),
.B1(n_91),
.B2(n_92),
.Y(n_86)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_89),
.B(n_125),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_90),
.B(n_123),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_90),
.B(n_191),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_91),
.A2(n_92),
.B1(n_138),
.B2(n_139),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_91),
.B(n_180),
.C(n_182),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_91),
.A2(n_92),
.B1(n_182),
.B2(n_210),
.Y(n_209)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_92),
.B(n_139),
.C(n_142),
.Y(n_314)
);

OAI21xp5_ASAP7_75t_SL g103 ( 
.A1(n_93),
.A2(n_104),
.B(n_105),
.Y(n_103)
);

AOI21xp33_ASAP7_75t_L g96 ( 
.A1(n_97),
.A2(n_102),
.B(n_106),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_97),
.B(n_103),
.Y(n_102)
);

CKINVDCx16_ASAP7_75t_R g111 ( 
.A(n_97),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_97),
.A2(n_103),
.B1(n_111),
.B2(n_155),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_97),
.B(n_224),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_L g280 ( 
.A1(n_97),
.A2(n_111),
.B1(n_224),
.B2(n_281),
.Y(n_280)
);

AOI21xp5_ASAP7_75t_L g97 ( 
.A1(n_98),
.A2(n_100),
.B(n_101),
.Y(n_97)
);

OR2x2_ASAP7_75t_L g119 ( 
.A(n_98),
.B(n_120),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_SL g159 ( 
.A1(n_98),
.A2(n_160),
.B(n_161),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_SL g216 ( 
.A(n_98),
.B(n_101),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_SL g252 ( 
.A(n_98),
.B(n_253),
.Y(n_252)
);

INVx5_ASAP7_75t_L g117 ( 
.A(n_100),
.Y(n_117)
);

INVxp67_ASAP7_75t_L g118 ( 
.A(n_101),
.Y(n_118)
);

XOR2xp5_ASAP7_75t_L g109 ( 
.A(n_102),
.B(n_110),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_103),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_105),
.B(n_165),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_105),
.B(n_228),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_108),
.B(n_112),
.C(n_113),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_108),
.A2(n_109),
.B1(n_112),
.B2(n_171),
.Y(n_170)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_112),
.Y(n_171)
);

XOR2xp5_ASAP7_75t_L g169 ( 
.A(n_113),
.B(n_170),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_114),
.B(n_122),
.C(n_126),
.Y(n_113)
);

XOR2xp5_ASAP7_75t_L g151 ( 
.A(n_114),
.B(n_152),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_115),
.B(n_121),
.Y(n_114)
);

XOR2xp5_ASAP7_75t_L g301 ( 
.A(n_115),
.B(n_121),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_116),
.B(n_119),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_116),
.B(n_251),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_117),
.B(n_118),
.Y(n_116)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_117),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g259 ( 
.A(n_117),
.B(n_254),
.Y(n_259)
);

OAI21xp5_ASAP7_75t_L g200 ( 
.A1(n_119),
.A2(n_160),
.B(n_201),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_119),
.B(n_259),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_120),
.B(n_163),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_122),
.A2(n_126),
.B1(n_127),
.B2(n_153),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_122),
.Y(n_153)
);

CKINVDCx14_ASAP7_75t_R g123 ( 
.A(n_124),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_124),
.B(n_184),
.Y(n_278)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_125),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_127),
.Y(n_126)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

NAND3xp33_ASAP7_75t_SL g146 ( 
.A(n_132),
.B(n_147),
.C(n_148),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_133),
.B(n_134),
.Y(n_132)
);

OR2x2_ASAP7_75t_L g310 ( 
.A(n_133),
.B(n_134),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_L g134 ( 
.A(n_135),
.B(n_145),
.Y(n_134)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_136),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_142),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_139),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_SL g190 ( 
.A(n_140),
.B(n_191),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g317 ( 
.A(n_143),
.Y(n_317)
);

OAI21xp5_ASAP7_75t_L g148 ( 
.A1(n_149),
.A2(n_172),
.B(n_309),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_169),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g309 ( 
.A(n_150),
.B(n_169),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_154),
.C(n_156),
.Y(n_150)
);

XOR2xp5_ASAP7_75t_L g307 ( 
.A(n_151),
.B(n_154),
.Y(n_307)
);

XOR2xp5_ASAP7_75t_L g306 ( 
.A(n_156),
.B(n_307),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_166),
.C(n_167),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_157),
.A2(n_158),
.B1(n_296),
.B2(n_297),
.Y(n_295)
);

CKINVDCx16_ASAP7_75t_R g157 ( 
.A(n_158),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_164),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_L g178 ( 
.A(n_159),
.B(n_164),
.Y(n_178)
);

INVxp67_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_162),
.B(n_216),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_162),
.B(n_252),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_165),
.B(n_239),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g297 ( 
.A1(n_166),
.A2(n_167),
.B1(n_298),
.B2(n_299),
.Y(n_297)
);

CKINVDCx14_ASAP7_75t_R g298 ( 
.A(n_166),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_L g315 ( 
.A1(n_166),
.A2(n_298),
.B1(n_316),
.B2(n_318),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_166),
.B(n_313),
.C(n_318),
.Y(n_323)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_167),
.Y(n_299)
);

AOI21xp5_ASAP7_75t_L g172 ( 
.A1(n_173),
.A2(n_304),
.B(n_308),
.Y(n_172)
);

A2O1A1Ixp33_ASAP7_75t_SL g173 ( 
.A1(n_174),
.A2(n_217),
.B(n_290),
.C(n_303),
.Y(n_173)
);

OR2x2_ASAP7_75t_L g174 ( 
.A(n_175),
.B(n_205),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_175),
.B(n_205),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_176),
.A2(n_177),
.B1(n_188),
.B2(n_204),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g177 ( 
.A1(n_178),
.A2(n_179),
.B1(n_186),
.B2(n_187),
.Y(n_177)
);

CKINVDCx16_ASAP7_75t_R g186 ( 
.A(n_178),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_178),
.B(n_187),
.C(n_204),
.Y(n_291)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_179),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_180),
.A2(n_181),
.B1(n_208),
.B2(n_209),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_181),
.Y(n_180)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_182),
.Y(n_210)
);

CKINVDCx14_ASAP7_75t_R g183 ( 
.A(n_184),
.Y(n_183)
);

INVxp67_ASAP7_75t_SL g192 ( 
.A(n_185),
.Y(n_192)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_188),
.Y(n_204)
);

XOR2xp5_ASAP7_75t_L g188 ( 
.A(n_189),
.B(n_196),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_190),
.A2(n_193),
.B1(n_194),
.B2(n_195),
.Y(n_189)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_190),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_190),
.B(n_195),
.C(n_196),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_193),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_200),
.Y(n_196)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_197),
.B(n_200),
.Y(n_211)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_206),
.B(n_211),
.C(n_212),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_206),
.A2(n_207),
.B1(n_231),
.B2(n_232),
.Y(n_230)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

XOR2xp5_ASAP7_75t_L g232 ( 
.A(n_211),
.B(n_212),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_213),
.B(n_214),
.C(n_215),
.Y(n_212)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_213),
.B(n_222),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_214),
.B(n_215),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_216),
.B(n_267),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_218),
.B(n_289),
.Y(n_217)
);

OAI21xp5_ASAP7_75t_L g218 ( 
.A1(n_219),
.A2(n_233),
.B(n_288),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_220),
.B(n_230),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_SL g288 ( 
.A(n_220),
.B(n_230),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_221),
.B(n_223),
.C(n_226),
.Y(n_220)
);

XOR2xp5_ASAP7_75t_L g285 ( 
.A(n_221),
.B(n_286),
.Y(n_285)
);

XOR2xp5_ASAP7_75t_L g286 ( 
.A(n_223),
.B(n_226),
.Y(n_286)
);

CKINVDCx16_ASAP7_75t_R g281 ( 
.A(n_224),
.Y(n_281)
);

INVxp33_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

CKINVDCx14_ASAP7_75t_R g231 ( 
.A(n_232),
.Y(n_231)
);

AOI21xp5_ASAP7_75t_L g233 ( 
.A1(n_234),
.A2(n_283),
.B(n_287),
.Y(n_233)
);

OAI21xp5_ASAP7_75t_SL g234 ( 
.A1(n_235),
.A2(n_274),
.B(n_282),
.Y(n_234)
);

AOI21xp5_ASAP7_75t_L g235 ( 
.A1(n_236),
.A2(n_256),
.B(n_273),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_237),
.B(n_243),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_SL g273 ( 
.A(n_237),
.B(n_243),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_238),
.B(n_240),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_238),
.A2(n_240),
.B1(n_241),
.B2(n_261),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_238),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_241),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_244),
.A2(n_245),
.B1(n_250),
.B2(n_255),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_L g245 ( 
.A1(n_246),
.A2(n_247),
.B1(n_248),
.B2(n_249),
.Y(n_245)
);

CKINVDCx14_ASAP7_75t_R g248 ( 
.A(n_246),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_246),
.B(n_249),
.C(n_255),
.Y(n_275)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_247),
.Y(n_249)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_250),
.Y(n_255)
);

INVxp67_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

CKINVDCx16_ASAP7_75t_R g253 ( 
.A(n_254),
.Y(n_253)
);

OAI21xp5_ASAP7_75t_SL g256 ( 
.A1(n_257),
.A2(n_262),
.B(n_272),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_258),
.B(n_260),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_SL g272 ( 
.A(n_258),
.B(n_260),
.Y(n_272)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_259),
.Y(n_267)
);

AOI21xp5_ASAP7_75t_L g262 ( 
.A1(n_263),
.A2(n_268),
.B(n_271),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_264),
.B(n_266),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_269),
.B(n_270),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_SL g271 ( 
.A(n_269),
.B(n_270),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_275),
.B(n_276),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_SL g282 ( 
.A(n_275),
.B(n_276),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_277),
.B(n_280),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_278),
.B(n_279),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_278),
.B(n_279),
.C(n_280),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_284),
.B(n_285),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_SL g287 ( 
.A(n_284),
.B(n_285),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_291),
.B(n_292),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_SL g303 ( 
.A(n_291),
.B(n_292),
.Y(n_303)
);

XOR2xp5_ASAP7_75t_L g292 ( 
.A(n_293),
.B(n_302),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_294),
.A2(n_295),
.B1(n_300),
.B2(n_301),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_294),
.B(n_301),
.C(n_302),
.Y(n_305)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_297),
.Y(n_296)
);

CKINVDCx16_ASAP7_75t_R g300 ( 
.A(n_301),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_305),
.B(n_306),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_SL g308 ( 
.A(n_305),
.B(n_306),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_312),
.B(n_320),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_SL g321 ( 
.A(n_312),
.B(n_320),
.Y(n_321)
);

AOI22xp33_ASAP7_75t_SL g312 ( 
.A1(n_313),
.A2(n_314),
.B1(n_315),
.B2(n_319),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_314),
.Y(n_313)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_315),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_316),
.Y(n_318)
);


endmodule