module fake_jpeg_24799_n_34 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_34);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_34;

wire n_13;
wire n_21;
wire n_33;
wire n_23;
wire n_27;
wire n_22;
wire n_14;
wire n_19;
wire n_20;
wire n_18;
wire n_30;
wire n_16;
wire n_24;
wire n_28;
wire n_26;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_32;
wire n_15;

BUFx5_ASAP7_75t_L g13 ( 
.A(n_11),
.Y(n_13)
);

INVx11_ASAP7_75t_L g14 ( 
.A(n_10),
.Y(n_14)
);

INVx3_ASAP7_75t_L g15 ( 
.A(n_1),
.Y(n_15)
);

INVx3_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

INVx8_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

INVx13_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

INVx3_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

AOI21xp33_ASAP7_75t_L g25 ( 
.A1(n_22),
.A2(n_23),
.B(n_4),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_20),
.B(n_0),
.Y(n_23)
);

AOI22xp33_ASAP7_75t_L g24 ( 
.A1(n_17),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_L g26 ( 
.A1(n_24),
.A2(n_21),
.B1(n_15),
.B2(n_16),
.Y(n_26)
);

INVxp67_ASAP7_75t_SL g27 ( 
.A(n_25),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_27),
.Y(n_28)
);

AOI22xp5_ASAP7_75t_L g29 ( 
.A1(n_28),
.A2(n_26),
.B1(n_22),
.B2(n_20),
.Y(n_29)
);

INVxp67_ASAP7_75t_L g30 ( 
.A(n_29),
.Y(n_30)
);

AO21x1_ASAP7_75t_L g31 ( 
.A1(n_30),
.A2(n_18),
.B(n_19),
.Y(n_31)
);

OAI21xp5_ASAP7_75t_SL g32 ( 
.A1(n_31),
.A2(n_18),
.B(n_19),
.Y(n_32)
);

INVxp67_ASAP7_75t_L g33 ( 
.A(n_32),
.Y(n_33)
);

A2O1A1Ixp33_ASAP7_75t_L g34 ( 
.A1(n_33),
.A2(n_14),
.B(n_7),
.C(n_8),
.Y(n_34)
);


endmodule