module fake_jpeg_16565_n_115 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_115);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_115;

wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

BUFx6f_ASAP7_75t_L g12 ( 
.A(n_7),
.Y(n_12)
);

BUFx12f_ASAP7_75t_L g13 ( 
.A(n_0),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_3),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_4),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_5),
.Y(n_17)
);

BUFx10_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_1),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_7),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_11),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_0),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_1),
.Y(n_23)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_26),
.Y(n_40)
);

AND2x2_ASAP7_75t_L g27 ( 
.A(n_16),
.B(n_0),
.Y(n_27)
);

AND2x2_ASAP7_75t_L g39 ( 
.A(n_27),
.B(n_23),
.Y(n_39)
);

INVx11_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

INVx11_ASAP7_75t_L g43 ( 
.A(n_28),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_15),
.Y(n_29)
);

BUFx2_ASAP7_75t_SL g44 ( 
.A(n_29),
.Y(n_44)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_30),
.B(n_32),
.Y(n_48)
);

INVx5_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

INVx2_ASAP7_75t_SL g41 ( 
.A(n_31),
.Y(n_41)
);

INVx6_ASAP7_75t_SL g32 ( 
.A(n_13),
.Y(n_32)
);

INVx5_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_33),
.B(n_34),
.Y(n_49)
);

INVx11_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_13),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_35),
.Y(n_50)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_12),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_36),
.Y(n_53)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_12),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_37),
.B(n_18),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g38 ( 
.A1(n_28),
.A2(n_24),
.B1(n_23),
.B2(n_22),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_L g67 ( 
.A1(n_38),
.A2(n_42),
.B1(n_20),
.B2(n_29),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_SL g68 ( 
.A(n_39),
.B(n_46),
.Y(n_68)
);

OAI22xp33_ASAP7_75t_SL g42 ( 
.A1(n_28),
.A2(n_34),
.B1(n_24),
.B2(n_19),
.Y(n_42)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_45),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_27),
.B(n_16),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_L g47 ( 
.A1(n_36),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_47),
.A2(n_52),
.B1(n_25),
.B2(n_20),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_27),
.B(n_22),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_51),
.B(n_21),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g52 ( 
.A1(n_30),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_52)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_54),
.B(n_64),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_L g55 ( 
.A1(n_38),
.A2(n_37),
.B1(n_33),
.B2(n_31),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_55),
.A2(n_61),
.B1(n_67),
.B2(n_53),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_51),
.B(n_17),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_SL g71 ( 
.A(n_56),
.B(n_57),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_46),
.B(n_25),
.Y(n_57)
);

OAI21xp5_ASAP7_75t_SL g58 ( 
.A1(n_39),
.A2(n_35),
.B(n_19),
.Y(n_58)
);

AOI21xp5_ASAP7_75t_L g80 ( 
.A1(n_58),
.A2(n_49),
.B(n_8),
.Y(n_80)
);

XNOR2xp5_ASAP7_75t_L g60 ( 
.A(n_45),
.B(n_35),
.Y(n_60)
);

MAJIxp5_ASAP7_75t_L g78 ( 
.A(n_60),
.B(n_26),
.C(n_29),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_62),
.B(n_4),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_48),
.B(n_21),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_SL g77 ( 
.A(n_63),
.B(n_66),
.Y(n_77)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_40),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_39),
.B(n_35),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_65),
.B(n_47),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_50),
.B(n_17),
.Y(n_66)
);

CKINVDCx16_ASAP7_75t_R g70 ( 
.A(n_58),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_SL g83 ( 
.A(n_70),
.B(n_75),
.Y(n_83)
);

INVxp67_ASAP7_75t_L g72 ( 
.A(n_65),
.Y(n_72)
);

INVx13_ASAP7_75t_L g90 ( 
.A(n_72),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_54),
.A2(n_53),
.B1(n_43),
.B2(n_41),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_73),
.A2(n_74),
.B1(n_76),
.B2(n_44),
.Y(n_87)
);

AOI21xp5_ASAP7_75t_SL g76 ( 
.A1(n_59),
.A2(n_50),
.B(n_52),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_78),
.B(n_80),
.C(n_61),
.Y(n_82)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_79),
.Y(n_85)
);

INVx6_ASAP7_75t_L g81 ( 
.A(n_69),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_81),
.B(n_43),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_82),
.B(n_88),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_77),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_84),
.B(n_86),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_76),
.Y(n_86)
);

CKINVDCx14_ASAP7_75t_R g95 ( 
.A(n_87),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_78),
.B(n_60),
.C(n_59),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_88),
.B(n_89),
.C(n_71),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_72),
.B(n_75),
.C(n_68),
.Y(n_89)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_87),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_91),
.B(n_94),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_86),
.A2(n_74),
.B1(n_64),
.B2(n_62),
.Y(n_93)
);

AOI21xp5_ASAP7_75t_L g100 ( 
.A1(n_93),
.A2(n_96),
.B(n_85),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_L g96 ( 
.A1(n_83),
.A2(n_80),
.B(n_68),
.Y(n_96)
);

MAJx2_ASAP7_75t_L g99 ( 
.A(n_97),
.B(n_98),
.C(n_89),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_L g107 ( 
.A1(n_99),
.A2(n_100),
.B(n_81),
.Y(n_107)
);

NOR3xp33_ASAP7_75t_SL g102 ( 
.A(n_96),
.B(n_84),
.C(n_85),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_102),
.B(n_103),
.Y(n_106)
);

AO21x1_ASAP7_75t_L g103 ( 
.A1(n_92),
.A2(n_82),
.B(n_90),
.Y(n_103)
);

XNOR2xp5_ASAP7_75t_SL g104 ( 
.A(n_101),
.B(n_98),
.Y(n_104)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_104),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_101),
.A2(n_95),
.B1(n_90),
.B2(n_93),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_105),
.B(n_26),
.Y(n_109)
);

AOI21xp5_ASAP7_75t_SL g108 ( 
.A1(n_107),
.A2(n_106),
.B(n_104),
.Y(n_108)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_108),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_109),
.B(n_40),
.Y(n_111)
);

AOI332xp33_ASAP7_75t_SL g113 ( 
.A1(n_111),
.A2(n_110),
.A3(n_18),
.B1(n_10),
.B2(n_11),
.B3(n_9),
.C1(n_6),
.C2(n_41),
.Y(n_113)
);

HB1xp67_ASAP7_75t_L g114 ( 
.A(n_113),
.Y(n_114)
);

AOI322xp5_ASAP7_75t_L g115 ( 
.A1(n_114),
.A2(n_112),
.A3(n_9),
.B1(n_6),
.B2(n_18),
.C1(n_41),
.C2(n_32),
.Y(n_115)
);


endmodule