module fake_jpeg_25379_n_332 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_332);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_332;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_145;
wire n_18;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

CKINVDCx16_ASAP7_75t_R g18 ( 
.A(n_6),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

INVx2_ASAP7_75t_SL g20 ( 
.A(n_10),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_7),
.B(n_12),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_2),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_12),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_8),
.Y(n_29)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_15),
.Y(n_31)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_15),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_25),
.Y(n_35)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_35),
.Y(n_53)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_25),
.Y(n_36)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_36),
.Y(n_54)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_25),
.Y(n_37)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_37),
.Y(n_57)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_25),
.Y(n_38)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_38),
.Y(n_59)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_25),
.Y(n_39)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_39),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_22),
.B(n_34),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_40),
.B(n_43),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_34),
.B(n_0),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_41),
.B(n_17),
.Y(n_47)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_25),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_42),
.Y(n_46)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_17),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_34),
.Y(n_44)
);

OR2x2_ASAP7_75t_L g48 ( 
.A(n_44),
.B(n_17),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_24),
.Y(n_45)
);

BUFx2_ASAP7_75t_L g62 ( 
.A(n_45),
.Y(n_62)
);

AND2x2_ASAP7_75t_L g68 ( 
.A(n_47),
.B(n_44),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_48),
.B(n_61),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_37),
.A2(n_33),
.B1(n_32),
.B2(n_24),
.Y(n_49)
);

INVxp67_ASAP7_75t_L g69 ( 
.A(n_49),
.Y(n_69)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_35),
.Y(n_50)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_50),
.Y(n_71)
);

INVx11_ASAP7_75t_L g52 ( 
.A(n_45),
.Y(n_52)
);

INVx8_ASAP7_75t_L g73 ( 
.A(n_52),
.Y(n_73)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_35),
.Y(n_55)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_55),
.Y(n_75)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_35),
.Y(n_56)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_56),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_41),
.A2(n_33),
.B1(n_32),
.B2(n_24),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_58),
.A2(n_20),
.B1(n_30),
.B2(n_16),
.Y(n_94)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_41),
.Y(n_61)
);

HB1xp67_ASAP7_75t_L g63 ( 
.A(n_45),
.Y(n_63)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_63),
.Y(n_74)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_35),
.Y(n_64)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_64),
.Y(n_82)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_45),
.Y(n_65)
);

INVx8_ASAP7_75t_L g87 ( 
.A(n_65),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_40),
.B(n_22),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_66),
.B(n_27),
.Y(n_76)
);

AOI21xp5_ASAP7_75t_L g67 ( 
.A1(n_51),
.A2(n_40),
.B(n_1),
.Y(n_67)
);

INVxp67_ASAP7_75t_L g99 ( 
.A(n_67),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g95 ( 
.A(n_68),
.B(n_76),
.Y(n_95)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_52),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_70),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g72 ( 
.A1(n_47),
.A2(n_61),
.B1(n_51),
.B2(n_43),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_72),
.A2(n_80),
.B1(n_86),
.B2(n_88),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_66),
.B(n_44),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_78),
.B(n_83),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_48),
.A2(n_43),
.B1(n_32),
.B2(n_33),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_L g81 ( 
.A1(n_58),
.A2(n_33),
.B1(n_32),
.B2(n_43),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_L g117 ( 
.A1(n_81),
.A2(n_36),
.B1(n_42),
.B2(n_20),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_48),
.B(n_39),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_60),
.B(n_39),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g98 ( 
.A(n_84),
.B(n_92),
.Y(n_98)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_62),
.Y(n_85)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_85),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_60),
.A2(n_43),
.B1(n_30),
.B2(n_39),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_53),
.A2(n_30),
.B1(n_38),
.B2(n_37),
.Y(n_88)
);

AND2x2_ASAP7_75t_L g89 ( 
.A(n_57),
.B(n_38),
.Y(n_89)
);

A2O1A1Ixp33_ASAP7_75t_L g97 ( 
.A1(n_89),
.A2(n_91),
.B(n_38),
.C(n_37),
.Y(n_97)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_62),
.Y(n_90)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_90),
.Y(n_101)
);

AND2x2_ASAP7_75t_L g91 ( 
.A(n_57),
.B(n_38),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_59),
.B(n_45),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_59),
.B(n_31),
.Y(n_93)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_93),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_94),
.A2(n_20),
.B1(n_64),
.B2(n_56),
.Y(n_118)
);

AND2x2_ASAP7_75t_L g135 ( 
.A(n_97),
.B(n_86),
.Y(n_135)
);

AND2x2_ASAP7_75t_SL g102 ( 
.A(n_72),
.B(n_36),
.Y(n_102)
);

OAI21xp5_ASAP7_75t_SL g131 ( 
.A1(n_102),
.A2(n_109),
.B(n_111),
.Y(n_131)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_87),
.Y(n_103)
);

INVx1_ASAP7_75t_SL g127 ( 
.A(n_103),
.Y(n_127)
);

CKINVDCx16_ASAP7_75t_R g106 ( 
.A(n_92),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_106),
.B(n_113),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_71),
.Y(n_107)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_107),
.Y(n_132)
);

AND2x4_ASAP7_75t_SL g109 ( 
.A(n_83),
.B(n_37),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_71),
.Y(n_110)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_110),
.Y(n_145)
);

AND2x2_ASAP7_75t_L g111 ( 
.A(n_78),
.B(n_79),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_68),
.A2(n_69),
.B1(n_80),
.B2(n_79),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_112),
.A2(n_116),
.B1(n_94),
.B2(n_42),
.Y(n_125)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_75),
.Y(n_113)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_84),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_114),
.B(n_115),
.Y(n_141)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_89),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_68),
.A2(n_53),
.B1(n_42),
.B2(n_36),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_117),
.A2(n_73),
.B1(n_50),
.B2(n_55),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_118),
.A2(n_82),
.B1(n_77),
.B2(n_73),
.Y(n_149)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_87),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_119),
.B(n_121),
.Y(n_151)
);

AOI22x1_ASAP7_75t_SL g120 ( 
.A1(n_67),
.A2(n_21),
.B1(n_42),
.B2(n_36),
.Y(n_120)
);

OAI21xp33_ASAP7_75t_SL g139 ( 
.A1(n_120),
.A2(n_70),
.B(n_85),
.Y(n_139)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_87),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_76),
.B(n_27),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_SL g146 ( 
.A(n_122),
.B(n_31),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_104),
.B(n_93),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_123),
.B(n_126),
.Y(n_160)
);

AOI21xp5_ASAP7_75t_L g124 ( 
.A1(n_115),
.A2(n_91),
.B(n_89),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_L g162 ( 
.A1(n_124),
.A2(n_135),
.B(n_142),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_125),
.A2(n_130),
.B1(n_138),
.B2(n_139),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_111),
.B(n_91),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_111),
.B(n_91),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_128),
.B(n_152),
.Y(n_182)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_98),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_129),
.B(n_140),
.Y(n_158)
);

XOR2xp5_ASAP7_75t_L g134 ( 
.A(n_112),
.B(n_88),
.Y(n_134)
);

XOR2xp5_ASAP7_75t_L g161 ( 
.A(n_134),
.B(n_99),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_107),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_136),
.Y(n_163)
);

AOI21x1_ASAP7_75t_L g137 ( 
.A1(n_120),
.A2(n_89),
.B(n_74),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_L g157 ( 
.A(n_137),
.B(n_118),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_108),
.A2(n_74),
.B1(n_65),
.B2(n_90),
.Y(n_138)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_98),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_SL g142 ( 
.A1(n_109),
.A2(n_16),
.B(n_23),
.Y(n_142)
);

OA21x2_ASAP7_75t_L g143 ( 
.A1(n_105),
.A2(n_46),
.B(n_54),
.Y(n_143)
);

OA21x2_ASAP7_75t_L g170 ( 
.A1(n_143),
.A2(n_121),
.B(n_119),
.Y(n_170)
);

CKINVDCx16_ASAP7_75t_R g144 ( 
.A(n_116),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_144),
.B(n_146),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_108),
.A2(n_82),
.B1(n_77),
.B2(n_75),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_147),
.A2(n_95),
.B1(n_105),
.B2(n_100),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_95),
.B(n_54),
.C(n_46),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_148),
.B(n_97),
.C(n_102),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_149),
.A2(n_102),
.B1(n_114),
.B2(n_100),
.Y(n_155)
);

NAND2xp33_ASAP7_75t_SL g150 ( 
.A(n_109),
.B(n_62),
.Y(n_150)
);

AND2x2_ASAP7_75t_L g184 ( 
.A(n_150),
.B(n_54),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_98),
.B(n_73),
.Y(n_152)
);

FAx1_ASAP7_75t_SL g153 ( 
.A(n_126),
.B(n_95),
.CI(n_109),
.CON(n_153),
.SN(n_153)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_153),
.B(n_167),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_155),
.A2(n_180),
.B1(n_130),
.B2(n_127),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_156),
.B(n_165),
.C(n_172),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_SL g192 ( 
.A1(n_157),
.A2(n_179),
.B(n_181),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_L g207 ( 
.A1(n_159),
.A2(n_173),
.B1(n_19),
.B2(n_29),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g190 ( 
.A(n_161),
.B(n_164),
.Y(n_190)
);

XOR2xp5_ASAP7_75t_L g164 ( 
.A(n_131),
.B(n_99),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_129),
.B(n_140),
.C(n_131),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_133),
.B(n_96),
.Y(n_166)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_166),
.Y(n_187)
);

INVx3_ASAP7_75t_L g167 ( 
.A(n_127),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_151),
.Y(n_168)
);

AOI22xp33_ASAP7_75t_SL g213 ( 
.A1(n_168),
.A2(n_171),
.B1(n_177),
.B2(n_178),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_133),
.B(n_96),
.Y(n_169)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_169),
.Y(n_200)
);

OAI22x1_ASAP7_75t_L g188 ( 
.A1(n_170),
.A2(n_143),
.B1(n_137),
.B2(n_150),
.Y(n_188)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_151),
.Y(n_171)
);

XOR2xp5_ASAP7_75t_L g172 ( 
.A(n_128),
.B(n_101),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_L g173 ( 
.A1(n_144),
.A2(n_149),
.B1(n_152),
.B2(n_123),
.Y(n_173)
);

BUFx6f_ASAP7_75t_L g174 ( 
.A(n_132),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_174),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_136),
.B(n_103),
.Y(n_175)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_175),
.Y(n_209)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_143),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_143),
.Y(n_178)
);

INVxp67_ASAP7_75t_L g179 ( 
.A(n_124),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_134),
.A2(n_135),
.B1(n_148),
.B2(n_125),
.Y(n_180)
);

INVxp67_ASAP7_75t_L g181 ( 
.A(n_141),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_146),
.B(n_101),
.Y(n_183)
);

INVxp67_ASAP7_75t_L g193 ( 
.A(n_183),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_SL g199 ( 
.A1(n_184),
.A2(n_16),
.B(n_28),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_141),
.B(n_113),
.C(n_46),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_185),
.B(n_110),
.C(n_145),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_188),
.A2(n_196),
.B1(n_197),
.B2(n_201),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_154),
.A2(n_135),
.B1(n_138),
.B2(n_147),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_189),
.A2(n_205),
.B1(n_206),
.B2(n_207),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_181),
.B(n_142),
.Y(n_191)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_191),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_180),
.A2(n_127),
.B1(n_132),
.B2(n_145),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_198),
.B(n_204),
.C(n_156),
.Y(n_218)
);

OAI21xp5_ASAP7_75t_L g225 ( 
.A1(n_199),
.A2(n_191),
.B(n_210),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_184),
.A2(n_20),
.B1(n_23),
.B2(n_28),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_160),
.B(n_26),
.Y(n_202)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_202),
.Y(n_231)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_185),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_203),
.B(n_211),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_172),
.B(n_17),
.C(n_19),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_184),
.A2(n_20),
.B1(n_23),
.B2(n_28),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_179),
.A2(n_31),
.B1(n_27),
.B2(n_29),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_154),
.A2(n_29),
.B1(n_26),
.B2(n_19),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_208),
.A2(n_210),
.B1(n_212),
.B2(n_18),
.Y(n_216)
);

AOI22x1_ASAP7_75t_L g210 ( 
.A1(n_170),
.A2(n_19),
.B1(n_21),
.B2(n_2),
.Y(n_210)
);

INVxp67_ASAP7_75t_L g211 ( 
.A(n_159),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_176),
.A2(n_26),
.B1(n_18),
.B2(n_21),
.Y(n_212)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_170),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_214),
.B(n_157),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_L g246 ( 
.A1(n_216),
.A2(n_235),
.B1(n_236),
.B2(n_238),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_194),
.B(n_161),
.Y(n_217)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_217),
.B(n_219),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g258 ( 
.A(n_218),
.B(n_230),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_194),
.B(n_165),
.Y(n_219)
);

HB1xp67_ASAP7_75t_SL g220 ( 
.A(n_188),
.Y(n_220)
);

AOI21xp5_ASAP7_75t_L g242 ( 
.A1(n_220),
.A2(n_232),
.B(n_199),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_190),
.B(n_164),
.C(n_162),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_221),
.B(n_203),
.C(n_187),
.Y(n_243)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_202),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_222),
.B(n_233),
.Y(n_247)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_190),
.B(n_162),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g257 ( 
.A(n_224),
.B(n_227),
.Y(n_257)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_225),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_SL g227 ( 
.A(n_186),
.B(n_160),
.Y(n_227)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_229),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_192),
.B(n_153),
.Y(n_230)
);

OAI21xp5_ASAP7_75t_SL g232 ( 
.A1(n_192),
.A2(n_158),
.B(n_182),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_198),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_SL g234 ( 
.A(n_204),
.B(n_182),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_234),
.B(n_240),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_189),
.A2(n_163),
.B1(n_167),
.B2(n_153),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_211),
.A2(n_174),
.B1(n_1),
.B2(n_2),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_197),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_237),
.B(n_239),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_210),
.A2(n_14),
.B1(n_13),
.B2(n_12),
.Y(n_238)
);

CKINVDCx14_ASAP7_75t_R g239 ( 
.A(n_208),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_SL g240 ( 
.A(n_196),
.B(n_14),
.Y(n_240)
);

OAI21xp5_ASAP7_75t_SL g269 ( 
.A1(n_242),
.A2(n_246),
.B(n_238),
.Y(n_269)
);

XOR2xp5_ASAP7_75t_L g267 ( 
.A(n_243),
.B(n_215),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_228),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_244),
.B(n_245),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_227),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_218),
.B(n_209),
.C(n_200),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_248),
.B(n_250),
.C(n_255),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_219),
.B(n_214),
.C(n_205),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_SL g252 ( 
.A(n_231),
.B(n_213),
.Y(n_252)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_252),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_217),
.B(n_212),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g263 ( 
.A(n_254),
.B(n_230),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_234),
.B(n_201),
.C(n_195),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_224),
.B(n_206),
.C(n_193),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_256),
.B(n_259),
.C(n_11),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_221),
.B(n_193),
.C(n_14),
.Y(n_259)
);

NOR2x1_ASAP7_75t_L g260 ( 
.A(n_216),
.B(n_235),
.Y(n_260)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_260),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_249),
.A2(n_223),
.B1(n_226),
.B2(n_240),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_262),
.B(n_274),
.C(n_259),
.Y(n_285)
);

XOR2xp5_ASAP7_75t_L g283 ( 
.A(n_263),
.B(n_267),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_251),
.A2(n_215),
.B1(n_225),
.B2(n_236),
.Y(n_265)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_265),
.Y(n_281)
);

AOI21xp5_ASAP7_75t_L g290 ( 
.A1(n_269),
.A2(n_272),
.B(n_276),
.Y(n_290)
);

XNOR2x1_ASAP7_75t_L g270 ( 
.A(n_257),
.B(n_13),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_SL g286 ( 
.A(n_270),
.B(n_261),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_260),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_271)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_271),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_253),
.A2(n_0),
.B1(n_3),
.B2(n_4),
.Y(n_272)
);

CKINVDCx16_ASAP7_75t_R g273 ( 
.A(n_247),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g293 ( 
.A(n_273),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_250),
.A2(n_0),
.B1(n_4),
.B2(n_5),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_248),
.Y(n_277)
);

AOI21xp5_ASAP7_75t_L g291 ( 
.A1(n_277),
.A2(n_278),
.B(n_258),
.Y(n_291)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_255),
.Y(n_278)
);

AOI21xp5_ASAP7_75t_SL g279 ( 
.A1(n_275),
.A2(n_261),
.B(n_256),
.Y(n_279)
);

OAI321xp33_ASAP7_75t_L g302 ( 
.A1(n_279),
.A2(n_10),
.A3(n_5),
.B1(n_6),
.B2(n_7),
.C(n_8),
.Y(n_302)
);

BUFx24_ASAP7_75t_SL g280 ( 
.A(n_267),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_280),
.B(n_287),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_264),
.B(n_241),
.C(n_243),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_SL g301 ( 
.A(n_282),
.B(n_285),
.Y(n_301)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_286),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_264),
.B(n_278),
.C(n_274),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_263),
.B(n_241),
.C(n_258),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_SL g304 ( 
.A(n_288),
.B(n_292),
.Y(n_304)
);

XOR2x2_ASAP7_75t_L g289 ( 
.A(n_270),
.B(n_257),
.Y(n_289)
);

OR2x2_ASAP7_75t_L g299 ( 
.A(n_289),
.B(n_272),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_291),
.B(n_262),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_266),
.B(n_10),
.C(n_5),
.Y(n_292)
);

AOI21xp5_ASAP7_75t_L g294 ( 
.A1(n_281),
.A2(n_268),
.B(n_269),
.Y(n_294)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_294),
.Y(n_314)
);

AOI21xp5_ASAP7_75t_L g296 ( 
.A1(n_293),
.A2(n_276),
.B(n_271),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_296),
.B(n_306),
.Y(n_307)
);

XOR2xp5_ASAP7_75t_L g297 ( 
.A(n_283),
.B(n_265),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_297),
.B(n_298),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_299),
.B(n_303),
.Y(n_310)
);

XOR2xp5_ASAP7_75t_L g300 ( 
.A(n_283),
.B(n_4),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_300),
.B(n_6),
.C(n_7),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_L g308 ( 
.A1(n_302),
.A2(n_284),
.B1(n_289),
.B2(n_8),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_290),
.B(n_4),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_SL g306 ( 
.A(n_282),
.B(n_5),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_308),
.B(n_316),
.Y(n_320)
);

AOI22xp5_ASAP7_75t_L g309 ( 
.A1(n_295),
.A2(n_279),
.B1(n_286),
.B2(n_288),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_SL g319 ( 
.A1(n_309),
.A2(n_313),
.B1(n_304),
.B2(n_301),
.Y(n_319)
);

INVx2_ASAP7_75t_L g311 ( 
.A(n_299),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_311),
.B(n_315),
.Y(n_317)
);

FAx1_ASAP7_75t_SL g315 ( 
.A(n_297),
.B(n_6),
.CI(n_9),
.CON(n_315),
.SN(n_315)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_305),
.B(n_9),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_311),
.B(n_300),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_318),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_SL g325 ( 
.A(n_319),
.B(n_321),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_310),
.B(n_9),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_314),
.B(n_9),
.C(n_309),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_322),
.B(n_323),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_307),
.B(n_312),
.C(n_310),
.Y(n_323)
);

HB1xp67_ASAP7_75t_L g327 ( 
.A(n_326),
.Y(n_327)
);

OAI21xp5_ASAP7_75t_SL g328 ( 
.A1(n_327),
.A2(n_325),
.B(n_317),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_328),
.B(n_324),
.C(n_320),
.Y(n_329)
);

OAI21xp5_ASAP7_75t_L g330 ( 
.A1(n_329),
.A2(n_317),
.B(n_315),
.Y(n_330)
);

XNOR2x2_ASAP7_75t_SL g331 ( 
.A(n_330),
.B(n_313),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_SL g332 ( 
.A(n_331),
.B(n_315),
.Y(n_332)
);


endmodule