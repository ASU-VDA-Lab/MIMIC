module real_jpeg_30402_n_8 (n_5, n_4, n_0, n_1, n_2, n_6, n_7, n_3, n_8);

input n_5;
input n_4;
input n_0;
input n_1;
input n_2;
input n_6;
input n_7;
input n_3;

output n_8;

wire n_17;
wire n_37;
wire n_21;
wire n_33;
wire n_35;
wire n_29;
wire n_10;
wire n_31;
wire n_9;
wire n_12;
wire n_24;
wire n_34;
wire n_28;
wire n_23;
wire n_11;
wire n_14;
wire n_25;
wire n_22;
wire n_18;
wire n_36;
wire n_27;
wire n_32;
wire n_20;
wire n_19;
wire n_26;
wire n_30;
wire n_16;
wire n_15;
wire n_13;

CKINVDCx5p33_ASAP7_75t_R g20 ( 
.A(n_0),
.Y(n_20)
);

AND2x2_ASAP7_75t_L g23 ( 
.A(n_0),
.B(n_1),
.Y(n_23)
);

AND2x2_ASAP7_75t_L g35 ( 
.A(n_0),
.B(n_36),
.Y(n_35)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_0),
.Y(n_37)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_1),
.Y(n_36)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_2),
.Y(n_13)
);

NAND2x1p5_ASAP7_75t_L g14 ( 
.A(n_2),
.B(n_15),
.Y(n_14)
);

AOI22xp5_ASAP7_75t_L g32 ( 
.A1(n_3),
.A2(n_9),
.B1(n_33),
.B2(n_37),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_4),
.B(n_19),
.Y(n_18)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

INVx2_ASAP7_75t_L g11 ( 
.A(n_6),
.Y(n_11)
);

AND2x2_ASAP7_75t_L g12 ( 
.A(n_7),
.B(n_13),
.Y(n_12)
);

INVx3_ASAP7_75t_L g15 ( 
.A(n_7),
.Y(n_15)
);

OAI221xp5_ASAP7_75t_L g8 ( 
.A1(n_9),
.A2(n_16),
.B1(n_27),
.B2(n_28),
.C(n_32),
.Y(n_8)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_9),
.B(n_24),
.Y(n_27)
);

INVx1_ASAP7_75t_L g9 ( 
.A(n_10),
.Y(n_9)
);

OA21x2_ASAP7_75t_L g10 ( 
.A1(n_11),
.A2(n_12),
.B(n_14),
.Y(n_10)
);

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_21),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_SL g17 ( 
.A(n_18),
.B(n_20),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_SL g34 ( 
.A(n_18),
.B(n_35),
.Y(n_34)
);

AND2x2_ASAP7_75t_L g26 ( 
.A(n_19),
.B(n_23),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_SL g29 ( 
.A(n_19),
.B(n_30),
.Y(n_29)
);

BUFx12_ASAP7_75t_L g31 ( 
.A(n_20),
.Y(n_31)
);

OAI21xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_24),
.B(n_25),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_23),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_26),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_29),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_34),
.Y(n_33)
);


endmodule