module fake_jpeg_24725_n_283 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_283);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_283;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_252;
wire n_251;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_272;
wire n_280;
wire n_171;
wire n_263;
wire n_119;
wire n_23;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_121;
wire n_99;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

INVx5_ASAP7_75t_L g16 ( 
.A(n_13),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_7),
.Y(n_20)
);

BUFx12_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

INVx13_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_12),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_7),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_13),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_11),
.Y(n_28)
);

INVx11_ASAP7_75t_SL g29 ( 
.A(n_1),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_6),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_1),
.B(n_12),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_20),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_33),
.B(n_37),
.Y(n_56)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_16),
.Y(n_34)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_34),
.Y(n_46)
);

BUFx12_ASAP7_75t_L g35 ( 
.A(n_30),
.Y(n_35)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_35),
.Y(n_54)
);

HB1xp67_ASAP7_75t_L g36 ( 
.A(n_30),
.Y(n_36)
);

INVx5_ASAP7_75t_L g47 ( 
.A(n_36),
.Y(n_47)
);

CKINVDCx14_ASAP7_75t_R g37 ( 
.A(n_30),
.Y(n_37)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_26),
.Y(n_38)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_38),
.Y(n_43)
);

INVx11_ASAP7_75t_L g39 ( 
.A(n_29),
.Y(n_39)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_39),
.Y(n_44)
);

INVx5_ASAP7_75t_L g40 ( 
.A(n_21),
.Y(n_40)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_40),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g41 ( 
.A1(n_38),
.A2(n_18),
.B1(n_16),
.B2(n_22),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_41),
.A2(n_42),
.B1(n_39),
.B2(n_34),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g42 ( 
.A1(n_38),
.A2(n_18),
.B1(n_16),
.B2(n_22),
.Y(n_42)
);

AND2x4_ASAP7_75t_L g45 ( 
.A(n_36),
.B(n_30),
.Y(n_45)
);

AND2x2_ASAP7_75t_L g62 ( 
.A(n_45),
.B(n_37),
.Y(n_62)
);

OAI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_34),
.A2(n_22),
.B1(n_19),
.B2(n_29),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_48),
.A2(n_34),
.B1(n_38),
.B2(n_40),
.Y(n_61)
);

INVx5_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_49),
.B(n_55),
.Y(n_65)
);

AOI21xp33_ASAP7_75t_SL g51 ( 
.A1(n_34),
.A2(n_30),
.B(n_26),
.Y(n_51)
);

XNOR2xp5_ASAP7_75t_L g88 ( 
.A(n_51),
.B(n_21),
.Y(n_88)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

INVx6_ASAP7_75t_L g82 ( 
.A(n_52),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_33),
.B(n_32),
.Y(n_53)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_53),
.Y(n_73)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_39),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_57),
.B(n_59),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_SL g58 ( 
.A(n_33),
.B(n_32),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_58),
.B(n_33),
.Y(n_63)
);

INVx2_ASAP7_75t_SL g59 ( 
.A(n_36),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_60),
.A2(n_83),
.B1(n_85),
.B2(n_42),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_61),
.A2(n_44),
.B1(n_50),
.B2(n_43),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_SL g95 ( 
.A1(n_62),
.A2(n_84),
.B(n_88),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_63),
.B(n_72),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_56),
.B(n_38),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_64),
.B(n_69),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_45),
.A2(n_19),
.B1(n_37),
.B2(n_17),
.Y(n_66)
);

AOI21xp5_ASAP7_75t_L g96 ( 
.A1(n_66),
.A2(n_67),
.B(n_25),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_45),
.A2(n_19),
.B1(n_40),
.B2(n_17),
.Y(n_67)
);

HB1xp67_ASAP7_75t_L g68 ( 
.A(n_45),
.Y(n_68)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_68),
.Y(n_90)
);

AND2x2_ASAP7_75t_SL g69 ( 
.A(n_45),
.B(n_35),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_58),
.B(n_31),
.Y(n_71)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_71),
.Y(n_98)
);

INVx5_ASAP7_75t_L g72 ( 
.A(n_55),
.Y(n_72)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_54),
.Y(n_74)
);

INVx6_ASAP7_75t_L g91 ( 
.A(n_74),
.Y(n_91)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_54),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_75),
.B(n_76),
.Y(n_106)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_56),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_46),
.B(n_31),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_77),
.Y(n_92)
);

INVx5_ASAP7_75t_L g78 ( 
.A(n_57),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_78),
.B(n_80),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_59),
.B(n_21),
.Y(n_79)
);

CKINVDCx16_ASAP7_75t_R g89 ( 
.A(n_79),
.Y(n_89)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_44),
.Y(n_80)
);

NOR2x1_ASAP7_75t_L g81 ( 
.A(n_51),
.B(n_40),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_81),
.A2(n_76),
.B1(n_62),
.B2(n_66),
.Y(n_110)
);

OA22x2_ASAP7_75t_L g83 ( 
.A1(n_41),
.A2(n_40),
.B1(n_35),
.B2(n_26),
.Y(n_83)
);

NAND2x1_ASAP7_75t_SL g84 ( 
.A(n_54),
.B(n_35),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_46),
.A2(n_39),
.B1(n_25),
.B2(n_28),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_59),
.B(n_21),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_86),
.B(n_87),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_47),
.B(n_21),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_82),
.Y(n_93)
);

INVxp33_ASAP7_75t_L g125 ( 
.A(n_93),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_85),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_94),
.B(n_97),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_SL g143 ( 
.A1(n_96),
.A2(n_108),
.B(n_95),
.Y(n_143)
);

INVx8_ASAP7_75t_L g97 ( 
.A(n_72),
.Y(n_97)
);

AND2x6_ASAP7_75t_L g100 ( 
.A(n_81),
.B(n_15),
.Y(n_100)
);

BUFx3_ASAP7_75t_L g140 ( 
.A(n_100),
.Y(n_140)
);

INVx6_ASAP7_75t_SL g101 ( 
.A(n_84),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_101),
.B(n_104),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_102),
.A2(n_110),
.B1(n_115),
.B2(n_62),
.Y(n_117)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_74),
.Y(n_104)
);

BUFx2_ASAP7_75t_L g105 ( 
.A(n_78),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_105),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_70),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_107),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_SL g108 ( 
.A1(n_88),
.A2(n_52),
.B(n_43),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_64),
.B(n_47),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_109),
.B(n_114),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_65),
.B(n_50),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_SL g120 ( 
.A(n_113),
.B(n_75),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_69),
.B(n_35),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_117),
.A2(n_100),
.B1(n_89),
.B2(n_92),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_109),
.B(n_69),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_119),
.B(n_136),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_120),
.B(n_121),
.Y(n_144)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_111),
.Y(n_121)
);

CKINVDCx14_ASAP7_75t_R g123 ( 
.A(n_99),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_123),
.B(n_127),
.Y(n_152)
);

AND2x2_ASAP7_75t_L g124 ( 
.A(n_114),
.B(n_60),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_L g153 ( 
.A1(n_124),
.A2(n_128),
.B(n_132),
.Y(n_153)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_106),
.Y(n_127)
);

AND2x4_ASAP7_75t_L g128 ( 
.A(n_101),
.B(n_84),
.Y(n_128)
);

OR2x2_ASAP7_75t_L g130 ( 
.A(n_94),
.B(n_83),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_SL g173 ( 
.A(n_130),
.B(n_133),
.Y(n_173)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_105),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_131),
.B(n_134),
.Y(n_163)
);

AND2x2_ASAP7_75t_L g132 ( 
.A(n_103),
.B(n_83),
.Y(n_132)
);

OR2x2_ASAP7_75t_L g133 ( 
.A(n_92),
.B(n_83),
.Y(n_133)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_112),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_90),
.A2(n_73),
.B1(n_82),
.B2(n_61),
.Y(n_135)
);

INVxp67_ASAP7_75t_L g168 ( 
.A(n_135),
.Y(n_168)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_105),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_115),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_137),
.B(n_138),
.Y(n_150)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_102),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_103),
.B(n_108),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_139),
.B(n_141),
.Y(n_155)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_93),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_95),
.B(n_73),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_142),
.B(n_35),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g158 ( 
.A1(n_143),
.A2(n_49),
.B1(n_98),
.B2(n_97),
.Y(n_158)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_118),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_146),
.B(n_151),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_139),
.B(n_90),
.C(n_96),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_147),
.B(n_149),
.C(n_156),
.Y(n_189)
);

OR2x2_ASAP7_75t_L g148 ( 
.A(n_129),
.B(n_107),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_SL g196 ( 
.A(n_148),
.B(n_127),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_143),
.B(n_116),
.C(n_142),
.Y(n_149)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_135),
.Y(n_151)
);

OAI21xp33_ASAP7_75t_SL g188 ( 
.A1(n_154),
.A2(n_167),
.B(n_133),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_116),
.B(n_89),
.C(n_98),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_126),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_157),
.B(n_169),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_158),
.A2(n_160),
.B1(n_170),
.B2(n_131),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_L g159 ( 
.A1(n_128),
.A2(n_27),
.B(n_28),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_L g178 ( 
.A(n_159),
.B(n_161),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_138),
.A2(n_97),
.B1(n_91),
.B2(n_80),
.Y(n_160)
);

XOR2xp5_ASAP7_75t_L g161 ( 
.A(n_119),
.B(n_35),
.Y(n_161)
);

NAND3xp33_ASAP7_75t_L g162 ( 
.A(n_140),
.B(n_15),
.C(n_14),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_162),
.B(n_154),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_164),
.B(n_166),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_132),
.B(n_91),
.Y(n_165)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_165),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g166 ( 
.A(n_128),
.B(n_104),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_L g167 ( 
.A1(n_128),
.A2(n_27),
.B(n_24),
.Y(n_167)
);

INVxp67_ASAP7_75t_SL g169 ( 
.A(n_125),
.Y(n_169)
);

OA22x2_ASAP7_75t_L g170 ( 
.A1(n_128),
.A2(n_93),
.B1(n_91),
.B2(n_24),
.Y(n_170)
);

AOI22xp33_ASAP7_75t_SL g171 ( 
.A1(n_122),
.A2(n_23),
.B1(n_20),
.B2(n_3),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_L g198 ( 
.A1(n_171),
.A2(n_23),
.B1(n_141),
.B2(n_3),
.Y(n_198)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_126),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_172),
.B(n_136),
.Y(n_191)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_152),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_174),
.B(n_185),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_176),
.B(n_187),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_168),
.A2(n_137),
.B1(n_140),
.B2(n_130),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_177),
.A2(n_168),
.B1(n_164),
.B2(n_165),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_163),
.B(n_122),
.Y(n_179)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_179),
.Y(n_200)
);

INVx4_ASAP7_75t_L g182 ( 
.A(n_148),
.Y(n_182)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_182),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_183),
.B(n_184),
.Y(n_209)
);

BUFx12_ASAP7_75t_L g184 ( 
.A(n_144),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_145),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_145),
.Y(n_187)
);

CKINVDCx16_ASAP7_75t_R g216 ( 
.A(n_188),
.Y(n_216)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_155),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_190),
.B(n_193),
.Y(n_217)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_191),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_155),
.B(n_134),
.Y(n_192)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_192),
.Y(n_205)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_150),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_156),
.B(n_121),
.Y(n_194)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_194),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_R g195 ( 
.A(n_159),
.B(n_132),
.Y(n_195)
);

AOI21xp5_ASAP7_75t_SL g210 ( 
.A1(n_195),
.A2(n_153),
.B(n_170),
.Y(n_210)
);

AOI21xp5_ASAP7_75t_L g219 ( 
.A1(n_196),
.A2(n_198),
.B(n_173),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_167),
.B(n_124),
.Y(n_197)
);

INVxp67_ASAP7_75t_L g199 ( 
.A(n_197),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_SL g235 ( 
.A(n_201),
.B(n_0),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g206 ( 
.A(n_189),
.B(n_149),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_206),
.B(n_213),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_189),
.B(n_161),
.C(n_147),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_208),
.B(n_211),
.C(n_212),
.Y(n_221)
);

AOI21xp5_ASAP7_75t_SL g231 ( 
.A1(n_210),
.A2(n_193),
.B(n_185),
.Y(n_231)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_180),
.B(n_153),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g212 ( 
.A(n_180),
.B(n_166),
.Y(n_212)
);

NAND3xp33_ASAP7_75t_L g213 ( 
.A(n_195),
.B(n_170),
.C(n_150),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_178),
.B(n_117),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_215),
.B(n_218),
.C(n_183),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_178),
.B(n_124),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_219),
.B(n_175),
.Y(n_223)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_202),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_220),
.B(n_224),
.Y(n_240)
);

AOI21xp5_ASAP7_75t_L g222 ( 
.A1(n_210),
.A2(n_182),
.B(n_181),
.Y(n_222)
);

AOI21xp5_ASAP7_75t_L g238 ( 
.A1(n_222),
.A2(n_231),
.B(n_199),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_223),
.A2(n_234),
.B1(n_205),
.B2(n_218),
.Y(n_239)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_217),
.Y(n_224)
);

INVx13_ASAP7_75t_L g226 ( 
.A(n_200),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_226),
.B(n_214),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_227),
.B(n_235),
.Y(n_249)
);

OR2x2_ASAP7_75t_L g228 ( 
.A(n_209),
.B(n_170),
.Y(n_228)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_228),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_208),
.B(n_181),
.C(n_190),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_229),
.B(n_232),
.C(n_206),
.Y(n_245)
);

HB1xp67_ASAP7_75t_L g230 ( 
.A(n_203),
.Y(n_230)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_230),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_207),
.B(n_186),
.C(n_184),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_204),
.B(n_184),
.Y(n_233)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_233),
.Y(n_246)
);

XNOR2x1_ASAP7_75t_L g234 ( 
.A(n_215),
.B(n_177),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_SL g236 ( 
.A(n_211),
.B(n_0),
.Y(n_236)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_236),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_234),
.A2(n_216),
.B1(n_199),
.B2(n_201),
.Y(n_237)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_237),
.Y(n_259)
);

AOI22xp33_ASAP7_75t_L g256 ( 
.A1(n_238),
.A2(n_231),
.B1(n_235),
.B2(n_4),
.Y(n_256)
);

XOR2xp5_ASAP7_75t_L g252 ( 
.A(n_239),
.B(n_237),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_241),
.B(n_228),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_226),
.B(n_212),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_244),
.B(n_245),
.C(n_248),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_221),
.B(n_0),
.C(n_2),
.Y(n_248)
);

BUFx4f_ASAP7_75t_SL g250 ( 
.A(n_243),
.Y(n_250)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_250),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_SL g262 ( 
.A(n_252),
.B(n_253),
.Y(n_262)
);

AND2x2_ASAP7_75t_L g254 ( 
.A(n_249),
.B(n_225),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_254),
.B(n_257),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_245),
.B(n_230),
.C(n_236),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_255),
.B(n_251),
.C(n_250),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_L g264 ( 
.A1(n_256),
.A2(n_239),
.B1(n_246),
.B2(n_248),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_242),
.B(n_2),
.Y(n_257)
);

AOI31xp67_ASAP7_75t_L g258 ( 
.A1(n_238),
.A2(n_2),
.A3(n_3),
.B(n_5),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_258),
.B(n_5),
.Y(n_268)
);

OAI21xp5_ASAP7_75t_SL g260 ( 
.A1(n_240),
.A2(n_5),
.B(n_6),
.Y(n_260)
);

OAI21xp5_ASAP7_75t_SL g261 ( 
.A1(n_260),
.A2(n_247),
.B(n_259),
.Y(n_261)
);

BUFx24_ASAP7_75t_SL g270 ( 
.A(n_261),
.Y(n_270)
);

INVxp67_ASAP7_75t_L g274 ( 
.A(n_264),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_266),
.B(n_267),
.C(n_256),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_250),
.B(n_249),
.C(n_6),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_268),
.B(n_7),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_269),
.B(n_267),
.C(n_265),
.Y(n_275)
);

OAI21xp5_ASAP7_75t_L g271 ( 
.A1(n_263),
.A2(n_254),
.B(n_8),
.Y(n_271)
);

AOI21xp5_ASAP7_75t_L g277 ( 
.A1(n_271),
.A2(n_273),
.B(n_8),
.Y(n_277)
);

NOR3xp33_ASAP7_75t_SL g278 ( 
.A(n_272),
.B(n_262),
.C(n_10),
.Y(n_278)
);

OAI21xp5_ASAP7_75t_L g273 ( 
.A1(n_266),
.A2(n_8),
.B(n_9),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_275),
.B(n_9),
.C(n_11),
.Y(n_280)
);

INVxp67_ASAP7_75t_L g276 ( 
.A(n_270),
.Y(n_276)
);

A2O1A1Ixp33_ASAP7_75t_L g279 ( 
.A1(n_276),
.A2(n_277),
.B(n_278),
.C(n_274),
.Y(n_279)
);

XOR2xp5_ASAP7_75t_L g281 ( 
.A(n_279),
.B(n_280),
.Y(n_281)
);

XOR2xp5_ASAP7_75t_L g282 ( 
.A(n_281),
.B(n_9),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_282),
.B(n_12),
.Y(n_283)
);


endmodule