module fake_netlist_5_1377_n_653 (n_137, n_91, n_82, n_122, n_142, n_10, n_140, n_24, n_124, n_86, n_136, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_60, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_125, n_35, n_128, n_73, n_17, n_92, n_19, n_120, n_135, n_30, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_29, n_79, n_131, n_47, n_25, n_53, n_8, n_44, n_40, n_34, n_100, n_62, n_138, n_71, n_109, n_112, n_85, n_95, n_119, n_59, n_26, n_133, n_55, n_99, n_2, n_3, n_49, n_20, n_6, n_39, n_54, n_12, n_67, n_121, n_36, n_76, n_87, n_27, n_64, n_77, n_102, n_106, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_134, n_32, n_41, n_104, n_103, n_56, n_51, n_63, n_97, n_141, n_11, n_7, n_15, n_48, n_50, n_52, n_88, n_110, n_653);

input n_137;
input n_91;
input n_82;
input n_122;
input n_142;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_60;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_125;
input n_35;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_120;
input n_135;
input n_30;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_29;
input n_79;
input n_131;
input n_47;
input n_25;
input n_53;
input n_8;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_71;
input n_109;
input n_112;
input n_85;
input n_95;
input n_119;
input n_59;
input n_26;
input n_133;
input n_55;
input n_99;
input n_2;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_27;
input n_64;
input n_77;
input n_102;
input n_106;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_134;
input n_32;
input n_41;
input n_104;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_11;
input n_7;
input n_15;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_653;

wire n_294;
wire n_431;
wire n_318;
wire n_380;
wire n_419;
wire n_611;
wire n_444;
wire n_642;
wire n_469;
wire n_615;
wire n_194;
wire n_316;
wire n_389;
wire n_549;
wire n_418;
wire n_248;
wire n_146;
wire n_315;
wire n_268;
wire n_523;
wire n_451;
wire n_532;
wire n_619;
wire n_408;
wire n_376;
wire n_503;
wire n_235;
wire n_226;
wire n_605;
wire n_515;
wire n_353;
wire n_351;
wire n_367;
wire n_620;
wire n_643;
wire n_452;
wire n_397;
wire n_493;
wire n_525;
wire n_483;
wire n_544;
wire n_155;
wire n_649;
wire n_552;
wire n_547;
wire n_564;
wire n_467;
wire n_423;
wire n_284;
wire n_245;
wire n_501;
wire n_280;
wire n_590;
wire n_629;
wire n_378;
wire n_551;
wire n_581;
wire n_382;
wire n_554;
wire n_254;
wire n_583;
wire n_302;
wire n_265;
wire n_526;
wire n_293;
wire n_372;
wire n_443;
wire n_244;
wire n_173;
wire n_198;
wire n_447;
wire n_247;
wire n_314;
wire n_368;
wire n_433;
wire n_604;
wire n_321;
wire n_292;
wire n_625;
wire n_621;
wire n_455;
wire n_417;
wire n_612;
wire n_212;
wire n_385;
wire n_498;
wire n_516;
wire n_507;
wire n_497;
wire n_606;
wire n_559;
wire n_275;
wire n_640;
wire n_252;
wire n_624;
wire n_295;
wire n_330;
wire n_508;
wire n_506;
wire n_610;
wire n_509;
wire n_568;
wire n_147;
wire n_373;
wire n_307;
wire n_633;
wire n_530;
wire n_150;
wire n_439;
wire n_556;
wire n_209;
wire n_259;
wire n_448;
wire n_375;
wire n_301;
wire n_576;
wire n_186;
wire n_537;
wire n_191;
wire n_587;
wire n_492;
wire n_563;
wire n_171;
wire n_153;
wire n_524;
wire n_399;
wire n_341;
wire n_204;
wire n_394;
wire n_250;
wire n_579;
wire n_548;
wire n_543;
wire n_260;
wire n_298;
wire n_650;
wire n_320;
wire n_518;
wire n_505;
wire n_286;
wire n_282;
wire n_331;
wire n_406;
wire n_519;
wire n_470;
wire n_325;
wire n_449;
wire n_546;
wire n_281;
wire n_240;
wire n_381;
wire n_189;
wire n_220;
wire n_291;
wire n_231;
wire n_257;
wire n_390;
wire n_456;
wire n_371;
wire n_481;
wire n_535;
wire n_152;
wire n_540;
wire n_317;
wire n_618;
wire n_323;
wire n_569;
wire n_195;
wire n_356;
wire n_227;
wire n_592;
wire n_271;
wire n_335;
wire n_370;
wire n_167;
wire n_234;
wire n_343;
wire n_308;
wire n_428;
wire n_379;
wire n_267;
wire n_514;
wire n_457;
wire n_570;
wire n_297;
wire n_156;
wire n_603;
wire n_225;
wire n_377;
wire n_484;
wire n_219;
wire n_442;
wire n_157;
wire n_192;
wire n_636;
wire n_600;
wire n_223;
wire n_392;
wire n_158;
wire n_264;
wire n_472;
wire n_454;
wire n_387;
wire n_374;
wire n_163;
wire n_276;
wire n_339;
wire n_185;
wire n_183;
wire n_243;
wire n_398;
wire n_396;
wire n_635;
wire n_347;
wire n_169;
wire n_522;
wire n_550;
wire n_255;
wire n_215;
wire n_350;
wire n_196;
wire n_459;
wire n_646;
wire n_211;
wire n_218;
wire n_400;
wire n_181;
wire n_436;
wire n_290;
wire n_580;
wire n_221;
wire n_178;
wire n_622;
wire n_386;
wire n_578;
wire n_287;
wire n_344;
wire n_555;
wire n_473;
wire n_422;
wire n_475;
wire n_415;
wire n_485;
wire n_496;
wire n_355;
wire n_486;
wire n_336;
wire n_584;
wire n_591;
wire n_145;
wire n_521;
wire n_614;
wire n_337;
wire n_430;
wire n_313;
wire n_631;
wire n_479;
wire n_528;
wire n_510;
wire n_216;
wire n_168;
wire n_395;
wire n_164;
wire n_432;
wire n_553;
wire n_311;
wire n_208;
wire n_214;
wire n_328;
wire n_299;
wire n_303;
wire n_369;
wire n_296;
wire n_613;
wire n_241;
wire n_637;
wire n_357;
wire n_598;
wire n_608;
wire n_184;
wire n_446;
wire n_445;
wire n_165;
wire n_468;
wire n_499;
wire n_213;
wire n_342;
wire n_482;
wire n_517;
wire n_588;
wire n_361;
wire n_464;
wire n_363;
wire n_413;
wire n_402;
wire n_638;
wire n_197;
wire n_573;
wire n_236;
wire n_388;
wire n_249;
wire n_304;
wire n_329;
wire n_203;
wire n_274;
wire n_577;
wire n_384;
wire n_582;
wire n_460;
wire n_277;
wire n_338;
wire n_149;
wire n_477;
wire n_461;
wire n_333;
wire n_571;
wire n_309;
wire n_512;
wire n_462;
wire n_322;
wire n_567;
wire n_258;
wire n_652;
wire n_151;
wire n_306;
wire n_458;
wire n_288;
wire n_188;
wire n_190;
wire n_201;
wire n_263;
wire n_471;
wire n_609;
wire n_224;
wire n_228;
wire n_283;
wire n_383;
wire n_474;
wire n_542;
wire n_463;
wire n_488;
wire n_595;
wire n_502;
wire n_239;
wire n_466;
wire n_420;
wire n_630;
wire n_489;
wire n_632;
wire n_617;
wire n_310;
wire n_593;
wire n_504;
wire n_511;
wire n_586;
wire n_465;
wire n_358;
wire n_362;
wire n_170;
wire n_332;
wire n_161;
wire n_273;
wire n_349;
wire n_585;
wire n_270;
wire n_616;
wire n_230;
wire n_601;
wire n_279;
wire n_253;
wire n_261;
wire n_174;
wire n_289;
wire n_627;
wire n_206;
wire n_172;
wire n_217;
wire n_440;
wire n_478;
wire n_545;
wire n_441;
wire n_450;
wire n_648;
wire n_312;
wire n_476;
wire n_429;
wire n_534;
wire n_345;
wire n_210;
wire n_494;
wire n_641;
wire n_628;
wire n_365;
wire n_176;
wire n_557;
wire n_182;
wire n_354;
wire n_575;
wire n_607;
wire n_480;
wire n_647;
wire n_237;
wire n_425;
wire n_513;
wire n_407;
wire n_527;
wire n_180;
wire n_560;
wire n_340;
wire n_207;
wire n_561;
wire n_346;
wire n_393;
wire n_229;
wire n_495;
wire n_487;
wire n_602;
wire n_574;
wire n_437;
wire n_177;
wire n_453;
wire n_403;
wire n_421;
wire n_623;
wire n_405;
wire n_359;
wire n_490;
wire n_326;
wire n_233;
wire n_404;
wire n_205;
wire n_366;
wire n_572;
wire n_246;
wire n_596;
wire n_179;
wire n_410;
wire n_558;
wire n_269;
wire n_529;
wire n_285;
wire n_412;
wire n_232;
wire n_327;
wire n_644;
wire n_202;
wire n_266;
wire n_272;
wire n_491;
wire n_427;
wire n_193;
wire n_251;
wire n_352;
wire n_160;
wire n_565;
wire n_426;
wire n_566;
wire n_520;
wire n_409;
wire n_589;
wire n_597;
wire n_500;
wire n_562;
wire n_154;
wire n_148;
wire n_300;
wire n_651;
wire n_435;
wire n_159;
wire n_334;
wire n_599;
wire n_541;
wire n_391;
wire n_434;
wire n_645;
wire n_539;
wire n_175;
wire n_538;
wire n_262;
wire n_238;
wire n_639;
wire n_411;
wire n_414;
wire n_319;
wire n_364;
wire n_536;
wire n_531;
wire n_242;
wire n_360;
wire n_594;
wire n_200;
wire n_162;
wire n_222;
wire n_438;
wire n_324;
wire n_634;
wire n_416;
wire n_199;
wire n_187;
wire n_401;
wire n_348;
wire n_166;
wire n_626;
wire n_424;
wire n_256;
wire n_305;
wire n_533;
wire n_278;

CKINVDCx5p33_ASAP7_75t_R g145 ( 
.A(n_47),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_85),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_9),
.Y(n_147)
);

BUFx3_ASAP7_75t_L g148 ( 
.A(n_102),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_134),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_131),
.Y(n_150)
);

CKINVDCx5p33_ASAP7_75t_R g151 ( 
.A(n_83),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_101),
.Y(n_152)
);

BUFx2_ASAP7_75t_L g153 ( 
.A(n_71),
.Y(n_153)
);

INVxp67_ASAP7_75t_L g154 ( 
.A(n_110),
.Y(n_154)
);

INVx1_ASAP7_75t_SL g155 ( 
.A(n_32),
.Y(n_155)
);

CKINVDCx16_ASAP7_75t_R g156 ( 
.A(n_26),
.Y(n_156)
);

CKINVDCx5p33_ASAP7_75t_R g157 ( 
.A(n_133),
.Y(n_157)
);

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_95),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_55),
.Y(n_159)
);

CKINVDCx5p33_ASAP7_75t_R g160 ( 
.A(n_6),
.Y(n_160)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_144),
.Y(n_161)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_100),
.Y(n_162)
);

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_105),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_141),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_16),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_115),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_35),
.Y(n_167)
);

BUFx2_ASAP7_75t_L g168 ( 
.A(n_121),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_90),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_92),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_20),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_126),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_41),
.Y(n_173)
);

BUFx10_ASAP7_75t_L g174 ( 
.A(n_33),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_123),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_89),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_34),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_103),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_74),
.Y(n_179)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_112),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_117),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_21),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_13),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_7),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_4),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_120),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_53),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_3),
.Y(n_188)
);

BUFx10_ASAP7_75t_L g189 ( 
.A(n_29),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_136),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_107),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_49),
.Y(n_192)
);

INVx1_ASAP7_75t_SL g193 ( 
.A(n_63),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_130),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_78),
.Y(n_195)
);

INVx2_ASAP7_75t_SL g196 ( 
.A(n_142),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_81),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_138),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_48),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_22),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_40),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_76),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_111),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_37),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_31),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_7),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_5),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_109),
.Y(n_208)
);

INVx1_ASAP7_75t_SL g209 ( 
.A(n_98),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_2),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_66),
.Y(n_211)
);

BUFx6f_ASAP7_75t_L g212 ( 
.A(n_0),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_12),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_13),
.Y(n_214)
);

AND2x2_ASAP7_75t_L g215 ( 
.A(n_153),
.B(n_0),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_156),
.B(n_1),
.Y(n_216)
);

HB1xp67_ASAP7_75t_L g217 ( 
.A(n_147),
.Y(n_217)
);

AND2x4_ASAP7_75t_L g218 ( 
.A(n_148),
.B(n_1),
.Y(n_218)
);

INVx5_ASAP7_75t_L g219 ( 
.A(n_212),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_212),
.Y(n_220)
);

BUFx3_ASAP7_75t_L g221 ( 
.A(n_174),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_161),
.B(n_2),
.Y(n_222)
);

INVx5_ASAP7_75t_L g223 ( 
.A(n_212),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_161),
.B(n_3),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_212),
.B(n_4),
.Y(n_225)
);

BUFx3_ASAP7_75t_L g226 ( 
.A(n_174),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_168),
.B(n_5),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_185),
.Y(n_228)
);

BUFx6f_ASAP7_75t_L g229 ( 
.A(n_148),
.Y(n_229)
);

INVx6_ASAP7_75t_L g230 ( 
.A(n_189),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_189),
.B(n_6),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_162),
.B(n_8),
.Y(n_232)
);

AND2x2_ASAP7_75t_L g233 ( 
.A(n_196),
.B(n_8),
.Y(n_233)
);

INVx5_ASAP7_75t_L g234 ( 
.A(n_162),
.Y(n_234)
);

INVx5_ASAP7_75t_L g235 ( 
.A(n_180),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_146),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_180),
.B(n_9),
.Y(n_237)
);

BUFx12f_ASAP7_75t_L g238 ( 
.A(n_160),
.Y(n_238)
);

INVx5_ASAP7_75t_L g239 ( 
.A(n_183),
.Y(n_239)
);

BUFx2_ASAP7_75t_L g240 ( 
.A(n_206),
.Y(n_240)
);

BUFx2_ASAP7_75t_L g241 ( 
.A(n_207),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_SL g242 ( 
.A(n_184),
.B(n_10),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_154),
.B(n_10),
.Y(n_243)
);

INVx5_ASAP7_75t_L g244 ( 
.A(n_210),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_188),
.Y(n_245)
);

BUFx12f_ASAP7_75t_L g246 ( 
.A(n_213),
.Y(n_246)
);

INVx3_ASAP7_75t_L g247 ( 
.A(n_214),
.Y(n_247)
);

HB1xp67_ASAP7_75t_L g248 ( 
.A(n_159),
.Y(n_248)
);

AND2x4_ASAP7_75t_L g249 ( 
.A(n_164),
.B(n_11),
.Y(n_249)
);

AND2x2_ASAP7_75t_L g250 ( 
.A(n_155),
.B(n_193),
.Y(n_250)
);

INVx5_ASAP7_75t_L g251 ( 
.A(n_145),
.Y(n_251)
);

BUFx12f_ASAP7_75t_L g252 ( 
.A(n_151),
.Y(n_252)
);

HB1xp67_ASAP7_75t_L g253 ( 
.A(n_165),
.Y(n_253)
);

NOR2x1_ASAP7_75t_L g254 ( 
.A(n_167),
.B(n_14),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_SL g255 ( 
.A(n_149),
.B(n_209),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_171),
.B(n_11),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_173),
.B(n_12),
.Y(n_257)
);

AND2x4_ASAP7_75t_L g258 ( 
.A(n_195),
.B(n_15),
.Y(n_258)
);

BUFx6f_ASAP7_75t_L g259 ( 
.A(n_197),
.Y(n_259)
);

INVx5_ASAP7_75t_L g260 ( 
.A(n_157),
.Y(n_260)
);

BUFx12f_ASAP7_75t_L g261 ( 
.A(n_158),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_220),
.Y(n_262)
);

OA22x2_ASAP7_75t_L g263 ( 
.A1(n_248),
.A2(n_198),
.B1(n_201),
.B2(n_205),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_250),
.B(n_202),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_251),
.B(n_163),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_229),
.Y(n_266)
);

OAI22xp33_ASAP7_75t_L g267 ( 
.A1(n_242),
.A2(n_149),
.B1(n_150),
.B2(n_152),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_229),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_255),
.A2(n_166),
.B1(n_177),
.B2(n_178),
.Y(n_269)
);

INVx5_ASAP7_75t_L g270 ( 
.A(n_230),
.Y(n_270)
);

OAI22xp33_ASAP7_75t_SL g271 ( 
.A1(n_216),
.A2(n_211),
.B1(n_208),
.B2(n_204),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_255),
.A2(n_203),
.B1(n_200),
.B2(n_199),
.Y(n_272)
);

INVx2_ASAP7_75t_SL g273 ( 
.A(n_230),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_227),
.A2(n_181),
.B1(n_192),
.B2(n_191),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_215),
.A2(n_231),
.B1(n_246),
.B2(n_238),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_229),
.Y(n_276)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_219),
.Y(n_277)
);

OAI22xp33_ASAP7_75t_L g278 ( 
.A1(n_242),
.A2(n_194),
.B1(n_190),
.B2(n_187),
.Y(n_278)
);

OAI22xp33_ASAP7_75t_L g279 ( 
.A1(n_243),
.A2(n_186),
.B1(n_182),
.B2(n_179),
.Y(n_279)
);

AO22x2_ASAP7_75t_L g280 ( 
.A1(n_218),
.A2(n_176),
.B1(n_175),
.B2(n_172),
.Y(n_280)
);

NAND2xp33_ASAP7_75t_SL g281 ( 
.A(n_233),
.B(n_169),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_L g282 ( 
.A1(n_240),
.A2(n_241),
.B1(n_256),
.B2(n_257),
.Y(n_282)
);

AO22x2_ASAP7_75t_L g283 ( 
.A1(n_218),
.A2(n_170),
.B1(n_18),
.B2(n_19),
.Y(n_283)
);

OAI22xp33_ASAP7_75t_L g284 ( 
.A1(n_243),
.A2(n_17),
.B1(n_23),
.B2(n_24),
.Y(n_284)
);

AO22x2_ASAP7_75t_L g285 ( 
.A1(n_249),
.A2(n_224),
.B1(n_237),
.B2(n_232),
.Y(n_285)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_219),
.Y(n_286)
);

AO22x2_ASAP7_75t_L g287 ( 
.A1(n_249),
.A2(n_25),
.B1(n_27),
.B2(n_28),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_247),
.B(n_30),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_247),
.A2(n_36),
.B1(n_38),
.B2(n_39),
.Y(n_289)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_219),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g291 ( 
.A1(n_221),
.A2(n_42),
.B1(n_43),
.B2(n_44),
.Y(n_291)
);

AND2x2_ASAP7_75t_L g292 ( 
.A(n_226),
.B(n_45),
.Y(n_292)
);

AND2x2_ASAP7_75t_L g293 ( 
.A(n_239),
.B(n_46),
.Y(n_293)
);

AND2x2_ASAP7_75t_L g294 ( 
.A(n_239),
.B(n_50),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_252),
.A2(n_51),
.B1(n_52),
.B2(n_54),
.Y(n_295)
);

OR2x6_ASAP7_75t_L g296 ( 
.A(n_217),
.B(n_56),
.Y(n_296)
);

INVx2_ASAP7_75t_SL g297 ( 
.A(n_239),
.Y(n_297)
);

AO22x2_ASAP7_75t_L g298 ( 
.A1(n_222),
.A2(n_57),
.B1(n_58),
.B2(n_59),
.Y(n_298)
);

OAI22xp33_ASAP7_75t_SL g299 ( 
.A1(n_222),
.A2(n_60),
.B1(n_61),
.B2(n_62),
.Y(n_299)
);

OA22x2_ASAP7_75t_L g300 ( 
.A1(n_248),
.A2(n_64),
.B1(n_65),
.B2(n_67),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_L g301 ( 
.A1(n_261),
.A2(n_68),
.B1(n_69),
.B2(n_70),
.Y(n_301)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_223),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_SL g303 ( 
.A1(n_236),
.A2(n_72),
.B1(n_73),
.B2(n_75),
.Y(n_303)
);

OAI22xp33_ASAP7_75t_L g304 ( 
.A1(n_224),
.A2(n_77),
.B1(n_79),
.B2(n_80),
.Y(n_304)
);

BUFx10_ASAP7_75t_L g305 ( 
.A(n_228),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_245),
.Y(n_306)
);

OAI22xp33_ASAP7_75t_L g307 ( 
.A1(n_232),
.A2(n_237),
.B1(n_253),
.B2(n_217),
.Y(n_307)
);

OAI22xp33_ASAP7_75t_SL g308 ( 
.A1(n_253),
.A2(n_82),
.B1(n_84),
.B2(n_86),
.Y(n_308)
);

AND2x2_ASAP7_75t_L g309 ( 
.A(n_244),
.B(n_87),
.Y(n_309)
);

INVx2_ASAP7_75t_L g310 ( 
.A(n_223),
.Y(n_310)
);

OAI22xp33_ASAP7_75t_R g311 ( 
.A1(n_225),
.A2(n_244),
.B1(n_258),
.B2(n_254),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_L g312 ( 
.A1(n_258),
.A2(n_88),
.B1(n_91),
.B2(n_93),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_306),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_266),
.Y(n_314)
);

XOR2xp5_ASAP7_75t_L g315 ( 
.A(n_269),
.B(n_94),
.Y(n_315)
);

NOR2xp67_ASAP7_75t_L g316 ( 
.A(n_270),
.B(n_251),
.Y(n_316)
);

INVx2_ASAP7_75t_L g317 ( 
.A(n_262),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_268),
.Y(n_318)
);

AND2x2_ASAP7_75t_L g319 ( 
.A(n_270),
.B(n_244),
.Y(n_319)
);

AND2x2_ASAP7_75t_L g320 ( 
.A(n_264),
.B(n_260),
.Y(n_320)
);

INVxp33_ASAP7_75t_L g321 ( 
.A(n_282),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_276),
.Y(n_322)
);

XNOR2xp5_ASAP7_75t_L g323 ( 
.A(n_267),
.B(n_96),
.Y(n_323)
);

INVx3_ASAP7_75t_L g324 ( 
.A(n_277),
.Y(n_324)
);

AND2x2_ASAP7_75t_SL g325 ( 
.A(n_312),
.B(n_225),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_275),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g327 ( 
.A(n_272),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_305),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_285),
.B(n_235),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_286),
.Y(n_330)
);

AND2x2_ASAP7_75t_SL g331 ( 
.A(n_288),
.B(n_259),
.Y(n_331)
);

AOI21xp5_ASAP7_75t_L g332 ( 
.A1(n_285),
.A2(n_235),
.B(n_234),
.Y(n_332)
);

INVxp33_ASAP7_75t_SL g333 ( 
.A(n_274),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_278),
.B(n_260),
.Y(n_334)
);

AND2x2_ASAP7_75t_L g335 ( 
.A(n_273),
.B(n_297),
.Y(n_335)
);

INVx2_ASAP7_75t_SL g336 ( 
.A(n_263),
.Y(n_336)
);

AND2x2_ASAP7_75t_L g337 ( 
.A(n_292),
.B(n_296),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_290),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_302),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_310),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_265),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_300),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_293),
.Y(n_343)
);

BUFx6f_ASAP7_75t_L g344 ( 
.A(n_294),
.Y(n_344)
);

CKINVDCx20_ASAP7_75t_R g345 ( 
.A(n_296),
.Y(n_345)
);

INVx2_ASAP7_75t_SL g346 ( 
.A(n_280),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_309),
.Y(n_347)
);

AND2x4_ASAP7_75t_SL g348 ( 
.A(n_295),
.B(n_259),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_298),
.Y(n_349)
);

XOR2xp5_ASAP7_75t_L g350 ( 
.A(n_280),
.B(n_97),
.Y(n_350)
);

XOR2xp5_ASAP7_75t_L g351 ( 
.A(n_283),
.B(n_99),
.Y(n_351)
);

INVxp67_ASAP7_75t_SL g352 ( 
.A(n_307),
.Y(n_352)
);

AND2x4_ASAP7_75t_L g353 ( 
.A(n_291),
.B(n_260),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_298),
.Y(n_354)
);

AND2x4_ASAP7_75t_L g355 ( 
.A(n_301),
.B(n_251),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_289),
.Y(n_356)
);

OR2x2_ASAP7_75t_L g357 ( 
.A(n_281),
.B(n_259),
.Y(n_357)
);

INVx2_ASAP7_75t_L g358 ( 
.A(n_287),
.Y(n_358)
);

INVxp33_ASAP7_75t_L g359 ( 
.A(n_283),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_271),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_287),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_308),
.Y(n_362)
);

AND2x2_ASAP7_75t_L g363 ( 
.A(n_311),
.B(n_235),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_299),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_303),
.Y(n_365)
);

NOR2xp33_ASAP7_75t_SL g366 ( 
.A(n_284),
.B(n_234),
.Y(n_366)
);

INVx2_ASAP7_75t_L g367 ( 
.A(n_304),
.Y(n_367)
);

CKINVDCx20_ASAP7_75t_R g368 ( 
.A(n_279),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_306),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_306),
.Y(n_370)
);

INVx2_ASAP7_75t_L g371 ( 
.A(n_262),
.Y(n_371)
);

AND2x2_ASAP7_75t_L g372 ( 
.A(n_270),
.B(n_234),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_306),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_306),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_306),
.Y(n_375)
);

AND2x4_ASAP7_75t_L g376 ( 
.A(n_296),
.B(n_104),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_306),
.Y(n_377)
);

AND2x2_ASAP7_75t_L g378 ( 
.A(n_342),
.B(n_106),
.Y(n_378)
);

AND2x2_ASAP7_75t_L g379 ( 
.A(n_343),
.B(n_108),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_331),
.B(n_347),
.Y(n_380)
);

INVx2_ASAP7_75t_L g381 ( 
.A(n_317),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_313),
.Y(n_382)
);

INVx2_ASAP7_75t_SL g383 ( 
.A(n_357),
.Y(n_383)
);

AND2x2_ASAP7_75t_L g384 ( 
.A(n_352),
.B(n_113),
.Y(n_384)
);

AND2x2_ASAP7_75t_SL g385 ( 
.A(n_325),
.B(n_114),
.Y(n_385)
);

INVx2_ASAP7_75t_SL g386 ( 
.A(n_329),
.Y(n_386)
);

BUFx3_ASAP7_75t_L g387 ( 
.A(n_369),
.Y(n_387)
);

INVx2_ASAP7_75t_SL g388 ( 
.A(n_329),
.Y(n_388)
);

HB1xp67_ASAP7_75t_L g389 ( 
.A(n_336),
.Y(n_389)
);

INVx4_ASAP7_75t_L g390 ( 
.A(n_344),
.Y(n_390)
);

INVx2_ASAP7_75t_L g391 ( 
.A(n_371),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_370),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_373),
.Y(n_393)
);

AND2x2_ASAP7_75t_L g394 ( 
.A(n_352),
.B(n_116),
.Y(n_394)
);

AND2x4_ASAP7_75t_L g395 ( 
.A(n_376),
.B(n_118),
.Y(n_395)
);

INVx2_ASAP7_75t_L g396 ( 
.A(n_374),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_331),
.B(n_119),
.Y(n_397)
);

INVx2_ASAP7_75t_L g398 ( 
.A(n_375),
.Y(n_398)
);

INVx2_ASAP7_75t_L g399 ( 
.A(n_377),
.Y(n_399)
);

INVx2_ASAP7_75t_SL g400 ( 
.A(n_335),
.Y(n_400)
);

AND2x4_ASAP7_75t_L g401 ( 
.A(n_376),
.B(n_339),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_344),
.B(n_122),
.Y(n_402)
);

INVx2_ASAP7_75t_L g403 ( 
.A(n_330),
.Y(n_403)
);

AND2x2_ASAP7_75t_L g404 ( 
.A(n_325),
.B(n_124),
.Y(n_404)
);

AND2x2_ASAP7_75t_L g405 ( 
.A(n_337),
.B(n_125),
.Y(n_405)
);

AND2x2_ASAP7_75t_L g406 ( 
.A(n_367),
.B(n_127),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_338),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_340),
.Y(n_408)
);

HB1xp67_ASAP7_75t_L g409 ( 
.A(n_346),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_344),
.B(n_128),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_314),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_SL g412 ( 
.A(n_341),
.B(n_129),
.Y(n_412)
);

AND2x4_ASAP7_75t_L g413 ( 
.A(n_324),
.B(n_132),
.Y(n_413)
);

INVx1_ASAP7_75t_SL g414 ( 
.A(n_328),
.Y(n_414)
);

AND2x2_ASAP7_75t_L g415 ( 
.A(n_363),
.B(n_364),
.Y(n_415)
);

AND2x4_ASAP7_75t_L g416 ( 
.A(n_324),
.B(n_143),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_318),
.Y(n_417)
);

INVx2_ASAP7_75t_L g418 ( 
.A(n_322),
.Y(n_418)
);

OAI21xp5_ASAP7_75t_L g419 ( 
.A1(n_362),
.A2(n_135),
.B(n_137),
.Y(n_419)
);

OAI21xp5_ASAP7_75t_L g420 ( 
.A1(n_334),
.A2(n_356),
.B(n_332),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_344),
.Y(n_421)
);

INVx1_ASAP7_75t_SL g422 ( 
.A(n_360),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_320),
.B(n_139),
.Y(n_423)
);

AND2x2_ASAP7_75t_L g424 ( 
.A(n_358),
.B(n_140),
.Y(n_424)
);

INVx3_ASAP7_75t_L g425 ( 
.A(n_353),
.Y(n_425)
);

OAI21xp5_ASAP7_75t_L g426 ( 
.A1(n_334),
.A2(n_332),
.B(n_354),
.Y(n_426)
);

OAI21xp5_ASAP7_75t_L g427 ( 
.A1(n_349),
.A2(n_333),
.B(n_359),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_348),
.B(n_353),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_361),
.Y(n_429)
);

AND2x4_ASAP7_75t_L g430 ( 
.A(n_355),
.B(n_365),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_323),
.Y(n_431)
);

INVxp67_ASAP7_75t_L g432 ( 
.A(n_315),
.Y(n_432)
);

NOR2xp33_ASAP7_75t_L g433 ( 
.A(n_321),
.B(n_368),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_355),
.B(n_366),
.Y(n_434)
);

AND2x2_ASAP7_75t_L g435 ( 
.A(n_359),
.B(n_321),
.Y(n_435)
);

INVx2_ASAP7_75t_L g436 ( 
.A(n_372),
.Y(n_436)
);

NOR2xp33_ASAP7_75t_SL g437 ( 
.A(n_326),
.B(n_368),
.Y(n_437)
);

HB1xp67_ASAP7_75t_L g438 ( 
.A(n_351),
.Y(n_438)
);

AND2x2_ASAP7_75t_L g439 ( 
.A(n_319),
.B(n_366),
.Y(n_439)
);

INVx3_ASAP7_75t_L g440 ( 
.A(n_350),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_L g441 ( 
.A(n_316),
.B(n_327),
.Y(n_441)
);

NOR2xp33_ASAP7_75t_L g442 ( 
.A(n_380),
.B(n_327),
.Y(n_442)
);

AND2x4_ASAP7_75t_L g443 ( 
.A(n_401),
.B(n_387),
.Y(n_443)
);

BUFx6f_ASAP7_75t_L g444 ( 
.A(n_401),
.Y(n_444)
);

BUFx3_ASAP7_75t_L g445 ( 
.A(n_389),
.Y(n_445)
);

INVx6_ASAP7_75t_L g446 ( 
.A(n_413),
.Y(n_446)
);

BUFx6f_ASAP7_75t_L g447 ( 
.A(n_401),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_411),
.Y(n_448)
);

AND2x2_ASAP7_75t_L g449 ( 
.A(n_435),
.B(n_345),
.Y(n_449)
);

NOR2xp33_ASAP7_75t_L g450 ( 
.A(n_435),
.B(n_326),
.Y(n_450)
);

INVx2_ASAP7_75t_L g451 ( 
.A(n_396),
.Y(n_451)
);

AND2x2_ASAP7_75t_SL g452 ( 
.A(n_385),
.B(n_345),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_411),
.Y(n_453)
);

NAND2x1p5_ASAP7_75t_L g454 ( 
.A(n_390),
.B(n_395),
.Y(n_454)
);

NAND2x1p5_ASAP7_75t_L g455 ( 
.A(n_390),
.B(n_395),
.Y(n_455)
);

AND2x4_ASAP7_75t_L g456 ( 
.A(n_387),
.B(n_425),
.Y(n_456)
);

AND2x4_ASAP7_75t_L g457 ( 
.A(n_425),
.B(n_430),
.Y(n_457)
);

BUFx3_ASAP7_75t_L g458 ( 
.A(n_409),
.Y(n_458)
);

BUFx2_ASAP7_75t_L g459 ( 
.A(n_430),
.Y(n_459)
);

NAND2x1p5_ASAP7_75t_L g460 ( 
.A(n_390),
.B(n_395),
.Y(n_460)
);

BUFx6f_ASAP7_75t_L g461 ( 
.A(n_413),
.Y(n_461)
);

OR2x6_ASAP7_75t_L g462 ( 
.A(n_430),
.B(n_428),
.Y(n_462)
);

BUFx8_ASAP7_75t_SL g463 ( 
.A(n_440),
.Y(n_463)
);

BUFx12f_ASAP7_75t_L g464 ( 
.A(n_415),
.Y(n_464)
);

INVx2_ASAP7_75t_L g465 ( 
.A(n_396),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_417),
.Y(n_466)
);

AND2x4_ASAP7_75t_L g467 ( 
.A(n_425),
.B(n_386),
.Y(n_467)
);

OR2x6_ASAP7_75t_L g468 ( 
.A(n_404),
.B(n_386),
.Y(n_468)
);

BUFx12f_ASAP7_75t_L g469 ( 
.A(n_415),
.Y(n_469)
);

HB1xp67_ASAP7_75t_L g470 ( 
.A(n_429),
.Y(n_470)
);

NOR2xp33_ASAP7_75t_SL g471 ( 
.A(n_385),
.B(n_419),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_L g472 ( 
.A(n_406),
.B(n_420),
.Y(n_472)
);

NOR2x1_ASAP7_75t_SL g473 ( 
.A(n_421),
.B(n_397),
.Y(n_473)
);

INVx2_ASAP7_75t_L g474 ( 
.A(n_398),
.Y(n_474)
);

NOR2xp33_ASAP7_75t_SL g475 ( 
.A(n_404),
.B(n_394),
.Y(n_475)
);

AND2x2_ASAP7_75t_L g476 ( 
.A(n_414),
.B(n_433),
.Y(n_476)
);

NOR2xp33_ASAP7_75t_L g477 ( 
.A(n_384),
.B(n_394),
.Y(n_477)
);

INVx3_ASAP7_75t_L g478 ( 
.A(n_421),
.Y(n_478)
);

BUFx4f_ASAP7_75t_L g479 ( 
.A(n_384),
.Y(n_479)
);

OR2x6_ASAP7_75t_L g480 ( 
.A(n_388),
.B(n_427),
.Y(n_480)
);

AND2x2_ASAP7_75t_L g481 ( 
.A(n_431),
.B(n_383),
.Y(n_481)
);

AND2x2_ASAP7_75t_L g482 ( 
.A(n_431),
.B(n_383),
.Y(n_482)
);

INVx2_ASAP7_75t_L g483 ( 
.A(n_398),
.Y(n_483)
);

BUFx4f_ASAP7_75t_L g484 ( 
.A(n_405),
.Y(n_484)
);

AND2x4_ASAP7_75t_L g485 ( 
.A(n_388),
.B(n_392),
.Y(n_485)
);

INVx3_ASAP7_75t_SL g486 ( 
.A(n_449),
.Y(n_486)
);

INVx4_ASAP7_75t_L g487 ( 
.A(n_461),
.Y(n_487)
);

BUFx8_ASAP7_75t_L g488 ( 
.A(n_464),
.Y(n_488)
);

BUFx3_ASAP7_75t_L g489 ( 
.A(n_469),
.Y(n_489)
);

NAND2x1p5_ASAP7_75t_L g490 ( 
.A(n_461),
.B(n_406),
.Y(n_490)
);

BUFx3_ASAP7_75t_L g491 ( 
.A(n_445),
.Y(n_491)
);

INVx3_ASAP7_75t_L g492 ( 
.A(n_461),
.Y(n_492)
);

INVx2_ASAP7_75t_L g493 ( 
.A(n_478),
.Y(n_493)
);

BUFx3_ASAP7_75t_L g494 ( 
.A(n_458),
.Y(n_494)
);

CKINVDCx5p33_ASAP7_75t_R g495 ( 
.A(n_463),
.Y(n_495)
);

AND2x4_ASAP7_75t_L g496 ( 
.A(n_457),
.B(n_405),
.Y(n_496)
);

OR2x2_ASAP7_75t_L g497 ( 
.A(n_476),
.B(n_422),
.Y(n_497)
);

AND2x2_ASAP7_75t_L g498 ( 
.A(n_477),
.B(n_378),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_470),
.Y(n_499)
);

BUFx6f_ASAP7_75t_L g500 ( 
.A(n_446),
.Y(n_500)
);

BUFx8_ASAP7_75t_L g501 ( 
.A(n_459),
.Y(n_501)
);

CKINVDCx5p33_ASAP7_75t_R g502 ( 
.A(n_463),
.Y(n_502)
);

BUFx3_ASAP7_75t_L g503 ( 
.A(n_457),
.Y(n_503)
);

INVx3_ASAP7_75t_L g504 ( 
.A(n_446),
.Y(n_504)
);

INVx2_ASAP7_75t_L g505 ( 
.A(n_451),
.Y(n_505)
);

NOR2xp33_ASAP7_75t_L g506 ( 
.A(n_442),
.B(n_477),
.Y(n_506)
);

BUFx2_ASAP7_75t_SL g507 ( 
.A(n_443),
.Y(n_507)
);

INVx2_ASAP7_75t_L g508 ( 
.A(n_465),
.Y(n_508)
);

CKINVDCx5p33_ASAP7_75t_R g509 ( 
.A(n_450),
.Y(n_509)
);

INVx3_ASAP7_75t_SL g510 ( 
.A(n_480),
.Y(n_510)
);

BUFx4_ASAP7_75t_SL g511 ( 
.A(n_480),
.Y(n_511)
);

INVx4_ASAP7_75t_L g512 ( 
.A(n_446),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_470),
.Y(n_513)
);

INVx1_ASAP7_75t_SL g514 ( 
.A(n_481),
.Y(n_514)
);

AOI22xp33_ASAP7_75t_L g515 ( 
.A1(n_506),
.A2(n_471),
.B1(n_452),
.B2(n_442),
.Y(n_515)
);

INVx2_ASAP7_75t_SL g516 ( 
.A(n_491),
.Y(n_516)
);

CKINVDCx5p33_ASAP7_75t_R g517 ( 
.A(n_495),
.Y(n_517)
);

BUFx6f_ASAP7_75t_L g518 ( 
.A(n_503),
.Y(n_518)
);

INVx2_ASAP7_75t_L g519 ( 
.A(n_493),
.Y(n_519)
);

INVx2_ASAP7_75t_L g520 ( 
.A(n_493),
.Y(n_520)
);

INVxp67_ASAP7_75t_SL g521 ( 
.A(n_490),
.Y(n_521)
);

CKINVDCx11_ASAP7_75t_R g522 ( 
.A(n_486),
.Y(n_522)
);

CKINVDCx5p33_ASAP7_75t_R g523 ( 
.A(n_495),
.Y(n_523)
);

BUFx8_ASAP7_75t_L g524 ( 
.A(n_491),
.Y(n_524)
);

AND2x2_ASAP7_75t_L g525 ( 
.A(n_514),
.B(n_450),
.Y(n_525)
);

CKINVDCx20_ASAP7_75t_R g526 ( 
.A(n_502),
.Y(n_526)
);

CKINVDCx20_ASAP7_75t_R g527 ( 
.A(n_502),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_499),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_513),
.Y(n_529)
);

OAI22x1_ASAP7_75t_L g530 ( 
.A1(n_509),
.A2(n_440),
.B1(n_438),
.B2(n_453),
.Y(n_530)
);

AOI22xp33_ASAP7_75t_L g531 ( 
.A1(n_498),
.A2(n_471),
.B1(n_479),
.B2(n_475),
.Y(n_531)
);

INVx5_ASAP7_75t_L g532 ( 
.A(n_500),
.Y(n_532)
);

INVx2_ASAP7_75t_L g533 ( 
.A(n_505),
.Y(n_533)
);

CKINVDCx11_ASAP7_75t_R g534 ( 
.A(n_486),
.Y(n_534)
);

AND2x2_ASAP7_75t_L g535 ( 
.A(n_497),
.B(n_482),
.Y(n_535)
);

OAI22xp5_ASAP7_75t_L g536 ( 
.A1(n_498),
.A2(n_479),
.B1(n_484),
.B2(n_472),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_505),
.Y(n_537)
);

INVx2_ASAP7_75t_L g538 ( 
.A(n_508),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_508),
.Y(n_539)
);

AOI22xp33_ASAP7_75t_L g540 ( 
.A1(n_497),
.A2(n_475),
.B1(n_480),
.B2(n_484),
.Y(n_540)
);

CKINVDCx6p67_ASAP7_75t_R g541 ( 
.A(n_494),
.Y(n_541)
);

INVx2_ASAP7_75t_SL g542 ( 
.A(n_524),
.Y(n_542)
);

HB1xp67_ASAP7_75t_L g543 ( 
.A(n_528),
.Y(n_543)
);

OAI21xp33_ASAP7_75t_L g544 ( 
.A1(n_515),
.A2(n_437),
.B(n_509),
.Y(n_544)
);

AOI22xp33_ASAP7_75t_L g545 ( 
.A1(n_525),
.A2(n_412),
.B1(n_472),
.B2(n_510),
.Y(n_545)
);

OAI21xp33_ASAP7_75t_SL g546 ( 
.A1(n_531),
.A2(n_426),
.B(n_379),
.Y(n_546)
);

CKINVDCx5p33_ASAP7_75t_R g547 ( 
.A(n_523),
.Y(n_547)
);

INVx2_ASAP7_75t_L g548 ( 
.A(n_533),
.Y(n_548)
);

HB1xp67_ASAP7_75t_L g549 ( 
.A(n_529),
.Y(n_549)
);

CKINVDCx6p67_ASAP7_75t_R g550 ( 
.A(n_541),
.Y(n_550)
);

AND2x2_ASAP7_75t_SL g551 ( 
.A(n_540),
.B(n_496),
.Y(n_551)
);

OAI22xp5_ASAP7_75t_L g552 ( 
.A1(n_535),
.A2(n_468),
.B1(n_490),
.B2(n_510),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_L g553 ( 
.A(n_516),
.B(n_485),
.Y(n_553)
);

BUFx6f_ASAP7_75t_L g554 ( 
.A(n_518),
.Y(n_554)
);

OAI22xp33_ASAP7_75t_L g555 ( 
.A1(n_530),
.A2(n_468),
.B1(n_448),
.B2(n_466),
.Y(n_555)
);

INVx2_ASAP7_75t_L g556 ( 
.A(n_533),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_537),
.Y(n_557)
);

OAI21xp5_ASAP7_75t_SL g558 ( 
.A1(n_536),
.A2(n_440),
.B(n_432),
.Y(n_558)
);

OAI22xp5_ASAP7_75t_L g559 ( 
.A1(n_521),
.A2(n_468),
.B1(n_490),
.B2(n_455),
.Y(n_559)
);

AOI22xp33_ASAP7_75t_SL g560 ( 
.A1(n_524),
.A2(n_501),
.B1(n_434),
.B2(n_488),
.Y(n_560)
);

AOI22xp33_ASAP7_75t_L g561 ( 
.A1(n_522),
.A2(n_496),
.B1(n_379),
.B2(n_462),
.Y(n_561)
);

AOI22xp33_ASAP7_75t_L g562 ( 
.A1(n_522),
.A2(n_496),
.B1(n_462),
.B2(n_399),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_539),
.Y(n_563)
);

AOI22xp33_ASAP7_75t_L g564 ( 
.A1(n_534),
.A2(n_462),
.B1(n_399),
.B2(n_393),
.Y(n_564)
);

AOI22xp33_ASAP7_75t_SL g565 ( 
.A1(n_524),
.A2(n_501),
.B1(n_488),
.B2(n_439),
.Y(n_565)
);

BUFx4f_ASAP7_75t_SL g566 ( 
.A(n_526),
.Y(n_566)
);

AOI22xp33_ASAP7_75t_L g567 ( 
.A1(n_534),
.A2(n_392),
.B1(n_393),
.B2(n_439),
.Y(n_567)
);

OAI22xp5_ASAP7_75t_L g568 ( 
.A1(n_518),
.A2(n_454),
.B1(n_460),
.B2(n_455),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_538),
.Y(n_569)
);

AOI22xp5_ASAP7_75t_L g570 ( 
.A1(n_526),
.A2(n_441),
.B1(n_443),
.B2(n_456),
.Y(n_570)
);

BUFx12f_ASAP7_75t_L g571 ( 
.A(n_517),
.Y(n_571)
);

BUFx12f_ASAP7_75t_L g572 ( 
.A(n_517),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_543),
.Y(n_573)
);

AOI22xp33_ASAP7_75t_L g574 ( 
.A1(n_544),
.A2(n_417),
.B1(n_418),
.B2(n_485),
.Y(n_574)
);

AOI22xp33_ASAP7_75t_L g575 ( 
.A1(n_551),
.A2(n_403),
.B1(n_456),
.B2(n_474),
.Y(n_575)
);

OAI221xp5_ASAP7_75t_L g576 ( 
.A1(n_558),
.A2(n_382),
.B1(n_489),
.B2(n_407),
.C(n_408),
.Y(n_576)
);

AOI22xp33_ASAP7_75t_L g577 ( 
.A1(n_555),
.A2(n_403),
.B1(n_483),
.B2(n_444),
.Y(n_577)
);

OAI22xp5_ASAP7_75t_L g578 ( 
.A1(n_567),
.A2(n_454),
.B1(n_460),
.B2(n_507),
.Y(n_578)
);

AOI22xp33_ASAP7_75t_L g579 ( 
.A1(n_546),
.A2(n_378),
.B1(n_381),
.B2(n_391),
.Y(n_579)
);

OAI221xp5_ASAP7_75t_L g580 ( 
.A1(n_570),
.A2(n_561),
.B1(n_545),
.B2(n_564),
.C(n_562),
.Y(n_580)
);

AOI22xp33_ASAP7_75t_L g581 ( 
.A1(n_555),
.A2(n_447),
.B1(n_444),
.B2(n_423),
.Y(n_581)
);

AOI22xp33_ASAP7_75t_L g582 ( 
.A1(n_552),
.A2(n_447),
.B1(n_444),
.B2(n_518),
.Y(n_582)
);

OAI22xp5_ASAP7_75t_L g583 ( 
.A1(n_565),
.A2(n_489),
.B1(n_518),
.B2(n_527),
.Y(n_583)
);

AND2x2_ASAP7_75t_L g584 ( 
.A(n_543),
.B(n_519),
.Y(n_584)
);

OAI222xp33_ASAP7_75t_L g585 ( 
.A1(n_565),
.A2(n_560),
.B1(n_566),
.B2(n_542),
.C1(n_553),
.C2(n_559),
.Y(n_585)
);

INVx2_ASAP7_75t_L g586 ( 
.A(n_548),
.Y(n_586)
);

AOI22xp5_ASAP7_75t_L g587 ( 
.A1(n_560),
.A2(n_527),
.B1(n_488),
.B2(n_447),
.Y(n_587)
);

AOI22xp33_ASAP7_75t_L g588 ( 
.A1(n_549),
.A2(n_416),
.B1(n_413),
.B2(n_391),
.Y(n_588)
);

AOI22xp33_ASAP7_75t_L g589 ( 
.A1(n_549),
.A2(n_416),
.B1(n_381),
.B2(n_424),
.Y(n_589)
);

AND2x2_ASAP7_75t_L g590 ( 
.A(n_554),
.B(n_520),
.Y(n_590)
);

AOI22xp33_ASAP7_75t_L g591 ( 
.A1(n_571),
.A2(n_572),
.B1(n_416),
.B2(n_424),
.Y(n_591)
);

OAI22xp5_ASAP7_75t_L g592 ( 
.A1(n_550),
.A2(n_494),
.B1(n_492),
.B2(n_512),
.Y(n_592)
);

AOI22xp33_ASAP7_75t_L g593 ( 
.A1(n_557),
.A2(n_500),
.B1(n_504),
.B2(n_492),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_L g594 ( 
.A(n_556),
.B(n_538),
.Y(n_594)
);

AND2x2_ASAP7_75t_L g595 ( 
.A(n_584),
.B(n_554),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_L g596 ( 
.A(n_573),
.B(n_563),
.Y(n_596)
);

NAND3xp33_ASAP7_75t_L g597 ( 
.A(n_576),
.B(n_574),
.C(n_580),
.Y(n_597)
);

AND2x2_ASAP7_75t_L g598 ( 
.A(n_590),
.B(n_554),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_L g599 ( 
.A(n_586),
.B(n_569),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_L g600 ( 
.A(n_594),
.B(n_519),
.Y(n_600)
);

OAI21xp5_ASAP7_75t_SL g601 ( 
.A1(n_585),
.A2(n_568),
.B(n_511),
.Y(n_601)
);

AND2x2_ASAP7_75t_L g602 ( 
.A(n_582),
.B(n_520),
.Y(n_602)
);

OA211x2_ASAP7_75t_L g603 ( 
.A1(n_579),
.A2(n_402),
.B(n_410),
.C(n_473),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_L g604 ( 
.A(n_574),
.B(n_547),
.Y(n_604)
);

AND2x2_ASAP7_75t_L g605 ( 
.A(n_583),
.B(n_532),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_L g606 ( 
.A(n_579),
.B(n_532),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_L g607 ( 
.A(n_581),
.B(n_532),
.Y(n_607)
);

AND2x2_ASAP7_75t_L g608 ( 
.A(n_587),
.B(n_532),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_L g609 ( 
.A(n_596),
.B(n_577),
.Y(n_609)
);

AOI22xp33_ASAP7_75t_L g610 ( 
.A1(n_597),
.A2(n_591),
.B1(n_589),
.B2(n_575),
.Y(n_610)
);

AND2x2_ASAP7_75t_L g611 ( 
.A(n_595),
.B(n_593),
.Y(n_611)
);

AO21x2_ASAP7_75t_L g612 ( 
.A1(n_596),
.A2(n_592),
.B(n_578),
.Y(n_612)
);

AOI22xp5_ASAP7_75t_SL g613 ( 
.A1(n_608),
.A2(n_487),
.B1(n_500),
.B2(n_512),
.Y(n_613)
);

NAND3xp33_ASAP7_75t_L g614 ( 
.A(n_601),
.B(n_588),
.C(n_532),
.Y(n_614)
);

BUFx3_ASAP7_75t_L g615 ( 
.A(n_598),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_599),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_616),
.Y(n_617)
);

AND2x4_ASAP7_75t_L g618 ( 
.A(n_615),
.B(n_605),
.Y(n_618)
);

NOR3xp33_ASAP7_75t_L g619 ( 
.A(n_614),
.B(n_604),
.C(n_607),
.Y(n_619)
);

NAND4xp75_ASAP7_75t_L g620 ( 
.A(n_609),
.B(n_603),
.C(n_602),
.D(n_607),
.Y(n_620)
);

NOR2xp33_ASAP7_75t_L g621 ( 
.A(n_615),
.B(n_600),
.Y(n_621)
);

INVx2_ASAP7_75t_L g622 ( 
.A(n_612),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_L g623 ( 
.A(n_612),
.B(n_606),
.Y(n_623)
);

HB1xp67_ASAP7_75t_L g624 ( 
.A(n_622),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_617),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_623),
.Y(n_626)
);

INVx2_ASAP7_75t_L g627 ( 
.A(n_618),
.Y(n_627)
);

XOR2x2_ASAP7_75t_L g628 ( 
.A(n_620),
.B(n_611),
.Y(n_628)
);

HB1xp67_ASAP7_75t_L g629 ( 
.A(n_625),
.Y(n_629)
);

INVx2_ASAP7_75t_SL g630 ( 
.A(n_627),
.Y(n_630)
);

INVx2_ASAP7_75t_L g631 ( 
.A(n_624),
.Y(n_631)
);

INVx1_ASAP7_75t_SL g632 ( 
.A(n_628),
.Y(n_632)
);

INVx1_ASAP7_75t_SL g633 ( 
.A(n_626),
.Y(n_633)
);

INVx1_ASAP7_75t_SL g634 ( 
.A(n_632),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_629),
.Y(n_635)
);

CKINVDCx16_ASAP7_75t_R g636 ( 
.A(n_632),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_635),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_634),
.Y(n_638)
);

INVxp67_ASAP7_75t_L g639 ( 
.A(n_638),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_639),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_640),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_L g642 ( 
.A(n_641),
.B(n_636),
.Y(n_642)
);

AND2x2_ASAP7_75t_L g643 ( 
.A(n_642),
.B(n_637),
.Y(n_643)
);

AOI211xp5_ASAP7_75t_L g644 ( 
.A1(n_643),
.A2(n_633),
.B(n_631),
.C(n_619),
.Y(n_644)
);

HB1xp67_ASAP7_75t_L g645 ( 
.A(n_644),
.Y(n_645)
);

AOI22xp5_ASAP7_75t_L g646 ( 
.A1(n_645),
.A2(n_630),
.B1(n_624),
.B2(n_618),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_646),
.Y(n_647)
);

OAI22xp5_ASAP7_75t_L g648 ( 
.A1(n_647),
.A2(n_610),
.B1(n_621),
.B2(n_613),
.Y(n_648)
);

AOI22xp5_ASAP7_75t_L g649 ( 
.A1(n_647),
.A2(n_400),
.B1(n_610),
.B2(n_429),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_649),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_648),
.Y(n_651)
);

AOI221xp5_ASAP7_75t_L g652 ( 
.A1(n_651),
.A2(n_400),
.B1(n_467),
.B2(n_436),
.C(n_500),
.Y(n_652)
);

AOI211xp5_ASAP7_75t_L g653 ( 
.A1(n_652),
.A2(n_650),
.B(n_467),
.C(n_436),
.Y(n_653)
);


endmodule