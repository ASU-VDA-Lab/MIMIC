module fake_netlist_6_1671_n_1952 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_161, n_68, n_166, n_28, n_184, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_178, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_180, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_181, n_76, n_36, n_182, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_175, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_104, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_173, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_35, n_183, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_171, n_31, n_57, n_169, n_53, n_51, n_44, n_56, n_1952);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_161;
input n_68;
input n_166;
input n_28;
input n_184;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_178;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_175;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_104;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_173;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_35;
input n_183;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_171;
input n_31;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1952;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_1853;
wire n_783;
wire n_1738;
wire n_798;
wire n_188;
wire n_1575;
wire n_1854;
wire n_1923;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1691;
wire n_1688;
wire n_1009;
wire n_1743;
wire n_1930;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_1844;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_1786;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_200;
wire n_447;
wire n_1803;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1867;
wire n_1704;
wire n_1078;
wire n_544;
wire n_250;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1903;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_616;
wire n_658;
wire n_1874;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1902;
wire n_1842;
wire n_1620;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1798;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_1820;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_1936;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_1894;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_1815;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1911;
wire n_1644;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_1918;
wire n_577;
wire n_1843;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1909;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_1907;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1762;
wire n_1910;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1876;
wire n_1895;
wire n_1697;
wire n_243;
wire n_979;
wire n_1873;
wire n_905;
wire n_1866;
wire n_1680;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1865;
wire n_1875;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_1950;
wire n_530;
wire n_1563;
wire n_1912;
wire n_277;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_1760;
wire n_1927;
wire n_210;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1926;
wire n_1175;
wire n_328;
wire n_1386;
wire n_1896;
wire n_429;
wire n_1747;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1802;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_1801;
wire n_1886;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_1813;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_1709;
wire n_1825;
wire n_1757;
wire n_1796;
wire n_1792;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_462;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_297;
wire n_595;
wire n_627;
wire n_1767;
wire n_1779;
wire n_524;
wire n_1465;
wire n_342;
wire n_1858;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1932;
wire n_1101;
wire n_1026;
wire n_1880;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_1839;
wire n_685;
wire n_1765;
wire n_353;
wire n_605;
wire n_1514;
wire n_1863;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_851;
wire n_682;
wire n_305;
wire n_996;
wire n_532;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_1913;
wire n_510;
wire n_837;
wire n_1488;
wire n_1808;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_1947;
wire n_536;
wire n_1788;
wire n_622;
wire n_1469;
wire n_1838;
wire n_1835;
wire n_1766;
wire n_1776;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_1771;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_1878;
wire n_899;
wire n_189;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_1577;
wire n_1181;
wire n_1822;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_1817;
wire n_927;
wire n_1849;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_552;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_216;
wire n_912;
wire n_1857;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_755;
wire n_1021;
wire n_931;
wire n_474;
wire n_527;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_1897;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_1942;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_1837;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_211;
wire n_1483;
wire n_1834;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_1787;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1919;
wire n_1080;
wire n_723;
wire n_1877;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1939;
wire n_1769;
wire n_1220;
wire n_1893;
wire n_556;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_1951;
wire n_444;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1773;
wire n_1775;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_1745;
wire n_914;
wire n_759;
wire n_1831;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_1901;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1892;
wire n_1933;
wire n_1135;
wire n_1179;
wire n_1169;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1917;
wire n_1580;
wire n_1425;
wire n_1881;
wire n_1281;
wire n_1267;
wire n_1806;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_1855;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_1832;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1594;
wire n_664;
wire n_1869;
wire n_1764;
wire n_1429;
wire n_1610;
wire n_1889;
wire n_435;
wire n_1905;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_1937;
wire n_465;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_186;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1934;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_1871;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_1859;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_1916;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1852;
wire n_1024;
wire n_1768;
wire n_198;
wire n_1847;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1841;
wire n_1639;
wire n_1623;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1818;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1686;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1943;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1938;
wire n_1262;
wire n_218;
wire n_1891;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_1870;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1827;
wire n_1361;
wire n_1864;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_370;
wire n_1695;
wire n_1828;
wire n_650;
wire n_1046;
wire n_1940;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1883;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_1823;
wire n_227;
wire n_1720;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_1795;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1845;
wire n_1489;
wire n_942;
wire n_1524;
wire n_543;
wire n_1920;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1946;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_1846;
wire n_533;
wire n_806;
wire n_959;
wire n_879;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_1782;
wire n_282;
wire n_1676;
wire n_833;
wire n_1830;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_1900;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_1086;
wire n_1066;
wire n_1948;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1906;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_1758;
wire n_1925;
wire n_737;
wire n_1318;
wire n_1914;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1373;
wire n_1292;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_1931;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_1941;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1794;
wire n_1236;
wire n_1559;
wire n_1725;
wire n_1928;
wire n_1872;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1746;
wire n_1325;
wire n_1002;
wire n_1741;
wire n_1949;
wire n_545;
wire n_489;
wire n_1804;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1860;
wire n_1904;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1908;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_187;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1800;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_1826;
wire n_566;
wire n_1023;
wire n_1882;
wire n_1118;
wire n_1076;
wire n_194;
wire n_1007;
wire n_1807;
wire n_1929;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1814;
wire n_1631;
wire n_591;
wire n_1377;
wire n_1879;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_680;
wire n_367;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1824;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_1810;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_1729;
wire n_669;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1785;
wire n_763;
wire n_1147;
wire n_1848;
wire n_360;
wire n_1754;
wire n_1506;
wire n_1652;
wire n_1812;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_1173;
wire n_1924;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_1174;
wire n_1944;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_1945;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_1922;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1821;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_185;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1525;
wire n_455;
wire n_1585;
wire n_1851;
wire n_363;
wire n_1799;
wire n_1090;
wire n_592;
wire n_1816;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_1829;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_1789;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1921;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_271;
wire n_404;
wire n_1884;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1819;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_1861;
wire n_373;
wire n_1632;
wire n_1890;
wire n_1805;
wire n_257;
wire n_1557;
wire n_1888;
wire n_1833;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_1850;
wire n_1898;
wire n_1868;
wire n_207;
wire n_1089;
wire n_1887;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_1836;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1899;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_1862;
wire n_1856;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_540;
wire n_1423;
wire n_1935;
wire n_457;
wire n_364;
wire n_1915;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_827;
wire n_531;
wire n_361;
wire n_1025;
wire n_336;
wire n_1885;
wire n_1013;
wire n_1259;
wire n_192;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

CKINVDCx16_ASAP7_75t_R g185 ( 
.A(n_38),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_42),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_117),
.Y(n_187)
);

BUFx6f_ASAP7_75t_L g188 ( 
.A(n_150),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_26),
.Y(n_189)
);

INVx1_ASAP7_75t_SL g190 ( 
.A(n_153),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_90),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_15),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_63),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_109),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_55),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_100),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_102),
.Y(n_197)
);

INVx3_ASAP7_75t_L g198 ( 
.A(n_51),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_38),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_111),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_34),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_15),
.Y(n_202)
);

BUFx6f_ASAP7_75t_L g203 ( 
.A(n_177),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_162),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_16),
.Y(n_205)
);

BUFx6f_ASAP7_75t_L g206 ( 
.A(n_91),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_95),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_53),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_152),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_48),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_69),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_74),
.Y(n_212)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_182),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_61),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_25),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_136),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_104),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_4),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_18),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_72),
.Y(n_220)
);

BUFx10_ASAP7_75t_L g221 ( 
.A(n_98),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_42),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_40),
.Y(n_223)
);

CKINVDCx16_ASAP7_75t_R g224 ( 
.A(n_6),
.Y(n_224)
);

INVxp67_ASAP7_75t_L g225 ( 
.A(n_130),
.Y(n_225)
);

BUFx6f_ASAP7_75t_L g226 ( 
.A(n_143),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_169),
.Y(n_227)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_39),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_26),
.Y(n_229)
);

BUFx10_ASAP7_75t_L g230 ( 
.A(n_87),
.Y(n_230)
);

BUFx3_ASAP7_75t_L g231 ( 
.A(n_166),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_184),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_59),
.Y(n_233)
);

BUFx3_ASAP7_75t_L g234 ( 
.A(n_140),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_7),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_171),
.Y(n_236)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_92),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_56),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_19),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_81),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_16),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_125),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_88),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_138),
.Y(n_244)
);

BUFx3_ASAP7_75t_L g245 ( 
.A(n_178),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_149),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_34),
.Y(n_247)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_137),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_103),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_39),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_160),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_148),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_124),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_58),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_146),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_28),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_122),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_49),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_101),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_57),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_37),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_1),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_25),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_52),
.Y(n_264)
);

HB1xp67_ASAP7_75t_L g265 ( 
.A(n_76),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_181),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_179),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_6),
.Y(n_268)
);

BUFx3_ASAP7_75t_L g269 ( 
.A(n_64),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_51),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_133),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_18),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_65),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_119),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_99),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_47),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_155),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_144),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_142),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_110),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_29),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_7),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_52),
.Y(n_283)
);

BUFx2_ASAP7_75t_L g284 ( 
.A(n_112),
.Y(n_284)
);

INVxp67_ASAP7_75t_L g285 ( 
.A(n_129),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_56),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_172),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_163),
.Y(n_288)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_126),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_24),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_131),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_156),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_49),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_79),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_31),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_145),
.Y(n_296)
);

INVxp67_ASAP7_75t_L g297 ( 
.A(n_94),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_154),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_97),
.Y(n_299)
);

INVx2_ASAP7_75t_L g300 ( 
.A(n_55),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_13),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_24),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_40),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_45),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_70),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_151),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_176),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_157),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_108),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_107),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_5),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_13),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_75),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_120),
.Y(n_314)
);

BUFx10_ASAP7_75t_L g315 ( 
.A(n_17),
.Y(n_315)
);

INVxp67_ASAP7_75t_L g316 ( 
.A(n_36),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_141),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_71),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_173),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_29),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_58),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g322 ( 
.A(n_57),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g323 ( 
.A(n_73),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_158),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_0),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_47),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_89),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g328 ( 
.A(n_165),
.Y(n_328)
);

BUFx3_ASAP7_75t_L g329 ( 
.A(n_83),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_44),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_32),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_167),
.Y(n_332)
);

INVxp67_ASAP7_75t_L g333 ( 
.A(n_50),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_3),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_32),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_82),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_105),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_20),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_86),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_175),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_23),
.Y(n_341)
);

BUFx10_ASAP7_75t_L g342 ( 
.A(n_50),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_132),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_35),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_19),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_11),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_164),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_84),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_65),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_33),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_64),
.Y(n_351)
);

CKINVDCx20_ASAP7_75t_R g352 ( 
.A(n_63),
.Y(n_352)
);

CKINVDCx20_ASAP7_75t_R g353 ( 
.A(n_183),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_161),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_5),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_48),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_54),
.Y(n_357)
);

BUFx3_ASAP7_75t_L g358 ( 
.A(n_2),
.Y(n_358)
);

CKINVDCx20_ASAP7_75t_R g359 ( 
.A(n_31),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_21),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_23),
.Y(n_361)
);

INVx1_ASAP7_75t_SL g362 ( 
.A(n_159),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_106),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_62),
.Y(n_364)
);

BUFx10_ASAP7_75t_L g365 ( 
.A(n_128),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_35),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_96),
.Y(n_367)
);

BUFx3_ASAP7_75t_L g368 ( 
.A(n_22),
.Y(n_368)
);

INVxp67_ASAP7_75t_L g369 ( 
.A(n_192),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_187),
.Y(n_370)
);

CKINVDCx20_ASAP7_75t_R g371 ( 
.A(n_209),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_191),
.Y(n_372)
);

CKINVDCx20_ASAP7_75t_R g373 ( 
.A(n_252),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_198),
.Y(n_374)
);

INVxp33_ASAP7_75t_SL g375 ( 
.A(n_186),
.Y(n_375)
);

CKINVDCx16_ASAP7_75t_R g376 ( 
.A(n_185),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_194),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_196),
.Y(n_378)
);

INVxp67_ASAP7_75t_L g379 ( 
.A(n_192),
.Y(n_379)
);

CKINVDCx20_ASAP7_75t_R g380 ( 
.A(n_323),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_197),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_200),
.Y(n_382)
);

CKINVDCx20_ASAP7_75t_R g383 ( 
.A(n_328),
.Y(n_383)
);

NOR2xp67_ASAP7_75t_L g384 ( 
.A(n_198),
.B(n_0),
.Y(n_384)
);

INVxp67_ASAP7_75t_SL g385 ( 
.A(n_265),
.Y(n_385)
);

CKINVDCx20_ASAP7_75t_R g386 ( 
.A(n_353),
.Y(n_386)
);

XNOR2xp5_ASAP7_75t_L g387 ( 
.A(n_199),
.B(n_1),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_204),
.Y(n_388)
);

INVxp33_ASAP7_75t_SL g389 ( 
.A(n_189),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_198),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_228),
.Y(n_391)
);

INVxp67_ASAP7_75t_L g392 ( 
.A(n_195),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_228),
.Y(n_393)
);

CKINVDCx20_ASAP7_75t_R g394 ( 
.A(n_207),
.Y(n_394)
);

INVx2_ASAP7_75t_L g395 ( 
.A(n_300),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_212),
.Y(n_396)
);

INVxp67_ASAP7_75t_SL g397 ( 
.A(n_284),
.Y(n_397)
);

CKINVDCx20_ASAP7_75t_R g398 ( 
.A(n_216),
.Y(n_398)
);

CKINVDCx16_ASAP7_75t_R g399 ( 
.A(n_185),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_217),
.Y(n_400)
);

CKINVDCx20_ASAP7_75t_R g401 ( 
.A(n_240),
.Y(n_401)
);

NOR2xp67_ASAP7_75t_L g402 ( 
.A(n_300),
.B(n_2),
.Y(n_402)
);

NOR2xp33_ASAP7_75t_L g403 ( 
.A(n_284),
.B(n_3),
.Y(n_403)
);

NOR2xp33_ASAP7_75t_L g404 ( 
.A(n_227),
.B(n_4),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_195),
.Y(n_405)
);

NOR2xp67_ASAP7_75t_L g406 ( 
.A(n_316),
.B(n_8),
.Y(n_406)
);

NOR2xp33_ASAP7_75t_L g407 ( 
.A(n_227),
.B(n_8),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_211),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_211),
.Y(n_409)
);

INVxp67_ASAP7_75t_L g410 ( 
.A(n_214),
.Y(n_410)
);

CKINVDCx20_ASAP7_75t_R g411 ( 
.A(n_242),
.Y(n_411)
);

INVxp67_ASAP7_75t_SL g412 ( 
.A(n_231),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_214),
.Y(n_413)
);

CKINVDCx20_ASAP7_75t_R g414 ( 
.A(n_246),
.Y(n_414)
);

CKINVDCx20_ASAP7_75t_R g415 ( 
.A(n_249),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_222),
.Y(n_416)
);

INVx2_ASAP7_75t_L g417 ( 
.A(n_232),
.Y(n_417)
);

NOR2xp67_ASAP7_75t_L g418 ( 
.A(n_333),
.B(n_9),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_251),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_222),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_233),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_259),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_267),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_271),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_233),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_238),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_238),
.Y(n_427)
);

HB1xp67_ASAP7_75t_L g428 ( 
.A(n_224),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_239),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_239),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_247),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_247),
.Y(n_432)
);

INVx2_ASAP7_75t_L g433 ( 
.A(n_232),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_256),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_274),
.Y(n_435)
);

HB1xp67_ASAP7_75t_L g436 ( 
.A(n_224),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_256),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_258),
.Y(n_438)
);

HB1xp67_ASAP7_75t_L g439 ( 
.A(n_193),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_258),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_262),
.Y(n_441)
);

BUFx2_ASAP7_75t_L g442 ( 
.A(n_269),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_275),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_277),
.Y(n_444)
);

BUFx6f_ASAP7_75t_L g445 ( 
.A(n_188),
.Y(n_445)
);

CKINVDCx20_ASAP7_75t_R g446 ( 
.A(n_278),
.Y(n_446)
);

NOR2xp33_ASAP7_75t_L g447 ( 
.A(n_236),
.B(n_9),
.Y(n_447)
);

NOR2xp33_ASAP7_75t_L g448 ( 
.A(n_236),
.B(n_10),
.Y(n_448)
);

CKINVDCx5p33_ASAP7_75t_R g449 ( 
.A(n_279),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_262),
.Y(n_450)
);

INVxp67_ASAP7_75t_L g451 ( 
.A(n_264),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_264),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_272),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_272),
.Y(n_454)
);

INVx2_ASAP7_75t_L g455 ( 
.A(n_243),
.Y(n_455)
);

CKINVDCx5p33_ASAP7_75t_R g456 ( 
.A(n_280),
.Y(n_456)
);

INVxp33_ASAP7_75t_SL g457 ( 
.A(n_201),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_273),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_273),
.Y(n_459)
);

CKINVDCx20_ASAP7_75t_R g460 ( 
.A(n_287),
.Y(n_460)
);

BUFx6f_ASAP7_75t_L g461 ( 
.A(n_445),
.Y(n_461)
);

NOR2xp33_ASAP7_75t_L g462 ( 
.A(n_403),
.B(n_225),
.Y(n_462)
);

CKINVDCx5p33_ASAP7_75t_R g463 ( 
.A(n_370),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_417),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_417),
.Y(n_465)
);

NOR2xp33_ASAP7_75t_L g466 ( 
.A(n_397),
.B(n_285),
.Y(n_466)
);

AND2x4_ASAP7_75t_L g467 ( 
.A(n_384),
.B(n_231),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_L g468 ( 
.A(n_412),
.B(n_291),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_374),
.B(n_296),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_433),
.Y(n_470)
);

NAND2xp33_ASAP7_75t_L g471 ( 
.A(n_433),
.B(n_188),
.Y(n_471)
);

INVx2_ASAP7_75t_L g472 ( 
.A(n_445),
.Y(n_472)
);

AND2x2_ASAP7_75t_L g473 ( 
.A(n_455),
.B(n_234),
.Y(n_473)
);

AND2x4_ASAP7_75t_L g474 ( 
.A(n_384),
.B(n_234),
.Y(n_474)
);

BUFx6f_ASAP7_75t_L g475 ( 
.A(n_445),
.Y(n_475)
);

INVx3_ASAP7_75t_L g476 ( 
.A(n_445),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_395),
.Y(n_477)
);

INVx2_ASAP7_75t_L g478 ( 
.A(n_445),
.Y(n_478)
);

INVx3_ASAP7_75t_L g479 ( 
.A(n_445),
.Y(n_479)
);

INVx2_ASAP7_75t_L g480 ( 
.A(n_455),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_395),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_L g482 ( 
.A(n_374),
.B(n_309),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_L g483 ( 
.A(n_390),
.B(n_313),
.Y(n_483)
);

BUFx6f_ASAP7_75t_L g484 ( 
.A(n_390),
.Y(n_484)
);

INVx2_ASAP7_75t_L g485 ( 
.A(n_391),
.Y(n_485)
);

INVx2_ASAP7_75t_L g486 ( 
.A(n_391),
.Y(n_486)
);

BUFx6f_ASAP7_75t_L g487 ( 
.A(n_393),
.Y(n_487)
);

OAI21x1_ASAP7_75t_L g488 ( 
.A1(n_405),
.A2(n_237),
.B(n_213),
.Y(n_488)
);

INVx2_ASAP7_75t_L g489 ( 
.A(n_393),
.Y(n_489)
);

BUFx2_ASAP7_75t_L g490 ( 
.A(n_428),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_405),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_408),
.Y(n_492)
);

NOR2xp33_ASAP7_75t_L g493 ( 
.A(n_375),
.B(n_297),
.Y(n_493)
);

NOR2xp33_ASAP7_75t_SL g494 ( 
.A(n_376),
.B(n_315),
.Y(n_494)
);

INVxp67_ASAP7_75t_L g495 ( 
.A(n_436),
.Y(n_495)
);

AND2x2_ASAP7_75t_L g496 ( 
.A(n_442),
.B(n_245),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_408),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_409),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_409),
.Y(n_499)
);

OAI21x1_ASAP7_75t_L g500 ( 
.A1(n_413),
.A2(n_237),
.B(n_213),
.Y(n_500)
);

OAI21x1_ASAP7_75t_L g501 ( 
.A1(n_413),
.A2(n_289),
.B(n_248),
.Y(n_501)
);

OAI21x1_ASAP7_75t_L g502 ( 
.A1(n_416),
.A2(n_289),
.B(n_248),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_L g503 ( 
.A(n_404),
.B(n_314),
.Y(n_503)
);

INVx2_ASAP7_75t_L g504 ( 
.A(n_416),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_420),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_420),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_L g507 ( 
.A(n_407),
.B(n_319),
.Y(n_507)
);

INVx3_ASAP7_75t_L g508 ( 
.A(n_421),
.Y(n_508)
);

BUFx3_ASAP7_75t_L g509 ( 
.A(n_421),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_425),
.Y(n_510)
);

AND2x4_ASAP7_75t_L g511 ( 
.A(n_402),
.B(n_245),
.Y(n_511)
);

INVx2_ASAP7_75t_L g512 ( 
.A(n_425),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_426),
.Y(n_513)
);

BUFx6f_ASAP7_75t_L g514 ( 
.A(n_426),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_447),
.B(n_324),
.Y(n_515)
);

AND2x4_ASAP7_75t_L g516 ( 
.A(n_402),
.B(n_329),
.Y(n_516)
);

AND2x2_ASAP7_75t_L g517 ( 
.A(n_442),
.B(n_329),
.Y(n_517)
);

INVx3_ASAP7_75t_L g518 ( 
.A(n_427),
.Y(n_518)
);

INVx2_ASAP7_75t_L g519 ( 
.A(n_427),
.Y(n_519)
);

NOR2xp33_ASAP7_75t_L g520 ( 
.A(n_389),
.B(n_457),
.Y(n_520)
);

INVx2_ASAP7_75t_L g521 ( 
.A(n_429),
.Y(n_521)
);

INVx2_ASAP7_75t_L g522 ( 
.A(n_429),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_L g523 ( 
.A(n_448),
.B(n_332),
.Y(n_523)
);

INVx3_ASAP7_75t_L g524 ( 
.A(n_430),
.Y(n_524)
);

BUFx12f_ASAP7_75t_L g525 ( 
.A(n_372),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_430),
.Y(n_526)
);

INVxp67_ASAP7_75t_L g527 ( 
.A(n_439),
.Y(n_527)
);

CKINVDCx5p33_ASAP7_75t_R g528 ( 
.A(n_377),
.Y(n_528)
);

INVx2_ASAP7_75t_L g529 ( 
.A(n_431),
.Y(n_529)
);

HB1xp67_ASAP7_75t_L g530 ( 
.A(n_418),
.Y(n_530)
);

NAND2xp33_ASAP7_75t_L g531 ( 
.A(n_431),
.B(n_188),
.Y(n_531)
);

INVx2_ASAP7_75t_L g532 ( 
.A(n_432),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_432),
.Y(n_533)
);

INVx2_ASAP7_75t_L g534 ( 
.A(n_434),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_434),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_437),
.Y(n_536)
);

CKINVDCx20_ASAP7_75t_R g537 ( 
.A(n_371),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_437),
.Y(n_538)
);

CKINVDCx5p33_ASAP7_75t_R g539 ( 
.A(n_378),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_SL g540 ( 
.A(n_462),
.B(n_381),
.Y(n_540)
);

NOR2xp33_ASAP7_75t_L g541 ( 
.A(n_462),
.B(n_382),
.Y(n_541)
);

INVx2_ASAP7_75t_L g542 ( 
.A(n_480),
.Y(n_542)
);

INVx4_ASAP7_75t_L g543 ( 
.A(n_461),
.Y(n_543)
);

BUFx3_ASAP7_75t_L g544 ( 
.A(n_509),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_509),
.Y(n_545)
);

NOR2xp33_ASAP7_75t_L g546 ( 
.A(n_503),
.B(n_388),
.Y(n_546)
);

AND2x2_ASAP7_75t_L g547 ( 
.A(n_530),
.B(n_385),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_L g548 ( 
.A(n_468),
.B(n_467),
.Y(n_548)
);

BUFx4f_ASAP7_75t_L g549 ( 
.A(n_514),
.Y(n_549)
);

INVx2_ASAP7_75t_L g550 ( 
.A(n_480),
.Y(n_550)
);

BUFx3_ASAP7_75t_L g551 ( 
.A(n_509),
.Y(n_551)
);

BUFx6f_ASAP7_75t_L g552 ( 
.A(n_461),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_L g553 ( 
.A(n_468),
.B(n_396),
.Y(n_553)
);

INVx2_ASAP7_75t_L g554 ( 
.A(n_480),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_509),
.Y(n_555)
);

INVx2_ASAP7_75t_L g556 ( 
.A(n_480),
.Y(n_556)
);

INVx2_ASAP7_75t_L g557 ( 
.A(n_485),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_491),
.Y(n_558)
);

OR2x6_ASAP7_75t_L g559 ( 
.A(n_525),
.B(n_418),
.Y(n_559)
);

INVx2_ASAP7_75t_L g560 ( 
.A(n_485),
.Y(n_560)
);

INVx2_ASAP7_75t_L g561 ( 
.A(n_514),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_L g562 ( 
.A(n_467),
.B(n_400),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_SL g563 ( 
.A(n_520),
.B(n_419),
.Y(n_563)
);

OR2x2_ASAP7_75t_L g564 ( 
.A(n_490),
.B(n_376),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_491),
.Y(n_565)
);

AND2x2_ASAP7_75t_L g566 ( 
.A(n_530),
.B(n_438),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_491),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_492),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_SL g569 ( 
.A(n_520),
.B(n_422),
.Y(n_569)
);

BUFx4f_ASAP7_75t_L g570 ( 
.A(n_514),
.Y(n_570)
);

NAND2xp33_ASAP7_75t_SL g571 ( 
.A(n_490),
.B(n_460),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_SL g572 ( 
.A(n_493),
.B(n_423),
.Y(n_572)
);

BUFx2_ASAP7_75t_L g573 ( 
.A(n_490),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_492),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_492),
.Y(n_575)
);

AOI22xp33_ASAP7_75t_L g576 ( 
.A1(n_503),
.A2(n_269),
.B1(n_368),
.B2(n_358),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_497),
.Y(n_577)
);

INVxp33_ASAP7_75t_L g578 ( 
.A(n_496),
.Y(n_578)
);

INVx2_ASAP7_75t_L g579 ( 
.A(n_514),
.Y(n_579)
);

AO21x2_ASAP7_75t_L g580 ( 
.A1(n_488),
.A2(n_501),
.B(n_500),
.Y(n_580)
);

NAND2xp5_ASAP7_75t_SL g581 ( 
.A(n_493),
.B(n_424),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_497),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_497),
.Y(n_583)
);

INVx1_ASAP7_75t_SL g584 ( 
.A(n_537),
.Y(n_584)
);

OAI22xp33_ASAP7_75t_L g585 ( 
.A1(n_494),
.A2(n_399),
.B1(n_406),
.B2(n_202),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_498),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_498),
.Y(n_587)
);

INVxp33_ASAP7_75t_L g588 ( 
.A(n_496),
.Y(n_588)
);

NAND3xp33_ASAP7_75t_L g589 ( 
.A(n_466),
.B(n_379),
.C(n_369),
.Y(n_589)
);

AND2x6_ASAP7_75t_L g590 ( 
.A(n_467),
.B(n_188),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_498),
.Y(n_591)
);

INVx4_ASAP7_75t_L g592 ( 
.A(n_461),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_505),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_L g594 ( 
.A(n_467),
.B(n_435),
.Y(n_594)
);

AOI22xp33_ASAP7_75t_L g595 ( 
.A1(n_507),
.A2(n_358),
.B1(n_368),
.B2(n_304),
.Y(n_595)
);

INVx2_ASAP7_75t_L g596 ( 
.A(n_514),
.Y(n_596)
);

AND2x2_ASAP7_75t_L g597 ( 
.A(n_473),
.B(n_438),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_505),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_L g599 ( 
.A(n_467),
.B(n_443),
.Y(n_599)
);

NAND3xp33_ASAP7_75t_L g600 ( 
.A(n_466),
.B(n_410),
.C(n_392),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_505),
.Y(n_601)
);

INVx2_ASAP7_75t_L g602 ( 
.A(n_514),
.Y(n_602)
);

NOR2xp33_ASAP7_75t_L g603 ( 
.A(n_507),
.B(n_444),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_506),
.Y(n_604)
);

OAI22xp5_ASAP7_75t_L g605 ( 
.A1(n_515),
.A2(n_394),
.B1(n_398),
.B2(n_446),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_506),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_L g607 ( 
.A(n_467),
.B(n_449),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_L g608 ( 
.A(n_474),
.B(n_456),
.Y(n_608)
);

INVx2_ASAP7_75t_SL g609 ( 
.A(n_496),
.Y(n_609)
);

AOI22xp33_ASAP7_75t_L g610 ( 
.A1(n_515),
.A2(n_523),
.B1(n_474),
.B2(n_517),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_506),
.Y(n_611)
);

CKINVDCx5p33_ASAP7_75t_R g612 ( 
.A(n_463),
.Y(n_612)
);

CKINVDCx5p33_ASAP7_75t_R g613 ( 
.A(n_528),
.Y(n_613)
);

INVx1_ASAP7_75t_SL g614 ( 
.A(n_537),
.Y(n_614)
);

INVx2_ASAP7_75t_L g615 ( 
.A(n_514),
.Y(n_615)
);

INVx3_ASAP7_75t_L g616 ( 
.A(n_461),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_L g617 ( 
.A(n_474),
.B(n_190),
.Y(n_617)
);

BUFx6f_ASAP7_75t_L g618 ( 
.A(n_461),
.Y(n_618)
);

AOI22xp33_ASAP7_75t_L g619 ( 
.A1(n_523),
.A2(n_344),
.B1(n_311),
.B2(n_304),
.Y(n_619)
);

NOR2xp33_ASAP7_75t_L g620 ( 
.A(n_527),
.B(n_401),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_SL g621 ( 
.A(n_494),
.B(n_399),
.Y(n_621)
);

CKINVDCx16_ASAP7_75t_R g622 ( 
.A(n_525),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_SL g623 ( 
.A(n_527),
.B(n_411),
.Y(n_623)
);

NOR2xp33_ASAP7_75t_L g624 ( 
.A(n_539),
.B(n_414),
.Y(n_624)
);

INVx3_ASAP7_75t_L g625 ( 
.A(n_461),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_L g626 ( 
.A(n_474),
.B(n_362),
.Y(n_626)
);

INVx2_ASAP7_75t_L g627 ( 
.A(n_485),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_510),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_L g629 ( 
.A(n_474),
.B(n_337),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_510),
.Y(n_630)
);

BUFx6f_ASAP7_75t_L g631 ( 
.A(n_461),
.Y(n_631)
);

INVx2_ASAP7_75t_L g632 ( 
.A(n_486),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_510),
.Y(n_633)
);

INVx2_ASAP7_75t_L g634 ( 
.A(n_486),
.Y(n_634)
);

INVxp67_ASAP7_75t_SL g635 ( 
.A(n_476),
.Y(n_635)
);

NOR2xp33_ASAP7_75t_L g636 ( 
.A(n_469),
.B(n_415),
.Y(n_636)
);

INVx2_ASAP7_75t_L g637 ( 
.A(n_486),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_513),
.Y(n_638)
);

AND2x2_ASAP7_75t_L g639 ( 
.A(n_473),
.B(n_517),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_513),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_513),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_526),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_L g643 ( 
.A(n_474),
.B(n_339),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_L g644 ( 
.A(n_469),
.B(n_340),
.Y(n_644)
);

INVx2_ASAP7_75t_L g645 ( 
.A(n_514),
.Y(n_645)
);

INVx2_ASAP7_75t_L g646 ( 
.A(n_514),
.Y(n_646)
);

OAI21xp33_ASAP7_75t_SL g647 ( 
.A1(n_488),
.A2(n_305),
.B(n_295),
.Y(n_647)
);

INVx3_ASAP7_75t_L g648 ( 
.A(n_461),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_L g649 ( 
.A(n_482),
.B(n_348),
.Y(n_649)
);

INVx2_ASAP7_75t_L g650 ( 
.A(n_486),
.Y(n_650)
);

BUFx2_ASAP7_75t_L g651 ( 
.A(n_495),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_526),
.Y(n_652)
);

CKINVDCx5p33_ASAP7_75t_R g653 ( 
.A(n_525),
.Y(n_653)
);

NOR2xp33_ASAP7_75t_L g654 ( 
.A(n_482),
.B(n_373),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_526),
.Y(n_655)
);

BUFx6f_ASAP7_75t_L g656 ( 
.A(n_461),
.Y(n_656)
);

INVxp67_ASAP7_75t_SL g657 ( 
.A(n_476),
.Y(n_657)
);

INVx2_ASAP7_75t_L g658 ( 
.A(n_489),
.Y(n_658)
);

INVx2_ASAP7_75t_L g659 ( 
.A(n_489),
.Y(n_659)
);

CKINVDCx14_ASAP7_75t_R g660 ( 
.A(n_525),
.Y(n_660)
);

AOI22xp33_ASAP7_75t_L g661 ( 
.A1(n_517),
.A2(n_305),
.B1(n_311),
.B2(n_318),
.Y(n_661)
);

BUFx6f_ASAP7_75t_L g662 ( 
.A(n_475),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_535),
.Y(n_663)
);

INVx2_ASAP7_75t_L g664 ( 
.A(n_489),
.Y(n_664)
);

AOI22xp33_ASAP7_75t_L g665 ( 
.A1(n_511),
.A2(n_318),
.B1(n_325),
.B2(n_331),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_535),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_535),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_L g668 ( 
.A(n_483),
.B(n_354),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_SL g669 ( 
.A(n_495),
.B(n_221),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_L g670 ( 
.A(n_483),
.B(n_511),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_L g671 ( 
.A(n_511),
.B(n_363),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_536),
.Y(n_672)
);

NOR2xp33_ASAP7_75t_L g673 ( 
.A(n_536),
.B(n_380),
.Y(n_673)
);

INVxp33_ASAP7_75t_L g674 ( 
.A(n_473),
.Y(n_674)
);

INVx2_ASAP7_75t_L g675 ( 
.A(n_487),
.Y(n_675)
);

XOR2xp5_ASAP7_75t_SL g676 ( 
.A(n_499),
.B(n_243),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_536),
.Y(n_677)
);

INVx2_ASAP7_75t_L g678 ( 
.A(n_487),
.Y(n_678)
);

INVx5_ASAP7_75t_L g679 ( 
.A(n_475),
.Y(n_679)
);

BUFx10_ASAP7_75t_L g680 ( 
.A(n_511),
.Y(n_680)
);

AOI22xp33_ASAP7_75t_L g681 ( 
.A1(n_511),
.A2(n_516),
.B1(n_524),
.B2(n_518),
.Y(n_681)
);

INVx2_ASAP7_75t_L g682 ( 
.A(n_489),
.Y(n_682)
);

BUFx6f_ASAP7_75t_L g683 ( 
.A(n_475),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_538),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_SL g685 ( 
.A(n_511),
.B(n_221),
.Y(n_685)
);

BUFx6f_ASAP7_75t_L g686 ( 
.A(n_475),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_L g687 ( 
.A(n_516),
.B(n_244),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_538),
.Y(n_688)
);

AOI22xp33_ASAP7_75t_L g689 ( 
.A1(n_516),
.A2(n_295),
.B1(n_325),
.B2(n_331),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_538),
.Y(n_690)
);

NOR2xp33_ASAP7_75t_L g691 ( 
.A(n_499),
.B(n_383),
.Y(n_691)
);

OR2x2_ASAP7_75t_L g692 ( 
.A(n_564),
.B(n_387),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_545),
.Y(n_693)
);

INVx2_ASAP7_75t_L g694 ( 
.A(n_558),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_L g695 ( 
.A(n_546),
.B(n_516),
.Y(n_695)
);

AOI22xp5_ASAP7_75t_L g696 ( 
.A1(n_603),
.A2(n_541),
.B1(n_636),
.B2(n_654),
.Y(n_696)
);

NOR2xp67_ASAP7_75t_L g697 ( 
.A(n_620),
.B(n_533),
.Y(n_697)
);

INVx2_ASAP7_75t_L g698 ( 
.A(n_558),
.Y(n_698)
);

NOR2xp33_ASAP7_75t_L g699 ( 
.A(n_540),
.B(n_386),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_L g700 ( 
.A(n_610),
.B(n_516),
.Y(n_700)
);

AND2x2_ASAP7_75t_L g701 ( 
.A(n_639),
.B(n_508),
.Y(n_701)
);

BUFx8_ASAP7_75t_L g702 ( 
.A(n_573),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_L g703 ( 
.A(n_548),
.B(n_516),
.Y(n_703)
);

NOR2xp33_ASAP7_75t_L g704 ( 
.A(n_578),
.B(n_205),
.Y(n_704)
);

NOR2xp33_ASAP7_75t_L g705 ( 
.A(n_588),
.B(n_208),
.Y(n_705)
);

NOR2xp33_ASAP7_75t_L g706 ( 
.A(n_553),
.B(n_210),
.Y(n_706)
);

NOR2xp33_ASAP7_75t_L g707 ( 
.A(n_674),
.B(n_215),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_L g708 ( 
.A(n_670),
.B(n_508),
.Y(n_708)
);

NOR3xp33_ASAP7_75t_L g709 ( 
.A(n_605),
.B(n_451),
.C(n_219),
.Y(n_709)
);

NOR2xp67_ASAP7_75t_L g710 ( 
.A(n_624),
.B(n_533),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_L g711 ( 
.A(n_639),
.B(n_508),
.Y(n_711)
);

AOI22xp5_ASAP7_75t_L g712 ( 
.A1(n_609),
.A2(n_673),
.B1(n_626),
.B2(n_617),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_545),
.Y(n_713)
);

BUFx6f_ASAP7_75t_SL g714 ( 
.A(n_559),
.Y(n_714)
);

INVx2_ASAP7_75t_L g715 ( 
.A(n_565),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_555),
.Y(n_716)
);

HB1xp67_ASAP7_75t_L g717 ( 
.A(n_573),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_L g718 ( 
.A(n_609),
.B(n_508),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_SL g719 ( 
.A(n_681),
.B(n_188),
.Y(n_719)
);

INVxp67_ASAP7_75t_L g720 ( 
.A(n_651),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_555),
.Y(n_721)
);

AOI22xp33_ASAP7_75t_L g722 ( 
.A1(n_687),
.A2(n_508),
.B1(n_518),
.B2(n_524),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_L g723 ( 
.A(n_565),
.B(n_508),
.Y(n_723)
);

BUFx12f_ASAP7_75t_L g724 ( 
.A(n_653),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_L g725 ( 
.A(n_567),
.B(n_518),
.Y(n_725)
);

OR2x6_ASAP7_75t_L g726 ( 
.A(n_559),
.B(n_244),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_597),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_597),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_L g729 ( 
.A(n_567),
.B(n_518),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_SL g730 ( 
.A(n_680),
.B(n_203),
.Y(n_730)
);

AND2x2_ASAP7_75t_L g731 ( 
.A(n_566),
.B(n_518),
.Y(n_731)
);

INVx2_ASAP7_75t_L g732 ( 
.A(n_568),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_SL g733 ( 
.A(n_680),
.B(n_203),
.Y(n_733)
);

INVx3_ASAP7_75t_L g734 ( 
.A(n_552),
.Y(n_734)
);

BUFx6f_ASAP7_75t_L g735 ( 
.A(n_544),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_SL g736 ( 
.A(n_680),
.B(n_203),
.Y(n_736)
);

BUFx2_ASAP7_75t_L g737 ( 
.A(n_564),
.Y(n_737)
);

BUFx3_ASAP7_75t_L g738 ( 
.A(n_544),
.Y(n_738)
);

INVx2_ASAP7_75t_L g739 ( 
.A(n_568),
.Y(n_739)
);

AOI22xp33_ASAP7_75t_L g740 ( 
.A1(n_574),
.A2(n_518),
.B1(n_524),
.B2(n_343),
.Y(n_740)
);

INVx2_ASAP7_75t_L g741 ( 
.A(n_574),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_575),
.Y(n_742)
);

NOR4xp25_ASAP7_75t_SL g743 ( 
.A(n_621),
.B(n_320),
.C(n_286),
.D(n_283),
.Y(n_743)
);

NOR2xp33_ASAP7_75t_L g744 ( 
.A(n_572),
.B(n_218),
.Y(n_744)
);

INVx2_ASAP7_75t_SL g745 ( 
.A(n_566),
.Y(n_745)
);

INVx5_ASAP7_75t_L g746 ( 
.A(n_680),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_575),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_577),
.Y(n_748)
);

NOR2xp33_ASAP7_75t_L g749 ( 
.A(n_581),
.B(n_220),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_L g750 ( 
.A(n_577),
.B(n_524),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_L g751 ( 
.A(n_582),
.B(n_524),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_582),
.Y(n_752)
);

INVx2_ASAP7_75t_L g753 ( 
.A(n_583),
.Y(n_753)
);

AND2x4_ASAP7_75t_L g754 ( 
.A(n_544),
.B(n_253),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_SL g755 ( 
.A(n_562),
.B(n_203),
.Y(n_755)
);

CKINVDCx5p33_ASAP7_75t_R g756 ( 
.A(n_612),
.Y(n_756)
);

AND2x2_ASAP7_75t_L g757 ( 
.A(n_547),
.B(n_524),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_583),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_SL g759 ( 
.A(n_594),
.B(n_203),
.Y(n_759)
);

BUFx2_ASAP7_75t_L g760 ( 
.A(n_651),
.Y(n_760)
);

NOR3xp33_ASAP7_75t_L g761 ( 
.A(n_623),
.B(n_235),
.C(n_223),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_586),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_586),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_587),
.Y(n_764)
);

OR2x6_ASAP7_75t_L g765 ( 
.A(n_559),
.B(n_253),
.Y(n_765)
);

AND2x4_ASAP7_75t_L g766 ( 
.A(n_551),
.B(n_255),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_587),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_L g768 ( 
.A(n_591),
.B(n_484),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_591),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_593),
.Y(n_770)
);

INVx3_ASAP7_75t_L g771 ( 
.A(n_552),
.Y(n_771)
);

NOR2xp67_ASAP7_75t_L g772 ( 
.A(n_613),
.B(n_387),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_SL g773 ( 
.A(n_599),
.B(n_206),
.Y(n_773)
);

BUFx3_ASAP7_75t_L g774 ( 
.A(n_551),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_593),
.Y(n_775)
);

AND2x2_ASAP7_75t_L g776 ( 
.A(n_547),
.B(n_504),
.Y(n_776)
);

NOR2xp33_ASAP7_75t_L g777 ( 
.A(n_563),
.B(n_241),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_L g778 ( 
.A(n_598),
.B(n_484),
.Y(n_778)
);

INVx2_ASAP7_75t_L g779 ( 
.A(n_598),
.Y(n_779)
);

INVxp67_ASAP7_75t_L g780 ( 
.A(n_691),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_L g781 ( 
.A(n_601),
.B(n_484),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_L g782 ( 
.A(n_601),
.B(n_484),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_L g783 ( 
.A(n_604),
.B(n_484),
.Y(n_783)
);

NAND2xp33_ASAP7_75t_L g784 ( 
.A(n_590),
.B(n_561),
.Y(n_784)
);

INVx2_ASAP7_75t_L g785 ( 
.A(n_604),
.Y(n_785)
);

INVx2_ASAP7_75t_L g786 ( 
.A(n_606),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_L g787 ( 
.A(n_606),
.B(n_484),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_611),
.Y(n_788)
);

INVx1_ASAP7_75t_L g789 ( 
.A(n_611),
.Y(n_789)
);

AOI22xp33_ASAP7_75t_L g790 ( 
.A1(n_628),
.A2(n_298),
.B1(n_255),
.B2(n_257),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_L g791 ( 
.A(n_628),
.B(n_484),
.Y(n_791)
);

INVx4_ASAP7_75t_L g792 ( 
.A(n_551),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_630),
.Y(n_793)
);

INVx3_ASAP7_75t_L g794 ( 
.A(n_552),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_L g795 ( 
.A(n_630),
.B(n_633),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_L g796 ( 
.A(n_633),
.B(n_484),
.Y(n_796)
);

INVx2_ASAP7_75t_L g797 ( 
.A(n_638),
.Y(n_797)
);

AO221x1_ASAP7_75t_L g798 ( 
.A1(n_585),
.A2(n_206),
.B1(n_226),
.B2(n_335),
.C(n_338),
.Y(n_798)
);

NOR2xp33_ASAP7_75t_L g799 ( 
.A(n_569),
.B(n_250),
.Y(n_799)
);

AOI22xp5_ASAP7_75t_L g800 ( 
.A1(n_607),
.A2(n_299),
.B1(n_367),
.B2(n_347),
.Y(n_800)
);

AND2x2_ASAP7_75t_L g801 ( 
.A(n_638),
.B(n_640),
.Y(n_801)
);

NOR2xp33_ASAP7_75t_L g802 ( 
.A(n_644),
.B(n_254),
.Y(n_802)
);

NOR2xp33_ASAP7_75t_L g803 ( 
.A(n_649),
.B(n_260),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_640),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_SL g805 ( 
.A(n_608),
.B(n_206),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_L g806 ( 
.A(n_641),
.B(n_484),
.Y(n_806)
);

INVx3_ASAP7_75t_L g807 ( 
.A(n_552),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_L g808 ( 
.A(n_641),
.B(n_504),
.Y(n_808)
);

INVx2_ASAP7_75t_SL g809 ( 
.A(n_642),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_L g810 ( 
.A(n_642),
.B(n_504),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_L g811 ( 
.A(n_652),
.B(n_504),
.Y(n_811)
);

OR2x2_ASAP7_75t_L g812 ( 
.A(n_584),
.B(n_440),
.Y(n_812)
);

AOI22xp33_ASAP7_75t_L g813 ( 
.A1(n_690),
.A2(n_299),
.B1(n_257),
.B2(n_266),
.Y(n_813)
);

INVx2_ASAP7_75t_L g814 ( 
.A(n_652),
.Y(n_814)
);

AND2x4_ASAP7_75t_SL g815 ( 
.A(n_559),
.B(n_221),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_SL g816 ( 
.A(n_668),
.B(n_629),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_655),
.Y(n_817)
);

AND2x2_ASAP7_75t_L g818 ( 
.A(n_655),
.B(n_512),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_L g819 ( 
.A(n_663),
.B(n_512),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_SL g820 ( 
.A(n_643),
.B(n_206),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_L g821 ( 
.A(n_663),
.B(n_512),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_SL g822 ( 
.A(n_666),
.B(n_206),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_L g823 ( 
.A(n_666),
.B(n_512),
.Y(n_823)
);

AOI22xp33_ASAP7_75t_L g824 ( 
.A1(n_667),
.A2(n_347),
.B1(n_336),
.B2(n_266),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_SL g825 ( 
.A(n_667),
.B(n_226),
.Y(n_825)
);

AND2x2_ASAP7_75t_L g826 ( 
.A(n_672),
.B(n_519),
.Y(n_826)
);

AOI22xp5_ASAP7_75t_L g827 ( 
.A1(n_685),
.A2(n_343),
.B1(n_288),
.B2(n_292),
.Y(n_827)
);

INVx2_ASAP7_75t_L g828 ( 
.A(n_672),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_677),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_SL g830 ( 
.A(n_677),
.B(n_226),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_SL g831 ( 
.A(n_684),
.B(n_226),
.Y(n_831)
);

INVx2_ASAP7_75t_SL g832 ( 
.A(n_684),
.Y(n_832)
);

A2O1A1Ixp33_ASAP7_75t_L g833 ( 
.A1(n_647),
.A2(n_488),
.B(n_502),
.C(n_501),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_L g834 ( 
.A(n_688),
.B(n_519),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_SL g835 ( 
.A(n_688),
.B(n_226),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_L g836 ( 
.A(n_690),
.B(n_519),
.Y(n_836)
);

NOR2xp33_ASAP7_75t_L g837 ( 
.A(n_669),
.B(n_589),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_L g838 ( 
.A(n_635),
.B(n_519),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_L g839 ( 
.A(n_657),
.B(n_521),
.Y(n_839)
);

INVxp67_ASAP7_75t_L g840 ( 
.A(n_589),
.Y(n_840)
);

A2O1A1Ixp33_ASAP7_75t_L g841 ( 
.A1(n_647),
.A2(n_500),
.B(n_502),
.C(n_501),
.Y(n_841)
);

INVx8_ASAP7_75t_L g842 ( 
.A(n_559),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_L g843 ( 
.A(n_671),
.B(n_521),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_SL g844 ( 
.A(n_561),
.B(n_487),
.Y(n_844)
);

NOR2xp33_ASAP7_75t_L g845 ( 
.A(n_600),
.B(n_261),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_557),
.Y(n_846)
);

OAI22xp5_ASAP7_75t_L g847 ( 
.A1(n_619),
.A2(n_298),
.B1(n_367),
.B2(n_336),
.Y(n_847)
);

INVx2_ASAP7_75t_L g848 ( 
.A(n_550),
.Y(n_848)
);

AND2x6_ASAP7_75t_SL g849 ( 
.A(n_614),
.B(n_335),
.Y(n_849)
);

NOR2xp33_ASAP7_75t_L g850 ( 
.A(n_600),
.B(n_263),
.Y(n_850)
);

AOI22xp33_ASAP7_75t_L g851 ( 
.A1(n_590),
.A2(n_689),
.B1(n_665),
.B2(n_661),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_L g852 ( 
.A(n_616),
.B(n_521),
.Y(n_852)
);

INVx1_ASAP7_75t_L g853 ( 
.A(n_557),
.Y(n_853)
);

NOR2xp33_ASAP7_75t_L g854 ( 
.A(n_571),
.B(n_268),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_SL g855 ( 
.A(n_561),
.B(n_487),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_SL g856 ( 
.A(n_579),
.B(n_487),
.Y(n_856)
);

INVx2_ASAP7_75t_L g857 ( 
.A(n_550),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_L g858 ( 
.A(n_616),
.B(n_521),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_L g859 ( 
.A(n_616),
.B(n_522),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_L g860 ( 
.A(n_616),
.B(n_522),
.Y(n_860)
);

INVx1_ASAP7_75t_L g861 ( 
.A(n_560),
.Y(n_861)
);

OAI21xp5_ASAP7_75t_L g862 ( 
.A1(n_703),
.A2(n_570),
.B(n_549),
.Y(n_862)
);

NOR2xp33_ASAP7_75t_L g863 ( 
.A(n_696),
.B(n_660),
.Y(n_863)
);

INVx2_ASAP7_75t_L g864 ( 
.A(n_694),
.Y(n_864)
);

HB1xp67_ASAP7_75t_L g865 ( 
.A(n_717),
.Y(n_865)
);

AOI21xp5_ASAP7_75t_L g866 ( 
.A1(n_695),
.A2(n_570),
.B(n_549),
.Y(n_866)
);

A2O1A1Ixp33_ASAP7_75t_L g867 ( 
.A1(n_837),
.A2(n_310),
.B(n_288),
.C(n_317),
.Y(n_867)
);

AO21x1_ASAP7_75t_L g868 ( 
.A1(n_700),
.A2(n_294),
.B(n_292),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_801),
.Y(n_869)
);

AOI21xp5_ASAP7_75t_L g870 ( 
.A1(n_708),
.A2(n_570),
.B(n_549),
.Y(n_870)
);

AOI21xp5_ASAP7_75t_L g871 ( 
.A1(n_843),
.A2(n_592),
.B(n_543),
.Y(n_871)
);

AOI21xp5_ASAP7_75t_L g872 ( 
.A1(n_816),
.A2(n_592),
.B(n_543),
.Y(n_872)
);

AOI33xp33_ASAP7_75t_L g873 ( 
.A1(n_727),
.A2(n_595),
.A3(n_576),
.B1(n_728),
.B2(n_357),
.B3(n_344),
.Y(n_873)
);

NOR2xp33_ASAP7_75t_L g874 ( 
.A(n_780),
.B(n_622),
.Y(n_874)
);

A2O1A1Ixp33_ASAP7_75t_L g875 ( 
.A1(n_845),
.A2(n_307),
.B(n_327),
.C(n_306),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_L g876 ( 
.A(n_776),
.B(n_625),
.Y(n_876)
);

AOI21xp5_ASAP7_75t_L g877 ( 
.A1(n_816),
.A2(n_592),
.B(n_543),
.Y(n_877)
);

AOI21xp5_ASAP7_75t_L g878 ( 
.A1(n_746),
.A2(n_592),
.B(n_543),
.Y(n_878)
);

AND2x4_ASAP7_75t_L g879 ( 
.A(n_745),
.B(n_440),
.Y(n_879)
);

AOI21xp5_ASAP7_75t_L g880 ( 
.A1(n_746),
.A2(n_618),
.B(n_552),
.Y(n_880)
);

NOR3xp33_ASAP7_75t_L g881 ( 
.A(n_737),
.B(n_622),
.C(n_306),
.Y(n_881)
);

AOI21xp5_ASAP7_75t_L g882 ( 
.A1(n_746),
.A2(n_631),
.B(n_618),
.Y(n_882)
);

INVx3_ASAP7_75t_L g883 ( 
.A(n_735),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_L g884 ( 
.A(n_776),
.B(n_625),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_L g885 ( 
.A(n_757),
.B(n_625),
.Y(n_885)
);

NOR2xp33_ASAP7_75t_L g886 ( 
.A(n_840),
.B(n_229),
.Y(n_886)
);

INVx3_ASAP7_75t_L g887 ( 
.A(n_735),
.Y(n_887)
);

AOI22xp5_ASAP7_75t_L g888 ( 
.A1(n_706),
.A2(n_590),
.B1(n_646),
.B2(n_596),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_SL g889 ( 
.A(n_746),
.B(n_618),
.Y(n_889)
);

NOR2xp33_ASAP7_75t_L g890 ( 
.A(n_720),
.B(n_321),
.Y(n_890)
);

O2A1O1Ixp5_ASAP7_75t_L g891 ( 
.A1(n_755),
.A2(n_646),
.B(n_602),
.C(n_615),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_L g892 ( 
.A(n_757),
.B(n_625),
.Y(n_892)
);

AOI21xp5_ASAP7_75t_L g893 ( 
.A1(n_746),
.A2(n_711),
.B(n_730),
.Y(n_893)
);

BUFx8_ASAP7_75t_L g894 ( 
.A(n_760),
.Y(n_894)
);

OAI22xp5_ASAP7_75t_L g895 ( 
.A1(n_712),
.A2(n_294),
.B1(n_317),
.B2(n_307),
.Y(n_895)
);

NAND2xp5_ASAP7_75t_L g896 ( 
.A(n_731),
.B(n_648),
.Y(n_896)
);

INVx1_ASAP7_75t_L g897 ( 
.A(n_801),
.Y(n_897)
);

AOI21x1_ASAP7_75t_L g898 ( 
.A1(n_730),
.A2(n_596),
.B(n_579),
.Y(n_898)
);

HB1xp67_ASAP7_75t_L g899 ( 
.A(n_701),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_L g900 ( 
.A(n_731),
.B(n_648),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_L g901 ( 
.A(n_802),
.B(n_648),
.Y(n_901)
);

AOI21xp5_ASAP7_75t_L g902 ( 
.A1(n_733),
.A2(n_631),
.B(n_618),
.Y(n_902)
);

INVx1_ASAP7_75t_L g903 ( 
.A(n_694),
.Y(n_903)
);

OR2x2_ASAP7_75t_L g904 ( 
.A(n_812),
.B(n_676),
.Y(n_904)
);

BUFx3_ASAP7_75t_L g905 ( 
.A(n_756),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_SL g906 ( 
.A(n_710),
.B(n_631),
.Y(n_906)
);

CKINVDCx5p33_ASAP7_75t_R g907 ( 
.A(n_756),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_L g908 ( 
.A(n_803),
.B(n_648),
.Y(n_908)
);

NAND3xp33_ASAP7_75t_L g909 ( 
.A(n_850),
.B(n_276),
.C(n_270),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_L g910 ( 
.A(n_701),
.B(n_631),
.Y(n_910)
);

AOI21xp5_ASAP7_75t_L g911 ( 
.A1(n_736),
.A2(n_662),
.B(n_656),
.Y(n_911)
);

AND2x4_ASAP7_75t_L g912 ( 
.A(n_738),
.B(n_441),
.Y(n_912)
);

AOI21xp5_ASAP7_75t_L g913 ( 
.A1(n_736),
.A2(n_662),
.B(n_656),
.Y(n_913)
);

AOI22xp5_ASAP7_75t_L g914 ( 
.A1(n_744),
.A2(n_590),
.B1(n_645),
.B2(n_579),
.Y(n_914)
);

INVxp67_ASAP7_75t_L g915 ( 
.A(n_812),
.Y(n_915)
);

NOR3xp33_ASAP7_75t_L g916 ( 
.A(n_699),
.B(n_854),
.C(n_749),
.Y(n_916)
);

AND2x2_ASAP7_75t_L g917 ( 
.A(n_707),
.B(n_315),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_L g918 ( 
.A(n_809),
.B(n_656),
.Y(n_918)
);

AOI21xp5_ASAP7_75t_L g919 ( 
.A1(n_792),
.A2(n_662),
.B(n_656),
.Y(n_919)
);

NAND2x1p5_ASAP7_75t_L g920 ( 
.A(n_792),
.B(n_656),
.Y(n_920)
);

NOR2xp33_ASAP7_75t_SL g921 ( 
.A(n_772),
.B(n_322),
.Y(n_921)
);

NOR2xp33_ASAP7_75t_L g922 ( 
.A(n_704),
.B(n_705),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_698),
.Y(n_923)
);

OR2x6_ASAP7_75t_L g924 ( 
.A(n_842),
.B(n_308),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_L g925 ( 
.A(n_809),
.B(n_662),
.Y(n_925)
);

OAI22xp33_ASAP7_75t_L g926 ( 
.A1(n_832),
.A2(n_352),
.B1(n_359),
.B2(n_310),
.Y(n_926)
);

INVx3_ASAP7_75t_L g927 ( 
.A(n_735),
.Y(n_927)
);

A2O1A1Ixp33_ASAP7_75t_L g928 ( 
.A1(n_777),
.A2(n_327),
.B(n_308),
.C(n_502),
.Y(n_928)
);

NOR2xp33_ASAP7_75t_L g929 ( 
.A(n_799),
.B(n_281),
.Y(n_929)
);

AND2x2_ASAP7_75t_L g930 ( 
.A(n_697),
.B(n_315),
.Y(n_930)
);

OAI22xp5_ASAP7_75t_L g931 ( 
.A1(n_832),
.A2(n_645),
.B1(n_596),
.B2(n_602),
.Y(n_931)
);

NAND2xp5_ASAP7_75t_L g932 ( 
.A(n_742),
.B(n_747),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_L g933 ( 
.A(n_748),
.B(n_662),
.Y(n_933)
);

INVx2_ASAP7_75t_L g934 ( 
.A(n_698),
.Y(n_934)
);

NAND2xp5_ASAP7_75t_L g935 ( 
.A(n_752),
.B(n_683),
.Y(n_935)
);

NAND2xp5_ASAP7_75t_L g936 ( 
.A(n_758),
.B(n_683),
.Y(n_936)
);

NAND2xp5_ASAP7_75t_L g937 ( 
.A(n_762),
.B(n_683),
.Y(n_937)
);

AOI21xp5_ASAP7_75t_L g938 ( 
.A1(n_792),
.A2(n_839),
.B(n_838),
.Y(n_938)
);

AOI21xp5_ASAP7_75t_L g939 ( 
.A1(n_718),
.A2(n_784),
.B(n_795),
.Y(n_939)
);

HB1xp67_ASAP7_75t_L g940 ( 
.A(n_738),
.Y(n_940)
);

INVxp67_ASAP7_75t_L g941 ( 
.A(n_754),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_L g942 ( 
.A(n_763),
.B(n_764),
.Y(n_942)
);

AOI21xp5_ASAP7_75t_L g943 ( 
.A1(n_784),
.A2(n_686),
.B(n_683),
.Y(n_943)
);

NAND2xp5_ASAP7_75t_L g944 ( 
.A(n_767),
.B(n_683),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_L g945 ( 
.A(n_769),
.B(n_686),
.Y(n_945)
);

INVxp67_ASAP7_75t_SL g946 ( 
.A(n_735),
.Y(n_946)
);

AND2x4_ASAP7_75t_L g947 ( 
.A(n_774),
.B(n_441),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_L g948 ( 
.A(n_770),
.B(n_686),
.Y(n_948)
);

NAND2xp5_ASAP7_75t_L g949 ( 
.A(n_775),
.B(n_686),
.Y(n_949)
);

AOI22xp5_ASAP7_75t_L g950 ( 
.A1(n_754),
.A2(n_590),
.B1(n_615),
.B2(n_646),
.Y(n_950)
);

AOI21xp5_ASAP7_75t_L g951 ( 
.A1(n_719),
.A2(n_686),
.B(n_679),
.Y(n_951)
);

AND2x2_ASAP7_75t_L g952 ( 
.A(n_709),
.B(n_342),
.Y(n_952)
);

AND2x2_ASAP7_75t_L g953 ( 
.A(n_692),
.B(n_342),
.Y(n_953)
);

AND2x2_ASAP7_75t_L g954 ( 
.A(n_692),
.B(n_342),
.Y(n_954)
);

BUFx3_ASAP7_75t_L g955 ( 
.A(n_702),
.Y(n_955)
);

A2O1A1Ixp33_ASAP7_75t_L g956 ( 
.A1(n_800),
.A2(n_827),
.B(n_851),
.C(n_789),
.Y(n_956)
);

INVx2_ASAP7_75t_L g957 ( 
.A(n_715),
.Y(n_957)
);

BUFx4f_ASAP7_75t_L g958 ( 
.A(n_724),
.Y(n_958)
);

INVx3_ASAP7_75t_L g959 ( 
.A(n_774),
.Y(n_959)
);

BUFx4f_ASAP7_75t_SL g960 ( 
.A(n_724),
.Y(n_960)
);

INVxp67_ASAP7_75t_L g961 ( 
.A(n_754),
.Y(n_961)
);

INVx1_ASAP7_75t_L g962 ( 
.A(n_715),
.Y(n_962)
);

OR2x2_ASAP7_75t_L g963 ( 
.A(n_766),
.B(n_676),
.Y(n_963)
);

INVxp67_ASAP7_75t_L g964 ( 
.A(n_766),
.Y(n_964)
);

NAND2xp5_ASAP7_75t_L g965 ( 
.A(n_788),
.B(n_602),
.Y(n_965)
);

AOI21xp33_ASAP7_75t_L g966 ( 
.A1(n_726),
.A2(n_326),
.B(n_290),
.Y(n_966)
);

NAND2xp5_ASAP7_75t_L g967 ( 
.A(n_793),
.B(n_615),
.Y(n_967)
);

INVxp67_ASAP7_75t_L g968 ( 
.A(n_766),
.Y(n_968)
);

OR2x6_ASAP7_75t_L g969 ( 
.A(n_842),
.B(n_338),
.Y(n_969)
);

BUFx12f_ASAP7_75t_L g970 ( 
.A(n_702),
.Y(n_970)
);

AOI21xp5_ASAP7_75t_L g971 ( 
.A1(n_719),
.A2(n_679),
.B(n_580),
.Y(n_971)
);

INVx1_ASAP7_75t_L g972 ( 
.A(n_732),
.Y(n_972)
);

AOI21x1_ASAP7_75t_L g973 ( 
.A1(n_755),
.A2(n_645),
.B(n_675),
.Y(n_973)
);

INVx1_ASAP7_75t_L g974 ( 
.A(n_732),
.Y(n_974)
);

NAND2xp5_ASAP7_75t_L g975 ( 
.A(n_804),
.B(n_627),
.Y(n_975)
);

A2O1A1Ixp33_ASAP7_75t_L g976 ( 
.A1(n_817),
.A2(n_500),
.B(n_678),
.C(n_675),
.Y(n_976)
);

OAI21xp5_ASAP7_75t_L g977 ( 
.A1(n_723),
.A2(n_682),
.B(n_627),
.Y(n_977)
);

INVx2_ASAP7_75t_L g978 ( 
.A(n_739),
.Y(n_978)
);

AOI21xp5_ASAP7_75t_L g979 ( 
.A1(n_759),
.A2(n_679),
.B(n_580),
.Y(n_979)
);

AOI21xp5_ASAP7_75t_L g980 ( 
.A1(n_759),
.A2(n_679),
.B(n_580),
.Y(n_980)
);

AOI21xp5_ASAP7_75t_L g981 ( 
.A1(n_773),
.A2(n_805),
.B(n_852),
.Y(n_981)
);

HB1xp67_ASAP7_75t_L g982 ( 
.A(n_829),
.Y(n_982)
);

INVx1_ASAP7_75t_SL g983 ( 
.A(n_849),
.Y(n_983)
);

AOI21xp5_ASAP7_75t_L g984 ( 
.A1(n_773),
.A2(n_679),
.B(n_678),
.Y(n_984)
);

NOR2xp33_ASAP7_75t_L g985 ( 
.A(n_693),
.B(n_282),
.Y(n_985)
);

AND2x2_ASAP7_75t_L g986 ( 
.A(n_761),
.B(n_342),
.Y(n_986)
);

NAND2xp5_ASAP7_75t_L g987 ( 
.A(n_739),
.B(n_632),
.Y(n_987)
);

OAI22xp5_ASAP7_75t_L g988 ( 
.A1(n_741),
.A2(n_675),
.B1(n_678),
.B2(n_682),
.Y(n_988)
);

NAND2xp5_ASAP7_75t_SL g989 ( 
.A(n_741),
.B(n_632),
.Y(n_989)
);

OAI321xp33_ASAP7_75t_L g990 ( 
.A1(n_847),
.A2(n_366),
.A3(n_351),
.B1(n_357),
.B2(n_364),
.C(n_452),
.Y(n_990)
);

OAI22xp5_ASAP7_75t_L g991 ( 
.A1(n_753),
.A2(n_650),
.B1(n_664),
.B2(n_659),
.Y(n_991)
);

NAND2xp5_ASAP7_75t_SL g992 ( 
.A(n_815),
.B(n_779),
.Y(n_992)
);

BUFx8_ASAP7_75t_L g993 ( 
.A(n_714),
.Y(n_993)
);

A2O1A1Ixp33_ASAP7_75t_L g994 ( 
.A1(n_713),
.A2(n_658),
.B(n_637),
.C(n_634),
.Y(n_994)
);

INVxp67_ASAP7_75t_L g995 ( 
.A(n_716),
.Y(n_995)
);

AOI21xp5_ASAP7_75t_L g996 ( 
.A1(n_858),
.A2(n_679),
.B(n_475),
.Y(n_996)
);

NAND2xp5_ASAP7_75t_L g997 ( 
.A(n_779),
.B(n_785),
.Y(n_997)
);

BUFx2_ASAP7_75t_SL g998 ( 
.A(n_714),
.Y(n_998)
);

AOI21xp5_ASAP7_75t_L g999 ( 
.A1(n_859),
.A2(n_475),
.B(n_471),
.Y(n_999)
);

AOI21xp5_ASAP7_75t_L g1000 ( 
.A1(n_860),
.A2(n_475),
.B(n_471),
.Y(n_1000)
);

INVx2_ASAP7_75t_SL g1001 ( 
.A(n_702),
.Y(n_1001)
);

OAI22xp5_ASAP7_75t_L g1002 ( 
.A1(n_785),
.A2(n_786),
.B1(n_814),
.B2(n_797),
.Y(n_1002)
);

AOI21xp5_ASAP7_75t_L g1003 ( 
.A1(n_820),
.A2(n_475),
.B(n_637),
.Y(n_1003)
);

NAND2xp5_ASAP7_75t_L g1004 ( 
.A(n_786),
.B(n_634),
.Y(n_1004)
);

AOI21xp5_ASAP7_75t_L g1005 ( 
.A1(n_820),
.A2(n_475),
.B(n_658),
.Y(n_1005)
);

INVx2_ASAP7_75t_L g1006 ( 
.A(n_797),
.Y(n_1006)
);

NAND2xp5_ASAP7_75t_L g1007 ( 
.A(n_814),
.B(n_542),
.Y(n_1007)
);

BUFx6f_ASAP7_75t_L g1008 ( 
.A(n_842),
.Y(n_1008)
);

INVx1_ASAP7_75t_L g1009 ( 
.A(n_828),
.Y(n_1009)
);

NAND2x1_ASAP7_75t_L g1010 ( 
.A(n_734),
.B(n_590),
.Y(n_1010)
);

INVx2_ASAP7_75t_SL g1011 ( 
.A(n_815),
.Y(n_1011)
);

AOI21xp5_ASAP7_75t_L g1012 ( 
.A1(n_734),
.A2(n_542),
.B(n_556),
.Y(n_1012)
);

NAND2xp5_ASAP7_75t_SL g1013 ( 
.A(n_842),
.B(n_221),
.Y(n_1013)
);

INVx2_ASAP7_75t_L g1014 ( 
.A(n_848),
.Y(n_1014)
);

NAND2xp5_ASAP7_75t_L g1015 ( 
.A(n_721),
.B(n_554),
.Y(n_1015)
);

NAND2xp5_ASAP7_75t_L g1016 ( 
.A(n_818),
.B(n_826),
.Y(n_1016)
);

INVx2_ASAP7_75t_L g1017 ( 
.A(n_848),
.Y(n_1017)
);

BUFx12f_ASAP7_75t_L g1018 ( 
.A(n_726),
.Y(n_1018)
);

AND2x2_ASAP7_75t_L g1019 ( 
.A(n_743),
.B(n_450),
.Y(n_1019)
);

O2A1O1Ixp33_ASAP7_75t_L g1020 ( 
.A1(n_822),
.A2(n_531),
.B(n_364),
.C(n_554),
.Y(n_1020)
);

INVx2_ASAP7_75t_L g1021 ( 
.A(n_857),
.Y(n_1021)
);

OAI21xp5_ASAP7_75t_L g1022 ( 
.A1(n_725),
.A2(n_590),
.B(n_478),
.Y(n_1022)
);

BUFx6f_ASAP7_75t_L g1023 ( 
.A(n_771),
.Y(n_1023)
);

NAND2xp5_ASAP7_75t_L g1024 ( 
.A(n_818),
.B(n_826),
.Y(n_1024)
);

BUFx6f_ASAP7_75t_L g1025 ( 
.A(n_771),
.Y(n_1025)
);

AOI21xp5_ASAP7_75t_L g1026 ( 
.A1(n_771),
.A2(n_479),
.B(n_476),
.Y(n_1026)
);

HB1xp67_ASAP7_75t_L g1027 ( 
.A(n_726),
.Y(n_1027)
);

AOI21xp5_ASAP7_75t_L g1028 ( 
.A1(n_794),
.A2(n_479),
.B(n_476),
.Y(n_1028)
);

BUFx6f_ASAP7_75t_L g1029 ( 
.A(n_794),
.Y(n_1029)
);

NAND2xp5_ASAP7_75t_SL g1030 ( 
.A(n_722),
.B(n_487),
.Y(n_1030)
);

OAI21xp5_ASAP7_75t_L g1031 ( 
.A1(n_729),
.A2(n_472),
.B(n_478),
.Y(n_1031)
);

NOR2xp33_ASAP7_75t_L g1032 ( 
.A(n_750),
.B(n_293),
.Y(n_1032)
);

O2A1O1Ixp33_ASAP7_75t_SL g1033 ( 
.A1(n_833),
.A2(n_470),
.B(n_464),
.C(n_465),
.Y(n_1033)
);

AOI21xp5_ASAP7_75t_L g1034 ( 
.A1(n_794),
.A2(n_479),
.B(n_476),
.Y(n_1034)
);

OAI22xp5_ASAP7_75t_L g1035 ( 
.A1(n_740),
.A2(n_349),
.B1(n_350),
.B2(n_301),
.Y(n_1035)
);

INVx4_ASAP7_75t_L g1036 ( 
.A(n_714),
.Y(n_1036)
);

OAI22xp5_ASAP7_75t_L g1037 ( 
.A1(n_726),
.A2(n_356),
.B1(n_360),
.B2(n_302),
.Y(n_1037)
);

AOI21xp5_ASAP7_75t_L g1038 ( 
.A1(n_807),
.A2(n_751),
.B(n_836),
.Y(n_1038)
);

NAND2xp5_ASAP7_75t_L g1039 ( 
.A(n_857),
.B(n_522),
.Y(n_1039)
);

NAND2xp5_ASAP7_75t_SL g1040 ( 
.A(n_790),
.B(n_230),
.Y(n_1040)
);

OAI22xp33_ASAP7_75t_L g1041 ( 
.A1(n_765),
.A2(n_810),
.B1(n_808),
.B2(n_811),
.Y(n_1041)
);

INVxp67_ASAP7_75t_L g1042 ( 
.A(n_765),
.Y(n_1042)
);

INVx1_ASAP7_75t_L g1043 ( 
.A(n_846),
.Y(n_1043)
);

NAND2xp5_ASAP7_75t_L g1044 ( 
.A(n_853),
.B(n_522),
.Y(n_1044)
);

AOI21x1_ASAP7_75t_L g1045 ( 
.A1(n_844),
.A2(n_472),
.B(n_478),
.Y(n_1045)
);

AND2x2_ASAP7_75t_L g1046 ( 
.A(n_765),
.B(n_450),
.Y(n_1046)
);

NAND2xp5_ASAP7_75t_L g1047 ( 
.A(n_861),
.B(n_529),
.Y(n_1047)
);

NAND2xp5_ASAP7_75t_L g1048 ( 
.A(n_899),
.B(n_819),
.Y(n_1048)
);

INVx3_ASAP7_75t_L g1049 ( 
.A(n_883),
.Y(n_1049)
);

NAND2xp5_ASAP7_75t_L g1050 ( 
.A(n_899),
.B(n_922),
.Y(n_1050)
);

AOI21xp5_ASAP7_75t_L g1051 ( 
.A1(n_1016),
.A2(n_833),
.B(n_841),
.Y(n_1051)
);

INVx4_ASAP7_75t_L g1052 ( 
.A(n_1008),
.Y(n_1052)
);

NAND2xp5_ASAP7_75t_L g1053 ( 
.A(n_922),
.B(n_821),
.Y(n_1053)
);

INVx1_ASAP7_75t_L g1054 ( 
.A(n_982),
.Y(n_1054)
);

INVx6_ASAP7_75t_L g1055 ( 
.A(n_894),
.Y(n_1055)
);

INVx1_ASAP7_75t_L g1056 ( 
.A(n_982),
.Y(n_1056)
);

NAND2xp5_ASAP7_75t_R g1057 ( 
.A(n_1001),
.B(n_765),
.Y(n_1057)
);

NAND2xp5_ASAP7_75t_L g1058 ( 
.A(n_1024),
.B(n_823),
.Y(n_1058)
);

AO21x2_ASAP7_75t_L g1059 ( 
.A1(n_1041),
.A2(n_798),
.B(n_841),
.Y(n_1059)
);

AOI22xp33_ASAP7_75t_L g1060 ( 
.A1(n_916),
.A2(n_929),
.B1(n_1019),
.B2(n_895),
.Y(n_1060)
);

AOI22xp33_ASAP7_75t_L g1061 ( 
.A1(n_916),
.A2(n_813),
.B1(n_824),
.B2(n_230),
.Y(n_1061)
);

INVx1_ASAP7_75t_L g1062 ( 
.A(n_903),
.Y(n_1062)
);

INVx1_ASAP7_75t_L g1063 ( 
.A(n_923),
.Y(n_1063)
);

NOR2xp33_ASAP7_75t_L g1064 ( 
.A(n_886),
.B(n_834),
.Y(n_1064)
);

NOR2xp33_ASAP7_75t_R g1065 ( 
.A(n_907),
.B(n_768),
.Y(n_1065)
);

A2O1A1Ixp33_ASAP7_75t_L g1066 ( 
.A1(n_956),
.A2(n_806),
.B(n_781),
.C(n_782),
.Y(n_1066)
);

OAI21x1_ASAP7_75t_L g1067 ( 
.A1(n_1045),
.A2(n_783),
.B(n_791),
.Y(n_1067)
);

BUFx12f_ASAP7_75t_L g1068 ( 
.A(n_894),
.Y(n_1068)
);

NAND3xp33_ASAP7_75t_L g1069 ( 
.A(n_890),
.B(n_303),
.C(n_361),
.Y(n_1069)
);

AOI21xp5_ASAP7_75t_L g1070 ( 
.A1(n_938),
.A2(n_908),
.B(n_901),
.Y(n_1070)
);

NOR2xp33_ASAP7_75t_L g1071 ( 
.A(n_886),
.B(n_778),
.Y(n_1071)
);

AOI21xp5_ASAP7_75t_L g1072 ( 
.A1(n_866),
.A2(n_796),
.B(n_787),
.Y(n_1072)
);

NOR2xp33_ASAP7_75t_L g1073 ( 
.A(n_915),
.B(n_844),
.Y(n_1073)
);

NOR2xp33_ASAP7_75t_R g1074 ( 
.A(n_960),
.B(n_312),
.Y(n_1074)
);

HB1xp67_ASAP7_75t_L g1075 ( 
.A(n_865),
.Y(n_1075)
);

BUFx8_ASAP7_75t_L g1076 ( 
.A(n_970),
.Y(n_1076)
);

BUFx6f_ASAP7_75t_L g1077 ( 
.A(n_1008),
.Y(n_1077)
);

NOR2xp33_ASAP7_75t_L g1078 ( 
.A(n_915),
.B(n_890),
.Y(n_1078)
);

INVx1_ASAP7_75t_L g1079 ( 
.A(n_962),
.Y(n_1079)
);

OAI221xp5_ASAP7_75t_L g1080 ( 
.A1(n_869),
.A2(n_355),
.B1(n_346),
.B2(n_345),
.C(n_341),
.Y(n_1080)
);

NOR2xp33_ASAP7_75t_L g1081 ( 
.A(n_865),
.B(n_855),
.Y(n_1081)
);

OAI21xp33_ASAP7_75t_L g1082 ( 
.A1(n_917),
.A2(n_921),
.B(n_985),
.Y(n_1082)
);

AOI22xp33_ASAP7_75t_L g1083 ( 
.A1(n_963),
.A2(n_1046),
.B1(n_941),
.B2(n_964),
.Y(n_1083)
);

NOR3xp33_ASAP7_75t_SL g1084 ( 
.A(n_926),
.B(n_334),
.C(n_330),
.Y(n_1084)
);

NAND2xp5_ASAP7_75t_SL g1085 ( 
.A(n_904),
.B(n_230),
.Y(n_1085)
);

NAND2xp5_ASAP7_75t_SL g1086 ( 
.A(n_930),
.B(n_230),
.Y(n_1086)
);

NAND2xp5_ASAP7_75t_L g1087 ( 
.A(n_897),
.B(n_855),
.Y(n_1087)
);

INVx1_ASAP7_75t_L g1088 ( 
.A(n_972),
.Y(n_1088)
);

NAND2xp5_ASAP7_75t_L g1089 ( 
.A(n_910),
.B(n_856),
.Y(n_1089)
);

AOI21xp5_ASAP7_75t_L g1090 ( 
.A1(n_862),
.A2(n_856),
.B(n_835),
.Y(n_1090)
);

NOR2xp33_ASAP7_75t_L g1091 ( 
.A(n_874),
.B(n_822),
.Y(n_1091)
);

HB1xp67_ASAP7_75t_L g1092 ( 
.A(n_940),
.Y(n_1092)
);

OAI22xp5_ASAP7_75t_L g1093 ( 
.A1(n_941),
.A2(n_835),
.B1(n_831),
.B2(n_830),
.Y(n_1093)
);

BUFx2_ASAP7_75t_L g1094 ( 
.A(n_905),
.Y(n_1094)
);

O2A1O1Ixp33_ASAP7_75t_L g1095 ( 
.A1(n_875),
.A2(n_831),
.B(n_830),
.C(n_825),
.Y(n_1095)
);

AOI21xp5_ASAP7_75t_L g1096 ( 
.A1(n_876),
.A2(n_825),
.B(n_479),
.Y(n_1096)
);

AOI21xp5_ASAP7_75t_L g1097 ( 
.A1(n_884),
.A2(n_531),
.B(n_478),
.Y(n_1097)
);

AOI21xp5_ASAP7_75t_L g1098 ( 
.A1(n_939),
.A2(n_465),
.B(n_464),
.Y(n_1098)
);

OAI21xp5_ASAP7_75t_L g1099 ( 
.A1(n_896),
.A2(n_465),
.B(n_464),
.Y(n_1099)
);

AOI21xp5_ASAP7_75t_L g1100 ( 
.A1(n_893),
.A2(n_871),
.B(n_919),
.Y(n_1100)
);

BUFx3_ASAP7_75t_L g1101 ( 
.A(n_958),
.Y(n_1101)
);

NAND2xp5_ASAP7_75t_L g1102 ( 
.A(n_932),
.B(n_942),
.Y(n_1102)
);

INVx1_ASAP7_75t_L g1103 ( 
.A(n_974),
.Y(n_1103)
);

O2A1O1Ixp33_ASAP7_75t_L g1104 ( 
.A1(n_926),
.A2(n_534),
.B(n_532),
.C(n_529),
.Y(n_1104)
);

NAND3xp33_ASAP7_75t_SL g1105 ( 
.A(n_881),
.B(n_459),
.C(n_452),
.Y(n_1105)
);

AOI21xp5_ASAP7_75t_L g1106 ( 
.A1(n_971),
.A2(n_470),
.B(n_532),
.Y(n_1106)
);

INVx1_ASAP7_75t_SL g1107 ( 
.A(n_953),
.Y(n_1107)
);

BUFx6f_ASAP7_75t_L g1108 ( 
.A(n_1008),
.Y(n_1108)
);

OR2x6_ASAP7_75t_SL g1109 ( 
.A(n_909),
.B(n_453),
.Y(n_1109)
);

AOI22xp33_ASAP7_75t_L g1110 ( 
.A1(n_961),
.A2(n_964),
.B1(n_968),
.B2(n_952),
.Y(n_1110)
);

AOI21xp5_ASAP7_75t_L g1111 ( 
.A1(n_885),
.A2(n_470),
.B(n_532),
.Y(n_1111)
);

AO21x2_ASAP7_75t_L g1112 ( 
.A1(n_1041),
.A2(n_481),
.B(n_477),
.Y(n_1112)
);

INVx2_ASAP7_75t_L g1113 ( 
.A(n_864),
.Y(n_1113)
);

INVx3_ASAP7_75t_L g1114 ( 
.A(n_883),
.Y(n_1114)
);

NOR2xp33_ASAP7_75t_L g1115 ( 
.A(n_874),
.B(n_365),
.Y(n_1115)
);

INVx1_ASAP7_75t_SL g1116 ( 
.A(n_954),
.Y(n_1116)
);

BUFx6f_ASAP7_75t_L g1117 ( 
.A(n_1008),
.Y(n_1117)
);

NOR2xp33_ASAP7_75t_R g1118 ( 
.A(n_960),
.B(n_77),
.Y(n_1118)
);

OAI22xp5_ASAP7_75t_L g1119 ( 
.A1(n_961),
.A2(n_534),
.B1(n_532),
.B2(n_529),
.Y(n_1119)
);

OAI22xp5_ASAP7_75t_L g1120 ( 
.A1(n_968),
.A2(n_534),
.B1(n_529),
.B2(n_477),
.Y(n_1120)
);

OAI22xp5_ASAP7_75t_L g1121 ( 
.A1(n_995),
.A2(n_534),
.B1(n_481),
.B2(n_487),
.Y(n_1121)
);

AO32x2_ASAP7_75t_L g1122 ( 
.A1(n_1002),
.A2(n_365),
.A3(n_11),
.B1(n_12),
.B2(n_14),
.Y(n_1122)
);

HB1xp67_ASAP7_75t_L g1123 ( 
.A(n_940),
.Y(n_1123)
);

A2O1A1Ixp33_ASAP7_75t_L g1124 ( 
.A1(n_1032),
.A2(n_459),
.B(n_458),
.C(n_454),
.Y(n_1124)
);

BUFx3_ASAP7_75t_L g1125 ( 
.A(n_958),
.Y(n_1125)
);

NOR2xp33_ASAP7_75t_L g1126 ( 
.A(n_863),
.B(n_995),
.Y(n_1126)
);

BUFx6f_ASAP7_75t_L g1127 ( 
.A(n_1023),
.Y(n_1127)
);

AOI21xp5_ASAP7_75t_L g1128 ( 
.A1(n_892),
.A2(n_481),
.B(n_487),
.Y(n_1128)
);

NAND2xp5_ASAP7_75t_L g1129 ( 
.A(n_900),
.B(n_487),
.Y(n_1129)
);

AOI21xp5_ASAP7_75t_L g1130 ( 
.A1(n_870),
.A2(n_458),
.B(n_454),
.Y(n_1130)
);

BUFx12f_ASAP7_75t_L g1131 ( 
.A(n_993),
.Y(n_1131)
);

BUFx2_ASAP7_75t_L g1132 ( 
.A(n_969),
.Y(n_1132)
);

INVx4_ASAP7_75t_L g1133 ( 
.A(n_959),
.Y(n_1133)
);

INVx1_ASAP7_75t_L g1134 ( 
.A(n_1009),
.Y(n_1134)
);

INVxp67_ASAP7_75t_SL g1135 ( 
.A(n_946),
.Y(n_1135)
);

AOI21xp5_ASAP7_75t_L g1136 ( 
.A1(n_872),
.A2(n_123),
.B(n_180),
.Y(n_1136)
);

CKINVDCx14_ASAP7_75t_R g1137 ( 
.A(n_955),
.Y(n_1137)
);

AOI22xp33_ASAP7_75t_SL g1138 ( 
.A1(n_863),
.A2(n_986),
.B1(n_993),
.B2(n_1018),
.Y(n_1138)
);

INVx1_ASAP7_75t_L g1139 ( 
.A(n_934),
.Y(n_1139)
);

BUFx2_ASAP7_75t_L g1140 ( 
.A(n_969),
.Y(n_1140)
);

OAI21xp5_ASAP7_75t_L g1141 ( 
.A1(n_1038),
.A2(n_365),
.B(n_174),
.Y(n_1141)
);

AOI21xp5_ASAP7_75t_L g1142 ( 
.A1(n_877),
.A2(n_118),
.B(n_170),
.Y(n_1142)
);

NOR2xp33_ASAP7_75t_L g1143 ( 
.A(n_985),
.B(n_365),
.Y(n_1143)
);

OAI21x1_ASAP7_75t_L g1144 ( 
.A1(n_973),
.A2(n_898),
.B(n_878),
.Y(n_1144)
);

AOI21xp5_ASAP7_75t_L g1145 ( 
.A1(n_946),
.A2(n_168),
.B(n_147),
.Y(n_1145)
);

NAND2xp5_ASAP7_75t_L g1146 ( 
.A(n_997),
.B(n_139),
.Y(n_1146)
);

INVx1_ASAP7_75t_SL g1147 ( 
.A(n_983),
.Y(n_1147)
);

OAI22x1_ASAP7_75t_L g1148 ( 
.A1(n_1042),
.A2(n_10),
.B1(n_12),
.B2(n_14),
.Y(n_1148)
);

AOI21xp5_ASAP7_75t_L g1149 ( 
.A1(n_918),
.A2(n_135),
.B(n_134),
.Y(n_1149)
);

NOR2xp33_ASAP7_75t_L g1150 ( 
.A(n_966),
.B(n_17),
.Y(n_1150)
);

NAND2xp5_ASAP7_75t_L g1151 ( 
.A(n_957),
.B(n_127),
.Y(n_1151)
);

NAND2xp5_ASAP7_75t_L g1152 ( 
.A(n_978),
.B(n_121),
.Y(n_1152)
);

INVx1_ASAP7_75t_L g1153 ( 
.A(n_1006),
.Y(n_1153)
);

A2O1A1Ixp33_ASAP7_75t_L g1154 ( 
.A1(n_1032),
.A2(n_20),
.B(n_21),
.C(n_22),
.Y(n_1154)
);

NAND2xp5_ASAP7_75t_L g1155 ( 
.A(n_879),
.B(n_116),
.Y(n_1155)
);

OAI21xp33_ASAP7_75t_SL g1156 ( 
.A1(n_992),
.A2(n_27),
.B(n_28),
.Y(n_1156)
);

AOI21xp5_ASAP7_75t_L g1157 ( 
.A1(n_925),
.A2(n_115),
.B(n_114),
.Y(n_1157)
);

INVx1_ASAP7_75t_L g1158 ( 
.A(n_1014),
.Y(n_1158)
);

INVx2_ASAP7_75t_L g1159 ( 
.A(n_1017),
.Y(n_1159)
);

NAND2xp5_ASAP7_75t_SL g1160 ( 
.A(n_879),
.B(n_113),
.Y(n_1160)
);

CKINVDCx14_ASAP7_75t_R g1161 ( 
.A(n_1036),
.Y(n_1161)
);

NAND2xp5_ASAP7_75t_L g1162 ( 
.A(n_1021),
.B(n_93),
.Y(n_1162)
);

AOI21xp5_ASAP7_75t_L g1163 ( 
.A1(n_943),
.A2(n_85),
.B(n_80),
.Y(n_1163)
);

NAND3xp33_ASAP7_75t_L g1164 ( 
.A(n_881),
.B(n_27),
.C(n_30),
.Y(n_1164)
);

NAND2xp5_ASAP7_75t_L g1165 ( 
.A(n_959),
.B(n_78),
.Y(n_1165)
);

OR2x6_ASAP7_75t_L g1166 ( 
.A(n_998),
.B(n_30),
.Y(n_1166)
);

OAI22xp5_ASAP7_75t_SL g1167 ( 
.A1(n_1042),
.A2(n_33),
.B1(n_36),
.B2(n_37),
.Y(n_1167)
);

INVx1_ASAP7_75t_L g1168 ( 
.A(n_1043),
.Y(n_1168)
);

NAND2x1_ASAP7_75t_L g1169 ( 
.A(n_887),
.B(n_41),
.Y(n_1169)
);

BUFx6f_ASAP7_75t_L g1170 ( 
.A(n_1023),
.Y(n_1170)
);

OAI22xp5_ASAP7_75t_L g1171 ( 
.A1(n_1027),
.A2(n_41),
.B1(n_43),
.B2(n_44),
.Y(n_1171)
);

AOI22xp33_ASAP7_75t_L g1172 ( 
.A1(n_912),
.A2(n_43),
.B1(n_45),
.B2(n_46),
.Y(n_1172)
);

INVx2_ASAP7_75t_L g1173 ( 
.A(n_912),
.Y(n_1173)
);

A2O1A1Ixp33_ASAP7_75t_L g1174 ( 
.A1(n_873),
.A2(n_981),
.B(n_947),
.C(n_928),
.Y(n_1174)
);

AND2x4_ASAP7_75t_L g1175 ( 
.A(n_1036),
.B(n_46),
.Y(n_1175)
);

AOI21xp5_ASAP7_75t_L g1176 ( 
.A1(n_979),
.A2(n_72),
.B(n_54),
.Y(n_1176)
);

NOR2xp33_ASAP7_75t_L g1177 ( 
.A(n_947),
.B(n_53),
.Y(n_1177)
);

INVx1_ASAP7_75t_L g1178 ( 
.A(n_975),
.Y(n_1178)
);

NAND2xp5_ASAP7_75t_SL g1179 ( 
.A(n_1011),
.B(n_59),
.Y(n_1179)
);

NAND2xp5_ASAP7_75t_SL g1180 ( 
.A(n_1027),
.B(n_60),
.Y(n_1180)
);

INVx1_ASAP7_75t_SL g1181 ( 
.A(n_969),
.Y(n_1181)
);

INVx6_ASAP7_75t_L g1182 ( 
.A(n_1023),
.Y(n_1182)
);

A2O1A1Ixp33_ASAP7_75t_L g1183 ( 
.A1(n_888),
.A2(n_60),
.B(n_61),
.C(n_62),
.Y(n_1183)
);

AND2x4_ASAP7_75t_L g1184 ( 
.A(n_924),
.B(n_66),
.Y(n_1184)
);

INVx2_ASAP7_75t_L g1185 ( 
.A(n_1007),
.Y(n_1185)
);

BUFx8_ASAP7_75t_SL g1186 ( 
.A(n_924),
.Y(n_1186)
);

INVx1_ASAP7_75t_L g1187 ( 
.A(n_1044),
.Y(n_1187)
);

NAND2xp5_ASAP7_75t_SL g1188 ( 
.A(n_1023),
.B(n_66),
.Y(n_1188)
);

A2O1A1Ixp33_ASAP7_75t_L g1189 ( 
.A1(n_914),
.A2(n_867),
.B(n_891),
.C(n_950),
.Y(n_1189)
);

BUFx8_ASAP7_75t_L g1190 ( 
.A(n_1025),
.Y(n_1190)
);

INVx1_ASAP7_75t_L g1191 ( 
.A(n_1047),
.Y(n_1191)
);

O2A1O1Ixp33_ASAP7_75t_L g1192 ( 
.A1(n_1013),
.A2(n_67),
.B(n_68),
.C(n_69),
.Y(n_1192)
);

OAI22xp5_ASAP7_75t_L g1193 ( 
.A1(n_933),
.A2(n_67),
.B1(n_68),
.B2(n_70),
.Y(n_1193)
);

BUFx6f_ASAP7_75t_L g1194 ( 
.A(n_1025),
.Y(n_1194)
);

NAND2xp5_ASAP7_75t_SL g1195 ( 
.A(n_1025),
.B(n_71),
.Y(n_1195)
);

AOI21xp5_ASAP7_75t_L g1196 ( 
.A1(n_980),
.A2(n_889),
.B(n_920),
.Y(n_1196)
);

BUFx3_ASAP7_75t_L g1197 ( 
.A(n_924),
.Y(n_1197)
);

NAND2xp5_ASAP7_75t_L g1198 ( 
.A(n_965),
.B(n_967),
.Y(n_1198)
);

INVx4_ASAP7_75t_L g1199 ( 
.A(n_1025),
.Y(n_1199)
);

BUFx2_ASAP7_75t_L g1200 ( 
.A(n_887),
.Y(n_1200)
);

NOR2xp33_ASAP7_75t_R g1201 ( 
.A(n_927),
.B(n_1029),
.Y(n_1201)
);

NAND2xp5_ASAP7_75t_SL g1202 ( 
.A(n_1029),
.B(n_927),
.Y(n_1202)
);

NAND2xp5_ASAP7_75t_SL g1203 ( 
.A(n_1029),
.B(n_1037),
.Y(n_1203)
);

NAND2xp5_ASAP7_75t_SL g1204 ( 
.A(n_1029),
.B(n_920),
.Y(n_1204)
);

INVx4_ASAP7_75t_L g1205 ( 
.A(n_1010),
.Y(n_1205)
);

NAND2xp5_ASAP7_75t_L g1206 ( 
.A(n_987),
.B(n_1004),
.Y(n_1206)
);

BUFx8_ASAP7_75t_L g1207 ( 
.A(n_990),
.Y(n_1207)
);

AND2x2_ASAP7_75t_L g1208 ( 
.A(n_1035),
.B(n_1040),
.Y(n_1208)
);

NAND2xp5_ASAP7_75t_SL g1209 ( 
.A(n_868),
.B(n_906),
.Y(n_1209)
);

NAND2xp5_ASAP7_75t_L g1210 ( 
.A(n_1015),
.B(n_944),
.Y(n_1210)
);

O2A1O1Ixp33_ASAP7_75t_L g1211 ( 
.A1(n_1033),
.A2(n_994),
.B(n_976),
.C(n_931),
.Y(n_1211)
);

AOI21xp5_ASAP7_75t_L g1212 ( 
.A1(n_1030),
.A2(n_1031),
.B(n_1022),
.Y(n_1212)
);

OAI22xp5_ASAP7_75t_L g1213 ( 
.A1(n_1102),
.A2(n_948),
.B1(n_936),
.B2(n_937),
.Y(n_1213)
);

AO31x2_ASAP7_75t_L g1214 ( 
.A1(n_1070),
.A2(n_1189),
.A3(n_1100),
.B(n_1174),
.Y(n_1214)
);

AOI221x1_ASAP7_75t_L g1215 ( 
.A1(n_1143),
.A2(n_988),
.B1(n_999),
.B2(n_1000),
.C(n_991),
.Y(n_1215)
);

OAI21xp5_ASAP7_75t_L g1216 ( 
.A1(n_1051),
.A2(n_891),
.B(n_977),
.Y(n_1216)
);

AOI21x1_ASAP7_75t_L g1217 ( 
.A1(n_1209),
.A2(n_989),
.B(n_889),
.Y(n_1217)
);

OAI21xp33_ASAP7_75t_L g1218 ( 
.A1(n_1150),
.A2(n_949),
.B(n_945),
.Y(n_1218)
);

BUFx3_ASAP7_75t_L g1219 ( 
.A(n_1094),
.Y(n_1219)
);

AOI21xp33_ASAP7_75t_L g1220 ( 
.A1(n_1060),
.A2(n_935),
.B(n_989),
.Y(n_1220)
);

NAND2xp5_ASAP7_75t_L g1221 ( 
.A(n_1050),
.B(n_1039),
.Y(n_1221)
);

NAND2xp5_ASAP7_75t_L g1222 ( 
.A(n_1050),
.B(n_1102),
.Y(n_1222)
);

INVx2_ASAP7_75t_SL g1223 ( 
.A(n_1075),
.Y(n_1223)
);

AOI22xp33_ASAP7_75t_SL g1224 ( 
.A1(n_1207),
.A2(n_951),
.B1(n_902),
.B2(n_911),
.Y(n_1224)
);

OAI21x1_ASAP7_75t_L g1225 ( 
.A1(n_1144),
.A2(n_996),
.B(n_882),
.Y(n_1225)
);

NOR2xp33_ASAP7_75t_L g1226 ( 
.A(n_1126),
.B(n_1030),
.Y(n_1226)
);

BUFx6f_ASAP7_75t_L g1227 ( 
.A(n_1077),
.Y(n_1227)
);

AOI21xp5_ASAP7_75t_L g1228 ( 
.A1(n_1212),
.A2(n_880),
.B(n_913),
.Y(n_1228)
);

INVx1_ASAP7_75t_L g1229 ( 
.A(n_1168),
.Y(n_1229)
);

OA21x2_ASAP7_75t_L g1230 ( 
.A1(n_1141),
.A2(n_1003),
.B(n_1005),
.Y(n_1230)
);

AOI21xp5_ASAP7_75t_L g1231 ( 
.A1(n_1198),
.A2(n_1012),
.B(n_984),
.Y(n_1231)
);

O2A1O1Ixp33_ASAP7_75t_L g1232 ( 
.A1(n_1082),
.A2(n_1020),
.B(n_1026),
.C(n_1028),
.Y(n_1232)
);

AOI21xp5_ASAP7_75t_SL g1233 ( 
.A1(n_1058),
.A2(n_1034),
.B(n_1198),
.Y(n_1233)
);

AO31x2_ASAP7_75t_L g1234 ( 
.A1(n_1066),
.A2(n_1072),
.A3(n_1090),
.B(n_1196),
.Y(n_1234)
);

INVx1_ASAP7_75t_SL g1235 ( 
.A(n_1092),
.Y(n_1235)
);

OAI22xp5_ASAP7_75t_L g1236 ( 
.A1(n_1053),
.A2(n_1061),
.B1(n_1058),
.B2(n_1083),
.Y(n_1236)
);

OAI21xp5_ASAP7_75t_L g1237 ( 
.A1(n_1211),
.A2(n_1053),
.B(n_1064),
.Y(n_1237)
);

AOI21xp5_ASAP7_75t_L g1238 ( 
.A1(n_1210),
.A2(n_1206),
.B(n_1099),
.Y(n_1238)
);

OR2x2_ASAP7_75t_L g1239 ( 
.A(n_1107),
.B(n_1116),
.Y(n_1239)
);

INVxp67_ASAP7_75t_SL g1240 ( 
.A(n_1135),
.Y(n_1240)
);

A2O1A1Ixp33_ASAP7_75t_L g1241 ( 
.A1(n_1115),
.A2(n_1091),
.B(n_1071),
.C(n_1208),
.Y(n_1241)
);

INVx2_ASAP7_75t_L g1242 ( 
.A(n_1159),
.Y(n_1242)
);

AOI221xp5_ASAP7_75t_SL g1243 ( 
.A1(n_1154),
.A2(n_1183),
.B1(n_1193),
.B2(n_1080),
.C(n_1176),
.Y(n_1243)
);

INVx1_ASAP7_75t_L g1244 ( 
.A(n_1062),
.Y(n_1244)
);

OR2x6_ASAP7_75t_L g1245 ( 
.A(n_1055),
.B(n_1101),
.Y(n_1245)
);

A2O1A1Ixp33_ASAP7_75t_L g1246 ( 
.A1(n_1078),
.A2(n_1084),
.B(n_1069),
.C(n_1155),
.Y(n_1246)
);

OAI21x1_ASAP7_75t_L g1247 ( 
.A1(n_1067),
.A2(n_1106),
.B(n_1098),
.Y(n_1247)
);

INVx1_ASAP7_75t_SL g1248 ( 
.A(n_1123),
.Y(n_1248)
);

NAND2xp5_ASAP7_75t_SL g1249 ( 
.A(n_1065),
.B(n_1110),
.Y(n_1249)
);

OAI21xp5_ASAP7_75t_L g1250 ( 
.A1(n_1097),
.A2(n_1128),
.B(n_1111),
.Y(n_1250)
);

INVx1_ASAP7_75t_L g1251 ( 
.A(n_1063),
.Y(n_1251)
);

AOI21xp5_ASAP7_75t_L g1252 ( 
.A1(n_1210),
.A2(n_1206),
.B(n_1146),
.Y(n_1252)
);

OAI21xp5_ASAP7_75t_L g1253 ( 
.A1(n_1130),
.A2(n_1096),
.B(n_1089),
.Y(n_1253)
);

AOI21xp5_ASAP7_75t_L g1254 ( 
.A1(n_1146),
.A2(n_1089),
.B(n_1129),
.Y(n_1254)
);

A2O1A1Ixp33_ASAP7_75t_L g1255 ( 
.A1(n_1155),
.A2(n_1192),
.B(n_1178),
.C(n_1156),
.Y(n_1255)
);

AND2x2_ASAP7_75t_L g1256 ( 
.A(n_1173),
.B(n_1177),
.Y(n_1256)
);

AOI221x1_ASAP7_75t_L g1257 ( 
.A1(n_1130),
.A2(n_1164),
.B1(n_1136),
.B2(n_1142),
.C(n_1148),
.Y(n_1257)
);

INVx2_ASAP7_75t_SL g1258 ( 
.A(n_1190),
.Y(n_1258)
);

OAI22xp5_ASAP7_75t_L g1259 ( 
.A1(n_1048),
.A2(n_1172),
.B1(n_1088),
.B2(n_1079),
.Y(n_1259)
);

A2O1A1Ixp33_ASAP7_75t_L g1260 ( 
.A1(n_1073),
.A2(n_1095),
.B(n_1080),
.C(n_1086),
.Y(n_1260)
);

AND2x4_ASAP7_75t_L g1261 ( 
.A(n_1197),
.B(n_1052),
.Y(n_1261)
);

OAI21x1_ASAP7_75t_L g1262 ( 
.A1(n_1129),
.A2(n_1162),
.B(n_1152),
.Y(n_1262)
);

NAND2xp33_ASAP7_75t_SL g1263 ( 
.A(n_1118),
.B(n_1077),
.Y(n_1263)
);

INVx1_ASAP7_75t_L g1264 ( 
.A(n_1103),
.Y(n_1264)
);

INVx4_ASAP7_75t_L g1265 ( 
.A(n_1077),
.Y(n_1265)
);

AO31x2_ASAP7_75t_L g1266 ( 
.A1(n_1093),
.A2(n_1119),
.A3(n_1120),
.B(n_1151),
.Y(n_1266)
);

AO31x2_ASAP7_75t_L g1267 ( 
.A1(n_1151),
.A2(n_1152),
.A3(n_1162),
.B(n_1124),
.Y(n_1267)
);

AOI21xp5_ASAP7_75t_L g1268 ( 
.A1(n_1203),
.A2(n_1185),
.B(n_1187),
.Y(n_1268)
);

O2A1O1Ixp33_ASAP7_75t_L g1269 ( 
.A1(n_1085),
.A2(n_1180),
.B(n_1179),
.C(n_1171),
.Y(n_1269)
);

NAND2xp5_ASAP7_75t_L g1270 ( 
.A(n_1048),
.B(n_1191),
.Y(n_1270)
);

AO31x2_ASAP7_75t_L g1271 ( 
.A1(n_1121),
.A2(n_1165),
.A3(n_1163),
.B(n_1112),
.Y(n_1271)
);

AO31x2_ASAP7_75t_L g1272 ( 
.A1(n_1165),
.A2(n_1112),
.A3(n_1134),
.B(n_1087),
.Y(n_1272)
);

NAND2xp5_ASAP7_75t_L g1273 ( 
.A(n_1087),
.B(n_1113),
.Y(n_1273)
);

NAND2xp5_ASAP7_75t_L g1274 ( 
.A(n_1081),
.B(n_1153),
.Y(n_1274)
);

AND2x4_ASAP7_75t_L g1275 ( 
.A(n_1052),
.B(n_1054),
.Y(n_1275)
);

OAI21x1_ASAP7_75t_L g1276 ( 
.A1(n_1204),
.A2(n_1202),
.B(n_1145),
.Y(n_1276)
);

OAI21x1_ASAP7_75t_L g1277 ( 
.A1(n_1149),
.A2(n_1157),
.B(n_1049),
.Y(n_1277)
);

OAI22xp5_ASAP7_75t_L g1278 ( 
.A1(n_1167),
.A2(n_1056),
.B1(n_1109),
.B2(n_1138),
.Y(n_1278)
);

INVx1_ASAP7_75t_L g1279 ( 
.A(n_1158),
.Y(n_1279)
);

BUFx10_ASAP7_75t_L g1280 ( 
.A(n_1055),
.Y(n_1280)
);

OA21x2_ASAP7_75t_L g1281 ( 
.A1(n_1139),
.A2(n_1195),
.B(n_1188),
.Y(n_1281)
);

BUFx2_ASAP7_75t_L g1282 ( 
.A(n_1190),
.Y(n_1282)
);

INVx1_ASAP7_75t_L g1283 ( 
.A(n_1200),
.Y(n_1283)
);

O2A1O1Ixp33_ASAP7_75t_SL g1284 ( 
.A1(n_1160),
.A2(n_1169),
.B(n_1104),
.C(n_1181),
.Y(n_1284)
);

AOI21xp5_ASAP7_75t_L g1285 ( 
.A1(n_1059),
.A2(n_1133),
.B(n_1205),
.Y(n_1285)
);

BUFx6f_ASAP7_75t_L g1286 ( 
.A(n_1108),
.Y(n_1286)
);

OAI21x1_ASAP7_75t_L g1287 ( 
.A1(n_1049),
.A2(n_1114),
.B(n_1105),
.Y(n_1287)
);

AOI21xp5_ASAP7_75t_L g1288 ( 
.A1(n_1059),
.A2(n_1205),
.B(n_1114),
.Y(n_1288)
);

NOR2xp33_ASAP7_75t_L g1289 ( 
.A(n_1147),
.B(n_1132),
.Y(n_1289)
);

OAI21x1_ASAP7_75t_L g1290 ( 
.A1(n_1057),
.A2(n_1201),
.B(n_1199),
.Y(n_1290)
);

AO31x2_ASAP7_75t_L g1291 ( 
.A1(n_1199),
.A2(n_1122),
.A3(n_1140),
.B(n_1207),
.Y(n_1291)
);

AOI21xp5_ASAP7_75t_L g1292 ( 
.A1(n_1108),
.A2(n_1117),
.B(n_1194),
.Y(n_1292)
);

HB1xp67_ASAP7_75t_L g1293 ( 
.A(n_1108),
.Y(n_1293)
);

BUFx6f_ASAP7_75t_L g1294 ( 
.A(n_1117),
.Y(n_1294)
);

AO21x2_ASAP7_75t_L g1295 ( 
.A1(n_1184),
.A2(n_1122),
.B(n_1175),
.Y(n_1295)
);

AND2x2_ASAP7_75t_L g1296 ( 
.A(n_1184),
.B(n_1175),
.Y(n_1296)
);

OAI22x1_ASAP7_75t_L g1297 ( 
.A1(n_1166),
.A2(n_1186),
.B1(n_1161),
.B2(n_1055),
.Y(n_1297)
);

NAND2xp5_ASAP7_75t_L g1298 ( 
.A(n_1117),
.B(n_1194),
.Y(n_1298)
);

OAI21x1_ASAP7_75t_L g1299 ( 
.A1(n_1182),
.A2(n_1127),
.B(n_1170),
.Y(n_1299)
);

BUFx2_ASAP7_75t_L g1300 ( 
.A(n_1137),
.Y(n_1300)
);

AOI21xp33_ASAP7_75t_L g1301 ( 
.A1(n_1166),
.A2(n_1127),
.B(n_1170),
.Y(n_1301)
);

AND2x4_ASAP7_75t_L g1302 ( 
.A(n_1125),
.B(n_1170),
.Y(n_1302)
);

OAI21x1_ASAP7_75t_L g1303 ( 
.A1(n_1182),
.A2(n_1166),
.B(n_1131),
.Y(n_1303)
);

CKINVDCx11_ASAP7_75t_R g1304 ( 
.A(n_1068),
.Y(n_1304)
);

INVx4_ASAP7_75t_L g1305 ( 
.A(n_1076),
.Y(n_1305)
);

INVx1_ASAP7_75t_L g1306 ( 
.A(n_1074),
.Y(n_1306)
);

NOR2xp67_ASAP7_75t_L g1307 ( 
.A(n_1076),
.B(n_712),
.Y(n_1307)
);

OAI22x1_ASAP7_75t_L g1308 ( 
.A1(n_1126),
.A2(n_696),
.B1(n_1143),
.B2(n_1150),
.Y(n_1308)
);

INVx2_ASAP7_75t_L g1309 ( 
.A(n_1168),
.Y(n_1309)
);

BUFx6f_ASAP7_75t_L g1310 ( 
.A(n_1077),
.Y(n_1310)
);

BUFx6f_ASAP7_75t_L g1311 ( 
.A(n_1077),
.Y(n_1311)
);

INVx1_ASAP7_75t_L g1312 ( 
.A(n_1168),
.Y(n_1312)
);

INVx2_ASAP7_75t_L g1313 ( 
.A(n_1168),
.Y(n_1313)
);

AO31x2_ASAP7_75t_L g1314 ( 
.A1(n_1070),
.A2(n_868),
.A3(n_928),
.B(n_1189),
.Y(n_1314)
);

AOI21xp5_ASAP7_75t_L g1315 ( 
.A1(n_1070),
.A2(n_746),
.B(n_695),
.Y(n_1315)
);

OA21x2_ASAP7_75t_L g1316 ( 
.A1(n_1070),
.A2(n_1141),
.B(n_1212),
.Y(n_1316)
);

AOI21xp5_ASAP7_75t_L g1317 ( 
.A1(n_1070),
.A2(n_746),
.B(n_695),
.Y(n_1317)
);

INVx4_ASAP7_75t_L g1318 ( 
.A(n_1077),
.Y(n_1318)
);

OAI21xp5_ASAP7_75t_L g1319 ( 
.A1(n_1051),
.A2(n_1212),
.B(n_1189),
.Y(n_1319)
);

OAI21xp5_ASAP7_75t_L g1320 ( 
.A1(n_1051),
.A2(n_1212),
.B(n_1189),
.Y(n_1320)
);

AO32x2_ASAP7_75t_L g1321 ( 
.A1(n_1193),
.A2(n_895),
.A3(n_1167),
.B1(n_1171),
.B2(n_1002),
.Y(n_1321)
);

INVx5_ASAP7_75t_L g1322 ( 
.A(n_1077),
.Y(n_1322)
);

AO31x2_ASAP7_75t_L g1323 ( 
.A1(n_1070),
.A2(n_868),
.A3(n_928),
.B(n_1189),
.Y(n_1323)
);

OAI22xp5_ASAP7_75t_L g1324 ( 
.A1(n_1102),
.A2(n_696),
.B1(n_1060),
.B2(n_1050),
.Y(n_1324)
);

OAI21x1_ASAP7_75t_L g1325 ( 
.A1(n_1144),
.A2(n_1100),
.B(n_1067),
.Y(n_1325)
);

AOI21xp5_ASAP7_75t_L g1326 ( 
.A1(n_1070),
.A2(n_746),
.B(n_695),
.Y(n_1326)
);

OAI21x1_ASAP7_75t_L g1327 ( 
.A1(n_1144),
.A2(n_1100),
.B(n_1067),
.Y(n_1327)
);

AND2x4_ASAP7_75t_L g1328 ( 
.A(n_1173),
.B(n_1036),
.Y(n_1328)
);

OAI21x1_ASAP7_75t_L g1329 ( 
.A1(n_1144),
.A2(n_1100),
.B(n_1067),
.Y(n_1329)
);

INVxp67_ASAP7_75t_L g1330 ( 
.A(n_1075),
.Y(n_1330)
);

NAND2xp5_ASAP7_75t_SL g1331 ( 
.A(n_1082),
.B(n_696),
.Y(n_1331)
);

AOI21xp5_ASAP7_75t_L g1332 ( 
.A1(n_1070),
.A2(n_746),
.B(n_695),
.Y(n_1332)
);

INVx2_ASAP7_75t_L g1333 ( 
.A(n_1168),
.Y(n_1333)
);

AND2x4_ASAP7_75t_L g1334 ( 
.A(n_1173),
.B(n_1036),
.Y(n_1334)
);

AOI21xp5_ASAP7_75t_L g1335 ( 
.A1(n_1070),
.A2(n_746),
.B(n_695),
.Y(n_1335)
);

NAND2xp5_ASAP7_75t_L g1336 ( 
.A(n_1050),
.B(n_696),
.Y(n_1336)
);

INVx1_ASAP7_75t_L g1337 ( 
.A(n_1168),
.Y(n_1337)
);

INVx2_ASAP7_75t_L g1338 ( 
.A(n_1168),
.Y(n_1338)
);

AOI21xp5_ASAP7_75t_L g1339 ( 
.A1(n_1070),
.A2(n_746),
.B(n_695),
.Y(n_1339)
);

BUFx8_ASAP7_75t_L g1340 ( 
.A(n_1068),
.Y(n_1340)
);

BUFx6f_ASAP7_75t_L g1341 ( 
.A(n_1077),
.Y(n_1341)
);

AOI21xp5_ASAP7_75t_L g1342 ( 
.A1(n_1070),
.A2(n_746),
.B(n_695),
.Y(n_1342)
);

AOI21x1_ASAP7_75t_L g1343 ( 
.A1(n_1209),
.A2(n_1196),
.B(n_1090),
.Y(n_1343)
);

INVx5_ASAP7_75t_L g1344 ( 
.A(n_1077),
.Y(n_1344)
);

NAND2xp33_ASAP7_75t_L g1345 ( 
.A(n_1060),
.B(n_916),
.Y(n_1345)
);

NAND2xp5_ASAP7_75t_L g1346 ( 
.A(n_1050),
.B(n_696),
.Y(n_1346)
);

OAI22xp5_ASAP7_75t_L g1347 ( 
.A1(n_1102),
.A2(n_696),
.B1(n_1060),
.B2(n_1050),
.Y(n_1347)
);

INVx2_ASAP7_75t_SL g1348 ( 
.A(n_1094),
.Y(n_1348)
);

BUFx3_ASAP7_75t_L g1349 ( 
.A(n_1094),
.Y(n_1349)
);

NOR2xp33_ASAP7_75t_SL g1350 ( 
.A(n_1207),
.B(n_756),
.Y(n_1350)
);

A2O1A1Ixp33_ASAP7_75t_L g1351 ( 
.A1(n_1143),
.A2(n_696),
.B(n_922),
.C(n_916),
.Y(n_1351)
);

BUFx2_ASAP7_75t_L g1352 ( 
.A(n_1075),
.Y(n_1352)
);

AOI21xp5_ASAP7_75t_L g1353 ( 
.A1(n_1070),
.A2(n_746),
.B(n_695),
.Y(n_1353)
);

INVx1_ASAP7_75t_L g1354 ( 
.A(n_1168),
.Y(n_1354)
);

HB1xp67_ASAP7_75t_L g1355 ( 
.A(n_1075),
.Y(n_1355)
);

NAND2xp5_ASAP7_75t_L g1356 ( 
.A(n_1050),
.B(n_696),
.Y(n_1356)
);

INVx1_ASAP7_75t_L g1357 ( 
.A(n_1168),
.Y(n_1357)
);

A2O1A1Ixp33_ASAP7_75t_L g1358 ( 
.A1(n_1143),
.A2(n_696),
.B(n_922),
.C(n_916),
.Y(n_1358)
);

BUFx4f_ASAP7_75t_L g1359 ( 
.A(n_1068),
.Y(n_1359)
);

A2O1A1Ixp33_ASAP7_75t_L g1360 ( 
.A1(n_1143),
.A2(n_696),
.B(n_922),
.C(n_916),
.Y(n_1360)
);

OAI21x1_ASAP7_75t_L g1361 ( 
.A1(n_1144),
.A2(n_1100),
.B(n_1067),
.Y(n_1361)
);

NAND3xp33_ASAP7_75t_SL g1362 ( 
.A(n_1143),
.B(n_696),
.C(n_916),
.Y(n_1362)
);

BUFx10_ASAP7_75t_L g1363 ( 
.A(n_1150),
.Y(n_1363)
);

AOI21xp5_ASAP7_75t_L g1364 ( 
.A1(n_1070),
.A2(n_746),
.B(n_695),
.Y(n_1364)
);

O2A1O1Ixp33_ASAP7_75t_L g1365 ( 
.A1(n_1143),
.A2(n_916),
.B(n_929),
.C(n_780),
.Y(n_1365)
);

OAI21x1_ASAP7_75t_L g1366 ( 
.A1(n_1144),
.A2(n_1100),
.B(n_1067),
.Y(n_1366)
);

INVx1_ASAP7_75t_L g1367 ( 
.A(n_1168),
.Y(n_1367)
);

AOI21xp5_ASAP7_75t_L g1368 ( 
.A1(n_1070),
.A2(n_746),
.B(n_695),
.Y(n_1368)
);

INVx1_ASAP7_75t_SL g1369 ( 
.A(n_1075),
.Y(n_1369)
);

AOI21xp5_ASAP7_75t_L g1370 ( 
.A1(n_1070),
.A2(n_746),
.B(n_695),
.Y(n_1370)
);

AO31x2_ASAP7_75t_L g1371 ( 
.A1(n_1070),
.A2(n_868),
.A3(n_928),
.B(n_1189),
.Y(n_1371)
);

OAI21x1_ASAP7_75t_L g1372 ( 
.A1(n_1144),
.A2(n_1100),
.B(n_1067),
.Y(n_1372)
);

OA21x2_ASAP7_75t_L g1373 ( 
.A1(n_1070),
.A2(n_1141),
.B(n_1212),
.Y(n_1373)
);

INVx6_ASAP7_75t_L g1374 ( 
.A(n_1280),
.Y(n_1374)
);

AOI22xp33_ASAP7_75t_L g1375 ( 
.A1(n_1345),
.A2(n_1362),
.B1(n_1308),
.B2(n_1331),
.Y(n_1375)
);

CKINVDCx5p33_ASAP7_75t_R g1376 ( 
.A(n_1304),
.Y(n_1376)
);

CKINVDCx20_ASAP7_75t_R g1377 ( 
.A(n_1340),
.Y(n_1377)
);

CKINVDCx5p33_ASAP7_75t_R g1378 ( 
.A(n_1340),
.Y(n_1378)
);

INVx6_ASAP7_75t_L g1379 ( 
.A(n_1280),
.Y(n_1379)
);

CKINVDCx6p67_ASAP7_75t_R g1380 ( 
.A(n_1245),
.Y(n_1380)
);

INVx2_ASAP7_75t_L g1381 ( 
.A(n_1309),
.Y(n_1381)
);

OAI22x1_ASAP7_75t_L g1382 ( 
.A1(n_1249),
.A2(n_1226),
.B1(n_1356),
.B2(n_1336),
.Y(n_1382)
);

INVx2_ASAP7_75t_L g1383 ( 
.A(n_1313),
.Y(n_1383)
);

BUFx4_ASAP7_75t_SL g1384 ( 
.A(n_1245),
.Y(n_1384)
);

INVx2_ASAP7_75t_L g1385 ( 
.A(n_1333),
.Y(n_1385)
);

AOI22xp33_ASAP7_75t_L g1386 ( 
.A1(n_1324),
.A2(n_1347),
.B1(n_1236),
.B2(n_1346),
.Y(n_1386)
);

INVx1_ASAP7_75t_L g1387 ( 
.A(n_1338),
.Y(n_1387)
);

INVx2_ASAP7_75t_SL g1388 ( 
.A(n_1219),
.Y(n_1388)
);

CKINVDCx5p33_ASAP7_75t_R g1389 ( 
.A(n_1359),
.Y(n_1389)
);

INVx2_ASAP7_75t_L g1390 ( 
.A(n_1242),
.Y(n_1390)
);

BUFx6f_ASAP7_75t_L g1391 ( 
.A(n_1322),
.Y(n_1391)
);

INVx1_ASAP7_75t_SL g1392 ( 
.A(n_1369),
.Y(n_1392)
);

CKINVDCx6p67_ASAP7_75t_R g1393 ( 
.A(n_1245),
.Y(n_1393)
);

OAI21xp33_ASAP7_75t_L g1394 ( 
.A1(n_1351),
.A2(n_1360),
.B(n_1358),
.Y(n_1394)
);

INVx6_ASAP7_75t_L g1395 ( 
.A(n_1322),
.Y(n_1395)
);

NAND2xp5_ASAP7_75t_L g1396 ( 
.A(n_1222),
.B(n_1270),
.Y(n_1396)
);

CKINVDCx11_ASAP7_75t_R g1397 ( 
.A(n_1305),
.Y(n_1397)
);

BUFx12f_ASAP7_75t_L g1398 ( 
.A(n_1305),
.Y(n_1398)
);

INVx6_ASAP7_75t_L g1399 ( 
.A(n_1322),
.Y(n_1399)
);

INVx1_ASAP7_75t_L g1400 ( 
.A(n_1229),
.Y(n_1400)
);

INVx1_ASAP7_75t_L g1401 ( 
.A(n_1312),
.Y(n_1401)
);

NAND2x1p5_ASAP7_75t_L g1402 ( 
.A(n_1344),
.B(n_1290),
.Y(n_1402)
);

INVx4_ASAP7_75t_L g1403 ( 
.A(n_1344),
.Y(n_1403)
);

CKINVDCx11_ASAP7_75t_R g1404 ( 
.A(n_1300),
.Y(n_1404)
);

OAI22xp5_ASAP7_75t_SL g1405 ( 
.A1(n_1278),
.A2(n_1297),
.B1(n_1306),
.B2(n_1289),
.Y(n_1405)
);

INVx6_ASAP7_75t_L g1406 ( 
.A(n_1344),
.Y(n_1406)
);

AOI22xp33_ASAP7_75t_L g1407 ( 
.A1(n_1324),
.A2(n_1347),
.B1(n_1236),
.B2(n_1237),
.Y(n_1407)
);

BUFx2_ASAP7_75t_SL g1408 ( 
.A(n_1349),
.Y(n_1408)
);

OAI22xp5_ASAP7_75t_L g1409 ( 
.A1(n_1241),
.A2(n_1365),
.B1(n_1240),
.B2(n_1270),
.Y(n_1409)
);

BUFx6f_ASAP7_75t_L g1410 ( 
.A(n_1227),
.Y(n_1410)
);

BUFx12f_ASAP7_75t_L g1411 ( 
.A(n_1282),
.Y(n_1411)
);

INVx6_ASAP7_75t_L g1412 ( 
.A(n_1265),
.Y(n_1412)
);

OAI22x1_ASAP7_75t_L g1413 ( 
.A1(n_1235),
.A2(n_1248),
.B1(n_1274),
.B2(n_1352),
.Y(n_1413)
);

INVx1_ASAP7_75t_L g1414 ( 
.A(n_1337),
.Y(n_1414)
);

BUFx3_ASAP7_75t_L g1415 ( 
.A(n_1348),
.Y(n_1415)
);

INVx1_ASAP7_75t_L g1416 ( 
.A(n_1354),
.Y(n_1416)
);

OAI21xp33_ASAP7_75t_L g1417 ( 
.A1(n_1350),
.A2(n_1260),
.B(n_1246),
.Y(n_1417)
);

INVx6_ASAP7_75t_L g1418 ( 
.A(n_1318),
.Y(n_1418)
);

AOI22xp33_ASAP7_75t_L g1419 ( 
.A1(n_1237),
.A2(n_1363),
.B1(n_1278),
.B2(n_1350),
.Y(n_1419)
);

AOI22xp5_ASAP7_75t_L g1420 ( 
.A1(n_1307),
.A2(n_1363),
.B1(n_1256),
.B2(n_1296),
.Y(n_1420)
);

AOI22xp33_ASAP7_75t_L g1421 ( 
.A1(n_1295),
.A2(n_1320),
.B1(n_1319),
.B2(n_1259),
.Y(n_1421)
);

AOI22xp5_ASAP7_75t_L g1422 ( 
.A1(n_1307),
.A2(n_1334),
.B1(n_1328),
.B2(n_1243),
.Y(n_1422)
);

CKINVDCx20_ASAP7_75t_R g1423 ( 
.A(n_1359),
.Y(n_1423)
);

OAI21xp33_ASAP7_75t_SL g1424 ( 
.A1(n_1273),
.A2(n_1274),
.B(n_1221),
.Y(n_1424)
);

INVx3_ASAP7_75t_L g1425 ( 
.A(n_1227),
.Y(n_1425)
);

NAND2xp5_ASAP7_75t_L g1426 ( 
.A(n_1273),
.B(n_1239),
.Y(n_1426)
);

INVx2_ASAP7_75t_L g1427 ( 
.A(n_1357),
.Y(n_1427)
);

AND2x4_ASAP7_75t_L g1428 ( 
.A(n_1302),
.B(n_1261),
.Y(n_1428)
);

INVx1_ASAP7_75t_L g1429 ( 
.A(n_1367),
.Y(n_1429)
);

INVx1_ASAP7_75t_L g1430 ( 
.A(n_1244),
.Y(n_1430)
);

AOI22xp33_ASAP7_75t_L g1431 ( 
.A1(n_1295),
.A2(n_1320),
.B1(n_1319),
.B2(n_1259),
.Y(n_1431)
);

AOI22xp33_ASAP7_75t_L g1432 ( 
.A1(n_1218),
.A2(n_1220),
.B1(n_1279),
.B2(n_1252),
.Y(n_1432)
);

INVx1_ASAP7_75t_SL g1433 ( 
.A(n_1248),
.Y(n_1433)
);

INVx4_ASAP7_75t_L g1434 ( 
.A(n_1227),
.Y(n_1434)
);

AOI22xp33_ASAP7_75t_L g1435 ( 
.A1(n_1218),
.A2(n_1220),
.B1(n_1264),
.B2(n_1251),
.Y(n_1435)
);

CKINVDCx8_ASAP7_75t_R g1436 ( 
.A(n_1302),
.Y(n_1436)
);

BUFx6f_ASAP7_75t_L g1437 ( 
.A(n_1286),
.Y(n_1437)
);

INVx3_ASAP7_75t_SL g1438 ( 
.A(n_1261),
.Y(n_1438)
);

INVx2_ASAP7_75t_L g1439 ( 
.A(n_1281),
.Y(n_1439)
);

BUFx4f_ASAP7_75t_SL g1440 ( 
.A(n_1258),
.Y(n_1440)
);

CKINVDCx20_ASAP7_75t_R g1441 ( 
.A(n_1263),
.Y(n_1441)
);

AOI22xp33_ASAP7_75t_SL g1442 ( 
.A1(n_1316),
.A2(n_1373),
.B1(n_1303),
.B2(n_1291),
.Y(n_1442)
);

BUFx3_ASAP7_75t_L g1443 ( 
.A(n_1223),
.Y(n_1443)
);

INVxp67_ASAP7_75t_L g1444 ( 
.A(n_1283),
.Y(n_1444)
);

INVx1_ASAP7_75t_L g1445 ( 
.A(n_1298),
.Y(n_1445)
);

AOI22xp5_ASAP7_75t_L g1446 ( 
.A1(n_1328),
.A2(n_1334),
.B1(n_1243),
.B2(n_1275),
.Y(n_1446)
);

AOI22xp33_ASAP7_75t_L g1447 ( 
.A1(n_1238),
.A2(n_1373),
.B1(n_1316),
.B2(n_1268),
.Y(n_1447)
);

BUFx5_ASAP7_75t_L g1448 ( 
.A(n_1343),
.Y(n_1448)
);

BUFx8_ASAP7_75t_L g1449 ( 
.A(n_1286),
.Y(n_1449)
);

INVx1_ASAP7_75t_L g1450 ( 
.A(n_1299),
.Y(n_1450)
);

OAI22xp5_ASAP7_75t_L g1451 ( 
.A1(n_1255),
.A2(n_1330),
.B1(n_1269),
.B2(n_1275),
.Y(n_1451)
);

AOI22xp33_ASAP7_75t_SL g1452 ( 
.A1(n_1291),
.A2(n_1321),
.B1(n_1216),
.B2(n_1213),
.Y(n_1452)
);

NAND2xp5_ASAP7_75t_L g1453 ( 
.A(n_1254),
.B(n_1301),
.Y(n_1453)
);

INVx2_ASAP7_75t_L g1454 ( 
.A(n_1287),
.Y(n_1454)
);

INVx1_ASAP7_75t_L g1455 ( 
.A(n_1291),
.Y(n_1455)
);

INVx6_ASAP7_75t_L g1456 ( 
.A(n_1286),
.Y(n_1456)
);

AOI22xp33_ASAP7_75t_L g1457 ( 
.A1(n_1301),
.A2(n_1213),
.B1(n_1253),
.B2(n_1216),
.Y(n_1457)
);

CKINVDCx6p67_ASAP7_75t_R g1458 ( 
.A(n_1294),
.Y(n_1458)
);

NAND2xp5_ASAP7_75t_L g1459 ( 
.A(n_1233),
.B(n_1293),
.Y(n_1459)
);

INVx6_ASAP7_75t_L g1460 ( 
.A(n_1294),
.Y(n_1460)
);

NAND2xp5_ASAP7_75t_L g1461 ( 
.A(n_1272),
.B(n_1214),
.Y(n_1461)
);

BUFx2_ASAP7_75t_L g1462 ( 
.A(n_1294),
.Y(n_1462)
);

AOI22xp33_ASAP7_75t_L g1463 ( 
.A1(n_1224),
.A2(n_1253),
.B1(n_1250),
.B2(n_1288),
.Y(n_1463)
);

AOI22xp33_ASAP7_75t_SL g1464 ( 
.A1(n_1321),
.A2(n_1230),
.B1(n_1250),
.B2(n_1257),
.Y(n_1464)
);

BUFx2_ASAP7_75t_SL g1465 ( 
.A(n_1310),
.Y(n_1465)
);

BUFx8_ASAP7_75t_SL g1466 ( 
.A(n_1310),
.Y(n_1466)
);

CKINVDCx11_ASAP7_75t_R g1467 ( 
.A(n_1311),
.Y(n_1467)
);

AOI22xp33_ASAP7_75t_L g1468 ( 
.A1(n_1321),
.A2(n_1230),
.B1(n_1262),
.B2(n_1231),
.Y(n_1468)
);

OAI22xp33_ASAP7_75t_L g1469 ( 
.A1(n_1215),
.A2(n_1285),
.B1(n_1217),
.B2(n_1311),
.Y(n_1469)
);

AOI22xp33_ASAP7_75t_SL g1470 ( 
.A1(n_1214),
.A2(n_1341),
.B1(n_1311),
.B2(n_1276),
.Y(n_1470)
);

INVx6_ASAP7_75t_L g1471 ( 
.A(n_1341),
.Y(n_1471)
);

INVx2_ASAP7_75t_SL g1472 ( 
.A(n_1341),
.Y(n_1472)
);

INVx3_ASAP7_75t_SL g1473 ( 
.A(n_1292),
.Y(n_1473)
);

BUFx6f_ASAP7_75t_L g1474 ( 
.A(n_1277),
.Y(n_1474)
);

BUFx4f_ASAP7_75t_SL g1475 ( 
.A(n_1284),
.Y(n_1475)
);

INVx6_ASAP7_75t_L g1476 ( 
.A(n_1272),
.Y(n_1476)
);

AOI22xp33_ASAP7_75t_L g1477 ( 
.A1(n_1228),
.A2(n_1326),
.B1(n_1370),
.B2(n_1368),
.Y(n_1477)
);

OAI22xp33_ASAP7_75t_L g1478 ( 
.A1(n_1315),
.A2(n_1339),
.B1(n_1335),
.B2(n_1332),
.Y(n_1478)
);

AOI22xp33_ASAP7_75t_L g1479 ( 
.A1(n_1317),
.A2(n_1342),
.B1(n_1353),
.B2(n_1364),
.Y(n_1479)
);

AOI22xp33_ASAP7_75t_L g1480 ( 
.A1(n_1247),
.A2(n_1372),
.B1(n_1325),
.B2(n_1366),
.Y(n_1480)
);

AOI22xp33_ASAP7_75t_L g1481 ( 
.A1(n_1327),
.A2(n_1361),
.B1(n_1329),
.B2(n_1225),
.Y(n_1481)
);

BUFx4_ASAP7_75t_R g1482 ( 
.A(n_1232),
.Y(n_1482)
);

AND2x2_ASAP7_75t_L g1483 ( 
.A(n_1314),
.B(n_1371),
.Y(n_1483)
);

INVx6_ASAP7_75t_L g1484 ( 
.A(n_1234),
.Y(n_1484)
);

INVxp67_ASAP7_75t_L g1485 ( 
.A(n_1314),
.Y(n_1485)
);

INVx1_ASAP7_75t_SL g1486 ( 
.A(n_1371),
.Y(n_1486)
);

BUFx6f_ASAP7_75t_L g1487 ( 
.A(n_1234),
.Y(n_1487)
);

NAND2xp33_ASAP7_75t_R g1488 ( 
.A(n_1314),
.B(n_1371),
.Y(n_1488)
);

AOI22xp33_ASAP7_75t_L g1489 ( 
.A1(n_1323),
.A2(n_1266),
.B1(n_1267),
.B2(n_1271),
.Y(n_1489)
);

BUFx3_ASAP7_75t_L g1490 ( 
.A(n_1323),
.Y(n_1490)
);

CKINVDCx16_ASAP7_75t_R g1491 ( 
.A(n_1267),
.Y(n_1491)
);

OAI22xp5_ASAP7_75t_L g1492 ( 
.A1(n_1266),
.A2(n_696),
.B1(n_1358),
.B2(n_1351),
.Y(n_1492)
);

BUFx10_ASAP7_75t_L g1493 ( 
.A(n_1271),
.Y(n_1493)
);

AOI22xp33_ASAP7_75t_SL g1494 ( 
.A1(n_1271),
.A2(n_494),
.B1(n_1345),
.B2(n_1143),
.Y(n_1494)
);

AOI22xp33_ASAP7_75t_L g1495 ( 
.A1(n_1345),
.A2(n_1362),
.B1(n_916),
.B2(n_1308),
.Y(n_1495)
);

AOI22xp33_ASAP7_75t_L g1496 ( 
.A1(n_1345),
.A2(n_1362),
.B1(n_916),
.B2(n_1308),
.Y(n_1496)
);

INVxp67_ASAP7_75t_L g1497 ( 
.A(n_1355),
.Y(n_1497)
);

AOI22xp33_ASAP7_75t_SL g1498 ( 
.A1(n_1345),
.A2(n_494),
.B1(n_1143),
.B2(n_1350),
.Y(n_1498)
);

INVx1_ASAP7_75t_L g1499 ( 
.A(n_1309),
.Y(n_1499)
);

AOI22xp33_ASAP7_75t_SL g1500 ( 
.A1(n_1345),
.A2(n_494),
.B1(n_1143),
.B2(n_1350),
.Y(n_1500)
);

AOI22xp33_ASAP7_75t_L g1501 ( 
.A1(n_1345),
.A2(n_1362),
.B1(n_916),
.B2(n_1308),
.Y(n_1501)
);

INVx1_ASAP7_75t_L g1502 ( 
.A(n_1309),
.Y(n_1502)
);

OAI22xp5_ASAP7_75t_L g1503 ( 
.A1(n_1351),
.A2(n_696),
.B1(n_1360),
.B2(n_1358),
.Y(n_1503)
);

CKINVDCx5p33_ASAP7_75t_R g1504 ( 
.A(n_1304),
.Y(n_1504)
);

CKINVDCx20_ASAP7_75t_R g1505 ( 
.A(n_1304),
.Y(n_1505)
);

INVx1_ASAP7_75t_L g1506 ( 
.A(n_1309),
.Y(n_1506)
);

INVx1_ASAP7_75t_L g1507 ( 
.A(n_1309),
.Y(n_1507)
);

AND2x2_ASAP7_75t_L g1508 ( 
.A(n_1386),
.B(n_1495),
.Y(n_1508)
);

OAI21x1_ASAP7_75t_L g1509 ( 
.A1(n_1481),
.A2(n_1480),
.B(n_1477),
.Y(n_1509)
);

OR2x2_ASAP7_75t_L g1510 ( 
.A(n_1491),
.B(n_1461),
.Y(n_1510)
);

AND2x2_ASAP7_75t_L g1511 ( 
.A(n_1386),
.B(n_1495),
.Y(n_1511)
);

OR2x2_ASAP7_75t_L g1512 ( 
.A(n_1421),
.B(n_1431),
.Y(n_1512)
);

INVx2_ASAP7_75t_L g1513 ( 
.A(n_1439),
.Y(n_1513)
);

BUFx3_ASAP7_75t_L g1514 ( 
.A(n_1374),
.Y(n_1514)
);

AOI22xp33_ASAP7_75t_L g1515 ( 
.A1(n_1394),
.A2(n_1498),
.B1(n_1500),
.B2(n_1503),
.Y(n_1515)
);

OAI21x1_ASAP7_75t_L g1516 ( 
.A1(n_1481),
.A2(n_1479),
.B(n_1447),
.Y(n_1516)
);

AOI21x1_ASAP7_75t_L g1517 ( 
.A1(n_1492),
.A2(n_1453),
.B(n_1409),
.Y(n_1517)
);

AOI21x1_ASAP7_75t_L g1518 ( 
.A1(n_1382),
.A2(n_1459),
.B(n_1454),
.Y(n_1518)
);

AND2x4_ASAP7_75t_L g1519 ( 
.A(n_1450),
.B(n_1490),
.Y(n_1519)
);

INVx8_ASAP7_75t_L g1520 ( 
.A(n_1466),
.Y(n_1520)
);

BUFx3_ASAP7_75t_L g1521 ( 
.A(n_1380),
.Y(n_1521)
);

INVx2_ASAP7_75t_L g1522 ( 
.A(n_1427),
.Y(n_1522)
);

BUFx3_ASAP7_75t_L g1523 ( 
.A(n_1374),
.Y(n_1523)
);

OR2x2_ASAP7_75t_L g1524 ( 
.A(n_1421),
.B(n_1431),
.Y(n_1524)
);

INVx2_ASAP7_75t_L g1525 ( 
.A(n_1400),
.Y(n_1525)
);

INVx1_ASAP7_75t_L g1526 ( 
.A(n_1455),
.Y(n_1526)
);

INVx2_ASAP7_75t_L g1527 ( 
.A(n_1401),
.Y(n_1527)
);

BUFx2_ASAP7_75t_SL g1528 ( 
.A(n_1391),
.Y(n_1528)
);

BUFx8_ASAP7_75t_L g1529 ( 
.A(n_1398),
.Y(n_1529)
);

BUFx3_ASAP7_75t_L g1530 ( 
.A(n_1393),
.Y(n_1530)
);

OAI21xp5_ASAP7_75t_L g1531 ( 
.A1(n_1496),
.A2(n_1501),
.B(n_1375),
.Y(n_1531)
);

AND2x2_ASAP7_75t_L g1532 ( 
.A(n_1496),
.B(n_1501),
.Y(n_1532)
);

OAI21x1_ASAP7_75t_L g1533 ( 
.A1(n_1468),
.A2(n_1463),
.B(n_1489),
.Y(n_1533)
);

INVx1_ASAP7_75t_L g1534 ( 
.A(n_1483),
.Y(n_1534)
);

OAI21x1_ASAP7_75t_L g1535 ( 
.A1(n_1468),
.A2(n_1489),
.B(n_1432),
.Y(n_1535)
);

INVx3_ASAP7_75t_L g1536 ( 
.A(n_1474),
.Y(n_1536)
);

OR2x2_ASAP7_75t_L g1537 ( 
.A(n_1407),
.B(n_1485),
.Y(n_1537)
);

AO31x2_ASAP7_75t_L g1538 ( 
.A1(n_1413),
.A2(n_1451),
.A3(n_1464),
.B(n_1488),
.Y(n_1538)
);

INVx2_ASAP7_75t_L g1539 ( 
.A(n_1414),
.Y(n_1539)
);

INVx2_ASAP7_75t_L g1540 ( 
.A(n_1416),
.Y(n_1540)
);

INVx2_ASAP7_75t_SL g1541 ( 
.A(n_1384),
.Y(n_1541)
);

INVx1_ASAP7_75t_L g1542 ( 
.A(n_1476),
.Y(n_1542)
);

OAI21xp5_ASAP7_75t_L g1543 ( 
.A1(n_1498),
.A2(n_1500),
.B(n_1407),
.Y(n_1543)
);

CKINVDCx5p33_ASAP7_75t_R g1544 ( 
.A(n_1376),
.Y(n_1544)
);

AO21x2_ASAP7_75t_L g1545 ( 
.A1(n_1478),
.A2(n_1469),
.B(n_1485),
.Y(n_1545)
);

INVx2_ASAP7_75t_L g1546 ( 
.A(n_1429),
.Y(n_1546)
);

CKINVDCx5p33_ASAP7_75t_R g1547 ( 
.A(n_1504),
.Y(n_1547)
);

INVx1_ASAP7_75t_L g1548 ( 
.A(n_1486),
.Y(n_1548)
);

OAI22xp33_ASAP7_75t_L g1549 ( 
.A1(n_1420),
.A2(n_1475),
.B1(n_1422),
.B2(n_1396),
.Y(n_1549)
);

INVx2_ASAP7_75t_L g1550 ( 
.A(n_1430),
.Y(n_1550)
);

INVx3_ASAP7_75t_L g1551 ( 
.A(n_1487),
.Y(n_1551)
);

AO21x2_ASAP7_75t_L g1552 ( 
.A1(n_1478),
.A2(n_1469),
.B(n_1417),
.Y(n_1552)
);

INVx1_ASAP7_75t_L g1553 ( 
.A(n_1484),
.Y(n_1553)
);

AO31x2_ASAP7_75t_L g1554 ( 
.A1(n_1464),
.A2(n_1452),
.A3(n_1493),
.B(n_1494),
.Y(n_1554)
);

AND2x2_ASAP7_75t_L g1555 ( 
.A(n_1457),
.B(n_1494),
.Y(n_1555)
);

OR2x6_ASAP7_75t_L g1556 ( 
.A(n_1402),
.B(n_1482),
.Y(n_1556)
);

INVx1_ASAP7_75t_L g1557 ( 
.A(n_1424),
.Y(n_1557)
);

INVx2_ASAP7_75t_L g1558 ( 
.A(n_1387),
.Y(n_1558)
);

INVx2_ASAP7_75t_L g1559 ( 
.A(n_1499),
.Y(n_1559)
);

INVx1_ASAP7_75t_L g1560 ( 
.A(n_1448),
.Y(n_1560)
);

AND2x4_ASAP7_75t_L g1561 ( 
.A(n_1446),
.B(n_1457),
.Y(n_1561)
);

INVx1_ASAP7_75t_L g1562 ( 
.A(n_1448),
.Y(n_1562)
);

AOI22xp33_ASAP7_75t_SL g1563 ( 
.A1(n_1475),
.A2(n_1405),
.B1(n_1419),
.B2(n_1441),
.Y(n_1563)
);

OR2x2_ASAP7_75t_L g1564 ( 
.A(n_1435),
.B(n_1426),
.Y(n_1564)
);

INVx2_ASAP7_75t_L g1565 ( 
.A(n_1502),
.Y(n_1565)
);

INVx2_ASAP7_75t_L g1566 ( 
.A(n_1506),
.Y(n_1566)
);

AND2x4_ASAP7_75t_L g1567 ( 
.A(n_1507),
.B(n_1383),
.Y(n_1567)
);

BUFx2_ASAP7_75t_L g1568 ( 
.A(n_1497),
.Y(n_1568)
);

INVx2_ASAP7_75t_L g1569 ( 
.A(n_1381),
.Y(n_1569)
);

INVx1_ASAP7_75t_L g1570 ( 
.A(n_1442),
.Y(n_1570)
);

NAND2xp5_ASAP7_75t_L g1571 ( 
.A(n_1445),
.B(n_1392),
.Y(n_1571)
);

OR2x2_ASAP7_75t_L g1572 ( 
.A(n_1435),
.B(n_1432),
.Y(n_1572)
);

AND2x2_ASAP7_75t_L g1573 ( 
.A(n_1442),
.B(n_1385),
.Y(n_1573)
);

AO21x2_ASAP7_75t_L g1574 ( 
.A1(n_1470),
.A2(n_1390),
.B(n_1444),
.Y(n_1574)
);

INVx1_ASAP7_75t_L g1575 ( 
.A(n_1470),
.Y(n_1575)
);

OR2x6_ASAP7_75t_L g1576 ( 
.A(n_1402),
.B(n_1408),
.Y(n_1576)
);

INVx2_ASAP7_75t_L g1577 ( 
.A(n_1444),
.Y(n_1577)
);

AO21x2_ASAP7_75t_L g1578 ( 
.A1(n_1497),
.A2(n_1473),
.B(n_1419),
.Y(n_1578)
);

INVx2_ASAP7_75t_L g1579 ( 
.A(n_1473),
.Y(n_1579)
);

INVx1_ASAP7_75t_L g1580 ( 
.A(n_1395),
.Y(n_1580)
);

AND2x2_ASAP7_75t_L g1581 ( 
.A(n_1428),
.B(n_1433),
.Y(n_1581)
);

NAND2xp5_ASAP7_75t_L g1582 ( 
.A(n_1428),
.B(n_1443),
.Y(n_1582)
);

INVx1_ASAP7_75t_L g1583 ( 
.A(n_1395),
.Y(n_1583)
);

AND2x2_ASAP7_75t_L g1584 ( 
.A(n_1462),
.B(n_1425),
.Y(n_1584)
);

INVx1_ASAP7_75t_L g1585 ( 
.A(n_1395),
.Y(n_1585)
);

AOI22xp33_ASAP7_75t_L g1586 ( 
.A1(n_1411),
.A2(n_1404),
.B1(n_1415),
.B2(n_1397),
.Y(n_1586)
);

INVx1_ASAP7_75t_L g1587 ( 
.A(n_1399),
.Y(n_1587)
);

INVx1_ASAP7_75t_L g1588 ( 
.A(n_1399),
.Y(n_1588)
);

AND2x2_ASAP7_75t_L g1589 ( 
.A(n_1425),
.B(n_1438),
.Y(n_1589)
);

INVx1_ASAP7_75t_L g1590 ( 
.A(n_1399),
.Y(n_1590)
);

NAND2xp5_ASAP7_75t_L g1591 ( 
.A(n_1388),
.B(n_1436),
.Y(n_1591)
);

CKINVDCx6p67_ASAP7_75t_R g1592 ( 
.A(n_1423),
.Y(n_1592)
);

INVx1_ASAP7_75t_L g1593 ( 
.A(n_1406),
.Y(n_1593)
);

OAI22xp5_ASAP7_75t_L g1594 ( 
.A1(n_1379),
.A2(n_1440),
.B1(n_1389),
.B2(n_1406),
.Y(n_1594)
);

INVx1_ASAP7_75t_L g1595 ( 
.A(n_1406),
.Y(n_1595)
);

INVx1_ASAP7_75t_L g1596 ( 
.A(n_1403),
.Y(n_1596)
);

INVx1_ASAP7_75t_L g1597 ( 
.A(n_1403),
.Y(n_1597)
);

INVx1_ASAP7_75t_L g1598 ( 
.A(n_1384),
.Y(n_1598)
);

INVx1_ASAP7_75t_L g1599 ( 
.A(n_1410),
.Y(n_1599)
);

OAI221xp5_ASAP7_75t_L g1600 ( 
.A1(n_1379),
.A2(n_1378),
.B1(n_1472),
.B2(n_1418),
.C(n_1412),
.Y(n_1600)
);

HB1xp67_ASAP7_75t_SL g1601 ( 
.A(n_1449),
.Y(n_1601)
);

OR2x6_ASAP7_75t_L g1602 ( 
.A(n_1556),
.B(n_1379),
.Y(n_1602)
);

AO21x2_ASAP7_75t_L g1603 ( 
.A1(n_1516),
.A2(n_1465),
.B(n_1458),
.Y(n_1603)
);

O2A1O1Ixp33_ASAP7_75t_SL g1604 ( 
.A1(n_1543),
.A2(n_1377),
.B(n_1505),
.C(n_1449),
.Y(n_1604)
);

A2O1A1Ixp33_ASAP7_75t_L g1605 ( 
.A1(n_1531),
.A2(n_1410),
.B(n_1437),
.C(n_1467),
.Y(n_1605)
);

OAI22xp5_ASAP7_75t_L g1606 ( 
.A1(n_1563),
.A2(n_1440),
.B1(n_1418),
.B2(n_1412),
.Y(n_1606)
);

INVx2_ASAP7_75t_L g1607 ( 
.A(n_1525),
.Y(n_1607)
);

OAI21xp5_ASAP7_75t_L g1608 ( 
.A1(n_1515),
.A2(n_1434),
.B(n_1418),
.Y(n_1608)
);

O2A1O1Ixp5_ASAP7_75t_L g1609 ( 
.A1(n_1517),
.A2(n_1434),
.B(n_1412),
.C(n_1456),
.Y(n_1609)
);

OR2x2_ASAP7_75t_L g1610 ( 
.A(n_1510),
.B(n_1437),
.Y(n_1610)
);

AOI22xp5_ASAP7_75t_SL g1611 ( 
.A1(n_1532),
.A2(n_1437),
.B1(n_1456),
.B2(n_1460),
.Y(n_1611)
);

OAI21xp5_ASAP7_75t_L g1612 ( 
.A1(n_1532),
.A2(n_1471),
.B(n_1456),
.Y(n_1612)
);

A2O1A1Ixp33_ASAP7_75t_L g1613 ( 
.A1(n_1555),
.A2(n_1511),
.B(n_1508),
.C(n_1561),
.Y(n_1613)
);

NAND2xp5_ASAP7_75t_L g1614 ( 
.A(n_1564),
.B(n_1460),
.Y(n_1614)
);

OA21x2_ASAP7_75t_L g1615 ( 
.A1(n_1535),
.A2(n_1516),
.B(n_1533),
.Y(n_1615)
);

NOR2xp33_ASAP7_75t_L g1616 ( 
.A(n_1549),
.B(n_1564),
.Y(n_1616)
);

INVx2_ASAP7_75t_L g1617 ( 
.A(n_1527),
.Y(n_1617)
);

AND2x2_ASAP7_75t_L g1618 ( 
.A(n_1581),
.B(n_1471),
.Y(n_1618)
);

OAI21xp5_ASAP7_75t_L g1619 ( 
.A1(n_1517),
.A2(n_1511),
.B(n_1508),
.Y(n_1619)
);

OR2x2_ASAP7_75t_L g1620 ( 
.A(n_1510),
.B(n_1534),
.Y(n_1620)
);

OR2x2_ASAP7_75t_L g1621 ( 
.A(n_1534),
.B(n_1577),
.Y(n_1621)
);

AOI221xp5_ASAP7_75t_L g1622 ( 
.A1(n_1555),
.A2(n_1561),
.B1(n_1557),
.B2(n_1568),
.C(n_1572),
.Y(n_1622)
);

AND2x4_ASAP7_75t_L g1623 ( 
.A(n_1519),
.B(n_1542),
.Y(n_1623)
);

NOR3xp33_ASAP7_75t_SL g1624 ( 
.A(n_1600),
.B(n_1594),
.C(n_1547),
.Y(n_1624)
);

OAI22xp5_ASAP7_75t_L g1625 ( 
.A1(n_1556),
.A2(n_1601),
.B1(n_1561),
.B2(n_1541),
.Y(n_1625)
);

NOR2x1_ASAP7_75t_SL g1626 ( 
.A(n_1556),
.B(n_1578),
.Y(n_1626)
);

O2A1O1Ixp33_ASAP7_75t_L g1627 ( 
.A1(n_1572),
.A2(n_1579),
.B(n_1571),
.C(n_1561),
.Y(n_1627)
);

BUFx2_ASAP7_75t_L g1628 ( 
.A(n_1514),
.Y(n_1628)
);

OR2x2_ASAP7_75t_L g1629 ( 
.A(n_1539),
.B(n_1540),
.Y(n_1629)
);

AND2x2_ASAP7_75t_L g1630 ( 
.A(n_1584),
.B(n_1578),
.Y(n_1630)
);

NAND2x1p5_ASAP7_75t_L g1631 ( 
.A(n_1579),
.B(n_1557),
.Y(n_1631)
);

OAI21x1_ASAP7_75t_SL g1632 ( 
.A1(n_1518),
.A2(n_1540),
.B(n_1550),
.Y(n_1632)
);

BUFx3_ASAP7_75t_L g1633 ( 
.A(n_1514),
.Y(n_1633)
);

BUFx6f_ASAP7_75t_L g1634 ( 
.A(n_1523),
.Y(n_1634)
);

AOI221xp5_ASAP7_75t_L g1635 ( 
.A1(n_1552),
.A2(n_1575),
.B1(n_1570),
.B2(n_1512),
.C(n_1524),
.Y(n_1635)
);

OAI21xp5_ASAP7_75t_L g1636 ( 
.A1(n_1518),
.A2(n_1509),
.B(n_1533),
.Y(n_1636)
);

OAI211xp5_ASAP7_75t_SL g1637 ( 
.A1(n_1586),
.A2(n_1598),
.B(n_1591),
.C(n_1582),
.Y(n_1637)
);

NOR2x1_ASAP7_75t_SL g1638 ( 
.A(n_1556),
.B(n_1578),
.Y(n_1638)
);

OAI21x1_ASAP7_75t_SL g1639 ( 
.A1(n_1546),
.A2(n_1550),
.B(n_1565),
.Y(n_1639)
);

NOR2xp33_ASAP7_75t_L g1640 ( 
.A(n_1556),
.B(n_1537),
.Y(n_1640)
);

OR2x2_ASAP7_75t_L g1641 ( 
.A(n_1546),
.B(n_1512),
.Y(n_1641)
);

OR2x2_ASAP7_75t_L g1642 ( 
.A(n_1524),
.B(n_1537),
.Y(n_1642)
);

NAND2xp5_ASAP7_75t_L g1643 ( 
.A(n_1567),
.B(n_1558),
.Y(n_1643)
);

OAI22xp5_ASAP7_75t_L g1644 ( 
.A1(n_1541),
.A2(n_1598),
.B1(n_1530),
.B2(n_1521),
.Y(n_1644)
);

NAND2xp5_ASAP7_75t_L g1645 ( 
.A(n_1567),
.B(n_1558),
.Y(n_1645)
);

OR2x2_ASAP7_75t_L g1646 ( 
.A(n_1573),
.B(n_1559),
.Y(n_1646)
);

AND2x2_ASAP7_75t_L g1647 ( 
.A(n_1573),
.B(n_1589),
.Y(n_1647)
);

CKINVDCx5p33_ASAP7_75t_R g1648 ( 
.A(n_1592),
.Y(n_1648)
);

AND2x2_ASAP7_75t_L g1649 ( 
.A(n_1566),
.B(n_1522),
.Y(n_1649)
);

AOI21xp5_ASAP7_75t_L g1650 ( 
.A1(n_1552),
.A2(n_1545),
.B(n_1576),
.Y(n_1650)
);

NOR2x1_ASAP7_75t_SL g1651 ( 
.A(n_1576),
.B(n_1574),
.Y(n_1651)
);

AND2x2_ASAP7_75t_L g1652 ( 
.A(n_1522),
.B(n_1538),
.Y(n_1652)
);

INVx5_ASAP7_75t_SL g1653 ( 
.A(n_1592),
.Y(n_1653)
);

OR2x6_ASAP7_75t_L g1654 ( 
.A(n_1576),
.B(n_1553),
.Y(n_1654)
);

AND2x2_ASAP7_75t_L g1655 ( 
.A(n_1538),
.B(n_1599),
.Y(n_1655)
);

O2A1O1Ixp33_ASAP7_75t_L g1656 ( 
.A1(n_1521),
.A2(n_1530),
.B(n_1583),
.C(n_1593),
.Y(n_1656)
);

OAI21xp5_ASAP7_75t_L g1657 ( 
.A1(n_1596),
.A2(n_1597),
.B(n_1593),
.Y(n_1657)
);

AO32x2_ASAP7_75t_L g1658 ( 
.A1(n_1554),
.A2(n_1538),
.A3(n_1570),
.B1(n_1575),
.B2(n_1574),
.Y(n_1658)
);

AND2x2_ASAP7_75t_L g1659 ( 
.A(n_1538),
.B(n_1599),
.Y(n_1659)
);

A2O1A1Ixp33_ASAP7_75t_L g1660 ( 
.A1(n_1538),
.A2(n_1530),
.B(n_1521),
.C(n_1554),
.Y(n_1660)
);

A2O1A1Ixp33_ASAP7_75t_L g1661 ( 
.A1(n_1538),
.A2(n_1554),
.B(n_1548),
.C(n_1545),
.Y(n_1661)
);

OR2x2_ASAP7_75t_L g1662 ( 
.A(n_1548),
.B(n_1513),
.Y(n_1662)
);

INVx1_ASAP7_75t_L g1663 ( 
.A(n_1607),
.Y(n_1663)
);

OAI22xp5_ASAP7_75t_L g1664 ( 
.A1(n_1605),
.A2(n_1576),
.B1(n_1523),
.B2(n_1590),
.Y(n_1664)
);

OR2x2_ASAP7_75t_L g1665 ( 
.A(n_1620),
.B(n_1554),
.Y(n_1665)
);

AND2x2_ASAP7_75t_L g1666 ( 
.A(n_1647),
.B(n_1630),
.Y(n_1666)
);

INVx1_ASAP7_75t_L g1667 ( 
.A(n_1617),
.Y(n_1667)
);

BUFx12f_ASAP7_75t_L g1668 ( 
.A(n_1648),
.Y(n_1668)
);

INVx1_ASAP7_75t_L g1669 ( 
.A(n_1617),
.Y(n_1669)
);

AND2x2_ASAP7_75t_L g1670 ( 
.A(n_1655),
.B(n_1554),
.Y(n_1670)
);

AND2x4_ASAP7_75t_L g1671 ( 
.A(n_1654),
.B(n_1551),
.Y(n_1671)
);

NOR2x1_ASAP7_75t_L g1672 ( 
.A(n_1633),
.B(n_1576),
.Y(n_1672)
);

NAND2xp5_ASAP7_75t_L g1673 ( 
.A(n_1619),
.B(n_1569),
.Y(n_1673)
);

OR2x2_ASAP7_75t_L g1674 ( 
.A(n_1646),
.B(n_1652),
.Y(n_1674)
);

OAI22xp5_ASAP7_75t_L g1675 ( 
.A1(n_1605),
.A2(n_1588),
.B1(n_1580),
.B2(n_1583),
.Y(n_1675)
);

AND2x2_ASAP7_75t_L g1676 ( 
.A(n_1659),
.B(n_1554),
.Y(n_1676)
);

AND2x2_ASAP7_75t_L g1677 ( 
.A(n_1658),
.B(n_1574),
.Y(n_1677)
);

AOI22xp33_ASAP7_75t_L g1678 ( 
.A1(n_1616),
.A2(n_1580),
.B1(n_1585),
.B2(n_1595),
.Y(n_1678)
);

OR2x2_ASAP7_75t_L g1679 ( 
.A(n_1641),
.B(n_1526),
.Y(n_1679)
);

BUFx2_ASAP7_75t_L g1680 ( 
.A(n_1631),
.Y(n_1680)
);

OR2x2_ASAP7_75t_L g1681 ( 
.A(n_1642),
.B(n_1526),
.Y(n_1681)
);

INVxp67_ASAP7_75t_SL g1682 ( 
.A(n_1614),
.Y(n_1682)
);

BUFx2_ASAP7_75t_L g1683 ( 
.A(n_1631),
.Y(n_1683)
);

AND2x2_ASAP7_75t_L g1684 ( 
.A(n_1658),
.B(n_1560),
.Y(n_1684)
);

INVx1_ASAP7_75t_L g1685 ( 
.A(n_1629),
.Y(n_1685)
);

OR2x2_ASAP7_75t_SL g1686 ( 
.A(n_1615),
.B(n_1588),
.Y(n_1686)
);

INVx1_ASAP7_75t_L g1687 ( 
.A(n_1621),
.Y(n_1687)
);

INVx1_ASAP7_75t_L g1688 ( 
.A(n_1662),
.Y(n_1688)
);

INVx1_ASAP7_75t_L g1689 ( 
.A(n_1643),
.Y(n_1689)
);

INVx2_ASAP7_75t_L g1690 ( 
.A(n_1649),
.Y(n_1690)
);

AND2x4_ASAP7_75t_SL g1691 ( 
.A(n_1602),
.B(n_1536),
.Y(n_1691)
);

AOI22xp33_ASAP7_75t_L g1692 ( 
.A1(n_1616),
.A2(n_1585),
.B1(n_1587),
.B2(n_1595),
.Y(n_1692)
);

AOI22xp5_ASAP7_75t_L g1693 ( 
.A1(n_1637),
.A2(n_1606),
.B1(n_1625),
.B2(n_1602),
.Y(n_1693)
);

NOR2xp33_ASAP7_75t_L g1694 ( 
.A(n_1637),
.B(n_1648),
.Y(n_1694)
);

INVx1_ASAP7_75t_L g1695 ( 
.A(n_1639),
.Y(n_1695)
);

AND2x2_ASAP7_75t_L g1696 ( 
.A(n_1658),
.B(n_1562),
.Y(n_1696)
);

INVx1_ASAP7_75t_L g1697 ( 
.A(n_1645),
.Y(n_1697)
);

INVx1_ASAP7_75t_L g1698 ( 
.A(n_1632),
.Y(n_1698)
);

AND2x2_ASAP7_75t_L g1699 ( 
.A(n_1666),
.B(n_1615),
.Y(n_1699)
);

NAND2xp5_ASAP7_75t_L g1700 ( 
.A(n_1697),
.B(n_1635),
.Y(n_1700)
);

INVx1_ASAP7_75t_SL g1701 ( 
.A(n_1680),
.Y(n_1701)
);

OAI221xp5_ASAP7_75t_SL g1702 ( 
.A1(n_1693),
.A2(n_1613),
.B1(n_1622),
.B2(n_1627),
.C(n_1661),
.Y(n_1702)
);

INVx2_ASAP7_75t_L g1703 ( 
.A(n_1684),
.Y(n_1703)
);

AND2x2_ASAP7_75t_L g1704 ( 
.A(n_1670),
.B(n_1651),
.Y(n_1704)
);

INVx1_ASAP7_75t_SL g1705 ( 
.A(n_1680),
.Y(n_1705)
);

HB1xp67_ASAP7_75t_L g1706 ( 
.A(n_1684),
.Y(n_1706)
);

INVxp67_ASAP7_75t_L g1707 ( 
.A(n_1698),
.Y(n_1707)
);

INVx4_ASAP7_75t_L g1708 ( 
.A(n_1668),
.Y(n_1708)
);

AND2x4_ASAP7_75t_L g1709 ( 
.A(n_1671),
.B(n_1654),
.Y(n_1709)
);

AOI22xp5_ASAP7_75t_L g1710 ( 
.A1(n_1694),
.A2(n_1613),
.B1(n_1640),
.B2(n_1664),
.Y(n_1710)
);

INVx1_ASAP7_75t_L g1711 ( 
.A(n_1663),
.Y(n_1711)
);

OAI21xp33_ASAP7_75t_L g1712 ( 
.A1(n_1677),
.A2(n_1624),
.B(n_1661),
.Y(n_1712)
);

AOI221xp5_ASAP7_75t_L g1713 ( 
.A1(n_1677),
.A2(n_1604),
.B1(n_1660),
.B2(n_1650),
.C(n_1624),
.Y(n_1713)
);

NAND2xp5_ASAP7_75t_L g1714 ( 
.A(n_1697),
.B(n_1660),
.Y(n_1714)
);

NOR2xp33_ASAP7_75t_L g1715 ( 
.A(n_1668),
.B(n_1644),
.Y(n_1715)
);

OAI322xp33_ASAP7_75t_L g1716 ( 
.A1(n_1665),
.A2(n_1681),
.A3(n_1673),
.B1(n_1679),
.B2(n_1689),
.C1(n_1676),
.C2(n_1670),
.Y(n_1716)
);

INVx2_ASAP7_75t_L g1717 ( 
.A(n_1696),
.Y(n_1717)
);

OAI21xp5_ASAP7_75t_L g1718 ( 
.A1(n_1675),
.A2(n_1636),
.B(n_1609),
.Y(n_1718)
);

AND2x4_ASAP7_75t_L g1719 ( 
.A(n_1671),
.B(n_1626),
.Y(n_1719)
);

AND2x4_ASAP7_75t_L g1720 ( 
.A(n_1671),
.B(n_1638),
.Y(n_1720)
);

AND4x1_ASAP7_75t_L g1721 ( 
.A(n_1672),
.B(n_1656),
.C(n_1608),
.D(n_1609),
.Y(n_1721)
);

INVx2_ASAP7_75t_L g1722 ( 
.A(n_1663),
.Y(n_1722)
);

AOI22xp33_ASAP7_75t_L g1723 ( 
.A1(n_1682),
.A2(n_1602),
.B1(n_1653),
.B2(n_1612),
.Y(n_1723)
);

INVx1_ASAP7_75t_SL g1724 ( 
.A(n_1683),
.Y(n_1724)
);

INVx1_ASAP7_75t_L g1725 ( 
.A(n_1667),
.Y(n_1725)
);

AND2x4_ASAP7_75t_L g1726 ( 
.A(n_1691),
.B(n_1603),
.Y(n_1726)
);

HB1xp67_ASAP7_75t_L g1727 ( 
.A(n_1667),
.Y(n_1727)
);

OR2x2_ASAP7_75t_L g1728 ( 
.A(n_1686),
.B(n_1603),
.Y(n_1728)
);

BUFx2_ASAP7_75t_L g1729 ( 
.A(n_1686),
.Y(n_1729)
);

AND2x2_ASAP7_75t_L g1730 ( 
.A(n_1690),
.B(n_1623),
.Y(n_1730)
);

OAI22xp5_ASAP7_75t_L g1731 ( 
.A1(n_1665),
.A2(n_1611),
.B1(n_1653),
.B2(n_1610),
.Y(n_1731)
);

AOI221xp5_ASAP7_75t_L g1732 ( 
.A1(n_1678),
.A2(n_1604),
.B1(n_1657),
.B2(n_1520),
.C(n_1628),
.Y(n_1732)
);

INVx1_ASAP7_75t_L g1733 ( 
.A(n_1669),
.Y(n_1733)
);

BUFx2_ASAP7_75t_L g1734 ( 
.A(n_1729),
.Y(n_1734)
);

INVx2_ASAP7_75t_L g1735 ( 
.A(n_1703),
.Y(n_1735)
);

XNOR2xp5_ASAP7_75t_L g1736 ( 
.A(n_1710),
.B(n_1618),
.Y(n_1736)
);

INVx1_ASAP7_75t_L g1737 ( 
.A(n_1711),
.Y(n_1737)
);

BUFx2_ASAP7_75t_L g1738 ( 
.A(n_1729),
.Y(n_1738)
);

OR2x2_ASAP7_75t_L g1739 ( 
.A(n_1706),
.B(n_1674),
.Y(n_1739)
);

INVx1_ASAP7_75t_L g1740 ( 
.A(n_1711),
.Y(n_1740)
);

INVx2_ASAP7_75t_L g1741 ( 
.A(n_1703),
.Y(n_1741)
);

INVx2_ASAP7_75t_L g1742 ( 
.A(n_1703),
.Y(n_1742)
);

NAND2xp5_ASAP7_75t_L g1743 ( 
.A(n_1700),
.B(n_1688),
.Y(n_1743)
);

NAND2xp5_ASAP7_75t_L g1744 ( 
.A(n_1700),
.B(n_1688),
.Y(n_1744)
);

OR2x2_ASAP7_75t_L g1745 ( 
.A(n_1706),
.B(n_1674),
.Y(n_1745)
);

NAND2xp5_ASAP7_75t_L g1746 ( 
.A(n_1714),
.B(n_1685),
.Y(n_1746)
);

NAND2xp5_ASAP7_75t_L g1747 ( 
.A(n_1714),
.B(n_1685),
.Y(n_1747)
);

INVx1_ASAP7_75t_L g1748 ( 
.A(n_1725),
.Y(n_1748)
);

NAND2xp5_ASAP7_75t_L g1749 ( 
.A(n_1707),
.B(n_1687),
.Y(n_1749)
);

AOI22xp33_ASAP7_75t_L g1750 ( 
.A1(n_1712),
.A2(n_1692),
.B1(n_1653),
.B2(n_1695),
.Y(n_1750)
);

NOR2x1_ASAP7_75t_L g1751 ( 
.A(n_1708),
.B(n_1695),
.Y(n_1751)
);

INVx2_ASAP7_75t_L g1752 ( 
.A(n_1717),
.Y(n_1752)
);

AND2x4_ASAP7_75t_L g1753 ( 
.A(n_1719),
.B(n_1720),
.Y(n_1753)
);

INVx1_ASAP7_75t_SL g1754 ( 
.A(n_1701),
.Y(n_1754)
);

INVx1_ASAP7_75t_L g1755 ( 
.A(n_1725),
.Y(n_1755)
);

INVx1_ASAP7_75t_L g1756 ( 
.A(n_1733),
.Y(n_1756)
);

INVx5_ASAP7_75t_L g1757 ( 
.A(n_1708),
.Y(n_1757)
);

INVx1_ASAP7_75t_L g1758 ( 
.A(n_1733),
.Y(n_1758)
);

AND2x4_ASAP7_75t_L g1759 ( 
.A(n_1719),
.B(n_1683),
.Y(n_1759)
);

INVx1_ASAP7_75t_L g1760 ( 
.A(n_1727),
.Y(n_1760)
);

INVx2_ASAP7_75t_L g1761 ( 
.A(n_1717),
.Y(n_1761)
);

INVx1_ASAP7_75t_L g1762 ( 
.A(n_1727),
.Y(n_1762)
);

OR2x2_ASAP7_75t_L g1763 ( 
.A(n_1728),
.B(n_1681),
.Y(n_1763)
);

INVx1_ASAP7_75t_L g1764 ( 
.A(n_1722),
.Y(n_1764)
);

BUFx2_ASAP7_75t_L g1765 ( 
.A(n_1719),
.Y(n_1765)
);

NAND2xp5_ASAP7_75t_L g1766 ( 
.A(n_1743),
.B(n_1710),
.Y(n_1766)
);

INVx1_ASAP7_75t_L g1767 ( 
.A(n_1737),
.Y(n_1767)
);

OR2x2_ASAP7_75t_L g1768 ( 
.A(n_1763),
.B(n_1728),
.Y(n_1768)
);

NAND2xp5_ASAP7_75t_L g1769 ( 
.A(n_1743),
.B(n_1712),
.Y(n_1769)
);

NAND2xp5_ASAP7_75t_L g1770 ( 
.A(n_1744),
.B(n_1730),
.Y(n_1770)
);

INVx2_ASAP7_75t_L g1771 ( 
.A(n_1735),
.Y(n_1771)
);

INVx2_ASAP7_75t_L g1772 ( 
.A(n_1735),
.Y(n_1772)
);

INVx1_ASAP7_75t_L g1773 ( 
.A(n_1737),
.Y(n_1773)
);

OR2x2_ASAP7_75t_L g1774 ( 
.A(n_1763),
.B(n_1728),
.Y(n_1774)
);

INVx1_ASAP7_75t_L g1775 ( 
.A(n_1740),
.Y(n_1775)
);

INVx1_ASAP7_75t_L g1776 ( 
.A(n_1740),
.Y(n_1776)
);

AND2x4_ASAP7_75t_L g1777 ( 
.A(n_1757),
.B(n_1719),
.Y(n_1777)
);

INVx1_ASAP7_75t_L g1778 ( 
.A(n_1748),
.Y(n_1778)
);

NAND2xp5_ASAP7_75t_L g1779 ( 
.A(n_1744),
.B(n_1730),
.Y(n_1779)
);

NAND2xp33_ASAP7_75t_R g1780 ( 
.A(n_1734),
.B(n_1544),
.Y(n_1780)
);

INVx1_ASAP7_75t_L g1781 ( 
.A(n_1748),
.Y(n_1781)
);

OR2x2_ASAP7_75t_L g1782 ( 
.A(n_1763),
.B(n_1699),
.Y(n_1782)
);

NAND2xp5_ASAP7_75t_L g1783 ( 
.A(n_1736),
.B(n_1730),
.Y(n_1783)
);

OR2x2_ASAP7_75t_L g1784 ( 
.A(n_1746),
.B(n_1699),
.Y(n_1784)
);

INVx1_ASAP7_75t_L g1785 ( 
.A(n_1755),
.Y(n_1785)
);

NOR2x1_ASAP7_75t_L g1786 ( 
.A(n_1751),
.B(n_1708),
.Y(n_1786)
);

INVx2_ASAP7_75t_L g1787 ( 
.A(n_1735),
.Y(n_1787)
);

HB1xp67_ASAP7_75t_L g1788 ( 
.A(n_1734),
.Y(n_1788)
);

INVx1_ASAP7_75t_L g1789 ( 
.A(n_1755),
.Y(n_1789)
);

NAND2xp5_ASAP7_75t_L g1790 ( 
.A(n_1736),
.B(n_1707),
.Y(n_1790)
);

HB1xp67_ASAP7_75t_L g1791 ( 
.A(n_1734),
.Y(n_1791)
);

NAND2xp5_ASAP7_75t_L g1792 ( 
.A(n_1736),
.B(n_1701),
.Y(n_1792)
);

AOI21xp5_ASAP7_75t_L g1793 ( 
.A1(n_1750),
.A2(n_1702),
.B(n_1718),
.Y(n_1793)
);

AND2x4_ASAP7_75t_L g1794 ( 
.A(n_1757),
.B(n_1719),
.Y(n_1794)
);

NAND2xp5_ASAP7_75t_L g1795 ( 
.A(n_1746),
.B(n_1705),
.Y(n_1795)
);

INVx1_ASAP7_75t_L g1796 ( 
.A(n_1756),
.Y(n_1796)
);

INVx1_ASAP7_75t_L g1797 ( 
.A(n_1756),
.Y(n_1797)
);

AND2x2_ASAP7_75t_L g1798 ( 
.A(n_1765),
.B(n_1704),
.Y(n_1798)
);

INVx1_ASAP7_75t_L g1799 ( 
.A(n_1758),
.Y(n_1799)
);

INVx1_ASAP7_75t_L g1800 ( 
.A(n_1758),
.Y(n_1800)
);

AND2x2_ASAP7_75t_L g1801 ( 
.A(n_1765),
.B(n_1704),
.Y(n_1801)
);

AND2x2_ASAP7_75t_L g1802 ( 
.A(n_1765),
.B(n_1704),
.Y(n_1802)
);

NAND2xp5_ASAP7_75t_L g1803 ( 
.A(n_1747),
.B(n_1705),
.Y(n_1803)
);

NAND3xp33_ASAP7_75t_L g1804 ( 
.A(n_1750),
.B(n_1702),
.C(n_1713),
.Y(n_1804)
);

INVx1_ASAP7_75t_L g1805 ( 
.A(n_1760),
.Y(n_1805)
);

INVx2_ASAP7_75t_L g1806 ( 
.A(n_1735),
.Y(n_1806)
);

INVx1_ASAP7_75t_L g1807 ( 
.A(n_1760),
.Y(n_1807)
);

INVx1_ASAP7_75t_L g1808 ( 
.A(n_1749),
.Y(n_1808)
);

INVx1_ASAP7_75t_L g1809 ( 
.A(n_1773),
.Y(n_1809)
);

INVx1_ASAP7_75t_L g1810 ( 
.A(n_1773),
.Y(n_1810)
);

INVx2_ASAP7_75t_L g1811 ( 
.A(n_1788),
.Y(n_1811)
);

NAND2xp5_ASAP7_75t_L g1812 ( 
.A(n_1769),
.B(n_1747),
.Y(n_1812)
);

INVx1_ASAP7_75t_SL g1813 ( 
.A(n_1791),
.Y(n_1813)
);

AND2x2_ASAP7_75t_L g1814 ( 
.A(n_1798),
.B(n_1801),
.Y(n_1814)
);

AND2x2_ASAP7_75t_L g1815 ( 
.A(n_1798),
.B(n_1738),
.Y(n_1815)
);

NAND4xp25_ASAP7_75t_L g1816 ( 
.A(n_1804),
.B(n_1713),
.C(n_1732),
.D(n_1718),
.Y(n_1816)
);

BUFx2_ASAP7_75t_L g1817 ( 
.A(n_1786),
.Y(n_1817)
);

AOI22xp33_ASAP7_75t_SL g1818 ( 
.A1(n_1793),
.A2(n_1738),
.B1(n_1757),
.B2(n_1708),
.Y(n_1818)
);

NAND2xp5_ASAP7_75t_L g1819 ( 
.A(n_1766),
.B(n_1738),
.Y(n_1819)
);

OR2x2_ASAP7_75t_L g1820 ( 
.A(n_1770),
.B(n_1779),
.Y(n_1820)
);

INVxp33_ASAP7_75t_L g1821 ( 
.A(n_1792),
.Y(n_1821)
);

INVx1_ASAP7_75t_L g1822 ( 
.A(n_1775),
.Y(n_1822)
);

NOR2xp33_ASAP7_75t_L g1823 ( 
.A(n_1790),
.B(n_1708),
.Y(n_1823)
);

AND2x2_ASAP7_75t_L g1824 ( 
.A(n_1801),
.B(n_1753),
.Y(n_1824)
);

OAI31xp33_ASAP7_75t_L g1825 ( 
.A1(n_1783),
.A2(n_1715),
.A3(n_1754),
.B(n_1731),
.Y(n_1825)
);

AND2x2_ASAP7_75t_L g1826 ( 
.A(n_1802),
.B(n_1753),
.Y(n_1826)
);

NAND2xp5_ASAP7_75t_L g1827 ( 
.A(n_1808),
.B(n_1762),
.Y(n_1827)
);

AND2x2_ASAP7_75t_L g1828 ( 
.A(n_1802),
.B(n_1753),
.Y(n_1828)
);

NAND2xp5_ASAP7_75t_L g1829 ( 
.A(n_1795),
.B(n_1754),
.Y(n_1829)
);

NAND2xp33_ASAP7_75t_SL g1830 ( 
.A(n_1780),
.B(n_1731),
.Y(n_1830)
);

OR2x2_ASAP7_75t_L g1831 ( 
.A(n_1803),
.B(n_1784),
.Y(n_1831)
);

OR2x2_ASAP7_75t_L g1832 ( 
.A(n_1784),
.B(n_1749),
.Y(n_1832)
);

AND2x2_ASAP7_75t_L g1833 ( 
.A(n_1777),
.B(n_1753),
.Y(n_1833)
);

INVx1_ASAP7_75t_L g1834 ( 
.A(n_1775),
.Y(n_1834)
);

AND2x2_ASAP7_75t_L g1835 ( 
.A(n_1777),
.B(n_1794),
.Y(n_1835)
);

INVx1_ASAP7_75t_L g1836 ( 
.A(n_1776),
.Y(n_1836)
);

AND2x2_ASAP7_75t_L g1837 ( 
.A(n_1777),
.B(n_1753),
.Y(n_1837)
);

AOI22xp5_ASAP7_75t_L g1838 ( 
.A1(n_1794),
.A2(n_1732),
.B1(n_1757),
.B2(n_1723),
.Y(n_1838)
);

NOR2x1_ASAP7_75t_L g1839 ( 
.A(n_1805),
.B(n_1751),
.Y(n_1839)
);

NAND2xp5_ASAP7_75t_L g1840 ( 
.A(n_1805),
.B(n_1762),
.Y(n_1840)
);

INVx2_ASAP7_75t_L g1841 ( 
.A(n_1771),
.Y(n_1841)
);

INVx1_ASAP7_75t_L g1842 ( 
.A(n_1776),
.Y(n_1842)
);

AND2x2_ASAP7_75t_L g1843 ( 
.A(n_1794),
.B(n_1759),
.Y(n_1843)
);

INVx2_ASAP7_75t_L g1844 ( 
.A(n_1771),
.Y(n_1844)
);

INVx1_ASAP7_75t_L g1845 ( 
.A(n_1809),
.Y(n_1845)
);

OAI322xp33_ASAP7_75t_L g1846 ( 
.A1(n_1819),
.A2(n_1774),
.A3(n_1768),
.B1(n_1807),
.B2(n_1782),
.C1(n_1778),
.C2(n_1799),
.Y(n_1846)
);

INVxp67_ASAP7_75t_L g1847 ( 
.A(n_1817),
.Y(n_1847)
);

OR2x2_ASAP7_75t_L g1848 ( 
.A(n_1813),
.B(n_1807),
.Y(n_1848)
);

NOR2xp33_ASAP7_75t_L g1849 ( 
.A(n_1816),
.B(n_1757),
.Y(n_1849)
);

OAI222xp33_ASAP7_75t_L g1850 ( 
.A1(n_1838),
.A2(n_1757),
.B1(n_1774),
.B2(n_1768),
.C1(n_1723),
.C2(n_1782),
.Y(n_1850)
);

INVx1_ASAP7_75t_L g1851 ( 
.A(n_1809),
.Y(n_1851)
);

INVx1_ASAP7_75t_L g1852 ( 
.A(n_1810),
.Y(n_1852)
);

INVx1_ASAP7_75t_L g1853 ( 
.A(n_1810),
.Y(n_1853)
);

NAND2xp5_ASAP7_75t_L g1854 ( 
.A(n_1821),
.B(n_1767),
.Y(n_1854)
);

INVx1_ASAP7_75t_L g1855 ( 
.A(n_1822),
.Y(n_1855)
);

INVx1_ASAP7_75t_L g1856 ( 
.A(n_1822),
.Y(n_1856)
);

NAND2xp5_ASAP7_75t_L g1857 ( 
.A(n_1819),
.B(n_1781),
.Y(n_1857)
);

OAI22xp5_ASAP7_75t_L g1858 ( 
.A1(n_1838),
.A2(n_1757),
.B1(n_1745),
.B2(n_1739),
.Y(n_1858)
);

OAI21xp33_ASAP7_75t_L g1859 ( 
.A1(n_1816),
.A2(n_1721),
.B(n_1785),
.Y(n_1859)
);

AND2x2_ASAP7_75t_L g1860 ( 
.A(n_1814),
.B(n_1757),
.Y(n_1860)
);

OAI33xp33_ASAP7_75t_L g1861 ( 
.A1(n_1827),
.A2(n_1800),
.A3(n_1799),
.B1(n_1778),
.B2(n_1797),
.B3(n_1796),
.Y(n_1861)
);

OAI211xp5_ASAP7_75t_L g1862 ( 
.A1(n_1818),
.A2(n_1757),
.B(n_1800),
.C(n_1789),
.Y(n_1862)
);

INVx2_ASAP7_75t_L g1863 ( 
.A(n_1815),
.Y(n_1863)
);

INVx2_ASAP7_75t_L g1864 ( 
.A(n_1815),
.Y(n_1864)
);

INVxp67_ASAP7_75t_SL g1865 ( 
.A(n_1839),
.Y(n_1865)
);

OR2x2_ASAP7_75t_L g1866 ( 
.A(n_1829),
.B(n_1739),
.Y(n_1866)
);

O2A1O1Ixp33_ASAP7_75t_L g1867 ( 
.A1(n_1825),
.A2(n_1716),
.B(n_1787),
.C(n_1772),
.Y(n_1867)
);

AOI22xp5_ASAP7_75t_L g1868 ( 
.A1(n_1830),
.A2(n_1720),
.B1(n_1759),
.B2(n_1726),
.Y(n_1868)
);

AOI22xp5_ASAP7_75t_L g1869 ( 
.A1(n_1823),
.A2(n_1720),
.B1(n_1759),
.B2(n_1726),
.Y(n_1869)
);

INVx1_ASAP7_75t_L g1870 ( 
.A(n_1834),
.Y(n_1870)
);

XNOR2xp5_ASAP7_75t_L g1871 ( 
.A(n_1835),
.B(n_1721),
.Y(n_1871)
);

NOR2xp33_ASAP7_75t_L g1872 ( 
.A(n_1859),
.B(n_1812),
.Y(n_1872)
);

NAND2xp5_ASAP7_75t_L g1873 ( 
.A(n_1849),
.B(n_1813),
.Y(n_1873)
);

INVx1_ASAP7_75t_L g1874 ( 
.A(n_1848),
.Y(n_1874)
);

INVx1_ASAP7_75t_L g1875 ( 
.A(n_1848),
.Y(n_1875)
);

INVx1_ASAP7_75t_L g1876 ( 
.A(n_1863),
.Y(n_1876)
);

OAI22xp33_ASAP7_75t_SL g1877 ( 
.A1(n_1865),
.A2(n_1817),
.B1(n_1839),
.B2(n_1811),
.Y(n_1877)
);

AND2x4_ASAP7_75t_L g1878 ( 
.A(n_1863),
.B(n_1811),
.Y(n_1878)
);

OAI32xp33_ASAP7_75t_L g1879 ( 
.A1(n_1849),
.A2(n_1858),
.A3(n_1864),
.B1(n_1847),
.B2(n_1812),
.Y(n_1879)
);

NOR2xp67_ASAP7_75t_L g1880 ( 
.A(n_1862),
.B(n_1811),
.Y(n_1880)
);

NAND2xp5_ASAP7_75t_L g1881 ( 
.A(n_1864),
.B(n_1814),
.Y(n_1881)
);

AOI321xp33_ASAP7_75t_L g1882 ( 
.A1(n_1865),
.A2(n_1835),
.A3(n_1825),
.B1(n_1843),
.B2(n_1831),
.C(n_1833),
.Y(n_1882)
);

OAI22xp5_ASAP7_75t_L g1883 ( 
.A1(n_1871),
.A2(n_1831),
.B1(n_1832),
.B2(n_1840),
.Y(n_1883)
);

INVx1_ASAP7_75t_L g1884 ( 
.A(n_1845),
.Y(n_1884)
);

NAND2xp5_ASAP7_75t_SL g1885 ( 
.A(n_1868),
.B(n_1843),
.Y(n_1885)
);

AOI221xp5_ASAP7_75t_SL g1886 ( 
.A1(n_1846),
.A2(n_1840),
.B1(n_1827),
.B2(n_1834),
.C(n_1842),
.Y(n_1886)
);

AOI22xp5_ASAP7_75t_L g1887 ( 
.A1(n_1860),
.A2(n_1833),
.B1(n_1837),
.B2(n_1828),
.Y(n_1887)
);

OAI31xp33_ASAP7_75t_L g1888 ( 
.A1(n_1850),
.A2(n_1837),
.A3(n_1826),
.B(n_1824),
.Y(n_1888)
);

INVx1_ASAP7_75t_L g1889 ( 
.A(n_1851),
.Y(n_1889)
);

AND2x4_ASAP7_75t_L g1890 ( 
.A(n_1860),
.B(n_1824),
.Y(n_1890)
);

INVx2_ASAP7_75t_L g1891 ( 
.A(n_1852),
.Y(n_1891)
);

INVxp67_ASAP7_75t_L g1892 ( 
.A(n_1854),
.Y(n_1892)
);

NOR2xp33_ASAP7_75t_L g1893 ( 
.A(n_1892),
.B(n_1866),
.Y(n_1893)
);

NAND2xp5_ASAP7_75t_L g1894 ( 
.A(n_1874),
.B(n_1853),
.Y(n_1894)
);

INVx1_ASAP7_75t_L g1895 ( 
.A(n_1878),
.Y(n_1895)
);

INVx1_ASAP7_75t_L g1896 ( 
.A(n_1878),
.Y(n_1896)
);

NAND2xp5_ASAP7_75t_L g1897 ( 
.A(n_1875),
.B(n_1855),
.Y(n_1897)
);

INVx1_ASAP7_75t_L g1898 ( 
.A(n_1876),
.Y(n_1898)
);

A2O1A1Ixp33_ASAP7_75t_L g1899 ( 
.A1(n_1882),
.A2(n_1867),
.B(n_1857),
.C(n_1869),
.Y(n_1899)
);

INVx1_ASAP7_75t_L g1900 ( 
.A(n_1881),
.Y(n_1900)
);

NAND2xp5_ASAP7_75t_L g1901 ( 
.A(n_1872),
.B(n_1856),
.Y(n_1901)
);

NAND2xp5_ASAP7_75t_L g1902 ( 
.A(n_1883),
.B(n_1870),
.Y(n_1902)
);

OR2x2_ASAP7_75t_L g1903 ( 
.A(n_1883),
.B(n_1820),
.Y(n_1903)
);

AOI22xp33_ASAP7_75t_L g1904 ( 
.A1(n_1888),
.A2(n_1861),
.B1(n_1820),
.B2(n_1828),
.Y(n_1904)
);

INVx2_ASAP7_75t_L g1905 ( 
.A(n_1890),
.Y(n_1905)
);

XNOR2x1_ASAP7_75t_L g1906 ( 
.A(n_1873),
.B(n_1826),
.Y(n_1906)
);

OR2x2_ASAP7_75t_L g1907 ( 
.A(n_1903),
.B(n_1891),
.Y(n_1907)
);

OR2x2_ASAP7_75t_L g1908 ( 
.A(n_1895),
.B(n_1885),
.Y(n_1908)
);

NAND3xp33_ASAP7_75t_SL g1909 ( 
.A(n_1899),
.B(n_1887),
.C(n_1877),
.Y(n_1909)
);

O2A1O1Ixp33_ASAP7_75t_L g1910 ( 
.A1(n_1902),
.A2(n_1879),
.B(n_1880),
.C(n_1884),
.Y(n_1910)
);

AOI21xp5_ASAP7_75t_L g1911 ( 
.A1(n_1901),
.A2(n_1889),
.B(n_1890),
.Y(n_1911)
);

AOI221xp5_ASAP7_75t_L g1912 ( 
.A1(n_1904),
.A2(n_1886),
.B1(n_1893),
.B2(n_1896),
.C(n_1905),
.Y(n_1912)
);

NAND3xp33_ASAP7_75t_L g1913 ( 
.A(n_1900),
.B(n_1886),
.C(n_1842),
.Y(n_1913)
);

NAND2xp5_ASAP7_75t_SL g1914 ( 
.A(n_1894),
.B(n_1832),
.Y(n_1914)
);

AOI21xp5_ASAP7_75t_L g1915 ( 
.A1(n_1906),
.A2(n_1836),
.B(n_1844),
.Y(n_1915)
);

NOR3xp33_ASAP7_75t_L g1916 ( 
.A(n_1894),
.B(n_1836),
.C(n_1844),
.Y(n_1916)
);

NAND2xp5_ASAP7_75t_SL g1917 ( 
.A(n_1897),
.B(n_1898),
.Y(n_1917)
);

OR2x2_ASAP7_75t_L g1918 ( 
.A(n_1907),
.B(n_1897),
.Y(n_1918)
);

AOI22xp33_ASAP7_75t_SL g1919 ( 
.A1(n_1913),
.A2(n_1520),
.B1(n_1529),
.B2(n_1841),
.Y(n_1919)
);

AOI211xp5_ASAP7_75t_L g1920 ( 
.A1(n_1909),
.A2(n_1844),
.B(n_1841),
.C(n_1716),
.Y(n_1920)
);

OAI211xp5_ASAP7_75t_SL g1921 ( 
.A1(n_1912),
.A2(n_1841),
.B(n_1806),
.C(n_1787),
.Y(n_1921)
);

AOI22xp5_ASAP7_75t_L g1922 ( 
.A1(n_1908),
.A2(n_1759),
.B1(n_1720),
.B2(n_1726),
.Y(n_1922)
);

NAND5xp2_ASAP7_75t_L g1923 ( 
.A(n_1910),
.B(n_1529),
.C(n_1520),
.D(n_1590),
.E(n_1587),
.Y(n_1923)
);

AOI21xp5_ASAP7_75t_L g1924 ( 
.A1(n_1923),
.A2(n_1917),
.B(n_1914),
.Y(n_1924)
);

INVxp67_ASAP7_75t_SL g1925 ( 
.A(n_1918),
.Y(n_1925)
);

OAI211xp5_ASAP7_75t_SL g1926 ( 
.A1(n_1919),
.A2(n_1911),
.B(n_1915),
.C(n_1916),
.Y(n_1926)
);

INVx1_ASAP7_75t_L g1927 ( 
.A(n_1921),
.Y(n_1927)
);

AOI221xp5_ASAP7_75t_L g1928 ( 
.A1(n_1920),
.A2(n_1806),
.B1(n_1772),
.B2(n_1724),
.C(n_1520),
.Y(n_1928)
);

NAND3xp33_ASAP7_75t_L g1929 ( 
.A(n_1922),
.B(n_1529),
.C(n_1596),
.Y(n_1929)
);

OAI221xp5_ASAP7_75t_L g1930 ( 
.A1(n_1919),
.A2(n_1724),
.B1(n_1739),
.B2(n_1745),
.C(n_1761),
.Y(n_1930)
);

NOR3xp33_ASAP7_75t_L g1931 ( 
.A(n_1925),
.B(n_1529),
.C(n_1520),
.Y(n_1931)
);

NOR2x1_ASAP7_75t_L g1932 ( 
.A(n_1926),
.B(n_1759),
.Y(n_1932)
);

INVx1_ASAP7_75t_L g1933 ( 
.A(n_1927),
.Y(n_1933)
);

INVx1_ASAP7_75t_L g1934 ( 
.A(n_1924),
.Y(n_1934)
);

NOR3xp33_ASAP7_75t_L g1935 ( 
.A(n_1928),
.B(n_1720),
.C(n_1726),
.Y(n_1935)
);

INVx1_ASAP7_75t_L g1936 ( 
.A(n_1930),
.Y(n_1936)
);

NOR2xp33_ASAP7_75t_L g1937 ( 
.A(n_1934),
.B(n_1929),
.Y(n_1937)
);

INVx1_ASAP7_75t_L g1938 ( 
.A(n_1933),
.Y(n_1938)
);

NAND4xp25_ASAP7_75t_L g1939 ( 
.A(n_1931),
.B(n_1633),
.C(n_1726),
.D(n_1709),
.Y(n_1939)
);

NAND2xp5_ASAP7_75t_L g1940 ( 
.A(n_1938),
.B(n_1932),
.Y(n_1940)
);

HB1xp67_ASAP7_75t_L g1941 ( 
.A(n_1940),
.Y(n_1941)
);

NAND2xp5_ASAP7_75t_L g1942 ( 
.A(n_1941),
.B(n_1936),
.Y(n_1942)
);

OAI22x1_ASAP7_75t_L g1943 ( 
.A1(n_1941),
.A2(n_1937),
.B1(n_1939),
.B2(n_1935),
.Y(n_1943)
);

OAI22x1_ASAP7_75t_SL g1944 ( 
.A1(n_1942),
.A2(n_1752),
.B1(n_1742),
.B2(n_1761),
.Y(n_1944)
);

OAI22xp5_ASAP7_75t_L g1945 ( 
.A1(n_1943),
.A2(n_1752),
.B1(n_1742),
.B2(n_1761),
.Y(n_1945)
);

AO21x2_ASAP7_75t_L g1946 ( 
.A1(n_1945),
.A2(n_1742),
.B(n_1761),
.Y(n_1946)
);

HB1xp67_ASAP7_75t_L g1947 ( 
.A(n_1944),
.Y(n_1947)
);

AOI221x1_ASAP7_75t_L g1948 ( 
.A1(n_1947),
.A2(n_1764),
.B1(n_1741),
.B2(n_1742),
.C(n_1752),
.Y(n_1948)
);

INVx1_ASAP7_75t_L g1949 ( 
.A(n_1948),
.Y(n_1949)
);

OAI22xp33_ASAP7_75t_L g1950 ( 
.A1(n_1949),
.A2(n_1946),
.B1(n_1741),
.B2(n_1752),
.Y(n_1950)
);

AOI221xp5_ASAP7_75t_L g1951 ( 
.A1(n_1950),
.A2(n_1946),
.B1(n_1764),
.B2(n_1741),
.C(n_1528),
.Y(n_1951)
);

AOI211xp5_ASAP7_75t_L g1952 ( 
.A1(n_1951),
.A2(n_1597),
.B(n_1634),
.C(n_1741),
.Y(n_1952)
);


endmodule