module fake_netlist_6_817_n_2072 (n_52, n_435, n_1, n_91, n_326, n_256, n_440, n_507, n_209, n_367, n_465, n_63, n_223, n_278, n_341, n_362, n_148, n_226, n_161, n_22, n_208, n_462, n_68, n_316, n_419, n_28, n_304, n_212, n_50, n_7, n_144, n_365, n_125, n_168, n_384, n_297, n_524, n_342, n_77, n_106, n_358, n_160, n_449, n_131, n_188, n_310, n_509, n_186, n_245, n_0, n_368, n_396, n_495, n_350, n_78, n_84, n_568, n_392, n_442, n_480, n_142, n_143, n_382, n_180, n_62, n_557, n_349, n_233, n_255, n_284, n_400, n_140, n_337, n_214, n_485, n_67, n_15, n_443, n_246, n_38, n_471, n_289, n_421, n_424, n_59, n_181, n_182, n_238, n_202, n_320, n_108, n_327, n_369, n_280, n_287, n_353, n_555, n_389, n_415, n_65, n_230, n_461, n_141, n_383, n_200, n_447, n_176, n_114, n_86, n_198, n_104, n_222, n_179, n_248, n_300, n_517, n_71, n_74, n_229, n_542, n_305, n_72, n_532, n_173, n_535, n_250, n_372, n_468, n_544, n_111, n_504, n_314, n_378, n_413, n_377, n_35, n_183, n_510, n_79, n_375, n_338, n_522, n_466, n_506, n_56, n_360, n_119, n_235, n_536, n_147, n_191, n_340, n_387, n_452, n_39, n_344, n_73, n_428, n_432, n_101, n_167, n_174, n_127, n_516, n_153, n_525, n_156, n_491, n_145, n_42, n_133, n_96, n_8, n_371, n_567, n_189, n_405, n_213, n_538, n_294, n_302, n_499, n_380, n_129, n_197, n_11, n_137, n_17, n_343, n_448, n_20, n_494, n_539, n_493, n_397, n_155, n_109, n_529, n_445, n_425, n_122, n_45, n_454, n_34, n_218, n_70, n_234, n_37, n_486, n_381, n_82, n_27, n_236, n_112, n_172, n_472, n_270, n_239, n_126, n_414, n_97, n_563, n_58, n_490, n_290, n_220, n_118, n_224, n_48, n_25, n_93, n_80, n_196, n_402, n_352, n_478, n_9, n_460, n_107, n_6, n_417, n_14, n_446, n_498, n_89, n_374, n_366, n_407, n_450, n_103, n_272, n_526, n_185, n_348, n_69, n_376, n_390, n_473, n_293, n_31, n_334, n_559, n_53, n_370, n_44, n_458, n_232, n_16, n_163, n_46, n_330, n_470, n_475, n_298, n_18, n_492, n_281, n_258, n_551, n_154, n_456, n_564, n_98, n_260, n_265, n_313, n_451, n_279, n_252, n_228, n_565, n_356, n_166, n_184, n_552, n_216, n_455, n_83, n_521, n_363, n_395, n_323, n_393, n_411, n_503, n_152, n_92, n_513, n_321, n_331, n_105, n_227, n_132, n_570, n_406, n_483, n_102, n_204, n_482, n_474, n_527, n_261, n_420, n_312, n_394, n_32, n_66, n_130, n_519, n_541, n_512, n_164, n_292, n_100, n_121, n_307, n_469, n_433, n_500, n_23, n_476, n_2, n_291, n_219, n_543, n_357, n_150, n_264, n_263, n_481, n_325, n_329, n_464, n_561, n_33, n_477, n_549, n_533, n_408, n_61, n_237, n_244, n_399, n_76, n_243, n_124, n_548, n_94, n_282, n_436, n_116, n_211, n_523, n_117, n_175, n_322, n_345, n_409, n_231, n_354, n_40, n_505, n_240, n_139, n_319, n_41, n_134, n_547, n_537, n_273, n_558, n_95, n_311, n_10, n_403, n_253, n_123, n_136, n_546, n_562, n_249, n_201, n_386, n_556, n_159, n_157, n_162, n_115, n_487, n_550, n_128, n_241, n_30, n_275, n_553, n_43, n_560, n_276, n_569, n_441, n_221, n_444, n_423, n_146, n_318, n_303, n_511, n_467, n_306, n_21, n_193, n_269, n_359, n_346, n_88, n_3, n_416, n_530, n_277, n_520, n_418, n_113, n_4, n_199, n_138, n_266, n_296, n_268, n_271, n_404, n_439, n_158, n_217, n_49, n_210, n_299, n_518, n_206, n_5, n_453, n_333, n_215, n_178, n_247, n_225, n_308, n_309, n_355, n_426, n_317, n_149, n_431, n_90, n_347, n_24, n_459, n_54, n_502, n_328, n_534, n_488, n_429, n_373, n_87, n_195, n_285, n_497, n_85, n_99, n_257, n_13, n_203, n_286, n_254, n_207, n_242, n_19, n_47, n_29, n_75, n_401, n_324, n_335, n_430, n_463, n_545, n_489, n_205, n_120, n_251, n_301, n_274, n_110, n_151, n_412, n_81, n_36, n_26, n_55, n_267, n_438, n_339, n_315, n_434, n_515, n_64, n_288, n_427, n_479, n_496, n_422, n_135, n_165, n_351, n_437, n_259, n_177, n_540, n_514, n_528, n_391, n_457, n_364, n_295, n_385, n_388, n_190, n_262, n_484, n_187, n_501, n_531, n_60, n_361, n_508, n_379, n_170, n_332, n_336, n_12, n_398, n_410, n_566, n_554, n_194, n_171, n_192, n_57, n_169, n_51, n_283, n_2072);

input n_52;
input n_435;
input n_1;
input n_91;
input n_326;
input n_256;
input n_440;
input n_507;
input n_209;
input n_367;
input n_465;
input n_63;
input n_223;
input n_278;
input n_341;
input n_362;
input n_148;
input n_226;
input n_161;
input n_22;
input n_208;
input n_462;
input n_68;
input n_316;
input n_419;
input n_28;
input n_304;
input n_212;
input n_50;
input n_7;
input n_144;
input n_365;
input n_125;
input n_168;
input n_384;
input n_297;
input n_524;
input n_342;
input n_77;
input n_106;
input n_358;
input n_160;
input n_449;
input n_131;
input n_188;
input n_310;
input n_509;
input n_186;
input n_245;
input n_0;
input n_368;
input n_396;
input n_495;
input n_350;
input n_78;
input n_84;
input n_568;
input n_392;
input n_442;
input n_480;
input n_142;
input n_143;
input n_382;
input n_180;
input n_62;
input n_557;
input n_349;
input n_233;
input n_255;
input n_284;
input n_400;
input n_140;
input n_337;
input n_214;
input n_485;
input n_67;
input n_15;
input n_443;
input n_246;
input n_38;
input n_471;
input n_289;
input n_421;
input n_424;
input n_59;
input n_181;
input n_182;
input n_238;
input n_202;
input n_320;
input n_108;
input n_327;
input n_369;
input n_280;
input n_287;
input n_353;
input n_555;
input n_389;
input n_415;
input n_65;
input n_230;
input n_461;
input n_141;
input n_383;
input n_200;
input n_447;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_222;
input n_179;
input n_248;
input n_300;
input n_517;
input n_71;
input n_74;
input n_229;
input n_542;
input n_305;
input n_72;
input n_532;
input n_173;
input n_535;
input n_250;
input n_372;
input n_468;
input n_544;
input n_111;
input n_504;
input n_314;
input n_378;
input n_413;
input n_377;
input n_35;
input n_183;
input n_510;
input n_79;
input n_375;
input n_338;
input n_522;
input n_466;
input n_506;
input n_56;
input n_360;
input n_119;
input n_235;
input n_536;
input n_147;
input n_191;
input n_340;
input n_387;
input n_452;
input n_39;
input n_344;
input n_73;
input n_428;
input n_432;
input n_101;
input n_167;
input n_174;
input n_127;
input n_516;
input n_153;
input n_525;
input n_156;
input n_491;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_371;
input n_567;
input n_189;
input n_405;
input n_213;
input n_538;
input n_294;
input n_302;
input n_499;
input n_380;
input n_129;
input n_197;
input n_11;
input n_137;
input n_17;
input n_343;
input n_448;
input n_20;
input n_494;
input n_539;
input n_493;
input n_397;
input n_155;
input n_109;
input n_529;
input n_445;
input n_425;
input n_122;
input n_45;
input n_454;
input n_34;
input n_218;
input n_70;
input n_234;
input n_37;
input n_486;
input n_381;
input n_82;
input n_27;
input n_236;
input n_112;
input n_172;
input n_472;
input n_270;
input n_239;
input n_126;
input n_414;
input n_97;
input n_563;
input n_58;
input n_490;
input n_290;
input n_220;
input n_118;
input n_224;
input n_48;
input n_25;
input n_93;
input n_80;
input n_196;
input n_402;
input n_352;
input n_478;
input n_9;
input n_460;
input n_107;
input n_6;
input n_417;
input n_14;
input n_446;
input n_498;
input n_89;
input n_374;
input n_366;
input n_407;
input n_450;
input n_103;
input n_272;
input n_526;
input n_185;
input n_348;
input n_69;
input n_376;
input n_390;
input n_473;
input n_293;
input n_31;
input n_334;
input n_559;
input n_53;
input n_370;
input n_44;
input n_458;
input n_232;
input n_16;
input n_163;
input n_46;
input n_330;
input n_470;
input n_475;
input n_298;
input n_18;
input n_492;
input n_281;
input n_258;
input n_551;
input n_154;
input n_456;
input n_564;
input n_98;
input n_260;
input n_265;
input n_313;
input n_451;
input n_279;
input n_252;
input n_228;
input n_565;
input n_356;
input n_166;
input n_184;
input n_552;
input n_216;
input n_455;
input n_83;
input n_521;
input n_363;
input n_395;
input n_323;
input n_393;
input n_411;
input n_503;
input n_152;
input n_92;
input n_513;
input n_321;
input n_331;
input n_105;
input n_227;
input n_132;
input n_570;
input n_406;
input n_483;
input n_102;
input n_204;
input n_482;
input n_474;
input n_527;
input n_261;
input n_420;
input n_312;
input n_394;
input n_32;
input n_66;
input n_130;
input n_519;
input n_541;
input n_512;
input n_164;
input n_292;
input n_100;
input n_121;
input n_307;
input n_469;
input n_433;
input n_500;
input n_23;
input n_476;
input n_2;
input n_291;
input n_219;
input n_543;
input n_357;
input n_150;
input n_264;
input n_263;
input n_481;
input n_325;
input n_329;
input n_464;
input n_561;
input n_33;
input n_477;
input n_549;
input n_533;
input n_408;
input n_61;
input n_237;
input n_244;
input n_399;
input n_76;
input n_243;
input n_124;
input n_548;
input n_94;
input n_282;
input n_436;
input n_116;
input n_211;
input n_523;
input n_117;
input n_175;
input n_322;
input n_345;
input n_409;
input n_231;
input n_354;
input n_40;
input n_505;
input n_240;
input n_139;
input n_319;
input n_41;
input n_134;
input n_547;
input n_537;
input n_273;
input n_558;
input n_95;
input n_311;
input n_10;
input n_403;
input n_253;
input n_123;
input n_136;
input n_546;
input n_562;
input n_249;
input n_201;
input n_386;
input n_556;
input n_159;
input n_157;
input n_162;
input n_115;
input n_487;
input n_550;
input n_128;
input n_241;
input n_30;
input n_275;
input n_553;
input n_43;
input n_560;
input n_276;
input n_569;
input n_441;
input n_221;
input n_444;
input n_423;
input n_146;
input n_318;
input n_303;
input n_511;
input n_467;
input n_306;
input n_21;
input n_193;
input n_269;
input n_359;
input n_346;
input n_88;
input n_3;
input n_416;
input n_530;
input n_277;
input n_520;
input n_418;
input n_113;
input n_4;
input n_199;
input n_138;
input n_266;
input n_296;
input n_268;
input n_271;
input n_404;
input n_439;
input n_158;
input n_217;
input n_49;
input n_210;
input n_299;
input n_518;
input n_206;
input n_5;
input n_453;
input n_333;
input n_215;
input n_178;
input n_247;
input n_225;
input n_308;
input n_309;
input n_355;
input n_426;
input n_317;
input n_149;
input n_431;
input n_90;
input n_347;
input n_24;
input n_459;
input n_54;
input n_502;
input n_328;
input n_534;
input n_488;
input n_429;
input n_373;
input n_87;
input n_195;
input n_285;
input n_497;
input n_85;
input n_99;
input n_257;
input n_13;
input n_203;
input n_286;
input n_254;
input n_207;
input n_242;
input n_19;
input n_47;
input n_29;
input n_75;
input n_401;
input n_324;
input n_335;
input n_430;
input n_463;
input n_545;
input n_489;
input n_205;
input n_120;
input n_251;
input n_301;
input n_274;
input n_110;
input n_151;
input n_412;
input n_81;
input n_36;
input n_26;
input n_55;
input n_267;
input n_438;
input n_339;
input n_315;
input n_434;
input n_515;
input n_64;
input n_288;
input n_427;
input n_479;
input n_496;
input n_422;
input n_135;
input n_165;
input n_351;
input n_437;
input n_259;
input n_177;
input n_540;
input n_514;
input n_528;
input n_391;
input n_457;
input n_364;
input n_295;
input n_385;
input n_388;
input n_190;
input n_262;
input n_484;
input n_187;
input n_501;
input n_531;
input n_60;
input n_361;
input n_508;
input n_379;
input n_170;
input n_332;
input n_336;
input n_12;
input n_398;
input n_410;
input n_566;
input n_554;
input n_194;
input n_171;
input n_192;
input n_57;
input n_169;
input n_51;
input n_283;

output n_2072;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_1212;
wire n_726;
wire n_700;
wire n_1307;
wire n_2003;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_1853;
wire n_783;
wire n_1738;
wire n_798;
wire n_1575;
wire n_1854;
wire n_1923;
wire n_1342;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_1739;
wire n_2051;
wire n_1380;
wire n_1402;
wire n_1688;
wire n_1691;
wire n_1975;
wire n_1009;
wire n_1743;
wire n_1930;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1991;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_1844;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_1786;
wire n_830;
wire n_873;
wire n_1371;
wire n_1285;
wire n_1985;
wire n_1803;
wire n_1172;
wire n_852;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1867;
wire n_1704;
wire n_1078;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_2019;
wire n_836;
wire n_1261;
wire n_945;
wire n_1649;
wire n_2018;
wire n_1903;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_616;
wire n_658;
wire n_1874;
wire n_1119;
wire n_2013;
wire n_1433;
wire n_1902;
wire n_1842;
wire n_1620;
wire n_2044;
wire n_1954;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1798;
wire n_1550;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_940;
wire n_770;
wire n_1781;
wire n_1971;
wire n_2058;
wire n_2004;
wire n_1106;
wire n_886;
wire n_1471;
wire n_953;
wire n_1094;
wire n_1345;
wire n_1820;
wire n_1421;
wire n_1936;
wire n_638;
wire n_1404;
wire n_1211;
wire n_887;
wire n_1660;
wire n_1961;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_1894;
wire n_1231;
wire n_1978;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_1815;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_1193;
wire n_1967;
wire n_1054;
wire n_1333;
wire n_1648;
wire n_1911;
wire n_1956;
wire n_1644;
wire n_2011;
wire n_1558;
wire n_1732;
wire n_699;
wire n_1986;
wire n_824;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_1918;
wire n_577;
wire n_1843;
wire n_619;
wire n_1367;
wire n_1336;
wire n_572;
wire n_813;
wire n_1909;
wire n_1481;
wire n_606;
wire n_1441;
wire n_818;
wire n_1309;
wire n_1123;
wire n_645;
wire n_1381;
wire n_1699;
wire n_916;
wire n_1970;
wire n_608;
wire n_630;
wire n_2059;
wire n_792;
wire n_1328;
wire n_1957;
wire n_1907;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_982;
wire n_1762;
wire n_1910;
wire n_1075;
wire n_932;
wire n_1876;
wire n_1895;
wire n_1697;
wire n_979;
wire n_1873;
wire n_905;
wire n_1866;
wire n_1680;
wire n_993;
wire n_689;
wire n_2031;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1988;
wire n_1278;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_2009;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_2068;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_1354;
wire n_586;
wire n_1875;
wire n_1865;
wire n_1701;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_1950;
wire n_1563;
wire n_1912;
wire n_1982;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_1335;
wire n_1760;
wire n_1927;
wire n_2028;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_1165;
wire n_702;
wire n_2008;
wire n_1926;
wire n_1175;
wire n_1386;
wire n_1896;
wire n_1747;
wire n_1012;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1977;
wire n_1802;
wire n_1504;
wire n_1655;
wire n_835;
wire n_928;
wire n_1214;
wire n_850;
wire n_690;
wire n_1886;
wire n_1801;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_1813;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_1124;
wire n_1624;
wire n_1965;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_1082;
wire n_1317;
wire n_593;
wire n_697;
wire n_687;
wire n_890;
wire n_637;
wire n_701;
wire n_950;
wire n_2036;
wire n_1709;
wire n_1825;
wire n_1757;
wire n_1796;
wire n_1792;
wire n_891;
wire n_2067;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_1987;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_1990;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_595;
wire n_627;
wire n_1767;
wire n_1779;
wire n_1465;
wire n_1858;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_673;
wire n_1969;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_1968;
wire n_898;
wire n_1952;
wire n_865;
wire n_925;
wire n_1932;
wire n_1101;
wire n_1026;
wire n_1880;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_1839;
wire n_685;
wire n_1765;
wire n_605;
wire n_1514;
wire n_1863;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_996;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_791;
wire n_1913;
wire n_837;
wire n_1488;
wire n_1808;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_1947;
wire n_1788;
wire n_1999;
wire n_622;
wire n_1469;
wire n_2060;
wire n_1838;
wire n_1835;
wire n_1776;
wire n_1766;
wire n_1959;
wire n_2002;
wire n_581;
wire n_765;
wire n_1492;
wire n_987;
wire n_1340;
wire n_1771;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_1878;
wire n_899;
wire n_738;
wire n_2012;
wire n_1304;
wire n_1035;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_2069;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_1577;
wire n_1181;
wire n_1822;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_1992;
wire n_648;
wire n_657;
wire n_1049;
wire n_2057;
wire n_1666;
wire n_1505;
wire n_803;
wire n_1717;
wire n_926;
wire n_1817;
wire n_927;
wire n_1849;
wire n_919;
wire n_1698;
wire n_929;
wire n_1228;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_912;
wire n_1857;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_1955;
wire n_755;
wire n_931;
wire n_1021;
wire n_683;
wire n_811;
wire n_1207;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_1250;
wire n_1137;
wire n_1897;
wire n_2064;
wire n_880;
wire n_2053;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_1942;
wire n_1966;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_1837;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_1440;
wire n_2063;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_1483;
wire n_1834;
wire n_1372;
wire n_1457;
wire n_1719;
wire n_1339;
wire n_1787;
wire n_1993;
wire n_1427;
wire n_1466;
wire n_1919;
wire n_1080;
wire n_723;
wire n_1877;
wire n_596;
wire n_1141;
wire n_1268;
wire n_1939;
wire n_2030;
wire n_1769;
wire n_1220;
wire n_1893;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_2025;
wire n_1125;
wire n_970;
wire n_1980;
wire n_642;
wire n_995;
wire n_1159;
wire n_1092;
wire n_1060;
wire n_1951;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_1286;
wire n_1775;
wire n_1773;
wire n_1053;
wire n_1681;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_775;
wire n_651;
wire n_1153;
wire n_1618;
wire n_1531;
wire n_1185;
wire n_1745;
wire n_914;
wire n_759;
wire n_1831;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_773;
wire n_1901;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1892;
wire n_1933;
wire n_1135;
wire n_1179;
wire n_1169;
wire n_1617;
wire n_1470;
wire n_1243;
wire n_848;
wire n_1096;
wire n_1091;
wire n_1917;
wire n_2000;
wire n_1580;
wire n_1425;
wire n_1881;
wire n_1267;
wire n_1281;
wire n_1806;
wire n_983;
wire n_2023;
wire n_1520;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_1731;
wire n_1855;
wire n_1636;
wire n_1437;
wire n_1832;
wire n_1645;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_2049;
wire n_1331;
wire n_613;
wire n_736;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_778;
wire n_1668;
wire n_1134;
wire n_1129;
wire n_602;
wire n_1696;
wire n_1995;
wire n_1594;
wire n_664;
wire n_1869;
wire n_1764;
wire n_1429;
wire n_1610;
wire n_1889;
wire n_1905;
wire n_2016;
wire n_793;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_1937;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_1744;
wire n_828;
wire n_607;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_952;
wire n_725;
wire n_999;
wire n_1254;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_724;
wire n_1934;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_1871;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_1549;
wire n_1510;
wire n_892;
wire n_768;
wire n_1468;
wire n_1859;
wire n_1095;
wire n_2024;
wire n_1595;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_1916;
wire n_597;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1852;
wire n_1024;
wire n_1768;
wire n_1847;
wire n_2052;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_923;
wire n_1409;
wire n_1841;
wire n_1639;
wire n_1623;
wire n_1015;
wire n_1503;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_1126;
wire n_1997;
wire n_710;
wire n_1108;
wire n_1818;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1960;
wire n_2061;
wire n_1686;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1943;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_1694;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_1983;
wire n_1938;
wire n_1262;
wire n_1891;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_2037;
wire n_782;
wire n_1539;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_1472;
wire n_2050;
wire n_1081;
wire n_1870;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_1827;
wire n_1361;
wire n_1864;
wire n_2006;
wire n_1491;
wire n_662;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_2017;
wire n_1695;
wire n_1828;
wire n_2046;
wire n_650;
wire n_1046;
wire n_1940;
wire n_1979;
wire n_1145;
wire n_1121;
wire n_1102;
wire n_1963;
wire n_972;
wire n_1405;
wire n_1406;
wire n_1332;
wire n_624;
wire n_962;
wire n_1041;
wire n_1569;
wire n_936;
wire n_1883;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_1222;
wire n_599;
wire n_776;
wire n_1823;
wire n_1974;
wire n_1720;
wire n_934;
wire n_1637;
wire n_1407;
wire n_1795;
wire n_1341;
wire n_1456;
wire n_1845;
wire n_1489;
wire n_942;
wire n_1524;
wire n_1964;
wire n_1920;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_2007;
wire n_2039;
wire n_1946;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_1640;
wire n_804;
wire n_1846;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_1343;
wire n_1522;
wire n_1782;
wire n_1676;
wire n_833;
wire n_1830;
wire n_1567;
wire n_1319;
wire n_707;
wire n_1900;
wire n_799;
wire n_1548;
wire n_1155;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_2021;
wire n_1086;
wire n_1066;
wire n_1948;
wire n_2026;
wire n_1282;
wire n_652;
wire n_1906;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_1758;
wire n_1925;
wire n_737;
wire n_1318;
wire n_1914;
wire n_1235;
wire n_1229;
wire n_1292;
wire n_1373;
wire n_1029;
wire n_1447;
wire n_2056;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_1248;
wire n_1556;
wire n_902;
wire n_1047;
wire n_1984;
wire n_1385;
wire n_1269;
wire n_1931;
wire n_672;
wire n_1257;
wire n_1751;
wire n_1375;
wire n_1941;
wire n_655;
wire n_706;
wire n_1045;
wire n_1794;
wire n_786;
wire n_1650;
wire n_1236;
wire n_1962;
wire n_1559;
wire n_1725;
wire n_1928;
wire n_1872;
wire n_834;
wire n_743;
wire n_766;
wire n_1741;
wire n_1325;
wire n_1002;
wire n_1746;
wire n_1949;
wire n_1804;
wire n_1727;
wire n_1019;
wire n_636;
wire n_2054;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_2062;
wire n_2041;
wire n_1477;
wire n_1360;
wire n_1860;
wire n_1904;
wire n_1200;
wire n_2070;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1908;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_1098;
wire n_1329;
wire n_2045;
wire n_817;
wire n_897;
wire n_846;
wire n_2066;
wire n_841;
wire n_1476;
wire n_1001;
wire n_1800;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_1191;
wire n_1826;
wire n_1023;
wire n_1882;
wire n_1076;
wire n_1118;
wire n_1007;
wire n_1807;
wire n_1929;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1814;
wire n_1631;
wire n_591;
wire n_1377;
wire n_1879;
wire n_853;
wire n_695;
wire n_1542;
wire n_875;
wire n_680;
wire n_1678;
wire n_661;
wire n_1716;
wire n_1256;
wire n_671;
wire n_1953;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_1976;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1824;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_1516;
wire n_1536;
wire n_2029;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_1074;
wire n_698;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_955;
wire n_1379;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_1810;
wire n_573;
wire n_769;
wire n_676;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_814;
wire n_1643;
wire n_2020;
wire n_1729;
wire n_669;
wire n_2048;
wire n_2005;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_691;
wire n_1408;
wire n_1196;
wire n_1598;
wire n_863;
wire n_601;
wire n_1283;
wire n_918;
wire n_748;
wire n_1848;
wire n_1114;
wire n_1785;
wire n_1147;
wire n_763;
wire n_1754;
wire n_1506;
wire n_1652;
wire n_1812;
wire n_957;
wire n_1994;
wire n_895;
wire n_866;
wire n_1227;
wire n_744;
wire n_971;
wire n_946;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_1173;
wire n_1924;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_1174;
wire n_1944;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_844;
wire n_1017;
wire n_1083;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_2022;
wire n_1945;
wire n_910;
wire n_1721;
wire n_1656;
wire n_1460;
wire n_911;
wire n_1464;
wire n_653;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_2034;
wire n_576;
wire n_1028;
wire n_1922;
wire n_2032;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_1973;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1821;
wire n_1104;
wire n_854;
wire n_1058;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_712;
wire n_1276;
wire n_2015;
wire n_1148;
wire n_1989;
wire n_1161;
wire n_1085;
wire n_2014;
wire n_2042;
wire n_1239;
wire n_771;
wire n_1584;
wire n_924;
wire n_1582;
wire n_1149;
wire n_1184;
wire n_719;
wire n_1972;
wire n_1525;
wire n_1585;
wire n_1851;
wire n_1799;
wire n_1090;
wire n_592;
wire n_1816;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_984;
wire n_1829;
wire n_2035;
wire n_1450;
wire n_1638;
wire n_868;
wire n_859;
wire n_2033;
wire n_735;
wire n_1789;
wire n_1770;
wire n_878;
wire n_620;
wire n_1218;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_1144;
wire n_2071;
wire n_985;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_980;
wire n_1306;
wire n_2010;
wire n_1651;
wire n_1198;
wire n_2047;
wire n_1609;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1998;
wire n_1574;
wire n_756;
wire n_1619;
wire n_1981;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_1552;
wire n_583;
wire n_1996;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_2043;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_849;
wire n_753;
wire n_1753;
wire n_973;
wire n_1921;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_2065;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_2001;
wire n_1884;
wire n_2040;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_1260;
wire n_1819;
wire n_2055;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_2038;
wire n_812;
wire n_1131;
wire n_1761;
wire n_1578;
wire n_1006;
wire n_1861;
wire n_1632;
wire n_1890;
wire n_1805;
wire n_1557;
wire n_1888;
wire n_1833;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_1850;
wire n_1898;
wire n_1868;
wire n_1089;
wire n_1887;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_1242;
wire n_1836;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_640;
wire n_1322;
wire n_965;
wire n_1899;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_1862;
wire n_1856;
wire n_1958;
wire n_784;
wire n_1059;
wire n_1197;
wire n_722;
wire n_862;
wire n_1423;
wire n_1935;
wire n_2027;
wire n_1915;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_827;
wire n_1025;
wire n_1885;
wire n_1013;
wire n_1259;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

INVx1_ASAP7_75t_L g571 ( 
.A(n_264),
.Y(n_571)
);

CKINVDCx5p33_ASAP7_75t_R g572 ( 
.A(n_250),
.Y(n_572)
);

CKINVDCx5p33_ASAP7_75t_R g573 ( 
.A(n_121),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_167),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_294),
.Y(n_575)
);

CKINVDCx5p33_ASAP7_75t_R g576 ( 
.A(n_331),
.Y(n_576)
);

CKINVDCx5p33_ASAP7_75t_R g577 ( 
.A(n_481),
.Y(n_577)
);

CKINVDCx5p33_ASAP7_75t_R g578 ( 
.A(n_545),
.Y(n_578)
);

CKINVDCx5p33_ASAP7_75t_R g579 ( 
.A(n_535),
.Y(n_579)
);

CKINVDCx5p33_ASAP7_75t_R g580 ( 
.A(n_489),
.Y(n_580)
);

CKINVDCx20_ASAP7_75t_R g581 ( 
.A(n_487),
.Y(n_581)
);

CKINVDCx5p33_ASAP7_75t_R g582 ( 
.A(n_200),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_281),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_520),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_526),
.Y(n_585)
);

BUFx5_ASAP7_75t_L g586 ( 
.A(n_527),
.Y(n_586)
);

CKINVDCx5p33_ASAP7_75t_R g587 ( 
.A(n_403),
.Y(n_587)
);

CKINVDCx5p33_ASAP7_75t_R g588 ( 
.A(n_519),
.Y(n_588)
);

CKINVDCx5p33_ASAP7_75t_R g589 ( 
.A(n_180),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_203),
.Y(n_590)
);

BUFx10_ASAP7_75t_L g591 ( 
.A(n_2),
.Y(n_591)
);

CKINVDCx5p33_ASAP7_75t_R g592 ( 
.A(n_52),
.Y(n_592)
);

CKINVDCx5p33_ASAP7_75t_R g593 ( 
.A(n_5),
.Y(n_593)
);

BUFx3_ASAP7_75t_L g594 ( 
.A(n_569),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_4),
.Y(n_595)
);

CKINVDCx16_ASAP7_75t_R g596 ( 
.A(n_292),
.Y(n_596)
);

CKINVDCx5p33_ASAP7_75t_R g597 ( 
.A(n_305),
.Y(n_597)
);

CKINVDCx5p33_ASAP7_75t_R g598 ( 
.A(n_289),
.Y(n_598)
);

CKINVDCx5p33_ASAP7_75t_R g599 ( 
.A(n_532),
.Y(n_599)
);

CKINVDCx5p33_ASAP7_75t_R g600 ( 
.A(n_272),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_211),
.Y(n_601)
);

INVx2_ASAP7_75t_SL g602 ( 
.A(n_541),
.Y(n_602)
);

CKINVDCx20_ASAP7_75t_R g603 ( 
.A(n_278),
.Y(n_603)
);

BUFx10_ASAP7_75t_L g604 ( 
.A(n_214),
.Y(n_604)
);

CKINVDCx5p33_ASAP7_75t_R g605 ( 
.A(n_4),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_469),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_301),
.Y(n_607)
);

CKINVDCx5p33_ASAP7_75t_R g608 ( 
.A(n_252),
.Y(n_608)
);

INVx2_ASAP7_75t_L g609 ( 
.A(n_216),
.Y(n_609)
);

INVx1_ASAP7_75t_SL g610 ( 
.A(n_505),
.Y(n_610)
);

CKINVDCx5p33_ASAP7_75t_R g611 ( 
.A(n_450),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_488),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_448),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_459),
.Y(n_614)
);

BUFx10_ASAP7_75t_L g615 ( 
.A(n_60),
.Y(n_615)
);

CKINVDCx5p33_ASAP7_75t_R g616 ( 
.A(n_521),
.Y(n_616)
);

CKINVDCx5p33_ASAP7_75t_R g617 ( 
.A(n_525),
.Y(n_617)
);

CKINVDCx20_ASAP7_75t_R g618 ( 
.A(n_391),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_539),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_540),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_500),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_536),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_538),
.Y(n_623)
);

CKINVDCx5p33_ASAP7_75t_R g624 ( 
.A(n_333),
.Y(n_624)
);

CKINVDCx5p33_ASAP7_75t_R g625 ( 
.A(n_113),
.Y(n_625)
);

CKINVDCx5p33_ASAP7_75t_R g626 ( 
.A(n_296),
.Y(n_626)
);

CKINVDCx20_ASAP7_75t_R g627 ( 
.A(n_232),
.Y(n_627)
);

INVx3_ASAP7_75t_L g628 ( 
.A(n_76),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_556),
.Y(n_629)
);

CKINVDCx5p33_ASAP7_75t_R g630 ( 
.A(n_68),
.Y(n_630)
);

CKINVDCx5p33_ASAP7_75t_R g631 ( 
.A(n_293),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_139),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_11),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_61),
.Y(n_634)
);

CKINVDCx5p33_ASAP7_75t_R g635 ( 
.A(n_63),
.Y(n_635)
);

CKINVDCx5p33_ASAP7_75t_R g636 ( 
.A(n_446),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_522),
.Y(n_637)
);

CKINVDCx5p33_ASAP7_75t_R g638 ( 
.A(n_51),
.Y(n_638)
);

CKINVDCx5p33_ASAP7_75t_R g639 ( 
.A(n_146),
.Y(n_639)
);

CKINVDCx5p33_ASAP7_75t_R g640 ( 
.A(n_7),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_534),
.Y(n_641)
);

CKINVDCx5p33_ASAP7_75t_R g642 ( 
.A(n_262),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_549),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_492),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_53),
.Y(n_645)
);

CKINVDCx5p33_ASAP7_75t_R g646 ( 
.A(n_473),
.Y(n_646)
);

CKINVDCx5p33_ASAP7_75t_R g647 ( 
.A(n_122),
.Y(n_647)
);

CKINVDCx20_ASAP7_75t_R g648 ( 
.A(n_185),
.Y(n_648)
);

CKINVDCx5p33_ASAP7_75t_R g649 ( 
.A(n_416),
.Y(n_649)
);

CKINVDCx5p33_ASAP7_75t_R g650 ( 
.A(n_373),
.Y(n_650)
);

BUFx6f_ASAP7_75t_L g651 ( 
.A(n_111),
.Y(n_651)
);

BUFx2_ASAP7_75t_L g652 ( 
.A(n_283),
.Y(n_652)
);

CKINVDCx5p33_ASAP7_75t_R g653 ( 
.A(n_524),
.Y(n_653)
);

INVxp67_ASAP7_75t_L g654 ( 
.A(n_436),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_102),
.Y(n_655)
);

CKINVDCx5p33_ASAP7_75t_R g656 ( 
.A(n_421),
.Y(n_656)
);

CKINVDCx5p33_ASAP7_75t_R g657 ( 
.A(n_222),
.Y(n_657)
);

CKINVDCx5p33_ASAP7_75t_R g658 ( 
.A(n_152),
.Y(n_658)
);

INVxp67_ASAP7_75t_L g659 ( 
.A(n_172),
.Y(n_659)
);

CKINVDCx5p33_ASAP7_75t_R g660 ( 
.A(n_362),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_273),
.Y(n_661)
);

CKINVDCx5p33_ASAP7_75t_R g662 ( 
.A(n_45),
.Y(n_662)
);

CKINVDCx5p33_ASAP7_75t_R g663 ( 
.A(n_503),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_173),
.Y(n_664)
);

CKINVDCx5p33_ASAP7_75t_R g665 ( 
.A(n_215),
.Y(n_665)
);

INVx1_ASAP7_75t_SL g666 ( 
.A(n_18),
.Y(n_666)
);

CKINVDCx5p33_ASAP7_75t_R g667 ( 
.A(n_523),
.Y(n_667)
);

HB1xp67_ASAP7_75t_L g668 ( 
.A(n_515),
.Y(n_668)
);

CKINVDCx5p33_ASAP7_75t_R g669 ( 
.A(n_86),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_235),
.Y(n_670)
);

CKINVDCx5p33_ASAP7_75t_R g671 ( 
.A(n_20),
.Y(n_671)
);

CKINVDCx5p33_ASAP7_75t_R g672 ( 
.A(n_455),
.Y(n_672)
);

CKINVDCx5p33_ASAP7_75t_R g673 ( 
.A(n_354),
.Y(n_673)
);

INVx2_ASAP7_75t_L g674 ( 
.A(n_249),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_433),
.Y(n_675)
);

CKINVDCx5p33_ASAP7_75t_R g676 ( 
.A(n_74),
.Y(n_676)
);

HB1xp67_ASAP7_75t_L g677 ( 
.A(n_491),
.Y(n_677)
);

CKINVDCx5p33_ASAP7_75t_R g678 ( 
.A(n_415),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_136),
.Y(n_679)
);

CKINVDCx5p33_ASAP7_75t_R g680 ( 
.A(n_375),
.Y(n_680)
);

CKINVDCx5p33_ASAP7_75t_R g681 ( 
.A(n_404),
.Y(n_681)
);

CKINVDCx5p33_ASAP7_75t_R g682 ( 
.A(n_15),
.Y(n_682)
);

INVx2_ASAP7_75t_L g683 ( 
.A(n_504),
.Y(n_683)
);

CKINVDCx5p33_ASAP7_75t_R g684 ( 
.A(n_224),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_288),
.Y(n_685)
);

BUFx10_ASAP7_75t_L g686 ( 
.A(n_547),
.Y(n_686)
);

CKINVDCx5p33_ASAP7_75t_R g687 ( 
.A(n_371),
.Y(n_687)
);

CKINVDCx5p33_ASAP7_75t_R g688 ( 
.A(n_382),
.Y(n_688)
);

CKINVDCx5p33_ASAP7_75t_R g689 ( 
.A(n_11),
.Y(n_689)
);

CKINVDCx5p33_ASAP7_75t_R g690 ( 
.A(n_542),
.Y(n_690)
);

CKINVDCx5p33_ASAP7_75t_R g691 ( 
.A(n_290),
.Y(n_691)
);

CKINVDCx5p33_ASAP7_75t_R g692 ( 
.A(n_406),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_320),
.Y(n_693)
);

INVx1_ASAP7_75t_SL g694 ( 
.A(n_160),
.Y(n_694)
);

CKINVDCx5p33_ASAP7_75t_R g695 ( 
.A(n_356),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_168),
.Y(n_696)
);

CKINVDCx5p33_ASAP7_75t_R g697 ( 
.A(n_18),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_322),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_280),
.Y(n_699)
);

CKINVDCx5p33_ASAP7_75t_R g700 ( 
.A(n_405),
.Y(n_700)
);

INVx2_ASAP7_75t_L g701 ( 
.A(n_386),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_313),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_530),
.Y(n_703)
);

CKINVDCx5p33_ASAP7_75t_R g704 ( 
.A(n_395),
.Y(n_704)
);

BUFx5_ASAP7_75t_L g705 ( 
.A(n_381),
.Y(n_705)
);

CKINVDCx20_ASAP7_75t_R g706 ( 
.A(n_101),
.Y(n_706)
);

CKINVDCx20_ASAP7_75t_R g707 ( 
.A(n_518),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_64),
.Y(n_708)
);

INVx1_ASAP7_75t_SL g709 ( 
.A(n_531),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_181),
.Y(n_710)
);

CKINVDCx5p33_ASAP7_75t_R g711 ( 
.A(n_226),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_140),
.Y(n_712)
);

CKINVDCx20_ASAP7_75t_R g713 ( 
.A(n_302),
.Y(n_713)
);

CKINVDCx20_ASAP7_75t_R g714 ( 
.A(n_513),
.Y(n_714)
);

INVx2_ASAP7_75t_L g715 ( 
.A(n_279),
.Y(n_715)
);

BUFx3_ASAP7_75t_L g716 ( 
.A(n_102),
.Y(n_716)
);

CKINVDCx5p33_ASAP7_75t_R g717 ( 
.A(n_368),
.Y(n_717)
);

CKINVDCx5p33_ASAP7_75t_R g718 ( 
.A(n_544),
.Y(n_718)
);

CKINVDCx5p33_ASAP7_75t_R g719 ( 
.A(n_287),
.Y(n_719)
);

INVx2_ASAP7_75t_L g720 ( 
.A(n_92),
.Y(n_720)
);

CKINVDCx5p33_ASAP7_75t_R g721 ( 
.A(n_468),
.Y(n_721)
);

CKINVDCx5p33_ASAP7_75t_R g722 ( 
.A(n_335),
.Y(n_722)
);

CKINVDCx5p33_ASAP7_75t_R g723 ( 
.A(n_457),
.Y(n_723)
);

BUFx3_ASAP7_75t_L g724 ( 
.A(n_251),
.Y(n_724)
);

CKINVDCx5p33_ASAP7_75t_R g725 ( 
.A(n_528),
.Y(n_725)
);

CKINVDCx5p33_ASAP7_75t_R g726 ( 
.A(n_149),
.Y(n_726)
);

CKINVDCx5p33_ASAP7_75t_R g727 ( 
.A(n_508),
.Y(n_727)
);

CKINVDCx5p33_ASAP7_75t_R g728 ( 
.A(n_550),
.Y(n_728)
);

CKINVDCx5p33_ASAP7_75t_R g729 ( 
.A(n_543),
.Y(n_729)
);

BUFx6f_ASAP7_75t_L g730 ( 
.A(n_533),
.Y(n_730)
);

INVx1_ASAP7_75t_SL g731 ( 
.A(n_430),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_546),
.Y(n_732)
);

CKINVDCx5p33_ASAP7_75t_R g733 ( 
.A(n_511),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_412),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_175),
.Y(n_735)
);

CKINVDCx5p33_ASAP7_75t_R g736 ( 
.A(n_24),
.Y(n_736)
);

CKINVDCx5p33_ASAP7_75t_R g737 ( 
.A(n_400),
.Y(n_737)
);

CKINVDCx5p33_ASAP7_75t_R g738 ( 
.A(n_559),
.Y(n_738)
);

HB1xp67_ASAP7_75t_L g739 ( 
.A(n_548),
.Y(n_739)
);

CKINVDCx5p33_ASAP7_75t_R g740 ( 
.A(n_26),
.Y(n_740)
);

CKINVDCx5p33_ASAP7_75t_R g741 ( 
.A(n_223),
.Y(n_741)
);

CKINVDCx5p33_ASAP7_75t_R g742 ( 
.A(n_228),
.Y(n_742)
);

CKINVDCx5p33_ASAP7_75t_R g743 ( 
.A(n_129),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_225),
.Y(n_744)
);

CKINVDCx5p33_ASAP7_75t_R g745 ( 
.A(n_529),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_537),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_628),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_628),
.Y(n_748)
);

CKINVDCx5p33_ASAP7_75t_R g749 ( 
.A(n_572),
.Y(n_749)
);

INVxp67_ASAP7_75t_SL g750 ( 
.A(n_668),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_651),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_651),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_651),
.Y(n_753)
);

CKINVDCx20_ASAP7_75t_R g754 ( 
.A(n_581),
.Y(n_754)
);

CKINVDCx14_ASAP7_75t_R g755 ( 
.A(n_652),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_716),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_595),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_633),
.Y(n_758)
);

CKINVDCx5p33_ASAP7_75t_R g759 ( 
.A(n_573),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_634),
.Y(n_760)
);

CKINVDCx5p33_ASAP7_75t_R g761 ( 
.A(n_576),
.Y(n_761)
);

INVxp67_ASAP7_75t_L g762 ( 
.A(n_591),
.Y(n_762)
);

CKINVDCx5p33_ASAP7_75t_R g763 ( 
.A(n_577),
.Y(n_763)
);

CKINVDCx5p33_ASAP7_75t_R g764 ( 
.A(n_578),
.Y(n_764)
);

CKINVDCx5p33_ASAP7_75t_R g765 ( 
.A(n_579),
.Y(n_765)
);

BUFx5_ASAP7_75t_L g766 ( 
.A(n_571),
.Y(n_766)
);

HB1xp67_ASAP7_75t_L g767 ( 
.A(n_592),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_645),
.Y(n_768)
);

CKINVDCx5p33_ASAP7_75t_R g769 ( 
.A(n_580),
.Y(n_769)
);

INVxp67_ASAP7_75t_SL g770 ( 
.A(n_677),
.Y(n_770)
);

INVx1_ASAP7_75t_SL g771 ( 
.A(n_666),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_655),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_708),
.Y(n_773)
);

CKINVDCx20_ASAP7_75t_R g774 ( 
.A(n_603),
.Y(n_774)
);

INVxp67_ASAP7_75t_SL g775 ( 
.A(n_739),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_574),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_575),
.Y(n_777)
);

INVxp67_ASAP7_75t_L g778 ( 
.A(n_591),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_583),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_584),
.Y(n_780)
);

CKINVDCx5p33_ASAP7_75t_R g781 ( 
.A(n_582),
.Y(n_781)
);

CKINVDCx5p33_ASAP7_75t_R g782 ( 
.A(n_587),
.Y(n_782)
);

INVx2_ASAP7_75t_SL g783 ( 
.A(n_615),
.Y(n_783)
);

BUFx6f_ASAP7_75t_L g784 ( 
.A(n_730),
.Y(n_784)
);

CKINVDCx20_ASAP7_75t_R g785 ( 
.A(n_618),
.Y(n_785)
);

INVxp67_ASAP7_75t_SL g786 ( 
.A(n_594),
.Y(n_786)
);

INVx2_ASAP7_75t_L g787 ( 
.A(n_586),
.Y(n_787)
);

CKINVDCx16_ASAP7_75t_R g788 ( 
.A(n_596),
.Y(n_788)
);

INVx1_ASAP7_75t_L g789 ( 
.A(n_585),
.Y(n_789)
);

CKINVDCx20_ASAP7_75t_R g790 ( 
.A(n_627),
.Y(n_790)
);

INVxp67_ASAP7_75t_SL g791 ( 
.A(n_724),
.Y(n_791)
);

CKINVDCx20_ASAP7_75t_R g792 ( 
.A(n_648),
.Y(n_792)
);

BUFx3_ASAP7_75t_L g793 ( 
.A(n_604),
.Y(n_793)
);

INVx1_ASAP7_75t_SL g794 ( 
.A(n_706),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_590),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_601),
.Y(n_796)
);

BUFx2_ASAP7_75t_L g797 ( 
.A(n_593),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_606),
.Y(n_798)
);

CKINVDCx5p33_ASAP7_75t_R g799 ( 
.A(n_588),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_607),
.Y(n_800)
);

INVxp67_ASAP7_75t_SL g801 ( 
.A(n_654),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_612),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_613),
.Y(n_803)
);

INVxp33_ASAP7_75t_SL g804 ( 
.A(n_605),
.Y(n_804)
);

BUFx3_ASAP7_75t_L g805 ( 
.A(n_604),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_614),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_619),
.Y(n_807)
);

CKINVDCx5p33_ASAP7_75t_R g808 ( 
.A(n_589),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_620),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_621),
.Y(n_810)
);

CKINVDCx5p33_ASAP7_75t_R g811 ( 
.A(n_597),
.Y(n_811)
);

INVxp33_ASAP7_75t_L g812 ( 
.A(n_720),
.Y(n_812)
);

CKINVDCx5p33_ASAP7_75t_R g813 ( 
.A(n_598),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_622),
.Y(n_814)
);

INVx3_ASAP7_75t_L g815 ( 
.A(n_615),
.Y(n_815)
);

INVx2_ASAP7_75t_L g816 ( 
.A(n_586),
.Y(n_816)
);

CKINVDCx20_ASAP7_75t_R g817 ( 
.A(n_707),
.Y(n_817)
);

CKINVDCx5p33_ASAP7_75t_R g818 ( 
.A(n_599),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_623),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_629),
.Y(n_820)
);

INVx1_ASAP7_75t_L g821 ( 
.A(n_632),
.Y(n_821)
);

INVx2_ASAP7_75t_L g822 ( 
.A(n_586),
.Y(n_822)
);

CKINVDCx5p33_ASAP7_75t_R g823 ( 
.A(n_600),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_637),
.Y(n_824)
);

CKINVDCx16_ASAP7_75t_R g825 ( 
.A(n_713),
.Y(n_825)
);

INVx1_ASAP7_75t_SL g826 ( 
.A(n_625),
.Y(n_826)
);

INVxp67_ASAP7_75t_SL g827 ( 
.A(n_659),
.Y(n_827)
);

BUFx6f_ASAP7_75t_L g828 ( 
.A(n_730),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_641),
.Y(n_829)
);

BUFx2_ASAP7_75t_L g830 ( 
.A(n_630),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_643),
.Y(n_831)
);

CKINVDCx5p33_ASAP7_75t_R g832 ( 
.A(n_608),
.Y(n_832)
);

INVxp67_ASAP7_75t_SL g833 ( 
.A(n_644),
.Y(n_833)
);

CKINVDCx5p33_ASAP7_75t_R g834 ( 
.A(n_611),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_661),
.Y(n_835)
);

CKINVDCx5p33_ASAP7_75t_R g836 ( 
.A(n_616),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_664),
.Y(n_837)
);

CKINVDCx5p33_ASAP7_75t_R g838 ( 
.A(n_617),
.Y(n_838)
);

HB1xp67_ASAP7_75t_L g839 ( 
.A(n_635),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_670),
.Y(n_840)
);

CKINVDCx20_ASAP7_75t_R g841 ( 
.A(n_714),
.Y(n_841)
);

INVx2_ASAP7_75t_L g842 ( 
.A(n_586),
.Y(n_842)
);

INVxp67_ASAP7_75t_SL g843 ( 
.A(n_675),
.Y(n_843)
);

INVxp33_ASAP7_75t_L g844 ( 
.A(n_679),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_685),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_693),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_696),
.Y(n_847)
);

AOI22xp5_ASAP7_75t_L g848 ( 
.A1(n_788),
.A2(n_638),
.B1(n_662),
.B2(n_640),
.Y(n_848)
);

BUFx2_ASAP7_75t_L g849 ( 
.A(n_762),
.Y(n_849)
);

OA21x2_ASAP7_75t_L g850 ( 
.A1(n_776),
.A2(n_699),
.B(n_698),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_751),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_752),
.Y(n_852)
);

INVx1_ASAP7_75t_L g853 ( 
.A(n_753),
.Y(n_853)
);

INVx5_ASAP7_75t_L g854 ( 
.A(n_784),
.Y(n_854)
);

OAI22xp5_ASAP7_75t_SL g855 ( 
.A1(n_755),
.A2(n_671),
.B1(n_676),
.B2(n_669),
.Y(n_855)
);

INVx5_ASAP7_75t_L g856 ( 
.A(n_784),
.Y(n_856)
);

BUFx2_ASAP7_75t_L g857 ( 
.A(n_778),
.Y(n_857)
);

INVx3_ASAP7_75t_L g858 ( 
.A(n_784),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_828),
.Y(n_859)
);

AOI22xp5_ASAP7_75t_L g860 ( 
.A1(n_750),
.A2(n_682),
.B1(n_697),
.B2(n_689),
.Y(n_860)
);

OA21x2_ASAP7_75t_L g861 ( 
.A1(n_777),
.A2(n_703),
.B(n_702),
.Y(n_861)
);

INVxp67_ASAP7_75t_L g862 ( 
.A(n_771),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_L g863 ( 
.A(n_749),
.B(n_602),
.Y(n_863)
);

AND2x4_ASAP7_75t_L g864 ( 
.A(n_786),
.B(n_609),
.Y(n_864)
);

INVx2_ASAP7_75t_L g865 ( 
.A(n_828),
.Y(n_865)
);

BUFx8_ASAP7_75t_L g866 ( 
.A(n_797),
.Y(n_866)
);

INVx3_ASAP7_75t_L g867 ( 
.A(n_828),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_L g868 ( 
.A(n_759),
.B(n_674),
.Y(n_868)
);

INVx2_ASAP7_75t_L g869 ( 
.A(n_766),
.Y(n_869)
);

INVx2_ASAP7_75t_L g870 ( 
.A(n_766),
.Y(n_870)
);

OA21x2_ASAP7_75t_L g871 ( 
.A1(n_779),
.A2(n_712),
.B(n_710),
.Y(n_871)
);

BUFx6f_ASAP7_75t_L g872 ( 
.A(n_757),
.Y(n_872)
);

INVx2_ASAP7_75t_L g873 ( 
.A(n_766),
.Y(n_873)
);

INVx3_ASAP7_75t_L g874 ( 
.A(n_787),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_L g875 ( 
.A(n_761),
.B(n_683),
.Y(n_875)
);

INVx1_ASAP7_75t_L g876 ( 
.A(n_780),
.Y(n_876)
);

INVx2_ASAP7_75t_L g877 ( 
.A(n_766),
.Y(n_877)
);

INVx2_ASAP7_75t_L g878 ( 
.A(n_766),
.Y(n_878)
);

BUFx3_ASAP7_75t_L g879 ( 
.A(n_756),
.Y(n_879)
);

INVx2_ASAP7_75t_L g880 ( 
.A(n_758),
.Y(n_880)
);

INVx3_ASAP7_75t_L g881 ( 
.A(n_816),
.Y(n_881)
);

CKINVDCx11_ASAP7_75t_R g882 ( 
.A(n_794),
.Y(n_882)
);

INVx2_ASAP7_75t_L g883 ( 
.A(n_760),
.Y(n_883)
);

AND2x2_ASAP7_75t_L g884 ( 
.A(n_826),
.B(n_791),
.Y(n_884)
);

INVx6_ASAP7_75t_L g885 ( 
.A(n_793),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_789),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_795),
.Y(n_887)
);

INVx1_ASAP7_75t_SL g888 ( 
.A(n_794),
.Y(n_888)
);

AND2x2_ASAP7_75t_L g889 ( 
.A(n_767),
.B(n_686),
.Y(n_889)
);

OAI22xp5_ASAP7_75t_L g890 ( 
.A1(n_770),
.A2(n_740),
.B1(n_736),
.B2(n_610),
.Y(n_890)
);

INVx1_ASAP7_75t_L g891 ( 
.A(n_796),
.Y(n_891)
);

INVx1_ASAP7_75t_L g892 ( 
.A(n_798),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_800),
.Y(n_893)
);

INVx1_ASAP7_75t_L g894 ( 
.A(n_802),
.Y(n_894)
);

INVx2_ASAP7_75t_L g895 ( 
.A(n_768),
.Y(n_895)
);

NAND2xp5_ASAP7_75t_SL g896 ( 
.A(n_771),
.B(n_686),
.Y(n_896)
);

INVx1_ASAP7_75t_L g897 ( 
.A(n_803),
.Y(n_897)
);

CKINVDCx11_ASAP7_75t_R g898 ( 
.A(n_754),
.Y(n_898)
);

INVx1_ASAP7_75t_L g899 ( 
.A(n_806),
.Y(n_899)
);

HB1xp67_ASAP7_75t_L g900 ( 
.A(n_805),
.Y(n_900)
);

INVx2_ASAP7_75t_L g901 ( 
.A(n_772),
.Y(n_901)
);

AOI22xp5_ASAP7_75t_L g902 ( 
.A1(n_775),
.A2(n_804),
.B1(n_827),
.B2(n_801),
.Y(n_902)
);

INVx1_ASAP7_75t_L g903 ( 
.A(n_807),
.Y(n_903)
);

BUFx3_ASAP7_75t_L g904 ( 
.A(n_763),
.Y(n_904)
);

INVx3_ASAP7_75t_L g905 ( 
.A(n_822),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_809),
.Y(n_906)
);

AND2x2_ASAP7_75t_L g907 ( 
.A(n_839),
.B(n_694),
.Y(n_907)
);

AND2x2_ASAP7_75t_L g908 ( 
.A(n_830),
.B(n_709),
.Y(n_908)
);

INVx1_ASAP7_75t_L g909 ( 
.A(n_810),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_L g910 ( 
.A(n_764),
.B(n_701),
.Y(n_910)
);

AOI22xp5_ASAP7_75t_L g911 ( 
.A1(n_783),
.A2(n_731),
.B1(n_624),
.B2(n_631),
.Y(n_911)
);

NOR2x1_ASAP7_75t_L g912 ( 
.A(n_814),
.B(n_732),
.Y(n_912)
);

AND2x4_ASAP7_75t_L g913 ( 
.A(n_815),
.B(n_715),
.Y(n_913)
);

BUFx3_ASAP7_75t_L g914 ( 
.A(n_765),
.Y(n_914)
);

OA21x2_ASAP7_75t_L g915 ( 
.A1(n_819),
.A2(n_821),
.B(n_820),
.Y(n_915)
);

AND2x2_ASAP7_75t_L g916 ( 
.A(n_812),
.B(n_626),
.Y(n_916)
);

BUFx3_ASAP7_75t_L g917 ( 
.A(n_769),
.Y(n_917)
);

AND2x6_ASAP7_75t_L g918 ( 
.A(n_842),
.B(n_730),
.Y(n_918)
);

INVx1_ASAP7_75t_L g919 ( 
.A(n_824),
.Y(n_919)
);

AND2x6_ASAP7_75t_L g920 ( 
.A(n_747),
.B(n_734),
.Y(n_920)
);

INVx2_ASAP7_75t_L g921 ( 
.A(n_773),
.Y(n_921)
);

NOR2xp33_ASAP7_75t_SL g922 ( 
.A(n_825),
.B(n_636),
.Y(n_922)
);

AND2x2_ASAP7_75t_SL g923 ( 
.A(n_815),
.B(n_735),
.Y(n_923)
);

INVx2_ASAP7_75t_L g924 ( 
.A(n_829),
.Y(n_924)
);

INVx1_ASAP7_75t_L g925 ( 
.A(n_831),
.Y(n_925)
);

INVx2_ASAP7_75t_L g926 ( 
.A(n_835),
.Y(n_926)
);

INVx3_ASAP7_75t_L g927 ( 
.A(n_748),
.Y(n_927)
);

NOR2xp33_ASAP7_75t_L g928 ( 
.A(n_781),
.B(n_744),
.Y(n_928)
);

NAND2xp5_ASAP7_75t_L g929 ( 
.A(n_782),
.B(n_746),
.Y(n_929)
);

BUFx6f_ASAP7_75t_L g930 ( 
.A(n_837),
.Y(n_930)
);

INVx6_ASAP7_75t_L g931 ( 
.A(n_844),
.Y(n_931)
);

INVx1_ASAP7_75t_L g932 ( 
.A(n_840),
.Y(n_932)
);

BUFx6f_ASAP7_75t_L g933 ( 
.A(n_845),
.Y(n_933)
);

NOR2xp33_ASAP7_75t_L g934 ( 
.A(n_868),
.B(n_799),
.Y(n_934)
);

NOR2xp33_ASAP7_75t_L g935 ( 
.A(n_875),
.B(n_808),
.Y(n_935)
);

INVx1_ASAP7_75t_L g936 ( 
.A(n_874),
.Y(n_936)
);

BUFx6f_ASAP7_75t_L g937 ( 
.A(n_930),
.Y(n_937)
);

INVx2_ASAP7_75t_L g938 ( 
.A(n_865),
.Y(n_938)
);

INVx2_ASAP7_75t_L g939 ( 
.A(n_858),
.Y(n_939)
);

INVx2_ASAP7_75t_L g940 ( 
.A(n_858),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_L g941 ( 
.A(n_884),
.B(n_811),
.Y(n_941)
);

INVx3_ASAP7_75t_L g942 ( 
.A(n_874),
.Y(n_942)
);

INVx1_ASAP7_75t_L g943 ( 
.A(n_876),
.Y(n_943)
);

NAND2xp5_ASAP7_75t_SL g944 ( 
.A(n_862),
.B(n_813),
.Y(n_944)
);

INVx3_ASAP7_75t_L g945 ( 
.A(n_881),
.Y(n_945)
);

INVx2_ASAP7_75t_L g946 ( 
.A(n_867),
.Y(n_946)
);

INVx2_ASAP7_75t_L g947 ( 
.A(n_867),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_SL g948 ( 
.A(n_923),
.B(n_818),
.Y(n_948)
);

INVx2_ASAP7_75t_L g949 ( 
.A(n_859),
.Y(n_949)
);

INVx2_ASAP7_75t_L g950 ( 
.A(n_851),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_L g951 ( 
.A(n_910),
.B(n_823),
.Y(n_951)
);

CKINVDCx20_ASAP7_75t_R g952 ( 
.A(n_898),
.Y(n_952)
);

NAND2xp5_ASAP7_75t_SL g953 ( 
.A(n_908),
.B(n_832),
.Y(n_953)
);

BUFx6f_ASAP7_75t_SL g954 ( 
.A(n_904),
.Y(n_954)
);

INVx2_ASAP7_75t_L g955 ( 
.A(n_852),
.Y(n_955)
);

BUFx6f_ASAP7_75t_L g956 ( 
.A(n_930),
.Y(n_956)
);

NAND2xp33_ASAP7_75t_L g957 ( 
.A(n_929),
.B(n_863),
.Y(n_957)
);

AND2x2_ASAP7_75t_L g958 ( 
.A(n_931),
.B(n_834),
.Y(n_958)
);

AND2x2_ASAP7_75t_SL g959 ( 
.A(n_922),
.B(n_774),
.Y(n_959)
);

INVx1_ASAP7_75t_L g960 ( 
.A(n_881),
.Y(n_960)
);

INVx1_ASAP7_75t_L g961 ( 
.A(n_886),
.Y(n_961)
);

INVx4_ASAP7_75t_L g962 ( 
.A(n_930),
.Y(n_962)
);

BUFx6f_ASAP7_75t_L g963 ( 
.A(n_933),
.Y(n_963)
);

INVx2_ASAP7_75t_SL g964 ( 
.A(n_931),
.Y(n_964)
);

INVx2_ASAP7_75t_L g965 ( 
.A(n_853),
.Y(n_965)
);

INVx1_ASAP7_75t_L g966 ( 
.A(n_887),
.Y(n_966)
);

INVx1_ASAP7_75t_L g967 ( 
.A(n_891),
.Y(n_967)
);

INVxp33_ASAP7_75t_L g968 ( 
.A(n_882),
.Y(n_968)
);

INVx2_ASAP7_75t_L g969 ( 
.A(n_924),
.Y(n_969)
);

NAND2xp5_ASAP7_75t_SL g970 ( 
.A(n_907),
.B(n_836),
.Y(n_970)
);

INVx1_ASAP7_75t_L g971 ( 
.A(n_892),
.Y(n_971)
);

INVx1_ASAP7_75t_L g972 ( 
.A(n_905),
.Y(n_972)
);

NAND2xp5_ASAP7_75t_SL g973 ( 
.A(n_916),
.B(n_838),
.Y(n_973)
);

INVx2_ASAP7_75t_L g974 ( 
.A(n_926),
.Y(n_974)
);

INVx2_ASAP7_75t_SL g975 ( 
.A(n_889),
.Y(n_975)
);

INVx1_ASAP7_75t_L g976 ( 
.A(n_893),
.Y(n_976)
);

INVx1_ASAP7_75t_L g977 ( 
.A(n_894),
.Y(n_977)
);

INVx1_ASAP7_75t_L g978 ( 
.A(n_897),
.Y(n_978)
);

INVx2_ASAP7_75t_L g979 ( 
.A(n_880),
.Y(n_979)
);

AOI22xp5_ASAP7_75t_L g980 ( 
.A1(n_902),
.A2(n_843),
.B1(n_833),
.B2(n_790),
.Y(n_980)
);

INVx4_ASAP7_75t_L g981 ( 
.A(n_933),
.Y(n_981)
);

BUFx4f_ASAP7_75t_L g982 ( 
.A(n_850),
.Y(n_982)
);

INVx2_ASAP7_75t_L g983 ( 
.A(n_883),
.Y(n_983)
);

INVx2_ASAP7_75t_L g984 ( 
.A(n_895),
.Y(n_984)
);

INVx1_ASAP7_75t_L g985 ( 
.A(n_905),
.Y(n_985)
);

INVx2_ASAP7_75t_L g986 ( 
.A(n_901),
.Y(n_986)
);

INVx2_ASAP7_75t_L g987 ( 
.A(n_921),
.Y(n_987)
);

AOI21x1_ASAP7_75t_L g988 ( 
.A1(n_869),
.A2(n_847),
.B(n_846),
.Y(n_988)
);

NAND2xp5_ASAP7_75t_L g989 ( 
.A(n_928),
.B(n_864),
.Y(n_989)
);

NOR3xp33_ASAP7_75t_L g990 ( 
.A(n_896),
.B(n_745),
.C(n_642),
.Y(n_990)
);

NAND2xp5_ASAP7_75t_L g991 ( 
.A(n_864),
.B(n_639),
.Y(n_991)
);

AND2x2_ASAP7_75t_L g992 ( 
.A(n_888),
.B(n_785),
.Y(n_992)
);

INVx2_ASAP7_75t_L g993 ( 
.A(n_933),
.Y(n_993)
);

INVx2_ASAP7_75t_L g994 ( 
.A(n_872),
.Y(n_994)
);

AND2x2_ASAP7_75t_L g995 ( 
.A(n_849),
.B(n_792),
.Y(n_995)
);

AND2x2_ASAP7_75t_L g996 ( 
.A(n_849),
.B(n_817),
.Y(n_996)
);

INVx3_ASAP7_75t_L g997 ( 
.A(n_854),
.Y(n_997)
);

INVx2_ASAP7_75t_L g998 ( 
.A(n_872),
.Y(n_998)
);

AND2x6_ASAP7_75t_L g999 ( 
.A(n_912),
.B(n_586),
.Y(n_999)
);

AND2x2_ASAP7_75t_L g1000 ( 
.A(n_857),
.B(n_841),
.Y(n_1000)
);

INVx1_ASAP7_75t_L g1001 ( 
.A(n_915),
.Y(n_1001)
);

INVx1_ASAP7_75t_L g1002 ( 
.A(n_915),
.Y(n_1002)
);

NOR2xp33_ASAP7_75t_L g1003 ( 
.A(n_911),
.B(n_722),
.Y(n_1003)
);

INVx2_ASAP7_75t_SL g1004 ( 
.A(n_885),
.Y(n_1004)
);

INVx1_ASAP7_75t_L g1005 ( 
.A(n_899),
.Y(n_1005)
);

INVx1_ASAP7_75t_L g1006 ( 
.A(n_903),
.Y(n_1006)
);

AND3x2_ASAP7_75t_L g1007 ( 
.A(n_857),
.B(n_705),
.C(n_0),
.Y(n_1007)
);

NAND2xp33_ASAP7_75t_L g1008 ( 
.A(n_920),
.B(n_705),
.Y(n_1008)
);

OR2x2_ASAP7_75t_L g1009 ( 
.A(n_890),
.B(n_723),
.Y(n_1009)
);

NAND2xp5_ASAP7_75t_L g1010 ( 
.A(n_920),
.B(n_646),
.Y(n_1010)
);

INVx2_ASAP7_75t_L g1011 ( 
.A(n_872),
.Y(n_1011)
);

INVx2_ASAP7_75t_L g1012 ( 
.A(n_906),
.Y(n_1012)
);

INVx2_ASAP7_75t_SL g1013 ( 
.A(n_885),
.Y(n_1013)
);

AND2x6_ASAP7_75t_L g1014 ( 
.A(n_870),
.B(n_705),
.Y(n_1014)
);

INVx1_ASAP7_75t_L g1015 ( 
.A(n_909),
.Y(n_1015)
);

NAND2xp33_ASAP7_75t_L g1016 ( 
.A(n_920),
.B(n_705),
.Y(n_1016)
);

NAND2xp5_ASAP7_75t_L g1017 ( 
.A(n_919),
.B(n_647),
.Y(n_1017)
);

INVx3_ASAP7_75t_L g1018 ( 
.A(n_854),
.Y(n_1018)
);

NAND2xp33_ASAP7_75t_L g1019 ( 
.A(n_918),
.B(n_705),
.Y(n_1019)
);

AO21x2_ASAP7_75t_L g1020 ( 
.A1(n_848),
.A2(n_650),
.B(n_649),
.Y(n_1020)
);

INVx2_ASAP7_75t_L g1021 ( 
.A(n_925),
.Y(n_1021)
);

INVx2_ASAP7_75t_L g1022 ( 
.A(n_932),
.Y(n_1022)
);

INVx1_ASAP7_75t_L g1023 ( 
.A(n_879),
.Y(n_1023)
);

INVx2_ASAP7_75t_L g1024 ( 
.A(n_927),
.Y(n_1024)
);

INVx3_ASAP7_75t_L g1025 ( 
.A(n_854),
.Y(n_1025)
);

CKINVDCx12_ASAP7_75t_R g1026 ( 
.A(n_855),
.Y(n_1026)
);

OR2x2_ASAP7_75t_L g1027 ( 
.A(n_860),
.B(n_733),
.Y(n_1027)
);

CKINVDCx20_ASAP7_75t_R g1028 ( 
.A(n_952),
.Y(n_1028)
);

INVx1_ASAP7_75t_L g1029 ( 
.A(n_1005),
.Y(n_1029)
);

AND2x2_ASAP7_75t_L g1030 ( 
.A(n_975),
.B(n_914),
.Y(n_1030)
);

INVx1_ASAP7_75t_L g1031 ( 
.A(n_1005),
.Y(n_1031)
);

CKINVDCx20_ASAP7_75t_R g1032 ( 
.A(n_992),
.Y(n_1032)
);

AND2x2_ASAP7_75t_L g1033 ( 
.A(n_958),
.B(n_917),
.Y(n_1033)
);

INVx1_ASAP7_75t_L g1034 ( 
.A(n_1006),
.Y(n_1034)
);

NOR2xp33_ASAP7_75t_L g1035 ( 
.A(n_941),
.B(n_900),
.Y(n_1035)
);

AND2x2_ASAP7_75t_L g1036 ( 
.A(n_989),
.B(n_964),
.Y(n_1036)
);

INVx1_ASAP7_75t_L g1037 ( 
.A(n_1006),
.Y(n_1037)
);

INVx2_ASAP7_75t_L g1038 ( 
.A(n_936),
.Y(n_1038)
);

INVx1_ASAP7_75t_L g1039 ( 
.A(n_1015),
.Y(n_1039)
);

INVx1_ASAP7_75t_L g1040 ( 
.A(n_1015),
.Y(n_1040)
);

INVx1_ASAP7_75t_L g1041 ( 
.A(n_943),
.Y(n_1041)
);

INVx1_ASAP7_75t_L g1042 ( 
.A(n_961),
.Y(n_1042)
);

CKINVDCx20_ASAP7_75t_R g1043 ( 
.A(n_995),
.Y(n_1043)
);

AND2x4_ASAP7_75t_L g1044 ( 
.A(n_1023),
.B(n_913),
.Y(n_1044)
);

INVx1_ASAP7_75t_L g1045 ( 
.A(n_966),
.Y(n_1045)
);

INVx1_ASAP7_75t_L g1046 ( 
.A(n_967),
.Y(n_1046)
);

INVx1_ASAP7_75t_L g1047 ( 
.A(n_971),
.Y(n_1047)
);

AND2x6_ASAP7_75t_L g1048 ( 
.A(n_1001),
.B(n_913),
.Y(n_1048)
);

INVx2_ASAP7_75t_SL g1049 ( 
.A(n_938),
.Y(n_1049)
);

INVx1_ASAP7_75t_L g1050 ( 
.A(n_976),
.Y(n_1050)
);

INVx4_ASAP7_75t_SL g1051 ( 
.A(n_954),
.Y(n_1051)
);

INVx1_ASAP7_75t_L g1052 ( 
.A(n_977),
.Y(n_1052)
);

AND2x4_ASAP7_75t_L g1053 ( 
.A(n_1012),
.B(n_927),
.Y(n_1053)
);

NOR2xp67_ASAP7_75t_L g1054 ( 
.A(n_1004),
.B(n_1013),
.Y(n_1054)
);

INVx1_ASAP7_75t_L g1055 ( 
.A(n_978),
.Y(n_1055)
);

INVx1_ASAP7_75t_L g1056 ( 
.A(n_1021),
.Y(n_1056)
);

INVxp67_ASAP7_75t_L g1057 ( 
.A(n_996),
.Y(n_1057)
);

INVx2_ASAP7_75t_L g1058 ( 
.A(n_936),
.Y(n_1058)
);

CKINVDCx16_ASAP7_75t_R g1059 ( 
.A(n_954),
.Y(n_1059)
);

INVx1_ASAP7_75t_L g1060 ( 
.A(n_1022),
.Y(n_1060)
);

INVx1_ASAP7_75t_L g1061 ( 
.A(n_969),
.Y(n_1061)
);

CKINVDCx5p33_ASAP7_75t_R g1062 ( 
.A(n_959),
.Y(n_1062)
);

NAND2xp5_ASAP7_75t_L g1063 ( 
.A(n_934),
.B(n_935),
.Y(n_1063)
);

AND2x4_ASAP7_75t_L g1064 ( 
.A(n_993),
.B(n_653),
.Y(n_1064)
);

AND2x2_ASAP7_75t_L g1065 ( 
.A(n_944),
.B(n_850),
.Y(n_1065)
);

INVx1_ASAP7_75t_L g1066 ( 
.A(n_974),
.Y(n_1066)
);

XOR2x2_ASAP7_75t_L g1067 ( 
.A(n_1003),
.B(n_1),
.Y(n_1067)
);

INVx1_ASAP7_75t_L g1068 ( 
.A(n_979),
.Y(n_1068)
);

NAND2xp5_ASAP7_75t_L g1069 ( 
.A(n_951),
.B(n_873),
.Y(n_1069)
);

INVx1_ASAP7_75t_L g1070 ( 
.A(n_983),
.Y(n_1070)
);

INVx1_ASAP7_75t_L g1071 ( 
.A(n_984),
.Y(n_1071)
);

INVx1_ASAP7_75t_L g1072 ( 
.A(n_986),
.Y(n_1072)
);

BUFx6f_ASAP7_75t_L g1073 ( 
.A(n_937),
.Y(n_1073)
);

INVx1_ASAP7_75t_L g1074 ( 
.A(n_987),
.Y(n_1074)
);

INVx1_ASAP7_75t_L g1075 ( 
.A(n_1024),
.Y(n_1075)
);

OAI21xp5_ASAP7_75t_L g1076 ( 
.A1(n_982),
.A2(n_1002),
.B(n_1001),
.Y(n_1076)
);

INVx1_ASAP7_75t_L g1077 ( 
.A(n_960),
.Y(n_1077)
);

INVx1_ASAP7_75t_L g1078 ( 
.A(n_960),
.Y(n_1078)
);

NAND2xp33_ASAP7_75t_R g1079 ( 
.A(n_1000),
.B(n_861),
.Y(n_1079)
);

INVx1_ASAP7_75t_L g1080 ( 
.A(n_972),
.Y(n_1080)
);

AND2x2_ASAP7_75t_L g1081 ( 
.A(n_970),
.B(n_861),
.Y(n_1081)
);

INVx1_ASAP7_75t_L g1082 ( 
.A(n_972),
.Y(n_1082)
);

AOI21xp5_ASAP7_75t_L g1083 ( 
.A1(n_982),
.A2(n_878),
.B(n_877),
.Y(n_1083)
);

OAI21xp5_ASAP7_75t_L g1084 ( 
.A1(n_1002),
.A2(n_871),
.B(n_918),
.Y(n_1084)
);

AOI21xp5_ASAP7_75t_L g1085 ( 
.A1(n_957),
.A2(n_991),
.B(n_1017),
.Y(n_1085)
);

NAND2xp5_ASAP7_75t_L g1086 ( 
.A(n_962),
.B(n_871),
.Y(n_1086)
);

INVx1_ASAP7_75t_L g1087 ( 
.A(n_985),
.Y(n_1087)
);

INVx2_ASAP7_75t_L g1088 ( 
.A(n_985),
.Y(n_1088)
);

INVxp67_ASAP7_75t_L g1089 ( 
.A(n_953),
.Y(n_1089)
);

AND2x4_ASAP7_75t_L g1090 ( 
.A(n_994),
.B(n_656),
.Y(n_1090)
);

INVx1_ASAP7_75t_L g1091 ( 
.A(n_950),
.Y(n_1091)
);

INVx1_ASAP7_75t_L g1092 ( 
.A(n_955),
.Y(n_1092)
);

NAND2xp5_ASAP7_75t_SL g1093 ( 
.A(n_937),
.B(n_866),
.Y(n_1093)
);

INVx2_ASAP7_75t_SL g1094 ( 
.A(n_939),
.Y(n_1094)
);

NAND2xp5_ASAP7_75t_SL g1095 ( 
.A(n_937),
.B(n_866),
.Y(n_1095)
);

INVx2_ASAP7_75t_L g1096 ( 
.A(n_988),
.Y(n_1096)
);

NOR2xp33_ASAP7_75t_SL g1097 ( 
.A(n_968),
.B(n_657),
.Y(n_1097)
);

INVx1_ASAP7_75t_L g1098 ( 
.A(n_965),
.Y(n_1098)
);

INVx1_ASAP7_75t_L g1099 ( 
.A(n_942),
.Y(n_1099)
);

AND2x2_ASAP7_75t_L g1100 ( 
.A(n_980),
.B(n_658),
.Y(n_1100)
);

INVx1_ASAP7_75t_L g1101 ( 
.A(n_942),
.Y(n_1101)
);

OR2x6_ASAP7_75t_L g1102 ( 
.A(n_973),
.B(n_0),
.Y(n_1102)
);

INVx1_ASAP7_75t_L g1103 ( 
.A(n_945),
.Y(n_1103)
);

INVx1_ASAP7_75t_L g1104 ( 
.A(n_945),
.Y(n_1104)
);

NAND2xp5_ASAP7_75t_L g1105 ( 
.A(n_962),
.B(n_918),
.Y(n_1105)
);

NAND2xp5_ASAP7_75t_L g1106 ( 
.A(n_981),
.B(n_660),
.Y(n_1106)
);

AND2x4_ASAP7_75t_L g1107 ( 
.A(n_998),
.B(n_663),
.Y(n_1107)
);

INVx2_ASAP7_75t_SL g1108 ( 
.A(n_940),
.Y(n_1108)
);

INVx1_ASAP7_75t_L g1109 ( 
.A(n_949),
.Y(n_1109)
);

INVx1_ASAP7_75t_L g1110 ( 
.A(n_946),
.Y(n_1110)
);

INVx1_ASAP7_75t_L g1111 ( 
.A(n_947),
.Y(n_1111)
);

INVx1_ASAP7_75t_L g1112 ( 
.A(n_1011),
.Y(n_1112)
);

NOR2xp33_ASAP7_75t_L g1113 ( 
.A(n_948),
.B(n_665),
.Y(n_1113)
);

XOR2xp5_ASAP7_75t_L g1114 ( 
.A(n_1027),
.B(n_667),
.Y(n_1114)
);

INVx1_ASAP7_75t_L g1115 ( 
.A(n_956),
.Y(n_1115)
);

INVx2_ASAP7_75t_L g1116 ( 
.A(n_956),
.Y(n_1116)
);

NOR2xp33_ASAP7_75t_L g1117 ( 
.A(n_1009),
.B(n_672),
.Y(n_1117)
);

INVx1_ASAP7_75t_L g1118 ( 
.A(n_956),
.Y(n_1118)
);

INVx1_ASAP7_75t_L g1119 ( 
.A(n_963),
.Y(n_1119)
);

INVx1_ASAP7_75t_L g1120 ( 
.A(n_963),
.Y(n_1120)
);

AND2x2_ASAP7_75t_L g1121 ( 
.A(n_963),
.B(n_673),
.Y(n_1121)
);

INVx1_ASAP7_75t_L g1122 ( 
.A(n_1014),
.Y(n_1122)
);

XOR2xp5_ASAP7_75t_L g1123 ( 
.A(n_1010),
.B(n_678),
.Y(n_1123)
);

CKINVDCx20_ASAP7_75t_R g1124 ( 
.A(n_1026),
.Y(n_1124)
);

INVx1_ASAP7_75t_L g1125 ( 
.A(n_1014),
.Y(n_1125)
);

INVx1_ASAP7_75t_L g1126 ( 
.A(n_1014),
.Y(n_1126)
);

OR2x6_ASAP7_75t_L g1127 ( 
.A(n_1033),
.B(n_981),
.Y(n_1127)
);

AOI22xp5_ASAP7_75t_L g1128 ( 
.A1(n_1063),
.A2(n_1020),
.B1(n_990),
.B2(n_1016),
.Y(n_1128)
);

INVx2_ASAP7_75t_L g1129 ( 
.A(n_1038),
.Y(n_1129)
);

NAND2x1_ASAP7_75t_L g1130 ( 
.A(n_1048),
.B(n_1014),
.Y(n_1130)
);

BUFx12f_ASAP7_75t_L g1131 ( 
.A(n_1102),
.Y(n_1131)
);

INVx8_ASAP7_75t_L g1132 ( 
.A(n_1073),
.Y(n_1132)
);

NAND2xp5_ASAP7_75t_L g1133 ( 
.A(n_1076),
.B(n_999),
.Y(n_1133)
);

NOR2xp33_ASAP7_75t_L g1134 ( 
.A(n_1035),
.B(n_1089),
.Y(n_1134)
);

NAND2xp5_ASAP7_75t_L g1135 ( 
.A(n_1069),
.B(n_999),
.Y(n_1135)
);

AOI22xp33_ASAP7_75t_L g1136 ( 
.A1(n_1081),
.A2(n_999),
.B1(n_1008),
.B2(n_1019),
.Y(n_1136)
);

NAND2xp5_ASAP7_75t_L g1137 ( 
.A(n_1029),
.B(n_999),
.Y(n_1137)
);

INVx2_ASAP7_75t_L g1138 ( 
.A(n_1058),
.Y(n_1138)
);

NAND2xp5_ASAP7_75t_L g1139 ( 
.A(n_1031),
.B(n_680),
.Y(n_1139)
);

OR2x6_ASAP7_75t_L g1140 ( 
.A(n_1102),
.B(n_1007),
.Y(n_1140)
);

AO22x1_ASAP7_75t_L g1141 ( 
.A1(n_1117),
.A2(n_684),
.B1(n_687),
.B2(n_681),
.Y(n_1141)
);

NAND2xp5_ASAP7_75t_L g1142 ( 
.A(n_1034),
.B(n_688),
.Y(n_1142)
);

INVx2_ASAP7_75t_L g1143 ( 
.A(n_1088),
.Y(n_1143)
);

NOR3xp33_ASAP7_75t_L g1144 ( 
.A(n_1057),
.B(n_741),
.C(n_738),
.Y(n_1144)
);

INVx2_ASAP7_75t_SL g1145 ( 
.A(n_1036),
.Y(n_1145)
);

INVx1_ASAP7_75t_L g1146 ( 
.A(n_1037),
.Y(n_1146)
);

INVx2_ASAP7_75t_L g1147 ( 
.A(n_1096),
.Y(n_1147)
);

INVx1_ASAP7_75t_L g1148 ( 
.A(n_1039),
.Y(n_1148)
);

BUFx3_ASAP7_75t_L g1149 ( 
.A(n_1028),
.Y(n_1149)
);

NAND2xp5_ASAP7_75t_L g1150 ( 
.A(n_1040),
.B(n_690),
.Y(n_1150)
);

INVx1_ASAP7_75t_L g1151 ( 
.A(n_1077),
.Y(n_1151)
);

NOR3xp33_ASAP7_75t_SL g1152 ( 
.A(n_1062),
.B(n_1079),
.C(n_1059),
.Y(n_1152)
);

NAND2xp5_ASAP7_75t_L g1153 ( 
.A(n_1065),
.B(n_691),
.Y(n_1153)
);

NAND2xp5_ASAP7_75t_L g1154 ( 
.A(n_1085),
.B(n_692),
.Y(n_1154)
);

NAND2xp5_ASAP7_75t_SL g1155 ( 
.A(n_1030),
.B(n_695),
.Y(n_1155)
);

AND2x4_ASAP7_75t_SL g1156 ( 
.A(n_1032),
.B(n_997),
.Y(n_1156)
);

INVx1_ASAP7_75t_L g1157 ( 
.A(n_1078),
.Y(n_1157)
);

NAND2xp5_ASAP7_75t_L g1158 ( 
.A(n_1041),
.B(n_700),
.Y(n_1158)
);

NAND2xp5_ASAP7_75t_SL g1159 ( 
.A(n_1113),
.B(n_704),
.Y(n_1159)
);

INVx1_ASAP7_75t_L g1160 ( 
.A(n_1080),
.Y(n_1160)
);

NOR3xp33_ASAP7_75t_L g1161 ( 
.A(n_1100),
.B(n_717),
.C(n_711),
.Y(n_1161)
);

INVx4_ASAP7_75t_L g1162 ( 
.A(n_1073),
.Y(n_1162)
);

AOI22xp5_ASAP7_75t_L g1163 ( 
.A1(n_1042),
.A2(n_719),
.B1(n_721),
.B2(n_718),
.Y(n_1163)
);

NAND2xp5_ASAP7_75t_SL g1164 ( 
.A(n_1045),
.B(n_725),
.Y(n_1164)
);

BUFx2_ASAP7_75t_L g1165 ( 
.A(n_1043),
.Y(n_1165)
);

INVx1_ASAP7_75t_L g1166 ( 
.A(n_1082),
.Y(n_1166)
);

AOI22xp5_ASAP7_75t_L g1167 ( 
.A1(n_1046),
.A2(n_727),
.B1(n_728),
.B2(n_726),
.Y(n_1167)
);

AND2x2_ASAP7_75t_L g1168 ( 
.A(n_1044),
.B(n_729),
.Y(n_1168)
);

NAND2xp5_ASAP7_75t_L g1169 ( 
.A(n_1047),
.B(n_737),
.Y(n_1169)
);

AOI22xp33_ASAP7_75t_L g1170 ( 
.A1(n_1048),
.A2(n_743),
.B1(n_742),
.B2(n_997),
.Y(n_1170)
);

INVx1_ASAP7_75t_L g1171 ( 
.A(n_1087),
.Y(n_1171)
);

NAND2xp5_ASAP7_75t_L g1172 ( 
.A(n_1050),
.B(n_1018),
.Y(n_1172)
);

NAND2xp5_ASAP7_75t_L g1173 ( 
.A(n_1052),
.B(n_1018),
.Y(n_1173)
);

INVx2_ASAP7_75t_L g1174 ( 
.A(n_1055),
.Y(n_1174)
);

NAND2xp5_ASAP7_75t_L g1175 ( 
.A(n_1099),
.B(n_1025),
.Y(n_1175)
);

NAND2xp5_ASAP7_75t_L g1176 ( 
.A(n_1101),
.B(n_1025),
.Y(n_1176)
);

NAND2xp5_ASAP7_75t_L g1177 ( 
.A(n_1103),
.B(n_856),
.Y(n_1177)
);

INVxp67_ASAP7_75t_L g1178 ( 
.A(n_1056),
.Y(n_1178)
);

NAND2x1_ASAP7_75t_L g1179 ( 
.A(n_1048),
.B(n_116),
.Y(n_1179)
);

NOR3x1_ASAP7_75t_L g1180 ( 
.A(n_1093),
.B(n_1),
.C(n_2),
.Y(n_1180)
);

INVxp67_ASAP7_75t_L g1181 ( 
.A(n_1060),
.Y(n_1181)
);

INVx1_ASAP7_75t_L g1182 ( 
.A(n_1061),
.Y(n_1182)
);

BUFx8_ASAP7_75t_L g1183 ( 
.A(n_1051),
.Y(n_1183)
);

INVx8_ASAP7_75t_L g1184 ( 
.A(n_1044),
.Y(n_1184)
);

AND2x2_ASAP7_75t_L g1185 ( 
.A(n_1123),
.B(n_3),
.Y(n_1185)
);

INVx1_ASAP7_75t_L g1186 ( 
.A(n_1066),
.Y(n_1186)
);

NAND2xp5_ASAP7_75t_L g1187 ( 
.A(n_1104),
.B(n_856),
.Y(n_1187)
);

AND2x4_ASAP7_75t_L g1188 ( 
.A(n_1054),
.B(n_117),
.Y(n_1188)
);

NOR2x2_ASAP7_75t_L g1189 ( 
.A(n_1067),
.B(n_3),
.Y(n_1189)
);

AND2x4_ASAP7_75t_L g1190 ( 
.A(n_1053),
.B(n_1091),
.Y(n_1190)
);

NAND2xp5_ASAP7_75t_L g1191 ( 
.A(n_1068),
.B(n_856),
.Y(n_1191)
);

NOR2xp33_ASAP7_75t_L g1192 ( 
.A(n_1114),
.B(n_5),
.Y(n_1192)
);

INVx2_ASAP7_75t_SL g1193 ( 
.A(n_1064),
.Y(n_1193)
);

INVx1_ASAP7_75t_L g1194 ( 
.A(n_1070),
.Y(n_1194)
);

NAND2xp5_ASAP7_75t_L g1195 ( 
.A(n_1071),
.B(n_6),
.Y(n_1195)
);

A2O1A1Ixp33_ASAP7_75t_L g1196 ( 
.A1(n_1084),
.A2(n_8),
.B(n_6),
.C(n_7),
.Y(n_1196)
);

NAND2xp5_ASAP7_75t_SL g1197 ( 
.A(n_1053),
.B(n_118),
.Y(n_1197)
);

INVx2_ASAP7_75t_L g1198 ( 
.A(n_1072),
.Y(n_1198)
);

AND2x6_ASAP7_75t_SL g1199 ( 
.A(n_1064),
.B(n_8),
.Y(n_1199)
);

NOR2xp67_ASAP7_75t_L g1200 ( 
.A(n_1094),
.B(n_119),
.Y(n_1200)
);

INVx2_ASAP7_75t_SL g1201 ( 
.A(n_1090),
.Y(n_1201)
);

INVx2_ASAP7_75t_L g1202 ( 
.A(n_1074),
.Y(n_1202)
);

INVx2_ASAP7_75t_L g1203 ( 
.A(n_1075),
.Y(n_1203)
);

OAI21xp5_ASAP7_75t_L g1204 ( 
.A1(n_1083),
.A2(n_123),
.B(n_120),
.Y(n_1204)
);

AO22x1_ASAP7_75t_L g1205 ( 
.A1(n_1090),
.A2(n_12),
.B1(n_9),
.B2(n_10),
.Y(n_1205)
);

AOI22xp33_ASAP7_75t_L g1206 ( 
.A1(n_1092),
.A2(n_12),
.B1(n_9),
.B2(n_10),
.Y(n_1206)
);

INVx1_ASAP7_75t_L g1207 ( 
.A(n_1146),
.Y(n_1207)
);

INVx4_ASAP7_75t_L g1208 ( 
.A(n_1132),
.Y(n_1208)
);

BUFx3_ASAP7_75t_L g1209 ( 
.A(n_1183),
.Y(n_1209)
);

INVx1_ASAP7_75t_L g1210 ( 
.A(n_1147),
.Y(n_1210)
);

NAND2xp5_ASAP7_75t_L g1211 ( 
.A(n_1134),
.B(n_1098),
.Y(n_1211)
);

INVx2_ASAP7_75t_L g1212 ( 
.A(n_1174),
.Y(n_1212)
);

BUFx6f_ASAP7_75t_L g1213 ( 
.A(n_1132),
.Y(n_1213)
);

NAND2xp5_ASAP7_75t_L g1214 ( 
.A(n_1148),
.B(n_1121),
.Y(n_1214)
);

OR2x2_ASAP7_75t_L g1215 ( 
.A(n_1165),
.B(n_1107),
.Y(n_1215)
);

INVx1_ASAP7_75t_L g1216 ( 
.A(n_1151),
.Y(n_1216)
);

INVx2_ASAP7_75t_L g1217 ( 
.A(n_1157),
.Y(n_1217)
);

A2O1A1Ixp33_ASAP7_75t_L g1218 ( 
.A1(n_1128),
.A2(n_1109),
.B(n_1086),
.C(n_1110),
.Y(n_1218)
);

NAND2xp5_ASAP7_75t_L g1219 ( 
.A(n_1145),
.B(n_1049),
.Y(n_1219)
);

NAND2xp5_ASAP7_75t_L g1220 ( 
.A(n_1160),
.B(n_1108),
.Y(n_1220)
);

INVx1_ASAP7_75t_SL g1221 ( 
.A(n_1156),
.Y(n_1221)
);

BUFx6f_ASAP7_75t_L g1222 ( 
.A(n_1149),
.Y(n_1222)
);

INVx2_ASAP7_75t_L g1223 ( 
.A(n_1166),
.Y(n_1223)
);

NAND2xp5_ASAP7_75t_L g1224 ( 
.A(n_1171),
.B(n_1107),
.Y(n_1224)
);

HB1xp67_ASAP7_75t_L g1225 ( 
.A(n_1190),
.Y(n_1225)
);

AOI22xp33_ASAP7_75t_L g1226 ( 
.A1(n_1161),
.A2(n_1111),
.B1(n_1112),
.B2(n_1116),
.Y(n_1226)
);

INVx1_ASAP7_75t_L g1227 ( 
.A(n_1182),
.Y(n_1227)
);

NAND2xp5_ASAP7_75t_L g1228 ( 
.A(n_1153),
.B(n_1106),
.Y(n_1228)
);

INVxp67_ASAP7_75t_L g1229 ( 
.A(n_1140),
.Y(n_1229)
);

HB1xp67_ASAP7_75t_L g1230 ( 
.A(n_1190),
.Y(n_1230)
);

A2O1A1Ixp33_ASAP7_75t_L g1231 ( 
.A1(n_1135),
.A2(n_1125),
.B(n_1126),
.C(n_1122),
.Y(n_1231)
);

INVx2_ASAP7_75t_L g1232 ( 
.A(n_1129),
.Y(n_1232)
);

INVx4_ASAP7_75t_L g1233 ( 
.A(n_1184),
.Y(n_1233)
);

INVx2_ASAP7_75t_L g1234 ( 
.A(n_1138),
.Y(n_1234)
);

NOR3xp33_ASAP7_75t_SL g1235 ( 
.A(n_1192),
.B(n_1095),
.C(n_1155),
.Y(n_1235)
);

INVx2_ASAP7_75t_L g1236 ( 
.A(n_1143),
.Y(n_1236)
);

OR2x2_ASAP7_75t_SL g1237 ( 
.A(n_1189),
.B(n_1124),
.Y(n_1237)
);

HB1xp67_ASAP7_75t_L g1238 ( 
.A(n_1127),
.Y(n_1238)
);

INVx1_ASAP7_75t_SL g1239 ( 
.A(n_1168),
.Y(n_1239)
);

CKINVDCx5p33_ASAP7_75t_R g1240 ( 
.A(n_1183),
.Y(n_1240)
);

INVx1_ASAP7_75t_L g1241 ( 
.A(n_1186),
.Y(n_1241)
);

INVx4_ASAP7_75t_L g1242 ( 
.A(n_1184),
.Y(n_1242)
);

BUFx2_ASAP7_75t_L g1243 ( 
.A(n_1127),
.Y(n_1243)
);

AND2x2_ASAP7_75t_L g1244 ( 
.A(n_1193),
.B(n_1051),
.Y(n_1244)
);

INVx2_ASAP7_75t_L g1245 ( 
.A(n_1198),
.Y(n_1245)
);

NAND2xp5_ASAP7_75t_L g1246 ( 
.A(n_1194),
.B(n_1115),
.Y(n_1246)
);

BUFx2_ASAP7_75t_L g1247 ( 
.A(n_1162),
.Y(n_1247)
);

INVx2_ASAP7_75t_L g1248 ( 
.A(n_1202),
.Y(n_1248)
);

BUFx6f_ASAP7_75t_L g1249 ( 
.A(n_1188),
.Y(n_1249)
);

BUFx3_ASAP7_75t_L g1250 ( 
.A(n_1131),
.Y(n_1250)
);

INVx1_ASAP7_75t_L g1251 ( 
.A(n_1203),
.Y(n_1251)
);

AOI22xp5_ASAP7_75t_L g1252 ( 
.A1(n_1201),
.A2(n_1118),
.B1(n_1120),
.B2(n_1119),
.Y(n_1252)
);

AND2x2_ASAP7_75t_L g1253 ( 
.A(n_1185),
.B(n_1097),
.Y(n_1253)
);

HB1xp67_ASAP7_75t_L g1254 ( 
.A(n_1178),
.Y(n_1254)
);

OAI221xp5_ASAP7_75t_L g1255 ( 
.A1(n_1181),
.A2(n_1105),
.B1(n_15),
.B2(n_13),
.C(n_14),
.Y(n_1255)
);

OR2x2_ASAP7_75t_L g1256 ( 
.A(n_1158),
.B(n_13),
.Y(n_1256)
);

INVxp67_ASAP7_75t_L g1257 ( 
.A(n_1140),
.Y(n_1257)
);

BUFx6f_ASAP7_75t_L g1258 ( 
.A(n_1188),
.Y(n_1258)
);

OAI22xp5_ASAP7_75t_L g1259 ( 
.A1(n_1136),
.A2(n_125),
.B1(n_126),
.B2(n_124),
.Y(n_1259)
);

HB1xp67_ASAP7_75t_L g1260 ( 
.A(n_1195),
.Y(n_1260)
);

AND2x6_ASAP7_75t_L g1261 ( 
.A(n_1180),
.B(n_127),
.Y(n_1261)
);

AND2x2_ASAP7_75t_L g1262 ( 
.A(n_1144),
.B(n_1152),
.Y(n_1262)
);

INVx2_ASAP7_75t_SL g1263 ( 
.A(n_1164),
.Y(n_1263)
);

INVx3_ASAP7_75t_L g1264 ( 
.A(n_1199),
.Y(n_1264)
);

NAND2x1p5_ASAP7_75t_L g1265 ( 
.A(n_1130),
.B(n_128),
.Y(n_1265)
);

NAND2xp5_ASAP7_75t_L g1266 ( 
.A(n_1139),
.B(n_14),
.Y(n_1266)
);

INVx3_ASAP7_75t_L g1267 ( 
.A(n_1179),
.Y(n_1267)
);

OR2x6_ASAP7_75t_L g1268 ( 
.A(n_1205),
.B(n_16),
.Y(n_1268)
);

AND2x2_ASAP7_75t_L g1269 ( 
.A(n_1169),
.B(n_16),
.Y(n_1269)
);

OR2x6_ASAP7_75t_L g1270 ( 
.A(n_1197),
.B(n_17),
.Y(n_1270)
);

NAND2xp5_ASAP7_75t_L g1271 ( 
.A(n_1142),
.B(n_17),
.Y(n_1271)
);

AND2x2_ASAP7_75t_L g1272 ( 
.A(n_1150),
.B(n_19),
.Y(n_1272)
);

BUFx6f_ASAP7_75t_L g1273 ( 
.A(n_1191),
.Y(n_1273)
);

NOR2xp33_ASAP7_75t_L g1274 ( 
.A(n_1159),
.B(n_19),
.Y(n_1274)
);

BUFx4f_ASAP7_75t_L g1275 ( 
.A(n_1206),
.Y(n_1275)
);

AO221x1_ASAP7_75t_L g1276 ( 
.A1(n_1196),
.A2(n_22),
.B1(n_20),
.B2(n_21),
.C(n_23),
.Y(n_1276)
);

INVx1_ASAP7_75t_L g1277 ( 
.A(n_1175),
.Y(n_1277)
);

INVx1_ASAP7_75t_L g1278 ( 
.A(n_1176),
.Y(n_1278)
);

NAND2xp5_ASAP7_75t_L g1279 ( 
.A(n_1172),
.B(n_21),
.Y(n_1279)
);

INVxp67_ASAP7_75t_L g1280 ( 
.A(n_1173),
.Y(n_1280)
);

NAND2xp5_ASAP7_75t_L g1281 ( 
.A(n_1141),
.B(n_22),
.Y(n_1281)
);

NAND2xp5_ASAP7_75t_L g1282 ( 
.A(n_1137),
.B(n_23),
.Y(n_1282)
);

INVx1_ASAP7_75t_L g1283 ( 
.A(n_1177),
.Y(n_1283)
);

OAI21x1_ASAP7_75t_L g1284 ( 
.A1(n_1267),
.A2(n_1204),
.B(n_1133),
.Y(n_1284)
);

NOR2xp33_ASAP7_75t_L g1285 ( 
.A(n_1211),
.B(n_1163),
.Y(n_1285)
);

OR2x2_ASAP7_75t_L g1286 ( 
.A(n_1215),
.B(n_1167),
.Y(n_1286)
);

AOI21x1_ASAP7_75t_L g1287 ( 
.A1(n_1282),
.A2(n_1154),
.B(n_1187),
.Y(n_1287)
);

INVx2_ASAP7_75t_L g1288 ( 
.A(n_1217),
.Y(n_1288)
);

OAI21x1_ASAP7_75t_SL g1289 ( 
.A1(n_1259),
.A2(n_1170),
.B(n_1200),
.Y(n_1289)
);

NAND2xp5_ASAP7_75t_SL g1290 ( 
.A(n_1275),
.B(n_24),
.Y(n_1290)
);

NAND3xp33_ASAP7_75t_L g1291 ( 
.A(n_1274),
.B(n_25),
.C(n_26),
.Y(n_1291)
);

BUFx3_ASAP7_75t_L g1292 ( 
.A(n_1213),
.Y(n_1292)
);

NAND2xp5_ASAP7_75t_L g1293 ( 
.A(n_1260),
.B(n_25),
.Y(n_1293)
);

OAI21x1_ASAP7_75t_L g1294 ( 
.A1(n_1265),
.A2(n_131),
.B(n_130),
.Y(n_1294)
);

AOI221x1_ASAP7_75t_L g1295 ( 
.A1(n_1231),
.A2(n_1218),
.B1(n_1281),
.B2(n_1228),
.C(n_1271),
.Y(n_1295)
);

OAI21x1_ASAP7_75t_L g1296 ( 
.A1(n_1246),
.A2(n_133),
.B(n_132),
.Y(n_1296)
);

AO31x2_ASAP7_75t_L g1297 ( 
.A1(n_1266),
.A2(n_135),
.A3(n_137),
.B(n_134),
.Y(n_1297)
);

INVx1_ASAP7_75t_L g1298 ( 
.A(n_1207),
.Y(n_1298)
);

NAND2x1p5_ASAP7_75t_L g1299 ( 
.A(n_1208),
.B(n_138),
.Y(n_1299)
);

AND2x4_ASAP7_75t_L g1300 ( 
.A(n_1233),
.B(n_570),
.Y(n_1300)
);

NAND2xp5_ASAP7_75t_L g1301 ( 
.A(n_1280),
.B(n_27),
.Y(n_1301)
);

AND2x2_ASAP7_75t_L g1302 ( 
.A(n_1253),
.B(n_1239),
.Y(n_1302)
);

OAI21x1_ASAP7_75t_L g1303 ( 
.A1(n_1210),
.A2(n_142),
.B(n_141),
.Y(n_1303)
);

AOI21x1_ASAP7_75t_SL g1304 ( 
.A1(n_1262),
.A2(n_27),
.B(n_28),
.Y(n_1304)
);

INVx3_ASAP7_75t_L g1305 ( 
.A(n_1213),
.Y(n_1305)
);

AO31x2_ASAP7_75t_L g1306 ( 
.A1(n_1279),
.A2(n_144),
.A3(n_145),
.B(n_143),
.Y(n_1306)
);

OAI21x1_ASAP7_75t_L g1307 ( 
.A1(n_1210),
.A2(n_148),
.B(n_147),
.Y(n_1307)
);

NAND2xp5_ASAP7_75t_L g1308 ( 
.A(n_1277),
.B(n_1278),
.Y(n_1308)
);

A2O1A1Ixp33_ASAP7_75t_L g1309 ( 
.A1(n_1269),
.A2(n_30),
.B(n_28),
.C(n_29),
.Y(n_1309)
);

BUFx3_ASAP7_75t_L g1310 ( 
.A(n_1222),
.Y(n_1310)
);

NAND2xp5_ASAP7_75t_L g1311 ( 
.A(n_1214),
.B(n_29),
.Y(n_1311)
);

OAI21x1_ASAP7_75t_L g1312 ( 
.A1(n_1226),
.A2(n_151),
.B(n_150),
.Y(n_1312)
);

INVx3_ASAP7_75t_L g1313 ( 
.A(n_1242),
.Y(n_1313)
);

NAND2xp5_ASAP7_75t_SL g1314 ( 
.A(n_1249),
.B(n_30),
.Y(n_1314)
);

AOI21x1_ASAP7_75t_SL g1315 ( 
.A1(n_1272),
.A2(n_31),
.B(n_32),
.Y(n_1315)
);

OAI21xp5_ASAP7_75t_L g1316 ( 
.A1(n_1224),
.A2(n_154),
.B(n_153),
.Y(n_1316)
);

OAI21xp5_ASAP7_75t_L g1317 ( 
.A1(n_1283),
.A2(n_156),
.B(n_155),
.Y(n_1317)
);

INVx2_ASAP7_75t_SL g1318 ( 
.A(n_1222),
.Y(n_1318)
);

AO21x1_ASAP7_75t_L g1319 ( 
.A1(n_1256),
.A2(n_31),
.B(n_32),
.Y(n_1319)
);

OAI21x1_ASAP7_75t_L g1320 ( 
.A1(n_1251),
.A2(n_158),
.B(n_157),
.Y(n_1320)
);

CKINVDCx20_ASAP7_75t_R g1321 ( 
.A(n_1237),
.Y(n_1321)
);

O2A1O1Ixp5_ASAP7_75t_L g1322 ( 
.A1(n_1227),
.A2(n_35),
.B(n_33),
.C(n_34),
.Y(n_1322)
);

AOI21xp5_ASAP7_75t_SL g1323 ( 
.A1(n_1249),
.A2(n_161),
.B(n_159),
.Y(n_1323)
);

OAI21x1_ASAP7_75t_L g1324 ( 
.A1(n_1232),
.A2(n_163),
.B(n_162),
.Y(n_1324)
);

INVx2_ASAP7_75t_L g1325 ( 
.A(n_1223),
.Y(n_1325)
);

BUFx6f_ASAP7_75t_L g1326 ( 
.A(n_1247),
.Y(n_1326)
);

INVx4_ASAP7_75t_L g1327 ( 
.A(n_1247),
.Y(n_1327)
);

BUFx2_ASAP7_75t_L g1328 ( 
.A(n_1225),
.Y(n_1328)
);

OAI21x1_ASAP7_75t_L g1329 ( 
.A1(n_1234),
.A2(n_165),
.B(n_164),
.Y(n_1329)
);

NAND2xp5_ASAP7_75t_L g1330 ( 
.A(n_1216),
.B(n_33),
.Y(n_1330)
);

OR2x2_ASAP7_75t_L g1331 ( 
.A(n_1230),
.B(n_34),
.Y(n_1331)
);

AND2x6_ASAP7_75t_L g1332 ( 
.A(n_1258),
.B(n_166),
.Y(n_1332)
);

AOI21xp5_ASAP7_75t_L g1333 ( 
.A1(n_1263),
.A2(n_170),
.B(n_169),
.Y(n_1333)
);

INVx1_ASAP7_75t_L g1334 ( 
.A(n_1241),
.Y(n_1334)
);

OAI21x1_ASAP7_75t_L g1335 ( 
.A1(n_1236),
.A2(n_1248),
.B(n_1245),
.Y(n_1335)
);

AOI21x1_ASAP7_75t_L g1336 ( 
.A1(n_1220),
.A2(n_174),
.B(n_171),
.Y(n_1336)
);

NOR2x1_ASAP7_75t_SL g1337 ( 
.A(n_1270),
.B(n_1258),
.Y(n_1337)
);

OAI21xp5_ASAP7_75t_L g1338 ( 
.A1(n_1212),
.A2(n_177),
.B(n_176),
.Y(n_1338)
);

NAND2xp5_ASAP7_75t_SL g1339 ( 
.A(n_1254),
.B(n_35),
.Y(n_1339)
);

INVx1_ASAP7_75t_L g1340 ( 
.A(n_1219),
.Y(n_1340)
);

INVxp67_ASAP7_75t_SL g1341 ( 
.A(n_1238),
.Y(n_1341)
);

NAND2xp5_ASAP7_75t_L g1342 ( 
.A(n_1270),
.B(n_36),
.Y(n_1342)
);

OAI21x1_ASAP7_75t_L g1343 ( 
.A1(n_1252),
.A2(n_179),
.B(n_178),
.Y(n_1343)
);

NAND2xp5_ASAP7_75t_L g1344 ( 
.A(n_1273),
.B(n_36),
.Y(n_1344)
);

INVx2_ASAP7_75t_SL g1345 ( 
.A(n_1244),
.Y(n_1345)
);

AOI21xp5_ASAP7_75t_L g1346 ( 
.A1(n_1243),
.A2(n_183),
.B(n_182),
.Y(n_1346)
);

INVx2_ASAP7_75t_L g1347 ( 
.A(n_1273),
.Y(n_1347)
);

INVx2_ASAP7_75t_L g1348 ( 
.A(n_1276),
.Y(n_1348)
);

A2O1A1Ixp33_ASAP7_75t_L g1349 ( 
.A1(n_1235),
.A2(n_1255),
.B(n_1243),
.C(n_1229),
.Y(n_1349)
);

NAND2xp5_ASAP7_75t_L g1350 ( 
.A(n_1261),
.B(n_37),
.Y(n_1350)
);

INVx1_ASAP7_75t_L g1351 ( 
.A(n_1276),
.Y(n_1351)
);

AO31x2_ASAP7_75t_L g1352 ( 
.A1(n_1261),
.A2(n_1268),
.A3(n_186),
.B(n_187),
.Y(n_1352)
);

INVx1_ASAP7_75t_L g1353 ( 
.A(n_1268),
.Y(n_1353)
);

AOI21xp5_ASAP7_75t_L g1354 ( 
.A1(n_1221),
.A2(n_188),
.B(n_184),
.Y(n_1354)
);

OAI21xp5_ASAP7_75t_L g1355 ( 
.A1(n_1261),
.A2(n_190),
.B(n_189),
.Y(n_1355)
);

NOR2xp33_ASAP7_75t_L g1356 ( 
.A(n_1257),
.B(n_37),
.Y(n_1356)
);

OAI21x1_ASAP7_75t_SL g1357 ( 
.A1(n_1209),
.A2(n_192),
.B(n_191),
.Y(n_1357)
);

AOI21xp5_ASAP7_75t_L g1358 ( 
.A1(n_1250),
.A2(n_194),
.B(n_193),
.Y(n_1358)
);

AOI21x1_ASAP7_75t_L g1359 ( 
.A1(n_1264),
.A2(n_568),
.B(n_196),
.Y(n_1359)
);

OAI22xp5_ASAP7_75t_L g1360 ( 
.A1(n_1240),
.A2(n_40),
.B1(n_38),
.B2(n_39),
.Y(n_1360)
);

A2O1A1Ixp33_ASAP7_75t_L g1361 ( 
.A1(n_1285),
.A2(n_40),
.B(n_38),
.C(n_39),
.Y(n_1361)
);

BUFx10_ASAP7_75t_L g1362 ( 
.A(n_1326),
.Y(n_1362)
);

OAI21x1_ASAP7_75t_L g1363 ( 
.A1(n_1284),
.A2(n_197),
.B(n_195),
.Y(n_1363)
);

INVx1_ASAP7_75t_SL g1364 ( 
.A(n_1302),
.Y(n_1364)
);

AO31x2_ASAP7_75t_L g1365 ( 
.A1(n_1295),
.A2(n_199),
.A3(n_201),
.B(n_198),
.Y(n_1365)
);

INVx2_ASAP7_75t_L g1366 ( 
.A(n_1288),
.Y(n_1366)
);

AOI21xp5_ASAP7_75t_L g1367 ( 
.A1(n_1289),
.A2(n_567),
.B(n_204),
.Y(n_1367)
);

OAI21x1_ASAP7_75t_SL g1368 ( 
.A1(n_1355),
.A2(n_41),
.B(n_42),
.Y(n_1368)
);

OAI21xp5_ASAP7_75t_L g1369 ( 
.A1(n_1349),
.A2(n_41),
.B(n_42),
.Y(n_1369)
);

INVx2_ASAP7_75t_L g1370 ( 
.A(n_1325),
.Y(n_1370)
);

NAND2xp5_ASAP7_75t_L g1371 ( 
.A(n_1308),
.B(n_43),
.Y(n_1371)
);

AOI21xp5_ASAP7_75t_L g1372 ( 
.A1(n_1289),
.A2(n_566),
.B(n_205),
.Y(n_1372)
);

BUFx6f_ASAP7_75t_L g1373 ( 
.A(n_1310),
.Y(n_1373)
);

OAI21x1_ASAP7_75t_L g1374 ( 
.A1(n_1324),
.A2(n_206),
.B(n_202),
.Y(n_1374)
);

AO31x2_ASAP7_75t_L g1375 ( 
.A1(n_1351),
.A2(n_208),
.A3(n_209),
.B(n_207),
.Y(n_1375)
);

BUFx6f_ASAP7_75t_L g1376 ( 
.A(n_1326),
.Y(n_1376)
);

OAI21x1_ASAP7_75t_L g1377 ( 
.A1(n_1329),
.A2(n_212),
.B(n_210),
.Y(n_1377)
);

O2A1O1Ixp5_ASAP7_75t_L g1378 ( 
.A1(n_1287),
.A2(n_45),
.B(n_43),
.C(n_44),
.Y(n_1378)
);

AOI21xp5_ASAP7_75t_L g1379 ( 
.A1(n_1338),
.A2(n_1317),
.B(n_1316),
.Y(n_1379)
);

AOI21xp5_ASAP7_75t_L g1380 ( 
.A1(n_1346),
.A2(n_217),
.B(n_213),
.Y(n_1380)
);

INVx5_ASAP7_75t_L g1381 ( 
.A(n_1305),
.Y(n_1381)
);

NAND2xp5_ASAP7_75t_L g1382 ( 
.A(n_1340),
.B(n_1311),
.Y(n_1382)
);

AO31x2_ASAP7_75t_L g1383 ( 
.A1(n_1348),
.A2(n_219),
.A3(n_220),
.B(n_218),
.Y(n_1383)
);

AOI21xp5_ASAP7_75t_L g1384 ( 
.A1(n_1333),
.A2(n_565),
.B(n_227),
.Y(n_1384)
);

AOI21xp5_ASAP7_75t_L g1385 ( 
.A1(n_1312),
.A2(n_564),
.B(n_229),
.Y(n_1385)
);

HB1xp67_ASAP7_75t_L g1386 ( 
.A(n_1328),
.Y(n_1386)
);

INVx1_ASAP7_75t_L g1387 ( 
.A(n_1298),
.Y(n_1387)
);

INVx2_ASAP7_75t_L g1388 ( 
.A(n_1334),
.Y(n_1388)
);

AO21x2_ASAP7_75t_L g1389 ( 
.A1(n_1343),
.A2(n_230),
.B(n_221),
.Y(n_1389)
);

OAI21x1_ASAP7_75t_L g1390 ( 
.A1(n_1303),
.A2(n_233),
.B(n_231),
.Y(n_1390)
);

CKINVDCx20_ASAP7_75t_R g1391 ( 
.A(n_1321),
.Y(n_1391)
);

AOI21xp5_ASAP7_75t_L g1392 ( 
.A1(n_1294),
.A2(n_563),
.B(n_236),
.Y(n_1392)
);

OAI21x1_ASAP7_75t_L g1393 ( 
.A1(n_1307),
.A2(n_237),
.B(n_234),
.Y(n_1393)
);

NAND2xp5_ASAP7_75t_L g1394 ( 
.A(n_1328),
.B(n_1301),
.Y(n_1394)
);

AOI21xp5_ASAP7_75t_SL g1395 ( 
.A1(n_1300),
.A2(n_239),
.B(n_238),
.Y(n_1395)
);

NAND3xp33_ASAP7_75t_SL g1396 ( 
.A(n_1290),
.B(n_44),
.C(n_46),
.Y(n_1396)
);

INVx1_ASAP7_75t_L g1397 ( 
.A(n_1335),
.Y(n_1397)
);

AOI21xp5_ASAP7_75t_L g1398 ( 
.A1(n_1354),
.A2(n_241),
.B(n_240),
.Y(n_1398)
);

INVx2_ASAP7_75t_SL g1399 ( 
.A(n_1292),
.Y(n_1399)
);

AOI21xp5_ASAP7_75t_L g1400 ( 
.A1(n_1320),
.A2(n_243),
.B(n_242),
.Y(n_1400)
);

AND2x4_ASAP7_75t_L g1401 ( 
.A(n_1318),
.B(n_244),
.Y(n_1401)
);

NAND2xp5_ASAP7_75t_L g1402 ( 
.A(n_1293),
.B(n_46),
.Y(n_1402)
);

AOI21xp5_ASAP7_75t_L g1403 ( 
.A1(n_1323),
.A2(n_246),
.B(n_245),
.Y(n_1403)
);

OR2x2_ASAP7_75t_L g1404 ( 
.A(n_1286),
.B(n_47),
.Y(n_1404)
);

OAI21x1_ASAP7_75t_L g1405 ( 
.A1(n_1296),
.A2(n_248),
.B(n_247),
.Y(n_1405)
);

NAND2xp5_ASAP7_75t_L g1406 ( 
.A(n_1337),
.B(n_1347),
.Y(n_1406)
);

NAND3xp33_ASAP7_75t_SL g1407 ( 
.A(n_1319),
.B(n_47),
.C(n_48),
.Y(n_1407)
);

NAND2xp5_ASAP7_75t_SL g1408 ( 
.A(n_1353),
.B(n_48),
.Y(n_1408)
);

OAI21xp5_ASAP7_75t_L g1409 ( 
.A1(n_1291),
.A2(n_49),
.B(n_50),
.Y(n_1409)
);

AO31x2_ASAP7_75t_L g1410 ( 
.A1(n_1309),
.A2(n_254),
.A3(n_255),
.B(n_253),
.Y(n_1410)
);

OAI21x1_ASAP7_75t_L g1411 ( 
.A1(n_1336),
.A2(n_257),
.B(n_256),
.Y(n_1411)
);

OAI22xp5_ASAP7_75t_L g1412 ( 
.A1(n_1341),
.A2(n_51),
.B1(n_49),
.B2(n_50),
.Y(n_1412)
);

OAI22x1_ASAP7_75t_L g1413 ( 
.A1(n_1342),
.A2(n_54),
.B1(n_52),
.B2(n_53),
.Y(n_1413)
);

AOI21xp5_ASAP7_75t_L g1414 ( 
.A1(n_1358),
.A2(n_259),
.B(n_258),
.Y(n_1414)
);

O2A1O1Ixp33_ASAP7_75t_L g1415 ( 
.A1(n_1339),
.A2(n_56),
.B(n_54),
.C(n_55),
.Y(n_1415)
);

OAI22xp5_ASAP7_75t_L g1416 ( 
.A1(n_1327),
.A2(n_57),
.B1(n_55),
.B2(n_56),
.Y(n_1416)
);

O2A1O1Ixp33_ASAP7_75t_SL g1417 ( 
.A1(n_1350),
.A2(n_59),
.B(n_57),
.C(n_58),
.Y(n_1417)
);

INVx1_ASAP7_75t_L g1418 ( 
.A(n_1330),
.Y(n_1418)
);

AOI21xp5_ASAP7_75t_L g1419 ( 
.A1(n_1322),
.A2(n_261),
.B(n_260),
.Y(n_1419)
);

AND2x2_ASAP7_75t_L g1420 ( 
.A(n_1344),
.B(n_58),
.Y(n_1420)
);

INVx1_ASAP7_75t_L g1421 ( 
.A(n_1331),
.Y(n_1421)
);

AO31x2_ASAP7_75t_L g1422 ( 
.A1(n_1304),
.A2(n_265),
.A3(n_266),
.B(n_263),
.Y(n_1422)
);

NAND2xp5_ASAP7_75t_SL g1423 ( 
.A(n_1345),
.B(n_59),
.Y(n_1423)
);

INVx1_ASAP7_75t_L g1424 ( 
.A(n_1297),
.Y(n_1424)
);

NAND2xp5_ASAP7_75t_L g1425 ( 
.A(n_1314),
.B(n_60),
.Y(n_1425)
);

AOI21xp5_ASAP7_75t_L g1426 ( 
.A1(n_1300),
.A2(n_268),
.B(n_267),
.Y(n_1426)
);

INVx1_ASAP7_75t_L g1427 ( 
.A(n_1297),
.Y(n_1427)
);

INVx2_ASAP7_75t_L g1428 ( 
.A(n_1359),
.Y(n_1428)
);

NOR2xp67_ASAP7_75t_L g1429 ( 
.A(n_1313),
.B(n_1356),
.Y(n_1429)
);

OAI21x1_ASAP7_75t_L g1430 ( 
.A1(n_1315),
.A2(n_270),
.B(n_269),
.Y(n_1430)
);

AOI22xp5_ASAP7_75t_L g1431 ( 
.A1(n_1332),
.A2(n_63),
.B1(n_61),
.B2(n_62),
.Y(n_1431)
);

OAI22x1_ASAP7_75t_L g1432 ( 
.A1(n_1299),
.A2(n_65),
.B1(n_62),
.B2(n_64),
.Y(n_1432)
);

AOI211x1_ASAP7_75t_L g1433 ( 
.A1(n_1360),
.A2(n_67),
.B(n_65),
.C(n_66),
.Y(n_1433)
);

OAI21x1_ASAP7_75t_L g1434 ( 
.A1(n_1357),
.A2(n_274),
.B(n_271),
.Y(n_1434)
);

AO31x2_ASAP7_75t_L g1435 ( 
.A1(n_1306),
.A2(n_276),
.A3(n_277),
.B(n_275),
.Y(n_1435)
);

OAI21x1_ASAP7_75t_L g1436 ( 
.A1(n_1306),
.A2(n_1352),
.B(n_1332),
.Y(n_1436)
);

OAI21x1_ASAP7_75t_L g1437 ( 
.A1(n_1352),
.A2(n_284),
.B(n_282),
.Y(n_1437)
);

OAI21x1_ASAP7_75t_L g1438 ( 
.A1(n_1332),
.A2(n_286),
.B(n_285),
.Y(n_1438)
);

INVx5_ASAP7_75t_L g1439 ( 
.A(n_1326),
.Y(n_1439)
);

AOI21xp5_ASAP7_75t_L g1440 ( 
.A1(n_1289),
.A2(n_295),
.B(n_291),
.Y(n_1440)
);

AOI22xp33_ASAP7_75t_L g1441 ( 
.A1(n_1285),
.A2(n_68),
.B1(n_66),
.B2(n_67),
.Y(n_1441)
);

AND2x2_ASAP7_75t_L g1442 ( 
.A(n_1302),
.B(n_69),
.Y(n_1442)
);

INVx1_ASAP7_75t_SL g1443 ( 
.A(n_1302),
.Y(n_1443)
);

OAI21x1_ASAP7_75t_L g1444 ( 
.A1(n_1284),
.A2(n_298),
.B(n_297),
.Y(n_1444)
);

OAI21x1_ASAP7_75t_L g1445 ( 
.A1(n_1284),
.A2(n_300),
.B(n_299),
.Y(n_1445)
);

OR2x2_ASAP7_75t_L g1446 ( 
.A(n_1302),
.B(n_69),
.Y(n_1446)
);

A2O1A1Ixp33_ASAP7_75t_L g1447 ( 
.A1(n_1285),
.A2(n_72),
.B(n_70),
.C(n_71),
.Y(n_1447)
);

AOI21xp5_ASAP7_75t_L g1448 ( 
.A1(n_1289),
.A2(n_304),
.B(n_303),
.Y(n_1448)
);

INVx1_ASAP7_75t_L g1449 ( 
.A(n_1298),
.Y(n_1449)
);

INVx3_ASAP7_75t_L g1450 ( 
.A(n_1326),
.Y(n_1450)
);

AOI21xp5_ASAP7_75t_L g1451 ( 
.A1(n_1289),
.A2(n_307),
.B(n_306),
.Y(n_1451)
);

OAI21x1_ASAP7_75t_L g1452 ( 
.A1(n_1284),
.A2(n_309),
.B(n_308),
.Y(n_1452)
);

INVx3_ASAP7_75t_L g1453 ( 
.A(n_1326),
.Y(n_1453)
);

INVx2_ASAP7_75t_L g1454 ( 
.A(n_1288),
.Y(n_1454)
);

OAI21x1_ASAP7_75t_L g1455 ( 
.A1(n_1284),
.A2(n_311),
.B(n_310),
.Y(n_1455)
);

INVx1_ASAP7_75t_L g1456 ( 
.A(n_1387),
.Y(n_1456)
);

INVx1_ASAP7_75t_L g1457 ( 
.A(n_1449),
.Y(n_1457)
);

INVx1_ASAP7_75t_L g1458 ( 
.A(n_1388),
.Y(n_1458)
);

BUFx8_ASAP7_75t_L g1459 ( 
.A(n_1373),
.Y(n_1459)
);

OAI22xp33_ASAP7_75t_L g1460 ( 
.A1(n_1431),
.A2(n_72),
.B1(n_70),
.B2(n_71),
.Y(n_1460)
);

BUFx2_ASAP7_75t_L g1461 ( 
.A(n_1386),
.Y(n_1461)
);

OAI22xp33_ASAP7_75t_L g1462 ( 
.A1(n_1369),
.A2(n_1409),
.B1(n_1396),
.B2(n_1379),
.Y(n_1462)
);

AND2x2_ASAP7_75t_L g1463 ( 
.A(n_1364),
.B(n_312),
.Y(n_1463)
);

AOI22xp33_ASAP7_75t_L g1464 ( 
.A1(n_1368),
.A2(n_75),
.B1(n_73),
.B2(n_74),
.Y(n_1464)
);

INVx6_ASAP7_75t_L g1465 ( 
.A(n_1439),
.Y(n_1465)
);

BUFx2_ASAP7_75t_L g1466 ( 
.A(n_1450),
.Y(n_1466)
);

NAND2xp5_ASAP7_75t_L g1467 ( 
.A(n_1382),
.B(n_73),
.Y(n_1467)
);

HB1xp67_ASAP7_75t_L g1468 ( 
.A(n_1394),
.Y(n_1468)
);

OAI22xp5_ASAP7_75t_L g1469 ( 
.A1(n_1418),
.A2(n_77),
.B1(n_75),
.B2(n_76),
.Y(n_1469)
);

CKINVDCx16_ASAP7_75t_R g1470 ( 
.A(n_1391),
.Y(n_1470)
);

INVx2_ASAP7_75t_L g1471 ( 
.A(n_1366),
.Y(n_1471)
);

AOI22xp33_ASAP7_75t_SL g1472 ( 
.A1(n_1412),
.A2(n_79),
.B1(n_77),
.B2(n_78),
.Y(n_1472)
);

INVx2_ASAP7_75t_L g1473 ( 
.A(n_1370),
.Y(n_1473)
);

INVx2_ASAP7_75t_L g1474 ( 
.A(n_1454),
.Y(n_1474)
);

OAI22xp33_ASAP7_75t_L g1475 ( 
.A1(n_1413),
.A2(n_80),
.B1(n_78),
.B2(n_79),
.Y(n_1475)
);

INVx8_ASAP7_75t_L g1476 ( 
.A(n_1439),
.Y(n_1476)
);

INVx4_ASAP7_75t_SL g1477 ( 
.A(n_1373),
.Y(n_1477)
);

INVx1_ASAP7_75t_L g1478 ( 
.A(n_1424),
.Y(n_1478)
);

HB1xp67_ASAP7_75t_L g1479 ( 
.A(n_1443),
.Y(n_1479)
);

AOI22xp33_ASAP7_75t_L g1480 ( 
.A1(n_1407),
.A2(n_82),
.B1(n_80),
.B2(n_81),
.Y(n_1480)
);

INVx1_ASAP7_75t_L g1481 ( 
.A(n_1427),
.Y(n_1481)
);

OAI22xp5_ASAP7_75t_L g1482 ( 
.A1(n_1429),
.A2(n_1441),
.B1(n_1406),
.B2(n_1404),
.Y(n_1482)
);

INVx1_ASAP7_75t_L g1483 ( 
.A(n_1397),
.Y(n_1483)
);

NAND2xp5_ASAP7_75t_L g1484 ( 
.A(n_1421),
.B(n_81),
.Y(n_1484)
);

AOI22xp33_ASAP7_75t_L g1485 ( 
.A1(n_1432),
.A2(n_84),
.B1(n_82),
.B2(n_83),
.Y(n_1485)
);

INVx1_ASAP7_75t_L g1486 ( 
.A(n_1371),
.Y(n_1486)
);

HB1xp67_ASAP7_75t_L g1487 ( 
.A(n_1453),
.Y(n_1487)
);

CKINVDCx5p33_ASAP7_75t_R g1488 ( 
.A(n_1376),
.Y(n_1488)
);

OAI22xp33_ASAP7_75t_L g1489 ( 
.A1(n_1402),
.A2(n_85),
.B1(n_83),
.B2(n_84),
.Y(n_1489)
);

INVx4_ASAP7_75t_L g1490 ( 
.A(n_1381),
.Y(n_1490)
);

OAI21xp5_ASAP7_75t_SL g1491 ( 
.A1(n_1361),
.A2(n_85),
.B(n_86),
.Y(n_1491)
);

AOI22xp33_ASAP7_75t_SL g1492 ( 
.A1(n_1416),
.A2(n_1425),
.B1(n_1372),
.B2(n_1367),
.Y(n_1492)
);

AOI22xp33_ASAP7_75t_L g1493 ( 
.A1(n_1408),
.A2(n_89),
.B1(n_87),
.B2(n_88),
.Y(n_1493)
);

INVx2_ASAP7_75t_L g1494 ( 
.A(n_1376),
.Y(n_1494)
);

INVx5_ASAP7_75t_L g1495 ( 
.A(n_1362),
.Y(n_1495)
);

INVx2_ASAP7_75t_L g1496 ( 
.A(n_1383),
.Y(n_1496)
);

INVx6_ASAP7_75t_L g1497 ( 
.A(n_1381),
.Y(n_1497)
);

OAI22xp5_ASAP7_75t_SL g1498 ( 
.A1(n_1433),
.A2(n_89),
.B1(n_87),
.B2(n_88),
.Y(n_1498)
);

INVx2_ASAP7_75t_L g1499 ( 
.A(n_1383),
.Y(n_1499)
);

INVx6_ASAP7_75t_L g1500 ( 
.A(n_1401),
.Y(n_1500)
);

INVx1_ASAP7_75t_L g1501 ( 
.A(n_1378),
.Y(n_1501)
);

CKINVDCx16_ASAP7_75t_R g1502 ( 
.A(n_1442),
.Y(n_1502)
);

OAI21xp5_ASAP7_75t_SL g1503 ( 
.A1(n_1447),
.A2(n_90),
.B(n_91),
.Y(n_1503)
);

BUFx8_ASAP7_75t_SL g1504 ( 
.A(n_1420),
.Y(n_1504)
);

INVx1_ASAP7_75t_L g1505 ( 
.A(n_1436),
.Y(n_1505)
);

CKINVDCx20_ASAP7_75t_R g1506 ( 
.A(n_1399),
.Y(n_1506)
);

INVx1_ASAP7_75t_L g1507 ( 
.A(n_1435),
.Y(n_1507)
);

AOI22xp33_ASAP7_75t_SL g1508 ( 
.A1(n_1440),
.A2(n_92),
.B1(n_90),
.B2(n_91),
.Y(n_1508)
);

BUFx4f_ASAP7_75t_SL g1509 ( 
.A(n_1446),
.Y(n_1509)
);

AND2x2_ASAP7_75t_L g1510 ( 
.A(n_1423),
.B(n_314),
.Y(n_1510)
);

INVx2_ASAP7_75t_SL g1511 ( 
.A(n_1438),
.Y(n_1511)
);

INVx1_ASAP7_75t_L g1512 ( 
.A(n_1435),
.Y(n_1512)
);

NAND2xp5_ASAP7_75t_L g1513 ( 
.A(n_1415),
.B(n_93),
.Y(n_1513)
);

INVx1_ASAP7_75t_SL g1514 ( 
.A(n_1448),
.Y(n_1514)
);

BUFx2_ASAP7_75t_L g1515 ( 
.A(n_1410),
.Y(n_1515)
);

BUFx3_ASAP7_75t_L g1516 ( 
.A(n_1434),
.Y(n_1516)
);

CKINVDCx11_ASAP7_75t_R g1517 ( 
.A(n_1428),
.Y(n_1517)
);

INVx2_ASAP7_75t_L g1518 ( 
.A(n_1365),
.Y(n_1518)
);

NAND2xp5_ASAP7_75t_L g1519 ( 
.A(n_1417),
.B(n_93),
.Y(n_1519)
);

BUFx2_ASAP7_75t_L g1520 ( 
.A(n_1410),
.Y(n_1520)
);

OAI21xp5_ASAP7_75t_SL g1521 ( 
.A1(n_1414),
.A2(n_1403),
.B(n_1380),
.Y(n_1521)
);

INVx2_ASAP7_75t_SL g1522 ( 
.A(n_1375),
.Y(n_1522)
);

BUFx8_ASAP7_75t_SL g1523 ( 
.A(n_1395),
.Y(n_1523)
);

CKINVDCx5p33_ASAP7_75t_R g1524 ( 
.A(n_1426),
.Y(n_1524)
);

INVx1_ASAP7_75t_L g1525 ( 
.A(n_1422),
.Y(n_1525)
);

NAND2xp5_ASAP7_75t_L g1526 ( 
.A(n_1451),
.B(n_94),
.Y(n_1526)
);

NAND2xp5_ASAP7_75t_L g1527 ( 
.A(n_1398),
.B(n_94),
.Y(n_1527)
);

INVx6_ASAP7_75t_L g1528 ( 
.A(n_1437),
.Y(n_1528)
);

NAND2xp5_ASAP7_75t_L g1529 ( 
.A(n_1419),
.B(n_95),
.Y(n_1529)
);

BUFx3_ASAP7_75t_L g1530 ( 
.A(n_1405),
.Y(n_1530)
);

AOI21xp33_ASAP7_75t_L g1531 ( 
.A1(n_1389),
.A2(n_95),
.B(n_96),
.Y(n_1531)
);

BUFx3_ASAP7_75t_L g1532 ( 
.A(n_1375),
.Y(n_1532)
);

AOI22xp33_ASAP7_75t_L g1533 ( 
.A1(n_1384),
.A2(n_98),
.B1(n_96),
.B2(n_97),
.Y(n_1533)
);

CKINVDCx5p33_ASAP7_75t_R g1534 ( 
.A(n_1392),
.Y(n_1534)
);

INVx1_ASAP7_75t_L g1535 ( 
.A(n_1422),
.Y(n_1535)
);

AND2x2_ASAP7_75t_L g1536 ( 
.A(n_1430),
.B(n_315),
.Y(n_1536)
);

INVx2_ASAP7_75t_L g1537 ( 
.A(n_1365),
.Y(n_1537)
);

INVx2_ASAP7_75t_L g1538 ( 
.A(n_1411),
.Y(n_1538)
);

INVx1_ASAP7_75t_L g1539 ( 
.A(n_1363),
.Y(n_1539)
);

CKINVDCx5p33_ASAP7_75t_R g1540 ( 
.A(n_1385),
.Y(n_1540)
);

BUFx12f_ASAP7_75t_L g1541 ( 
.A(n_1444),
.Y(n_1541)
);

BUFx3_ASAP7_75t_L g1542 ( 
.A(n_1445),
.Y(n_1542)
);

INVx1_ASAP7_75t_L g1543 ( 
.A(n_1452),
.Y(n_1543)
);

BUFx3_ASAP7_75t_L g1544 ( 
.A(n_1455),
.Y(n_1544)
);

BUFx12f_ASAP7_75t_L g1545 ( 
.A(n_1400),
.Y(n_1545)
);

OAI22xp5_ASAP7_75t_L g1546 ( 
.A1(n_1390),
.A2(n_99),
.B1(n_97),
.B2(n_98),
.Y(n_1546)
);

INVx5_ASAP7_75t_L g1547 ( 
.A(n_1393),
.Y(n_1547)
);

INVx1_ASAP7_75t_L g1548 ( 
.A(n_1374),
.Y(n_1548)
);

BUFx4f_ASAP7_75t_SL g1549 ( 
.A(n_1377),
.Y(n_1549)
);

AOI22xp33_ASAP7_75t_L g1550 ( 
.A1(n_1369),
.A2(n_101),
.B1(n_99),
.B2(n_100),
.Y(n_1550)
);

OAI22xp33_ASAP7_75t_L g1551 ( 
.A1(n_1431),
.A2(n_104),
.B1(n_100),
.B2(n_103),
.Y(n_1551)
);

OAI21xp5_ASAP7_75t_SL g1552 ( 
.A1(n_1369),
.A2(n_103),
.B(n_104),
.Y(n_1552)
);

AOI22xp33_ASAP7_75t_SL g1553 ( 
.A1(n_1369),
.A2(n_107),
.B1(n_105),
.B2(n_106),
.Y(n_1553)
);

CKINVDCx11_ASAP7_75t_R g1554 ( 
.A(n_1391),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_1456),
.Y(n_1555)
);

INVx1_ASAP7_75t_L g1556 ( 
.A(n_1478),
.Y(n_1556)
);

INVx1_ASAP7_75t_L g1557 ( 
.A(n_1481),
.Y(n_1557)
);

INVx1_ASAP7_75t_L g1558 ( 
.A(n_1483),
.Y(n_1558)
);

BUFx2_ASAP7_75t_L g1559 ( 
.A(n_1461),
.Y(n_1559)
);

AOI22xp33_ASAP7_75t_L g1560 ( 
.A1(n_1462),
.A2(n_107),
.B1(n_105),
.B2(n_106),
.Y(n_1560)
);

INVx2_ASAP7_75t_L g1561 ( 
.A(n_1458),
.Y(n_1561)
);

INVx1_ASAP7_75t_L g1562 ( 
.A(n_1457),
.Y(n_1562)
);

INVxp33_ASAP7_75t_L g1563 ( 
.A(n_1554),
.Y(n_1563)
);

INVx3_ASAP7_75t_L g1564 ( 
.A(n_1497),
.Y(n_1564)
);

INVx2_ASAP7_75t_L g1565 ( 
.A(n_1471),
.Y(n_1565)
);

INVx1_ASAP7_75t_L g1566 ( 
.A(n_1468),
.Y(n_1566)
);

INVxp67_ASAP7_75t_L g1567 ( 
.A(n_1479),
.Y(n_1567)
);

INVx3_ASAP7_75t_L g1568 ( 
.A(n_1497),
.Y(n_1568)
);

INVx1_ASAP7_75t_L g1569 ( 
.A(n_1507),
.Y(n_1569)
);

AND2x2_ASAP7_75t_L g1570 ( 
.A(n_1502),
.B(n_1486),
.Y(n_1570)
);

BUFx6f_ASAP7_75t_SL g1571 ( 
.A(n_1490),
.Y(n_1571)
);

NAND2xp5_ASAP7_75t_L g1572 ( 
.A(n_1473),
.B(n_108),
.Y(n_1572)
);

INVx1_ASAP7_75t_L g1573 ( 
.A(n_1512),
.Y(n_1573)
);

INVx1_ASAP7_75t_L g1574 ( 
.A(n_1474),
.Y(n_1574)
);

INVx1_ASAP7_75t_L g1575 ( 
.A(n_1525),
.Y(n_1575)
);

HB1xp67_ASAP7_75t_L g1576 ( 
.A(n_1487),
.Y(n_1576)
);

INVx3_ASAP7_75t_L g1577 ( 
.A(n_1465),
.Y(n_1577)
);

INVx2_ASAP7_75t_L g1578 ( 
.A(n_1505),
.Y(n_1578)
);

AOI21x1_ASAP7_75t_L g1579 ( 
.A1(n_1529),
.A2(n_108),
.B(n_109),
.Y(n_1579)
);

INVx2_ASAP7_75t_L g1580 ( 
.A(n_1496),
.Y(n_1580)
);

INVx1_ASAP7_75t_L g1581 ( 
.A(n_1535),
.Y(n_1581)
);

INVx1_ASAP7_75t_L g1582 ( 
.A(n_1515),
.Y(n_1582)
);

INVx2_ASAP7_75t_L g1583 ( 
.A(n_1499),
.Y(n_1583)
);

INVx3_ASAP7_75t_L g1584 ( 
.A(n_1465),
.Y(n_1584)
);

INVx3_ASAP7_75t_L g1585 ( 
.A(n_1476),
.Y(n_1585)
);

INVx1_ASAP7_75t_L g1586 ( 
.A(n_1520),
.Y(n_1586)
);

OAI21x1_ASAP7_75t_L g1587 ( 
.A1(n_1539),
.A2(n_317),
.B(n_316),
.Y(n_1587)
);

INVx1_ASAP7_75t_L g1588 ( 
.A(n_1501),
.Y(n_1588)
);

INVx1_ASAP7_75t_L g1589 ( 
.A(n_1518),
.Y(n_1589)
);

INVx1_ASAP7_75t_L g1590 ( 
.A(n_1537),
.Y(n_1590)
);

NAND2xp5_ASAP7_75t_L g1591 ( 
.A(n_1467),
.B(n_109),
.Y(n_1591)
);

BUFx6f_ASAP7_75t_L g1592 ( 
.A(n_1476),
.Y(n_1592)
);

BUFx3_ASAP7_75t_L g1593 ( 
.A(n_1459),
.Y(n_1593)
);

AND2x4_ASAP7_75t_L g1594 ( 
.A(n_1466),
.B(n_318),
.Y(n_1594)
);

BUFx2_ASAP7_75t_L g1595 ( 
.A(n_1459),
.Y(n_1595)
);

AOI22xp33_ASAP7_75t_SL g1596 ( 
.A1(n_1498),
.A2(n_112),
.B1(n_110),
.B2(n_111),
.Y(n_1596)
);

INVx1_ASAP7_75t_L g1597 ( 
.A(n_1522),
.Y(n_1597)
);

OAI22xp5_ASAP7_75t_L g1598 ( 
.A1(n_1550),
.A2(n_113),
.B1(n_110),
.B2(n_112),
.Y(n_1598)
);

INVx2_ASAP7_75t_L g1599 ( 
.A(n_1494),
.Y(n_1599)
);

AOI21x1_ASAP7_75t_L g1600 ( 
.A1(n_1526),
.A2(n_114),
.B(n_115),
.Y(n_1600)
);

OA21x2_ASAP7_75t_L g1601 ( 
.A1(n_1543),
.A2(n_1531),
.B(n_1548),
.Y(n_1601)
);

INVx2_ASAP7_75t_L g1602 ( 
.A(n_1538),
.Y(n_1602)
);

INVx2_ASAP7_75t_L g1603 ( 
.A(n_1511),
.Y(n_1603)
);

INVx1_ASAP7_75t_L g1604 ( 
.A(n_1532),
.Y(n_1604)
);

INVx1_ASAP7_75t_L g1605 ( 
.A(n_1484),
.Y(n_1605)
);

INVx1_ASAP7_75t_L g1606 ( 
.A(n_1519),
.Y(n_1606)
);

INVx2_ASAP7_75t_L g1607 ( 
.A(n_1528),
.Y(n_1607)
);

INVx3_ASAP7_75t_L g1608 ( 
.A(n_1495),
.Y(n_1608)
);

INVx1_ASAP7_75t_L g1609 ( 
.A(n_1516),
.Y(n_1609)
);

INVx1_ASAP7_75t_L g1610 ( 
.A(n_1530),
.Y(n_1610)
);

OAI21xp5_ASAP7_75t_L g1611 ( 
.A1(n_1552),
.A2(n_321),
.B(n_319),
.Y(n_1611)
);

NAND2xp5_ASAP7_75t_L g1612 ( 
.A(n_1482),
.B(n_114),
.Y(n_1612)
);

INVx1_ASAP7_75t_L g1613 ( 
.A(n_1528),
.Y(n_1613)
);

AND2x2_ASAP7_75t_L g1614 ( 
.A(n_1463),
.B(n_115),
.Y(n_1614)
);

INVx2_ASAP7_75t_L g1615 ( 
.A(n_1542),
.Y(n_1615)
);

OR2x2_ASAP7_75t_L g1616 ( 
.A(n_1470),
.B(n_323),
.Y(n_1616)
);

INVx1_ASAP7_75t_L g1617 ( 
.A(n_1544),
.Y(n_1617)
);

AOI21x1_ASAP7_75t_L g1618 ( 
.A1(n_1546),
.A2(n_1527),
.B(n_1513),
.Y(n_1618)
);

INVx1_ASAP7_75t_L g1619 ( 
.A(n_1536),
.Y(n_1619)
);

INVx2_ASAP7_75t_SL g1620 ( 
.A(n_1488),
.Y(n_1620)
);

INVx1_ASAP7_75t_SL g1621 ( 
.A(n_1509),
.Y(n_1621)
);

INVx1_ASAP7_75t_L g1622 ( 
.A(n_1517),
.Y(n_1622)
);

NAND2xp5_ASAP7_75t_L g1623 ( 
.A(n_1524),
.B(n_1553),
.Y(n_1623)
);

INVx2_ASAP7_75t_L g1624 ( 
.A(n_1547),
.Y(n_1624)
);

BUFx3_ASAP7_75t_L g1625 ( 
.A(n_1506),
.Y(n_1625)
);

OAI21xp5_ASAP7_75t_L g1626 ( 
.A1(n_1492),
.A2(n_324),
.B(n_325),
.Y(n_1626)
);

OAI21x1_ASAP7_75t_L g1627 ( 
.A1(n_1521),
.A2(n_326),
.B(n_327),
.Y(n_1627)
);

INVx1_ASAP7_75t_L g1628 ( 
.A(n_1549),
.Y(n_1628)
);

A2O1A1Ixp33_ASAP7_75t_L g1629 ( 
.A1(n_1491),
.A2(n_330),
.B(n_328),
.C(n_329),
.Y(n_1629)
);

INVx3_ASAP7_75t_L g1630 ( 
.A(n_1495),
.Y(n_1630)
);

INVx2_ASAP7_75t_L g1631 ( 
.A(n_1547),
.Y(n_1631)
);

INVx2_ASAP7_75t_L g1632 ( 
.A(n_1547),
.Y(n_1632)
);

AOI22xp33_ASAP7_75t_L g1633 ( 
.A1(n_1460),
.A2(n_1551),
.B1(n_1508),
.B2(n_1480),
.Y(n_1633)
);

INVx1_ASAP7_75t_L g1634 ( 
.A(n_1540),
.Y(n_1634)
);

CKINVDCx12_ASAP7_75t_R g1635 ( 
.A(n_1510),
.Y(n_1635)
);

INVx1_ASAP7_75t_L g1636 ( 
.A(n_1541),
.Y(n_1636)
);

INVx2_ASAP7_75t_L g1637 ( 
.A(n_1500),
.Y(n_1637)
);

INVx1_ASAP7_75t_L g1638 ( 
.A(n_1534),
.Y(n_1638)
);

INVx1_ASAP7_75t_L g1639 ( 
.A(n_1469),
.Y(n_1639)
);

BUFx2_ASAP7_75t_L g1640 ( 
.A(n_1495),
.Y(n_1640)
);

INVx2_ASAP7_75t_L g1641 ( 
.A(n_1500),
.Y(n_1641)
);

INVx1_ASAP7_75t_L g1642 ( 
.A(n_1514),
.Y(n_1642)
);

AND2x2_ASAP7_75t_L g1643 ( 
.A(n_1464),
.B(n_562),
.Y(n_1643)
);

INVx1_ASAP7_75t_L g1644 ( 
.A(n_1489),
.Y(n_1644)
);

AND2x2_ASAP7_75t_L g1645 ( 
.A(n_1477),
.B(n_332),
.Y(n_1645)
);

INVx3_ASAP7_75t_L g1646 ( 
.A(n_1545),
.Y(n_1646)
);

INVx1_ASAP7_75t_L g1647 ( 
.A(n_1477),
.Y(n_1647)
);

INVx2_ASAP7_75t_L g1648 ( 
.A(n_1523),
.Y(n_1648)
);

BUFx3_ASAP7_75t_L g1649 ( 
.A(n_1504),
.Y(n_1649)
);

AND2x2_ASAP7_75t_L g1650 ( 
.A(n_1485),
.B(n_561),
.Y(n_1650)
);

INVx1_ASAP7_75t_L g1651 ( 
.A(n_1503),
.Y(n_1651)
);

BUFx3_ASAP7_75t_L g1652 ( 
.A(n_1475),
.Y(n_1652)
);

OAI22xp5_ASAP7_75t_SL g1653 ( 
.A1(n_1472),
.A2(n_337),
.B1(n_334),
.B2(n_336),
.Y(n_1653)
);

HB1xp67_ASAP7_75t_L g1654 ( 
.A(n_1533),
.Y(n_1654)
);

INVx1_ASAP7_75t_L g1655 ( 
.A(n_1493),
.Y(n_1655)
);

AO31x2_ASAP7_75t_L g1656 ( 
.A1(n_1525),
.A2(n_340),
.A3(n_338),
.B(n_339),
.Y(n_1656)
);

INVx1_ASAP7_75t_L g1657 ( 
.A(n_1456),
.Y(n_1657)
);

NAND2xp5_ASAP7_75t_L g1658 ( 
.A(n_1468),
.B(n_341),
.Y(n_1658)
);

INVx1_ASAP7_75t_L g1659 ( 
.A(n_1478),
.Y(n_1659)
);

AND2x2_ASAP7_75t_L g1660 ( 
.A(n_1468),
.B(n_560),
.Y(n_1660)
);

INVx2_ASAP7_75t_L g1661 ( 
.A(n_1458),
.Y(n_1661)
);

OAI21x1_ASAP7_75t_L g1662 ( 
.A1(n_1496),
.A2(n_342),
.B(n_343),
.Y(n_1662)
);

INVx1_ASAP7_75t_L g1663 ( 
.A(n_1478),
.Y(n_1663)
);

INVx2_ASAP7_75t_L g1664 ( 
.A(n_1458),
.Y(n_1664)
);

INVx1_ASAP7_75t_SL g1665 ( 
.A(n_1509),
.Y(n_1665)
);

INVx2_ASAP7_75t_L g1666 ( 
.A(n_1458),
.Y(n_1666)
);

HB1xp67_ASAP7_75t_L g1667 ( 
.A(n_1461),
.Y(n_1667)
);

AND2x2_ASAP7_75t_L g1668 ( 
.A(n_1468),
.B(n_344),
.Y(n_1668)
);

INVx1_ASAP7_75t_L g1669 ( 
.A(n_1556),
.Y(n_1669)
);

INVx1_ASAP7_75t_L g1670 ( 
.A(n_1556),
.Y(n_1670)
);

AND2x4_ASAP7_75t_L g1671 ( 
.A(n_1607),
.B(n_345),
.Y(n_1671)
);

INVx2_ASAP7_75t_L g1672 ( 
.A(n_1561),
.Y(n_1672)
);

OR2x2_ASAP7_75t_L g1673 ( 
.A(n_1566),
.B(n_346),
.Y(n_1673)
);

OA21x2_ASAP7_75t_L g1674 ( 
.A1(n_1588),
.A2(n_558),
.B(n_347),
.Y(n_1674)
);

INVx2_ASAP7_75t_L g1675 ( 
.A(n_1661),
.Y(n_1675)
);

INVx2_ASAP7_75t_L g1676 ( 
.A(n_1664),
.Y(n_1676)
);

INVx1_ASAP7_75t_L g1677 ( 
.A(n_1557),
.Y(n_1677)
);

INVx2_ASAP7_75t_L g1678 ( 
.A(n_1666),
.Y(n_1678)
);

BUFx4f_ASAP7_75t_SL g1679 ( 
.A(n_1625),
.Y(n_1679)
);

OR2x2_ASAP7_75t_L g1680 ( 
.A(n_1667),
.B(n_348),
.Y(n_1680)
);

BUFx6f_ASAP7_75t_L g1681 ( 
.A(n_1592),
.Y(n_1681)
);

AO21x2_ASAP7_75t_L g1682 ( 
.A1(n_1624),
.A2(n_349),
.B(n_350),
.Y(n_1682)
);

INVx3_ASAP7_75t_L g1683 ( 
.A(n_1608),
.Y(n_1683)
);

AND2x2_ASAP7_75t_L g1684 ( 
.A(n_1559),
.B(n_351),
.Y(n_1684)
);

AND2x4_ASAP7_75t_L g1685 ( 
.A(n_1615),
.B(n_352),
.Y(n_1685)
);

INVx2_ASAP7_75t_L g1686 ( 
.A(n_1555),
.Y(n_1686)
);

CKINVDCx5p33_ASAP7_75t_R g1687 ( 
.A(n_1649),
.Y(n_1687)
);

HB1xp67_ASAP7_75t_L g1688 ( 
.A(n_1576),
.Y(n_1688)
);

AO21x2_ASAP7_75t_L g1689 ( 
.A1(n_1631),
.A2(n_353),
.B(n_355),
.Y(n_1689)
);

INVx1_ASAP7_75t_L g1690 ( 
.A(n_1562),
.Y(n_1690)
);

BUFx2_ASAP7_75t_L g1691 ( 
.A(n_1567),
.Y(n_1691)
);

HB1xp67_ASAP7_75t_L g1692 ( 
.A(n_1642),
.Y(n_1692)
);

OA21x2_ASAP7_75t_L g1693 ( 
.A1(n_1575),
.A2(n_357),
.B(n_358),
.Y(n_1693)
);

INVx4_ASAP7_75t_L g1694 ( 
.A(n_1646),
.Y(n_1694)
);

INVx1_ASAP7_75t_L g1695 ( 
.A(n_1557),
.Y(n_1695)
);

INVx1_ASAP7_75t_L g1696 ( 
.A(n_1659),
.Y(n_1696)
);

INVx1_ASAP7_75t_L g1697 ( 
.A(n_1659),
.Y(n_1697)
);

AND2x2_ASAP7_75t_L g1698 ( 
.A(n_1570),
.B(n_1622),
.Y(n_1698)
);

INVxp67_ASAP7_75t_L g1699 ( 
.A(n_1605),
.Y(n_1699)
);

NAND2xp5_ASAP7_75t_L g1700 ( 
.A(n_1606),
.B(n_359),
.Y(n_1700)
);

HB1xp67_ASAP7_75t_L g1701 ( 
.A(n_1582),
.Y(n_1701)
);

BUFx6f_ASAP7_75t_L g1702 ( 
.A(n_1592),
.Y(n_1702)
);

NAND2xp5_ASAP7_75t_L g1703 ( 
.A(n_1574),
.B(n_360),
.Y(n_1703)
);

AO21x2_ASAP7_75t_L g1704 ( 
.A1(n_1632),
.A2(n_361),
.B(n_363),
.Y(n_1704)
);

AO21x2_ASAP7_75t_L g1705 ( 
.A1(n_1581),
.A2(n_364),
.B(n_365),
.Y(n_1705)
);

INVx2_ASAP7_75t_L g1706 ( 
.A(n_1657),
.Y(n_1706)
);

NOR2xp33_ASAP7_75t_L g1707 ( 
.A(n_1634),
.B(n_366),
.Y(n_1707)
);

INVx1_ASAP7_75t_L g1708 ( 
.A(n_1562),
.Y(n_1708)
);

INVx1_ASAP7_75t_L g1709 ( 
.A(n_1663),
.Y(n_1709)
);

OAI21x1_ASAP7_75t_L g1710 ( 
.A1(n_1627),
.A2(n_367),
.B(n_369),
.Y(n_1710)
);

AND3x2_ASAP7_75t_L g1711 ( 
.A(n_1595),
.B(n_370),
.C(n_372),
.Y(n_1711)
);

AND2x2_ASAP7_75t_L g1712 ( 
.A(n_1637),
.B(n_374),
.Y(n_1712)
);

INVxp67_ASAP7_75t_SL g1713 ( 
.A(n_1586),
.Y(n_1713)
);

BUFx2_ASAP7_75t_L g1714 ( 
.A(n_1636),
.Y(n_1714)
);

OR2x6_ASAP7_75t_L g1715 ( 
.A(n_1646),
.B(n_376),
.Y(n_1715)
);

AND2x2_ASAP7_75t_L g1716 ( 
.A(n_1641),
.B(n_377),
.Y(n_1716)
);

INVx2_ASAP7_75t_L g1717 ( 
.A(n_1565),
.Y(n_1717)
);

NAND2xp5_ASAP7_75t_L g1718 ( 
.A(n_1638),
.B(n_378),
.Y(n_1718)
);

INVx1_ASAP7_75t_L g1719 ( 
.A(n_1663),
.Y(n_1719)
);

BUFx3_ASAP7_75t_L g1720 ( 
.A(n_1593),
.Y(n_1720)
);

AND2x2_ASAP7_75t_L g1721 ( 
.A(n_1609),
.B(n_379),
.Y(n_1721)
);

AND2x2_ASAP7_75t_L g1722 ( 
.A(n_1610),
.B(n_380),
.Y(n_1722)
);

OA21x2_ASAP7_75t_L g1723 ( 
.A1(n_1569),
.A2(n_557),
.B(n_383),
.Y(n_1723)
);

HB1xp67_ASAP7_75t_L g1724 ( 
.A(n_1558),
.Y(n_1724)
);

HB1xp67_ASAP7_75t_L g1725 ( 
.A(n_1558),
.Y(n_1725)
);

INVx1_ASAP7_75t_L g1726 ( 
.A(n_1573),
.Y(n_1726)
);

AND2x2_ASAP7_75t_L g1727 ( 
.A(n_1617),
.B(n_384),
.Y(n_1727)
);

AO21x2_ASAP7_75t_L g1728 ( 
.A1(n_1597),
.A2(n_385),
.B(n_387),
.Y(n_1728)
);

NAND2xp5_ASAP7_75t_L g1729 ( 
.A(n_1619),
.B(n_388),
.Y(n_1729)
);

INVx1_ASAP7_75t_L g1730 ( 
.A(n_1578),
.Y(n_1730)
);

INVx2_ASAP7_75t_SL g1731 ( 
.A(n_1564),
.Y(n_1731)
);

INVx2_ASAP7_75t_L g1732 ( 
.A(n_1599),
.Y(n_1732)
);

INVx2_ASAP7_75t_L g1733 ( 
.A(n_1589),
.Y(n_1733)
);

INVx1_ASAP7_75t_L g1734 ( 
.A(n_1590),
.Y(n_1734)
);

INVx1_ASAP7_75t_L g1735 ( 
.A(n_1580),
.Y(n_1735)
);

BUFx2_ASAP7_75t_L g1736 ( 
.A(n_1628),
.Y(n_1736)
);

INVx4_ASAP7_75t_L g1737 ( 
.A(n_1608),
.Y(n_1737)
);

NAND2xp5_ASAP7_75t_L g1738 ( 
.A(n_1644),
.B(n_389),
.Y(n_1738)
);

NAND2xp5_ASAP7_75t_L g1739 ( 
.A(n_1651),
.B(n_390),
.Y(n_1739)
);

INVx2_ASAP7_75t_SL g1740 ( 
.A(n_1564),
.Y(n_1740)
);

OA21x2_ASAP7_75t_L g1741 ( 
.A1(n_1604),
.A2(n_1603),
.B(n_1602),
.Y(n_1741)
);

AND2x2_ASAP7_75t_L g1742 ( 
.A(n_1568),
.B(n_1621),
.Y(n_1742)
);

INVx2_ASAP7_75t_L g1743 ( 
.A(n_1583),
.Y(n_1743)
);

INVx1_ASAP7_75t_L g1744 ( 
.A(n_1604),
.Y(n_1744)
);

INVx2_ASAP7_75t_L g1745 ( 
.A(n_1640),
.Y(n_1745)
);

AND2x4_ASAP7_75t_L g1746 ( 
.A(n_1745),
.B(n_1613),
.Y(n_1746)
);

BUFx6f_ASAP7_75t_L g1747 ( 
.A(n_1681),
.Y(n_1747)
);

AND2x2_ASAP7_75t_L g1748 ( 
.A(n_1688),
.B(n_1563),
.Y(n_1748)
);

HB1xp67_ASAP7_75t_L g1749 ( 
.A(n_1741),
.Y(n_1749)
);

HB1xp67_ASAP7_75t_L g1750 ( 
.A(n_1741),
.Y(n_1750)
);

AND2x2_ASAP7_75t_L g1751 ( 
.A(n_1691),
.B(n_1665),
.Y(n_1751)
);

INVx1_ASAP7_75t_L g1752 ( 
.A(n_1724),
.Y(n_1752)
);

AND2x2_ASAP7_75t_L g1753 ( 
.A(n_1692),
.B(n_1568),
.Y(n_1753)
);

NAND2xp5_ASAP7_75t_L g1754 ( 
.A(n_1699),
.B(n_1601),
.Y(n_1754)
);

AND2x2_ASAP7_75t_L g1755 ( 
.A(n_1714),
.B(n_1577),
.Y(n_1755)
);

INVx2_ASAP7_75t_L g1756 ( 
.A(n_1686),
.Y(n_1756)
);

AND2x2_ASAP7_75t_L g1757 ( 
.A(n_1698),
.B(n_1577),
.Y(n_1757)
);

AND2x2_ASAP7_75t_L g1758 ( 
.A(n_1736),
.B(n_1584),
.Y(n_1758)
);

INVx2_ASAP7_75t_L g1759 ( 
.A(n_1706),
.Y(n_1759)
);

AND2x2_ASAP7_75t_L g1760 ( 
.A(n_1683),
.B(n_1584),
.Y(n_1760)
);

NAND2xp5_ASAP7_75t_L g1761 ( 
.A(n_1725),
.B(n_1601),
.Y(n_1761)
);

INVx1_ASAP7_75t_L g1762 ( 
.A(n_1669),
.Y(n_1762)
);

NOR2x1_ASAP7_75t_L g1763 ( 
.A(n_1694),
.B(n_1630),
.Y(n_1763)
);

OR2x2_ASAP7_75t_L g1764 ( 
.A(n_1701),
.B(n_1713),
.Y(n_1764)
);

INVx1_ASAP7_75t_L g1765 ( 
.A(n_1669),
.Y(n_1765)
);

INVx2_ASAP7_75t_SL g1766 ( 
.A(n_1720),
.Y(n_1766)
);

INVxp67_ASAP7_75t_SL g1767 ( 
.A(n_1670),
.Y(n_1767)
);

AND2x2_ASAP7_75t_L g1768 ( 
.A(n_1683),
.B(n_1648),
.Y(n_1768)
);

OR2x2_ASAP7_75t_L g1769 ( 
.A(n_1730),
.B(n_1616),
.Y(n_1769)
);

AND2x2_ASAP7_75t_L g1770 ( 
.A(n_1694),
.B(n_1620),
.Y(n_1770)
);

OR2x2_ASAP7_75t_L g1771 ( 
.A(n_1730),
.B(n_1612),
.Y(n_1771)
);

BUFx3_ASAP7_75t_L g1772 ( 
.A(n_1681),
.Y(n_1772)
);

AND2x2_ASAP7_75t_L g1773 ( 
.A(n_1672),
.B(n_1675),
.Y(n_1773)
);

INVx2_ASAP7_75t_L g1774 ( 
.A(n_1732),
.Y(n_1774)
);

AND2x2_ASAP7_75t_L g1775 ( 
.A(n_1676),
.B(n_1630),
.Y(n_1775)
);

NAND2xp5_ASAP7_75t_L g1776 ( 
.A(n_1678),
.B(n_1591),
.Y(n_1776)
);

NAND2xp5_ASAP7_75t_L g1777 ( 
.A(n_1717),
.B(n_1618),
.Y(n_1777)
);

INVx1_ASAP7_75t_L g1778 ( 
.A(n_1670),
.Y(n_1778)
);

CKINVDCx14_ASAP7_75t_R g1779 ( 
.A(n_1687),
.Y(n_1779)
);

INVx1_ASAP7_75t_L g1780 ( 
.A(n_1677),
.Y(n_1780)
);

HB1xp67_ASAP7_75t_L g1781 ( 
.A(n_1677),
.Y(n_1781)
);

AND2x2_ASAP7_75t_L g1782 ( 
.A(n_1737),
.B(n_1585),
.Y(n_1782)
);

INVx1_ASAP7_75t_L g1783 ( 
.A(n_1695),
.Y(n_1783)
);

NOR2x1_ASAP7_75t_SL g1784 ( 
.A(n_1728),
.B(n_1592),
.Y(n_1784)
);

INVx2_ASAP7_75t_L g1785 ( 
.A(n_1695),
.Y(n_1785)
);

AND2x2_ASAP7_75t_L g1786 ( 
.A(n_1737),
.B(n_1585),
.Y(n_1786)
);

INVxp33_ASAP7_75t_L g1787 ( 
.A(n_1707),
.Y(n_1787)
);

INVx1_ASAP7_75t_L g1788 ( 
.A(n_1696),
.Y(n_1788)
);

INVx2_ASAP7_75t_L g1789 ( 
.A(n_1696),
.Y(n_1789)
);

AND2x2_ASAP7_75t_L g1790 ( 
.A(n_1731),
.B(n_1647),
.Y(n_1790)
);

NAND2xp5_ASAP7_75t_L g1791 ( 
.A(n_1697),
.B(n_1639),
.Y(n_1791)
);

INVx1_ASAP7_75t_L g1792 ( 
.A(n_1697),
.Y(n_1792)
);

AND2x2_ASAP7_75t_L g1793 ( 
.A(n_1740),
.B(n_1614),
.Y(n_1793)
);

HB1xp67_ASAP7_75t_L g1794 ( 
.A(n_1744),
.Y(n_1794)
);

INVx1_ASAP7_75t_L g1795 ( 
.A(n_1690),
.Y(n_1795)
);

INVx2_ASAP7_75t_L g1796 ( 
.A(n_1708),
.Y(n_1796)
);

BUFx2_ASAP7_75t_L g1797 ( 
.A(n_1744),
.Y(n_1797)
);

INVxp67_ASAP7_75t_R g1798 ( 
.A(n_1742),
.Y(n_1798)
);

NAND2xp5_ASAP7_75t_L g1799 ( 
.A(n_1709),
.B(n_1572),
.Y(n_1799)
);

BUFx2_ASAP7_75t_L g1800 ( 
.A(n_1681),
.Y(n_1800)
);

INVx1_ASAP7_75t_L g1801 ( 
.A(n_1719),
.Y(n_1801)
);

INVx1_ASAP7_75t_L g1802 ( 
.A(n_1726),
.Y(n_1802)
);

INVx1_ASAP7_75t_L g1803 ( 
.A(n_1734),
.Y(n_1803)
);

AND2x2_ASAP7_75t_L g1804 ( 
.A(n_1743),
.B(n_1668),
.Y(n_1804)
);

AND2x2_ASAP7_75t_L g1805 ( 
.A(n_1735),
.B(n_1660),
.Y(n_1805)
);

AND2x2_ASAP7_75t_L g1806 ( 
.A(n_1735),
.B(n_1594),
.Y(n_1806)
);

INVx3_ASAP7_75t_L g1807 ( 
.A(n_1702),
.Y(n_1807)
);

HB1xp67_ASAP7_75t_L g1808 ( 
.A(n_1734),
.Y(n_1808)
);

AND2x2_ASAP7_75t_L g1809 ( 
.A(n_1733),
.B(n_1594),
.Y(n_1809)
);

AND2x2_ASAP7_75t_L g1810 ( 
.A(n_1798),
.B(n_1748),
.Y(n_1810)
);

HB1xp67_ASAP7_75t_L g1811 ( 
.A(n_1749),
.Y(n_1811)
);

AND2x2_ASAP7_75t_L g1812 ( 
.A(n_1760),
.B(n_1702),
.Y(n_1812)
);

OR2x2_ASAP7_75t_L g1813 ( 
.A(n_1764),
.B(n_1673),
.Y(n_1813)
);

INVx1_ASAP7_75t_L g1814 ( 
.A(n_1808),
.Y(n_1814)
);

AND2x2_ASAP7_75t_L g1815 ( 
.A(n_1753),
.B(n_1702),
.Y(n_1815)
);

INVx2_ASAP7_75t_L g1816 ( 
.A(n_1749),
.Y(n_1816)
);

INVx1_ASAP7_75t_L g1817 ( 
.A(n_1808),
.Y(n_1817)
);

BUFx3_ASAP7_75t_L g1818 ( 
.A(n_1772),
.Y(n_1818)
);

AND2x2_ASAP7_75t_L g1819 ( 
.A(n_1782),
.B(n_1684),
.Y(n_1819)
);

BUFx3_ASAP7_75t_L g1820 ( 
.A(n_1772),
.Y(n_1820)
);

BUFx2_ASAP7_75t_L g1821 ( 
.A(n_1763),
.Y(n_1821)
);

INVx1_ASAP7_75t_L g1822 ( 
.A(n_1781),
.Y(n_1822)
);

INVx3_ASAP7_75t_L g1823 ( 
.A(n_1747),
.Y(n_1823)
);

NAND2xp5_ASAP7_75t_L g1824 ( 
.A(n_1777),
.B(n_1693),
.Y(n_1824)
);

INVx2_ASAP7_75t_L g1825 ( 
.A(n_1785),
.Y(n_1825)
);

INVx3_ASAP7_75t_L g1826 ( 
.A(n_1747),
.Y(n_1826)
);

INVx4_ASAP7_75t_L g1827 ( 
.A(n_1747),
.Y(n_1827)
);

AND2x2_ASAP7_75t_L g1828 ( 
.A(n_1786),
.B(n_1693),
.Y(n_1828)
);

BUFx2_ASAP7_75t_L g1829 ( 
.A(n_1800),
.Y(n_1829)
);

AND2x4_ASAP7_75t_SL g1830 ( 
.A(n_1758),
.B(n_1715),
.Y(n_1830)
);

INVx1_ASAP7_75t_L g1831 ( 
.A(n_1781),
.Y(n_1831)
);

INVx1_ASAP7_75t_L g1832 ( 
.A(n_1794),
.Y(n_1832)
);

HB1xp67_ASAP7_75t_L g1833 ( 
.A(n_1750),
.Y(n_1833)
);

AND2x4_ASAP7_75t_L g1834 ( 
.A(n_1752),
.B(n_1680),
.Y(n_1834)
);

INVx1_ASAP7_75t_L g1835 ( 
.A(n_1794),
.Y(n_1835)
);

INVx1_ASAP7_75t_L g1836 ( 
.A(n_1762),
.Y(n_1836)
);

HB1xp67_ASAP7_75t_L g1837 ( 
.A(n_1750),
.Y(n_1837)
);

BUFx2_ASAP7_75t_L g1838 ( 
.A(n_1746),
.Y(n_1838)
);

INVx2_ASAP7_75t_L g1839 ( 
.A(n_1785),
.Y(n_1839)
);

AND2x2_ASAP7_75t_L g1840 ( 
.A(n_1768),
.B(n_1723),
.Y(n_1840)
);

INVx1_ASAP7_75t_L g1841 ( 
.A(n_1765),
.Y(n_1841)
);

BUFx3_ASAP7_75t_L g1842 ( 
.A(n_1747),
.Y(n_1842)
);

BUFx6f_ASAP7_75t_L g1843 ( 
.A(n_1807),
.Y(n_1843)
);

INVxp67_ASAP7_75t_SL g1844 ( 
.A(n_1761),
.Y(n_1844)
);

AND2x4_ASAP7_75t_L g1845 ( 
.A(n_1746),
.B(n_1721),
.Y(n_1845)
);

INVx1_ASAP7_75t_SL g1846 ( 
.A(n_1797),
.Y(n_1846)
);

INVx1_ASAP7_75t_L g1847 ( 
.A(n_1778),
.Y(n_1847)
);

AND2x2_ASAP7_75t_L g1848 ( 
.A(n_1810),
.B(n_1755),
.Y(n_1848)
);

INVx1_ASAP7_75t_L g1849 ( 
.A(n_1836),
.Y(n_1849)
);

INVx1_ASAP7_75t_L g1850 ( 
.A(n_1841),
.Y(n_1850)
);

NAND4xp25_ASAP7_75t_L g1851 ( 
.A(n_1824),
.B(n_1596),
.C(n_1633),
.D(n_1560),
.Y(n_1851)
);

INVx2_ASAP7_75t_L g1852 ( 
.A(n_1842),
.Y(n_1852)
);

HB1xp67_ASAP7_75t_L g1853 ( 
.A(n_1846),
.Y(n_1853)
);

AND2x2_ASAP7_75t_L g1854 ( 
.A(n_1829),
.B(n_1770),
.Y(n_1854)
);

AND2x2_ASAP7_75t_L g1855 ( 
.A(n_1838),
.B(n_1757),
.Y(n_1855)
);

AND2x2_ASAP7_75t_L g1856 ( 
.A(n_1812),
.B(n_1793),
.Y(n_1856)
);

INVx2_ASAP7_75t_L g1857 ( 
.A(n_1842),
.Y(n_1857)
);

INVx1_ASAP7_75t_L g1858 ( 
.A(n_1847),
.Y(n_1858)
);

AND2x2_ASAP7_75t_L g1859 ( 
.A(n_1815),
.B(n_1751),
.Y(n_1859)
);

INVx1_ASAP7_75t_L g1860 ( 
.A(n_1811),
.Y(n_1860)
);

NAND2xp5_ASAP7_75t_L g1861 ( 
.A(n_1844),
.B(n_1754),
.Y(n_1861)
);

OR2x2_ASAP7_75t_L g1862 ( 
.A(n_1813),
.B(n_1777),
.Y(n_1862)
);

HB1xp67_ASAP7_75t_L g1863 ( 
.A(n_1846),
.Y(n_1863)
);

INVx2_ASAP7_75t_L g1864 ( 
.A(n_1823),
.Y(n_1864)
);

OR2x2_ASAP7_75t_L g1865 ( 
.A(n_1824),
.B(n_1754),
.Y(n_1865)
);

AND2x2_ASAP7_75t_L g1866 ( 
.A(n_1840),
.B(n_1775),
.Y(n_1866)
);

OR2x2_ASAP7_75t_L g1867 ( 
.A(n_1844),
.B(n_1771),
.Y(n_1867)
);

INVx4_ASAP7_75t_L g1868 ( 
.A(n_1827),
.Y(n_1868)
);

NAND2xp5_ASAP7_75t_L g1869 ( 
.A(n_1814),
.B(n_1802),
.Y(n_1869)
);

NAND2xp5_ASAP7_75t_L g1870 ( 
.A(n_1817),
.B(n_1822),
.Y(n_1870)
);

HB1xp67_ASAP7_75t_L g1871 ( 
.A(n_1811),
.Y(n_1871)
);

INVx1_ASAP7_75t_L g1872 ( 
.A(n_1833),
.Y(n_1872)
);

NAND2xp5_ASAP7_75t_L g1873 ( 
.A(n_1831),
.B(n_1832),
.Y(n_1873)
);

INVx1_ASAP7_75t_L g1874 ( 
.A(n_1833),
.Y(n_1874)
);

AND2x2_ASAP7_75t_L g1875 ( 
.A(n_1818),
.B(n_1790),
.Y(n_1875)
);

AND2x2_ASAP7_75t_L g1876 ( 
.A(n_1818),
.B(n_1805),
.Y(n_1876)
);

AND2x2_ASAP7_75t_L g1877 ( 
.A(n_1820),
.B(n_1804),
.Y(n_1877)
);

INVx1_ASAP7_75t_L g1878 ( 
.A(n_1837),
.Y(n_1878)
);

INVx2_ASAP7_75t_L g1879 ( 
.A(n_1823),
.Y(n_1879)
);

AND2x2_ASAP7_75t_L g1880 ( 
.A(n_1820),
.B(n_1807),
.Y(n_1880)
);

OR2x6_ASAP7_75t_L g1881 ( 
.A(n_1821),
.B(n_1715),
.Y(n_1881)
);

AOI22xp5_ASAP7_75t_L g1882 ( 
.A1(n_1851),
.A2(n_1652),
.B1(n_1834),
.B2(n_1828),
.Y(n_1882)
);

INVx2_ASAP7_75t_L g1883 ( 
.A(n_1868),
.Y(n_1883)
);

INVx3_ASAP7_75t_L g1884 ( 
.A(n_1868),
.Y(n_1884)
);

AND2x2_ASAP7_75t_L g1885 ( 
.A(n_1848),
.B(n_1827),
.Y(n_1885)
);

INVx2_ASAP7_75t_L g1886 ( 
.A(n_1880),
.Y(n_1886)
);

OR2x2_ASAP7_75t_L g1887 ( 
.A(n_1862),
.B(n_1776),
.Y(n_1887)
);

AND2x2_ASAP7_75t_L g1888 ( 
.A(n_1852),
.B(n_1826),
.Y(n_1888)
);

AND2x4_ASAP7_75t_SL g1889 ( 
.A(n_1881),
.B(n_1845),
.Y(n_1889)
);

NAND2xp5_ASAP7_75t_L g1890 ( 
.A(n_1853),
.B(n_1834),
.Y(n_1890)
);

NAND2xp5_ASAP7_75t_L g1891 ( 
.A(n_1863),
.B(n_1776),
.Y(n_1891)
);

INVx1_ASAP7_75t_L g1892 ( 
.A(n_1871),
.Y(n_1892)
);

OR2x2_ASAP7_75t_L g1893 ( 
.A(n_1867),
.B(n_1769),
.Y(n_1893)
);

AND2x2_ASAP7_75t_L g1894 ( 
.A(n_1857),
.B(n_1826),
.Y(n_1894)
);

INVx1_ASAP7_75t_L g1895 ( 
.A(n_1849),
.Y(n_1895)
);

INVx1_ASAP7_75t_L g1896 ( 
.A(n_1860),
.Y(n_1896)
);

INVx2_ASAP7_75t_L g1897 ( 
.A(n_1854),
.Y(n_1897)
);

AND2x4_ASAP7_75t_L g1898 ( 
.A(n_1881),
.B(n_1859),
.Y(n_1898)
);

HB1xp67_ASAP7_75t_L g1899 ( 
.A(n_1872),
.Y(n_1899)
);

OAI21xp33_ASAP7_75t_L g1900 ( 
.A1(n_1851),
.A2(n_1787),
.B(n_1623),
.Y(n_1900)
);

AND2x2_ASAP7_75t_L g1901 ( 
.A(n_1855),
.B(n_1845),
.Y(n_1901)
);

INVx2_ASAP7_75t_L g1902 ( 
.A(n_1875),
.Y(n_1902)
);

NAND2xp5_ASAP7_75t_L g1903 ( 
.A(n_1900),
.B(n_1864),
.Y(n_1903)
);

NAND2xp5_ASAP7_75t_L g1904 ( 
.A(n_1897),
.B(n_1879),
.Y(n_1904)
);

OAI221xp5_ASAP7_75t_L g1905 ( 
.A1(n_1882),
.A2(n_1881),
.B1(n_1865),
.B2(n_1861),
.C(n_1873),
.Y(n_1905)
);

OAI22xp33_ASAP7_75t_SL g1906 ( 
.A1(n_1884),
.A2(n_1861),
.B1(n_1878),
.B2(n_1874),
.Y(n_1906)
);

NOR2xp33_ASAP7_75t_L g1907 ( 
.A(n_1883),
.B(n_1779),
.Y(n_1907)
);

OAI22xp33_ASAP7_75t_L g1908 ( 
.A1(n_1890),
.A2(n_1787),
.B1(n_1873),
.B2(n_1870),
.Y(n_1908)
);

INVx2_ASAP7_75t_SL g1909 ( 
.A(n_1889),
.Y(n_1909)
);

NAND2xp5_ASAP7_75t_L g1910 ( 
.A(n_1902),
.B(n_1850),
.Y(n_1910)
);

NAND2xp33_ASAP7_75t_SL g1911 ( 
.A(n_1898),
.B(n_1884),
.Y(n_1911)
);

NAND2xp33_ASAP7_75t_SL g1912 ( 
.A(n_1898),
.B(n_1877),
.Y(n_1912)
);

NAND2xp5_ASAP7_75t_L g1913 ( 
.A(n_1892),
.B(n_1858),
.Y(n_1913)
);

NOR2xp33_ASAP7_75t_L g1914 ( 
.A(n_1886),
.B(n_1779),
.Y(n_1914)
);

OAI22xp33_ASAP7_75t_L g1915 ( 
.A1(n_1891),
.A2(n_1870),
.B1(n_1843),
.B2(n_1837),
.Y(n_1915)
);

INVx1_ASAP7_75t_L g1916 ( 
.A(n_1899),
.Y(n_1916)
);

NOR2xp33_ASAP7_75t_L g1917 ( 
.A(n_1907),
.B(n_1901),
.Y(n_1917)
);

OR2x2_ASAP7_75t_L g1918 ( 
.A(n_1903),
.B(n_1892),
.Y(n_1918)
);

INVx1_ASAP7_75t_SL g1919 ( 
.A(n_1911),
.Y(n_1919)
);

NAND2xp5_ASAP7_75t_L g1920 ( 
.A(n_1916),
.B(n_1888),
.Y(n_1920)
);

OR2x2_ASAP7_75t_L g1921 ( 
.A(n_1904),
.B(n_1893),
.Y(n_1921)
);

NAND2xp5_ASAP7_75t_L g1922 ( 
.A(n_1909),
.B(n_1894),
.Y(n_1922)
);

NOR2xp33_ASAP7_75t_SL g1923 ( 
.A(n_1914),
.B(n_1885),
.Y(n_1923)
);

INVx1_ASAP7_75t_L g1924 ( 
.A(n_1913),
.Y(n_1924)
);

INVx1_ASAP7_75t_L g1925 ( 
.A(n_1910),
.Y(n_1925)
);

NAND2xp5_ASAP7_75t_L g1926 ( 
.A(n_1906),
.B(n_1895),
.Y(n_1926)
);

INVx1_ASAP7_75t_L g1927 ( 
.A(n_1912),
.Y(n_1927)
);

INVx1_ASAP7_75t_L g1928 ( 
.A(n_1908),
.Y(n_1928)
);

INVx2_ASAP7_75t_L g1929 ( 
.A(n_1905),
.Y(n_1929)
);

INVx1_ASAP7_75t_L g1930 ( 
.A(n_1921),
.Y(n_1930)
);

INVx2_ASAP7_75t_L g1931 ( 
.A(n_1922),
.Y(n_1931)
);

INVx1_ASAP7_75t_SL g1932 ( 
.A(n_1919),
.Y(n_1932)
);

AND2x2_ASAP7_75t_L g1933 ( 
.A(n_1927),
.B(n_1896),
.Y(n_1933)
);

INVx3_ASAP7_75t_L g1934 ( 
.A(n_1918),
.Y(n_1934)
);

NAND2x1_ASAP7_75t_SL g1935 ( 
.A(n_1928),
.B(n_1896),
.Y(n_1935)
);

NAND2xp5_ASAP7_75t_L g1936 ( 
.A(n_1929),
.B(n_1915),
.Y(n_1936)
);

INVx1_ASAP7_75t_L g1937 ( 
.A(n_1920),
.Y(n_1937)
);

OAI22xp5_ASAP7_75t_L g1938 ( 
.A1(n_1926),
.A2(n_1887),
.B1(n_1830),
.B2(n_1766),
.Y(n_1938)
);

XNOR2xp5_ASAP7_75t_L g1939 ( 
.A(n_1925),
.B(n_1830),
.Y(n_1939)
);

INVx2_ASAP7_75t_L g1940 ( 
.A(n_1924),
.Y(n_1940)
);

INVx1_ASAP7_75t_L g1941 ( 
.A(n_1933),
.Y(n_1941)
);

AOI222xp33_ASAP7_75t_L g1942 ( 
.A1(n_1934),
.A2(n_1917),
.B1(n_1923),
.B2(n_1611),
.C1(n_1598),
.C2(n_1816),
.Y(n_1942)
);

OAI221xp5_ASAP7_75t_SL g1943 ( 
.A1(n_1932),
.A2(n_1629),
.B1(n_1816),
.B2(n_1869),
.C(n_1739),
.Y(n_1943)
);

OAI22xp33_ASAP7_75t_L g1944 ( 
.A1(n_1936),
.A2(n_1843),
.B1(n_1869),
.B2(n_1679),
.Y(n_1944)
);

OAI33xp33_ASAP7_75t_L g1945 ( 
.A1(n_1937),
.A2(n_1835),
.A3(n_1761),
.B1(n_1799),
.B2(n_1653),
.B3(n_1791),
.Y(n_1945)
);

NAND2xp5_ASAP7_75t_L g1946 ( 
.A(n_1935),
.B(n_1876),
.Y(n_1946)
);

OAI22xp33_ASAP7_75t_L g1947 ( 
.A1(n_1930),
.A2(n_1843),
.B1(n_1654),
.B2(n_1626),
.Y(n_1947)
);

AND2x2_ASAP7_75t_L g1948 ( 
.A(n_1931),
.B(n_1856),
.Y(n_1948)
);

INVx1_ASAP7_75t_L g1949 ( 
.A(n_1940),
.Y(n_1949)
);

NAND2xp5_ASAP7_75t_L g1950 ( 
.A(n_1935),
.B(n_1939),
.Y(n_1950)
);

OAI22xp33_ASAP7_75t_L g1951 ( 
.A1(n_1938),
.A2(n_1843),
.B1(n_1799),
.B2(n_1767),
.Y(n_1951)
);

NAND2xp5_ASAP7_75t_L g1952 ( 
.A(n_1941),
.B(n_1866),
.Y(n_1952)
);

AOI221xp5_ASAP7_75t_L g1953 ( 
.A1(n_1945),
.A2(n_1655),
.B1(n_1738),
.B2(n_1700),
.C(n_1650),
.Y(n_1953)
);

O2A1O1Ixp33_ASAP7_75t_L g1954 ( 
.A1(n_1950),
.A2(n_1718),
.B(n_1643),
.C(n_1728),
.Y(n_1954)
);

OAI21xp5_ASAP7_75t_SL g1955 ( 
.A1(n_1942),
.A2(n_1711),
.B(n_1645),
.Y(n_1955)
);

NAND2xp5_ASAP7_75t_L g1956 ( 
.A(n_1946),
.B(n_1825),
.Y(n_1956)
);

AOI221xp5_ASAP7_75t_L g1957 ( 
.A1(n_1943),
.A2(n_1791),
.B1(n_1571),
.B2(n_1767),
.C(n_1801),
.Y(n_1957)
);

OAI221xp5_ASAP7_75t_SL g1958 ( 
.A1(n_1951),
.A2(n_1944),
.B1(n_1949),
.B2(n_1947),
.C(n_1948),
.Y(n_1958)
);

INVx1_ASAP7_75t_L g1959 ( 
.A(n_1941),
.Y(n_1959)
);

XNOR2xp5_ASAP7_75t_L g1960 ( 
.A(n_1950),
.B(n_1600),
.Y(n_1960)
);

CKINVDCx20_ASAP7_75t_R g1961 ( 
.A(n_1959),
.Y(n_1961)
);

INVx1_ASAP7_75t_L g1962 ( 
.A(n_1952),
.Y(n_1962)
);

INVxp33_ASAP7_75t_SL g1963 ( 
.A(n_1960),
.Y(n_1963)
);

INVxp33_ASAP7_75t_SL g1964 ( 
.A(n_1955),
.Y(n_1964)
);

XNOR2xp5_ASAP7_75t_L g1965 ( 
.A(n_1957),
.B(n_1579),
.Y(n_1965)
);

INVx2_ASAP7_75t_L g1966 ( 
.A(n_1956),
.Y(n_1966)
);

AND2x2_ASAP7_75t_L g1967 ( 
.A(n_1953),
.B(n_1819),
.Y(n_1967)
);

INVx2_ASAP7_75t_L g1968 ( 
.A(n_1958),
.Y(n_1968)
);

INVxp67_ASAP7_75t_L g1969 ( 
.A(n_1954),
.Y(n_1969)
);

INVx1_ASAP7_75t_L g1970 ( 
.A(n_1952),
.Y(n_1970)
);

NOR2xp33_ASAP7_75t_L g1971 ( 
.A(n_1958),
.B(n_1571),
.Y(n_1971)
);

INVx1_ASAP7_75t_SL g1972 ( 
.A(n_1959),
.Y(n_1972)
);

INVx2_ASAP7_75t_L g1973 ( 
.A(n_1959),
.Y(n_1973)
);

AND2x2_ASAP7_75t_L g1974 ( 
.A(n_1971),
.B(n_1839),
.Y(n_1974)
);

NAND4xp75_ASAP7_75t_L g1975 ( 
.A(n_1968),
.B(n_1674),
.C(n_1723),
.D(n_1716),
.Y(n_1975)
);

AND2x2_ASAP7_75t_L g1976 ( 
.A(n_1967),
.B(n_1839),
.Y(n_1976)
);

AOI22xp33_ASAP7_75t_L g1977 ( 
.A1(n_1964),
.A2(n_1963),
.B1(n_1961),
.B2(n_1962),
.Y(n_1977)
);

NOR3xp33_ASAP7_75t_L g1978 ( 
.A(n_1970),
.B(n_1658),
.C(n_1729),
.Y(n_1978)
);

NAND2xp5_ASAP7_75t_L g1979 ( 
.A(n_1972),
.B(n_1973),
.Y(n_1979)
);

INVx1_ASAP7_75t_L g1980 ( 
.A(n_1972),
.Y(n_1980)
);

NAND2xp5_ASAP7_75t_SL g1981 ( 
.A(n_1969),
.B(n_1685),
.Y(n_1981)
);

NAND2xp5_ASAP7_75t_L g1982 ( 
.A(n_1966),
.B(n_1795),
.Y(n_1982)
);

NOR3xp33_ASAP7_75t_L g1983 ( 
.A(n_1979),
.B(n_1965),
.C(n_1712),
.Y(n_1983)
);

NOR3xp33_ASAP7_75t_L g1984 ( 
.A(n_1980),
.B(n_1703),
.C(n_1722),
.Y(n_1984)
);

AOI211xp5_ASAP7_75t_L g1985 ( 
.A1(n_1981),
.A2(n_1727),
.B(n_1671),
.C(n_1685),
.Y(n_1985)
);

OAI321xp33_ASAP7_75t_L g1986 ( 
.A1(n_1977),
.A2(n_1784),
.A3(n_1806),
.B1(n_1803),
.B2(n_1809),
.C(n_1792),
.Y(n_1986)
);

NAND2xp5_ASAP7_75t_L g1987 ( 
.A(n_1976),
.B(n_1774),
.Y(n_1987)
);

AOI221xp5_ASAP7_75t_L g1988 ( 
.A1(n_1974),
.A2(n_1982),
.B1(n_1978),
.B2(n_1975),
.C(n_1705),
.Y(n_1988)
);

OAI211xp5_ASAP7_75t_L g1989 ( 
.A1(n_1977),
.A2(n_1674),
.B(n_1587),
.C(n_1710),
.Y(n_1989)
);

AND2x2_ASAP7_75t_L g1990 ( 
.A(n_1983),
.B(n_1773),
.Y(n_1990)
);

AND2x2_ASAP7_75t_L g1991 ( 
.A(n_1987),
.B(n_1756),
.Y(n_1991)
);

OAI211xp5_ASAP7_75t_L g1992 ( 
.A1(n_1988),
.A2(n_1788),
.B(n_1783),
.C(n_1780),
.Y(n_1992)
);

AOI221xp5_ASAP7_75t_L g1993 ( 
.A1(n_1986),
.A2(n_1705),
.B1(n_1671),
.B2(n_1689),
.C(n_1704),
.Y(n_1993)
);

NOR5xp2_ASAP7_75t_L g1994 ( 
.A(n_1989),
.B(n_1656),
.C(n_1689),
.D(n_1682),
.E(n_1704),
.Y(n_1994)
);

NAND4xp25_ASAP7_75t_L g1995 ( 
.A(n_1984),
.B(n_1635),
.C(n_1759),
.D(n_1796),
.Y(n_1995)
);

NAND4xp75_ASAP7_75t_L g1996 ( 
.A(n_1985),
.B(n_1682),
.C(n_1789),
.D(n_1656),
.Y(n_1996)
);

AOI322xp5_ASAP7_75t_L g1997 ( 
.A1(n_1983),
.A2(n_1656),
.A3(n_1662),
.B1(n_394),
.B2(n_396),
.C1(n_397),
.C2(n_398),
.Y(n_1997)
);

OR3x1_ASAP7_75t_L g1998 ( 
.A(n_1986),
.B(n_392),
.C(n_393),
.Y(n_1998)
);

OAI222xp33_ASAP7_75t_R g1999 ( 
.A1(n_1983),
.A2(n_555),
.B1(n_401),
.B2(n_402),
.C1(n_407),
.C2(n_408),
.Y(n_1999)
);

NAND5xp2_ASAP7_75t_L g2000 ( 
.A(n_1988),
.B(n_399),
.C(n_409),
.D(n_410),
.E(n_411),
.Y(n_2000)
);

NAND2x1p5_ASAP7_75t_L g2001 ( 
.A(n_1990),
.B(n_413),
.Y(n_2001)
);

OAI211xp5_ASAP7_75t_L g2002 ( 
.A1(n_1992),
.A2(n_414),
.B(n_417),
.C(n_418),
.Y(n_2002)
);

INVx1_ASAP7_75t_L g2003 ( 
.A(n_1998),
.Y(n_2003)
);

NAND5xp2_ASAP7_75t_L g2004 ( 
.A(n_1991),
.B(n_1997),
.C(n_1999),
.D(n_2000),
.E(n_1993),
.Y(n_2004)
);

HB1xp67_ASAP7_75t_L g2005 ( 
.A(n_1996),
.Y(n_2005)
);

AND2x4_ASAP7_75t_L g2006 ( 
.A(n_1995),
.B(n_419),
.Y(n_2006)
);

NOR2xp67_ASAP7_75t_SL g2007 ( 
.A(n_1994),
.B(n_420),
.Y(n_2007)
);

AND3x2_ASAP7_75t_L g2008 ( 
.A(n_1999),
.B(n_422),
.C(n_423),
.Y(n_2008)
);

INVx2_ASAP7_75t_L g2009 ( 
.A(n_1996),
.Y(n_2009)
);

OA22x2_ASAP7_75t_L g2010 ( 
.A1(n_1992),
.A2(n_424),
.B1(n_425),
.B2(n_426),
.Y(n_2010)
);

NOR3xp33_ASAP7_75t_SL g2011 ( 
.A(n_2000),
.B(n_554),
.C(n_427),
.Y(n_2011)
);

NAND4xp75_ASAP7_75t_L g2012 ( 
.A(n_1990),
.B(n_428),
.C(n_429),
.D(n_431),
.Y(n_2012)
);

INVxp67_ASAP7_75t_L g2013 ( 
.A(n_2000),
.Y(n_2013)
);

INVx2_ASAP7_75t_L g2014 ( 
.A(n_1996),
.Y(n_2014)
);

NOR3xp33_ASAP7_75t_SL g2015 ( 
.A(n_2003),
.B(n_2002),
.C(n_2004),
.Y(n_2015)
);

OA22x2_ASAP7_75t_L g2016 ( 
.A1(n_2008),
.A2(n_432),
.B1(n_434),
.B2(n_435),
.Y(n_2016)
);

NAND2xp33_ASAP7_75t_SL g2017 ( 
.A(n_2007),
.B(n_553),
.Y(n_2017)
);

CKINVDCx20_ASAP7_75t_R g2018 ( 
.A(n_2013),
.Y(n_2018)
);

XNOR2xp5_ASAP7_75t_L g2019 ( 
.A(n_2011),
.B(n_437),
.Y(n_2019)
);

OR2x2_ASAP7_75t_L g2020 ( 
.A(n_2001),
.B(n_438),
.Y(n_2020)
);

NAND2xp5_ASAP7_75t_L g2021 ( 
.A(n_2006),
.B(n_439),
.Y(n_2021)
);

NAND2xp5_ASAP7_75t_L g2022 ( 
.A(n_2005),
.B(n_440),
.Y(n_2022)
);

INVx2_ASAP7_75t_L g2023 ( 
.A(n_2012),
.Y(n_2023)
);

AOI22xp5_ASAP7_75t_L g2024 ( 
.A1(n_2009),
.A2(n_441),
.B1(n_442),
.B2(n_443),
.Y(n_2024)
);

NAND2xp5_ASAP7_75t_L g2025 ( 
.A(n_2014),
.B(n_444),
.Y(n_2025)
);

INVxp67_ASAP7_75t_SL g2026 ( 
.A(n_2010),
.Y(n_2026)
);

HB1xp67_ASAP7_75t_L g2027 ( 
.A(n_2001),
.Y(n_2027)
);

INVx2_ASAP7_75t_L g2028 ( 
.A(n_2001),
.Y(n_2028)
);

NAND4xp75_ASAP7_75t_L g2029 ( 
.A(n_2003),
.B(n_445),
.C(n_447),
.D(n_449),
.Y(n_2029)
);

OR2x2_ASAP7_75t_L g2030 ( 
.A(n_2004),
.B(n_451),
.Y(n_2030)
);

INVx1_ASAP7_75t_L g2031 ( 
.A(n_2003),
.Y(n_2031)
);

NOR2x1_ASAP7_75t_L g2032 ( 
.A(n_2012),
.B(n_452),
.Y(n_2032)
);

INVx1_ASAP7_75t_SL g2033 ( 
.A(n_2020),
.Y(n_2033)
);

INVx2_ASAP7_75t_L g2034 ( 
.A(n_2029),
.Y(n_2034)
);

INVx1_ASAP7_75t_SL g2035 ( 
.A(n_2017),
.Y(n_2035)
);

INVx2_ASAP7_75t_L g2036 ( 
.A(n_2028),
.Y(n_2036)
);

INVx2_ASAP7_75t_L g2037 ( 
.A(n_2030),
.Y(n_2037)
);

AOI222xp33_ASAP7_75t_L g2038 ( 
.A1(n_2031),
.A2(n_453),
.B1(n_454),
.B2(n_456),
.C1(n_458),
.C2(n_460),
.Y(n_2038)
);

INVx2_ASAP7_75t_L g2039 ( 
.A(n_2019),
.Y(n_2039)
);

OAI211xp5_ASAP7_75t_L g2040 ( 
.A1(n_2026),
.A2(n_2022),
.B(n_2025),
.C(n_2032),
.Y(n_2040)
);

NAND2xp5_ASAP7_75t_L g2041 ( 
.A(n_2027),
.B(n_461),
.Y(n_2041)
);

HB1xp67_ASAP7_75t_L g2042 ( 
.A(n_2016),
.Y(n_2042)
);

BUFx2_ASAP7_75t_L g2043 ( 
.A(n_2018),
.Y(n_2043)
);

AOI22xp5_ASAP7_75t_L g2044 ( 
.A1(n_2023),
.A2(n_462),
.B1(n_463),
.B2(n_464),
.Y(n_2044)
);

XNOR2xp5_ASAP7_75t_L g2045 ( 
.A(n_2015),
.B(n_465),
.Y(n_2045)
);

AOI22xp5_ASAP7_75t_L g2046 ( 
.A1(n_2043),
.A2(n_2021),
.B1(n_2024),
.B2(n_470),
.Y(n_2046)
);

AO22x2_ASAP7_75t_L g2047 ( 
.A1(n_2036),
.A2(n_466),
.B1(n_467),
.B2(n_471),
.Y(n_2047)
);

OR2x2_ASAP7_75t_L g2048 ( 
.A(n_2037),
.B(n_2035),
.Y(n_2048)
);

INVx1_ASAP7_75t_L g2049 ( 
.A(n_2045),
.Y(n_2049)
);

BUFx2_ASAP7_75t_L g2050 ( 
.A(n_2042),
.Y(n_2050)
);

INVx1_ASAP7_75t_L g2051 ( 
.A(n_2041),
.Y(n_2051)
);

OAI22xp33_ASAP7_75t_L g2052 ( 
.A1(n_2034),
.A2(n_472),
.B1(n_474),
.B2(n_475),
.Y(n_2052)
);

OAI22x1_ASAP7_75t_L g2053 ( 
.A1(n_2033),
.A2(n_476),
.B1(n_477),
.B2(n_478),
.Y(n_2053)
);

AOI31xp33_ASAP7_75t_L g2054 ( 
.A1(n_2040),
.A2(n_552),
.A3(n_480),
.B(n_482),
.Y(n_2054)
);

AOI21xp33_ASAP7_75t_SL g2055 ( 
.A1(n_2054),
.A2(n_2039),
.B(n_2038),
.Y(n_2055)
);

OAI22xp5_ASAP7_75t_L g2056 ( 
.A1(n_2050),
.A2(n_2044),
.B1(n_483),
.B2(n_484),
.Y(n_2056)
);

OAI22xp5_ASAP7_75t_SL g2057 ( 
.A1(n_2049),
.A2(n_479),
.B1(n_485),
.B2(n_486),
.Y(n_2057)
);

AOI22xp5_ASAP7_75t_L g2058 ( 
.A1(n_2046),
.A2(n_551),
.B1(n_493),
.B2(n_494),
.Y(n_2058)
);

OAI22xp5_ASAP7_75t_L g2059 ( 
.A1(n_2058),
.A2(n_2048),
.B1(n_2051),
.B2(n_2052),
.Y(n_2059)
);

OAI22xp5_ASAP7_75t_SL g2060 ( 
.A1(n_2057),
.A2(n_2053),
.B1(n_2047),
.B2(n_496),
.Y(n_2060)
);

INVx1_ASAP7_75t_L g2061 ( 
.A(n_2060),
.Y(n_2061)
);

INVx1_ASAP7_75t_L g2062 ( 
.A(n_2059),
.Y(n_2062)
);

INVx1_ASAP7_75t_L g2063 ( 
.A(n_2062),
.Y(n_2063)
);

AOI21xp5_ASAP7_75t_L g2064 ( 
.A1(n_2061),
.A2(n_2055),
.B(n_2056),
.Y(n_2064)
);

AOI22xp33_ASAP7_75t_L g2065 ( 
.A1(n_2063),
.A2(n_2047),
.B1(n_495),
.B2(n_497),
.Y(n_2065)
);

AOI22xp33_ASAP7_75t_L g2066 ( 
.A1(n_2064),
.A2(n_490),
.B1(n_498),
.B2(n_499),
.Y(n_2066)
);

NAND2xp5_ASAP7_75t_SL g2067 ( 
.A(n_2065),
.B(n_2066),
.Y(n_2067)
);

AOI21xp5_ASAP7_75t_L g2068 ( 
.A1(n_2065),
.A2(n_501),
.B(n_502),
.Y(n_2068)
);

OR2x6_ASAP7_75t_L g2069 ( 
.A(n_2067),
.B(n_506),
.Y(n_2069)
);

OR2x6_ASAP7_75t_L g2070 ( 
.A(n_2068),
.B(n_507),
.Y(n_2070)
);

AOI221xp5_ASAP7_75t_L g2071 ( 
.A1(n_2070),
.A2(n_509),
.B1(n_510),
.B2(n_512),
.C(n_514),
.Y(n_2071)
);

AOI211xp5_ASAP7_75t_L g2072 ( 
.A1(n_2071),
.A2(n_2069),
.B(n_516),
.C(n_517),
.Y(n_2072)
);


endmodule