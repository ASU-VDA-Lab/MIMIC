module fake_netlist_6_2431_n_873 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_161, n_68, n_166, n_28, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_178, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_180, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_181, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_175, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_104, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_173, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_171, n_31, n_57, n_169, n_53, n_51, n_44, n_56, n_873);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_161;
input n_68;
input n_166;
input n_28;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_178;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_181;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_175;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_104;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_173;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_171;
input n_31;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_873;

wire n_591;
wire n_435;
wire n_793;
wire n_326;
wire n_801;
wire n_256;
wire n_853;
wire n_440;
wire n_587;
wire n_695;
wire n_507;
wire n_580;
wire n_762;
wire n_209;
wire n_367;
wire n_465;
wire n_680;
wire n_741;
wire n_760;
wire n_590;
wire n_625;
wire n_661;
wire n_223;
wire n_278;
wire n_341;
wire n_362;
wire n_226;
wire n_828;
wire n_208;
wire n_462;
wire n_607;
wire n_671;
wire n_726;
wire n_316;
wire n_419;
wire n_304;
wire n_212;
wire n_700;
wire n_694;
wire n_740;
wire n_578;
wire n_703;
wire n_365;
wire n_384;
wire n_297;
wire n_595;
wire n_627;
wire n_524;
wire n_342;
wire n_820;
wire n_783;
wire n_725;
wire n_358;
wire n_751;
wire n_449;
wire n_749;
wire n_798;
wire n_188;
wire n_310;
wire n_509;
wire n_186;
wire n_245;
wire n_368;
wire n_575;
wire n_677;
wire n_805;
wire n_396;
wire n_495;
wire n_815;
wire n_350;
wire n_585;
wire n_732;
wire n_568;
wire n_392;
wire n_840;
wire n_442;
wire n_480;
wire n_724;
wire n_382;
wire n_673;
wire n_628;
wire n_557;
wire n_823;
wire n_349;
wire n_643;
wire n_233;
wire n_617;
wire n_698;
wire n_845;
wire n_255;
wire n_807;
wire n_739;
wire n_284;
wire n_400;
wire n_337;
wire n_865;
wire n_214;
wire n_485;
wire n_443;
wire n_246;
wire n_768;
wire n_471;
wire n_289;
wire n_421;
wire n_781;
wire n_424;
wire n_789;
wire n_615;
wire n_182;
wire n_238;
wire n_573;
wire n_769;
wire n_202;
wire n_320;
wire n_639;
wire n_676;
wire n_327;
wire n_794;
wire n_727;
wire n_369;
wire n_597;
wire n_685;
wire n_280;
wire n_287;
wire n_832;
wire n_353;
wire n_610;
wire n_555;
wire n_389;
wire n_814;
wire n_415;
wire n_830;
wire n_230;
wire n_605;
wire n_461;
wire n_383;
wire n_826;
wire n_669;
wire n_200;
wire n_447;
wire n_872;
wire n_198;
wire n_222;
wire n_300;
wire n_248;
wire n_517;
wire n_718;
wire n_747;
wire n_852;
wire n_667;
wire n_229;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_621;
wire n_305;
wire n_721;
wire n_750;
wire n_532;
wire n_742;
wire n_535;
wire n_691;
wire n_250;
wire n_372;
wire n_468;
wire n_544;
wire n_504;
wire n_314;
wire n_378;
wire n_413;
wire n_377;
wire n_791;
wire n_183;
wire n_510;
wire n_837;
wire n_836;
wire n_863;
wire n_375;
wire n_601;
wire n_338;
wire n_522;
wire n_466;
wire n_704;
wire n_748;
wire n_506;
wire n_763;
wire n_360;
wire n_603;
wire n_235;
wire n_536;
wire n_866;
wire n_622;
wire n_191;
wire n_340;
wire n_710;
wire n_387;
wire n_452;
wire n_616;
wire n_658;
wire n_744;
wire n_344;
wire n_581;
wire n_428;
wire n_761;
wire n_785;
wire n_746;
wire n_609;
wire n_765;
wire n_432;
wire n_641;
wire n_822;
wire n_693;
wire n_631;
wire n_516;
wire n_720;
wire n_758;
wire n_525;
wire n_842;
wire n_611;
wire n_491;
wire n_656;
wire n_772;
wire n_843;
wire n_797;
wire n_666;
wire n_371;
wire n_795;
wire n_770;
wire n_567;
wire n_189;
wire n_738;
wire n_405;
wire n_213;
wire n_538;
wire n_294;
wire n_302;
wire n_499;
wire n_380;
wire n_838;
wire n_705;
wire n_647;
wire n_197;
wire n_343;
wire n_844;
wire n_448;
wire n_494;
wire n_539;
wire n_493;
wire n_397;
wire n_614;
wire n_529;
wire n_445;
wire n_425;
wire n_684;
wire n_454;
wire n_218;
wire n_638;
wire n_234;
wire n_486;
wire n_381;
wire n_236;
wire n_653;
wire n_752;
wire n_713;
wire n_648;
wire n_657;
wire n_576;
wire n_472;
wire n_270;
wire n_239;
wire n_414;
wire n_563;
wire n_782;
wire n_490;
wire n_803;
wire n_290;
wire n_220;
wire n_809;
wire n_224;
wire n_839;
wire n_734;
wire n_708;
wire n_196;
wire n_402;
wire n_352;
wire n_668;
wire n_478;
wire n_626;
wire n_574;
wire n_779;
wire n_800;
wire n_460;
wire n_854;
wire n_417;
wire n_446;
wire n_498;
wire n_662;
wire n_374;
wire n_659;
wire n_709;
wire n_870;
wire n_366;
wire n_777;
wire n_407;
wire n_450;
wire n_808;
wire n_867;
wire n_272;
wire n_526;
wire n_185;
wire n_712;
wire n_348;
wire n_711;
wire n_579;
wire n_376;
wire n_390;
wire n_473;
wire n_293;
wire n_334;
wire n_559;
wire n_370;
wire n_458;
wire n_232;
wire n_650;
wire n_717;
wire n_330;
wire n_771;
wire n_470;
wire n_475;
wire n_298;
wire n_492;
wire n_281;
wire n_258;
wire n_551;
wire n_699;
wire n_456;
wire n_564;
wire n_260;
wire n_265;
wire n_313;
wire n_451;
wire n_624;
wire n_824;
wire n_279;
wire n_686;
wire n_796;
wire n_252;
wire n_757;
wire n_228;
wire n_565;
wire n_594;
wire n_719;
wire n_356;
wire n_577;
wire n_184;
wire n_552;
wire n_619;
wire n_216;
wire n_455;
wire n_521;
wire n_363;
wire n_572;
wire n_395;
wire n_813;
wire n_592;
wire n_745;
wire n_654;
wire n_323;
wire n_829;
wire n_606;
wire n_393;
wire n_818;
wire n_411;
wire n_503;
wire n_716;
wire n_623;
wire n_599;
wire n_513;
wire n_855;
wire n_776;
wire n_321;
wire n_645;
wire n_331;
wire n_227;
wire n_868;
wire n_570;
wire n_731;
wire n_859;
wire n_406;
wire n_483;
wire n_735;
wire n_204;
wire n_482;
wire n_755;
wire n_527;
wire n_474;
wire n_261;
wire n_608;
wire n_620;
wire n_420;
wire n_683;
wire n_630;
wire n_312;
wire n_394;
wire n_519;
wire n_541;
wire n_512;
wire n_292;
wire n_307;
wire n_469;
wire n_433;
wire n_500;
wire n_792;
wire n_476;
wire n_714;
wire n_291;
wire n_219;
wire n_543;
wire n_357;
wire n_264;
wire n_263;
wire n_589;
wire n_860;
wire n_481;
wire n_788;
wire n_819;
wire n_821;
wire n_325;
wire n_767;
wire n_804;
wire n_329;
wire n_464;
wire n_600;
wire n_831;
wire n_802;
wire n_561;
wire n_477;
wire n_549;
wire n_533;
wire n_408;
wire n_806;
wire n_864;
wire n_237;
wire n_584;
wire n_244;
wire n_399;
wire n_243;
wire n_548;
wire n_282;
wire n_436;
wire n_833;
wire n_211;
wire n_523;
wire n_322;
wire n_707;
wire n_345;
wire n_409;
wire n_231;
wire n_354;
wire n_689;
wire n_799;
wire n_505;
wire n_240;
wire n_756;
wire n_319;
wire n_547;
wire n_537;
wire n_273;
wire n_558;
wire n_810;
wire n_635;
wire n_787;
wire n_311;
wire n_403;
wire n_723;
wire n_253;
wire n_634;
wire n_583;
wire n_596;
wire n_546;
wire n_562;
wire n_249;
wire n_201;
wire n_386;
wire n_764;
wire n_556;
wire n_692;
wire n_733;
wire n_754;
wire n_487;
wire n_550;
wire n_241;
wire n_275;
wire n_553;
wire n_652;
wire n_849;
wire n_560;
wire n_753;
wire n_642;
wire n_276;
wire n_569;
wire n_441;
wire n_221;
wire n_811;
wire n_444;
wire n_586;
wire n_423;
wire n_737;
wire n_318;
wire n_303;
wire n_511;
wire n_715;
wire n_467;
wire n_306;
wire n_193;
wire n_269;
wire n_359;
wire n_346;
wire n_416;
wire n_530;
wire n_277;
wire n_520;
wire n_418;
wire n_618;
wire n_790;
wire n_582;
wire n_199;
wire n_266;
wire n_296;
wire n_861;
wire n_674;
wire n_857;
wire n_871;
wire n_775;
wire n_571;
wire n_268;
wire n_271;
wire n_404;
wire n_651;
wire n_439;
wire n_217;
wire n_210;
wire n_299;
wire n_518;
wire n_206;
wire n_679;
wire n_453;
wire n_612;
wire n_633;
wire n_665;
wire n_333;
wire n_588;
wire n_215;
wire n_247;
wire n_225;
wire n_308;
wire n_309;
wire n_759;
wire n_355;
wire n_426;
wire n_317;
wire n_632;
wire n_702;
wire n_431;
wire n_347;
wire n_812;
wire n_459;
wire n_502;
wire n_328;
wire n_672;
wire n_534;
wire n_488;
wire n_429;
wire n_373;
wire n_195;
wire n_497;
wire n_285;
wire n_780;
wire n_773;
wire n_675;
wire n_257;
wire n_730;
wire n_655;
wire n_706;
wire n_786;
wire n_670;
wire n_286;
wire n_203;
wire n_254;
wire n_207;
wire n_834;
wire n_242;
wire n_835;
wire n_690;
wire n_850;
wire n_401;
wire n_324;
wire n_743;
wire n_766;
wire n_816;
wire n_335;
wire n_430;
wire n_463;
wire n_545;
wire n_489;
wire n_205;
wire n_604;
wire n_848;
wire n_251;
wire n_301;
wire n_274;
wire n_636;
wire n_825;
wire n_728;
wire n_681;
wire n_729;
wire n_774;
wire n_412;
wire n_640;
wire n_660;
wire n_267;
wire n_438;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_515;
wire n_288;
wire n_427;
wire n_479;
wire n_598;
wire n_496;
wire n_422;
wire n_696;
wire n_688;
wire n_722;
wire n_862;
wire n_351;
wire n_869;
wire n_437;
wire n_259;
wire n_540;
wire n_593;
wire n_514;
wire n_646;
wire n_528;
wire n_391;
wire n_457;
wire n_687;
wire n_697;
wire n_364;
wire n_637;
wire n_295;
wire n_385;
wire n_701;
wire n_817;
wire n_629;
wire n_388;
wire n_190;
wire n_858;
wire n_262;
wire n_484;
wire n_613;
wire n_736;
wire n_187;
wire n_846;
wire n_501;
wire n_841;
wire n_531;
wire n_827;
wire n_361;
wire n_508;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_332;
wire n_336;
wire n_398;
wire n_410;
wire n_566;
wire n_554;
wire n_602;
wire n_194;
wire n_664;
wire n_678;
wire n_192;
wire n_649;
wire n_283;

INVx1_ASAP7_75t_L g182 ( 
.A(n_83),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_181),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_173),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_134),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_27),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_18),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_8),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_22),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_96),
.Y(n_190)
);

BUFx3_ASAP7_75t_L g191 ( 
.A(n_104),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_68),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_32),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_30),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_112),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_165),
.Y(n_196)
);

BUFx6f_ASAP7_75t_L g197 ( 
.A(n_9),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_109),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_73),
.Y(n_199)
);

CKINVDCx14_ASAP7_75t_R g200 ( 
.A(n_148),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_174),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_82),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_84),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_62),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_124),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_151),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_125),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_152),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_114),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_2),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_72),
.Y(n_211)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_180),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_51),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_85),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_10),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_177),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_156),
.Y(n_217)
);

BUFx3_ASAP7_75t_L g218 ( 
.A(n_158),
.Y(n_218)
);

BUFx3_ASAP7_75t_L g219 ( 
.A(n_36),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_175),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_113),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_2),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_92),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_117),
.Y(n_224)
);

CKINVDCx16_ASAP7_75t_R g225 ( 
.A(n_127),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_172),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_128),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_166),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_119),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_31),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_57),
.Y(n_231)
);

INVx1_ASAP7_75t_SL g232 ( 
.A(n_44),
.Y(n_232)
);

BUFx6f_ASAP7_75t_L g233 ( 
.A(n_26),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_139),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_28),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_176),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_78),
.Y(n_237)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_41),
.Y(n_238)
);

INVxp67_ASAP7_75t_SL g239 ( 
.A(n_131),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_130),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_4),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_162),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_43),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_150),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_50),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_100),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_65),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_22),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_21),
.Y(n_249)
);

INVx1_ASAP7_75t_SL g250 ( 
.A(n_90),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_138),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_107),
.Y(n_252)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_63),
.Y(n_253)
);

BUFx6f_ASAP7_75t_L g254 ( 
.A(n_146),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_47),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_6),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_46),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_197),
.Y(n_258)
);

INVx2_ASAP7_75t_SL g259 ( 
.A(n_197),
.Y(n_259)
);

BUFx6f_ASAP7_75t_L g260 ( 
.A(n_254),
.Y(n_260)
);

HB1xp67_ASAP7_75t_L g261 ( 
.A(n_186),
.Y(n_261)
);

HB1xp67_ASAP7_75t_L g262 ( 
.A(n_215),
.Y(n_262)
);

BUFx2_ASAP7_75t_L g263 ( 
.A(n_241),
.Y(n_263)
);

BUFx6f_ASAP7_75t_L g264 ( 
.A(n_254),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_SL g265 ( 
.A(n_225),
.B(n_0),
.Y(n_265)
);

AND2x2_ASAP7_75t_L g266 ( 
.A(n_200),
.B(n_0),
.Y(n_266)
);

BUFx6f_ASAP7_75t_L g267 ( 
.A(n_254),
.Y(n_267)
);

AND2x4_ASAP7_75t_L g268 ( 
.A(n_191),
.B(n_29),
.Y(n_268)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_197),
.Y(n_269)
);

HB1xp67_ASAP7_75t_L g270 ( 
.A(n_248),
.Y(n_270)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_197),
.Y(n_271)
);

AND2x6_ASAP7_75t_L g272 ( 
.A(n_254),
.B(n_33),
.Y(n_272)
);

BUFx12f_ASAP7_75t_L g273 ( 
.A(n_249),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_212),
.B(n_1),
.Y(n_274)
);

BUFx6f_ASAP7_75t_L g275 ( 
.A(n_191),
.Y(n_275)
);

BUFx8_ASAP7_75t_L g276 ( 
.A(n_233),
.Y(n_276)
);

AND2x4_ASAP7_75t_L g277 ( 
.A(n_218),
.B(n_34),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_212),
.B(n_1),
.Y(n_278)
);

BUFx2_ASAP7_75t_L g279 ( 
.A(n_256),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_238),
.B(n_3),
.Y(n_280)
);

INVx4_ASAP7_75t_L g281 ( 
.A(n_218),
.Y(n_281)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_233),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_SL g283 ( 
.A(n_233),
.B(n_3),
.Y(n_283)
);

INVx5_ASAP7_75t_L g284 ( 
.A(n_219),
.Y(n_284)
);

BUFx6f_ASAP7_75t_L g285 ( 
.A(n_219),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_238),
.B(n_4),
.Y(n_286)
);

AND2x2_ASAP7_75t_L g287 ( 
.A(n_200),
.B(n_5),
.Y(n_287)
);

BUFx6f_ASAP7_75t_L g288 ( 
.A(n_253),
.Y(n_288)
);

BUFx6f_ASAP7_75t_L g289 ( 
.A(n_253),
.Y(n_289)
);

AND2x2_ASAP7_75t_L g290 ( 
.A(n_233),
.B(n_5),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_232),
.B(n_6),
.Y(n_291)
);

BUFx6f_ASAP7_75t_L g292 ( 
.A(n_182),
.Y(n_292)
);

BUFx3_ASAP7_75t_L g293 ( 
.A(n_185),
.Y(n_293)
);

BUFx8_ASAP7_75t_L g294 ( 
.A(n_193),
.Y(n_294)
);

INVx5_ASAP7_75t_L g295 ( 
.A(n_239),
.Y(n_295)
);

BUFx3_ASAP7_75t_L g296 ( 
.A(n_195),
.Y(n_296)
);

BUFx6f_ASAP7_75t_L g297 ( 
.A(n_199),
.Y(n_297)
);

BUFx6f_ASAP7_75t_L g298 ( 
.A(n_201),
.Y(n_298)
);

HB1xp67_ASAP7_75t_L g299 ( 
.A(n_187),
.Y(n_299)
);

AND2x4_ASAP7_75t_L g300 ( 
.A(n_205),
.B(n_35),
.Y(n_300)
);

AND2x4_ASAP7_75t_L g301 ( 
.A(n_206),
.B(n_37),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_250),
.B(n_7),
.Y(n_302)
);

INVx5_ASAP7_75t_L g303 ( 
.A(n_183),
.Y(n_303)
);

HB1xp67_ASAP7_75t_L g304 ( 
.A(n_188),
.Y(n_304)
);

AND2x4_ASAP7_75t_L g305 ( 
.A(n_217),
.B(n_38),
.Y(n_305)
);

AND2x2_ASAP7_75t_L g306 ( 
.A(n_189),
.B(n_7),
.Y(n_306)
);

INVx2_ASAP7_75t_L g307 ( 
.A(n_210),
.Y(n_307)
);

INVx4_ASAP7_75t_L g308 ( 
.A(n_184),
.Y(n_308)
);

AND2x4_ASAP7_75t_L g309 ( 
.A(n_223),
.B(n_39),
.Y(n_309)
);

INVx3_ASAP7_75t_L g310 ( 
.A(n_260),
.Y(n_310)
);

OAI22xp33_ASAP7_75t_SL g311 ( 
.A1(n_265),
.A2(n_224),
.B1(n_229),
.B2(n_231),
.Y(n_311)
);

OAI22xp33_ASAP7_75t_SL g312 ( 
.A1(n_283),
.A2(n_240),
.B1(n_243),
.B2(n_245),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_L g313 ( 
.A1(n_266),
.A2(n_230),
.B1(n_235),
.B2(n_228),
.Y(n_313)
);

INVx1_ASAP7_75t_SL g314 ( 
.A(n_263),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_258),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_308),
.B(n_190),
.Y(n_316)
);

OAI22xp33_ASAP7_75t_SL g317 ( 
.A1(n_283),
.A2(n_257),
.B1(n_255),
.B2(n_252),
.Y(n_317)
);

AO22x2_ASAP7_75t_L g318 ( 
.A1(n_266),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_SL g319 ( 
.A1(n_291),
.A2(n_222),
.B1(n_230),
.B2(n_235),
.Y(n_319)
);

AND2x2_ASAP7_75t_L g320 ( 
.A(n_261),
.B(n_192),
.Y(n_320)
);

INVx2_ASAP7_75t_L g321 ( 
.A(n_269),
.Y(n_321)
);

AO22x2_ASAP7_75t_L g322 ( 
.A1(n_287),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_322)
);

OAI22xp5_ASAP7_75t_SL g323 ( 
.A1(n_302),
.A2(n_211),
.B1(n_246),
.B2(n_247),
.Y(n_323)
);

INVxp33_ASAP7_75t_L g324 ( 
.A(n_262),
.Y(n_324)
);

OAI22xp33_ASAP7_75t_R g325 ( 
.A1(n_270),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_325)
);

BUFx10_ASAP7_75t_L g326 ( 
.A(n_274),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_269),
.Y(n_327)
);

AO22x2_ASAP7_75t_L g328 ( 
.A1(n_287),
.A2(n_14),
.B1(n_15),
.B2(n_16),
.Y(n_328)
);

AOI22xp5_ASAP7_75t_L g329 ( 
.A1(n_273),
.A2(n_251),
.B1(n_244),
.B2(n_242),
.Y(n_329)
);

INVx3_ASAP7_75t_L g330 ( 
.A(n_260),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_271),
.Y(n_331)
);

OAI22xp33_ASAP7_75t_SL g332 ( 
.A1(n_268),
.A2(n_237),
.B1(n_236),
.B2(n_234),
.Y(n_332)
);

INVx2_ASAP7_75t_L g333 ( 
.A(n_271),
.Y(n_333)
);

AND2x4_ASAP7_75t_L g334 ( 
.A(n_268),
.B(n_194),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_308),
.B(n_196),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_282),
.Y(n_336)
);

AOI22xp5_ASAP7_75t_L g337 ( 
.A1(n_273),
.A2(n_227),
.B1(n_226),
.B2(n_221),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_282),
.Y(n_338)
);

INVx2_ASAP7_75t_L g339 ( 
.A(n_260),
.Y(n_339)
);

INVx2_ASAP7_75t_L g340 ( 
.A(n_260),
.Y(n_340)
);

AND2x2_ASAP7_75t_L g341 ( 
.A(n_263),
.B(n_198),
.Y(n_341)
);

OAI22xp5_ASAP7_75t_SL g342 ( 
.A1(n_279),
.A2(n_220),
.B1(n_216),
.B2(n_214),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_288),
.Y(n_343)
);

OAI22xp33_ASAP7_75t_L g344 ( 
.A1(n_278),
.A2(n_286),
.B1(n_279),
.B2(n_299),
.Y(n_344)
);

OAI22xp5_ASAP7_75t_L g345 ( 
.A1(n_280),
.A2(n_277),
.B1(n_268),
.B2(n_306),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_288),
.Y(n_346)
);

OAI22xp33_ASAP7_75t_R g347 ( 
.A1(n_304),
.A2(n_14),
.B1(n_15),
.B2(n_16),
.Y(n_347)
);

AOI22xp5_ASAP7_75t_L g348 ( 
.A1(n_277),
.A2(n_213),
.B1(n_209),
.B2(n_208),
.Y(n_348)
);

OAI22xp33_ASAP7_75t_SL g349 ( 
.A1(n_277),
.A2(n_207),
.B1(n_204),
.B2(n_203),
.Y(n_349)
);

INVx2_ASAP7_75t_L g350 ( 
.A(n_267),
.Y(n_350)
);

AOI22xp5_ASAP7_75t_L g351 ( 
.A1(n_300),
.A2(n_202),
.B1(n_18),
.B2(n_19),
.Y(n_351)
);

AO22x2_ASAP7_75t_L g352 ( 
.A1(n_290),
.A2(n_17),
.B1(n_19),
.B2(n_20),
.Y(n_352)
);

AO22x2_ASAP7_75t_L g353 ( 
.A1(n_290),
.A2(n_17),
.B1(n_20),
.B2(n_21),
.Y(n_353)
);

AOI22xp5_ASAP7_75t_L g354 ( 
.A1(n_300),
.A2(n_23),
.B1(n_24),
.B2(n_25),
.Y(n_354)
);

AO22x2_ASAP7_75t_L g355 ( 
.A1(n_306),
.A2(n_23),
.B1(n_24),
.B2(n_25),
.Y(n_355)
);

OAI22xp33_ASAP7_75t_L g356 ( 
.A1(n_281),
.A2(n_26),
.B1(n_27),
.B2(n_40),
.Y(n_356)
);

OAI22xp33_ASAP7_75t_SL g357 ( 
.A1(n_281),
.A2(n_42),
.B1(n_45),
.B2(n_48),
.Y(n_357)
);

AO22x2_ASAP7_75t_L g358 ( 
.A1(n_300),
.A2(n_49),
.B1(n_52),
.B2(n_53),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_288),
.Y(n_359)
);

INVx2_ASAP7_75t_L g360 ( 
.A(n_267),
.Y(n_360)
);

AOI22x1_ASAP7_75t_SL g361 ( 
.A1(n_281),
.A2(n_54),
.B1(n_55),
.B2(n_56),
.Y(n_361)
);

AND2x2_ASAP7_75t_L g362 ( 
.A(n_308),
.B(n_58),
.Y(n_362)
);

INVx2_ASAP7_75t_L g363 ( 
.A(n_267),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_L g364 ( 
.A(n_301),
.B(n_59),
.Y(n_364)
);

AOI22xp5_ASAP7_75t_L g365 ( 
.A1(n_301),
.A2(n_60),
.B1(n_61),
.B2(n_64),
.Y(n_365)
);

XOR2xp5_ASAP7_75t_L g366 ( 
.A(n_313),
.B(n_301),
.Y(n_366)
);

INVx2_ASAP7_75t_L g367 ( 
.A(n_310),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_343),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_346),
.Y(n_369)
);

AND2x6_ASAP7_75t_L g370 ( 
.A(n_364),
.B(n_305),
.Y(n_370)
);

NOR2xp33_ASAP7_75t_L g371 ( 
.A(n_345),
.B(n_275),
.Y(n_371)
);

INVxp33_ASAP7_75t_L g372 ( 
.A(n_324),
.Y(n_372)
);

AND2x4_ASAP7_75t_L g373 ( 
.A(n_334),
.B(n_305),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_359),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_310),
.Y(n_375)
);

CKINVDCx20_ASAP7_75t_R g376 ( 
.A(n_314),
.Y(n_376)
);

AND2x4_ASAP7_75t_L g377 ( 
.A(n_334),
.B(n_305),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_SL g378 ( 
.A(n_317),
.B(n_309),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_330),
.Y(n_379)
);

INVxp33_ASAP7_75t_L g380 ( 
.A(n_319),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_330),
.Y(n_381)
);

INVxp67_ASAP7_75t_L g382 ( 
.A(n_341),
.Y(n_382)
);

NOR2xp33_ASAP7_75t_L g383 ( 
.A(n_344),
.B(n_275),
.Y(n_383)
);

AND2x2_ASAP7_75t_L g384 ( 
.A(n_320),
.B(n_293),
.Y(n_384)
);

NAND2x1p5_ASAP7_75t_L g385 ( 
.A(n_365),
.B(n_309),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_342),
.Y(n_386)
);

INVx2_ASAP7_75t_L g387 ( 
.A(n_339),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_315),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_SL g389 ( 
.A(n_311),
.B(n_309),
.Y(n_389)
);

NOR2xp33_ASAP7_75t_L g390 ( 
.A(n_326),
.B(n_275),
.Y(n_390)
);

AND2x4_ASAP7_75t_L g391 ( 
.A(n_351),
.B(n_275),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_321),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_333),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_340),
.Y(n_394)
);

INVx2_ASAP7_75t_L g395 ( 
.A(n_350),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_360),
.Y(n_396)
);

CKINVDCx20_ASAP7_75t_R g397 ( 
.A(n_323),
.Y(n_397)
);

BUFx6f_ASAP7_75t_L g398 ( 
.A(n_363),
.Y(n_398)
);

AND2x2_ASAP7_75t_L g399 ( 
.A(n_326),
.B(n_293),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_327),
.Y(n_400)
);

XOR2xp5_ASAP7_75t_L g401 ( 
.A(n_329),
.B(n_66),
.Y(n_401)
);

AND2x2_ASAP7_75t_L g402 ( 
.A(n_316),
.B(n_335),
.Y(n_402)
);

NOR2xp33_ASAP7_75t_L g403 ( 
.A(n_348),
.B(n_285),
.Y(n_403)
);

AND2x2_ASAP7_75t_L g404 ( 
.A(n_337),
.B(n_296),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_331),
.Y(n_405)
);

BUFx2_ASAP7_75t_L g406 ( 
.A(n_318),
.Y(n_406)
);

AND2x2_ASAP7_75t_L g407 ( 
.A(n_336),
.B(n_296),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_338),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_312),
.Y(n_409)
);

INVx2_ASAP7_75t_L g410 ( 
.A(n_362),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_354),
.Y(n_411)
);

AOI21xp5_ASAP7_75t_L g412 ( 
.A1(n_332),
.A2(n_259),
.B(n_349),
.Y(n_412)
);

NOR2x1_ASAP7_75t_L g413 ( 
.A(n_356),
.B(n_307),
.Y(n_413)
);

XOR2xp5_ASAP7_75t_L g414 ( 
.A(n_361),
.B(n_67),
.Y(n_414)
);

OAI21xp5_ASAP7_75t_L g415 ( 
.A1(n_357),
.A2(n_272),
.B(n_295),
.Y(n_415)
);

XOR2xp5_ASAP7_75t_L g416 ( 
.A(n_358),
.B(n_69),
.Y(n_416)
);

HB1xp67_ASAP7_75t_L g417 ( 
.A(n_318),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_358),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_352),
.Y(n_419)
);

AOI21xp5_ASAP7_75t_L g420 ( 
.A1(n_352),
.A2(n_259),
.B(n_288),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_353),
.Y(n_421)
);

NOR2xp33_ASAP7_75t_L g422 ( 
.A(n_322),
.B(n_285),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_353),
.Y(n_423)
);

NOR2xp33_ASAP7_75t_L g424 ( 
.A(n_322),
.B(n_285),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_328),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_328),
.Y(n_426)
);

AND2x2_ASAP7_75t_L g427 ( 
.A(n_355),
.B(n_284),
.Y(n_427)
);

NOR2xp33_ASAP7_75t_L g428 ( 
.A(n_355),
.B(n_285),
.Y(n_428)
);

XOR2x2_ASAP7_75t_L g429 ( 
.A(n_347),
.B(n_294),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_325),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_347),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_343),
.Y(n_432)
);

NOR2xp33_ASAP7_75t_L g433 ( 
.A(n_345),
.B(n_303),
.Y(n_433)
);

NOR2xp33_ASAP7_75t_L g434 ( 
.A(n_345),
.B(n_303),
.Y(n_434)
);

AND2x2_ASAP7_75t_L g435 ( 
.A(n_384),
.B(n_307),
.Y(n_435)
);

INVx1_ASAP7_75t_SL g436 ( 
.A(n_376),
.Y(n_436)
);

AND2x2_ASAP7_75t_L g437 ( 
.A(n_373),
.B(n_289),
.Y(n_437)
);

OAI21xp5_ASAP7_75t_L g438 ( 
.A1(n_371),
.A2(n_433),
.B(n_434),
.Y(n_438)
);

INVx2_ASAP7_75t_L g439 ( 
.A(n_400),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_371),
.B(n_295),
.Y(n_440)
);

AND2x2_ASAP7_75t_L g441 ( 
.A(n_373),
.B(n_377),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_402),
.B(n_295),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_377),
.B(n_295),
.Y(n_443)
);

AND2x2_ASAP7_75t_L g444 ( 
.A(n_382),
.B(n_289),
.Y(n_444)
);

AND2x2_ASAP7_75t_SL g445 ( 
.A(n_433),
.B(n_289),
.Y(n_445)
);

BUFx6f_ASAP7_75t_L g446 ( 
.A(n_398),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_387),
.Y(n_447)
);

INVxp67_ASAP7_75t_L g448 ( 
.A(n_399),
.Y(n_448)
);

AND2x4_ASAP7_75t_L g449 ( 
.A(n_409),
.B(n_272),
.Y(n_449)
);

NOR2xp67_ASAP7_75t_L g450 ( 
.A(n_410),
.B(n_295),
.Y(n_450)
);

AND2x2_ASAP7_75t_L g451 ( 
.A(n_382),
.B(n_289),
.Y(n_451)
);

INVx1_ASAP7_75t_SL g452 ( 
.A(n_372),
.Y(n_452)
);

INVx2_ASAP7_75t_L g453 ( 
.A(n_405),
.Y(n_453)
);

INVx2_ASAP7_75t_L g454 ( 
.A(n_408),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_L g455 ( 
.A(n_385),
.B(n_303),
.Y(n_455)
);

AND2x2_ASAP7_75t_L g456 ( 
.A(n_383),
.B(n_297),
.Y(n_456)
);

OR2x2_ASAP7_75t_L g457 ( 
.A(n_411),
.B(n_297),
.Y(n_457)
);

AND2x2_ASAP7_75t_L g458 ( 
.A(n_383),
.B(n_413),
.Y(n_458)
);

NOR2xp33_ASAP7_75t_L g459 ( 
.A(n_390),
.B(n_303),
.Y(n_459)
);

BUFx6f_ASAP7_75t_L g460 ( 
.A(n_398),
.Y(n_460)
);

HB1xp67_ASAP7_75t_L g461 ( 
.A(n_390),
.Y(n_461)
);

INVx2_ASAP7_75t_L g462 ( 
.A(n_395),
.Y(n_462)
);

INVx2_ASAP7_75t_L g463 ( 
.A(n_392),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_L g464 ( 
.A(n_385),
.B(n_370),
.Y(n_464)
);

AND2x4_ASAP7_75t_SL g465 ( 
.A(n_391),
.B(n_297),
.Y(n_465)
);

INVx2_ASAP7_75t_L g466 ( 
.A(n_393),
.Y(n_466)
);

INVx2_ASAP7_75t_SL g467 ( 
.A(n_391),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_394),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_370),
.B(n_303),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_396),
.Y(n_470)
);

AND2x2_ASAP7_75t_L g471 ( 
.A(n_427),
.B(n_297),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_388),
.Y(n_472)
);

BUFx3_ASAP7_75t_L g473 ( 
.A(n_407),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_370),
.B(n_292),
.Y(n_474)
);

INVx1_ASAP7_75t_SL g475 ( 
.A(n_404),
.Y(n_475)
);

AND2x2_ASAP7_75t_L g476 ( 
.A(n_403),
.B(n_298),
.Y(n_476)
);

OAI21xp5_ASAP7_75t_L g477 ( 
.A1(n_434),
.A2(n_272),
.B(n_284),
.Y(n_477)
);

INVx2_ASAP7_75t_L g478 ( 
.A(n_398),
.Y(n_478)
);

NOR2xp33_ASAP7_75t_L g479 ( 
.A(n_403),
.B(n_294),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_L g480 ( 
.A(n_370),
.B(n_292),
.Y(n_480)
);

AOI22xp5_ASAP7_75t_L g481 ( 
.A1(n_422),
.A2(n_298),
.B1(n_292),
.B2(n_272),
.Y(n_481)
);

HB1xp67_ASAP7_75t_L g482 ( 
.A(n_422),
.Y(n_482)
);

OAI21xp5_ASAP7_75t_L g483 ( 
.A1(n_389),
.A2(n_272),
.B(n_284),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_L g484 ( 
.A(n_370),
.B(n_292),
.Y(n_484)
);

INVxp67_ASAP7_75t_L g485 ( 
.A(n_366),
.Y(n_485)
);

AND2x2_ASAP7_75t_L g486 ( 
.A(n_424),
.B(n_298),
.Y(n_486)
);

INVx3_ASAP7_75t_L g487 ( 
.A(n_367),
.Y(n_487)
);

NOR2xp33_ASAP7_75t_L g488 ( 
.A(n_378),
.B(n_294),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_L g489 ( 
.A(n_368),
.B(n_292),
.Y(n_489)
);

INVx2_ASAP7_75t_L g490 ( 
.A(n_369),
.Y(n_490)
);

INVx4_ASAP7_75t_L g491 ( 
.A(n_374),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_432),
.Y(n_492)
);

NOR2xp33_ASAP7_75t_L g493 ( 
.A(n_424),
.B(n_276),
.Y(n_493)
);

AND2x2_ASAP7_75t_SL g494 ( 
.A(n_418),
.B(n_298),
.Y(n_494)
);

INVx3_ASAP7_75t_L g495 ( 
.A(n_375),
.Y(n_495)
);

INVx2_ASAP7_75t_L g496 ( 
.A(n_379),
.Y(n_496)
);

INVx2_ASAP7_75t_L g497 ( 
.A(n_381),
.Y(n_497)
);

INVx2_ASAP7_75t_L g498 ( 
.A(n_419),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_L g499 ( 
.A(n_420),
.B(n_276),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_420),
.B(n_276),
.Y(n_500)
);

CKINVDCx5p33_ASAP7_75t_R g501 ( 
.A(n_386),
.Y(n_501)
);

INVx3_ASAP7_75t_SL g502 ( 
.A(n_397),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_421),
.Y(n_503)
);

BUFx6f_ASAP7_75t_L g504 ( 
.A(n_423),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_425),
.Y(n_505)
);

OR2x6_ASAP7_75t_L g506 ( 
.A(n_467),
.B(n_406),
.Y(n_506)
);

INVx2_ASAP7_75t_L g507 ( 
.A(n_495),
.Y(n_507)
);

AND2x2_ASAP7_75t_L g508 ( 
.A(n_435),
.B(n_428),
.Y(n_508)
);

INVx2_ASAP7_75t_L g509 ( 
.A(n_495),
.Y(n_509)
);

INVx3_ASAP7_75t_L g510 ( 
.A(n_478),
.Y(n_510)
);

AND2x2_ASAP7_75t_L g511 ( 
.A(n_435),
.B(n_428),
.Y(n_511)
);

INVx2_ASAP7_75t_L g512 ( 
.A(n_495),
.Y(n_512)
);

OR2x6_ASAP7_75t_L g513 ( 
.A(n_467),
.B(n_412),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_492),
.Y(n_514)
);

AND2x4_ASAP7_75t_L g515 ( 
.A(n_441),
.B(n_412),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_L g516 ( 
.A(n_438),
.B(n_426),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_492),
.Y(n_517)
);

NOR2xp33_ASAP7_75t_L g518 ( 
.A(n_458),
.B(n_380),
.Y(n_518)
);

BUFx3_ASAP7_75t_L g519 ( 
.A(n_504),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_L g520 ( 
.A(n_456),
.B(n_417),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_437),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_437),
.Y(n_522)
);

AND2x2_ASAP7_75t_L g523 ( 
.A(n_475),
.B(n_430),
.Y(n_523)
);

AND2x2_ASAP7_75t_L g524 ( 
.A(n_475),
.B(n_417),
.Y(n_524)
);

BUFx3_ASAP7_75t_L g525 ( 
.A(n_504),
.Y(n_525)
);

AND2x4_ASAP7_75t_L g526 ( 
.A(n_441),
.B(n_415),
.Y(n_526)
);

AND2x2_ASAP7_75t_L g527 ( 
.A(n_458),
.B(n_431),
.Y(n_527)
);

INVx4_ASAP7_75t_L g528 ( 
.A(n_446),
.Y(n_528)
);

INVx2_ASAP7_75t_L g529 ( 
.A(n_462),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_472),
.Y(n_530)
);

HB1xp67_ASAP7_75t_L g531 ( 
.A(n_452),
.Y(n_531)
);

AND2x6_ASAP7_75t_L g532 ( 
.A(n_464),
.B(n_416),
.Y(n_532)
);

AND2x2_ASAP7_75t_L g533 ( 
.A(n_473),
.B(n_429),
.Y(n_533)
);

BUFx12f_ASAP7_75t_L g534 ( 
.A(n_501),
.Y(n_534)
);

NOR2xp33_ASAP7_75t_L g535 ( 
.A(n_482),
.B(n_401),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_472),
.Y(n_536)
);

INVx3_ASAP7_75t_L g537 ( 
.A(n_478),
.Y(n_537)
);

INVx2_ASAP7_75t_L g538 ( 
.A(n_462),
.Y(n_538)
);

OR2x6_ASAP7_75t_L g539 ( 
.A(n_448),
.B(n_414),
.Y(n_539)
);

AND2x2_ASAP7_75t_L g540 ( 
.A(n_473),
.B(n_284),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_439),
.Y(n_541)
);

BUFx6f_ASAP7_75t_L g542 ( 
.A(n_504),
.Y(n_542)
);

BUFx4f_ASAP7_75t_L g543 ( 
.A(n_504),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_L g544 ( 
.A(n_456),
.B(n_284),
.Y(n_544)
);

NAND2x1p5_ASAP7_75t_L g545 ( 
.A(n_504),
.B(n_264),
.Y(n_545)
);

NOR2xp33_ASAP7_75t_L g546 ( 
.A(n_461),
.B(n_70),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_439),
.Y(n_547)
);

CKINVDCx8_ASAP7_75t_R g548 ( 
.A(n_501),
.Y(n_548)
);

NAND2x1p5_ASAP7_75t_L g549 ( 
.A(n_446),
.B(n_264),
.Y(n_549)
);

OR2x2_ASAP7_75t_L g550 ( 
.A(n_436),
.B(n_71),
.Y(n_550)
);

AND2x2_ASAP7_75t_L g551 ( 
.A(n_444),
.B(n_267),
.Y(n_551)
);

BUFx8_ASAP7_75t_L g552 ( 
.A(n_498),
.Y(n_552)
);

CKINVDCx8_ASAP7_75t_R g553 ( 
.A(n_479),
.Y(n_553)
);

AND2x2_ASAP7_75t_SL g554 ( 
.A(n_445),
.B(n_272),
.Y(n_554)
);

BUFx6f_ASAP7_75t_L g555 ( 
.A(n_446),
.Y(n_555)
);

BUFx6f_ASAP7_75t_L g556 ( 
.A(n_446),
.Y(n_556)
);

NAND2x1p5_ASAP7_75t_L g557 ( 
.A(n_446),
.B(n_460),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_L g558 ( 
.A(n_445),
.B(n_476),
.Y(n_558)
);

NOR2xp33_ASAP7_75t_L g559 ( 
.A(n_457),
.B(n_74),
.Y(n_559)
);

AND2x2_ASAP7_75t_L g560 ( 
.A(n_444),
.B(n_451),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_L g561 ( 
.A(n_445),
.B(n_264),
.Y(n_561)
);

INVx4_ASAP7_75t_L g562 ( 
.A(n_460),
.Y(n_562)
);

OR2x2_ASAP7_75t_L g563 ( 
.A(n_457),
.B(n_75),
.Y(n_563)
);

BUFx6f_ASAP7_75t_L g564 ( 
.A(n_460),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_453),
.Y(n_565)
);

NOR2x1_ASAP7_75t_R g566 ( 
.A(n_534),
.B(n_498),
.Y(n_566)
);

NAND2x1p5_ASAP7_75t_L g567 ( 
.A(n_543),
.B(n_460),
.Y(n_567)
);

INVx2_ASAP7_75t_SL g568 ( 
.A(n_531),
.Y(n_568)
);

INVx2_ASAP7_75t_L g569 ( 
.A(n_529),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_SL g570 ( 
.A(n_518),
.B(n_465),
.Y(n_570)
);

BUFx3_ASAP7_75t_L g571 ( 
.A(n_531),
.Y(n_571)
);

INVx3_ASAP7_75t_L g572 ( 
.A(n_528),
.Y(n_572)
);

BUFx6f_ASAP7_75t_L g573 ( 
.A(n_555),
.Y(n_573)
);

INVx3_ASAP7_75t_L g574 ( 
.A(n_528),
.Y(n_574)
);

NAND2x1p5_ASAP7_75t_L g575 ( 
.A(n_543),
.B(n_460),
.Y(n_575)
);

NAND2x1p5_ASAP7_75t_L g576 ( 
.A(n_519),
.B(n_491),
.Y(n_576)
);

INVx1_ASAP7_75t_SL g577 ( 
.A(n_523),
.Y(n_577)
);

INVxp67_ASAP7_75t_SL g578 ( 
.A(n_542),
.Y(n_578)
);

BUFx8_ASAP7_75t_L g579 ( 
.A(n_534),
.Y(n_579)
);

BUFx3_ASAP7_75t_L g580 ( 
.A(n_548),
.Y(n_580)
);

BUFx4f_ASAP7_75t_L g581 ( 
.A(n_506),
.Y(n_581)
);

BUFx3_ASAP7_75t_L g582 ( 
.A(n_548),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_514),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_517),
.Y(n_584)
);

INVx3_ASAP7_75t_L g585 ( 
.A(n_528),
.Y(n_585)
);

INVxp67_ASAP7_75t_SL g586 ( 
.A(n_542),
.Y(n_586)
);

BUFx6f_ASAP7_75t_L g587 ( 
.A(n_555),
.Y(n_587)
);

INVx5_ASAP7_75t_L g588 ( 
.A(n_542),
.Y(n_588)
);

OR2x2_ASAP7_75t_L g589 ( 
.A(n_518),
.B(n_485),
.Y(n_589)
);

INVx2_ASAP7_75t_L g590 ( 
.A(n_529),
.Y(n_590)
);

BUFx4_ASAP7_75t_SL g591 ( 
.A(n_506),
.Y(n_591)
);

BUFx4f_ASAP7_75t_SL g592 ( 
.A(n_552),
.Y(n_592)
);

INVx6_ASAP7_75t_SL g593 ( 
.A(n_539),
.Y(n_593)
);

INVx5_ASAP7_75t_L g594 ( 
.A(n_542),
.Y(n_594)
);

NOR2xp33_ASAP7_75t_L g595 ( 
.A(n_553),
.B(n_502),
.Y(n_595)
);

NAND2x1p5_ASAP7_75t_L g596 ( 
.A(n_519),
.B(n_491),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_L g597 ( 
.A(n_560),
.B(n_476),
.Y(n_597)
);

CKINVDCx20_ASAP7_75t_R g598 ( 
.A(n_553),
.Y(n_598)
);

BUFx3_ASAP7_75t_L g599 ( 
.A(n_552),
.Y(n_599)
);

INVx2_ASAP7_75t_SL g600 ( 
.A(n_550),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_530),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_536),
.Y(n_602)
);

INVx1_ASAP7_75t_SL g603 ( 
.A(n_524),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_L g604 ( 
.A(n_516),
.B(n_486),
.Y(n_604)
);

NOR2xp33_ASAP7_75t_L g605 ( 
.A(n_527),
.B(n_494),
.Y(n_605)
);

CKINVDCx16_ASAP7_75t_R g606 ( 
.A(n_539),
.Y(n_606)
);

BUFx2_ASAP7_75t_SL g607 ( 
.A(n_515),
.Y(n_607)
);

BUFx6f_ASAP7_75t_L g608 ( 
.A(n_555),
.Y(n_608)
);

BUFx4_ASAP7_75t_SL g609 ( 
.A(n_506),
.Y(n_609)
);

INVx2_ASAP7_75t_L g610 ( 
.A(n_538),
.Y(n_610)
);

INVx3_ASAP7_75t_SL g611 ( 
.A(n_539),
.Y(n_611)
);

OAI22xp33_ASAP7_75t_L g612 ( 
.A1(n_520),
.A2(n_481),
.B1(n_503),
.B2(n_505),
.Y(n_612)
);

INVx6_ASAP7_75t_L g613 ( 
.A(n_552),
.Y(n_613)
);

INVx3_ASAP7_75t_L g614 ( 
.A(n_555),
.Y(n_614)
);

BUFx12f_ASAP7_75t_L g615 ( 
.A(n_515),
.Y(n_615)
);

NAND2x1p5_ASAP7_75t_L g616 ( 
.A(n_525),
.B(n_491),
.Y(n_616)
);

INVx2_ASAP7_75t_L g617 ( 
.A(n_569),
.Y(n_617)
);

INVx2_ASAP7_75t_L g618 ( 
.A(n_590),
.Y(n_618)
);

INVx3_ASAP7_75t_L g619 ( 
.A(n_572),
.Y(n_619)
);

AOI22xp5_ASAP7_75t_L g620 ( 
.A1(n_605),
.A2(n_535),
.B1(n_532),
.B2(n_515),
.Y(n_620)
);

OAI22xp5_ASAP7_75t_L g621 ( 
.A1(n_605),
.A2(n_558),
.B1(n_525),
.B2(n_554),
.Y(n_621)
);

CKINVDCx11_ASAP7_75t_R g622 ( 
.A(n_611),
.Y(n_622)
);

BUFx2_ASAP7_75t_L g623 ( 
.A(n_571),
.Y(n_623)
);

NAND2x1p5_ASAP7_75t_L g624 ( 
.A(n_588),
.B(n_562),
.Y(n_624)
);

INVx8_ASAP7_75t_L g625 ( 
.A(n_588),
.Y(n_625)
);

BUFx6f_ASAP7_75t_L g626 ( 
.A(n_573),
.Y(n_626)
);

OAI22xp5_ASAP7_75t_L g627 ( 
.A1(n_607),
.A2(n_554),
.B1(n_465),
.B2(n_526),
.Y(n_627)
);

AOI22xp33_ASAP7_75t_L g628 ( 
.A1(n_589),
.A2(n_532),
.B1(n_511),
.B2(n_508),
.Y(n_628)
);

BUFx6f_ASAP7_75t_L g629 ( 
.A(n_573),
.Y(n_629)
);

BUFx12f_ASAP7_75t_L g630 ( 
.A(n_579),
.Y(n_630)
);

INVx6_ASAP7_75t_L g631 ( 
.A(n_579),
.Y(n_631)
);

BUFx12f_ASAP7_75t_L g632 ( 
.A(n_613),
.Y(n_632)
);

NAND2x1p5_ASAP7_75t_L g633 ( 
.A(n_588),
.B(n_562),
.Y(n_633)
);

OAI22xp33_ASAP7_75t_L g634 ( 
.A1(n_577),
.A2(n_502),
.B1(n_535),
.B2(n_563),
.Y(n_634)
);

CKINVDCx20_ASAP7_75t_R g635 ( 
.A(n_598),
.Y(n_635)
);

INVx6_ASAP7_75t_L g636 ( 
.A(n_613),
.Y(n_636)
);

AOI22xp33_ASAP7_75t_L g637 ( 
.A1(n_615),
.A2(n_532),
.B1(n_526),
.B2(n_533),
.Y(n_637)
);

INVx4_ASAP7_75t_L g638 ( 
.A(n_588),
.Y(n_638)
);

INVx2_ASAP7_75t_L g639 ( 
.A(n_610),
.Y(n_639)
);

INVx2_ASAP7_75t_SL g640 ( 
.A(n_568),
.Y(n_640)
);

AOI22xp33_ASAP7_75t_L g641 ( 
.A1(n_570),
.A2(n_532),
.B1(n_526),
.B2(n_513),
.Y(n_641)
);

AOI22xp5_ASAP7_75t_L g642 ( 
.A1(n_577),
.A2(n_532),
.B1(n_486),
.B2(n_521),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_583),
.Y(n_643)
);

CKINVDCx11_ASAP7_75t_R g644 ( 
.A(n_611),
.Y(n_644)
);

OAI22xp5_ASAP7_75t_L g645 ( 
.A1(n_603),
.A2(n_546),
.B1(n_559),
.B2(n_513),
.Y(n_645)
);

INVx1_ASAP7_75t_SL g646 ( 
.A(n_603),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_584),
.Y(n_647)
);

INVx6_ASAP7_75t_L g648 ( 
.A(n_613),
.Y(n_648)
);

BUFx6f_ASAP7_75t_L g649 ( 
.A(n_573),
.Y(n_649)
);

BUFx2_ASAP7_75t_SL g650 ( 
.A(n_580),
.Y(n_650)
);

CKINVDCx11_ASAP7_75t_R g651 ( 
.A(n_606),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_601),
.Y(n_652)
);

INVx6_ASAP7_75t_L g653 ( 
.A(n_582),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_602),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_604),
.Y(n_655)
);

CKINVDCx11_ASAP7_75t_R g656 ( 
.A(n_599),
.Y(n_656)
);

BUFx3_ASAP7_75t_L g657 ( 
.A(n_592),
.Y(n_657)
);

OAI22xp5_ASAP7_75t_L g658 ( 
.A1(n_604),
.A2(n_546),
.B1(n_559),
.B2(n_513),
.Y(n_658)
);

OAI21xp33_ASAP7_75t_L g659 ( 
.A1(n_600),
.A2(n_488),
.B(n_493),
.Y(n_659)
);

OAI22xp5_ASAP7_75t_L g660 ( 
.A1(n_620),
.A2(n_595),
.B1(n_581),
.B2(n_592),
.Y(n_660)
);

OAI22xp5_ASAP7_75t_L g661 ( 
.A1(n_628),
.A2(n_581),
.B1(n_596),
.B2(n_616),
.Y(n_661)
);

AOI22xp33_ASAP7_75t_SL g662 ( 
.A1(n_645),
.A2(n_477),
.B1(n_597),
.B2(n_494),
.Y(n_662)
);

AND2x2_ASAP7_75t_L g663 ( 
.A(n_655),
.B(n_541),
.Y(n_663)
);

AOI22xp33_ASAP7_75t_L g664 ( 
.A1(n_634),
.A2(n_593),
.B1(n_597),
.B2(n_522),
.Y(n_664)
);

OAI21xp5_ASAP7_75t_SL g665 ( 
.A1(n_637),
.A2(n_481),
.B(n_499),
.Y(n_665)
);

AOI22xp33_ASAP7_75t_L g666 ( 
.A1(n_659),
.A2(n_593),
.B1(n_454),
.B2(n_453),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_L g667 ( 
.A(n_655),
.B(n_451),
.Y(n_667)
);

INVx5_ASAP7_75t_SL g668 ( 
.A(n_626),
.Y(n_668)
);

AOI211xp5_ASAP7_75t_L g669 ( 
.A1(n_658),
.A2(n_502),
.B(n_566),
.C(n_612),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_643),
.Y(n_670)
);

AOI22xp33_ASAP7_75t_L g671 ( 
.A1(n_641),
.A2(n_454),
.B1(n_547),
.B2(n_565),
.Y(n_671)
);

AOI22xp33_ASAP7_75t_L g672 ( 
.A1(n_642),
.A2(n_442),
.B1(n_463),
.B2(n_466),
.Y(n_672)
);

INVx4_ASAP7_75t_L g673 ( 
.A(n_625),
.Y(n_673)
);

AOI22xp33_ASAP7_75t_L g674 ( 
.A1(n_642),
.A2(n_466),
.B1(n_463),
.B2(n_490),
.Y(n_674)
);

AOI22xp5_ASAP7_75t_L g675 ( 
.A1(n_635),
.A2(n_540),
.B1(n_500),
.B2(n_471),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_L g676 ( 
.A(n_646),
.B(n_471),
.Y(n_676)
);

BUFx2_ASAP7_75t_L g677 ( 
.A(n_623),
.Y(n_677)
);

AND2x2_ASAP7_75t_L g678 ( 
.A(n_643),
.B(n_538),
.Y(n_678)
);

AOI22xp33_ASAP7_75t_L g679 ( 
.A1(n_622),
.A2(n_490),
.B1(n_496),
.B2(n_497),
.Y(n_679)
);

INVx2_ASAP7_75t_L g680 ( 
.A(n_647),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_647),
.Y(n_681)
);

INVx3_ASAP7_75t_L g682 ( 
.A(n_638),
.Y(n_682)
);

INVx2_ASAP7_75t_SL g683 ( 
.A(n_625),
.Y(n_683)
);

OAI21xp5_ASAP7_75t_SL g684 ( 
.A1(n_627),
.A2(n_621),
.B(n_612),
.Y(n_684)
);

AOI22xp33_ASAP7_75t_SL g685 ( 
.A1(n_650),
.A2(n_494),
.B1(n_616),
.B2(n_576),
.Y(n_685)
);

AND2x2_ASAP7_75t_L g686 ( 
.A(n_652),
.B(n_578),
.Y(n_686)
);

AND2x2_ASAP7_75t_L g687 ( 
.A(n_652),
.B(n_578),
.Y(n_687)
);

AND2x2_ASAP7_75t_L g688 ( 
.A(n_654),
.B(n_586),
.Y(n_688)
);

HB1xp67_ASAP7_75t_L g689 ( 
.A(n_640),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_654),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_617),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_618),
.Y(n_692)
);

AOI22xp33_ASAP7_75t_L g693 ( 
.A1(n_644),
.A2(n_496),
.B1(n_497),
.B2(n_470),
.Y(n_693)
);

AOI22xp33_ASAP7_75t_L g694 ( 
.A1(n_651),
.A2(n_470),
.B1(n_468),
.B2(n_447),
.Y(n_694)
);

BUFx3_ASAP7_75t_L g695 ( 
.A(n_653),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_639),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_626),
.Y(n_697)
);

HB1xp67_ASAP7_75t_L g698 ( 
.A(n_653),
.Y(n_698)
);

AND2x2_ASAP7_75t_L g699 ( 
.A(n_619),
.B(n_586),
.Y(n_699)
);

INVx1_ASAP7_75t_SL g700 ( 
.A(n_656),
.Y(n_700)
);

OAI222xp33_ASAP7_75t_L g701 ( 
.A1(n_619),
.A2(n_596),
.B1(n_576),
.B2(n_561),
.C1(n_440),
.C2(n_468),
.Y(n_701)
);

OAI22xp5_ASAP7_75t_L g702 ( 
.A1(n_636),
.A2(n_567),
.B1(n_575),
.B2(n_594),
.Y(n_702)
);

OAI222xp33_ASAP7_75t_L g703 ( 
.A1(n_638),
.A2(n_567),
.B1(n_575),
.B2(n_509),
.C1(n_512),
.C2(n_507),
.Y(n_703)
);

AOI22xp33_ASAP7_75t_L g704 ( 
.A1(n_632),
.A2(n_447),
.B1(n_487),
.B2(n_551),
.Y(n_704)
);

INVx4_ASAP7_75t_SL g705 ( 
.A(n_636),
.Y(n_705)
);

INVx4_ASAP7_75t_L g706 ( 
.A(n_626),
.Y(n_706)
);

BUFx3_ASAP7_75t_L g707 ( 
.A(n_648),
.Y(n_707)
);

AOI22xp33_ASAP7_75t_SL g708 ( 
.A1(n_631),
.A2(n_609),
.B1(n_591),
.B2(n_483),
.Y(n_708)
);

BUFx2_ASAP7_75t_L g709 ( 
.A(n_629),
.Y(n_709)
);

AOI22xp33_ASAP7_75t_L g710 ( 
.A1(n_648),
.A2(n_487),
.B1(n_450),
.B2(n_449),
.Y(n_710)
);

AOI22xp33_ASAP7_75t_L g711 ( 
.A1(n_657),
.A2(n_487),
.B1(n_450),
.B2(n_449),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_629),
.Y(n_712)
);

AOI22xp33_ASAP7_75t_L g713 ( 
.A1(n_662),
.A2(n_664),
.B1(n_660),
.B2(n_675),
.Y(n_713)
);

AOI22xp33_ASAP7_75t_L g714 ( 
.A1(n_666),
.A2(n_631),
.B1(n_630),
.B2(n_512),
.Y(n_714)
);

AOI22xp33_ASAP7_75t_SL g715 ( 
.A1(n_661),
.A2(n_455),
.B1(n_572),
.B2(n_574),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_681),
.Y(n_716)
);

AOI22xp33_ASAP7_75t_SL g717 ( 
.A1(n_677),
.A2(n_574),
.B1(n_585),
.B2(n_594),
.Y(n_717)
);

AOI22xp33_ASAP7_75t_L g718 ( 
.A1(n_677),
.A2(n_480),
.B1(n_484),
.B2(n_474),
.Y(n_718)
);

AOI22xp33_ASAP7_75t_L g719 ( 
.A1(n_694),
.A2(n_708),
.B1(n_693),
.B2(n_679),
.Y(n_719)
);

AOI22xp33_ASAP7_75t_L g720 ( 
.A1(n_685),
.A2(n_544),
.B1(n_459),
.B2(n_449),
.Y(n_720)
);

AND2x2_ASAP7_75t_SL g721 ( 
.A(n_669),
.B(n_587),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_681),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_L g723 ( 
.A(n_691),
.B(n_692),
.Y(n_723)
);

AOI22xp33_ASAP7_75t_SL g724 ( 
.A1(n_702),
.A2(n_585),
.B1(n_594),
.B2(n_609),
.Y(n_724)
);

AOI22xp33_ASAP7_75t_L g725 ( 
.A1(n_671),
.A2(n_449),
.B1(n_507),
.B2(n_509),
.Y(n_725)
);

OA21x2_ASAP7_75t_L g726 ( 
.A1(n_684),
.A2(n_701),
.B(n_665),
.Y(n_726)
);

AOI22xp33_ASAP7_75t_L g727 ( 
.A1(n_689),
.A2(n_537),
.B1(n_510),
.B2(n_443),
.Y(n_727)
);

AOI22xp33_ASAP7_75t_L g728 ( 
.A1(n_672),
.A2(n_510),
.B1(n_537),
.B2(n_629),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_670),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_L g730 ( 
.A(n_696),
.B(n_649),
.Y(n_730)
);

NAND2xp33_ASAP7_75t_SL g731 ( 
.A(n_698),
.B(n_591),
.Y(n_731)
);

INVx2_ASAP7_75t_L g732 ( 
.A(n_680),
.Y(n_732)
);

OAI22xp5_ASAP7_75t_L g733 ( 
.A1(n_704),
.A2(n_633),
.B1(n_624),
.B2(n_594),
.Y(n_733)
);

OAI22xp5_ASAP7_75t_L g734 ( 
.A1(n_711),
.A2(n_503),
.B1(n_505),
.B2(n_545),
.Y(n_734)
);

OAI22xp5_ASAP7_75t_L g735 ( 
.A1(n_676),
.A2(n_545),
.B1(n_614),
.B2(n_649),
.Y(n_735)
);

OAI22xp5_ASAP7_75t_L g736 ( 
.A1(n_674),
.A2(n_614),
.B1(n_649),
.B2(n_557),
.Y(n_736)
);

AOI22xp33_ASAP7_75t_L g737 ( 
.A1(n_663),
.A2(n_469),
.B1(n_608),
.B2(n_587),
.Y(n_737)
);

OAI221xp5_ASAP7_75t_L g738 ( 
.A1(n_710),
.A2(n_489),
.B1(n_557),
.B2(n_564),
.C(n_556),
.Y(n_738)
);

AOI221xp5_ASAP7_75t_L g739 ( 
.A1(n_667),
.A2(n_264),
.B1(n_587),
.B2(n_608),
.C(n_556),
.Y(n_739)
);

NAND3xp33_ASAP7_75t_L g740 ( 
.A(n_663),
.B(n_608),
.C(n_564),
.Y(n_740)
);

OAI222xp33_ASAP7_75t_L g741 ( 
.A1(n_690),
.A2(n_549),
.B1(n_77),
.B2(n_79),
.C1(n_80),
.C2(n_81),
.Y(n_741)
);

OAI22xp5_ASAP7_75t_L g742 ( 
.A1(n_695),
.A2(n_564),
.B1(n_556),
.B2(n_549),
.Y(n_742)
);

OAI22xp5_ASAP7_75t_L g743 ( 
.A1(n_695),
.A2(n_564),
.B1(n_556),
.B2(n_264),
.Y(n_743)
);

AOI22xp33_ASAP7_75t_L g744 ( 
.A1(n_680),
.A2(n_76),
.B1(n_86),
.B2(n_87),
.Y(n_744)
);

AOI22xp33_ASAP7_75t_L g745 ( 
.A1(n_707),
.A2(n_88),
.B1(n_89),
.B2(n_91),
.Y(n_745)
);

AND2x2_ASAP7_75t_L g746 ( 
.A(n_686),
.B(n_687),
.Y(n_746)
);

AOI22xp33_ASAP7_75t_L g747 ( 
.A1(n_707),
.A2(n_93),
.B1(n_94),
.B2(n_95),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_L g748 ( 
.A(n_686),
.B(n_97),
.Y(n_748)
);

OAI221xp5_ASAP7_75t_L g749 ( 
.A1(n_700),
.A2(n_98),
.B1(n_99),
.B2(n_101),
.C(n_102),
.Y(n_749)
);

NAND3xp33_ASAP7_75t_L g750 ( 
.A(n_687),
.B(n_103),
.C(n_105),
.Y(n_750)
);

AOI22xp33_ASAP7_75t_L g751 ( 
.A1(n_678),
.A2(n_179),
.B1(n_108),
.B2(n_110),
.Y(n_751)
);

AOI22xp33_ASAP7_75t_L g752 ( 
.A1(n_678),
.A2(n_106),
.B1(n_111),
.B2(n_115),
.Y(n_752)
);

NAND3xp33_ASAP7_75t_L g753 ( 
.A(n_688),
.B(n_116),
.C(n_118),
.Y(n_753)
);

AOI22xp33_ASAP7_75t_L g754 ( 
.A1(n_688),
.A2(n_178),
.B1(n_121),
.B2(n_122),
.Y(n_754)
);

INVx2_ASAP7_75t_L g755 ( 
.A(n_699),
.Y(n_755)
);

OAI221xp5_ASAP7_75t_SL g756 ( 
.A1(n_713),
.A2(n_719),
.B1(n_754),
.B2(n_749),
.C(n_752),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_L g757 ( 
.A(n_746),
.B(n_699),
.Y(n_757)
);

NAND3xp33_ASAP7_75t_L g758 ( 
.A(n_713),
.B(n_712),
.C(n_697),
.Y(n_758)
);

NAND3xp33_ASAP7_75t_L g759 ( 
.A(n_754),
.B(n_712),
.C(n_706),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_SL g760 ( 
.A(n_721),
.B(n_682),
.Y(n_760)
);

NOR3xp33_ASAP7_75t_L g761 ( 
.A(n_750),
.B(n_673),
.C(n_682),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_L g762 ( 
.A(n_755),
.B(n_709),
.Y(n_762)
);

OAI21xp33_ASAP7_75t_L g763 ( 
.A1(n_751),
.A2(n_683),
.B(n_682),
.Y(n_763)
);

AND2x2_ASAP7_75t_L g764 ( 
.A(n_716),
.B(n_709),
.Y(n_764)
);

NAND3xp33_ASAP7_75t_L g765 ( 
.A(n_751),
.B(n_706),
.C(n_673),
.Y(n_765)
);

NAND3xp33_ASAP7_75t_L g766 ( 
.A(n_752),
.B(n_706),
.C(n_673),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_L g767 ( 
.A(n_723),
.B(n_705),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_L g768 ( 
.A(n_729),
.B(n_705),
.Y(n_768)
);

AND2x2_ASAP7_75t_L g769 ( 
.A(n_722),
.B(n_668),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_732),
.Y(n_770)
);

AOI221xp5_ASAP7_75t_L g771 ( 
.A1(n_741),
.A2(n_683),
.B1(n_703),
.B2(n_705),
.C(n_129),
.Y(n_771)
);

AND2x2_ASAP7_75t_L g772 ( 
.A(n_726),
.B(n_668),
.Y(n_772)
);

AND2x2_ASAP7_75t_L g773 ( 
.A(n_726),
.B(n_668),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_L g774 ( 
.A(n_726),
.B(n_730),
.Y(n_774)
);

OAI21xp33_ASAP7_75t_L g775 ( 
.A1(n_714),
.A2(n_705),
.B(n_123),
.Y(n_775)
);

AOI211xp5_ASAP7_75t_SL g776 ( 
.A1(n_733),
.A2(n_668),
.B(n_126),
.C(n_132),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_L g777 ( 
.A(n_748),
.B(n_120),
.Y(n_777)
);

AND2x2_ASAP7_75t_L g778 ( 
.A(n_721),
.B(n_133),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_L g779 ( 
.A(n_715),
.B(n_135),
.Y(n_779)
);

NAND3xp33_ASAP7_75t_L g780 ( 
.A(n_753),
.B(n_136),
.C(n_137),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_L g781 ( 
.A(n_714),
.B(n_140),
.Y(n_781)
);

AND2x2_ASAP7_75t_L g782 ( 
.A(n_737),
.B(n_141),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_L g783 ( 
.A(n_724),
.B(n_142),
.Y(n_783)
);

AND2x2_ASAP7_75t_L g784 ( 
.A(n_720),
.B(n_143),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_L g785 ( 
.A(n_735),
.B(n_144),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_L g786 ( 
.A(n_718),
.B(n_145),
.Y(n_786)
);

HB1xp67_ASAP7_75t_L g787 ( 
.A(n_764),
.Y(n_787)
);

INVx2_ASAP7_75t_SL g788 ( 
.A(n_764),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_L g789 ( 
.A(n_774),
.B(n_757),
.Y(n_789)
);

AO21x2_ASAP7_75t_L g790 ( 
.A1(n_761),
.A2(n_740),
.B(n_738),
.Y(n_790)
);

AND2x2_ASAP7_75t_L g791 ( 
.A(n_773),
.B(n_717),
.Y(n_791)
);

AND2x2_ASAP7_75t_L g792 ( 
.A(n_773),
.B(n_739),
.Y(n_792)
);

OA211x2_ASAP7_75t_L g793 ( 
.A1(n_771),
.A2(n_763),
.B(n_775),
.C(n_760),
.Y(n_793)
);

AND2x4_ASAP7_75t_L g794 ( 
.A(n_769),
.B(n_747),
.Y(n_794)
);

OR2x2_ASAP7_75t_L g795 ( 
.A(n_762),
.B(n_731),
.Y(n_795)
);

OR2x2_ASAP7_75t_L g796 ( 
.A(n_770),
.B(n_742),
.Y(n_796)
);

NAND3xp33_ASAP7_75t_L g797 ( 
.A(n_756),
.B(n_744),
.C(n_745),
.Y(n_797)
);

AND2x4_ASAP7_75t_L g798 ( 
.A(n_769),
.B(n_727),
.Y(n_798)
);

NOR2x1_ASAP7_75t_SL g799 ( 
.A(n_760),
.B(n_743),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_L g800 ( 
.A(n_767),
.B(n_734),
.Y(n_800)
);

AND2x2_ASAP7_75t_L g801 ( 
.A(n_772),
.B(n_736),
.Y(n_801)
);

INVx3_ASAP7_75t_L g802 ( 
.A(n_768),
.Y(n_802)
);

NAND3xp33_ASAP7_75t_L g803 ( 
.A(n_758),
.B(n_725),
.C(n_728),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_L g804 ( 
.A(n_759),
.B(n_778),
.Y(n_804)
);

NAND4xp75_ASAP7_75t_L g805 ( 
.A(n_778),
.B(n_147),
.C(n_149),
.D(n_153),
.Y(n_805)
);

AND2x2_ASAP7_75t_L g806 ( 
.A(n_787),
.B(n_776),
.Y(n_806)
);

XNOR2xp5_ASAP7_75t_L g807 ( 
.A(n_793),
.B(n_765),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_788),
.Y(n_808)
);

AND2x2_ASAP7_75t_L g809 ( 
.A(n_788),
.B(n_766),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_789),
.Y(n_810)
);

BUFx2_ASAP7_75t_L g811 ( 
.A(n_802),
.Y(n_811)
);

INVx2_ASAP7_75t_L g812 ( 
.A(n_802),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_802),
.Y(n_813)
);

NAND4xp75_ASAP7_75t_L g814 ( 
.A(n_792),
.B(n_784),
.C(n_779),
.D(n_782),
.Y(n_814)
);

NAND4xp75_ASAP7_75t_L g815 ( 
.A(n_792),
.B(n_784),
.C(n_782),
.D(n_783),
.Y(n_815)
);

INVxp67_ASAP7_75t_L g816 ( 
.A(n_804),
.Y(n_816)
);

INVx2_ASAP7_75t_L g817 ( 
.A(n_796),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_817),
.Y(n_818)
);

XOR2x2_ASAP7_75t_L g819 ( 
.A(n_807),
.B(n_797),
.Y(n_819)
);

XOR2x2_ASAP7_75t_L g820 ( 
.A(n_807),
.B(n_795),
.Y(n_820)
);

INVx2_ASAP7_75t_L g821 ( 
.A(n_817),
.Y(n_821)
);

INVx1_ASAP7_75t_SL g822 ( 
.A(n_809),
.Y(n_822)
);

INVx2_ASAP7_75t_L g823 ( 
.A(n_821),
.Y(n_823)
);

BUFx3_ASAP7_75t_L g824 ( 
.A(n_820),
.Y(n_824)
);

INVx2_ASAP7_75t_L g825 ( 
.A(n_821),
.Y(n_825)
);

AOI22x1_ASAP7_75t_L g826 ( 
.A1(n_819),
.A2(n_806),
.B1(n_795),
.B2(n_809),
.Y(n_826)
);

AOI22xp5_ASAP7_75t_SL g827 ( 
.A1(n_822),
.A2(n_806),
.B1(n_816),
.B2(n_811),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_823),
.Y(n_828)
);

INVx2_ASAP7_75t_SL g829 ( 
.A(n_827),
.Y(n_829)
);

INVx2_ASAP7_75t_L g830 ( 
.A(n_825),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_830),
.Y(n_831)
);

AND4x1_ASAP7_75t_L g832 ( 
.A(n_828),
.B(n_824),
.C(n_826),
.D(n_780),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_831),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_832),
.Y(n_834)
);

INVxp67_ASAP7_75t_L g835 ( 
.A(n_832),
.Y(n_835)
);

AOI22xp33_ASAP7_75t_L g836 ( 
.A1(n_834),
.A2(n_829),
.B1(n_826),
.B2(n_830),
.Y(n_836)
);

INVxp67_ASAP7_75t_SL g837 ( 
.A(n_835),
.Y(n_837)
);

NOR4xp25_ASAP7_75t_L g838 ( 
.A(n_833),
.B(n_829),
.C(n_822),
.D(n_818),
.Y(n_838)
);

AOI22xp5_ASAP7_75t_L g839 ( 
.A1(n_835),
.A2(n_814),
.B1(n_815),
.B2(n_805),
.Y(n_839)
);

AOI22xp33_ASAP7_75t_L g840 ( 
.A1(n_834),
.A2(n_790),
.B1(n_794),
.B2(n_798),
.Y(n_840)
);

INVxp67_ASAP7_75t_SL g841 ( 
.A(n_835),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_837),
.Y(n_842)
);

AOI22xp5_ASAP7_75t_L g843 ( 
.A1(n_836),
.A2(n_810),
.B1(n_790),
.B2(n_791),
.Y(n_843)
);

INVx2_ASAP7_75t_L g844 ( 
.A(n_841),
.Y(n_844)
);

NOR2x1_ASAP7_75t_L g845 ( 
.A(n_838),
.B(n_811),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_839),
.Y(n_846)
);

AOI22xp5_ASAP7_75t_L g847 ( 
.A1(n_840),
.A2(n_790),
.B1(n_791),
.B2(n_800),
.Y(n_847)
);

AOI22xp5_ASAP7_75t_L g848 ( 
.A1(n_836),
.A2(n_794),
.B1(n_803),
.B2(n_813),
.Y(n_848)
);

INVx2_ASAP7_75t_SL g849 ( 
.A(n_844),
.Y(n_849)
);

OAI22xp5_ASAP7_75t_L g850 ( 
.A1(n_848),
.A2(n_808),
.B1(n_812),
.B2(n_794),
.Y(n_850)
);

OAI211xp5_ASAP7_75t_L g851 ( 
.A1(n_845),
.A2(n_781),
.B(n_786),
.C(n_785),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_842),
.Y(n_852)
);

AO22x2_ASAP7_75t_L g853 ( 
.A1(n_846),
.A2(n_843),
.B1(n_847),
.B2(n_812),
.Y(n_853)
);

NAND4xp75_ASAP7_75t_L g854 ( 
.A(n_845),
.B(n_777),
.C(n_801),
.D(n_799),
.Y(n_854)
);

INVx2_ASAP7_75t_L g855 ( 
.A(n_849),
.Y(n_855)
);

INVx2_ASAP7_75t_L g856 ( 
.A(n_852),
.Y(n_856)
);

HB1xp67_ASAP7_75t_L g857 ( 
.A(n_854),
.Y(n_857)
);

OA22x2_ASAP7_75t_L g858 ( 
.A1(n_850),
.A2(n_798),
.B1(n_801),
.B2(n_796),
.Y(n_858)
);

INVx3_ASAP7_75t_L g859 ( 
.A(n_853),
.Y(n_859)
);

INVx1_ASAP7_75t_L g860 ( 
.A(n_851),
.Y(n_860)
);

INVx1_ASAP7_75t_L g861 ( 
.A(n_855),
.Y(n_861)
);

INVxp67_ASAP7_75t_SL g862 ( 
.A(n_859),
.Y(n_862)
);

CKINVDCx20_ASAP7_75t_R g863 ( 
.A(n_857),
.Y(n_863)
);

AOI22xp5_ASAP7_75t_L g864 ( 
.A1(n_860),
.A2(n_798),
.B1(n_155),
.B2(n_157),
.Y(n_864)
);

AOI22xp5_ASAP7_75t_L g865 ( 
.A1(n_860),
.A2(n_154),
.B1(n_159),
.B2(n_160),
.Y(n_865)
);

INVx2_ASAP7_75t_L g866 ( 
.A(n_863),
.Y(n_866)
);

OR2x2_ASAP7_75t_SL g867 ( 
.A(n_861),
.B(n_856),
.Y(n_867)
);

AOI22xp33_ASAP7_75t_L g868 ( 
.A1(n_866),
.A2(n_862),
.B1(n_858),
.B2(n_864),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_868),
.Y(n_869)
);

OAI22xp33_ASAP7_75t_L g870 ( 
.A1(n_869),
.A2(n_865),
.B1(n_867),
.B2(n_164),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_870),
.Y(n_871)
);

AOI221xp5_ASAP7_75t_L g872 ( 
.A1(n_871),
.A2(n_161),
.B1(n_163),
.B2(n_167),
.C(n_168),
.Y(n_872)
);

AOI211xp5_ASAP7_75t_L g873 ( 
.A1(n_872),
.A2(n_169),
.B(n_170),
.C(n_171),
.Y(n_873)
);


endmodule