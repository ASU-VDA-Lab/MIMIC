module real_aes_2909_n_398 (n_76, n_113, n_187, n_90, n_257, n_390, n_65, n_74, n_185, n_285, n_30, n_222, n_61, n_20, n_287, n_357, n_386, n_64, n_254, n_207, n_10, n_83, n_181, n_362, n_124, n_191, n_209, n_299, n_322, n_328, n_19, n_40, n_318, n_355, n_239, n_100, n_54, n_112, n_319, n_364, n_35, n_42, n_329, n_132, n_131, n_144, n_169, n_242, n_376, n_308, n_172, n_341, n_232, n_6, n_69, n_317, n_353, n_321, n_73, n_320, n_77, n_260, n_37, n_97, n_186, n_138, n_379, n_374, n_26, n_235, n_378, n_245, n_161, n_189, n_271, n_2, n_145, n_227, n_92, n_330, n_388, n_395, n_332, n_292, n_116, n_94, n_289, n_280, n_333, n_213, n_356, n_184, n_28, n_372, n_202, n_56, n_370, n_34, n_98, n_384, n_121, n_352, n_125, n_216, n_82, n_327, n_47, n_106, n_32, n_263, n_230, n_51, n_248, n_301, n_27, n_343, n_369, n_174, n_18, n_104, n_211, n_281, n_173, n_234, n_284, n_153, n_316, n_75, n_178, n_298, n_49, n_43, n_297, n_383, n_9, n_119, n_310, n_164, n_231, n_44, n_102, n_122, n_141, n_128, n_111, n_167, n_80, n_179, n_12, n_68, n_129, n_345, n_304, n_381, n_311, n_324, n_25, n_278, n_236, n_367, n_267, n_218, n_48, n_204, n_339, n_89, n_277, n_331, n_93, n_182, n_363, n_323, n_199, n_350, n_142, n_223, n_67, n_368, n_250, n_85, n_45, n_5, n_244, n_118, n_139, n_87, n_171, n_78, n_146, n_17, n_226, n_255, n_286, n_120, n_261, n_238, n_391, n_360, n_58, n_165, n_361, n_246, n_176, n_163, n_29, n_52, n_251, n_220, n_387, n_197, n_296, n_3, n_41, n_256, n_71, n_302, n_351, n_126, n_200, n_115, n_96, n_110, n_392, n_150, n_147, n_288, n_23, n_334, n_274, n_160, n_303, n_95, n_188, n_269, n_201, n_306, n_158, n_4, n_366, n_346, n_193, n_397, n_293, n_162, n_358, n_385, n_275, n_214, n_46, n_109, n_59, n_203, n_81, n_133, n_377, n_273, n_114, n_276, n_295, n_382, n_265, n_354, n_154, n_127, n_326, n_24, n_217, n_55, n_62, n_291, n_148, n_88, n_159, n_11, n_108, n_373, n_60, n_233, n_290, n_365, n_155, n_243, n_268, n_136, n_157, n_282, n_389, n_101, n_309, n_344, n_229, n_107, n_33, n_53, n_36, n_149, n_190, n_262, n_134, n_349, n_336, n_195, n_300, n_252, n_283, n_314, n_249, n_221, n_156, n_359, n_57, n_66, n_21, n_31, n_8, n_312, n_183, n_266, n_205, n_335, n_177, n_313, n_22, n_140, n_219, n_180, n_212, n_210, n_325, n_338, n_371, n_103, n_166, n_224, n_151, n_130, n_253, n_99, n_15, n_72, n_152, n_198, n_7, n_228, n_272, n_196, n_347, n_315, n_123, n_279, n_79, n_270, n_305, n_117, n_208, n_215, n_135, n_70, n_50, n_170, n_86, n_375, n_340, n_13, n_380, n_394, n_168, n_175, n_241, n_105, n_84, n_294, n_393, n_258, n_206, n_307, n_396, n_342, n_348, n_14, n_194, n_137, n_225, n_16, n_39, n_337, n_247, n_240, n_38, n_259, n_143, n_192, n_0, n_264, n_63, n_1, n_237, n_91, n_398);
input n_76;
input n_113;
input n_187;
input n_90;
input n_257;
input n_390;
input n_65;
input n_74;
input n_185;
input n_285;
input n_30;
input n_222;
input n_61;
input n_20;
input n_287;
input n_357;
input n_386;
input n_64;
input n_254;
input n_207;
input n_10;
input n_83;
input n_181;
input n_362;
input n_124;
input n_191;
input n_209;
input n_299;
input n_322;
input n_328;
input n_19;
input n_40;
input n_318;
input n_355;
input n_239;
input n_100;
input n_54;
input n_112;
input n_319;
input n_364;
input n_35;
input n_42;
input n_329;
input n_132;
input n_131;
input n_144;
input n_169;
input n_242;
input n_376;
input n_308;
input n_172;
input n_341;
input n_232;
input n_6;
input n_69;
input n_317;
input n_353;
input n_321;
input n_73;
input n_320;
input n_77;
input n_260;
input n_37;
input n_97;
input n_186;
input n_138;
input n_379;
input n_374;
input n_26;
input n_235;
input n_378;
input n_245;
input n_161;
input n_189;
input n_271;
input n_2;
input n_145;
input n_227;
input n_92;
input n_330;
input n_388;
input n_395;
input n_332;
input n_292;
input n_116;
input n_94;
input n_289;
input n_280;
input n_333;
input n_213;
input n_356;
input n_184;
input n_28;
input n_372;
input n_202;
input n_56;
input n_370;
input n_34;
input n_98;
input n_384;
input n_121;
input n_352;
input n_125;
input n_216;
input n_82;
input n_327;
input n_47;
input n_106;
input n_32;
input n_263;
input n_230;
input n_51;
input n_248;
input n_301;
input n_27;
input n_343;
input n_369;
input n_174;
input n_18;
input n_104;
input n_211;
input n_281;
input n_173;
input n_234;
input n_284;
input n_153;
input n_316;
input n_75;
input n_178;
input n_298;
input n_49;
input n_43;
input n_297;
input n_383;
input n_9;
input n_119;
input n_310;
input n_164;
input n_231;
input n_44;
input n_102;
input n_122;
input n_141;
input n_128;
input n_111;
input n_167;
input n_80;
input n_179;
input n_12;
input n_68;
input n_129;
input n_345;
input n_304;
input n_381;
input n_311;
input n_324;
input n_25;
input n_278;
input n_236;
input n_367;
input n_267;
input n_218;
input n_48;
input n_204;
input n_339;
input n_89;
input n_277;
input n_331;
input n_93;
input n_182;
input n_363;
input n_323;
input n_199;
input n_350;
input n_142;
input n_223;
input n_67;
input n_368;
input n_250;
input n_85;
input n_45;
input n_5;
input n_244;
input n_118;
input n_139;
input n_87;
input n_171;
input n_78;
input n_146;
input n_17;
input n_226;
input n_255;
input n_286;
input n_120;
input n_261;
input n_238;
input n_391;
input n_360;
input n_58;
input n_165;
input n_361;
input n_246;
input n_176;
input n_163;
input n_29;
input n_52;
input n_251;
input n_220;
input n_387;
input n_197;
input n_296;
input n_3;
input n_41;
input n_256;
input n_71;
input n_302;
input n_351;
input n_126;
input n_200;
input n_115;
input n_96;
input n_110;
input n_392;
input n_150;
input n_147;
input n_288;
input n_23;
input n_334;
input n_274;
input n_160;
input n_303;
input n_95;
input n_188;
input n_269;
input n_201;
input n_306;
input n_158;
input n_4;
input n_366;
input n_346;
input n_193;
input n_397;
input n_293;
input n_162;
input n_358;
input n_385;
input n_275;
input n_214;
input n_46;
input n_109;
input n_59;
input n_203;
input n_81;
input n_133;
input n_377;
input n_273;
input n_114;
input n_276;
input n_295;
input n_382;
input n_265;
input n_354;
input n_154;
input n_127;
input n_326;
input n_24;
input n_217;
input n_55;
input n_62;
input n_291;
input n_148;
input n_88;
input n_159;
input n_11;
input n_108;
input n_373;
input n_60;
input n_233;
input n_290;
input n_365;
input n_155;
input n_243;
input n_268;
input n_136;
input n_157;
input n_282;
input n_389;
input n_101;
input n_309;
input n_344;
input n_229;
input n_107;
input n_33;
input n_53;
input n_36;
input n_149;
input n_190;
input n_262;
input n_134;
input n_349;
input n_336;
input n_195;
input n_300;
input n_252;
input n_283;
input n_314;
input n_249;
input n_221;
input n_156;
input n_359;
input n_57;
input n_66;
input n_21;
input n_31;
input n_8;
input n_312;
input n_183;
input n_266;
input n_205;
input n_335;
input n_177;
input n_313;
input n_22;
input n_140;
input n_219;
input n_180;
input n_212;
input n_210;
input n_325;
input n_338;
input n_371;
input n_103;
input n_166;
input n_224;
input n_151;
input n_130;
input n_253;
input n_99;
input n_15;
input n_72;
input n_152;
input n_198;
input n_7;
input n_228;
input n_272;
input n_196;
input n_347;
input n_315;
input n_123;
input n_279;
input n_79;
input n_270;
input n_305;
input n_117;
input n_208;
input n_215;
input n_135;
input n_70;
input n_50;
input n_170;
input n_86;
input n_375;
input n_340;
input n_13;
input n_380;
input n_394;
input n_168;
input n_175;
input n_241;
input n_105;
input n_84;
input n_294;
input n_393;
input n_258;
input n_206;
input n_307;
input n_396;
input n_342;
input n_348;
input n_14;
input n_194;
input n_137;
input n_225;
input n_16;
input n_39;
input n_337;
input n_247;
input n_240;
input n_38;
input n_259;
input n_143;
input n_192;
input n_0;
input n_264;
input n_63;
input n_1;
input n_237;
input n_91;
output n_398;
wire n_480;
wire n_1073;
wire n_476;
wire n_758;
wire n_599;
wire n_436;
wire n_887;
wire n_684;
wire n_1066;
wire n_1096;
wire n_821;
wire n_830;
wire n_624;
wire n_1018;
wire n_980;
wire n_800;
wire n_778;
wire n_618;
wire n_1106;
wire n_522;
wire n_1092;
wire n_838;
wire n_933;
wire n_485;
wire n_822;
wire n_846;
wire n_750;
wire n_631;
wire n_943;
wire n_977;
wire n_503;
wire n_635;
wire n_673;
wire n_792;
wire n_518;
wire n_905;
wire n_1067;
wire n_878;
wire n_665;
wire n_991;
wire n_667;
wire n_1114;
wire n_577;
wire n_1004;
wire n_580;
wire n_469;
wire n_987;
wire n_759;
wire n_979;
wire n_445;
wire n_1065;
wire n_596;
wire n_592;
wire n_540;
wire n_1064;
wire n_1075;
wire n_657;
wire n_900;
wire n_718;
wire n_841;
wire n_669;
wire n_1091;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_421;
wire n_555;
wire n_766;
wire n_852;
wire n_1113;
wire n_974;
wire n_919;
wire n_1089;
wire n_857;
wire n_461;
wire n_1047;
wire n_1016;
wire n_908;
wire n_549;
wire n_571;
wire n_694;
wire n_491;
wire n_923;
wire n_894;
wire n_1034;
wire n_952;
wire n_429;
wire n_1110;
wire n_752;
wire n_448;
wire n_545;
wire n_556;
wire n_593;
wire n_460;
wire n_937;
wire n_773;
wire n_989;
wire n_401;
wire n_538;
wire n_431;
wire n_1044;
wire n_963;
wire n_865;
wire n_666;
wire n_551;
wire n_884;
wire n_537;
wire n_560;
wire n_660;
wire n_1094;
wire n_814;
wire n_944;
wire n_886;
wire n_594;
wire n_856;
wire n_983;
wire n_767;
wire n_696;
wire n_889;
wire n_955;
wire n_975;
wire n_704;
wire n_941;
wire n_453;
wire n_932;
wire n_647;
wire n_948;
wire n_399;
wire n_700;
wire n_1021;
wire n_677;
wire n_958;
wire n_1046;
wire n_591;
wire n_775;
wire n_763;
wire n_1093;
wire n_1109;
wire n_870;
wire n_961;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_415;
wire n_572;
wire n_519;
wire n_815;
wire n_564;
wire n_638;
wire n_1116;
wire n_573;
wire n_510;
wire n_1099;
wire n_709;
wire n_786;
wire n_512;
wire n_795;
wire n_816;
wire n_539;
wire n_400;
wire n_626;
wire n_625;
wire n_953;
wire n_462;
wire n_615;
wire n_990;
wire n_550;
wire n_966;
wire n_1108;
wire n_670;
wire n_818;
wire n_716;
wire n_918;
wire n_883;
wire n_478;
wire n_584;
wire n_896;
wire n_408;
wire n_553;
wire n_892;
wire n_528;
wire n_1078;
wire n_495;
wire n_578;
wire n_994;
wire n_1072;
wire n_938;
wire n_744;
wire n_935;
wire n_824;
wire n_1098;
wire n_467;
wire n_875;
wire n_951;
wire n_774;
wire n_992;
wire n_813;
wire n_791;
wire n_981;
wire n_466;
wire n_559;
wire n_636;
wire n_872;
wire n_976;
wire n_1049;
wire n_906;
wire n_477;
wire n_515;
wire n_984;
wire n_1019;
wire n_680;
wire n_595;
wire n_1086;
wire n_726;
wire n_1070;
wire n_517;
wire n_683;
wire n_780;
wire n_904;
wire n_840;
wire n_570;
wire n_675;
wire n_931;
wire n_920;
wire n_530;
wire n_835;
wire n_535;
wire n_732;
wire n_834;
wire n_882;
wire n_784;
wire n_496;
wire n_693;
wire n_962;
wire n_1082;
wire n_468;
wire n_746;
wire n_532;
wire n_656;
wire n_755;
wire n_1025;
wire n_409;
wire n_860;
wire n_748;
wire n_781;
wire n_523;
wire n_909;
wire n_996;
wire n_439;
wire n_1062;
wire n_576;
wire n_924;
wire n_956;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_874;
wire n_801;
wire n_529;
wire n_1115;
wire n_455;
wire n_504;
wire n_725;
wire n_960;
wire n_671;
wire n_1081;
wire n_973;
wire n_1084;
wire n_659;
wire n_547;
wire n_682;
wire n_634;
wire n_903;
wire n_454;
wire n_812;
wire n_782;
wire n_443;
wire n_565;
wire n_817;
wire n_760;
wire n_608;
wire n_925;
wire n_534;
wire n_708;
wire n_1029;
wire n_1020;
wire n_457;
wire n_885;
wire n_1059;
wire n_950;
wire n_993;
wire n_493;
wire n_664;
wire n_819;
wire n_737;
wire n_1013;
wire n_1017;
wire n_581;
wire n_610;
wire n_936;
wire n_1035;
wire n_620;
wire n_582;
wire n_641;
wire n_1063;
wire n_828;
wire n_808;
wire n_770;
wire n_940;
wire n_745;
wire n_722;
wire n_867;
wire n_1100;
wire n_688;
wire n_609;
wire n_425;
wire n_1042;
wire n_879;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_1006;
wire n_690;
wire n_629;
wire n_1053;
wire n_499;
wire n_508;
wire n_706;
wire n_901;
wire n_561;
wire n_970;
wire n_947;
wire n_876;
wire n_1112;
wire n_437;
wire n_428;
wire n_405;
wire n_621;
wire n_783;
wire n_1107;
wire n_1012;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_769;
wire n_505;
wire n_527;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_1054;
wire n_672;
wire n_567;
wire n_916;
wire n_406;
wire n_1050;
wire n_426;
wire n_602;
wire n_617;
wire n_402;
wire n_552;
wire n_733;
wire n_658;
wire n_676;
wire n_986;
wire n_1083;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_880;
wire n_1031;
wire n_1037;
wire n_1103;
wire n_1008;
wire n_807;
wire n_1011;
wire n_416;
wire n_790;
wire n_895;
wire n_832;
wire n_410;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_913;
wire n_999;
wire n_619;
wire n_1095;
wire n_1060;
wire n_859;
wire n_695;
wire n_685;
wire n_881;
wire n_1080;
wire n_917;
wire n_632;
wire n_768;
wire n_412;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_985;
wire n_1077;
wire n_488;
wire n_501;
wire n_1041;
wire n_1111;
wire n_910;
wire n_869;
wire n_613;
wire n_642;
wire n_957;
wire n_995;
wire n_954;
wire n_702;
wire n_969;
wire n_912;
wire n_1009;
wire n_1007;
wire n_464;
wire n_945;
wire n_604;
wire n_734;
wire n_898;
wire n_848;
wire n_562;
wire n_1022;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_756;
wire n_569;
wire n_997;
wire n_563;
wire n_785;
wire n_891;
wire n_430;
wire n_568;
wire n_413;
wire n_471;
wire n_902;
wire n_1105;
wire n_853;
wire n_810;
wire n_843;
wire n_1079;
wire n_579;
wire n_1033;
wire n_699;
wire n_1003;
wire n_533;
wire n_1000;
wire n_1028;
wire n_727;
wire n_1014;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_914;
wire n_536;
wire n_707;
wire n_622;
wire n_470;
wire n_851;
wire n_915;
wire n_1002;
wire n_934;
wire n_494;
wire n_1001;
wire n_711;
wire n_864;
wire n_1027;
wire n_1058;
wire n_927;
wire n_1038;
wire n_965;
wire n_723;
wire n_662;
wire n_1085;
wire n_845;
wire n_850;
wire n_1043;
wire n_720;
wire n_968;
wire n_972;
wire n_435;
wire n_1026;
wire n_511;
wire n_484;
wire n_893;
wire n_492;
wire n_1068;
wire n_509;
wire n_407;
wire n_419;
wire n_730;
wire n_1023;
wire n_643;
wire n_747;
wire n_486;
wire n_930;
wire n_1057;
wire n_411;
wire n_697;
wire n_978;
wire n_907;
wire n_847;
wire n_779;
wire n_481;
wire n_691;
wire n_498;
wire n_765;
wire n_826;
wire n_648;
wire n_589;
wire n_628;
wire n_1005;
wire n_939;
wire n_487;
wire n_831;
wire n_653;
wire n_526;
wire n_637;
wire n_899;
wire n_928;
wire n_692;
wire n_544;
wire n_789;
wire n_1087;
wire n_1051;
wire n_738;
wire n_701;
wire n_827;
wire n_809;
wire n_482;
wire n_633;
wire n_520;
wire n_679;
wire n_922;
wire n_926;
wire n_942;
wire n_1048;
wire n_472;
wire n_971;
wire n_866;
wire n_452;
wire n_787;
wire n_1052;
wire n_1071;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_1097;
wire n_715;
wire n_959;
wire n_946;
wire n_420;
wire n_612;
wire n_858;
wire n_873;
wire n_438;
wire n_764;
wire n_794;
wire n_741;
wire n_753;
wire n_623;
wire n_1032;
wire n_446;
wire n_721;
wire n_681;
wire n_982;
wire n_456;
wire n_717;
wire n_1090;
wire n_712;
wire n_433;
wire n_516;
wire n_627;
wire n_739;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_524;
wire n_861;
wire n_705;
wire n_762;
wire n_575;
wire n_479;
wire n_442;
wire n_825;
wire n_698;
wire n_740;
wire n_541;
wire n_839;
wire n_546;
wire n_587;
wire n_639;
wire n_1010;
wire n_811;
wire n_1015;
wire n_459;
wire n_558;
wire n_863;
wire n_998;
wire n_724;
wire n_440;
wire n_525;
wire n_1074;
wire n_644;
wire n_674;
wire n_836;
wire n_888;
wire n_793;
wire n_1056;
wire n_583;
wire n_833;
wire n_414;
wire n_757;
wire n_929;
wire n_686;
wire n_776;
wire n_803;
wire n_890;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_949;
wire n_614;
wire n_586;
wire n_911;
wire n_772;
wire n_450;
wire n_788;
wire n_441;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_967;
wire n_837;
wire n_1045;
wire n_871;
wire n_474;
wire n_829;
wire n_1030;
wire n_988;
wire n_1055;
wire n_1088;
wire n_921;
wire n_597;
wire n_640;
wire n_483;
wire n_611;
wire n_1036;
wire n_687;
wire n_729;
wire n_844;
wire n_646;
wire n_650;
wire n_710;
wire n_743;
wire n_823;
wire n_652;
wire n_703;
wire n_1040;
wire n_500;
wire n_1101;
wire n_601;
wire n_661;
wire n_463;
wire n_1076;
wire n_804;
wire n_1102;
wire n_447;
wire n_603;
wire n_403;
wire n_854;
wire n_424;
wire n_877;
wire n_802;
wire n_868;
wire n_1039;
wire n_574;
wire n_1069;
wire n_1024;
wire n_842;
wire n_1104;
wire n_849;
wire n_1061;
wire n_475;
wire n_554;
wire n_897;
wire n_855;
wire n_798;
wire n_668;
wire n_797;
wire n_862;
AOI22xp33_ASAP7_75t_L g1035 ( .A1(n_0), .A2(n_346), .B1(n_603), .B2(n_762), .Y(n_1035) );
AOI22xp33_ASAP7_75t_L g977 ( .A1(n_1), .A2(n_233), .B1(n_609), .B2(n_610), .Y(n_977) );
CKINVDCx20_ASAP7_75t_R g752 ( .A(n_2), .Y(n_752) );
AOI22xp33_ASAP7_75t_L g814 ( .A1(n_3), .A2(n_87), .B1(n_518), .B2(n_815), .Y(n_814) );
AOI22xp5_ASAP7_75t_L g889 ( .A1(n_4), .A2(n_209), .B1(n_675), .B2(n_720), .Y(n_889) );
NAND2xp5_ASAP7_75t_L g1028 ( .A(n_5), .B(n_844), .Y(n_1028) );
AOI22xp5_ASAP7_75t_L g438 ( .A1(n_6), .A2(n_51), .B1(n_439), .B2(n_443), .Y(n_438) );
AOI22xp5_ASAP7_75t_L g557 ( .A1(n_7), .A2(n_105), .B1(n_558), .B2(n_560), .Y(n_557) );
AOI22xp33_ASAP7_75t_SL g916 ( .A1(n_8), .A2(n_344), .B1(n_475), .B2(n_534), .Y(n_916) );
AOI22xp33_ASAP7_75t_L g894 ( .A1(n_9), .A2(n_202), .B1(n_469), .B2(n_472), .Y(n_894) );
AOI22xp33_ASAP7_75t_L g648 ( .A1(n_10), .A2(n_301), .B1(n_519), .B2(n_649), .Y(n_648) );
AOI22xp33_ASAP7_75t_L g740 ( .A1(n_11), .A2(n_383), .B1(n_629), .B2(n_741), .Y(n_740) );
AOI22xp33_ASAP7_75t_L g566 ( .A1(n_12), .A2(n_258), .B1(n_567), .B2(n_569), .Y(n_566) );
AOI22xp33_ASAP7_75t_L g767 ( .A1(n_13), .A2(n_218), .B1(n_605), .B2(n_606), .Y(n_767) );
AOI22xp33_ASAP7_75t_L g536 ( .A1(n_14), .A2(n_83), .B1(n_470), .B2(n_472), .Y(n_536) );
AOI22xp33_ASAP7_75t_SL g780 ( .A1(n_15), .A2(n_86), .B1(n_528), .B2(n_598), .Y(n_780) );
AOI22xp33_ASAP7_75t_L g465 ( .A1(n_16), .A2(n_109), .B1(n_466), .B2(n_469), .Y(n_465) );
AOI22xp33_ASAP7_75t_L g531 ( .A1(n_17), .A2(n_342), .B1(n_477), .B2(n_532), .Y(n_531) );
AOI22xp33_ASAP7_75t_L g944 ( .A1(n_18), .A2(n_263), .B1(n_707), .B2(n_945), .Y(n_944) );
AOI22xp33_ASAP7_75t_L g717 ( .A1(n_19), .A2(n_88), .B1(n_718), .B2(n_720), .Y(n_717) );
AOI22xp33_ASAP7_75t_L g781 ( .A1(n_20), .A2(n_234), .B1(n_594), .B2(n_782), .Y(n_781) );
AOI22xp33_ASAP7_75t_L g654 ( .A1(n_21), .A2(n_193), .B1(n_517), .B2(n_575), .Y(n_654) );
AOI22xp33_ASAP7_75t_L g736 ( .A1(n_22), .A2(n_366), .B1(n_726), .B2(n_737), .Y(n_736) );
AOI22xp33_ASAP7_75t_L g498 ( .A1(n_23), .A2(n_155), .B1(n_429), .B2(n_499), .Y(n_498) );
AOI22xp33_ASAP7_75t_L g524 ( .A1(n_24), .A2(n_62), .B1(n_497), .B2(n_525), .Y(n_524) );
AO222x2_ASAP7_75t_L g755 ( .A1(n_25), .A2(n_150), .B1(n_259), .B2(n_540), .C1(n_542), .C2(n_543), .Y(n_755) );
CKINVDCx20_ASAP7_75t_R g924 ( .A(n_26), .Y(n_924) );
CKINVDCx20_ASAP7_75t_R g925 ( .A(n_27), .Y(n_925) );
AOI22xp33_ASAP7_75t_L g758 ( .A1(n_28), .A2(n_353), .B1(n_594), .B2(n_595), .Y(n_758) );
INVx1_ASAP7_75t_SL g417 ( .A(n_29), .Y(n_417) );
NOR2xp33_ASAP7_75t_L g1053 ( .A(n_29), .B(n_44), .Y(n_1053) );
AOI22xp33_ASAP7_75t_L g625 ( .A1(n_30), .A2(n_361), .B1(n_477), .B2(n_481), .Y(n_625) );
CKINVDCx20_ASAP7_75t_R g774 ( .A(n_31), .Y(n_774) );
AOI22xp5_ASAP7_75t_L g508 ( .A1(n_32), .A2(n_187), .B1(n_509), .B2(n_510), .Y(n_508) );
AOI22xp33_ASAP7_75t_SL g989 ( .A1(n_33), .A2(n_142), .B1(n_448), .B2(n_665), .Y(n_989) );
NAND2xp5_ASAP7_75t_L g743 ( .A(n_34), .B(n_410), .Y(n_743) );
AOI22xp33_ASAP7_75t_L g1039 ( .A1(n_35), .A2(n_311), .B1(n_605), .B2(n_606), .Y(n_1039) );
AOI22x1_ASAP7_75t_L g788 ( .A1(n_36), .A2(n_211), .B1(n_570), .B2(n_605), .Y(n_788) );
AOI22xp33_ASAP7_75t_L g593 ( .A1(n_37), .A2(n_127), .B1(n_594), .B2(n_595), .Y(n_593) );
AOI22xp33_ASAP7_75t_L g1012 ( .A1(n_38), .A2(n_232), .B1(n_479), .B2(n_718), .Y(n_1012) );
AOI22xp33_ASAP7_75t_L g628 ( .A1(n_39), .A2(n_229), .B1(n_429), .B2(n_629), .Y(n_628) );
OA22x2_ASAP7_75t_L g838 ( .A1(n_40), .A2(n_839), .B1(n_840), .B2(n_866), .Y(n_838) );
CKINVDCx20_ASAP7_75t_R g866 ( .A(n_40), .Y(n_866) );
AOI22xp33_ASAP7_75t_L g1111 ( .A1(n_41), .A2(n_297), .B1(n_507), .B2(n_1112), .Y(n_1111) );
AOI22xp33_ASAP7_75t_L g527 ( .A1(n_42), .A2(n_201), .B1(n_528), .B2(n_529), .Y(n_527) );
AOI22xp33_ASAP7_75t_L g734 ( .A1(n_43), .A2(n_345), .B1(n_466), .B2(n_677), .Y(n_734) );
AO22x2_ASAP7_75t_L g419 ( .A1(n_44), .A2(n_374), .B1(n_416), .B2(n_420), .Y(n_419) );
AOI22xp33_ASAP7_75t_L g795 ( .A1(n_45), .A2(n_225), .B1(n_458), .B2(n_519), .Y(n_795) );
AOI22xp33_ASAP7_75t_L g998 ( .A1(n_46), .A2(n_185), .B1(n_723), .B2(n_800), .Y(n_998) );
AOI22xp33_ASAP7_75t_L g1105 ( .A1(n_47), .A2(n_376), .B1(n_469), .B2(n_726), .Y(n_1105) );
AOI22xp33_ASAP7_75t_L g496 ( .A1(n_48), .A2(n_54), .B1(n_452), .B2(n_497), .Y(n_496) );
AOI22xp33_ASAP7_75t_L g951 ( .A1(n_49), .A2(n_158), .B1(n_677), .B2(n_952), .Y(n_951) );
AOI22xp33_ASAP7_75t_L g796 ( .A1(n_50), .A2(n_302), .B1(n_461), .B2(n_466), .Y(n_796) );
NAND2xp5_ASAP7_75t_L g1015 ( .A(n_52), .B(n_1016), .Y(n_1015) );
INVx1_ASAP7_75t_L g418 ( .A(n_53), .Y(n_418) );
AOI22xp33_ASAP7_75t_L g953 ( .A1(n_55), .A2(n_253), .B1(n_479), .B2(n_954), .Y(n_953) );
AOI22xp33_ASAP7_75t_L g428 ( .A1(n_56), .A2(n_317), .B1(n_429), .B2(n_434), .Y(n_428) );
AOI22xp33_ASAP7_75t_L g476 ( .A1(n_57), .A2(n_315), .B1(n_477), .B2(n_479), .Y(n_476) );
AOI22xp33_ASAP7_75t_SL g911 ( .A1(n_58), .A2(n_149), .B1(n_538), .B2(n_912), .Y(n_911) );
CKINVDCx20_ASAP7_75t_R g705 ( .A(n_59), .Y(n_705) );
AOI22xp5_ASAP7_75t_L g973 ( .A1(n_60), .A2(n_369), .B1(n_912), .B2(n_956), .Y(n_973) );
AOI22xp33_ASAP7_75t_L g537 ( .A1(n_61), .A2(n_324), .B1(n_474), .B2(n_538), .Y(n_537) );
AOI22xp5_ASAP7_75t_L g662 ( .A1(n_63), .A2(n_269), .B1(n_439), .B2(n_663), .Y(n_662) );
AOI22xp33_ASAP7_75t_L g1077 ( .A1(n_64), .A2(n_181), .B1(n_581), .B2(n_1078), .Y(n_1077) );
AOI22xp33_ASAP7_75t_L g679 ( .A1(n_65), .A2(n_227), .B1(n_469), .B2(n_680), .Y(n_679) );
NAND2xp5_ASAP7_75t_L g409 ( .A(n_66), .B(n_410), .Y(n_409) );
AO22x2_ASAP7_75t_L g426 ( .A1(n_67), .A2(n_206), .B1(n_416), .B2(n_427), .Y(n_426) );
AOI22xp33_ASAP7_75t_L g516 ( .A1(n_68), .A2(n_330), .B1(n_517), .B2(n_519), .Y(n_516) );
AOI22xp33_ASAP7_75t_L g576 ( .A1(n_69), .A2(n_90), .B1(n_515), .B2(n_577), .Y(n_576) );
AOI22xp33_ASAP7_75t_L g798 ( .A1(n_70), .A2(n_257), .B1(n_477), .B2(n_479), .Y(n_798) );
AOI22xp33_ASAP7_75t_L g620 ( .A1(n_71), .A2(n_152), .B1(n_509), .B2(n_621), .Y(n_620) );
AOI22xp33_ASAP7_75t_L g447 ( .A1(n_72), .A2(n_367), .B1(n_448), .B2(n_452), .Y(n_447) );
AOI22xp33_ASAP7_75t_L g986 ( .A1(n_73), .A2(n_119), .B1(n_778), .B2(n_987), .Y(n_986) );
AOI22xp33_ASAP7_75t_L g1083 ( .A1(n_74), .A2(n_249), .B1(n_563), .B2(n_970), .Y(n_1083) );
AOI22xp33_ASAP7_75t_L g1032 ( .A1(n_75), .A2(n_172), .B1(n_528), .B2(n_598), .Y(n_1032) );
AOI22xp33_ASAP7_75t_L g821 ( .A1(n_76), .A2(n_309), .B1(n_653), .B2(n_822), .Y(n_821) );
AOI22xp5_ASAP7_75t_L g789 ( .A1(n_77), .A2(n_176), .B1(n_606), .B2(n_612), .Y(n_789) );
AOI22xp33_ASAP7_75t_L g995 ( .A1(n_78), .A2(n_339), .B1(n_570), .B2(n_822), .Y(n_995) );
AOI22xp5_ASAP7_75t_L g676 ( .A1(n_79), .A2(n_216), .B1(n_466), .B2(n_677), .Y(n_676) );
AOI22xp33_ASAP7_75t_SL g913 ( .A1(n_80), .A2(n_347), .B1(n_718), .B2(n_914), .Y(n_913) );
AOI22xp5_ASAP7_75t_L g1036 ( .A1(n_81), .A2(n_166), .B1(n_570), .B2(n_723), .Y(n_1036) );
AOI22xp33_ASAP7_75t_SL g761 ( .A1(n_82), .A2(n_124), .B1(n_603), .B2(n_762), .Y(n_761) );
AOI22xp33_ASAP7_75t_L g1108 ( .A1(n_84), .A2(n_214), .B1(n_429), .B2(n_434), .Y(n_1108) );
AOI22xp33_ASAP7_75t_L g611 ( .A1(n_85), .A2(n_306), .B1(n_612), .B2(n_613), .Y(n_611) );
AOI22xp33_ASAP7_75t_L g1029 ( .A1(n_89), .A2(n_271), .B1(n_542), .B2(n_778), .Y(n_1029) );
AOI221xp5_ASAP7_75t_L g861 ( .A1(n_91), .A2(n_375), .B1(n_515), .B2(n_818), .C(n_862), .Y(n_861) );
AOI22xp33_ASAP7_75t_L g955 ( .A1(n_92), .A2(n_112), .B1(n_815), .B2(n_956), .Y(n_955) );
AOI222xp33_ASAP7_75t_L g1113 ( .A1(n_93), .A2(n_156), .B1(n_248), .B2(n_707), .C1(n_806), .C2(n_825), .Y(n_1113) );
NAND2xp5_ASAP7_75t_L g876 ( .A(n_94), .B(n_825), .Y(n_876) );
AOI22xp33_ASAP7_75t_SL g710 ( .A1(n_95), .A2(n_207), .B1(n_525), .B2(n_711), .Y(n_710) );
AOI22xp33_ASAP7_75t_L g1092 ( .A1(n_96), .A2(n_295), .B1(n_815), .B2(n_1093), .Y(n_1092) );
OAI22x1_ASAP7_75t_L g906 ( .A1(n_97), .A2(n_907), .B1(n_908), .B2(n_932), .Y(n_906) );
INVx1_ASAP7_75t_L g932 ( .A(n_97), .Y(n_932) );
AOI22xp5_ASAP7_75t_L g733 ( .A1(n_98), .A2(n_256), .B1(n_458), .B2(n_474), .Y(n_733) );
AOI22xp33_ASAP7_75t_L g645 ( .A1(n_99), .A2(n_387), .B1(n_439), .B2(n_443), .Y(n_645) );
AOI22xp33_ASAP7_75t_L g820 ( .A1(n_100), .A2(n_245), .B1(n_481), .B2(n_718), .Y(n_820) );
AOI22xp5_ASAP7_75t_L g803 ( .A1(n_101), .A2(n_325), .B1(n_741), .B2(n_804), .Y(n_803) );
AOI22xp5_ASAP7_75t_L g502 ( .A1(n_102), .A2(n_299), .B1(n_503), .B2(n_507), .Y(n_502) );
AOI22xp33_ASAP7_75t_L g681 ( .A1(n_103), .A2(n_143), .B1(n_682), .B2(n_683), .Y(n_681) );
AOI22xp33_ASAP7_75t_L g712 ( .A1(n_104), .A2(n_341), .B1(n_499), .B2(n_564), .Y(n_712) );
AOI22xp5_ASAP7_75t_L g1031 ( .A1(n_106), .A2(n_250), .B1(n_558), .B2(n_782), .Y(n_1031) );
AOI22xp5_ASAP7_75t_L g875 ( .A1(n_107), .A2(n_252), .B1(n_631), .B2(n_701), .Y(n_875) );
INVx1_ASAP7_75t_L g845 ( .A(n_108), .Y(n_845) );
AOI22xp33_ASAP7_75t_L g471 ( .A1(n_110), .A2(n_273), .B1(n_472), .B2(n_474), .Y(n_471) );
AOI222xp33_ASAP7_75t_L g805 ( .A1(n_111), .A2(n_189), .B1(n_359), .B2(n_443), .C1(n_492), .C2(n_806), .Y(n_805) );
AOI22xp33_ASAP7_75t_L g596 ( .A1(n_113), .A2(n_168), .B1(n_597), .B2(n_598), .Y(n_596) );
AOI22xp33_ASAP7_75t_L g562 ( .A1(n_114), .A2(n_292), .B1(n_434), .B2(n_563), .Y(n_562) );
AOI22xp33_ASAP7_75t_L g917 ( .A1(n_115), .A2(n_141), .B1(n_918), .B2(n_919), .Y(n_917) );
AOI22xp33_ASAP7_75t_L g571 ( .A1(n_116), .A2(n_255), .B1(n_532), .B2(n_572), .Y(n_571) );
AOI22xp5_ASAP7_75t_L g817 ( .A1(n_117), .A2(n_208), .B1(n_818), .B2(n_819), .Y(n_817) );
AOI22xp33_ASAP7_75t_L g928 ( .A1(n_118), .A2(n_226), .B1(n_711), .B2(n_929), .Y(n_928) );
AOI22xp33_ASAP7_75t_L g997 ( .A1(n_120), .A2(n_351), .B1(n_461), .B2(n_956), .Y(n_997) );
NAND2xp5_ASAP7_75t_L g940 ( .A(n_121), .B(n_941), .Y(n_940) );
AO22x2_ASAP7_75t_L g423 ( .A1(n_122), .A2(n_304), .B1(n_416), .B2(n_424), .Y(n_423) );
AOI22xp33_ASAP7_75t_L g643 ( .A1(n_123), .A2(n_323), .B1(n_499), .B2(n_644), .Y(n_643) );
CKINVDCx20_ASAP7_75t_R g854 ( .A(n_125), .Y(n_854) );
OAI22x1_ASAP7_75t_L g521 ( .A1(n_126), .A2(n_522), .B1(n_544), .B2(n_545), .Y(n_521) );
CKINVDCx16_ASAP7_75t_R g545 ( .A(n_126), .Y(n_545) );
AO21x2_ASAP7_75t_L g809 ( .A1(n_128), .A2(n_810), .B(n_832), .Y(n_809) );
NOR2xp33_ASAP7_75t_L g832 ( .A(n_128), .B(n_812), .Y(n_832) );
AOI22xp33_ASAP7_75t_L g828 ( .A1(n_129), .A2(n_133), .B1(n_579), .B2(n_581), .Y(n_828) );
AOI22xp33_ASAP7_75t_L g652 ( .A1(n_130), .A2(n_288), .B1(n_513), .B2(n_653), .Y(n_652) );
AOI22xp33_ASAP7_75t_L g1013 ( .A1(n_131), .A2(n_392), .B1(n_510), .B2(n_956), .Y(n_1013) );
AOI22xp33_ASAP7_75t_L g1110 ( .A1(n_132), .A2(n_241), .B1(n_461), .B2(n_892), .Y(n_1110) );
AOI22xp33_ASAP7_75t_L g739 ( .A1(n_134), .A2(n_265), .B1(n_665), .B2(n_666), .Y(n_739) );
AOI22xp33_ASAP7_75t_L g947 ( .A1(n_135), .A2(n_286), .B1(n_948), .B2(n_949), .Y(n_947) );
AOI22xp33_ASAP7_75t_L g715 ( .A1(n_136), .A2(n_268), .B1(n_677), .B2(n_716), .Y(n_715) );
INVx1_ASAP7_75t_L g807 ( .A(n_137), .Y(n_807) );
AOI22xp33_ASAP7_75t_L g601 ( .A1(n_138), .A2(n_365), .B1(n_602), .B2(n_603), .Y(n_601) );
OA22x2_ASAP7_75t_L g869 ( .A1(n_139), .A2(n_870), .B1(n_871), .B2(n_872), .Y(n_869) );
INVx1_ASAP7_75t_L g870 ( .A(n_139), .Y(n_870) );
AOI22xp33_ASAP7_75t_L g608 ( .A1(n_140), .A2(n_221), .B1(n_609), .B2(n_610), .Y(n_608) );
AOI22xp33_ASAP7_75t_L g725 ( .A1(n_144), .A2(n_254), .B1(n_470), .B2(n_726), .Y(n_725) );
AOI22xp33_ASAP7_75t_L g891 ( .A1(n_145), .A2(n_182), .B1(n_892), .B2(n_893), .Y(n_891) );
CKINVDCx20_ASAP7_75t_R g1040 ( .A(n_146), .Y(n_1040) );
AOI22xp33_ASAP7_75t_L g622 ( .A1(n_147), .A2(n_243), .B1(n_513), .B2(n_623), .Y(n_622) );
OA22x2_ASAP7_75t_L g936 ( .A1(n_148), .A2(n_937), .B1(n_938), .B2(n_958), .Y(n_936) );
CKINVDCx20_ASAP7_75t_R g937 ( .A(n_148), .Y(n_937) );
AOI22xp5_ASAP7_75t_L g670 ( .A1(n_151), .A2(n_180), .B1(n_429), .B2(n_671), .Y(n_670) );
AOI22xp5_ASAP7_75t_L g763 ( .A1(n_153), .A2(n_165), .B1(n_612), .B2(n_613), .Y(n_763) );
AOI22xp5_ASAP7_75t_L g664 ( .A1(n_154), .A2(n_348), .B1(n_665), .B2(n_666), .Y(n_664) );
CKINVDCx20_ASAP7_75t_R g878 ( .A(n_157), .Y(n_878) );
CKINVDCx20_ASAP7_75t_R g857 ( .A(n_159), .Y(n_857) );
AOI22xp33_ASAP7_75t_L g826 ( .A1(n_160), .A2(n_190), .B1(n_804), .B2(n_827), .Y(n_826) );
AOI22xp5_ASAP7_75t_L g457 ( .A1(n_161), .A2(n_238), .B1(n_458), .B2(n_461), .Y(n_457) );
AOI22xp5_ASAP7_75t_L g742 ( .A1(n_162), .A2(n_264), .B1(n_439), .B2(n_631), .Y(n_742) );
NAND2xp5_ASAP7_75t_L g848 ( .A(n_163), .B(n_582), .Y(n_848) );
BUFx2_ASAP7_75t_R g1097 ( .A(n_164), .Y(n_1097) );
AOI22xp33_ASAP7_75t_L g533 ( .A1(n_167), .A2(n_235), .B1(n_461), .B2(n_534), .Y(n_533) );
AOI22xp5_ASAP7_75t_L g888 ( .A1(n_169), .A2(n_393), .B1(n_677), .B2(n_716), .Y(n_888) );
NAND2xp5_ASAP7_75t_L g966 ( .A(n_170), .B(n_825), .Y(n_966) );
AOI22xp33_ASAP7_75t_L g974 ( .A1(n_171), .A2(n_307), .B1(n_481), .B2(n_675), .Y(n_974) );
NAND2xp5_ASAP7_75t_L g640 ( .A(n_173), .B(n_641), .Y(n_640) );
AOI22xp33_ASAP7_75t_L g957 ( .A1(n_174), .A2(n_200), .B1(n_623), .B2(n_822), .Y(n_957) );
AOI22xp33_ASAP7_75t_SL g994 ( .A1(n_175), .A2(n_337), .B1(n_477), .B2(n_651), .Y(n_994) );
AOI22xp33_ASAP7_75t_L g1104 ( .A1(n_177), .A2(n_310), .B1(n_458), .B2(n_519), .Y(n_1104) );
AOI22xp33_ASAP7_75t_SL g1090 ( .A1(n_178), .A2(n_251), .B1(n_567), .B2(n_819), .Y(n_1090) );
AOI22xp33_ASAP7_75t_L g1095 ( .A1(n_179), .A2(n_356), .B1(n_653), .B2(n_918), .Y(n_1095) );
AOI22xp33_ASAP7_75t_L g722 ( .A1(n_183), .A2(n_368), .B1(n_723), .B2(n_724), .Y(n_722) );
CKINVDCx20_ASAP7_75t_R g703 ( .A(n_184), .Y(n_703) );
AOI22xp33_ASAP7_75t_SL g1086 ( .A1(n_186), .A2(n_260), .B1(n_1087), .B2(n_1089), .Y(n_1086) );
AOI22xp33_ASAP7_75t_L g851 ( .A1(n_188), .A2(n_289), .B1(n_434), .B2(n_564), .Y(n_851) );
CKINVDCx20_ASAP7_75t_R g883 ( .A(n_191), .Y(n_883) );
NAND2xp5_ASAP7_75t_L g627 ( .A(n_192), .B(n_492), .Y(n_627) );
AOI22xp5_ASAP7_75t_L g1020 ( .A1(n_194), .A2(n_394), .B1(n_579), .B2(n_707), .Y(n_1020) );
CKINVDCx20_ASAP7_75t_R g847 ( .A(n_195), .Y(n_847) );
CKINVDCx20_ASAP7_75t_R g584 ( .A(n_196), .Y(n_584) );
AOI22xp33_ASAP7_75t_L g802 ( .A1(n_197), .A2(n_222), .B1(n_497), .B2(n_665), .Y(n_802) );
AOI22xp33_ASAP7_75t_L g632 ( .A1(n_198), .A2(n_283), .B1(n_452), .B2(n_497), .Y(n_632) );
AOI22xp33_ASAP7_75t_L g646 ( .A1(n_199), .A2(n_277), .B1(n_452), .B2(n_497), .Y(n_646) );
CKINVDCx20_ASAP7_75t_R g880 ( .A(n_203), .Y(n_880) );
AOI22xp33_ASAP7_75t_L g574 ( .A1(n_204), .A2(n_396), .B1(n_509), .B2(n_575), .Y(n_574) );
AOI22xp33_ASAP7_75t_L g1018 ( .A1(n_205), .A2(n_272), .B1(n_563), .B2(n_970), .Y(n_1018) );
INVx1_ASAP7_75t_L g1052 ( .A(n_206), .Y(n_1052) );
AOI22xp33_ASAP7_75t_L g604 ( .A1(n_210), .A2(n_247), .B1(n_605), .B2(n_606), .Y(n_604) );
AOI22xp33_ASAP7_75t_L g785 ( .A1(n_212), .A2(n_278), .B1(n_603), .B2(n_762), .Y(n_785) );
CKINVDCx20_ASAP7_75t_R g860 ( .A(n_213), .Y(n_860) );
AOI22xp33_ASAP7_75t_L g931 ( .A1(n_215), .A2(n_331), .B1(n_804), .B2(n_827), .Y(n_931) );
XNOR2xp5_ASAP7_75t_L g768 ( .A(n_217), .B(n_769), .Y(n_768) );
XNOR2xp5_ASAP7_75t_L g791 ( .A(n_217), .B(n_769), .Y(n_791) );
CKINVDCx20_ASAP7_75t_R g859 ( .A(n_219), .Y(n_859) );
AOI22xp5_ASAP7_75t_L g968 ( .A1(n_220), .A2(n_377), .B1(n_497), .B2(n_525), .Y(n_968) );
OAI22xp5_ASAP7_75t_L g405 ( .A1(n_223), .A2(n_406), .B1(n_407), .B2(n_483), .Y(n_405) );
INVxp67_ASAP7_75t_L g483 ( .A(n_223), .Y(n_483) );
CKINVDCx20_ASAP7_75t_R g863 ( .A(n_224), .Y(n_863) );
AOI22xp33_ASAP7_75t_L g1007 ( .A1(n_228), .A2(n_298), .B1(n_1008), .B2(n_1009), .Y(n_1007) );
AOI22xp33_ASAP7_75t_L g1010 ( .A1(n_230), .A2(n_333), .B1(n_623), .B2(n_822), .Y(n_1010) );
OA22x2_ASAP7_75t_L g729 ( .A1(n_231), .A2(n_730), .B1(n_731), .B2(n_744), .Y(n_729) );
INVxp67_ASAP7_75t_L g744 ( .A(n_231), .Y(n_744) );
OA22x2_ASAP7_75t_L g746 ( .A1(n_231), .A2(n_730), .B1(n_731), .B2(n_744), .Y(n_746) );
INVx2_ASAP7_75t_L g1065 ( .A(n_236), .Y(n_1065) );
AOI22xp33_ASAP7_75t_L g765 ( .A1(n_237), .A2(n_388), .B1(n_610), .B2(n_766), .Y(n_765) );
OA22x2_ASAP7_75t_L g658 ( .A1(n_239), .A2(n_659), .B1(n_685), .B2(n_686), .Y(n_658) );
CKINVDCx20_ASAP7_75t_R g685 ( .A(n_239), .Y(n_685) );
AOI22xp33_ASAP7_75t_SL g512 ( .A1(n_240), .A2(n_293), .B1(n_513), .B2(n_515), .Y(n_512) );
AOI22xp33_ASAP7_75t_L g799 ( .A1(n_242), .A2(n_266), .B1(n_680), .B2(n_800), .Y(n_799) );
CKINVDCx20_ASAP7_75t_R g922 ( .A(n_244), .Y(n_922) );
INVx1_ASAP7_75t_L g1076 ( .A(n_246), .Y(n_1076) );
AOI22xp33_ASAP7_75t_L g674 ( .A1(n_261), .A2(n_300), .B1(n_507), .B2(n_675), .Y(n_674) );
CKINVDCx20_ASAP7_75t_R g864 ( .A(n_262), .Y(n_864) );
CKINVDCx16_ASAP7_75t_R g614 ( .A(n_267), .Y(n_614) );
AOI22xp33_ASAP7_75t_L g990 ( .A1(n_270), .A2(n_358), .B1(n_943), .B2(n_991), .Y(n_990) );
AOI22xp5_ASAP7_75t_L g591 ( .A1(n_274), .A2(n_355), .B1(n_542), .B2(n_543), .Y(n_591) );
CKINVDCx20_ASAP7_75t_R g772 ( .A(n_275), .Y(n_772) );
AOI22xp33_ASAP7_75t_L g850 ( .A1(n_276), .A2(n_322), .B1(n_497), .B2(n_525), .Y(n_850) );
AOI22xp5_ASAP7_75t_L g494 ( .A1(n_279), .A2(n_290), .B1(n_439), .B2(n_443), .Y(n_494) );
AOI22xp33_ASAP7_75t_L g942 ( .A1(n_280), .A2(n_336), .B1(n_629), .B2(n_943), .Y(n_942) );
AOI22xp33_ASAP7_75t_SL g757 ( .A1(n_281), .A2(n_303), .B1(n_597), .B2(n_598), .Y(n_757) );
AO22x2_ASAP7_75t_L g616 ( .A1(n_282), .A2(n_617), .B1(n_633), .B2(n_634), .Y(n_616) );
CKINVDCx20_ASAP7_75t_R g633 ( .A(n_282), .Y(n_633) );
AOI22xp33_ASAP7_75t_L g786 ( .A1(n_284), .A2(n_397), .B1(n_609), .B2(n_610), .Y(n_786) );
NAND2xp5_ASAP7_75t_L g824 ( .A(n_285), .B(n_825), .Y(n_824) );
AOI22xp5_ASAP7_75t_L g965 ( .A1(n_287), .A2(n_320), .B1(n_443), .B2(n_701), .Y(n_965) );
AOI22x1_ASAP7_75t_L g486 ( .A1(n_291), .A2(n_487), .B1(n_488), .B2(n_520), .Y(n_486) );
INVx1_ASAP7_75t_L g520 ( .A(n_291), .Y(n_520) );
XNOR2x1_ASAP7_75t_L g548 ( .A(n_291), .B(n_488), .Y(n_548) );
AOI22xp5_ASAP7_75t_L g976 ( .A1(n_294), .A2(n_373), .B1(n_474), .B2(n_538), .Y(n_976) );
OA22x2_ASAP7_75t_L g1002 ( .A1(n_296), .A2(n_1003), .B1(n_1004), .B2(n_1005), .Y(n_1002) );
INVx1_ASAP7_75t_L g1003 ( .A(n_296), .Y(n_1003) );
NOR2xp33_ASAP7_75t_L g1050 ( .A(n_304), .B(n_1051), .Y(n_1050) );
AOI22xp33_ASAP7_75t_L g630 ( .A1(n_305), .A2(n_371), .B1(n_439), .B2(n_631), .Y(n_630) );
AOI222xp33_ASAP7_75t_L g539 ( .A1(n_308), .A2(n_321), .B1(n_354), .B2(n_540), .C1(n_541), .C2(n_543), .Y(n_539) );
NAND2xp5_ASAP7_75t_L g668 ( .A(n_312), .B(n_410), .Y(n_668) );
AOI22xp33_ASAP7_75t_L g1080 ( .A1(n_313), .A2(n_360), .B1(n_525), .B2(n_1081), .Y(n_1080) );
AOI22xp33_ASAP7_75t_L g650 ( .A1(n_314), .A2(n_395), .B1(n_477), .B2(n_651), .Y(n_650) );
CKINVDCx20_ASAP7_75t_R g708 ( .A(n_316), .Y(n_708) );
CKINVDCx20_ASAP7_75t_R g776 ( .A(n_318), .Y(n_776) );
AOI22xp33_ASAP7_75t_L g829 ( .A1(n_319), .A2(n_349), .B1(n_560), .B2(n_830), .Y(n_829) );
CKINVDCx20_ASAP7_75t_R g493 ( .A(n_326), .Y(n_493) );
AOI22xp5_ASAP7_75t_L g735 ( .A1(n_327), .A2(n_338), .B1(n_572), .B2(n_651), .Y(n_735) );
INVx1_ASAP7_75t_L g727 ( .A(n_328), .Y(n_727) );
INVx3_ASAP7_75t_L g416 ( .A(n_329), .Y(n_416) );
AOI22xp33_ASAP7_75t_L g1038 ( .A1(n_332), .A2(n_340), .B1(n_610), .B2(n_766), .Y(n_1038) );
AOI222xp33_ASAP7_75t_L g578 ( .A1(n_334), .A2(n_372), .B1(n_384), .B2(n_410), .C1(n_579), .C2(n_581), .Y(n_578) );
OAI22x1_ASAP7_75t_L g637 ( .A1(n_335), .A2(n_638), .B1(n_655), .B2(n_656), .Y(n_637) );
INVx1_ASAP7_75t_L g656 ( .A(n_335), .Y(n_656) );
CKINVDCx20_ASAP7_75t_R g978 ( .A(n_343), .Y(n_978) );
AOI22xp5_ASAP7_75t_L g1019 ( .A1(n_350), .A2(n_380), .B1(n_525), .B2(n_830), .Y(n_1019) );
AOI22xp33_ASAP7_75t_L g619 ( .A1(n_352), .A2(n_385), .B1(n_466), .B2(n_519), .Y(n_619) );
CKINVDCx20_ASAP7_75t_R g985 ( .A(n_357), .Y(n_985) );
CKINVDCx20_ASAP7_75t_R g885 ( .A(n_362), .Y(n_885) );
INVx1_ASAP7_75t_L g981 ( .A(n_363), .Y(n_981) );
AOI22xp33_ASAP7_75t_L g969 ( .A1(n_364), .A2(n_391), .B1(n_429), .B2(n_970), .Y(n_969) );
AOI22xp33_ASAP7_75t_L g1107 ( .A1(n_370), .A2(n_382), .B1(n_497), .B2(n_665), .Y(n_1107) );
INVx1_ASAP7_75t_L g1047 ( .A(n_378), .Y(n_1047) );
NAND2xp5_ASAP7_75t_SL g1064 ( .A(n_378), .B(n_1065), .Y(n_1064) );
INVx1_ASAP7_75t_L g1066 ( .A(n_379), .Y(n_1066) );
INVx1_ASAP7_75t_L g1048 ( .A(n_381), .Y(n_1048) );
AND2x2_ASAP7_75t_R g1114 ( .A(n_381), .B(n_1047), .Y(n_1114) );
INVxp67_ASAP7_75t_L g1063 ( .A(n_386), .Y(n_1063) );
NAND2xp5_ASAP7_75t_L g590 ( .A(n_389), .B(n_540), .Y(n_590) );
XOR2xp5_ASAP7_75t_L g1100 ( .A(n_390), .B(n_1101), .Y(n_1100) );
AOI21xp5_ASAP7_75t_L g398 ( .A1(n_399), .A2(n_1054), .B(n_1057), .Y(n_398) );
AOI21xp33_ASAP7_75t_L g399 ( .A1(n_400), .A2(n_903), .B(n_1044), .Y(n_399) );
INVx1_ASAP7_75t_L g1056 ( .A(n_400), .Y(n_1056) );
AOI22xp5_ASAP7_75t_L g400 ( .A1(n_401), .A2(n_692), .B1(n_901), .B2(n_902), .Y(n_400) );
INVx1_ASAP7_75t_L g901 ( .A(n_401), .Y(n_901) );
AOI22xp5_ASAP7_75t_L g401 ( .A1(n_402), .A2(n_551), .B1(n_690), .B2(n_691), .Y(n_401) );
INVx2_ASAP7_75t_L g690 ( .A(n_402), .Y(n_690) );
INVx2_ASAP7_75t_SL g402 ( .A(n_403), .Y(n_402) );
OA22x2_ASAP7_75t_L g403 ( .A1(n_404), .A2(n_484), .B1(n_549), .B2(n_550), .Y(n_403) );
HB1xp67_ASAP7_75t_SL g404 ( .A(n_405), .Y(n_404) );
INVx2_ASAP7_75t_L g549 ( .A(n_405), .Y(n_549) );
INVx1_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
NOR2xp67_ASAP7_75t_L g407 ( .A(n_408), .B(n_456), .Y(n_407) );
NAND4xp25_ASAP7_75t_L g408 ( .A(n_409), .B(n_428), .C(n_438), .D(n_447), .Y(n_408) );
HB1xp67_ASAP7_75t_L g941 ( .A(n_410), .Y(n_941) );
INVx3_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
INVx4_ASAP7_75t_SL g492 ( .A(n_411), .Y(n_492) );
INVx3_ASAP7_75t_SL g642 ( .A(n_411), .Y(n_642) );
INVx3_ASAP7_75t_L g825 ( .A(n_411), .Y(n_825) );
INVx4_ASAP7_75t_SL g844 ( .A(n_411), .Y(n_844) );
BUFx2_ASAP7_75t_L g923 ( .A(n_411), .Y(n_923) );
INVx6_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
AND2x2_ASAP7_75t_L g412 ( .A(n_413), .B(n_421), .Y(n_412) );
AND2x4_ASAP7_75t_L g436 ( .A(n_413), .B(n_437), .Y(n_436) );
AND2x4_ASAP7_75t_L g453 ( .A(n_413), .B(n_454), .Y(n_453) );
AND2x2_ASAP7_75t_L g529 ( .A(n_413), .B(n_437), .Y(n_529) );
AND2x4_ASAP7_75t_L g540 ( .A(n_413), .B(n_421), .Y(n_540) );
AND2x2_ASAP7_75t_L g595 ( .A(n_413), .B(n_454), .Y(n_595) );
AND2x2_ASAP7_75t_L g598 ( .A(n_413), .B(n_437), .Y(n_598) );
AND2x2_ASAP7_75t_L g782 ( .A(n_413), .B(n_454), .Y(n_782) );
AND2x2_ASAP7_75t_L g413 ( .A(n_414), .B(n_419), .Y(n_413) );
INVx2_ASAP7_75t_L g433 ( .A(n_414), .Y(n_433) );
AND2x2_ASAP7_75t_L g441 ( .A(n_414), .B(n_442), .Y(n_441) );
HB1xp67_ASAP7_75t_L g446 ( .A(n_414), .Y(n_446) );
OAI22x1_ASAP7_75t_L g414 ( .A1(n_415), .A2(n_416), .B1(n_417), .B2(n_418), .Y(n_414) );
INVx1_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
INVx1_ASAP7_75t_L g420 ( .A(n_416), .Y(n_420) );
INVx2_ASAP7_75t_L g424 ( .A(n_416), .Y(n_424) );
INVx1_ASAP7_75t_L g427 ( .A(n_416), .Y(n_427) );
AND2x2_ASAP7_75t_L g432 ( .A(n_419), .B(n_433), .Y(n_432) );
INVx2_ASAP7_75t_L g442 ( .A(n_419), .Y(n_442) );
BUFx2_ASAP7_75t_L g482 ( .A(n_419), .Y(n_482) );
AND2x2_ASAP7_75t_L g460 ( .A(n_421), .B(n_432), .Y(n_460) );
AND2x4_ASAP7_75t_L g468 ( .A(n_421), .B(n_464), .Y(n_468) );
AND2x4_ASAP7_75t_L g473 ( .A(n_421), .B(n_441), .Y(n_473) );
AND2x6_ASAP7_75t_L g605 ( .A(n_421), .B(n_432), .Y(n_605) );
AND2x2_ASAP7_75t_L g609 ( .A(n_421), .B(n_441), .Y(n_609) );
AND2x2_ASAP7_75t_L g612 ( .A(n_421), .B(n_464), .Y(n_612) );
AND2x2_ASAP7_75t_L g766 ( .A(n_421), .B(n_441), .Y(n_766) );
AND2x4_ASAP7_75t_L g421 ( .A(n_422), .B(n_425), .Y(n_421) );
INVx1_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
AND2x4_ASAP7_75t_L g431 ( .A(n_423), .B(n_425), .Y(n_431) );
AND2x2_ASAP7_75t_L g445 ( .A(n_423), .B(n_426), .Y(n_445) );
INVx1_ASAP7_75t_L g451 ( .A(n_423), .Y(n_451) );
INVxp67_ASAP7_75t_L g437 ( .A(n_425), .Y(n_437) );
INVx2_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
AND2x2_ASAP7_75t_L g450 ( .A(n_426), .B(n_451), .Y(n_450) );
BUFx3_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
BUFx6f_ASAP7_75t_L g564 ( .A(n_430), .Y(n_564) );
BUFx2_ASAP7_75t_L g741 ( .A(n_430), .Y(n_741) );
BUFx2_ASAP7_75t_L g943 ( .A(n_430), .Y(n_943) );
AND2x4_ASAP7_75t_L g430 ( .A(n_431), .B(n_432), .Y(n_430) );
AND2x2_ASAP7_75t_L g440 ( .A(n_431), .B(n_441), .Y(n_440) );
AND2x4_ASAP7_75t_L g475 ( .A(n_431), .B(n_464), .Y(n_475) );
AND2x2_ASAP7_75t_L g528 ( .A(n_431), .B(n_432), .Y(n_528) );
AND2x4_ASAP7_75t_L g542 ( .A(n_431), .B(n_441), .Y(n_542) );
AND2x2_ASAP7_75t_L g597 ( .A(n_431), .B(n_432), .Y(n_597) );
AND2x2_ASAP7_75t_L g613 ( .A(n_431), .B(n_464), .Y(n_613) );
AND2x2_ASAP7_75t_L g478 ( .A(n_432), .B(n_450), .Y(n_478) );
AND2x2_ASAP7_75t_L g602 ( .A(n_432), .B(n_450), .Y(n_602) );
AND2x2_ASAP7_75t_SL g762 ( .A(n_432), .B(n_450), .Y(n_762) );
AND2x4_ASAP7_75t_L g464 ( .A(n_433), .B(n_442), .Y(n_464) );
INVx2_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
INVx2_ASAP7_75t_SL g499 ( .A(n_435), .Y(n_499) );
INVx1_ASAP7_75t_L g629 ( .A(n_435), .Y(n_629) );
INVx2_ASAP7_75t_SL g671 ( .A(n_435), .Y(n_671) );
INVx2_ASAP7_75t_L g804 ( .A(n_435), .Y(n_804) );
OAI22xp5_ASAP7_75t_L g882 ( .A1(n_435), .A2(n_883), .B1(n_884), .B2(n_885), .Y(n_882) );
INVx2_ASAP7_75t_L g970 ( .A(n_435), .Y(n_970) );
INVx2_ASAP7_75t_L g991 ( .A(n_435), .Y(n_991) );
INVx6_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
BUFx5_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
BUFx3_ASAP7_75t_L g580 ( .A(n_440), .Y(n_580) );
INVx2_ASAP7_75t_L g702 ( .A(n_440), .Y(n_702) );
BUFx3_ASAP7_75t_L g946 ( .A(n_440), .Y(n_946) );
AND2x2_ASAP7_75t_L g449 ( .A(n_441), .B(n_450), .Y(n_449) );
AND2x4_ASAP7_75t_L g594 ( .A(n_441), .B(n_450), .Y(n_594) );
BUFx3_ASAP7_75t_L g707 ( .A(n_443), .Y(n_707) );
INVx2_ASAP7_75t_L g926 ( .A(n_443), .Y(n_926) );
BUFx12f_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
INVx3_ASAP7_75t_L g583 ( .A(n_444), .Y(n_583) );
AND2x2_ASAP7_75t_L g444 ( .A(n_445), .B(n_446), .Y(n_444) );
AND2x4_ASAP7_75t_L g470 ( .A(n_445), .B(n_464), .Y(n_470) );
AND2x4_ASAP7_75t_L g481 ( .A(n_445), .B(n_482), .Y(n_481) );
AND2x2_ASAP7_75t_SL g543 ( .A(n_445), .B(n_446), .Y(n_543) );
AND2x4_ASAP7_75t_L g603 ( .A(n_445), .B(n_482), .Y(n_603) );
AND2x4_ASAP7_75t_L g610 ( .A(n_445), .B(n_464), .Y(n_610) );
AND2x2_ASAP7_75t_SL g778 ( .A(n_445), .B(n_446), .Y(n_778) );
INVx1_ASAP7_75t_L g879 ( .A(n_448), .Y(n_879) );
HB1xp67_ASAP7_75t_L g948 ( .A(n_448), .Y(n_948) );
BUFx6f_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
BUFx6f_ASAP7_75t_L g497 ( .A(n_449), .Y(n_497) );
INVx3_ASAP7_75t_L g559 ( .A(n_449), .Y(n_559) );
AND2x4_ASAP7_75t_L g463 ( .A(n_450), .B(n_464), .Y(n_463) );
AND2x6_ASAP7_75t_L g606 ( .A(n_450), .B(n_464), .Y(n_606) );
HB1xp67_ASAP7_75t_L g455 ( .A(n_451), .Y(n_455) );
BUFx4f_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
INVx2_ASAP7_75t_L g526 ( .A(n_453), .Y(n_526) );
BUFx3_ASAP7_75t_L g561 ( .A(n_453), .Y(n_561) );
BUFx6f_ASAP7_75t_SL g665 ( .A(n_453), .Y(n_665) );
INVx1_ASAP7_75t_L g930 ( .A(n_453), .Y(n_930) );
INVx1_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
NAND4xp25_ASAP7_75t_L g456 ( .A(n_457), .B(n_465), .C(n_471), .D(n_476), .Y(n_456) );
INVx2_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
INVx2_ASAP7_75t_SL g509 ( .A(n_459), .Y(n_509) );
INVx2_ASAP7_75t_SL g649 ( .A(n_459), .Y(n_649) );
INVx2_ASAP7_75t_L g682 ( .A(n_459), .Y(n_682) );
INVx3_ASAP7_75t_L g956 ( .A(n_459), .Y(n_956) );
INVx3_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
BUFx2_ASAP7_75t_L g534 ( .A(n_460), .Y(n_534) );
BUFx2_ASAP7_75t_L g716 ( .A(n_460), .Y(n_716) );
INVx2_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
INVx2_ASAP7_75t_SL g510 ( .A(n_462), .Y(n_510) );
INVx2_ASAP7_75t_L g575 ( .A(n_462), .Y(n_575) );
INVx1_ASAP7_75t_SL g621 ( .A(n_462), .Y(n_621) );
INVx2_ASAP7_75t_L g677 ( .A(n_462), .Y(n_677) );
INVx2_ASAP7_75t_L g819 ( .A(n_462), .Y(n_819) );
HB1xp67_ASAP7_75t_L g865 ( .A(n_462), .Y(n_865) );
INVx2_ASAP7_75t_SL g912 ( .A(n_462), .Y(n_912) );
INVx8_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
BUFx2_ASAP7_75t_L g1008 ( .A(n_466), .Y(n_1008) );
INVx2_ASAP7_75t_SL g466 ( .A(n_467), .Y(n_466) );
INVx4_ASAP7_75t_L g518 ( .A(n_467), .Y(n_518) );
INVx2_ASAP7_75t_L g538 ( .A(n_467), .Y(n_538) );
INVx3_ASAP7_75t_SL g723 ( .A(n_467), .Y(n_723) );
INVx2_ASAP7_75t_SL g892 ( .A(n_467), .Y(n_892) );
INVx8_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
BUFx3_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
BUFx2_ASAP7_75t_SL g515 ( .A(n_470), .Y(n_515) );
INVx2_ASAP7_75t_L g624 ( .A(n_470), .Y(n_624) );
BUFx2_ASAP7_75t_SL g653 ( .A(n_470), .Y(n_653) );
BUFx3_ASAP7_75t_L g800 ( .A(n_470), .Y(n_800) );
BUFx3_ASAP7_75t_L g472 ( .A(n_473), .Y(n_472) );
INVx6_ASAP7_75t_L g514 ( .A(n_473), .Y(n_514) );
BUFx3_ASAP7_75t_L g822 ( .A(n_473), .Y(n_822) );
HB1xp67_ASAP7_75t_L g724 ( .A(n_474), .Y(n_724) );
BUFx6f_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
BUFx3_ASAP7_75t_L g519 ( .A(n_475), .Y(n_519) );
BUFx6f_ASAP7_75t_L g570 ( .A(n_475), .Y(n_570) );
INVx2_ASAP7_75t_L g684 ( .A(n_475), .Y(n_684) );
BUFx6f_ASAP7_75t_L g477 ( .A(n_478), .Y(n_477) );
INVx2_ASAP7_75t_L g506 ( .A(n_478), .Y(n_506) );
BUFx3_ASAP7_75t_L g675 ( .A(n_478), .Y(n_675) );
INVx2_ASAP7_75t_L g479 ( .A(n_480), .Y(n_479) );
INVx3_ASAP7_75t_L g507 ( .A(n_480), .Y(n_507) );
OAI22xp33_ASAP7_75t_L g853 ( .A1(n_480), .A2(n_854), .B1(n_855), .B2(n_857), .Y(n_853) );
INVx2_ASAP7_75t_L g914 ( .A(n_480), .Y(n_914) );
INVx2_ASAP7_75t_L g1089 ( .A(n_480), .Y(n_1089) );
INVx5_ASAP7_75t_SL g480 ( .A(n_481), .Y(n_480) );
BUFx2_ASAP7_75t_L g532 ( .A(n_481), .Y(n_532) );
BUFx2_ASAP7_75t_L g651 ( .A(n_481), .Y(n_651) );
BUFx3_ASAP7_75t_L g720 ( .A(n_481), .Y(n_720) );
INVx2_ASAP7_75t_L g550 ( .A(n_484), .Y(n_550) );
AO22x2_ASAP7_75t_L g484 ( .A1(n_485), .A2(n_521), .B1(n_546), .B2(n_547), .Y(n_484) );
INVx1_ASAP7_75t_L g485 ( .A(n_486), .Y(n_485) );
INVx2_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
AND2x4_ASAP7_75t_L g488 ( .A(n_489), .B(n_500), .Y(n_488) );
NOR2xp67_ASAP7_75t_L g489 ( .A(n_490), .B(n_495), .Y(n_489) );
OAI21xp5_ASAP7_75t_SL g490 ( .A1(n_491), .A2(n_493), .B(n_494), .Y(n_490) );
INVx1_ASAP7_75t_L g491 ( .A(n_492), .Y(n_491) );
NAND2xp5_ASAP7_75t_L g495 ( .A(n_496), .B(n_498), .Y(n_495) );
BUFx6f_ASAP7_75t_SL g711 ( .A(n_497), .Y(n_711) );
NOR2x1_ASAP7_75t_L g500 ( .A(n_501), .B(n_511), .Y(n_500) );
NAND2xp5_ASAP7_75t_L g501 ( .A(n_502), .B(n_508), .Y(n_501) );
INVx1_ASAP7_75t_L g503 ( .A(n_504), .Y(n_503) );
INVx1_ASAP7_75t_L g856 ( .A(n_504), .Y(n_856) );
INVx1_ASAP7_75t_L g504 ( .A(n_505), .Y(n_504) );
BUFx6f_ASAP7_75t_L g572 ( .A(n_505), .Y(n_572) );
INVx1_ASAP7_75t_L g1088 ( .A(n_505), .Y(n_1088) );
INVx2_ASAP7_75t_L g505 ( .A(n_506), .Y(n_505) );
INVx1_ASAP7_75t_L g719 ( .A(n_506), .Y(n_719) );
NAND2xp5_ASAP7_75t_L g511 ( .A(n_512), .B(n_516), .Y(n_511) );
INVx2_ASAP7_75t_L g513 ( .A(n_514), .Y(n_513) );
INVx2_ASAP7_75t_L g577 ( .A(n_514), .Y(n_577) );
INVx2_ASAP7_75t_L g680 ( .A(n_514), .Y(n_680) );
INVx3_ASAP7_75t_L g726 ( .A(n_514), .Y(n_726) );
OAI22xp5_ASAP7_75t_L g862 ( .A1(n_514), .A2(n_863), .B1(n_864), .B2(n_865), .Y(n_862) );
INVx1_ASAP7_75t_SL g918 ( .A(n_514), .Y(n_918) );
BUFx6f_ASAP7_75t_L g517 ( .A(n_518), .Y(n_517) );
INVx2_ASAP7_75t_L g568 ( .A(n_518), .Y(n_568) );
BUFx2_ASAP7_75t_L g1009 ( .A(n_519), .Y(n_1009) );
INVx2_ASAP7_75t_L g546 ( .A(n_521), .Y(n_546) );
NAND4xp25_ASAP7_75t_SL g522 ( .A(n_523), .B(n_530), .C(n_535), .D(n_539), .Y(n_522) );
AND4x1_ASAP7_75t_L g544 ( .A(n_523), .B(n_530), .C(n_535), .D(n_539), .Y(n_544) );
AND2x2_ASAP7_75t_L g523 ( .A(n_524), .B(n_527), .Y(n_523) );
INVx2_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
AND2x2_ASAP7_75t_L g530 ( .A(n_531), .B(n_533), .Y(n_530) );
INVx2_ASAP7_75t_L g1094 ( .A(n_534), .Y(n_1094) );
AND2x2_ASAP7_75t_L g535 ( .A(n_536), .B(n_537), .Y(n_535) );
INVx2_ASAP7_75t_SL g773 ( .A(n_540), .Y(n_773) );
HB1xp67_ASAP7_75t_L g541 ( .A(n_542), .Y(n_541) );
INVx1_ASAP7_75t_SL g775 ( .A(n_542), .Y(n_775) );
INVx1_ASAP7_75t_L g547 ( .A(n_548), .Y(n_547) );
INVx1_ASAP7_75t_L g691 ( .A(n_551), .Y(n_691) );
AOI22xp5_ASAP7_75t_L g551 ( .A1(n_552), .A2(n_615), .B1(n_688), .B2(n_689), .Y(n_551) );
INVx1_ASAP7_75t_L g688 ( .A(n_552), .Y(n_688) );
OA22x2_ASAP7_75t_L g552 ( .A1(n_553), .A2(n_554), .B1(n_585), .B2(n_586), .Y(n_552) );
INVx2_ASAP7_75t_SL g553 ( .A(n_554), .Y(n_553) );
XNOR2x1_ASAP7_75t_L g554 ( .A(n_555), .B(n_584), .Y(n_554) );
NAND4xp75_ASAP7_75t_L g555 ( .A(n_556), .B(n_565), .C(n_573), .D(n_578), .Y(n_555) );
AND2x2_ASAP7_75t_L g556 ( .A(n_557), .B(n_562), .Y(n_556) );
INVx2_ASAP7_75t_SL g1082 ( .A(n_558), .Y(n_1082) );
INVx4_ASAP7_75t_L g558 ( .A(n_559), .Y(n_558) );
INVx2_ASAP7_75t_L g666 ( .A(n_559), .Y(n_666) );
INVx1_ASAP7_75t_L g831 ( .A(n_559), .Y(n_831) );
BUFx6f_ASAP7_75t_SL g560 ( .A(n_561), .Y(n_560) );
BUFx2_ASAP7_75t_L g563 ( .A(n_564), .Y(n_563) );
BUFx4f_ASAP7_75t_SL g644 ( .A(n_564), .Y(n_644) );
BUFx2_ASAP7_75t_L g827 ( .A(n_564), .Y(n_827) );
INVx1_ASAP7_75t_L g884 ( .A(n_564), .Y(n_884) );
AND2x2_ASAP7_75t_L g565 ( .A(n_566), .B(n_571), .Y(n_565) );
INVx1_ASAP7_75t_L g567 ( .A(n_568), .Y(n_567) );
OAI22xp33_ASAP7_75t_L g858 ( .A1(n_568), .A2(n_816), .B1(n_859), .B2(n_860), .Y(n_858) );
BUFx6f_ASAP7_75t_L g569 ( .A(n_570), .Y(n_569) );
INVx2_ASAP7_75t_L g816 ( .A(n_570), .Y(n_816) );
AND2x2_ASAP7_75t_L g573 ( .A(n_574), .B(n_576), .Y(n_573) );
INVx1_ASAP7_75t_L g846 ( .A(n_579), .Y(n_846) );
BUFx6f_ASAP7_75t_SL g579 ( .A(n_580), .Y(n_579) );
BUFx6f_ASAP7_75t_L g581 ( .A(n_582), .Y(n_581) );
INVx3_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
INVx2_ASAP7_75t_L g631 ( .A(n_583), .Y(n_631) );
INVx2_ASAP7_75t_L g663 ( .A(n_583), .Y(n_663) );
INVx2_ASAP7_75t_L g585 ( .A(n_586), .Y(n_585) );
AO22x2_ASAP7_75t_L g868 ( .A1(n_586), .A2(n_869), .B1(n_895), .B2(n_896), .Y(n_868) );
INVx1_ASAP7_75t_L g896 ( .A(n_586), .Y(n_896) );
XOR2x2_ASAP7_75t_L g586 ( .A(n_587), .B(n_614), .Y(n_586) );
NAND2x1p5_ASAP7_75t_L g587 ( .A(n_588), .B(n_599), .Y(n_587) );
NOR2x1_ASAP7_75t_L g588 ( .A(n_589), .B(n_592), .Y(n_588) );
NAND2xp5_ASAP7_75t_L g589 ( .A(n_590), .B(n_591), .Y(n_589) );
NAND2xp5_ASAP7_75t_L g592 ( .A(n_593), .B(n_596), .Y(n_592) );
NOR2x1_ASAP7_75t_L g599 ( .A(n_600), .B(n_607), .Y(n_599) );
NAND2xp5_ASAP7_75t_L g600 ( .A(n_601), .B(n_604), .Y(n_600) );
NAND2xp5_ASAP7_75t_L g607 ( .A(n_608), .B(n_611), .Y(n_607) );
INVx1_ASAP7_75t_L g689 ( .A(n_615), .Y(n_689) );
XNOR2xp5_ASAP7_75t_L g615 ( .A(n_616), .B(n_635), .Y(n_615) );
INVx1_ASAP7_75t_SL g634 ( .A(n_617), .Y(n_634) );
NOR2x1_ASAP7_75t_L g617 ( .A(n_618), .B(n_626), .Y(n_617) );
NAND4xp25_ASAP7_75t_L g618 ( .A(n_619), .B(n_620), .C(n_622), .D(n_625), .Y(n_618) );
INVx2_ASAP7_75t_SL g623 ( .A(n_624), .Y(n_623) );
INVx2_ASAP7_75t_SL g737 ( .A(n_624), .Y(n_737) );
NAND4xp25_ASAP7_75t_SL g626 ( .A(n_627), .B(n_628), .C(n_630), .D(n_632), .Y(n_626) );
AO22x2_ASAP7_75t_L g635 ( .A1(n_636), .A2(n_637), .B1(n_657), .B2(n_658), .Y(n_635) );
INVx1_ASAP7_75t_L g636 ( .A(n_637), .Y(n_636) );
INVx1_ASAP7_75t_L g655 ( .A(n_638), .Y(n_655) );
OR2x2_ASAP7_75t_L g638 ( .A(n_639), .B(n_647), .Y(n_638) );
NAND4xp25_ASAP7_75t_L g639 ( .A(n_640), .B(n_643), .C(n_645), .D(n_646), .Y(n_639) );
INVx3_ASAP7_75t_L g704 ( .A(n_641), .Y(n_704) );
BUFx6f_ASAP7_75t_L g641 ( .A(n_642), .Y(n_641) );
INVx2_ASAP7_75t_L g1017 ( .A(n_642), .Y(n_1017) );
NAND4xp25_ASAP7_75t_L g647 ( .A(n_648), .B(n_650), .C(n_652), .D(n_654), .Y(n_647) );
INVx2_ASAP7_75t_L g657 ( .A(n_658), .Y(n_657) );
NAND2xp5_ASAP7_75t_L g659 ( .A(n_660), .B(n_672), .Y(n_659) );
NOR3xp33_ASAP7_75t_L g660 ( .A(n_661), .B(n_667), .C(n_669), .Y(n_660) );
NOR4xp25_ASAP7_75t_L g686 ( .A(n_661), .B(n_673), .C(n_678), .D(n_687), .Y(n_686) );
NAND2xp5_ASAP7_75t_L g661 ( .A(n_662), .B(n_664), .Y(n_661) );
INVxp67_ASAP7_75t_L g881 ( .A(n_665), .Y(n_881) );
BUFx2_ASAP7_75t_SL g949 ( .A(n_665), .Y(n_949) );
INVxp67_ASAP7_75t_L g667 ( .A(n_668), .Y(n_667) );
NAND2xp5_ASAP7_75t_L g687 ( .A(n_668), .B(n_670), .Y(n_687) );
INVxp67_ASAP7_75t_SL g669 ( .A(n_670), .Y(n_669) );
NOR2xp33_ASAP7_75t_L g672 ( .A(n_673), .B(n_678), .Y(n_672) );
NAND2xp5_ASAP7_75t_L g673 ( .A(n_674), .B(n_676), .Y(n_673) );
BUFx2_ASAP7_75t_L g954 ( .A(n_675), .Y(n_954) );
NAND2xp5_ASAP7_75t_L g678 ( .A(n_679), .B(n_681), .Y(n_678) );
INVx2_ASAP7_75t_L g683 ( .A(n_684), .Y(n_683) );
INVx1_ASAP7_75t_L g893 ( .A(n_684), .Y(n_893) );
INVx2_ASAP7_75t_L g902 ( .A(n_692), .Y(n_902) );
XNOR2x1_ASAP7_75t_L g692 ( .A(n_693), .B(n_835), .Y(n_692) );
OA22x2_ASAP7_75t_L g693 ( .A1(n_694), .A2(n_747), .B1(n_748), .B2(n_834), .Y(n_693) );
INVx1_ASAP7_75t_L g834 ( .A(n_694), .Y(n_834) );
OAI22xp5_ASAP7_75t_L g694 ( .A1(n_695), .A2(n_728), .B1(n_745), .B2(n_746), .Y(n_694) );
INVx3_ASAP7_75t_L g745 ( .A(n_695), .Y(n_745) );
XOR2x2_ASAP7_75t_L g695 ( .A(n_696), .B(n_727), .Y(n_695) );
NAND2xp5_ASAP7_75t_SL g696 ( .A(n_697), .B(n_713), .Y(n_696) );
NOR2x1_ASAP7_75t_L g697 ( .A(n_698), .B(n_709), .Y(n_697) );
OAI222xp33_ASAP7_75t_L g698 ( .A1(n_699), .A2(n_703), .B1(n_704), .B2(n_705), .C1(n_706), .C2(n_708), .Y(n_698) );
INVx1_ASAP7_75t_L g699 ( .A(n_700), .Y(n_699) );
HB1xp67_ASAP7_75t_L g700 ( .A(n_701), .Y(n_700) );
INVx2_ASAP7_75t_L g701 ( .A(n_702), .Y(n_701) );
INVx1_ASAP7_75t_L g806 ( .A(n_702), .Y(n_806) );
INVx2_ASAP7_75t_L g1078 ( .A(n_702), .Y(n_1078) );
INVx1_ASAP7_75t_L g706 ( .A(n_707), .Y(n_706) );
NAND2xp5_ASAP7_75t_L g709 ( .A(n_710), .B(n_712), .Y(n_709) );
NOR2xp33_ASAP7_75t_L g713 ( .A(n_714), .B(n_721), .Y(n_713) );
NAND2xp5_ASAP7_75t_L g714 ( .A(n_715), .B(n_717), .Y(n_714) );
BUFx3_ASAP7_75t_L g818 ( .A(n_716), .Y(n_818) );
BUFx6f_ASAP7_75t_L g718 ( .A(n_719), .Y(n_718) );
NAND2xp5_ASAP7_75t_L g721 ( .A(n_722), .B(n_725), .Y(n_721) );
INVx1_ASAP7_75t_L g728 ( .A(n_729), .Y(n_728) );
INVx2_ASAP7_75t_SL g730 ( .A(n_731), .Y(n_730) );
NOR2x1_ASAP7_75t_L g731 ( .A(n_732), .B(n_738), .Y(n_731) );
NAND4xp25_ASAP7_75t_SL g732 ( .A(n_733), .B(n_734), .C(n_735), .D(n_736), .Y(n_732) );
NAND4xp25_ASAP7_75t_L g738 ( .A(n_739), .B(n_740), .C(n_742), .D(n_743), .Y(n_738) );
INVx2_ASAP7_75t_L g747 ( .A(n_748), .Y(n_747) );
AOI22x1_ASAP7_75t_L g748 ( .A1(n_749), .A2(n_808), .B1(n_809), .B2(n_833), .Y(n_748) );
INVx2_ASAP7_75t_L g833 ( .A(n_749), .Y(n_833) );
XNOR2x1_ASAP7_75t_L g749 ( .A(n_750), .B(n_792), .Y(n_749) );
OAI21xp5_ASAP7_75t_L g750 ( .A1(n_751), .A2(n_768), .B(n_790), .Y(n_750) );
NAND2xp5_ASAP7_75t_L g790 ( .A(n_751), .B(n_791), .Y(n_790) );
XNOR2x1_ASAP7_75t_L g751 ( .A(n_752), .B(n_753), .Y(n_751) );
AND2x2_ASAP7_75t_L g753 ( .A(n_754), .B(n_759), .Y(n_753) );
NOR2xp33_ASAP7_75t_L g754 ( .A(n_755), .B(n_756), .Y(n_754) );
NAND2xp5_ASAP7_75t_L g756 ( .A(n_757), .B(n_758), .Y(n_756) );
NOR2xp33_ASAP7_75t_L g759 ( .A(n_760), .B(n_764), .Y(n_759) );
NAND2xp5_ASAP7_75t_L g760 ( .A(n_761), .B(n_763), .Y(n_760) );
NAND2xp5_ASAP7_75t_L g764 ( .A(n_765), .B(n_767), .Y(n_764) );
NAND2x1p5_ASAP7_75t_L g769 ( .A(n_770), .B(n_783), .Y(n_769) );
NOR2x1_ASAP7_75t_L g770 ( .A(n_771), .B(n_779), .Y(n_770) );
OAI222xp33_ASAP7_75t_L g771 ( .A1(n_772), .A2(n_773), .B1(n_774), .B2(n_775), .C1(n_776), .C2(n_777), .Y(n_771) );
OAI21xp5_ASAP7_75t_SL g984 ( .A1(n_773), .A2(n_985), .B(n_986), .Y(n_984) );
INVx1_ASAP7_75t_L g987 ( .A(n_775), .Y(n_987) );
INVxp67_ASAP7_75t_L g777 ( .A(n_778), .Y(n_777) );
NAND2xp5_ASAP7_75t_L g779 ( .A(n_780), .B(n_781), .Y(n_779) );
NOR2x1_ASAP7_75t_L g783 ( .A(n_784), .B(n_787), .Y(n_783) );
NAND2xp5_ASAP7_75t_L g784 ( .A(n_785), .B(n_786), .Y(n_784) );
NAND2xp5_ASAP7_75t_L g787 ( .A(n_788), .B(n_789), .Y(n_787) );
HB1xp67_ASAP7_75t_L g899 ( .A(n_791), .Y(n_899) );
XOR2x2_ASAP7_75t_L g792 ( .A(n_793), .B(n_807), .Y(n_792) );
NAND4xp75_ASAP7_75t_L g793 ( .A(n_794), .B(n_797), .C(n_801), .D(n_805), .Y(n_793) );
AND2x2_ASAP7_75t_L g794 ( .A(n_795), .B(n_796), .Y(n_794) );
AND2x2_ASAP7_75t_L g797 ( .A(n_798), .B(n_799), .Y(n_797) );
BUFx6f_ASAP7_75t_L g919 ( .A(n_800), .Y(n_919) );
AND2x2_ASAP7_75t_L g801 ( .A(n_802), .B(n_803), .Y(n_801) );
INVx2_ASAP7_75t_L g808 ( .A(n_809), .Y(n_808) );
INVx1_ASAP7_75t_L g810 ( .A(n_811), .Y(n_810) );
INVx1_ASAP7_75t_L g811 ( .A(n_812), .Y(n_811) );
NOR2xp33_ASAP7_75t_L g812 ( .A(n_813), .B(n_823), .Y(n_812) );
NAND4xp25_ASAP7_75t_SL g813 ( .A(n_814), .B(n_817), .C(n_820), .D(n_821), .Y(n_813) );
INVx2_ASAP7_75t_L g815 ( .A(n_816), .Y(n_815) );
NAND4xp25_ASAP7_75t_SL g823 ( .A(n_824), .B(n_826), .C(n_828), .D(n_829), .Y(n_823) );
BUFx3_ASAP7_75t_L g830 ( .A(n_831), .Y(n_830) );
OAI22xp5_ASAP7_75t_L g835 ( .A1(n_836), .A2(n_837), .B1(n_867), .B2(n_900), .Y(n_835) );
INVx1_ASAP7_75t_L g836 ( .A(n_837), .Y(n_836) );
INVx1_ASAP7_75t_L g837 ( .A(n_838), .Y(n_837) );
INVx2_ASAP7_75t_L g839 ( .A(n_840), .Y(n_839) );
AND3x2_ASAP7_75t_L g840 ( .A(n_841), .B(n_852), .C(n_861), .Y(n_840) );
NOR2xp33_ASAP7_75t_L g841 ( .A(n_842), .B(n_849), .Y(n_841) );
OAI221xp5_ASAP7_75t_L g842 ( .A1(n_843), .A2(n_845), .B1(n_846), .B2(n_847), .C(n_848), .Y(n_842) );
INVx1_ASAP7_75t_SL g843 ( .A(n_844), .Y(n_843) );
OAI222xp33_ASAP7_75t_L g921 ( .A1(n_846), .A2(n_922), .B1(n_923), .B2(n_924), .C1(n_925), .C2(n_926), .Y(n_921) );
NAND2xp5_ASAP7_75t_L g849 ( .A(n_850), .B(n_851), .Y(n_849) );
NOR2xp33_ASAP7_75t_L g852 ( .A(n_853), .B(n_858), .Y(n_852) );
INVx1_ASAP7_75t_L g855 ( .A(n_856), .Y(n_855) );
INVx2_ASAP7_75t_L g900 ( .A(n_867), .Y(n_900) );
XNOR2x1_ASAP7_75t_L g867 ( .A(n_868), .B(n_897), .Y(n_867) );
INVx1_ASAP7_75t_L g895 ( .A(n_869), .Y(n_895) );
INVx2_ASAP7_75t_L g871 ( .A(n_872), .Y(n_871) );
AND2x2_ASAP7_75t_L g872 ( .A(n_873), .B(n_886), .Y(n_872) );
NOR3xp33_ASAP7_75t_L g873 ( .A(n_874), .B(n_877), .C(n_882), .Y(n_873) );
NAND2xp5_ASAP7_75t_L g874 ( .A(n_875), .B(n_876), .Y(n_874) );
OAI22xp5_ASAP7_75t_L g877 ( .A1(n_878), .A2(n_879), .B1(n_880), .B2(n_881), .Y(n_877) );
NOR2xp33_ASAP7_75t_L g886 ( .A(n_887), .B(n_890), .Y(n_886) );
NAND2xp5_ASAP7_75t_L g887 ( .A(n_888), .B(n_889), .Y(n_887) );
NAND2xp5_ASAP7_75t_L g890 ( .A(n_891), .B(n_894), .Y(n_890) );
BUFx2_ASAP7_75t_L g952 ( .A(n_892), .Y(n_952) );
INVx2_ASAP7_75t_L g897 ( .A(n_898), .Y(n_897) );
INVx2_ASAP7_75t_L g898 ( .A(n_899), .Y(n_898) );
INVx1_ASAP7_75t_L g1055 ( .A(n_903), .Y(n_1055) );
AOI22xp33_ASAP7_75t_SL g903 ( .A1(n_904), .A2(n_905), .B1(n_933), .B2(n_1043), .Y(n_903) );
INVx2_ASAP7_75t_L g904 ( .A(n_905), .Y(n_904) );
BUFx3_ASAP7_75t_L g905 ( .A(n_906), .Y(n_905) );
INVx2_ASAP7_75t_L g907 ( .A(n_908), .Y(n_907) );
AND2x4_ASAP7_75t_L g908 ( .A(n_909), .B(n_920), .Y(n_908) );
NOR2x1_ASAP7_75t_L g909 ( .A(n_910), .B(n_915), .Y(n_909) );
NAND2xp5_ASAP7_75t_L g910 ( .A(n_911), .B(n_913), .Y(n_910) );
NAND2xp5_ASAP7_75t_L g915 ( .A(n_916), .B(n_917), .Y(n_915) );
NOR2x1_ASAP7_75t_L g920 ( .A(n_921), .B(n_927), .Y(n_920) );
NAND2xp5_ASAP7_75t_L g927 ( .A(n_928), .B(n_931), .Y(n_927) );
INVx2_ASAP7_75t_SL g929 ( .A(n_930), .Y(n_929) );
INVx1_ASAP7_75t_L g1043 ( .A(n_933), .Y(n_1043) );
AOI22xp5_ASAP7_75t_L g933 ( .A1(n_934), .A2(n_1000), .B1(n_1041), .B2(n_1042), .Y(n_933) );
INVx2_ASAP7_75t_L g1041 ( .A(n_934), .Y(n_1041) );
AOI22x1_ASAP7_75t_SL g934 ( .A1(n_935), .A2(n_936), .B1(n_959), .B2(n_999), .Y(n_934) );
INVx1_ASAP7_75t_L g935 ( .A(n_936), .Y(n_935) );
INVx1_ASAP7_75t_L g958 ( .A(n_938), .Y(n_958) );
OR2x2_ASAP7_75t_L g938 ( .A(n_939), .B(n_950), .Y(n_938) );
NAND4xp25_ASAP7_75t_SL g939 ( .A(n_940), .B(n_942), .C(n_944), .D(n_947), .Y(n_939) );
BUFx6f_ASAP7_75t_L g945 ( .A(n_946), .Y(n_945) );
NAND4xp25_ASAP7_75t_L g950 ( .A(n_951), .B(n_953), .C(n_955), .D(n_957), .Y(n_950) );
INVx2_ASAP7_75t_L g999 ( .A(n_959), .Y(n_999) );
OA22x2_ASAP7_75t_L g959 ( .A1(n_960), .A2(n_961), .B1(n_979), .B2(n_980), .Y(n_959) );
INVx2_ASAP7_75t_L g960 ( .A(n_961), .Y(n_960) );
XOR2x2_ASAP7_75t_L g961 ( .A(n_962), .B(n_978), .Y(n_961) );
NAND2x1p5_ASAP7_75t_L g962 ( .A(n_963), .B(n_971), .Y(n_962) );
NOR2x1_ASAP7_75t_L g963 ( .A(n_964), .B(n_967), .Y(n_963) );
NAND2xp5_ASAP7_75t_L g964 ( .A(n_965), .B(n_966), .Y(n_964) );
NAND2xp5_ASAP7_75t_L g967 ( .A(n_968), .B(n_969), .Y(n_967) );
NOR2x1_ASAP7_75t_L g971 ( .A(n_972), .B(n_975), .Y(n_971) );
NAND2xp5_ASAP7_75t_L g972 ( .A(n_973), .B(n_974), .Y(n_972) );
NAND2xp5_ASAP7_75t_L g975 ( .A(n_976), .B(n_977), .Y(n_975) );
OAI22xp5_ASAP7_75t_L g1022 ( .A1(n_979), .A2(n_980), .B1(n_1023), .B2(n_1024), .Y(n_1022) );
INVx2_ASAP7_75t_SL g979 ( .A(n_980), .Y(n_979) );
XNOR2x1_ASAP7_75t_L g980 ( .A(n_981), .B(n_982), .Y(n_980) );
NAND2x1_ASAP7_75t_L g982 ( .A(n_983), .B(n_992), .Y(n_982) );
NOR2xp67_ASAP7_75t_L g983 ( .A(n_984), .B(n_988), .Y(n_983) );
NAND2xp5_ASAP7_75t_L g988 ( .A(n_989), .B(n_990), .Y(n_988) );
NOR2xp33_ASAP7_75t_L g992 ( .A(n_993), .B(n_996), .Y(n_992) );
NAND2xp5_ASAP7_75t_L g993 ( .A(n_994), .B(n_995), .Y(n_993) );
NAND2xp5_ASAP7_75t_L g996 ( .A(n_997), .B(n_998), .Y(n_996) );
INVx3_ASAP7_75t_L g1042 ( .A(n_1000), .Y(n_1042) );
OA22x2_ASAP7_75t_L g1000 ( .A1(n_1001), .A2(n_1002), .B1(n_1021), .B2(n_1022), .Y(n_1000) );
INVx1_ASAP7_75t_L g1001 ( .A(n_1002), .Y(n_1001) );
INVx1_ASAP7_75t_L g1004 ( .A(n_1005), .Y(n_1004) );
NOR3x1_ASAP7_75t_SL g1005 ( .A(n_1006), .B(n_1011), .C(n_1014), .Y(n_1005) );
NAND2xp5_ASAP7_75t_L g1006 ( .A(n_1007), .B(n_1010), .Y(n_1006) );
NAND2xp5_ASAP7_75t_L g1011 ( .A(n_1012), .B(n_1013), .Y(n_1011) );
NAND4xp25_ASAP7_75t_SL g1014 ( .A(n_1015), .B(n_1018), .C(n_1019), .D(n_1020), .Y(n_1014) );
INVx2_ASAP7_75t_L g1016 ( .A(n_1017), .Y(n_1016) );
OAI21xp5_ASAP7_75t_SL g1075 ( .A1(n_1017), .A2(n_1076), .B(n_1077), .Y(n_1075) );
INVx1_ASAP7_75t_L g1021 ( .A(n_1022), .Y(n_1021) );
INVx1_ASAP7_75t_SL g1023 ( .A(n_1024), .Y(n_1023) );
XOR2x2_ASAP7_75t_L g1024 ( .A(n_1025), .B(n_1040), .Y(n_1024) );
NAND2xp5_ASAP7_75t_SL g1025 ( .A(n_1026), .B(n_1033), .Y(n_1025) );
NOR2xp33_ASAP7_75t_L g1026 ( .A(n_1027), .B(n_1030), .Y(n_1026) );
NAND2xp5_ASAP7_75t_L g1027 ( .A(n_1028), .B(n_1029), .Y(n_1027) );
NAND2xp5_ASAP7_75t_L g1030 ( .A(n_1031), .B(n_1032), .Y(n_1030) );
NOR2xp33_ASAP7_75t_L g1033 ( .A(n_1034), .B(n_1037), .Y(n_1033) );
NAND2xp5_ASAP7_75t_L g1034 ( .A(n_1035), .B(n_1036), .Y(n_1034) );
NAND2xp5_ASAP7_75t_L g1037 ( .A(n_1038), .B(n_1039), .Y(n_1037) );
INVx2_ASAP7_75t_SL g1044 ( .A(n_1045), .Y(n_1044) );
AND2x2_ASAP7_75t_L g1045 ( .A(n_1046), .B(n_1049), .Y(n_1045) );
NAND2xp5_ASAP7_75t_L g1099 ( .A(n_1046), .B(n_1050), .Y(n_1099) );
NOR2xp33_ASAP7_75t_L g1046 ( .A(n_1047), .B(n_1048), .Y(n_1046) );
INVx1_ASAP7_75t_L g1061 ( .A(n_1048), .Y(n_1061) );
INVx1_ASAP7_75t_L g1049 ( .A(n_1050), .Y(n_1049) );
NAND2xp5_ASAP7_75t_L g1051 ( .A(n_1052), .B(n_1053), .Y(n_1051) );
NAND2xp5_ASAP7_75t_L g1054 ( .A(n_1055), .B(n_1056), .Y(n_1054) );
OAI21xp5_ASAP7_75t_L g1057 ( .A1(n_1058), .A2(n_1066), .B(n_1067), .Y(n_1057) );
CKINVDCx20_ASAP7_75t_R g1058 ( .A(n_1059), .Y(n_1058) );
AND2x4_ASAP7_75t_SL g1059 ( .A(n_1060), .B(n_1062), .Y(n_1059) );
INVx1_ASAP7_75t_L g1060 ( .A(n_1061), .Y(n_1060) );
OR2x2_ASAP7_75t_L g1116 ( .A(n_1061), .B(n_1062), .Y(n_1116) );
NOR2xp33_ASAP7_75t_L g1062 ( .A(n_1063), .B(n_1064), .Y(n_1062) );
AOI222xp33_ASAP7_75t_L g1067 ( .A1(n_1068), .A2(n_1097), .B1(n_1098), .B2(n_1100), .C1(n_1114), .C2(n_1115), .Y(n_1067) );
INVx2_ASAP7_75t_L g1068 ( .A(n_1069), .Y(n_1068) );
INVx2_ASAP7_75t_L g1069 ( .A(n_1070), .Y(n_1069) );
INVx1_ASAP7_75t_L g1070 ( .A(n_1071), .Y(n_1070) );
AOI22x1_ASAP7_75t_L g1071 ( .A1(n_1072), .A2(n_1073), .B1(n_1096), .B2(n_1097), .Y(n_1071) );
INVx2_ASAP7_75t_L g1072 ( .A(n_1073), .Y(n_1072) );
AND2x2_ASAP7_75t_L g1073 ( .A(n_1074), .B(n_1084), .Y(n_1073) );
NOR2xp33_ASAP7_75t_L g1074 ( .A(n_1075), .B(n_1079), .Y(n_1074) );
NAND2xp5_ASAP7_75t_L g1079 ( .A(n_1080), .B(n_1083), .Y(n_1079) );
INVx1_ASAP7_75t_L g1081 ( .A(n_1082), .Y(n_1081) );
NOR2x1_ASAP7_75t_L g1084 ( .A(n_1085), .B(n_1091), .Y(n_1084) );
NAND2xp5_ASAP7_75t_L g1085 ( .A(n_1086), .B(n_1090), .Y(n_1085) );
INVx1_ASAP7_75t_L g1087 ( .A(n_1088), .Y(n_1087) );
INVx1_ASAP7_75t_L g1112 ( .A(n_1088), .Y(n_1112) );
NAND2xp5_ASAP7_75t_L g1091 ( .A(n_1092), .B(n_1095), .Y(n_1091) );
INVx2_ASAP7_75t_L g1093 ( .A(n_1094), .Y(n_1093) );
INVx1_ASAP7_75t_L g1096 ( .A(n_1097), .Y(n_1096) );
CKINVDCx6p67_ASAP7_75t_R g1098 ( .A(n_1099), .Y(n_1098) );
HB1xp67_ASAP7_75t_L g1101 ( .A(n_1102), .Y(n_1101) );
NAND4xp75_ASAP7_75t_L g1102 ( .A(n_1103), .B(n_1106), .C(n_1109), .D(n_1113), .Y(n_1102) );
AND2x2_ASAP7_75t_L g1103 ( .A(n_1104), .B(n_1105), .Y(n_1103) );
AND2x2_ASAP7_75t_L g1106 ( .A(n_1107), .B(n_1108), .Y(n_1106) );
AND2x2_ASAP7_75t_L g1109 ( .A(n_1110), .B(n_1111), .Y(n_1109) );
CKINVDCx20_ASAP7_75t_R g1115 ( .A(n_1116), .Y(n_1115) );
endmodule