module fake_ibex_683_n_3008 (n_151, n_85, n_507, n_540, n_395, n_84, n_64, n_171, n_103, n_529, n_389, n_204, n_274, n_387, n_130, n_177, n_76, n_273, n_309, n_330, n_9, n_328, n_293, n_341, n_372, n_124, n_37, n_256, n_418, n_193, n_510, n_446, n_108, n_350, n_165, n_452, n_86, n_70, n_255, n_175, n_398, n_59, n_28, n_125, n_304, n_191, n_5, n_62, n_71, n_153, n_545, n_194, n_249, n_334, n_312, n_478, n_239, n_94, n_134, n_432, n_371, n_403, n_423, n_357, n_88, n_412, n_457, n_494, n_142, n_226, n_336, n_258, n_40, n_90, n_17, n_74, n_449, n_547, n_176, n_58, n_43, n_216, n_33, n_421, n_475, n_166, n_163, n_500, n_542, n_114, n_236, n_34, n_376, n_377, n_531, n_15, n_556, n_24, n_189, n_498, n_280, n_317, n_340, n_375, n_105, n_187, n_1, n_154, n_182, n_196, n_326, n_327, n_89, n_50, n_144, n_170, n_270, n_346, n_383, n_113, n_117, n_417, n_471, n_265, n_504, n_158, n_259, n_276, n_339, n_470, n_210, n_348, n_220, n_91, n_481, n_287, n_54, n_243, n_19, n_497, n_228, n_147, n_552, n_251, n_384, n_373, n_458, n_244, n_73, n_343, n_310, n_426, n_323, n_469, n_143, n_106, n_386, n_549, n_8, n_224, n_183, n_533, n_508, n_67, n_453, n_333, n_110, n_306, n_400, n_47, n_550, n_169, n_10, n_21, n_242, n_278, n_316, n_16, n_404, n_60, n_557, n_7, n_109, n_127, n_121, n_527, n_465, n_48, n_325, n_57, n_301, n_496, n_434, n_296, n_120, n_168, n_526, n_155, n_315, n_441, n_13, n_122, n_523, n_116, n_370, n_431, n_0, n_289, n_12, n_515, n_150, n_286, n_321, n_133, n_51, n_215, n_279, n_49, n_374, n_235, n_464, n_538, n_22, n_136, n_261, n_521, n_459, n_30, n_518, n_367, n_221, n_437, n_355, n_474, n_407, n_102, n_490, n_52, n_448, n_99, n_466, n_269, n_156, n_126, n_530, n_356, n_25, n_104, n_45, n_420, n_483, n_543, n_141, n_487, n_222, n_186, n_524, n_349, n_454, n_295, n_331, n_230, n_96, n_185, n_388, n_536, n_352, n_290, n_174, n_467, n_427, n_157, n_219, n_246, n_31, n_442, n_146, n_207, n_438, n_167, n_128, n_253, n_208, n_234, n_3, n_152, n_300, n_145, n_65, n_358, n_205, n_488, n_139, n_514, n_429, n_275, n_541, n_98, n_129, n_267, n_245, n_229, n_209, n_472, n_347, n_473, n_445, n_335, n_413, n_82, n_263, n_27, n_353, n_359, n_299, n_87, n_262, n_433, n_75, n_439, n_137, n_338, n_173, n_477, n_363, n_402, n_180, n_369, n_201, n_14, n_351, n_368, n_456, n_257, n_77, n_44, n_401, n_553, n_554, n_66, n_305, n_307, n_192, n_140, n_484, n_480, n_416, n_365, n_4, n_6, n_539, n_100, n_179, n_354, n_206, n_392, n_516, n_548, n_329, n_447, n_26, n_188, n_200, n_444, n_506, n_546, n_199, n_495, n_410, n_308, n_463, n_411, n_135, n_520, n_512, n_283, n_366, n_397, n_111, n_36, n_18, n_322, n_53, n_227, n_499, n_115, n_11, n_248, n_92, n_451, n_101, n_190, n_138, n_409, n_214, n_238, n_332, n_517, n_211, n_218, n_314, n_132, n_277, n_555, n_337, n_522, n_479, n_534, n_225, n_360, n_272, n_511, n_23, n_468, n_223, n_381, n_525, n_535, n_382, n_502, n_532, n_95, n_405, n_415, n_285, n_288, n_247, n_320, n_379, n_551, n_55, n_291, n_318, n_63, n_161, n_237, n_29, n_203, n_268, n_440, n_148, n_2, n_342, n_233, n_385, n_414, n_430, n_118, n_378, n_486, n_422, n_164, n_38, n_198, n_264, n_217, n_324, n_391, n_537, n_78, n_20, n_69, n_390, n_544, n_39, n_178, n_509, n_303, n_362, n_93, n_505, n_162, n_482, n_240, n_282, n_61, n_501, n_266, n_42, n_294, n_112, n_485, n_46, n_284, n_80, n_172, n_250, n_493, n_460, n_476, n_461, n_313, n_519, n_345, n_408, n_119, n_361, n_455, n_419, n_72, n_319, n_195, n_513, n_212, n_311, n_406, n_97, n_197, n_528, n_181, n_131, n_123, n_260, n_462, n_302, n_450, n_443, n_344, n_393, n_436, n_428, n_491, n_297, n_435, n_41, n_252, n_396, n_83, n_32, n_107, n_149, n_489, n_399, n_254, n_213, n_424, n_271, n_241, n_68, n_503, n_292, n_394, n_79, n_81, n_35, n_364, n_159, n_202, n_231, n_298, n_160, n_184, n_56, n_492, n_232, n_380, n_281, n_425, n_3008);

input n_151;
input n_85;
input n_507;
input n_540;
input n_395;
input n_84;
input n_64;
input n_171;
input n_103;
input n_529;
input n_389;
input n_204;
input n_274;
input n_387;
input n_130;
input n_177;
input n_76;
input n_273;
input n_309;
input n_330;
input n_9;
input n_328;
input n_293;
input n_341;
input n_372;
input n_124;
input n_37;
input n_256;
input n_418;
input n_193;
input n_510;
input n_446;
input n_108;
input n_350;
input n_165;
input n_452;
input n_86;
input n_70;
input n_255;
input n_175;
input n_398;
input n_59;
input n_28;
input n_125;
input n_304;
input n_191;
input n_5;
input n_62;
input n_71;
input n_153;
input n_545;
input n_194;
input n_249;
input n_334;
input n_312;
input n_478;
input n_239;
input n_94;
input n_134;
input n_432;
input n_371;
input n_403;
input n_423;
input n_357;
input n_88;
input n_412;
input n_457;
input n_494;
input n_142;
input n_226;
input n_336;
input n_258;
input n_40;
input n_90;
input n_17;
input n_74;
input n_449;
input n_547;
input n_176;
input n_58;
input n_43;
input n_216;
input n_33;
input n_421;
input n_475;
input n_166;
input n_163;
input n_500;
input n_542;
input n_114;
input n_236;
input n_34;
input n_376;
input n_377;
input n_531;
input n_15;
input n_556;
input n_24;
input n_189;
input n_498;
input n_280;
input n_317;
input n_340;
input n_375;
input n_105;
input n_187;
input n_1;
input n_154;
input n_182;
input n_196;
input n_326;
input n_327;
input n_89;
input n_50;
input n_144;
input n_170;
input n_270;
input n_346;
input n_383;
input n_113;
input n_117;
input n_417;
input n_471;
input n_265;
input n_504;
input n_158;
input n_259;
input n_276;
input n_339;
input n_470;
input n_210;
input n_348;
input n_220;
input n_91;
input n_481;
input n_287;
input n_54;
input n_243;
input n_19;
input n_497;
input n_228;
input n_147;
input n_552;
input n_251;
input n_384;
input n_373;
input n_458;
input n_244;
input n_73;
input n_343;
input n_310;
input n_426;
input n_323;
input n_469;
input n_143;
input n_106;
input n_386;
input n_549;
input n_8;
input n_224;
input n_183;
input n_533;
input n_508;
input n_67;
input n_453;
input n_333;
input n_110;
input n_306;
input n_400;
input n_47;
input n_550;
input n_169;
input n_10;
input n_21;
input n_242;
input n_278;
input n_316;
input n_16;
input n_404;
input n_60;
input n_557;
input n_7;
input n_109;
input n_127;
input n_121;
input n_527;
input n_465;
input n_48;
input n_325;
input n_57;
input n_301;
input n_496;
input n_434;
input n_296;
input n_120;
input n_168;
input n_526;
input n_155;
input n_315;
input n_441;
input n_13;
input n_122;
input n_523;
input n_116;
input n_370;
input n_431;
input n_0;
input n_289;
input n_12;
input n_515;
input n_150;
input n_286;
input n_321;
input n_133;
input n_51;
input n_215;
input n_279;
input n_49;
input n_374;
input n_235;
input n_464;
input n_538;
input n_22;
input n_136;
input n_261;
input n_521;
input n_459;
input n_30;
input n_518;
input n_367;
input n_221;
input n_437;
input n_355;
input n_474;
input n_407;
input n_102;
input n_490;
input n_52;
input n_448;
input n_99;
input n_466;
input n_269;
input n_156;
input n_126;
input n_530;
input n_356;
input n_25;
input n_104;
input n_45;
input n_420;
input n_483;
input n_543;
input n_141;
input n_487;
input n_222;
input n_186;
input n_524;
input n_349;
input n_454;
input n_295;
input n_331;
input n_230;
input n_96;
input n_185;
input n_388;
input n_536;
input n_352;
input n_290;
input n_174;
input n_467;
input n_427;
input n_157;
input n_219;
input n_246;
input n_31;
input n_442;
input n_146;
input n_207;
input n_438;
input n_167;
input n_128;
input n_253;
input n_208;
input n_234;
input n_3;
input n_152;
input n_300;
input n_145;
input n_65;
input n_358;
input n_205;
input n_488;
input n_139;
input n_514;
input n_429;
input n_275;
input n_541;
input n_98;
input n_129;
input n_267;
input n_245;
input n_229;
input n_209;
input n_472;
input n_347;
input n_473;
input n_445;
input n_335;
input n_413;
input n_82;
input n_263;
input n_27;
input n_353;
input n_359;
input n_299;
input n_87;
input n_262;
input n_433;
input n_75;
input n_439;
input n_137;
input n_338;
input n_173;
input n_477;
input n_363;
input n_402;
input n_180;
input n_369;
input n_201;
input n_14;
input n_351;
input n_368;
input n_456;
input n_257;
input n_77;
input n_44;
input n_401;
input n_553;
input n_554;
input n_66;
input n_305;
input n_307;
input n_192;
input n_140;
input n_484;
input n_480;
input n_416;
input n_365;
input n_4;
input n_6;
input n_539;
input n_100;
input n_179;
input n_354;
input n_206;
input n_392;
input n_516;
input n_548;
input n_329;
input n_447;
input n_26;
input n_188;
input n_200;
input n_444;
input n_506;
input n_546;
input n_199;
input n_495;
input n_410;
input n_308;
input n_463;
input n_411;
input n_135;
input n_520;
input n_512;
input n_283;
input n_366;
input n_397;
input n_111;
input n_36;
input n_18;
input n_322;
input n_53;
input n_227;
input n_499;
input n_115;
input n_11;
input n_248;
input n_92;
input n_451;
input n_101;
input n_190;
input n_138;
input n_409;
input n_214;
input n_238;
input n_332;
input n_517;
input n_211;
input n_218;
input n_314;
input n_132;
input n_277;
input n_555;
input n_337;
input n_522;
input n_479;
input n_534;
input n_225;
input n_360;
input n_272;
input n_511;
input n_23;
input n_468;
input n_223;
input n_381;
input n_525;
input n_535;
input n_382;
input n_502;
input n_532;
input n_95;
input n_405;
input n_415;
input n_285;
input n_288;
input n_247;
input n_320;
input n_379;
input n_551;
input n_55;
input n_291;
input n_318;
input n_63;
input n_161;
input n_237;
input n_29;
input n_203;
input n_268;
input n_440;
input n_148;
input n_2;
input n_342;
input n_233;
input n_385;
input n_414;
input n_430;
input n_118;
input n_378;
input n_486;
input n_422;
input n_164;
input n_38;
input n_198;
input n_264;
input n_217;
input n_324;
input n_391;
input n_537;
input n_78;
input n_20;
input n_69;
input n_390;
input n_544;
input n_39;
input n_178;
input n_509;
input n_303;
input n_362;
input n_93;
input n_505;
input n_162;
input n_482;
input n_240;
input n_282;
input n_61;
input n_501;
input n_266;
input n_42;
input n_294;
input n_112;
input n_485;
input n_46;
input n_284;
input n_80;
input n_172;
input n_250;
input n_493;
input n_460;
input n_476;
input n_461;
input n_313;
input n_519;
input n_345;
input n_408;
input n_119;
input n_361;
input n_455;
input n_419;
input n_72;
input n_319;
input n_195;
input n_513;
input n_212;
input n_311;
input n_406;
input n_97;
input n_197;
input n_528;
input n_181;
input n_131;
input n_123;
input n_260;
input n_462;
input n_302;
input n_450;
input n_443;
input n_344;
input n_393;
input n_436;
input n_428;
input n_491;
input n_297;
input n_435;
input n_41;
input n_252;
input n_396;
input n_83;
input n_32;
input n_107;
input n_149;
input n_489;
input n_399;
input n_254;
input n_213;
input n_424;
input n_271;
input n_241;
input n_68;
input n_503;
input n_292;
input n_394;
input n_79;
input n_81;
input n_35;
input n_364;
input n_159;
input n_202;
input n_231;
input n_298;
input n_160;
input n_184;
input n_56;
input n_492;
input n_232;
input n_380;
input n_281;
input n_425;

output n_3008;

wire n_1084;
wire n_2594;
wire n_1474;
wire n_1295;
wire n_1983;
wire n_2804;
wire n_992;
wire n_1582;
wire n_2201;
wire n_2512;
wire n_766;
wire n_2960;
wire n_2175;
wire n_2071;
wire n_2796;
wire n_1110;
wire n_2607;
wire n_1382;
wire n_2569;
wire n_2949;
wire n_1998;
wire n_2840;
wire n_1596;
wire n_926;
wire n_1079;
wire n_2835;
wire n_1100;
wire n_845;
wire n_2177;
wire n_1930;
wire n_2123;
wire n_1234;
wire n_2047;
wire n_1594;
wire n_1944;
wire n_2235;
wire n_1802;
wire n_2498;
wire n_773;
wire n_2038;
wire n_2504;
wire n_1469;
wire n_821;
wire n_2017;
wire n_1227;
wire n_873;
wire n_962;
wire n_1080;
wire n_909;
wire n_862;
wire n_2290;
wire n_957;
wire n_1652;
wire n_969;
wire n_678;
wire n_1859;
wire n_1954;
wire n_2183;
wire n_2074;
wire n_2897;
wire n_1883;
wire n_1125;
wire n_733;
wire n_2687;
wire n_2037;
wire n_622;
wire n_1226;
wire n_1034;
wire n_2383;
wire n_1765;
wire n_872;
wire n_2392;
wire n_1873;
wire n_1619;
wire n_1666;
wire n_2640;
wire n_2682;
wire n_930;
wire n_1044;
wire n_1492;
wire n_1134;
wire n_1478;
wire n_1684;
wire n_1796;
wire n_1614;
wire n_2374;
wire n_2598;
wire n_1722;
wire n_911;
wire n_2023;
wire n_652;
wire n_781;
wire n_2720;
wire n_802;
wire n_2335;
wire n_1233;
wire n_2322;
wire n_2955;
wire n_2276;
wire n_1045;
wire n_2989;
wire n_1856;
wire n_963;
wire n_1782;
wire n_2230;
wire n_2889;
wire n_2139;
wire n_2847;
wire n_1308;
wire n_1138;
wire n_2943;
wire n_708;
wire n_1096;
wire n_2151;
wire n_2391;
wire n_1391;
wire n_667;
wire n_884;
wire n_2396;
wire n_850;
wire n_1971;
wire n_2485;
wire n_2479;
wire n_879;
wire n_2179;
wire n_1957;
wire n_2188;
wire n_723;
wire n_1144;
wire n_2359;
wire n_2360;
wire n_2506;
wire n_1392;
wire n_2158;
wire n_1268;
wire n_2571;
wire n_739;
wire n_2724;
wire n_2475;
wire n_853;
wire n_948;
wire n_2799;
wire n_1752;
wire n_1829;
wire n_1338;
wire n_1730;
wire n_875;
wire n_1307;
wire n_1327;
wire n_2644;
wire n_876;
wire n_711;
wire n_1840;
wire n_2837;
wire n_671;
wire n_989;
wire n_1908;
wire n_1668;
wire n_2343;
wire n_2605;
wire n_2887;
wire n_1641;
wire n_829;
wire n_2565;
wire n_825;
wire n_1480;
wire n_1463;
wire n_1823;
wire n_1681;
wire n_2921;
wire n_939;
wire n_1636;
wire n_1687;
wire n_655;
wire n_2192;
wire n_1766;
wire n_1922;
wire n_2032;
wire n_2820;
wire n_641;
wire n_1937;
wire n_2311;
wire n_893;
wire n_1654;
wire n_2995;
wire n_1258;
wire n_1344;
wire n_2208;
wire n_2198;
wire n_1929;
wire n_2707;
wire n_1749;
wire n_1680;
wire n_835;
wire n_1981;
wire n_1195;
wire n_2918;
wire n_824;
wire n_1945;
wire n_2638;
wire n_694;
wire n_787;
wire n_2860;
wire n_2448;
wire n_614;
wire n_2015;
wire n_2537;
wire n_1130;
wire n_2643;
wire n_1228;
wire n_2998;
wire n_2336;
wire n_2163;
wire n_1081;
wire n_2354;
wire n_1155;
wire n_1292;
wire n_2432;
wire n_2873;
wire n_1576;
wire n_1664;
wire n_2273;
wire n_852;
wire n_1427;
wire n_1133;
wire n_2421;
wire n_1926;
wire n_904;
wire n_2363;
wire n_2814;
wire n_2003;
wire n_1970;
wire n_2621;
wire n_1778;
wire n_646;
wire n_2558;
wire n_2953;
wire n_2922;
wire n_2347;
wire n_2839;
wire n_1030;
wire n_1698;
wire n_1094;
wire n_2462;
wire n_1496;
wire n_2333;
wire n_715;
wire n_1910;
wire n_1663;
wire n_2436;
wire n_1214;
wire n_1274;
wire n_2705;
wire n_2527;
wire n_1606;
wire n_769;
wire n_1595;
wire n_2164;
wire n_1509;
wire n_1618;
wire n_1648;
wire n_2944;
wire n_1886;
wire n_2269;
wire n_857;
wire n_765;
wire n_1070;
wire n_1841;
wire n_2472;
wire n_777;
wire n_2685;
wire n_2846;
wire n_1955;
wire n_917;
wire n_2249;
wire n_2413;
wire n_2362;
wire n_968;
wire n_2822;
wire n_1253;
wire n_1306;
wire n_1484;
wire n_2686;
wire n_1493;
wire n_2597;
wire n_1313;
wire n_2774;
wire n_558;
wire n_2090;
wire n_666;
wire n_2260;
wire n_2812;
wire n_2753;
wire n_1638;
wire n_2215;
wire n_1071;
wire n_1449;
wire n_1723;
wire n_1960;
wire n_2663;
wire n_793;
wire n_937;
wire n_2595;
wire n_2116;
wire n_1645;
wire n_973;
wire n_1038;
wire n_2280;
wire n_618;
wire n_1943;
wire n_1863;
wire n_2844;
wire n_1269;
wire n_2393;
wire n_2773;
wire n_662;
wire n_2906;
wire n_979;
wire n_1309;
wire n_1999;
wire n_1316;
wire n_1562;
wire n_1215;
wire n_629;
wire n_2777;
wire n_2480;
wire n_1445;
wire n_573;
wire n_2283;
wire n_2806;
wire n_2813;
wire n_2147;
wire n_1716;
wire n_1466;
wire n_1412;
wire n_1672;
wire n_1007;
wire n_2253;
wire n_643;
wire n_1276;
wire n_1637;
wire n_841;
wire n_2900;
wire n_772;
wire n_810;
wire n_1401;
wire n_1817;
wire n_2951;
wire n_2145;
wire n_2122;
wire n_1588;
wire n_2216;
wire n_1301;
wire n_2579;
wire n_2876;
wire n_2242;
wire n_869;
wire n_1620;
wire n_1561;
wire n_718;
wire n_2370;
wire n_2025;
wire n_1078;
wire n_2247;
wire n_1219;
wire n_713;
wire n_1865;
wire n_1252;
wire n_2022;
wire n_2730;
wire n_1170;
wire n_1927;
wire n_605;
wire n_2373;
wire n_630;
wire n_1869;
wire n_567;
wire n_2275;
wire n_1853;
wire n_2980;
wire n_2189;
wire n_2482;
wire n_745;
wire n_2767;
wire n_2826;
wire n_2899;
wire n_2112;
wire n_1753;
wire n_564;
wire n_562;
wire n_1322;
wire n_2008;
wire n_1305;
wire n_2088;
wire n_795;
wire n_592;
wire n_1248;
wire n_2762;
wire n_2171;
wire n_762;
wire n_1388;
wire n_2859;
wire n_800;
wire n_2564;
wire n_706;
wire n_784;
wire n_684;
wire n_1653;
wire n_1375;
wire n_1356;
wire n_894;
wire n_1118;
wire n_692;
wire n_2591;
wire n_1881;
wire n_1969;
wire n_709;
wire n_1296;
wire n_971;
wire n_1326;
wire n_702;
wire n_1350;
wire n_906;
wire n_2957;
wire n_2586;
wire n_1093;
wire n_1764;
wire n_2412;
wire n_2783;
wire n_978;
wire n_899;
wire n_579;
wire n_1799;
wire n_1019;
wire n_902;
wire n_1689;
wire n_1250;
wire n_2550;
wire n_1190;
wire n_1304;
wire n_744;
wire n_563;
wire n_2541;
wire n_1506;
wire n_881;
wire n_2987;
wire n_1702;
wire n_734;
wire n_1558;
wire n_2750;
wire n_1650;
wire n_1520;
wire n_1073;
wire n_1453;
wire n_1108;
wire n_2722;
wire n_2509;
wire n_2727;
wire n_1794;
wire n_1423;
wire n_1239;
wire n_2399;
wire n_1370;
wire n_2719;
wire n_1209;
wire n_1708;
wire n_2213;
wire n_2723;
wire n_1616;
wire n_729;
wire n_1569;
wire n_2664;
wire n_1434;
wire n_603;
wire n_1649;
wire n_2389;
wire n_1936;
wire n_2114;
wire n_1717;
wire n_2107;
wire n_1609;
wire n_2257;
wire n_1613;
wire n_820;
wire n_805;
wire n_1988;
wire n_670;
wire n_1132;
wire n_892;
wire n_1467;
wire n_1803;
wire n_2401;
wire n_1787;
wire n_2782;
wire n_2511;
wire n_1281;
wire n_1447;
wire n_2166;
wire n_2451;
wire n_2150;
wire n_695;
wire n_1549;
wire n_639;
wire n_2631;
wire n_1867;
wire n_1531;
wire n_2919;
wire n_1332;
wire n_2660;
wire n_2661;
wire n_2292;
wire n_2334;
wire n_1424;
wire n_2444;
wire n_2350;
wire n_1742;
wire n_2625;
wire n_1818;
wire n_870;
wire n_2199;
wire n_1709;
wire n_1610;
wire n_2219;
wire n_1298;
wire n_1844;
wire n_1387;
wire n_2649;
wire n_609;
wire n_1040;
wire n_2203;
wire n_2693;
wire n_1159;
wire n_1368;
wire n_2281;
wire n_1154;
wire n_2539;
wire n_2431;
wire n_1701;
wire n_2084;
wire n_1243;
wire n_2387;
wire n_2646;
wire n_2397;
wire n_1121;
wire n_693;
wire n_2746;
wire n_2256;
wire n_606;
wire n_737;
wire n_2445;
wire n_2729;
wire n_1571;
wire n_1980;
wire n_2529;
wire n_2019;
wire n_1407;
wire n_1235;
wire n_1821;
wire n_1003;
wire n_889;
wire n_2708;
wire n_2748;
wire n_816;
wire n_1058;
wire n_1835;
wire n_1862;
wire n_2224;
wire n_2697;
wire n_2470;
wire n_2355;
wire n_2890;
wire n_2731;
wire n_1543;
wire n_823;
wire n_2233;
wire n_2499;
wire n_1504;
wire n_1519;
wire n_1425;
wire n_1781;
wire n_2069;
wire n_2602;
wire n_1441;
wire n_2028;
wire n_1924;
wire n_2856;
wire n_1921;
wire n_657;
wire n_1156;
wire n_2857;
wire n_1293;
wire n_1360;
wire n_749;
wire n_1555;
wire n_1394;
wire n_1347;
wire n_819;
wire n_2070;
wire n_1042;
wire n_822;
wire n_1888;
wire n_743;
wire n_754;
wire n_1786;
wire n_2033;
wire n_1319;
wire n_1553;
wire n_1041;
wire n_2766;
wire n_2828;
wire n_1964;
wire n_1090;
wire n_1196;
wire n_1182;
wire n_1271;
wire n_2416;
wire n_2786;
wire n_1731;
wire n_1905;
wire n_2962;
wire n_1031;
wire n_2879;
wire n_2958;
wire n_2052;
wire n_981;
wire n_2425;
wire n_2800;
wire n_3006;
wire n_2118;
wire n_2259;
wire n_2162;
wire n_2236;
wire n_2377;
wire n_2718;
wire n_2577;
wire n_1591;
wire n_583;
wire n_2289;
wire n_2288;
wire n_2841;
wire n_1671;
wire n_1795;
wire n_1409;
wire n_1015;
wire n_663;
wire n_2744;
wire n_2101;
wire n_2795;
wire n_1377;
wire n_2473;
wire n_1583;
wire n_1521;
wire n_2632;
wire n_1152;
wire n_2456;
wire n_2924;
wire n_2264;
wire n_2076;
wire n_1036;
wire n_974;
wire n_2599;
wire n_1831;
wire n_608;
wire n_864;
wire n_1987;
wire n_959;
wire n_1106;
wire n_1312;
wire n_1129;
wire n_1244;
wire n_1733;
wire n_1634;
wire n_2853;
wire n_1932;
wire n_1452;
wire n_1552;
wire n_1318;
wire n_1508;
wire n_2217;
wire n_738;
wire n_1217;
wire n_2866;
wire n_2655;
wire n_2454;
wire n_1715;
wire n_1189;
wire n_761;
wire n_748;
wire n_1713;
wire n_901;
wire n_1577;
wire n_2036;
wire n_1255;
wire n_2829;
wire n_2968;
wire n_2740;
wire n_1700;
wire n_2623;
wire n_2622;
wire n_2819;
wire n_1218;
wire n_2178;
wire n_1181;
wire n_1140;
wire n_1985;
wire n_1772;
wire n_2858;
wire n_1056;
wire n_2626;
wire n_1283;
wire n_3007;
wire n_1446;
wire n_2404;
wire n_1487;
wire n_2789;
wire n_2603;
wire n_840;
wire n_1203;
wire n_1421;
wire n_561;
wire n_2821;
wire n_2424;
wire n_846;
wire n_1793;
wire n_1237;
wire n_2573;
wire n_2390;
wire n_2880;
wire n_2423;
wire n_859;
wire n_965;
wire n_1109;
wire n_2741;
wire n_2793;
wire n_1633;
wire n_2580;
wire n_1711;
wire n_1051;
wire n_1008;
wire n_2964;
wire n_2375;
wire n_1498;
wire n_2312;
wire n_2572;
wire n_2946;
wire n_1053;
wire n_1656;
wire n_1207;
wire n_1076;
wire n_1735;
wire n_2063;
wire n_1032;
wire n_936;
wire n_1884;
wire n_2176;
wire n_1825;
wire n_2805;
wire n_1589;
wire n_2717;
wire n_2204;
wire n_2863;
wire n_2575;
wire n_1210;
wire n_2319;
wire n_591;
wire n_2877;
wire n_1933;
wire n_2522;
wire n_1996;
wire n_1510;
wire n_1201;
wire n_1842;
wire n_2852;
wire n_2132;
wire n_1246;
wire n_1677;
wire n_732;
wire n_1236;
wire n_832;
wire n_2297;
wire n_2780;
wire n_1792;
wire n_1712;
wire n_1984;
wire n_590;
wire n_1568;
wire n_2885;
wire n_1877;
wire n_1184;
wire n_1477;
wire n_2080;
wire n_2220;
wire n_2585;
wire n_1724;
wire n_2554;
wire n_2838;
wire n_1364;
wire n_1540;
wire n_1676;
wire n_1013;
wire n_2468;
wire n_929;
wire n_637;
wire n_1136;
wire n_1890;
wire n_1075;
wire n_1249;
wire n_1918;
wire n_574;
wire n_2606;
wire n_2549;
wire n_2461;
wire n_2006;
wire n_2440;
wire n_1229;
wire n_1440;
wire n_1490;
wire n_2152;
wire n_907;
wire n_1179;
wire n_1990;
wire n_1153;
wire n_1751;
wire n_669;
wire n_2787;
wire n_2467;
wire n_2146;
wire n_2341;
wire n_1737;
wire n_2779;
wire n_1117;
wire n_1273;
wire n_2547;
wire n_2930;
wire n_2616;
wire n_1748;
wire n_2662;
wire n_1083;
wire n_1014;
wire n_724;
wire n_2883;
wire n_938;
wire n_1178;
wire n_2935;
wire n_878;
wire n_2441;
wire n_2358;
wire n_2490;
wire n_594;
wire n_2361;
wire n_1464;
wire n_1566;
wire n_944;
wire n_3003;
wire n_1848;
wire n_623;
wire n_2062;
wire n_2277;
wire n_585;
wire n_2650;
wire n_1982;
wire n_2252;
wire n_2888;
wire n_2339;
wire n_1334;
wire n_1963;
wire n_1695;
wire n_1418;
wire n_2999;
wire n_2402;
wire n_1137;
wire n_2552;
wire n_2910;
wire n_660;
wire n_2590;
wire n_1977;
wire n_2294;
wire n_1200;
wire n_2295;
wire n_2530;
wire n_2379;
wire n_1120;
wire n_2300;
wire n_2792;
wire n_576;
wire n_1602;
wire n_2965;
wire n_1776;
wire n_2372;
wire n_2382;
wire n_1852;
wire n_1522;
wire n_2523;
wire n_2557;
wire n_1279;
wire n_2505;
wire n_931;
wire n_607;
wire n_827;
wire n_2481;
wire n_1064;
wire n_1408;
wire n_2832;
wire n_1028;
wire n_1264;
wire n_2808;
wire n_2287;
wire n_2954;
wire n_2102;
wire n_1935;
wire n_2046;
wire n_1146;
wire n_2785;
wire n_2751;
wire n_705;
wire n_2142;
wire n_1548;
wire n_2977;
wire n_1682;
wire n_1608;
wire n_1009;
wire n_1260;
wire n_589;
wire n_1896;
wire n_1704;
wire n_2160;
wire n_2699;
wire n_2234;
wire n_847;
wire n_2991;
wire n_1436;
wire n_2600;
wire n_1069;
wire n_1485;
wire n_2239;
wire n_1465;
wire n_1352;
wire n_1171;
wire n_1126;
wire n_1232;
wire n_1979;
wire n_2328;
wire n_2715;
wire n_679;
wire n_1345;
wire n_2434;
wire n_696;
wire n_837;
wire n_1590;
wire n_2332;
wire n_640;
wire n_2971;
wire n_954;
wire n_1628;
wire n_725;
wire n_1773;
wire n_596;
wire n_2133;
wire n_1545;
wire n_2369;
wire n_1471;
wire n_1738;
wire n_998;
wire n_1115;
wire n_1395;
wire n_1729;
wire n_2551;
wire n_801;
wire n_2823;
wire n_2094;
wire n_2613;
wire n_1479;
wire n_2306;
wire n_1046;
wire n_2419;
wire n_2934;
wire n_2807;
wire n_882;
wire n_942;
wire n_1627;
wire n_1431;
wire n_651;
wire n_721;
wire n_2525;
wire n_814;
wire n_1864;
wire n_943;
wire n_2568;
wire n_2629;
wire n_1086;
wire n_1523;
wire n_2197;
wire n_1756;
wire n_2010;
wire n_2097;
wire n_2733;
wire n_2241;
wire n_1470;
wire n_2098;
wire n_2109;
wire n_1761;
wire n_2648;
wire n_2458;
wire n_1836;
wire n_2398;
wire n_1593;
wire n_986;
wire n_1420;
wire n_2651;
wire n_1750;
wire n_1775;
wire n_2833;
wire n_1699;
wire n_927;
wire n_1563;
wire n_615;
wire n_2905;
wire n_803;
wire n_2570;
wire n_1875;
wire n_1615;
wire n_2184;
wire n_2418;
wire n_1087;
wire n_757;
wire n_1539;
wire n_712;
wire n_1400;
wire n_1599;
wire n_1806;
wire n_2711;
wire n_2842;
wire n_650;
wire n_2635;
wire n_2469;
wire n_1575;
wire n_2209;
wire n_1448;
wire n_2077;
wire n_2520;
wire n_817;
wire n_2193;
wire n_2612;
wire n_2095;
wire n_2486;
wire n_2628;
wire n_2395;
wire n_951;
wire n_2521;
wire n_2908;
wire n_2053;
wire n_2752;
wire n_1580;
wire n_2124;
wire n_1574;
wire n_780;
wire n_2200;
wire n_1705;
wire n_633;
wire n_2304;
wire n_1746;
wire n_726;
wire n_1439;
wire n_2263;
wire n_2212;
wire n_2352;
wire n_2716;
wire n_863;
wire n_597;
wire n_2185;
wire n_1832;
wire n_1128;
wire n_2476;
wire n_2376;
wire n_2979;
wire n_1266;
wire n_1300;
wire n_2781;
wire n_807;
wire n_741;
wire n_2460;
wire n_2170;
wire n_1785;
wire n_1870;
wire n_2484;
wire n_2721;
wire n_1405;
wire n_2884;
wire n_997;
wire n_2308;
wire n_2986;
wire n_1428;
wire n_2691;
wire n_2243;
wire n_2400;
wire n_2903;
wire n_891;
wire n_2507;
wire n_2759;
wire n_1528;
wire n_1495;
wire n_2463;
wire n_2654;
wire n_717;
wire n_2975;
wire n_1357;
wire n_2503;
wire n_2478;
wire n_2794;
wire n_1512;
wire n_2496;
wire n_668;
wire n_2974;
wire n_871;
wire n_2990;
wire n_2923;
wire n_1339;
wire n_1544;
wire n_1426;
wire n_2365;
wire n_2245;
wire n_1315;
wire n_1413;
wire n_2464;
wire n_811;
wire n_808;
wire n_945;
wire n_2925;
wire n_2270;
wire n_1706;
wire n_1560;
wire n_1592;
wire n_2776;
wire n_1461;
wire n_2695;
wire n_2630;
wire n_903;
wire n_1967;
wire n_2340;
wire n_2117;
wire n_1095;
wire n_1328;
wire n_1265;
wire n_2488;
wire n_1378;
wire n_2042;
wire n_1048;
wire n_774;
wire n_2459;
wire n_1925;
wire n_2439;
wire n_2106;
wire n_588;
wire n_1430;
wire n_2414;
wire n_1251;
wire n_1247;
wire n_2450;
wire n_836;
wire n_1475;
wire n_2465;
wire n_1263;
wire n_1185;
wire n_1683;
wire n_1122;
wire n_2765;
wire n_890;
wire n_628;
wire n_874;
wire n_1505;
wire n_2941;
wire n_1163;
wire n_677;
wire n_1514;
wire n_964;
wire n_2728;
wire n_2948;
wire n_916;
wire n_2298;
wire n_2771;
wire n_2936;
wire n_895;
wire n_687;
wire n_1035;
wire n_2427;
wire n_2045;
wire n_2985;
wire n_1535;
wire n_751;
wire n_2190;
wire n_1127;
wire n_932;
wire n_1972;
wire n_2772;
wire n_2778;
wire n_947;
wire n_1004;
wire n_831;
wire n_778;
wire n_1898;
wire n_1254;
wire n_1148;
wire n_1667;
wire n_1104;
wire n_1845;
wire n_1011;
wire n_2205;
wire n_2684;
wire n_2875;
wire n_2524;
wire n_1437;
wire n_2747;
wire n_626;
wire n_1707;
wire n_1941;
wire n_2422;
wire n_2064;
wire n_1679;
wire n_2342;
wire n_2755;
wire n_2301;
wire n_1497;
wire n_2002;
wire n_2055;
wire n_2385;
wire n_2545;
wire n_1578;
wire n_2050;
wire n_1143;
wire n_1783;
wire n_2712;
wire n_2584;
wire n_972;
wire n_1815;
wire n_2500;
wire n_601;
wire n_610;
wire n_1917;
wire n_1444;
wire n_920;
wire n_664;
wire n_2442;
wire n_1067;
wire n_2763;
wire n_2788;
wire n_994;
wire n_2000;
wire n_2089;
wire n_1857;
wire n_2761;
wire n_1920;
wire n_2696;
wire n_887;
wire n_1162;
wire n_1997;
wire n_2578;
wire n_2745;
wire n_1894;
wire n_2110;
wire n_2904;
wire n_2896;
wire n_2997;
wire n_634;
wire n_991;
wire n_961;
wire n_1223;
wire n_1349;
wire n_1331;
wire n_2127;
wire n_1323;
wire n_578;
wire n_1739;
wire n_1777;
wire n_1353;
wire n_2386;
wire n_1429;
wire n_2029;
wire n_2026;
wire n_1546;
wire n_1432;
wire n_2103;
wire n_1950;
wire n_1320;
wire n_996;
wire n_915;
wire n_2238;
wire n_2619;
wire n_1174;
wire n_1874;
wire n_1834;
wire n_2862;
wire n_1727;
wire n_1286;
wire n_1657;
wire n_1741;
wire n_1294;
wire n_1601;
wire n_900;
wire n_1351;
wire n_2933;
wire n_2138;
wire n_647;
wire n_1380;
wire n_1367;
wire n_1291;
wire n_2895;
wire n_1914;
wire n_1458;
wire n_1694;
wire n_1460;
wire n_2041;
wire n_2271;
wire n_2356;
wire n_1830;
wire n_2261;
wire n_1629;
wire n_2994;
wire n_2011;
wire n_2620;
wire n_1826;
wire n_1855;
wire n_1662;
wire n_2187;
wire n_2105;
wire n_1340;
wire n_2694;
wire n_2562;
wire n_2642;
wire n_2647;
wire n_1626;
wire n_674;
wire n_2223;
wire n_1660;
wire n_1850;
wire n_1643;
wire n_1670;
wire n_1789;
wire n_2415;
wire n_2344;
wire n_2317;
wire n_2556;
wire n_1112;
wire n_1267;
wire n_2384;
wire n_2683;
wire n_1384;
wire n_1376;
wire n_1537;
wire n_1858;
wire n_2815;
wire n_1816;
wire n_2446;
wire n_1612;
wire n_703;
wire n_2318;
wire n_1172;
wire n_2659;
wire n_1099;
wire n_598;
wire n_2141;
wire n_2902;
wire n_2909;
wire n_1422;
wire n_1527;
wire n_1055;
wire n_1524;
wire n_673;
wire n_798;
wire n_2849;
wire n_2947;
wire n_1754;
wire n_1177;
wire n_1025;
wire n_1991;
wire n_2566;
wire n_2679;
wire n_2210;
wire n_1517;
wire n_690;
wire n_2502;
wire n_1225;
wire n_1962;
wire n_2346;
wire n_982;
wire n_1624;
wire n_785;
wire n_1952;
wire n_2180;
wire n_3002;
wire n_2087;
wire n_2920;
wire n_604;
wire n_1598;
wire n_2952;
wire n_2617;
wire n_977;
wire n_2878;
wire n_1895;
wire n_2250;
wire n_719;
wire n_1491;
wire n_1860;
wire n_2831;
wire n_716;
wire n_1810;
wire n_1763;
wire n_923;
wire n_642;
wire n_1607;
wire n_2865;
wire n_2075;
wire n_2959;
wire n_1625;
wire n_2610;
wire n_2420;
wire n_2380;
wire n_2240;
wire n_933;
wire n_2221;
wire n_1774;
wire n_1797;
wire n_2516;
wire n_2120;
wire n_1037;
wire n_1899;
wire n_2031;
wire n_1348;
wire n_838;
wire n_1289;
wire n_2892;
wire n_1021;
wire n_746;
wire n_1557;
wire n_1188;
wire n_1567;
wire n_2007;
wire n_742;
wire n_1191;
wire n_2004;
wire n_2024;
wire n_2086;
wire n_1503;
wire n_1052;
wire n_789;
wire n_1942;
wire n_656;
wire n_602;
wire n_2309;
wire n_842;
wire n_2274;
wire n_2698;
wire n_767;
wire n_1617;
wire n_1839;
wire n_1587;
wire n_2330;
wire n_2639;
wire n_2555;
wire n_636;
wire n_1259;
wire n_2108;
wire n_2535;
wire n_595;
wire n_1001;
wire n_2945;
wire n_570;
wire n_2143;
wire n_2410;
wire n_1396;
wire n_2916;
wire n_1224;
wire n_1923;
wire n_2196;
wire n_2739;
wire n_2611;
wire n_1538;
wire n_2528;
wire n_2548;
wire n_2709;
wire n_2633;
wire n_1017;
wire n_2244;
wire n_730;
wire n_2604;
wire n_2351;
wire n_2437;
wire n_2049;
wire n_1456;
wire n_1889;
wire n_625;
wire n_2113;
wire n_619;
wire n_2665;
wire n_1124;
wire n_611;
wire n_1690;
wire n_2688;
wire n_2881;
wire n_1673;
wire n_2018;
wire n_922;
wire n_2817;
wire n_1790;
wire n_993;
wire n_851;
wire n_2085;
wire n_2581;
wire n_1725;
wire n_2809;
wire n_2149;
wire n_2237;
wire n_2320;
wire n_2268;
wire n_1135;
wire n_2255;
wire n_2001;
wire n_1820;
wire n_1800;
wire n_2758;
wire n_613;
wire n_659;
wire n_1494;
wire n_1550;
wire n_2060;
wire n_1066;
wire n_2214;
wire n_1169;
wire n_648;
wire n_571;
wire n_1726;
wire n_1946;
wire n_1938;
wire n_830;
wire n_1241;
wire n_2589;
wire n_1072;
wire n_2194;
wire n_1231;
wire n_1173;
wire n_2736;
wire n_1208;
wire n_1604;
wire n_1639;
wire n_2735;
wire n_2845;
wire n_826;
wire n_1976;
wire n_2154;
wire n_2035;
wire n_1337;
wire n_2732;
wire n_2984;
wire n_1906;
wire n_3004;
wire n_1647;
wire n_1901;
wire n_839;
wire n_768;
wire n_1278;
wire n_2059;
wire n_796;
wire n_797;
wire n_1006;
wire n_2956;
wire n_1238;
wire n_1415;
wire n_976;
wire n_1710;
wire n_1063;
wire n_2153;
wire n_2452;
wire n_1270;
wire n_2891;
wire n_834;
wire n_2457;
wire n_2144;
wire n_1476;
wire n_935;
wire n_1603;
wire n_925;
wire n_2592;
wire n_1054;
wire n_2027;
wire n_2072;
wire n_2737;
wire n_2012;
wire n_722;
wire n_2251;
wire n_2963;
wire n_1644;
wire n_1406;
wire n_1489;
wire n_1880;
wire n_1993;
wire n_2137;
wire n_804;
wire n_1455;
wire n_1642;
wire n_1871;
wire n_2182;
wire n_2868;
wire n_2447;
wire n_2818;
wire n_1057;
wire n_1473;
wire n_2125;
wire n_2426;
wire n_2894;
wire n_1403;
wire n_2181;
wire n_2587;
wire n_1149;
wire n_1176;
wire n_1502;
wire n_1605;
wire n_868;
wire n_2099;
wire n_1202;
wire n_1065;
wire n_1897;
wire n_2477;
wire n_1457;
wire n_905;
wire n_2159;
wire n_975;
wire n_675;
wire n_624;
wire n_934;
wire n_775;
wire n_950;
wire n_2700;
wire n_685;
wire n_1222;
wire n_1630;
wire n_2286;
wire n_1879;
wire n_1959;
wire n_2563;
wire n_1198;
wire n_2206;
wire n_1311;
wire n_1261;
wire n_2299;
wire n_2078;
wire n_2265;
wire n_776;
wire n_1114;
wire n_1167;
wire n_818;
wire n_2677;
wire n_2531;
wire n_2315;
wire n_2157;
wire n_1282;
wire n_2067;
wire n_2517;
wire n_1321;
wire n_700;
wire n_1779;
wire n_2489;
wire n_1770;
wire n_1107;
wire n_1846;
wire n_2211;
wire n_1573;
wire n_2950;
wire n_815;
wire n_919;
wire n_2272;
wire n_1956;
wire n_681;
wire n_2608;
wire n_2983;
wire n_1718;
wire n_2225;
wire n_2546;
wire n_1411;
wire n_2825;
wire n_1139;
wire n_858;
wire n_1018;
wire n_2345;
wire n_1324;
wire n_1669;
wire n_1501;
wire n_2742;
wire n_782;
wire n_616;
wire n_1885;
wire n_1740;
wire n_1989;
wire n_1838;
wire n_833;
wire n_2680;
wire n_1343;
wire n_1801;
wire n_1371;
wire n_1513;
wire n_728;
wire n_3001;
wire n_2861;
wire n_2976;
wire n_2161;
wire n_2191;
wire n_2329;
wire n_1788;
wire n_2093;
wire n_2348;
wire n_786;
wire n_2675;
wire n_2417;
wire n_2576;
wire n_2043;
wire n_2366;
wire n_1621;
wire n_2338;
wire n_1919;
wire n_1342;
wire n_752;
wire n_2756;
wire n_2893;
wire n_2009;
wire n_2248;
wire n_958;
wire n_1175;
wire n_1416;
wire n_1659;
wire n_2850;
wire n_1221;
wire n_1047;
wire n_1878;
wire n_1515;
wire n_1374;
wire n_2851;
wire n_2438;
wire n_1435;
wire n_1688;
wire n_792;
wire n_2973;
wire n_1314;
wire n_1433;
wire n_2567;
wire n_575;
wire n_1242;
wire n_1119;
wire n_2229;
wire n_2810;
wire n_2867;
wire n_1085;
wire n_2388;
wire n_2981;
wire n_2222;
wire n_1907;
wire n_885;
wire n_1530;
wire n_877;
wire n_2871;
wire n_2135;
wire n_1088;
wire n_896;
wire n_2764;
wire n_2624;
wire n_1813;
wire n_1451;
wire n_1005;
wire n_1102;
wire n_631;
wire n_794;
wire n_2471;
wire n_1288;
wire n_1275;
wire n_985;
wire n_1165;
wire n_897;
wire n_1622;
wire n_2757;
wire n_2714;
wire n_2669;
wire n_697;
wire n_2869;
wire n_1105;
wire n_1459;
wire n_912;
wire n_2898;
wire n_2232;
wire n_2455;
wire n_2121;
wire n_1893;
wire n_2519;
wire n_1570;
wire n_2231;
wire n_2874;
wire n_701;
wire n_995;
wire n_2278;
wire n_1000;
wire n_2284;
wire n_1931;
wire n_2433;
wire n_2803;
wire n_2816;
wire n_1256;
wire n_2798;
wire n_587;
wire n_1303;
wire n_1994;
wire n_1771;
wire n_1526;
wire n_764;
wire n_1507;
wire n_1206;
wire n_1809;
wire n_855;
wire n_2367;
wire n_812;
wire n_2658;
wire n_1961;
wire n_2553;
wire n_1050;
wire n_2218;
wire n_2667;
wire n_599;
wire n_1769;
wire n_2130;
wire n_1060;
wire n_1372;
wire n_1847;
wire n_756;
wire n_1565;
wire n_1257;
wire n_2325;
wire n_2864;
wire n_1632;
wire n_2406;
wire n_688;
wire n_1542;
wire n_946;
wire n_1586;
wire n_707;
wire n_1362;
wire n_1547;
wire n_1097;
wire n_2518;
wire n_2784;
wire n_1909;
wire n_2543;
wire n_2381;
wire n_621;
wire n_2313;
wire n_956;
wire n_790;
wire n_2495;
wire n_2992;
wire n_1541;
wire n_2703;
wire n_1812;
wire n_1951;
wire n_586;
wire n_1330;
wire n_638;
wire n_1697;
wire n_2128;
wire n_2574;
wire n_1872;
wire n_1940;
wire n_2690;
wire n_593;
wire n_1747;
wire n_1212;
wire n_1887;
wire n_1199;
wire n_2020;
wire n_1978;
wire n_2508;
wire n_2540;
wire n_1767;
wire n_1939;
wire n_2428;
wire n_1768;
wire n_1443;
wire n_2068;
wire n_2636;
wire n_2672;
wire n_1585;
wire n_1861;
wire n_2316;
wire n_1564;
wire n_1995;
wire n_1631;
wire n_2593;
wire n_1623;
wire n_2911;
wire n_861;
wire n_1828;
wire n_2364;
wire n_1389;
wire n_1131;
wire n_2641;
wire n_1798;
wire n_727;
wire n_1077;
wire n_1554;
wire n_1481;
wire n_1584;
wire n_2021;
wire n_1928;
wire n_2713;
wire n_828;
wire n_2938;
wire n_1438;
wire n_1973;
wire n_2314;
wire n_2939;
wire n_2156;
wire n_2494;
wire n_753;
wire n_2126;
wire n_747;
wire n_645;
wire n_1147;
wire n_1363;
wire n_2228;
wire n_1691;
wire n_1098;
wire n_584;
wire n_1366;
wire n_1518;
wire n_1187;
wire n_1361;
wire n_2034;
wire n_1693;
wire n_698;
wire n_2790;
wire n_2872;
wire n_2411;
wire n_2081;
wire n_1892;
wire n_1061;
wire n_2266;
wire n_2993;
wire n_682;
wire n_2061;
wire n_1373;
wire n_2449;
wire n_1686;
wire n_2131;
wire n_2526;
wire n_2830;
wire n_1302;
wire n_2083;
wire n_886;
wire n_2119;
wire n_1010;
wire n_883;
wire n_2207;
wire n_2044;
wire n_2542;
wire n_755;
wire n_2091;
wire n_2843;
wire n_1029;
wire n_2394;
wire n_770;
wire n_1572;
wire n_1635;
wire n_2827;
wire n_941;
wire n_1245;
wire n_1317;
wire n_2615;
wire n_2487;
wire n_2701;
wire n_2929;
wire n_632;
wire n_1329;
wire n_2409;
wire n_2637;
wire n_2337;
wire n_854;
wire n_2405;
wire n_2601;
wire n_2513;
wire n_1297;
wire n_714;
wire n_1369;
wire n_1912;
wire n_1734;
wire n_1876;
wire n_2666;
wire n_2323;
wire n_740;
wire n_1811;
wire n_928;
wire n_898;
wire n_1285;
wire n_967;
wire n_2561;
wire n_736;
wire n_2913;
wire n_2491;
wire n_1529;
wire n_1381;
wire n_1824;
wire n_2254;
wire n_1597;
wire n_1161;
wire n_1103;
wire n_1486;
wire n_1068;
wire n_617;
wire n_1833;
wire n_2914;
wire n_2371;
wire n_914;
wire n_1986;
wire n_2882;
wire n_1024;
wire n_1141;
wire n_1949;
wire n_1197;
wire n_2493;
wire n_2429;
wire n_2408;
wire n_1168;
wire n_865;
wire n_3000;
wire n_2115;
wire n_2013;
wire n_2140;
wire n_2134;
wire n_569;
wire n_2483;
wire n_2305;
wire n_600;
wire n_1556;
wire n_1192;
wire n_1646;
wire n_1290;
wire n_2514;
wire n_2466;
wire n_1759;
wire n_2048;
wire n_2760;
wire n_987;
wire n_750;
wire n_1299;
wire n_2942;
wire n_2096;
wire n_2129;
wire n_665;
wire n_1101;
wire n_2532;
wire n_2079;
wire n_2296;
wire n_1720;
wire n_880;
wire n_654;
wire n_2671;
wire n_1911;
wire n_2293;
wire n_731;
wire n_1336;
wire n_2734;
wire n_2870;
wire n_1166;
wire n_758;
wire n_720;
wire n_1390;
wire n_710;
wire n_2775;
wire n_1023;
wire n_568;
wire n_1358;
wire n_813;
wire n_2310;
wire n_1211;
wire n_1397;
wire n_2674;
wire n_1284;
wire n_2005;
wire n_1359;
wire n_1116;
wire n_2811;
wire n_1758;
wire n_791;
wire n_1532;
wire n_2848;
wire n_1419;
wire n_580;
wire n_2689;
wire n_1784;
wire n_1685;
wire n_1992;
wire n_1082;
wire n_1213;
wire n_2596;
wire n_2801;
wire n_980;
wire n_1193;
wire n_849;
wire n_1488;
wire n_2928;
wire n_2227;
wire n_2652;
wire n_1074;
wire n_759;
wire n_1379;
wire n_1721;
wire n_2972;
wire n_2627;
wire n_1827;
wire n_953;
wire n_1180;
wire n_1462;
wire n_2326;
wire n_1866;
wire n_1220;
wire n_1398;
wire n_2111;
wire n_2169;
wire n_1262;
wire n_1904;
wire n_2966;
wire n_1692;
wire n_2501;
wire n_2051;
wire n_1012;
wire n_1805;
wire n_960;
wire n_689;
wire n_1022;
wire n_1760;
wire n_676;
wire n_1240;
wire n_2173;
wire n_1183;
wire n_1204;
wire n_1151;
wire n_2824;
wire n_1814;
wire n_771;
wire n_2982;
wire n_999;
wire n_2634;
wire n_1092;
wire n_1808;
wire n_560;
wire n_2768;
wire n_2668;
wire n_1658;
wire n_1386;
wire n_2588;
wire n_2931;
wire n_2492;
wire n_910;
wire n_2291;
wire n_635;
wire n_844;
wire n_2172;
wire n_1728;
wire n_1020;
wire n_1142;
wire n_1385;
wire n_783;
wire n_2927;
wire n_1062;
wire n_1230;
wire n_1027;
wire n_1516;
wire n_2533;
wire n_1499;
wire n_1500;
wire n_2155;
wire n_2706;
wire n_1868;
wire n_966;
wire n_2303;
wire n_2104;
wire n_949;
wire n_704;
wire n_2148;
wire n_2357;
wire n_2618;
wire n_2653;
wire n_2855;
wire n_924;
wire n_2937;
wire n_2331;
wire n_1600;
wire n_1661;
wire n_2967;
wire n_1965;
wire n_3005;
wire n_1757;
wire n_699;
wire n_2136;
wire n_2403;
wire n_918;
wire n_2056;
wire n_1913;
wire n_672;
wire n_2702;
wire n_2054;
wire n_1039;
wire n_2226;
wire n_2407;
wire n_2791;
wire n_1043;
wire n_1402;
wire n_2267;
wire n_735;
wire n_1450;
wire n_2082;
wire n_2302;
wire n_2560;
wire n_2453;
wire n_2092;
wire n_566;
wire n_581;
wire n_1472;
wire n_1365;
wire n_2443;
wire n_2802;
wire n_2797;
wire n_2279;
wire n_1089;
wire n_1536;
wire n_1049;
wire n_1719;
wire n_2066;
wire n_1158;
wire n_1974;
wire n_2988;
wire n_763;
wire n_1882;
wire n_2770;
wire n_2961;
wire n_2704;
wire n_2996;
wire n_1915;
wire n_2836;
wire n_940;
wire n_1762;
wire n_2534;
wire n_1404;
wire n_788;
wire n_1736;
wire n_2907;
wire n_1160;
wire n_1442;
wire n_658;
wire n_1948;
wire n_2168;
wire n_1216;
wire n_2681;
wire n_1891;
wire n_1026;
wire n_2886;
wire n_1454;
wire n_1033;
wire n_627;
wire n_990;
wire n_1383;
wire n_1968;
wire n_2057;
wire n_2609;
wire n_2378;
wire n_888;
wire n_2749;
wire n_1325;
wire n_2754;
wire n_2014;
wire n_582;
wire n_1483;
wire n_1703;
wire n_653;
wire n_1205;
wire n_1822;
wire n_843;
wire n_1953;
wire n_1059;
wire n_2969;
wire n_799;
wire n_2692;
wire n_691;
wire n_1804;
wire n_1581;
wire n_1837;
wire n_1744;
wire n_1975;
wire n_1414;
wire n_2324;
wire n_2246;
wire n_2738;
wire n_1002;
wire n_1851;
wire n_1755;
wire n_2195;
wire n_2940;
wire n_1111;
wire n_1819;
wire n_1341;
wire n_1807;
wire n_2670;
wire n_2645;
wire n_2202;
wire n_1310;
wire n_1745;
wire n_1714;
wire n_612;
wire n_1958;
wire n_1611;
wire n_2559;
wire n_2262;
wire n_955;
wire n_1333;
wire n_1916;
wire n_2726;
wire n_2917;
wire n_2073;
wire n_952;
wire n_1675;
wire n_1947;
wire n_2165;
wire n_1640;
wire n_2016;
wire n_1551;
wire n_1145;
wire n_1533;
wire n_2307;
wire n_2515;
wire n_1511;
wire n_1791;
wire n_1113;
wire n_1651;
wire n_1966;
wire n_2058;
wire n_2678;
wire n_1468;
wire n_2327;
wire n_2656;
wire n_913;
wire n_2353;
wire n_1164;
wire n_2258;
wire n_1732;
wire n_2167;
wire n_1354;
wire n_2039;
wire n_1277;
wire n_1696;
wire n_1016;
wire n_680;
wire n_1355;
wire n_809;
wire n_2544;
wire n_856;
wire n_779;
wire n_2538;
wire n_2582;
wire n_1559;
wire n_2321;
wire n_2915;
wire n_1579;
wire n_1280;
wire n_2854;
wire n_2932;
wire n_1335;
wire n_2285;
wire n_1934;
wire n_1900;
wire n_2040;
wire n_2174;
wire n_1843;
wire n_2186;
wire n_2510;
wire n_2030;
wire n_2614;
wire n_2435;
wire n_1665;
wire n_2583;
wire n_1091;
wire n_1678;
wire n_1780;
wire n_2725;
wire n_1287;
wire n_2769;
wire n_1482;
wire n_860;
wire n_1525;
wire n_848;
wire n_661;
wire n_2100;
wire n_2349;
wire n_1902;
wire n_2536;
wire n_2474;
wire n_1194;
wire n_1150;
wire n_683;
wire n_620;
wire n_1399;
wire n_1903;
wire n_1674;
wire n_1849;
wire n_686;
wire n_572;
wire n_867;
wire n_983;
wire n_1417;
wire n_644;
wire n_577;
wire n_2282;
wire n_970;
wire n_2430;
wire n_2673;
wire n_921;
wire n_2676;
wire n_2926;
wire n_1534;
wire n_2912;
wire n_908;
wire n_1346;
wire n_565;
wire n_2834;
wire n_1123;
wire n_2710;
wire n_1272;
wire n_2497;
wire n_1393;
wire n_2970;
wire n_984;
wire n_1655;
wire n_2978;
wire n_1410;
wire n_988;
wire n_2368;
wire n_760;
wire n_1157;
wire n_806;
wire n_2657;
wire n_1186;
wire n_2065;
wire n_2901;
wire n_1743;
wire n_2743;
wire n_649;
wire n_1854;
wire n_866;
wire n_559;

INVx1_ASAP7_75t_L g558 ( 
.A(n_379),
.Y(n_558)
);

INVx2_ASAP7_75t_L g559 ( 
.A(n_129),
.Y(n_559)
);

CKINVDCx5p33_ASAP7_75t_R g560 ( 
.A(n_394),
.Y(n_560)
);

CKINVDCx5p33_ASAP7_75t_R g561 ( 
.A(n_296),
.Y(n_561)
);

CKINVDCx5p33_ASAP7_75t_R g562 ( 
.A(n_158),
.Y(n_562)
);

CKINVDCx5p33_ASAP7_75t_R g563 ( 
.A(n_194),
.Y(n_563)
);

CKINVDCx20_ASAP7_75t_R g564 ( 
.A(n_484),
.Y(n_564)
);

CKINVDCx5p33_ASAP7_75t_R g565 ( 
.A(n_150),
.Y(n_565)
);

CKINVDCx5p33_ASAP7_75t_R g566 ( 
.A(n_456),
.Y(n_566)
);

CKINVDCx5p33_ASAP7_75t_R g567 ( 
.A(n_425),
.Y(n_567)
);

CKINVDCx5p33_ASAP7_75t_R g568 ( 
.A(n_342),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_219),
.Y(n_569)
);

CKINVDCx5p33_ASAP7_75t_R g570 ( 
.A(n_508),
.Y(n_570)
);

CKINVDCx5p33_ASAP7_75t_R g571 ( 
.A(n_497),
.Y(n_571)
);

CKINVDCx5p33_ASAP7_75t_R g572 ( 
.A(n_416),
.Y(n_572)
);

CKINVDCx5p33_ASAP7_75t_R g573 ( 
.A(n_542),
.Y(n_573)
);

CKINVDCx5p33_ASAP7_75t_R g574 ( 
.A(n_513),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_504),
.Y(n_575)
);

CKINVDCx20_ASAP7_75t_R g576 ( 
.A(n_60),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_130),
.Y(n_577)
);

CKINVDCx5p33_ASAP7_75t_R g578 ( 
.A(n_507),
.Y(n_578)
);

CKINVDCx5p33_ASAP7_75t_R g579 ( 
.A(n_206),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_51),
.Y(n_580)
);

CKINVDCx5p33_ASAP7_75t_R g581 ( 
.A(n_190),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_398),
.Y(n_582)
);

CKINVDCx16_ASAP7_75t_R g583 ( 
.A(n_491),
.Y(n_583)
);

CKINVDCx5p33_ASAP7_75t_R g584 ( 
.A(n_135),
.Y(n_584)
);

CKINVDCx5p33_ASAP7_75t_R g585 ( 
.A(n_151),
.Y(n_585)
);

CKINVDCx20_ASAP7_75t_R g586 ( 
.A(n_274),
.Y(n_586)
);

CKINVDCx5p33_ASAP7_75t_R g587 ( 
.A(n_264),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_232),
.Y(n_588)
);

CKINVDCx5p33_ASAP7_75t_R g589 ( 
.A(n_461),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_130),
.Y(n_590)
);

CKINVDCx5p33_ASAP7_75t_R g591 ( 
.A(n_544),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_347),
.Y(n_592)
);

INVx2_ASAP7_75t_L g593 ( 
.A(n_188),
.Y(n_593)
);

BUFx3_ASAP7_75t_L g594 ( 
.A(n_359),
.Y(n_594)
);

CKINVDCx5p33_ASAP7_75t_R g595 ( 
.A(n_144),
.Y(n_595)
);

INVx2_ASAP7_75t_SL g596 ( 
.A(n_494),
.Y(n_596)
);

CKINVDCx5p33_ASAP7_75t_R g597 ( 
.A(n_329),
.Y(n_597)
);

CKINVDCx5p33_ASAP7_75t_R g598 ( 
.A(n_36),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_475),
.Y(n_599)
);

BUFx10_ASAP7_75t_L g600 ( 
.A(n_323),
.Y(n_600)
);

BUFx3_ASAP7_75t_L g601 ( 
.A(n_22),
.Y(n_601)
);

CKINVDCx5p33_ASAP7_75t_R g602 ( 
.A(n_405),
.Y(n_602)
);

CKINVDCx5p33_ASAP7_75t_R g603 ( 
.A(n_428),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_235),
.Y(n_604)
);

CKINVDCx5p33_ASAP7_75t_R g605 ( 
.A(n_250),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_16),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_362),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_454),
.Y(n_608)
);

CKINVDCx5p33_ASAP7_75t_R g609 ( 
.A(n_96),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_102),
.Y(n_610)
);

CKINVDCx5p33_ASAP7_75t_R g611 ( 
.A(n_314),
.Y(n_611)
);

INVx2_ASAP7_75t_L g612 ( 
.A(n_498),
.Y(n_612)
);

BUFx10_ASAP7_75t_L g613 ( 
.A(n_362),
.Y(n_613)
);

CKINVDCx5p33_ASAP7_75t_R g614 ( 
.A(n_409),
.Y(n_614)
);

CKINVDCx5p33_ASAP7_75t_R g615 ( 
.A(n_418),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_546),
.Y(n_616)
);

CKINVDCx20_ASAP7_75t_R g617 ( 
.A(n_144),
.Y(n_617)
);

CKINVDCx5p33_ASAP7_75t_R g618 ( 
.A(n_124),
.Y(n_618)
);

CKINVDCx5p33_ASAP7_75t_R g619 ( 
.A(n_286),
.Y(n_619)
);

CKINVDCx5p33_ASAP7_75t_R g620 ( 
.A(n_458),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_223),
.Y(n_621)
);

CKINVDCx5p33_ASAP7_75t_R g622 ( 
.A(n_549),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_224),
.Y(n_623)
);

INVx2_ASAP7_75t_SL g624 ( 
.A(n_169),
.Y(n_624)
);

CKINVDCx5p33_ASAP7_75t_R g625 ( 
.A(n_318),
.Y(n_625)
);

CKINVDCx20_ASAP7_75t_R g626 ( 
.A(n_556),
.Y(n_626)
);

CKINVDCx5p33_ASAP7_75t_R g627 ( 
.A(n_444),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_310),
.Y(n_628)
);

CKINVDCx5p33_ASAP7_75t_R g629 ( 
.A(n_43),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_223),
.Y(n_630)
);

CKINVDCx20_ASAP7_75t_R g631 ( 
.A(n_43),
.Y(n_631)
);

CKINVDCx5p33_ASAP7_75t_R g632 ( 
.A(n_31),
.Y(n_632)
);

CKINVDCx5p33_ASAP7_75t_R g633 ( 
.A(n_373),
.Y(n_633)
);

INVx2_ASAP7_75t_L g634 ( 
.A(n_471),
.Y(n_634)
);

INVxp67_ASAP7_75t_L g635 ( 
.A(n_247),
.Y(n_635)
);

CKINVDCx5p33_ASAP7_75t_R g636 ( 
.A(n_496),
.Y(n_636)
);

BUFx10_ASAP7_75t_L g637 ( 
.A(n_243),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_417),
.Y(n_638)
);

CKINVDCx5p33_ASAP7_75t_R g639 ( 
.A(n_259),
.Y(n_639)
);

CKINVDCx5p33_ASAP7_75t_R g640 ( 
.A(n_11),
.Y(n_640)
);

BUFx10_ASAP7_75t_L g641 ( 
.A(n_10),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_242),
.Y(n_642)
);

CKINVDCx5p33_ASAP7_75t_R g643 ( 
.A(n_263),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_325),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_495),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_139),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_474),
.Y(n_647)
);

CKINVDCx5p33_ASAP7_75t_R g648 ( 
.A(n_396),
.Y(n_648)
);

CKINVDCx5p33_ASAP7_75t_R g649 ( 
.A(n_411),
.Y(n_649)
);

CKINVDCx5p33_ASAP7_75t_R g650 ( 
.A(n_227),
.Y(n_650)
);

CKINVDCx5p33_ASAP7_75t_R g651 ( 
.A(n_73),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_258),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_156),
.Y(n_653)
);

BUFx3_ASAP7_75t_L g654 ( 
.A(n_287),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_46),
.Y(n_655)
);

CKINVDCx16_ASAP7_75t_R g656 ( 
.A(n_352),
.Y(n_656)
);

BUFx10_ASAP7_75t_L g657 ( 
.A(n_85),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_11),
.Y(n_658)
);

CKINVDCx5p33_ASAP7_75t_R g659 ( 
.A(n_88),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_473),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_4),
.Y(n_661)
);

CKINVDCx5p33_ASAP7_75t_R g662 ( 
.A(n_436),
.Y(n_662)
);

CKINVDCx5p33_ASAP7_75t_R g663 ( 
.A(n_81),
.Y(n_663)
);

CKINVDCx5p33_ASAP7_75t_R g664 ( 
.A(n_550),
.Y(n_664)
);

CKINVDCx5p33_ASAP7_75t_R g665 ( 
.A(n_392),
.Y(n_665)
);

CKINVDCx5p33_ASAP7_75t_R g666 ( 
.A(n_91),
.Y(n_666)
);

CKINVDCx5p33_ASAP7_75t_R g667 ( 
.A(n_259),
.Y(n_667)
);

HB1xp67_ASAP7_75t_L g668 ( 
.A(n_512),
.Y(n_668)
);

CKINVDCx5p33_ASAP7_75t_R g669 ( 
.A(n_506),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_49),
.Y(n_670)
);

BUFx10_ASAP7_75t_L g671 ( 
.A(n_102),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_19),
.Y(n_672)
);

CKINVDCx5p33_ASAP7_75t_R g673 ( 
.A(n_162),
.Y(n_673)
);

CKINVDCx5p33_ASAP7_75t_R g674 ( 
.A(n_268),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_118),
.Y(n_675)
);

CKINVDCx5p33_ASAP7_75t_R g676 ( 
.A(n_327),
.Y(n_676)
);

CKINVDCx5p33_ASAP7_75t_R g677 ( 
.A(n_334),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_244),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_47),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_3),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_369),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_77),
.Y(n_682)
);

CKINVDCx5p33_ASAP7_75t_R g683 ( 
.A(n_519),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_280),
.Y(n_684)
);

BUFx6f_ASAP7_75t_L g685 ( 
.A(n_235),
.Y(n_685)
);

CKINVDCx5p33_ASAP7_75t_R g686 ( 
.A(n_413),
.Y(n_686)
);

CKINVDCx5p33_ASAP7_75t_R g687 ( 
.A(n_322),
.Y(n_687)
);

CKINVDCx5p33_ASAP7_75t_R g688 ( 
.A(n_357),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_91),
.Y(n_689)
);

CKINVDCx5p33_ASAP7_75t_R g690 ( 
.A(n_101),
.Y(n_690)
);

CKINVDCx5p33_ASAP7_75t_R g691 ( 
.A(n_25),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_121),
.Y(n_692)
);

BUFx3_ASAP7_75t_L g693 ( 
.A(n_490),
.Y(n_693)
);

CKINVDCx20_ASAP7_75t_R g694 ( 
.A(n_459),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_122),
.Y(n_695)
);

BUFx2_ASAP7_75t_SL g696 ( 
.A(n_127),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_1),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_9),
.Y(n_698)
);

CKINVDCx5p33_ASAP7_75t_R g699 ( 
.A(n_388),
.Y(n_699)
);

INVx1_ASAP7_75t_SL g700 ( 
.A(n_329),
.Y(n_700)
);

CKINVDCx5p33_ASAP7_75t_R g701 ( 
.A(n_419),
.Y(n_701)
);

CKINVDCx5p33_ASAP7_75t_R g702 ( 
.A(n_452),
.Y(n_702)
);

CKINVDCx20_ASAP7_75t_R g703 ( 
.A(n_54),
.Y(n_703)
);

CKINVDCx20_ASAP7_75t_R g704 ( 
.A(n_476),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_31),
.Y(n_705)
);

CKINVDCx16_ASAP7_75t_R g706 ( 
.A(n_172),
.Y(n_706)
);

CKINVDCx5p33_ASAP7_75t_R g707 ( 
.A(n_70),
.Y(n_707)
);

INVx1_ASAP7_75t_SL g708 ( 
.A(n_149),
.Y(n_708)
);

CKINVDCx20_ASAP7_75t_R g709 ( 
.A(n_40),
.Y(n_709)
);

INVx1_ASAP7_75t_SL g710 ( 
.A(n_446),
.Y(n_710)
);

CKINVDCx14_ASAP7_75t_R g711 ( 
.A(n_25),
.Y(n_711)
);

INVx1_ASAP7_75t_SL g712 ( 
.A(n_156),
.Y(n_712)
);

CKINVDCx5p33_ASAP7_75t_R g713 ( 
.A(n_477),
.Y(n_713)
);

CKINVDCx5p33_ASAP7_75t_R g714 ( 
.A(n_438),
.Y(n_714)
);

CKINVDCx5p33_ASAP7_75t_R g715 ( 
.A(n_538),
.Y(n_715)
);

BUFx2_ASAP7_75t_L g716 ( 
.A(n_167),
.Y(n_716)
);

BUFx10_ASAP7_75t_L g717 ( 
.A(n_389),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_50),
.Y(n_718)
);

INVx2_ASAP7_75t_L g719 ( 
.A(n_152),
.Y(n_719)
);

CKINVDCx14_ASAP7_75t_R g720 ( 
.A(n_499),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_274),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_360),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_400),
.Y(n_723)
);

CKINVDCx5p33_ASAP7_75t_R g724 ( 
.A(n_505),
.Y(n_724)
);

CKINVDCx20_ASAP7_75t_R g725 ( 
.A(n_384),
.Y(n_725)
);

BUFx6f_ASAP7_75t_L g726 ( 
.A(n_524),
.Y(n_726)
);

CKINVDCx5p33_ASAP7_75t_R g727 ( 
.A(n_232),
.Y(n_727)
);

INVx2_ASAP7_75t_SL g728 ( 
.A(n_161),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_540),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_246),
.Y(n_730)
);

CKINVDCx5p33_ASAP7_75t_R g731 ( 
.A(n_331),
.Y(n_731)
);

CKINVDCx5p33_ASAP7_75t_R g732 ( 
.A(n_397),
.Y(n_732)
);

INVx1_ASAP7_75t_SL g733 ( 
.A(n_478),
.Y(n_733)
);

CKINVDCx5p33_ASAP7_75t_R g734 ( 
.A(n_358),
.Y(n_734)
);

CKINVDCx5p33_ASAP7_75t_R g735 ( 
.A(n_220),
.Y(n_735)
);

BUFx3_ASAP7_75t_L g736 ( 
.A(n_177),
.Y(n_736)
);

CKINVDCx5p33_ASAP7_75t_R g737 ( 
.A(n_393),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_386),
.Y(n_738)
);

INVx1_ASAP7_75t_SL g739 ( 
.A(n_406),
.Y(n_739)
);

CKINVDCx5p33_ASAP7_75t_R g740 ( 
.A(n_276),
.Y(n_740)
);

CKINVDCx5p33_ASAP7_75t_R g741 ( 
.A(n_46),
.Y(n_741)
);

CKINVDCx20_ASAP7_75t_R g742 ( 
.A(n_260),
.Y(n_742)
);

CKINVDCx5p33_ASAP7_75t_R g743 ( 
.A(n_224),
.Y(n_743)
);

CKINVDCx5p33_ASAP7_75t_R g744 ( 
.A(n_128),
.Y(n_744)
);

CKINVDCx5p33_ASAP7_75t_R g745 ( 
.A(n_153),
.Y(n_745)
);

BUFx5_ASAP7_75t_L g746 ( 
.A(n_41),
.Y(n_746)
);

CKINVDCx20_ASAP7_75t_R g747 ( 
.A(n_415),
.Y(n_747)
);

CKINVDCx5p33_ASAP7_75t_R g748 ( 
.A(n_207),
.Y(n_748)
);

INVx2_ASAP7_75t_SL g749 ( 
.A(n_57),
.Y(n_749)
);

INVx2_ASAP7_75t_L g750 ( 
.A(n_399),
.Y(n_750)
);

CKINVDCx5p33_ASAP7_75t_R g751 ( 
.A(n_16),
.Y(n_751)
);

CKINVDCx5p33_ASAP7_75t_R g752 ( 
.A(n_429),
.Y(n_752)
);

CKINVDCx5p33_ASAP7_75t_R g753 ( 
.A(n_146),
.Y(n_753)
);

CKINVDCx5p33_ASAP7_75t_R g754 ( 
.A(n_128),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_225),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_120),
.Y(n_756)
);

CKINVDCx5p33_ASAP7_75t_R g757 ( 
.A(n_22),
.Y(n_757)
);

CKINVDCx5p33_ASAP7_75t_R g758 ( 
.A(n_404),
.Y(n_758)
);

BUFx3_ASAP7_75t_L g759 ( 
.A(n_311),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_182),
.Y(n_760)
);

INVx2_ASAP7_75t_L g761 ( 
.A(n_236),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_137),
.Y(n_762)
);

CKINVDCx5p33_ASAP7_75t_R g763 ( 
.A(n_106),
.Y(n_763)
);

CKINVDCx5p33_ASAP7_75t_R g764 ( 
.A(n_332),
.Y(n_764)
);

CKINVDCx5p33_ASAP7_75t_R g765 ( 
.A(n_100),
.Y(n_765)
);

CKINVDCx5p33_ASAP7_75t_R g766 ( 
.A(n_23),
.Y(n_766)
);

INVx2_ASAP7_75t_L g767 ( 
.A(n_276),
.Y(n_767)
);

INVx2_ASAP7_75t_L g768 ( 
.A(n_124),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_213),
.Y(n_769)
);

INVx2_ASAP7_75t_SL g770 ( 
.A(n_181),
.Y(n_770)
);

BUFx2_ASAP7_75t_L g771 ( 
.A(n_301),
.Y(n_771)
);

CKINVDCx5p33_ASAP7_75t_R g772 ( 
.A(n_383),
.Y(n_772)
);

CKINVDCx20_ASAP7_75t_R g773 ( 
.A(n_283),
.Y(n_773)
);

CKINVDCx5p33_ASAP7_75t_R g774 ( 
.A(n_402),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_50),
.Y(n_775)
);

BUFx2_ASAP7_75t_L g776 ( 
.A(n_313),
.Y(n_776)
);

CKINVDCx5p33_ASAP7_75t_R g777 ( 
.A(n_238),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_186),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_209),
.Y(n_779)
);

CKINVDCx5p33_ASAP7_75t_R g780 ( 
.A(n_184),
.Y(n_780)
);

CKINVDCx20_ASAP7_75t_R g781 ( 
.A(n_76),
.Y(n_781)
);

CKINVDCx20_ASAP7_75t_R g782 ( 
.A(n_412),
.Y(n_782)
);

CKINVDCx5p33_ASAP7_75t_R g783 ( 
.A(n_108),
.Y(n_783)
);

INVx1_ASAP7_75t_L g784 ( 
.A(n_364),
.Y(n_784)
);

CKINVDCx5p33_ASAP7_75t_R g785 ( 
.A(n_79),
.Y(n_785)
);

CKINVDCx5p33_ASAP7_75t_R g786 ( 
.A(n_175),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_20),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_387),
.Y(n_788)
);

CKINVDCx20_ASAP7_75t_R g789 ( 
.A(n_427),
.Y(n_789)
);

CKINVDCx5p33_ASAP7_75t_R g790 ( 
.A(n_137),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_57),
.Y(n_791)
);

CKINVDCx5p33_ASAP7_75t_R g792 ( 
.A(n_216),
.Y(n_792)
);

CKINVDCx20_ASAP7_75t_R g793 ( 
.A(n_391),
.Y(n_793)
);

INVx1_ASAP7_75t_SL g794 ( 
.A(n_375),
.Y(n_794)
);

CKINVDCx5p33_ASAP7_75t_R g795 ( 
.A(n_466),
.Y(n_795)
);

CKINVDCx5p33_ASAP7_75t_R g796 ( 
.A(n_335),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_172),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_49),
.Y(n_798)
);

CKINVDCx20_ASAP7_75t_R g799 ( 
.A(n_86),
.Y(n_799)
);

BUFx3_ASAP7_75t_L g800 ( 
.A(n_10),
.Y(n_800)
);

BUFx2_ASAP7_75t_L g801 ( 
.A(n_482),
.Y(n_801)
);

CKINVDCx5p33_ASAP7_75t_R g802 ( 
.A(n_138),
.Y(n_802)
);

CKINVDCx5p33_ASAP7_75t_R g803 ( 
.A(n_501),
.Y(n_803)
);

CKINVDCx5p33_ASAP7_75t_R g804 ( 
.A(n_173),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_129),
.Y(n_805)
);

INVx2_ASAP7_75t_L g806 ( 
.A(n_222),
.Y(n_806)
);

CKINVDCx5p33_ASAP7_75t_R g807 ( 
.A(n_502),
.Y(n_807)
);

CKINVDCx5p33_ASAP7_75t_R g808 ( 
.A(n_17),
.Y(n_808)
);

CKINVDCx5p33_ASAP7_75t_R g809 ( 
.A(n_434),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_191),
.Y(n_810)
);

CKINVDCx5p33_ASAP7_75t_R g811 ( 
.A(n_545),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_435),
.Y(n_812)
);

CKINVDCx5p33_ASAP7_75t_R g813 ( 
.A(n_18),
.Y(n_813)
);

CKINVDCx5p33_ASAP7_75t_R g814 ( 
.A(n_443),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_190),
.Y(n_815)
);

CKINVDCx5p33_ASAP7_75t_R g816 ( 
.A(n_535),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_140),
.Y(n_817)
);

CKINVDCx5p33_ASAP7_75t_R g818 ( 
.A(n_366),
.Y(n_818)
);

CKINVDCx20_ASAP7_75t_R g819 ( 
.A(n_151),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_343),
.Y(n_820)
);

CKINVDCx20_ASAP7_75t_R g821 ( 
.A(n_271),
.Y(n_821)
);

CKINVDCx5p33_ASAP7_75t_R g822 ( 
.A(n_252),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_510),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_472),
.Y(n_824)
);

CKINVDCx20_ASAP7_75t_R g825 ( 
.A(n_307),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_228),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_500),
.Y(n_827)
);

CKINVDCx5p33_ASAP7_75t_R g828 ( 
.A(n_395),
.Y(n_828)
);

CKINVDCx5p33_ASAP7_75t_R g829 ( 
.A(n_155),
.Y(n_829)
);

CKINVDCx5p33_ASAP7_75t_R g830 ( 
.A(n_367),
.Y(n_830)
);

CKINVDCx5p33_ASAP7_75t_R g831 ( 
.A(n_332),
.Y(n_831)
);

CKINVDCx5p33_ASAP7_75t_R g832 ( 
.A(n_227),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_234),
.Y(n_833)
);

BUFx3_ASAP7_75t_L g834 ( 
.A(n_243),
.Y(n_834)
);

CKINVDCx5p33_ASAP7_75t_R g835 ( 
.A(n_78),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_468),
.Y(n_836)
);

CKINVDCx5p33_ASAP7_75t_R g837 ( 
.A(n_511),
.Y(n_837)
);

INVx2_ASAP7_75t_SL g838 ( 
.A(n_176),
.Y(n_838)
);

CKINVDCx16_ASAP7_75t_R g839 ( 
.A(n_207),
.Y(n_839)
);

CKINVDCx5p33_ASAP7_75t_R g840 ( 
.A(n_273),
.Y(n_840)
);

BUFx6f_ASAP7_75t_L g841 ( 
.A(n_263),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_162),
.Y(n_842)
);

BUFx2_ASAP7_75t_SL g843 ( 
.A(n_30),
.Y(n_843)
);

INVx1_ASAP7_75t_SL g844 ( 
.A(n_206),
.Y(n_844)
);

BUFx10_ASAP7_75t_L g845 ( 
.A(n_230),
.Y(n_845)
);

BUFx10_ASAP7_75t_L g846 ( 
.A(n_226),
.Y(n_846)
);

BUFx6f_ASAP7_75t_L g847 ( 
.A(n_522),
.Y(n_847)
);

INVx1_ASAP7_75t_L g848 ( 
.A(n_552),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_503),
.Y(n_849)
);

CKINVDCx5p33_ASAP7_75t_R g850 ( 
.A(n_59),
.Y(n_850)
);

CKINVDCx5p33_ASAP7_75t_R g851 ( 
.A(n_244),
.Y(n_851)
);

CKINVDCx5p33_ASAP7_75t_R g852 ( 
.A(n_448),
.Y(n_852)
);

INVx1_ASAP7_75t_L g853 ( 
.A(n_368),
.Y(n_853)
);

INVx2_ASAP7_75t_L g854 ( 
.A(n_303),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_229),
.Y(n_855)
);

CKINVDCx5p33_ASAP7_75t_R g856 ( 
.A(n_229),
.Y(n_856)
);

CKINVDCx5p33_ASAP7_75t_R g857 ( 
.A(n_449),
.Y(n_857)
);

INVx2_ASAP7_75t_L g858 ( 
.A(n_423),
.Y(n_858)
);

INVx1_ASAP7_75t_SL g859 ( 
.A(n_169),
.Y(n_859)
);

CKINVDCx5p33_ASAP7_75t_R g860 ( 
.A(n_381),
.Y(n_860)
);

INVx1_ASAP7_75t_L g861 ( 
.A(n_114),
.Y(n_861)
);

INVx1_ASAP7_75t_L g862 ( 
.A(n_369),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_297),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_71),
.Y(n_864)
);

CKINVDCx5p33_ASAP7_75t_R g865 ( 
.A(n_340),
.Y(n_865)
);

CKINVDCx5p33_ASAP7_75t_R g866 ( 
.A(n_526),
.Y(n_866)
);

CKINVDCx5p33_ASAP7_75t_R g867 ( 
.A(n_359),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_321),
.Y(n_868)
);

CKINVDCx5p33_ASAP7_75t_R g869 ( 
.A(n_131),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_37),
.Y(n_870)
);

CKINVDCx5p33_ASAP7_75t_R g871 ( 
.A(n_469),
.Y(n_871)
);

BUFx2_ASAP7_75t_L g872 ( 
.A(n_509),
.Y(n_872)
);

CKINVDCx5p33_ASAP7_75t_R g873 ( 
.A(n_492),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_306),
.Y(n_874)
);

CKINVDCx5p33_ASAP7_75t_R g875 ( 
.A(n_307),
.Y(n_875)
);

BUFx3_ASAP7_75t_L g876 ( 
.A(n_205),
.Y(n_876)
);

CKINVDCx5p33_ASAP7_75t_R g877 ( 
.A(n_390),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_131),
.Y(n_878)
);

CKINVDCx5p33_ASAP7_75t_R g879 ( 
.A(n_493),
.Y(n_879)
);

CKINVDCx5p33_ASAP7_75t_R g880 ( 
.A(n_179),
.Y(n_880)
);

CKINVDCx5p33_ASAP7_75t_R g881 ( 
.A(n_231),
.Y(n_881)
);

CKINVDCx5p33_ASAP7_75t_R g882 ( 
.A(n_316),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_179),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_189),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_485),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_385),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_101),
.Y(n_887)
);

INVx2_ASAP7_75t_L g888 ( 
.A(n_66),
.Y(n_888)
);

CKINVDCx5p33_ASAP7_75t_R g889 ( 
.A(n_370),
.Y(n_889)
);

BUFx3_ASAP7_75t_L g890 ( 
.A(n_336),
.Y(n_890)
);

INVx1_ASAP7_75t_L g891 ( 
.A(n_305),
.Y(n_891)
);

CKINVDCx5p33_ASAP7_75t_R g892 ( 
.A(n_366),
.Y(n_892)
);

INVx2_ASAP7_75t_SL g893 ( 
.A(n_348),
.Y(n_893)
);

INVx1_ASAP7_75t_L g894 ( 
.A(n_83),
.Y(n_894)
);

CKINVDCx5p33_ASAP7_75t_R g895 ( 
.A(n_79),
.Y(n_895)
);

CKINVDCx5p33_ASAP7_75t_R g896 ( 
.A(n_528),
.Y(n_896)
);

BUFx6f_ASAP7_75t_L g897 ( 
.A(n_311),
.Y(n_897)
);

INVx1_ASAP7_75t_L g898 ( 
.A(n_378),
.Y(n_898)
);

INVx2_ASAP7_75t_L g899 ( 
.A(n_17),
.Y(n_899)
);

INVx1_ASAP7_75t_L g900 ( 
.A(n_178),
.Y(n_900)
);

CKINVDCx5p33_ASAP7_75t_R g901 ( 
.A(n_426),
.Y(n_901)
);

CKINVDCx5p33_ASAP7_75t_R g902 ( 
.A(n_455),
.Y(n_902)
);

CKINVDCx5p33_ASAP7_75t_R g903 ( 
.A(n_47),
.Y(n_903)
);

CKINVDCx5p33_ASAP7_75t_R g904 ( 
.A(n_273),
.Y(n_904)
);

CKINVDCx5p33_ASAP7_75t_R g905 ( 
.A(n_408),
.Y(n_905)
);

CKINVDCx5p33_ASAP7_75t_R g906 ( 
.A(n_29),
.Y(n_906)
);

CKINVDCx20_ASAP7_75t_R g907 ( 
.A(n_555),
.Y(n_907)
);

CKINVDCx5p33_ASAP7_75t_R g908 ( 
.A(n_119),
.Y(n_908)
);

CKINVDCx20_ASAP7_75t_R g909 ( 
.A(n_533),
.Y(n_909)
);

CKINVDCx20_ASAP7_75t_R g910 ( 
.A(n_75),
.Y(n_910)
);

CKINVDCx5p33_ASAP7_75t_R g911 ( 
.A(n_221),
.Y(n_911)
);

CKINVDCx20_ASAP7_75t_R g912 ( 
.A(n_403),
.Y(n_912)
);

CKINVDCx20_ASAP7_75t_R g913 ( 
.A(n_656),
.Y(n_913)
);

INVx1_ASAP7_75t_L g914 ( 
.A(n_668),
.Y(n_914)
);

CKINVDCx5p33_ASAP7_75t_R g915 ( 
.A(n_711),
.Y(n_915)
);

CKINVDCx14_ASAP7_75t_R g916 ( 
.A(n_720),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_624),
.Y(n_917)
);

INVx1_ASAP7_75t_L g918 ( 
.A(n_624),
.Y(n_918)
);

INVx1_ASAP7_75t_L g919 ( 
.A(n_728),
.Y(n_919)
);

CKINVDCx20_ASAP7_75t_R g920 ( 
.A(n_706),
.Y(n_920)
);

CKINVDCx20_ASAP7_75t_R g921 ( 
.A(n_839),
.Y(n_921)
);

HB1xp67_ASAP7_75t_L g922 ( 
.A(n_716),
.Y(n_922)
);

INVxp33_ASAP7_75t_SL g923 ( 
.A(n_561),
.Y(n_923)
);

NOR2xp33_ASAP7_75t_L g924 ( 
.A(n_596),
.B(n_0),
.Y(n_924)
);

INVx1_ASAP7_75t_L g925 ( 
.A(n_728),
.Y(n_925)
);

CKINVDCx5p33_ASAP7_75t_R g926 ( 
.A(n_564),
.Y(n_926)
);

HB1xp67_ASAP7_75t_L g927 ( 
.A(n_771),
.Y(n_927)
);

INVx1_ASAP7_75t_L g928 ( 
.A(n_749),
.Y(n_928)
);

INVx1_ASAP7_75t_L g929 ( 
.A(n_749),
.Y(n_929)
);

INVx1_ASAP7_75t_L g930 ( 
.A(n_770),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_770),
.Y(n_931)
);

CKINVDCx5p33_ASAP7_75t_R g932 ( 
.A(n_626),
.Y(n_932)
);

CKINVDCx20_ASAP7_75t_R g933 ( 
.A(n_576),
.Y(n_933)
);

CKINVDCx20_ASAP7_75t_R g934 ( 
.A(n_586),
.Y(n_934)
);

INVx1_ASAP7_75t_L g935 ( 
.A(n_838),
.Y(n_935)
);

NOR2xp33_ASAP7_75t_L g936 ( 
.A(n_596),
.B(n_0),
.Y(n_936)
);

INVxp33_ASAP7_75t_L g937 ( 
.A(n_776),
.Y(n_937)
);

CKINVDCx5p33_ASAP7_75t_R g938 ( 
.A(n_583),
.Y(n_938)
);

NOR2xp33_ASAP7_75t_L g939 ( 
.A(n_801),
.B(n_1),
.Y(n_939)
);

AND2x2_ASAP7_75t_L g940 ( 
.A(n_872),
.B(n_2),
.Y(n_940)
);

HB1xp67_ASAP7_75t_L g941 ( 
.A(n_561),
.Y(n_941)
);

CKINVDCx16_ASAP7_75t_R g942 ( 
.A(n_600),
.Y(n_942)
);

CKINVDCx20_ASAP7_75t_R g943 ( 
.A(n_617),
.Y(n_943)
);

CKINVDCx5p33_ASAP7_75t_R g944 ( 
.A(n_912),
.Y(n_944)
);

NOR2xp67_ASAP7_75t_L g945 ( 
.A(n_838),
.B(n_2),
.Y(n_945)
);

INVx1_ASAP7_75t_L g946 ( 
.A(n_893),
.Y(n_946)
);

NOR2xp67_ASAP7_75t_L g947 ( 
.A(n_893),
.B(n_635),
.Y(n_947)
);

INVx1_ASAP7_75t_L g948 ( 
.A(n_594),
.Y(n_948)
);

CKINVDCx20_ASAP7_75t_R g949 ( 
.A(n_631),
.Y(n_949)
);

CKINVDCx20_ASAP7_75t_R g950 ( 
.A(n_703),
.Y(n_950)
);

INVx1_ASAP7_75t_L g951 ( 
.A(n_601),
.Y(n_951)
);

CKINVDCx16_ASAP7_75t_R g952 ( 
.A(n_600),
.Y(n_952)
);

INVxp67_ASAP7_75t_SL g953 ( 
.A(n_654),
.Y(n_953)
);

CKINVDCx20_ASAP7_75t_R g954 ( 
.A(n_709),
.Y(n_954)
);

INVx1_ASAP7_75t_L g955 ( 
.A(n_654),
.Y(n_955)
);

CKINVDCx5p33_ASAP7_75t_R g956 ( 
.A(n_694),
.Y(n_956)
);

CKINVDCx5p33_ASAP7_75t_R g957 ( 
.A(n_704),
.Y(n_957)
);

INVxp67_ASAP7_75t_SL g958 ( 
.A(n_736),
.Y(n_958)
);

CKINVDCx20_ASAP7_75t_R g959 ( 
.A(n_742),
.Y(n_959)
);

CKINVDCx20_ASAP7_75t_R g960 ( 
.A(n_773),
.Y(n_960)
);

INVx1_ASAP7_75t_L g961 ( 
.A(n_736),
.Y(n_961)
);

CKINVDCx5p33_ASAP7_75t_R g962 ( 
.A(n_725),
.Y(n_962)
);

INVxp67_ASAP7_75t_SL g963 ( 
.A(n_759),
.Y(n_963)
);

CKINVDCx20_ASAP7_75t_R g964 ( 
.A(n_781),
.Y(n_964)
);

INVxp67_ASAP7_75t_SL g965 ( 
.A(n_800),
.Y(n_965)
);

CKINVDCx5p33_ASAP7_75t_R g966 ( 
.A(n_562),
.Y(n_966)
);

INVx1_ASAP7_75t_L g967 ( 
.A(n_800),
.Y(n_967)
);

INVx1_ASAP7_75t_L g968 ( 
.A(n_834),
.Y(n_968)
);

HB1xp67_ASAP7_75t_L g969 ( 
.A(n_562),
.Y(n_969)
);

CKINVDCx16_ASAP7_75t_R g970 ( 
.A(n_600),
.Y(n_970)
);

CKINVDCx20_ASAP7_75t_R g971 ( 
.A(n_799),
.Y(n_971)
);

CKINVDCx5p33_ASAP7_75t_R g972 ( 
.A(n_747),
.Y(n_972)
);

INVxp33_ASAP7_75t_SL g973 ( 
.A(n_563),
.Y(n_973)
);

CKINVDCx20_ASAP7_75t_R g974 ( 
.A(n_819),
.Y(n_974)
);

INVx1_ASAP7_75t_L g975 ( 
.A(n_876),
.Y(n_975)
);

CKINVDCx20_ASAP7_75t_R g976 ( 
.A(n_821),
.Y(n_976)
);

CKINVDCx5p33_ASAP7_75t_R g977 ( 
.A(n_782),
.Y(n_977)
);

INVx1_ASAP7_75t_L g978 ( 
.A(n_876),
.Y(n_978)
);

INVx1_ASAP7_75t_L g979 ( 
.A(n_890),
.Y(n_979)
);

HB1xp67_ASAP7_75t_L g980 ( 
.A(n_563),
.Y(n_980)
);

INVx1_ASAP7_75t_L g981 ( 
.A(n_890),
.Y(n_981)
);

CKINVDCx20_ASAP7_75t_R g982 ( 
.A(n_825),
.Y(n_982)
);

INVx1_ASAP7_75t_L g983 ( 
.A(n_559),
.Y(n_983)
);

CKINVDCx5p33_ASAP7_75t_R g984 ( 
.A(n_789),
.Y(n_984)
);

AND2x2_ASAP7_75t_L g985 ( 
.A(n_613),
.B(n_3),
.Y(n_985)
);

CKINVDCx5p33_ASAP7_75t_R g986 ( 
.A(n_793),
.Y(n_986)
);

CKINVDCx5p33_ASAP7_75t_R g987 ( 
.A(n_907),
.Y(n_987)
);

CKINVDCx5p33_ASAP7_75t_R g988 ( 
.A(n_909),
.Y(n_988)
);

CKINVDCx5p33_ASAP7_75t_R g989 ( 
.A(n_560),
.Y(n_989)
);

INVx1_ASAP7_75t_L g990 ( 
.A(n_559),
.Y(n_990)
);

INVx2_ASAP7_75t_L g991 ( 
.A(n_746),
.Y(n_991)
);

CKINVDCx5p33_ASAP7_75t_R g992 ( 
.A(n_560),
.Y(n_992)
);

INVx1_ASAP7_75t_L g993 ( 
.A(n_593),
.Y(n_993)
);

CKINVDCx5p33_ASAP7_75t_R g994 ( 
.A(n_566),
.Y(n_994)
);

CKINVDCx5p33_ASAP7_75t_R g995 ( 
.A(n_566),
.Y(n_995)
);

INVx1_ASAP7_75t_L g996 ( 
.A(n_719),
.Y(n_996)
);

NOR2xp33_ASAP7_75t_L g997 ( 
.A(n_558),
.B(n_4),
.Y(n_997)
);

CKINVDCx5p33_ASAP7_75t_R g998 ( 
.A(n_567),
.Y(n_998)
);

NOR2xp33_ASAP7_75t_L g999 ( 
.A(n_575),
.B(n_5),
.Y(n_999)
);

CKINVDCx5p33_ASAP7_75t_R g1000 ( 
.A(n_567),
.Y(n_1000)
);

CKINVDCx20_ASAP7_75t_R g1001 ( 
.A(n_910),
.Y(n_1001)
);

INVx1_ASAP7_75t_L g1002 ( 
.A(n_719),
.Y(n_1002)
);

INVx1_ASAP7_75t_L g1003 ( 
.A(n_761),
.Y(n_1003)
);

INVx1_ASAP7_75t_L g1004 ( 
.A(n_761),
.Y(n_1004)
);

NOR2xp33_ASAP7_75t_L g1005 ( 
.A(n_582),
.B(n_5),
.Y(n_1005)
);

NAND2xp5_ASAP7_75t_L g1006 ( 
.A(n_565),
.B(n_6),
.Y(n_1006)
);

INVx1_ASAP7_75t_L g1007 ( 
.A(n_767),
.Y(n_1007)
);

NAND2xp5_ASAP7_75t_L g1008 ( 
.A(n_565),
.B(n_6),
.Y(n_1008)
);

INVx1_ASAP7_75t_L g1009 ( 
.A(n_767),
.Y(n_1009)
);

NOR2xp33_ASAP7_75t_L g1010 ( 
.A(n_599),
.B(n_7),
.Y(n_1010)
);

INVx1_ASAP7_75t_L g1011 ( 
.A(n_768),
.Y(n_1011)
);

INVx1_ASAP7_75t_L g1012 ( 
.A(n_768),
.Y(n_1012)
);

INVx1_ASAP7_75t_L g1013 ( 
.A(n_806),
.Y(n_1013)
);

INVxp67_ASAP7_75t_L g1014 ( 
.A(n_613),
.Y(n_1014)
);

CKINVDCx14_ASAP7_75t_R g1015 ( 
.A(n_717),
.Y(n_1015)
);

NOR2xp33_ASAP7_75t_L g1016 ( 
.A(n_608),
.B(n_7),
.Y(n_1016)
);

BUFx3_ASAP7_75t_L g1017 ( 
.A(n_693),
.Y(n_1017)
);

INVxp33_ASAP7_75t_SL g1018 ( 
.A(n_568),
.Y(n_1018)
);

NOR2xp33_ASAP7_75t_L g1019 ( 
.A(n_616),
.B(n_8),
.Y(n_1019)
);

CKINVDCx5p33_ASAP7_75t_R g1020 ( 
.A(n_570),
.Y(n_1020)
);

INVx1_ASAP7_75t_L g1021 ( 
.A(n_806),
.Y(n_1021)
);

INVx1_ASAP7_75t_L g1022 ( 
.A(n_854),
.Y(n_1022)
);

BUFx3_ASAP7_75t_L g1023 ( 
.A(n_693),
.Y(n_1023)
);

INVx1_ASAP7_75t_L g1024 ( 
.A(n_854),
.Y(n_1024)
);

INVx1_ASAP7_75t_L g1025 ( 
.A(n_888),
.Y(n_1025)
);

INVx1_ASAP7_75t_L g1026 ( 
.A(n_888),
.Y(n_1026)
);

CKINVDCx20_ASAP7_75t_R g1027 ( 
.A(n_911),
.Y(n_1027)
);

CKINVDCx20_ASAP7_75t_R g1028 ( 
.A(n_911),
.Y(n_1028)
);

CKINVDCx20_ASAP7_75t_R g1029 ( 
.A(n_568),
.Y(n_1029)
);

CKINVDCx5p33_ASAP7_75t_R g1030 ( 
.A(n_570),
.Y(n_1030)
);

CKINVDCx5p33_ASAP7_75t_R g1031 ( 
.A(n_571),
.Y(n_1031)
);

CKINVDCx5p33_ASAP7_75t_R g1032 ( 
.A(n_571),
.Y(n_1032)
);

CKINVDCx5p33_ASAP7_75t_R g1033 ( 
.A(n_572),
.Y(n_1033)
);

INVx1_ASAP7_75t_L g1034 ( 
.A(n_899),
.Y(n_1034)
);

NOR2xp33_ASAP7_75t_L g1035 ( 
.A(n_638),
.B(n_8),
.Y(n_1035)
);

NOR2xp67_ASAP7_75t_L g1036 ( 
.A(n_899),
.B(n_569),
.Y(n_1036)
);

CKINVDCx5p33_ASAP7_75t_R g1037 ( 
.A(n_572),
.Y(n_1037)
);

NOR2xp33_ASAP7_75t_L g1038 ( 
.A(n_645),
.B(n_9),
.Y(n_1038)
);

INVxp33_ASAP7_75t_SL g1039 ( 
.A(n_579),
.Y(n_1039)
);

INVx1_ASAP7_75t_L g1040 ( 
.A(n_746),
.Y(n_1040)
);

CKINVDCx5p33_ASAP7_75t_R g1041 ( 
.A(n_579),
.Y(n_1041)
);

CKINVDCx20_ASAP7_75t_R g1042 ( 
.A(n_908),
.Y(n_1042)
);

INVx1_ASAP7_75t_L g1043 ( 
.A(n_746),
.Y(n_1043)
);

INVx2_ASAP7_75t_L g1044 ( 
.A(n_991),
.Y(n_1044)
);

BUFx6f_ASAP7_75t_L g1045 ( 
.A(n_991),
.Y(n_1045)
);

INVx1_ASAP7_75t_L g1046 ( 
.A(n_917),
.Y(n_1046)
);

INVx1_ASAP7_75t_L g1047 ( 
.A(n_918),
.Y(n_1047)
);

INVx2_ASAP7_75t_L g1048 ( 
.A(n_1040),
.Y(n_1048)
);

NAND2xp5_ASAP7_75t_L g1049 ( 
.A(n_914),
.B(n_581),
.Y(n_1049)
);

AND2x4_ASAP7_75t_L g1050 ( 
.A(n_919),
.B(n_577),
.Y(n_1050)
);

INVx3_ASAP7_75t_L g1051 ( 
.A(n_1017),
.Y(n_1051)
);

INVx2_ASAP7_75t_L g1052 ( 
.A(n_1043),
.Y(n_1052)
);

INVx1_ASAP7_75t_L g1053 ( 
.A(n_925),
.Y(n_1053)
);

INVx2_ASAP7_75t_L g1054 ( 
.A(n_1023),
.Y(n_1054)
);

INVx3_ASAP7_75t_L g1055 ( 
.A(n_928),
.Y(n_1055)
);

INVx2_ASAP7_75t_L g1056 ( 
.A(n_1023),
.Y(n_1056)
);

BUFx6f_ASAP7_75t_L g1057 ( 
.A(n_983),
.Y(n_1057)
);

NAND2xp5_ASAP7_75t_SL g1058 ( 
.A(n_924),
.B(n_612),
.Y(n_1058)
);

INVx1_ASAP7_75t_L g1059 ( 
.A(n_929),
.Y(n_1059)
);

INVx1_ASAP7_75t_L g1060 ( 
.A(n_930),
.Y(n_1060)
);

INVx2_ASAP7_75t_L g1061 ( 
.A(n_990),
.Y(n_1061)
);

AND2x4_ASAP7_75t_L g1062 ( 
.A(n_931),
.B(n_580),
.Y(n_1062)
);

INVx2_ASAP7_75t_L g1063 ( 
.A(n_993),
.Y(n_1063)
);

NAND2xp5_ASAP7_75t_SL g1064 ( 
.A(n_936),
.B(n_612),
.Y(n_1064)
);

INVx1_ASAP7_75t_L g1065 ( 
.A(n_935),
.Y(n_1065)
);

INVx1_ASAP7_75t_L g1066 ( 
.A(n_946),
.Y(n_1066)
);

INVx2_ASAP7_75t_L g1067 ( 
.A(n_996),
.Y(n_1067)
);

AND2x2_ASAP7_75t_L g1068 ( 
.A(n_922),
.B(n_637),
.Y(n_1068)
);

INVx1_ASAP7_75t_L g1069 ( 
.A(n_948),
.Y(n_1069)
);

BUFx2_ASAP7_75t_L g1070 ( 
.A(n_966),
.Y(n_1070)
);

AND2x6_ASAP7_75t_L g1071 ( 
.A(n_940),
.B(n_634),
.Y(n_1071)
);

INVx1_ASAP7_75t_L g1072 ( 
.A(n_951),
.Y(n_1072)
);

BUFx2_ASAP7_75t_L g1073 ( 
.A(n_966),
.Y(n_1073)
);

INVx2_ASAP7_75t_L g1074 ( 
.A(n_1002),
.Y(n_1074)
);

AOI22xp5_ASAP7_75t_L g1075 ( 
.A1(n_923),
.A2(n_585),
.B1(n_587),
.B2(n_584),
.Y(n_1075)
);

INVx2_ASAP7_75t_L g1076 ( 
.A(n_1003),
.Y(n_1076)
);

INVx1_ASAP7_75t_L g1077 ( 
.A(n_955),
.Y(n_1077)
);

INVx1_ASAP7_75t_L g1078 ( 
.A(n_961),
.Y(n_1078)
);

BUFx6f_ASAP7_75t_L g1079 ( 
.A(n_1004),
.Y(n_1079)
);

INVx1_ASAP7_75t_L g1080 ( 
.A(n_967),
.Y(n_1080)
);

INVx1_ASAP7_75t_L g1081 ( 
.A(n_968),
.Y(n_1081)
);

INVx6_ASAP7_75t_L g1082 ( 
.A(n_942),
.Y(n_1082)
);

INVx1_ASAP7_75t_L g1083 ( 
.A(n_975),
.Y(n_1083)
);

INVx2_ASAP7_75t_L g1084 ( 
.A(n_1007),
.Y(n_1084)
);

INVx2_ASAP7_75t_L g1085 ( 
.A(n_1009),
.Y(n_1085)
);

INVx1_ASAP7_75t_L g1086 ( 
.A(n_978),
.Y(n_1086)
);

INVx2_ASAP7_75t_L g1087 ( 
.A(n_1011),
.Y(n_1087)
);

OA21x2_ASAP7_75t_L g1088 ( 
.A1(n_979),
.A2(n_750),
.B(n_634),
.Y(n_1088)
);

INVx2_ASAP7_75t_L g1089 ( 
.A(n_1012),
.Y(n_1089)
);

INVx2_ASAP7_75t_L g1090 ( 
.A(n_1013),
.Y(n_1090)
);

INVx3_ASAP7_75t_L g1091 ( 
.A(n_981),
.Y(n_1091)
);

INVx1_ASAP7_75t_L g1092 ( 
.A(n_953),
.Y(n_1092)
);

INVx1_ASAP7_75t_L g1093 ( 
.A(n_958),
.Y(n_1093)
);

INVx2_ASAP7_75t_L g1094 ( 
.A(n_1021),
.Y(n_1094)
);

INVx2_ASAP7_75t_L g1095 ( 
.A(n_1022),
.Y(n_1095)
);

CKINVDCx5p33_ASAP7_75t_R g1096 ( 
.A(n_923),
.Y(n_1096)
);

HB1xp67_ASAP7_75t_L g1097 ( 
.A(n_969),
.Y(n_1097)
);

HB1xp67_ASAP7_75t_L g1098 ( 
.A(n_980),
.Y(n_1098)
);

INVx2_ASAP7_75t_L g1099 ( 
.A(n_1024),
.Y(n_1099)
);

INVx3_ASAP7_75t_L g1100 ( 
.A(n_1025),
.Y(n_1100)
);

AND2x2_ASAP7_75t_L g1101 ( 
.A(n_927),
.B(n_637),
.Y(n_1101)
);

INVx1_ASAP7_75t_L g1102 ( 
.A(n_963),
.Y(n_1102)
);

INVx2_ASAP7_75t_L g1103 ( 
.A(n_1026),
.Y(n_1103)
);

INVx1_ASAP7_75t_L g1104 ( 
.A(n_965),
.Y(n_1104)
);

INVx2_ASAP7_75t_L g1105 ( 
.A(n_1034),
.Y(n_1105)
);

NAND2xp5_ASAP7_75t_L g1106 ( 
.A(n_1015),
.B(n_584),
.Y(n_1106)
);

INVx3_ASAP7_75t_L g1107 ( 
.A(n_985),
.Y(n_1107)
);

INVx2_ASAP7_75t_L g1108 ( 
.A(n_997),
.Y(n_1108)
);

OA21x2_ASAP7_75t_L g1109 ( 
.A1(n_999),
.A2(n_858),
.B(n_750),
.Y(n_1109)
);

NAND2xp5_ASAP7_75t_SL g1110 ( 
.A(n_947),
.B(n_858),
.Y(n_1110)
);

INVx2_ASAP7_75t_L g1111 ( 
.A(n_1005),
.Y(n_1111)
);

NAND2xp5_ASAP7_75t_L g1112 ( 
.A(n_973),
.B(n_1039),
.Y(n_1112)
);

OAI21x1_ASAP7_75t_L g1113 ( 
.A1(n_1006),
.A2(n_660),
.B(n_647),
.Y(n_1113)
);

AND2x4_ASAP7_75t_L g1114 ( 
.A(n_1036),
.B(n_588),
.Y(n_1114)
);

BUFx6f_ASAP7_75t_L g1115 ( 
.A(n_1010),
.Y(n_1115)
);

INVx2_ASAP7_75t_L g1116 ( 
.A(n_1016),
.Y(n_1116)
);

INVx2_ASAP7_75t_L g1117 ( 
.A(n_1019),
.Y(n_1117)
);

NAND2xp5_ASAP7_75t_L g1118 ( 
.A(n_973),
.B(n_585),
.Y(n_1118)
);

NAND2xp5_ASAP7_75t_SL g1119 ( 
.A(n_945),
.B(n_723),
.Y(n_1119)
);

INVx1_ASAP7_75t_L g1120 ( 
.A(n_1035),
.Y(n_1120)
);

INVx1_ASAP7_75t_L g1121 ( 
.A(n_1038),
.Y(n_1121)
);

BUFx6f_ASAP7_75t_L g1122 ( 
.A(n_1008),
.Y(n_1122)
);

INVx1_ASAP7_75t_L g1123 ( 
.A(n_939),
.Y(n_1123)
);

BUFx6f_ASAP7_75t_L g1124 ( 
.A(n_989),
.Y(n_1124)
);

INVx2_ASAP7_75t_L g1125 ( 
.A(n_1014),
.Y(n_1125)
);

INVx2_ASAP7_75t_L g1126 ( 
.A(n_992),
.Y(n_1126)
);

NOR2xp33_ASAP7_75t_L g1127 ( 
.A(n_1018),
.B(n_729),
.Y(n_1127)
);

AND2x2_ASAP7_75t_L g1128 ( 
.A(n_952),
.B(n_637),
.Y(n_1128)
);

INVx1_ASAP7_75t_L g1129 ( 
.A(n_994),
.Y(n_1129)
);

INVx1_ASAP7_75t_L g1130 ( 
.A(n_995),
.Y(n_1130)
);

INVx1_ASAP7_75t_L g1131 ( 
.A(n_998),
.Y(n_1131)
);

AND2x4_ASAP7_75t_L g1132 ( 
.A(n_1041),
.B(n_590),
.Y(n_1132)
);

NAND2xp5_ASAP7_75t_L g1133 ( 
.A(n_1018),
.B(n_587),
.Y(n_1133)
);

BUFx6f_ASAP7_75t_L g1134 ( 
.A(n_1000),
.Y(n_1134)
);

NOR2xp33_ASAP7_75t_L g1135 ( 
.A(n_1039),
.B(n_738),
.Y(n_1135)
);

AND2x2_ASAP7_75t_L g1136 ( 
.A(n_970),
.B(n_641),
.Y(n_1136)
);

INVx2_ASAP7_75t_L g1137 ( 
.A(n_1020),
.Y(n_1137)
);

BUFx6f_ASAP7_75t_L g1138 ( 
.A(n_1030),
.Y(n_1138)
);

INVx1_ASAP7_75t_L g1139 ( 
.A(n_1031),
.Y(n_1139)
);

NAND2xp5_ASAP7_75t_L g1140 ( 
.A(n_1032),
.B(n_595),
.Y(n_1140)
);

NAND2xp5_ASAP7_75t_L g1141 ( 
.A(n_1033),
.B(n_595),
.Y(n_1141)
);

HB1xp67_ASAP7_75t_L g1142 ( 
.A(n_1041),
.Y(n_1142)
);

BUFx6f_ASAP7_75t_L g1143 ( 
.A(n_1037),
.Y(n_1143)
);

INVx1_ASAP7_75t_L g1144 ( 
.A(n_916),
.Y(n_1144)
);

BUFx6f_ASAP7_75t_L g1145 ( 
.A(n_915),
.Y(n_1145)
);

NAND2xp5_ASAP7_75t_L g1146 ( 
.A(n_915),
.B(n_597),
.Y(n_1146)
);

INVx1_ASAP7_75t_L g1147 ( 
.A(n_938),
.Y(n_1147)
);

INVx1_ASAP7_75t_L g1148 ( 
.A(n_938),
.Y(n_1148)
);

INVx1_ASAP7_75t_L g1149 ( 
.A(n_1027),
.Y(n_1149)
);

INVx1_ASAP7_75t_L g1150 ( 
.A(n_1027),
.Y(n_1150)
);

INVx6_ASAP7_75t_L g1151 ( 
.A(n_1028),
.Y(n_1151)
);

INVx1_ASAP7_75t_L g1152 ( 
.A(n_1028),
.Y(n_1152)
);

AND2x4_ASAP7_75t_L g1153 ( 
.A(n_1029),
.B(n_592),
.Y(n_1153)
);

INVx4_ASAP7_75t_L g1154 ( 
.A(n_926),
.Y(n_1154)
);

NOR2xp33_ASAP7_75t_L g1155 ( 
.A(n_1029),
.B(n_788),
.Y(n_1155)
);

AND2x4_ASAP7_75t_L g1156 ( 
.A(n_1042),
.B(n_604),
.Y(n_1156)
);

INVx2_ASAP7_75t_L g1157 ( 
.A(n_1042),
.Y(n_1157)
);

INVx1_ASAP7_75t_L g1158 ( 
.A(n_932),
.Y(n_1158)
);

HB1xp67_ASAP7_75t_L g1159 ( 
.A(n_944),
.Y(n_1159)
);

XNOR2x2_ASAP7_75t_L g1160 ( 
.A(n_933),
.B(n_700),
.Y(n_1160)
);

BUFx6f_ASAP7_75t_L g1161 ( 
.A(n_956),
.Y(n_1161)
);

INVx1_ASAP7_75t_L g1162 ( 
.A(n_957),
.Y(n_1162)
);

INVx1_ASAP7_75t_L g1163 ( 
.A(n_962),
.Y(n_1163)
);

INVx1_ASAP7_75t_L g1164 ( 
.A(n_972),
.Y(n_1164)
);

INVxp67_ASAP7_75t_L g1165 ( 
.A(n_977),
.Y(n_1165)
);

INVx2_ASAP7_75t_L g1166 ( 
.A(n_913),
.Y(n_1166)
);

INVx1_ASAP7_75t_L g1167 ( 
.A(n_984),
.Y(n_1167)
);

INVx1_ASAP7_75t_L g1168 ( 
.A(n_986),
.Y(n_1168)
);

HB1xp67_ASAP7_75t_L g1169 ( 
.A(n_987),
.Y(n_1169)
);

NAND2xp5_ASAP7_75t_L g1170 ( 
.A(n_988),
.B(n_597),
.Y(n_1170)
);

INVx1_ASAP7_75t_L g1171 ( 
.A(n_913),
.Y(n_1171)
);

INVx1_ASAP7_75t_L g1172 ( 
.A(n_920),
.Y(n_1172)
);

HB1xp67_ASAP7_75t_L g1173 ( 
.A(n_920),
.Y(n_1173)
);

BUFx6f_ASAP7_75t_L g1174 ( 
.A(n_921),
.Y(n_1174)
);

INVx1_ASAP7_75t_L g1175 ( 
.A(n_921),
.Y(n_1175)
);

INVx1_ASAP7_75t_L g1176 ( 
.A(n_933),
.Y(n_1176)
);

AND2x4_ASAP7_75t_L g1177 ( 
.A(n_934),
.B(n_606),
.Y(n_1177)
);

INVx1_ASAP7_75t_L g1178 ( 
.A(n_934),
.Y(n_1178)
);

INVx1_ASAP7_75t_L g1179 ( 
.A(n_943),
.Y(n_1179)
);

INVx1_ASAP7_75t_L g1180 ( 
.A(n_943),
.Y(n_1180)
);

INVx2_ASAP7_75t_L g1181 ( 
.A(n_949),
.Y(n_1181)
);

BUFx6f_ASAP7_75t_L g1182 ( 
.A(n_949),
.Y(n_1182)
);

AND2x4_ASAP7_75t_L g1183 ( 
.A(n_950),
.B(n_607),
.Y(n_1183)
);

NOR2xp33_ASAP7_75t_SL g1184 ( 
.A(n_954),
.B(n_573),
.Y(n_1184)
);

OAI22xp5_ASAP7_75t_SL g1185 ( 
.A1(n_954),
.A2(n_908),
.B1(n_605),
.B2(n_609),
.Y(n_1185)
);

NAND2xp5_ASAP7_75t_L g1186 ( 
.A(n_959),
.B(n_598),
.Y(n_1186)
);

CKINVDCx5p33_ASAP7_75t_R g1187 ( 
.A(n_959),
.Y(n_1187)
);

NAND2xp5_ASAP7_75t_L g1188 ( 
.A(n_960),
.B(n_598),
.Y(n_1188)
);

INVx1_ASAP7_75t_L g1189 ( 
.A(n_960),
.Y(n_1189)
);

OA21x2_ASAP7_75t_L g1190 ( 
.A1(n_964),
.A2(n_823),
.B(n_812),
.Y(n_1190)
);

INVx4_ASAP7_75t_L g1191 ( 
.A(n_964),
.Y(n_1191)
);

NAND2xp5_ASAP7_75t_L g1192 ( 
.A(n_971),
.B(n_605),
.Y(n_1192)
);

INVx2_ASAP7_75t_L g1193 ( 
.A(n_971),
.Y(n_1193)
);

NOR2xp33_ASAP7_75t_L g1194 ( 
.A(n_974),
.B(n_824),
.Y(n_1194)
);

CKINVDCx8_ASAP7_75t_R g1195 ( 
.A(n_974),
.Y(n_1195)
);

HB1xp67_ASAP7_75t_L g1196 ( 
.A(n_1001),
.Y(n_1196)
);

INVx1_ASAP7_75t_L g1197 ( 
.A(n_976),
.Y(n_1197)
);

INVx2_ASAP7_75t_L g1198 ( 
.A(n_976),
.Y(n_1198)
);

INVx2_ASAP7_75t_L g1199 ( 
.A(n_982),
.Y(n_1199)
);

BUFx6f_ASAP7_75t_L g1200 ( 
.A(n_982),
.Y(n_1200)
);

INVx3_ASAP7_75t_L g1201 ( 
.A(n_1001),
.Y(n_1201)
);

INVx3_ASAP7_75t_L g1202 ( 
.A(n_1017),
.Y(n_1202)
);

INVx1_ASAP7_75t_L g1203 ( 
.A(n_917),
.Y(n_1203)
);

INVx1_ASAP7_75t_L g1204 ( 
.A(n_917),
.Y(n_1204)
);

BUFx6f_ASAP7_75t_L g1205 ( 
.A(n_991),
.Y(n_1205)
);

INVx2_ASAP7_75t_L g1206 ( 
.A(n_991),
.Y(n_1206)
);

HB1xp67_ASAP7_75t_L g1207 ( 
.A(n_941),
.Y(n_1207)
);

INVxp67_ASAP7_75t_L g1208 ( 
.A(n_941),
.Y(n_1208)
);

AND2x2_ASAP7_75t_L g1209 ( 
.A(n_937),
.B(n_641),
.Y(n_1209)
);

INVx2_ASAP7_75t_L g1210 ( 
.A(n_991),
.Y(n_1210)
);

NAND2xp5_ASAP7_75t_L g1211 ( 
.A(n_914),
.B(n_609),
.Y(n_1211)
);

NAND2xp5_ASAP7_75t_L g1212 ( 
.A(n_914),
.B(n_611),
.Y(n_1212)
);

HB1xp67_ASAP7_75t_L g1213 ( 
.A(n_941),
.Y(n_1213)
);

INVx1_ASAP7_75t_L g1214 ( 
.A(n_917),
.Y(n_1214)
);

INVx1_ASAP7_75t_L g1215 ( 
.A(n_917),
.Y(n_1215)
);

AND2x4_ASAP7_75t_L g1216 ( 
.A(n_917),
.B(n_610),
.Y(n_1216)
);

BUFx6f_ASAP7_75t_L g1217 ( 
.A(n_991),
.Y(n_1217)
);

INVx2_ASAP7_75t_L g1218 ( 
.A(n_991),
.Y(n_1218)
);

INVx1_ASAP7_75t_L g1219 ( 
.A(n_917),
.Y(n_1219)
);

INVx3_ASAP7_75t_L g1220 ( 
.A(n_1017),
.Y(n_1220)
);

BUFx6f_ASAP7_75t_L g1221 ( 
.A(n_991),
.Y(n_1221)
);

BUFx2_ASAP7_75t_L g1222 ( 
.A(n_966),
.Y(n_1222)
);

NAND2xp33_ASAP7_75t_SL g1223 ( 
.A(n_985),
.B(n_573),
.Y(n_1223)
);

NAND2xp5_ASAP7_75t_SL g1224 ( 
.A(n_1040),
.B(n_827),
.Y(n_1224)
);

INVx1_ASAP7_75t_L g1225 ( 
.A(n_917),
.Y(n_1225)
);

INVx1_ASAP7_75t_L g1226 ( 
.A(n_917),
.Y(n_1226)
);

INVx1_ASAP7_75t_L g1227 ( 
.A(n_917),
.Y(n_1227)
);

AND2x2_ASAP7_75t_L g1228 ( 
.A(n_937),
.B(n_657),
.Y(n_1228)
);

BUFx6f_ASAP7_75t_L g1229 ( 
.A(n_991),
.Y(n_1229)
);

NAND2xp5_ASAP7_75t_L g1230 ( 
.A(n_914),
.B(n_618),
.Y(n_1230)
);

INVx2_ASAP7_75t_L g1231 ( 
.A(n_991),
.Y(n_1231)
);

INVx1_ASAP7_75t_L g1232 ( 
.A(n_917),
.Y(n_1232)
);

AND2x4_ASAP7_75t_L g1233 ( 
.A(n_917),
.B(n_621),
.Y(n_1233)
);

INVx3_ASAP7_75t_L g1234 ( 
.A(n_917),
.Y(n_1234)
);

INVxp67_ASAP7_75t_L g1235 ( 
.A(n_941),
.Y(n_1235)
);

OAI21x1_ASAP7_75t_L g1236 ( 
.A1(n_991),
.A2(n_848),
.B(n_836),
.Y(n_1236)
);

INVx1_ASAP7_75t_L g1237 ( 
.A(n_917),
.Y(n_1237)
);

INVx1_ASAP7_75t_L g1238 ( 
.A(n_917),
.Y(n_1238)
);

INVx1_ASAP7_75t_L g1239 ( 
.A(n_917),
.Y(n_1239)
);

INVx1_ASAP7_75t_L g1240 ( 
.A(n_917),
.Y(n_1240)
);

INVx1_ASAP7_75t_L g1241 ( 
.A(n_917),
.Y(n_1241)
);

INVx2_ASAP7_75t_L g1242 ( 
.A(n_991),
.Y(n_1242)
);

NAND2xp5_ASAP7_75t_L g1243 ( 
.A(n_914),
.B(n_618),
.Y(n_1243)
);

INVx2_ASAP7_75t_L g1244 ( 
.A(n_991),
.Y(n_1244)
);

NAND2xp33_ASAP7_75t_L g1245 ( 
.A(n_915),
.B(n_746),
.Y(n_1245)
);

OAI21x1_ASAP7_75t_L g1246 ( 
.A1(n_991),
.A2(n_885),
.B(n_849),
.Y(n_1246)
);

INVx2_ASAP7_75t_L g1247 ( 
.A(n_991),
.Y(n_1247)
);

INVx2_ASAP7_75t_L g1248 ( 
.A(n_1236),
.Y(n_1248)
);

INVx1_ASAP7_75t_L g1249 ( 
.A(n_1055),
.Y(n_1249)
);

NOR2xp33_ASAP7_75t_L g1250 ( 
.A(n_1092),
.B(n_717),
.Y(n_1250)
);

INVx2_ASAP7_75t_L g1251 ( 
.A(n_1236),
.Y(n_1251)
);

NAND3xp33_ASAP7_75t_L g1252 ( 
.A(n_1075),
.B(n_625),
.C(n_619),
.Y(n_1252)
);

OAI22xp5_ASAP7_75t_L g1253 ( 
.A1(n_1112),
.A2(n_625),
.B1(n_629),
.B2(n_619),
.Y(n_1253)
);

NOR2xp33_ASAP7_75t_L g1254 ( 
.A(n_1093),
.B(n_717),
.Y(n_1254)
);

INVx1_ASAP7_75t_L g1255 ( 
.A(n_1055),
.Y(n_1255)
);

AND2x2_ASAP7_75t_L g1256 ( 
.A(n_1209),
.B(n_657),
.Y(n_1256)
);

NAND2xp5_ASAP7_75t_L g1257 ( 
.A(n_1102),
.B(n_574),
.Y(n_1257)
);

NAND2xp5_ASAP7_75t_SL g1258 ( 
.A(n_1122),
.B(n_898),
.Y(n_1258)
);

NAND2xp5_ASAP7_75t_L g1259 ( 
.A(n_1104),
.B(n_574),
.Y(n_1259)
);

BUFx2_ASAP7_75t_L g1260 ( 
.A(n_1096),
.Y(n_1260)
);

INVx1_ASAP7_75t_SL g1261 ( 
.A(n_1082),
.Y(n_1261)
);

INVx1_ASAP7_75t_L g1262 ( 
.A(n_1234),
.Y(n_1262)
);

BUFx2_ASAP7_75t_L g1263 ( 
.A(n_1096),
.Y(n_1263)
);

INVxp33_ASAP7_75t_L g1264 ( 
.A(n_1097),
.Y(n_1264)
);

NAND2xp5_ASAP7_75t_SL g1265 ( 
.A(n_1122),
.B(n_1115),
.Y(n_1265)
);

CKINVDCx5p33_ASAP7_75t_R g1266 ( 
.A(n_1187),
.Y(n_1266)
);

NAND2xp5_ASAP7_75t_SL g1267 ( 
.A(n_1122),
.B(n_886),
.Y(n_1267)
);

NAND2xp5_ASAP7_75t_L g1268 ( 
.A(n_1120),
.B(n_578),
.Y(n_1268)
);

BUFx10_ASAP7_75t_L g1269 ( 
.A(n_1082),
.Y(n_1269)
);

INVx2_ASAP7_75t_SL g1270 ( 
.A(n_1082),
.Y(n_1270)
);

AOI22xp5_ASAP7_75t_L g1271 ( 
.A1(n_1132),
.A2(n_734),
.B1(n_735),
.B2(n_629),
.Y(n_1271)
);

NAND2xp5_ASAP7_75t_SL g1272 ( 
.A(n_1122),
.B(n_726),
.Y(n_1272)
);

NOR2xp33_ASAP7_75t_L g1273 ( 
.A(n_1125),
.B(n_1123),
.Y(n_1273)
);

OR2x2_ASAP7_75t_L g1274 ( 
.A(n_1186),
.B(n_734),
.Y(n_1274)
);

NAND2xp5_ASAP7_75t_SL g1275 ( 
.A(n_1115),
.B(n_1113),
.Y(n_1275)
);

AND3x1_ASAP7_75t_L g1276 ( 
.A(n_1184),
.B(n_628),
.C(n_623),
.Y(n_1276)
);

NAND2xp5_ASAP7_75t_L g1277 ( 
.A(n_1121),
.B(n_589),
.Y(n_1277)
);

NAND2xp5_ASAP7_75t_SL g1278 ( 
.A(n_1115),
.B(n_726),
.Y(n_1278)
);

OAI22xp5_ASAP7_75t_L g1279 ( 
.A1(n_1049),
.A2(n_840),
.B1(n_850),
.B2(n_735),
.Y(n_1279)
);

AND2x6_ASAP7_75t_L g1280 ( 
.A(n_1128),
.B(n_726),
.Y(n_1280)
);

INVx1_ASAP7_75t_L g1281 ( 
.A(n_1234),
.Y(n_1281)
);

INVx1_ASAP7_75t_L g1282 ( 
.A(n_1046),
.Y(n_1282)
);

AOI22xp33_ASAP7_75t_L g1283 ( 
.A1(n_1108),
.A2(n_746),
.B1(n_642),
.B2(n_644),
.Y(n_1283)
);

NAND2xp33_ASAP7_75t_L g1284 ( 
.A(n_1071),
.B(n_746),
.Y(n_1284)
);

INVx1_ASAP7_75t_L g1285 ( 
.A(n_1047),
.Y(n_1285)
);

BUFx3_ASAP7_75t_L g1286 ( 
.A(n_1051),
.Y(n_1286)
);

BUFx6f_ASAP7_75t_L g1287 ( 
.A(n_1246),
.Y(n_1287)
);

BUFx6f_ASAP7_75t_SL g1288 ( 
.A(n_1191),
.Y(n_1288)
);

INVx2_ASAP7_75t_SL g1289 ( 
.A(n_1228),
.Y(n_1289)
);

INVx4_ASAP7_75t_L g1290 ( 
.A(n_1051),
.Y(n_1290)
);

AOI22xp33_ASAP7_75t_L g1291 ( 
.A1(n_1108),
.A2(n_746),
.B1(n_646),
.B2(n_652),
.Y(n_1291)
);

INVx2_ASAP7_75t_L g1292 ( 
.A(n_1051),
.Y(n_1292)
);

CKINVDCx5p33_ASAP7_75t_R g1293 ( 
.A(n_1187),
.Y(n_1293)
);

OR2x2_ASAP7_75t_L g1294 ( 
.A(n_1188),
.B(n_840),
.Y(n_1294)
);

INVx2_ASAP7_75t_L g1295 ( 
.A(n_1202),
.Y(n_1295)
);

NOR2xp33_ASAP7_75t_L g1296 ( 
.A(n_1125),
.B(n_589),
.Y(n_1296)
);

BUFx3_ASAP7_75t_L g1297 ( 
.A(n_1202),
.Y(n_1297)
);

INVx1_ASAP7_75t_L g1298 ( 
.A(n_1053),
.Y(n_1298)
);

BUFx2_ASAP7_75t_L g1299 ( 
.A(n_1070),
.Y(n_1299)
);

NOR2xp33_ASAP7_75t_L g1300 ( 
.A(n_1111),
.B(n_591),
.Y(n_1300)
);

CKINVDCx20_ASAP7_75t_R g1301 ( 
.A(n_1185),
.Y(n_1301)
);

OAI22x1_ASAP7_75t_L g1302 ( 
.A1(n_1191),
.A2(n_851),
.B1(n_856),
.B2(n_850),
.Y(n_1302)
);

INVxp67_ASAP7_75t_L g1303 ( 
.A(n_1097),
.Y(n_1303)
);

AND2x6_ASAP7_75t_L g1304 ( 
.A(n_1136),
.B(n_726),
.Y(n_1304)
);

INVx2_ASAP7_75t_L g1305 ( 
.A(n_1202),
.Y(n_1305)
);

INVx2_ASAP7_75t_L g1306 ( 
.A(n_1220),
.Y(n_1306)
);

NAND2xp5_ASAP7_75t_L g1307 ( 
.A(n_1111),
.B(n_591),
.Y(n_1307)
);

INVx3_ASAP7_75t_L g1308 ( 
.A(n_1057),
.Y(n_1308)
);

NOR2xp33_ASAP7_75t_L g1309 ( 
.A(n_1116),
.B(n_602),
.Y(n_1309)
);

INVx2_ASAP7_75t_SL g1310 ( 
.A(n_1098),
.Y(n_1310)
);

NOR2xp33_ASAP7_75t_L g1311 ( 
.A(n_1116),
.B(n_602),
.Y(n_1311)
);

NOR2xp33_ASAP7_75t_L g1312 ( 
.A(n_1117),
.B(n_603),
.Y(n_1312)
);

NAND2xp5_ASAP7_75t_L g1313 ( 
.A(n_1117),
.B(n_603),
.Y(n_1313)
);

INVx1_ASAP7_75t_L g1314 ( 
.A(n_1059),
.Y(n_1314)
);

INVx2_ASAP7_75t_L g1315 ( 
.A(n_1220),
.Y(n_1315)
);

INVx1_ASAP7_75t_L g1316 ( 
.A(n_1060),
.Y(n_1316)
);

INVx2_ASAP7_75t_L g1317 ( 
.A(n_1220),
.Y(n_1317)
);

AND2x2_ASAP7_75t_L g1318 ( 
.A(n_1098),
.B(n_671),
.Y(n_1318)
);

INVx2_ASAP7_75t_L g1319 ( 
.A(n_1088),
.Y(n_1319)
);

INVx2_ASAP7_75t_L g1320 ( 
.A(n_1088),
.Y(n_1320)
);

NOR2x1p5_ASAP7_75t_L g1321 ( 
.A(n_1154),
.B(n_851),
.Y(n_1321)
);

INVx2_ASAP7_75t_L g1322 ( 
.A(n_1054),
.Y(n_1322)
);

INVxp67_ASAP7_75t_SL g1323 ( 
.A(n_1088),
.Y(n_1323)
);

INVx5_ASAP7_75t_L g1324 ( 
.A(n_1045),
.Y(n_1324)
);

INVx2_ASAP7_75t_L g1325 ( 
.A(n_1054),
.Y(n_1325)
);

AOI22xp33_ASAP7_75t_L g1326 ( 
.A1(n_1109),
.A2(n_653),
.B1(n_655),
.B2(n_630),
.Y(n_1326)
);

INVx1_ASAP7_75t_L g1327 ( 
.A(n_1065),
.Y(n_1327)
);

AOI22xp33_ASAP7_75t_L g1328 ( 
.A1(n_1109),
.A2(n_661),
.B1(n_670),
.B2(n_658),
.Y(n_1328)
);

NOR2xp33_ASAP7_75t_L g1329 ( 
.A(n_1127),
.B(n_614),
.Y(n_1329)
);

INVx2_ASAP7_75t_L g1330 ( 
.A(n_1056),
.Y(n_1330)
);

INVx1_ASAP7_75t_L g1331 ( 
.A(n_1066),
.Y(n_1331)
);

INVx1_ASAP7_75t_L g1332 ( 
.A(n_1203),
.Y(n_1332)
);

NAND2xp5_ASAP7_75t_L g1333 ( 
.A(n_1050),
.B(n_1062),
.Y(n_1333)
);

AOI22xp5_ASAP7_75t_L g1334 ( 
.A1(n_1132),
.A2(n_865),
.B1(n_867),
.B2(n_856),
.Y(n_1334)
);

INVx4_ASAP7_75t_L g1335 ( 
.A(n_1145),
.Y(n_1335)
);

AOI22xp33_ASAP7_75t_L g1336 ( 
.A1(n_1109),
.A2(n_1071),
.B1(n_1061),
.B2(n_1067),
.Y(n_1336)
);

NAND2xp5_ASAP7_75t_L g1337 ( 
.A(n_1050),
.B(n_614),
.Y(n_1337)
);

INVx1_ASAP7_75t_L g1338 ( 
.A(n_1204),
.Y(n_1338)
);

NOR2xp33_ASAP7_75t_L g1339 ( 
.A(n_1127),
.B(n_615),
.Y(n_1339)
);

INVx1_ASAP7_75t_L g1340 ( 
.A(n_1214),
.Y(n_1340)
);

AO21x2_ASAP7_75t_L g1341 ( 
.A1(n_1113),
.A2(n_1224),
.B(n_1064),
.Y(n_1341)
);

INVx1_ASAP7_75t_SL g1342 ( 
.A(n_1073),
.Y(n_1342)
);

HB1xp67_ASAP7_75t_L g1343 ( 
.A(n_1207),
.Y(n_1343)
);

INVx1_ASAP7_75t_L g1344 ( 
.A(n_1215),
.Y(n_1344)
);

INVx5_ASAP7_75t_L g1345 ( 
.A(n_1045),
.Y(n_1345)
);

AO22x2_ASAP7_75t_L g1346 ( 
.A1(n_1153),
.A2(n_843),
.B1(n_696),
.B2(n_675),
.Y(n_1346)
);

NAND2xp5_ASAP7_75t_L g1347 ( 
.A(n_1050),
.B(n_615),
.Y(n_1347)
);

INVx1_ASAP7_75t_L g1348 ( 
.A(n_1219),
.Y(n_1348)
);

NOR2xp33_ASAP7_75t_L g1349 ( 
.A(n_1135),
.B(n_620),
.Y(n_1349)
);

OR2x6_ASAP7_75t_L g1350 ( 
.A(n_1154),
.B(n_672),
.Y(n_1350)
);

NAND2xp5_ASAP7_75t_SL g1351 ( 
.A(n_1115),
.B(n_726),
.Y(n_1351)
);

NAND2xp5_ASAP7_75t_L g1352 ( 
.A(n_1062),
.B(n_1216),
.Y(n_1352)
);

NOR2xp33_ASAP7_75t_L g1353 ( 
.A(n_1135),
.B(n_620),
.Y(n_1353)
);

BUFx4f_ASAP7_75t_L g1354 ( 
.A(n_1145),
.Y(n_1354)
);

OR2x2_ASAP7_75t_L g1355 ( 
.A(n_1192),
.B(n_865),
.Y(n_1355)
);

AND2x4_ASAP7_75t_L g1356 ( 
.A(n_1126),
.B(n_1137),
.Y(n_1356)
);

NAND2xp5_ASAP7_75t_L g1357 ( 
.A(n_1062),
.B(n_622),
.Y(n_1357)
);

INVx1_ASAP7_75t_L g1358 ( 
.A(n_1225),
.Y(n_1358)
);

NAND2xp5_ASAP7_75t_L g1359 ( 
.A(n_1216),
.B(n_622),
.Y(n_1359)
);

NAND2xp5_ASAP7_75t_SL g1360 ( 
.A(n_1048),
.B(n_847),
.Y(n_1360)
);

NOR2xp33_ASAP7_75t_L g1361 ( 
.A(n_1216),
.B(n_627),
.Y(n_1361)
);

INVx1_ASAP7_75t_L g1362 ( 
.A(n_1226),
.Y(n_1362)
);

NOR2xp33_ASAP7_75t_L g1363 ( 
.A(n_1233),
.B(n_627),
.Y(n_1363)
);

INVx3_ASAP7_75t_L g1364 ( 
.A(n_1079),
.Y(n_1364)
);

BUFx4f_ASAP7_75t_L g1365 ( 
.A(n_1145),
.Y(n_1365)
);

BUFx4f_ASAP7_75t_L g1366 ( 
.A(n_1145),
.Y(n_1366)
);

AOI22xp33_ASAP7_75t_L g1367 ( 
.A1(n_1071),
.A2(n_678),
.B1(n_680),
.B2(n_679),
.Y(n_1367)
);

AND2x6_ASAP7_75t_L g1368 ( 
.A(n_1132),
.B(n_847),
.Y(n_1368)
);

INVx2_ASAP7_75t_L g1369 ( 
.A(n_1079),
.Y(n_1369)
);

NAND2xp5_ASAP7_75t_L g1370 ( 
.A(n_1233),
.B(n_732),
.Y(n_1370)
);

INVx3_ASAP7_75t_L g1371 ( 
.A(n_1079),
.Y(n_1371)
);

NAND2xp5_ASAP7_75t_L g1372 ( 
.A(n_1233),
.B(n_732),
.Y(n_1372)
);

BUFx3_ASAP7_75t_L g1373 ( 
.A(n_1071),
.Y(n_1373)
);

INVxp67_ASAP7_75t_SL g1374 ( 
.A(n_1107),
.Y(n_1374)
);

INVx5_ASAP7_75t_L g1375 ( 
.A(n_1045),
.Y(n_1375)
);

INVx1_ASAP7_75t_L g1376 ( 
.A(n_1227),
.Y(n_1376)
);

OAI22xp5_ASAP7_75t_L g1377 ( 
.A1(n_1211),
.A2(n_875),
.B1(n_880),
.B2(n_869),
.Y(n_1377)
);

NAND3xp33_ASAP7_75t_L g1378 ( 
.A(n_1155),
.B(n_881),
.C(n_880),
.Y(n_1378)
);

INVx2_ASAP7_75t_L g1379 ( 
.A(n_1061),
.Y(n_1379)
);

INVx1_ASAP7_75t_SL g1380 ( 
.A(n_1222),
.Y(n_1380)
);

INVx4_ASAP7_75t_L g1381 ( 
.A(n_1124),
.Y(n_1381)
);

INVx2_ASAP7_75t_L g1382 ( 
.A(n_1063),
.Y(n_1382)
);

BUFx10_ASAP7_75t_L g1383 ( 
.A(n_1155),
.Y(n_1383)
);

CKINVDCx8_ASAP7_75t_R g1384 ( 
.A(n_1182),
.Y(n_1384)
);

NOR2xp33_ASAP7_75t_L g1385 ( 
.A(n_1212),
.B(n_852),
.Y(n_1385)
);

INVx4_ASAP7_75t_L g1386 ( 
.A(n_1124),
.Y(n_1386)
);

NAND2xp5_ASAP7_75t_SL g1387 ( 
.A(n_1048),
.B(n_847),
.Y(n_1387)
);

INVx2_ASAP7_75t_L g1388 ( 
.A(n_1063),
.Y(n_1388)
);

AND2x2_ASAP7_75t_L g1389 ( 
.A(n_1207),
.B(n_671),
.Y(n_1389)
);

AND2x2_ASAP7_75t_L g1390 ( 
.A(n_1213),
.B(n_671),
.Y(n_1390)
);

CKINVDCx11_ASAP7_75t_R g1391 ( 
.A(n_1195),
.Y(n_1391)
);

INVx4_ASAP7_75t_L g1392 ( 
.A(n_1124),
.Y(n_1392)
);

AND2x6_ASAP7_75t_L g1393 ( 
.A(n_1126),
.B(n_847),
.Y(n_1393)
);

NAND2xp5_ASAP7_75t_L g1394 ( 
.A(n_1071),
.B(n_857),
.Y(n_1394)
);

INVx2_ASAP7_75t_SL g1395 ( 
.A(n_1213),
.Y(n_1395)
);

AND2x2_ASAP7_75t_L g1396 ( 
.A(n_1068),
.B(n_845),
.Y(n_1396)
);

AND2x2_ASAP7_75t_L g1397 ( 
.A(n_1101),
.B(n_845),
.Y(n_1397)
);

BUFx10_ASAP7_75t_L g1398 ( 
.A(n_1124),
.Y(n_1398)
);

INVx1_ASAP7_75t_L g1399 ( 
.A(n_1232),
.Y(n_1399)
);

INVx5_ASAP7_75t_L g1400 ( 
.A(n_1045),
.Y(n_1400)
);

HB1xp67_ASAP7_75t_L g1401 ( 
.A(n_1142),
.Y(n_1401)
);

OR2x6_ASAP7_75t_L g1402 ( 
.A(n_1154),
.B(n_681),
.Y(n_1402)
);

NOR2xp33_ASAP7_75t_L g1403 ( 
.A(n_1230),
.B(n_860),
.Y(n_1403)
);

NAND2xp33_ASAP7_75t_L g1404 ( 
.A(n_1137),
.B(n_866),
.Y(n_1404)
);

AND2x6_ASAP7_75t_L g1405 ( 
.A(n_1134),
.B(n_847),
.Y(n_1405)
);

AOI22xp5_ASAP7_75t_L g1406 ( 
.A1(n_1223),
.A2(n_889),
.B1(n_892),
.B2(n_882),
.Y(n_1406)
);

INVx2_ASAP7_75t_SL g1407 ( 
.A(n_1118),
.Y(n_1407)
);

INVx2_ASAP7_75t_L g1408 ( 
.A(n_1067),
.Y(n_1408)
);

NOR2x1p5_ASAP7_75t_L g1409 ( 
.A(n_1201),
.B(n_882),
.Y(n_1409)
);

CKINVDCx5p33_ASAP7_75t_R g1410 ( 
.A(n_1195),
.Y(n_1410)
);

INVx2_ASAP7_75t_L g1411 ( 
.A(n_1074),
.Y(n_1411)
);

INVx2_ASAP7_75t_L g1412 ( 
.A(n_1074),
.Y(n_1412)
);

NOR2xp33_ASAP7_75t_L g1413 ( 
.A(n_1243),
.B(n_866),
.Y(n_1413)
);

BUFx3_ASAP7_75t_L g1414 ( 
.A(n_1134),
.Y(n_1414)
);

BUFx2_ASAP7_75t_L g1415 ( 
.A(n_1142),
.Y(n_1415)
);

NAND2xp5_ASAP7_75t_SL g1416 ( 
.A(n_1052),
.B(n_871),
.Y(n_1416)
);

OR2x6_ASAP7_75t_L g1417 ( 
.A(n_1161),
.B(n_682),
.Y(n_1417)
);

NAND2xp5_ASAP7_75t_L g1418 ( 
.A(n_1100),
.B(n_1237),
.Y(n_1418)
);

INVx1_ASAP7_75t_L g1419 ( 
.A(n_1238),
.Y(n_1419)
);

BUFx6f_ASAP7_75t_L g1420 ( 
.A(n_1205),
.Y(n_1420)
);

INVx3_ASAP7_75t_L g1421 ( 
.A(n_1100),
.Y(n_1421)
);

INVxp67_ASAP7_75t_SL g1422 ( 
.A(n_1076),
.Y(n_1422)
);

BUFx6f_ASAP7_75t_L g1423 ( 
.A(n_1205),
.Y(n_1423)
);

BUFx3_ASAP7_75t_L g1424 ( 
.A(n_1134),
.Y(n_1424)
);

INVx2_ASAP7_75t_L g1425 ( 
.A(n_1076),
.Y(n_1425)
);

OR2x2_ASAP7_75t_L g1426 ( 
.A(n_1208),
.B(n_889),
.Y(n_1426)
);

INVx4_ASAP7_75t_SL g1427 ( 
.A(n_1134),
.Y(n_1427)
);

INVx1_ASAP7_75t_L g1428 ( 
.A(n_1239),
.Y(n_1428)
);

INVx1_ASAP7_75t_L g1429 ( 
.A(n_1240),
.Y(n_1429)
);

BUFx6f_ASAP7_75t_L g1430 ( 
.A(n_1205),
.Y(n_1430)
);

INVx1_ASAP7_75t_L g1431 ( 
.A(n_1241),
.Y(n_1431)
);

AND2x2_ASAP7_75t_L g1432 ( 
.A(n_1235),
.B(n_1133),
.Y(n_1432)
);

INVx3_ASAP7_75t_L g1433 ( 
.A(n_1091),
.Y(n_1433)
);

INVx4_ASAP7_75t_L g1434 ( 
.A(n_1138),
.Y(n_1434)
);

OR2x2_ASAP7_75t_L g1435 ( 
.A(n_1159),
.B(n_1169),
.Y(n_1435)
);

INVx3_ASAP7_75t_L g1436 ( 
.A(n_1091),
.Y(n_1436)
);

AOI22xp33_ASAP7_75t_L g1437 ( 
.A1(n_1084),
.A2(n_689),
.B1(n_692),
.B2(n_684),
.Y(n_1437)
);

NAND2xp5_ASAP7_75t_L g1438 ( 
.A(n_1058),
.B(n_871),
.Y(n_1438)
);

AND2x4_ASAP7_75t_L g1439 ( 
.A(n_1129),
.B(n_695),
.Y(n_1439)
);

NOR2x1p5_ASAP7_75t_L g1440 ( 
.A(n_1201),
.B(n_892),
.Y(n_1440)
);

INVx1_ASAP7_75t_SL g1441 ( 
.A(n_1151),
.Y(n_1441)
);

NOR2xp33_ASAP7_75t_L g1442 ( 
.A(n_1119),
.B(n_873),
.Y(n_1442)
);

INVx2_ASAP7_75t_L g1443 ( 
.A(n_1084),
.Y(n_1443)
);

INVxp33_ASAP7_75t_L g1444 ( 
.A(n_1194),
.Y(n_1444)
);

NAND3xp33_ASAP7_75t_L g1445 ( 
.A(n_1140),
.B(n_903),
.C(n_895),
.Y(n_1445)
);

NAND2xp5_ASAP7_75t_SL g1446 ( 
.A(n_1052),
.B(n_877),
.Y(n_1446)
);

BUFx6f_ASAP7_75t_L g1447 ( 
.A(n_1205),
.Y(n_1447)
);

INVx1_ASAP7_75t_L g1448 ( 
.A(n_1085),
.Y(n_1448)
);

BUFx6f_ASAP7_75t_L g1449 ( 
.A(n_1217),
.Y(n_1449)
);

NAND2xp5_ASAP7_75t_L g1450 ( 
.A(n_1069),
.B(n_879),
.Y(n_1450)
);

NAND3xp33_ASAP7_75t_L g1451 ( 
.A(n_1141),
.B(n_903),
.C(n_895),
.Y(n_1451)
);

AND2x4_ASAP7_75t_L g1452 ( 
.A(n_1130),
.B(n_697),
.Y(n_1452)
);

INVx1_ASAP7_75t_L g1453 ( 
.A(n_1087),
.Y(n_1453)
);

INVx1_ASAP7_75t_L g1454 ( 
.A(n_1087),
.Y(n_1454)
);

NAND2xp5_ASAP7_75t_SL g1455 ( 
.A(n_1217),
.B(n_896),
.Y(n_1455)
);

AND2x2_ASAP7_75t_SL g1456 ( 
.A(n_1190),
.B(n_685),
.Y(n_1456)
);

INVxp67_ASAP7_75t_L g1457 ( 
.A(n_1223),
.Y(n_1457)
);

INVx2_ASAP7_75t_L g1458 ( 
.A(n_1089),
.Y(n_1458)
);

AOI22xp33_ASAP7_75t_L g1459 ( 
.A1(n_1090),
.A2(n_698),
.B1(n_718),
.B2(n_705),
.Y(n_1459)
);

INVx1_ASAP7_75t_L g1460 ( 
.A(n_1090),
.Y(n_1460)
);

NOR3xp33_ASAP7_75t_L g1461 ( 
.A(n_1194),
.B(n_712),
.C(n_708),
.Y(n_1461)
);

INVx1_ASAP7_75t_L g1462 ( 
.A(n_1094),
.Y(n_1462)
);

INVx1_ASAP7_75t_L g1463 ( 
.A(n_1094),
.Y(n_1463)
);

AND2x2_ASAP7_75t_SL g1464 ( 
.A(n_1190),
.B(n_1245),
.Y(n_1464)
);

INVx1_ASAP7_75t_L g1465 ( 
.A(n_1095),
.Y(n_1465)
);

NOR2xp33_ASAP7_75t_SL g1466 ( 
.A(n_1165),
.B(n_904),
.Y(n_1466)
);

INVx1_ASAP7_75t_L g1467 ( 
.A(n_1095),
.Y(n_1467)
);

INVx2_ASAP7_75t_SL g1468 ( 
.A(n_1106),
.Y(n_1468)
);

INVx4_ASAP7_75t_L g1469 ( 
.A(n_1138),
.Y(n_1469)
);

INVx3_ASAP7_75t_L g1470 ( 
.A(n_1099),
.Y(n_1470)
);

NAND3xp33_ASAP7_75t_L g1471 ( 
.A(n_1146),
.B(n_906),
.C(n_904),
.Y(n_1471)
);

INVx2_ASAP7_75t_SL g1472 ( 
.A(n_1138),
.Y(n_1472)
);

BUFx10_ASAP7_75t_L g1473 ( 
.A(n_1138),
.Y(n_1473)
);

INVx4_ASAP7_75t_L g1474 ( 
.A(n_1143),
.Y(n_1474)
);

NAND2xp5_ASAP7_75t_L g1475 ( 
.A(n_1072),
.B(n_901),
.Y(n_1475)
);

INVx2_ASAP7_75t_L g1476 ( 
.A(n_1103),
.Y(n_1476)
);

NAND2xp5_ASAP7_75t_SL g1477 ( 
.A(n_1217),
.B(n_901),
.Y(n_1477)
);

AOI22xp5_ASAP7_75t_L g1478 ( 
.A1(n_1147),
.A2(n_906),
.B1(n_633),
.B2(n_639),
.Y(n_1478)
);

INVx4_ASAP7_75t_L g1479 ( 
.A(n_1143),
.Y(n_1479)
);

NOR2x1p5_ASAP7_75t_L g1480 ( 
.A(n_1201),
.B(n_632),
.Y(n_1480)
);

INVx1_ASAP7_75t_L g1481 ( 
.A(n_1103),
.Y(n_1481)
);

INVx2_ASAP7_75t_L g1482 ( 
.A(n_1105),
.Y(n_1482)
);

NAND2xp5_ASAP7_75t_L g1483 ( 
.A(n_1077),
.B(n_902),
.Y(n_1483)
);

INVx2_ASAP7_75t_L g1484 ( 
.A(n_1105),
.Y(n_1484)
);

NAND2xp5_ASAP7_75t_SL g1485 ( 
.A(n_1221),
.B(n_1229),
.Y(n_1485)
);

CKINVDCx20_ASAP7_75t_R g1486 ( 
.A(n_1151),
.Y(n_1486)
);

AOI22xp33_ASAP7_75t_L g1487 ( 
.A1(n_1078),
.A2(n_721),
.B1(n_730),
.B2(n_722),
.Y(n_1487)
);

AOI22xp33_ASAP7_75t_L g1488 ( 
.A1(n_1080),
.A2(n_755),
.B1(n_760),
.B2(n_756),
.Y(n_1488)
);

INVx1_ASAP7_75t_L g1489 ( 
.A(n_1081),
.Y(n_1489)
);

INVx2_ASAP7_75t_SL g1490 ( 
.A(n_1143),
.Y(n_1490)
);

AND2x2_ASAP7_75t_L g1491 ( 
.A(n_1153),
.B(n_845),
.Y(n_1491)
);

BUFx6f_ASAP7_75t_L g1492 ( 
.A(n_1221),
.Y(n_1492)
);

INVx3_ASAP7_75t_L g1493 ( 
.A(n_1083),
.Y(n_1493)
);

AOI22xp33_ASAP7_75t_L g1494 ( 
.A1(n_1086),
.A2(n_762),
.B1(n_775),
.B2(n_769),
.Y(n_1494)
);

BUFx6f_ASAP7_75t_L g1495 ( 
.A(n_1229),
.Y(n_1495)
);

BUFx3_ASAP7_75t_L g1496 ( 
.A(n_1143),
.Y(n_1496)
);

BUFx3_ASAP7_75t_L g1497 ( 
.A(n_1114),
.Y(n_1497)
);

INVx1_ASAP7_75t_L g1498 ( 
.A(n_1114),
.Y(n_1498)
);

OAI22xp33_ASAP7_75t_L g1499 ( 
.A1(n_1190),
.A2(n_779),
.B1(n_784),
.B2(n_778),
.Y(n_1499)
);

INVx1_ASAP7_75t_L g1500 ( 
.A(n_1114),
.Y(n_1500)
);

INVx1_ASAP7_75t_L g1501 ( 
.A(n_1110),
.Y(n_1501)
);

BUFx3_ASAP7_75t_L g1502 ( 
.A(n_1229),
.Y(n_1502)
);

AND2x4_ASAP7_75t_L g1503 ( 
.A(n_1131),
.B(n_787),
.Y(n_1503)
);

BUFx6f_ASAP7_75t_SL g1504 ( 
.A(n_1174),
.Y(n_1504)
);

NOR2xp33_ASAP7_75t_L g1505 ( 
.A(n_1407),
.B(n_1139),
.Y(n_1505)
);

OR2x2_ASAP7_75t_L g1506 ( 
.A(n_1342),
.B(n_1196),
.Y(n_1506)
);

NOR2xp33_ASAP7_75t_L g1507 ( 
.A(n_1444),
.B(n_1148),
.Y(n_1507)
);

NOR2xp33_ASAP7_75t_L g1508 ( 
.A(n_1444),
.B(n_1170),
.Y(n_1508)
);

NAND2xp5_ASAP7_75t_L g1509 ( 
.A(n_1333),
.B(n_1153),
.Y(n_1509)
);

NAND2xp5_ASAP7_75t_L g1510 ( 
.A(n_1352),
.B(n_1329),
.Y(n_1510)
);

INVx2_ASAP7_75t_L g1511 ( 
.A(n_1421),
.Y(n_1511)
);

AOI22xp5_ASAP7_75t_L g1512 ( 
.A1(n_1303),
.A2(n_1156),
.B1(n_1245),
.B2(n_1183),
.Y(n_1512)
);

INVx1_ASAP7_75t_L g1513 ( 
.A(n_1374),
.Y(n_1513)
);

INVx1_ASAP7_75t_L g1514 ( 
.A(n_1374),
.Y(n_1514)
);

NOR2xp33_ASAP7_75t_SL g1515 ( 
.A(n_1380),
.B(n_1159),
.Y(n_1515)
);

NAND2xp5_ASAP7_75t_L g1516 ( 
.A(n_1339),
.B(n_1110),
.Y(n_1516)
);

AOI22xp33_ASAP7_75t_L g1517 ( 
.A1(n_1456),
.A2(n_1464),
.B1(n_1273),
.B2(n_1499),
.Y(n_1517)
);

INVx1_ASAP7_75t_SL g1518 ( 
.A(n_1299),
.Y(n_1518)
);

BUFx6f_ASAP7_75t_SL g1519 ( 
.A(n_1269),
.Y(n_1519)
);

INVx1_ASAP7_75t_L g1520 ( 
.A(n_1418),
.Y(n_1520)
);

AND2x2_ASAP7_75t_L g1521 ( 
.A(n_1343),
.B(n_1169),
.Y(n_1521)
);

BUFx3_ASAP7_75t_L g1522 ( 
.A(n_1269),
.Y(n_1522)
);

NAND3xp33_ASAP7_75t_SL g1523 ( 
.A(n_1461),
.B(n_905),
.C(n_844),
.Y(n_1523)
);

NAND2xp5_ASAP7_75t_SL g1524 ( 
.A(n_1499),
.B(n_1044),
.Y(n_1524)
);

NAND2xp5_ASAP7_75t_L g1525 ( 
.A(n_1349),
.B(n_1224),
.Y(n_1525)
);

AND2x2_ASAP7_75t_L g1526 ( 
.A(n_1343),
.B(n_1303),
.Y(n_1526)
);

INVx1_ASAP7_75t_L g1527 ( 
.A(n_1282),
.Y(n_1527)
);

NAND2xp5_ASAP7_75t_L g1528 ( 
.A(n_1353),
.B(n_1177),
.Y(n_1528)
);

INVx2_ASAP7_75t_L g1529 ( 
.A(n_1421),
.Y(n_1529)
);

OAI22xp5_ASAP7_75t_L g1530 ( 
.A1(n_1422),
.A2(n_1157),
.B1(n_1162),
.B2(n_1158),
.Y(n_1530)
);

INVx1_ASAP7_75t_L g1531 ( 
.A(n_1285),
.Y(n_1531)
);

NAND2xp5_ASAP7_75t_L g1532 ( 
.A(n_1353),
.B(n_1177),
.Y(n_1532)
);

NAND2xp5_ASAP7_75t_L g1533 ( 
.A(n_1300),
.B(n_1183),
.Y(n_1533)
);

AOI22xp5_ASAP7_75t_L g1534 ( 
.A1(n_1432),
.A2(n_1183),
.B1(n_1163),
.B2(n_1167),
.Y(n_1534)
);

OR2x2_ASAP7_75t_L g1535 ( 
.A(n_1435),
.B(n_1196),
.Y(n_1535)
);

INVx1_ASAP7_75t_L g1536 ( 
.A(n_1298),
.Y(n_1536)
);

INVxp67_ASAP7_75t_L g1537 ( 
.A(n_1401),
.Y(n_1537)
);

BUFx3_ASAP7_75t_L g1538 ( 
.A(n_1384),
.Y(n_1538)
);

BUFx2_ASAP7_75t_L g1539 ( 
.A(n_1415),
.Y(n_1539)
);

INVx3_ASAP7_75t_L g1540 ( 
.A(n_1286),
.Y(n_1540)
);

NOR2xp33_ASAP7_75t_L g1541 ( 
.A(n_1457),
.B(n_1164),
.Y(n_1541)
);

AOI22xp5_ASAP7_75t_L g1542 ( 
.A1(n_1310),
.A2(n_1395),
.B1(n_1264),
.B2(n_1401),
.Y(n_1542)
);

NAND2xp5_ASAP7_75t_L g1543 ( 
.A(n_1300),
.B(n_1144),
.Y(n_1543)
);

INVx1_ASAP7_75t_L g1544 ( 
.A(n_1314),
.Y(n_1544)
);

BUFx2_ASAP7_75t_L g1545 ( 
.A(n_1260),
.Y(n_1545)
);

NAND2xp5_ASAP7_75t_L g1546 ( 
.A(n_1309),
.B(n_640),
.Y(n_1546)
);

NAND2xp5_ASAP7_75t_L g1547 ( 
.A(n_1311),
.B(n_643),
.Y(n_1547)
);

NAND2xp5_ASAP7_75t_L g1548 ( 
.A(n_1311),
.B(n_1312),
.Y(n_1548)
);

NAND2xp5_ASAP7_75t_SL g1549 ( 
.A(n_1287),
.B(n_1206),
.Y(n_1549)
);

O2A1O1Ixp33_ASAP7_75t_L g1550 ( 
.A1(n_1461),
.A2(n_1157),
.B(n_1150),
.C(n_1152),
.Y(n_1550)
);

NAND2xp5_ASAP7_75t_L g1551 ( 
.A(n_1312),
.B(n_650),
.Y(n_1551)
);

NAND2xp5_ASAP7_75t_L g1552 ( 
.A(n_1273),
.B(n_1422),
.Y(n_1552)
);

OR2x2_ASAP7_75t_L g1553 ( 
.A(n_1264),
.B(n_1181),
.Y(n_1553)
);

OAI22xp5_ASAP7_75t_L g1554 ( 
.A1(n_1323),
.A2(n_1168),
.B1(n_1151),
.B2(n_1166),
.Y(n_1554)
);

INVx3_ASAP7_75t_L g1555 ( 
.A(n_1286),
.Y(n_1555)
);

INVx2_ASAP7_75t_L g1556 ( 
.A(n_1470),
.Y(n_1556)
);

INVx2_ASAP7_75t_L g1557 ( 
.A(n_1470),
.Y(n_1557)
);

AOI22xp33_ASAP7_75t_L g1558 ( 
.A1(n_1326),
.A2(n_791),
.B1(n_798),
.B2(n_797),
.Y(n_1558)
);

AND2x2_ASAP7_75t_L g1559 ( 
.A(n_1263),
.B(n_1149),
.Y(n_1559)
);

NAND2xp5_ASAP7_75t_L g1560 ( 
.A(n_1385),
.B(n_651),
.Y(n_1560)
);

NOR2xp33_ASAP7_75t_L g1561 ( 
.A(n_1457),
.B(n_1166),
.Y(n_1561)
);

INVx1_ASAP7_75t_L g1562 ( 
.A(n_1316),
.Y(n_1562)
);

NAND2xp5_ASAP7_75t_L g1563 ( 
.A(n_1385),
.B(n_659),
.Y(n_1563)
);

O2A1O1Ixp33_ASAP7_75t_L g1564 ( 
.A1(n_1279),
.A2(n_1172),
.B(n_1175),
.C(n_1171),
.Y(n_1564)
);

INVx1_ASAP7_75t_L g1565 ( 
.A(n_1327),
.Y(n_1565)
);

INVx2_ASAP7_75t_L g1566 ( 
.A(n_1433),
.Y(n_1566)
);

NOR2xp33_ASAP7_75t_L g1567 ( 
.A(n_1468),
.B(n_1161),
.Y(n_1567)
);

INVx1_ASAP7_75t_L g1568 ( 
.A(n_1331),
.Y(n_1568)
);

NAND2xp5_ASAP7_75t_L g1569 ( 
.A(n_1403),
.B(n_663),
.Y(n_1569)
);

INVx2_ASAP7_75t_L g1570 ( 
.A(n_1433),
.Y(n_1570)
);

INVx1_ASAP7_75t_L g1571 ( 
.A(n_1332),
.Y(n_1571)
);

INVx1_ASAP7_75t_L g1572 ( 
.A(n_1338),
.Y(n_1572)
);

OAI22xp5_ASAP7_75t_L g1573 ( 
.A1(n_1336),
.A2(n_1367),
.B1(n_1328),
.B2(n_1326),
.Y(n_1573)
);

NAND2xp5_ASAP7_75t_L g1574 ( 
.A(n_1403),
.B(n_666),
.Y(n_1574)
);

NAND2xp5_ASAP7_75t_L g1575 ( 
.A(n_1413),
.B(n_667),
.Y(n_1575)
);

NAND2xp33_ASAP7_75t_L g1576 ( 
.A(n_1368),
.B(n_1161),
.Y(n_1576)
);

INVx1_ASAP7_75t_L g1577 ( 
.A(n_1340),
.Y(n_1577)
);

NAND2xp5_ASAP7_75t_L g1578 ( 
.A(n_1413),
.B(n_673),
.Y(n_1578)
);

NAND2xp5_ASAP7_75t_SL g1579 ( 
.A(n_1287),
.B(n_1206),
.Y(n_1579)
);

INVx2_ASAP7_75t_SL g1580 ( 
.A(n_1350),
.Y(n_1580)
);

INVx2_ASAP7_75t_L g1581 ( 
.A(n_1436),
.Y(n_1581)
);

BUFx3_ASAP7_75t_L g1582 ( 
.A(n_1414),
.Y(n_1582)
);

NAND2xp5_ASAP7_75t_SL g1583 ( 
.A(n_1287),
.B(n_1210),
.Y(n_1583)
);

NAND2xp5_ASAP7_75t_L g1584 ( 
.A(n_1296),
.B(n_674),
.Y(n_1584)
);

INVx2_ASAP7_75t_SL g1585 ( 
.A(n_1350),
.Y(n_1585)
);

INVx2_ASAP7_75t_SL g1586 ( 
.A(n_1350),
.Y(n_1586)
);

INVx2_ASAP7_75t_L g1587 ( 
.A(n_1436),
.Y(n_1587)
);

A2O1A1Ixp33_ASAP7_75t_L g1588 ( 
.A1(n_1344),
.A2(n_1218),
.B(n_1231),
.C(n_1210),
.Y(n_1588)
);

HB1xp67_ASAP7_75t_L g1589 ( 
.A(n_1417),
.Y(n_1589)
);

NOR2xp67_ASAP7_75t_L g1590 ( 
.A(n_1302),
.B(n_1173),
.Y(n_1590)
);

INVx1_ASAP7_75t_L g1591 ( 
.A(n_1348),
.Y(n_1591)
);

BUFx8_ASAP7_75t_L g1592 ( 
.A(n_1288),
.Y(n_1592)
);

OAI22xp5_ASAP7_75t_L g1593 ( 
.A1(n_1336),
.A2(n_1193),
.B1(n_1199),
.B2(n_1198),
.Y(n_1593)
);

AOI22xp5_ASAP7_75t_L g1594 ( 
.A1(n_1396),
.A2(n_1193),
.B1(n_1199),
.B2(n_1198),
.Y(n_1594)
);

OAI22xp33_ASAP7_75t_SL g1595 ( 
.A1(n_1466),
.A2(n_1160),
.B1(n_1178),
.B2(n_1176),
.Y(n_1595)
);

NAND2xp5_ASAP7_75t_SL g1596 ( 
.A(n_1287),
.B(n_1218),
.Y(n_1596)
);

INVx3_ASAP7_75t_L g1597 ( 
.A(n_1297),
.Y(n_1597)
);

INVx2_ASAP7_75t_L g1598 ( 
.A(n_1493),
.Y(n_1598)
);

INVx2_ASAP7_75t_L g1599 ( 
.A(n_1297),
.Y(n_1599)
);

NAND2xp5_ASAP7_75t_SL g1600 ( 
.A(n_1248),
.B(n_1231),
.Y(n_1600)
);

INVx4_ASAP7_75t_L g1601 ( 
.A(n_1368),
.Y(n_1601)
);

INVxp67_ASAP7_75t_L g1602 ( 
.A(n_1368),
.Y(n_1602)
);

BUFx3_ASAP7_75t_L g1603 ( 
.A(n_1414),
.Y(n_1603)
);

NAND2xp5_ASAP7_75t_L g1604 ( 
.A(n_1361),
.B(n_676),
.Y(n_1604)
);

NAND2xp5_ASAP7_75t_L g1605 ( 
.A(n_1361),
.B(n_677),
.Y(n_1605)
);

INVx2_ASAP7_75t_SL g1606 ( 
.A(n_1402),
.Y(n_1606)
);

OAI221xp5_ASAP7_75t_L g1607 ( 
.A1(n_1271),
.A2(n_1173),
.B1(n_1189),
.B2(n_1180),
.C(n_1179),
.Y(n_1607)
);

NAND2xp5_ASAP7_75t_L g1608 ( 
.A(n_1363),
.B(n_687),
.Y(n_1608)
);

INVx1_ASAP7_75t_L g1609 ( 
.A(n_1358),
.Y(n_1609)
);

NAND2xp5_ASAP7_75t_L g1610 ( 
.A(n_1363),
.B(n_688),
.Y(n_1610)
);

AOI22xp33_ASAP7_75t_L g1611 ( 
.A1(n_1328),
.A2(n_805),
.B1(n_815),
.B2(n_810),
.Y(n_1611)
);

AND2x2_ASAP7_75t_L g1612 ( 
.A(n_1318),
.B(n_1174),
.Y(n_1612)
);

OAI22x1_ASAP7_75t_R g1613 ( 
.A1(n_1301),
.A2(n_1197),
.B1(n_1200),
.B2(n_1182),
.Y(n_1613)
);

NAND2xp5_ASAP7_75t_L g1614 ( 
.A(n_1307),
.B(n_690),
.Y(n_1614)
);

OAI22xp5_ASAP7_75t_L g1615 ( 
.A1(n_1367),
.A2(n_1174),
.B1(n_820),
.B2(n_826),
.Y(n_1615)
);

INVx2_ASAP7_75t_L g1616 ( 
.A(n_1249),
.Y(n_1616)
);

NOR2xp33_ASAP7_75t_L g1617 ( 
.A(n_1356),
.B(n_691),
.Y(n_1617)
);

INVxp33_ASAP7_75t_L g1618 ( 
.A(n_1426),
.Y(n_1618)
);

NAND2xp5_ASAP7_75t_L g1619 ( 
.A(n_1313),
.B(n_707),
.Y(n_1619)
);

AND2x2_ASAP7_75t_L g1620 ( 
.A(n_1389),
.B(n_1182),
.Y(n_1620)
);

OR2x2_ASAP7_75t_L g1621 ( 
.A(n_1261),
.B(n_1182),
.Y(n_1621)
);

OAI22xp5_ASAP7_75t_L g1622 ( 
.A1(n_1373),
.A2(n_833),
.B1(n_842),
.B2(n_817),
.Y(n_1622)
);

BUFx6f_ASAP7_75t_L g1623 ( 
.A(n_1502),
.Y(n_1623)
);

NAND2xp5_ASAP7_75t_L g1624 ( 
.A(n_1362),
.B(n_1376),
.Y(n_1624)
);

OR2x2_ASAP7_75t_L g1625 ( 
.A(n_1441),
.B(n_1200),
.Y(n_1625)
);

NOR3xp33_ASAP7_75t_L g1626 ( 
.A(n_1378),
.B(n_1252),
.C(n_1471),
.Y(n_1626)
);

O2A1O1Ixp33_ASAP7_75t_L g1627 ( 
.A1(n_1377),
.A2(n_853),
.B(n_861),
.C(n_855),
.Y(n_1627)
);

INVx2_ASAP7_75t_L g1628 ( 
.A(n_1255),
.Y(n_1628)
);

BUFx6f_ASAP7_75t_L g1629 ( 
.A(n_1502),
.Y(n_1629)
);

INVx4_ASAP7_75t_L g1630 ( 
.A(n_1368),
.Y(n_1630)
);

BUFx6f_ASAP7_75t_L g1631 ( 
.A(n_1319),
.Y(n_1631)
);

AOI221xp5_ASAP7_75t_L g1632 ( 
.A1(n_1253),
.A2(n_1200),
.B1(n_862),
.B2(n_868),
.C(n_864),
.Y(n_1632)
);

NAND2xp5_ASAP7_75t_SL g1633 ( 
.A(n_1248),
.B(n_1242),
.Y(n_1633)
);

AO22x1_ASAP7_75t_L g1634 ( 
.A1(n_1266),
.A2(n_1200),
.B1(n_727),
.B2(n_731),
.Y(n_1634)
);

AOI21xp5_ASAP7_75t_L g1635 ( 
.A1(n_1275),
.A2(n_1247),
.B(n_1244),
.Y(n_1635)
);

INVx1_ASAP7_75t_L g1636 ( 
.A(n_1399),
.Y(n_1636)
);

INVx2_ASAP7_75t_L g1637 ( 
.A(n_1262),
.Y(n_1637)
);

BUFx8_ASAP7_75t_L g1638 ( 
.A(n_1288),
.Y(n_1638)
);

AND2x6_ASAP7_75t_L g1639 ( 
.A(n_1373),
.B(n_1244),
.Y(n_1639)
);

INVx2_ASAP7_75t_L g1640 ( 
.A(n_1281),
.Y(n_1640)
);

NAND2xp5_ASAP7_75t_SL g1641 ( 
.A(n_1251),
.B(n_1319),
.Y(n_1641)
);

AND2x4_ASAP7_75t_L g1642 ( 
.A(n_1402),
.B(n_863),
.Y(n_1642)
);

INVx2_ASAP7_75t_L g1643 ( 
.A(n_1292),
.Y(n_1643)
);

INVx2_ASAP7_75t_L g1644 ( 
.A(n_1295),
.Y(n_1644)
);

A2O1A1Ixp33_ASAP7_75t_L g1645 ( 
.A1(n_1419),
.A2(n_874),
.B(n_878),
.C(n_870),
.Y(n_1645)
);

NOR2xp33_ASAP7_75t_L g1646 ( 
.A(n_1356),
.B(n_740),
.Y(n_1646)
);

INVx2_ASAP7_75t_L g1647 ( 
.A(n_1305),
.Y(n_1647)
);

INVx2_ASAP7_75t_L g1648 ( 
.A(n_1306),
.Y(n_1648)
);

INVx3_ASAP7_75t_L g1649 ( 
.A(n_1290),
.Y(n_1649)
);

INVx2_ASAP7_75t_L g1650 ( 
.A(n_1315),
.Y(n_1650)
);

OA21x2_ASAP7_75t_L g1651 ( 
.A1(n_1251),
.A2(n_1247),
.B(n_884),
.Y(n_1651)
);

O2A1O1Ixp33_ASAP7_75t_L g1652 ( 
.A1(n_1274),
.A2(n_887),
.B(n_891),
.C(n_883),
.Y(n_1652)
);

NAND2xp5_ASAP7_75t_L g1653 ( 
.A(n_1428),
.B(n_1429),
.Y(n_1653)
);

INVx1_ASAP7_75t_L g1654 ( 
.A(n_1431),
.Y(n_1654)
);

NAND2xp5_ASAP7_75t_L g1655 ( 
.A(n_1337),
.B(n_741),
.Y(n_1655)
);

BUFx6f_ASAP7_75t_L g1656 ( 
.A(n_1320),
.Y(n_1656)
);

INVx3_ASAP7_75t_L g1657 ( 
.A(n_1290),
.Y(n_1657)
);

NAND2xp5_ASAP7_75t_L g1658 ( 
.A(n_1347),
.B(n_743),
.Y(n_1658)
);

AND2x2_ASAP7_75t_L g1659 ( 
.A(n_1390),
.B(n_846),
.Y(n_1659)
);

NAND2xp5_ASAP7_75t_L g1660 ( 
.A(n_1357),
.B(n_744),
.Y(n_1660)
);

NOR2xp67_ASAP7_75t_L g1661 ( 
.A(n_1406),
.B(n_12),
.Y(n_1661)
);

NAND3xp33_ASAP7_75t_L g1662 ( 
.A(n_1404),
.B(n_748),
.C(n_745),
.Y(n_1662)
);

NOR2xp33_ASAP7_75t_L g1663 ( 
.A(n_1289),
.B(n_751),
.Y(n_1663)
);

NOR3xp33_ASAP7_75t_L g1664 ( 
.A(n_1445),
.B(n_859),
.C(n_794),
.Y(n_1664)
);

INVx2_ASAP7_75t_L g1665 ( 
.A(n_1317),
.Y(n_1665)
);

NAND2xp5_ASAP7_75t_L g1666 ( 
.A(n_1359),
.B(n_753),
.Y(n_1666)
);

AOI22xp33_ASAP7_75t_L g1667 ( 
.A1(n_1489),
.A2(n_900),
.B1(n_894),
.B2(n_841),
.Y(n_1667)
);

INVxp67_ASAP7_75t_L g1668 ( 
.A(n_1417),
.Y(n_1668)
);

INVx8_ASAP7_75t_L g1669 ( 
.A(n_1402),
.Y(n_1669)
);

AOI22xp5_ASAP7_75t_L g1670 ( 
.A1(n_1397),
.A2(n_757),
.B1(n_763),
.B2(n_754),
.Y(n_1670)
);

NOR2xp33_ASAP7_75t_R g1671 ( 
.A(n_1391),
.B(n_764),
.Y(n_1671)
);

NOR2xp33_ASAP7_75t_L g1672 ( 
.A(n_1294),
.B(n_765),
.Y(n_1672)
);

INVx1_ASAP7_75t_L g1673 ( 
.A(n_1497),
.Y(n_1673)
);

NAND2xp5_ASAP7_75t_L g1674 ( 
.A(n_1370),
.B(n_766),
.Y(n_1674)
);

AND2x6_ASAP7_75t_L g1675 ( 
.A(n_1320),
.B(n_685),
.Y(n_1675)
);

BUFx3_ASAP7_75t_L g1676 ( 
.A(n_1424),
.Y(n_1676)
);

INVx1_ASAP7_75t_L g1677 ( 
.A(n_1497),
.Y(n_1677)
);

INVx2_ASAP7_75t_L g1678 ( 
.A(n_1379),
.Y(n_1678)
);

CKINVDCx5p33_ASAP7_75t_R g1679 ( 
.A(n_1391),
.Y(n_1679)
);

OAI21xp5_ASAP7_75t_L g1680 ( 
.A1(n_1275),
.A2(n_733),
.B(n_710),
.Y(n_1680)
);

NAND2xp5_ASAP7_75t_SL g1681 ( 
.A(n_1276),
.B(n_636),
.Y(n_1681)
);

OR2x6_ASAP7_75t_SL g1682 ( 
.A(n_1410),
.B(n_777),
.Y(n_1682)
);

INVx2_ASAP7_75t_L g1683 ( 
.A(n_1382),
.Y(n_1683)
);

INVx2_ASAP7_75t_L g1684 ( 
.A(n_1388),
.Y(n_1684)
);

INVxp67_ASAP7_75t_L g1685 ( 
.A(n_1417),
.Y(n_1685)
);

INVxp67_ASAP7_75t_L g1686 ( 
.A(n_1280),
.Y(n_1686)
);

INVx1_ASAP7_75t_L g1687 ( 
.A(n_1498),
.Y(n_1687)
);

AO22x2_ASAP7_75t_L g1688 ( 
.A1(n_1265),
.A2(n_739),
.B1(n_846),
.B2(n_14),
.Y(n_1688)
);

INVx3_ASAP7_75t_L g1689 ( 
.A(n_1335),
.Y(n_1689)
);

INVxp67_ASAP7_75t_L g1690 ( 
.A(n_1280),
.Y(n_1690)
);

NAND2xp5_ASAP7_75t_L g1691 ( 
.A(n_1372),
.B(n_780),
.Y(n_1691)
);

INVx3_ASAP7_75t_L g1692 ( 
.A(n_1335),
.Y(n_1692)
);

NAND2xp5_ASAP7_75t_L g1693 ( 
.A(n_1268),
.B(n_783),
.Y(n_1693)
);

INVx1_ASAP7_75t_L g1694 ( 
.A(n_1500),
.Y(n_1694)
);

INVx1_ASAP7_75t_L g1695 ( 
.A(n_1448),
.Y(n_1695)
);

NAND2xp5_ASAP7_75t_SL g1696 ( 
.A(n_1439),
.B(n_648),
.Y(n_1696)
);

NAND2xp5_ASAP7_75t_SL g1697 ( 
.A(n_1439),
.B(n_649),
.Y(n_1697)
);

NAND2xp5_ASAP7_75t_L g1698 ( 
.A(n_1277),
.B(n_785),
.Y(n_1698)
);

NAND2xp5_ASAP7_75t_SL g1699 ( 
.A(n_1452),
.B(n_662),
.Y(n_1699)
);

AND2x4_ASAP7_75t_L g1700 ( 
.A(n_1321),
.B(n_685),
.Y(n_1700)
);

INVx2_ASAP7_75t_L g1701 ( 
.A(n_1408),
.Y(n_1701)
);

INVx1_ASAP7_75t_L g1702 ( 
.A(n_1453),
.Y(n_1702)
);

INVx1_ASAP7_75t_L g1703 ( 
.A(n_1454),
.Y(n_1703)
);

INVx2_ASAP7_75t_L g1704 ( 
.A(n_1411),
.Y(n_1704)
);

NAND2xp5_ASAP7_75t_L g1705 ( 
.A(n_1257),
.B(n_786),
.Y(n_1705)
);

NOR2xp33_ASAP7_75t_L g1706 ( 
.A(n_1355),
.B(n_790),
.Y(n_1706)
);

NAND2xp5_ASAP7_75t_L g1707 ( 
.A(n_1259),
.B(n_792),
.Y(n_1707)
);

NAND2xp5_ASAP7_75t_SL g1708 ( 
.A(n_1452),
.B(n_664),
.Y(n_1708)
);

INVx1_ASAP7_75t_L g1709 ( 
.A(n_1460),
.Y(n_1709)
);

NAND2xp5_ASAP7_75t_L g1710 ( 
.A(n_1503),
.B(n_796),
.Y(n_1710)
);

OR2x2_ASAP7_75t_L g1711 ( 
.A(n_1334),
.B(n_802),
.Y(n_1711)
);

INVx1_ASAP7_75t_L g1712 ( 
.A(n_1462),
.Y(n_1712)
);

NOR2xp33_ASAP7_75t_L g1713 ( 
.A(n_1256),
.B(n_804),
.Y(n_1713)
);

INVx1_ASAP7_75t_L g1714 ( 
.A(n_1463),
.Y(n_1714)
);

NAND2xp5_ASAP7_75t_SL g1715 ( 
.A(n_1503),
.B(n_665),
.Y(n_1715)
);

NAND2xp5_ASAP7_75t_SL g1716 ( 
.A(n_1420),
.B(n_669),
.Y(n_1716)
);

INVxp67_ASAP7_75t_L g1717 ( 
.A(n_1280),
.Y(n_1717)
);

INVx2_ASAP7_75t_L g1718 ( 
.A(n_1412),
.Y(n_1718)
);

AND2x2_ASAP7_75t_L g1719 ( 
.A(n_1491),
.B(n_846),
.Y(n_1719)
);

NAND2xp5_ASAP7_75t_SL g1720 ( 
.A(n_1420),
.B(n_683),
.Y(n_1720)
);

INVx1_ASAP7_75t_L g1721 ( 
.A(n_1465),
.Y(n_1721)
);

INVx1_ASAP7_75t_L g1722 ( 
.A(n_1467),
.Y(n_1722)
);

INVx1_ASAP7_75t_L g1723 ( 
.A(n_1481),
.Y(n_1723)
);

AND2x2_ASAP7_75t_L g1724 ( 
.A(n_1383),
.B(n_808),
.Y(n_1724)
);

NAND2xp5_ASAP7_75t_SL g1725 ( 
.A(n_1420),
.B(n_686),
.Y(n_1725)
);

AND2x2_ASAP7_75t_L g1726 ( 
.A(n_1383),
.B(n_813),
.Y(n_1726)
);

INVx2_ASAP7_75t_L g1727 ( 
.A(n_1425),
.Y(n_1727)
);

NAND2xp5_ASAP7_75t_SL g1728 ( 
.A(n_1423),
.B(n_699),
.Y(n_1728)
);

AND2x4_ASAP7_75t_L g1729 ( 
.A(n_1480),
.B(n_685),
.Y(n_1729)
);

INVx2_ASAP7_75t_L g1730 ( 
.A(n_1443),
.Y(n_1730)
);

NAND2xp5_ASAP7_75t_L g1731 ( 
.A(n_1450),
.B(n_818),
.Y(n_1731)
);

NAND2xp5_ASAP7_75t_SL g1732 ( 
.A(n_1423),
.B(n_701),
.Y(n_1732)
);

INVx2_ASAP7_75t_L g1733 ( 
.A(n_1458),
.Y(n_1733)
);

NAND2xp5_ASAP7_75t_SL g1734 ( 
.A(n_1423),
.B(n_702),
.Y(n_1734)
);

NAND2xp5_ASAP7_75t_L g1735 ( 
.A(n_1475),
.B(n_822),
.Y(n_1735)
);

OAI22xp5_ASAP7_75t_L g1736 ( 
.A1(n_1283),
.A2(n_829),
.B1(n_831),
.B2(n_830),
.Y(n_1736)
);

NAND2xp5_ASAP7_75t_L g1737 ( 
.A(n_1483),
.B(n_832),
.Y(n_1737)
);

NAND2xp5_ASAP7_75t_SL g1738 ( 
.A(n_1430),
.B(n_713),
.Y(n_1738)
);

INVx1_ASAP7_75t_L g1739 ( 
.A(n_1476),
.Y(n_1739)
);

NAND2xp5_ASAP7_75t_SL g1740 ( 
.A(n_1430),
.B(n_714),
.Y(n_1740)
);

INVx3_ASAP7_75t_L g1741 ( 
.A(n_1424),
.Y(n_1741)
);

HB1xp67_ASAP7_75t_L g1742 ( 
.A(n_1346),
.Y(n_1742)
);

BUFx6f_ASAP7_75t_SL g1743 ( 
.A(n_1270),
.Y(n_1743)
);

INVx1_ASAP7_75t_L g1744 ( 
.A(n_1482),
.Y(n_1744)
);

INVx2_ASAP7_75t_L g1745 ( 
.A(n_1484),
.Y(n_1745)
);

NAND2xp5_ASAP7_75t_L g1746 ( 
.A(n_1250),
.B(n_835),
.Y(n_1746)
);

AOI21xp5_ASAP7_75t_L g1747 ( 
.A1(n_1265),
.A2(n_724),
.B(n_715),
.Y(n_1747)
);

INVx1_ASAP7_75t_L g1748 ( 
.A(n_1346),
.Y(n_1748)
);

AOI22xp33_ASAP7_75t_L g1749 ( 
.A1(n_1284),
.A2(n_841),
.B1(n_897),
.B2(n_685),
.Y(n_1749)
);

INVx1_ASAP7_75t_L g1750 ( 
.A(n_1346),
.Y(n_1750)
);

INVx3_ASAP7_75t_L g1751 ( 
.A(n_1496),
.Y(n_1751)
);

BUFx3_ASAP7_75t_L g1752 ( 
.A(n_1496),
.Y(n_1752)
);

NAND2xp5_ASAP7_75t_L g1753 ( 
.A(n_1254),
.B(n_737),
.Y(n_1753)
);

NAND2xp5_ASAP7_75t_SL g1754 ( 
.A(n_1430),
.B(n_752),
.Y(n_1754)
);

NAND2xp5_ASAP7_75t_SL g1755 ( 
.A(n_1430),
.B(n_758),
.Y(n_1755)
);

INVx1_ASAP7_75t_L g1756 ( 
.A(n_1258),
.Y(n_1756)
);

INVx8_ASAP7_75t_L g1757 ( 
.A(n_1504),
.Y(n_1757)
);

HB1xp67_ASAP7_75t_L g1758 ( 
.A(n_1504),
.Y(n_1758)
);

NAND2xp5_ASAP7_75t_L g1759 ( 
.A(n_1404),
.B(n_772),
.Y(n_1759)
);

AND2x2_ASAP7_75t_L g1760 ( 
.A(n_1478),
.B(n_841),
.Y(n_1760)
);

INVxp33_ASAP7_75t_L g1761 ( 
.A(n_1409),
.Y(n_1761)
);

NAND3xp33_ASAP7_75t_L g1762 ( 
.A(n_1451),
.B(n_795),
.C(n_774),
.Y(n_1762)
);

NOR2xp67_ASAP7_75t_L g1763 ( 
.A(n_1293),
.B(n_12),
.Y(n_1763)
);

NAND2xp5_ASAP7_75t_SL g1764 ( 
.A(n_1447),
.B(n_803),
.Y(n_1764)
);

INVx1_ASAP7_75t_L g1765 ( 
.A(n_1267),
.Y(n_1765)
);

INVx1_ASAP7_75t_L g1766 ( 
.A(n_1267),
.Y(n_1766)
);

INVx1_ASAP7_75t_L g1767 ( 
.A(n_1501),
.Y(n_1767)
);

INVx2_ASAP7_75t_L g1768 ( 
.A(n_1322),
.Y(n_1768)
);

AND2x2_ASAP7_75t_L g1769 ( 
.A(n_1440),
.B(n_841),
.Y(n_1769)
);

OAI22xp33_ASAP7_75t_L g1770 ( 
.A1(n_1438),
.A2(n_897),
.B1(n_841),
.B2(n_809),
.Y(n_1770)
);

NAND2xp5_ASAP7_75t_L g1771 ( 
.A(n_1416),
.B(n_807),
.Y(n_1771)
);

INVx1_ASAP7_75t_L g1772 ( 
.A(n_1325),
.Y(n_1772)
);

INVx2_ASAP7_75t_SL g1773 ( 
.A(n_1398),
.Y(n_1773)
);

AO22x2_ASAP7_75t_L g1774 ( 
.A1(n_1427),
.A2(n_15),
.B1(n_13),
.B2(n_14),
.Y(n_1774)
);

NOR2xp33_ASAP7_75t_L g1775 ( 
.A(n_1442),
.B(n_811),
.Y(n_1775)
);

AND2x2_ASAP7_75t_L g1776 ( 
.A(n_1487),
.B(n_897),
.Y(n_1776)
);

AOI22xp5_ASAP7_75t_L g1777 ( 
.A1(n_1280),
.A2(n_816),
.B1(n_828),
.B2(n_814),
.Y(n_1777)
);

OR2x6_ASAP7_75t_L g1778 ( 
.A(n_1381),
.B(n_897),
.Y(n_1778)
);

NAND2xp5_ASAP7_75t_L g1779 ( 
.A(n_1416),
.B(n_837),
.Y(n_1779)
);

INVx1_ASAP7_75t_L g1780 ( 
.A(n_1330),
.Y(n_1780)
);

BUFx5_ASAP7_75t_L g1781 ( 
.A(n_1405),
.Y(n_1781)
);

INVx2_ASAP7_75t_L g1782 ( 
.A(n_1308),
.Y(n_1782)
);

NAND2xp5_ASAP7_75t_SL g1783 ( 
.A(n_1447),
.B(n_557),
.Y(n_1783)
);

NAND2xp5_ASAP7_75t_L g1784 ( 
.A(n_1446),
.B(n_13),
.Y(n_1784)
);

INVx2_ASAP7_75t_SL g1785 ( 
.A(n_1398),
.Y(n_1785)
);

NOR2xp33_ASAP7_75t_L g1786 ( 
.A(n_1442),
.B(n_15),
.Y(n_1786)
);

NAND2xp33_ASAP7_75t_SL g1787 ( 
.A(n_1381),
.B(n_18),
.Y(n_1787)
);

CKINVDCx5p33_ASAP7_75t_R g1788 ( 
.A(n_1486),
.Y(n_1788)
);

INVx6_ASAP7_75t_L g1789 ( 
.A(n_1473),
.Y(n_1789)
);

NAND2xp5_ASAP7_75t_L g1790 ( 
.A(n_1446),
.B(n_19),
.Y(n_1790)
);

NAND2xp5_ASAP7_75t_L g1791 ( 
.A(n_1283),
.B(n_1291),
.Y(n_1791)
);

NAND2xp33_ASAP7_75t_L g1792 ( 
.A(n_1405),
.B(n_377),
.Y(n_1792)
);

AOI21xp33_ASAP7_75t_L g1793 ( 
.A1(n_1786),
.A2(n_1284),
.B(n_1472),
.Y(n_1793)
);

NOR3xp33_ASAP7_75t_L g1794 ( 
.A(n_1607),
.B(n_1392),
.C(n_1386),
.Y(n_1794)
);

AOI21xp5_ASAP7_75t_L g1795 ( 
.A1(n_1641),
.A2(n_1485),
.B(n_1351),
.Y(n_1795)
);

BUFx6f_ASAP7_75t_L g1796 ( 
.A(n_1631),
.Y(n_1796)
);

INVx3_ASAP7_75t_L g1797 ( 
.A(n_1789),
.Y(n_1797)
);

AOI21xp5_ASAP7_75t_L g1798 ( 
.A1(n_1600),
.A2(n_1278),
.B(n_1272),
.Y(n_1798)
);

NAND2xp5_ASAP7_75t_SL g1799 ( 
.A(n_1515),
.B(n_1354),
.Y(n_1799)
);

NAND2xp5_ASAP7_75t_L g1800 ( 
.A(n_1520),
.B(n_1527),
.Y(n_1800)
);

NAND2xp5_ASAP7_75t_L g1801 ( 
.A(n_1531),
.B(n_1341),
.Y(n_1801)
);

AND2x2_ASAP7_75t_L g1802 ( 
.A(n_1526),
.B(n_1537),
.Y(n_1802)
);

NAND2xp5_ASAP7_75t_L g1803 ( 
.A(n_1536),
.B(n_1341),
.Y(n_1803)
);

NAND2xp5_ASAP7_75t_L g1804 ( 
.A(n_1544),
.B(n_1487),
.Y(n_1804)
);

AOI21xp5_ASAP7_75t_L g1805 ( 
.A1(n_1600),
.A2(n_1278),
.B(n_1272),
.Y(n_1805)
);

INVx3_ASAP7_75t_L g1806 ( 
.A(n_1789),
.Y(n_1806)
);

AOI21xp5_ASAP7_75t_L g1807 ( 
.A1(n_1633),
.A2(n_1477),
.B(n_1455),
.Y(n_1807)
);

INVx2_ASAP7_75t_SL g1808 ( 
.A(n_1757),
.Y(n_1808)
);

NOR2xp33_ASAP7_75t_L g1809 ( 
.A(n_1618),
.B(n_1486),
.Y(n_1809)
);

INVx2_ASAP7_75t_L g1810 ( 
.A(n_1651),
.Y(n_1810)
);

NOR2xp33_ASAP7_75t_SL g1811 ( 
.A(n_1669),
.B(n_1301),
.Y(n_1811)
);

AND2x2_ASAP7_75t_L g1812 ( 
.A(n_1537),
.B(n_1488),
.Y(n_1812)
);

INVx1_ASAP7_75t_L g1813 ( 
.A(n_1562),
.Y(n_1813)
);

NAND2xp5_ASAP7_75t_SL g1814 ( 
.A(n_1542),
.B(n_1354),
.Y(n_1814)
);

A2O1A1Ixp33_ASAP7_75t_L g1815 ( 
.A1(n_1548),
.A2(n_1490),
.B(n_1365),
.C(n_1366),
.Y(n_1815)
);

NAND2xp5_ASAP7_75t_L g1816 ( 
.A(n_1565),
.B(n_1568),
.Y(n_1816)
);

OAI22xp5_ASAP7_75t_L g1817 ( 
.A1(n_1552),
.A2(n_1394),
.B1(n_1366),
.B2(n_1365),
.Y(n_1817)
);

INVx2_ASAP7_75t_L g1818 ( 
.A(n_1571),
.Y(n_1818)
);

INVx2_ASAP7_75t_L g1819 ( 
.A(n_1572),
.Y(n_1819)
);

OAI21xp5_ASAP7_75t_L g1820 ( 
.A1(n_1525),
.A2(n_1477),
.B(n_1455),
.Y(n_1820)
);

A2O1A1Ixp33_ASAP7_75t_L g1821 ( 
.A1(n_1786),
.A2(n_1550),
.B(n_1510),
.C(n_1507),
.Y(n_1821)
);

OR2x2_ASAP7_75t_L g1822 ( 
.A(n_1518),
.B(n_1488),
.Y(n_1822)
);

NOR2xp67_ASAP7_75t_L g1823 ( 
.A(n_1679),
.B(n_1386),
.Y(n_1823)
);

NAND2xp5_ASAP7_75t_SL g1824 ( 
.A(n_1580),
.B(n_1473),
.Y(n_1824)
);

BUFx3_ASAP7_75t_L g1825 ( 
.A(n_1592),
.Y(n_1825)
);

NAND2xp5_ASAP7_75t_L g1826 ( 
.A(n_1577),
.B(n_1494),
.Y(n_1826)
);

OR2x6_ASAP7_75t_L g1827 ( 
.A(n_1669),
.B(n_1392),
.Y(n_1827)
);

INVx1_ASAP7_75t_L g1828 ( 
.A(n_1591),
.Y(n_1828)
);

AND2x6_ASAP7_75t_L g1829 ( 
.A(n_1631),
.B(n_1364),
.Y(n_1829)
);

NAND2xp5_ASAP7_75t_L g1830 ( 
.A(n_1508),
.B(n_1494),
.Y(n_1830)
);

NAND2xp5_ASAP7_75t_L g1831 ( 
.A(n_1508),
.B(n_1437),
.Y(n_1831)
);

BUFx6f_ASAP7_75t_L g1832 ( 
.A(n_1631),
.Y(n_1832)
);

O2A1O1Ixp33_ASAP7_75t_L g1833 ( 
.A1(n_1528),
.A2(n_1459),
.B(n_1437),
.C(n_1387),
.Y(n_1833)
);

OAI21xp5_ASAP7_75t_L g1834 ( 
.A1(n_1635),
.A2(n_1588),
.B(n_1791),
.Y(n_1834)
);

NAND2xp5_ASAP7_75t_L g1835 ( 
.A(n_1532),
.B(n_1459),
.Y(n_1835)
);

INVx4_ASAP7_75t_L g1836 ( 
.A(n_1669),
.Y(n_1836)
);

BUFx6f_ASAP7_75t_L g1837 ( 
.A(n_1631),
.Y(n_1837)
);

NAND2xp5_ASAP7_75t_L g1838 ( 
.A(n_1521),
.B(n_1304),
.Y(n_1838)
);

INVx2_ASAP7_75t_L g1839 ( 
.A(n_1609),
.Y(n_1839)
);

NAND2xp5_ASAP7_75t_L g1840 ( 
.A(n_1533),
.B(n_1304),
.Y(n_1840)
);

INVx4_ASAP7_75t_L g1841 ( 
.A(n_1757),
.Y(n_1841)
);

NOR2xp33_ASAP7_75t_L g1842 ( 
.A(n_1506),
.B(n_1535),
.Y(n_1842)
);

NOR2xp67_ASAP7_75t_L g1843 ( 
.A(n_1758),
.B(n_1434),
.Y(n_1843)
);

AOI21xp5_ASAP7_75t_L g1844 ( 
.A1(n_1549),
.A2(n_1583),
.B(n_1579),
.Y(n_1844)
);

OAI22xp5_ASAP7_75t_L g1845 ( 
.A1(n_1517),
.A2(n_1469),
.B1(n_1474),
.B2(n_1434),
.Y(n_1845)
);

OAI21xp5_ASAP7_75t_L g1846 ( 
.A1(n_1516),
.A2(n_1369),
.B(n_1364),
.Y(n_1846)
);

INVx1_ASAP7_75t_L g1847 ( 
.A(n_1636),
.Y(n_1847)
);

AOI21xp5_ASAP7_75t_L g1848 ( 
.A1(n_1579),
.A2(n_1596),
.B(n_1583),
.Y(n_1848)
);

NAND2xp5_ASAP7_75t_L g1849 ( 
.A(n_1509),
.B(n_1304),
.Y(n_1849)
);

INVx2_ASAP7_75t_L g1850 ( 
.A(n_1654),
.Y(n_1850)
);

AOI21xp5_ASAP7_75t_L g1851 ( 
.A1(n_1596),
.A2(n_1360),
.B(n_1447),
.Y(n_1851)
);

BUFx12f_ASAP7_75t_L g1852 ( 
.A(n_1592),
.Y(n_1852)
);

NAND2xp5_ASAP7_75t_SL g1853 ( 
.A(n_1585),
.B(n_1469),
.Y(n_1853)
);

INVxp67_ASAP7_75t_L g1854 ( 
.A(n_1539),
.Y(n_1854)
);

NAND2xp5_ASAP7_75t_SL g1855 ( 
.A(n_1586),
.B(n_1474),
.Y(n_1855)
);

AND2x4_ASAP7_75t_L g1856 ( 
.A(n_1606),
.B(n_1427),
.Y(n_1856)
);

O2A1O1Ixp5_ASAP7_75t_L g1857 ( 
.A1(n_1680),
.A2(n_1681),
.B(n_1524),
.C(n_1770),
.Y(n_1857)
);

AOI21xp5_ASAP7_75t_L g1858 ( 
.A1(n_1624),
.A2(n_1492),
.B(n_1449),
.Y(n_1858)
);

NOR2xp33_ASAP7_75t_L g1859 ( 
.A(n_1545),
.B(n_1479),
.Y(n_1859)
);

AND2x2_ASAP7_75t_L g1860 ( 
.A(n_1672),
.B(n_1479),
.Y(n_1860)
);

AND2x4_ASAP7_75t_L g1861 ( 
.A(n_1522),
.B(n_1427),
.Y(n_1861)
);

INVx1_ASAP7_75t_L g1862 ( 
.A(n_1653),
.Y(n_1862)
);

AOI22xp5_ASAP7_75t_L g1863 ( 
.A1(n_1559),
.A2(n_1304),
.B1(n_1371),
.B2(n_1393),
.Y(n_1863)
);

INVx3_ASAP7_75t_L g1864 ( 
.A(n_1789),
.Y(n_1864)
);

NAND2xp5_ASAP7_75t_L g1865 ( 
.A(n_1561),
.B(n_1324),
.Y(n_1865)
);

AND2x2_ASAP7_75t_L g1866 ( 
.A(n_1672),
.B(n_1324),
.Y(n_1866)
);

CKINVDCx20_ASAP7_75t_R g1867 ( 
.A(n_1638),
.Y(n_1867)
);

NOR2xp33_ASAP7_75t_L g1868 ( 
.A(n_1534),
.B(n_1371),
.Y(n_1868)
);

BUFx6f_ASAP7_75t_L g1869 ( 
.A(n_1656),
.Y(n_1869)
);

NOR2xp33_ASAP7_75t_L g1870 ( 
.A(n_1711),
.B(n_1324),
.Y(n_1870)
);

NAND2xp5_ASAP7_75t_L g1871 ( 
.A(n_1561),
.B(n_1324),
.Y(n_1871)
);

OAI21xp5_ASAP7_75t_L g1872 ( 
.A1(n_1756),
.A2(n_1375),
.B(n_1345),
.Y(n_1872)
);

A2O1A1Ixp33_ASAP7_75t_L g1873 ( 
.A1(n_1541),
.A2(n_1375),
.B(n_1400),
.C(n_1345),
.Y(n_1873)
);

NAND2xp5_ASAP7_75t_L g1874 ( 
.A(n_1512),
.B(n_1541),
.Y(n_1874)
);

NAND2xp5_ASAP7_75t_SL g1875 ( 
.A(n_1668),
.B(n_1345),
.Y(n_1875)
);

NAND2xp5_ASAP7_75t_SL g1876 ( 
.A(n_1668),
.B(n_1400),
.Y(n_1876)
);

INVx3_ASAP7_75t_L g1877 ( 
.A(n_1649),
.Y(n_1877)
);

A2O1A1Ixp33_ASAP7_75t_L g1878 ( 
.A1(n_1652),
.A2(n_1400),
.B(n_1495),
.C(n_1393),
.Y(n_1878)
);

NOR2x1_ASAP7_75t_R g1879 ( 
.A(n_1788),
.B(n_1393),
.Y(n_1879)
);

NAND2xp5_ASAP7_75t_L g1880 ( 
.A(n_1505),
.B(n_1495),
.Y(n_1880)
);

NAND2xp5_ASAP7_75t_L g1881 ( 
.A(n_1659),
.B(n_20),
.Y(n_1881)
);

OAI21xp5_ASAP7_75t_L g1882 ( 
.A1(n_1765),
.A2(n_382),
.B(n_380),
.Y(n_1882)
);

NOR3xp33_ASAP7_75t_L g1883 ( 
.A(n_1523),
.B(n_21),
.C(n_23),
.Y(n_1883)
);

INVx4_ASAP7_75t_L g1884 ( 
.A(n_1757),
.Y(n_1884)
);

NAND2xp5_ASAP7_75t_L g1885 ( 
.A(n_1558),
.B(n_21),
.Y(n_1885)
);

NAND2xp5_ASAP7_75t_L g1886 ( 
.A(n_1558),
.B(n_24),
.Y(n_1886)
);

A2O1A1Ixp33_ASAP7_75t_L g1887 ( 
.A1(n_1627),
.A2(n_27),
.B(n_24),
.C(n_26),
.Y(n_1887)
);

NAND2xp5_ASAP7_75t_L g1888 ( 
.A(n_1611),
.B(n_26),
.Y(n_1888)
);

A2O1A1Ixp33_ASAP7_75t_L g1889 ( 
.A1(n_1706),
.A2(n_29),
.B(n_27),
.C(n_28),
.Y(n_1889)
);

INVx1_ASAP7_75t_L g1890 ( 
.A(n_1687),
.Y(n_1890)
);

NAND2xp5_ASAP7_75t_L g1891 ( 
.A(n_1513),
.B(n_28),
.Y(n_1891)
);

OAI21xp5_ASAP7_75t_L g1892 ( 
.A1(n_1766),
.A2(n_407),
.B(n_401),
.Y(n_1892)
);

OAI21xp5_ASAP7_75t_L g1893 ( 
.A1(n_1739),
.A2(n_414),
.B(n_410),
.Y(n_1893)
);

BUFx6f_ASAP7_75t_L g1894 ( 
.A(n_1656),
.Y(n_1894)
);

OAI21xp5_ASAP7_75t_L g1895 ( 
.A1(n_1744),
.A2(n_421),
.B(n_420),
.Y(n_1895)
);

AOI21xp5_ASAP7_75t_L g1896 ( 
.A1(n_1524),
.A2(n_424),
.B(n_422),
.Y(n_1896)
);

NAND2xp5_ASAP7_75t_L g1897 ( 
.A(n_1514),
.B(n_1573),
.Y(n_1897)
);

NAND2xp5_ASAP7_75t_L g1898 ( 
.A(n_1611),
.B(n_32),
.Y(n_1898)
);

NAND2xp5_ASAP7_75t_L g1899 ( 
.A(n_1517),
.B(n_1748),
.Y(n_1899)
);

NOR2xp33_ASAP7_75t_L g1900 ( 
.A(n_1696),
.B(n_33),
.Y(n_1900)
);

OAI21xp5_ASAP7_75t_L g1901 ( 
.A1(n_1678),
.A2(n_431),
.B(n_430),
.Y(n_1901)
);

INVx1_ASAP7_75t_L g1902 ( 
.A(n_1694),
.Y(n_1902)
);

AND3x2_ASAP7_75t_L g1903 ( 
.A(n_1742),
.B(n_34),
.C(n_35),
.Y(n_1903)
);

NAND2xp5_ASAP7_75t_L g1904 ( 
.A(n_1750),
.B(n_35),
.Y(n_1904)
);

AOI21xp5_ASAP7_75t_L g1905 ( 
.A1(n_1614),
.A2(n_433),
.B(n_432),
.Y(n_1905)
);

INVx11_ASAP7_75t_L g1906 ( 
.A(n_1638),
.Y(n_1906)
);

NOR2xp33_ASAP7_75t_L g1907 ( 
.A(n_1696),
.B(n_36),
.Y(n_1907)
);

OAI21xp5_ASAP7_75t_L g1908 ( 
.A1(n_1683),
.A2(n_439),
.B(n_437),
.Y(n_1908)
);

OAI21xp5_ASAP7_75t_L g1909 ( 
.A1(n_1684),
.A2(n_441),
.B(n_440),
.Y(n_1909)
);

OAI21xp5_ASAP7_75t_L g1910 ( 
.A1(n_1701),
.A2(n_445),
.B(n_442),
.Y(n_1910)
);

OAI21xp5_ASAP7_75t_L g1911 ( 
.A1(n_1704),
.A2(n_450),
.B(n_447),
.Y(n_1911)
);

AOI21xp5_ASAP7_75t_L g1912 ( 
.A1(n_1619),
.A2(n_453),
.B(n_451),
.Y(n_1912)
);

NAND2xp5_ASAP7_75t_L g1913 ( 
.A(n_1695),
.B(n_37),
.Y(n_1913)
);

O2A1O1Ixp5_ASAP7_75t_L g1914 ( 
.A1(n_1681),
.A2(n_1770),
.B(n_1720),
.C(n_1725),
.Y(n_1914)
);

OAI22xp5_ASAP7_75t_L g1915 ( 
.A1(n_1685),
.A2(n_40),
.B1(n_38),
.B2(n_39),
.Y(n_1915)
);

A2O1A1Ixp33_ASAP7_75t_L g1916 ( 
.A1(n_1784),
.A2(n_41),
.B(n_38),
.C(n_39),
.Y(n_1916)
);

AOI22xp5_ASAP7_75t_L g1917 ( 
.A1(n_1713),
.A2(n_1742),
.B1(n_1719),
.B2(n_1685),
.Y(n_1917)
);

INVx2_ASAP7_75t_L g1918 ( 
.A(n_1616),
.Y(n_1918)
);

NOR2xp67_ASAP7_75t_L g1919 ( 
.A(n_1758),
.B(n_42),
.Y(n_1919)
);

NOR2xp33_ASAP7_75t_L g1920 ( 
.A(n_1697),
.B(n_42),
.Y(n_1920)
);

HB1xp67_ASAP7_75t_L g1921 ( 
.A(n_1589),
.Y(n_1921)
);

NAND2xp5_ASAP7_75t_L g1922 ( 
.A(n_1702),
.B(n_44),
.Y(n_1922)
);

NAND2xp5_ASAP7_75t_L g1923 ( 
.A(n_1703),
.B(n_45),
.Y(n_1923)
);

AOI21xp5_ASAP7_75t_L g1924 ( 
.A1(n_1598),
.A2(n_1698),
.B(n_1693),
.Y(n_1924)
);

NAND2xp5_ASAP7_75t_SL g1925 ( 
.A(n_1589),
.B(n_45),
.Y(n_1925)
);

NAND2xp5_ASAP7_75t_L g1926 ( 
.A(n_1709),
.B(n_48),
.Y(n_1926)
);

NAND2xp5_ASAP7_75t_L g1927 ( 
.A(n_1712),
.B(n_51),
.Y(n_1927)
);

INVx2_ASAP7_75t_L g1928 ( 
.A(n_1628),
.Y(n_1928)
);

NAND2xp5_ASAP7_75t_SL g1929 ( 
.A(n_1777),
.B(n_52),
.Y(n_1929)
);

AND2x2_ASAP7_75t_L g1930 ( 
.A(n_1724),
.B(n_52),
.Y(n_1930)
);

INVx2_ASAP7_75t_L g1931 ( 
.A(n_1637),
.Y(n_1931)
);

OAI21xp5_ASAP7_75t_L g1932 ( 
.A1(n_1718),
.A2(n_460),
.B(n_457),
.Y(n_1932)
);

OAI21xp5_ASAP7_75t_L g1933 ( 
.A1(n_1727),
.A2(n_463),
.B(n_462),
.Y(n_1933)
);

NAND2xp5_ASAP7_75t_L g1934 ( 
.A(n_1714),
.B(n_53),
.Y(n_1934)
);

NAND2xp5_ASAP7_75t_L g1935 ( 
.A(n_1721),
.B(n_53),
.Y(n_1935)
);

BUFx3_ASAP7_75t_L g1936 ( 
.A(n_1538),
.Y(n_1936)
);

AOI21xp5_ASAP7_75t_L g1937 ( 
.A1(n_1705),
.A2(n_465),
.B(n_464),
.Y(n_1937)
);

OAI21xp5_ASAP7_75t_L g1938 ( 
.A1(n_1730),
.A2(n_470),
.B(n_467),
.Y(n_1938)
);

NAND2xp5_ASAP7_75t_L g1939 ( 
.A(n_1722),
.B(n_1723),
.Y(n_1939)
);

NAND2xp5_ASAP7_75t_L g1940 ( 
.A(n_1767),
.B(n_54),
.Y(n_1940)
);

NAND2xp5_ASAP7_75t_SL g1941 ( 
.A(n_1601),
.B(n_1630),
.Y(n_1941)
);

NAND2xp5_ASAP7_75t_L g1942 ( 
.A(n_1626),
.B(n_55),
.Y(n_1942)
);

AND2x2_ASAP7_75t_L g1943 ( 
.A(n_1726),
.B(n_55),
.Y(n_1943)
);

AOI21xp5_ASAP7_75t_L g1944 ( 
.A1(n_1707),
.A2(n_480),
.B(n_479),
.Y(n_1944)
);

BUFx3_ASAP7_75t_L g1945 ( 
.A(n_1682),
.Y(n_1945)
);

AOI22xp5_ASAP7_75t_L g1946 ( 
.A1(n_1713),
.A2(n_59),
.B1(n_56),
.B2(n_58),
.Y(n_1946)
);

NAND2xp5_ASAP7_75t_SL g1947 ( 
.A(n_1601),
.B(n_56),
.Y(n_1947)
);

NAND2xp5_ASAP7_75t_L g1948 ( 
.A(n_1626),
.B(n_58),
.Y(n_1948)
);

AOI21xp5_ASAP7_75t_L g1949 ( 
.A1(n_1731),
.A2(n_483),
.B(n_481),
.Y(n_1949)
);

NAND2xp5_ASAP7_75t_L g1950 ( 
.A(n_1640),
.B(n_61),
.Y(n_1950)
);

AOI21xp5_ASAP7_75t_L g1951 ( 
.A1(n_1735),
.A2(n_487),
.B(n_486),
.Y(n_1951)
);

INVx1_ASAP7_75t_L g1952 ( 
.A(n_1553),
.Y(n_1952)
);

INVx2_ASAP7_75t_L g1953 ( 
.A(n_1733),
.Y(n_1953)
);

BUFx3_ASAP7_75t_L g1954 ( 
.A(n_1773),
.Y(n_1954)
);

NAND2xp5_ASAP7_75t_L g1955 ( 
.A(n_1593),
.B(n_61),
.Y(n_1955)
);

NAND3xp33_ASAP7_75t_L g1956 ( 
.A(n_1664),
.B(n_62),
.C(n_63),
.Y(n_1956)
);

AOI21xp5_ASAP7_75t_L g1957 ( 
.A1(n_1737),
.A2(n_489),
.B(n_488),
.Y(n_1957)
);

NAND2xp5_ASAP7_75t_L g1958 ( 
.A(n_1612),
.B(n_62),
.Y(n_1958)
);

NAND2xp5_ASAP7_75t_L g1959 ( 
.A(n_1620),
.B(n_63),
.Y(n_1959)
);

INVx1_ASAP7_75t_L g1960 ( 
.A(n_1776),
.Y(n_1960)
);

BUFx12f_ASAP7_75t_L g1961 ( 
.A(n_1621),
.Y(n_1961)
);

NAND2xp5_ASAP7_75t_SL g1962 ( 
.A(n_1630),
.B(n_1642),
.Y(n_1962)
);

OAI21xp5_ASAP7_75t_L g1963 ( 
.A1(n_1745),
.A2(n_1780),
.B(n_1772),
.Y(n_1963)
);

NAND2xp5_ASAP7_75t_L g1964 ( 
.A(n_1645),
.B(n_64),
.Y(n_1964)
);

INVx1_ASAP7_75t_L g1965 ( 
.A(n_1760),
.Y(n_1965)
);

INVx1_ASAP7_75t_L g1966 ( 
.A(n_1769),
.Y(n_1966)
);

NAND2xp5_ASAP7_75t_L g1967 ( 
.A(n_1645),
.B(n_64),
.Y(n_1967)
);

NAND2xp5_ASAP7_75t_L g1968 ( 
.A(n_1543),
.B(n_65),
.Y(n_1968)
);

NAND2xp5_ASAP7_75t_L g1969 ( 
.A(n_1642),
.B(n_65),
.Y(n_1969)
);

O2A1O1Ixp33_ASAP7_75t_L g1970 ( 
.A1(n_1595),
.A2(n_68),
.B(n_66),
.C(n_67),
.Y(n_1970)
);

AOI21xp5_ASAP7_75t_L g1971 ( 
.A1(n_1656),
.A2(n_515),
.B(n_514),
.Y(n_1971)
);

NAND2xp5_ASAP7_75t_L g1972 ( 
.A(n_1530),
.B(n_67),
.Y(n_1972)
);

AND2x6_ASAP7_75t_L g1973 ( 
.A(n_1656),
.B(n_516),
.Y(n_1973)
);

NAND2xp5_ASAP7_75t_L g1974 ( 
.A(n_1594),
.B(n_68),
.Y(n_1974)
);

INVx4_ASAP7_75t_L g1975 ( 
.A(n_1519),
.Y(n_1975)
);

NAND2xp5_ASAP7_75t_L g1976 ( 
.A(n_1546),
.B(n_69),
.Y(n_1976)
);

AND2x2_ASAP7_75t_L g1977 ( 
.A(n_1617),
.B(n_69),
.Y(n_1977)
);

NAND2xp5_ASAP7_75t_SL g1978 ( 
.A(n_1785),
.B(n_1567),
.Y(n_1978)
);

O2A1O1Ixp5_ASAP7_75t_L g1979 ( 
.A1(n_1716),
.A2(n_518),
.B(n_520),
.C(n_517),
.Y(n_1979)
);

O2A1O1Ixp33_ASAP7_75t_L g1980 ( 
.A1(n_1523),
.A2(n_1615),
.B(n_1554),
.C(n_1564),
.Y(n_1980)
);

NOR3xp33_ASAP7_75t_L g1981 ( 
.A(n_1634),
.B(n_70),
.C(n_72),
.Y(n_1981)
);

NAND2xp5_ASAP7_75t_L g1982 ( 
.A(n_1547),
.B(n_72),
.Y(n_1982)
);

NAND2xp5_ASAP7_75t_L g1983 ( 
.A(n_1551),
.B(n_73),
.Y(n_1983)
);

AOI21xp5_ASAP7_75t_L g1984 ( 
.A1(n_1655),
.A2(n_523),
.B(n_521),
.Y(n_1984)
);

NAND2xp5_ASAP7_75t_L g1985 ( 
.A(n_1632),
.B(n_74),
.Y(n_1985)
);

A2O1A1Ixp33_ASAP7_75t_L g1986 ( 
.A1(n_1790),
.A2(n_77),
.B(n_74),
.C(n_75),
.Y(n_1986)
);

INVx1_ASAP7_75t_L g1987 ( 
.A(n_1673),
.Y(n_1987)
);

AOI21xp5_ASAP7_75t_L g1988 ( 
.A1(n_1658),
.A2(n_527),
.B(n_525),
.Y(n_1988)
);

NAND2xp5_ASAP7_75t_L g1989 ( 
.A(n_1560),
.B(n_78),
.Y(n_1989)
);

NAND2xp5_ASAP7_75t_L g1990 ( 
.A(n_1563),
.B(n_80),
.Y(n_1990)
);

AOI21xp5_ASAP7_75t_L g1991 ( 
.A1(n_1660),
.A2(n_530),
.B(n_529),
.Y(n_1991)
);

OAI21xp5_ASAP7_75t_L g1992 ( 
.A1(n_1768),
.A2(n_532),
.B(n_531),
.Y(n_1992)
);

AOI21xp5_ASAP7_75t_L g1993 ( 
.A1(n_1666),
.A2(n_1691),
.B(n_1674),
.Y(n_1993)
);

NAND2xp5_ASAP7_75t_L g1994 ( 
.A(n_1569),
.B(n_80),
.Y(n_1994)
);

NAND2xp5_ASAP7_75t_L g1995 ( 
.A(n_1574),
.B(n_81),
.Y(n_1995)
);

AND2x2_ASAP7_75t_L g1996 ( 
.A(n_1617),
.B(n_82),
.Y(n_1996)
);

NAND2xp5_ASAP7_75t_L g1997 ( 
.A(n_1575),
.B(n_82),
.Y(n_1997)
);

AOI21xp5_ASAP7_75t_L g1998 ( 
.A1(n_1759),
.A2(n_536),
.B(n_534),
.Y(n_1998)
);

NOR2xp33_ASAP7_75t_L g1999 ( 
.A(n_1697),
.B(n_83),
.Y(n_1999)
);

OAI21xp5_ASAP7_75t_L g2000 ( 
.A1(n_1643),
.A2(n_539),
.B(n_537),
.Y(n_2000)
);

NOR2xp67_ASAP7_75t_L g2001 ( 
.A(n_1590),
.B(n_84),
.Y(n_2001)
);

INVx2_ASAP7_75t_SL g2002 ( 
.A(n_1671),
.Y(n_2002)
);

INVx2_ASAP7_75t_L g2003 ( 
.A(n_1644),
.Y(n_2003)
);

AOI21xp5_ASAP7_75t_L g2004 ( 
.A1(n_1584),
.A2(n_543),
.B(n_541),
.Y(n_2004)
);

INVx1_ASAP7_75t_L g2005 ( 
.A(n_1677),
.Y(n_2005)
);

NAND2xp5_ASAP7_75t_L g2006 ( 
.A(n_1578),
.B(n_84),
.Y(n_2006)
);

NOR2xp33_ASAP7_75t_SL g2007 ( 
.A(n_1519),
.B(n_85),
.Y(n_2007)
);

BUFx3_ASAP7_75t_L g2008 ( 
.A(n_1625),
.Y(n_2008)
);

AO21x1_ASAP7_75t_L g2009 ( 
.A1(n_1787),
.A2(n_548),
.B(n_547),
.Y(n_2009)
);

AND2x2_ASAP7_75t_L g2010 ( 
.A(n_1646),
.B(n_1670),
.Y(n_2010)
);

INVxp67_ASAP7_75t_L g2011 ( 
.A(n_1646),
.Y(n_2011)
);

NAND2xp5_ASAP7_75t_L g2012 ( 
.A(n_1567),
.B(n_86),
.Y(n_2012)
);

NAND2xp5_ASAP7_75t_L g2013 ( 
.A(n_1729),
.B(n_1700),
.Y(n_2013)
);

NAND2xp5_ASAP7_75t_L g2014 ( 
.A(n_1729),
.B(n_87),
.Y(n_2014)
);

AO21x1_ASAP7_75t_L g2015 ( 
.A1(n_1783),
.A2(n_553),
.B(n_551),
.Y(n_2015)
);

INVx1_ASAP7_75t_L g2016 ( 
.A(n_1688),
.Y(n_2016)
);

NAND2xp5_ASAP7_75t_L g2017 ( 
.A(n_1700),
.B(n_87),
.Y(n_2017)
);

INVx2_ASAP7_75t_L g2018 ( 
.A(n_1647),
.Y(n_2018)
);

INVx2_ASAP7_75t_SL g2019 ( 
.A(n_1671),
.Y(n_2019)
);

AOI21xp5_ASAP7_75t_L g2020 ( 
.A1(n_1771),
.A2(n_554),
.B(n_89),
.Y(n_2020)
);

O2A1O1Ixp33_ASAP7_75t_L g2021 ( 
.A1(n_1604),
.A2(n_92),
.B(n_89),
.C(n_90),
.Y(n_2021)
);

BUFx4f_ASAP7_75t_L g2022 ( 
.A(n_1778),
.Y(n_2022)
);

AOI21xp5_ASAP7_75t_L g2023 ( 
.A1(n_1779),
.A2(n_90),
.B(n_92),
.Y(n_2023)
);

NAND2xp5_ASAP7_75t_L g2024 ( 
.A(n_1605),
.B(n_93),
.Y(n_2024)
);

INVx1_ASAP7_75t_L g2025 ( 
.A(n_1688),
.Y(n_2025)
);

INVx1_ASAP7_75t_L g2026 ( 
.A(n_1688),
.Y(n_2026)
);

OAI21xp5_ASAP7_75t_L g2027 ( 
.A1(n_1648),
.A2(n_94),
.B(n_95),
.Y(n_2027)
);

NAND2xp5_ASAP7_75t_L g2028 ( 
.A(n_1608),
.B(n_95),
.Y(n_2028)
);

INVx5_ASAP7_75t_L g2029 ( 
.A(n_1778),
.Y(n_2029)
);

OAI21xp5_ASAP7_75t_L g2030 ( 
.A1(n_1650),
.A2(n_96),
.B(n_97),
.Y(n_2030)
);

OAI21xp33_ASAP7_75t_L g2031 ( 
.A1(n_1663),
.A2(n_97),
.B(n_98),
.Y(n_2031)
);

INVx2_ASAP7_75t_L g2032 ( 
.A(n_1665),
.Y(n_2032)
);

BUFx2_ASAP7_75t_L g2033 ( 
.A(n_1778),
.Y(n_2033)
);

NAND2xp5_ASAP7_75t_L g2034 ( 
.A(n_1775),
.B(n_98),
.Y(n_2034)
);

NAND2xp5_ASAP7_75t_L g2035 ( 
.A(n_1775),
.B(n_99),
.Y(n_2035)
);

BUFx3_ASAP7_75t_L g2036 ( 
.A(n_1582),
.Y(n_2036)
);

O2A1O1Ixp5_ASAP7_75t_L g2037 ( 
.A1(n_1720),
.A2(n_105),
.B(n_103),
.C(n_104),
.Y(n_2037)
);

AOI21xp5_ASAP7_75t_L g2038 ( 
.A1(n_1556),
.A2(n_107),
.B(n_108),
.Y(n_2038)
);

AOI21xp5_ASAP7_75t_L g2039 ( 
.A1(n_1557),
.A2(n_107),
.B(n_109),
.Y(n_2039)
);

INVx3_ASAP7_75t_L g2040 ( 
.A(n_1649),
.Y(n_2040)
);

BUFx2_ASAP7_75t_SL g2041 ( 
.A(n_1743),
.Y(n_2041)
);

NAND2xp5_ASAP7_75t_L g2042 ( 
.A(n_1511),
.B(n_109),
.Y(n_2042)
);

OR2x2_ASAP7_75t_L g2043 ( 
.A(n_1710),
.B(n_110),
.Y(n_2043)
);

NAND3xp33_ASAP7_75t_SL g2044 ( 
.A(n_1664),
.B(n_110),
.C(n_111),
.Y(n_2044)
);

NAND2xp5_ASAP7_75t_L g2045 ( 
.A(n_1529),
.B(n_111),
.Y(n_2045)
);

INVx1_ASAP7_75t_L g2046 ( 
.A(n_1774),
.Y(n_2046)
);

INVx1_ASAP7_75t_L g2047 ( 
.A(n_1774),
.Y(n_2047)
);

NAND2xp5_ASAP7_75t_SL g2048 ( 
.A(n_1657),
.B(n_112),
.Y(n_2048)
);

AND2x2_ASAP7_75t_L g2049 ( 
.A(n_1663),
.B(n_112),
.Y(n_2049)
);

AOI21xp5_ASAP7_75t_L g2050 ( 
.A1(n_1753),
.A2(n_113),
.B(n_114),
.Y(n_2050)
);

NAND2xp5_ASAP7_75t_L g2051 ( 
.A(n_1566),
.B(n_1570),
.Y(n_2051)
);

OAI22xp5_ASAP7_75t_L g2052 ( 
.A1(n_1774),
.A2(n_117),
.B1(n_115),
.B2(n_116),
.Y(n_2052)
);

HB1xp67_ASAP7_75t_L g2053 ( 
.A(n_1661),
.Y(n_2053)
);

BUFx2_ASAP7_75t_L g2054 ( 
.A(n_1603),
.Y(n_2054)
);

OAI21xp5_ASAP7_75t_L g2055 ( 
.A1(n_1662),
.A2(n_116),
.B(n_118),
.Y(n_2055)
);

AOI21xp5_ASAP7_75t_L g2056 ( 
.A1(n_1746),
.A2(n_119),
.B(n_120),
.Y(n_2056)
);

AOI21xp5_ASAP7_75t_L g2057 ( 
.A1(n_1610),
.A2(n_123),
.B(n_125),
.Y(n_2057)
);

INVx1_ASAP7_75t_L g2058 ( 
.A(n_1581),
.Y(n_2058)
);

INVx2_ASAP7_75t_L g2059 ( 
.A(n_1741),
.Y(n_2059)
);

AOI21xp5_ASAP7_75t_L g2060 ( 
.A1(n_1782),
.A2(n_123),
.B(n_125),
.Y(n_2060)
);

NAND2xp5_ASAP7_75t_L g2061 ( 
.A(n_1587),
.B(n_126),
.Y(n_2061)
);

NAND2xp5_ASAP7_75t_L g2062 ( 
.A(n_1667),
.B(n_126),
.Y(n_2062)
);

NAND2xp5_ASAP7_75t_L g2063 ( 
.A(n_1699),
.B(n_132),
.Y(n_2063)
);

NAND2xp5_ASAP7_75t_L g2064 ( 
.A(n_1699),
.B(n_133),
.Y(n_2064)
);

INVx3_ASAP7_75t_L g2065 ( 
.A(n_1657),
.Y(n_2065)
);

BUFx8_ASAP7_75t_L g2066 ( 
.A(n_1743),
.Y(n_2066)
);

NOR2xp33_ASAP7_75t_L g2067 ( 
.A(n_1708),
.B(n_133),
.Y(n_2067)
);

BUFx6f_ASAP7_75t_L g2068 ( 
.A(n_1623),
.Y(n_2068)
);

AOI21xp5_ASAP7_75t_L g2069 ( 
.A1(n_1725),
.A2(n_134),
.B(n_135),
.Y(n_2069)
);

NAND2xp5_ASAP7_75t_L g2070 ( 
.A(n_1667),
.B(n_134),
.Y(n_2070)
);

NAND2xp5_ASAP7_75t_SL g2071 ( 
.A(n_1676),
.B(n_136),
.Y(n_2071)
);

INVx1_ASAP7_75t_L g2072 ( 
.A(n_1622),
.Y(n_2072)
);

OR2x2_ASAP7_75t_L g2073 ( 
.A(n_1708),
.B(n_136),
.Y(n_2073)
);

OAI21xp5_ASAP7_75t_L g2074 ( 
.A1(n_1762),
.A2(n_138),
.B(n_139),
.Y(n_2074)
);

OAI22xp5_ASAP7_75t_L g2075 ( 
.A1(n_1686),
.A2(n_142),
.B1(n_140),
.B2(n_141),
.Y(n_2075)
);

NAND2xp5_ASAP7_75t_L g2076 ( 
.A(n_1715),
.B(n_141),
.Y(n_2076)
);

NAND2xp5_ASAP7_75t_SL g2077 ( 
.A(n_1752),
.B(n_142),
.Y(n_2077)
);

INVx2_ASAP7_75t_L g2078 ( 
.A(n_1741),
.Y(n_2078)
);

NAND2x1p5_ASAP7_75t_L g2079 ( 
.A(n_1689),
.B(n_143),
.Y(n_2079)
);

A2O1A1Ixp33_ASAP7_75t_L g2080 ( 
.A1(n_1749),
.A2(n_1763),
.B(n_1555),
.C(n_1597),
.Y(n_2080)
);

NAND2xp5_ASAP7_75t_L g2081 ( 
.A(n_1715),
.B(n_143),
.Y(n_2081)
);

OAI21xp5_ASAP7_75t_L g2082 ( 
.A1(n_1749),
.A2(n_145),
.B(n_146),
.Y(n_2082)
);

CKINVDCx10_ASAP7_75t_R g2083 ( 
.A(n_1613),
.Y(n_2083)
);

INVx1_ASAP7_75t_L g2084 ( 
.A(n_1689),
.Y(n_2084)
);

A2O1A1Ixp33_ASAP7_75t_L g2085 ( 
.A1(n_1540),
.A2(n_149),
.B(n_147),
.C(n_148),
.Y(n_2085)
);

NAND2xp5_ASAP7_75t_L g2086 ( 
.A(n_1599),
.B(n_152),
.Y(n_2086)
);

A2O1A1Ixp33_ASAP7_75t_L g2087 ( 
.A1(n_1540),
.A2(n_155),
.B(n_153),
.C(n_154),
.Y(n_2087)
);

NAND3xp33_ASAP7_75t_SL g2088 ( 
.A(n_1761),
.B(n_154),
.C(n_157),
.Y(n_2088)
);

BUFx6f_ASAP7_75t_L g2089 ( 
.A(n_1623),
.Y(n_2089)
);

AND2x2_ASAP7_75t_L g2090 ( 
.A(n_1736),
.B(n_159),
.Y(n_2090)
);

AND2x2_ASAP7_75t_L g2091 ( 
.A(n_1692),
.B(n_159),
.Y(n_2091)
);

NAND2xp5_ASAP7_75t_L g2092 ( 
.A(n_1639),
.B(n_160),
.Y(n_2092)
);

NOR2xp33_ASAP7_75t_L g2093 ( 
.A(n_1555),
.B(n_160),
.Y(n_2093)
);

AOI21xp5_ASAP7_75t_L g2094 ( 
.A1(n_1728),
.A2(n_161),
.B(n_163),
.Y(n_2094)
);

NAND2xp5_ASAP7_75t_L g2095 ( 
.A(n_1639),
.B(n_163),
.Y(n_2095)
);

AOI21xp5_ASAP7_75t_L g2096 ( 
.A1(n_1732),
.A2(n_164),
.B(n_165),
.Y(n_2096)
);

NAND2xp5_ASAP7_75t_L g2097 ( 
.A(n_1597),
.B(n_165),
.Y(n_2097)
);

NAND2xp5_ASAP7_75t_L g2098 ( 
.A(n_1639),
.B(n_166),
.Y(n_2098)
);

OAI22xp5_ASAP7_75t_L g2099 ( 
.A1(n_1686),
.A2(n_166),
.B1(n_167),
.B2(n_168),
.Y(n_2099)
);

AOI22xp5_ASAP7_75t_L g2100 ( 
.A1(n_1639),
.A2(n_168),
.B1(n_170),
.B2(n_171),
.Y(n_2100)
);

AND2x2_ASAP7_75t_L g2101 ( 
.A(n_1842),
.B(n_170),
.Y(n_2101)
);

NAND2xp5_ASAP7_75t_L g2102 ( 
.A(n_1862),
.B(n_1751),
.Y(n_2102)
);

NOR2xp33_ASAP7_75t_L g2103 ( 
.A(n_2011),
.B(n_1732),
.Y(n_2103)
);

INVx1_ASAP7_75t_L g2104 ( 
.A(n_1818),
.Y(n_2104)
);

NOR2xp33_ASAP7_75t_R g2105 ( 
.A(n_1867),
.B(n_1576),
.Y(n_2105)
);

AOI21xp33_ASAP7_75t_L g2106 ( 
.A1(n_1980),
.A2(n_1738),
.B(n_1734),
.Y(n_2106)
);

A2O1A1Ixp33_ASAP7_75t_L g2107 ( 
.A1(n_1993),
.A2(n_1747),
.B(n_1751),
.C(n_1690),
.Y(n_2107)
);

OA22x2_ASAP7_75t_L g2108 ( 
.A1(n_1917),
.A2(n_1903),
.B1(n_2053),
.B2(n_1946),
.Y(n_2108)
);

OR2x6_ASAP7_75t_L g2109 ( 
.A(n_1827),
.B(n_1602),
.Y(n_2109)
);

AOI21xp5_ASAP7_75t_L g2110 ( 
.A1(n_1858),
.A2(n_1754),
.B(n_1740),
.Y(n_2110)
);

AOI22xp33_ASAP7_75t_L g2111 ( 
.A1(n_2010),
.A2(n_1874),
.B1(n_1812),
.B2(n_1830),
.Y(n_2111)
);

INVx3_ASAP7_75t_L g2112 ( 
.A(n_2022),
.Y(n_2112)
);

NAND3xp33_ASAP7_75t_SL g2113 ( 
.A(n_2007),
.B(n_1754),
.C(n_1740),
.Y(n_2113)
);

NOR2xp33_ASAP7_75t_L g2114 ( 
.A(n_1822),
.B(n_1755),
.Y(n_2114)
);

NAND3xp33_ASAP7_75t_SL g2115 ( 
.A(n_1811),
.B(n_1883),
.C(n_1970),
.Y(n_2115)
);

INVx1_ASAP7_75t_L g2116 ( 
.A(n_1819),
.Y(n_2116)
);

BUFx12f_ASAP7_75t_L g2117 ( 
.A(n_1852),
.Y(n_2117)
);

NAND2xp5_ASAP7_75t_SL g2118 ( 
.A(n_2022),
.B(n_1623),
.Y(n_2118)
);

BUFx10_ASAP7_75t_L g2119 ( 
.A(n_1861),
.Y(n_2119)
);

INVxp67_ASAP7_75t_L g2120 ( 
.A(n_1802),
.Y(n_2120)
);

NAND2x1p5_ASAP7_75t_L g2121 ( 
.A(n_1841),
.B(n_1623),
.Y(n_2121)
);

BUFx2_ASAP7_75t_L g2122 ( 
.A(n_1961),
.Y(n_2122)
);

AOI21xp5_ASAP7_75t_L g2123 ( 
.A1(n_1844),
.A2(n_1764),
.B(n_1755),
.Y(n_2123)
);

NOR3xp33_ASAP7_75t_L g2124 ( 
.A(n_2088),
.B(n_1717),
.C(n_1690),
.Y(n_2124)
);

NAND2xp5_ASAP7_75t_SL g2125 ( 
.A(n_2029),
.B(n_1629),
.Y(n_2125)
);

NAND2xp5_ASAP7_75t_L g2126 ( 
.A(n_1831),
.B(n_1717),
.Y(n_2126)
);

NAND2xp5_ASAP7_75t_SL g2127 ( 
.A(n_2029),
.B(n_1800),
.Y(n_2127)
);

BUFx4_ASAP7_75t_SL g2128 ( 
.A(n_1825),
.Y(n_2128)
);

BUFx3_ASAP7_75t_L g2129 ( 
.A(n_2066),
.Y(n_2129)
);

INVx1_ASAP7_75t_L g2130 ( 
.A(n_1839),
.Y(n_2130)
);

NOR2xp33_ASAP7_75t_L g2131 ( 
.A(n_1854),
.B(n_1602),
.Y(n_2131)
);

NOR2xp33_ASAP7_75t_L g2132 ( 
.A(n_1809),
.B(n_1629),
.Y(n_2132)
);

NAND2xp5_ASAP7_75t_L g2133 ( 
.A(n_1800),
.B(n_1629),
.Y(n_2133)
);

INVx2_ASAP7_75t_SL g2134 ( 
.A(n_1906),
.Y(n_2134)
);

BUFx6f_ASAP7_75t_L g2135 ( 
.A(n_1796),
.Y(n_2135)
);

NAND2xp5_ASAP7_75t_L g2136 ( 
.A(n_1952),
.B(n_2072),
.Y(n_2136)
);

INVx1_ASAP7_75t_L g2137 ( 
.A(n_1850),
.Y(n_2137)
);

AOI22xp5_ASAP7_75t_L g2138 ( 
.A1(n_1835),
.A2(n_1675),
.B1(n_1792),
.B2(n_1781),
.Y(n_2138)
);

CKINVDCx5p33_ASAP7_75t_R g2139 ( 
.A(n_2066),
.Y(n_2139)
);

NAND2xp5_ASAP7_75t_L g2140 ( 
.A(n_1804),
.B(n_1675),
.Y(n_2140)
);

INVx2_ASAP7_75t_SL g2141 ( 
.A(n_1841),
.Y(n_2141)
);

O2A1O1Ixp33_ASAP7_75t_L g2142 ( 
.A1(n_1821),
.A2(n_1675),
.B(n_173),
.C(n_174),
.Y(n_2142)
);

AND2x4_ASAP7_75t_L g2143 ( 
.A(n_1836),
.B(n_1675),
.Y(n_2143)
);

AOI21xp5_ASAP7_75t_L g2144 ( 
.A1(n_1848),
.A2(n_1675),
.B(n_1781),
.Y(n_2144)
);

O2A1O1Ixp33_ASAP7_75t_L g2145 ( 
.A1(n_1889),
.A2(n_171),
.B(n_174),
.C(n_175),
.Y(n_2145)
);

AOI21xp5_ASAP7_75t_L g2146 ( 
.A1(n_1834),
.A2(n_1781),
.B(n_176),
.Y(n_2146)
);

OR2x2_ASAP7_75t_L g2147 ( 
.A(n_1836),
.B(n_1816),
.Y(n_2147)
);

CKINVDCx6p67_ASAP7_75t_R g2148 ( 
.A(n_1945),
.Y(n_2148)
);

NAND3xp33_ASAP7_75t_L g2149 ( 
.A(n_1981),
.B(n_1781),
.C(n_180),
.Y(n_2149)
);

NAND2xp5_ASAP7_75t_SL g2150 ( 
.A(n_2033),
.B(n_180),
.Y(n_2150)
);

NAND2xp5_ASAP7_75t_L g2151 ( 
.A(n_1804),
.B(n_181),
.Y(n_2151)
);

INVx2_ASAP7_75t_L g2152 ( 
.A(n_1810),
.Y(n_2152)
);

BUFx12f_ASAP7_75t_L g2153 ( 
.A(n_1975),
.Y(n_2153)
);

INVx1_ASAP7_75t_L g2154 ( 
.A(n_1813),
.Y(n_2154)
);

OAI21xp5_ASAP7_75t_L g2155 ( 
.A1(n_1857),
.A2(n_182),
.B(n_183),
.Y(n_2155)
);

NAND2xp5_ASAP7_75t_L g2156 ( 
.A(n_1826),
.B(n_183),
.Y(n_2156)
);

NAND2xp5_ASAP7_75t_L g2157 ( 
.A(n_1826),
.B(n_184),
.Y(n_2157)
);

AOI22xp5_ASAP7_75t_L g2158 ( 
.A1(n_2016),
.A2(n_185),
.B1(n_186),
.B2(n_187),
.Y(n_2158)
);

BUFx3_ASAP7_75t_L g2159 ( 
.A(n_1884),
.Y(n_2159)
);

INVx4_ASAP7_75t_L g2160 ( 
.A(n_1884),
.Y(n_2160)
);

NAND2xp5_ASAP7_75t_SL g2161 ( 
.A(n_1843),
.B(n_185),
.Y(n_2161)
);

AND2x2_ASAP7_75t_L g2162 ( 
.A(n_1930),
.B(n_187),
.Y(n_2162)
);

INVx1_ASAP7_75t_L g2163 ( 
.A(n_1828),
.Y(n_2163)
);

INVx2_ASAP7_75t_L g2164 ( 
.A(n_1847),
.Y(n_2164)
);

CKINVDCx5p33_ASAP7_75t_R g2165 ( 
.A(n_2083),
.Y(n_2165)
);

O2A1O1Ixp5_ASAP7_75t_L g2166 ( 
.A1(n_1914),
.A2(n_188),
.B(n_189),
.C(n_191),
.Y(n_2166)
);

INVx1_ASAP7_75t_L g2167 ( 
.A(n_1816),
.Y(n_2167)
);

NOR2xp33_ASAP7_75t_L g2168 ( 
.A(n_2002),
.B(n_2019),
.Y(n_2168)
);

NAND2xp5_ASAP7_75t_L g2169 ( 
.A(n_1939),
.B(n_192),
.Y(n_2169)
);

BUFx6f_ASAP7_75t_L g2170 ( 
.A(n_1796),
.Y(n_2170)
);

INVx1_ASAP7_75t_L g2171 ( 
.A(n_1913),
.Y(n_2171)
);

A2O1A1Ixp33_ASAP7_75t_L g2172 ( 
.A1(n_1924),
.A2(n_192),
.B(n_193),
.C(n_194),
.Y(n_2172)
);

A2O1A1Ixp33_ASAP7_75t_SL g2173 ( 
.A1(n_2074),
.A2(n_193),
.B(n_195),
.C(n_196),
.Y(n_2173)
);

NOR2xp33_ASAP7_75t_L g2174 ( 
.A(n_1859),
.B(n_195),
.Y(n_2174)
);

INVx3_ASAP7_75t_L g2175 ( 
.A(n_1856),
.Y(n_2175)
);

A2O1A1Ixp33_ASAP7_75t_SL g2176 ( 
.A1(n_2055),
.A2(n_196),
.B(n_197),
.C(n_198),
.Y(n_2176)
);

OAI22xp5_ASAP7_75t_SL g2177 ( 
.A1(n_2079),
.A2(n_197),
.B1(n_198),
.B2(n_199),
.Y(n_2177)
);

A2O1A1Ixp33_ASAP7_75t_L g2178 ( 
.A1(n_1833),
.A2(n_199),
.B(n_200),
.C(n_201),
.Y(n_2178)
);

NAND2xp5_ASAP7_75t_L g2179 ( 
.A(n_1939),
.B(n_200),
.Y(n_2179)
);

NAND2xp5_ASAP7_75t_L g2180 ( 
.A(n_1890),
.B(n_1902),
.Y(n_2180)
);

NAND2xp5_ASAP7_75t_SL g2181 ( 
.A(n_1794),
.B(n_1860),
.Y(n_2181)
);

OAI22xp5_ASAP7_75t_L g2182 ( 
.A1(n_2034),
.A2(n_201),
.B1(n_202),
.B2(n_203),
.Y(n_2182)
);

O2A1O1Ixp5_ASAP7_75t_L g2183 ( 
.A1(n_1799),
.A2(n_2080),
.B(n_1814),
.C(n_2035),
.Y(n_2183)
);

NAND2xp5_ASAP7_75t_L g2184 ( 
.A(n_1977),
.B(n_202),
.Y(n_2184)
);

INVx2_ASAP7_75t_L g2185 ( 
.A(n_1918),
.Y(n_2185)
);

AND2x4_ASAP7_75t_L g2186 ( 
.A(n_1827),
.B(n_203),
.Y(n_2186)
);

INVx5_ASAP7_75t_L g2187 ( 
.A(n_1827),
.Y(n_2187)
);

CKINVDCx11_ASAP7_75t_R g2188 ( 
.A(n_1975),
.Y(n_2188)
);

OAI22xp5_ASAP7_75t_SL g2189 ( 
.A1(n_2079),
.A2(n_376),
.B1(n_205),
.B2(n_208),
.Y(n_2189)
);

NAND2xp5_ASAP7_75t_L g2190 ( 
.A(n_1996),
.B(n_204),
.Y(n_2190)
);

O2A1O1Ixp5_ASAP7_75t_L g2191 ( 
.A1(n_2034),
.A2(n_204),
.B(n_208),
.C(n_209),
.Y(n_2191)
);

AOI21xp5_ASAP7_75t_L g2192 ( 
.A1(n_1795),
.A2(n_210),
.B(n_211),
.Y(n_2192)
);

OAI22xp5_ASAP7_75t_L g2193 ( 
.A1(n_2035),
.A2(n_212),
.B1(n_213),
.B2(n_214),
.Y(n_2193)
);

AND2x4_ASAP7_75t_L g2194 ( 
.A(n_1808),
.B(n_212),
.Y(n_2194)
);

AOI21xp5_ASAP7_75t_L g2195 ( 
.A1(n_1798),
.A2(n_214),
.B(n_215),
.Y(n_2195)
);

OR2x6_ASAP7_75t_L g2196 ( 
.A(n_2041),
.B(n_215),
.Y(n_2196)
);

NAND2xp5_ASAP7_75t_L g2197 ( 
.A(n_1943),
.B(n_216),
.Y(n_2197)
);

NAND2xp5_ASAP7_75t_L g2198 ( 
.A(n_2049),
.B(n_217),
.Y(n_2198)
);

AO22x1_ASAP7_75t_L g2199 ( 
.A1(n_2052),
.A2(n_218),
.B1(n_219),
.B2(n_220),
.Y(n_2199)
);

BUFx2_ASAP7_75t_R g2200 ( 
.A(n_1936),
.Y(n_2200)
);

O2A1O1Ixp33_ASAP7_75t_L g2201 ( 
.A1(n_1887),
.A2(n_218),
.B(n_221),
.C(n_222),
.Y(n_2201)
);

O2A1O1Ixp33_ASAP7_75t_L g2202 ( 
.A1(n_1881),
.A2(n_225),
.B(n_226),
.C(n_228),
.Y(n_2202)
);

OAI22xp5_ASAP7_75t_L g2203 ( 
.A1(n_1968),
.A2(n_230),
.B1(n_231),
.B2(n_233),
.Y(n_2203)
);

CKINVDCx5p33_ASAP7_75t_R g2204 ( 
.A(n_1954),
.Y(n_2204)
);

INVx4_ASAP7_75t_L g2205 ( 
.A(n_1861),
.Y(n_2205)
);

NAND2xp5_ASAP7_75t_SL g2206 ( 
.A(n_1863),
.B(n_233),
.Y(n_2206)
);

NAND2xp5_ASAP7_75t_L g2207 ( 
.A(n_1921),
.B(n_234),
.Y(n_2207)
);

BUFx6f_ASAP7_75t_L g2208 ( 
.A(n_1796),
.Y(n_2208)
);

NOR3xp33_ASAP7_75t_SL g2209 ( 
.A(n_2044),
.B(n_236),
.C(n_237),
.Y(n_2209)
);

HB1xp67_ASAP7_75t_L g2210 ( 
.A(n_2008),
.Y(n_2210)
);

NOR2xp33_ASAP7_75t_L g2211 ( 
.A(n_2043),
.B(n_237),
.Y(n_2211)
);

NAND2xp5_ASAP7_75t_L g2212 ( 
.A(n_1968),
.B(n_238),
.Y(n_2212)
);

BUFx6f_ASAP7_75t_L g2213 ( 
.A(n_1832),
.Y(n_2213)
);

BUFx6f_ASAP7_75t_L g2214 ( 
.A(n_1832),
.Y(n_2214)
);

O2A1O1Ixp33_ASAP7_75t_L g2215 ( 
.A1(n_2076),
.A2(n_239),
.B(n_240),
.C(n_241),
.Y(n_2215)
);

NOR2xp33_ASAP7_75t_L g2216 ( 
.A(n_2073),
.B(n_239),
.Y(n_2216)
);

AOI21xp5_ASAP7_75t_L g2217 ( 
.A1(n_1805),
.A2(n_240),
.B(n_241),
.Y(n_2217)
);

INVx1_ASAP7_75t_L g2218 ( 
.A(n_1913),
.Y(n_2218)
);

NAND2xp5_ASAP7_75t_L g2219 ( 
.A(n_1899),
.B(n_1868),
.Y(n_2219)
);

NAND2xp5_ASAP7_75t_L g2220 ( 
.A(n_1899),
.B(n_242),
.Y(n_2220)
);

AOI21xp5_ASAP7_75t_L g2221 ( 
.A1(n_1851),
.A2(n_245),
.B(n_246),
.Y(n_2221)
);

BUFx2_ASAP7_75t_L g2222 ( 
.A(n_2054),
.Y(n_2222)
);

A2O1A1Ixp33_ASAP7_75t_SL g2223 ( 
.A1(n_1900),
.A2(n_248),
.B(n_249),
.C(n_250),
.Y(n_2223)
);

BUFx3_ASAP7_75t_L g2224 ( 
.A(n_2036),
.Y(n_2224)
);

AOI21xp5_ASAP7_75t_L g2225 ( 
.A1(n_1897),
.A2(n_248),
.B(n_249),
.Y(n_2225)
);

AND2x4_ASAP7_75t_L g2226 ( 
.A(n_1962),
.B(n_251),
.Y(n_2226)
);

NAND2xp5_ASAP7_75t_SL g2227 ( 
.A(n_1856),
.B(n_253),
.Y(n_2227)
);

INVx4_ASAP7_75t_L g2228 ( 
.A(n_1797),
.Y(n_2228)
);

A2O1A1Ixp33_ASAP7_75t_SL g2229 ( 
.A1(n_1907),
.A2(n_1999),
.B(n_2067),
.C(n_1920),
.Y(n_2229)
);

INVx2_ASAP7_75t_L g2230 ( 
.A(n_1928),
.Y(n_2230)
);

AND2x4_ASAP7_75t_L g2231 ( 
.A(n_1823),
.B(n_254),
.Y(n_2231)
);

INVx1_ASAP7_75t_L g2232 ( 
.A(n_1922),
.Y(n_2232)
);

OAI22xp5_ASAP7_75t_L g2233 ( 
.A1(n_1960),
.A2(n_254),
.B1(n_255),
.B2(n_256),
.Y(n_2233)
);

AOI22xp33_ASAP7_75t_L g2234 ( 
.A1(n_2090),
.A2(n_255),
.B1(n_256),
.B2(n_257),
.Y(n_2234)
);

BUFx6f_ASAP7_75t_SL g2235 ( 
.A(n_2025),
.Y(n_2235)
);

AOI21xp5_ASAP7_75t_L g2236 ( 
.A1(n_1897),
.A2(n_258),
.B(n_260),
.Y(n_2236)
);

AND2x2_ASAP7_75t_L g2237 ( 
.A(n_1931),
.B(n_261),
.Y(n_2237)
);

NOR2xp33_ASAP7_75t_L g2238 ( 
.A(n_1870),
.B(n_261),
.Y(n_2238)
);

INVx1_ASAP7_75t_L g2239 ( 
.A(n_1922),
.Y(n_2239)
);

INVx2_ASAP7_75t_L g2240 ( 
.A(n_1953),
.Y(n_2240)
);

O2A1O1Ixp33_ASAP7_75t_L g2241 ( 
.A1(n_2076),
.A2(n_262),
.B(n_264),
.C(n_265),
.Y(n_2241)
);

BUFx6f_ASAP7_75t_L g2242 ( 
.A(n_1832),
.Y(n_2242)
);

NAND2xp5_ASAP7_75t_SL g2243 ( 
.A(n_1898),
.B(n_262),
.Y(n_2243)
);

CKINVDCx5p33_ASAP7_75t_R g2244 ( 
.A(n_1915),
.Y(n_2244)
);

NOR2xp67_ASAP7_75t_L g2245 ( 
.A(n_2046),
.B(n_265),
.Y(n_2245)
);

AOI21xp5_ASAP7_75t_L g2246 ( 
.A1(n_1801),
.A2(n_266),
.B(n_267),
.Y(n_2246)
);

OAI21xp33_ASAP7_75t_SL g2247 ( 
.A1(n_1801),
.A2(n_266),
.B(n_267),
.Y(n_2247)
);

O2A1O1Ixp33_ASAP7_75t_L g2248 ( 
.A1(n_2081),
.A2(n_268),
.B(n_269),
.C(n_270),
.Y(n_2248)
);

AOI21xp5_ASAP7_75t_L g2249 ( 
.A1(n_1803),
.A2(n_269),
.B(n_270),
.Y(n_2249)
);

NOR2xp33_ASAP7_75t_R g2250 ( 
.A(n_1797),
.B(n_271),
.Y(n_2250)
);

AND2x2_ASAP7_75t_L g2251 ( 
.A(n_1987),
.B(n_2005),
.Y(n_2251)
);

INVx1_ASAP7_75t_L g2252 ( 
.A(n_1923),
.Y(n_2252)
);

NAND2xp5_ASAP7_75t_L g2253 ( 
.A(n_1974),
.B(n_272),
.Y(n_2253)
);

INVx1_ASAP7_75t_L g2254 ( 
.A(n_1923),
.Y(n_2254)
);

NOR3xp33_ASAP7_75t_SL g2255 ( 
.A(n_1956),
.B(n_275),
.C(n_277),
.Y(n_2255)
);

INVx2_ASAP7_75t_L g2256 ( 
.A(n_2003),
.Y(n_2256)
);

NOR2xp33_ASAP7_75t_R g2257 ( 
.A(n_1806),
.B(n_277),
.Y(n_2257)
);

INVxp67_ASAP7_75t_SL g2258 ( 
.A(n_1879),
.Y(n_2258)
);

INVx1_ASAP7_75t_L g2259 ( 
.A(n_1926),
.Y(n_2259)
);

O2A1O1Ixp33_ASAP7_75t_SL g2260 ( 
.A1(n_1878),
.A2(n_1873),
.B(n_1941),
.C(n_1815),
.Y(n_2260)
);

INVx4_ASAP7_75t_L g2261 ( 
.A(n_1806),
.Y(n_2261)
);

NOR2xp33_ASAP7_75t_L g2262 ( 
.A(n_2081),
.B(n_278),
.Y(n_2262)
);

OAI21xp5_ASAP7_75t_L g2263 ( 
.A1(n_1820),
.A2(n_279),
.B(n_281),
.Y(n_2263)
);

AOI22xp5_ASAP7_75t_L g2264 ( 
.A1(n_2026),
.A2(n_1898),
.B1(n_2047),
.B2(n_1985),
.Y(n_2264)
);

AOI21xp5_ASAP7_75t_L g2265 ( 
.A1(n_1803),
.A2(n_281),
.B(n_282),
.Y(n_2265)
);

NAND2xp5_ASAP7_75t_SL g2266 ( 
.A(n_1919),
.B(n_283),
.Y(n_2266)
);

NAND2xp5_ASAP7_75t_SL g2267 ( 
.A(n_1866),
.B(n_284),
.Y(n_2267)
);

NAND2xp5_ASAP7_75t_SL g2268 ( 
.A(n_2068),
.B(n_285),
.Y(n_2268)
);

BUFx6f_ASAP7_75t_L g2269 ( 
.A(n_1837),
.Y(n_2269)
);

AND2x2_ASAP7_75t_L g2270 ( 
.A(n_1964),
.B(n_287),
.Y(n_2270)
);

NOR2xp33_ASAP7_75t_L g2271 ( 
.A(n_1969),
.B(n_288),
.Y(n_2271)
);

NAND2xp5_ASAP7_75t_L g2272 ( 
.A(n_1972),
.B(n_288),
.Y(n_2272)
);

NAND2xp5_ASAP7_75t_L g2273 ( 
.A(n_1885),
.B(n_289),
.Y(n_2273)
);

BUFx3_ASAP7_75t_L g2274 ( 
.A(n_1864),
.Y(n_2274)
);

INVx2_ASAP7_75t_L g2275 ( 
.A(n_2018),
.Y(n_2275)
);

NOR2xp33_ASAP7_75t_L g2276 ( 
.A(n_1838),
.B(n_2063),
.Y(n_2276)
);

OAI22xp5_ASAP7_75t_L g2277 ( 
.A1(n_1958),
.A2(n_289),
.B1(n_290),
.B2(n_291),
.Y(n_2277)
);

AOI22xp33_ASAP7_75t_L g2278 ( 
.A1(n_1925),
.A2(n_290),
.B1(n_291),
.B2(n_292),
.Y(n_2278)
);

O2A1O1Ixp33_ASAP7_75t_L g2279 ( 
.A1(n_2064),
.A2(n_292),
.B(n_293),
.C(n_294),
.Y(n_2279)
);

AND2x4_ASAP7_75t_L g2280 ( 
.A(n_1864),
.B(n_293),
.Y(n_2280)
);

A2O1A1Ixp33_ASAP7_75t_L g2281 ( 
.A1(n_2031),
.A2(n_294),
.B(n_295),
.C(n_296),
.Y(n_2281)
);

OR2x6_ASAP7_75t_L g2282 ( 
.A(n_2013),
.B(n_297),
.Y(n_2282)
);

INVx2_ASAP7_75t_L g2283 ( 
.A(n_2032),
.Y(n_2283)
);

NAND2xp5_ASAP7_75t_L g2284 ( 
.A(n_1886),
.B(n_1888),
.Y(n_2284)
);

NAND2xp5_ASAP7_75t_L g2285 ( 
.A(n_1891),
.B(n_1958),
.Y(n_2285)
);

OAI22xp5_ASAP7_75t_SL g2286 ( 
.A1(n_1964),
.A2(n_298),
.B1(n_299),
.B2(n_300),
.Y(n_2286)
);

BUFx3_ASAP7_75t_L g2287 ( 
.A(n_1829),
.Y(n_2287)
);

INVx1_ASAP7_75t_L g2288 ( 
.A(n_1926),
.Y(n_2288)
);

HB1xp67_ASAP7_75t_L g2289 ( 
.A(n_2091),
.Y(n_2289)
);

INVx1_ASAP7_75t_SL g2290 ( 
.A(n_2098),
.Y(n_2290)
);

INVx1_ASAP7_75t_L g2291 ( 
.A(n_1927),
.Y(n_2291)
);

NAND2xp5_ASAP7_75t_SL g2292 ( 
.A(n_2068),
.B(n_301),
.Y(n_2292)
);

BUFx12f_ASAP7_75t_L g2293 ( 
.A(n_1973),
.Y(n_2293)
);

NOR3xp33_ASAP7_75t_SL g2294 ( 
.A(n_1916),
.B(n_1986),
.C(n_1948),
.Y(n_2294)
);

NAND2xp5_ASAP7_75t_L g2295 ( 
.A(n_1891),
.B(n_1959),
.Y(n_2295)
);

OR2x2_ASAP7_75t_L g2296 ( 
.A(n_1927),
.B(n_302),
.Y(n_2296)
);

NAND2xp5_ASAP7_75t_SL g2297 ( 
.A(n_2068),
.B(n_302),
.Y(n_2297)
);

A2O1A1Ixp33_ASAP7_75t_L g2298 ( 
.A1(n_2057),
.A2(n_303),
.B(n_304),
.C(n_305),
.Y(n_2298)
);

BUFx3_ASAP7_75t_L g2299 ( 
.A(n_1829),
.Y(n_2299)
);

INVx1_ASAP7_75t_SL g2300 ( 
.A(n_2098),
.Y(n_2300)
);

BUFx2_ASAP7_75t_L g2301 ( 
.A(n_1963),
.Y(n_2301)
);

NAND2xp5_ASAP7_75t_L g2302 ( 
.A(n_1959),
.B(n_304),
.Y(n_2302)
);

HB1xp67_ASAP7_75t_L g2303 ( 
.A(n_2097),
.Y(n_2303)
);

INVx2_ASAP7_75t_L g2304 ( 
.A(n_1950),
.Y(n_2304)
);

BUFx6f_ASAP7_75t_L g2305 ( 
.A(n_1837),
.Y(n_2305)
);

BUFx12f_ASAP7_75t_L g2306 ( 
.A(n_1973),
.Y(n_2306)
);

INVx1_ASAP7_75t_L g2307 ( 
.A(n_1934),
.Y(n_2307)
);

NAND2xp5_ASAP7_75t_L g2308 ( 
.A(n_1934),
.B(n_306),
.Y(n_2308)
);

NAND2x1p5_ASAP7_75t_L g2309 ( 
.A(n_2089),
.B(n_308),
.Y(n_2309)
);

O2A1O1Ixp5_ASAP7_75t_L g2310 ( 
.A1(n_1793),
.A2(n_308),
.B(n_309),
.C(n_310),
.Y(n_2310)
);

BUFx6f_ASAP7_75t_L g2311 ( 
.A(n_1837),
.Y(n_2311)
);

NOR2xp33_ASAP7_75t_L g2312 ( 
.A(n_2024),
.B(n_2028),
.Y(n_2312)
);

AOI22xp33_ASAP7_75t_L g2313 ( 
.A1(n_1965),
.A2(n_309),
.B1(n_312),
.B2(n_313),
.Y(n_2313)
);

INVx3_ASAP7_75t_SL g2314 ( 
.A(n_1824),
.Y(n_2314)
);

NOR2xp67_ASAP7_75t_SL g2315 ( 
.A(n_2082),
.B(n_312),
.Y(n_2315)
);

A2O1A1Ixp33_ASAP7_75t_L g2316 ( 
.A1(n_2021),
.A2(n_314),
.B(n_315),
.C(n_316),
.Y(n_2316)
);

AND2x4_ASAP7_75t_L g2317 ( 
.A(n_1877),
.B(n_315),
.Y(n_2317)
);

INVx2_ASAP7_75t_L g2318 ( 
.A(n_1935),
.Y(n_2318)
);

A2O1A1Ixp33_ASAP7_75t_L g2319 ( 
.A1(n_2056),
.A2(n_317),
.B(n_319),
.C(n_320),
.Y(n_2319)
);

AND2x4_ASAP7_75t_L g2320 ( 
.A(n_1877),
.B(n_321),
.Y(n_2320)
);

NAND2xp5_ASAP7_75t_L g2321 ( 
.A(n_1989),
.B(n_324),
.Y(n_2321)
);

INVx3_ASAP7_75t_SL g2322 ( 
.A(n_1875),
.Y(n_2322)
);

AOI21xp5_ASAP7_75t_L g2323 ( 
.A1(n_1807),
.A2(n_326),
.B(n_327),
.Y(n_2323)
);

OAI21xp33_ASAP7_75t_SL g2324 ( 
.A1(n_2027),
.A2(n_328),
.B(n_330),
.Y(n_2324)
);

A2O1A1Ixp33_ASAP7_75t_L g2325 ( 
.A1(n_2050),
.A2(n_328),
.B(n_330),
.C(n_331),
.Y(n_2325)
);

BUFx6f_ASAP7_75t_L g2326 ( 
.A(n_1869),
.Y(n_2326)
);

NAND2xp5_ASAP7_75t_SL g2327 ( 
.A(n_2089),
.B(n_333),
.Y(n_2327)
);

INVx4_ASAP7_75t_L g2328 ( 
.A(n_1829),
.Y(n_2328)
);

NOR3xp33_ASAP7_75t_SL g2329 ( 
.A(n_1942),
.B(n_333),
.C(n_334),
.Y(n_2329)
);

INVx1_ASAP7_75t_L g2330 ( 
.A(n_1940),
.Y(n_2330)
);

AOI222xp33_ASAP7_75t_L g2331 ( 
.A1(n_1967),
.A2(n_335),
.B1(n_336),
.B2(n_337),
.C1(n_338),
.C2(n_339),
.Y(n_2331)
);

BUFx6f_ASAP7_75t_L g2332 ( 
.A(n_1869),
.Y(n_2332)
);

CKINVDCx14_ASAP7_75t_R g2333 ( 
.A(n_2075),
.Y(n_2333)
);

BUFx3_ASAP7_75t_L g2334 ( 
.A(n_1829),
.Y(n_2334)
);

CKINVDCx5p33_ASAP7_75t_R g2335 ( 
.A(n_2099),
.Y(n_2335)
);

OAI22xp5_ASAP7_75t_L g2336 ( 
.A1(n_1955),
.A2(n_337),
.B1(n_338),
.B2(n_339),
.Y(n_2336)
);

OAI21xp33_ASAP7_75t_L g2337 ( 
.A1(n_1942),
.A2(n_341),
.B(n_342),
.Y(n_2337)
);

NOR2xp33_ASAP7_75t_L g2338 ( 
.A(n_1978),
.B(n_1966),
.Y(n_2338)
);

NOR2xp33_ASAP7_75t_L g2339 ( 
.A(n_1990),
.B(n_344),
.Y(n_2339)
);

OAI22x1_ASAP7_75t_L g2340 ( 
.A1(n_2100),
.A2(n_345),
.B1(n_346),
.B2(n_347),
.Y(n_2340)
);

AOI22xp5_ASAP7_75t_L g2341 ( 
.A1(n_1967),
.A2(n_348),
.B1(n_349),
.B2(n_350),
.Y(n_2341)
);

INVx1_ASAP7_75t_L g2342 ( 
.A(n_1940),
.Y(n_2342)
);

O2A1O1Ixp33_ASAP7_75t_L g2343 ( 
.A1(n_1994),
.A2(n_349),
.B(n_351),
.C(n_352),
.Y(n_2343)
);

O2A1O1Ixp33_ASAP7_75t_L g2344 ( 
.A1(n_1995),
.A2(n_351),
.B(n_353),
.C(n_354),
.Y(n_2344)
);

OAI22xp5_ASAP7_75t_L g2345 ( 
.A1(n_2012),
.A2(n_353),
.B1(n_354),
.B2(n_355),
.Y(n_2345)
);

AOI21xp5_ASAP7_75t_L g2346 ( 
.A1(n_1793),
.A2(n_356),
.B(n_357),
.Y(n_2346)
);

NAND2x1_ASAP7_75t_L g2347 ( 
.A(n_2328),
.B(n_1973),
.Y(n_2347)
);

NAND2xp5_ASAP7_75t_L g2348 ( 
.A(n_2111),
.B(n_1997),
.Y(n_2348)
);

INVx2_ASAP7_75t_L g2349 ( 
.A(n_2152),
.Y(n_2349)
);

OAI221xp5_ASAP7_75t_L g2350 ( 
.A1(n_2229),
.A2(n_2006),
.B1(n_1976),
.B2(n_1983),
.C(n_1982),
.Y(n_2350)
);

AND2x2_ASAP7_75t_L g2351 ( 
.A(n_2101),
.B(n_2058),
.Y(n_2351)
);

NOR2xp33_ASAP7_75t_L g2352 ( 
.A(n_2333),
.B(n_2071),
.Y(n_2352)
);

AOI21xp5_ASAP7_75t_L g2353 ( 
.A1(n_2138),
.A2(n_2144),
.B(n_2260),
.Y(n_2353)
);

AOI21xp5_ASAP7_75t_L g2354 ( 
.A1(n_2285),
.A2(n_1894),
.B(n_1893),
.Y(n_2354)
);

AND2x2_ASAP7_75t_L g2355 ( 
.A(n_2147),
.B(n_2001),
.Y(n_2355)
);

INVx1_ASAP7_75t_L g2356 ( 
.A(n_2154),
.Y(n_2356)
);

OAI22xp5_ASAP7_75t_L g2357 ( 
.A1(n_2282),
.A2(n_2167),
.B1(n_2335),
.B2(n_2186),
.Y(n_2357)
);

NAND2xp5_ASAP7_75t_L g2358 ( 
.A(n_2120),
.B(n_1904),
.Y(n_2358)
);

BUFx6f_ASAP7_75t_L g2359 ( 
.A(n_2159),
.Y(n_2359)
);

INVx1_ASAP7_75t_L g2360 ( 
.A(n_2163),
.Y(n_2360)
);

O2A1O1Ixp33_ASAP7_75t_SL g2361 ( 
.A1(n_2118),
.A2(n_2085),
.B(n_2087),
.C(n_1947),
.Y(n_2361)
);

HB1xp67_ASAP7_75t_L g2362 ( 
.A(n_2210),
.Y(n_2362)
);

AOI21xp5_ASAP7_75t_L g2363 ( 
.A1(n_2295),
.A2(n_1894),
.B(n_1895),
.Y(n_2363)
);

INVx2_ASAP7_75t_SL g2364 ( 
.A(n_2128),
.Y(n_2364)
);

INVx1_ASAP7_75t_L g2365 ( 
.A(n_2251),
.Y(n_2365)
);

AO31x2_ASAP7_75t_L g2366 ( 
.A1(n_2140),
.A2(n_2009),
.A3(n_2146),
.B(n_2301),
.Y(n_2366)
);

A2O1A1Ixp33_ASAP7_75t_L g2367 ( 
.A1(n_2247),
.A2(n_2324),
.B(n_2312),
.C(n_2201),
.Y(n_2367)
);

NAND2xp5_ASAP7_75t_L g2368 ( 
.A(n_2219),
.B(n_1904),
.Y(n_2368)
);

NAND2xp5_ASAP7_75t_L g2369 ( 
.A(n_2180),
.B(n_1948),
.Y(n_2369)
);

INVxp67_ASAP7_75t_L g2370 ( 
.A(n_2222),
.Y(n_2370)
);

INVxp67_ASAP7_75t_SL g2371 ( 
.A(n_2133),
.Y(n_2371)
);

AOI21xp5_ASAP7_75t_L g2372 ( 
.A1(n_2110),
.A2(n_1910),
.B(n_1901),
.Y(n_2372)
);

INVx3_ASAP7_75t_L g2373 ( 
.A(n_2160),
.Y(n_2373)
);

AO31x2_ASAP7_75t_L g2374 ( 
.A1(n_2178),
.A2(n_2015),
.A3(n_1896),
.B(n_1845),
.Y(n_2374)
);

INVx1_ASAP7_75t_L g2375 ( 
.A(n_2164),
.Y(n_2375)
);

AND2x4_ASAP7_75t_L g2376 ( 
.A(n_2187),
.B(n_2040),
.Y(n_2376)
);

A2O1A1Ixp33_ASAP7_75t_L g2377 ( 
.A1(n_2247),
.A2(n_2030),
.B(n_2023),
.C(n_2037),
.Y(n_2377)
);

A2O1A1Ixp33_ASAP7_75t_L g2378 ( 
.A1(n_2324),
.A2(n_2093),
.B(n_2096),
.C(n_2094),
.Y(n_2378)
);

INVx1_ASAP7_75t_L g2379 ( 
.A(n_2104),
.Y(n_2379)
);

AOI21xp5_ASAP7_75t_L g2380 ( 
.A1(n_2107),
.A2(n_1911),
.B(n_1908),
.Y(n_2380)
);

INVx2_ASAP7_75t_L g2381 ( 
.A(n_2116),
.Y(n_2381)
);

AO21x1_ASAP7_75t_L g2382 ( 
.A1(n_2155),
.A2(n_2077),
.B(n_2048),
.Y(n_2382)
);

INVxp67_ASAP7_75t_SL g2383 ( 
.A(n_2289),
.Y(n_2383)
);

NAND2xp33_ASAP7_75t_L g2384 ( 
.A(n_2187),
.B(n_1973),
.Y(n_2384)
);

AO21x2_ASAP7_75t_L g2385 ( 
.A1(n_2245),
.A2(n_1882),
.B(n_1892),
.Y(n_2385)
);

INVx1_ASAP7_75t_L g2386 ( 
.A(n_2130),
.Y(n_2386)
);

NOR2xp33_ASAP7_75t_L g2387 ( 
.A(n_2244),
.B(n_2014),
.Y(n_2387)
);

NOR2x1_ASAP7_75t_SL g2388 ( 
.A(n_2293),
.B(n_2097),
.Y(n_2388)
);

INVx6_ASAP7_75t_L g2389 ( 
.A(n_2117),
.Y(n_2389)
);

INVx2_ASAP7_75t_L g2390 ( 
.A(n_2137),
.Y(n_2390)
);

A2O1A1Ixp33_ASAP7_75t_L g2391 ( 
.A1(n_2145),
.A2(n_2069),
.B(n_2020),
.C(n_2070),
.Y(n_2391)
);

OR2x6_ASAP7_75t_L g2392 ( 
.A(n_2160),
.B(n_2038),
.Y(n_2392)
);

NAND2xp5_ASAP7_75t_L g2393 ( 
.A(n_2136),
.B(n_2062),
.Y(n_2393)
);

INVx1_ASAP7_75t_L g2394 ( 
.A(n_2185),
.Y(n_2394)
);

INVx1_ASAP7_75t_L g2395 ( 
.A(n_2230),
.Y(n_2395)
);

INVx1_ASAP7_75t_L g2396 ( 
.A(n_2240),
.Y(n_2396)
);

AOI21xp5_ASAP7_75t_L g2397 ( 
.A1(n_2123),
.A2(n_1938),
.B(n_1933),
.Y(n_2397)
);

BUFx2_ASAP7_75t_L g2398 ( 
.A(n_2105),
.Y(n_2398)
);

BUFx2_ASAP7_75t_L g2399 ( 
.A(n_2205),
.Y(n_2399)
);

CKINVDCx5p33_ASAP7_75t_R g2400 ( 
.A(n_2139),
.Y(n_2400)
);

AND2x4_ASAP7_75t_L g2401 ( 
.A(n_2187),
.B(n_2040),
.Y(n_2401)
);

INVx3_ASAP7_75t_SL g2402 ( 
.A(n_2129),
.Y(n_2402)
);

CKINVDCx5p33_ASAP7_75t_R g2403 ( 
.A(n_2165),
.Y(n_2403)
);

AOI21xp5_ASAP7_75t_L g2404 ( 
.A1(n_2106),
.A2(n_1992),
.B(n_1909),
.Y(n_2404)
);

AOI22xp33_ASAP7_75t_SL g2405 ( 
.A1(n_2250),
.A2(n_1973),
.B1(n_2092),
.B2(n_2095),
.Y(n_2405)
);

A2O1A1Ixp33_ASAP7_75t_L g2406 ( 
.A1(n_2142),
.A2(n_2039),
.B(n_2060),
.C(n_1944),
.Y(n_2406)
);

AND2x4_ASAP7_75t_L g2407 ( 
.A(n_2112),
.B(n_2065),
.Y(n_2407)
);

NAND2xp5_ASAP7_75t_SL g2408 ( 
.A(n_2226),
.B(n_1932),
.Y(n_2408)
);

AOI21xp5_ASAP7_75t_L g2409 ( 
.A1(n_2183),
.A2(n_2000),
.B(n_2004),
.Y(n_2409)
);

BUFx6f_ASAP7_75t_L g2410 ( 
.A(n_2135),
.Y(n_2410)
);

CKINVDCx5p33_ASAP7_75t_R g2411 ( 
.A(n_2188),
.Y(n_2411)
);

AOI21xp5_ASAP7_75t_L g2412 ( 
.A1(n_2284),
.A2(n_1880),
.B(n_1840),
.Y(n_2412)
);

O2A1O1Ixp33_ASAP7_75t_SL g2413 ( 
.A1(n_2127),
.A2(n_1929),
.B(n_2017),
.C(n_1876),
.Y(n_2413)
);

OAI21xp5_ASAP7_75t_L g2414 ( 
.A1(n_2166),
.A2(n_2211),
.B(n_2339),
.Y(n_2414)
);

AOI22xp5_ASAP7_75t_L g2415 ( 
.A1(n_2108),
.A2(n_1849),
.B1(n_2045),
.B2(n_2042),
.Y(n_2415)
);

OAI21xp5_ASAP7_75t_L g2416 ( 
.A1(n_2294),
.A2(n_1817),
.B(n_2086),
.Y(n_2416)
);

BUFx2_ASAP7_75t_L g2417 ( 
.A(n_2205),
.Y(n_2417)
);

AND2x2_ASAP7_75t_L g2418 ( 
.A(n_2162),
.B(n_358),
.Y(n_2418)
);

CKINVDCx16_ASAP7_75t_R g2419 ( 
.A(n_2196),
.Y(n_2419)
);

AO21x2_ASAP7_75t_L g2420 ( 
.A1(n_2245),
.A2(n_2115),
.B(n_2181),
.Y(n_2420)
);

BUFx2_ASAP7_75t_R g2421 ( 
.A(n_2204),
.Y(n_2421)
);

BUFx2_ASAP7_75t_L g2422 ( 
.A(n_2112),
.Y(n_2422)
);

AOI21xp5_ASAP7_75t_L g2423 ( 
.A1(n_2304),
.A2(n_1912),
.B(n_1905),
.Y(n_2423)
);

BUFx10_ASAP7_75t_L g2424 ( 
.A(n_2134),
.Y(n_2424)
);

NOR2xp33_ASAP7_75t_SL g2425 ( 
.A(n_2200),
.B(n_1829),
.Y(n_2425)
);

INVx1_ASAP7_75t_L g2426 ( 
.A(n_2256),
.Y(n_2426)
);

INVxp67_ASAP7_75t_SL g2427 ( 
.A(n_2306),
.Y(n_2427)
);

INVx1_ASAP7_75t_L g2428 ( 
.A(n_2275),
.Y(n_2428)
);

INVxp67_ASAP7_75t_SL g2429 ( 
.A(n_2303),
.Y(n_2429)
);

O2A1O1Ixp33_ASAP7_75t_SL g2430 ( 
.A1(n_2281),
.A2(n_1871),
.B(n_1865),
.C(n_2061),
.Y(n_2430)
);

A2O1A1Ixp33_ASAP7_75t_L g2431 ( 
.A1(n_2337),
.A2(n_2238),
.B(n_2209),
.C(n_2262),
.Y(n_2431)
);

INVx1_ASAP7_75t_L g2432 ( 
.A(n_2283),
.Y(n_2432)
);

NAND2xp5_ASAP7_75t_L g2433 ( 
.A(n_2171),
.B(n_2045),
.Y(n_2433)
);

INVx1_ASAP7_75t_L g2434 ( 
.A(n_2237),
.Y(n_2434)
);

OAI21xp5_ASAP7_75t_L g2435 ( 
.A1(n_2191),
.A2(n_2310),
.B(n_2316),
.Y(n_2435)
);

AOI21xp5_ASAP7_75t_L g2436 ( 
.A1(n_2318),
.A2(n_1951),
.B(n_1937),
.Y(n_2436)
);

OAI21x1_ASAP7_75t_L g2437 ( 
.A1(n_2125),
.A2(n_1971),
.B(n_1979),
.Y(n_2437)
);

OAI21xp5_ASAP7_75t_L g2438 ( 
.A1(n_2243),
.A2(n_1957),
.B(n_1949),
.Y(n_2438)
);

OR2x2_ASAP7_75t_L g2439 ( 
.A(n_2282),
.B(n_2051),
.Y(n_2439)
);

BUFx3_ASAP7_75t_L g2440 ( 
.A(n_2224),
.Y(n_2440)
);

A2O1A1Ixp33_ASAP7_75t_L g2441 ( 
.A1(n_2315),
.A2(n_1991),
.B(n_1984),
.C(n_1988),
.Y(n_2441)
);

NOR2xp33_ASAP7_75t_L g2442 ( 
.A(n_2122),
.B(n_2084),
.Y(n_2442)
);

AOI21xp5_ASAP7_75t_L g2443 ( 
.A1(n_2218),
.A2(n_1998),
.B(n_1872),
.Y(n_2443)
);

AND2x2_ASAP7_75t_L g2444 ( 
.A(n_2194),
.B(n_360),
.Y(n_2444)
);

NAND2xp5_ASAP7_75t_L g2445 ( 
.A(n_2232),
.B(n_2051),
.Y(n_2445)
);

BUFx6f_ASAP7_75t_L g2446 ( 
.A(n_2135),
.Y(n_2446)
);

BUFx12f_ASAP7_75t_L g2447 ( 
.A(n_2153),
.Y(n_2447)
);

AOI21xp5_ASAP7_75t_L g2448 ( 
.A1(n_2239),
.A2(n_1846),
.B(n_2078),
.Y(n_2448)
);

OAI22xp5_ASAP7_75t_L g2449 ( 
.A1(n_2196),
.A2(n_2065),
.B1(n_2059),
.B2(n_1855),
.Y(n_2449)
);

NAND2xp5_ASAP7_75t_L g2450 ( 
.A(n_2252),
.B(n_2254),
.Y(n_2450)
);

A2O1A1Ixp33_ASAP7_75t_L g2451 ( 
.A1(n_2263),
.A2(n_1853),
.B(n_363),
.C(n_364),
.Y(n_2451)
);

AOI221xp5_ASAP7_75t_L g2452 ( 
.A1(n_2336),
.A2(n_361),
.B1(n_363),
.B2(n_365),
.C(n_367),
.Y(n_2452)
);

O2A1O1Ixp33_ASAP7_75t_SL g2453 ( 
.A1(n_2113),
.A2(n_361),
.B(n_365),
.C(n_368),
.Y(n_2453)
);

INVx3_ASAP7_75t_L g2454 ( 
.A(n_2143),
.Y(n_2454)
);

NAND2xp5_ASAP7_75t_L g2455 ( 
.A(n_2259),
.B(n_376),
.Y(n_2455)
);

NOR2xp33_ASAP7_75t_L g2456 ( 
.A(n_2103),
.B(n_370),
.Y(n_2456)
);

AO32x2_ASAP7_75t_L g2457 ( 
.A1(n_2286),
.A2(n_371),
.A3(n_372),
.B1(n_373),
.B2(n_374),
.Y(n_2457)
);

AOI21xp5_ASAP7_75t_L g2458 ( 
.A1(n_2288),
.A2(n_371),
.B(n_372),
.Y(n_2458)
);

AOI21xp5_ASAP7_75t_L g2459 ( 
.A1(n_2291),
.A2(n_374),
.B(n_375),
.Y(n_2459)
);

AOI21xp5_ASAP7_75t_L g2460 ( 
.A1(n_2307),
.A2(n_2342),
.B(n_2330),
.Y(n_2460)
);

OAI21xp5_ASAP7_75t_L g2461 ( 
.A1(n_2149),
.A2(n_2272),
.B(n_2216),
.Y(n_2461)
);

AOI21xp5_ASAP7_75t_L g2462 ( 
.A1(n_2212),
.A2(n_2173),
.B(n_2176),
.Y(n_2462)
);

OAI22x1_ASAP7_75t_L g2463 ( 
.A1(n_2341),
.A2(n_2158),
.B1(n_2231),
.B2(n_2226),
.Y(n_2463)
);

AOI21xp5_ASAP7_75t_L g2464 ( 
.A1(n_2126),
.A2(n_2302),
.B(n_2156),
.Y(n_2464)
);

OR2x2_ASAP7_75t_L g2465 ( 
.A(n_2169),
.B(n_2179),
.Y(n_2465)
);

AOI21xp5_ASAP7_75t_L g2466 ( 
.A1(n_2151),
.A2(n_2157),
.B(n_2276),
.Y(n_2466)
);

INVx2_ASAP7_75t_L g2467 ( 
.A(n_2102),
.Y(n_2467)
);

INVx1_ASAP7_75t_L g2468 ( 
.A(n_2280),
.Y(n_2468)
);

AO31x2_ASAP7_75t_L g2469 ( 
.A1(n_2172),
.A2(n_2340),
.A3(n_2220),
.B(n_2346),
.Y(n_2469)
);

AOI21xp5_ASAP7_75t_L g2470 ( 
.A1(n_2290),
.A2(n_2300),
.B(n_2206),
.Y(n_2470)
);

AOI21x1_ASAP7_75t_L g2471 ( 
.A1(n_2199),
.A2(n_2266),
.B(n_2161),
.Y(n_2471)
);

CKINVDCx20_ASAP7_75t_R g2472 ( 
.A(n_2148),
.Y(n_2472)
);

CKINVDCx11_ASAP7_75t_R g2473 ( 
.A(n_2196),
.Y(n_2473)
);

BUFx10_ASAP7_75t_L g2474 ( 
.A(n_2141),
.Y(n_2474)
);

O2A1O1Ixp33_ASAP7_75t_SL g2475 ( 
.A1(n_2223),
.A2(n_2325),
.B(n_2298),
.C(n_2319),
.Y(n_2475)
);

INVx2_ASAP7_75t_L g2476 ( 
.A(n_2270),
.Y(n_2476)
);

INVx2_ASAP7_75t_L g2477 ( 
.A(n_2296),
.Y(n_2477)
);

AOI21xp5_ASAP7_75t_L g2478 ( 
.A1(n_2308),
.A2(n_2321),
.B(n_2273),
.Y(n_2478)
);

INVx2_ASAP7_75t_L g2479 ( 
.A(n_2317),
.Y(n_2479)
);

AOI21xp5_ASAP7_75t_L g2480 ( 
.A1(n_2253),
.A2(n_2114),
.B(n_2242),
.Y(n_2480)
);

OR2x2_ASAP7_75t_L g2481 ( 
.A(n_2207),
.B(n_2280),
.Y(n_2481)
);

AOI21xp5_ASAP7_75t_L g2482 ( 
.A1(n_2135),
.A2(n_2305),
.B(n_2242),
.Y(n_2482)
);

OAI21xp5_ASAP7_75t_SL g2483 ( 
.A1(n_2331),
.A2(n_2341),
.B(n_2231),
.Y(n_2483)
);

INVx2_ASAP7_75t_L g2484 ( 
.A(n_2317),
.Y(n_2484)
);

OAI21xp5_ASAP7_75t_L g2485 ( 
.A1(n_2271),
.A2(n_2225),
.B(n_2236),
.Y(n_2485)
);

OAI21xp5_ASAP7_75t_L g2486 ( 
.A1(n_2198),
.A2(n_2184),
.B(n_2190),
.Y(n_2486)
);

HB1xp67_ASAP7_75t_L g2487 ( 
.A(n_2320),
.Y(n_2487)
);

AOI21x1_ASAP7_75t_L g2488 ( 
.A1(n_2267),
.A2(n_2143),
.B(n_2327),
.Y(n_2488)
);

BUFx2_ASAP7_75t_R g2489 ( 
.A(n_2322),
.Y(n_2489)
);

NOR2xp33_ASAP7_75t_SL g2490 ( 
.A(n_2328),
.B(n_2258),
.Y(n_2490)
);

AOI21xp5_ASAP7_75t_L g2491 ( 
.A1(n_2170),
.A2(n_2242),
.B(n_2208),
.Y(n_2491)
);

NOR2xp33_ASAP7_75t_L g2492 ( 
.A(n_2132),
.B(n_2314),
.Y(n_2492)
);

NAND2xp5_ASAP7_75t_L g2493 ( 
.A(n_2338),
.B(n_2174),
.Y(n_2493)
);

AOI21xp5_ASAP7_75t_L g2494 ( 
.A1(n_2170),
.A2(n_2213),
.B(n_2208),
.Y(n_2494)
);

O2A1O1Ixp5_ASAP7_75t_SL g2495 ( 
.A1(n_2268),
.A2(n_2292),
.B(n_2297),
.C(n_2150),
.Y(n_2495)
);

AND2x2_ASAP7_75t_L g2496 ( 
.A(n_2329),
.B(n_2257),
.Y(n_2496)
);

AOI22xp33_ASAP7_75t_L g2497 ( 
.A1(n_2463),
.A2(n_2177),
.B1(n_2189),
.B2(n_2286),
.Y(n_2497)
);

BUFx10_ASAP7_75t_L g2498 ( 
.A(n_2364),
.Y(n_2498)
);

INVx3_ASAP7_75t_L g2499 ( 
.A(n_2373),
.Y(n_2499)
);

AOI22xp5_ASAP7_75t_L g2500 ( 
.A1(n_2483),
.A2(n_2177),
.B1(n_2189),
.B2(n_2158),
.Y(n_2500)
);

CKINVDCx11_ASAP7_75t_R g2501 ( 
.A(n_2447),
.Y(n_2501)
);

INVx4_ASAP7_75t_L g2502 ( 
.A(n_2373),
.Y(n_2502)
);

AOI22xp33_ASAP7_75t_SL g2503 ( 
.A1(n_2357),
.A2(n_2235),
.B1(n_2320),
.B2(n_2309),
.Y(n_2503)
);

BUFx3_ASAP7_75t_L g2504 ( 
.A(n_2359),
.Y(n_2504)
);

INVx1_ASAP7_75t_L g2505 ( 
.A(n_2356),
.Y(n_2505)
);

BUFx12f_ASAP7_75t_L g2506 ( 
.A(n_2389),
.Y(n_2506)
);

INVx1_ASAP7_75t_L g2507 ( 
.A(n_2360),
.Y(n_2507)
);

INVx6_ASAP7_75t_L g2508 ( 
.A(n_2474),
.Y(n_2508)
);

CKINVDCx11_ASAP7_75t_R g2509 ( 
.A(n_2402),
.Y(n_2509)
);

OAI22xp5_ASAP7_75t_L g2510 ( 
.A1(n_2419),
.A2(n_2264),
.B1(n_2234),
.B2(n_2255),
.Y(n_2510)
);

INVx1_ASAP7_75t_SL g2511 ( 
.A(n_2399),
.Y(n_2511)
);

AOI22xp33_ASAP7_75t_L g2512 ( 
.A1(n_2473),
.A2(n_2496),
.B1(n_2456),
.B2(n_2461),
.Y(n_2512)
);

AOI22xp33_ASAP7_75t_L g2513 ( 
.A1(n_2493),
.A2(n_2235),
.B1(n_2193),
.B2(n_2182),
.Y(n_2513)
);

OR2x2_ASAP7_75t_L g2514 ( 
.A(n_2365),
.B(n_2175),
.Y(n_2514)
);

OAI22xp5_ASAP7_75t_L g2515 ( 
.A1(n_2367),
.A2(n_2313),
.B1(n_2203),
.B2(n_2277),
.Y(n_2515)
);

BUFx6f_ASAP7_75t_L g2516 ( 
.A(n_2359),
.Y(n_2516)
);

INVx2_ASAP7_75t_SL g2517 ( 
.A(n_2474),
.Y(n_2517)
);

OAI22xp33_ASAP7_75t_L g2518 ( 
.A1(n_2425),
.A2(n_2109),
.B1(n_2233),
.B2(n_2227),
.Y(n_2518)
);

INVx4_ASAP7_75t_L g2519 ( 
.A(n_2359),
.Y(n_2519)
);

INVx5_ASAP7_75t_L g2520 ( 
.A(n_2389),
.Y(n_2520)
);

INVx1_ASAP7_75t_L g2521 ( 
.A(n_2379),
.Y(n_2521)
);

AOI22xp33_ASAP7_75t_SL g2522 ( 
.A1(n_2487),
.A2(n_2175),
.B1(n_2334),
.B2(n_2299),
.Y(n_2522)
);

OAI22xp5_ASAP7_75t_L g2523 ( 
.A1(n_2405),
.A2(n_2278),
.B1(n_2109),
.B2(n_2265),
.Y(n_2523)
);

BUFx2_ASAP7_75t_L g2524 ( 
.A(n_2362),
.Y(n_2524)
);

OAI22xp5_ASAP7_75t_L g2525 ( 
.A1(n_2439),
.A2(n_2109),
.B1(n_2249),
.B2(n_2246),
.Y(n_2525)
);

INVx11_ASAP7_75t_L g2526 ( 
.A(n_2472),
.Y(n_2526)
);

INVx6_ASAP7_75t_L g2527 ( 
.A(n_2424),
.Y(n_2527)
);

INVx1_ASAP7_75t_L g2528 ( 
.A(n_2386),
.Y(n_2528)
);

BUFx2_ASAP7_75t_SL g2529 ( 
.A(n_2424),
.Y(n_2529)
);

INVx1_ASAP7_75t_L g2530 ( 
.A(n_2375),
.Y(n_2530)
);

BUFx6f_ASAP7_75t_L g2531 ( 
.A(n_2410),
.Y(n_2531)
);

AOI22xp33_ASAP7_75t_SL g2532 ( 
.A1(n_2388),
.A2(n_2287),
.B1(n_2345),
.B2(n_2119),
.Y(n_2532)
);

INVx1_ASAP7_75t_L g2533 ( 
.A(n_2381),
.Y(n_2533)
);

INVx1_ASAP7_75t_L g2534 ( 
.A(n_2390),
.Y(n_2534)
);

HB1xp67_ASAP7_75t_L g2535 ( 
.A(n_2429),
.Y(n_2535)
);

CKINVDCx11_ASAP7_75t_R g2536 ( 
.A(n_2440),
.Y(n_2536)
);

INVx4_ASAP7_75t_L g2537 ( 
.A(n_2417),
.Y(n_2537)
);

INVx1_ASAP7_75t_L g2538 ( 
.A(n_2394),
.Y(n_2538)
);

AOI22xp33_ASAP7_75t_L g2539 ( 
.A1(n_2348),
.A2(n_2197),
.B1(n_2124),
.B2(n_2323),
.Y(n_2539)
);

AOI22xp33_ASAP7_75t_L g2540 ( 
.A1(n_2352),
.A2(n_2192),
.B1(n_2195),
.B2(n_2217),
.Y(n_2540)
);

INVx2_ASAP7_75t_L g2541 ( 
.A(n_2349),
.Y(n_2541)
);

CKINVDCx11_ASAP7_75t_R g2542 ( 
.A(n_2398),
.Y(n_2542)
);

AOI22xp33_ASAP7_75t_L g2543 ( 
.A1(n_2414),
.A2(n_2131),
.B1(n_2221),
.B2(n_2228),
.Y(n_2543)
);

OAI22xp5_ASAP7_75t_SL g2544 ( 
.A1(n_2411),
.A2(n_2261),
.B1(n_2228),
.B2(n_2168),
.Y(n_2544)
);

OAI22xp5_ASAP7_75t_L g2545 ( 
.A1(n_2369),
.A2(n_2248),
.B1(n_2241),
.B2(n_2215),
.Y(n_2545)
);

BUFx3_ASAP7_75t_L g2546 ( 
.A(n_2400),
.Y(n_2546)
);

AOI22xp33_ASAP7_75t_SL g2547 ( 
.A1(n_2388),
.A2(n_2119),
.B1(n_2261),
.B2(n_2274),
.Y(n_2547)
);

INVx3_ASAP7_75t_L g2548 ( 
.A(n_2347),
.Y(n_2548)
);

INVxp67_ASAP7_75t_SL g2549 ( 
.A(n_2384),
.Y(n_2549)
);

OAI22xp5_ASAP7_75t_L g2550 ( 
.A1(n_2431),
.A2(n_2202),
.B1(n_2344),
.B2(n_2343),
.Y(n_2550)
);

AOI22xp33_ASAP7_75t_L g2551 ( 
.A1(n_2355),
.A2(n_2121),
.B1(n_2170),
.B2(n_2208),
.Y(n_2551)
);

BUFx6f_ASAP7_75t_L g2552 ( 
.A(n_2410),
.Y(n_2552)
);

AOI22xp33_ASAP7_75t_SL g2553 ( 
.A1(n_2449),
.A2(n_2213),
.B1(n_2214),
.B2(n_2269),
.Y(n_2553)
);

INVx1_ASAP7_75t_L g2554 ( 
.A(n_2395),
.Y(n_2554)
);

NAND2x1p5_ASAP7_75t_L g2555 ( 
.A(n_2376),
.B(n_2213),
.Y(n_2555)
);

CKINVDCx11_ASAP7_75t_R g2556 ( 
.A(n_2403),
.Y(n_2556)
);

HB1xp67_ASAP7_75t_L g2557 ( 
.A(n_2383),
.Y(n_2557)
);

INVx2_ASAP7_75t_L g2558 ( 
.A(n_2396),
.Y(n_2558)
);

OAI22xp5_ASAP7_75t_L g2559 ( 
.A1(n_2415),
.A2(n_2279),
.B1(n_2332),
.B2(n_2214),
.Y(n_2559)
);

INVx2_ASAP7_75t_L g2560 ( 
.A(n_2426),
.Y(n_2560)
);

BUFx4_ASAP7_75t_SL g2561 ( 
.A(n_2489),
.Y(n_2561)
);

INVx6_ASAP7_75t_L g2562 ( 
.A(n_2376),
.Y(n_2562)
);

INVx1_ASAP7_75t_L g2563 ( 
.A(n_2428),
.Y(n_2563)
);

CKINVDCx11_ASAP7_75t_R g2564 ( 
.A(n_2421),
.Y(n_2564)
);

OR2x2_ASAP7_75t_L g2565 ( 
.A(n_2370),
.B(n_2214),
.Y(n_2565)
);

CKINVDCx11_ASAP7_75t_R g2566 ( 
.A(n_2422),
.Y(n_2566)
);

OAI22xp5_ASAP7_75t_L g2567 ( 
.A1(n_2481),
.A2(n_2451),
.B1(n_2484),
.B2(n_2479),
.Y(n_2567)
);

HB1xp67_ASAP7_75t_L g2568 ( 
.A(n_2432),
.Y(n_2568)
);

BUFx4f_ASAP7_75t_SL g2569 ( 
.A(n_2454),
.Y(n_2569)
);

INVx2_ASAP7_75t_L g2570 ( 
.A(n_2467),
.Y(n_2570)
);

BUFx6f_ASAP7_75t_L g2571 ( 
.A(n_2410),
.Y(n_2571)
);

AOI22xp33_ASAP7_75t_L g2572 ( 
.A1(n_2476),
.A2(n_2269),
.B1(n_2305),
.B2(n_2311),
.Y(n_2572)
);

INVx1_ASAP7_75t_L g2573 ( 
.A(n_2450),
.Y(n_2573)
);

INVx2_ASAP7_75t_L g2574 ( 
.A(n_2445),
.Y(n_2574)
);

INVx5_ASAP7_75t_L g2575 ( 
.A(n_2446),
.Y(n_2575)
);

BUFx12f_ASAP7_75t_L g2576 ( 
.A(n_2444),
.Y(n_2576)
);

INVx1_ASAP7_75t_L g2577 ( 
.A(n_2477),
.Y(n_2577)
);

BUFx2_ASAP7_75t_SL g2578 ( 
.A(n_2427),
.Y(n_2578)
);

OAI22xp5_ASAP7_75t_L g2579 ( 
.A1(n_2393),
.A2(n_2269),
.B1(n_2311),
.B2(n_2326),
.Y(n_2579)
);

INVx1_ASAP7_75t_L g2580 ( 
.A(n_2434),
.Y(n_2580)
);

INVx8_ASAP7_75t_L g2581 ( 
.A(n_2401),
.Y(n_2581)
);

INVx1_ASAP7_75t_L g2582 ( 
.A(n_2351),
.Y(n_2582)
);

CKINVDCx5p33_ASAP7_75t_R g2583 ( 
.A(n_2442),
.Y(n_2583)
);

INVx1_ASAP7_75t_L g2584 ( 
.A(n_2455),
.Y(n_2584)
);

BUFx12f_ASAP7_75t_L g2585 ( 
.A(n_2407),
.Y(n_2585)
);

CKINVDCx11_ASAP7_75t_R g2586 ( 
.A(n_2392),
.Y(n_2586)
);

OAI22xp5_ASAP7_75t_L g2587 ( 
.A1(n_2368),
.A2(n_2408),
.B1(n_2433),
.B2(n_2465),
.Y(n_2587)
);

BUFx3_ASAP7_75t_L g2588 ( 
.A(n_2401),
.Y(n_2588)
);

INVx2_ASAP7_75t_L g2589 ( 
.A(n_2446),
.Y(n_2589)
);

INVx1_ASAP7_75t_L g2590 ( 
.A(n_2468),
.Y(n_2590)
);

BUFx6f_ASAP7_75t_SL g2591 ( 
.A(n_2407),
.Y(n_2591)
);

OAI22xp33_ASAP7_75t_L g2592 ( 
.A1(n_2490),
.A2(n_2326),
.B1(n_2332),
.B2(n_2392),
.Y(n_2592)
);

OAI22xp5_ASAP7_75t_L g2593 ( 
.A1(n_2358),
.A2(n_2326),
.B1(n_2377),
.B2(n_2466),
.Y(n_2593)
);

INVx1_ASAP7_75t_L g2594 ( 
.A(n_2460),
.Y(n_2594)
);

BUFx2_ASAP7_75t_L g2595 ( 
.A(n_2454),
.Y(n_2595)
);

BUFx8_ASAP7_75t_SL g2596 ( 
.A(n_2418),
.Y(n_2596)
);

NAND2x1p5_ASAP7_75t_L g2597 ( 
.A(n_2446),
.B(n_2492),
.Y(n_2597)
);

BUFx4_ASAP7_75t_SL g2598 ( 
.A(n_2457),
.Y(n_2598)
);

BUFx2_ASAP7_75t_L g2599 ( 
.A(n_2371),
.Y(n_2599)
);

INVx4_ASAP7_75t_L g2600 ( 
.A(n_2420),
.Y(n_2600)
);

NAND2xp5_ASAP7_75t_L g2601 ( 
.A(n_2387),
.B(n_2478),
.Y(n_2601)
);

AOI22xp33_ASAP7_75t_SL g2602 ( 
.A1(n_2485),
.A2(n_2416),
.B1(n_2350),
.B2(n_2435),
.Y(n_2602)
);

INVx1_ASAP7_75t_L g2603 ( 
.A(n_2457),
.Y(n_2603)
);

CKINVDCx20_ASAP7_75t_R g2604 ( 
.A(n_2480),
.Y(n_2604)
);

AOI22xp33_ASAP7_75t_L g2605 ( 
.A1(n_2452),
.A2(n_2382),
.B1(n_2486),
.B2(n_2464),
.Y(n_2605)
);

INVx1_ASAP7_75t_L g2606 ( 
.A(n_2457),
.Y(n_2606)
);

INVx1_ASAP7_75t_L g2607 ( 
.A(n_2471),
.Y(n_2607)
);

BUFx2_ASAP7_75t_SL g2608 ( 
.A(n_2482),
.Y(n_2608)
);

INVx5_ASAP7_75t_L g2609 ( 
.A(n_2491),
.Y(n_2609)
);

INVx1_ASAP7_75t_L g2610 ( 
.A(n_2448),
.Y(n_2610)
);

CKINVDCx5p33_ASAP7_75t_R g2611 ( 
.A(n_2458),
.Y(n_2611)
);

NAND2xp5_ASAP7_75t_L g2612 ( 
.A(n_2587),
.B(n_2603),
.Y(n_2612)
);

INVx3_ASAP7_75t_L g2613 ( 
.A(n_2548),
.Y(n_2613)
);

AO21x2_ASAP7_75t_L g2614 ( 
.A1(n_2593),
.A2(n_2353),
.B(n_2380),
.Y(n_2614)
);

INVx2_ASAP7_75t_L g2615 ( 
.A(n_2610),
.Y(n_2615)
);

INVx1_ASAP7_75t_L g2616 ( 
.A(n_2594),
.Y(n_2616)
);

INVx2_ASAP7_75t_SL g2617 ( 
.A(n_2502),
.Y(n_2617)
);

OAI21xp33_ASAP7_75t_SL g2618 ( 
.A1(n_2497),
.A2(n_2502),
.B(n_2500),
.Y(n_2618)
);

AO21x2_ASAP7_75t_L g2619 ( 
.A1(n_2607),
.A2(n_2404),
.B(n_2372),
.Y(n_2619)
);

INVx1_ASAP7_75t_L g2620 ( 
.A(n_2505),
.Y(n_2620)
);

INVx1_ASAP7_75t_L g2621 ( 
.A(n_2507),
.Y(n_2621)
);

BUFx3_ASAP7_75t_L g2622 ( 
.A(n_2581),
.Y(n_2622)
);

HB1xp67_ASAP7_75t_L g2623 ( 
.A(n_2535),
.Y(n_2623)
);

NAND2xp5_ASAP7_75t_L g2624 ( 
.A(n_2587),
.B(n_2606),
.Y(n_2624)
);

INVx1_ASAP7_75t_L g2625 ( 
.A(n_2521),
.Y(n_2625)
);

AND2x2_ASAP7_75t_L g2626 ( 
.A(n_2582),
.B(n_2366),
.Y(n_2626)
);

INVx1_ASAP7_75t_L g2627 ( 
.A(n_2528),
.Y(n_2627)
);

INVxp33_ASAP7_75t_L g2628 ( 
.A(n_2509),
.Y(n_2628)
);

INVx6_ASAP7_75t_L g2629 ( 
.A(n_2575),
.Y(n_2629)
);

OAI22xp5_ASAP7_75t_L g2630 ( 
.A1(n_2500),
.A2(n_2378),
.B1(n_2470),
.B2(n_2459),
.Y(n_2630)
);

AND2x4_ASAP7_75t_L g2631 ( 
.A(n_2548),
.B(n_2549),
.Y(n_2631)
);

HB1xp67_ASAP7_75t_L g2632 ( 
.A(n_2557),
.Y(n_2632)
);

HB1xp67_ASAP7_75t_L g2633 ( 
.A(n_2599),
.Y(n_2633)
);

CKINVDCx5p33_ASAP7_75t_R g2634 ( 
.A(n_2501),
.Y(n_2634)
);

BUFx2_ASAP7_75t_L g2635 ( 
.A(n_2537),
.Y(n_2635)
);

INVx2_ASAP7_75t_L g2636 ( 
.A(n_2541),
.Y(n_2636)
);

AOI22xp33_ASAP7_75t_L g2637 ( 
.A1(n_2510),
.A2(n_2462),
.B1(n_2412),
.B2(n_2438),
.Y(n_2637)
);

AND2x4_ASAP7_75t_L g2638 ( 
.A(n_2600),
.B(n_2366),
.Y(n_2638)
);

INVx2_ASAP7_75t_L g2639 ( 
.A(n_2558),
.Y(n_2639)
);

INVx2_ASAP7_75t_L g2640 ( 
.A(n_2560),
.Y(n_2640)
);

OAI21x1_ASAP7_75t_L g2641 ( 
.A1(n_2579),
.A2(n_2437),
.B(n_2494),
.Y(n_2641)
);

AOI21x1_ASAP7_75t_L g2642 ( 
.A1(n_2559),
.A2(n_2409),
.B(n_2488),
.Y(n_2642)
);

INVx1_ASAP7_75t_L g2643 ( 
.A(n_2530),
.Y(n_2643)
);

BUFx6f_ASAP7_75t_L g2644 ( 
.A(n_2531),
.Y(n_2644)
);

INVx1_ASAP7_75t_L g2645 ( 
.A(n_2538),
.Y(n_2645)
);

INVx2_ASAP7_75t_L g2646 ( 
.A(n_2554),
.Y(n_2646)
);

INVx1_ASAP7_75t_L g2647 ( 
.A(n_2563),
.Y(n_2647)
);

INVx1_ASAP7_75t_L g2648 ( 
.A(n_2533),
.Y(n_2648)
);

AND2x4_ASAP7_75t_L g2649 ( 
.A(n_2600),
.B(n_2366),
.Y(n_2649)
);

INVx1_ASAP7_75t_L g2650 ( 
.A(n_2534),
.Y(n_2650)
);

NOR2xp33_ASAP7_75t_L g2651 ( 
.A(n_2583),
.B(n_2453),
.Y(n_2651)
);

AOI22xp33_ASAP7_75t_L g2652 ( 
.A1(n_2510),
.A2(n_2443),
.B1(n_2385),
.B2(n_2363),
.Y(n_2652)
);

INVx3_ASAP7_75t_L g2653 ( 
.A(n_2609),
.Y(n_2653)
);

INVx3_ASAP7_75t_L g2654 ( 
.A(n_2609),
.Y(n_2654)
);

AND2x2_ASAP7_75t_L g2655 ( 
.A(n_2580),
.B(n_2469),
.Y(n_2655)
);

INVx1_ASAP7_75t_L g2656 ( 
.A(n_2590),
.Y(n_2656)
);

INVx1_ASAP7_75t_L g2657 ( 
.A(n_2570),
.Y(n_2657)
);

NOR2xp33_ASAP7_75t_L g2658 ( 
.A(n_2596),
.B(n_2475),
.Y(n_2658)
);

INVx1_ASAP7_75t_L g2659 ( 
.A(n_2568),
.Y(n_2659)
);

INVx3_ASAP7_75t_L g2660 ( 
.A(n_2609),
.Y(n_2660)
);

AND2x2_ASAP7_75t_L g2661 ( 
.A(n_2577),
.B(n_2469),
.Y(n_2661)
);

OAI21x1_ASAP7_75t_L g2662 ( 
.A1(n_2525),
.A2(n_2397),
.B(n_2354),
.Y(n_2662)
);

OAI21xp5_ASAP7_75t_L g2663 ( 
.A1(n_2545),
.A2(n_2391),
.B(n_2495),
.Y(n_2663)
);

INVx2_ASAP7_75t_SL g2664 ( 
.A(n_2537),
.Y(n_2664)
);

CKINVDCx5p33_ASAP7_75t_R g2665 ( 
.A(n_2526),
.Y(n_2665)
);

INVx2_ASAP7_75t_L g2666 ( 
.A(n_2589),
.Y(n_2666)
);

INVx1_ASAP7_75t_L g2667 ( 
.A(n_2574),
.Y(n_2667)
);

BUFx8_ASAP7_75t_SL g2668 ( 
.A(n_2506),
.Y(n_2668)
);

OA21x2_ASAP7_75t_L g2669 ( 
.A1(n_2605),
.A2(n_2601),
.B(n_2436),
.Y(n_2669)
);

INVx1_ASAP7_75t_L g2670 ( 
.A(n_2573),
.Y(n_2670)
);

INVx2_ASAP7_75t_L g2671 ( 
.A(n_2531),
.Y(n_2671)
);

AND2x4_ASAP7_75t_L g2672 ( 
.A(n_2531),
.B(n_2374),
.Y(n_2672)
);

AND2x2_ASAP7_75t_L g2673 ( 
.A(n_2602),
.B(n_2469),
.Y(n_2673)
);

INVx1_ASAP7_75t_L g2674 ( 
.A(n_2598),
.Y(n_2674)
);

INVx1_ASAP7_75t_L g2675 ( 
.A(n_2514),
.Y(n_2675)
);

INVx1_ASAP7_75t_L g2676 ( 
.A(n_2608),
.Y(n_2676)
);

INVx1_ASAP7_75t_L g2677 ( 
.A(n_2595),
.Y(n_2677)
);

INVx1_ASAP7_75t_L g2678 ( 
.A(n_2499),
.Y(n_2678)
);

INVx2_ASAP7_75t_L g2679 ( 
.A(n_2552),
.Y(n_2679)
);

INVxp67_ASAP7_75t_L g2680 ( 
.A(n_2635),
.Y(n_2680)
);

AND2x2_ASAP7_75t_L g2681 ( 
.A(n_2626),
.B(n_2524),
.Y(n_2681)
);

OR2x2_ASAP7_75t_L g2682 ( 
.A(n_2623),
.B(n_2511),
.Y(n_2682)
);

AND2x2_ASAP7_75t_L g2683 ( 
.A(n_2626),
.B(n_2604),
.Y(n_2683)
);

INVx1_ASAP7_75t_L g2684 ( 
.A(n_2646),
.Y(n_2684)
);

OR2x6_ASAP7_75t_L g2685 ( 
.A(n_2674),
.B(n_2581),
.Y(n_2685)
);

AND2x2_ASAP7_75t_L g2686 ( 
.A(n_2655),
.B(n_2584),
.Y(n_2686)
);

AND2x2_ASAP7_75t_L g2687 ( 
.A(n_2655),
.B(n_2586),
.Y(n_2687)
);

OA21x2_ASAP7_75t_L g2688 ( 
.A1(n_2662),
.A2(n_2559),
.B(n_2539),
.Y(n_2688)
);

INVx1_ASAP7_75t_L g2689 ( 
.A(n_2646),
.Y(n_2689)
);

AND2x2_ASAP7_75t_L g2690 ( 
.A(n_2661),
.B(n_2511),
.Y(n_2690)
);

AND2x4_ASAP7_75t_L g2691 ( 
.A(n_2672),
.B(n_2552),
.Y(n_2691)
);

AND2x2_ASAP7_75t_L g2692 ( 
.A(n_2661),
.B(n_2597),
.Y(n_2692)
);

AOI22xp5_ASAP7_75t_L g2693 ( 
.A1(n_2618),
.A2(n_2518),
.B1(n_2515),
.B2(n_2513),
.Y(n_2693)
);

INVx2_ASAP7_75t_L g2694 ( 
.A(n_2615),
.Y(n_2694)
);

CKINVDCx5p33_ASAP7_75t_R g2695 ( 
.A(n_2668),
.Y(n_2695)
);

NAND2xp5_ASAP7_75t_L g2696 ( 
.A(n_2612),
.B(n_2545),
.Y(n_2696)
);

AND2x2_ASAP7_75t_L g2697 ( 
.A(n_2615),
.B(n_2597),
.Y(n_2697)
);

OAI22xp5_ASAP7_75t_L g2698 ( 
.A1(n_2622),
.A2(n_2503),
.B1(n_2532),
.B2(n_2553),
.Y(n_2698)
);

OR2x2_ASAP7_75t_L g2699 ( 
.A(n_2632),
.B(n_2565),
.Y(n_2699)
);

AOI21xp5_ASAP7_75t_L g2700 ( 
.A1(n_2663),
.A2(n_2592),
.B(n_2430),
.Y(n_2700)
);

AND2x4_ASAP7_75t_L g2701 ( 
.A(n_2672),
.B(n_2552),
.Y(n_2701)
);

AND2x2_ASAP7_75t_L g2702 ( 
.A(n_2615),
.B(n_2571),
.Y(n_2702)
);

OAI21x1_ASAP7_75t_L g2703 ( 
.A1(n_2642),
.A2(n_2525),
.B(n_2423),
.Y(n_2703)
);

OAI21xp5_ASAP7_75t_L g2704 ( 
.A1(n_2618),
.A2(n_2550),
.B(n_2515),
.Y(n_2704)
);

OR2x2_ASAP7_75t_L g2705 ( 
.A(n_2659),
.B(n_2517),
.Y(n_2705)
);

OAI21xp5_ASAP7_75t_L g2706 ( 
.A1(n_2663),
.A2(n_2550),
.B(n_2523),
.Y(n_2706)
);

AND2x2_ASAP7_75t_L g2707 ( 
.A(n_2639),
.B(n_2571),
.Y(n_2707)
);

INVx1_ASAP7_75t_L g2708 ( 
.A(n_2646),
.Y(n_2708)
);

NAND3xp33_ASAP7_75t_L g2709 ( 
.A(n_2637),
.B(n_2512),
.C(n_2566),
.Y(n_2709)
);

AND2x2_ASAP7_75t_L g2710 ( 
.A(n_2639),
.B(n_2571),
.Y(n_2710)
);

NAND2xp5_ASAP7_75t_L g2711 ( 
.A(n_2612),
.B(n_2567),
.Y(n_2711)
);

AND2x2_ASAP7_75t_L g2712 ( 
.A(n_2639),
.B(n_2499),
.Y(n_2712)
);

AND2x4_ASAP7_75t_L g2713 ( 
.A(n_2672),
.B(n_2516),
.Y(n_2713)
);

AND2x2_ASAP7_75t_L g2714 ( 
.A(n_2640),
.B(n_2516),
.Y(n_2714)
);

INVx1_ASAP7_75t_L g2715 ( 
.A(n_2640),
.Y(n_2715)
);

INVx3_ASAP7_75t_L g2716 ( 
.A(n_2653),
.Y(n_2716)
);

NOR2xp33_ASAP7_75t_L g2717 ( 
.A(n_2628),
.B(n_2520),
.Y(n_2717)
);

NAND2xp5_ASAP7_75t_L g2718 ( 
.A(n_2624),
.B(n_2611),
.Y(n_2718)
);

AND2x2_ASAP7_75t_SL g2719 ( 
.A(n_2635),
.B(n_2519),
.Y(n_2719)
);

NAND2x1p5_ASAP7_75t_L g2720 ( 
.A(n_2622),
.B(n_2575),
.Y(n_2720)
);

NAND2xp5_ASAP7_75t_L g2721 ( 
.A(n_2696),
.B(n_2624),
.Y(n_2721)
);

INVx1_ASAP7_75t_SL g2722 ( 
.A(n_2719),
.Y(n_2722)
);

INVx1_ASAP7_75t_L g2723 ( 
.A(n_2684),
.Y(n_2723)
);

AOI211xp5_ASAP7_75t_SL g2724 ( 
.A1(n_2698),
.A2(n_2673),
.B(n_2630),
.C(n_2658),
.Y(n_2724)
);

OR2x2_ASAP7_75t_L g2725 ( 
.A(n_2682),
.B(n_2659),
.Y(n_2725)
);

AND2x2_ASAP7_75t_L g2726 ( 
.A(n_2686),
.B(n_2673),
.Y(n_2726)
);

INVxp67_ASAP7_75t_SL g2727 ( 
.A(n_2680),
.Y(n_2727)
);

INVx3_ASAP7_75t_L g2728 ( 
.A(n_2716),
.Y(n_2728)
);

NAND2xp5_ASAP7_75t_L g2729 ( 
.A(n_2696),
.B(n_2633),
.Y(n_2729)
);

INVx2_ASAP7_75t_SL g2730 ( 
.A(n_2719),
.Y(n_2730)
);

INVx1_ASAP7_75t_L g2731 ( 
.A(n_2684),
.Y(n_2731)
);

INVx1_ASAP7_75t_L g2732 ( 
.A(n_2689),
.Y(n_2732)
);

NAND2xp5_ASAP7_75t_L g2733 ( 
.A(n_2686),
.B(n_2670),
.Y(n_2733)
);

OR2x2_ASAP7_75t_L g2734 ( 
.A(n_2682),
.B(n_2675),
.Y(n_2734)
);

INVx1_ASAP7_75t_L g2735 ( 
.A(n_2689),
.Y(n_2735)
);

OR2x2_ASAP7_75t_L g2736 ( 
.A(n_2699),
.B(n_2675),
.Y(n_2736)
);

NAND2xp5_ASAP7_75t_L g2737 ( 
.A(n_2711),
.B(n_2670),
.Y(n_2737)
);

NAND2xp5_ASAP7_75t_L g2738 ( 
.A(n_2711),
.B(n_2667),
.Y(n_2738)
);

INVx1_ASAP7_75t_L g2739 ( 
.A(n_2708),
.Y(n_2739)
);

AND2x2_ASAP7_75t_L g2740 ( 
.A(n_2690),
.B(n_2672),
.Y(n_2740)
);

HB1xp67_ASAP7_75t_L g2741 ( 
.A(n_2699),
.Y(n_2741)
);

AND2x2_ASAP7_75t_L g2742 ( 
.A(n_2690),
.B(n_2638),
.Y(n_2742)
);

AOI22xp33_ASAP7_75t_SL g2743 ( 
.A1(n_2719),
.A2(n_2674),
.B1(n_2617),
.B2(n_2664),
.Y(n_2743)
);

INVx2_ASAP7_75t_SL g2744 ( 
.A(n_2685),
.Y(n_2744)
);

INVx1_ASAP7_75t_L g2745 ( 
.A(n_2708),
.Y(n_2745)
);

INVx1_ASAP7_75t_L g2746 ( 
.A(n_2715),
.Y(n_2746)
);

AND2x2_ASAP7_75t_L g2747 ( 
.A(n_2681),
.B(n_2638),
.Y(n_2747)
);

INVxp67_ASAP7_75t_SL g2748 ( 
.A(n_2716),
.Y(n_2748)
);

OAI222xp33_ASAP7_75t_L g2749 ( 
.A1(n_2685),
.A2(n_2664),
.B1(n_2617),
.B2(n_2630),
.C1(n_2652),
.C2(n_2676),
.Y(n_2749)
);

INVx1_ASAP7_75t_L g2750 ( 
.A(n_2715),
.Y(n_2750)
);

INVx1_ASAP7_75t_L g2751 ( 
.A(n_2694),
.Y(n_2751)
);

AND2x2_ASAP7_75t_L g2752 ( 
.A(n_2681),
.B(n_2638),
.Y(n_2752)
);

INVx1_ASAP7_75t_L g2753 ( 
.A(n_2694),
.Y(n_2753)
);

AND2x2_ASAP7_75t_L g2754 ( 
.A(n_2683),
.B(n_2638),
.Y(n_2754)
);

AND2x2_ASAP7_75t_L g2755 ( 
.A(n_2683),
.B(n_2649),
.Y(n_2755)
);

INVx2_ASAP7_75t_L g2756 ( 
.A(n_2751),
.Y(n_2756)
);

BUFx2_ASAP7_75t_L g2757 ( 
.A(n_2744),
.Y(n_2757)
);

OAI322xp33_ASAP7_75t_L g2758 ( 
.A1(n_2721),
.A2(n_2693),
.A3(n_2718),
.B1(n_2698),
.B2(n_2705),
.C1(n_2717),
.C2(n_2709),
.Y(n_2758)
);

OR2x2_ASAP7_75t_L g2759 ( 
.A(n_2729),
.B(n_2725),
.Y(n_2759)
);

INVx1_ASAP7_75t_L g2760 ( 
.A(n_2723),
.Y(n_2760)
);

INVxp67_ASAP7_75t_L g2761 ( 
.A(n_2727),
.Y(n_2761)
);

OR2x2_ASAP7_75t_L g2762 ( 
.A(n_2725),
.B(n_2705),
.Y(n_2762)
);

AND2x2_ASAP7_75t_L g2763 ( 
.A(n_2726),
.B(n_2687),
.Y(n_2763)
);

NAND2xp5_ASAP7_75t_L g2764 ( 
.A(n_2737),
.B(n_2718),
.Y(n_2764)
);

INVx2_ASAP7_75t_L g2765 ( 
.A(n_2751),
.Y(n_2765)
);

INVx2_ASAP7_75t_L g2766 ( 
.A(n_2753),
.Y(n_2766)
);

INVx2_ASAP7_75t_L g2767 ( 
.A(n_2753),
.Y(n_2767)
);

AND2x2_ASAP7_75t_L g2768 ( 
.A(n_2726),
.B(n_2687),
.Y(n_2768)
);

INVx1_ASAP7_75t_L g2769 ( 
.A(n_2723),
.Y(n_2769)
);

AND2x4_ASAP7_75t_L g2770 ( 
.A(n_2728),
.B(n_2716),
.Y(n_2770)
);

NAND2xp5_ASAP7_75t_L g2771 ( 
.A(n_2738),
.B(n_2669),
.Y(n_2771)
);

AND2x2_ASAP7_75t_L g2772 ( 
.A(n_2742),
.B(n_2688),
.Y(n_2772)
);

AND2x2_ASAP7_75t_L g2773 ( 
.A(n_2742),
.B(n_2740),
.Y(n_2773)
);

OR2x2_ASAP7_75t_L g2774 ( 
.A(n_2741),
.B(n_2669),
.Y(n_2774)
);

INVx2_ASAP7_75t_L g2775 ( 
.A(n_2731),
.Y(n_2775)
);

NAND2xp33_ASAP7_75t_SL g2776 ( 
.A(n_2744),
.B(n_2695),
.Y(n_2776)
);

OAI221xp5_ASAP7_75t_L g2777 ( 
.A1(n_2724),
.A2(n_2704),
.B1(n_2693),
.B2(n_2706),
.C(n_2709),
.Y(n_2777)
);

AOI22xp33_ASAP7_75t_L g2778 ( 
.A1(n_2754),
.A2(n_2704),
.B1(n_2706),
.B2(n_2651),
.Y(n_2778)
);

INVx2_ASAP7_75t_L g2779 ( 
.A(n_2731),
.Y(n_2779)
);

INVx2_ASAP7_75t_L g2780 ( 
.A(n_2732),
.Y(n_2780)
);

AND2x2_ASAP7_75t_L g2781 ( 
.A(n_2747),
.B(n_2752),
.Y(n_2781)
);

INVx1_ASAP7_75t_L g2782 ( 
.A(n_2732),
.Y(n_2782)
);

INVx1_ASAP7_75t_L g2783 ( 
.A(n_2735),
.Y(n_2783)
);

AND2x2_ASAP7_75t_L g2784 ( 
.A(n_2740),
.B(n_2688),
.Y(n_2784)
);

AND2x2_ASAP7_75t_L g2785 ( 
.A(n_2747),
.B(n_2688),
.Y(n_2785)
);

AND2x2_ASAP7_75t_L g2786 ( 
.A(n_2752),
.B(n_2692),
.Y(n_2786)
);

OR2x2_ASAP7_75t_L g2787 ( 
.A(n_2734),
.B(n_2669),
.Y(n_2787)
);

INVx1_ASAP7_75t_L g2788 ( 
.A(n_2735),
.Y(n_2788)
);

AO21x2_ASAP7_75t_L g2789 ( 
.A1(n_2749),
.A2(n_2700),
.B(n_2619),
.Y(n_2789)
);

OAI221xp5_ASAP7_75t_L g2790 ( 
.A1(n_2743),
.A2(n_2529),
.B1(n_2578),
.B2(n_2520),
.C(n_2508),
.Y(n_2790)
);

INVx4_ASAP7_75t_L g2791 ( 
.A(n_2730),
.Y(n_2791)
);

HB1xp67_ASAP7_75t_L g2792 ( 
.A(n_2746),
.Y(n_2792)
);

INVx1_ASAP7_75t_L g2793 ( 
.A(n_2792),
.Y(n_2793)
);

NOR2x1_ASAP7_75t_L g2794 ( 
.A(n_2790),
.B(n_2622),
.Y(n_2794)
);

OR2x2_ASAP7_75t_L g2795 ( 
.A(n_2787),
.B(n_2734),
.Y(n_2795)
);

AND2x2_ASAP7_75t_L g2796 ( 
.A(n_2757),
.B(n_2754),
.Y(n_2796)
);

AND2x2_ASAP7_75t_L g2797 ( 
.A(n_2757),
.B(n_2755),
.Y(n_2797)
);

AND2x2_ASAP7_75t_L g2798 ( 
.A(n_2784),
.B(n_2772),
.Y(n_2798)
);

INVx1_ASAP7_75t_L g2799 ( 
.A(n_2792),
.Y(n_2799)
);

INVx1_ASAP7_75t_L g2800 ( 
.A(n_2775),
.Y(n_2800)
);

OAI22xp5_ASAP7_75t_L g2801 ( 
.A1(n_2777),
.A2(n_2730),
.B1(n_2722),
.B2(n_2685),
.Y(n_2801)
);

NAND2xp5_ASAP7_75t_L g2802 ( 
.A(n_2761),
.B(n_2733),
.Y(n_2802)
);

HB1xp67_ASAP7_75t_L g2803 ( 
.A(n_2761),
.Y(n_2803)
);

INVx1_ASAP7_75t_L g2804 ( 
.A(n_2759),
.Y(n_2804)
);

INVx1_ASAP7_75t_L g2805 ( 
.A(n_2775),
.Y(n_2805)
);

NAND2xp5_ASAP7_75t_L g2806 ( 
.A(n_2764),
.B(n_2755),
.Y(n_2806)
);

AND2x2_ASAP7_75t_L g2807 ( 
.A(n_2784),
.B(n_2736),
.Y(n_2807)
);

NAND2xp5_ASAP7_75t_L g2808 ( 
.A(n_2764),
.B(n_2736),
.Y(n_2808)
);

OR2x2_ASAP7_75t_L g2809 ( 
.A(n_2787),
.B(n_2746),
.Y(n_2809)
);

BUFx3_ASAP7_75t_L g2810 ( 
.A(n_2790),
.Y(n_2810)
);

INVxp67_ASAP7_75t_SL g2811 ( 
.A(n_2774),
.Y(n_2811)
);

INVx1_ASAP7_75t_L g2812 ( 
.A(n_2759),
.Y(n_2812)
);

OR2x2_ASAP7_75t_L g2813 ( 
.A(n_2809),
.B(n_2771),
.Y(n_2813)
);

INVx1_ASAP7_75t_L g2814 ( 
.A(n_2803),
.Y(n_2814)
);

NAND2xp5_ASAP7_75t_L g2815 ( 
.A(n_2804),
.B(n_2778),
.Y(n_2815)
);

INVx1_ASAP7_75t_L g2816 ( 
.A(n_2812),
.Y(n_2816)
);

NAND4xp25_ASAP7_75t_SL g2817 ( 
.A(n_2794),
.B(n_2777),
.C(n_2776),
.D(n_2758),
.Y(n_2817)
);

NOR2xp33_ASAP7_75t_L g2818 ( 
.A(n_2810),
.B(n_2758),
.Y(n_2818)
);

INVx2_ASAP7_75t_L g2819 ( 
.A(n_2809),
.Y(n_2819)
);

INVx1_ASAP7_75t_L g2820 ( 
.A(n_2808),
.Y(n_2820)
);

AO22x1_ASAP7_75t_L g2821 ( 
.A1(n_2810),
.A2(n_2520),
.B1(n_2634),
.B2(n_2791),
.Y(n_2821)
);

AND2x2_ASAP7_75t_L g2822 ( 
.A(n_2807),
.B(n_2798),
.Y(n_2822)
);

INVx1_ASAP7_75t_L g2823 ( 
.A(n_2802),
.Y(n_2823)
);

INVx1_ASAP7_75t_L g2824 ( 
.A(n_2795),
.Y(n_2824)
);

INVx3_ASAP7_75t_L g2825 ( 
.A(n_2795),
.Y(n_2825)
);

INVx1_ASAP7_75t_L g2826 ( 
.A(n_2793),
.Y(n_2826)
);

INVx1_ASAP7_75t_L g2827 ( 
.A(n_2793),
.Y(n_2827)
);

AND2x2_ASAP7_75t_L g2828 ( 
.A(n_2807),
.B(n_2784),
.Y(n_2828)
);

INVx1_ASAP7_75t_L g2829 ( 
.A(n_2799),
.Y(n_2829)
);

NOR5xp2_ASAP7_75t_L g2830 ( 
.A(n_2811),
.B(n_2748),
.C(n_2789),
.D(n_2676),
.E(n_2783),
.Y(n_2830)
);

INVx3_ASAP7_75t_R g2831 ( 
.A(n_2801),
.Y(n_2831)
);

AND2x2_ASAP7_75t_L g2832 ( 
.A(n_2798),
.B(n_2772),
.Y(n_2832)
);

AND2x2_ASAP7_75t_L g2833 ( 
.A(n_2796),
.B(n_2772),
.Y(n_2833)
);

AND2x2_ASAP7_75t_L g2834 ( 
.A(n_2796),
.B(n_2785),
.Y(n_2834)
);

INVx2_ASAP7_75t_L g2835 ( 
.A(n_2825),
.Y(n_2835)
);

INVx1_ASAP7_75t_SL g2836 ( 
.A(n_2814),
.Y(n_2836)
);

OAI21xp33_ASAP7_75t_L g2837 ( 
.A1(n_2817),
.A2(n_2818),
.B(n_2815),
.Y(n_2837)
);

NAND2xp5_ASAP7_75t_L g2838 ( 
.A(n_2823),
.B(n_2785),
.Y(n_2838)
);

OR2x2_ASAP7_75t_L g2839 ( 
.A(n_2824),
.B(n_2771),
.Y(n_2839)
);

AND2x2_ASAP7_75t_L g2840 ( 
.A(n_2822),
.B(n_2797),
.Y(n_2840)
);

OR2x2_ASAP7_75t_L g2841 ( 
.A(n_2813),
.B(n_2799),
.Y(n_2841)
);

INVx2_ASAP7_75t_L g2842 ( 
.A(n_2825),
.Y(n_2842)
);

INVx1_ASAP7_75t_L g2843 ( 
.A(n_2825),
.Y(n_2843)
);

NOR2x1_ASAP7_75t_L g2844 ( 
.A(n_2826),
.B(n_2546),
.Y(n_2844)
);

NAND2xp5_ASAP7_75t_L g2845 ( 
.A(n_2820),
.B(n_2785),
.Y(n_2845)
);

AND2x2_ASAP7_75t_L g2846 ( 
.A(n_2822),
.B(n_2797),
.Y(n_2846)
);

INVx1_ASAP7_75t_L g2847 ( 
.A(n_2816),
.Y(n_2847)
);

NOR2x1p5_ASAP7_75t_L g2848 ( 
.A(n_2831),
.B(n_2791),
.Y(n_2848)
);

INVx2_ASAP7_75t_SL g2849 ( 
.A(n_2821),
.Y(n_2849)
);

INVx2_ASAP7_75t_L g2850 ( 
.A(n_2819),
.Y(n_2850)
);

AND2x2_ASAP7_75t_L g2851 ( 
.A(n_2833),
.B(n_2763),
.Y(n_2851)
);

INVx1_ASAP7_75t_SL g2852 ( 
.A(n_2836),
.Y(n_2852)
);

INVx1_ASAP7_75t_L g2853 ( 
.A(n_2843),
.Y(n_2853)
);

AND2x4_ASAP7_75t_L g2854 ( 
.A(n_2844),
.B(n_2819),
.Y(n_2854)
);

OAI22xp33_ASAP7_75t_SL g2855 ( 
.A1(n_2849),
.A2(n_2831),
.B1(n_2829),
.B2(n_2827),
.Y(n_2855)
);

OAI22xp5_ASAP7_75t_L g2856 ( 
.A1(n_2848),
.A2(n_2849),
.B1(n_2837),
.B2(n_2838),
.Y(n_2856)
);

INVxp67_ASAP7_75t_SL g2857 ( 
.A(n_2835),
.Y(n_2857)
);

INVx1_ASAP7_75t_SL g2858 ( 
.A(n_2835),
.Y(n_2858)
);

OAI21xp5_ASAP7_75t_L g2859 ( 
.A1(n_2842),
.A2(n_2834),
.B(n_2833),
.Y(n_2859)
);

INVx1_ASAP7_75t_L g2860 ( 
.A(n_2842),
.Y(n_2860)
);

AOI22xp5_ASAP7_75t_L g2861 ( 
.A1(n_2840),
.A2(n_2821),
.B1(n_2789),
.B2(n_2834),
.Y(n_2861)
);

INVx1_ASAP7_75t_L g2862 ( 
.A(n_2850),
.Y(n_2862)
);

NAND2xp5_ASAP7_75t_L g2863 ( 
.A(n_2840),
.B(n_2832),
.Y(n_2863)
);

NAND2xp5_ASAP7_75t_SL g2864 ( 
.A(n_2850),
.B(n_2791),
.Y(n_2864)
);

AOI22x1_ASAP7_75t_L g2865 ( 
.A1(n_2847),
.A2(n_2665),
.B1(n_2841),
.B2(n_2846),
.Y(n_2865)
);

OAI221xp5_ASAP7_75t_L g2866 ( 
.A1(n_2841),
.A2(n_2791),
.B1(n_2813),
.B2(n_2774),
.C(n_2832),
.Y(n_2866)
);

INVx1_ASAP7_75t_L g2867 ( 
.A(n_2839),
.Y(n_2867)
);

INVxp67_ASAP7_75t_SL g2868 ( 
.A(n_2857),
.Y(n_2868)
);

INVx2_ASAP7_75t_L g2869 ( 
.A(n_2862),
.Y(n_2869)
);

INVx1_ASAP7_75t_L g2870 ( 
.A(n_2852),
.Y(n_2870)
);

AOI22xp33_ASAP7_75t_L g2871 ( 
.A1(n_2852),
.A2(n_2846),
.B1(n_2789),
.B2(n_2845),
.Y(n_2871)
);

INVx1_ASAP7_75t_SL g2872 ( 
.A(n_2858),
.Y(n_2872)
);

INVxp67_ASAP7_75t_L g2873 ( 
.A(n_2856),
.Y(n_2873)
);

OAI221xp5_ASAP7_75t_L g2874 ( 
.A1(n_2865),
.A2(n_2851),
.B1(n_2700),
.B2(n_2527),
.C(n_2828),
.Y(n_2874)
);

INVx1_ASAP7_75t_L g2875 ( 
.A(n_2860),
.Y(n_2875)
);

NAND2xp5_ASAP7_75t_SL g2876 ( 
.A(n_2855),
.B(n_2498),
.Y(n_2876)
);

NOR3xp33_ASAP7_75t_SL g2877 ( 
.A(n_2866),
.B(n_2853),
.C(n_2864),
.Y(n_2877)
);

NAND2xp5_ASAP7_75t_L g2878 ( 
.A(n_2867),
.B(n_2851),
.Y(n_2878)
);

O2A1O1Ixp5_ASAP7_75t_L g2879 ( 
.A1(n_2859),
.A2(n_2854),
.B(n_2863),
.C(n_2861),
.Y(n_2879)
);

AND2x2_ASAP7_75t_L g2880 ( 
.A(n_2854),
.B(n_2828),
.Y(n_2880)
);

OAI22xp5_ASAP7_75t_L g2881 ( 
.A1(n_2852),
.A2(n_2806),
.B1(n_2763),
.B2(n_2768),
.Y(n_2881)
);

AOI21xp33_ASAP7_75t_L g2882 ( 
.A1(n_2852),
.A2(n_2789),
.B(n_2504),
.Y(n_2882)
);

NAND2xp5_ASAP7_75t_SL g2883 ( 
.A(n_2873),
.B(n_2498),
.Y(n_2883)
);

INVx1_ASAP7_75t_L g2884 ( 
.A(n_2868),
.Y(n_2884)
);

INVx1_ASAP7_75t_SL g2885 ( 
.A(n_2872),
.Y(n_2885)
);

INVx1_ASAP7_75t_L g2886 ( 
.A(n_2870),
.Y(n_2886)
);

XOR2x2_ASAP7_75t_L g2887 ( 
.A(n_2876),
.B(n_2561),
.Y(n_2887)
);

INVx1_ASAP7_75t_L g2888 ( 
.A(n_2869),
.Y(n_2888)
);

OR2x2_ASAP7_75t_L g2889 ( 
.A(n_2878),
.B(n_2762),
.Y(n_2889)
);

INVx1_ASAP7_75t_L g2890 ( 
.A(n_2869),
.Y(n_2890)
);

INVxp33_ASAP7_75t_L g2891 ( 
.A(n_2876),
.Y(n_2891)
);

XOR2x2_ASAP7_75t_L g2892 ( 
.A(n_2874),
.B(n_2564),
.Y(n_2892)
);

O2A1O1Ixp33_ASAP7_75t_L g2893 ( 
.A1(n_2879),
.A2(n_2875),
.B(n_2877),
.C(n_2882),
.Y(n_2893)
);

INVx1_ASAP7_75t_L g2894 ( 
.A(n_2880),
.Y(n_2894)
);

NAND2xp5_ASAP7_75t_L g2895 ( 
.A(n_2881),
.B(n_2768),
.Y(n_2895)
);

INVx1_ASAP7_75t_L g2896 ( 
.A(n_2871),
.Y(n_2896)
);

INVxp67_ASAP7_75t_SL g2897 ( 
.A(n_2871),
.Y(n_2897)
);

AOI22xp5_ASAP7_75t_L g2898 ( 
.A1(n_2873),
.A2(n_2542),
.B1(n_2556),
.B2(n_2536),
.Y(n_2898)
);

OAI211xp5_ASAP7_75t_L g2899 ( 
.A1(n_2873),
.A2(n_2547),
.B(n_2830),
.C(n_2519),
.Y(n_2899)
);

AOI222xp33_ASAP7_75t_L g2900 ( 
.A1(n_2873),
.A2(n_2576),
.B1(n_2800),
.B2(n_2805),
.C1(n_2527),
.C2(n_2770),
.Y(n_2900)
);

INVx1_ASAP7_75t_L g2901 ( 
.A(n_2884),
.Y(n_2901)
);

NAND2xp5_ASAP7_75t_L g2902 ( 
.A(n_2885),
.B(n_2800),
.Y(n_2902)
);

NOR2x1_ASAP7_75t_L g2903 ( 
.A(n_2885),
.B(n_2805),
.Y(n_2903)
);

OAI211xp5_ASAP7_75t_L g2904 ( 
.A1(n_2893),
.A2(n_2540),
.B(n_2543),
.C(n_2522),
.Y(n_2904)
);

NAND2xp5_ASAP7_75t_L g2905 ( 
.A(n_2897),
.B(n_2760),
.Y(n_2905)
);

NAND2xp5_ASAP7_75t_SL g2906 ( 
.A(n_2891),
.B(n_2770),
.Y(n_2906)
);

NAND2xp5_ASAP7_75t_L g2907 ( 
.A(n_2894),
.B(n_2896),
.Y(n_2907)
);

NAND4xp25_ASAP7_75t_L g2908 ( 
.A(n_2900),
.B(n_2523),
.C(n_2551),
.D(n_2770),
.Y(n_2908)
);

AOI211xp5_ASAP7_75t_L g2909 ( 
.A1(n_2883),
.A2(n_2544),
.B(n_2770),
.C(n_2516),
.Y(n_2909)
);

XOR2x2_ASAP7_75t_L g2910 ( 
.A(n_2887),
.B(n_2892),
.Y(n_2910)
);

NAND2xp5_ASAP7_75t_L g2911 ( 
.A(n_2886),
.B(n_2760),
.Y(n_2911)
);

HB1xp67_ASAP7_75t_L g2912 ( 
.A(n_2888),
.Y(n_2912)
);

NAND4xp25_ASAP7_75t_L g2913 ( 
.A(n_2898),
.B(n_2762),
.C(n_2508),
.D(n_2588),
.Y(n_2913)
);

INVx1_ASAP7_75t_SL g2914 ( 
.A(n_2890),
.Y(n_2914)
);

NAND2xp5_ASAP7_75t_L g2915 ( 
.A(n_2895),
.B(n_2769),
.Y(n_2915)
);

AOI211xp5_ASAP7_75t_L g2916 ( 
.A1(n_2914),
.A2(n_2899),
.B(n_2889),
.C(n_2544),
.Y(n_2916)
);

NOR2xp33_ASAP7_75t_R g2917 ( 
.A(n_2901),
.B(n_2585),
.Y(n_2917)
);

OAI211xp5_ASAP7_75t_L g2918 ( 
.A1(n_2907),
.A2(n_2728),
.B(n_2688),
.C(n_2575),
.Y(n_2918)
);

AOI221xp5_ASAP7_75t_L g2919 ( 
.A1(n_2912),
.A2(n_2902),
.B1(n_2905),
.B2(n_2911),
.C(n_2906),
.Y(n_2919)
);

AOI22xp5_ASAP7_75t_L g2920 ( 
.A1(n_2910),
.A2(n_2913),
.B1(n_2904),
.B2(n_2909),
.Y(n_2920)
);

NAND5xp2_ASAP7_75t_L g2921 ( 
.A(n_2915),
.B(n_2720),
.C(n_2642),
.D(n_2555),
.E(n_2572),
.Y(n_2921)
);

NOR2x1_ASAP7_75t_L g2922 ( 
.A(n_2903),
.B(n_2685),
.Y(n_2922)
);

AND2x4_ASAP7_75t_L g2923 ( 
.A(n_2908),
.B(n_2685),
.Y(n_2923)
);

AOI221xp5_ASAP7_75t_L g2924 ( 
.A1(n_2914),
.A2(n_2728),
.B1(n_2783),
.B2(n_2782),
.C(n_2769),
.Y(n_2924)
);

OAI222xp33_ASAP7_75t_L g2925 ( 
.A1(n_2914),
.A2(n_2720),
.B1(n_2569),
.B2(n_2728),
.C1(n_2773),
.C2(n_2781),
.Y(n_2925)
);

OAI221xp5_ASAP7_75t_SL g2926 ( 
.A1(n_2914),
.A2(n_2716),
.B1(n_2773),
.B2(n_2781),
.C(n_2786),
.Y(n_2926)
);

AOI221xp5_ASAP7_75t_SL g2927 ( 
.A1(n_2914),
.A2(n_2773),
.B1(n_2786),
.B2(n_2782),
.C(n_2788),
.Y(n_2927)
);

OAI21x1_ASAP7_75t_SL g2928 ( 
.A1(n_2920),
.A2(n_2669),
.B(n_2780),
.Y(n_2928)
);

NAND3xp33_ASAP7_75t_L g2929 ( 
.A(n_2919),
.B(n_2788),
.C(n_2780),
.Y(n_2929)
);

OAI22xp5_ASAP7_75t_L g2930 ( 
.A1(n_2916),
.A2(n_2720),
.B1(n_2629),
.B2(n_2562),
.Y(n_2930)
);

OAI211xp5_ASAP7_75t_L g2931 ( 
.A1(n_2917),
.A2(n_2922),
.B(n_2927),
.C(n_2924),
.Y(n_2931)
);

OAI211xp5_ASAP7_75t_SL g2932 ( 
.A1(n_2918),
.A2(n_2441),
.B(n_2406),
.C(n_2653),
.Y(n_2932)
);

AOI221xp5_ASAP7_75t_L g2933 ( 
.A1(n_2923),
.A2(n_2361),
.B1(n_2413),
.B2(n_2625),
.C(n_2627),
.Y(n_2933)
);

OAI21xp33_ASAP7_75t_SL g2934 ( 
.A1(n_2926),
.A2(n_2703),
.B(n_2779),
.Y(n_2934)
);

OAI211xp5_ASAP7_75t_SL g2935 ( 
.A1(n_2921),
.A2(n_2660),
.B(n_2653),
.C(n_2654),
.Y(n_2935)
);

AOI321xp33_ASAP7_75t_L g2936 ( 
.A1(n_2925),
.A2(n_2631),
.A3(n_2713),
.B1(n_2677),
.B2(n_2701),
.C(n_2691),
.Y(n_2936)
);

AOI211x1_ASAP7_75t_SL g2937 ( 
.A1(n_2927),
.A2(n_2780),
.B(n_2779),
.C(n_2775),
.Y(n_2937)
);

AOI221xp5_ASAP7_75t_L g2938 ( 
.A1(n_2919),
.A2(n_2627),
.B1(n_2625),
.B2(n_2621),
.C(n_2620),
.Y(n_2938)
);

AOI221xp5_ASAP7_75t_L g2939 ( 
.A1(n_2919),
.A2(n_2620),
.B1(n_2621),
.B2(n_2591),
.C(n_2779),
.Y(n_2939)
);

AOI21xp5_ASAP7_75t_L g2940 ( 
.A1(n_2919),
.A2(n_2766),
.B(n_2765),
.Y(n_2940)
);

AO22x2_ASAP7_75t_L g2941 ( 
.A1(n_2923),
.A2(n_2767),
.B1(n_2766),
.B2(n_2765),
.Y(n_2941)
);

OAI22xp5_ASAP7_75t_L g2942 ( 
.A1(n_2931),
.A2(n_2629),
.B1(n_2562),
.B2(n_2591),
.Y(n_2942)
);

INVx2_ASAP7_75t_SL g2943 ( 
.A(n_2930),
.Y(n_2943)
);

INVx2_ASAP7_75t_L g2944 ( 
.A(n_2941),
.Y(n_2944)
);

INVx2_ASAP7_75t_L g2945 ( 
.A(n_2941),
.Y(n_2945)
);

INVx1_ASAP7_75t_L g2946 ( 
.A(n_2928),
.Y(n_2946)
);

AOI22xp5_ASAP7_75t_L g2947 ( 
.A1(n_2935),
.A2(n_2629),
.B1(n_2581),
.B2(n_2631),
.Y(n_2947)
);

OR2x2_ASAP7_75t_L g2948 ( 
.A(n_2929),
.B(n_2756),
.Y(n_2948)
);

INVx2_ASAP7_75t_L g2949 ( 
.A(n_2936),
.Y(n_2949)
);

NOR2xp33_ASAP7_75t_L g2950 ( 
.A(n_2934),
.B(n_2629),
.Y(n_2950)
);

OAI22xp5_ASAP7_75t_L g2951 ( 
.A1(n_2939),
.A2(n_2629),
.B1(n_2766),
.B2(n_2765),
.Y(n_2951)
);

NOR2x1_ASAP7_75t_L g2952 ( 
.A(n_2940),
.B(n_2756),
.Y(n_2952)
);

NAND4xp75_ASAP7_75t_L g2953 ( 
.A(n_2933),
.B(n_2677),
.C(n_2678),
.D(n_2667),
.Y(n_2953)
);

NOR2x1p5_ASAP7_75t_L g2954 ( 
.A(n_2937),
.B(n_2613),
.Y(n_2954)
);

INVx1_ASAP7_75t_L g2955 ( 
.A(n_2932),
.Y(n_2955)
);

AND2x4_ASAP7_75t_L g2956 ( 
.A(n_2938),
.B(n_2767),
.Y(n_2956)
);

NAND4xp75_ASAP7_75t_L g2957 ( 
.A(n_2933),
.B(n_2678),
.C(n_2712),
.D(n_2647),
.Y(n_2957)
);

OR2x2_ASAP7_75t_L g2958 ( 
.A(n_2943),
.B(n_2767),
.Y(n_2958)
);

AOI32xp33_ASAP7_75t_L g2959 ( 
.A1(n_2955),
.A2(n_2631),
.A3(n_2660),
.B1(n_2654),
.B2(n_2653),
.Y(n_2959)
);

CKINVDCx12_ASAP7_75t_R g2960 ( 
.A(n_2949),
.Y(n_2960)
);

AND2x4_ASAP7_75t_L g2961 ( 
.A(n_2946),
.B(n_2954),
.Y(n_2961)
);

NAND2xp5_ASAP7_75t_L g2962 ( 
.A(n_2950),
.B(n_2756),
.Y(n_2962)
);

NOR3xp33_ASAP7_75t_L g2963 ( 
.A(n_2942),
.B(n_2654),
.C(n_2660),
.Y(n_2963)
);

INVx2_ASAP7_75t_L g2964 ( 
.A(n_2948),
.Y(n_2964)
);

NAND2xp5_ASAP7_75t_L g2965 ( 
.A(n_2944),
.B(n_2645),
.Y(n_2965)
);

NAND3xp33_ASAP7_75t_L g2966 ( 
.A(n_2945),
.B(n_2645),
.C(n_2647),
.Y(n_2966)
);

NAND3x1_ASAP7_75t_SL g2967 ( 
.A(n_2952),
.B(n_2953),
.C(n_2957),
.Y(n_2967)
);

AND2x2_ASAP7_75t_L g2968 ( 
.A(n_2956),
.B(n_2692),
.Y(n_2968)
);

AOI221xp5_ASAP7_75t_L g2969 ( 
.A1(n_2956),
.A2(n_2643),
.B1(n_2648),
.B2(n_2650),
.C(n_2654),
.Y(n_2969)
);

NOR4xp75_ASAP7_75t_L g2970 ( 
.A(n_2951),
.B(n_2613),
.C(n_2660),
.D(n_2714),
.Y(n_2970)
);

NOR2x1_ASAP7_75t_L g2971 ( 
.A(n_2947),
.B(n_2613),
.Y(n_2971)
);

NAND2xp5_ASAP7_75t_L g2972 ( 
.A(n_2961),
.B(n_2643),
.Y(n_2972)
);

AOI22xp5_ASAP7_75t_L g2973 ( 
.A1(n_2960),
.A2(n_2631),
.B1(n_2713),
.B2(n_2701),
.Y(n_2973)
);

NOR2xp33_ASAP7_75t_L g2974 ( 
.A(n_2964),
.B(n_2613),
.Y(n_2974)
);

AOI21xp5_ASAP7_75t_L g2975 ( 
.A1(n_2965),
.A2(n_2619),
.B(n_2650),
.Y(n_2975)
);

OAI211xp5_ASAP7_75t_SL g2976 ( 
.A1(n_2958),
.A2(n_2648),
.B(n_2750),
.C(n_2739),
.Y(n_2976)
);

AOI22xp5_ASAP7_75t_L g2977 ( 
.A1(n_2962),
.A2(n_2713),
.B1(n_2691),
.B2(n_2701),
.Y(n_2977)
);

XNOR2x1_ASAP7_75t_L g2978 ( 
.A(n_2970),
.B(n_2555),
.Y(n_2978)
);

OAI22xp5_ASAP7_75t_L g2979 ( 
.A1(n_2971),
.A2(n_2713),
.B1(n_2691),
.B2(n_2701),
.Y(n_2979)
);

XNOR2xp5_ASAP7_75t_L g2980 ( 
.A(n_2967),
.B(n_2691),
.Y(n_2980)
);

INVxp67_ASAP7_75t_SL g2981 ( 
.A(n_2966),
.Y(n_2981)
);

INVx4_ASAP7_75t_L g2982 ( 
.A(n_2980),
.Y(n_2982)
);

OAI22xp5_ASAP7_75t_L g2983 ( 
.A1(n_2974),
.A2(n_2968),
.B1(n_2959),
.B2(n_2969),
.Y(n_2983)
);

OA22x2_ASAP7_75t_L g2984 ( 
.A1(n_2981),
.A2(n_2963),
.B1(n_2750),
.B2(n_2745),
.Y(n_2984)
);

OAI22xp5_ASAP7_75t_L g2985 ( 
.A1(n_2978),
.A2(n_2745),
.B1(n_2739),
.B2(n_2671),
.Y(n_2985)
);

INVx1_ASAP7_75t_L g2986 ( 
.A(n_2972),
.Y(n_2986)
);

AOI22xp5_ASAP7_75t_L g2987 ( 
.A1(n_2973),
.A2(n_2619),
.B1(n_2649),
.B2(n_2614),
.Y(n_2987)
);

AO22x2_ASAP7_75t_L g2988 ( 
.A1(n_2975),
.A2(n_2656),
.B1(n_2671),
.B2(n_2679),
.Y(n_2988)
);

OAI22xp5_ASAP7_75t_L g2989 ( 
.A1(n_2977),
.A2(n_2671),
.B1(n_2679),
.B2(n_2656),
.Y(n_2989)
);

OAI221xp5_ASAP7_75t_L g2990 ( 
.A1(n_2982),
.A2(n_2976),
.B1(n_2979),
.B2(n_2644),
.C(n_2679),
.Y(n_2990)
);

NAND2xp5_ASAP7_75t_L g2991 ( 
.A(n_2986),
.B(n_2644),
.Y(n_2991)
);

INVx4_ASAP7_75t_L g2992 ( 
.A(n_2984),
.Y(n_2992)
);

OAI22x1_ASAP7_75t_L g2993 ( 
.A1(n_2987),
.A2(n_2649),
.B1(n_2712),
.B2(n_2714),
.Y(n_2993)
);

INVx1_ASAP7_75t_L g2994 ( 
.A(n_2988),
.Y(n_2994)
);

INVx1_ASAP7_75t_L g2995 ( 
.A(n_2983),
.Y(n_2995)
);

O2A1O1Ixp33_ASAP7_75t_L g2996 ( 
.A1(n_2995),
.A2(n_2985),
.B(n_2989),
.C(n_2649),
.Y(n_2996)
);

OAI22xp5_ASAP7_75t_SL g2997 ( 
.A1(n_2992),
.A2(n_2644),
.B1(n_2657),
.B2(n_2640),
.Y(n_2997)
);

AOI22x1_ASAP7_75t_L g2998 ( 
.A1(n_2994),
.A2(n_2644),
.B1(n_2707),
.B2(n_2710),
.Y(n_2998)
);

AOI22xp5_ASAP7_75t_L g2999 ( 
.A1(n_2991),
.A2(n_2990),
.B1(n_2993),
.B2(n_2619),
.Y(n_2999)
);

OA21x2_ASAP7_75t_L g3000 ( 
.A1(n_2999),
.A2(n_2703),
.B(n_2641),
.Y(n_3000)
);

INVx2_ASAP7_75t_L g3001 ( 
.A(n_2998),
.Y(n_3001)
);

OAI21xp33_ASAP7_75t_L g3002 ( 
.A1(n_2996),
.A2(n_2710),
.B(n_2707),
.Y(n_3002)
);

AOI22xp33_ASAP7_75t_L g3003 ( 
.A1(n_3002),
.A2(n_2997),
.B1(n_2644),
.B2(n_2697),
.Y(n_3003)
);

AOI22x1_ASAP7_75t_L g3004 ( 
.A1(n_3003),
.A2(n_3001),
.B1(n_3000),
.B2(n_2644),
.Y(n_3004)
);

INVx2_ASAP7_75t_L g3005 ( 
.A(n_3004),
.Y(n_3005)
);

OAI22xp33_ASAP7_75t_L g3006 ( 
.A1(n_3004),
.A2(n_2657),
.B1(n_2666),
.B2(n_2636),
.Y(n_3006)
);

OAI221xp5_ASAP7_75t_R g3007 ( 
.A1(n_3005),
.A2(n_3006),
.B1(n_2697),
.B2(n_2702),
.C(n_2703),
.Y(n_3007)
);

AOI211xp5_ASAP7_75t_L g3008 ( 
.A1(n_3007),
.A2(n_2702),
.B(n_2694),
.C(n_2616),
.Y(n_3008)
);


endmodule