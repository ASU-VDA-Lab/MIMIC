module real_jpeg_3221_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_78;
wire n_83;
wire n_249;
wire n_166;
wire n_176;
wire n_221;
wire n_215;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_237;
wire n_174;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_243;
wire n_255;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_13;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_188;
wire n_139;
wire n_142;
wire n_175;
wire n_238;
wire n_76;
wire n_67;
wire n_79;
wire n_178;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_44;
wire n_28;
wire n_267;
wire n_208;
wire n_62;
wire n_239;
wire n_162;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_172;
wire n_160;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_262;
wire n_222;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_192;
wire n_203;
wire n_100;
wire n_198;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_258;
wire n_205;
wire n_195;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_204;
wire n_158;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_241;
wire n_103;
wire n_225;
wire n_259;
wire n_232;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_167;
wire n_213;
wire n_244;
wire n_179;
wire n_216;
wire n_133;
wire n_202;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_102;
wire n_81;
wire n_85;
wire n_181;
wire n_101;
wire n_256;
wire n_182;
wire n_253;
wire n_96;
wire n_89;
wire n_16;

INVx2_ASAP7_75t_L g47 ( 
.A(n_0),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g102 ( 
.A(n_1),
.Y(n_102)
);

OAI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_2),
.A2(n_33),
.B1(n_34),
.B2(n_60),
.Y(n_59)
);

CKINVDCx14_ASAP7_75t_R g60 ( 
.A(n_2),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_2),
.A2(n_52),
.B1(n_54),
.B2(n_60),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_2),
.A2(n_46),
.B1(n_48),
.B2(n_60),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g37 ( 
.A1(n_3),
.A2(n_24),
.B1(n_25),
.B2(n_38),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_3),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_3),
.A2(n_33),
.B1(n_34),
.B2(n_38),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_3),
.A2(n_38),
.B1(n_52),
.B2(n_54),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_3),
.A2(n_38),
.B1(n_46),
.B2(n_48),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_3),
.B(n_30),
.C(n_34),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_3),
.B(n_32),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_3),
.B(n_52),
.C(n_64),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_3),
.B(n_102),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_3),
.B(n_44),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_3),
.B(n_45),
.C(n_48),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_3),
.B(n_67),
.Y(n_245)
);

BUFx4f_ASAP7_75t_L g64 ( 
.A(n_4),
.Y(n_64)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

AOI22xp33_ASAP7_75t_L g23 ( 
.A1(n_6),
.A2(n_24),
.B1(n_25),
.B2(n_28),
.Y(n_23)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

OAI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_6),
.A2(n_28),
.B1(n_33),
.B2(n_34),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_6),
.A2(n_28),
.B1(n_52),
.B2(n_54),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_6),
.A2(n_28),
.B1(n_46),
.B2(n_48),
.Y(n_170)
);

BUFx16f_ASAP7_75t_L g45 ( 
.A(n_7),
.Y(n_45)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_8),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

OAI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_10),
.A2(n_52),
.B1(n_54),
.B2(n_56),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_10),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g68 ( 
.A1(n_10),
.A2(n_33),
.B1(n_34),
.B2(n_56),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_10),
.A2(n_46),
.B1(n_48),
.B2(n_56),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_11),
.Y(n_53)
);

XOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_115),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_SL g13 ( 
.A(n_14),
.B(n_114),
.Y(n_13)
);

INVxp67_ASAP7_75t_L g14 ( 
.A(n_15),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_SL g15 ( 
.A(n_16),
.B(n_80),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_16),
.B(n_80),
.Y(n_114)
);

XNOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_74),
.Y(n_16)
);

OAI22xp5_ASAP7_75t_SL g17 ( 
.A1(n_18),
.A2(n_19),
.B1(n_70),
.B2(n_73),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

AOI22xp5_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_21),
.B1(n_39),
.B2(n_40),
.Y(n_19)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_20),
.B(n_127),
.C(n_128),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_20),
.A2(n_21),
.B1(n_127),
.B2(n_143),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_20),
.A2(n_21),
.B1(n_91),
.B2(n_172),
.Y(n_171)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_21),
.B(n_91),
.C(n_164),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_29),
.B1(n_32),
.B2(n_37),
.Y(n_21)
);

INVxp67_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

OA21x2_ASAP7_75t_L g70 ( 
.A1(n_23),
.A2(n_71),
.B(n_72),
.Y(n_70)
);

O2A1O1Ixp33_ASAP7_75t_L g29 ( 
.A1(n_24),
.A2(n_30),
.B(n_31),
.C(n_32),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_24),
.B(n_30),
.Y(n_31)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_25),
.B(n_167),
.Y(n_166)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_29),
.B(n_37),
.Y(n_72)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_29),
.Y(n_113)
);

AO22x1_ASAP7_75t_SL g32 ( 
.A1(n_30),
.A2(n_33),
.B1(n_34),
.B2(n_36),
.Y(n_32)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_30),
.Y(n_36)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_32),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g63 ( 
.A1(n_33),
.A2(n_34),
.B1(n_64),
.B2(n_65),
.Y(n_63)
);

INVx2_ASAP7_75t_SL g33 ( 
.A(n_34),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_34),
.B(n_221),
.Y(n_220)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_37),
.B(n_112),
.Y(n_111)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_SL g40 ( 
.A1(n_41),
.A2(n_57),
.B1(n_58),
.B2(n_69),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_41),
.Y(n_69)
);

MAJIxp5_ASAP7_75t_L g74 ( 
.A(n_41),
.B(n_70),
.C(n_75),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_41),
.A2(n_69),
.B1(n_75),
.B2(n_84),
.Y(n_83)
);

AND2x2_ASAP7_75t_SL g41 ( 
.A(n_42),
.B(n_55),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_43),
.B(n_50),
.Y(n_42)
);

OAI21xp5_ASAP7_75t_L g105 ( 
.A1(n_43),
.A2(n_89),
.B(n_106),
.Y(n_105)
);

OA22x2_ASAP7_75t_L g131 ( 
.A1(n_43),
.A2(n_50),
.B1(n_108),
.B2(n_132),
.Y(n_131)
);

OA22x2_ASAP7_75t_L g153 ( 
.A1(n_43),
.A2(n_50),
.B1(n_108),
.B2(n_132),
.Y(n_153)
);

AOI21xp5_ASAP7_75t_L g180 ( 
.A1(n_43),
.A2(n_50),
.B(n_108),
.Y(n_180)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

OR2x2_ASAP7_75t_L g50 ( 
.A(n_44),
.B(n_51),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_44),
.A2(n_55),
.B1(n_88),
.B2(n_90),
.Y(n_87)
);

AO22x1_ASAP7_75t_SL g44 ( 
.A1(n_45),
.A2(n_46),
.B1(n_48),
.B2(n_49),
.Y(n_44)
);

INVx11_ASAP7_75t_L g49 ( 
.A(n_45),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_L g51 ( 
.A1(n_45),
.A2(n_49),
.B1(n_52),
.B2(n_54),
.Y(n_51)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_46),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_46),
.B(n_102),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_48),
.B(n_231),
.Y(n_230)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_50),
.Y(n_90)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_52),
.Y(n_54)
);

AOI22x1_ASAP7_75t_L g66 ( 
.A1(n_52),
.A2(n_54),
.B1(n_64),
.B2(n_65),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_52),
.B(n_238),
.Y(n_237)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

CKINVDCx16_ASAP7_75t_R g57 ( 
.A(n_58),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g58 ( 
.A1(n_59),
.A2(n_61),
.B1(n_67),
.B2(n_68),
.Y(n_58)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_59),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_61),
.A2(n_67),
.B1(n_92),
.B2(n_93),
.Y(n_91)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_62),
.B(n_79),
.Y(n_78)
);

AOI21xp5_ASAP7_75t_L g154 ( 
.A1(n_62),
.A2(n_66),
.B(n_79),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_63),
.B(n_66),
.Y(n_62)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_64),
.Y(n_65)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_66),
.Y(n_67)
);

OAI21xp5_ASAP7_75t_L g75 ( 
.A1(n_66),
.A2(n_76),
.B(n_77),
.Y(n_75)
);

AO21x1_ASAP7_75t_L g127 ( 
.A1(n_67),
.A2(n_78),
.B(n_92),
.Y(n_127)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_70),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_70),
.A2(n_73),
.B1(n_82),
.B2(n_83),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_70),
.A2(n_73),
.B1(n_183),
.B2(n_184),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_70),
.A2(n_73),
.B1(n_154),
.B2(n_201),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_71),
.B(n_113),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_73),
.B(n_147),
.C(n_154),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_73),
.B(n_127),
.C(n_180),
.Y(n_179)
);

CKINVDCx14_ASAP7_75t_R g84 ( 
.A(n_75),
.Y(n_84)
);

INVxp67_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVxp67_ASAP7_75t_L g93 ( 
.A(n_79),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_81),
.B(n_85),
.C(n_94),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_81),
.A2(n_85),
.B1(n_86),
.B2(n_119),
.Y(n_118)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_81),
.Y(n_119)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_86),
.Y(n_85)
);

OAI21xp5_ASAP7_75t_L g125 ( 
.A1(n_86),
.A2(n_87),
.B(n_91),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_91),
.Y(n_86)
);

INVxp67_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_90),
.B(n_107),
.Y(n_106)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_91),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_91),
.B(n_188),
.C(n_189),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_91),
.A2(n_172),
.B1(n_214),
.B2(n_217),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_L g117 ( 
.A(n_94),
.B(n_118),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_L g94 ( 
.A1(n_95),
.A2(n_109),
.B(n_110),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_95),
.A2(n_96),
.B1(n_122),
.B2(n_123),
.Y(n_121)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_105),
.Y(n_96)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_97),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_97),
.A2(n_109),
.B1(n_110),
.B2(n_111),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_97),
.A2(n_105),
.B1(n_109),
.B2(n_145),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_98),
.B(n_104),
.Y(n_97)
);

INVxp33_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_99),
.B(n_151),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_100),
.B(n_103),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_100),
.A2(n_103),
.B1(n_104),
.B2(n_134),
.Y(n_133)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_101),
.B(n_151),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_101),
.A2(n_102),
.B1(n_151),
.B2(n_170),
.Y(n_169)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_102),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_SL g149 ( 
.A1(n_103),
.A2(n_134),
.B(n_150),
.Y(n_149)
);

OA21x2_ASAP7_75t_L g189 ( 
.A1(n_103),
.A2(n_150),
.B(n_190),
.Y(n_189)
);

CKINVDCx16_ASAP7_75t_R g145 ( 
.A(n_105),
.Y(n_145)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

CKINVDCx16_ASAP7_75t_R g110 ( 
.A(n_111),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_L g115 ( 
.A1(n_116),
.A2(n_135),
.B(n_268),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_117),
.B(n_120),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_117),
.B(n_120),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_121),
.B(n_124),
.C(n_126),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_121),
.A2(n_124),
.B1(n_125),
.B2(n_157),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_121),
.Y(n_157)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

XNOR2xp5_ASAP7_75t_L g155 ( 
.A(n_126),
.B(n_156),
.Y(n_155)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_127),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_127),
.A2(n_143),
.B1(n_180),
.B2(n_185),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_127),
.A2(n_143),
.B1(n_152),
.B2(n_153),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_127),
.B(n_152),
.C(n_253),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_128),
.A2(n_129),
.B1(n_141),
.B2(n_142),
.Y(n_140)
);

CKINVDCx16_ASAP7_75t_R g128 ( 
.A(n_129),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_133),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g203 ( 
.A1(n_130),
.A2(n_131),
.B1(n_133),
.B2(n_204),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_L g244 ( 
.A1(n_130),
.A2(n_131),
.B1(n_245),
.B2(n_246),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_L g257 ( 
.A1(n_130),
.A2(n_131),
.B1(n_218),
.B2(n_258),
.Y(n_257)
);

INVx1_ASAP7_75t_SL g130 ( 
.A(n_131),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_131),
.B(n_213),
.C(n_218),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_131),
.B(n_169),
.C(n_245),
.Y(n_250)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_133),
.Y(n_204)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

HB1xp67_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_L g137 ( 
.A1(n_138),
.A2(n_158),
.B(n_267),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_155),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_139),
.B(n_155),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_144),
.C(n_146),
.Y(n_139)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_140),
.B(n_144),
.Y(n_265)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_146),
.B(n_265),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_147),
.A2(n_148),
.B1(n_199),
.B2(n_200),
.Y(n_198)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_152),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_149),
.A2(n_152),
.B1(n_153),
.B2(n_177),
.Y(n_176)
);

CKINVDCx16_ASAP7_75t_R g177 ( 
.A(n_149),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_152),
.A2(n_153),
.B1(n_237),
.B2(n_239),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_152),
.B(n_239),
.Y(n_247)
);

INVx1_ASAP7_75t_SL g152 ( 
.A(n_153),
.Y(n_152)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_154),
.Y(n_201)
);

AOI21xp5_ASAP7_75t_L g158 ( 
.A1(n_159),
.A2(n_262),
.B(n_266),
.Y(n_158)
);

OAI211xp5_ASAP7_75t_L g159 ( 
.A1(n_160),
.A2(n_191),
.B(n_205),
.C(n_206),
.Y(n_159)
);

OR2x2_ASAP7_75t_L g160 ( 
.A(n_161),
.B(n_181),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_161),
.B(n_181),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_162),
.A2(n_163),
.B1(n_173),
.B2(n_174),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_162),
.B(n_176),
.C(n_178),
.Y(n_193)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_SL g163 ( 
.A(n_164),
.B(n_171),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_165),
.B(n_168),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g186 ( 
.A1(n_165),
.A2(n_166),
.B1(n_168),
.B2(n_169),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_166),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_168),
.A2(n_169),
.B1(n_243),
.B2(n_244),
.Y(n_242)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g232 ( 
.A(n_169),
.B(n_233),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_169),
.B(n_233),
.Y(n_234)
);

INVxp67_ASAP7_75t_L g190 ( 
.A(n_170),
.Y(n_190)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_175),
.A2(n_176),
.B1(n_178),
.B2(n_179),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_180),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_182),
.B(n_186),
.C(n_187),
.Y(n_181)
);

XOR2xp5_ASAP7_75t_L g210 ( 
.A(n_182),
.B(n_211),
.Y(n_210)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_186),
.B(n_187),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_188),
.A2(n_189),
.B1(n_215),
.B2(n_216),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_188),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_189),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_189),
.B(n_230),
.Y(n_229)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

NAND3xp33_ASAP7_75t_SL g206 ( 
.A(n_192),
.B(n_207),
.C(n_208),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_193),
.B(n_194),
.Y(n_192)
);

OR2x2_ASAP7_75t_L g205 ( 
.A(n_193),
.B(n_194),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_L g194 ( 
.A(n_195),
.B(n_196),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_195),
.B(n_197),
.C(n_203),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_197),
.A2(n_198),
.B1(n_202),
.B2(n_203),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_L g208 ( 
.A1(n_209),
.A2(n_224),
.B(n_261),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_SL g209 ( 
.A(n_210),
.B(n_212),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_210),
.B(n_212),
.Y(n_261)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_213),
.B(n_257),
.Y(n_256)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_214),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_216),
.B(n_236),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_216),
.B(n_236),
.Y(n_240)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_218),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_219),
.B(n_222),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_L g253 ( 
.A1(n_219),
.A2(n_220),
.B1(n_222),
.B2(n_223),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_220),
.Y(n_219)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

AOI21xp5_ASAP7_75t_SL g224 ( 
.A1(n_225),
.A2(n_255),
.B(n_260),
.Y(n_224)
);

OAI21xp5_ASAP7_75t_SL g225 ( 
.A1(n_226),
.A2(n_249),
.B(n_254),
.Y(n_225)
);

AOI21xp5_ASAP7_75t_L g226 ( 
.A1(n_227),
.A2(n_241),
.B(n_248),
.Y(n_226)
);

OAI21xp5_ASAP7_75t_L g227 ( 
.A1(n_228),
.A2(n_235),
.B(n_240),
.Y(n_227)
);

AOI21xp5_ASAP7_75t_L g228 ( 
.A1(n_229),
.A2(n_232),
.B(n_234),
.Y(n_228)
);

CKINVDCx16_ASAP7_75t_R g239 ( 
.A(n_237),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_242),
.B(n_247),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_242),
.B(n_247),
.Y(n_248)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_245),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_250),
.B(n_251),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_250),
.B(n_251),
.Y(n_254)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_252),
.B(n_253),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_SL g255 ( 
.A(n_256),
.B(n_259),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_256),
.B(n_259),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_263),
.B(n_264),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_263),
.B(n_264),
.Y(n_266)
);


endmodule