module fake_jpeg_870_n_233 (n_13, n_21, n_53, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_51, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_52, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_233);

input n_13;
input n_21;
input n_53;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_51;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_52;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_233;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_127;
wire n_76;
wire n_154;
wire n_205;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_155;
wire n_207;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_223;
wire n_171;
wire n_119;
wire n_69;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_143;
wire n_202;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_139;
wire n_61;
wire n_172;
wire n_173;
wire n_232;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_91;
wire n_54;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_149;
wire n_157;
wire n_87;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_96;

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_47),
.Y(n_54)
);

BUFx10_ASAP7_75t_L g55 ( 
.A(n_23),
.Y(n_55)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_53),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_4),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_34),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_17),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_5),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_43),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_45),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_41),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_46),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_2),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_6),
.Y(n_66)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_30),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_7),
.Y(n_68)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_9),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_29),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_11),
.Y(n_71)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_51),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_39),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_40),
.Y(n_74)
);

INVxp67_ASAP7_75t_L g75 ( 
.A(n_19),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_21),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_14),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_20),
.Y(n_78)
);

BUFx5_ASAP7_75t_L g79 ( 
.A(n_12),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_59),
.B(n_0),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_80),
.B(n_75),
.Y(n_100)
);

INVx5_ASAP7_75t_L g81 ( 
.A(n_67),
.Y(n_81)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_81),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_70),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_82),
.Y(n_89)
);

BUFx3_ASAP7_75t_L g83 ( 
.A(n_75),
.Y(n_83)
);

INVxp67_ASAP7_75t_SL g93 ( 
.A(n_83),
.Y(n_93)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_69),
.Y(n_84)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_84),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_70),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_85),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_73),
.Y(n_86)
);

INVx5_ASAP7_75t_L g88 ( 
.A(n_86),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_73),
.Y(n_87)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_87),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_81),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_90),
.B(n_54),
.Y(n_105)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_84),
.Y(n_91)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_91),
.Y(n_107)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_83),
.Y(n_92)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_92),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_SL g95 ( 
.A(n_82),
.B(n_60),
.Y(n_95)
);

OR2x2_ASAP7_75t_L g118 ( 
.A(n_95),
.B(n_100),
.Y(n_118)
);

INVx4_ASAP7_75t_L g97 ( 
.A(n_85),
.Y(n_97)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_97),
.Y(n_101)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_96),
.Y(n_102)
);

INVx4_ASAP7_75t_L g138 ( 
.A(n_102),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_L g103 ( 
.A1(n_91),
.A2(n_87),
.B1(n_86),
.B2(n_69),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_103),
.A2(n_72),
.B1(n_55),
.B2(n_79),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_98),
.A2(n_78),
.B1(n_77),
.B2(n_65),
.Y(n_104)
);

AND2x2_ASAP7_75t_L g121 ( 
.A(n_104),
.B(n_105),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_98),
.A2(n_78),
.B1(n_77),
.B2(n_56),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_106),
.A2(n_94),
.B1(n_67),
.B2(n_65),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_95),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_108),
.B(n_110),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_88),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_88),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_111),
.B(n_113),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_90),
.B(n_63),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_112),
.B(n_115),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_89),
.Y(n_113)
);

BUFx2_ASAP7_75t_L g114 ( 
.A(n_96),
.Y(n_114)
);

INVx3_ASAP7_75t_SL g139 ( 
.A(n_114),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_99),
.B(n_63),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_99),
.B(n_58),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_116),
.B(n_119),
.Y(n_135)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_97),
.Y(n_117)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_117),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_89),
.B(n_58),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_112),
.B(n_92),
.C(n_93),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_123),
.B(n_140),
.C(n_139),
.Y(n_158)
);

AND2x2_ASAP7_75t_L g124 ( 
.A(n_115),
.B(n_116),
.Y(n_124)
);

XNOR2xp5_ASAP7_75t_L g164 ( 
.A(n_124),
.B(n_127),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_125),
.A2(n_128),
.B1(n_131),
.B2(n_142),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_106),
.A2(n_119),
.B1(n_104),
.B2(n_118),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_126),
.A2(n_133),
.B1(n_55),
.B2(n_79),
.Y(n_144)
);

XOR2xp5_ASAP7_75t_SL g127 ( 
.A(n_118),
.B(n_109),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_105),
.A2(n_94),
.B1(n_57),
.B2(n_68),
.Y(n_128)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_107),
.Y(n_130)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_130),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_101),
.A2(n_57),
.B1(n_68),
.B2(n_56),
.Y(n_131)
);

INVx5_ASAP7_75t_L g132 ( 
.A(n_102),
.Y(n_132)
);

BUFx2_ASAP7_75t_L g150 ( 
.A(n_132),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_107),
.A2(n_64),
.B1(n_76),
.B2(n_71),
.Y(n_133)
);

AOI31xp33_ASAP7_75t_L g134 ( 
.A1(n_109),
.A2(n_64),
.A3(n_72),
.B(n_74),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_134),
.B(n_49),
.Y(n_152)
);

MAJx2_ASAP7_75t_L g136 ( 
.A(n_114),
.B(n_66),
.C(n_62),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_136),
.B(n_127),
.C(n_133),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_L g140 ( 
.A(n_117),
.B(n_55),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_101),
.B(n_61),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_141),
.B(n_1),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_143),
.B(n_152),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_144),
.A2(n_155),
.B1(n_161),
.B2(n_10),
.Y(n_170)
);

INVx6_ASAP7_75t_L g145 ( 
.A(n_137),
.Y(n_145)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_145),
.Y(n_172)
);

AO22x1_ASAP7_75t_SL g146 ( 
.A1(n_121),
.A2(n_55),
.B1(n_52),
.B2(n_50),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_146),
.B(n_13),
.Y(n_179)
);

OR2x2_ASAP7_75t_L g147 ( 
.A(n_129),
.B(n_0),
.Y(n_147)
);

CKINVDCx14_ASAP7_75t_R g176 ( 
.A(n_147),
.Y(n_176)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_120),
.Y(n_149)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_149),
.Y(n_175)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_138),
.Y(n_151)
);

INVxp67_ASAP7_75t_SL g167 ( 
.A(n_151),
.Y(n_167)
);

INVxp67_ASAP7_75t_L g153 ( 
.A(n_139),
.Y(n_153)
);

INVxp67_ASAP7_75t_L g180 ( 
.A(n_153),
.Y(n_180)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_138),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_154),
.B(n_159),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_122),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_156),
.B(n_160),
.Y(n_177)
);

INVxp33_ASAP7_75t_L g157 ( 
.A(n_121),
.Y(n_157)
);

INVx4_ASAP7_75t_SL g187 ( 
.A(n_157),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_158),
.B(n_44),
.C(n_42),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_135),
.B(n_3),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g160 ( 
.A(n_132),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_124),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_123),
.B(n_7),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_SL g178 ( 
.A(n_162),
.B(n_13),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_136),
.B(n_8),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_163),
.B(n_14),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_140),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_SL g174 ( 
.A1(n_166),
.A2(n_11),
.B(n_12),
.Y(n_174)
);

AND2x6_ASAP7_75t_L g168 ( 
.A(n_164),
.B(n_48),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_168),
.B(n_170),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_169),
.B(n_173),
.C(n_183),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g194 ( 
.A(n_174),
.B(n_178),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_179),
.A2(n_182),
.B1(n_153),
.B2(n_150),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_SL g193 ( 
.A1(n_181),
.A2(n_185),
.B(n_18),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_157),
.A2(n_15),
.B1(n_16),
.B2(n_17),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_145),
.B(n_26),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_183),
.A2(n_186),
.B1(n_16),
.B2(n_18),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_150),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_184),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_147),
.B(n_15),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_165),
.A2(n_158),
.B1(n_146),
.B2(n_148),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_188),
.B(n_180),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_187),
.A2(n_146),
.B1(n_160),
.B2(n_28),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_SL g203 ( 
.A1(n_189),
.A2(n_199),
.B(n_179),
.Y(n_203)
);

XOR2xp5_ASAP7_75t_L g190 ( 
.A(n_186),
.B(n_25),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_190),
.B(n_192),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_L g211 ( 
.A1(n_191),
.A2(n_198),
.B1(n_170),
.B2(n_167),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g192 ( 
.A(n_169),
.B(n_27),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_193),
.B(n_196),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_187),
.B(n_31),
.C(n_37),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_197),
.B(n_35),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_172),
.A2(n_19),
.B1(n_20),
.B2(n_21),
.Y(n_198)
);

AOI21xp5_ASAP7_75t_L g199 ( 
.A1(n_176),
.A2(n_33),
.B(n_36),
.Y(n_199)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_200),
.Y(n_201)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_201),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_202),
.A2(n_209),
.B1(n_211),
.B2(n_190),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_203),
.B(n_208),
.C(n_192),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_195),
.B(n_171),
.Y(n_205)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_205),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_196),
.B(n_177),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_L g216 ( 
.A(n_207),
.B(n_210),
.Y(n_216)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_197),
.Y(n_209)
);

OAI21xp5_ASAP7_75t_SL g210 ( 
.A1(n_189),
.A2(n_182),
.B(n_180),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g223 ( 
.A(n_213),
.B(n_217),
.Y(n_223)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_215),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_204),
.B(n_194),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_SL g218 ( 
.A(n_204),
.B(n_175),
.Y(n_218)
);

OAI21xp5_ASAP7_75t_SL g220 ( 
.A1(n_218),
.A2(n_219),
.B(n_203),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_206),
.B(n_174),
.C(n_168),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_220),
.B(n_216),
.C(n_221),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_214),
.A2(n_210),
.B1(n_23),
.B2(n_24),
.Y(n_222)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_222),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_224),
.B(n_223),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_226),
.B(n_225),
.Y(n_227)
);

OAI21xp5_ASAP7_75t_SL g228 ( 
.A1(n_227),
.A2(n_212),
.B(n_222),
.Y(n_228)
);

NAND3xp33_ASAP7_75t_SL g229 ( 
.A(n_228),
.B(n_218),
.C(n_24),
.Y(n_229)
);

AND2x2_ASAP7_75t_L g230 ( 
.A(n_229),
.B(n_22),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_230),
.Y(n_231)
);

AOI21xp5_ASAP7_75t_L g232 ( 
.A1(n_231),
.A2(n_32),
.B(n_38),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_232),
.B(n_22),
.Y(n_233)
);


endmodule