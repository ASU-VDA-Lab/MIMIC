module real_jpeg_24003_n_10 (n_5, n_4, n_8, n_0, n_1, n_2, n_6, n_7, n_3, n_9, n_10);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_2;
input n_6;
input n_7;
input n_3;
input n_9;

output n_10;

wire n_108;
wire n_54;
wire n_37;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_104;
wire n_64;
wire n_11;
wire n_47;
wire n_131;
wire n_22;
wire n_87;
wire n_40;
wire n_105;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_140;
wire n_126;
wire n_13;
wire n_113;
wire n_120;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_142;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_147;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_62;
wire n_121;
wire n_106;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_69;
wire n_31;
wire n_137;
wire n_129;
wire n_135;
wire n_134;
wire n_72;
wire n_100;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_117;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_30;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_12;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_128;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_101;
wire n_96;
wire n_89;
wire n_16;

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_1),
.Y(n_58)
);

BUFx8_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

BUFx10_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_SL g28 ( 
.A1(n_4),
.A2(n_29),
.B1(n_30),
.B2(n_31),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_4),
.Y(n_30)
);

AOI22xp33_ASAP7_75t_SL g42 ( 
.A1(n_4),
.A2(n_23),
.B1(n_25),
.B2(n_30),
.Y(n_42)
);

OAI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_4),
.A2(n_30),
.B1(n_48),
.B2(n_50),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_4),
.A2(n_30),
.B1(n_77),
.B2(n_78),
.Y(n_76)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_5),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_6),
.B(n_21),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_L g37 ( 
.A1(n_6),
.A2(n_29),
.B1(n_31),
.B2(n_38),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_6),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_SL g52 ( 
.A1(n_6),
.A2(n_23),
.B1(n_25),
.B2(n_38),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_6),
.A2(n_38),
.B1(n_48),
.B2(n_50),
.Y(n_62)
);

MAJIxp5_ASAP7_75t_L g66 ( 
.A(n_6),
.B(n_45),
.C(n_48),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_6),
.A2(n_38),
.B1(n_77),
.B2(n_81),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_6),
.B(n_22),
.C(n_25),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_6),
.B(n_29),
.C(n_58),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_6),
.B(n_32),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_6),
.B(n_61),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_6),
.B(n_51),
.Y(n_134)
);

INVx13_ASAP7_75t_L g77 ( 
.A(n_7),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_L g83 ( 
.A1(n_7),
.A2(n_22),
.B1(n_26),
.B2(n_77),
.Y(n_83)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_8),
.Y(n_49)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_9),
.Y(n_36)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_9),
.Y(n_105)
);

XNOR2xp5_ASAP7_75t_L g10 ( 
.A(n_11),
.B(n_108),
.Y(n_10)
);

NAND2xp5_ASAP7_75t_SL g11 ( 
.A(n_12),
.B(n_107),
.Y(n_11)
);

INVxp67_ASAP7_75t_L g12 ( 
.A(n_13),
.Y(n_12)
);

NOR2xp33_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_71),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_14),
.B(n_71),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_54),
.C(n_63),
.Y(n_14)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_15),
.A2(n_16),
.B1(n_147),
.B2(n_149),
.Y(n_146)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_16),
.Y(n_15)
);

OAI22xp5_ASAP7_75t_SL g16 ( 
.A1(n_17),
.A2(n_18),
.B1(n_40),
.B2(n_53),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_18),
.Y(n_17)
);

AOI22xp5_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_20),
.B1(n_27),
.B2(n_39),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_20),
.Y(n_19)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_20),
.B(n_27),
.C(n_40),
.Y(n_96)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_21),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_21),
.B(n_83),
.Y(n_82)
);

AO22x1_ASAP7_75t_SL g21 ( 
.A1(n_22),
.A2(n_23),
.B1(n_25),
.B2(n_26),
.Y(n_21)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_22),
.Y(n_26)
);

INVx3_ASAP7_75t_SL g25 ( 
.A(n_23),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_L g44 ( 
.A1(n_23),
.A2(n_25),
.B1(n_45),
.B2(n_46),
.Y(n_44)
);

CKINVDCx6p67_ASAP7_75t_R g23 ( 
.A(n_24),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_25),
.B(n_66),
.Y(n_65)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_27),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_SL g122 ( 
.A(n_27),
.B(n_123),
.Y(n_122)
);

AOI21xp5_ASAP7_75t_L g27 ( 
.A1(n_28),
.A2(n_32),
.B(n_34),
.Y(n_27)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_28),
.A2(n_69),
.B1(n_103),
.B2(n_104),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_29),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_29),
.B(n_36),
.Y(n_35)
);

OA22x2_ASAP7_75t_L g60 ( 
.A1(n_29),
.A2(n_31),
.B1(n_58),
.B2(n_59),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_29),
.B(n_124),
.Y(n_123)
);

INVx3_ASAP7_75t_SL g32 ( 
.A(n_33),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_33),
.B(n_35),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_35),
.B(n_37),
.Y(n_34)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_35),
.Y(n_103)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_37),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_39),
.B(n_113),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_39),
.B(n_113),
.Y(n_128)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g40 ( 
.A1(n_41),
.A2(n_43),
.B1(n_51),
.B2(n_52),
.Y(n_40)
);

INVxp67_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

OAI21xp5_ASAP7_75t_L g86 ( 
.A1(n_42),
.A2(n_47),
.B(n_87),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_43),
.B(n_52),
.Y(n_87)
);

AND2x2_ASAP7_75t_L g43 ( 
.A(n_44),
.B(n_47),
.Y(n_43)
);

INVx5_ASAP7_75t_L g46 ( 
.A(n_45),
.Y(n_46)
);

OA22x2_ASAP7_75t_SL g47 ( 
.A1(n_45),
.A2(n_46),
.B1(n_48),
.B2(n_50),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_47),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_48),
.Y(n_50)
);

OAI22xp33_ASAP7_75t_L g57 ( 
.A1(n_48),
.A2(n_50),
.B1(n_58),
.B2(n_59),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_48),
.B(n_118),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_54),
.A2(n_134),
.B1(n_135),
.B2(n_136),
.Y(n_133)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_54),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_54),
.B(n_102),
.C(n_134),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_54),
.A2(n_63),
.B1(n_135),
.B2(n_148),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g54 ( 
.A1(n_55),
.A2(n_56),
.B1(n_61),
.B2(n_62),
.Y(n_54)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_55),
.Y(n_115)
);

INVxp67_ASAP7_75t_L g90 ( 
.A(n_56),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_56),
.B(n_62),
.Y(n_116)
);

AND2x2_ASAP7_75t_L g56 ( 
.A(n_57),
.B(n_60),
.Y(n_56)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_58),
.Y(n_59)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_60),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_60),
.B(n_90),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_L g114 ( 
.A1(n_60),
.A2(n_115),
.B(n_116),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_62),
.B(n_89),
.Y(n_88)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_63),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_64),
.B(n_67),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_64),
.A2(n_65),
.B1(n_67),
.B2(n_68),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_65),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_68),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_69),
.B(n_70),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_72),
.A2(n_73),
.B1(n_94),
.B2(n_95),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_74),
.A2(n_84),
.B1(n_85),
.B2(n_93),
.Y(n_73)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_74),
.Y(n_93)
);

OAI21xp5_ASAP7_75t_L g74 ( 
.A1(n_75),
.A2(n_76),
.B(n_79),
.Y(n_74)
);

INVx6_ASAP7_75t_L g78 ( 
.A(n_77),
.Y(n_78)
);

INVx8_ASAP7_75t_L g81 ( 
.A(n_77),
.Y(n_81)
);

INVx8_ASAP7_75t_L g99 ( 
.A(n_77),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_80),
.B(n_82),
.Y(n_79)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_86),
.A2(n_88),
.B1(n_91),
.B2(n_92),
.Y(n_85)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_86),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_86),
.A2(n_91),
.B1(n_114),
.B2(n_119),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_86),
.B(n_114),
.C(n_142),
.Y(n_145)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_88),
.Y(n_92)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

XOR2xp5_ASAP7_75t_L g95 ( 
.A(n_96),
.B(n_97),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_98),
.A2(n_101),
.B1(n_102),
.B2(n_106),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_98),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_100),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_101),
.A2(n_102),
.B1(n_132),
.B2(n_133),
.Y(n_131)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_102),
.B(n_126),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_102),
.B(n_126),
.Y(n_127)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

AOI21xp5_ASAP7_75t_L g108 ( 
.A1(n_109),
.A2(n_144),
.B(n_150),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_SL g109 ( 
.A1(n_110),
.A2(n_138),
.B(n_143),
.Y(n_109)
);

AOI21xp5_ASAP7_75t_L g110 ( 
.A1(n_111),
.A2(n_129),
.B(n_137),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_SL g111 ( 
.A1(n_112),
.A2(n_121),
.B(n_128),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_114),
.A2(n_117),
.B1(n_119),
.B2(n_120),
.Y(n_113)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_114),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_114),
.B(n_120),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_117),
.Y(n_120)
);

AOI21xp5_ASAP7_75t_L g121 ( 
.A1(n_122),
.A2(n_125),
.B(n_127),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_131),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_SL g137 ( 
.A(n_130),
.B(n_131),
.Y(n_137)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_134),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_140),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_139),
.B(n_140),
.Y(n_143)
);

XOR2xp5_ASAP7_75t_L g140 ( 
.A(n_141),
.B(n_142),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_146),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_SL g150 ( 
.A(n_145),
.B(n_146),
.Y(n_150)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_147),
.Y(n_149)
);


endmodule