module fake_jpeg_20091_n_107 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_107);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_107;

wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_106;
wire n_44;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_100;
wire n_82;
wire n_96;

INVx1_ASAP7_75t_L g35 ( 
.A(n_28),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_9),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_10),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_31),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_6),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_32),
.Y(n_40)
);

BUFx5_ASAP7_75t_L g41 ( 
.A(n_25),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_19),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_27),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_24),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_23),
.Y(n_45)
);

BUFx5_ASAP7_75t_L g46 ( 
.A(n_13),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_7),
.Y(n_47)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_30),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_21),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_37),
.B(n_0),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_50),
.B(n_53),
.Y(n_59)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_48),
.Y(n_51)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_51),
.Y(n_60)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_41),
.Y(n_52)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_52),
.Y(n_63)
);

BUFx4f_ASAP7_75t_SL g53 ( 
.A(n_41),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_46),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_54),
.Y(n_67)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_48),
.Y(n_55)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_55),
.Y(n_61)
);

INVx6_ASAP7_75t_SL g56 ( 
.A(n_46),
.Y(n_56)
);

INVx2_ASAP7_75t_SL g58 ( 
.A(n_56),
.Y(n_58)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_51),
.Y(n_57)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_57),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_56),
.A2(n_38),
.B1(n_39),
.B2(n_47),
.Y(n_62)
);

CKINVDCx14_ASAP7_75t_R g74 ( 
.A(n_62),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_L g64 ( 
.A1(n_55),
.A2(n_49),
.B1(n_42),
.B2(n_43),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_64),
.B(n_65),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_L g65 ( 
.A1(n_52),
.A2(n_40),
.B1(n_36),
.B2(n_35),
.Y(n_65)
);

BUFx12f_ASAP7_75t_L g66 ( 
.A(n_51),
.Y(n_66)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_66),
.Y(n_72)
);

A2O1A1Ixp33_ASAP7_75t_L g68 ( 
.A1(n_59),
.A2(n_0),
.B(n_1),
.C(n_2),
.Y(n_68)
);

AOI21xp5_ASAP7_75t_SL g88 ( 
.A1(n_68),
.A2(n_71),
.B(n_3),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_59),
.B(n_44),
.Y(n_69)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_69),
.Y(n_81)
);

AOI21xp5_ASAP7_75t_L g71 ( 
.A1(n_63),
.A2(n_45),
.B(n_17),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_67),
.B(n_16),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_73),
.B(n_78),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g75 ( 
.A(n_66),
.B(n_18),
.C(n_33),
.Y(n_75)
);

AND2x2_ASAP7_75t_L g87 ( 
.A(n_75),
.B(n_22),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_60),
.B(n_1),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_76),
.B(n_77),
.Y(n_85)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_61),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_58),
.B(n_15),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_64),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_79),
.Y(n_82)
);

INVxp67_ASAP7_75t_L g83 ( 
.A(n_78),
.Y(n_83)
);

INVx1_ASAP7_75t_SL g90 ( 
.A(n_83),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_80),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_84),
.A2(n_73),
.B1(n_86),
.B2(n_85),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_87),
.B(n_88),
.Y(n_91)
);

AND2x2_ASAP7_75t_L g89 ( 
.A(n_74),
.B(n_5),
.Y(n_89)
);

INVxp67_ASAP7_75t_L g93 ( 
.A(n_89),
.Y(n_93)
);

OAI21xp5_ASAP7_75t_SL g96 ( 
.A1(n_92),
.A2(n_94),
.B(n_90),
.Y(n_96)
);

INVxp67_ASAP7_75t_L g94 ( 
.A(n_86),
.Y(n_94)
);

XNOR2xp5_ASAP7_75t_SL g95 ( 
.A(n_91),
.B(n_82),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_95),
.B(n_96),
.C(n_81),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_93),
.Y(n_97)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_97),
.Y(n_99)
);

HB1xp67_ASAP7_75t_L g100 ( 
.A(n_98),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_100),
.A2(n_99),
.B1(n_70),
.B2(n_72),
.Y(n_101)
);

XNOR2xp5_ASAP7_75t_L g102 ( 
.A(n_101),
.B(n_8),
.Y(n_102)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_102),
.Y(n_103)
);

XOR2xp5_ASAP7_75t_L g104 ( 
.A(n_103),
.B(n_11),
.Y(n_104)
);

OAI21xp5_ASAP7_75t_L g105 ( 
.A1(n_104),
.A2(n_12),
.B(n_14),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_L g106 ( 
.A1(n_105),
.A2(n_34),
.B1(n_26),
.B2(n_29),
.Y(n_106)
);

XNOR2xp5_ASAP7_75t_L g107 ( 
.A(n_106),
.B(n_20),
.Y(n_107)
);


endmodule