module fake_jpeg_23664_n_304 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_304);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_304;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_182;
wire n_19;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_228;
wire n_178;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_288;
wire n_272;
wire n_284;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_301;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_298;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_145;
wire n_20;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_303;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_240;
wire n_212;
wire n_294;
wire n_299;
wire n_211;
wire n_300;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_302;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_297;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_4),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_11),
.Y(n_14)
);

INVx4_ASAP7_75t_L g15 ( 
.A(n_10),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

INVx8_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

INVx8_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

CKINVDCx16_ASAP7_75t_R g21 ( 
.A(n_9),
.Y(n_21)
);

CKINVDCx16_ASAP7_75t_R g22 ( 
.A(n_7),
.Y(n_22)
);

INVx8_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

INVx3_ASAP7_75t_R g24 ( 
.A(n_1),
.Y(n_24)
);

INVx11_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_11),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_19),
.Y(n_28)
);

INVx11_ASAP7_75t_L g38 ( 
.A(n_28),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_24),
.Y(n_29)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_29),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_27),
.B(n_12),
.Y(n_30)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_30),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_26),
.Y(n_31)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_31),
.Y(n_50)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_25),
.Y(n_32)
);

HB1xp67_ASAP7_75t_L g48 ( 
.A(n_32),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_24),
.Y(n_33)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_33),
.Y(n_41)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_19),
.Y(n_34)
);

INVx4_ASAP7_75t_SL g44 ( 
.A(n_34),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_24),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_35),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_24),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_36),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_24),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_37),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_31),
.Y(n_40)
);

INVx5_ASAP7_75t_L g60 ( 
.A(n_40),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_L g47 ( 
.A1(n_28),
.A2(n_19),
.B1(n_15),
.B2(n_23),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_47),
.A2(n_25),
.B1(n_15),
.B2(n_23),
.Y(n_71)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_32),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_49),
.B(n_14),
.Y(n_78)
);

INVxp67_ASAP7_75t_L g51 ( 
.A(n_29),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_51),
.B(n_53),
.Y(n_59)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_34),
.Y(n_52)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_52),
.Y(n_58)
);

CKINVDCx16_ASAP7_75t_R g53 ( 
.A(n_29),
.Y(n_53)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_33),
.Y(n_54)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_54),
.Y(n_62)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_33),
.Y(n_55)
);

INVx5_ASAP7_75t_L g66 ( 
.A(n_55),
.Y(n_66)
);

INVx2_ASAP7_75t_SL g56 ( 
.A(n_35),
.Y(n_56)
);

CKINVDCx16_ASAP7_75t_R g74 ( 
.A(n_56),
.Y(n_74)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_42),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_57),
.B(n_61),
.Y(n_80)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_42),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_44),
.A2(n_19),
.B1(n_15),
.B2(n_25),
.Y(n_63)
);

OAI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_63),
.A2(n_72),
.B1(n_23),
.B2(n_18),
.Y(n_96)
);

INVxp67_ASAP7_75t_L g64 ( 
.A(n_48),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_64),
.B(n_67),
.Y(n_81)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_38),
.Y(n_65)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_65),
.Y(n_86)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_52),
.Y(n_67)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_42),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_68),
.B(n_69),
.Y(n_92)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_50),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_40),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_70),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_71),
.A2(n_49),
.B1(n_41),
.B2(n_23),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_44),
.A2(n_15),
.B1(n_25),
.B2(n_21),
.Y(n_72)
);

BUFx3_ASAP7_75t_L g73 ( 
.A(n_50),
.Y(n_73)
);

INVx8_ASAP7_75t_L g94 ( 
.A(n_73),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_46),
.Y(n_75)
);

BUFx2_ASAP7_75t_L g98 ( 
.A(n_75),
.Y(n_98)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_38),
.Y(n_76)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_76),
.Y(n_91)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_44),
.Y(n_77)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_77),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_78),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g79 ( 
.A(n_59),
.B(n_39),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_79),
.B(n_82),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_SL g82 ( 
.A(n_69),
.B(n_39),
.Y(n_82)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_66),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_83),
.B(n_84),
.Y(n_111)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_73),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g85 ( 
.A(n_74),
.B(n_24),
.Y(n_85)
);

OAI21xp5_ASAP7_75t_SL g105 ( 
.A1(n_85),
.A2(n_87),
.B(n_101),
.Y(n_105)
);

AND2x2_ASAP7_75t_L g87 ( 
.A(n_57),
.B(n_24),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_88),
.A2(n_95),
.B1(n_77),
.B2(n_76),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_64),
.B(n_51),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_89),
.B(n_93),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_58),
.B(n_53),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_66),
.A2(n_55),
.B1(n_41),
.B2(n_56),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_L g119 ( 
.A1(n_96),
.A2(n_18),
.B1(n_60),
.B2(n_22),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_58),
.B(n_17),
.C(n_26),
.Y(n_99)
);

XNOR2xp5_ASAP7_75t_L g107 ( 
.A(n_99),
.B(n_17),
.Y(n_107)
);

OAI21xp5_ASAP7_75t_SL g101 ( 
.A1(n_62),
.A2(n_17),
.B(n_26),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_88),
.A2(n_54),
.B1(n_68),
.B2(n_61),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_103),
.A2(n_118),
.B1(n_123),
.B2(n_92),
.Y(n_130)
);

INVx5_ASAP7_75t_L g104 ( 
.A(n_83),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_104),
.B(n_106),
.Y(n_136)
);

INVx13_ASAP7_75t_L g106 ( 
.A(n_83),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_107),
.B(n_109),
.C(n_112),
.Y(n_137)
);

INVx13_ASAP7_75t_L g108 ( 
.A(n_84),
.Y(n_108)
);

INVxp67_ASAP7_75t_L g140 ( 
.A(n_108),
.Y(n_140)
);

NAND2xp33_ASAP7_75t_SL g109 ( 
.A(n_101),
.B(n_17),
.Y(n_109)
);

OAI21xp33_ASAP7_75t_L g110 ( 
.A1(n_97),
.A2(n_17),
.B(n_10),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_110),
.B(n_114),
.Y(n_132)
);

NOR2xp67_ASAP7_75t_SL g112 ( 
.A(n_96),
.B(n_17),
.Y(n_112)
);

HB1xp67_ASAP7_75t_L g113 ( 
.A(n_98),
.Y(n_113)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_113),
.Y(n_126)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_80),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_L g127 ( 
.A1(n_115),
.A2(n_112),
.B1(n_87),
.B2(n_104),
.Y(n_127)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_80),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_116),
.B(n_87),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_95),
.A2(n_65),
.B1(n_18),
.B2(n_17),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_119),
.A2(n_89),
.B1(n_92),
.B2(n_91),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_90),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_120),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_97),
.B(n_45),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_121),
.B(n_123),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_L g122 ( 
.A(n_99),
.B(n_37),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_122),
.B(n_100),
.C(n_86),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_93),
.B(n_43),
.Y(n_123)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_94),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_124),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_94),
.B(n_60),
.Y(n_125)
);

INVxp67_ASAP7_75t_L g144 ( 
.A(n_125),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_127),
.A2(n_94),
.B1(n_106),
.B2(n_108),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_128),
.A2(n_130),
.B1(n_133),
.B2(n_142),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_117),
.B(n_82),
.Y(n_131)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_131),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_105),
.A2(n_109),
.B1(n_117),
.B2(n_116),
.Y(n_133)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_135),
.Y(n_161)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_111),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_138),
.B(n_139),
.Y(n_151)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_121),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_105),
.A2(n_87),
.B1(n_85),
.B2(n_81),
.Y(n_142)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_103),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_143),
.B(n_149),
.Y(n_164)
);

XOR2xp5_ASAP7_75t_L g170 ( 
.A(n_145),
.B(n_150),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_114),
.A2(n_85),
.B1(n_81),
.B2(n_100),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_146),
.A2(n_130),
.B1(n_128),
.B2(n_143),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_102),
.B(n_122),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_147),
.B(n_148),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_107),
.B(n_85),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_SL g149 ( 
.A(n_120),
.B(n_79),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_115),
.B(n_91),
.C(n_86),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_134),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_154),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_155),
.A2(n_145),
.B1(n_138),
.B2(n_126),
.Y(n_199)
);

AND2x6_ASAP7_75t_L g156 ( 
.A(n_133),
.B(n_124),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_SL g177 ( 
.A1(n_156),
.A2(n_158),
.B(n_160),
.Y(n_177)
);

INVxp67_ASAP7_75t_L g157 ( 
.A(n_136),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_157),
.B(n_166),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_SL g158 ( 
.A1(n_142),
.A2(n_118),
.B(n_90),
.Y(n_158)
);

AND2x2_ASAP7_75t_L g160 ( 
.A(n_146),
.B(n_106),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_162),
.A2(n_176),
.B1(n_150),
.B2(n_144),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_L g163 ( 
.A1(n_132),
.A2(n_14),
.B(n_16),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_SL g180 ( 
.A1(n_163),
.A2(n_165),
.B(n_168),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_SL g165 ( 
.A1(n_137),
.A2(n_108),
.B(n_16),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_134),
.B(n_98),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_131),
.B(n_46),
.Y(n_167)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_167),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_136),
.B(n_98),
.Y(n_168)
);

INVxp67_ASAP7_75t_L g169 ( 
.A(n_127),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_169),
.B(n_162),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_141),
.B(n_56),
.Y(n_171)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_171),
.Y(n_188)
);

INVx13_ASAP7_75t_L g172 ( 
.A(n_140),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_SL g197 ( 
.A1(n_172),
.A2(n_173),
.B1(n_153),
.B2(n_21),
.Y(n_197)
);

AOI21xp5_ASAP7_75t_L g173 ( 
.A1(n_137),
.A2(n_16),
.B(n_13),
.Y(n_173)
);

AND2x2_ASAP7_75t_L g174 ( 
.A(n_129),
.B(n_0),
.Y(n_174)
);

AND2x2_ASAP7_75t_L g192 ( 
.A(n_174),
.B(n_175),
.Y(n_192)
);

AND2x2_ASAP7_75t_L g175 ( 
.A(n_129),
.B(n_0),
.Y(n_175)
);

OAI32xp33_ASAP7_75t_L g176 ( 
.A1(n_148),
.A2(n_14),
.A3(n_36),
.B1(n_35),
.B2(n_20),
.Y(n_176)
);

OA21x2_ASAP7_75t_SL g179 ( 
.A1(n_165),
.A2(n_132),
.B(n_147),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_SL g206 ( 
.A(n_179),
.B(n_173),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_L g204 ( 
.A1(n_181),
.A2(n_197),
.B1(n_198),
.B2(n_201),
.Y(n_204)
);

BUFx6f_ASAP7_75t_L g182 ( 
.A(n_172),
.Y(n_182)
);

BUFx2_ASAP7_75t_L g213 ( 
.A(n_182),
.Y(n_213)
);

CKINVDCx16_ASAP7_75t_R g183 ( 
.A(n_168),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_183),
.B(n_191),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_154),
.B(n_141),
.Y(n_184)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_184),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_172),
.B(n_126),
.Y(n_185)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_185),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_SL g189 ( 
.A(n_164),
.B(n_149),
.Y(n_189)
);

CKINVDCx14_ASAP7_75t_R g209 ( 
.A(n_189),
.Y(n_209)
);

INVxp67_ASAP7_75t_L g190 ( 
.A(n_171),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_190),
.B(n_193),
.Y(n_222)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_151),
.Y(n_191)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_151),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_167),
.Y(n_194)
);

OAI22xp33_ASAP7_75t_SL g212 ( 
.A1(n_194),
.A2(n_196),
.B1(n_199),
.B2(n_200),
.Y(n_212)
);

AOI21xp5_ASAP7_75t_SL g195 ( 
.A1(n_164),
.A2(n_139),
.B(n_135),
.Y(n_195)
);

AOI21xp5_ASAP7_75t_SL g218 ( 
.A1(n_195),
.A2(n_163),
.B(n_160),
.Y(n_218)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_174),
.Y(n_196)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_174),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_156),
.A2(n_18),
.B1(n_27),
.B2(n_13),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_199),
.B(n_170),
.C(n_159),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_202),
.B(n_211),
.C(n_214),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g203 ( 
.A(n_177),
.B(n_170),
.Y(n_203)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_203),
.B(n_205),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_SL g205 ( 
.A(n_198),
.B(n_152),
.Y(n_205)
);

CKINVDCx14_ASAP7_75t_R g238 ( 
.A(n_206),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_SL g207 ( 
.A(n_177),
.B(n_152),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_SL g234 ( 
.A(n_207),
.B(n_219),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_186),
.B(n_159),
.C(n_161),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g214 ( 
.A(n_180),
.B(n_155),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_180),
.B(n_158),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_215),
.B(n_192),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_L g216 ( 
.A1(n_201),
.A2(n_153),
.B1(n_161),
.B2(n_160),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_216),
.A2(n_221),
.B1(n_176),
.B2(n_27),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_187),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_217),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_218),
.A2(n_200),
.B1(n_196),
.B2(n_194),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_SL g219 ( 
.A(n_195),
.B(n_192),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_L g221 ( 
.A1(n_191),
.A2(n_193),
.B1(n_187),
.B2(n_189),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_202),
.B(n_203),
.C(n_211),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_224),
.B(n_228),
.C(n_231),
.Y(n_244)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_222),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_225),
.B(n_46),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_226),
.A2(n_230),
.B1(n_239),
.B2(n_22),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_227),
.B(n_240),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_207),
.B(n_186),
.C(n_178),
.Y(n_228)
);

HB1xp67_ASAP7_75t_L g229 ( 
.A(n_213),
.Y(n_229)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_229),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_209),
.A2(n_190),
.B1(n_188),
.B2(n_192),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_222),
.B(n_188),
.C(n_175),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_214),
.B(n_175),
.C(n_182),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_232),
.B(n_236),
.C(n_241),
.Y(n_248)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_235),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_219),
.B(n_75),
.C(n_45),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_204),
.A2(n_208),
.B1(n_210),
.B2(n_220),
.Y(n_237)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_237),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_205),
.A2(n_13),
.B1(n_22),
.B2(n_21),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_212),
.B(n_45),
.C(n_43),
.Y(n_241)
);

AOI221xp5_ASAP7_75t_L g242 ( 
.A1(n_234),
.A2(n_215),
.B1(n_218),
.B2(n_213),
.C(n_11),
.Y(n_242)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_242),
.Y(n_269)
);

XOR2xp5_ASAP7_75t_L g267 ( 
.A(n_243),
.B(n_250),
.Y(n_267)
);

AOI21xp5_ASAP7_75t_L g245 ( 
.A1(n_228),
.A2(n_12),
.B(n_9),
.Y(n_245)
);

AOI21xp5_ASAP7_75t_L g261 ( 
.A1(n_245),
.A2(n_251),
.B(n_20),
.Y(n_261)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_246),
.Y(n_271)
);

INVx13_ASAP7_75t_L g249 ( 
.A(n_234),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_249),
.B(n_2),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_223),
.B(n_20),
.Y(n_250)
);

FAx1_ASAP7_75t_SL g253 ( 
.A(n_231),
.B(n_20),
.CI(n_36),
.CON(n_253),
.SN(n_253)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_253),
.B(n_256),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_240),
.B(n_9),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_254),
.B(n_0),
.C(n_1),
.Y(n_260)
);

HB1xp67_ASAP7_75t_L g256 ( 
.A(n_233),
.Y(n_256)
);

OAI21xp33_ASAP7_75t_L g257 ( 
.A1(n_232),
.A2(n_0),
.B(n_1),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_257),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_270)
);

AOI21xp5_ASAP7_75t_SL g258 ( 
.A1(n_255),
.A2(n_236),
.B(n_238),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_258),
.B(n_264),
.Y(n_273)
);

AOI31xp33_ASAP7_75t_L g259 ( 
.A1(n_257),
.A2(n_223),
.A3(n_241),
.B(n_224),
.Y(n_259)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_259),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_260),
.B(n_263),
.C(n_3),
.Y(n_279)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_261),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_244),
.B(n_43),
.C(n_2),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_262),
.B(n_244),
.C(n_247),
.Y(n_275)
);

AOI21xp5_ASAP7_75t_L g263 ( 
.A1(n_248),
.A2(n_1),
.B(n_2),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_248),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_265),
.B(n_270),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_252),
.B(n_3),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_266),
.B(n_254),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_272),
.B(n_280),
.Y(n_286)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_267),
.B(n_243),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_SL g288 ( 
.A(n_274),
.B(n_277),
.Y(n_288)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_275),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_268),
.B(n_253),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_267),
.B(n_250),
.C(n_249),
.Y(n_278)
);

OAI21xp5_ASAP7_75t_SL g287 ( 
.A1(n_278),
.A2(n_265),
.B(n_269),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_SL g283 ( 
.A(n_279),
.B(n_270),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_262),
.B(n_5),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_283),
.B(n_285),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_SL g285 ( 
.A(n_275),
.B(n_258),
.Y(n_285)
);

XOR2xp5_ASAP7_75t_L g291 ( 
.A(n_287),
.B(n_278),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_282),
.B(n_273),
.Y(n_289)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_289),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_SL g290 ( 
.A(n_276),
.B(n_271),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_290),
.B(n_286),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_291),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_289),
.A2(n_281),
.B1(n_274),
.B2(n_260),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_293),
.B(n_295),
.Y(n_298)
);

HB1xp67_ASAP7_75t_L g297 ( 
.A(n_291),
.Y(n_297)
);

AOI322xp5_ASAP7_75t_L g299 ( 
.A1(n_297),
.A2(n_288),
.A3(n_294),
.B1(n_292),
.B2(n_284),
.C1(n_6),
.C2(n_8),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_299),
.B(n_298),
.C(n_296),
.Y(n_300)
);

NAND3xp33_ASAP7_75t_L g301 ( 
.A(n_300),
.B(n_6),
.C(n_7),
.Y(n_301)
);

AOI21xp5_ASAP7_75t_SL g302 ( 
.A1(n_301),
.A2(n_6),
.B(n_8),
.Y(n_302)
);

XOR2xp5_ASAP7_75t_L g303 ( 
.A(n_302),
.B(n_8),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_L g304 ( 
.A(n_303),
.B(n_8),
.Y(n_304)
);


endmodule