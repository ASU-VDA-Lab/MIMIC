module fake_jpeg_11188_n_43 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_43);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;

output n_43;

wire n_13;
wire n_21;
wire n_33;
wire n_10;
wire n_23;
wire n_27;
wire n_22;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

CKINVDCx20_ASAP7_75t_R g7 ( 
.A(n_3),
.Y(n_7)
);

INVx1_ASAP7_75t_L g8 ( 
.A(n_5),
.Y(n_8)
);

BUFx12f_ASAP7_75t_L g9 ( 
.A(n_5),
.Y(n_9)
);

INVx4_ASAP7_75t_L g10 ( 
.A(n_2),
.Y(n_10)
);

BUFx3_ASAP7_75t_L g11 ( 
.A(n_6),
.Y(n_11)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_2),
.Y(n_12)
);

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_0),
.Y(n_13)
);

INVx2_ASAP7_75t_L g14 ( 
.A(n_0),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_13),
.Y(n_15)
);

INVx5_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

INVx1_ASAP7_75t_SL g16 ( 
.A(n_9),
.Y(n_16)
);

OR2x2_ASAP7_75t_L g27 ( 
.A(n_16),
.B(n_17),
.Y(n_27)
);

INVx6_ASAP7_75t_SL g17 ( 
.A(n_9),
.Y(n_17)
);

INVx6_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_18),
.Y(n_26)
);

INVx11_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

AOI22xp33_ASAP7_75t_L g20 ( 
.A1(n_14),
.A2(n_1),
.B1(n_6),
.B2(n_4),
.Y(n_20)
);

OAI22xp5_ASAP7_75t_SL g22 ( 
.A1(n_20),
.A2(n_11),
.B1(n_8),
.B2(n_12),
.Y(n_22)
);

INVx5_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

AOI21xp5_ASAP7_75t_L g25 ( 
.A1(n_21),
.A2(n_1),
.B(n_4),
.Y(n_25)
);

AOI22xp5_ASAP7_75t_L g24 ( 
.A1(n_18),
.A2(n_11),
.B1(n_7),
.B2(n_1),
.Y(n_24)
);

AOI21xp5_ASAP7_75t_L g29 ( 
.A1(n_24),
.A2(n_25),
.B(n_19),
.Y(n_29)
);

CKINVDCx16_ASAP7_75t_R g28 ( 
.A(n_27),
.Y(n_28)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_28),
.Y(n_32)
);

AOI22xp33_ASAP7_75t_L g31 ( 
.A1(n_29),
.A2(n_22),
.B1(n_19),
.B2(n_18),
.Y(n_31)
);

HB1xp67_ASAP7_75t_L g30 ( 
.A(n_29),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_30),
.B(n_21),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_31),
.B(n_23),
.Y(n_35)
);

AND2x2_ASAP7_75t_SL g33 ( 
.A(n_32),
.B(n_24),
.Y(n_33)
);

OAI21xp5_ASAP7_75t_SL g36 ( 
.A1(n_33),
.A2(n_35),
.B(n_30),
.Y(n_36)
);

OR2x2_ASAP7_75t_L g37 ( 
.A(n_34),
.B(n_23),
.Y(n_37)
);

AOI21xp5_ASAP7_75t_L g40 ( 
.A1(n_36),
.A2(n_26),
.B(n_15),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_SL g41 ( 
.A1(n_37),
.A2(n_26),
.B1(n_38),
.B2(n_32),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_SL g38 ( 
.A(n_33),
.B(n_15),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_38),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_40),
.B(n_41),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_42),
.B(n_39),
.Y(n_43)
);


endmodule