module fake_jpeg_5646_n_206 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_206);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_206;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_9),
.Y(n_15)
);

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_12),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_7),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_13),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_3),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_6),
.Y(n_25)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

BUFx16f_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_6),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_5),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_18),
.B(n_24),
.Y(n_31)
);

AND2x2_ASAP7_75t_L g53 ( 
.A(n_31),
.B(n_37),
.Y(n_53)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_19),
.Y(n_32)
);

INVx11_ASAP7_75t_L g47 ( 
.A(n_32),
.Y(n_47)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_19),
.Y(n_33)
);

INVx11_ASAP7_75t_L g55 ( 
.A(n_33),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_15),
.B(n_0),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_34),
.B(n_21),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_16),
.Y(n_35)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_35),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_27),
.Y(n_36)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_36),
.Y(n_60)
);

AND2x2_ASAP7_75t_SL g37 ( 
.A(n_27),
.B(n_0),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_27),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_38),
.B(n_39),
.Y(n_44)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_27),
.Y(n_39)
);

INVx5_ASAP7_75t_L g40 ( 
.A(n_19),
.Y(n_40)
);

HB1xp67_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_16),
.Y(n_41)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_41),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_31),
.B(n_18),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_42),
.B(n_51),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g43 ( 
.A1(n_37),
.A2(n_26),
.B1(n_28),
.B2(n_33),
.Y(n_43)
);

INVxp67_ASAP7_75t_L g74 ( 
.A(n_43),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_37),
.B(n_18),
.Y(n_46)
);

OAI21xp33_ASAP7_75t_L g62 ( 
.A1(n_46),
.A2(n_56),
.B(n_58),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_36),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_49),
.Y(n_77)
);

OA22x2_ASAP7_75t_L g50 ( 
.A1(n_40),
.A2(n_28),
.B1(n_26),
.B2(n_16),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_50),
.A2(n_55),
.B1(n_46),
.B2(n_41),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_38),
.B(n_24),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_52),
.B(n_21),
.Y(n_71)
);

OR2x2_ASAP7_75t_SL g56 ( 
.A(n_36),
.B(n_22),
.Y(n_56)
);

NAND2xp33_ASAP7_75t_SL g57 ( 
.A(n_32),
.B(n_30),
.Y(n_57)
);

A2O1A1Ixp33_ASAP7_75t_L g66 ( 
.A1(n_57),
.A2(n_25),
.B(n_20),
.C(n_30),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_35),
.B(n_17),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_33),
.B(n_17),
.Y(n_59)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_59),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_54),
.B(n_26),
.Y(n_63)
);

CKINVDCx14_ASAP7_75t_R g97 ( 
.A(n_63),
.Y(n_97)
);

INVx5_ASAP7_75t_L g64 ( 
.A(n_50),
.Y(n_64)
);

INVxp67_ASAP7_75t_L g91 ( 
.A(n_64),
.Y(n_91)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_50),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_65),
.B(n_78),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_66),
.B(n_70),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_51),
.B(n_23),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_67),
.B(n_68),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_47),
.B(n_23),
.Y(n_68)
);

MAJx2_ASAP7_75t_L g69 ( 
.A(n_53),
.B(n_57),
.C(n_50),
.Y(n_69)
);

XOR2xp5_ASAP7_75t_L g89 ( 
.A(n_69),
.B(n_59),
.Y(n_89)
);

CKINVDCx16_ASAP7_75t_R g70 ( 
.A(n_44),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_71),
.B(n_79),
.Y(n_90)
);

INVx5_ASAP7_75t_L g72 ( 
.A(n_50),
.Y(n_72)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_72),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_42),
.B(n_28),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_75),
.B(n_48),
.Y(n_80)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_76),
.B(n_16),
.Y(n_100)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_47),
.Y(n_78)
);

CKINVDCx16_ASAP7_75t_R g79 ( 
.A(n_44),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_80),
.B(n_84),
.Y(n_119)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_78),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_81),
.B(n_82),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_65),
.A2(n_55),
.B1(n_60),
.B2(n_47),
.Y(n_82)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_77),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_83),
.B(n_85),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_75),
.B(n_61),
.Y(n_84)
);

OR2x2_ASAP7_75t_L g85 ( 
.A(n_64),
.B(n_53),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_74),
.A2(n_55),
.B1(n_48),
.B2(n_53),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_86),
.A2(n_93),
.B1(n_94),
.B2(n_100),
.Y(n_115)
);

XNOR2xp5_ASAP7_75t_SL g103 ( 
.A(n_89),
.B(n_99),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_74),
.A2(n_56),
.B1(n_60),
.B2(n_49),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_72),
.A2(n_60),
.B1(n_58),
.B2(n_39),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_66),
.B(n_73),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_95),
.B(n_98),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_73),
.B(n_52),
.Y(n_98)
);

AND2x2_ASAP7_75t_SL g99 ( 
.A(n_69),
.B(n_36),
.Y(n_99)
);

INVx13_ASAP7_75t_L g102 ( 
.A(n_99),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_102),
.B(n_105),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_80),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_104),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_99),
.A2(n_76),
.B1(n_61),
.B2(n_77),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_83),
.B(n_79),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_SL g133 ( 
.A(n_107),
.B(n_112),
.Y(n_133)
);

AND2x6_ASAP7_75t_L g108 ( 
.A(n_99),
.B(n_62),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_108),
.B(n_93),
.C(n_90),
.Y(n_128)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_84),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_109),
.B(n_110),
.Y(n_134)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_92),
.Y(n_110)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_94),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_111),
.B(n_113),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_97),
.B(n_70),
.Y(n_112)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_87),
.Y(n_113)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_87),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_116),
.B(n_118),
.Y(n_135)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_81),
.Y(n_117)
);

INVxp33_ASAP7_75t_L g121 ( 
.A(n_117),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_95),
.B(n_45),
.Y(n_118)
);

AND2x2_ASAP7_75t_L g120 ( 
.A(n_105),
.B(n_89),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_L g152 ( 
.A1(n_120),
.A2(n_127),
.B(n_98),
.Y(n_152)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_117),
.Y(n_123)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_123),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_119),
.B(n_109),
.Y(n_125)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_125),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_119),
.B(n_86),
.Y(n_126)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_126),
.Y(n_144)
);

NAND2x1_ASAP7_75t_SL g127 ( 
.A(n_108),
.B(n_85),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_SL g145 ( 
.A1(n_128),
.A2(n_102),
.B(n_116),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_104),
.B(n_100),
.Y(n_130)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_130),
.Y(n_146)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_106),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_131),
.B(n_132),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_114),
.Y(n_132)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_101),
.Y(n_136)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_136),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_103),
.B(n_85),
.C(n_100),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_137),
.B(n_103),
.C(n_113),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_L g161 ( 
.A(n_139),
.B(n_148),
.Y(n_161)
);

XOR2xp5_ASAP7_75t_L g140 ( 
.A(n_127),
.B(n_115),
.Y(n_140)
);

XOR2xp5_ASAP7_75t_L g158 ( 
.A(n_140),
.B(n_142),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_L g142 ( 
.A(n_127),
.B(n_115),
.Y(n_142)
);

AOI21xp5_ASAP7_75t_L g159 ( 
.A1(n_145),
.A2(n_130),
.B(n_126),
.Y(n_159)
);

CKINVDCx16_ASAP7_75t_R g147 ( 
.A(n_134),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_147),
.B(n_151),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_137),
.B(n_111),
.C(n_110),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_128),
.B(n_90),
.C(n_45),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_L g164 ( 
.A(n_149),
.B(n_152),
.Y(n_164)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_125),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_L g153 ( 
.A(n_122),
.B(n_88),
.Y(n_153)
);

BUFx24_ASAP7_75t_SL g160 ( 
.A(n_153),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_138),
.B(n_124),
.Y(n_155)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_155),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_146),
.A2(n_124),
.B1(n_129),
.B2(n_131),
.Y(n_156)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_156),
.Y(n_168)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_149),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_157),
.B(n_165),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_L g169 ( 
.A1(n_159),
.A2(n_139),
.B(n_141),
.Y(n_169)
);

OAI22xp33_ASAP7_75t_L g162 ( 
.A1(n_142),
.A2(n_135),
.B1(n_132),
.B2(n_91),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_162),
.A2(n_150),
.B1(n_152),
.B2(n_153),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_144),
.A2(n_136),
.B1(n_120),
.B2(n_133),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_163),
.B(n_120),
.Y(n_172)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_140),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_148),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_166),
.B(n_96),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_169),
.B(n_173),
.C(n_174),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_170),
.B(n_161),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_SL g181 ( 
.A(n_172),
.B(n_170),
.Y(n_181)
);

XOR2xp5_ASAP7_75t_L g173 ( 
.A(n_158),
.B(n_88),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_158),
.B(n_143),
.C(n_121),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_175),
.B(n_176),
.C(n_177),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_L g176 ( 
.A1(n_154),
.A2(n_22),
.B(n_15),
.Y(n_176)
);

MAJx2_ASAP7_75t_L g177 ( 
.A(n_164),
.B(n_16),
.C(n_123),
.Y(n_177)
);

O2A1O1Ixp33_ASAP7_75t_L g178 ( 
.A1(n_171),
.A2(n_162),
.B(n_164),
.C(n_161),
.Y(n_178)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_178),
.Y(n_188)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_175),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_180),
.B(n_1),
.Y(n_192)
);

O2A1O1Ixp33_ASAP7_75t_SL g193 ( 
.A1(n_181),
.A2(n_182),
.B(n_186),
.C(n_10),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_167),
.B(n_143),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_184),
.B(n_1),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_173),
.B(n_160),
.C(n_29),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_185),
.B(n_14),
.C(n_12),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g186 ( 
.A1(n_168),
.A2(n_25),
.B1(n_20),
.B2(n_29),
.Y(n_186)
);

AO21x1_ASAP7_75t_L g187 ( 
.A1(n_178),
.A2(n_177),
.B(n_14),
.Y(n_187)
);

BUFx24_ASAP7_75t_SL g194 ( 
.A(n_187),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_189),
.B(n_190),
.Y(n_195)
);

NOR3xp33_ASAP7_75t_L g191 ( 
.A(n_183),
.B(n_11),
.C(n_10),
.Y(n_191)
);

AO21x1_ASAP7_75t_L g197 ( 
.A1(n_191),
.A2(n_11),
.B(n_3),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_192),
.B(n_184),
.C(n_179),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_193),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_198)
);

FAx1_ASAP7_75t_SL g199 ( 
.A(n_196),
.B(n_189),
.CI(n_188),
.CON(n_199),
.SN(n_199)
);

AO21x1_ASAP7_75t_SL g202 ( 
.A1(n_197),
.A2(n_8),
.B(n_2),
.Y(n_202)
);

INVxp67_ASAP7_75t_L g200 ( 
.A(n_198),
.Y(n_200)
);

AND2x2_ASAP7_75t_L g204 ( 
.A(n_199),
.B(n_201),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_L g201 ( 
.A1(n_195),
.A2(n_194),
.B(n_4),
.Y(n_201)
);

OAI311xp33_ASAP7_75t_L g203 ( 
.A1(n_202),
.A2(n_2),
.A3(n_5),
.B1(n_8),
.C1(n_200),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_203),
.B(n_5),
.C(n_8),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_L g206 ( 
.A(n_205),
.B(n_204),
.Y(n_206)
);


endmodule