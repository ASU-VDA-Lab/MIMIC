module fake_jpeg_7913_n_204 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_204);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_204;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_4),
.Y(n_14)
);

INVx11_ASAP7_75t_L g15 ( 
.A(n_1),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_3),
.Y(n_16)
);

BUFx3_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_9),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_10),
.Y(n_24)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_11),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_4),
.Y(n_28)
);

INVx11_ASAP7_75t_L g29 ( 
.A(n_15),
.Y(n_29)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_29),
.Y(n_47)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_17),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_30),
.B(n_34),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_17),
.Y(n_31)
);

INVx5_ASAP7_75t_L g51 ( 
.A(n_31),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_32),
.Y(n_44)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_23),
.Y(n_33)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_33),
.Y(n_49)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_17),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_15),
.Y(n_35)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_35),
.Y(n_40)
);

INVx11_ASAP7_75t_L g36 ( 
.A(n_23),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_36),
.B(n_37),
.Y(n_41)
);

INVx11_ASAP7_75t_L g37 ( 
.A(n_23),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_22),
.Y(n_38)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_38),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_L g42 ( 
.A1(n_33),
.A2(n_19),
.B1(n_25),
.B2(n_20),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_L g75 ( 
.A1(n_42),
.A2(n_37),
.B1(n_30),
.B2(n_26),
.Y(n_75)
);

BUFx12_ASAP7_75t_L g45 ( 
.A(n_38),
.Y(n_45)
);

CKINVDCx14_ASAP7_75t_R g70 ( 
.A(n_45),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_34),
.B(n_27),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_SL g67 ( 
.A(n_46),
.B(n_53),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_33),
.A2(n_14),
.B1(n_16),
.B2(n_28),
.Y(n_48)
);

AOI21xp5_ASAP7_75t_L g76 ( 
.A1(n_48),
.A2(n_50),
.B(n_26),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_33),
.A2(n_14),
.B1(n_16),
.B2(n_28),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_33),
.A2(n_19),
.B1(n_25),
.B2(n_18),
.Y(n_52)
);

OAI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_52),
.A2(n_54),
.B1(n_36),
.B2(n_37),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_SL g53 ( 
.A(n_30),
.B(n_27),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_36),
.A2(n_20),
.B1(n_18),
.B2(n_21),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_32),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_55),
.B(n_29),
.Y(n_60)
);

AOI32xp33_ASAP7_75t_L g56 ( 
.A1(n_49),
.A2(n_31),
.A3(n_38),
.B1(n_29),
.B2(n_32),
.Y(n_56)
);

A2O1A1Ixp33_ASAP7_75t_L g84 ( 
.A1(n_56),
.A2(n_58),
.B(n_76),
.C(n_42),
.Y(n_84)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_51),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_57),
.B(n_61),
.Y(n_79)
);

AND2x4_ASAP7_75t_L g58 ( 
.A(n_47),
.B(n_29),
.Y(n_58)
);

INVx5_ASAP7_75t_L g59 ( 
.A(n_51),
.Y(n_59)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_59),
.Y(n_85)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_60),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_53),
.B(n_21),
.Y(n_61)
);

OAI22xp33_ASAP7_75t_L g93 ( 
.A1(n_62),
.A2(n_63),
.B1(n_75),
.B2(n_44),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_51),
.A2(n_36),
.B1(n_37),
.B2(n_24),
.Y(n_63)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_47),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_64),
.B(n_66),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_39),
.B(n_35),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_65),
.B(n_55),
.Y(n_81)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_41),
.Y(n_66)
);

INVxp67_ASAP7_75t_L g68 ( 
.A(n_39),
.Y(n_68)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_68),
.Y(n_80)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_41),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_69),
.B(n_71),
.Y(n_97)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_45),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_48),
.B(n_24),
.Y(n_72)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_72),
.Y(n_89)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_46),
.Y(n_73)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_73),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_50),
.B(n_22),
.Y(n_74)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_74),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_60),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_77),
.B(n_64),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_81),
.B(n_83),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_68),
.B(n_43),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_84),
.A2(n_93),
.B1(n_49),
.B2(n_44),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_65),
.B(n_43),
.Y(n_86)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_86),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_72),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_87),
.B(n_92),
.Y(n_110)
);

NOR2x1_ASAP7_75t_L g88 ( 
.A(n_58),
.B(n_56),
.Y(n_88)
);

NOR2x1_ASAP7_75t_L g107 ( 
.A(n_88),
.B(n_76),
.Y(n_107)
);

AND2x2_ASAP7_75t_SL g92 ( 
.A(n_58),
.B(n_40),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_66),
.B(n_34),
.Y(n_94)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_94),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_67),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_95),
.B(n_99),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_69),
.B(n_34),
.Y(n_96)
);

XOR2xp5_ASAP7_75t_L g112 ( 
.A(n_96),
.B(n_98),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_73),
.B(n_34),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_58),
.B(n_40),
.C(n_38),
.Y(n_99)
);

AOI21xp5_ASAP7_75t_L g101 ( 
.A1(n_88),
.A2(n_58),
.B(n_59),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_SL g133 ( 
.A1(n_101),
.A2(n_90),
.B(n_34),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_82),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_103),
.B(n_104),
.Y(n_128)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_97),
.Y(n_104)
);

INVxp67_ASAP7_75t_L g106 ( 
.A(n_79),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_106),
.B(n_109),
.Y(n_132)
);

AO21x1_ASAP7_75t_L g134 ( 
.A1(n_107),
.A2(n_31),
.B(n_22),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_108),
.A2(n_93),
.B1(n_80),
.B2(n_86),
.Y(n_126)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_85),
.Y(n_109)
);

AND2x6_ASAP7_75t_L g111 ( 
.A(n_92),
.B(n_67),
.Y(n_111)
);

A2O1A1O1Ixp25_ASAP7_75t_L g131 ( 
.A1(n_111),
.A2(n_90),
.B(n_96),
.C(n_22),
.D(n_31),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_84),
.A2(n_49),
.B1(n_44),
.B2(n_70),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_113),
.A2(n_116),
.B1(n_99),
.B2(n_83),
.Y(n_122)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_114),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_91),
.A2(n_71),
.B1(n_32),
.B2(n_35),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_85),
.B(n_45),
.Y(n_117)
);

INVxp67_ASAP7_75t_L g125 ( 
.A(n_117),
.Y(n_125)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_98),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_118),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_78),
.B(n_45),
.Y(n_119)
);

INVxp33_ASAP7_75t_L g135 ( 
.A(n_119),
.Y(n_135)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_94),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_SL g123 ( 
.A1(n_120),
.A2(n_78),
.B(n_81),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_122),
.A2(n_126),
.B1(n_130),
.B2(n_102),
.Y(n_148)
);

AOI21xp5_ASAP7_75t_L g140 ( 
.A1(n_123),
.A2(n_133),
.B(n_137),
.Y(n_140)
);

AO22x1_ASAP7_75t_L g124 ( 
.A1(n_107),
.A2(n_92),
.B1(n_113),
.B2(n_101),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_124),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_110),
.A2(n_91),
.B1(n_87),
.B2(n_89),
.Y(n_129)
);

INVxp67_ASAP7_75t_L g155 ( 
.A(n_129),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_115),
.A2(n_89),
.B1(n_80),
.B2(n_95),
.Y(n_130)
);

XNOR2xp5_ASAP7_75t_L g141 ( 
.A(n_131),
.B(n_100),
.Y(n_141)
);

AOI222xp33_ASAP7_75t_L g151 ( 
.A1(n_134),
.A2(n_26),
.B1(n_106),
.B2(n_111),
.C1(n_34),
.C2(n_35),
.Y(n_151)
);

INVx3_ASAP7_75t_L g136 ( 
.A(n_109),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_136),
.B(n_138),
.Y(n_147)
);

AOI21xp5_ASAP7_75t_L g137 ( 
.A1(n_120),
.A2(n_57),
.B(n_38),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_116),
.Y(n_138)
);

XOR2xp5_ASAP7_75t_L g139 ( 
.A(n_112),
.B(n_34),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_139),
.B(n_105),
.C(n_112),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_141),
.B(n_145),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_SL g142 ( 
.A(n_128),
.B(n_102),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_142),
.B(n_143),
.Y(n_167)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_132),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_SL g144 ( 
.A(n_122),
.B(n_100),
.Y(n_144)
);

XOR2xp5_ASAP7_75t_L g163 ( 
.A(n_144),
.B(n_134),
.Y(n_163)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_137),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_146),
.B(n_139),
.C(n_133),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_148),
.A2(n_151),
.B1(n_152),
.B2(n_129),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_SL g149 ( 
.A(n_121),
.B(n_105),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_SL g160 ( 
.A(n_149),
.B(n_135),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_130),
.A2(n_118),
.B1(n_35),
.B2(n_32),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_136),
.B(n_135),
.Y(n_153)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_153),
.Y(n_159)
);

OAI32xp33_ASAP7_75t_L g154 ( 
.A1(n_124),
.A2(n_0),
.A3(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_154)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_154),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_156),
.B(n_165),
.C(n_140),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_158),
.A2(n_162),
.B1(n_155),
.B2(n_1),
.Y(n_176)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_160),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_150),
.A2(n_131),
.B1(n_127),
.B2(n_124),
.Y(n_162)
);

XOR2xp5_ASAP7_75t_L g173 ( 
.A(n_163),
.B(n_151),
.Y(n_173)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_147),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_SL g169 ( 
.A1(n_164),
.A2(n_166),
.B(n_159),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_146),
.B(n_125),
.C(n_8),
.Y(n_165)
);

INVxp67_ASAP7_75t_L g166 ( 
.A(n_152),
.Y(n_166)
);

OR2x2_ASAP7_75t_L g184 ( 
.A(n_169),
.B(n_2),
.Y(n_184)
);

FAx1_ASAP7_75t_SL g170 ( 
.A(n_156),
.B(n_144),
.CI(n_148),
.CON(n_170),
.SN(n_170)
);

OAI31xp33_ASAP7_75t_L g180 ( 
.A1(n_170),
.A2(n_158),
.A3(n_166),
.B(n_9),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_L g171 ( 
.A(n_165),
.B(n_141),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_L g182 ( 
.A(n_171),
.B(n_175),
.Y(n_182)
);

XOR2xp5_ASAP7_75t_L g179 ( 
.A(n_172),
.B(n_173),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_163),
.B(n_155),
.C(n_125),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g185 ( 
.A(n_174),
.B(n_177),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g175 ( 
.A(n_157),
.B(n_154),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_176),
.B(n_0),
.Y(n_183)
);

XOR2xp5_ASAP7_75t_L g177 ( 
.A(n_162),
.B(n_8),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_SL g178 ( 
.A1(n_168),
.A2(n_161),
.B(n_167),
.Y(n_178)
);

AOI21xp5_ASAP7_75t_L g192 ( 
.A1(n_178),
.A2(n_180),
.B(n_13),
.Y(n_192)
);

INVxp67_ASAP7_75t_SL g181 ( 
.A(n_174),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_181),
.B(n_183),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_184),
.B(n_2),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_181),
.A2(n_172),
.B1(n_177),
.B2(n_170),
.Y(n_187)
);

INVxp67_ASAP7_75t_L g194 ( 
.A(n_187),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_188),
.B(n_189),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_184),
.B(n_182),
.Y(n_189)
);

AND2x2_ASAP7_75t_L g190 ( 
.A(n_185),
.B(n_173),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_190),
.B(n_191),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_179),
.B(n_11),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_SL g197 ( 
.A1(n_192),
.A2(n_12),
.B(n_13),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_SL g193 ( 
.A(n_186),
.B(n_12),
.Y(n_193)
);

NOR3xp33_ASAP7_75t_L g198 ( 
.A(n_193),
.B(n_186),
.C(n_6),
.Y(n_198)
);

AOI21xp5_ASAP7_75t_L g199 ( 
.A1(n_197),
.A2(n_190),
.B(n_6),
.Y(n_199)
);

AOI21xp5_ASAP7_75t_L g203 ( 
.A1(n_198),
.A2(n_200),
.B(n_6),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_199),
.B(n_201),
.C(n_195),
.Y(n_202)
);

INVxp67_ASAP7_75t_L g200 ( 
.A(n_196),
.Y(n_200)
);

AOI21xp5_ASAP7_75t_L g201 ( 
.A1(n_194),
.A2(n_7),
.B(n_5),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_202),
.B(n_203),
.Y(n_204)
);


endmodule