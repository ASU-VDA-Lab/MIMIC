module fake_jpeg_2847_n_690 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_690);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_690;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_657;
wire n_27;
wire n_664;
wire n_365;
wire n_179;
wire n_620;
wire n_686;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_678;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_417;
wire n_362;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_635;
wire n_517;
wire n_629;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_643;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_647;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_641;
wire n_48;
wire n_465;
wire n_638;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_623;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_637;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_672;
wire n_309;
wire n_624;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_606;
wire n_496;
wire n_166;
wire n_688;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_646;
wire n_319;
wire n_689;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_663;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_393;
wire n_349;
wire n_234;
wire n_530;
wire n_634;
wire n_23;
wire n_69;
wire n_658;
wire n_195;
wire n_450;
wire n_557;
wire n_681;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_666;
wire n_639;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_645;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_622;
wire n_463;
wire n_667;
wire n_92;
wire n_332;
wire n_640;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_653;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_626;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_668;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_682;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_642;
wire n_101;
wire n_226;
wire n_509;
wire n_644;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_656;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_649;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_679;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_615;
wire n_598;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_662;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_676;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_648;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_670;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_683;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_631;
wire n_433;
wire n_636;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_650;
wire n_218;
wire n_63;
wire n_652;
wire n_599;
wire n_239;
wire n_674;
wire n_243;
wire n_481;
wire n_628;
wire n_619;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_419;
wire n_378;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_655;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_684;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_680;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_625;
wire n_147;
wire n_449;
wire n_627;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_659;
wire n_125;
wire n_661;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_687;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_673;
wire n_58;
wire n_41;
wire n_613;
wire n_630;
wire n_266;
wire n_548;
wire n_665;
wire n_72;
wire n_512;
wire n_654;
wire n_445;
wire n_443;
wire n_677;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_671;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_669;
wire n_524;
wire n_402;
wire n_563;
wire n_685;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_660;
wire n_373;
wire n_633;
wire n_112;
wire n_632;
wire n_616;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_651;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_675;
wire n_335;
wire n_120;
wire n_621;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx8_ASAP7_75t_L g20 ( 
.A(n_15),
.Y(n_20)
);

INVx6_ASAP7_75t_SL g21 ( 
.A(n_0),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_12),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_17),
.Y(n_23)
);

BUFx10_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_0),
.Y(n_25)
);

INVx11_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_12),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_16),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_12),
.Y(n_34)
);

INVx11_ASAP7_75t_SL g35 ( 
.A(n_17),
.Y(n_35)
);

BUFx16f_ASAP7_75t_L g36 ( 
.A(n_8),
.Y(n_36)
);

HB1xp67_ASAP7_75t_L g37 ( 
.A(n_17),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_14),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_2),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_10),
.Y(n_40)
);

BUFx4f_ASAP7_75t_SL g41 ( 
.A(n_2),
.Y(n_41)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_3),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_3),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_16),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_18),
.Y(n_45)
);

INVxp67_ASAP7_75t_L g46 ( 
.A(n_2),
.Y(n_46)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_9),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_1),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_13),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_13),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_6),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_7),
.Y(n_52)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_4),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_17),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_5),
.Y(n_55)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_11),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_9),
.Y(n_57)
);

AND2x2_ASAP7_75t_SL g58 ( 
.A(n_33),
.B(n_9),
.Y(n_58)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_58),
.B(n_39),
.C(n_52),
.Y(n_177)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_23),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g166 ( 
.A(n_59),
.Y(n_166)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_34),
.Y(n_60)
);

INVx4_ASAP7_75t_SL g151 ( 
.A(n_60),
.Y(n_151)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_33),
.Y(n_61)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_61),
.Y(n_134)
);

AND2x2_ASAP7_75t_L g62 ( 
.A(n_33),
.B(n_9),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_62),
.B(n_74),
.Y(n_149)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_21),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g192 ( 
.A(n_63),
.Y(n_192)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_21),
.Y(n_64)
);

INVx5_ASAP7_75t_L g144 ( 
.A(n_64),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_46),
.B(n_8),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_65),
.B(n_96),
.Y(n_195)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_47),
.Y(n_66)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_66),
.Y(n_138)
);

BUFx12f_ASAP7_75t_L g67 ( 
.A(n_21),
.Y(n_67)
);

INVx5_ASAP7_75t_L g145 ( 
.A(n_67),
.Y(n_145)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_47),
.Y(n_68)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_68),
.Y(n_154)
);

BUFx12_ASAP7_75t_L g69 ( 
.A(n_36),
.Y(n_69)
);

BUFx12f_ASAP7_75t_L g136 ( 
.A(n_69),
.Y(n_136)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_30),
.Y(n_70)
);

INVx3_ASAP7_75t_L g140 ( 
.A(n_70),
.Y(n_140)
);

BUFx12f_ASAP7_75t_L g71 ( 
.A(n_35),
.Y(n_71)
);

INVx5_ASAP7_75t_L g147 ( 
.A(n_71),
.Y(n_147)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_34),
.Y(n_72)
);

INVx3_ASAP7_75t_L g158 ( 
.A(n_72),
.Y(n_158)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_23),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g168 ( 
.A(n_73),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_SL g74 ( 
.A(n_22),
.B(n_8),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_23),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g172 ( 
.A(n_75),
.Y(n_172)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_34),
.Y(n_76)
);

INVx3_ASAP7_75t_L g167 ( 
.A(n_76),
.Y(n_167)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_47),
.Y(n_77)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_77),
.Y(n_137)
);

BUFx12f_ASAP7_75t_L g78 ( 
.A(n_35),
.Y(n_78)
);

INVx5_ASAP7_75t_L g150 ( 
.A(n_78),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_23),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g205 ( 
.A(n_79),
.Y(n_205)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_45),
.Y(n_80)
);

INVx3_ASAP7_75t_L g190 ( 
.A(n_80),
.Y(n_190)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_32),
.Y(n_81)
);

INVx6_ASAP7_75t_L g143 ( 
.A(n_81),
.Y(n_143)
);

BUFx12f_ASAP7_75t_L g82 ( 
.A(n_36),
.Y(n_82)
);

INVx5_ASAP7_75t_L g189 ( 
.A(n_82),
.Y(n_189)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_32),
.Y(n_83)
);

INVx6_ASAP7_75t_L g155 ( 
.A(n_83),
.Y(n_155)
);

BUFx5_ASAP7_75t_L g84 ( 
.A(n_36),
.Y(n_84)
);

INVx4_ASAP7_75t_L g183 ( 
.A(n_84),
.Y(n_183)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_30),
.Y(n_85)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_85),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_32),
.Y(n_86)
);

INVx6_ASAP7_75t_L g165 ( 
.A(n_86),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_32),
.Y(n_87)
);

INVx8_ASAP7_75t_L g139 ( 
.A(n_87),
.Y(n_139)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_30),
.Y(n_88)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_88),
.Y(n_170)
);

CKINVDCx16_ASAP7_75t_R g89 ( 
.A(n_41),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_89),
.B(n_121),
.Y(n_152)
);

INVx5_ASAP7_75t_L g90 ( 
.A(n_20),
.Y(n_90)
);

BUFx3_ASAP7_75t_L g194 ( 
.A(n_90),
.Y(n_194)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_44),
.Y(n_91)
);

BUFx12f_ASAP7_75t_L g146 ( 
.A(n_91),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_44),
.Y(n_92)
);

BUFx12f_ASAP7_75t_L g153 ( 
.A(n_92),
.Y(n_153)
);

INVx11_ASAP7_75t_L g93 ( 
.A(n_43),
.Y(n_93)
);

INVx11_ASAP7_75t_L g133 ( 
.A(n_93),
.Y(n_133)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_56),
.Y(n_94)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_94),
.Y(n_174)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_45),
.Y(n_95)
);

INVx3_ASAP7_75t_L g193 ( 
.A(n_95),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_27),
.B(n_10),
.Y(n_96)
);

INVx11_ASAP7_75t_L g97 ( 
.A(n_43),
.Y(n_97)
);

INVx4_ASAP7_75t_L g142 ( 
.A(n_97),
.Y(n_142)
);

BUFx5_ASAP7_75t_L g98 ( 
.A(n_36),
.Y(n_98)
);

INVx4_ASAP7_75t_L g188 ( 
.A(n_98),
.Y(n_188)
);

INVx8_ASAP7_75t_L g99 ( 
.A(n_43),
.Y(n_99)
);

INVx5_ASAP7_75t_L g208 ( 
.A(n_99),
.Y(n_208)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_27),
.Y(n_100)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_100),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_44),
.Y(n_101)
);

BUFx12f_ASAP7_75t_L g169 ( 
.A(n_101),
.Y(n_169)
);

INVx11_ASAP7_75t_L g102 ( 
.A(n_43),
.Y(n_102)
);

INVx4_ASAP7_75t_L g157 ( 
.A(n_102),
.Y(n_157)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_45),
.Y(n_103)
);

INVx3_ASAP7_75t_L g198 ( 
.A(n_103),
.Y(n_198)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_29),
.Y(n_104)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_104),
.Y(n_175)
);

BUFx12f_ASAP7_75t_L g105 ( 
.A(n_36),
.Y(n_105)
);

INVx4_ASAP7_75t_L g197 ( 
.A(n_105),
.Y(n_197)
);

INVx5_ASAP7_75t_L g106 ( 
.A(n_20),
.Y(n_106)
);

INVx4_ASAP7_75t_L g200 ( 
.A(n_106),
.Y(n_200)
);

BUFx3_ASAP7_75t_L g107 ( 
.A(n_20),
.Y(n_107)
);

INVx4_ASAP7_75t_L g206 ( 
.A(n_107),
.Y(n_206)
);

BUFx3_ASAP7_75t_L g108 ( 
.A(n_56),
.Y(n_108)
);

INVx4_ASAP7_75t_L g207 ( 
.A(n_108),
.Y(n_207)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_44),
.Y(n_109)
);

BUFx12f_ASAP7_75t_L g201 ( 
.A(n_109),
.Y(n_201)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_49),
.Y(n_110)
);

INVx4_ASAP7_75t_L g164 ( 
.A(n_110),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_49),
.Y(n_111)
);

INVx4_ASAP7_75t_L g178 ( 
.A(n_111),
.Y(n_178)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_43),
.Y(n_112)
);

INVx3_ASAP7_75t_L g199 ( 
.A(n_112),
.Y(n_199)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_56),
.Y(n_113)
);

INVx3_ASAP7_75t_L g227 ( 
.A(n_113),
.Y(n_227)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_40),
.Y(n_114)
);

HB1xp67_ASAP7_75t_L g228 ( 
.A(n_114),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_29),
.B(n_10),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_115),
.B(n_124),
.Y(n_221)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_40),
.Y(n_116)
);

INVx4_ASAP7_75t_L g216 ( 
.A(n_116),
.Y(n_216)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_49),
.Y(n_117)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_117),
.Y(n_180)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_49),
.Y(n_118)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_118),
.Y(n_184)
);

INVx6_ASAP7_75t_L g119 ( 
.A(n_31),
.Y(n_119)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_119),
.Y(n_186)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_50),
.Y(n_120)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_120),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_SL g121 ( 
.A(n_22),
.B(n_10),
.Y(n_121)
);

INVx8_ASAP7_75t_L g122 ( 
.A(n_40),
.Y(n_122)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_122),
.Y(n_203)
);

BUFx3_ASAP7_75t_L g123 ( 
.A(n_31),
.Y(n_123)
);

INVx1_ASAP7_75t_SL g212 ( 
.A(n_123),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_50),
.B(n_19),
.Y(n_124)
);

INVx4_ASAP7_75t_L g125 ( 
.A(n_40),
.Y(n_125)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_125),
.Y(n_210)
);

INVx13_ASAP7_75t_L g126 ( 
.A(n_41),
.Y(n_126)
);

INVx13_ASAP7_75t_L g202 ( 
.A(n_126),
.Y(n_202)
);

HB1xp67_ASAP7_75t_L g127 ( 
.A(n_40),
.Y(n_127)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_127),
.Y(n_217)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_31),
.Y(n_128)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_128),
.Y(n_220)
);

BUFx12f_ASAP7_75t_SL g129 ( 
.A(n_24),
.Y(n_129)
);

INVx6_ASAP7_75t_SL g231 ( 
.A(n_129),
.Y(n_231)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_31),
.Y(n_130)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_130),
.Y(n_222)
);

INVx11_ASAP7_75t_L g131 ( 
.A(n_41),
.Y(n_131)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_131),
.Y(n_234)
);

INVx13_ASAP7_75t_L g132 ( 
.A(n_41),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_132),
.Y(n_156)
);

AOI22xp33_ASAP7_75t_SL g135 ( 
.A1(n_131),
.A2(n_37),
.B1(n_26),
.B2(n_25),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g252 ( 
.A1(n_135),
.A2(n_159),
.B1(n_160),
.B2(n_163),
.Y(n_252)
);

OA22x2_ASAP7_75t_L g148 ( 
.A1(n_58),
.A2(n_37),
.B1(n_42),
.B2(n_53),
.Y(n_148)
);

AND2x2_ASAP7_75t_L g259 ( 
.A(n_148),
.B(n_177),
.Y(n_259)
);

AOI22xp33_ASAP7_75t_L g159 ( 
.A1(n_128),
.A2(n_41),
.B1(n_26),
.B2(n_25),
.Y(n_159)
);

AOI22xp33_ASAP7_75t_L g160 ( 
.A1(n_130),
.A2(n_83),
.B1(n_81),
.B2(n_79),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_64),
.B(n_57),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_SL g285 ( 
.A(n_162),
.B(n_171),
.Y(n_285)
);

AOI22xp33_ASAP7_75t_SL g163 ( 
.A1(n_63),
.A2(n_26),
.B1(n_54),
.B2(n_55),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_64),
.B(n_57),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_62),
.A2(n_54),
.B1(n_28),
.B2(n_38),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_173),
.A2(n_179),
.B1(n_187),
.B2(n_204),
.Y(n_236)
);

OAI22xp33_ASAP7_75t_SL g179 ( 
.A1(n_59),
.A2(n_28),
.B1(n_38),
.B2(n_52),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_67),
.B(n_55),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_181),
.B(n_182),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_67),
.B(n_51),
.Y(n_182)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_127),
.Y(n_185)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_185),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_73),
.A2(n_53),
.B1(n_42),
.B2(n_48),
.Y(n_187)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_70),
.Y(n_191)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_191),
.Y(n_267)
);

AOI22xp33_ASAP7_75t_SL g196 ( 
.A1(n_71),
.A2(n_51),
.B1(n_48),
.B2(n_39),
.Y(n_196)
);

AOI22xp33_ASAP7_75t_SL g248 ( 
.A1(n_196),
.A2(n_209),
.B1(n_78),
.B2(n_102),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_75),
.A2(n_53),
.B1(n_42),
.B2(n_24),
.Y(n_204)
);

AOI22xp33_ASAP7_75t_SL g209 ( 
.A1(n_71),
.A2(n_24),
.B1(n_11),
.B2(n_13),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_82),
.B(n_19),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_211),
.B(n_214),
.Y(n_282)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_125),
.Y(n_213)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_213),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_82),
.B(n_19),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_108),
.Y(n_215)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_215),
.Y(n_286)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_119),
.Y(n_218)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_218),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_105),
.B(n_19),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_219),
.B(n_233),
.Y(n_260)
);

AO22x1_ASAP7_75t_SL g223 ( 
.A1(n_105),
.A2(n_24),
.B1(n_18),
.B2(n_16),
.Y(n_223)
);

AND2x2_ASAP7_75t_L g288 ( 
.A(n_223),
.B(n_3),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_86),
.B(n_18),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_SL g243 ( 
.A(n_224),
.B(n_230),
.Y(n_243)
);

AOI22xp33_ASAP7_75t_L g225 ( 
.A1(n_87),
.A2(n_24),
.B1(n_1),
.B2(n_2),
.Y(n_225)
);

OAI22xp33_ASAP7_75t_SL g272 ( 
.A1(n_225),
.A2(n_226),
.B1(n_232),
.B2(n_118),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_90),
.A2(n_24),
.B1(n_18),
.B2(n_16),
.Y(n_226)
);

AND2x2_ASAP7_75t_L g229 ( 
.A(n_99),
.B(n_14),
.Y(n_229)
);

OAI21xp33_ASAP7_75t_L g276 ( 
.A1(n_229),
.A2(n_3),
.B(n_4),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_107),
.B(n_15),
.Y(n_230)
);

AOI22xp33_ASAP7_75t_L g232 ( 
.A1(n_91),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_78),
.B(n_15),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_L g235 ( 
.A1(n_92),
.A2(n_15),
.B1(n_14),
.B2(n_11),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_235),
.A2(n_179),
.B1(n_229),
.B2(n_176),
.Y(n_269)
);

INVxp67_ASAP7_75t_L g237 ( 
.A(n_231),
.Y(n_237)
);

INVxp67_ASAP7_75t_L g338 ( 
.A(n_237),
.Y(n_338)
);

INVx5_ASAP7_75t_L g238 ( 
.A(n_147),
.Y(n_238)
);

INVx4_ASAP7_75t_L g362 ( 
.A(n_238),
.Y(n_362)
);

BUFx3_ASAP7_75t_L g239 ( 
.A(n_150),
.Y(n_239)
);

INVx4_ASAP7_75t_L g383 ( 
.A(n_239),
.Y(n_383)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_186),
.Y(n_240)
);

INVx2_ASAP7_75t_L g330 ( 
.A(n_240),
.Y(n_330)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_217),
.Y(n_241)
);

INVx2_ASAP7_75t_L g332 ( 
.A(n_241),
.Y(n_332)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_220),
.Y(n_242)
);

INVx2_ASAP7_75t_L g357 ( 
.A(n_242),
.Y(n_357)
);

INVx4_ASAP7_75t_L g245 ( 
.A(n_234),
.Y(n_245)
);

INVx3_ASAP7_75t_L g349 ( 
.A(n_245),
.Y(n_349)
);

INVx5_ASAP7_75t_L g246 ( 
.A(n_189),
.Y(n_246)
);

INVx3_ASAP7_75t_L g389 ( 
.A(n_246),
.Y(n_389)
);

INVx11_ASAP7_75t_L g247 ( 
.A(n_146),
.Y(n_247)
);

INVx5_ASAP7_75t_SL g371 ( 
.A(n_247),
.Y(n_371)
);

INVxp67_ASAP7_75t_L g347 ( 
.A(n_248),
.Y(n_347)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_222),
.Y(n_249)
);

INVx2_ASAP7_75t_L g364 ( 
.A(n_249),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_SL g250 ( 
.A(n_221),
.B(n_123),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_SL g360 ( 
.A(n_250),
.B(n_258),
.Y(n_360)
);

INVx8_ASAP7_75t_L g251 ( 
.A(n_136),
.Y(n_251)
);

INVx2_ASAP7_75t_L g372 ( 
.A(n_251),
.Y(n_372)
);

INVx3_ASAP7_75t_L g253 ( 
.A(n_208),
.Y(n_253)
);

INVx2_ASAP7_75t_SL g370 ( 
.A(n_253),
.Y(n_370)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_180),
.Y(n_254)
);

INVx2_ASAP7_75t_L g385 ( 
.A(n_254),
.Y(n_385)
);

INVxp67_ASAP7_75t_L g255 ( 
.A(n_228),
.Y(n_255)
);

INVxp67_ASAP7_75t_L g359 ( 
.A(n_255),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_152),
.B(n_0),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_256),
.B(n_264),
.Y(n_331)
);

INVx5_ASAP7_75t_L g257 ( 
.A(n_136),
.Y(n_257)
);

BUFx6f_ASAP7_75t_L g345 ( 
.A(n_257),
.Y(n_345)
);

CKINVDCx16_ASAP7_75t_R g258 ( 
.A(n_202),
.Y(n_258)
);

HB1xp67_ASAP7_75t_L g261 ( 
.A(n_190),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g336 ( 
.A(n_261),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_156),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g368 ( 
.A(n_262),
.Y(n_368)
);

AOI22xp33_ASAP7_75t_SL g263 ( 
.A1(n_137),
.A2(n_97),
.B1(n_93),
.B2(n_122),
.Y(n_263)
);

AOI22xp33_ASAP7_75t_SL g329 ( 
.A1(n_263),
.A2(n_291),
.B1(n_298),
.B2(n_302),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_141),
.B(n_1),
.Y(n_264)
);

BUFx6f_ASAP7_75t_L g266 ( 
.A(n_166),
.Y(n_266)
);

BUFx6f_ASAP7_75t_L g365 ( 
.A(n_266),
.Y(n_365)
);

AOI21xp5_ASAP7_75t_L g268 ( 
.A1(n_135),
.A2(n_132),
.B(n_126),
.Y(n_268)
);

AOI21xp5_ASAP7_75t_L g384 ( 
.A1(n_268),
.A2(n_301),
.B(n_237),
.Y(n_384)
);

OAI22xp5_ASAP7_75t_L g340 ( 
.A1(n_269),
.A2(n_225),
.B1(n_232),
.B2(n_209),
.Y(n_340)
);

CKINVDCx14_ASAP7_75t_R g270 ( 
.A(n_202),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_SL g377 ( 
.A(n_270),
.B(n_273),
.Y(n_377)
);

INVx1_ASAP7_75t_SL g271 ( 
.A(n_151),
.Y(n_271)
);

AND2x2_ASAP7_75t_L g355 ( 
.A(n_271),
.B(n_276),
.Y(n_355)
);

AOI22xp5_ASAP7_75t_SL g326 ( 
.A1(n_272),
.A2(n_288),
.B1(n_317),
.B2(n_322),
.Y(n_326)
);

CKINVDCx16_ASAP7_75t_R g273 ( 
.A(n_228),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_144),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_SL g378 ( 
.A(n_274),
.B(n_277),
.Y(n_378)
);

INVx6_ASAP7_75t_L g275 ( 
.A(n_166),
.Y(n_275)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_275),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_SL g277 ( 
.A(n_149),
.B(n_117),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_145),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_278),
.B(n_279),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_195),
.B(n_111),
.Y(n_279)
);

INVx13_ASAP7_75t_L g280 ( 
.A(n_136),
.Y(n_280)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_280),
.Y(n_328)
);

INVx4_ASAP7_75t_SL g281 ( 
.A(n_193),
.Y(n_281)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_281),
.Y(n_334)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_184),
.Y(n_284)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_284),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_175),
.B(n_3),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_289),
.B(n_293),
.Y(n_348)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_134),
.Y(n_290)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_290),
.Y(n_344)
);

INVx11_ASAP7_75t_L g291 ( 
.A(n_146),
.Y(n_291)
);

INVx3_ASAP7_75t_L g292 ( 
.A(n_197),
.Y(n_292)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_292),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_148),
.B(n_4),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_148),
.B(n_4),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_294),
.B(n_311),
.Y(n_354)
);

INVx3_ASAP7_75t_SL g295 ( 
.A(n_151),
.Y(n_295)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_295),
.Y(n_380)
);

INVx2_ASAP7_75t_L g296 ( 
.A(n_138),
.Y(n_296)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_296),
.Y(n_381)
);

INVx2_ASAP7_75t_L g297 ( 
.A(n_154),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g351 ( 
.A(n_297),
.B(n_299),
.Y(n_351)
);

AOI22xp33_ASAP7_75t_SL g298 ( 
.A1(n_198),
.A2(n_110),
.B1(n_109),
.B2(n_101),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g299 ( 
.A(n_168),
.Y(n_299)
);

INVx6_ASAP7_75t_L g300 ( 
.A(n_172),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g356 ( 
.A(n_300),
.B(n_303),
.Y(n_356)
);

AOI21xp5_ASAP7_75t_L g301 ( 
.A1(n_163),
.A2(n_69),
.B(n_14),
.Y(n_301)
);

INVx2_ASAP7_75t_SL g302 ( 
.A(n_194),
.Y(n_302)
);

INVx2_ASAP7_75t_L g303 ( 
.A(n_203),
.Y(n_303)
);

AOI22xp33_ASAP7_75t_SL g304 ( 
.A1(n_227),
.A2(n_158),
.B1(n_167),
.B2(n_200),
.Y(n_304)
);

AOI22xp33_ASAP7_75t_SL g343 ( 
.A1(n_304),
.A2(n_312),
.B1(n_313),
.B2(n_315),
.Y(n_343)
);

INVx4_ASAP7_75t_L g305 ( 
.A(n_133),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g358 ( 
.A(n_305),
.B(n_306),
.Y(n_358)
);

INVx2_ASAP7_75t_L g306 ( 
.A(n_168),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_161),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g363 ( 
.A(n_307),
.B(n_308),
.Y(n_363)
);

INVxp67_ASAP7_75t_L g308 ( 
.A(n_210),
.Y(n_308)
);

INVx2_ASAP7_75t_L g309 ( 
.A(n_143),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g367 ( 
.A(n_309),
.B(n_310),
.Y(n_367)
);

INVx5_ASAP7_75t_L g310 ( 
.A(n_192),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_223),
.B(n_5),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_143),
.Y(n_312)
);

INVx3_ASAP7_75t_L g313 ( 
.A(n_212),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_170),
.B(n_69),
.C(n_6),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_314),
.B(n_183),
.C(n_188),
.Y(n_337)
);

INVxp67_ASAP7_75t_L g315 ( 
.A(n_199),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_174),
.Y(n_316)
);

AOI22xp33_ASAP7_75t_SL g369 ( 
.A1(n_316),
.A2(n_318),
.B1(n_319),
.B2(n_321),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_192),
.B(n_5),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_140),
.Y(n_318)
);

INVx2_ASAP7_75t_L g319 ( 
.A(n_155),
.Y(n_319)
);

AOI22xp5_ASAP7_75t_SL g320 ( 
.A1(n_206),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_320)
);

NOR2x1_ASAP7_75t_L g350 ( 
.A(n_320),
.B(n_323),
.Y(n_350)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_155),
.Y(n_321)
);

INVx4_ASAP7_75t_L g322 ( 
.A(n_133),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g323 ( 
.A(n_165),
.Y(n_323)
);

INVxp67_ASAP7_75t_L g324 ( 
.A(n_196),
.Y(n_324)
);

AOI22xp5_ASAP7_75t_SL g388 ( 
.A1(n_324),
.A2(n_325),
.B1(n_271),
.B2(n_295),
.Y(n_388)
);

INVx2_ASAP7_75t_L g325 ( 
.A(n_165),
.Y(n_325)
);

AOI22xp33_ASAP7_75t_L g333 ( 
.A1(n_252),
.A2(n_159),
.B1(n_160),
.B2(n_164),
.Y(n_333)
);

OAI22xp5_ASAP7_75t_L g421 ( 
.A1(n_333),
.A2(n_342),
.B1(n_361),
.B2(n_382),
.Y(n_421)
);

MAJIxp5_ASAP7_75t_L g396 ( 
.A(n_337),
.B(n_387),
.C(n_315),
.Y(n_396)
);

AOI22xp5_ASAP7_75t_L g391 ( 
.A1(n_340),
.A2(n_346),
.B1(n_352),
.B2(n_353),
.Y(n_391)
);

OAI21xp5_ASAP7_75t_L g341 ( 
.A1(n_324),
.A2(n_216),
.B(n_194),
.Y(n_341)
);

OAI21xp5_ASAP7_75t_SL g416 ( 
.A1(n_341),
.A2(n_384),
.B(n_386),
.Y(n_416)
);

AOI22x1_ASAP7_75t_L g342 ( 
.A1(n_293),
.A2(n_139),
.B1(n_153),
.B2(n_201),
.Y(n_342)
);

OAI22xp5_ASAP7_75t_SL g346 ( 
.A1(n_294),
.A2(n_164),
.B1(n_178),
.B2(n_205),
.Y(n_346)
);

OAI22xp5_ASAP7_75t_SL g352 ( 
.A1(n_269),
.A2(n_178),
.B1(n_172),
.B2(n_205),
.Y(n_352)
);

OAI22xp5_ASAP7_75t_L g353 ( 
.A1(n_311),
.A2(n_236),
.B1(n_259),
.B2(n_288),
.Y(n_353)
);

AOI22xp5_ASAP7_75t_L g361 ( 
.A1(n_236),
.A2(n_139),
.B1(n_216),
.B2(n_207),
.Y(n_361)
);

AOI32xp33_ASAP7_75t_L g366 ( 
.A1(n_260),
.A2(n_157),
.A3(n_142),
.B1(n_201),
.B2(n_153),
.Y(n_366)
);

NOR2xp33_ASAP7_75t_L g398 ( 
.A(n_366),
.B(n_262),
.Y(n_398)
);

OAI22xp5_ASAP7_75t_L g373 ( 
.A1(n_259),
.A2(n_146),
.B1(n_169),
.B2(n_153),
.Y(n_373)
);

AOI22xp5_ASAP7_75t_L g394 ( 
.A1(n_373),
.A2(n_376),
.B1(n_379),
.B2(n_281),
.Y(n_394)
);

OAI22xp33_ASAP7_75t_SL g375 ( 
.A1(n_301),
.A2(n_142),
.B1(n_157),
.B2(n_169),
.Y(n_375)
);

AOI22xp33_ASAP7_75t_L g417 ( 
.A1(n_375),
.A2(n_247),
.B1(n_310),
.B2(n_257),
.Y(n_417)
);

OAI22xp5_ASAP7_75t_SL g376 ( 
.A1(n_259),
.A2(n_201),
.B1(n_169),
.B2(n_7),
.Y(n_376)
);

OAI22xp5_ASAP7_75t_SL g379 ( 
.A1(n_288),
.A2(n_7),
.B1(n_5),
.B2(n_6),
.Y(n_379)
);

AOI22xp33_ASAP7_75t_L g382 ( 
.A1(n_268),
.A2(n_6),
.B1(n_7),
.B2(n_289),
.Y(n_382)
);

OAI21xp5_ASAP7_75t_L g386 ( 
.A1(n_282),
.A2(n_256),
.B(n_264),
.Y(n_386)
);

MAJIxp5_ASAP7_75t_L g387 ( 
.A(n_244),
.B(n_314),
.C(n_265),
.Y(n_387)
);

AND2x2_ASAP7_75t_L g411 ( 
.A(n_388),
.B(n_302),
.Y(n_411)
);

CKINVDCx20_ASAP7_75t_R g390 ( 
.A(n_351),
.Y(n_390)
);

NOR2xp33_ASAP7_75t_L g450 ( 
.A(n_390),
.B(n_392),
.Y(n_450)
);

OAI21xp33_ASAP7_75t_L g392 ( 
.A1(n_355),
.A2(n_285),
.B(n_243),
.Y(n_392)
);

AOI22xp33_ASAP7_75t_SL g393 ( 
.A1(n_347),
.A2(n_253),
.B1(n_302),
.B2(n_291),
.Y(n_393)
);

AOI22xp33_ASAP7_75t_SL g476 ( 
.A1(n_393),
.A2(n_417),
.B1(n_338),
.B2(n_383),
.Y(n_476)
);

AOI22xp5_ASAP7_75t_L g457 ( 
.A1(n_394),
.A2(n_406),
.B1(n_410),
.B2(n_434),
.Y(n_457)
);

AOI22xp5_ASAP7_75t_L g395 ( 
.A1(n_353),
.A2(n_325),
.B1(n_319),
.B2(n_309),
.Y(n_395)
);

OAI22xp5_ASAP7_75t_L g460 ( 
.A1(n_395),
.A2(n_429),
.B1(n_432),
.B2(n_438),
.Y(n_460)
);

MAJIxp5_ASAP7_75t_L g466 ( 
.A(n_396),
.B(n_397),
.C(n_404),
.Y(n_466)
);

XOR2xp5_ASAP7_75t_L g397 ( 
.A(n_387),
.B(n_286),
.Y(n_397)
);

INVxp67_ASAP7_75t_L g472 ( 
.A(n_398),
.Y(n_472)
);

INVx2_ASAP7_75t_L g399 ( 
.A(n_370),
.Y(n_399)
);

INVx2_ASAP7_75t_SL g459 ( 
.A(n_399),
.Y(n_459)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_356),
.Y(n_400)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_400),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_348),
.B(n_354),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_401),
.B(n_405),
.Y(n_442)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_335),
.Y(n_402)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_402),
.Y(n_444)
);

CKINVDCx20_ASAP7_75t_R g403 ( 
.A(n_363),
.Y(n_403)
);

NOR2xp33_ASAP7_75t_L g452 ( 
.A(n_403),
.B(n_418),
.Y(n_452)
);

MAJIxp5_ASAP7_75t_SL g404 ( 
.A(n_348),
.B(n_320),
.C(n_283),
.Y(n_404)
);

AO22x1_ASAP7_75t_SL g405 ( 
.A1(n_340),
.A2(n_290),
.B1(n_297),
.B2(n_296),
.Y(n_405)
);

OAI22xp5_ASAP7_75t_SL g406 ( 
.A1(n_326),
.A2(n_306),
.B1(n_300),
.B2(n_275),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_354),
.B(n_240),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_407),
.B(n_409),
.Y(n_458)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_335),
.Y(n_408)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_408),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_331),
.B(n_249),
.Y(n_409)
);

OAI22xp5_ASAP7_75t_SL g410 ( 
.A1(n_326),
.A2(n_284),
.B1(n_242),
.B2(n_254),
.Y(n_410)
);

INVx1_ASAP7_75t_SL g480 ( 
.A(n_411),
.Y(n_480)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_344),
.Y(n_412)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_412),
.Y(n_446)
);

MAJIxp5_ASAP7_75t_L g413 ( 
.A(n_337),
.B(n_267),
.C(n_287),
.Y(n_413)
);

XNOR2xp5_ASAP7_75t_L g441 ( 
.A(n_413),
.B(n_426),
.Y(n_441)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_344),
.Y(n_414)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_414),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_331),
.B(n_303),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_415),
.B(n_424),
.Y(n_462)
);

AOI32xp33_ASAP7_75t_L g418 ( 
.A1(n_386),
.A2(n_245),
.A3(n_241),
.B1(n_255),
.B2(n_308),
.Y(n_418)
);

AOI21xp5_ASAP7_75t_L g419 ( 
.A1(n_384),
.A2(n_322),
.B(n_305),
.Y(n_419)
);

CKINVDCx16_ASAP7_75t_R g465 ( 
.A(n_419),
.Y(n_465)
);

AOI21xp5_ASAP7_75t_L g420 ( 
.A1(n_341),
.A2(n_292),
.B(n_280),
.Y(n_420)
);

CKINVDCx16_ASAP7_75t_R g481 ( 
.A(n_420),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_SL g422 ( 
.A(n_339),
.B(n_313),
.Y(n_422)
);

NOR2xp33_ASAP7_75t_L g464 ( 
.A(n_422),
.B(n_430),
.Y(n_464)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_381),
.Y(n_423)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_423),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_SL g424 ( 
.A(n_378),
.B(n_266),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_381),
.Y(n_425)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_425),
.Y(n_453)
);

XOR2xp5_ASAP7_75t_L g426 ( 
.A(n_360),
.B(n_246),
.Y(n_426)
);

AOI22xp33_ASAP7_75t_L g427 ( 
.A1(n_368),
.A2(n_238),
.B1(n_239),
.B2(n_251),
.Y(n_427)
);

AOI22xp33_ASAP7_75t_L g447 ( 
.A1(n_427),
.A2(n_328),
.B1(n_334),
.B2(n_338),
.Y(n_447)
);

OAI32xp33_ASAP7_75t_L g428 ( 
.A1(n_350),
.A2(n_346),
.A3(n_342),
.B1(n_376),
.B2(n_347),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_428),
.B(n_431),
.Y(n_474)
);

AOI22xp5_ASAP7_75t_L g429 ( 
.A1(n_361),
.A2(n_352),
.B1(n_373),
.B2(n_342),
.Y(n_429)
);

CKINVDCx20_ASAP7_75t_R g430 ( 
.A(n_367),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_350),
.B(n_368),
.Y(n_431)
);

AOI22xp5_ASAP7_75t_L g432 ( 
.A1(n_350),
.A2(n_379),
.B1(n_355),
.B2(n_366),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_355),
.B(n_336),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g479 ( 
.A(n_433),
.B(n_437),
.Y(n_479)
);

OAI22xp5_ASAP7_75t_L g434 ( 
.A1(n_388),
.A2(n_329),
.B1(n_343),
.B2(n_369),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_380),
.Y(n_435)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_435),
.Y(n_463)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_380),
.Y(n_436)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_436),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_SL g437 ( 
.A(n_336),
.B(n_377),
.Y(n_437)
);

AOI22xp5_ASAP7_75t_L g438 ( 
.A1(n_327),
.A2(n_358),
.B1(n_370),
.B2(n_334),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_L g439 ( 
.A(n_370),
.B(n_327),
.Y(n_439)
);

XNOR2xp5_ASAP7_75t_L g461 ( 
.A(n_439),
.B(n_395),
.Y(n_461)
);

CKINVDCx20_ASAP7_75t_R g440 ( 
.A(n_439),
.Y(n_440)
);

NOR2xp33_ASAP7_75t_L g484 ( 
.A(n_440),
.B(n_451),
.Y(n_484)
);

AOI22xp33_ASAP7_75t_L g518 ( 
.A1(n_447),
.A2(n_467),
.B1(n_399),
.B2(n_412),
.Y(n_518)
);

CKINVDCx20_ASAP7_75t_R g451 ( 
.A(n_438),
.Y(n_451)
);

OAI22x1_ASAP7_75t_SL g454 ( 
.A1(n_432),
.A2(n_362),
.B1(n_389),
.B2(n_328),
.Y(n_454)
);

AOI22xp5_ASAP7_75t_L g489 ( 
.A1(n_454),
.A2(n_469),
.B1(n_470),
.B2(n_478),
.Y(n_489)
);

INVx6_ASAP7_75t_L g455 ( 
.A(n_430),
.Y(n_455)
);

INVx3_ASAP7_75t_SL g502 ( 
.A(n_455),
.Y(n_502)
);

XOR2xp5_ASAP7_75t_L g456 ( 
.A(n_397),
.B(n_374),
.Y(n_456)
);

MAJIxp5_ASAP7_75t_L g504 ( 
.A(n_456),
.B(n_396),
.C(n_413),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_L g485 ( 
.A(n_461),
.B(n_405),
.Y(n_485)
);

AOI22xp33_ASAP7_75t_L g467 ( 
.A1(n_421),
.A2(n_389),
.B1(n_362),
.B2(n_374),
.Y(n_467)
);

OAI22xp5_ASAP7_75t_L g468 ( 
.A1(n_391),
.A2(n_365),
.B1(n_330),
.B2(n_364),
.Y(n_468)
);

OAI22xp5_ASAP7_75t_L g507 ( 
.A1(n_468),
.A2(n_394),
.B1(n_425),
.B2(n_423),
.Y(n_507)
);

OAI22xp5_ASAP7_75t_SL g469 ( 
.A1(n_391),
.A2(n_365),
.B1(n_385),
.B2(n_364),
.Y(n_469)
);

OAI22xp5_ASAP7_75t_SL g470 ( 
.A1(n_429),
.A2(n_365),
.B1(n_385),
.B2(n_357),
.Y(n_470)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_402),
.Y(n_473)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_473),
.Y(n_488)
);

CKINVDCx20_ASAP7_75t_R g475 ( 
.A(n_437),
.Y(n_475)
);

NOR2xp33_ASAP7_75t_L g491 ( 
.A(n_475),
.B(n_479),
.Y(n_491)
);

INVxp67_ASAP7_75t_L g493 ( 
.A(n_476),
.Y(n_493)
);

AOI22xp5_ASAP7_75t_L g477 ( 
.A1(n_421),
.A2(n_371),
.B1(n_349),
.B2(n_332),
.Y(n_477)
);

OAI22xp5_ASAP7_75t_SL g498 ( 
.A1(n_477),
.A2(n_482),
.B1(n_436),
.B2(n_435),
.Y(n_498)
);

OAI22xp5_ASAP7_75t_SL g478 ( 
.A1(n_401),
.A2(n_357),
.B1(n_330),
.B2(n_332),
.Y(n_478)
);

AOI22xp5_ASAP7_75t_L g482 ( 
.A1(n_407),
.A2(n_371),
.B1(n_349),
.B2(n_372),
.Y(n_482)
);

AOI22xp33_ASAP7_75t_SL g483 ( 
.A1(n_434),
.A2(n_372),
.B1(n_383),
.B2(n_345),
.Y(n_483)
);

OAI21xp5_ASAP7_75t_SL g492 ( 
.A1(n_483),
.A2(n_420),
.B(n_419),
.Y(n_492)
);

XNOR2xp5_ASAP7_75t_SL g554 ( 
.A(n_485),
.B(n_501),
.Y(n_554)
);

BUFx3_ASAP7_75t_L g486 ( 
.A(n_455),
.Y(n_486)
);

NOR2xp33_ASAP7_75t_L g542 ( 
.A(n_486),
.B(n_494),
.Y(n_542)
);

CKINVDCx20_ASAP7_75t_R g487 ( 
.A(n_455),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_L g549 ( 
.A(n_487),
.B(n_490),
.Y(n_549)
);

CKINVDCx20_ASAP7_75t_R g490 ( 
.A(n_464),
.Y(n_490)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_491),
.Y(n_533)
);

AO21x1_ASAP7_75t_L g558 ( 
.A1(n_492),
.A2(n_503),
.B(n_506),
.Y(n_558)
);

NAND3xp33_ASAP7_75t_L g494 ( 
.A(n_450),
.B(n_403),
.C(n_390),
.Y(n_494)
);

AOI22xp5_ASAP7_75t_L g495 ( 
.A1(n_460),
.A2(n_406),
.B1(n_431),
.B2(n_410),
.Y(n_495)
);

OAI22xp5_ASAP7_75t_SL g530 ( 
.A1(n_495),
.A2(n_518),
.B1(n_522),
.B2(n_477),
.Y(n_530)
);

CKINVDCx20_ASAP7_75t_R g496 ( 
.A(n_478),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_L g550 ( 
.A(n_496),
.B(n_498),
.Y(n_550)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_463),
.Y(n_497)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_497),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_L g499 ( 
.A(n_475),
.B(n_440),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_L g561 ( 
.A(n_499),
.B(n_500),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_458),
.B(n_415),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_L g501 ( 
.A(n_458),
.B(n_442),
.Y(n_501)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_501),
.Y(n_536)
);

XNOR2x2_ASAP7_75t_L g503 ( 
.A(n_474),
.B(n_479),
.Y(n_503)
);

MAJIxp5_ASAP7_75t_L g526 ( 
.A(n_504),
.B(n_515),
.C(n_516),
.Y(n_526)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_463),
.Y(n_505)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_505),
.Y(n_553)
);

OR2x2_ASAP7_75t_L g506 ( 
.A(n_474),
.B(n_404),
.Y(n_506)
);

AOI22xp5_ASAP7_75t_L g531 ( 
.A1(n_507),
.A2(n_512),
.B1(n_517),
.B2(n_457),
.Y(n_531)
);

CKINVDCx20_ASAP7_75t_R g508 ( 
.A(n_482),
.Y(n_508)
);

NOR2xp33_ASAP7_75t_L g555 ( 
.A(n_508),
.B(n_511),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_L g509 ( 
.A(n_442),
.B(n_409),
.Y(n_509)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_509),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_L g510 ( 
.A(n_462),
.B(n_400),
.Y(n_510)
);

XOR2x1_ASAP7_75t_L g562 ( 
.A(n_510),
.B(n_520),
.Y(n_562)
);

AO21x1_ASAP7_75t_L g511 ( 
.A1(n_452),
.A2(n_416),
.B(n_472),
.Y(n_511)
);

OAI22xp5_ASAP7_75t_L g512 ( 
.A1(n_460),
.A2(n_428),
.B1(n_426),
.B2(n_405),
.Y(n_512)
);

HB1xp67_ASAP7_75t_L g513 ( 
.A(n_443),
.Y(n_513)
);

CKINVDCx20_ASAP7_75t_R g528 ( 
.A(n_513),
.Y(n_528)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_471),
.Y(n_514)
);

CKINVDCx20_ASAP7_75t_R g540 ( 
.A(n_514),
.Y(n_540)
);

MAJIxp5_ASAP7_75t_L g515 ( 
.A(n_456),
.B(n_416),
.C(n_433),
.Y(n_515)
);

MAJIxp5_ASAP7_75t_L g516 ( 
.A(n_441),
.B(n_424),
.C(n_405),
.Y(n_516)
);

OAI22xp5_ASAP7_75t_SL g517 ( 
.A1(n_451),
.A2(n_411),
.B1(n_418),
.B2(n_408),
.Y(n_517)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_471),
.Y(n_519)
);

CKINVDCx20_ASAP7_75t_R g543 ( 
.A(n_519),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_L g520 ( 
.A(n_462),
.B(n_414),
.Y(n_520)
);

NAND2xp33_ASAP7_75t_SL g521 ( 
.A(n_480),
.B(n_411),
.Y(n_521)
);

XOR2xp5_ASAP7_75t_L g525 ( 
.A(n_521),
.B(n_461),
.Y(n_525)
);

AOI22xp5_ASAP7_75t_L g522 ( 
.A1(n_454),
.A2(n_371),
.B1(n_345),
.B2(n_359),
.Y(n_522)
);

A2O1A1O1Ixp25_ASAP7_75t_L g523 ( 
.A1(n_466),
.A2(n_345),
.B(n_359),
.C(n_472),
.D(n_480),
.Y(n_523)
);

XNOR2xp5_ASAP7_75t_L g529 ( 
.A(n_523),
.B(n_466),
.Y(n_529)
);

NOR2xp33_ASAP7_75t_L g524 ( 
.A(n_443),
.B(n_448),
.Y(n_524)
);

CKINVDCx20_ASAP7_75t_R g545 ( 
.A(n_524),
.Y(n_545)
);

AND2x2_ASAP7_75t_L g573 ( 
.A(n_525),
.B(n_530),
.Y(n_573)
);

XOR2xp5_ASAP7_75t_L g527 ( 
.A(n_515),
.B(n_441),
.Y(n_527)
);

XOR2xp5_ASAP7_75t_L g588 ( 
.A(n_527),
.B(n_539),
.Y(n_588)
);

XOR2x2_ASAP7_75t_L g591 ( 
.A(n_529),
.B(n_521),
.Y(n_591)
);

OAI22xp5_ASAP7_75t_SL g569 ( 
.A1(n_531),
.A2(n_532),
.B1(n_537),
.B2(n_538),
.Y(n_569)
);

AOI22xp5_ASAP7_75t_L g532 ( 
.A1(n_512),
.A2(n_465),
.B1(n_470),
.B2(n_457),
.Y(n_532)
);

OAI22xp5_ASAP7_75t_SL g535 ( 
.A1(n_484),
.A2(n_465),
.B1(n_481),
.B2(n_446),
.Y(n_535)
);

AOI22xp5_ASAP7_75t_L g578 ( 
.A1(n_535),
.A2(n_544),
.B1(n_488),
.B2(n_519),
.Y(n_578)
);

AOI22xp5_ASAP7_75t_L g537 ( 
.A1(n_517),
.A2(n_469),
.B1(n_468),
.B2(n_481),
.Y(n_537)
);

AOI22xp5_ASAP7_75t_L g538 ( 
.A1(n_484),
.A2(n_444),
.B1(n_445),
.B2(n_446),
.Y(n_538)
);

XNOR2xp5_ASAP7_75t_L g539 ( 
.A(n_504),
.B(n_444),
.Y(n_539)
);

XOR2xp5_ASAP7_75t_L g541 ( 
.A(n_503),
.B(n_445),
.Y(n_541)
);

XOR2xp5_ASAP7_75t_L g590 ( 
.A(n_541),
.B(n_548),
.Y(n_590)
);

OAI22xp5_ASAP7_75t_SL g544 ( 
.A1(n_509),
.A2(n_473),
.B1(n_449),
.B2(n_453),
.Y(n_544)
);

MAJIxp5_ASAP7_75t_L g546 ( 
.A(n_516),
.B(n_448),
.C(n_449),
.Y(n_546)
);

MAJIxp5_ASAP7_75t_L g585 ( 
.A(n_546),
.B(n_556),
.C(n_488),
.Y(n_585)
);

AOI22xp5_ASAP7_75t_L g547 ( 
.A1(n_485),
.A2(n_453),
.B1(n_459),
.B2(n_508),
.Y(n_547)
);

OAI22xp5_ASAP7_75t_SL g583 ( 
.A1(n_547),
.A2(n_557),
.B1(n_559),
.B2(n_500),
.Y(n_583)
);

XNOR2xp5_ASAP7_75t_L g548 ( 
.A(n_503),
.B(n_459),
.Y(n_548)
);

XOR2xp5_ASAP7_75t_L g551 ( 
.A(n_510),
.B(n_459),
.Y(n_551)
);

XOR2xp5_ASAP7_75t_L g593 ( 
.A(n_551),
.B(n_552),
.Y(n_593)
);

XOR2xp5_ASAP7_75t_L g552 ( 
.A(n_506),
.B(n_511),
.Y(n_552)
);

HB1xp67_ASAP7_75t_L g568 ( 
.A(n_554),
.Y(n_568)
);

XOR2xp5_ASAP7_75t_L g556 ( 
.A(n_506),
.B(n_511),
.Y(n_556)
);

AOI22xp5_ASAP7_75t_L g557 ( 
.A1(n_496),
.A2(n_499),
.B1(n_507),
.B2(n_495),
.Y(n_557)
);

AOI22xp5_ASAP7_75t_L g559 ( 
.A1(n_498),
.A2(n_491),
.B1(n_487),
.B2(n_520),
.Y(n_559)
);

INVxp33_ASAP7_75t_L g563 ( 
.A(n_549),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_L g598 ( 
.A(n_563),
.B(n_577),
.Y(n_598)
);

OAI21xp5_ASAP7_75t_SL g564 ( 
.A1(n_555),
.A2(n_492),
.B(n_523),
.Y(n_564)
);

OAI21xp5_ASAP7_75t_SL g595 ( 
.A1(n_564),
.A2(n_558),
.B(n_532),
.Y(n_595)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_549),
.Y(n_565)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_565),
.Y(n_597)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_538),
.Y(n_566)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_566),
.Y(n_600)
);

INVxp67_ASAP7_75t_SL g567 ( 
.A(n_542),
.Y(n_567)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_567),
.Y(n_606)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_533),
.Y(n_570)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_570),
.Y(n_594)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_544),
.Y(n_571)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_571),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_SL g572 ( 
.A(n_539),
.B(n_490),
.Y(n_572)
);

NOR2xp33_ASAP7_75t_L g610 ( 
.A(n_572),
.B(n_576),
.Y(n_610)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_534),
.Y(n_574)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_574),
.Y(n_611)
);

AOI22x1_ASAP7_75t_L g575 ( 
.A1(n_530),
.A2(n_502),
.B1(n_486),
.B2(n_493),
.Y(n_575)
);

OAI22xp5_ASAP7_75t_L g596 ( 
.A1(n_575),
.A2(n_578),
.B1(n_584),
.B2(n_586),
.Y(n_596)
);

NOR2xp33_ASAP7_75t_L g576 ( 
.A(n_546),
.B(n_524),
.Y(n_576)
);

INVxp33_ASAP7_75t_L g577 ( 
.A(n_559),
.Y(n_577)
);

XNOR2xp5_ASAP7_75t_SL g579 ( 
.A(n_529),
.B(n_523),
.Y(n_579)
);

XOR2xp5_ASAP7_75t_L g619 ( 
.A(n_579),
.B(n_591),
.Y(n_619)
);

CKINVDCx20_ASAP7_75t_R g580 ( 
.A(n_561),
.Y(n_580)
);

NOR2xp33_ASAP7_75t_L g617 ( 
.A(n_580),
.B(n_589),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_L g581 ( 
.A(n_545),
.B(n_502),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_L g605 ( 
.A(n_581),
.B(n_582),
.Y(n_605)
);

INVxp33_ASAP7_75t_L g582 ( 
.A(n_550),
.Y(n_582)
);

AOI22xp5_ASAP7_75t_L g602 ( 
.A1(n_583),
.A2(n_550),
.B1(n_536),
.B2(n_551),
.Y(n_602)
);

AOI22xp5_ASAP7_75t_L g584 ( 
.A1(n_531),
.A2(n_489),
.B1(n_502),
.B2(n_522),
.Y(n_584)
);

XNOR2xp5_ASAP7_75t_L g599 ( 
.A(n_585),
.B(n_591),
.Y(n_599)
);

AOI22xp5_ASAP7_75t_L g586 ( 
.A1(n_557),
.A2(n_489),
.B1(n_497),
.B2(n_505),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_L g587 ( 
.A(n_561),
.B(n_514),
.Y(n_587)
);

INVx2_ASAP7_75t_L g612 ( 
.A(n_587),
.Y(n_612)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_553),
.Y(n_589)
);

HB1xp67_ASAP7_75t_L g592 ( 
.A(n_562),
.Y(n_592)
);

OAI22xp5_ASAP7_75t_L g608 ( 
.A1(n_592),
.A2(n_541),
.B1(n_548),
.B2(n_556),
.Y(n_608)
);

AOI21x1_ASAP7_75t_SL g621 ( 
.A1(n_595),
.A2(n_613),
.B(n_573),
.Y(n_621)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_602),
.Y(n_630)
);

OAI22xp5_ASAP7_75t_SL g603 ( 
.A1(n_577),
.A2(n_560),
.B1(n_547),
.B2(n_537),
.Y(n_603)
);

INVxp67_ASAP7_75t_L g628 ( 
.A(n_603),
.Y(n_628)
);

XNOR2xp5_ASAP7_75t_L g604 ( 
.A(n_588),
.B(n_552),
.Y(n_604)
);

NOR2xp33_ASAP7_75t_L g623 ( 
.A(n_604),
.B(n_618),
.Y(n_623)
);

MAJIxp5_ASAP7_75t_L g607 ( 
.A(n_588),
.B(n_526),
.C(n_527),
.Y(n_607)
);

MAJIxp5_ASAP7_75t_L g624 ( 
.A(n_607),
.B(n_614),
.C(n_615),
.Y(n_624)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_608),
.Y(n_627)
);

AOI22xp5_ASAP7_75t_L g609 ( 
.A1(n_569),
.A2(n_535),
.B1(n_525),
.B2(n_562),
.Y(n_609)
);

INVx2_ASAP7_75t_L g632 ( 
.A(n_609),
.Y(n_632)
);

OAI21xp5_ASAP7_75t_SL g613 ( 
.A1(n_564),
.A2(n_558),
.B(n_540),
.Y(n_613)
);

MAJIxp5_ASAP7_75t_L g614 ( 
.A(n_585),
.B(n_526),
.C(n_554),
.Y(n_614)
);

MAJIxp5_ASAP7_75t_L g615 ( 
.A(n_593),
.B(n_528),
.C(n_543),
.Y(n_615)
);

MAJIxp5_ASAP7_75t_L g616 ( 
.A(n_593),
.B(n_579),
.C(n_590),
.Y(n_616)
);

MAJIxp5_ASAP7_75t_L g625 ( 
.A(n_616),
.B(n_568),
.C(n_570),
.Y(n_625)
);

XNOR2xp5_ASAP7_75t_L g618 ( 
.A(n_590),
.B(n_573),
.Y(n_618)
);

XOR2xp5_ASAP7_75t_SL g635 ( 
.A(n_619),
.B(n_578),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_L g620 ( 
.A(n_605),
.B(n_563),
.Y(n_620)
);

CKINVDCx20_ASAP7_75t_R g643 ( 
.A(n_620),
.Y(n_643)
);

OAI21xp5_ASAP7_75t_L g645 ( 
.A1(n_621),
.A2(n_613),
.B(n_598),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_L g622 ( 
.A(n_605),
.B(n_581),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_L g649 ( 
.A(n_622),
.B(n_629),
.Y(n_649)
);

XNOR2xp5_ASAP7_75t_L g646 ( 
.A(n_625),
.B(n_631),
.Y(n_646)
);

MAJIxp5_ASAP7_75t_L g626 ( 
.A(n_614),
.B(n_573),
.C(n_582),
.Y(n_626)
);

MAJIxp5_ASAP7_75t_L g644 ( 
.A(n_626),
.B(n_636),
.C(n_638),
.Y(n_644)
);

FAx1_ASAP7_75t_SL g629 ( 
.A(n_616),
.B(n_619),
.CI(n_583),
.CON(n_629),
.SN(n_629)
);

XOR2xp5_ASAP7_75t_L g631 ( 
.A(n_604),
.B(n_569),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_L g633 ( 
.A(n_617),
.B(n_587),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_L g651 ( 
.A(n_633),
.B(n_637),
.Y(n_651)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_594),
.Y(n_634)
);

NOR2xp33_ASAP7_75t_L g642 ( 
.A(n_634),
.B(n_639),
.Y(n_642)
);

XOR2xp5_ASAP7_75t_L g650 ( 
.A(n_635),
.B(n_603),
.Y(n_650)
);

MAJIxp5_ASAP7_75t_L g636 ( 
.A(n_607),
.B(n_565),
.C(n_586),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_L g637 ( 
.A(n_598),
.B(n_584),
.Y(n_637)
);

MAJIxp5_ASAP7_75t_L g638 ( 
.A(n_615),
.B(n_575),
.C(n_599),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_594),
.Y(n_639)
);

MAJIxp5_ASAP7_75t_L g640 ( 
.A(n_599),
.B(n_575),
.C(n_618),
.Y(n_640)
);

MAJIxp5_ASAP7_75t_L g647 ( 
.A(n_640),
.B(n_641),
.C(n_601),
.Y(n_647)
);

MAJIxp5_ASAP7_75t_L g641 ( 
.A(n_609),
.B(n_610),
.C(n_595),
.Y(n_641)
);

OR2x2_ASAP7_75t_L g661 ( 
.A(n_645),
.B(n_650),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_L g665 ( 
.A(n_647),
.B(n_648),
.Y(n_665)
);

MAJIxp5_ASAP7_75t_L g648 ( 
.A(n_636),
.B(n_624),
.C(n_626),
.Y(n_648)
);

OAI22xp5_ASAP7_75t_SL g652 ( 
.A1(n_628),
.A2(n_600),
.B1(n_601),
.B2(n_597),
.Y(n_652)
);

AOI22xp5_ASAP7_75t_L g668 ( 
.A1(n_652),
.A2(n_658),
.B1(n_637),
.B2(n_632),
.Y(n_668)
);

NOR2xp33_ASAP7_75t_L g653 ( 
.A(n_641),
.B(n_606),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_L g669 ( 
.A(n_653),
.B(n_654),
.Y(n_669)
);

MAJIxp5_ASAP7_75t_L g654 ( 
.A(n_624),
.B(n_596),
.C(n_602),
.Y(n_654)
);

NOR2xp67_ASAP7_75t_L g655 ( 
.A(n_625),
.B(n_612),
.Y(n_655)
);

AOI21x1_ASAP7_75t_L g666 ( 
.A1(n_655),
.A2(n_630),
.B(n_640),
.Y(n_666)
);

CKINVDCx5p33_ASAP7_75t_R g656 ( 
.A(n_620),
.Y(n_656)
);

OAI21xp5_ASAP7_75t_L g670 ( 
.A1(n_656),
.A2(n_657),
.B(n_635),
.Y(n_670)
);

AOI21xp5_ASAP7_75t_L g657 ( 
.A1(n_622),
.A2(n_612),
.B(n_611),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_L g658 ( 
.A(n_633),
.B(n_611),
.Y(n_658)
);

MAJIxp5_ASAP7_75t_L g659 ( 
.A(n_648),
.B(n_631),
.C(n_627),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_L g672 ( 
.A(n_659),
.B(n_660),
.Y(n_672)
);

MAJIxp5_ASAP7_75t_L g660 ( 
.A(n_644),
.B(n_638),
.C(n_628),
.Y(n_660)
);

NOR2xp33_ASAP7_75t_SL g662 ( 
.A(n_642),
.B(n_658),
.Y(n_662)
);

NOR2xp33_ASAP7_75t_L g673 ( 
.A(n_662),
.B(n_643),
.Y(n_673)
);

NOR2xp33_ASAP7_75t_L g663 ( 
.A(n_647),
.B(n_630),
.Y(n_663)
);

AOI21xp5_ASAP7_75t_L g676 ( 
.A1(n_663),
.A2(n_664),
.B(n_666),
.Y(n_676)
);

OAI21xp5_ASAP7_75t_SL g664 ( 
.A1(n_649),
.A2(n_645),
.B(n_621),
.Y(n_664)
);

MAJIxp5_ASAP7_75t_L g667 ( 
.A(n_644),
.B(n_632),
.C(n_623),
.Y(n_667)
);

MAJIxp5_ASAP7_75t_L g671 ( 
.A(n_667),
.B(n_646),
.C(n_654),
.Y(n_671)
);

XOR2xp5_ASAP7_75t_L g674 ( 
.A(n_668),
.B(n_670),
.Y(n_674)
);

NOR2xp67_ASAP7_75t_SL g679 ( 
.A(n_671),
.B(n_660),
.Y(n_679)
);

NOR2xp33_ASAP7_75t_SL g683 ( 
.A(n_673),
.B(n_675),
.Y(n_683)
);

NOR2xp33_ASAP7_75t_L g675 ( 
.A(n_667),
.B(n_649),
.Y(n_675)
);

NOR2xp33_ASAP7_75t_L g677 ( 
.A(n_669),
.B(n_651),
.Y(n_677)
);

AOI21xp5_ASAP7_75t_L g682 ( 
.A1(n_677),
.A2(n_678),
.B(n_646),
.Y(n_682)
);

OAI21xp5_ASAP7_75t_SL g678 ( 
.A1(n_665),
.A2(n_670),
.B(n_661),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_L g685 ( 
.A(n_679),
.B(n_680),
.Y(n_685)
);

NOR2xp33_ASAP7_75t_L g680 ( 
.A(n_671),
.B(n_661),
.Y(n_680)
);

AOI21x1_ASAP7_75t_L g681 ( 
.A1(n_676),
.A2(n_659),
.B(n_651),
.Y(n_681)
);

AOI21xp5_ASAP7_75t_L g684 ( 
.A1(n_681),
.A2(n_682),
.B(n_672),
.Y(n_684)
);

AOI21xp5_ASAP7_75t_L g686 ( 
.A1(n_684),
.A2(n_683),
.B(n_674),
.Y(n_686)
);

MAJIxp5_ASAP7_75t_L g687 ( 
.A(n_686),
.B(n_685),
.C(n_674),
.Y(n_687)
);

AOI21xp5_ASAP7_75t_L g688 ( 
.A1(n_687),
.A2(n_657),
.B(n_652),
.Y(n_688)
);

XOR2xp5_ASAP7_75t_L g689 ( 
.A(n_688),
.B(n_650),
.Y(n_689)
);

AOI22xp33_ASAP7_75t_L g690 ( 
.A1(n_689),
.A2(n_629),
.B1(n_656),
.B2(n_687),
.Y(n_690)
);


endmodule