module fake_netlist_6_2210_n_119 (n_16, n_1, n_9, n_8, n_18, n_10, n_21, n_24, n_6, n_15, n_27, n_3, n_14, n_0, n_4, n_22, n_26, n_13, n_11, n_28, n_17, n_23, n_12, n_20, n_7, n_30, n_2, n_5, n_19, n_29, n_25, n_119);

input n_16;
input n_1;
input n_9;
input n_8;
input n_18;
input n_10;
input n_21;
input n_24;
input n_6;
input n_15;
input n_27;
input n_3;
input n_14;
input n_0;
input n_4;
input n_22;
input n_26;
input n_13;
input n_11;
input n_28;
input n_17;
input n_23;
input n_12;
input n_20;
input n_7;
input n_30;
input n_2;
input n_5;
input n_19;
input n_29;
input n_25;

output n_119;

wire n_52;
wire n_91;
wire n_46;
wire n_88;
wire n_98;
wire n_113;
wire n_63;
wire n_39;
wire n_73;
wire n_68;
wire n_50;
wire n_49;
wire n_83;
wire n_101;
wire n_77;
wire n_106;
wire n_92;
wire n_42;
wire n_96;
wire n_90;
wire n_105;
wire n_54;
wire n_102;
wire n_87;
wire n_32;
wire n_66;
wire n_99;
wire n_85;
wire n_78;
wire n_84;
wire n_100;
wire n_47;
wire n_62;
wire n_75;
wire n_109;
wire n_45;
wire n_34;
wire n_70;
wire n_37;
wire n_67;
wire n_33;
wire n_82;
wire n_38;
wire n_110;
wire n_61;
wire n_112;
wire n_81;
wire n_59;
wire n_76;
wire n_36;
wire n_55;
wire n_94;
wire n_97;
wire n_108;
wire n_58;
wire n_116;
wire n_64;
wire n_117;
wire n_118;
wire n_48;
wire n_65;
wire n_93;
wire n_40;
wire n_80;
wire n_41;
wire n_114;
wire n_86;
wire n_104;
wire n_95;
wire n_107;
wire n_71;
wire n_74;
wire n_72;
wire n_89;
wire n_103;
wire n_111;
wire n_60;
wire n_35;
wire n_115;
wire n_69;
wire n_79;
wire n_43;
wire n_31;
wire n_57;
wire n_53;
wire n_51;
wire n_44;
wire n_56;

INVx1_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_L g33 ( 
.A1(n_11),
.A2(n_16),
.B1(n_13),
.B2(n_6),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_26),
.Y(n_34)
);

AND2x2_ASAP7_75t_L g35 ( 
.A(n_5),
.B(n_4),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_8),
.Y(n_36)
);

BUFx2_ASAP7_75t_L g37 ( 
.A(n_29),
.Y(n_37)
);

HB1xp67_ASAP7_75t_L g38 ( 
.A(n_27),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_6),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_20),
.B(n_15),
.Y(n_40)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_5),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_2),
.Y(n_42)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_9),
.Y(n_43)
);

AND2x6_ASAP7_75t_L g44 ( 
.A(n_14),
.B(n_24),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_7),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_18),
.B(n_1),
.Y(n_46)
);

INVxp67_ASAP7_75t_L g47 ( 
.A(n_4),
.Y(n_47)
);

AND2x2_ASAP7_75t_L g48 ( 
.A(n_1),
.B(n_21),
.Y(n_48)
);

AND2x2_ASAP7_75t_L g49 ( 
.A(n_10),
.B(n_17),
.Y(n_49)
);

AND2x4_ASAP7_75t_L g50 ( 
.A(n_25),
.B(n_28),
.Y(n_50)
);

BUFx2_ASAP7_75t_L g51 ( 
.A(n_3),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_22),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_12),
.Y(n_53)
);

HB1xp67_ASAP7_75t_L g54 ( 
.A(n_30),
.Y(n_54)
);

BUFx6f_ASAP7_75t_SL g55 ( 
.A(n_41),
.Y(n_55)
);

NOR3xp33_ASAP7_75t_L g56 ( 
.A(n_41),
.B(n_0),
.C(n_19),
.Y(n_56)
);

NAND2xp33_ASAP7_75t_L g57 ( 
.A(n_35),
.B(n_0),
.Y(n_57)
);

NAND2xp33_ASAP7_75t_L g58 ( 
.A(n_42),
.B(n_23),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_42),
.Y(n_59)
);

OR2x2_ASAP7_75t_L g60 ( 
.A(n_51),
.B(n_47),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_38),
.B(n_54),
.Y(n_61)
);

NAND2xp33_ASAP7_75t_L g62 ( 
.A(n_42),
.B(n_48),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_38),
.B(n_54),
.Y(n_63)
);

INVx1_ASAP7_75t_SL g64 ( 
.A(n_34),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_37),
.B(n_53),
.Y(n_65)
);

INVx2_ASAP7_75t_SL g66 ( 
.A(n_32),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_42),
.B(n_43),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_43),
.B(n_50),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_59),
.Y(n_69)
);

INVx1_ASAP7_75t_SL g70 ( 
.A(n_64),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_63),
.B(n_36),
.Y(n_71)
);

AND2x2_ASAP7_75t_L g72 ( 
.A(n_65),
.B(n_31),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_66),
.Y(n_73)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_55),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_67),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_68),
.Y(n_76)
);

BUFx3_ASAP7_75t_L g77 ( 
.A(n_60),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_63),
.A2(n_46),
.B1(n_34),
.B2(n_49),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_61),
.B(n_50),
.Y(n_79)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_69),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_76),
.Y(n_81)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_69),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_76),
.B(n_68),
.Y(n_83)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_69),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_69),
.Y(n_85)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_69),
.Y(n_86)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_73),
.Y(n_87)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_73),
.Y(n_88)
);

BUFx3_ASAP7_75t_L g89 ( 
.A(n_75),
.Y(n_89)
);

OAI21xp33_ASAP7_75t_SL g90 ( 
.A1(n_79),
.A2(n_46),
.B(n_39),
.Y(n_90)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_84),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_83),
.B(n_72),
.Y(n_92)
);

OR2x2_ASAP7_75t_L g93 ( 
.A(n_89),
.B(n_70),
.Y(n_93)
);

OR2x2_ASAP7_75t_L g94 ( 
.A(n_89),
.B(n_77),
.Y(n_94)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_88),
.Y(n_95)
);

AND2x2_ASAP7_75t_L g96 ( 
.A(n_83),
.B(n_72),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_81),
.B(n_77),
.Y(n_97)
);

AND2x2_ASAP7_75t_L g98 ( 
.A(n_96),
.B(n_92),
.Y(n_98)
);

OR2x2_ASAP7_75t_L g99 ( 
.A(n_93),
.B(n_78),
.Y(n_99)
);

AND2x4_ASAP7_75t_L g100 ( 
.A(n_95),
.B(n_87),
.Y(n_100)
);

INVx1_ASAP7_75t_SL g101 ( 
.A(n_94),
.Y(n_101)
);

HB1xp67_ASAP7_75t_L g102 ( 
.A(n_101),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_99),
.Y(n_103)
);

OAI31xp33_ASAP7_75t_L g104 ( 
.A1(n_99),
.A2(n_92),
.A3(n_71),
.B(n_97),
.Y(n_104)
);

AO21x1_ASAP7_75t_L g105 ( 
.A1(n_98),
.A2(n_57),
.B(n_62),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_103),
.A2(n_98),
.B1(n_90),
.B2(n_100),
.Y(n_106)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_102),
.Y(n_107)
);

AOI21xp5_ASAP7_75t_L g108 ( 
.A1(n_104),
.A2(n_91),
.B(n_100),
.Y(n_108)
);

NOR3xp33_ASAP7_75t_L g109 ( 
.A(n_105),
.B(n_74),
.C(n_75),
.Y(n_109)
);

AOI322xp5_ASAP7_75t_L g110 ( 
.A1(n_107),
.A2(n_47),
.A3(n_56),
.B1(n_52),
.B2(n_45),
.C1(n_88),
.C2(n_58),
.Y(n_110)
);

AOI222xp33_ASAP7_75t_L g111 ( 
.A1(n_106),
.A2(n_33),
.B1(n_44),
.B2(n_100),
.C1(n_40),
.C2(n_74),
.Y(n_111)
);

NAND4xp75_ASAP7_75t_L g112 ( 
.A(n_111),
.B(n_105),
.C(n_108),
.D(n_109),
.Y(n_112)
);

AOI21xp5_ASAP7_75t_L g113 ( 
.A1(n_110),
.A2(n_91),
.B(n_82),
.Y(n_113)
);

OAI311xp33_ASAP7_75t_L g114 ( 
.A1(n_111),
.A2(n_74),
.A3(n_85),
.B1(n_84),
.C1(n_44),
.Y(n_114)
);

XOR2xp5_ASAP7_75t_L g115 ( 
.A(n_112),
.B(n_113),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_114),
.A2(n_80),
.B1(n_82),
.B2(n_86),
.Y(n_116)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_116),
.Y(n_117)
);

AOI21xp5_ASAP7_75t_L g118 ( 
.A1(n_117),
.A2(n_44),
.B(n_115),
.Y(n_118)
);

OR2x6_ASAP7_75t_L g119 ( 
.A(n_118),
.B(n_44),
.Y(n_119)
);


endmodule