module fake_jpeg_4034_n_137 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_137);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_137;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_6),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_5),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_4),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g15 ( 
.A(n_0),
.B(n_4),
.Y(n_15)
);

INVx3_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

BUFx8_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

INVx11_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_3),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_0),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_6),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_8),
.Y(n_25)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_22),
.Y(n_26)
);

INVx5_ASAP7_75t_L g37 ( 
.A(n_26),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_SL g27 ( 
.A(n_15),
.B(n_23),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_SL g41 ( 
.A(n_27),
.B(n_33),
.Y(n_41)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_22),
.Y(n_28)
);

BUFx8_ASAP7_75t_L g44 ( 
.A(n_28),
.Y(n_44)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_22),
.Y(n_29)
);

BUFx16f_ASAP7_75t_L g45 ( 
.A(n_29),
.Y(n_45)
);

INVx4_ASAP7_75t_SL g30 ( 
.A(n_17),
.Y(n_30)
);

OR2x2_ASAP7_75t_SL g34 ( 
.A(n_30),
.B(n_32),
.Y(n_34)
);

INVx3_ASAP7_75t_SL g31 ( 
.A(n_17),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_31),
.Y(n_42)
);

AND2x2_ASAP7_75t_L g32 ( 
.A(n_17),
.B(n_1),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_16),
.B(n_14),
.Y(n_33)
);

AOI22xp33_ASAP7_75t_SL g35 ( 
.A1(n_30),
.A2(n_16),
.B1(n_18),
.B2(n_21),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_L g51 ( 
.A1(n_35),
.A2(n_38),
.B1(n_40),
.B2(n_39),
.Y(n_51)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_28),
.Y(n_36)
);

INVx5_ASAP7_75t_L g59 ( 
.A(n_36),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_L g38 ( 
.A1(n_32),
.A2(n_16),
.B1(n_25),
.B2(n_18),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_32),
.B(n_13),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_39),
.B(n_32),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_L g40 ( 
.A1(n_32),
.A2(n_25),
.B1(n_18),
.B2(n_21),
.Y(n_40)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_28),
.Y(n_43)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_43),
.Y(n_50)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_37),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_46),
.B(n_47),
.Y(n_68)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_37),
.Y(n_47)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_45),
.Y(n_48)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_48),
.Y(n_67)
);

AND2x2_ASAP7_75t_L g69 ( 
.A(n_49),
.B(n_30),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g60 ( 
.A1(n_51),
.A2(n_54),
.B1(n_27),
.B2(n_19),
.Y(n_60)
);

AOI21xp5_ASAP7_75t_L g52 ( 
.A1(n_34),
.A2(n_33),
.B(n_30),
.Y(n_52)
);

OAI21xp5_ASAP7_75t_SL g75 ( 
.A1(n_52),
.A2(n_31),
.B(n_29),
.Y(n_75)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_45),
.Y(n_53)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_53),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g54 ( 
.A1(n_41),
.A2(n_33),
.B1(n_27),
.B2(n_12),
.Y(n_54)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_45),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_SL g63 ( 
.A(n_55),
.B(n_56),
.Y(n_63)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_44),
.Y(n_56)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_42),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_SL g72 ( 
.A(n_57),
.B(n_58),
.Y(n_72)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_44),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_60),
.B(n_73),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_50),
.B(n_52),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_SL g78 ( 
.A(n_61),
.B(n_69),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_47),
.B(n_34),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_62),
.B(n_74),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_59),
.B(n_19),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_64),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_SL g65 ( 
.A(n_59),
.B(n_30),
.C(n_31),
.Y(n_65)
);

OAI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_65),
.A2(n_29),
.B1(n_36),
.B2(n_43),
.Y(n_76)
);

XNOR2xp5_ASAP7_75t_L g66 ( 
.A(n_46),
.B(n_31),
.Y(n_66)
);

XOR2xp5_ASAP7_75t_L g88 ( 
.A(n_66),
.B(n_75),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_53),
.B(n_24),
.Y(n_71)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_71),
.Y(n_77)
);

O2A1O1Ixp33_ASAP7_75t_L g73 ( 
.A1(n_57),
.A2(n_31),
.B(n_28),
.C(n_29),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_55),
.B(n_44),
.Y(n_74)
);

AND2x2_ASAP7_75t_L g96 ( 
.A(n_76),
.B(n_65),
.Y(n_96)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_68),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_79),
.B(n_80),
.Y(n_93)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_72),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_63),
.B(n_42),
.Y(n_82)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_82),
.Y(n_97)
);

HB1xp67_ASAP7_75t_L g84 ( 
.A(n_70),
.Y(n_84)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_84),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_69),
.A2(n_42),
.B1(n_12),
.B2(n_23),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g91 ( 
.A(n_85),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_69),
.B(n_17),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_87),
.B(n_66),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_75),
.A2(n_26),
.B1(n_20),
.B2(n_24),
.Y(n_89)
);

INVxp67_ASAP7_75t_L g95 ( 
.A(n_89),
.Y(n_95)
);

OAI21xp5_ASAP7_75t_L g90 ( 
.A1(n_87),
.A2(n_62),
.B(n_60),
.Y(n_90)
);

AOI21xp5_ASAP7_75t_L g104 ( 
.A1(n_90),
.A2(n_81),
.B(n_89),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_92),
.B(n_85),
.Y(n_105)
);

XNOR2xp5_ASAP7_75t_L g94 ( 
.A(n_88),
.B(n_74),
.Y(n_94)
);

XOR2xp5_ASAP7_75t_L g107 ( 
.A(n_94),
.B(n_99),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_96),
.A2(n_77),
.B1(n_83),
.B2(n_26),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_88),
.B(n_67),
.C(n_73),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_86),
.B(n_26),
.C(n_15),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_100),
.B(n_101),
.Y(n_111)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_86),
.Y(n_101)
);

OAI21xp33_ASAP7_75t_L g102 ( 
.A1(n_96),
.A2(n_78),
.B(n_99),
.Y(n_102)
);

OAI21xp5_ASAP7_75t_SL g114 ( 
.A1(n_102),
.A2(n_104),
.B(n_108),
.Y(n_114)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_93),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_SL g112 ( 
.A(n_103),
.B(n_105),
.Y(n_112)
);

A2O1A1O1Ixp25_ASAP7_75t_L g106 ( 
.A1(n_95),
.A2(n_80),
.B(n_77),
.C(n_83),
.D(n_79),
.Y(n_106)
);

XNOR2xp5_ASAP7_75t_L g113 ( 
.A(n_106),
.B(n_95),
.Y(n_113)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_100),
.Y(n_108)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_98),
.Y(n_109)
);

NAND2xp33_ASAP7_75t_SL g118 ( 
.A(n_109),
.B(n_1),
.Y(n_118)
);

FAx1_ASAP7_75t_SL g116 ( 
.A(n_110),
.B(n_91),
.CI(n_14),
.CON(n_116),
.SN(n_116)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_113),
.B(n_116),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_107),
.B(n_97),
.C(n_91),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_115),
.B(n_107),
.C(n_17),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_110),
.A2(n_20),
.B1(n_13),
.B2(n_14),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_117),
.B(n_118),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_112),
.B(n_111),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_119),
.B(n_113),
.Y(n_125)
);

AOI21xp5_ASAP7_75t_L g120 ( 
.A1(n_114),
.A2(n_102),
.B(n_106),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_120),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_122),
.B(n_124),
.C(n_116),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_115),
.B(n_14),
.C(n_7),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_L g130 ( 
.A1(n_125),
.A2(n_126),
.B(n_127),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_123),
.A2(n_114),
.B1(n_116),
.B2(n_117),
.Y(n_126)
);

AOI21xp5_ASAP7_75t_SL g128 ( 
.A1(n_121),
.A2(n_10),
.B(n_9),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_L g132 ( 
.A1(n_128),
.A2(n_129),
.B(n_9),
.Y(n_132)
);

AOI21xp33_ASAP7_75t_L g131 ( 
.A1(n_125),
.A2(n_7),
.B(n_8),
.Y(n_131)
);

AOI21xp5_ASAP7_75t_L g133 ( 
.A1(n_131),
.A2(n_2),
.B(n_3),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_132),
.B(n_6),
.Y(n_134)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_133),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_L g136 ( 
.A1(n_135),
.A2(n_130),
.B(n_134),
.Y(n_136)
);

XOR2xp5_ASAP7_75t_L g137 ( 
.A(n_136),
.B(n_2),
.Y(n_137)
);


endmodule