module fake_jpeg_25697_n_200 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_200);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_200;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

INVx2_ASAP7_75t_L g15 ( 
.A(n_11),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_9),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_5),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_2),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_10),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_13),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_2),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_7),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_12),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_10),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_21),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_32),
.B(n_34),
.Y(n_43)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_24),
.Y(n_33)
);

INVx8_ASAP7_75t_L g55 ( 
.A(n_33),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_15),
.B(n_0),
.Y(n_34)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_21),
.Y(n_35)
);

INVx2_ASAP7_75t_SL g53 ( 
.A(n_35),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_15),
.Y(n_36)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_36),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_15),
.Y(n_37)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_37),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_16),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_38),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_21),
.B(n_0),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_39),
.B(n_41),
.Y(n_42)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_21),
.Y(n_40)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_40),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_16),
.B(n_0),
.Y(n_41)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_36),
.Y(n_46)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_46),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_38),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_47),
.B(n_19),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g49 ( 
.A1(n_39),
.A2(n_18),
.B1(n_30),
.B2(n_28),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_49),
.A2(n_51),
.B1(n_17),
.B2(n_23),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_L g51 ( 
.A1(n_32),
.A2(n_18),
.B1(n_30),
.B2(n_28),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_41),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_52),
.B(n_20),
.Y(n_71)
);

AND2x2_ASAP7_75t_L g54 ( 
.A(n_36),
.B(n_25),
.Y(n_54)
);

MAJIxp5_ASAP7_75t_L g59 ( 
.A(n_54),
.B(n_37),
.C(n_36),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_52),
.A2(n_33),
.B1(n_19),
.B2(n_27),
.Y(n_56)
);

INVxp67_ASAP7_75t_L g94 ( 
.A(n_56),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_44),
.B(n_34),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_57),
.B(n_60),
.Y(n_81)
);

AND2x2_ASAP7_75t_SL g58 ( 
.A(n_50),
.B(n_37),
.Y(n_58)
);

AND2x2_ASAP7_75t_L g95 ( 
.A(n_58),
.B(n_59),
.Y(n_95)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_55),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_44),
.B(n_26),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_61),
.B(n_66),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_55),
.A2(n_33),
.B1(n_27),
.B2(n_23),
.Y(n_62)
);

CKINVDCx16_ASAP7_75t_R g85 ( 
.A(n_62),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_63),
.B(n_80),
.Y(n_103)
);

OA22x2_ASAP7_75t_L g64 ( 
.A1(n_46),
.A2(n_35),
.B1(n_32),
.B2(n_40),
.Y(n_64)
);

AO21x1_ASAP7_75t_L g101 ( 
.A1(n_64),
.A2(n_65),
.B(n_75),
.Y(n_101)
);

OR2x4_ASAP7_75t_L g65 ( 
.A(n_49),
.B(n_37),
.Y(n_65)
);

INVxp67_ASAP7_75t_L g66 ( 
.A(n_43),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_47),
.B(n_29),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_67),
.B(n_72),
.Y(n_89)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_45),
.Y(n_69)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_69),
.Y(n_84)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_55),
.Y(n_70)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_70),
.Y(n_102)
);

OAI21xp33_ASAP7_75t_L g100 ( 
.A1(n_71),
.A2(n_17),
.B(n_31),
.Y(n_100)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_54),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_43),
.B(n_29),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_73),
.B(n_74),
.Y(n_90)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_45),
.Y(n_74)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_42),
.B(n_25),
.Y(n_75)
);

CKINVDCx14_ASAP7_75t_R g76 ( 
.A(n_42),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_76),
.B(n_77),
.Y(n_91)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_48),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_54),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_78),
.B(n_79),
.Y(n_99)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_54),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_72),
.A2(n_40),
.B1(n_35),
.B2(n_48),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_82),
.A2(n_93),
.B1(n_98),
.B2(n_92),
.Y(n_112)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_64),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_83),
.B(n_87),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_66),
.B(n_50),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_86),
.B(n_75),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_58),
.Y(n_87)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_64),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_92),
.B(n_96),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_78),
.A2(n_46),
.B1(n_53),
.B2(n_20),
.Y(n_93)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_64),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_71),
.B(n_26),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_97),
.B(n_100),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_65),
.A2(n_53),
.B1(n_20),
.B2(n_17),
.Y(n_98)
);

XOR2xp5_ASAP7_75t_L g106 ( 
.A(n_99),
.B(n_80),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_106),
.B(n_119),
.C(n_103),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_81),
.B(n_79),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_SL g127 ( 
.A(n_107),
.B(n_110),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_109),
.B(n_111),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_81),
.B(n_58),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_86),
.B(n_99),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_112),
.A2(n_91),
.B1(n_89),
.B2(n_82),
.Y(n_137)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_102),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_113),
.B(n_115),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_83),
.A2(n_59),
.B1(n_60),
.B2(n_75),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_114),
.A2(n_116),
.B1(n_53),
.B2(n_68),
.Y(n_142)
);

BUFx3_ASAP7_75t_L g115 ( 
.A(n_102),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_96),
.A2(n_85),
.B1(n_94),
.B2(n_101),
.Y(n_116)
);

INVx5_ASAP7_75t_L g117 ( 
.A(n_84),
.Y(n_117)
);

BUFx2_ASAP7_75t_L g125 ( 
.A(n_117),
.Y(n_125)
);

CKINVDCx16_ASAP7_75t_R g118 ( 
.A(n_88),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_118),
.B(n_120),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_L g119 ( 
.A(n_101),
.B(n_31),
.Y(n_119)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_88),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_90),
.B(n_70),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_SL g130 ( 
.A(n_121),
.B(n_91),
.Y(n_130)
);

CKINVDCx16_ASAP7_75t_R g122 ( 
.A(n_90),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_122),
.B(n_124),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_95),
.A2(n_101),
.B1(n_85),
.B2(n_98),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_123),
.A2(n_53),
.B1(n_69),
.B2(n_74),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_95),
.B(n_77),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_130),
.B(n_135),
.Y(n_148)
);

MAJx2_ASAP7_75t_L g150 ( 
.A(n_132),
.B(n_22),
.C(n_24),
.Y(n_150)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_108),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_133),
.B(n_134),
.Y(n_151)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_104),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_SL g135 ( 
.A(n_111),
.B(n_103),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_124),
.B(n_95),
.C(n_87),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_136),
.B(n_138),
.C(n_25),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_137),
.A2(n_142),
.B1(n_1),
.B2(n_2),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_106),
.B(n_89),
.C(n_93),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_L g139 ( 
.A1(n_109),
.A2(n_84),
.B(n_68),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_L g145 ( 
.A1(n_139),
.A2(n_141),
.B(n_115),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_140),
.B(n_1),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_L g141 ( 
.A1(n_120),
.A2(n_123),
.B(n_116),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_112),
.A2(n_119),
.B1(n_105),
.B2(n_113),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_143),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_L g164 ( 
.A(n_144),
.B(n_145),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_136),
.B(n_117),
.C(n_25),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_146),
.B(n_147),
.C(n_149),
.Y(n_167)
);

XOR2xp5_ASAP7_75t_L g147 ( 
.A(n_138),
.B(n_22),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_141),
.B(n_24),
.C(n_22),
.Y(n_149)
);

XNOR2x1_ASAP7_75t_L g162 ( 
.A(n_150),
.B(n_147),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_152),
.A2(n_135),
.B1(n_133),
.B2(n_127),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_134),
.B(n_1),
.Y(n_153)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_153),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_SL g169 ( 
.A1(n_154),
.A2(n_126),
.B(n_143),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_126),
.B(n_3),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_155),
.B(n_156),
.Y(n_168)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_128),
.Y(n_156)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_157),
.Y(n_160)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_125),
.Y(n_158)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_158),
.Y(n_161)
);

MAJx2_ASAP7_75t_L g173 ( 
.A(n_162),
.B(n_149),
.C(n_150),
.Y(n_173)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_163),
.Y(n_178)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_151),
.Y(n_165)
);

AOI21xp5_ASAP7_75t_L g175 ( 
.A1(n_165),
.A2(n_169),
.B(n_155),
.Y(n_175)
);

BUFx12_ASAP7_75t_L g166 ( 
.A(n_146),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_166),
.B(n_144),
.C(n_145),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_170),
.B(n_177),
.Y(n_184)
);

OAI22xp33_ASAP7_75t_L g171 ( 
.A1(n_160),
.A2(n_151),
.B1(n_129),
.B2(n_131),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_171),
.A2(n_166),
.B1(n_125),
.B2(n_6),
.Y(n_185)
);

XOR2xp5_ASAP7_75t_L g172 ( 
.A(n_167),
.B(n_132),
.Y(n_172)
);

XOR2xp5_ASAP7_75t_L g181 ( 
.A(n_172),
.B(n_173),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_L g174 ( 
.A1(n_167),
.A2(n_148),
.B(n_153),
.Y(n_174)
);

AOI21xp5_ASAP7_75t_L g180 ( 
.A1(n_174),
.A2(n_168),
.B(n_162),
.Y(n_180)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_175),
.Y(n_179)
);

O2A1O1Ixp33_ASAP7_75t_L g176 ( 
.A1(n_169),
.A2(n_139),
.B(n_157),
.C(n_142),
.Y(n_176)
);

OAI31xp33_ASAP7_75t_L g182 ( 
.A1(n_176),
.A2(n_159),
.A3(n_168),
.B(n_164),
.Y(n_182)
);

AOI21xp5_ASAP7_75t_L g177 ( 
.A1(n_164),
.A2(n_140),
.B(n_4),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_180),
.B(n_166),
.C(n_14),
.Y(n_188)
);

A2O1A1Ixp33_ASAP7_75t_L g186 ( 
.A1(n_182),
.A2(n_171),
.B(n_176),
.C(n_173),
.Y(n_186)
);

AOI21xp5_ASAP7_75t_L g183 ( 
.A1(n_178),
.A2(n_159),
.B(n_161),
.Y(n_183)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_183),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_185),
.B(n_179),
.Y(n_190)
);

AOI21xp5_ASAP7_75t_L g193 ( 
.A1(n_186),
.A2(n_187),
.B(n_5),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_188),
.B(n_181),
.C(n_182),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_SL g189 ( 
.A(n_184),
.B(n_13),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_189),
.B(n_190),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_191),
.B(n_192),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g192 ( 
.A(n_186),
.B(n_181),
.Y(n_192)
);

OAI321xp33_ASAP7_75t_L g196 ( 
.A1(n_193),
.A2(n_3),
.A3(n_7),
.B1(n_8),
.B2(n_9),
.C(n_10),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_SL g197 ( 
.A1(n_196),
.A2(n_194),
.B(n_8),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_197),
.B(n_198),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_195),
.B(n_192),
.C(n_7),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_199),
.B(n_8),
.Y(n_200)
);


endmodule