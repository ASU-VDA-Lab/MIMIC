module fake_jpeg_12566_n_567 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_567);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_567;

wire n_529;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_19;
wire n_182;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_547;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_384;
wire n_296;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_1),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_17),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_17),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_15),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_15),
.Y(n_26)
);

BUFx24_ASAP7_75t_L g27 ( 
.A(n_18),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

BUFx4f_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_17),
.Y(n_30)
);

BUFx8_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_5),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_7),
.B(n_4),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_3),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_13),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_7),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_6),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_16),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_14),
.Y(n_40)
);

CKINVDCx16_ASAP7_75t_R g41 ( 
.A(n_12),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_14),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_7),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_11),
.Y(n_44)
);

BUFx5_ASAP7_75t_L g45 ( 
.A(n_3),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_10),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_15),
.Y(n_47)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_18),
.Y(n_48)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_4),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_10),
.Y(n_50)
);

INVx8_ASAP7_75t_L g51 ( 
.A(n_8),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_8),
.Y(n_52)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_10),
.Y(n_53)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_31),
.Y(n_54)
);

INVx5_ASAP7_75t_L g109 ( 
.A(n_54),
.Y(n_109)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_49),
.Y(n_55)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_55),
.Y(n_114)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_43),
.Y(n_56)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_56),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_34),
.B(n_18),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_57),
.B(n_107),
.Y(n_111)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_30),
.Y(n_58)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_58),
.Y(n_123)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_49),
.Y(n_59)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_59),
.Y(n_119)
);

BUFx5_ASAP7_75t_L g60 ( 
.A(n_45),
.Y(n_60)
);

BUFx5_ASAP7_75t_L g125 ( 
.A(n_60),
.Y(n_125)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_20),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_61),
.Y(n_118)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_43),
.Y(n_62)
);

BUFx12f_ASAP7_75t_L g153 ( 
.A(n_62),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_20),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_63),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_20),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_64),
.Y(n_136)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_24),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g143 ( 
.A(n_65),
.Y(n_143)
);

CKINVDCx16_ASAP7_75t_R g66 ( 
.A(n_27),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_66),
.B(n_86),
.Y(n_120)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_30),
.Y(n_67)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_67),
.Y(n_137)
);

INVx11_ASAP7_75t_L g68 ( 
.A(n_27),
.Y(n_68)
);

INVx11_ASAP7_75t_L g110 ( 
.A(n_68),
.Y(n_110)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_47),
.Y(n_69)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_69),
.Y(n_163)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_27),
.Y(n_70)
);

BUFx2_ASAP7_75t_L g128 ( 
.A(n_70),
.Y(n_128)
);

INVx6_ASAP7_75t_L g71 ( 
.A(n_24),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g146 ( 
.A(n_71),
.Y(n_146)
);

BUFx12_ASAP7_75t_L g72 ( 
.A(n_27),
.Y(n_72)
);

BUFx4f_ASAP7_75t_SL g144 ( 
.A(n_72),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_24),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g149 ( 
.A(n_73),
.Y(n_149)
);

INVx8_ASAP7_75t_L g74 ( 
.A(n_45),
.Y(n_74)
);

BUFx2_ASAP7_75t_L g154 ( 
.A(n_74),
.Y(n_154)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_22),
.Y(n_75)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_75),
.Y(n_124)
);

INVx6_ASAP7_75t_L g76 ( 
.A(n_28),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g168 ( 
.A(n_76),
.Y(n_168)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_43),
.Y(n_77)
);

INVx3_ASAP7_75t_L g156 ( 
.A(n_77),
.Y(n_156)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_22),
.Y(n_78)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_78),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_23),
.B(n_16),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g140 ( 
.A(n_79),
.B(n_90),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_28),
.Y(n_80)
);

INVx6_ASAP7_75t_L g139 ( 
.A(n_80),
.Y(n_139)
);

INVx5_ASAP7_75t_L g81 ( 
.A(n_25),
.Y(n_81)
);

INVx5_ASAP7_75t_L g115 ( 
.A(n_81),
.Y(n_115)
);

INVx1_ASAP7_75t_SL g82 ( 
.A(n_43),
.Y(n_82)
);

INVx4_ASAP7_75t_SL g171 ( 
.A(n_82),
.Y(n_171)
);

BUFx4f_ASAP7_75t_L g83 ( 
.A(n_31),
.Y(n_83)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_83),
.Y(n_152)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_47),
.Y(n_84)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_84),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_28),
.Y(n_85)
);

INVx6_ASAP7_75t_L g158 ( 
.A(n_85),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_34),
.Y(n_86)
);

CKINVDCx16_ASAP7_75t_R g87 ( 
.A(n_25),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_87),
.B(n_91),
.Y(n_121)
);

INVx6_ASAP7_75t_L g88 ( 
.A(n_40),
.Y(n_88)
);

INVx3_ASAP7_75t_SL g122 ( 
.A(n_88),
.Y(n_122)
);

BUFx12f_ASAP7_75t_L g89 ( 
.A(n_31),
.Y(n_89)
);

INVx5_ASAP7_75t_L g164 ( 
.A(n_89),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_23),
.B(n_16),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_26),
.Y(n_91)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_29),
.Y(n_92)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_92),
.Y(n_155)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_25),
.Y(n_93)
);

INVx4_ASAP7_75t_L g116 ( 
.A(n_93),
.Y(n_116)
);

BUFx2_ASAP7_75t_R g94 ( 
.A(n_41),
.Y(n_94)
);

INVx13_ASAP7_75t_L g162 ( 
.A(n_94),
.Y(n_162)
);

INVx5_ASAP7_75t_L g95 ( 
.A(n_48),
.Y(n_95)
);

INVx4_ASAP7_75t_L g130 ( 
.A(n_95),
.Y(n_130)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_29),
.Y(n_96)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_96),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_26),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_97),
.B(n_100),
.Y(n_157)
);

BUFx12f_ASAP7_75t_L g98 ( 
.A(n_31),
.Y(n_98)
);

INVx4_ASAP7_75t_L g135 ( 
.A(n_98),
.Y(n_135)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_29),
.Y(n_99)
);

INVx4_ASAP7_75t_L g141 ( 
.A(n_99),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_39),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_40),
.Y(n_101)
);

INVx8_ASAP7_75t_L g117 ( 
.A(n_101),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_39),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_102),
.B(n_42),
.Y(n_159)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_48),
.Y(n_103)
);

INVx4_ASAP7_75t_L g148 ( 
.A(n_103),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_19),
.B(n_0),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_SL g150 ( 
.A(n_104),
.B(n_106),
.Y(n_150)
);

BUFx12_ASAP7_75t_L g105 ( 
.A(n_41),
.Y(n_105)
);

BUFx8_ASAP7_75t_L g170 ( 
.A(n_105),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_19),
.B(n_0),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_48),
.B(n_0),
.Y(n_107)
);

BUFx3_ASAP7_75t_L g108 ( 
.A(n_32),
.Y(n_108)
);

BUFx12f_ASAP7_75t_L g165 ( 
.A(n_108),
.Y(n_165)
);

A2O1A1Ixp33_ASAP7_75t_L g113 ( 
.A1(n_94),
.A2(n_105),
.B(n_68),
.C(n_46),
.Y(n_113)
);

OR2x2_ASAP7_75t_L g185 ( 
.A(n_113),
.B(n_77),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_61),
.A2(n_40),
.B1(n_52),
.B2(n_37),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_126),
.A2(n_33),
.B1(n_35),
.B2(n_46),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_93),
.B(n_38),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_127),
.B(n_132),
.Y(n_193)
);

CKINVDCx16_ASAP7_75t_R g129 ( 
.A(n_105),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_129),
.B(n_131),
.Y(n_176)
);

CKINVDCx16_ASAP7_75t_R g131 ( 
.A(n_72),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_103),
.B(n_38),
.Y(n_132)
);

INVx8_ASAP7_75t_L g133 ( 
.A(n_60),
.Y(n_133)
);

INVx5_ASAP7_75t_L g182 ( 
.A(n_133),
.Y(n_182)
);

AND2x2_ASAP7_75t_SL g138 ( 
.A(n_54),
.B(n_98),
.Y(n_138)
);

AND2x2_ASAP7_75t_L g200 ( 
.A(n_138),
.B(n_98),
.Y(n_200)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_70),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_145),
.B(n_159),
.Y(n_180)
);

BUFx5_ASAP7_75t_L g147 ( 
.A(n_72),
.Y(n_147)
);

BUFx3_ASAP7_75t_L g174 ( 
.A(n_147),
.Y(n_174)
);

INVx8_ASAP7_75t_L g151 ( 
.A(n_63),
.Y(n_151)
);

INVx4_ASAP7_75t_L g188 ( 
.A(n_151),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_SL g160 ( 
.A(n_54),
.B(n_42),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_SL g232 ( 
.A(n_160),
.B(n_161),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_82),
.B(n_37),
.Y(n_161)
);

INVx11_ASAP7_75t_L g166 ( 
.A(n_83),
.Y(n_166)
);

INVxp67_ASAP7_75t_L g177 ( 
.A(n_166),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_SL g167 ( 
.A(n_89),
.B(n_52),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_SL g234 ( 
.A(n_167),
.B(n_5),
.Y(n_234)
);

INVx11_ASAP7_75t_L g173 ( 
.A(n_83),
.Y(n_173)
);

CKINVDCx16_ASAP7_75t_R g226 ( 
.A(n_173),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_111),
.B(n_36),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_SL g256 ( 
.A(n_175),
.B(n_183),
.Y(n_256)
);

AOI22xp33_ASAP7_75t_SL g178 ( 
.A1(n_133),
.A2(n_53),
.B1(n_51),
.B2(n_89),
.Y(n_178)
);

INVxp67_ASAP7_75t_L g242 ( 
.A(n_178),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_150),
.A2(n_65),
.B1(n_76),
.B2(n_71),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_179),
.A2(n_222),
.B1(n_227),
.B2(n_209),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_113),
.B(n_44),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_181),
.B(n_184),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_140),
.B(n_44),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_123),
.B(n_36),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_SL g287 ( 
.A1(n_185),
.A2(n_220),
.B(n_125),
.Y(n_287)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_137),
.Y(n_186)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_186),
.Y(n_250)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_163),
.Y(n_187)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_187),
.Y(n_254)
);

INVx1_ASAP7_75t_SL g189 ( 
.A(n_138),
.Y(n_189)
);

INVx1_ASAP7_75t_SL g247 ( 
.A(n_189),
.Y(n_247)
);

AOI22xp33_ASAP7_75t_L g190 ( 
.A1(n_117),
.A2(n_88),
.B1(n_101),
.B2(n_64),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g237 ( 
.A1(n_190),
.A2(n_191),
.B1(n_202),
.B2(n_213),
.Y(n_237)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_141),
.Y(n_192)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_192),
.Y(n_270)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_141),
.Y(n_194)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_194),
.Y(n_276)
);

BUFx3_ASAP7_75t_L g195 ( 
.A(n_153),
.Y(n_195)
);

INVx4_ASAP7_75t_L g263 ( 
.A(n_195),
.Y(n_263)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_155),
.Y(n_196)
);

INVx2_ASAP7_75t_L g281 ( 
.A(n_196),
.Y(n_281)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_169),
.Y(n_197)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_197),
.Y(n_286)
);

INVx2_ASAP7_75t_SL g198 ( 
.A(n_166),
.Y(n_198)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_198),
.Y(n_261)
);

BUFx6f_ASAP7_75t_L g199 ( 
.A(n_134),
.Y(n_199)
);

BUFx6f_ASAP7_75t_L g240 ( 
.A(n_199),
.Y(n_240)
);

AND2x2_ASAP7_75t_L g251 ( 
.A(n_200),
.B(n_209),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_157),
.B(n_56),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g275 ( 
.A(n_201),
.B(n_203),
.Y(n_275)
);

AOI22xp33_ASAP7_75t_L g202 ( 
.A1(n_117),
.A2(n_85),
.B1(n_80),
.B2(n_73),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_120),
.B(n_95),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_121),
.B(n_81),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_204),
.B(n_206),
.Y(n_241)
);

INVx4_ASAP7_75t_L g205 ( 
.A(n_135),
.Y(n_205)
);

BUFx2_ASAP7_75t_L g239 ( 
.A(n_205),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_172),
.B(n_62),
.Y(n_206)
);

INVx4_ASAP7_75t_L g207 ( 
.A(n_135),
.Y(n_207)
);

BUFx2_ASAP7_75t_L g285 ( 
.A(n_207),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_124),
.A2(n_108),
.B1(n_53),
.B2(n_51),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_208),
.A2(n_231),
.B1(n_149),
.B2(n_118),
.Y(n_267)
);

AND2x2_ASAP7_75t_SL g209 ( 
.A(n_114),
.B(n_32),
.Y(n_209)
);

BUFx6f_ASAP7_75t_L g210 ( 
.A(n_134),
.Y(n_210)
);

INVx6_ASAP7_75t_L g273 ( 
.A(n_210),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_119),
.B(n_35),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_211),
.B(n_218),
.Y(n_259)
);

AND2x2_ASAP7_75t_L g212 ( 
.A(n_171),
.B(n_32),
.Y(n_212)
);

AND2x2_ASAP7_75t_L g266 ( 
.A(n_212),
.B(n_224),
.Y(n_266)
);

AOI22xp33_ASAP7_75t_L g213 ( 
.A1(n_151),
.A2(n_33),
.B1(n_21),
.B2(n_51),
.Y(n_213)
);

AOI22xp33_ASAP7_75t_SL g214 ( 
.A1(n_154),
.A2(n_53),
.B1(n_74),
.B2(n_21),
.Y(n_214)
);

AOI22xp33_ASAP7_75t_SL g255 ( 
.A1(n_214),
.A2(n_128),
.B1(n_110),
.B2(n_153),
.Y(n_255)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_122),
.Y(n_215)
);

HB1xp67_ASAP7_75t_L g249 ( 
.A(n_215),
.Y(n_249)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_152),
.Y(n_216)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_216),
.Y(n_271)
);

AOI22xp33_ASAP7_75t_L g217 ( 
.A1(n_139),
.A2(n_50),
.B1(n_29),
.B2(n_32),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_L g252 ( 
.A1(n_217),
.A2(n_221),
.B1(n_128),
.B2(n_164),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_173),
.Y(n_218)
);

INVx4_ASAP7_75t_L g219 ( 
.A(n_165),
.Y(n_219)
);

INVx4_ASAP7_75t_L g290 ( 
.A(n_219),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_154),
.A2(n_50),
.B1(n_32),
.B2(n_3),
.Y(n_220)
);

AOI22xp33_ASAP7_75t_L g221 ( 
.A1(n_139),
.A2(n_50),
.B1(n_2),
.B2(n_3),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_142),
.A2(n_1),
.B1(n_2),
.B2(n_4),
.Y(n_222)
);

BUFx6f_ASAP7_75t_L g223 ( 
.A(n_136),
.Y(n_223)
);

INVx3_ASAP7_75t_L g238 ( 
.A(n_223),
.Y(n_238)
);

AND2x2_ASAP7_75t_L g224 ( 
.A(n_171),
.B(n_1),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_116),
.B(n_1),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_225),
.B(n_234),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_122),
.A2(n_14),
.B1(n_6),
.B2(n_7),
.Y(n_227)
);

INVx4_ASAP7_75t_L g228 ( 
.A(n_165),
.Y(n_228)
);

INVx3_ASAP7_75t_L g265 ( 
.A(n_228),
.Y(n_265)
);

INVx6_ASAP7_75t_L g229 ( 
.A(n_136),
.Y(n_229)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_229),
.Y(n_278)
);

INVx4_ASAP7_75t_L g230 ( 
.A(n_165),
.Y(n_230)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_230),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_158),
.A2(n_5),
.B1(n_6),
.B2(n_8),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_158),
.B(n_5),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_233),
.B(n_8),
.Y(n_248)
);

INVx4_ASAP7_75t_L g235 ( 
.A(n_109),
.Y(n_235)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_235),
.Y(n_274)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_112),
.Y(n_236)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_236),
.Y(n_280)
);

AND2x2_ASAP7_75t_L g307 ( 
.A(n_243),
.B(n_245),
.Y(n_307)
);

O2A1O1Ixp33_ASAP7_75t_L g245 ( 
.A1(n_181),
.A2(n_110),
.B(n_162),
.C(n_145),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_180),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_246),
.B(n_257),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_SL g301 ( 
.A(n_248),
.B(n_258),
.Y(n_301)
);

AND2x2_ASAP7_75t_L g320 ( 
.A(n_252),
.B(n_264),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_193),
.B(n_143),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_253),
.B(n_269),
.Y(n_293)
);

AOI22xp33_ASAP7_75t_SL g334 ( 
.A1(n_255),
.A2(n_198),
.B1(n_174),
.B2(n_235),
.Y(n_334)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_184),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g258 ( 
.A(n_189),
.B(n_156),
.Y(n_258)
);

BUFx12_ASAP7_75t_L g260 ( 
.A(n_219),
.Y(n_260)
);

INVx13_ASAP7_75t_L g297 ( 
.A(n_260),
.Y(n_297)
);

OAI22xp33_ASAP7_75t_SL g262 ( 
.A1(n_185),
.A2(n_143),
.B1(n_168),
.B2(n_146),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_262),
.A2(n_267),
.B1(n_291),
.B2(n_200),
.Y(n_304)
);

OA22x2_ASAP7_75t_L g264 ( 
.A1(n_208),
.A2(n_146),
.B1(n_168),
.B2(n_118),
.Y(n_264)
);

AOI22xp33_ASAP7_75t_L g268 ( 
.A1(n_227),
.A2(n_148),
.B1(n_116),
.B2(n_149),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_SL g330 ( 
.A1(n_268),
.A2(n_198),
.B1(n_215),
.B2(n_177),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_233),
.B(n_148),
.Y(n_269)
);

INVx2_ASAP7_75t_SL g277 ( 
.A(n_182),
.Y(n_277)
);

INVx2_ASAP7_75t_L g296 ( 
.A(n_277),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_176),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_282),
.B(n_284),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_209),
.B(n_162),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_SL g328 ( 
.A(n_283),
.B(n_170),
.Y(n_328)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_212),
.Y(n_284)
);

OR2x2_ASAP7_75t_L g298 ( 
.A(n_287),
.B(n_182),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_232),
.B(n_130),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_SL g336 ( 
.A(n_288),
.B(n_144),
.Y(n_336)
);

INVx13_ASAP7_75t_L g289 ( 
.A(n_226),
.Y(n_289)
);

INVx13_ASAP7_75t_L g303 ( 
.A(n_289),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_L g291 ( 
.A1(n_191),
.A2(n_115),
.B1(n_130),
.B2(n_170),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g292 ( 
.A(n_249),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_292),
.B(n_306),
.Y(n_350)
);

BUFx10_ASAP7_75t_L g294 ( 
.A(n_289),
.Y(n_294)
);

INVx2_ASAP7_75t_SL g379 ( 
.A(n_294),
.Y(n_379)
);

OAI21xp5_ASAP7_75t_SL g371 ( 
.A1(n_298),
.A2(n_177),
.B(n_144),
.Y(n_371)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_261),
.Y(n_299)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_299),
.Y(n_341)
);

INVxp67_ASAP7_75t_L g300 ( 
.A(n_275),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_SL g351 ( 
.A(n_300),
.B(n_309),
.Y(n_351)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_261),
.Y(n_302)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_302),
.Y(n_360)
);

OAI22xp5_ASAP7_75t_L g349 ( 
.A1(n_304),
.A2(n_339),
.B1(n_277),
.B2(n_264),
.Y(n_349)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_281),
.Y(n_305)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_305),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_248),
.B(n_224),
.Y(n_306)
);

INVx13_ASAP7_75t_L g308 ( 
.A(n_260),
.Y(n_308)
);

INVxp67_ASAP7_75t_L g353 ( 
.A(n_308),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_259),
.B(n_236),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_281),
.Y(n_310)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_310),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_256),
.B(n_192),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_311),
.B(n_315),
.Y(n_356)
);

INVxp67_ASAP7_75t_L g312 ( 
.A(n_241),
.Y(n_312)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_312),
.Y(n_370)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_286),
.Y(n_313)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_313),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_269),
.B(n_224),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_286),
.Y(n_316)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_316),
.Y(n_346)
);

INVxp67_ASAP7_75t_L g317 ( 
.A(n_251),
.Y(n_317)
);

BUFx2_ASAP7_75t_L g345 ( 
.A(n_317),
.Y(n_345)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_280),
.Y(n_318)
);

INVx2_ASAP7_75t_L g373 ( 
.A(n_318),
.Y(n_373)
);

OAI22xp33_ASAP7_75t_SL g319 ( 
.A1(n_243),
.A2(n_220),
.B1(n_231),
.B2(n_188),
.Y(n_319)
);

AOI22xp5_ASAP7_75t_L g342 ( 
.A1(n_319),
.A2(n_242),
.B1(n_237),
.B2(n_251),
.Y(n_342)
);

INVx13_ASAP7_75t_L g321 ( 
.A(n_260),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g355 ( 
.A(n_321),
.Y(n_355)
);

INVx2_ASAP7_75t_L g322 ( 
.A(n_278),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_322),
.B(n_323),
.Y(n_361)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_271),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_253),
.B(n_194),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_324),
.B(n_326),
.Y(n_366)
);

AOI21xp5_ASAP7_75t_L g325 ( 
.A1(n_287),
.A2(n_200),
.B(n_212),
.Y(n_325)
);

AOI21xp5_ASAP7_75t_L g381 ( 
.A1(n_325),
.A2(n_298),
.B(n_307),
.Y(n_381)
);

INVx1_ASAP7_75t_SL g326 ( 
.A(n_239),
.Y(n_326)
);

INVx4_ASAP7_75t_L g327 ( 
.A(n_273),
.Y(n_327)
);

AOI22xp33_ASAP7_75t_SL g358 ( 
.A1(n_327),
.A2(n_333),
.B1(n_334),
.B2(n_336),
.Y(n_358)
);

XNOR2xp5_ASAP7_75t_L g343 ( 
.A(n_328),
.B(n_258),
.Y(n_343)
);

AND2x6_ASAP7_75t_L g329 ( 
.A(n_244),
.B(n_245),
.Y(n_329)
);

AOI32xp33_ASAP7_75t_L g357 ( 
.A1(n_329),
.A2(n_170),
.A3(n_279),
.B1(n_254),
.B2(n_153),
.Y(n_357)
);

AOI22xp33_ASAP7_75t_L g374 ( 
.A1(n_330),
.A2(n_337),
.B1(n_238),
.B2(n_285),
.Y(n_374)
);

INVxp67_ASAP7_75t_L g331 ( 
.A(n_251),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_331),
.B(n_332),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_244),
.B(n_222),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_270),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g335 ( 
.A(n_250),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g359 ( 
.A(n_335),
.Y(n_359)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_270),
.Y(n_337)
);

OR2x2_ASAP7_75t_L g338 ( 
.A(n_283),
.B(n_207),
.Y(n_338)
);

OAI21xp5_ASAP7_75t_L g365 ( 
.A1(n_338),
.A2(n_325),
.B(n_328),
.Y(n_365)
);

AOI22xp33_ASAP7_75t_L g339 ( 
.A1(n_267),
.A2(n_188),
.B1(n_229),
.B2(n_196),
.Y(n_339)
);

INVx13_ASAP7_75t_L g340 ( 
.A(n_263),
.Y(n_340)
);

CKINVDCx20_ASAP7_75t_R g377 ( 
.A(n_340),
.Y(n_377)
);

OR2x2_ASAP7_75t_L g405 ( 
.A(n_342),
.B(n_371),
.Y(n_405)
);

XOR2xp5_ASAP7_75t_L g407 ( 
.A(n_343),
.B(n_365),
.Y(n_407)
);

OAI22xp5_ASAP7_75t_SL g344 ( 
.A1(n_304),
.A2(n_242),
.B1(n_264),
.B2(n_247),
.Y(n_344)
);

AOI22xp5_ASAP7_75t_L g385 ( 
.A1(n_344),
.A2(n_349),
.B1(n_375),
.B2(n_380),
.Y(n_385)
);

XNOR2xp5_ASAP7_75t_L g347 ( 
.A(n_301),
.B(n_247),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_L g387 ( 
.A(n_347),
.B(n_348),
.C(n_352),
.Y(n_387)
);

XNOR2xp5_ASAP7_75t_L g348 ( 
.A(n_301),
.B(n_266),
.Y(n_348)
);

XNOR2xp5_ASAP7_75t_L g352 ( 
.A(n_293),
.B(n_266),
.Y(n_352)
);

AOI22xp5_ASAP7_75t_L g354 ( 
.A1(n_307),
.A2(n_266),
.B1(n_264),
.B2(n_277),
.Y(n_354)
);

OAI22xp5_ASAP7_75t_SL g399 ( 
.A1(n_354),
.A2(n_363),
.B1(n_383),
.B2(n_342),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_SL g386 ( 
.A(n_357),
.B(n_378),
.Y(n_386)
);

OAI32xp33_ASAP7_75t_L g362 ( 
.A1(n_332),
.A2(n_197),
.A3(n_278),
.B1(n_274),
.B2(n_276),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_362),
.B(n_324),
.Y(n_392)
);

AOI22xp5_ASAP7_75t_L g363 ( 
.A1(n_307),
.A2(n_238),
.B1(n_273),
.B2(n_240),
.Y(n_363)
);

MAJIxp5_ASAP7_75t_L g364 ( 
.A(n_338),
.B(n_272),
.C(n_276),
.Y(n_364)
);

MAJIxp5_ASAP7_75t_L g391 ( 
.A(n_364),
.B(n_382),
.C(n_338),
.Y(n_391)
);

OAI21xp5_ASAP7_75t_L g368 ( 
.A1(n_298),
.A2(n_265),
.B(n_285),
.Y(n_368)
);

OAI21xp5_ASAP7_75t_L g394 ( 
.A1(n_368),
.A2(n_381),
.B(n_294),
.Y(n_394)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_374),
.Y(n_388)
);

OAI22xp5_ASAP7_75t_L g375 ( 
.A1(n_295),
.A2(n_210),
.B1(n_223),
.B2(n_199),
.Y(n_375)
);

CKINVDCx20_ASAP7_75t_R g378 ( 
.A(n_294),
.Y(n_378)
);

OAI22xp5_ASAP7_75t_SL g380 ( 
.A1(n_293),
.A2(n_240),
.B1(n_265),
.B2(n_239),
.Y(n_380)
);

XNOR2xp5_ASAP7_75t_L g382 ( 
.A(n_315),
.B(n_290),
.Y(n_382)
);

AOI22xp5_ASAP7_75t_L g383 ( 
.A1(n_320),
.A2(n_290),
.B1(n_263),
.B2(n_205),
.Y(n_383)
);

AOI22x1_ASAP7_75t_L g384 ( 
.A1(n_344),
.A2(n_320),
.B1(n_329),
.B2(n_330),
.Y(n_384)
);

OAI22xp5_ASAP7_75t_L g430 ( 
.A1(n_384),
.A2(n_389),
.B1(n_392),
.B2(n_383),
.Y(n_430)
);

AOI22xp5_ASAP7_75t_L g389 ( 
.A1(n_376),
.A2(n_320),
.B1(n_302),
.B2(n_299),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_361),
.Y(n_390)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_390),
.Y(n_429)
);

XNOR2xp5_ASAP7_75t_L g428 ( 
.A(n_391),
.B(n_414),
.Y(n_428)
);

MAJIxp5_ASAP7_75t_L g393 ( 
.A(n_365),
.B(n_352),
.C(n_348),
.Y(n_393)
);

MAJIxp5_ASAP7_75t_L g441 ( 
.A(n_393),
.B(n_404),
.C(n_408),
.Y(n_441)
);

OAI21xp5_ASAP7_75t_L g434 ( 
.A1(n_394),
.A2(n_358),
.B(n_353),
.Y(n_434)
);

OAI21xp5_ASAP7_75t_L g395 ( 
.A1(n_381),
.A2(n_336),
.B(n_314),
.Y(n_395)
);

INVxp67_ASAP7_75t_L g422 ( 
.A(n_395),
.Y(n_422)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_361),
.Y(n_396)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_396),
.Y(n_438)
);

A2O1A1O1Ixp25_ASAP7_75t_L g397 ( 
.A1(n_376),
.A2(n_306),
.B(n_309),
.C(n_311),
.D(n_294),
.Y(n_397)
);

MAJIxp5_ASAP7_75t_SL g423 ( 
.A(n_397),
.B(n_364),
.C(n_368),
.Y(n_423)
);

NOR2xp33_ASAP7_75t_L g398 ( 
.A(n_359),
.B(n_335),
.Y(n_398)
);

NOR2xp33_ASAP7_75t_SL g424 ( 
.A(n_398),
.B(n_415),
.Y(n_424)
);

AOI22xp5_ASAP7_75t_L g447 ( 
.A1(n_399),
.A2(n_401),
.B1(n_403),
.B2(n_420),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_350),
.B(n_292),
.Y(n_400)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_400),
.Y(n_446)
);

OAI22xp5_ASAP7_75t_SL g401 ( 
.A1(n_354),
.A2(n_322),
.B1(n_296),
.B2(n_323),
.Y(n_401)
);

OAI21xp5_ASAP7_75t_L g402 ( 
.A1(n_371),
.A2(n_294),
.B(n_318),
.Y(n_402)
);

INVxp67_ASAP7_75t_L g448 ( 
.A(n_402),
.Y(n_448)
);

OAI22xp5_ASAP7_75t_SL g403 ( 
.A1(n_350),
.A2(n_296),
.B1(n_327),
.B2(n_305),
.Y(n_403)
);

MAJIxp5_ASAP7_75t_L g404 ( 
.A(n_343),
.B(n_337),
.C(n_333),
.Y(n_404)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_373),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_406),
.B(n_410),
.Y(n_432)
);

XOR2xp5_ASAP7_75t_L g408 ( 
.A(n_382),
.B(n_316),
.Y(n_408)
);

CKINVDCx14_ASAP7_75t_R g409 ( 
.A(n_351),
.Y(n_409)
);

NOR2xp33_ASAP7_75t_L g427 ( 
.A(n_409),
.B(n_345),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_366),
.B(n_313),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_366),
.B(n_310),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_411),
.B(n_412),
.Y(n_443)
);

INVx2_ASAP7_75t_L g412 ( 
.A(n_379),
.Y(n_412)
);

INVx13_ASAP7_75t_L g413 ( 
.A(n_353),
.Y(n_413)
);

CKINVDCx20_ASAP7_75t_R g437 ( 
.A(n_413),
.Y(n_437)
);

XOR2xp5_ASAP7_75t_L g414 ( 
.A(n_347),
.B(n_303),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_SL g415 ( 
.A(n_370),
.B(n_326),
.Y(n_415)
);

NOR2xp33_ASAP7_75t_L g416 ( 
.A(n_356),
.B(n_195),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_SL g425 ( 
.A(n_416),
.B(n_417),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_SL g417 ( 
.A(n_356),
.B(n_230),
.Y(n_417)
);

NOR2xp33_ASAP7_75t_L g418 ( 
.A(n_355),
.B(n_228),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_SL g450 ( 
.A(n_418),
.B(n_419),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_SL g419 ( 
.A(n_345),
.B(n_303),
.Y(n_419)
);

OAI22xp5_ASAP7_75t_SL g420 ( 
.A1(n_363),
.A2(n_303),
.B1(n_321),
.B2(n_308),
.Y(n_420)
);

OAI22xp5_ASAP7_75t_SL g421 ( 
.A1(n_405),
.A2(n_392),
.B1(n_389),
.B2(n_385),
.Y(n_421)
);

AOI22xp5_ASAP7_75t_L g466 ( 
.A1(n_421),
.A2(n_430),
.B1(n_452),
.B2(n_388),
.Y(n_466)
);

HB1xp67_ASAP7_75t_L g457 ( 
.A(n_423),
.Y(n_457)
);

CKINVDCx16_ASAP7_75t_R g426 ( 
.A(n_400),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_SL g458 ( 
.A(n_426),
.B(n_435),
.Y(n_458)
);

NAND3xp33_ASAP7_75t_L g473 ( 
.A(n_427),
.B(n_433),
.C(n_444),
.Y(n_473)
);

XNOR2xp5_ASAP7_75t_L g431 ( 
.A(n_387),
.B(n_341),
.Y(n_431)
);

XOR2xp5_ASAP7_75t_L g481 ( 
.A(n_431),
.B(n_440),
.Y(n_481)
);

NOR2xp33_ASAP7_75t_L g433 ( 
.A(n_404),
.B(n_360),
.Y(n_433)
);

NOR2xp33_ASAP7_75t_L g476 ( 
.A(n_434),
.B(n_439),
.Y(n_476)
);

CKINVDCx16_ASAP7_75t_R g435 ( 
.A(n_410),
.Y(n_435)
);

INVx8_ASAP7_75t_L g436 ( 
.A(n_413),
.Y(n_436)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_436),
.Y(n_454)
);

OAI21xp5_ASAP7_75t_L g439 ( 
.A1(n_405),
.A2(n_380),
.B(n_346),
.Y(n_439)
);

XNOR2xp5_ASAP7_75t_L g440 ( 
.A(n_387),
.B(n_372),
.Y(n_440)
);

OAI21xp5_ASAP7_75t_L g442 ( 
.A1(n_394),
.A2(n_346),
.B(n_367),
.Y(n_442)
);

HB1xp67_ASAP7_75t_L g474 ( 
.A(n_442),
.Y(n_474)
);

NOR2xp33_ASAP7_75t_L g444 ( 
.A(n_395),
.B(n_377),
.Y(n_444)
);

MAJx2_ASAP7_75t_L g445 ( 
.A(n_393),
.B(n_391),
.C(n_407),
.Y(n_445)
);

XNOR2xp5_ASAP7_75t_L g459 ( 
.A(n_445),
.B(n_451),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_403),
.B(n_362),
.Y(n_449)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_449),
.Y(n_460)
);

OAI21xp5_ASAP7_75t_L g451 ( 
.A1(n_402),
.A2(n_369),
.B(n_379),
.Y(n_451)
);

OAI22xp5_ASAP7_75t_SL g452 ( 
.A1(n_385),
.A2(n_373),
.B1(n_379),
.B2(n_340),
.Y(n_452)
);

OAI21xp5_ASAP7_75t_SL g453 ( 
.A1(n_386),
.A2(n_321),
.B(n_308),
.Y(n_453)
);

XNOR2xp5_ASAP7_75t_L g463 ( 
.A(n_453),
.B(n_414),
.Y(n_463)
);

MAJIxp5_ASAP7_75t_L g455 ( 
.A(n_441),
.B(n_407),
.C(n_408),
.Y(n_455)
);

MAJIxp5_ASAP7_75t_L g484 ( 
.A(n_455),
.B(n_468),
.C(n_479),
.Y(n_484)
);

OAI22x1_ASAP7_75t_SL g456 ( 
.A1(n_447),
.A2(n_384),
.B1(n_396),
.B2(n_390),
.Y(n_456)
);

AOI22xp5_ASAP7_75t_L g482 ( 
.A1(n_456),
.A2(n_448),
.B1(n_438),
.B2(n_429),
.Y(n_482)
);

BUFx24_ASAP7_75t_SL g461 ( 
.A(n_424),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_SL g500 ( 
.A(n_461),
.B(n_469),
.Y(n_500)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_446),
.Y(n_462)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_462),
.Y(n_491)
);

INVx1_ASAP7_75t_SL g483 ( 
.A(n_463),
.Y(n_483)
);

AOI22xp5_ASAP7_75t_L g464 ( 
.A1(n_421),
.A2(n_399),
.B1(n_401),
.B2(n_384),
.Y(n_464)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_464),
.Y(n_495)
);

OAI22xp5_ASAP7_75t_SL g465 ( 
.A1(n_447),
.A2(n_388),
.B1(n_411),
.B2(n_397),
.Y(n_465)
);

HB1xp67_ASAP7_75t_L g487 ( 
.A(n_465),
.Y(n_487)
);

HB1xp67_ASAP7_75t_L g490 ( 
.A(n_466),
.Y(n_490)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_446),
.Y(n_467)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_467),
.Y(n_497)
);

MAJIxp5_ASAP7_75t_L g468 ( 
.A(n_441),
.B(n_406),
.C(n_420),
.Y(n_468)
);

CKINVDCx20_ASAP7_75t_R g469 ( 
.A(n_432),
.Y(n_469)
);

OAI22xp5_ASAP7_75t_SL g470 ( 
.A1(n_449),
.A2(n_412),
.B1(n_340),
.B2(n_174),
.Y(n_470)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_470),
.Y(n_499)
);

XNOR2xp5_ASAP7_75t_L g471 ( 
.A(n_431),
.B(n_297),
.Y(n_471)
);

XOR2xp5_ASAP7_75t_L g485 ( 
.A(n_471),
.B(n_472),
.Y(n_485)
);

XNOR2xp5_ASAP7_75t_L g472 ( 
.A(n_440),
.B(n_428),
.Y(n_472)
);

BUFx24_ASAP7_75t_SL g475 ( 
.A(n_422),
.Y(n_475)
);

CKINVDCx20_ASAP7_75t_R g489 ( 
.A(n_475),
.Y(n_489)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_432),
.Y(n_477)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_477),
.Y(n_503)
);

CKINVDCx20_ASAP7_75t_R g478 ( 
.A(n_443),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_L g498 ( 
.A(n_478),
.B(n_480),
.Y(n_498)
);

MAJIxp5_ASAP7_75t_L g479 ( 
.A(n_445),
.B(n_297),
.C(n_11),
.Y(n_479)
);

AOI22xp5_ASAP7_75t_L g480 ( 
.A1(n_439),
.A2(n_297),
.B1(n_11),
.B2(n_12),
.Y(n_480)
);

OAI22xp5_ASAP7_75t_SL g506 ( 
.A1(n_482),
.A2(n_496),
.B1(n_502),
.B2(n_480),
.Y(n_506)
);

CKINVDCx16_ASAP7_75t_R g486 ( 
.A(n_474),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_SL g517 ( 
.A(n_486),
.B(n_488),
.Y(n_517)
);

MAJIxp5_ASAP7_75t_L g488 ( 
.A(n_472),
.B(n_428),
.C(n_423),
.Y(n_488)
);

XOR2xp5_ASAP7_75t_L g492 ( 
.A(n_459),
.B(n_422),
.Y(n_492)
);

XNOR2xp5_ASAP7_75t_SL g513 ( 
.A(n_492),
.B(n_504),
.Y(n_513)
);

MAJIxp5_ASAP7_75t_L g493 ( 
.A(n_468),
.B(n_448),
.C(n_442),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_SL g521 ( 
.A(n_493),
.B(n_501),
.Y(n_521)
);

OAI21xp5_ASAP7_75t_SL g494 ( 
.A1(n_476),
.A2(n_429),
.B(n_438),
.Y(n_494)
);

AOI21xp5_ASAP7_75t_L g511 ( 
.A1(n_494),
.A2(n_437),
.B(n_425),
.Y(n_511)
);

AOI22xp5_ASAP7_75t_L g496 ( 
.A1(n_460),
.A2(n_456),
.B1(n_434),
.B2(n_457),
.Y(n_496)
);

MAJIxp5_ASAP7_75t_L g501 ( 
.A(n_481),
.B(n_451),
.C(n_453),
.Y(n_501)
);

AOI22xp5_ASAP7_75t_L g502 ( 
.A1(n_464),
.A2(n_452),
.B1(n_443),
.B2(n_437),
.Y(n_502)
);

XOR2xp5_ASAP7_75t_L g504 ( 
.A(n_459),
.B(n_450),
.Y(n_504)
);

MAJIxp5_ASAP7_75t_L g505 ( 
.A(n_484),
.B(n_455),
.C(n_481),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_SL g531 ( 
.A(n_505),
.B(n_509),
.Y(n_531)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_506),
.Y(n_523)
);

AOI22xp33_ASAP7_75t_SL g507 ( 
.A1(n_499),
.A2(n_487),
.B1(n_490),
.B2(n_495),
.Y(n_507)
);

OAI22xp5_ASAP7_75t_L g527 ( 
.A1(n_507),
.A2(n_520),
.B1(n_496),
.B2(n_482),
.Y(n_527)
);

CKINVDCx20_ASAP7_75t_R g508 ( 
.A(n_498),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_L g537 ( 
.A(n_508),
.B(n_516),
.Y(n_537)
);

MAJIxp5_ASAP7_75t_L g509 ( 
.A(n_484),
.B(n_471),
.C(n_463),
.Y(n_509)
);

MAJIxp5_ASAP7_75t_L g510 ( 
.A(n_493),
.B(n_479),
.C(n_458),
.Y(n_510)
);

MAJIxp5_ASAP7_75t_L g526 ( 
.A(n_510),
.B(n_485),
.C(n_492),
.Y(n_526)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_511),
.Y(n_536)
);

NOR2xp33_ASAP7_75t_L g512 ( 
.A(n_489),
.B(n_473),
.Y(n_512)
);

NOR2xp33_ASAP7_75t_SL g535 ( 
.A(n_512),
.B(n_514),
.Y(n_535)
);

NOR2xp33_ASAP7_75t_L g514 ( 
.A(n_500),
.B(n_454),
.Y(n_514)
);

NOR2xp33_ASAP7_75t_SL g515 ( 
.A(n_488),
.B(n_436),
.Y(n_515)
);

NOR2xp33_ASAP7_75t_L g524 ( 
.A(n_515),
.B(n_522),
.Y(n_524)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_498),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_L g518 ( 
.A(n_494),
.B(n_9),
.Y(n_518)
);

XNOR2xp5_ASAP7_75t_L g534 ( 
.A(n_518),
.B(n_519),
.Y(n_534)
);

OAI22xp5_ASAP7_75t_SL g519 ( 
.A1(n_495),
.A2(n_9),
.B1(n_11),
.B2(n_12),
.Y(n_519)
);

AOI22xp5_ASAP7_75t_SL g520 ( 
.A1(n_501),
.A2(n_9),
.B1(n_12),
.B2(n_13),
.Y(n_520)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_491),
.Y(n_522)
);

NOR2xp33_ASAP7_75t_L g525 ( 
.A(n_517),
.B(n_504),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_L g545 ( 
.A(n_525),
.B(n_526),
.Y(n_545)
);

AOI22xp5_ASAP7_75t_L g542 ( 
.A1(n_527),
.A2(n_530),
.B1(n_519),
.B2(n_518),
.Y(n_542)
);

MAJIxp5_ASAP7_75t_L g528 ( 
.A(n_521),
.B(n_485),
.C(n_483),
.Y(n_528)
);

MAJIxp5_ASAP7_75t_L g538 ( 
.A(n_528),
.B(n_532),
.C(n_510),
.Y(n_538)
);

AND2x2_ASAP7_75t_L g529 ( 
.A(n_509),
.B(n_483),
.Y(n_529)
);

INVxp67_ASAP7_75t_L g541 ( 
.A(n_529),
.Y(n_541)
);

BUFx10_ASAP7_75t_L g530 ( 
.A(n_511),
.Y(n_530)
);

MAJIxp5_ASAP7_75t_L g532 ( 
.A(n_505),
.B(n_502),
.C(n_503),
.Y(n_532)
);

OAI21xp5_ASAP7_75t_SL g533 ( 
.A1(n_516),
.A2(n_497),
.B(n_9),
.Y(n_533)
);

XNOR2xp5_ASAP7_75t_L g543 ( 
.A(n_533),
.B(n_522),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_L g549 ( 
.A(n_538),
.B(n_539),
.Y(n_549)
);

MAJIxp5_ASAP7_75t_L g539 ( 
.A(n_531),
.B(n_513),
.C(n_506),
.Y(n_539)
);

MAJIxp5_ASAP7_75t_L g540 ( 
.A(n_532),
.B(n_513),
.C(n_508),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_L g555 ( 
.A(n_540),
.B(n_542),
.Y(n_555)
);

NOR2xp33_ASAP7_75t_L g550 ( 
.A(n_543),
.B(n_547),
.Y(n_550)
);

MAJIxp5_ASAP7_75t_L g544 ( 
.A(n_529),
.B(n_520),
.C(n_13),
.Y(n_544)
);

MAJIxp5_ASAP7_75t_L g551 ( 
.A(n_544),
.B(n_534),
.C(n_533),
.Y(n_551)
);

NOR2xp33_ASAP7_75t_L g546 ( 
.A(n_535),
.B(n_13),
.Y(n_546)
);

CKINVDCx20_ASAP7_75t_R g554 ( 
.A(n_546),
.Y(n_554)
);

NOR2xp33_ASAP7_75t_L g547 ( 
.A(n_536),
.B(n_524),
.Y(n_547)
);

XOR2xp5_ASAP7_75t_L g548 ( 
.A(n_528),
.B(n_526),
.Y(n_548)
);

XOR2xp5_ASAP7_75t_L g552 ( 
.A(n_548),
.B(n_523),
.Y(n_552)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_551),
.Y(n_558)
);

OR2x2_ASAP7_75t_L g559 ( 
.A(n_552),
.B(n_553),
.Y(n_559)
);

MAJIxp5_ASAP7_75t_L g553 ( 
.A(n_548),
.B(n_537),
.C(n_530),
.Y(n_553)
);

OAI21x1_ASAP7_75t_L g556 ( 
.A1(n_550),
.A2(n_545),
.B(n_530),
.Y(n_556)
);

NOR2xp33_ASAP7_75t_L g560 ( 
.A(n_556),
.B(n_557),
.Y(n_560)
);

INVxp67_ASAP7_75t_L g557 ( 
.A(n_549),
.Y(n_557)
);

INVxp67_ASAP7_75t_L g561 ( 
.A(n_559),
.Y(n_561)
);

BUFx24_ASAP7_75t_SL g562 ( 
.A(n_561),
.Y(n_562)
);

INVxp67_ASAP7_75t_L g563 ( 
.A(n_562),
.Y(n_563)
);

AOI322xp5_ASAP7_75t_L g564 ( 
.A1(n_563),
.A2(n_560),
.A3(n_558),
.B1(n_554),
.B2(n_541),
.C1(n_553),
.C2(n_555),
.Y(n_564)
);

FAx1_ASAP7_75t_SL g565 ( 
.A(n_564),
.B(n_540),
.CI(n_537),
.CON(n_565),
.SN(n_565)
);

MAJIxp5_ASAP7_75t_L g566 ( 
.A(n_565),
.B(n_541),
.C(n_552),
.Y(n_566)
);

AO21x1_ASAP7_75t_L g567 ( 
.A1(n_566),
.A2(n_565),
.B(n_534),
.Y(n_567)
);


endmodule