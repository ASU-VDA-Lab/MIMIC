module real_jpeg_29701_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_68;
wire n_146;
wire n_83;
wire n_78;
wire n_166;
wire n_176;
wire n_215;
wire n_221;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_200;
wire n_164;
wire n_140;
wire n_126;
wire n_214;
wire n_120;
wire n_113;
wire n_155;
wire n_199;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_188;
wire n_139;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_208;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_172;
wire n_160;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_203;
wire n_192;
wire n_100;
wire n_198;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_110;
wire n_61;
wire n_205;
wire n_195;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_103;
wire n_225;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_185;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_97;
wire n_75;
wire n_187;
wire n_34;
wire n_190;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_216;
wire n_128;
wire n_167;
wire n_179;
wire n_202;
wire n_213;
wire n_133;
wire n_138;
wire n_25;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;

INVx11_ASAP7_75t_L g38 ( 
.A(n_0),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_1),
.A2(n_29),
.B1(n_59),
.B2(n_63),
.Y(n_62)
);

CKINVDCx16_ASAP7_75t_R g63 ( 
.A(n_1),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_1),
.A2(n_30),
.B1(n_63),
.B2(n_73),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_SL g168 ( 
.A1(n_1),
.A2(n_35),
.B1(n_41),
.B2(n_63),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_1),
.A2(n_55),
.B1(n_56),
.B2(n_63),
.Y(n_200)
);

AOI22xp33_ASAP7_75t_L g66 ( 
.A1(n_2),
.A2(n_29),
.B1(n_59),
.B2(n_67),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_2),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_2),
.A2(n_30),
.B1(n_67),
.B2(n_73),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_L g102 ( 
.A1(n_2),
.A2(n_55),
.B1(n_56),
.B2(n_67),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_2),
.A2(n_35),
.B1(n_41),
.B2(n_67),
.Y(n_171)
);

BUFx12_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_4),
.A2(n_55),
.B1(n_56),
.B2(n_88),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_4),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_4),
.A2(n_29),
.B1(n_59),
.B2(n_88),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_L g145 ( 
.A1(n_4),
.A2(n_35),
.B1(n_41),
.B2(n_88),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_5),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_SL g46 ( 
.A1(n_6),
.A2(n_35),
.B1(n_41),
.B2(n_47),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_6),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_L g129 ( 
.A1(n_6),
.A2(n_47),
.B1(n_55),
.B2(n_56),
.Y(n_129)
);

BUFx10_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_8),
.A2(n_30),
.B1(n_72),
.B2(n_73),
.Y(n_71)
);

CKINVDCx16_ASAP7_75t_R g72 ( 
.A(n_8),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_L g109 ( 
.A1(n_8),
.A2(n_29),
.B1(n_59),
.B2(n_72),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_SL g166 ( 
.A1(n_8),
.A2(n_55),
.B1(n_56),
.B2(n_72),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_SL g176 ( 
.A1(n_8),
.A2(n_35),
.B1(n_41),
.B2(n_72),
.Y(n_176)
);

AOI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_9),
.A2(n_35),
.B1(n_41),
.B2(n_127),
.Y(n_126)
);

CKINVDCx16_ASAP7_75t_R g127 ( 
.A(n_9),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_SL g40 ( 
.A1(n_10),
.A2(n_35),
.B1(n_41),
.B2(n_42),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_10),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_L g95 ( 
.A1(n_10),
.A2(n_42),
.B1(n_55),
.B2(n_56),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_L g84 ( 
.A1(n_11),
.A2(n_35),
.B1(n_41),
.B2(n_85),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_11),
.Y(n_85)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

AOI21xp5_ASAP7_75t_L g28 ( 
.A1(n_12),
.A2(n_27),
.B(n_29),
.Y(n_28)
);

OAI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_12),
.A2(n_25),
.B1(n_30),
.B2(n_73),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_12),
.B(n_56),
.Y(n_156)
);

A2O1A1O1Ixp25_ASAP7_75t_L g158 ( 
.A1(n_12),
.A2(n_56),
.B(n_90),
.C(n_156),
.D(n_159),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_12),
.B(n_53),
.Y(n_163)
);

OAI21xp33_ASAP7_75t_L g186 ( 
.A1(n_12),
.A2(n_34),
.B(n_169),
.Y(n_186)
);

A2O1A1O1Ixp25_ASAP7_75t_L g196 ( 
.A1(n_12),
.A2(n_52),
.B(n_59),
.C(n_65),
.D(n_197),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_12),
.B(n_59),
.Y(n_197)
);

INVx11_ASAP7_75t_L g92 ( 
.A(n_13),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_13),
.A2(n_35),
.B1(n_41),
.B2(n_92),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_13),
.B(n_35),
.Y(n_157)
);

BUFx24_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_15),
.A2(n_54),
.B1(n_55),
.B2(n_56),
.Y(n_53)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_15),
.Y(n_54)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_15),
.Y(n_58)
);

INVx11_ASAP7_75t_SL g37 ( 
.A(n_16),
.Y(n_37)
);

XOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_135),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_133),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_110),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_SL g134 ( 
.A(n_20),
.B(n_110),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_81),
.C(n_97),
.Y(n_20)
);

XNOR2xp5_ASAP7_75t_L g147 ( 
.A(n_21),
.B(n_148),
.Y(n_147)
);

XOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_48),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_22),
.B(n_49),
.C(n_80),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_31),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_23),
.A2(n_24),
.B1(n_31),
.B2(n_32),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_24),
.Y(n_23)
);

A2O1A1Ixp33_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_26),
.B(n_28),
.C(n_30),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_SL g146 ( 
.A(n_25),
.B(n_74),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_SL g181 ( 
.A(n_25),
.B(n_96),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_25),
.B(n_38),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_26),
.A2(n_27),
.B1(n_29),
.B2(n_59),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_L g78 ( 
.A1(n_26),
.A2(n_27),
.B1(n_30),
.B2(n_73),
.Y(n_78)
);

CKINVDCx14_ASAP7_75t_R g26 ( 
.A(n_27),
.Y(n_26)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_29),
.A2(n_58),
.B1(n_59),
.B2(n_60),
.Y(n_57)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_29),
.Y(n_59)
);

AOI32xp33_ASAP7_75t_L g204 ( 
.A1(n_29),
.A2(n_56),
.A3(n_197),
.B1(n_205),
.B2(n_206),
.Y(n_204)
);

INVx13_ASAP7_75t_L g73 ( 
.A(n_30),
.Y(n_73)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

AOI22xp5_ASAP7_75t_L g32 ( 
.A1(n_33),
.A2(n_39),
.B1(n_43),
.B2(n_46),
.Y(n_32)
);

AOI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_33),
.A2(n_43),
.B1(n_175),
.B2(n_177),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_34),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_34),
.A2(n_38),
.B1(n_83),
.B2(n_84),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_34),
.A2(n_84),
.B1(n_125),
.B2(n_126),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_34),
.A2(n_40),
.B1(n_44),
.B2(n_145),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_L g167 ( 
.A1(n_34),
.A2(n_168),
.B(n_169),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_34),
.B(n_171),
.Y(n_184)
);

NAND2x1_ASAP7_75t_SL g34 ( 
.A(n_35),
.B(n_38),
.Y(n_34)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_35),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx11_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx11_ASAP7_75t_L g45 ( 
.A(n_38),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_40),
.Y(n_39)
);

AOI32xp33_ASAP7_75t_L g155 ( 
.A1(n_41),
.A2(n_55),
.A3(n_92),
.B1(n_156),
.B2(n_157),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_SL g187 ( 
.A(n_41),
.B(n_188),
.Y(n_187)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

OAI21xp5_ASAP7_75t_SL g182 ( 
.A1(n_44),
.A2(n_176),
.B(n_183),
.Y(n_182)
);

INVx11_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx5_ASAP7_75t_SL g125 ( 
.A(n_45),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_45),
.B(n_170),
.Y(n_169)
);

AOI21xp5_ASAP7_75t_L g202 ( 
.A1(n_45),
.A2(n_184),
.B(n_203),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_46),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g48 ( 
.A1(n_49),
.A2(n_50),
.B1(n_69),
.B2(n_80),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_50),
.Y(n_49)
);

OAI21xp5_ASAP7_75t_SL g50 ( 
.A1(n_51),
.A2(n_61),
.B(n_64),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_52),
.A2(n_53),
.B1(n_62),
.B2(n_108),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_52),
.B(n_122),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_SL g52 ( 
.A(n_53),
.B(n_57),
.Y(n_52)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_53),
.Y(n_68)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_54),
.Y(n_60)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_55),
.Y(n_56)
);

NAND2xp33_ASAP7_75t_SL g206 ( 
.A(n_55),
.B(n_60),
.Y(n_206)
);

O2A1O1Ixp33_ASAP7_75t_L g90 ( 
.A1(n_56),
.A2(n_91),
.B(n_93),
.C(n_94),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_56),
.B(n_91),
.Y(n_93)
);

INVx6_ASAP7_75t_L g205 ( 
.A(n_60),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_62),
.Y(n_61)
);

INVxp67_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_66),
.B(n_68),
.Y(n_65)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_66),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_L g119 ( 
.A1(n_68),
.A2(n_120),
.B(n_121),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_L g143 ( 
.A1(n_68),
.A2(n_109),
.B(n_121),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_69),
.Y(n_80)
);

OAI21xp5_ASAP7_75t_L g69 ( 
.A1(n_70),
.A2(n_74),
.B(n_76),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_71),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_71),
.A2(n_75),
.B1(n_77),
.B2(n_117),
.Y(n_116)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g77 ( 
.A(n_75),
.B(n_78),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_75),
.B(n_79),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_77),
.B(n_79),
.Y(n_76)
);

AOI21xp5_ASAP7_75t_L g103 ( 
.A1(n_77),
.A2(n_104),
.B(n_105),
.Y(n_103)
);

XNOR2xp5_ASAP7_75t_L g148 ( 
.A(n_81),
.B(n_97),
.Y(n_148)
);

XOR2xp5_ASAP7_75t_L g81 ( 
.A(n_82),
.B(n_86),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_82),
.B(n_86),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_87),
.A2(n_89),
.B1(n_95),
.B2(n_96),
.Y(n_86)
);

OAI21xp5_ASAP7_75t_SL g99 ( 
.A1(n_87),
.A2(n_96),
.B(n_100),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_89),
.A2(n_95),
.B1(n_96),
.B2(n_129),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_SL g215 ( 
.A1(n_89),
.A2(n_216),
.B(n_217),
.Y(n_215)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_90),
.B(n_101),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_90),
.A2(n_94),
.B1(n_199),
.B2(n_200),
.Y(n_198)
);

INVx11_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_94),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_96),
.B(n_102),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_L g165 ( 
.A1(n_96),
.A2(n_100),
.B(n_166),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_98),
.B(n_103),
.C(n_107),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_98),
.A2(n_99),
.B1(n_107),
.B2(n_140),
.Y(n_139)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

CKINVDCx16_ASAP7_75t_R g101 ( 
.A(n_102),
.Y(n_101)
);

XNOR2xp5_ASAP7_75t_SL g138 ( 
.A(n_103),
.B(n_139),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_106),
.Y(n_105)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_107),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_109),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_111),
.A2(n_130),
.B1(n_131),
.B2(n_132),
.Y(n_110)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_111),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_SL g111 ( 
.A(n_112),
.B(n_123),
.Y(n_111)
);

XNOR2xp5_ASAP7_75t_SL g112 ( 
.A(n_113),
.B(n_114),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_115),
.A2(n_116),
.B1(n_118),
.B2(n_119),
.Y(n_114)
);

CKINVDCx14_ASAP7_75t_R g115 ( 
.A(n_116),
.Y(n_115)
);

CKINVDCx14_ASAP7_75t_R g118 ( 
.A(n_119),
.Y(n_118)
);

XNOR2xp5_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_128),
.Y(n_123)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_130),
.Y(n_132)
);

INVxp67_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_L g135 ( 
.A1(n_136),
.A2(n_149),
.B(n_224),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_147),
.Y(n_136)
);

AND2x2_ASAP7_75t_L g225 ( 
.A(n_137),
.B(n_147),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_141),
.C(n_142),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_138),
.B(n_222),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_141),
.B(n_142),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_143),
.B(n_144),
.C(n_146),
.Y(n_142)
);

XNOR2xp5_ASAP7_75t_SL g211 ( 
.A(n_143),
.B(n_212),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g212 ( 
.A(n_144),
.B(n_146),
.Y(n_212)
);

CKINVDCx16_ASAP7_75t_R g203 ( 
.A(n_145),
.Y(n_203)
);

AOI21xp5_ASAP7_75t_L g149 ( 
.A1(n_150),
.A2(n_219),
.B(n_223),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_SL g150 ( 
.A1(n_151),
.A2(n_208),
.B(n_218),
.Y(n_150)
);

AOI21xp5_ASAP7_75t_L g151 ( 
.A1(n_152),
.A2(n_192),
.B(n_207),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_SL g152 ( 
.A1(n_153),
.A2(n_172),
.B(n_191),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_160),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_154),
.B(n_160),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_158),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_L g178 ( 
.A(n_155),
.B(n_158),
.Y(n_178)
);

INVxp67_ASAP7_75t_L g217 ( 
.A(n_159),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g160 ( 
.A(n_161),
.B(n_167),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_162),
.A2(n_163),
.B1(n_164),
.B2(n_165),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_162),
.B(n_165),
.C(n_167),
.Y(n_193)
);

CKINVDCx16_ASAP7_75t_R g162 ( 
.A(n_163),
.Y(n_162)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_166),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_168),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_171),
.Y(n_170)
);

AOI21xp5_ASAP7_75t_L g172 ( 
.A1(n_173),
.A2(n_179),
.B(n_190),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_178),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_SL g190 ( 
.A(n_174),
.B(n_178),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_176),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_SL g179 ( 
.A1(n_180),
.A2(n_185),
.B(n_189),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_182),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_181),
.B(n_182),
.Y(n_189)
);

INVxp67_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_186),
.B(n_187),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_193),
.B(n_194),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_SL g207 ( 
.A(n_193),
.B(n_194),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_L g194 ( 
.A(n_195),
.B(n_201),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_198),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_196),
.B(n_198),
.C(n_201),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_200),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_SL g201 ( 
.A(n_202),
.B(n_204),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_202),
.B(n_204),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_209),
.B(n_210),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_209),
.B(n_210),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g210 ( 
.A(n_211),
.B(n_213),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_211),
.B(n_214),
.C(n_215),
.Y(n_220)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_214),
.B(n_215),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_220),
.B(n_221),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_SL g223 ( 
.A(n_220),
.B(n_221),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_225),
.Y(n_224)
);


endmodule