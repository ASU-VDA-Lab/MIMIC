module fake_jpeg_7723_n_139 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_139);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_139;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_57;
wire n_21;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_7),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_6),
.Y(n_13)
);

INVx4_ASAP7_75t_L g14 ( 
.A(n_11),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_0),
.Y(n_15)
);

INVx3_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

INVx4_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

INVx6_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_2),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_5),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_11),
.Y(n_22)
);

BUFx16f_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_1),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_10),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_18),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_SL g38 ( 
.A(n_27),
.B(n_33),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_23),
.Y(n_28)
);

INVx2_ASAP7_75t_SL g44 ( 
.A(n_28),
.Y(n_44)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_29),
.B(n_30),
.Y(n_39)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_23),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_31),
.B(n_32),
.Y(n_43)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_23),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_18),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_12),
.B(n_0),
.Y(n_34)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_34),
.Y(n_42)
);

INVx11_ASAP7_75t_L g35 ( 
.A(n_15),
.Y(n_35)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_35),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_L g36 ( 
.A1(n_27),
.A2(n_18),
.B1(n_16),
.B2(n_17),
.Y(n_36)
);

AOI22xp33_ASAP7_75t_L g54 ( 
.A1(n_36),
.A2(n_16),
.B1(n_17),
.B2(n_29),
.Y(n_54)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_34),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_40),
.B(n_45),
.Y(n_52)
);

AND2x2_ASAP7_75t_L g41 ( 
.A(n_32),
.B(n_23),
.Y(n_41)
);

AOI21xp5_ASAP7_75t_L g60 ( 
.A1(n_41),
.A2(n_46),
.B(n_26),
.Y(n_60)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_35),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_33),
.A2(n_16),
.B1(n_17),
.B2(n_14),
.Y(n_46)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_47),
.B(n_49),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_32),
.Y(n_48)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_48),
.Y(n_51)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_28),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_50),
.B(n_58),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_42),
.B(n_25),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_SL g68 ( 
.A(n_53),
.B(n_20),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_54),
.A2(n_61),
.B1(n_63),
.B2(n_30),
.Y(n_65)
);

MAJIxp5_ASAP7_75t_L g55 ( 
.A(n_43),
.B(n_31),
.C(n_23),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_55),
.B(n_41),
.Y(n_64)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_36),
.Y(n_56)
);

BUFx2_ASAP7_75t_SL g66 ( 
.A(n_56),
.Y(n_66)
);

OAI21xp5_ASAP7_75t_SL g57 ( 
.A1(n_39),
.A2(n_31),
.B(n_26),
.Y(n_57)
);

INVxp67_ASAP7_75t_L g67 ( 
.A(n_57),
.Y(n_67)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_37),
.Y(n_58)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_37),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_59),
.B(n_60),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_42),
.A2(n_26),
.B1(n_21),
.B2(n_29),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_45),
.A2(n_21),
.B1(n_29),
.B2(n_30),
.Y(n_63)
);

XOR2xp5_ASAP7_75t_L g85 ( 
.A(n_64),
.B(n_44),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_65),
.A2(n_75),
.B1(n_51),
.B2(n_24),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_68),
.B(n_69),
.Y(n_89)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_62),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_52),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_70),
.B(n_72),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_SL g72 ( 
.A(n_50),
.B(n_20),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_55),
.B(n_41),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_73),
.B(n_15),
.Y(n_87)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_58),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_74),
.B(n_77),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_56),
.A2(n_47),
.B1(n_21),
.B2(n_15),
.Y(n_75)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_59),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_57),
.Y(n_78)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_78),
.Y(n_81)
);

OAI21xp5_ASAP7_75t_L g79 ( 
.A1(n_67),
.A2(n_60),
.B(n_19),
.Y(n_79)
);

XOR2xp5_ASAP7_75t_L g94 ( 
.A(n_79),
.B(n_85),
.Y(n_94)
);

INVx13_ASAP7_75t_L g80 ( 
.A(n_74),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_80),
.B(n_83),
.Y(n_98)
);

OA21x2_ASAP7_75t_L g83 ( 
.A1(n_78),
.A2(n_15),
.B(n_28),
.Y(n_83)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_71),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_84),
.B(n_87),
.Y(n_102)
);

OAI21xp5_ASAP7_75t_L g86 ( 
.A1(n_67),
.A2(n_24),
.B(n_19),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_86),
.B(n_88),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_64),
.B(n_51),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_90),
.A2(n_75),
.B1(n_70),
.B2(n_66),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_91),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_92),
.B(n_95),
.Y(n_107)
);

CKINVDCx16_ASAP7_75t_R g95 ( 
.A(n_82),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_80),
.Y(n_96)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_96),
.Y(n_106)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_89),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_97),
.B(n_99),
.Y(n_104)
);

OAI22x1_ASAP7_75t_L g100 ( 
.A1(n_83),
.A2(n_76),
.B1(n_65),
.B2(n_73),
.Y(n_100)
);

AOI21xp5_ASAP7_75t_L g109 ( 
.A1(n_100),
.A2(n_83),
.B(n_81),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_84),
.B(n_72),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_101),
.B(n_103),
.Y(n_110)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_88),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_94),
.B(n_85),
.C(n_87),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_105),
.B(n_112),
.Y(n_114)
);

XNOR2xp5_ASAP7_75t_SL g108 ( 
.A(n_94),
.B(n_79),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_108),
.A2(n_113),
.B1(n_103),
.B2(n_93),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_109),
.A2(n_44),
.B1(n_25),
.B2(n_22),
.Y(n_117)
);

XOR2xp5_ASAP7_75t_L g111 ( 
.A(n_100),
.B(n_86),
.Y(n_111)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_111),
.Y(n_119)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_102),
.Y(n_112)
);

OAI32xp33_ASAP7_75t_L g113 ( 
.A1(n_93),
.A2(n_81),
.A3(n_90),
.B1(n_69),
.B2(n_77),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_SL g126 ( 
.A(n_115),
.B(n_113),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_104),
.A2(n_98),
.B1(n_96),
.B2(n_12),
.Y(n_116)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_116),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_117),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_108),
.A2(n_22),
.B1(n_13),
.B2(n_48),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_118),
.B(n_120),
.C(n_110),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_107),
.A2(n_13),
.B1(n_44),
.B2(n_3),
.Y(n_120)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_122),
.Y(n_128)
);

HB1xp67_ASAP7_75t_L g124 ( 
.A(n_114),
.Y(n_124)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_124),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_119),
.B(n_105),
.C(n_111),
.Y(n_125)
);

XNOR2xp5_ASAP7_75t_L g129 ( 
.A(n_125),
.B(n_126),
.Y(n_129)
);

AND2x2_ASAP7_75t_L g127 ( 
.A(n_121),
.B(n_115),
.Y(n_127)
);

AOI322xp5_ASAP7_75t_L g132 ( 
.A1(n_127),
.A2(n_128),
.A3(n_130),
.B1(n_129),
.B2(n_106),
.C1(n_8),
.C2(n_9),
.Y(n_132)
);

O2A1O1Ixp33_ASAP7_75t_L g131 ( 
.A1(n_127),
.A2(n_123),
.B(n_116),
.C(n_118),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_131),
.B(n_2),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_132),
.B(n_133),
.C(n_0),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_128),
.B(n_8),
.C(n_10),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_134),
.B(n_135),
.C(n_2),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_136),
.B(n_3),
.Y(n_137)
);

AOI21xp5_ASAP7_75t_L g138 ( 
.A1(n_137),
.A2(n_3),
.B(n_4),
.Y(n_138)
);

XOR2xp5_ASAP7_75t_L g139 ( 
.A(n_138),
.B(n_4),
.Y(n_139)
);


endmodule