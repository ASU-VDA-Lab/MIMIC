module real_aes_1345_n_270 (n_17, n_28, n_226, n_76, n_202, n_255, n_149, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_257, n_261, n_262, n_238, n_65, n_47, n_74, n_106, n_58, n_185, n_134, n_32, n_30, n_263, n_230, n_165, n_51, n_195, n_246, n_248, n_252, n_176, n_27, n_163, n_222, n_249, n_61, n_29, n_20, n_52, n_221, n_174, n_156, n_57, n_64, n_66, n_254, n_18, n_207, n_104, n_21, n_31, n_8, n_251, n_183, n_266, n_205, n_220, n_211, n_10, n_177, n_83, n_181, n_197, n_124, n_22, n_173, n_191, n_209, n_3, n_41, n_140, n_234, n_153, n_75, n_178, n_219, n_256, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_239, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_224, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_253, n_35, n_42, n_147, n_150, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_95, n_131, n_144, n_164, n_231, n_169, n_242, n_44, n_102, n_188, n_269, n_152, n_198, n_201, n_122, n_7, n_228, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_232, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_69, n_46, n_109, n_59, n_25, n_203, n_236, n_73, n_77, n_218, n_81, n_133, n_48, n_267, n_260, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_138, n_50, n_114, n_89, n_170, n_26, n_235, n_265, n_86, n_93, n_182, n_154, n_127, n_199, n_245, n_161, n_189, n_13, n_24, n_217, n_2, n_142, n_55, n_168, n_175, n_241, n_145, n_62, n_105, n_223, n_84, n_227, n_67, n_92, n_33, n_206, n_258, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_225, n_16, n_250, n_116, n_94, n_229, n_39, n_5, n_45, n_60, n_233, n_240, n_247, n_38, n_259, n_155, n_243, n_118, n_143, n_139, n_244, n_192, n_213, n_268, n_136, n_87, n_171, n_0, n_157, n_78, n_264, n_101, n_63, n_1, n_146, n_237, n_107, n_184, n_53, n_36, n_270);
input n_17;
input n_28;
input n_226;
input n_76;
input n_202;
input n_255;
input n_149;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_257;
input n_261;
input n_262;
input n_238;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_134;
input n_32;
input n_30;
input n_263;
input n_230;
input n_165;
input n_51;
input n_195;
input n_246;
input n_248;
input n_252;
input n_176;
input n_27;
input n_163;
input n_222;
input n_249;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_254;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_251;
input n_183;
input n_266;
input n_205;
input n_220;
input n_211;
input n_10;
input n_177;
input n_83;
input n_181;
input n_197;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_3;
input n_41;
input n_140;
input n_234;
input n_153;
input n_75;
input n_178;
input n_219;
input n_256;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_239;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_224;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_253;
input n_35;
input n_42;
input n_147;
input n_150;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_95;
input n_131;
input n_144;
input n_164;
input n_231;
input n_169;
input n_242;
input n_44;
input n_102;
input n_188;
input n_269;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_228;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_232;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_69;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_236;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_267;
input n_260;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_138;
input n_50;
input n_114;
input n_89;
input n_170;
input n_26;
input n_235;
input n_265;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_245;
input n_161;
input n_189;
input n_13;
input n_24;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_241;
input n_145;
input n_62;
input n_105;
input n_223;
input n_84;
input n_227;
input n_67;
input n_92;
input n_33;
input n_206;
input n_258;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_225;
input n_16;
input n_250;
input n_116;
input n_94;
input n_229;
input n_39;
input n_5;
input n_45;
input n_60;
input n_233;
input n_240;
input n_247;
input n_38;
input n_259;
input n_155;
input n_243;
input n_118;
input n_143;
input n_139;
input n_244;
input n_192;
input n_213;
input n_268;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_264;
input n_101;
input n_63;
input n_1;
input n_146;
input n_237;
input n_107;
input n_184;
input n_53;
input n_36;
output n_270;
wire n_480;
wire n_476;
wire n_758;
wire n_599;
wire n_436;
wire n_684;
wire n_390;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_522;
wire n_485;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_362;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_766;
wire n_461;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_537;
wire n_666;
wire n_560;
wire n_660;
wire n_594;
wire n_767;
wire n_696;
wire n_704;
wire n_453;
wire n_379;
wire n_374;
wire n_647;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_775;
wire n_763;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_415;
wire n_572;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_578;
wire n_528;
wire n_372;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_352;
wire n_467;
wire n_327;
wire n_774;
wire n_466;
wire n_559;
wire n_636;
wire n_477;
wire n_515;
wire n_680;
wire n_595;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_570;
wire n_675;
wire n_530;
wire n_535;
wire n_732;
wire n_281;
wire n_496;
wire n_693;
wire n_468;
wire n_746;
wire n_284;
wire n_316;
wire n_532;
wire n_656;
wire n_755;
wire n_409;
wire n_748;
wire n_781;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_310;
wire n_725;
wire n_455;
wire n_504;
wire n_671;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_443;
wire n_565;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_457;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_664;
wire n_278;
wire n_367;
wire n_737;
wire n_581;
wire n_610;
wire n_620;
wire n_582;
wire n_641;
wire n_770;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_363;
wire n_417;
wire n_754;
wire n_449;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_561;
wire n_437;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_505;
wire n_527;
wire n_434;
wire n_502;
wire n_769;
wire n_600;
wire n_731;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_733;
wire n_402;
wire n_552;
wire n_602;
wire n_617;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_286;
wire n_416;
wire n_410;
wire n_751;
wire n_490;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_361;
wire n_632;
wire n_768;
wire n_412;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_642;
wire n_613;
wire n_387;
wire n_296;
wire n_702;
wire n_302;
wire n_464;
wire n_351;
wire n_604;
wire n_734;
wire n_392;
wire n_562;
wire n_288;
wire n_713;
wire n_404;
wire n_598;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_274;
wire n_569;
wire n_303;
wire n_563;
wire n_430;
wire n_568;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_397;
wire n_293;
wire n_358;
wire n_385;
wire n_275;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_536;
wire n_707;
wire n_622;
wire n_470;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_720;
wire n_354;
wire n_435;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_481;
wire n_498;
wire n_691;
wire n_765;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_692;
wire n_544;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_482;
wire n_633;
wire n_520;
wire n_679;
wire n_472;
wire n_452;
wire n_630;
wire n_689;
wire n_715;
wire n_420;
wire n_349;
wire n_336;
wire n_612;
wire n_438;
wire n_764;
wire n_300;
wire n_741;
wire n_283;
wire n_314;
wire n_753;
wire n_623;
wire n_446;
wire n_721;
wire n_681;
wire n_456;
wire n_359;
wire n_717;
wire n_312;
wire n_712;
wire n_433;
wire n_335;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_524;
wire n_705;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_541;
wire n_546;
wire n_587;
wire n_639;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_272;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_279;
wire n_686;
wire n_776;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_441;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_375;
wire n_597;
wire n_640;
wire n_340;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_743;
wire n_393;
wire n_294;
wire n_652;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_424;
wire n_574;
wire n_337;
wire n_475;
wire n_554;
wire n_668;
AOI22xp33_ASAP7_75t_L g509 ( .A1(n_0), .A2(n_223), .B1(n_305), .B2(n_510), .Y(n_509) );
AO222x2_ASAP7_75t_SL g387 ( .A1(n_1), .A2(n_31), .B1(n_145), .B2(n_363), .C1(n_388), .C2(n_391), .Y(n_387) );
CKINVDCx20_ASAP7_75t_R g700 ( .A(n_2), .Y(n_700) );
AOI22xp33_ASAP7_75t_L g770 ( .A1(n_3), .A2(n_92), .B1(n_410), .B2(n_460), .Y(n_770) );
AOI22xp5_ASAP7_75t_L g767 ( .A1(n_4), .A2(n_231), .B1(n_709), .B2(n_768), .Y(n_767) );
AOI22xp33_ASAP7_75t_L g673 ( .A1(n_5), .A2(n_227), .B1(n_334), .B2(n_335), .Y(n_673) );
AOI22xp5_ASAP7_75t_L g530 ( .A1(n_6), .A2(n_243), .B1(n_427), .B2(n_531), .Y(n_530) );
AOI22xp33_ASAP7_75t_L g399 ( .A1(n_7), .A2(n_23), .B1(n_400), .B2(n_402), .Y(n_399) );
AO22x2_ASAP7_75t_L g295 ( .A1(n_8), .A2(n_177), .B1(n_296), .B2(n_297), .Y(n_295) );
INVx1_ASAP7_75t_L g729 ( .A(n_8), .Y(n_729) );
AOI22xp33_ASAP7_75t_L g573 ( .A1(n_9), .A2(n_221), .B1(n_427), .B2(n_531), .Y(n_573) );
AOI22xp33_ASAP7_75t_L g565 ( .A1(n_10), .A2(n_63), .B1(n_396), .B2(n_398), .Y(n_565) );
AOI22xp33_ASAP7_75t_L g675 ( .A1(n_11), .A2(n_252), .B1(n_330), .B2(n_341), .Y(n_675) );
AOI22xp33_ASAP7_75t_L g564 ( .A1(n_12), .A2(n_100), .B1(n_388), .B2(n_393), .Y(n_564) );
AOI22xp33_ASAP7_75t_L g666 ( .A1(n_13), .A2(n_160), .B1(n_413), .B2(n_417), .Y(n_666) );
OA22x2_ASAP7_75t_L g286 ( .A1(n_14), .A2(n_287), .B1(n_288), .B2(n_289), .Y(n_286) );
INVx1_ASAP7_75t_L g287 ( .A(n_14), .Y(n_287) );
AOI22xp33_ASAP7_75t_SL g762 ( .A1(n_15), .A2(n_19), .B1(n_741), .B2(n_742), .Y(n_762) );
AOI22xp5_ASAP7_75t_L g340 ( .A1(n_16), .A2(n_26), .B1(n_341), .B2(n_342), .Y(n_340) );
AOI22xp5_ASAP7_75t_L g366 ( .A1(n_17), .A2(n_84), .B1(n_367), .B2(n_370), .Y(n_366) );
AOI22xp33_ASAP7_75t_L g746 ( .A1(n_18), .A2(n_39), .B1(n_457), .B2(n_709), .Y(n_746) );
AO22x2_ASAP7_75t_L g309 ( .A1(n_20), .A2(n_65), .B1(n_296), .B2(n_310), .Y(n_309) );
NOR2xp33_ASAP7_75t_L g727 ( .A(n_20), .B(n_728), .Y(n_727) );
AOI22xp33_ASAP7_75t_L g616 ( .A1(n_21), .A2(n_148), .B1(n_334), .B2(n_342), .Y(n_616) );
AO222x2_ASAP7_75t_SL g445 ( .A1(n_22), .A2(n_143), .B1(n_249), .B2(n_375), .C1(n_446), .C2(n_447), .Y(n_445) );
AOI22xp5_ASAP7_75t_L g514 ( .A1(n_24), .A2(n_129), .B1(n_358), .B2(n_515), .Y(n_514) );
AOI22xp33_ASAP7_75t_L g674 ( .A1(n_25), .A2(n_201), .B1(n_337), .B2(n_339), .Y(n_674) );
AOI22xp33_ASAP7_75t_L g487 ( .A1(n_27), .A2(n_62), .B1(n_488), .B2(n_489), .Y(n_487) );
AOI22xp33_ASAP7_75t_L g535 ( .A1(n_28), .A2(n_132), .B1(n_536), .B2(n_538), .Y(n_535) );
AOI22xp33_ASAP7_75t_L g740 ( .A1(n_29), .A2(n_52), .B1(n_741), .B2(n_742), .Y(n_740) );
AOI22xp33_ASAP7_75t_L g517 ( .A1(n_30), .A2(n_81), .B1(n_413), .B2(n_416), .Y(n_517) );
AOI22xp5_ASAP7_75t_L g329 ( .A1(n_32), .A2(n_58), .B1(n_330), .B2(n_331), .Y(n_329) );
AOI222xp33_ASAP7_75t_L g291 ( .A1(n_33), .A2(n_224), .B1(n_259), .B2(n_292), .C1(n_305), .C2(n_311), .Y(n_291) );
AOI22xp33_ASAP7_75t_L g737 ( .A1(n_34), .A2(n_253), .B1(n_460), .B2(n_538), .Y(n_737) );
AOI22xp33_ASAP7_75t_L g518 ( .A1(n_35), .A2(n_268), .B1(n_334), .B2(n_335), .Y(n_518) );
AOI22xp33_ASAP7_75t_L g615 ( .A1(n_36), .A2(n_232), .B1(n_335), .B2(n_341), .Y(n_615) );
AOI22xp5_ASAP7_75t_L g333 ( .A1(n_37), .A2(n_116), .B1(n_334), .B2(n_335), .Y(n_333) );
AOI22xp5_ASAP7_75t_L g479 ( .A1(n_38), .A2(n_156), .B1(n_444), .B2(n_480), .Y(n_479) );
AOI22xp33_ASAP7_75t_L g609 ( .A1(n_40), .A2(n_113), .B1(n_305), .B2(n_510), .Y(n_609) );
CKINVDCx20_ASAP7_75t_R g702 ( .A(n_41), .Y(n_702) );
AOI22xp33_ASAP7_75t_L g357 ( .A1(n_42), .A2(n_181), .B1(n_334), .B2(n_358), .Y(n_357) );
AOI22xp33_ASAP7_75t_L g682 ( .A1(n_43), .A2(n_169), .B1(n_319), .B2(n_508), .Y(n_682) );
AOI22xp33_ASAP7_75t_SL g712 ( .A1(n_44), .A2(n_53), .B1(n_465), .B2(n_713), .Y(n_712) );
AOI22xp33_ASAP7_75t_L g657 ( .A1(n_45), .A2(n_192), .B1(n_482), .B2(n_563), .Y(n_657) );
AOI22xp33_ASAP7_75t_L g546 ( .A1(n_46), .A2(n_139), .B1(n_547), .B2(n_548), .Y(n_546) );
AOI22xp5_ASAP7_75t_L g771 ( .A1(n_47), .A2(n_131), .B1(n_423), .B2(n_772), .Y(n_771) );
AOI22xp5_ASAP7_75t_L g490 ( .A1(n_48), .A2(n_102), .B1(n_420), .B2(n_491), .Y(n_490) );
AOI22xp33_ASAP7_75t_L g635 ( .A1(n_49), .A2(n_258), .B1(n_410), .B2(n_636), .Y(n_635) );
AOI22xp33_ASAP7_75t_L g660 ( .A1(n_50), .A2(n_74), .B1(n_638), .B2(n_661), .Y(n_660) );
AOI22xp33_ASAP7_75t_SL g323 ( .A1(n_51), .A2(n_262), .B1(n_324), .B2(n_327), .Y(n_323) );
AOI22xp5_ASAP7_75t_L g763 ( .A1(n_54), .A2(n_220), .B1(n_547), .B2(n_548), .Y(n_763) );
AOI22xp33_ASAP7_75t_L g766 ( .A1(n_55), .A2(n_248), .B1(n_451), .B2(n_462), .Y(n_766) );
AOI22xp33_ASAP7_75t_L g459 ( .A1(n_56), .A2(n_141), .B1(n_460), .B2(n_462), .Y(n_459) );
AOI22xp33_ASAP7_75t_SL g759 ( .A1(n_57), .A2(n_267), .B1(n_626), .B2(n_760), .Y(n_759) );
AOI22xp33_ASAP7_75t_L g348 ( .A1(n_59), .A2(n_196), .B1(n_335), .B2(n_349), .Y(n_348) );
AOI22xp33_ASAP7_75t_L g395 ( .A1(n_60), .A2(n_97), .B1(n_396), .B2(n_398), .Y(n_395) );
AOI22xp33_ASAP7_75t_L g676 ( .A1(n_61), .A2(n_120), .B1(n_331), .B2(n_461), .Y(n_676) );
AOI22xp5_ASAP7_75t_L g605 ( .A1(n_64), .A2(n_80), .B1(n_327), .B2(n_505), .Y(n_605) );
AOI22xp33_ASAP7_75t_L g654 ( .A1(n_66), .A2(n_137), .B1(n_397), .B2(n_626), .Y(n_654) );
AOI22xp33_ASAP7_75t_L g450 ( .A1(n_67), .A2(n_98), .B1(n_451), .B2(n_453), .Y(n_450) );
AOI22xp5_ASAP7_75t_L g336 ( .A1(n_68), .A2(n_261), .B1(n_337), .B2(n_339), .Y(n_336) );
XNOR2x2_ASAP7_75t_L g619 ( .A(n_69), .B(n_620), .Y(n_619) );
AOI22xp33_ASAP7_75t_L g628 ( .A1(n_70), .A2(n_187), .B1(n_389), .B2(n_629), .Y(n_628) );
NAND2xp5_ASAP7_75t_L g630 ( .A(n_71), .B(n_596), .Y(n_630) );
AOI22xp33_ASAP7_75t_L g350 ( .A1(n_72), .A2(n_157), .B1(n_331), .B2(n_351), .Y(n_350) );
AOI22xp33_ASAP7_75t_L g708 ( .A1(n_73), .A2(n_153), .B1(n_457), .B2(n_709), .Y(n_708) );
AOI22xp33_ASAP7_75t_L g667 ( .A1(n_75), .A2(n_218), .B1(n_406), .B2(n_515), .Y(n_667) );
AOI22xp33_ASAP7_75t_L g738 ( .A1(n_76), .A2(n_121), .B1(n_533), .B2(n_534), .Y(n_738) );
AOI22xp33_ASAP7_75t_L g481 ( .A1(n_77), .A2(n_103), .B1(n_482), .B2(n_483), .Y(n_481) );
INVx3_ASAP7_75t_L g296 ( .A(n_78), .Y(n_296) );
AOI22xp33_ASAP7_75t_L g439 ( .A1(n_79), .A2(n_265), .B1(n_367), .B2(n_440), .Y(n_439) );
AOI22xp33_ASAP7_75t_L g745 ( .A1(n_82), .A2(n_230), .B1(n_464), .B2(n_465), .Y(n_745) );
CKINVDCx20_ASAP7_75t_R g411 ( .A(n_83), .Y(n_411) );
AOI22xp33_ASAP7_75t_SL g707 ( .A1(n_85), .A2(n_236), .B1(n_451), .B2(n_534), .Y(n_707) );
AOI22xp33_ASAP7_75t_L g587 ( .A1(n_86), .A2(n_165), .B1(n_330), .B2(n_331), .Y(n_587) );
NAND2xp5_ASAP7_75t_L g696 ( .A(n_87), .B(n_626), .Y(n_696) );
AOI22xp33_ASAP7_75t_L g743 ( .A1(n_88), .A2(n_108), .B1(n_444), .B2(n_547), .Y(n_743) );
OA22x2_ASAP7_75t_L g525 ( .A1(n_89), .A2(n_526), .B1(n_527), .B2(n_528), .Y(n_525) );
INVx1_ASAP7_75t_L g526 ( .A(n_89), .Y(n_526) );
NAND2xp5_ASAP7_75t_SL g566 ( .A(n_90), .B(n_543), .Y(n_566) );
CKINVDCx20_ASAP7_75t_R g694 ( .A(n_91), .Y(n_694) );
AO22x1_ASAP7_75t_L g622 ( .A1(n_93), .A2(n_138), .B1(n_440), .B2(n_623), .Y(n_622) );
AOI22xp33_ASAP7_75t_L g532 ( .A1(n_94), .A2(n_117), .B1(n_533), .B2(n_534), .Y(n_532) );
INVx1_ASAP7_75t_SL g301 ( .A(n_95), .Y(n_301) );
NOR2xp33_ASAP7_75t_L g730 ( .A(n_95), .B(n_118), .Y(n_730) );
AOI222xp33_ASAP7_75t_L g747 ( .A1(n_96), .A2(n_109), .B1(n_226), .B2(n_396), .C1(n_398), .C2(n_477), .Y(n_747) );
INVx2_ASAP7_75t_L g277 ( .A(n_99), .Y(n_277) );
AOI22xp5_ASAP7_75t_L g372 ( .A1(n_101), .A2(n_217), .B1(n_373), .B2(n_375), .Y(n_372) );
XOR2x2_ASAP7_75t_L g582 ( .A(n_104), .B(n_583), .Y(n_582) );
AOI22xp33_ASAP7_75t_L g613 ( .A1(n_105), .A2(n_263), .B1(n_331), .B2(n_351), .Y(n_613) );
AOI22xp33_ASAP7_75t_L g639 ( .A1(n_106), .A2(n_200), .B1(n_640), .B2(n_641), .Y(n_639) );
CKINVDCx20_ASAP7_75t_R g653 ( .A(n_107), .Y(n_653) );
AOI22xp5_ASAP7_75t_L g561 ( .A1(n_110), .A2(n_124), .B1(n_400), .B2(n_562), .Y(n_561) );
AOI22xp33_ASAP7_75t_L g412 ( .A1(n_111), .A2(n_269), .B1(n_413), .B2(n_415), .Y(n_412) );
AOI22xp33_ASAP7_75t_L g574 ( .A1(n_112), .A2(n_126), .B1(n_536), .B2(n_575), .Y(n_574) );
AOI22xp33_ASAP7_75t_L g426 ( .A1(n_114), .A2(n_211), .B1(n_427), .B2(n_430), .Y(n_426) );
XNOR2x1_ASAP7_75t_SL g753 ( .A(n_115), .B(n_754), .Y(n_753) );
INVx1_ASAP7_75t_L g781 ( .A(n_115), .Y(n_781) );
AO22x2_ASAP7_75t_L g303 ( .A1(n_118), .A2(n_184), .B1(n_296), .B2(n_304), .Y(n_303) );
NAND2xp5_ASAP7_75t_L g606 ( .A(n_119), .B(n_311), .Y(n_606) );
AOI22xp33_ASAP7_75t_L g442 ( .A1(n_122), .A2(n_247), .B1(n_443), .B2(n_444), .Y(n_442) );
NAND2xp5_ASAP7_75t_L g362 ( .A(n_123), .B(n_363), .Y(n_362) );
AOI22xp33_ASAP7_75t_SL g656 ( .A1(n_125), .A2(n_152), .B1(n_480), .B2(n_629), .Y(n_656) );
AOI22xp33_ASAP7_75t_L g504 ( .A1(n_127), .A2(n_210), .B1(n_327), .B2(n_505), .Y(n_504) );
AOI22xp33_ASAP7_75t_L g455 ( .A1(n_128), .A2(n_140), .B1(n_456), .B2(n_457), .Y(n_455) );
CKINVDCx20_ASAP7_75t_R g668 ( .A(n_130), .Y(n_668) );
CKINVDCx20_ASAP7_75t_R g503 ( .A(n_133), .Y(n_503) );
INVx1_ASAP7_75t_L g302 ( .A(n_134), .Y(n_302) );
AOI22xp33_ASAP7_75t_SL g513 ( .A1(n_135), .A2(n_197), .B1(n_337), .B2(n_353), .Y(n_513) );
AOI22xp33_ASAP7_75t_L g549 ( .A1(n_136), .A2(n_164), .B1(n_396), .B2(n_398), .Y(n_549) );
AOI22xp5_ASAP7_75t_L g732 ( .A1(n_142), .A2(n_733), .B1(n_734), .B2(n_748), .Y(n_732) );
CKINVDCx20_ASAP7_75t_R g748 ( .A(n_142), .Y(n_748) );
XNOR2xp5_ASAP7_75t_L g689 ( .A(n_144), .B(n_690), .Y(n_689) );
AOI22xp5_ASAP7_75t_L g486 ( .A1(n_146), .A2(n_172), .B1(n_337), .B2(n_339), .Y(n_486) );
AOI22xp33_ASAP7_75t_L g592 ( .A1(n_147), .A2(n_228), .B1(n_367), .B2(n_508), .Y(n_592) );
CKINVDCx20_ASAP7_75t_R g758 ( .A(n_149), .Y(n_758) );
AOI22xp5_ASAP7_75t_L g352 ( .A1(n_150), .A2(n_257), .B1(n_353), .B2(n_355), .Y(n_352) );
NAND2xp5_ASAP7_75t_L g678 ( .A(n_151), .B(n_596), .Y(n_678) );
AOI22xp33_ASAP7_75t_L g588 ( .A1(n_154), .A2(n_214), .B1(n_349), .B2(n_493), .Y(n_588) );
AOI22xp33_ASAP7_75t_SL g507 ( .A1(n_155), .A2(n_254), .B1(n_319), .B2(n_508), .Y(n_507) );
AOI22xp33_ASAP7_75t_L g586 ( .A1(n_158), .A2(n_175), .B1(n_337), .B2(n_339), .Y(n_586) );
AOI22xp33_ASAP7_75t_L g612 ( .A1(n_159), .A2(n_188), .B1(n_337), .B2(n_339), .Y(n_612) );
AO22x2_ASAP7_75t_L g436 ( .A1(n_161), .A2(n_437), .B1(n_466), .B2(n_467), .Y(n_436) );
INVx1_ASAP7_75t_L g467 ( .A(n_161), .Y(n_467) );
AOI22xp5_ASAP7_75t_L g568 ( .A1(n_162), .A2(n_212), .B1(n_569), .B2(n_572), .Y(n_568) );
AOI22xp33_ASAP7_75t_L g550 ( .A1(n_163), .A2(n_235), .B1(n_551), .B2(n_553), .Y(n_550) );
AOI22xp33_ASAP7_75t_L g492 ( .A1(n_166), .A2(n_190), .B1(n_493), .B2(n_494), .Y(n_492) );
AO22x1_ASAP7_75t_L g624 ( .A1(n_167), .A2(n_246), .B1(n_625), .B2(n_626), .Y(n_624) );
AOI22xp33_ASAP7_75t_L g539 ( .A1(n_168), .A2(n_203), .B1(n_464), .B2(n_540), .Y(n_539) );
AOI22xp5_ASAP7_75t_L g608 ( .A1(n_170), .A2(n_202), .B1(n_315), .B2(n_319), .Y(n_608) );
CKINVDCx20_ASAP7_75t_R g704 ( .A(n_171), .Y(n_704) );
AOI22xp5_ASAP7_75t_L g314 ( .A1(n_173), .A2(n_245), .B1(n_315), .B2(n_319), .Y(n_314) );
AOI22xp33_ASAP7_75t_L g463 ( .A1(n_174), .A2(n_193), .B1(n_464), .B2(n_465), .Y(n_463) );
AOI22xp33_ASAP7_75t_L g662 ( .A1(n_176), .A2(n_205), .B1(n_663), .B2(n_664), .Y(n_662) );
AOI22xp33_ASAP7_75t_SL g590 ( .A1(n_178), .A2(n_239), .B1(n_447), .B2(n_591), .Y(n_590) );
AOI22xp33_ASAP7_75t_L g637 ( .A1(n_179), .A2(n_244), .B1(n_457), .B2(n_638), .Y(n_637) );
AOI22xp5_ASAP7_75t_L g632 ( .A1(n_180), .A2(n_222), .B1(n_633), .B2(n_634), .Y(n_632) );
INVx1_ASAP7_75t_L g617 ( .A(n_182), .Y(n_617) );
NAND2xp5_ASAP7_75t_L g542 ( .A(n_183), .B(n_543), .Y(n_542) );
AOI22xp33_ASAP7_75t_L g714 ( .A1(n_185), .A2(n_229), .B1(n_464), .B2(n_715), .Y(n_714) );
AOI22xp33_ASAP7_75t_L g577 ( .A1(n_186), .A2(n_198), .B1(n_462), .B2(n_578), .Y(n_577) );
AOI22xp33_ASAP7_75t_L g679 ( .A1(n_189), .A2(n_241), .B1(n_324), .B2(n_327), .Y(n_679) );
NAND2xp5_ASAP7_75t_L g595 ( .A(n_191), .B(n_596), .Y(n_595) );
CKINVDCx20_ASAP7_75t_R g407 ( .A(n_194), .Y(n_407) );
NAND2xp5_ASAP7_75t_L g476 ( .A(n_195), .B(n_477), .Y(n_476) );
AO21x2_ASAP7_75t_L g384 ( .A1(n_199), .A2(n_385), .B(n_432), .Y(n_384) );
INVx1_ASAP7_75t_L g434 ( .A(n_199), .Y(n_434) );
XOR2x2_ASAP7_75t_L g558 ( .A(n_204), .B(n_559), .Y(n_558) );
NAND2xp5_ASAP7_75t_SL g278 ( .A(n_206), .B(n_279), .Y(n_278) );
INVx1_ASAP7_75t_L g725 ( .A(n_206), .Y(n_725) );
AOI22xp33_ASAP7_75t_L g594 ( .A1(n_207), .A2(n_240), .B1(n_292), .B2(n_305), .Y(n_594) );
AO22x2_ASAP7_75t_L g670 ( .A1(n_208), .A2(n_671), .B1(n_683), .B2(n_684), .Y(n_670) );
CKINVDCx20_ASAP7_75t_R g683 ( .A(n_208), .Y(n_683) );
AOI22xp33_ASAP7_75t_L g478 ( .A1(n_209), .A2(n_250), .B1(n_373), .B2(n_375), .Y(n_478) );
AOI22xp33_ASAP7_75t_L g419 ( .A1(n_213), .A2(n_225), .B1(n_420), .B2(n_423), .Y(n_419) );
AOI211xp5_ASAP7_75t_L g270 ( .A1(n_215), .A2(n_271), .B(n_280), .C(n_731), .Y(n_270) );
INVx1_ASAP7_75t_L g274 ( .A(n_216), .Y(n_274) );
AND2x2_ASAP7_75t_R g750 ( .A(n_216), .B(n_725), .Y(n_750) );
CKINVDCx20_ASAP7_75t_R g693 ( .A(n_219), .Y(n_693) );
INVxp67_ASAP7_75t_L g279 ( .A(n_233), .Y(n_279) );
XNOR2x1_ASAP7_75t_L g473 ( .A(n_234), .B(n_474), .Y(n_473) );
INVx1_ASAP7_75t_L g519 ( .A(n_237), .Y(n_519) );
AOI22xp5_ASAP7_75t_L g378 ( .A1(n_238), .A2(n_266), .B1(n_292), .B2(n_305), .Y(n_378) );
AOI22xp33_ASAP7_75t_L g585 ( .A1(n_242), .A2(n_251), .B1(n_334), .B2(n_335), .Y(n_585) );
AOI22xp33_ASAP7_75t_L g680 ( .A1(n_255), .A2(n_260), .B1(n_292), .B2(n_681), .Y(n_680) );
CKINVDCx20_ASAP7_75t_R g698 ( .A(n_256), .Y(n_698) );
OA22x2_ASAP7_75t_L g343 ( .A1(n_264), .A2(n_344), .B1(n_345), .B2(n_379), .Y(n_343) );
INVx1_ASAP7_75t_L g379 ( .A(n_264), .Y(n_379) );
BUFx2_ASAP7_75t_L g271 ( .A(n_272), .Y(n_271) );
NOR2x1_ASAP7_75t_R g272 ( .A(n_273), .B(n_275), .Y(n_272) );
OR2x2_ASAP7_75t_L g780 ( .A(n_273), .B(n_276), .Y(n_780) );
INVx1_ASAP7_75t_L g273 ( .A(n_274), .Y(n_273) );
NOR2xp33_ASAP7_75t_L g724 ( .A(n_274), .B(n_725), .Y(n_724) );
INVx1_ASAP7_75t_L g275 ( .A(n_276), .Y(n_275) );
NOR2xp33_ASAP7_75t_L g276 ( .A(n_277), .B(n_278), .Y(n_276) );
AOI221xp5_ASAP7_75t_L g280 ( .A1(n_281), .A2(n_522), .B1(n_720), .B2(n_721), .C(n_722), .Y(n_280) );
INVx1_ASAP7_75t_L g721 ( .A(n_281), .Y(n_721) );
XNOR2xp5_ASAP7_75t_L g281 ( .A(n_282), .B(n_470), .Y(n_281) );
AOI22xp5_ASAP7_75t_L g282 ( .A1(n_283), .A2(n_284), .B1(n_382), .B2(n_469), .Y(n_282) );
INVx1_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
HB1xp67_ASAP7_75t_L g284 ( .A(n_285), .Y(n_284) );
OAI22xp33_ASAP7_75t_SL g285 ( .A1(n_286), .A2(n_343), .B1(n_380), .B2(n_381), .Y(n_285) );
INVx1_ASAP7_75t_L g380 ( .A(n_286), .Y(n_380) );
INVx2_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
NOR2x1_ASAP7_75t_L g289 ( .A(n_290), .B(n_328), .Y(n_289) );
NAND3xp33_ASAP7_75t_L g290 ( .A(n_291), .B(n_314), .C(n_323), .Y(n_290) );
AND2x2_ASAP7_75t_L g292 ( .A(n_293), .B(n_298), .Y(n_292) );
AND2x4_ASAP7_75t_L g393 ( .A(n_293), .B(n_298), .Y(n_393) );
AND2x2_ASAP7_75t_L g510 ( .A(n_293), .B(n_298), .Y(n_510) );
INVxp67_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
AND2x4_ASAP7_75t_L g308 ( .A(n_294), .B(n_309), .Y(n_308) );
AND2x4_ASAP7_75t_L g312 ( .A(n_294), .B(n_313), .Y(n_312) );
INVx2_ASAP7_75t_L g294 ( .A(n_295), .Y(n_294) );
AND2x2_ASAP7_75t_L g320 ( .A(n_295), .B(n_318), .Y(n_320) );
AND2x2_ASAP7_75t_L g326 ( .A(n_295), .B(n_309), .Y(n_326) );
INVx1_ASAP7_75t_L g297 ( .A(n_296), .Y(n_297) );
OAI22x1_ASAP7_75t_L g299 ( .A1(n_296), .A2(n_300), .B1(n_301), .B2(n_302), .Y(n_299) );
INVx1_ASAP7_75t_L g300 ( .A(n_296), .Y(n_300) );
INVx1_ASAP7_75t_L g304 ( .A(n_296), .Y(n_304) );
INVx2_ASAP7_75t_L g310 ( .A(n_296), .Y(n_310) );
AND2x4_ASAP7_75t_L g311 ( .A(n_298), .B(n_312), .Y(n_311) );
AND2x2_ASAP7_75t_L g315 ( .A(n_298), .B(n_316), .Y(n_315) );
AND2x2_ASAP7_75t_L g365 ( .A(n_298), .B(n_312), .Y(n_365) );
AND2x4_ASAP7_75t_L g371 ( .A(n_298), .B(n_316), .Y(n_371) );
AND2x2_ASAP7_75t_L g508 ( .A(n_298), .B(n_316), .Y(n_508) );
AND2x2_ASAP7_75t_L g298 ( .A(n_299), .B(n_303), .Y(n_298) );
INVx2_ASAP7_75t_L g307 ( .A(n_299), .Y(n_307) );
AND2x2_ASAP7_75t_L g321 ( .A(n_299), .B(n_322), .Y(n_321) );
HB1xp67_ASAP7_75t_L g325 ( .A(n_299), .Y(n_325) );
AND2x2_ASAP7_75t_L g306 ( .A(n_303), .B(n_307), .Y(n_306) );
INVx2_ASAP7_75t_L g322 ( .A(n_303), .Y(n_322) );
BUFx2_ASAP7_75t_L g338 ( .A(n_303), .Y(n_338) );
AND2x2_ASAP7_75t_L g305 ( .A(n_306), .B(n_308), .Y(n_305) );
AND2x6_ASAP7_75t_L g335 ( .A(n_306), .B(n_312), .Y(n_335) );
AND2x2_ASAP7_75t_L g339 ( .A(n_306), .B(n_320), .Y(n_339) );
AND2x2_ASAP7_75t_L g354 ( .A(n_306), .B(n_320), .Y(n_354) );
AND2x4_ASAP7_75t_L g390 ( .A(n_306), .B(n_308), .Y(n_390) );
AND2x2_ASAP7_75t_L g422 ( .A(n_306), .B(n_312), .Y(n_422) );
AND2x2_ASAP7_75t_L g681 ( .A(n_306), .B(n_308), .Y(n_681) );
AND2x4_ASAP7_75t_L g332 ( .A(n_307), .B(n_322), .Y(n_332) );
AND2x4_ASAP7_75t_L g327 ( .A(n_308), .B(n_321), .Y(n_327) );
AND2x2_ASAP7_75t_L g341 ( .A(n_308), .B(n_332), .Y(n_341) );
AND2x4_ASAP7_75t_L g349 ( .A(n_308), .B(n_332), .Y(n_349) );
AND2x2_ASAP7_75t_L g374 ( .A(n_308), .B(n_321), .Y(n_374) );
INVx1_ASAP7_75t_L g313 ( .A(n_309), .Y(n_313) );
INVx1_ASAP7_75t_L g318 ( .A(n_309), .Y(n_318) );
INVx2_ASAP7_75t_SL g502 ( .A(n_311), .Y(n_502) );
AND2x2_ASAP7_75t_L g330 ( .A(n_312), .B(n_321), .Y(n_330) );
AND2x2_ASAP7_75t_L g342 ( .A(n_312), .B(n_332), .Y(n_342) );
AND2x2_ASAP7_75t_L g351 ( .A(n_312), .B(n_321), .Y(n_351) );
AND2x4_ASAP7_75t_L g360 ( .A(n_312), .B(n_332), .Y(n_360) );
AND2x4_ASAP7_75t_L g414 ( .A(n_312), .B(n_321), .Y(n_414) );
INVx1_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
HB1xp67_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
AND2x4_ASAP7_75t_L g319 ( .A(n_320), .B(n_321), .Y(n_319) );
AND2x6_ASAP7_75t_L g334 ( .A(n_320), .B(n_332), .Y(n_334) );
AND2x2_ASAP7_75t_L g369 ( .A(n_320), .B(n_321), .Y(n_369) );
AND2x4_ASAP7_75t_L g425 ( .A(n_320), .B(n_332), .Y(n_425) );
AND2x2_ASAP7_75t_SL g324 ( .A(n_325), .B(n_326), .Y(n_324) );
AND2x2_ASAP7_75t_L g377 ( .A(n_325), .B(n_326), .Y(n_377) );
AND2x2_ASAP7_75t_SL g505 ( .A(n_325), .B(n_326), .Y(n_505) );
AND2x4_ASAP7_75t_L g331 ( .A(n_326), .B(n_332), .Y(n_331) );
AND2x4_ASAP7_75t_L g337 ( .A(n_326), .B(n_338), .Y(n_337) );
AND2x4_ASAP7_75t_L g356 ( .A(n_326), .B(n_338), .Y(n_356) );
AND2x4_ASAP7_75t_L g417 ( .A(n_326), .B(n_332), .Y(n_417) );
NAND4xp25_ASAP7_75t_L g328 ( .A(n_329), .B(n_333), .C(n_336), .D(n_340), .Y(n_328) );
INVx2_ASAP7_75t_L g381 ( .A(n_343), .Y(n_381) );
INVx1_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
NOR2xp67_ASAP7_75t_L g345 ( .A(n_346), .B(n_361), .Y(n_345) );
NAND3xp33_ASAP7_75t_L g346 ( .A(n_347), .B(n_352), .C(n_357), .Y(n_346) );
AND2x2_ASAP7_75t_L g347 ( .A(n_348), .B(n_350), .Y(n_347) );
BUFx3_ASAP7_75t_L g410 ( .A(n_349), .Y(n_410) );
INVx2_ASAP7_75t_L g454 ( .A(n_349), .Y(n_454) );
BUFx6f_ASAP7_75t_L g515 ( .A(n_349), .Y(n_515) );
BUFx6f_ASAP7_75t_L g717 ( .A(n_349), .Y(n_717) );
BUFx3_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
INVx2_ASAP7_75t_L g429 ( .A(n_354), .Y(n_429) );
BUFx6f_ASAP7_75t_L g456 ( .A(n_354), .Y(n_456) );
BUFx2_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
INVx5_ASAP7_75t_SL g431 ( .A(n_356), .Y(n_431) );
BUFx2_ASAP7_75t_L g768 ( .A(n_356), .Y(n_768) );
INVx3_ASAP7_75t_SL g358 ( .A(n_359), .Y(n_358) );
INVx2_ASAP7_75t_L g406 ( .A(n_359), .Y(n_406) );
INVx4_ASAP7_75t_L g461 ( .A(n_359), .Y(n_461) );
INVx3_ASAP7_75t_L g493 ( .A(n_359), .Y(n_493) );
INVx2_ASAP7_75t_SL g636 ( .A(n_359), .Y(n_636) );
INVx2_ASAP7_75t_SL g713 ( .A(n_359), .Y(n_713) );
INVx8_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
NAND4xp25_ASAP7_75t_L g361 ( .A(n_362), .B(n_366), .C(n_372), .D(n_378), .Y(n_361) );
INVx3_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
INVx3_ASAP7_75t_L g446 ( .A(n_364), .Y(n_446) );
INVx4_ASAP7_75t_SL g477 ( .A(n_364), .Y(n_477) );
INVx3_ASAP7_75t_SL g545 ( .A(n_364), .Y(n_545) );
INVx4_ASAP7_75t_SL g596 ( .A(n_364), .Y(n_596) );
INVx6_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
INVx2_ASAP7_75t_SL g552 ( .A(n_367), .Y(n_552) );
INVx4_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
INVx1_ASAP7_75t_L g401 ( .A(n_368), .Y(n_401) );
INVx2_ASAP7_75t_L g623 ( .A(n_368), .Y(n_623) );
INVx3_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
BUFx6f_ASAP7_75t_L g482 ( .A(n_369), .Y(n_482) );
BUFx6f_ASAP7_75t_L g741 ( .A(n_369), .Y(n_741) );
BUFx2_ASAP7_75t_SL g402 ( .A(n_370), .Y(n_402) );
BUFx6f_ASAP7_75t_SL g370 ( .A(n_371), .Y(n_370) );
INVx2_ASAP7_75t_L g441 ( .A(n_371), .Y(n_441) );
INVx1_ASAP7_75t_L g484 ( .A(n_371), .Y(n_484) );
BUFx3_ASAP7_75t_L g563 ( .A(n_371), .Y(n_563) );
BUFx4f_ASAP7_75t_L g742 ( .A(n_371), .Y(n_742) );
BUFx3_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
BUFx3_ASAP7_75t_L g397 ( .A(n_374), .Y(n_397) );
INVx2_ASAP7_75t_L g448 ( .A(n_374), .Y(n_448) );
BUFx5_ASAP7_75t_L g760 ( .A(n_374), .Y(n_760) );
BUFx6f_ASAP7_75t_L g398 ( .A(n_375), .Y(n_398) );
INVx3_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
INVx2_ASAP7_75t_L g591 ( .A(n_376), .Y(n_591) );
INVx3_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
BUFx12f_ASAP7_75t_L g626 ( .A(n_377), .Y(n_626) );
INVx1_ASAP7_75t_L g469 ( .A(n_382), .Y(n_469) );
AOI22xp33_ASAP7_75t_SL g382 ( .A1(n_383), .A2(n_384), .B1(n_435), .B2(n_468), .Y(n_382) );
INVx1_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
NAND3xp33_ASAP7_75t_L g385 ( .A(n_386), .B(n_403), .C(n_418), .Y(n_385) );
NOR2xp33_ASAP7_75t_L g386 ( .A(n_387), .B(n_394), .Y(n_386) );
NOR4xp25_ASAP7_75t_L g432 ( .A(n_387), .B(n_394), .C(n_404), .D(n_433), .Y(n_432) );
BUFx2_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
BUFx4f_ASAP7_75t_SL g547 ( .A(n_389), .Y(n_547) );
BUFx6f_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
BUFx3_ASAP7_75t_L g443 ( .A(n_390), .Y(n_443) );
BUFx2_ASAP7_75t_L g480 ( .A(n_390), .Y(n_480) );
INVx2_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
INVx2_ASAP7_75t_SL g444 ( .A(n_392), .Y(n_444) );
INVx2_ASAP7_75t_L g548 ( .A(n_392), .Y(n_548) );
INVx2_ASAP7_75t_L g629 ( .A(n_392), .Y(n_629) );
OAI22xp33_ASAP7_75t_L g701 ( .A1(n_392), .A2(n_702), .B1(n_703), .B2(n_704), .Y(n_701) );
INVx6_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
NAND2xp5_ASAP7_75t_L g394 ( .A(n_395), .B(n_399), .Y(n_394) );
BUFx6f_ASAP7_75t_SL g396 ( .A(n_397), .Y(n_396) );
INVx1_ASAP7_75t_L g695 ( .A(n_397), .Y(n_695) );
INVx1_ASAP7_75t_L g699 ( .A(n_400), .Y(n_699) );
BUFx3_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
INVxp67_ASAP7_75t_SL g403 ( .A(n_404), .Y(n_403) );
OAI221xp5_ASAP7_75t_SL g404 ( .A1(n_405), .A2(n_407), .B1(n_408), .B2(n_411), .C(n_412), .Y(n_404) );
INVx1_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
INVx1_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
BUFx2_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
BUFx3_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
INVx6_ASAP7_75t_L g452 ( .A(n_414), .Y(n_452) );
BUFx3_ASAP7_75t_L g488 ( .A(n_414), .Y(n_488) );
BUFx6f_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
BUFx3_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
BUFx2_ASAP7_75t_SL g462 ( .A(n_417), .Y(n_462) );
BUFx3_ASAP7_75t_L g489 ( .A(n_417), .Y(n_489) );
BUFx2_ASAP7_75t_SL g534 ( .A(n_417), .Y(n_534) );
INVx2_ASAP7_75t_L g642 ( .A(n_417), .Y(n_642) );
NAND2xp5_ASAP7_75t_SL g433 ( .A(n_418), .B(n_434), .Y(n_433) );
AND2x2_ASAP7_75t_L g418 ( .A(n_419), .B(n_426), .Y(n_418) );
INVx3_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
INVx2_ASAP7_75t_SL g464 ( .A(n_421), .Y(n_464) );
INVx2_ASAP7_75t_L g633 ( .A(n_421), .Y(n_633) );
INVx2_ASAP7_75t_SL g772 ( .A(n_421), .Y(n_772) );
INVx3_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
BUFx2_ASAP7_75t_L g571 ( .A(n_422), .Y(n_571) );
BUFx2_ASAP7_75t_L g663 ( .A(n_422), .Y(n_663) );
INVx2_ASAP7_75t_SL g423 ( .A(n_424), .Y(n_423) );
INVx1_ASAP7_75t_SL g465 ( .A(n_424), .Y(n_465) );
INVx2_ASAP7_75t_L g494 ( .A(n_424), .Y(n_494) );
INVx2_ASAP7_75t_L g540 ( .A(n_424), .Y(n_540) );
INVx2_ASAP7_75t_L g572 ( .A(n_424), .Y(n_572) );
INVx2_ASAP7_75t_L g634 ( .A(n_424), .Y(n_634) );
INVx2_ASAP7_75t_L g664 ( .A(n_424), .Y(n_664) );
INVx8_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
BUFx6f_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
INVx1_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
INVx1_ASAP7_75t_L g638 ( .A(n_429), .Y(n_638) );
INVx2_ASAP7_75t_L g710 ( .A(n_429), .Y(n_710) );
INVx2_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
INVx3_ASAP7_75t_L g457 ( .A(n_431), .Y(n_457) );
INVx2_ASAP7_75t_L g531 ( .A(n_431), .Y(n_531) );
INVx2_ASAP7_75t_L g661 ( .A(n_431), .Y(n_661) );
INVx2_ASAP7_75t_SL g435 ( .A(n_436), .Y(n_435) );
HB1xp67_ASAP7_75t_L g468 ( .A(n_436), .Y(n_468) );
INVx1_ASAP7_75t_SL g466 ( .A(n_437), .Y(n_466) );
NOR4xp75_ASAP7_75t_L g437 ( .A(n_438), .B(n_445), .C(n_449), .D(n_458), .Y(n_437) );
NAND2xp5_ASAP7_75t_L g438 ( .A(n_439), .B(n_442), .Y(n_438) );
INVx2_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
BUFx2_ASAP7_75t_L g554 ( .A(n_441), .Y(n_554) );
INVx2_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
INVx1_ASAP7_75t_L g625 ( .A(n_448), .Y(n_625) );
NAND2xp5_ASAP7_75t_L g449 ( .A(n_450), .B(n_455), .Y(n_449) );
INVx2_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
INVx2_ASAP7_75t_L g533 ( .A(n_452), .Y(n_533) );
INVx1_ASAP7_75t_SL g578 ( .A(n_452), .Y(n_578) );
INVx2_ASAP7_75t_L g640 ( .A(n_452), .Y(n_640) );
INVx1_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
INVx1_ASAP7_75t_L g491 ( .A(n_454), .Y(n_491) );
NAND2xp5_ASAP7_75t_L g458 ( .A(n_459), .B(n_463), .Y(n_458) );
BUFx6f_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
INVx2_ASAP7_75t_L g537 ( .A(n_461), .Y(n_537) );
OAI22xp5_ASAP7_75t_L g470 ( .A1(n_471), .A2(n_495), .B1(n_520), .B2(n_521), .Y(n_470) );
INVx2_ASAP7_75t_L g520 ( .A(n_471), .Y(n_520) );
BUFx3_ASAP7_75t_L g471 ( .A(n_472), .Y(n_471) );
INVx1_ASAP7_75t_L g472 ( .A(n_473), .Y(n_472) );
OR2x2_ASAP7_75t_L g474 ( .A(n_475), .B(n_485), .Y(n_474) );
NAND4xp25_ASAP7_75t_L g475 ( .A(n_476), .B(n_478), .C(n_479), .D(n_481), .Y(n_475) );
INVx2_ASAP7_75t_SL g483 ( .A(n_484), .Y(n_483) );
NAND4xp25_ASAP7_75t_L g485 ( .A(n_486), .B(n_487), .C(n_490), .D(n_492), .Y(n_485) );
INVx1_ASAP7_75t_L g521 ( .A(n_495), .Y(n_521) );
INVx1_ASAP7_75t_L g495 ( .A(n_496), .Y(n_495) );
INVx2_ASAP7_75t_L g496 ( .A(n_497), .Y(n_496) );
INVx1_ASAP7_75t_L g497 ( .A(n_498), .Y(n_497) );
XOR2x2_ASAP7_75t_L g498 ( .A(n_499), .B(n_519), .Y(n_498) );
NAND2x1_ASAP7_75t_L g499 ( .A(n_500), .B(n_511), .Y(n_499) );
NOR2xp33_ASAP7_75t_L g500 ( .A(n_501), .B(n_506), .Y(n_500) );
OAI21xp5_ASAP7_75t_SL g501 ( .A1(n_502), .A2(n_503), .B(n_504), .Y(n_501) );
NAND2xp5_ASAP7_75t_L g506 ( .A(n_507), .B(n_509), .Y(n_506) );
NOR2x1_ASAP7_75t_L g511 ( .A(n_512), .B(n_516), .Y(n_511) );
NAND2xp5_ASAP7_75t_L g512 ( .A(n_513), .B(n_514), .Y(n_512) );
BUFx6f_ASAP7_75t_L g538 ( .A(n_515), .Y(n_538) );
INVx2_ASAP7_75t_L g576 ( .A(n_515), .Y(n_576) );
NAND2xp5_ASAP7_75t_L g516 ( .A(n_517), .B(n_518), .Y(n_516) );
INVxp67_ASAP7_75t_SL g720 ( .A(n_522), .Y(n_720) );
XOR2xp5_ASAP7_75t_L g522 ( .A(n_523), .B(n_597), .Y(n_522) );
AOI22xp5_ASAP7_75t_L g523 ( .A1(n_524), .A2(n_525), .B1(n_555), .B2(n_556), .Y(n_523) );
INVx2_ASAP7_75t_SL g524 ( .A(n_525), .Y(n_524) );
INVx1_ASAP7_75t_L g527 ( .A(n_528), .Y(n_527) );
NOR2x1_ASAP7_75t_L g528 ( .A(n_529), .B(n_541), .Y(n_528) );
NAND4xp25_ASAP7_75t_L g529 ( .A(n_530), .B(n_532), .C(n_535), .D(n_539), .Y(n_529) );
INVx1_ASAP7_75t_L g536 ( .A(n_537), .Y(n_536) );
NAND4xp25_ASAP7_75t_SL g541 ( .A(n_542), .B(n_546), .C(n_549), .D(n_550), .Y(n_541) );
INVx2_ASAP7_75t_L g543 ( .A(n_544), .Y(n_543) );
OAI21xp33_ASAP7_75t_SL g652 ( .A1(n_544), .A2(n_653), .B(n_654), .Y(n_652) );
OAI221xp5_ASAP7_75t_L g692 ( .A1(n_544), .A2(n_693), .B1(n_694), .B2(n_695), .C(n_696), .Y(n_692) );
INVx2_ASAP7_75t_L g544 ( .A(n_545), .Y(n_544) );
INVx1_ASAP7_75t_L g703 ( .A(n_547), .Y(n_703) );
INVx1_ASAP7_75t_L g551 ( .A(n_552), .Y(n_551) );
INVx3_ASAP7_75t_L g553 ( .A(n_554), .Y(n_553) );
OAI22xp5_ASAP7_75t_L g697 ( .A1(n_554), .A2(n_698), .B1(n_699), .B2(n_700), .Y(n_697) );
INVx1_ASAP7_75t_L g555 ( .A(n_556), .Y(n_555) );
OAI22xp5_ASAP7_75t_SL g556 ( .A1(n_557), .A2(n_558), .B1(n_579), .B2(n_580), .Y(n_556) );
INVx4_ASAP7_75t_L g557 ( .A(n_558), .Y(n_557) );
NOR2x1_ASAP7_75t_L g559 ( .A(n_560), .B(n_567), .Y(n_559) );
NAND4xp25_ASAP7_75t_L g560 ( .A(n_561), .B(n_564), .C(n_565), .D(n_566), .Y(n_560) );
BUFx6f_ASAP7_75t_SL g562 ( .A(n_563), .Y(n_562) );
NAND4xp25_ASAP7_75t_L g567 ( .A(n_568), .B(n_573), .C(n_574), .D(n_577), .Y(n_567) );
INVx2_ASAP7_75t_L g569 ( .A(n_570), .Y(n_569) );
INVx2_ASAP7_75t_L g570 ( .A(n_571), .Y(n_570) );
INVx2_ASAP7_75t_L g575 ( .A(n_576), .Y(n_575) );
INVx1_ASAP7_75t_SL g579 ( .A(n_580), .Y(n_579) );
INVx1_ASAP7_75t_L g580 ( .A(n_581), .Y(n_580) );
OAI22xp5_ASAP7_75t_L g688 ( .A1(n_581), .A2(n_582), .B1(n_689), .B2(n_718), .Y(n_688) );
INVx2_ASAP7_75t_L g581 ( .A(n_582), .Y(n_581) );
NOR3xp33_ASAP7_75t_L g583 ( .A(n_584), .B(n_589), .C(n_593), .Y(n_583) );
NAND4xp25_ASAP7_75t_L g584 ( .A(n_585), .B(n_586), .C(n_587), .D(n_588), .Y(n_584) );
NAND2xp5_ASAP7_75t_L g589 ( .A(n_590), .B(n_592), .Y(n_589) );
NAND2xp5_ASAP7_75t_L g593 ( .A(n_594), .B(n_595), .Y(n_593) );
INVx1_ASAP7_75t_SL g757 ( .A(n_596), .Y(n_757) );
OAI22xp5_ASAP7_75t_L g597 ( .A1(n_598), .A2(n_644), .B1(n_645), .B2(n_719), .Y(n_597) );
INVx1_ASAP7_75t_L g719 ( .A(n_598), .Y(n_719) );
INVx1_ASAP7_75t_L g598 ( .A(n_599), .Y(n_598) );
INVx1_ASAP7_75t_L g599 ( .A(n_600), .Y(n_599) );
OAI22xp5_ASAP7_75t_L g600 ( .A1(n_601), .A2(n_618), .B1(n_619), .B2(n_643), .Y(n_600) );
INVx3_ASAP7_75t_SL g643 ( .A(n_601), .Y(n_643) );
XOR2x2_ASAP7_75t_L g601 ( .A(n_602), .B(n_617), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g602 ( .A(n_603), .B(n_610), .Y(n_602) );
NOR2xp33_ASAP7_75t_L g603 ( .A(n_604), .B(n_607), .Y(n_603) );
NAND2xp5_ASAP7_75t_SL g604 ( .A(n_605), .B(n_606), .Y(n_604) );
NAND2xp5_ASAP7_75t_L g607 ( .A(n_608), .B(n_609), .Y(n_607) );
NOR2xp33_ASAP7_75t_L g610 ( .A(n_611), .B(n_614), .Y(n_610) );
NAND2xp5_ASAP7_75t_L g611 ( .A(n_612), .B(n_613), .Y(n_611) );
NAND2xp5_ASAP7_75t_L g614 ( .A(n_615), .B(n_616), .Y(n_614) );
INVx1_ASAP7_75t_SL g618 ( .A(n_619), .Y(n_618) );
NAND2xp5_ASAP7_75t_L g620 ( .A(n_621), .B(n_631), .Y(n_620) );
NOR3xp33_ASAP7_75t_L g621 ( .A(n_622), .B(n_624), .C(n_627), .Y(n_621) );
NAND2xp5_ASAP7_75t_SL g627 ( .A(n_628), .B(n_630), .Y(n_627) );
AND4x1_ASAP7_75t_L g631 ( .A(n_632), .B(n_635), .C(n_637), .D(n_639), .Y(n_631) );
INVx2_ASAP7_75t_SL g641 ( .A(n_642), .Y(n_641) );
INVx1_ASAP7_75t_L g644 ( .A(n_645), .Y(n_644) );
AOI22xp5_ASAP7_75t_L g645 ( .A1(n_646), .A2(n_647), .B1(n_686), .B2(n_687), .Y(n_645) );
INVx1_ASAP7_75t_SL g646 ( .A(n_647), .Y(n_646) );
INVx1_ASAP7_75t_L g647 ( .A(n_648), .Y(n_647) );
OAI22x1_ASAP7_75t_L g648 ( .A1(n_649), .A2(n_669), .B1(n_670), .B2(n_685), .Y(n_648) );
INVx2_ASAP7_75t_L g685 ( .A(n_649), .Y(n_685) );
XNOR2x1_ASAP7_75t_L g649 ( .A(n_650), .B(n_668), .Y(n_649) );
AND2x2_ASAP7_75t_L g650 ( .A(n_651), .B(n_658), .Y(n_650) );
NOR2xp33_ASAP7_75t_L g651 ( .A(n_652), .B(n_655), .Y(n_651) );
NAND2xp5_ASAP7_75t_L g655 ( .A(n_656), .B(n_657), .Y(n_655) );
NOR2xp33_ASAP7_75t_L g658 ( .A(n_659), .B(n_665), .Y(n_658) );
NAND2xp5_ASAP7_75t_L g659 ( .A(n_660), .B(n_662), .Y(n_659) );
NAND2xp5_ASAP7_75t_L g665 ( .A(n_666), .B(n_667), .Y(n_665) );
INVx3_ASAP7_75t_L g669 ( .A(n_670), .Y(n_669) );
INVx1_ASAP7_75t_L g684 ( .A(n_671), .Y(n_684) );
NOR2xp67_ASAP7_75t_L g671 ( .A(n_672), .B(n_677), .Y(n_671) );
NAND4xp25_ASAP7_75t_L g672 ( .A(n_673), .B(n_674), .C(n_675), .D(n_676), .Y(n_672) );
NAND4xp25_ASAP7_75t_SL g677 ( .A(n_678), .B(n_679), .C(n_680), .D(n_682), .Y(n_677) );
INVx1_ASAP7_75t_SL g686 ( .A(n_687), .Y(n_686) );
INVx1_ASAP7_75t_L g687 ( .A(n_688), .Y(n_687) );
INVx1_ASAP7_75t_L g718 ( .A(n_689), .Y(n_718) );
NAND2xp5_ASAP7_75t_L g690 ( .A(n_691), .B(n_705), .Y(n_690) );
NOR3xp33_ASAP7_75t_L g691 ( .A(n_692), .B(n_697), .C(n_701), .Y(n_691) );
NOR2xp33_ASAP7_75t_L g705 ( .A(n_706), .B(n_711), .Y(n_705) );
NAND2xp5_ASAP7_75t_L g706 ( .A(n_707), .B(n_708), .Y(n_706) );
BUFx6f_ASAP7_75t_L g709 ( .A(n_710), .Y(n_709) );
NAND2xp5_ASAP7_75t_L g711 ( .A(n_712), .B(n_714), .Y(n_711) );
INVx1_ASAP7_75t_L g715 ( .A(n_716), .Y(n_715) );
INVx1_ASAP7_75t_L g716 ( .A(n_717), .Y(n_716) );
INVx1_ASAP7_75t_SL g722 ( .A(n_723), .Y(n_722) );
AND2x2_ASAP7_75t_L g723 ( .A(n_724), .B(n_726), .Y(n_723) );
NAND2xp5_ASAP7_75t_L g777 ( .A(n_724), .B(n_727), .Y(n_777) );
INVx1_ASAP7_75t_L g726 ( .A(n_727), .Y(n_726) );
NAND2xp5_ASAP7_75t_L g728 ( .A(n_729), .B(n_730), .Y(n_728) );
OAI222xp33_ASAP7_75t_L g731 ( .A1(n_732), .A2(n_749), .B1(n_751), .B2(n_773), .C1(n_778), .C2(n_781), .Y(n_731) );
INVx1_ASAP7_75t_L g733 ( .A(n_734), .Y(n_733) );
HB1xp67_ASAP7_75t_L g734 ( .A(n_735), .Y(n_734) );
NAND4xp75_ASAP7_75t_SL g735 ( .A(n_736), .B(n_739), .C(n_744), .D(n_747), .Y(n_735) );
AND2x2_ASAP7_75t_L g736 ( .A(n_737), .B(n_738), .Y(n_736) );
AND2x2_ASAP7_75t_L g739 ( .A(n_740), .B(n_743), .Y(n_739) );
AND2x2_ASAP7_75t_L g744 ( .A(n_745), .B(n_746), .Y(n_744) );
INVx1_ASAP7_75t_L g749 ( .A(n_750), .Y(n_749) );
INVx1_ASAP7_75t_L g751 ( .A(n_752), .Y(n_751) );
HB1xp67_ASAP7_75t_L g752 ( .A(n_753), .Y(n_752) );
AND2x2_ASAP7_75t_L g754 ( .A(n_755), .B(n_764), .Y(n_754) );
NOR2xp33_ASAP7_75t_L g755 ( .A(n_756), .B(n_761), .Y(n_755) );
OAI21xp33_ASAP7_75t_L g756 ( .A1(n_757), .A2(n_758), .B(n_759), .Y(n_756) );
NAND2xp5_ASAP7_75t_L g761 ( .A(n_762), .B(n_763), .Y(n_761) );
NOR2xp33_ASAP7_75t_L g764 ( .A(n_765), .B(n_769), .Y(n_764) );
NAND2xp5_ASAP7_75t_L g765 ( .A(n_766), .B(n_767), .Y(n_765) );
NAND2xp5_ASAP7_75t_L g769 ( .A(n_770), .B(n_771), .Y(n_769) );
CKINVDCx20_ASAP7_75t_R g773 ( .A(n_774), .Y(n_773) );
CKINVDCx20_ASAP7_75t_R g774 ( .A(n_775), .Y(n_774) );
CKINVDCx20_ASAP7_75t_R g775 ( .A(n_776), .Y(n_775) );
CKINVDCx6p67_ASAP7_75t_R g776 ( .A(n_777), .Y(n_776) );
CKINVDCx20_ASAP7_75t_R g778 ( .A(n_779), .Y(n_778) );
CKINVDCx20_ASAP7_75t_R g779 ( .A(n_780), .Y(n_779) );
endmodule