module real_aes_467_n_98 (n_17, n_28, n_76, n_56, n_34, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_43, n_96, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_98);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_98;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_564;
wire n_519;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_178;
wire n_409;
wire n_748;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_449;
wire n_182;
wire n_363;
wire n_417;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_527;
wire n_434;
wire n_502;
wire n_505;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_404;
wire n_288;
wire n_598;
wire n_713;
wire n_735;
wire n_728;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_101;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_633;
wire n_520;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_420;
wire n_336;
wire n_349;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_314;
wire n_283;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_717;
wire n_456;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_99;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_719;
wire n_465;
wire n_473;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_743;
wire n_105;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
NAND2xp5_ASAP7_75t_SL g452 ( .A(n_0), .B(n_138), .Y(n_452) );
AOI21xp5_ASAP7_75t_L g482 ( .A1(n_1), .A2(n_146), .B(n_483), .Y(n_482) );
NAND2xp5_ASAP7_75t_L g730 ( .A(n_2), .B(n_731), .Y(n_730) );
NAND2xp5_ASAP7_75t_L g215 ( .A(n_3), .B(n_138), .Y(n_215) );
NAND2xp5_ASAP7_75t_L g177 ( .A(n_4), .B(n_165), .Y(n_177) );
NAND2xp5_ASAP7_75t_SL g463 ( .A(n_5), .B(n_165), .Y(n_463) );
INVx1_ASAP7_75t_L g134 ( .A(n_6), .Y(n_134) );
NAND2xp5_ASAP7_75t_L g492 ( .A(n_7), .B(n_165), .Y(n_492) );
CKINVDCx16_ASAP7_75t_R g731 ( .A(n_8), .Y(n_731) );
NAND2xp33_ASAP7_75t_L g533 ( .A(n_9), .B(n_163), .Y(n_533) );
AND2x2_ASAP7_75t_L g168 ( .A(n_10), .B(n_169), .Y(n_168) );
AND2x2_ASAP7_75t_L g179 ( .A(n_11), .B(n_180), .Y(n_179) );
INVx2_ASAP7_75t_L g125 ( .A(n_12), .Y(n_125) );
AOI221x1_ASAP7_75t_L g438 ( .A1(n_13), .A2(n_24), .B1(n_138), .B2(n_146), .C(n_439), .Y(n_438) );
NAND2xp5_ASAP7_75t_L g234 ( .A(n_14), .B(n_165), .Y(n_234) );
CKINVDCx16_ASAP7_75t_R g107 ( .A(n_15), .Y(n_107) );
NAND2xp5_ASAP7_75t_SL g529 ( .A(n_16), .B(n_138), .Y(n_529) );
AO21x2_ASAP7_75t_L g527 ( .A1(n_17), .A2(n_180), .B(n_528), .Y(n_527) );
NAND2xp5_ASAP7_75t_L g442 ( .A(n_18), .B(n_123), .Y(n_442) );
NAND2xp5_ASAP7_75t_L g516 ( .A(n_19), .B(n_165), .Y(n_516) );
AO21x1_ASAP7_75t_L g458 ( .A1(n_20), .A2(n_138), .B(n_459), .Y(n_458) );
NAND2xp5_ASAP7_75t_SL g219 ( .A(n_21), .B(n_138), .Y(n_219) );
INVx1_ASAP7_75t_L g110 ( .A(n_22), .Y(n_110) );
AOI22xp33_ASAP7_75t_L g128 ( .A1(n_23), .A2(n_87), .B1(n_129), .B2(n_138), .Y(n_128) );
NAND2x1_ASAP7_75t_L g450 ( .A(n_25), .B(n_165), .Y(n_450) );
NAND2x1_ASAP7_75t_L g491 ( .A(n_26), .B(n_163), .Y(n_491) );
OR2x2_ASAP7_75t_L g126 ( .A(n_27), .B(n_84), .Y(n_126) );
OA21x2_ASAP7_75t_L g158 ( .A1(n_27), .A2(n_84), .B(n_125), .Y(n_158) );
NAND2xp5_ASAP7_75t_L g485 ( .A(n_28), .B(n_163), .Y(n_485) );
NAND2xp5_ASAP7_75t_L g532 ( .A(n_29), .B(n_165), .Y(n_532) );
AO21x2_ASAP7_75t_L g229 ( .A1(n_30), .A2(n_169), .B(n_230), .Y(n_229) );
NAND2xp5_ASAP7_75t_L g462 ( .A(n_31), .B(n_163), .Y(n_462) );
AOI21xp5_ASAP7_75t_L g174 ( .A1(n_32), .A2(n_146), .B(n_175), .Y(n_174) );
NAND2xp5_ASAP7_75t_L g214 ( .A(n_33), .B(n_165), .Y(n_214) );
AOI21xp5_ASAP7_75t_L g469 ( .A1(n_34), .A2(n_146), .B(n_470), .Y(n_469) );
AND2x2_ASAP7_75t_L g136 ( .A(n_35), .B(n_137), .Y(n_136) );
AND2x2_ASAP7_75t_L g144 ( .A(n_35), .B(n_134), .Y(n_144) );
INVx1_ASAP7_75t_L g150 ( .A(n_35), .Y(n_150) );
OR2x6_ASAP7_75t_L g108 ( .A(n_36), .B(n_109), .Y(n_108) );
NAND2xp5_ASAP7_75t_SL g473 ( .A(n_37), .B(n_138), .Y(n_473) );
NAND2xp5_ASAP7_75t_L g178 ( .A(n_38), .B(n_138), .Y(n_178) );
NAND2xp5_ASAP7_75t_L g204 ( .A(n_39), .B(n_165), .Y(n_204) );
CKINVDCx20_ASAP7_75t_R g520 ( .A(n_40), .Y(n_520) );
NAND2xp5_ASAP7_75t_L g471 ( .A(n_41), .B(n_163), .Y(n_471) );
NAND2xp5_ASAP7_75t_L g187 ( .A(n_42), .B(n_138), .Y(n_187) );
AOI21xp5_ASAP7_75t_L g160 ( .A1(n_43), .A2(n_146), .B(n_161), .Y(n_160) );
AOI21xp5_ASAP7_75t_L g489 ( .A1(n_44), .A2(n_146), .B(n_490), .Y(n_489) );
NAND2xp5_ASAP7_75t_L g191 ( .A(n_45), .B(n_163), .Y(n_191) );
NAND2xp5_ASAP7_75t_L g451 ( .A(n_46), .B(n_163), .Y(n_451) );
NAND2xp5_ASAP7_75t_SL g231 ( .A(n_47), .B(n_138), .Y(n_231) );
INVx1_ASAP7_75t_L g132 ( .A(n_48), .Y(n_132) );
INVx1_ASAP7_75t_L g141 ( .A(n_48), .Y(n_141) );
NAND2xp5_ASAP7_75t_L g164 ( .A(n_49), .B(n_165), .Y(n_164) );
AND2x2_ASAP7_75t_L g199 ( .A(n_50), .B(n_123), .Y(n_199) );
NAND2xp5_ASAP7_75t_L g162 ( .A(n_51), .B(n_163), .Y(n_162) );
CKINVDCx20_ASAP7_75t_R g742 ( .A(n_52), .Y(n_742) );
NAND2xp5_ASAP7_75t_L g441 ( .A(n_53), .B(n_165), .Y(n_441) );
NAND2xp5_ASAP7_75t_L g213 ( .A(n_54), .B(n_163), .Y(n_213) );
AOI21xp5_ASAP7_75t_L g448 ( .A1(n_55), .A2(n_146), .B(n_449), .Y(n_448) );
NAND2xp5_ASAP7_75t_SL g167 ( .A(n_56), .B(n_138), .Y(n_167) );
AOI222xp33_ASAP7_75t_L g98 ( .A1(n_57), .A2(n_99), .B1(n_724), .B2(n_735), .C1(n_743), .C2(n_745), .Y(n_98) );
OAI22xp5_ASAP7_75t_L g737 ( .A1(n_57), .A2(n_112), .B1(n_719), .B2(n_738), .Y(n_737) );
CKINVDCx20_ASAP7_75t_R g738 ( .A(n_57), .Y(n_738) );
NAND2xp5_ASAP7_75t_SL g201 ( .A(n_58), .B(n_138), .Y(n_201) );
AOI21xp5_ASAP7_75t_L g211 ( .A1(n_59), .A2(n_146), .B(n_212), .Y(n_211) );
AND2x2_ASAP7_75t_L g225 ( .A(n_60), .B(n_124), .Y(n_225) );
AO21x1_ASAP7_75t_L g460 ( .A1(n_61), .A2(n_146), .B(n_461), .Y(n_460) );
NAND2xp5_ASAP7_75t_SL g481 ( .A(n_62), .B(n_138), .Y(n_481) );
NAND2xp5_ASAP7_75t_L g205 ( .A(n_63), .B(n_163), .Y(n_205) );
NAND2xp5_ASAP7_75t_SL g493 ( .A(n_64), .B(n_138), .Y(n_493) );
NAND2xp5_ASAP7_75t_L g235 ( .A(n_65), .B(n_163), .Y(n_235) );
AOI22xp5_ASAP7_75t_L g145 ( .A1(n_66), .A2(n_91), .B1(n_146), .B2(n_148), .Y(n_145) );
NAND2xp5_ASAP7_75t_L g222 ( .A(n_67), .B(n_165), .Y(n_222) );
AND2x2_ASAP7_75t_L g474 ( .A(n_68), .B(n_124), .Y(n_474) );
INVx1_ASAP7_75t_L g137 ( .A(n_69), .Y(n_137) );
INVx1_ASAP7_75t_L g143 ( .A(n_69), .Y(n_143) );
AND2x2_ASAP7_75t_L g494 ( .A(n_70), .B(n_169), .Y(n_494) );
NAND2xp5_ASAP7_75t_L g176 ( .A(n_71), .B(n_163), .Y(n_176) );
AOI21xp5_ASAP7_75t_L g202 ( .A1(n_72), .A2(n_146), .B(n_203), .Y(n_202) );
AOI21xp5_ASAP7_75t_L g188 ( .A1(n_73), .A2(n_146), .B(n_189), .Y(n_188) );
AOI21xp5_ASAP7_75t_L g232 ( .A1(n_74), .A2(n_146), .B(n_233), .Y(n_232) );
AND2x2_ASAP7_75t_L g216 ( .A(n_75), .B(n_124), .Y(n_216) );
NAND2xp5_ASAP7_75t_SL g122 ( .A(n_76), .B(n_123), .Y(n_122) );
INVx1_ASAP7_75t_L g111 ( .A(n_77), .Y(n_111) );
AND2x2_ASAP7_75t_L g479 ( .A(n_78), .B(n_169), .Y(n_479) );
NAND2xp5_ASAP7_75t_SL g518 ( .A(n_79), .B(n_138), .Y(n_518) );
AND2x2_ASAP7_75t_L g192 ( .A(n_80), .B(n_180), .Y(n_192) );
AOI22xp33_ASAP7_75t_L g716 ( .A1(n_81), .A2(n_100), .B1(n_717), .B2(n_722), .Y(n_716) );
AND2x2_ASAP7_75t_L g459 ( .A(n_82), .B(n_206), .Y(n_459) );
INVx1_ASAP7_75t_L g100 ( .A(n_83), .Y(n_100) );
AND2x2_ASAP7_75t_L g453 ( .A(n_85), .B(n_169), .Y(n_453) );
NAND2xp5_ASAP7_75t_L g517 ( .A(n_86), .B(n_163), .Y(n_517) );
NAND2xp5_ASAP7_75t_L g472 ( .A(n_88), .B(n_165), .Y(n_472) );
NAND2xp5_ASAP7_75t_L g440 ( .A(n_89), .B(n_163), .Y(n_440) );
AOI21xp5_ASAP7_75t_L g514 ( .A1(n_90), .A2(n_146), .B(n_515), .Y(n_514) );
AOI21xp5_ASAP7_75t_L g220 ( .A1(n_92), .A2(n_146), .B(n_221), .Y(n_220) );
NAND2xp5_ASAP7_75t_L g190 ( .A(n_93), .B(n_165), .Y(n_190) );
NAND2xp5_ASAP7_75t_L g484 ( .A(n_94), .B(n_165), .Y(n_484) );
BUFx2_ASAP7_75t_L g224 ( .A(n_95), .Y(n_224) );
BUFx2_ASAP7_75t_L g732 ( .A(n_96), .Y(n_732) );
BUFx2_ASAP7_75t_SL g749 ( .A(n_96), .Y(n_749) );
AOI21xp5_ASAP7_75t_L g530 ( .A1(n_97), .A2(n_146), .B(n_531), .Y(n_530) );
OAI21xp5_ASAP7_75t_L g99 ( .A1(n_100), .A2(n_101), .B(n_716), .Y(n_99) );
INVx1_ASAP7_75t_L g101 ( .A(n_102), .Y(n_101) );
OAI22xp5_ASAP7_75t_L g102 ( .A1(n_103), .A2(n_112), .B1(n_431), .B2(n_711), .Y(n_102) );
CKINVDCx6p67_ASAP7_75t_R g103 ( .A(n_104), .Y(n_103) );
CKINVDCx11_ASAP7_75t_R g718 ( .A(n_104), .Y(n_718) );
INVx3_ASAP7_75t_SL g104 ( .A(n_105), .Y(n_104) );
CKINVDCx5p33_ASAP7_75t_R g105 ( .A(n_106), .Y(n_105) );
AND2x6_ASAP7_75t_SL g106 ( .A(n_107), .B(n_108), .Y(n_106) );
OR2x6_ASAP7_75t_SL g714 ( .A(n_107), .B(n_715), .Y(n_714) );
OR2x2_ASAP7_75t_L g723 ( .A(n_107), .B(n_108), .Y(n_723) );
NAND2xp5_ASAP7_75t_L g734 ( .A(n_107), .B(n_715), .Y(n_734) );
CKINVDCx5p33_ASAP7_75t_R g715 ( .A(n_108), .Y(n_715) );
NAND2xp5_ASAP7_75t_L g109 ( .A(n_110), .B(n_111), .Y(n_109) );
INVx4_ASAP7_75t_L g719 ( .A(n_112), .Y(n_719) );
OR2x6_ASAP7_75t_L g112 ( .A(n_113), .B(n_368), .Y(n_112) );
NAND3xp33_ASAP7_75t_L g113 ( .A(n_114), .B(n_284), .C(n_321), .Y(n_113) );
NOR3xp33_ASAP7_75t_L g114 ( .A(n_115), .B(n_252), .C(n_267), .Y(n_114) );
OAI221xp5_ASAP7_75t_L g115 ( .A1(n_116), .A2(n_196), .B1(n_226), .B2(n_238), .C(n_239), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
NAND2xp5_ASAP7_75t_SL g117 ( .A(n_118), .B(n_181), .Y(n_117) );
OAI22xp33_ASAP7_75t_SL g312 ( .A1(n_118), .A2(n_276), .B1(n_313), .B2(n_316), .Y(n_312) );
OR2x2_ASAP7_75t_L g118 ( .A(n_119), .B(n_153), .Y(n_118) );
OAI21xp33_ASAP7_75t_SL g322 ( .A1(n_119), .A2(n_323), .B(n_329), .Y(n_322) );
OR2x2_ASAP7_75t_L g351 ( .A(n_119), .B(n_183), .Y(n_351) );
AND2x2_ASAP7_75t_L g352 ( .A(n_119), .B(n_271), .Y(n_352) );
INVx2_ASAP7_75t_L g383 ( .A(n_119), .Y(n_383) );
INVx2_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
NAND2xp5_ASAP7_75t_L g364 ( .A(n_120), .B(n_243), .Y(n_364) );
INVx2_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
OR2x2_ASAP7_75t_L g238 ( .A(n_121), .B(n_156), .Y(n_238) );
BUFx3_ASAP7_75t_L g264 ( .A(n_121), .Y(n_264) );
AND2x2_ASAP7_75t_L g400 ( .A(n_121), .B(n_401), .Y(n_400) );
AND2x2_ASAP7_75t_L g423 ( .A(n_121), .B(n_184), .Y(n_423) );
AND2x4_ASAP7_75t_L g121 ( .A(n_122), .B(n_127), .Y(n_121) );
AND2x4_ASAP7_75t_L g195 ( .A(n_122), .B(n_127), .Y(n_195) );
AO21x2_ASAP7_75t_L g127 ( .A1(n_123), .A2(n_128), .B(n_145), .Y(n_127) );
CKINVDCx5p33_ASAP7_75t_R g172 ( .A(n_123), .Y(n_172) );
AOI21xp5_ASAP7_75t_L g186 ( .A1(n_123), .A2(n_187), .B(n_188), .Y(n_186) );
OA21x2_ASAP7_75t_L g437 ( .A1(n_123), .A2(n_438), .B(n_442), .Y(n_437) );
AOI21xp5_ASAP7_75t_L g480 ( .A1(n_123), .A2(n_481), .B(n_482), .Y(n_480) );
OA21x2_ASAP7_75t_L g581 ( .A1(n_123), .A2(n_438), .B(n_442), .Y(n_581) );
BUFx6f_ASAP7_75t_L g123 ( .A(n_124), .Y(n_123) );
AND2x2_ASAP7_75t_SL g124 ( .A(n_125), .B(n_126), .Y(n_124) );
AND2x4_ASAP7_75t_L g206 ( .A(n_125), .B(n_126), .Y(n_206) );
AND2x4_ASAP7_75t_L g129 ( .A(n_130), .B(n_135), .Y(n_129) );
AND2x2_ASAP7_75t_L g130 ( .A(n_131), .B(n_133), .Y(n_130) );
INVx2_ASAP7_75t_L g131 ( .A(n_132), .Y(n_131) );
AND2x2_ASAP7_75t_L g147 ( .A(n_132), .B(n_134), .Y(n_147) );
AND2x4_ASAP7_75t_L g165 ( .A(n_132), .B(n_142), .Y(n_165) );
HB1xp67_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
BUFx3_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
AND2x6_ASAP7_75t_L g146 ( .A(n_136), .B(n_147), .Y(n_146) );
INVx2_ASAP7_75t_L g152 ( .A(n_137), .Y(n_152) );
AND2x6_ASAP7_75t_L g163 ( .A(n_137), .B(n_140), .Y(n_163) );
AND2x4_ASAP7_75t_L g138 ( .A(n_139), .B(n_144), .Y(n_138) );
AND2x4_ASAP7_75t_L g139 ( .A(n_140), .B(n_142), .Y(n_139) );
INVx2_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
INVx2_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
INVx5_ASAP7_75t_L g166 ( .A(n_144), .Y(n_166) );
AND2x4_ASAP7_75t_L g148 ( .A(n_147), .B(n_149), .Y(n_148) );
NOR2x1p5_ASAP7_75t_L g149 ( .A(n_150), .B(n_151), .Y(n_149) );
INVx3_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
INVx1_ASAP7_75t_SL g153 ( .A(n_154), .Y(n_153) );
NAND2xp5_ASAP7_75t_L g343 ( .A(n_154), .B(n_184), .Y(n_343) );
INVx1_ASAP7_75t_L g380 ( .A(n_154), .Y(n_380) );
AND2x2_ASAP7_75t_L g154 ( .A(n_155), .B(n_170), .Y(n_154) );
AND2x2_ASAP7_75t_L g194 ( .A(n_155), .B(n_195), .Y(n_194) );
INVx1_ASAP7_75t_L g401 ( .A(n_155), .Y(n_401) );
INVx2_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
INVx2_ASAP7_75t_L g244 ( .A(n_156), .Y(n_244) );
AND2x2_ASAP7_75t_L g245 ( .A(n_156), .B(n_170), .Y(n_245) );
AND2x2_ASAP7_75t_L g266 ( .A(n_156), .B(n_185), .Y(n_266) );
AND2x2_ASAP7_75t_L g348 ( .A(n_156), .B(n_171), .Y(n_348) );
AO21x2_ASAP7_75t_L g156 ( .A1(n_157), .A2(n_159), .B(n_168), .Y(n_156) );
INVx4_ASAP7_75t_L g169 ( .A(n_157), .Y(n_169) );
INVx3_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
BUFx4f_ASAP7_75t_L g180 ( .A(n_158), .Y(n_180) );
NAND2xp5_ASAP7_75t_L g159 ( .A(n_160), .B(n_167), .Y(n_159) );
AOI21xp5_ASAP7_75t_L g161 ( .A1(n_162), .A2(n_164), .B(n_166), .Y(n_161) );
NAND2xp5_ASAP7_75t_L g223 ( .A(n_163), .B(n_224), .Y(n_223) );
AOI21xp5_ASAP7_75t_L g175 ( .A1(n_166), .A2(n_176), .B(n_177), .Y(n_175) );
AOI21xp5_ASAP7_75t_L g189 ( .A1(n_166), .A2(n_190), .B(n_191), .Y(n_189) );
AOI21xp5_ASAP7_75t_L g203 ( .A1(n_166), .A2(n_204), .B(n_205), .Y(n_203) );
AOI21xp5_ASAP7_75t_L g212 ( .A1(n_166), .A2(n_213), .B(n_214), .Y(n_212) );
AOI21xp5_ASAP7_75t_L g221 ( .A1(n_166), .A2(n_222), .B(n_223), .Y(n_221) );
AOI21xp5_ASAP7_75t_L g233 ( .A1(n_166), .A2(n_234), .B(n_235), .Y(n_233) );
AOI21xp5_ASAP7_75t_L g439 ( .A1(n_166), .A2(n_440), .B(n_441), .Y(n_439) );
AOI21xp5_ASAP7_75t_L g449 ( .A1(n_166), .A2(n_450), .B(n_451), .Y(n_449) );
AOI21xp5_ASAP7_75t_L g461 ( .A1(n_166), .A2(n_462), .B(n_463), .Y(n_461) );
AOI21xp5_ASAP7_75t_L g470 ( .A1(n_166), .A2(n_471), .B(n_472), .Y(n_470) );
AOI21xp5_ASAP7_75t_L g483 ( .A1(n_166), .A2(n_484), .B(n_485), .Y(n_483) );
AOI21xp5_ASAP7_75t_L g490 ( .A1(n_166), .A2(n_491), .B(n_492), .Y(n_490) );
AOI21xp5_ASAP7_75t_L g515 ( .A1(n_166), .A2(n_516), .B(n_517), .Y(n_515) );
AOI21xp5_ASAP7_75t_L g531 ( .A1(n_166), .A2(n_532), .B(n_533), .Y(n_531) );
INVx3_ASAP7_75t_L g209 ( .A(n_169), .Y(n_209) );
AND2x4_ASAP7_75t_SL g241 ( .A(n_170), .B(n_185), .Y(n_241) );
INVx1_ASAP7_75t_L g272 ( .A(n_170), .Y(n_272) );
INVx2_ASAP7_75t_L g280 ( .A(n_170), .Y(n_280) );
HB1xp67_ASAP7_75t_L g304 ( .A(n_170), .Y(n_304) );
INVx3_ASAP7_75t_L g170 ( .A(n_171), .Y(n_170) );
HB1xp67_ASAP7_75t_L g193 ( .A(n_171), .Y(n_193) );
AOI21x1_ASAP7_75t_L g171 ( .A1(n_172), .A2(n_173), .B(n_179), .Y(n_171) );
AO21x2_ASAP7_75t_L g487 ( .A1(n_172), .A2(n_488), .B(n_494), .Y(n_487) );
NAND2xp5_ASAP7_75t_L g173 ( .A(n_174), .B(n_178), .Y(n_173) );
AOI21xp5_ASAP7_75t_L g218 ( .A1(n_180), .A2(n_219), .B(n_220), .Y(n_218) );
NAND2xp5_ASAP7_75t_L g181 ( .A(n_182), .B(n_194), .Y(n_181) );
AND2x2_ASAP7_75t_L g419 ( .A(n_182), .B(n_282), .Y(n_419) );
INVx1_ASAP7_75t_L g182 ( .A(n_183), .Y(n_182) );
NAND2xp5_ASAP7_75t_L g183 ( .A(n_184), .B(n_193), .Y(n_183) );
NAND2x1p5_ASAP7_75t_L g278 ( .A(n_184), .B(n_279), .Y(n_278) );
AND2x2_ASAP7_75t_L g330 ( .A(n_184), .B(n_245), .Y(n_330) );
AND2x2_ASAP7_75t_L g347 ( .A(n_184), .B(n_348), .Y(n_347) );
INVx4_ASAP7_75t_L g184 ( .A(n_185), .Y(n_184) );
AND2x4_ASAP7_75t_L g271 ( .A(n_185), .B(n_272), .Y(n_271) );
INVx1_ASAP7_75t_L g287 ( .A(n_185), .Y(n_287) );
AND2x2_ASAP7_75t_L g331 ( .A(n_185), .B(n_332), .Y(n_331) );
OR2x2_ASAP7_75t_L g338 ( .A(n_185), .B(n_339), .Y(n_338) );
NOR2x1_ASAP7_75t_L g353 ( .A(n_185), .B(n_244), .Y(n_353) );
BUFx2_ASAP7_75t_L g363 ( .A(n_185), .Y(n_363) );
AND2x2_ASAP7_75t_L g388 ( .A(n_185), .B(n_348), .Y(n_388) );
AND2x2_ASAP7_75t_L g409 ( .A(n_185), .B(n_410), .Y(n_409) );
OR2x6_ASAP7_75t_L g185 ( .A(n_186), .B(n_192), .Y(n_185) );
INVx1_ASAP7_75t_L g340 ( .A(n_193), .Y(n_340) );
NAND2xp5_ASAP7_75t_SL g286 ( .A(n_194), .B(n_287), .Y(n_286) );
AND2x2_ASAP7_75t_L g370 ( .A(n_194), .B(n_241), .Y(n_370) );
INVx3_ASAP7_75t_L g277 ( .A(n_195), .Y(n_277) );
AND2x2_ASAP7_75t_L g410 ( .A(n_195), .B(n_332), .Y(n_410) );
INVx1_ASAP7_75t_SL g196 ( .A(n_197), .Y(n_196) );
AOI22xp5_ASAP7_75t_L g239 ( .A1(n_197), .A2(n_240), .B1(n_245), .B2(n_246), .Y(n_239) );
AND2x2_ASAP7_75t_L g197 ( .A(n_198), .B(n_207), .Y(n_197) );
INVx4_ASAP7_75t_L g237 ( .A(n_198), .Y(n_237) );
INVx2_ASAP7_75t_L g274 ( .A(n_198), .Y(n_274) );
NAND2x1_ASAP7_75t_L g300 ( .A(n_198), .B(n_217), .Y(n_300) );
OR2x2_ASAP7_75t_L g315 ( .A(n_198), .B(n_250), .Y(n_315) );
OR2x2_ASAP7_75t_SL g342 ( .A(n_198), .B(n_314), .Y(n_342) );
AND2x2_ASAP7_75t_L g355 ( .A(n_198), .B(n_229), .Y(n_355) );
HB1xp67_ASAP7_75t_L g376 ( .A(n_198), .Y(n_376) );
OR2x6_ASAP7_75t_L g198 ( .A(n_199), .B(n_200), .Y(n_198) );
AOI21xp5_ASAP7_75t_L g200 ( .A1(n_201), .A2(n_202), .B(n_206), .Y(n_200) );
AOI21xp5_ASAP7_75t_L g230 ( .A1(n_206), .A2(n_231), .B(n_232), .Y(n_230) );
NAND2xp5_ASAP7_75t_L g464 ( .A(n_206), .B(n_465), .Y(n_464) );
INVx1_ASAP7_75t_SL g512 ( .A(n_206), .Y(n_512) );
AOI21xp5_ASAP7_75t_L g528 ( .A1(n_206), .A2(n_529), .B(n_530), .Y(n_528) );
INVx2_ASAP7_75t_L g255 ( .A(n_207), .Y(n_255) );
AND2x2_ASAP7_75t_L g387 ( .A(n_207), .B(n_361), .Y(n_387) );
NOR2x1_ASAP7_75t_SL g207 ( .A(n_208), .B(n_217), .Y(n_207) );
AND2x2_ASAP7_75t_L g228 ( .A(n_208), .B(n_229), .Y(n_228) );
AND2x2_ASAP7_75t_L g404 ( .A(n_208), .B(n_327), .Y(n_404) );
AO21x1_ASAP7_75t_SL g208 ( .A1(n_209), .A2(n_210), .B(n_216), .Y(n_208) );
AO21x2_ASAP7_75t_L g251 ( .A1(n_209), .A2(n_210), .B(n_216), .Y(n_251) );
AO21x2_ASAP7_75t_L g446 ( .A1(n_209), .A2(n_447), .B(n_453), .Y(n_446) );
AO21x2_ASAP7_75t_L g467 ( .A1(n_209), .A2(n_468), .B(n_474), .Y(n_467) );
AO21x2_ASAP7_75t_L g501 ( .A1(n_209), .A2(n_468), .B(n_474), .Y(n_501) );
AO21x2_ASAP7_75t_L g505 ( .A1(n_209), .A2(n_447), .B(n_453), .Y(n_505) );
NAND2xp5_ASAP7_75t_L g210 ( .A(n_211), .B(n_215), .Y(n_210) );
OR2x2_ASAP7_75t_L g236 ( .A(n_217), .B(n_237), .Y(n_236) );
AND2x2_ASAP7_75t_L g247 ( .A(n_217), .B(n_237), .Y(n_247) );
AND2x2_ASAP7_75t_L g293 ( .A(n_217), .B(n_250), .Y(n_293) );
OR2x2_ASAP7_75t_L g314 ( .A(n_217), .B(n_229), .Y(n_314) );
INVx2_ASAP7_75t_SL g320 ( .A(n_217), .Y(n_320) );
AND2x2_ASAP7_75t_L g326 ( .A(n_217), .B(n_327), .Y(n_326) );
AND2x2_ASAP7_75t_L g336 ( .A(n_217), .B(n_319), .Y(n_336) );
BUFx2_ASAP7_75t_L g358 ( .A(n_217), .Y(n_358) );
OR2x6_ASAP7_75t_L g217 ( .A(n_218), .B(n_225), .Y(n_217) );
INVx2_ASAP7_75t_L g405 ( .A(n_226), .Y(n_405) );
OR2x2_ASAP7_75t_L g226 ( .A(n_227), .B(n_236), .Y(n_226) );
OR2x2_ASAP7_75t_L g430 ( .A(n_227), .B(n_274), .Y(n_430) );
INVx2_ASAP7_75t_SL g227 ( .A(n_228), .Y(n_227) );
NAND2xp5_ASAP7_75t_L g296 ( .A(n_228), .B(n_237), .Y(n_296) );
AND2x2_ASAP7_75t_L g367 ( .A(n_228), .B(n_247), .Y(n_367) );
INVx1_ASAP7_75t_L g249 ( .A(n_229), .Y(n_249) );
HB1xp67_ASAP7_75t_L g258 ( .A(n_229), .Y(n_258) );
INVx1_ASAP7_75t_L g291 ( .A(n_229), .Y(n_291) );
INVx2_ASAP7_75t_L g327 ( .A(n_229), .Y(n_327) );
NOR2xp67_ASAP7_75t_L g257 ( .A(n_237), .B(n_258), .Y(n_257) );
BUFx2_ASAP7_75t_L g317 ( .A(n_237), .Y(n_317) );
INVx2_ASAP7_75t_SL g393 ( .A(n_238), .Y(n_393) );
AOI22xp33_ASAP7_75t_L g294 ( .A1(n_240), .A2(n_295), .B1(n_297), .B2(n_301), .Y(n_294) );
AND2x2_ASAP7_75t_SL g240 ( .A(n_241), .B(n_242), .Y(n_240) );
AND2x2_ASAP7_75t_L g421 ( .A(n_241), .B(n_277), .Y(n_421) );
INVx1_ASAP7_75t_L g242 ( .A(n_243), .Y(n_242) );
NOR2xp33_ASAP7_75t_L g366 ( .A(n_243), .B(n_287), .Y(n_366) );
INVx1_ASAP7_75t_L g243 ( .A(n_244), .Y(n_243) );
AND2x2_ASAP7_75t_L g332 ( .A(n_244), .B(n_280), .Y(n_332) );
NAND2xp5_ASAP7_75t_L g381 ( .A(n_245), .B(n_382), .Y(n_381) );
INVx1_ASAP7_75t_L g275 ( .A(n_246), .Y(n_275) );
AOI221xp5_ASAP7_75t_L g389 ( .A1(n_246), .A2(n_390), .B1(n_394), .B2(n_396), .C(n_398), .Y(n_389) );
AND2x2_ASAP7_75t_L g246 ( .A(n_247), .B(n_248), .Y(n_246) );
AND2x2_ASAP7_75t_L g259 ( .A(n_247), .B(n_260), .Y(n_259) );
INVxp67_ASAP7_75t_SL g283 ( .A(n_247), .Y(n_283) );
NAND2xp5_ASAP7_75t_L g345 ( .A(n_247), .B(n_290), .Y(n_345) );
INVx1_ASAP7_75t_SL g341 ( .A(n_248), .Y(n_341) );
AOI221xp5_ASAP7_75t_SL g369 ( .A1(n_248), .A2(n_259), .B1(n_370), .B2(n_371), .C(n_374), .Y(n_369) );
AOI322xp5_ASAP7_75t_L g402 ( .A1(n_248), .A2(n_320), .A3(n_347), .B1(n_403), .B2(n_405), .C1(n_406), .C2(n_409), .Y(n_402) );
AND2x2_ASAP7_75t_L g248 ( .A(n_249), .B(n_250), .Y(n_248) );
BUFx2_ASAP7_75t_L g269 ( .A(n_249), .Y(n_269) );
HB1xp67_ASAP7_75t_L g261 ( .A(n_250), .Y(n_261) );
INVx2_ASAP7_75t_L g319 ( .A(n_250), .Y(n_319) );
AND2x2_ASAP7_75t_L g360 ( .A(n_250), .B(n_361), .Y(n_360) );
INVx3_ASAP7_75t_L g250 ( .A(n_251), .Y(n_250) );
OA21x2_ASAP7_75t_SL g252 ( .A1(n_253), .A2(n_259), .B(n_262), .Y(n_252) );
AOI211xp5_ASAP7_75t_L g422 ( .A1(n_253), .A2(n_423), .B(n_424), .C(n_428), .Y(n_422) );
INVx1_ASAP7_75t_SL g253 ( .A(n_254), .Y(n_253) );
OR2x2_ASAP7_75t_L g254 ( .A(n_255), .B(n_256), .Y(n_254) );
OR2x2_ASAP7_75t_L g311 ( .A(n_255), .B(n_273), .Y(n_311) );
OR2x2_ASAP7_75t_L g395 ( .A(n_255), .B(n_290), .Y(n_395) );
INVx1_ASAP7_75t_L g256 ( .A(n_257), .Y(n_256) );
AND2x2_ASAP7_75t_L g335 ( .A(n_257), .B(n_336), .Y(n_335) );
INVx1_ASAP7_75t_L g413 ( .A(n_260), .Y(n_413) );
INVx1_ASAP7_75t_L g260 ( .A(n_261), .Y(n_260) );
INVx1_ASAP7_75t_L g299 ( .A(n_261), .Y(n_299) );
INVx1_ASAP7_75t_SL g262 ( .A(n_263), .Y(n_262) );
OR2x2_ASAP7_75t_L g263 ( .A(n_264), .B(n_265), .Y(n_263) );
OR2x2_ASAP7_75t_L g268 ( .A(n_264), .B(n_269), .Y(n_268) );
INVx1_ASAP7_75t_L g265 ( .A(n_266), .Y(n_265) );
AND2x2_ASAP7_75t_L g303 ( .A(n_266), .B(n_304), .Y(n_303) );
OAI322xp33_ASAP7_75t_L g267 ( .A1(n_268), .A2(n_270), .A3(n_273), .B1(n_275), .B2(n_276), .C1(n_281), .C2(n_283), .Y(n_267) );
INVx1_ASAP7_75t_L g309 ( .A(n_268), .Y(n_309) );
OR2x2_ASAP7_75t_L g281 ( .A(n_270), .B(n_282), .Y(n_281) );
NAND2xp5_ASAP7_75t_L g407 ( .A(n_270), .B(n_408), .Y(n_407) );
INVx2_ASAP7_75t_L g270 ( .A(n_271), .Y(n_270) );
INVx2_ASAP7_75t_L g273 ( .A(n_274), .Y(n_273) );
AND2x2_ASAP7_75t_L g292 ( .A(n_274), .B(n_293), .Y(n_292) );
OAI32xp33_ASAP7_75t_L g337 ( .A1(n_274), .A2(n_338), .A3(n_341), .B1(n_342), .B2(n_343), .Y(n_337) );
OR2x2_ASAP7_75t_L g276 ( .A(n_277), .B(n_278), .Y(n_276) );
INVx2_ASAP7_75t_L g282 ( .A(n_277), .Y(n_282) );
NAND2xp5_ASAP7_75t_L g339 ( .A(n_277), .B(n_340), .Y(n_339) );
NOR2x1_ASAP7_75t_L g379 ( .A(n_277), .B(n_380), .Y(n_379) );
AND2x2_ASAP7_75t_L g403 ( .A(n_277), .B(n_404), .Y(n_403) );
INVx1_ASAP7_75t_L g324 ( .A(n_278), .Y(n_324) );
INVx1_ASAP7_75t_SL g279 ( .A(n_280), .Y(n_279) );
NAND2xp5_ASAP7_75t_L g416 ( .A(n_282), .B(n_348), .Y(n_416) );
NOR2xp33_ASAP7_75t_L g284 ( .A(n_285), .B(n_305), .Y(n_284) );
OAI21xp33_ASAP7_75t_L g285 ( .A1(n_286), .A2(n_288), .B(n_294), .Y(n_285) );
INVx1_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
AND2x4_ASAP7_75t_SL g289 ( .A(n_290), .B(n_292), .Y(n_289) );
INVx3_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
AND2x2_ASAP7_75t_L g354 ( .A(n_293), .B(n_355), .Y(n_354) );
INVx1_ASAP7_75t_SL g295 ( .A(n_296), .Y(n_295) );
OAI22xp5_ASAP7_75t_L g417 ( .A1(n_296), .A2(n_316), .B1(n_418), .B2(n_420), .Y(n_417) );
INVx1_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
A2O1A1Ixp33_ASAP7_75t_L g344 ( .A1(n_298), .A2(n_345), .B(n_346), .C(n_349), .Y(n_344) );
OR2x2_ASAP7_75t_L g298 ( .A(n_299), .B(n_300), .Y(n_298) );
INVx3_ASAP7_75t_L g426 ( .A(n_300), .Y(n_426) );
INVx2_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
INVx1_ASAP7_75t_L g302 ( .A(n_303), .Y(n_302) );
INVx2_ASAP7_75t_L g307 ( .A(n_304), .Y(n_307) );
AO21x1_ASAP7_75t_L g305 ( .A1(n_306), .A2(n_308), .B(n_312), .Y(n_305) );
HB1xp67_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
INVx2_ASAP7_75t_L g372 ( .A(n_307), .Y(n_372) );
AND2x2_ASAP7_75t_L g308 ( .A(n_309), .B(n_310), .Y(n_308) );
INVx1_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
NOR2xp33_ASAP7_75t_L g398 ( .A(n_313), .B(n_399), .Y(n_398) );
OR2x2_ASAP7_75t_L g313 ( .A(n_314), .B(n_315), .Y(n_313) );
INVx1_ASAP7_75t_L g328 ( .A(n_315), .Y(n_328) );
OR2x2_ASAP7_75t_L g316 ( .A(n_317), .B(n_318), .Y(n_316) );
INVx1_ASAP7_75t_L g385 ( .A(n_318), .Y(n_385) );
NAND2xp5_ASAP7_75t_L g318 ( .A(n_319), .B(n_320), .Y(n_318) );
NOR3xp33_ASAP7_75t_L g321 ( .A(n_322), .B(n_344), .C(n_356), .Y(n_321) );
NAND2xp5_ASAP7_75t_L g323 ( .A(n_324), .B(n_325), .Y(n_323) );
OAI21xp5_ASAP7_75t_SL g386 ( .A1(n_325), .A2(n_387), .B(n_388), .Y(n_386) );
AND2x4_ASAP7_75t_L g325 ( .A(n_326), .B(n_328), .Y(n_325) );
INVx1_ASAP7_75t_L g361 ( .A(n_327), .Y(n_361) );
O2A1O1Ixp5_ASAP7_75t_SL g329 ( .A1(n_330), .A2(n_331), .B(n_333), .C(n_337), .Y(n_329) );
INVx1_ASAP7_75t_L g333 ( .A(n_334), .Y(n_333) );
INVx2_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
HB1xp67_ASAP7_75t_L g429 ( .A(n_339), .Y(n_429) );
INVx2_ASAP7_75t_L g414 ( .A(n_342), .Y(n_414) );
AOI21xp33_ASAP7_75t_L g428 ( .A1(n_343), .A2(n_429), .B(n_430), .Y(n_428) );
INVx1_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
INVx1_ASAP7_75t_L g408 ( .A(n_348), .Y(n_408) );
OAI31xp33_ASAP7_75t_L g349 ( .A1(n_350), .A2(n_352), .A3(n_353), .B(n_354), .Y(n_349) );
INVx1_ASAP7_75t_SL g350 ( .A(n_351), .Y(n_350) );
INVx1_ASAP7_75t_L g427 ( .A(n_355), .Y(n_427) );
OAI21xp5_ASAP7_75t_L g356 ( .A1(n_357), .A2(n_362), .B(n_365), .Y(n_356) );
NAND2xp5_ASAP7_75t_L g357 ( .A(n_358), .B(n_359), .Y(n_357) );
BUFx2_ASAP7_75t_SL g359 ( .A(n_360), .Y(n_359) );
INVx1_ASAP7_75t_L g377 ( .A(n_360), .Y(n_377) );
AOI21xp33_ASAP7_75t_SL g424 ( .A1(n_362), .A2(n_425), .B(n_427), .Y(n_424) );
OR2x2_ASAP7_75t_L g362 ( .A(n_363), .B(n_364), .Y(n_362) );
INVx2_ASAP7_75t_L g392 ( .A(n_363), .Y(n_392) );
NAND2xp5_ASAP7_75t_L g397 ( .A(n_363), .B(n_383), .Y(n_397) );
NAND2xp5_ASAP7_75t_L g399 ( .A(n_363), .B(n_400), .Y(n_399) );
INVx2_ASAP7_75t_L g373 ( .A(n_364), .Y(n_373) );
NAND2xp5_ASAP7_75t_L g365 ( .A(n_366), .B(n_367), .Y(n_365) );
NAND5xp2_ASAP7_75t_L g368 ( .A(n_369), .B(n_389), .C(n_402), .D(n_411), .E(n_422), .Y(n_368) );
AND2x2_ASAP7_75t_L g371 ( .A(n_372), .B(n_373), .Y(n_371) );
OAI221xp5_ASAP7_75t_L g374 ( .A1(n_375), .A2(n_378), .B1(n_381), .B2(n_384), .C(n_386), .Y(n_374) );
OR2x2_ASAP7_75t_L g375 ( .A(n_376), .B(n_377), .Y(n_375) );
INVx1_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
INVxp67_ASAP7_75t_SL g382 ( .A(n_383), .Y(n_382) );
INVx1_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
INVxp67_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
NAND2xp5_ASAP7_75t_L g391 ( .A(n_392), .B(n_393), .Y(n_391) );
INVx1_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
INVx1_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
INVx1_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
AOI21xp5_ASAP7_75t_L g411 ( .A1(n_412), .A2(n_415), .B(n_417), .Y(n_411) );
AND2x4_ASAP7_75t_L g412 ( .A(n_413), .B(n_414), .Y(n_412) );
INVx1_ASAP7_75t_SL g415 ( .A(n_416), .Y(n_415) );
INVx1_ASAP7_75t_SL g418 ( .A(n_419), .Y(n_418) );
INVxp67_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
INVx1_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
INVx3_ASAP7_75t_L g721 ( .A(n_431), .Y(n_721) );
NAND4xp75_ASAP7_75t_L g431 ( .A(n_432), .B(n_621), .C(n_661), .D(n_690), .Y(n_431) );
NOR2x1_ASAP7_75t_L g432 ( .A(n_433), .B(n_583), .Y(n_432) );
NAND2xp5_ASAP7_75t_L g433 ( .A(n_434), .B(n_540), .Y(n_433) );
AOI21xp5_ASAP7_75t_L g434 ( .A1(n_435), .A2(n_475), .B(n_495), .Y(n_434) );
AND2x2_ASAP7_75t_SL g435 ( .A(n_436), .B(n_443), .Y(n_435) );
AND2x4_ASAP7_75t_L g539 ( .A(n_436), .B(n_500), .Y(n_539) );
INVx1_ASAP7_75t_SL g592 ( .A(n_436), .Y(n_592) );
AOI21xp33_ASAP7_75t_L g627 ( .A1(n_436), .A2(n_628), .B(n_631), .Y(n_627) );
A2O1A1Ixp33_ASAP7_75t_SL g631 ( .A1(n_436), .A2(n_632), .B(n_633), .C(n_634), .Y(n_631) );
NAND2x1_ASAP7_75t_L g672 ( .A(n_436), .B(n_673), .Y(n_672) );
NAND2xp5_ASAP7_75t_L g694 ( .A(n_436), .B(n_633), .Y(n_694) );
INVx2_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
INVx2_ASAP7_75t_L g498 ( .A(n_437), .Y(n_498) );
HB1xp67_ASAP7_75t_L g571 ( .A(n_437), .Y(n_571) );
AND2x2_ASAP7_75t_L g443 ( .A(n_444), .B(n_454), .Y(n_443) );
AND2x2_ASAP7_75t_L g563 ( .A(n_444), .B(n_564), .Y(n_563) );
AND2x2_ASAP7_75t_L g644 ( .A(n_444), .B(n_500), .Y(n_644) );
INVx1_ASAP7_75t_L g704 ( .A(n_444), .Y(n_704) );
BUFx2_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
AND2x2_ASAP7_75t_L g548 ( .A(n_445), .B(n_466), .Y(n_548) );
AND2x2_ASAP7_75t_L g673 ( .A(n_445), .B(n_467), .Y(n_673) );
AND2x2_ASAP7_75t_L g678 ( .A(n_445), .B(n_638), .Y(n_678) );
INVx2_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
INVxp67_ASAP7_75t_L g554 ( .A(n_446), .Y(n_554) );
BUFx3_ASAP7_75t_L g587 ( .A(n_446), .Y(n_587) );
AND2x2_ASAP7_75t_L g633 ( .A(n_446), .B(n_467), .Y(n_633) );
NAND2xp5_ASAP7_75t_L g447 ( .A(n_448), .B(n_452), .Y(n_447) );
AND2x2_ASAP7_75t_L g618 ( .A(n_454), .B(n_497), .Y(n_618) );
AND2x2_ASAP7_75t_L g454 ( .A(n_455), .B(n_466), .Y(n_454) );
AND2x4_ASAP7_75t_L g500 ( .A(n_455), .B(n_501), .Y(n_500) );
OR2x2_ASAP7_75t_L g610 ( .A(n_455), .B(n_594), .Y(n_610) );
AND2x2_ASAP7_75t_SL g653 ( .A(n_455), .B(n_581), .Y(n_653) );
INVx2_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
BUFx2_ASAP7_75t_L g589 ( .A(n_456), .Y(n_589) );
INVx2_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
INVx2_ASAP7_75t_L g550 ( .A(n_457), .Y(n_550) );
OAI21x1_ASAP7_75t_SL g457 ( .A1(n_458), .A2(n_460), .B(n_464), .Y(n_457) );
INVx1_ASAP7_75t_L g465 ( .A(n_459), .Y(n_465) );
NAND2xp5_ASAP7_75t_L g553 ( .A(n_466), .B(n_550), .Y(n_553) );
AND2x2_ASAP7_75t_L g638 ( .A(n_466), .B(n_581), .Y(n_638) );
INVx2_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
AND2x2_ASAP7_75t_L g635 ( .A(n_467), .B(n_498), .Y(n_635) );
AND2x2_ASAP7_75t_L g655 ( .A(n_467), .B(n_581), .Y(n_655) );
NAND2xp5_ASAP7_75t_SL g468 ( .A(n_469), .B(n_473), .Y(n_468) );
NAND2xp5_ASAP7_75t_L g573 ( .A(n_475), .B(n_544), .Y(n_573) );
AOI221xp5_ASAP7_75t_L g666 ( .A1(n_475), .A2(n_667), .B1(n_668), .B2(n_669), .C(n_671), .Y(n_666) );
INVx2_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
OAI332xp33_ASAP7_75t_L g700 ( .A1(n_476), .A2(n_560), .A3(n_567), .B1(n_626), .B2(n_701), .B3(n_702), .C1(n_703), .C2(n_705), .Y(n_700) );
NAND2x1p5_ASAP7_75t_L g476 ( .A(n_477), .B(n_486), .Y(n_476) );
AND2x2_ASAP7_75t_L g506 ( .A(n_477), .B(n_487), .Y(n_506) );
AND2x2_ASAP7_75t_L g523 ( .A(n_477), .B(n_524), .Y(n_523) );
INVx4_ASAP7_75t_L g535 ( .A(n_477), .Y(n_535) );
AND2x2_ASAP7_75t_SL g595 ( .A(n_477), .B(n_536), .Y(n_595) );
INVx5_ASAP7_75t_L g477 ( .A(n_478), .Y(n_477) );
NOR2x1_ASAP7_75t_SL g557 ( .A(n_478), .B(n_524), .Y(n_557) );
NAND2xp5_ASAP7_75t_L g561 ( .A(n_478), .B(n_486), .Y(n_561) );
AND2x2_ASAP7_75t_L g568 ( .A(n_478), .B(n_487), .Y(n_568) );
BUFx2_ASAP7_75t_L g603 ( .A(n_478), .Y(n_603) );
AND2x2_ASAP7_75t_L g658 ( .A(n_478), .B(n_527), .Y(n_658) );
OR2x6_ASAP7_75t_L g478 ( .A(n_479), .B(n_480), .Y(n_478) );
OR2x2_ASAP7_75t_L g526 ( .A(n_486), .B(n_527), .Y(n_526) );
AND2x4_ASAP7_75t_L g536 ( .A(n_486), .B(n_537), .Y(n_536) );
INVx2_ASAP7_75t_L g576 ( .A(n_486), .Y(n_576) );
AND2x2_ASAP7_75t_L g646 ( .A(n_486), .B(n_545), .Y(n_646) );
AND2x2_ASAP7_75t_L g659 ( .A(n_486), .B(n_660), .Y(n_659) );
NAND2xp5_ASAP7_75t_L g677 ( .A(n_486), .B(n_660), .Y(n_677) );
INVx4_ASAP7_75t_L g486 ( .A(n_487), .Y(n_486) );
HB1xp67_ASAP7_75t_L g543 ( .A(n_487), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g488 ( .A(n_489), .B(n_493), .Y(n_488) );
OAI32xp33_ASAP7_75t_L g495 ( .A1(n_496), .A2(n_502), .A3(n_507), .B1(n_521), .B2(n_538), .Y(n_495) );
INVx2_ASAP7_75t_L g604 ( .A(n_496), .Y(n_604) );
OR2x2_ASAP7_75t_L g496 ( .A(n_497), .B(n_499), .Y(n_496) );
INVx1_ASAP7_75t_L g615 ( .A(n_497), .Y(n_615) );
BUFx2_ASAP7_75t_L g497 ( .A(n_498), .Y(n_497) );
AND2x4_ASAP7_75t_L g549 ( .A(n_498), .B(n_550), .Y(n_549) );
AND2x2_ASAP7_75t_L g682 ( .A(n_498), .B(n_587), .Y(n_682) );
INVx2_ASAP7_75t_L g499 ( .A(n_500), .Y(n_499) );
INVx2_ASAP7_75t_L g594 ( .A(n_501), .Y(n_594) );
INVx1_ASAP7_75t_L g502 ( .A(n_503), .Y(n_502) );
AND2x2_ASAP7_75t_L g503 ( .A(n_504), .B(n_506), .Y(n_503) );
INVx2_ASAP7_75t_L g582 ( .A(n_504), .Y(n_582) );
NAND2xp5_ASAP7_75t_L g624 ( .A(n_504), .B(n_625), .Y(n_624) );
BUFx2_ASAP7_75t_L g504 ( .A(n_505), .Y(n_504) );
AND2x4_ASAP7_75t_SL g593 ( .A(n_505), .B(n_594), .Y(n_593) );
INVx1_ASAP7_75t_L g670 ( .A(n_505), .Y(n_670) );
AND2x2_ASAP7_75t_L g688 ( .A(n_505), .B(n_550), .Y(n_688) );
INVx1_ASAP7_75t_L g507 ( .A(n_508), .Y(n_507) );
NOR2xp67_ASAP7_75t_SL g632 ( .A(n_508), .B(n_561), .Y(n_632) );
INVx2_ASAP7_75t_L g508 ( .A(n_509), .Y(n_508) );
NAND2xp5_ASAP7_75t_L g630 ( .A(n_509), .B(n_543), .Y(n_630) );
INVx2_ASAP7_75t_L g509 ( .A(n_510), .Y(n_509) );
AND2x2_ASAP7_75t_L g706 ( .A(n_510), .B(n_576), .Y(n_706) );
INVx1_ASAP7_75t_L g510 ( .A(n_511), .Y(n_510) );
INVx1_ASAP7_75t_L g537 ( .A(n_511), .Y(n_537) );
INVx2_ASAP7_75t_L g578 ( .A(n_511), .Y(n_578) );
AO21x2_ASAP7_75t_L g511 ( .A1(n_512), .A2(n_513), .B(n_519), .Y(n_511) );
NOR2xp33_ASAP7_75t_L g519 ( .A(n_512), .B(n_520), .Y(n_519) );
AO21x2_ASAP7_75t_L g524 ( .A1(n_512), .A2(n_513), .B(n_519), .Y(n_524) );
NAND2xp5_ASAP7_75t_L g513 ( .A(n_514), .B(n_518), .Y(n_513) );
NOR2xp33_ASAP7_75t_L g521 ( .A(n_522), .B(n_534), .Y(n_521) );
NAND2xp5_ASAP7_75t_L g665 ( .A(n_522), .B(n_580), .Y(n_665) );
AND2x4_ASAP7_75t_L g522 ( .A(n_523), .B(n_525), .Y(n_522) );
AND3x2_ASAP7_75t_L g620 ( .A(n_523), .B(n_567), .C(n_576), .Y(n_620) );
AND2x2_ASAP7_75t_L g544 ( .A(n_524), .B(n_545), .Y(n_544) );
NAND2xp5_ASAP7_75t_L g601 ( .A(n_524), .B(n_527), .Y(n_601) );
INVx2_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
OR2x2_ASAP7_75t_L g555 ( .A(n_526), .B(n_556), .Y(n_555) );
INVx2_ASAP7_75t_L g545 ( .A(n_527), .Y(n_545) );
INVx1_ASAP7_75t_L g560 ( .A(n_527), .Y(n_560) );
BUFx3_ASAP7_75t_L g567 ( .A(n_527), .Y(n_567) );
AND2x2_ASAP7_75t_L g577 ( .A(n_527), .B(n_578), .Y(n_577) );
AND2x2_ASAP7_75t_L g534 ( .A(n_535), .B(n_536), .Y(n_534) );
AND2x4_ASAP7_75t_L g586 ( .A(n_535), .B(n_587), .Y(n_586) );
NAND2xp5_ASAP7_75t_L g629 ( .A(n_535), .B(n_545), .Y(n_629) );
AND2x2_ASAP7_75t_L g585 ( .A(n_536), .B(n_560), .Y(n_585) );
INVx2_ASAP7_75t_L g612 ( .A(n_536), .Y(n_612) );
INVx1_ASAP7_75t_SL g538 ( .A(n_539), .Y(n_538) );
AOI211xp5_ASAP7_75t_L g540 ( .A1(n_541), .A2(n_546), .B(n_551), .C(n_572), .Y(n_540) );
OAI21xp5_ASAP7_75t_L g692 ( .A1(n_541), .A2(n_668), .B(n_693), .Y(n_692) );
INVx1_ASAP7_75t_L g541 ( .A(n_542), .Y(n_541) );
NAND2xp5_ASAP7_75t_L g542 ( .A(n_543), .B(n_544), .Y(n_542) );
NAND2xp5_ASAP7_75t_L g602 ( .A(n_544), .B(n_603), .Y(n_602) );
AOI211xp5_ASAP7_75t_SL g622 ( .A1(n_544), .A2(n_623), .B(n_627), .C(n_636), .Y(n_622) );
AND2x2_ASAP7_75t_L g608 ( .A(n_545), .B(n_568), .Y(n_608) );
OR2x2_ASAP7_75t_L g611 ( .A(n_545), .B(n_612), .Y(n_611) );
INVx1_ASAP7_75t_SL g546 ( .A(n_547), .Y(n_546) );
NAND2xp5_ASAP7_75t_L g547 ( .A(n_548), .B(n_549), .Y(n_547) );
NAND2xp5_ASAP7_75t_SL g698 ( .A(n_548), .B(n_653), .Y(n_698) );
NAND2xp5_ASAP7_75t_SL g607 ( .A(n_549), .B(n_594), .Y(n_607) );
AOI221xp5_ASAP7_75t_L g663 ( .A1(n_549), .A2(n_575), .B1(n_655), .B2(n_658), .C(n_664), .Y(n_663) );
AND2x4_ASAP7_75t_L g580 ( .A(n_550), .B(n_581), .Y(n_580) );
OR2x2_ASAP7_75t_L g626 ( .A(n_550), .B(n_581), .Y(n_626) );
OAI221xp5_ASAP7_75t_SL g551 ( .A1(n_552), .A2(n_555), .B1(n_558), .B2(n_562), .C(n_565), .Y(n_551) );
AND2x2_ASAP7_75t_L g697 ( .A(n_552), .B(n_698), .Y(n_697) );
OR2x2_ASAP7_75t_L g552 ( .A(n_553), .B(n_554), .Y(n_552) );
INVx1_ASAP7_75t_L g564 ( .A(n_553), .Y(n_564) );
INVx1_ASAP7_75t_L g650 ( .A(n_554), .Y(n_650) );
NOR2xp33_ASAP7_75t_L g671 ( .A(n_555), .B(n_672), .Y(n_671) );
INVx1_ASAP7_75t_L g556 ( .A(n_557), .Y(n_556) );
AND2x2_ASAP7_75t_L g569 ( .A(n_557), .B(n_560), .Y(n_569) );
AND2x2_ASAP7_75t_L g645 ( .A(n_557), .B(n_646), .Y(n_645) );
OR2x2_ASAP7_75t_L g558 ( .A(n_559), .B(n_561), .Y(n_558) );
INVx1_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
INVx1_ASAP7_75t_SL g562 ( .A(n_563), .Y(n_562) );
AND2x2_ASAP7_75t_L g570 ( .A(n_564), .B(n_571), .Y(n_570) );
OAI21xp5_ASAP7_75t_SL g565 ( .A1(n_566), .A2(n_569), .B(n_570), .Y(n_565) );
INVx1_ASAP7_75t_L g689 ( .A(n_566), .Y(n_689) );
AND2x2_ASAP7_75t_L g566 ( .A(n_567), .B(n_568), .Y(n_566) );
AND2x2_ASAP7_75t_L g668 ( .A(n_567), .B(n_595), .Y(n_668) );
AND2x2_ASAP7_75t_SL g641 ( .A(n_568), .B(n_577), .Y(n_641) );
AOI21xp33_ASAP7_75t_L g572 ( .A1(n_573), .A2(n_574), .B(n_579), .Y(n_572) );
OAI22xp33_ASAP7_75t_L g609 ( .A1(n_573), .A2(n_607), .B1(n_610), .B2(n_611), .Y(n_609) );
INVx1_ASAP7_75t_L g679 ( .A(n_573), .Y(n_679) );
INVx1_ASAP7_75t_L g574 ( .A(n_575), .Y(n_574) );
AND2x2_ASAP7_75t_L g575 ( .A(n_576), .B(n_577), .Y(n_575) );
INVx1_ASAP7_75t_L g599 ( .A(n_576), .Y(n_599) );
INVx1_ASAP7_75t_L g660 ( .A(n_578), .Y(n_660) );
NAND2xp5_ASAP7_75t_SL g579 ( .A(n_580), .B(n_582), .Y(n_579) );
NAND2xp5_ASAP7_75t_SL g701 ( .A(n_580), .B(n_650), .Y(n_701) );
AND2x2_ASAP7_75t_L g669 ( .A(n_581), .B(n_670), .Y(n_669) );
OAI211xp5_ASAP7_75t_L g662 ( .A1(n_582), .A2(n_663), .B(n_666), .C(n_674), .Y(n_662) );
NAND2xp5_ASAP7_75t_L g583 ( .A(n_584), .B(n_605), .Y(n_583) );
AOI322xp5_ASAP7_75t_L g584 ( .A1(n_585), .A2(n_586), .A3(n_588), .B1(n_590), .B2(n_595), .C1(n_596), .C2(n_604), .Y(n_584) );
CKINVDCx16_ASAP7_75t_R g702 ( .A(n_586), .Y(n_702) );
AND2x2_ASAP7_75t_L g652 ( .A(n_587), .B(n_653), .Y(n_652) );
INVx1_ASAP7_75t_SL g686 ( .A(n_587), .Y(n_686) );
INVx1_ASAP7_75t_L g588 ( .A(n_589), .Y(n_588) );
NOR2xp33_ASAP7_75t_SL g637 ( .A(n_589), .B(n_638), .Y(n_637) );
AND2x2_ASAP7_75t_SL g643 ( .A(n_589), .B(n_635), .Y(n_643) );
AND2x2_ASAP7_75t_L g667 ( .A(n_589), .B(n_633), .Y(n_667) );
INVx1_ASAP7_75t_L g590 ( .A(n_591), .Y(n_590) );
NAND2xp5_ASAP7_75t_L g591 ( .A(n_592), .B(n_593), .Y(n_591) );
INVx1_ASAP7_75t_L g639 ( .A(n_593), .Y(n_639) );
NAND2xp33_ASAP7_75t_SL g596 ( .A(n_597), .B(n_602), .Y(n_596) );
INVx1_ASAP7_75t_L g597 ( .A(n_598), .Y(n_597) );
AOI221xp5_ASAP7_75t_SL g642 ( .A1(n_598), .A2(n_643), .B1(n_644), .B2(n_645), .C(n_647), .Y(n_642) );
AND2x2_ASAP7_75t_L g598 ( .A(n_599), .B(n_600), .Y(n_598) );
INVxp67_ASAP7_75t_SL g600 ( .A(n_601), .Y(n_600) );
INVx1_ASAP7_75t_L g709 ( .A(n_601), .Y(n_709) );
AOI211xp5_ASAP7_75t_L g605 ( .A1(n_606), .A2(n_608), .B(n_609), .C(n_613), .Y(n_605) );
INVx1_ASAP7_75t_L g606 ( .A(n_607), .Y(n_606) );
INVx1_ASAP7_75t_SL g684 ( .A(n_608), .Y(n_684) );
INVx1_ASAP7_75t_L g616 ( .A(n_610), .Y(n_616) );
OR2x2_ASAP7_75t_L g703 ( .A(n_610), .B(n_704), .Y(n_703) );
INVx2_ASAP7_75t_SL g699 ( .A(n_611), .Y(n_699) );
AOI21xp33_ASAP7_75t_L g613 ( .A1(n_614), .A2(n_617), .B(n_619), .Y(n_613) );
NAND2xp5_ASAP7_75t_L g614 ( .A(n_615), .B(n_616), .Y(n_614) );
NAND2xp5_ASAP7_75t_L g710 ( .A(n_615), .B(n_633), .Y(n_710) );
INVx1_ASAP7_75t_SL g617 ( .A(n_618), .Y(n_617) );
INVx2_ASAP7_75t_L g619 ( .A(n_620), .Y(n_619) );
AND2x2_ASAP7_75t_L g621 ( .A(n_622), .B(n_642), .Y(n_621) );
INVx1_ASAP7_75t_SL g623 ( .A(n_624), .Y(n_623) );
NAND2xp5_ASAP7_75t_L g648 ( .A(n_625), .B(n_649), .Y(n_648) );
INVx1_ASAP7_75t_SL g625 ( .A(n_626), .Y(n_625) );
OR2x2_ASAP7_75t_L g628 ( .A(n_629), .B(n_630), .Y(n_628) );
OR2x2_ASAP7_75t_L g676 ( .A(n_629), .B(n_677), .Y(n_676) );
INVx1_ASAP7_75t_L g634 ( .A(n_635), .Y(n_634) );
AOI21xp33_ASAP7_75t_SL g636 ( .A1(n_637), .A2(n_639), .B(n_640), .Y(n_636) );
INVx2_ASAP7_75t_SL g640 ( .A(n_641), .Y(n_640) );
AOI31xp33_ASAP7_75t_L g647 ( .A1(n_648), .A2(n_651), .A3(n_654), .B(n_656), .Y(n_647) );
INVx1_ASAP7_75t_L g649 ( .A(n_650), .Y(n_649) );
INVx1_ASAP7_75t_L g651 ( .A(n_652), .Y(n_651) );
NAND2xp5_ASAP7_75t_L g685 ( .A(n_653), .B(n_686), .Y(n_685) );
INVx1_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
INVx1_ASAP7_75t_SL g656 ( .A(n_657), .Y(n_656) );
AND2x4_ASAP7_75t_L g657 ( .A(n_658), .B(n_659), .Y(n_657) );
INVx1_ASAP7_75t_L g661 ( .A(n_662), .Y(n_661) );
INVx1_ASAP7_75t_L g664 ( .A(n_665), .Y(n_664) );
AOI221xp5_ASAP7_75t_L g674 ( .A1(n_675), .A2(n_678), .B1(n_679), .B2(n_680), .C(n_683), .Y(n_674) );
INVx1_ASAP7_75t_L g675 ( .A(n_676), .Y(n_675) );
INVxp67_ASAP7_75t_L g680 ( .A(n_681), .Y(n_680) );
INVx1_ASAP7_75t_L g681 ( .A(n_682), .Y(n_681) );
OAI22xp5_ASAP7_75t_L g683 ( .A1(n_684), .A2(n_685), .B1(n_687), .B2(n_689), .Y(n_683) );
CKINVDCx16_ASAP7_75t_R g687 ( .A(n_688), .Y(n_687) );
NOR3xp33_ASAP7_75t_L g690 ( .A(n_691), .B(n_700), .C(n_707), .Y(n_690) );
NAND2xp5_ASAP7_75t_SL g691 ( .A(n_692), .B(n_695), .Y(n_691) );
INVx1_ASAP7_75t_L g693 ( .A(n_694), .Y(n_693) );
NAND2xp5_ASAP7_75t_L g695 ( .A(n_696), .B(n_699), .Y(n_695) );
INVxp67_ASAP7_75t_L g696 ( .A(n_697), .Y(n_696) );
INVx1_ASAP7_75t_SL g705 ( .A(n_706), .Y(n_705) );
NOR2xp33_ASAP7_75t_L g707 ( .A(n_708), .B(n_710), .Y(n_707) );
INVx1_ASAP7_75t_L g708 ( .A(n_709), .Y(n_708) );
BUFx4f_ASAP7_75t_SL g711 ( .A(n_712), .Y(n_711) );
CKINVDCx20_ASAP7_75t_R g712 ( .A(n_713), .Y(n_712) );
INVx1_ASAP7_75t_SL g720 ( .A(n_713), .Y(n_720) );
CKINVDCx11_ASAP7_75t_R g713 ( .A(n_714), .Y(n_713) );
OAI22xp5_ASAP7_75t_L g717 ( .A1(n_718), .A2(n_719), .B1(n_720), .B2(n_721), .Y(n_717) );
INVx3_ASAP7_75t_L g722 ( .A(n_723), .Y(n_722) );
INVx1_ASAP7_75t_SL g724 ( .A(n_725), .Y(n_724) );
INVx1_ASAP7_75t_L g725 ( .A(n_726), .Y(n_725) );
AND2x2_ASAP7_75t_L g726 ( .A(n_727), .B(n_733), .Y(n_726) );
INVxp67_ASAP7_75t_L g727 ( .A(n_728), .Y(n_727) );
NAND2xp5_ASAP7_75t_SL g728 ( .A(n_729), .B(n_732), .Y(n_728) );
INVx2_ASAP7_75t_L g729 ( .A(n_730), .Y(n_729) );
OR2x2_ASAP7_75t_SL g744 ( .A(n_730), .B(n_732), .Y(n_744) );
AOI21xp5_ASAP7_75t_L g746 ( .A1(n_730), .A2(n_747), .B(n_750), .Y(n_746) );
BUFx2_ASAP7_75t_L g733 ( .A(n_734), .Y(n_733) );
BUFx3_ASAP7_75t_L g740 ( .A(n_734), .Y(n_740) );
BUFx2_ASAP7_75t_L g751 ( .A(n_734), .Y(n_751) );
INVxp67_ASAP7_75t_L g735 ( .A(n_736), .Y(n_735) );
AOI21xp5_ASAP7_75t_L g736 ( .A1(n_737), .A2(n_739), .B(n_741), .Y(n_736) );
NOR2xp33_ASAP7_75t_SL g741 ( .A(n_739), .B(n_742), .Y(n_741) );
HB1xp67_ASAP7_75t_L g739 ( .A(n_740), .Y(n_739) );
CKINVDCx9p33_ASAP7_75t_R g743 ( .A(n_744), .Y(n_743) );
INVx1_ASAP7_75t_SL g745 ( .A(n_746), .Y(n_745) );
CKINVDCx11_ASAP7_75t_R g747 ( .A(n_748), .Y(n_747) );
CKINVDCx8_ASAP7_75t_R g748 ( .A(n_749), .Y(n_748) );
INVx2_ASAP7_75t_L g750 ( .A(n_751), .Y(n_750) );
endmodule