module real_aes_14757_n_78 (n_17, n_28, n_76, n_56, n_34, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_43, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_44, n_7, n_4, n_6, n_12, n_68, n_69, n_46, n_59, n_25, n_73, n_77, n_48, n_37, n_70, n_50, n_26, n_13, n_24, n_2, n_55, n_62, n_67, n_33, n_14, n_11, n_16, n_39, n_5, n_45, n_60, n_38, n_0, n_63, n_1, n_53, n_36, n_78);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_43;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_44;
input n_7;
input n_4;
input n_6;
input n_12;
input n_68;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_48;
input n_37;
input n_70;
input n_50;
input n_26;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_67;
input n_33;
input n_14;
input n_11;
input n_16;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_0;
input n_63;
input n_1;
input n_53;
input n_36;
output n_78;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_90;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_83;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_364;
wire n_421;
wire n_319;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_551;
wire n_320;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_97;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_92;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_94;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_98;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_82;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_656;
wire n_532;
wire n_178;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_310;
wire n_119;
wire n_455;
wire n_504;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_80;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_339;
wire n_398;
wire n_89;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_93;
wire n_182;
wire n_449;
wire n_363;
wire n_417;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_561;
wire n_142;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_527;
wire n_502;
wire n_434;
wire n_505;
wire n_600;
wire n_250;
wire n_85;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_87;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_96;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_95;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_81;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_720;
wire n_265;
wire n_354;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_419;
wire n_217;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_88;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_633;
wire n_679;
wire n_520;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_456;
wire n_359;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_103;
wire n_541;
wire n_166;
wire n_224;
wire n_546;
wire n_151;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_99;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_79;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_86;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_84;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
wire n_91;
CKINVDCx5p33_ASAP7_75t_R g673 ( .A(n_0), .Y(n_673) );
OA21x2_ASAP7_75t_L g99 ( .A1(n_1), .A2(n_47), .B(n_100), .Y(n_99) );
INVx1_ASAP7_75t_L g151 ( .A(n_1), .Y(n_151) );
NAND2xp5_ASAP7_75t_SL g238 ( .A(n_2), .B(n_103), .Y(n_238) );
INVx1_ASAP7_75t_L g674 ( .A(n_2), .Y(n_674) );
NAND2xp5_ASAP7_75t_SL g137 ( .A(n_3), .B(n_138), .Y(n_137) );
AOI221xp5_ASAP7_75t_L g517 ( .A1(n_4), .A2(n_61), .B1(n_518), .B2(n_522), .C(n_527), .Y(n_517) );
AOI22xp33_ASAP7_75t_L g602 ( .A1(n_4), .A2(n_46), .B1(n_577), .B2(n_603), .Y(n_602) );
INVx1_ASAP7_75t_L g535 ( .A(n_5), .Y(n_535) );
OAI221xp5_ASAP7_75t_L g631 ( .A1(n_5), .A2(n_9), .B1(n_632), .B2(n_633), .C(n_638), .Y(n_631) );
AOI221xp5_ASAP7_75t_L g536 ( .A1(n_6), .A2(n_62), .B1(n_518), .B2(n_537), .C(n_538), .Y(n_536) );
INVxp67_ASAP7_75t_SL g655 ( .A(n_6), .Y(n_655) );
HB1xp67_ASAP7_75t_L g683 ( .A(n_7), .Y(n_683) );
NAND2xp5_ASAP7_75t_L g140 ( .A(n_8), .B(n_116), .Y(n_140) );
INVx1_ASAP7_75t_L g534 ( .A(n_9), .Y(n_534) );
BUFx3_ASAP7_75t_L g575 ( .A(n_10), .Y(n_575) );
NAND2xp5_ASAP7_75t_L g115 ( .A(n_11), .B(n_116), .Y(n_115) );
INVx3_ASAP7_75t_L g566 ( .A(n_12), .Y(n_566) );
INVx2_ASAP7_75t_L g584 ( .A(n_13), .Y(n_584) );
INVx1_ASAP7_75t_L g621 ( .A(n_13), .Y(n_621) );
NAND2xp5_ASAP7_75t_L g187 ( .A(n_14), .B(n_160), .Y(n_187) );
NAND2xp5_ASAP7_75t_L g241 ( .A(n_15), .B(n_130), .Y(n_241) );
NAND2xp5_ASAP7_75t_L g236 ( .A(n_16), .B(n_237), .Y(n_236) );
CKINVDCx5p33_ASAP7_75t_R g170 ( .A(n_17), .Y(n_170) );
BUFx3_ASAP7_75t_L g105 ( .A(n_18), .Y(n_105) );
INVx1_ASAP7_75t_L g132 ( .A(n_18), .Y(n_132) );
NAND2xp5_ASAP7_75t_L g229 ( .A(n_19), .B(n_208), .Y(n_229) );
CKINVDCx5p33_ASAP7_75t_R g128 ( .A(n_20), .Y(n_128) );
OAI22xp5_ASAP7_75t_L g678 ( .A1(n_21), .A2(n_67), .B1(n_679), .B2(n_680), .Y(n_678) );
CKINVDCx5p33_ASAP7_75t_R g679 ( .A(n_21), .Y(n_679) );
BUFx10_ASAP7_75t_L g695 ( .A(n_22), .Y(n_695) );
INVx1_ASAP7_75t_L g494 ( .A(n_23), .Y(n_494) );
AOI22xp33_ASAP7_75t_L g592 ( .A1(n_23), .A2(n_61), .B1(n_593), .B2(n_596), .Y(n_592) );
NAND2xp5_ASAP7_75t_SL g224 ( .A(n_24), .B(n_225), .Y(n_224) );
INVx1_ASAP7_75t_L g708 ( .A(n_24), .Y(n_708) );
CKINVDCx5p33_ASAP7_75t_R g162 ( .A(n_25), .Y(n_162) );
OAI22xp5_ASAP7_75t_L g682 ( .A1(n_25), .A2(n_162), .B1(n_683), .B2(n_684), .Y(n_682) );
NAND2xp5_ASAP7_75t_SL g102 ( .A(n_26), .B(n_103), .Y(n_102) );
NAND2xp5_ASAP7_75t_SL g228 ( .A(n_27), .B(n_225), .Y(n_228) );
AOI22xp5_ASAP7_75t_L g715 ( .A1(n_27), .A2(n_490), .B1(n_716), .B2(n_720), .Y(n_715) );
AND2x2_ASAP7_75t_L g498 ( .A(n_28), .B(n_499), .Y(n_498) );
INVx1_ASAP7_75t_L g529 ( .A(n_28), .Y(n_529) );
AND2x2_ASAP7_75t_L g543 ( .A(n_28), .B(n_40), .Y(n_543) );
OAI22xp33_ASAP7_75t_L g559 ( .A1(n_29), .A2(n_35), .B1(n_560), .B2(n_561), .Y(n_559) );
AOI22xp33_ASAP7_75t_L g576 ( .A1(n_29), .A2(n_58), .B1(n_577), .B2(n_585), .Y(n_576) );
NAND2xp5_ASAP7_75t_L g207 ( .A(n_30), .B(n_208), .Y(n_207) );
NAND2xp33_ASAP7_75t_L g242 ( .A(n_31), .B(n_117), .Y(n_242) );
A2O1A1Ixp33_ASAP7_75t_L g156 ( .A1(n_32), .A2(n_157), .B(n_159), .C(n_163), .Y(n_156) );
INVx1_ASAP7_75t_L g96 ( .A(n_33), .Y(n_96) );
INVx2_ASAP7_75t_L g502 ( .A(n_34), .Y(n_502) );
AOI22xp33_ASAP7_75t_L g606 ( .A1(n_35), .A2(n_51), .B1(n_593), .B2(n_607), .Y(n_606) );
XNOR2xp5_ASAP7_75t_L g489 ( .A(n_36), .B(n_490), .Y(n_489) );
NAND2xp5_ASAP7_75t_L g226 ( .A(n_37), .B(n_212), .Y(n_226) );
NAND2xp5_ASAP7_75t_SL g185 ( .A(n_38), .B(n_186), .Y(n_185) );
NAND2xp5_ASAP7_75t_L g113 ( .A(n_39), .B(n_114), .Y(n_113) );
INVx2_ASAP7_75t_L g499 ( .A(n_40), .Y(n_499) );
NAND2xp5_ASAP7_75t_L g539 ( .A(n_40), .B(n_529), .Y(n_539) );
AO221x1_ASAP7_75t_L g249 ( .A1(n_41), .A2(n_68), .B1(n_172), .B2(n_225), .C(n_250), .Y(n_249) );
NAND2xp5_ASAP7_75t_SL g133 ( .A(n_42), .B(n_108), .Y(n_133) );
AND2x4_ASAP7_75t_L g95 ( .A(n_43), .B(n_96), .Y(n_95) );
HB1xp67_ASAP7_75t_L g665 ( .A(n_43), .Y(n_665) );
NAND3xp33_ASAP7_75t_L g213 ( .A(n_44), .B(n_163), .C(n_214), .Y(n_213) );
INVx1_ASAP7_75t_L g583 ( .A(n_45), .Y(n_583) );
INVx1_ASAP7_75t_L g590 ( .A(n_45), .Y(n_590) );
INVxp67_ASAP7_75t_SL g503 ( .A(n_46), .Y(n_503) );
INVx1_ASAP7_75t_L g150 ( .A(n_47), .Y(n_150) );
INVx1_ASAP7_75t_L g100 ( .A(n_48), .Y(n_100) );
CKINVDCx5p33_ASAP7_75t_R g167 ( .A(n_49), .Y(n_167) );
A2O1A1Ixp33_ASAP7_75t_L g176 ( .A1(n_50), .A2(n_177), .B(n_178), .C(n_180), .Y(n_176) );
INVxp67_ASAP7_75t_SL g516 ( .A(n_51), .Y(n_516) );
INVx2_ASAP7_75t_L g179 ( .A(n_52), .Y(n_179) );
NAND2xp5_ASAP7_75t_L g142 ( .A(n_53), .B(n_98), .Y(n_142) );
AOI22xp5_ASAP7_75t_L g668 ( .A1(n_54), .A2(n_669), .B1(n_670), .B2(n_671), .Y(n_668) );
INVx3_ASAP7_75t_L g669 ( .A(n_54), .Y(n_669) );
INVx1_ASAP7_75t_L g558 ( .A(n_55), .Y(n_558) );
OAI21xp5_ASAP7_75t_L g641 ( .A1(n_55), .A2(n_642), .B(n_645), .Y(n_641) );
OAI211xp5_ASAP7_75t_L g540 ( .A1(n_56), .A2(n_541), .B(n_546), .C(n_551), .Y(n_540) );
INVx1_ASAP7_75t_L g624 ( .A(n_56), .Y(n_624) );
NAND2xp5_ASAP7_75t_L g106 ( .A(n_57), .B(n_107), .Y(n_106) );
INVxp67_ASAP7_75t_SL g512 ( .A(n_58), .Y(n_512) );
AND2x2_ASAP7_75t_L g120 ( .A(n_59), .B(n_98), .Y(n_120) );
INVx1_ASAP7_75t_L g257 ( .A(n_60), .Y(n_257) );
INVxp33_ASAP7_75t_SL g616 ( .A(n_62), .Y(n_616) );
OAI22xp33_ASAP7_75t_L g253 ( .A1(n_63), .A2(n_66), .B1(n_103), .B2(n_160), .Y(n_253) );
NAND2xp5_ASAP7_75t_L g210 ( .A(n_64), .B(n_163), .Y(n_210) );
INVx1_ASAP7_75t_L g554 ( .A(n_65), .Y(n_554) );
INVx1_ASAP7_75t_L g680 ( .A(n_67), .Y(n_680) );
AND2x2_ASAP7_75t_L g189 ( .A(n_69), .B(n_190), .Y(n_189) );
INVx1_ASAP7_75t_L g110 ( .A(n_70), .Y(n_110) );
BUFx3_ASAP7_75t_L g135 ( .A(n_70), .Y(n_135) );
INVx1_ASAP7_75t_L g182 ( .A(n_70), .Y(n_182) );
NAND2xp5_ASAP7_75t_SL g219 ( .A(n_71), .B(n_220), .Y(n_219) );
NAND2xp5_ASAP7_75t_L g173 ( .A(n_72), .B(n_174), .Y(n_173) );
AND2x2_ASAP7_75t_L g501 ( .A(n_73), .B(n_502), .Y(n_501) );
INVx2_ASAP7_75t_L g508 ( .A(n_73), .Y(n_508) );
INVxp67_ASAP7_75t_SL g525 ( .A(n_73), .Y(n_525) );
NAND2xp5_ASAP7_75t_SL g206 ( .A(n_74), .B(n_108), .Y(n_206) );
NAND2xp5_ASAP7_75t_L g243 ( .A(n_75), .B(n_98), .Y(n_243) );
INVx2_ASAP7_75t_L g573 ( .A(n_76), .Y(n_573) );
CKINVDCx5p33_ASAP7_75t_R g216 ( .A(n_77), .Y(n_216) );
AOI21xp33_ASAP7_75t_SL g78 ( .A1(n_79), .A2(n_478), .B(n_488), .Y(n_78) );
INVx1_ASAP7_75t_L g79 ( .A(n_80), .Y(n_79) );
INVx1_ASAP7_75t_L g80 ( .A(n_81), .Y(n_80) );
NAND4xp75_ASAP7_75t_L g81 ( .A(n_82), .B(n_344), .C(n_398), .D(n_443), .Y(n_81) );
AND2x2_ASAP7_75t_L g82 ( .A(n_83), .B(n_329), .Y(n_82) );
NOR3xp33_ASAP7_75t_L g83 ( .A(n_84), .B(n_275), .C(n_310), .Y(n_83) );
OAI21xp5_ASAP7_75t_L g84 ( .A1(n_85), .A2(n_200), .B(n_244), .Y(n_84) );
NOR2x1_ASAP7_75t_L g85 ( .A(n_86), .B(n_194), .Y(n_85) );
NOR2xp33_ASAP7_75t_SL g86 ( .A(n_87), .B(n_143), .Y(n_86) );
OR2x2_ASAP7_75t_L g422 ( .A(n_87), .B(n_386), .Y(n_422) );
INVx1_ASAP7_75t_L g433 ( .A(n_87), .Y(n_433) );
OR2x2_ASAP7_75t_L g87 ( .A(n_88), .B(n_121), .Y(n_87) );
AND2x2_ASAP7_75t_L g199 ( .A(n_88), .B(n_175), .Y(n_199) );
NAND2xp5_ASAP7_75t_L g271 ( .A(n_88), .B(n_272), .Y(n_271) );
NAND2xp5_ASAP7_75t_L g395 ( .A(n_88), .B(n_274), .Y(n_395) );
INVx2_ASAP7_75t_L g88 ( .A(n_89), .Y(n_88) );
AND2x2_ASAP7_75t_L g296 ( .A(n_89), .B(n_175), .Y(n_296) );
INVx2_ASAP7_75t_L g89 ( .A(n_90), .Y(n_89) );
OR2x2_ASAP7_75t_L g320 ( .A(n_90), .B(n_175), .Y(n_320) );
INVx1_ASAP7_75t_L g324 ( .A(n_90), .Y(n_324) );
AND2x2_ASAP7_75t_L g343 ( .A(n_90), .B(n_123), .Y(n_343) );
AND2x2_ASAP7_75t_L g377 ( .A(n_90), .B(n_122), .Y(n_377) );
NAND2x1p5_ASAP7_75t_L g90 ( .A(n_91), .B(n_111), .Y(n_90) );
NAND2x1_ASAP7_75t_L g91 ( .A(n_92), .B(n_101), .Y(n_91) );
AOI21x1_ASAP7_75t_L g111 ( .A1(n_92), .A2(n_112), .B(n_120), .Y(n_111) );
O2A1O1Ixp5_ASAP7_75t_L g204 ( .A1(n_92), .A2(n_205), .B(n_209), .C(n_215), .Y(n_204) );
AND2x4_ASAP7_75t_L g92 ( .A(n_93), .B(n_97), .Y(n_92) );
AOI21xp33_ASAP7_75t_L g192 ( .A1(n_93), .A2(n_189), .B(n_193), .Y(n_192) );
OAI21xp5_ASAP7_75t_L g234 ( .A1(n_93), .A2(n_235), .B(n_240), .Y(n_234) );
INVx2_ASAP7_75t_L g93 ( .A(n_94), .Y(n_93) );
NOR2xp33_ASAP7_75t_L g230 ( .A(n_94), .B(n_98), .Y(n_230) );
NOR2xp33_ASAP7_75t_R g254 ( .A(n_94), .B(n_255), .Y(n_254) );
INVx3_ASAP7_75t_L g94 ( .A(n_95), .Y(n_94) );
BUFx6f_ASAP7_75t_SL g141 ( .A(n_95), .Y(n_141) );
INVx2_ASAP7_75t_L g154 ( .A(n_95), .Y(n_154) );
INVx1_ASAP7_75t_L g483 ( .A(n_95), .Y(n_483) );
HB1xp67_ASAP7_75t_L g663 ( .A(n_96), .Y(n_663) );
INVx2_ASAP7_75t_L g97 ( .A(n_98), .Y(n_97) );
INVxp67_ASAP7_75t_SL g221 ( .A(n_98), .Y(n_221) );
INVx1_ASAP7_75t_L g233 ( .A(n_98), .Y(n_233) );
BUFx6f_ASAP7_75t_L g98 ( .A(n_99), .Y(n_98) );
BUFx2_ASAP7_75t_L g125 ( .A(n_99), .Y(n_125) );
INVx1_ASAP7_75t_L g191 ( .A(n_99), .Y(n_191) );
INVx1_ASAP7_75t_L g152 ( .A(n_100), .Y(n_152) );
AOI21xp5_ASAP7_75t_SL g101 ( .A1(n_102), .A2(n_106), .B(n_109), .Y(n_101) );
INVx2_ASAP7_75t_L g103 ( .A(n_104), .Y(n_103) );
INVx2_ASAP7_75t_L g108 ( .A(n_104), .Y(n_108) );
INVx2_ASAP7_75t_L g114 ( .A(n_104), .Y(n_114) );
INVx2_ASAP7_75t_L g104 ( .A(n_105), .Y(n_104) );
BUFx6f_ASAP7_75t_L g117 ( .A(n_105), .Y(n_117) );
BUFx6f_ASAP7_75t_L g161 ( .A(n_105), .Y(n_161) );
INVx2_ASAP7_75t_SL g107 ( .A(n_108), .Y(n_107) );
INVx2_ASAP7_75t_SL g487 ( .A(n_109), .Y(n_487) );
BUFx3_ASAP7_75t_L g109 ( .A(n_110), .Y(n_109) );
INVx1_ASAP7_75t_L g119 ( .A(n_110), .Y(n_119) );
AOI21xp5_ASAP7_75t_L g112 ( .A1(n_113), .A2(n_115), .B(n_118), .Y(n_112) );
INVx2_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
INVx3_ASAP7_75t_L g208 ( .A(n_117), .Y(n_208) );
INVx2_ASAP7_75t_L g212 ( .A(n_117), .Y(n_212) );
INVx3_ASAP7_75t_L g250 ( .A(n_117), .Y(n_250) );
AOI21xp5_ASAP7_75t_L g136 ( .A1(n_118), .A2(n_137), .B(n_140), .Y(n_136) );
INVx1_ASAP7_75t_L g188 ( .A(n_118), .Y(n_188) );
BUFx10_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
AND2x2_ASAP7_75t_L g325 ( .A(n_121), .B(n_272), .Y(n_325) );
AND2x2_ASAP7_75t_L g397 ( .A(n_121), .B(n_146), .Y(n_397) );
OR2x2_ASAP7_75t_L g458 ( .A(n_121), .B(n_309), .Y(n_458) );
INVx2_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
INVx1_ASAP7_75t_L g262 ( .A(n_122), .Y(n_262) );
INVx1_ASAP7_75t_L g286 ( .A(n_122), .Y(n_286) );
INVx2_ASAP7_75t_L g122 ( .A(n_123), .Y(n_122) );
INVxp33_ASAP7_75t_L g419 ( .A(n_123), .Y(n_419) );
OAI21x1_ASAP7_75t_L g123 ( .A1(n_124), .A2(n_126), .B(n_142), .Y(n_123) );
BUFx3_ASAP7_75t_L g124 ( .A(n_125), .Y(n_124) );
INVxp67_ASAP7_75t_L g193 ( .A(n_125), .Y(n_193) );
OAI21x1_ASAP7_75t_L g126 ( .A1(n_127), .A2(n_136), .B(n_141), .Y(n_126) );
O2A1O1Ixp5_ASAP7_75t_L g127 ( .A1(n_128), .A2(n_129), .B(n_133), .C(n_134), .Y(n_127) );
INVx2_ASAP7_75t_L g129 ( .A(n_130), .Y(n_129) );
INVx2_ASAP7_75t_L g158 ( .A(n_130), .Y(n_158) );
NOR2xp33_ASAP7_75t_L g169 ( .A(n_130), .B(n_170), .Y(n_169) );
INVx3_ASAP7_75t_L g130 ( .A(n_131), .Y(n_130) );
BUFx6f_ASAP7_75t_L g225 ( .A(n_131), .Y(n_225) );
INVx2_ASAP7_75t_L g131 ( .A(n_132), .Y(n_131) );
BUFx6f_ASAP7_75t_L g139 ( .A(n_132), .Y(n_139) );
AOI21xp5_ASAP7_75t_L g205 ( .A1(n_134), .A2(n_206), .B(n_207), .Y(n_205) );
AOI21xp5_ASAP7_75t_L g227 ( .A1(n_134), .A2(n_228), .B(n_229), .Y(n_227) );
INVx1_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
INVx2_ASAP7_75t_L g163 ( .A(n_135), .Y(n_163) );
INVx2_ASAP7_75t_L g172 ( .A(n_135), .Y(n_172) );
INVx2_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
INVx1_ASAP7_75t_L g168 ( .A(n_139), .Y(n_168) );
INVx2_ASAP7_75t_L g186 ( .A(n_139), .Y(n_186) );
INVx2_ASAP7_75t_L g214 ( .A(n_139), .Y(n_214) );
INVx1_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
AND2x2_ASAP7_75t_L g342 ( .A(n_144), .B(n_343), .Y(n_342) );
AND2x2_ASAP7_75t_L g144 ( .A(n_145), .B(n_175), .Y(n_144) );
INVx2_ASAP7_75t_L g274 ( .A(n_145), .Y(n_274) );
OR2x2_ASAP7_75t_L g308 ( .A(n_145), .B(n_309), .Y(n_308) );
AND2x2_ASAP7_75t_L g366 ( .A(n_145), .B(n_309), .Y(n_366) );
AND2x2_ASAP7_75t_L g463 ( .A(n_145), .B(n_419), .Y(n_463) );
INVx3_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
NAND2xp5_ASAP7_75t_L g288 ( .A(n_146), .B(n_289), .Y(n_288) );
AO21x2_ASAP7_75t_L g146 ( .A1(n_147), .A2(n_155), .B(n_164), .Y(n_146) );
AO21x1_ASAP7_75t_SL g198 ( .A1(n_147), .A2(n_155), .B(n_164), .Y(n_198) );
INVxp67_ASAP7_75t_SL g147 ( .A(n_148), .Y(n_147) );
OAI21x1_ASAP7_75t_SL g164 ( .A1(n_148), .A2(n_165), .B(n_173), .Y(n_164) );
NAND2xp5_ASAP7_75t_L g148 ( .A(n_149), .B(n_153), .Y(n_148) );
INVx2_ASAP7_75t_L g174 ( .A(n_149), .Y(n_174) );
AO21x2_ASAP7_75t_L g149 ( .A1(n_150), .A2(n_151), .B(n_152), .Y(n_149) );
AOI21x1_ASAP7_75t_L g255 ( .A1(n_150), .A2(n_151), .B(n_152), .Y(n_255) );
INVx2_ASAP7_75t_SL g153 ( .A(n_154), .Y(n_153) );
INVx1_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
INVx2_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
NOR2xp33_ASAP7_75t_L g159 ( .A(n_160), .B(n_162), .Y(n_159) );
INVx2_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
INVx2_ASAP7_75t_L g237 ( .A(n_161), .Y(n_237) );
OAI21xp5_ASAP7_75t_L g165 ( .A1(n_166), .A2(n_169), .B(n_171), .Y(n_165) );
NOR2xp33_ASAP7_75t_L g166 ( .A(n_167), .B(n_168), .Y(n_166) );
INVx1_ASAP7_75t_L g177 ( .A(n_168), .Y(n_177) );
AOI21xp5_ASAP7_75t_L g223 ( .A1(n_171), .A2(n_224), .B(n_226), .Y(n_223) );
INVx1_ASAP7_75t_L g171 ( .A(n_172), .Y(n_171) );
INVx1_ASAP7_75t_L g272 ( .A(n_175), .Y(n_272) );
INVx1_ASAP7_75t_L g289 ( .A(n_175), .Y(n_289) );
INVx2_ASAP7_75t_L g309 ( .A(n_175), .Y(n_309) );
AO21x2_ASAP7_75t_L g175 ( .A1(n_176), .A2(n_183), .B(n_192), .Y(n_175) );
NOR2xp67_ASAP7_75t_L g178 ( .A(n_177), .B(n_179), .Y(n_178) );
INVx1_ASAP7_75t_L g180 ( .A(n_181), .Y(n_180) );
AOI21xp5_ASAP7_75t_L g240 ( .A1(n_181), .A2(n_241), .B(n_242), .Y(n_240) );
BUFx3_ASAP7_75t_L g181 ( .A(n_182), .Y(n_181) );
INVx2_ASAP7_75t_L g239 ( .A(n_182), .Y(n_239) );
AOI21xp5_ASAP7_75t_L g183 ( .A1(n_184), .A2(n_188), .B(n_189), .Y(n_183) );
NAND2xp5_ASAP7_75t_L g184 ( .A(n_185), .B(n_187), .Y(n_184) );
INVx2_ASAP7_75t_L g486 ( .A(n_186), .Y(n_486) );
INVx2_ASAP7_75t_L g190 ( .A(n_191), .Y(n_190) );
NOR2xp33_ASAP7_75t_L g215 ( .A(n_193), .B(n_216), .Y(n_215) );
INVx2_ASAP7_75t_L g194 ( .A(n_195), .Y(n_194) );
INVx2_ASAP7_75t_L g195 ( .A(n_196), .Y(n_195) );
OAI21xp5_ASAP7_75t_L g363 ( .A1(n_196), .A2(n_364), .B(n_367), .Y(n_363) );
AND2x4_ASAP7_75t_L g196 ( .A(n_197), .B(n_199), .Y(n_196) );
AND2x2_ASAP7_75t_L g360 ( .A(n_197), .B(n_312), .Y(n_360) );
INVx5_ASAP7_75t_L g386 ( .A(n_197), .Y(n_386) );
AND2x4_ASAP7_75t_SL g410 ( .A(n_197), .B(n_411), .Y(n_410) );
AND2x2_ASAP7_75t_L g437 ( .A(n_197), .B(n_350), .Y(n_437) );
NAND2xp5_ASAP7_75t_L g471 ( .A(n_197), .B(n_421), .Y(n_471) );
OR2x2_ASAP7_75t_L g474 ( .A(n_197), .B(n_458), .Y(n_474) );
BUFx6f_ASAP7_75t_L g197 ( .A(n_198), .Y(n_197) );
INVxp67_ASAP7_75t_L g407 ( .A(n_198), .Y(n_407) );
NAND2xp5_ASAP7_75t_L g260 ( .A(n_199), .B(n_261), .Y(n_260) );
AND2x2_ASAP7_75t_L g466 ( .A(n_199), .B(n_386), .Y(n_466) );
OAI22xp5_ASAP7_75t_L g347 ( .A1(n_200), .A2(n_348), .B1(n_352), .B2(n_355), .Y(n_347) );
INVx2_ASAP7_75t_L g200 ( .A(n_201), .Y(n_200) );
AND2x2_ASAP7_75t_L g201 ( .A(n_202), .B(n_217), .Y(n_201) );
NOR2x1_ASAP7_75t_SL g245 ( .A(n_202), .B(n_246), .Y(n_245) );
BUFx2_ASAP7_75t_SL g202 ( .A(n_203), .Y(n_202) );
INVx2_ASAP7_75t_L g279 ( .A(n_203), .Y(n_279) );
NAND2xp5_ASAP7_75t_L g282 ( .A(n_203), .B(n_283), .Y(n_282) );
INVx1_ASAP7_75t_L g362 ( .A(n_203), .Y(n_362) );
AND2x2_ASAP7_75t_L g404 ( .A(n_203), .B(n_231), .Y(n_404) );
INVx2_ASAP7_75t_L g203 ( .A(n_204), .Y(n_203) );
OAI21xp5_ASAP7_75t_L g209 ( .A1(n_210), .A2(n_211), .B(n_213), .Y(n_209) );
INVx2_ASAP7_75t_L g211 ( .A(n_212), .Y(n_211) );
AND2x4_ASAP7_75t_SL g303 ( .A(n_217), .B(n_304), .Y(n_303) );
NAND2xp5_ASAP7_75t_L g311 ( .A(n_217), .B(n_312), .Y(n_311) );
AND2x2_ASAP7_75t_L g361 ( .A(n_217), .B(n_362), .Y(n_361) );
AND2x2_ASAP7_75t_L g217 ( .A(n_218), .B(n_231), .Y(n_217) );
INVx3_ASAP7_75t_L g267 ( .A(n_218), .Y(n_267) );
OR2x2_ASAP7_75t_L g299 ( .A(n_218), .B(n_248), .Y(n_299) );
HB1xp67_ASAP7_75t_L g327 ( .A(n_218), .Y(n_327) );
AND2x2_ASAP7_75t_L g424 ( .A(n_218), .B(n_247), .Y(n_424) );
NOR2xp33_ASAP7_75t_L g447 ( .A(n_218), .B(n_231), .Y(n_447) );
AND2x4_ASAP7_75t_L g218 ( .A(n_219), .B(n_222), .Y(n_218) );
INVx1_ASAP7_75t_L g220 ( .A(n_221), .Y(n_220) );
OAI21xp5_ASAP7_75t_L g222 ( .A1(n_223), .A2(n_227), .B(n_230), .Y(n_222) );
INVx1_ASAP7_75t_L g247 ( .A(n_231), .Y(n_247) );
HB1xp67_ASAP7_75t_L g268 ( .A(n_231), .Y(n_268) );
INVx1_ASAP7_75t_L g283 ( .A(n_231), .Y(n_283) );
INVx1_ASAP7_75t_L g315 ( .A(n_231), .Y(n_315) );
OA21x2_ASAP7_75t_L g231 ( .A1(n_232), .A2(n_234), .B(n_243), .Y(n_231) );
INVx1_ASAP7_75t_SL g232 ( .A(n_233), .Y(n_232) );
AOI21xp5_ASAP7_75t_L g235 ( .A1(n_236), .A2(n_238), .B(n_239), .Y(n_235) );
INVx2_ASAP7_75t_L g252 ( .A(n_239), .Y(n_252) );
AOI22xp5_ASAP7_75t_L g244 ( .A1(n_245), .A2(n_259), .B1(n_263), .B2(n_269), .Y(n_244) );
NAND2xp5_ASAP7_75t_L g388 ( .A(n_245), .B(n_327), .Y(n_388) );
OR2x2_ASAP7_75t_L g368 ( .A(n_246), .B(n_316), .Y(n_368) );
OR2x2_ASAP7_75t_L g246 ( .A(n_247), .B(n_248), .Y(n_246) );
AND2x2_ASAP7_75t_L g277 ( .A(n_248), .B(n_278), .Y(n_277) );
INVx2_ASAP7_75t_SL g304 ( .A(n_248), .Y(n_304) );
BUFx3_ASAP7_75t_L g312 ( .A(n_248), .Y(n_312) );
AND2x2_ASAP7_75t_L g393 ( .A(n_248), .B(n_267), .Y(n_393) );
AND2x2_ASAP7_75t_L g448 ( .A(n_248), .B(n_279), .Y(n_448) );
AND2x2_ASAP7_75t_L g453 ( .A(n_248), .B(n_266), .Y(n_453) );
AO31x2_ASAP7_75t_L g248 ( .A1(n_249), .A2(n_251), .A3(n_254), .B(n_256), .Y(n_248) );
NAND2xp5_ASAP7_75t_L g251 ( .A(n_252), .B(n_253), .Y(n_251) );
INVx2_ASAP7_75t_L g258 ( .A(n_255), .Y(n_258) );
NOR2xp33_ASAP7_75t_L g256 ( .A(n_257), .B(n_258), .Y(n_256) );
AOI22xp33_ASAP7_75t_L g439 ( .A1(n_259), .A2(n_440), .B1(n_441), .B2(n_442), .Y(n_439) );
INVx2_ASAP7_75t_SL g259 ( .A(n_260), .Y(n_259) );
OR2x2_ASAP7_75t_L g333 ( .A(n_261), .B(n_334), .Y(n_333) );
NOR2xp33_ASAP7_75t_SL g449 ( .A(n_261), .B(n_450), .Y(n_449) );
INVx2_ASAP7_75t_L g261 ( .A(n_262), .Y(n_261) );
OR2x2_ASAP7_75t_L g292 ( .A(n_262), .B(n_271), .Y(n_292) );
AND2x4_ASAP7_75t_SL g318 ( .A(n_262), .B(n_319), .Y(n_318) );
NAND2xp5_ASAP7_75t_L g365 ( .A(n_262), .B(n_366), .Y(n_365) );
BUFx2_ASAP7_75t_L g379 ( .A(n_262), .Y(n_379) );
HB1xp67_ASAP7_75t_L g263 ( .A(n_264), .Y(n_263) );
AND2x2_ASAP7_75t_L g264 ( .A(n_265), .B(n_268), .Y(n_264) );
INVx1_ASAP7_75t_L g265 ( .A(n_266), .Y(n_265) );
AND2x2_ASAP7_75t_L g354 ( .A(n_266), .B(n_304), .Y(n_354) );
INVx1_ASAP7_75t_L g403 ( .A(n_266), .Y(n_403) );
INVx2_ASAP7_75t_L g266 ( .A(n_267), .Y(n_266) );
NAND2xp5_ASAP7_75t_L g316 ( .A(n_267), .B(n_279), .Y(n_316) );
OR2x2_ASAP7_75t_L g339 ( .A(n_268), .B(n_278), .Y(n_339) );
INVx1_ASAP7_75t_L g269 ( .A(n_270), .Y(n_269) );
OR2x2_ASAP7_75t_L g270 ( .A(n_271), .B(n_273), .Y(n_270) );
INVx1_ASAP7_75t_L g356 ( .A(n_271), .Y(n_356) );
OR2x2_ASAP7_75t_L g381 ( .A(n_271), .B(n_375), .Y(n_381) );
BUFx2_ASAP7_75t_SL g273 ( .A(n_274), .Y(n_273) );
INVx2_ASAP7_75t_L g375 ( .A(n_274), .Y(n_375) );
NAND3xp33_ASAP7_75t_SL g275 ( .A(n_276), .B(n_290), .C(n_300), .Y(n_275) );
OAI21xp33_ASAP7_75t_L g276 ( .A1(n_277), .A2(n_280), .B(n_284), .Y(n_276) );
AND2x4_ASAP7_75t_L g423 ( .A(n_277), .B(n_424), .Y(n_423) );
AND2x2_ASAP7_75t_L g335 ( .A(n_278), .B(n_303), .Y(n_335) );
INVx1_ASAP7_75t_L g391 ( .A(n_278), .Y(n_391) );
INVx2_ASAP7_75t_L g278 ( .A(n_279), .Y(n_278) );
INVx2_ASAP7_75t_L g280 ( .A(n_281), .Y(n_280) );
BUFx2_ASAP7_75t_L g281 ( .A(n_282), .Y(n_281) );
OR2x2_ASAP7_75t_L g298 ( .A(n_282), .B(n_299), .Y(n_298) );
INVx2_ASAP7_75t_L g328 ( .A(n_282), .Y(n_328) );
AOI22xp5_ASAP7_75t_L g445 ( .A1(n_284), .A2(n_446), .B1(n_449), .B2(n_451), .Y(n_445) );
AND2x2_ASAP7_75t_L g284 ( .A(n_285), .B(n_287), .Y(n_284) );
OR2x2_ASAP7_75t_L g294 ( .A(n_285), .B(n_295), .Y(n_294) );
INVx1_ASAP7_75t_L g307 ( .A(n_285), .Y(n_307) );
INVx1_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
OR2x2_ASAP7_75t_L g412 ( .A(n_286), .B(n_320), .Y(n_412) );
AND2x2_ASAP7_75t_L g421 ( .A(n_286), .B(n_324), .Y(n_421) );
INVx1_ASAP7_75t_L g334 ( .A(n_287), .Y(n_334) );
INVx1_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
OAI21xp5_ASAP7_75t_L g290 ( .A1(n_291), .A2(n_293), .B(n_297), .Y(n_290) );
INVxp67_ASAP7_75t_SL g291 ( .A(n_292), .Y(n_291) );
INVx2_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
INVx1_ASAP7_75t_L g295 ( .A(n_296), .Y(n_295) );
AND2x4_ASAP7_75t_L g380 ( .A(n_296), .B(n_375), .Y(n_380) );
INVx1_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
INVx2_ASAP7_75t_L g411 ( .A(n_299), .Y(n_411) );
NAND2xp5_ASAP7_75t_L g300 ( .A(n_301), .B(n_305), .Y(n_300) );
INVxp67_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
INVx2_ASAP7_75t_L g302 ( .A(n_303), .Y(n_302) );
NAND2xp5_ASAP7_75t_L g314 ( .A(n_304), .B(n_315), .Y(n_314) );
INVx1_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
OR2x2_ASAP7_75t_L g306 ( .A(n_307), .B(n_308), .Y(n_306) );
NAND2xp5_ASAP7_75t_L g455 ( .A(n_308), .B(n_456), .Y(n_455) );
INVx1_ASAP7_75t_L g349 ( .A(n_309), .Y(n_349) );
AND2x2_ASAP7_75t_L g418 ( .A(n_309), .B(n_419), .Y(n_418) );
A2O1A1Ixp33_ASAP7_75t_L g310 ( .A1(n_311), .A2(n_313), .B(n_317), .C(n_321), .Y(n_310) );
INVx1_ASAP7_75t_L g428 ( .A(n_312), .Y(n_428) );
INVx1_ASAP7_75t_L g441 ( .A(n_313), .Y(n_441) );
OR2x2_ASAP7_75t_L g313 ( .A(n_314), .B(n_316), .Y(n_313) );
INVx2_ASAP7_75t_L g414 ( .A(n_315), .Y(n_414) );
INVx2_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
INVx1_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
INVx2_ASAP7_75t_L g387 ( .A(n_320), .Y(n_387) );
NAND2xp5_ASAP7_75t_L g321 ( .A(n_322), .B(n_326), .Y(n_321) );
AND2x4_ASAP7_75t_L g322 ( .A(n_323), .B(n_325), .Y(n_322) );
OA21x2_ASAP7_75t_L g357 ( .A1(n_323), .A2(n_358), .B(n_363), .Y(n_357) );
INVx1_ASAP7_75t_L g457 ( .A(n_323), .Y(n_457) );
INVx3_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
INVx2_ASAP7_75t_L g426 ( .A(n_326), .Y(n_426) );
AND2x2_ASAP7_75t_L g326 ( .A(n_327), .B(n_328), .Y(n_326) );
NOR2xp33_ASAP7_75t_L g336 ( .A(n_327), .B(n_337), .Y(n_336) );
A2O1A1Ixp33_ASAP7_75t_L g329 ( .A1(n_330), .A2(n_335), .B(n_336), .C(n_340), .Y(n_329) );
INVxp67_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
NAND2xp5_ASAP7_75t_L g340 ( .A(n_331), .B(n_341), .Y(n_340) );
INVx1_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
INVx1_ASAP7_75t_L g332 ( .A(n_333), .Y(n_332) );
INVx2_ASAP7_75t_L g464 ( .A(n_335), .Y(n_464) );
INVx1_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
AOI22xp5_ASAP7_75t_L g465 ( .A1(n_338), .A2(n_466), .B1(n_467), .B2(n_470), .Y(n_465) );
INVx1_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
OR2x6_ASAP7_75t_L g352 ( .A(n_339), .B(n_353), .Y(n_352) );
OR2x2_ASAP7_75t_L g427 ( .A(n_339), .B(n_428), .Y(n_427) );
INVx1_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
INVx4_ASAP7_75t_L g351 ( .A(n_343), .Y(n_351) );
NOR2x1p5_ASAP7_75t_L g344 ( .A(n_345), .B(n_369), .Y(n_344) );
NAND2x1_ASAP7_75t_L g345 ( .A(n_346), .B(n_357), .Y(n_345) );
INVx1_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
INVx1_ASAP7_75t_L g460 ( .A(n_348), .Y(n_460) );
NAND2x1_ASAP7_75t_L g348 ( .A(n_349), .B(n_350), .Y(n_348) );
INVx1_ASAP7_75t_L g450 ( .A(n_349), .Y(n_450) );
INVx6_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
OAI22xp5_ASAP7_75t_L g389 ( .A1(n_352), .A2(n_390), .B1(n_394), .B2(n_396), .Y(n_389) );
INVx1_ASAP7_75t_L g401 ( .A(n_352), .Y(n_401) );
INVx1_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
HB1xp67_ASAP7_75t_L g382 ( .A(n_354), .Y(n_382) );
INVx1_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
INVxp33_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
AND2x2_ASAP7_75t_L g359 ( .A(n_360), .B(n_361), .Y(n_359) );
NAND2xp5_ASAP7_75t_L g477 ( .A(n_360), .B(n_372), .Y(n_477) );
INVx2_ASAP7_75t_L g373 ( .A(n_362), .Y(n_373) );
AND2x2_ASAP7_75t_L g435 ( .A(n_362), .B(n_393), .Y(n_435) );
INVx1_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
INVx1_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
INVx2_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
AOI211x1_ASAP7_75t_L g370 ( .A1(n_371), .A2(n_382), .B(n_383), .C(n_389), .Y(n_370) );
OAI211xp5_ASAP7_75t_L g371 ( .A1(n_372), .A2(n_374), .B(n_378), .C(n_381), .Y(n_371) );
INVx1_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
INVx1_ASAP7_75t_L g440 ( .A(n_374), .Y(n_440) );
OR2x2_ASAP7_75t_L g374 ( .A(n_375), .B(n_376), .Y(n_374) );
INVx1_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
AND2x2_ASAP7_75t_L g406 ( .A(n_377), .B(n_407), .Y(n_406) );
NAND2x1_ASAP7_75t_SL g378 ( .A(n_379), .B(n_380), .Y(n_378) );
NOR2xp33_ASAP7_75t_L g383 ( .A(n_384), .B(n_388), .Y(n_383) );
INVx1_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
AND2x2_ASAP7_75t_L g385 ( .A(n_386), .B(n_387), .Y(n_385) );
NAND2xp5_ASAP7_75t_L g420 ( .A(n_386), .B(n_421), .Y(n_420) );
AND2x2_ASAP7_75t_L g432 ( .A(n_386), .B(n_433), .Y(n_432) );
INVx1_ASAP7_75t_L g442 ( .A(n_390), .Y(n_442) );
OR2x2_ASAP7_75t_L g390 ( .A(n_391), .B(n_392), .Y(n_390) );
AND2x2_ASAP7_75t_L g469 ( .A(n_391), .B(n_453), .Y(n_469) );
INVx2_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
AND2x4_ASAP7_75t_L g459 ( .A(n_393), .B(n_404), .Y(n_459) );
HB1xp67_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
INVx1_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
NOR2x1_ASAP7_75t_L g398 ( .A(n_399), .B(n_430), .Y(n_398) );
NAND2xp5_ASAP7_75t_L g399 ( .A(n_400), .B(n_415), .Y(n_399) );
O2A1O1Ixp33_ASAP7_75t_SL g400 ( .A1(n_401), .A2(n_402), .B(n_405), .C(n_408), .Y(n_400) );
INVx1_ASAP7_75t_L g438 ( .A(n_402), .Y(n_438) );
AND2x2_ASAP7_75t_L g402 ( .A(n_403), .B(n_404), .Y(n_402) );
HB1xp67_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
NOR3xp33_ASAP7_75t_L g408 ( .A(n_409), .B(n_412), .C(n_413), .Y(n_408) );
INVx2_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
HB1xp67_ASAP7_75t_L g429 ( .A(n_412), .Y(n_429) );
NAND2xp5_ASAP7_75t_L g452 ( .A(n_413), .B(n_453), .Y(n_452) );
INVx2_ASAP7_75t_SL g413 ( .A(n_414), .Y(n_413) );
AOI21xp5_ASAP7_75t_L g415 ( .A1(n_416), .A2(n_423), .B(n_425), .Y(n_415) );
NAND3xp33_ASAP7_75t_SL g416 ( .A(n_417), .B(n_420), .C(n_422), .Y(n_416) );
INVx1_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
AOI22xp5_ASAP7_75t_L g472 ( .A1(n_421), .A2(n_473), .B1(n_475), .B2(n_476), .Y(n_472) );
AND2x4_ASAP7_75t_L g475 ( .A(n_424), .B(n_448), .Y(n_475) );
AOI21xp5_ASAP7_75t_L g425 ( .A1(n_426), .A2(n_427), .B(n_429), .Y(n_425) );
OAI221xp5_ASAP7_75t_L g430 ( .A1(n_431), .A2(n_434), .B1(n_436), .B2(n_438), .C(n_439), .Y(n_430) );
INVx1_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
INVx2_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
AOI22xp5_ASAP7_75t_L g454 ( .A1(n_435), .A2(n_455), .B1(n_459), .B2(n_460), .Y(n_454) );
INVxp67_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
NOR2x1_ASAP7_75t_SL g443 ( .A(n_444), .B(n_461), .Y(n_443) );
NAND2xp5_ASAP7_75t_L g444 ( .A(n_445), .B(n_454), .Y(n_444) );
AND2x4_ASAP7_75t_L g446 ( .A(n_447), .B(n_448), .Y(n_446) );
INVx1_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
AND2x2_ASAP7_75t_L g456 ( .A(n_457), .B(n_458), .Y(n_456) );
OAI211xp5_ASAP7_75t_L g461 ( .A1(n_462), .A2(n_464), .B(n_465), .C(n_472), .Y(n_461) );
INVx1_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
INVx1_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
INVx1_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
INVx2_ASAP7_75t_L g470 ( .A(n_471), .Y(n_470) );
INVx1_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
INVxp67_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
BUFx2_ASAP7_75t_L g478 ( .A(n_479), .Y(n_478) );
NOR2x1_ASAP7_75t_L g479 ( .A(n_480), .B(n_484), .Y(n_479) );
INVx1_ASAP7_75t_SL g480 ( .A(n_481), .Y(n_480) );
BUFx2_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
INVx1_ASAP7_75t_L g482 ( .A(n_483), .Y(n_482) );
AO21x2_ASAP7_75t_L g722 ( .A1(n_484), .A2(n_662), .B(n_723), .Y(n_722) );
NAND2xp5_ASAP7_75t_L g484 ( .A(n_485), .B(n_487), .Y(n_484) );
INVx1_ASAP7_75t_L g485 ( .A(n_486), .Y(n_485) );
OAI221xp5_ASAP7_75t_L g488 ( .A1(n_489), .A2(n_490), .B1(n_656), .B2(n_666), .C(n_715), .Y(n_488) );
OA21x2_ASAP7_75t_L g490 ( .A1(n_491), .A2(n_563), .B(n_567), .Y(n_490) );
NOR3xp33_ASAP7_75t_L g491 ( .A(n_492), .B(n_540), .C(n_559), .Y(n_491) );
NAND3xp33_ASAP7_75t_SL g492 ( .A(n_493), .B(n_509), .C(n_530), .Y(n_492) );
AOI22xp33_ASAP7_75t_L g493 ( .A1(n_494), .A2(n_495), .B1(n_503), .B2(n_504), .Y(n_493) );
AND2x4_ASAP7_75t_L g495 ( .A(n_496), .B(n_500), .Y(n_495) );
AND2x2_ASAP7_75t_L g504 ( .A(n_496), .B(n_505), .Y(n_504) );
INVx1_ASAP7_75t_L g496 ( .A(n_497), .Y(n_496) );
OR2x2_ASAP7_75t_L g560 ( .A(n_497), .B(n_544), .Y(n_560) );
INVx1_ASAP7_75t_L g562 ( .A(n_497), .Y(n_562) );
INVx1_ASAP7_75t_L g497 ( .A(n_498), .Y(n_497) );
AND2x2_ASAP7_75t_L g528 ( .A(n_499), .B(n_529), .Y(n_528) );
BUFx4f_ASAP7_75t_L g500 ( .A(n_501), .Y(n_500) );
BUFx6f_ASAP7_75t_L g511 ( .A(n_501), .Y(n_511) );
INVx2_ASAP7_75t_L g507 ( .A(n_502), .Y(n_507) );
INVx2_ASAP7_75t_L g520 ( .A(n_502), .Y(n_520) );
NAND2xp5_ASAP7_75t_L g545 ( .A(n_502), .B(n_508), .Y(n_545) );
BUFx6f_ASAP7_75t_L g505 ( .A(n_506), .Y(n_505) );
INVx5_ASAP7_75t_L g515 ( .A(n_506), .Y(n_515) );
AND2x4_ASAP7_75t_L g506 ( .A(n_507), .B(n_508), .Y(n_506) );
INVx1_ASAP7_75t_L g526 ( .A(n_507), .Y(n_526) );
INVx2_ASAP7_75t_L g521 ( .A(n_508), .Y(n_521) );
OAI221xp5_ASAP7_75t_L g509 ( .A1(n_510), .A2(n_512), .B1(n_513), .B2(n_516), .C(n_517), .Y(n_509) );
INVx3_ASAP7_75t_L g510 ( .A(n_511), .Y(n_510) );
BUFx12f_ASAP7_75t_SL g533 ( .A(n_511), .Y(n_533) );
OAI221xp5_ASAP7_75t_L g530 ( .A1(n_513), .A2(n_531), .B1(n_534), .B2(n_535), .C(n_536), .Y(n_530) );
INVx2_ASAP7_75t_SL g513 ( .A(n_514), .Y(n_513) );
INVx4_ASAP7_75t_L g514 ( .A(n_515), .Y(n_514) );
NAND2x1p5_ASAP7_75t_L g561 ( .A(n_518), .B(n_562), .Y(n_561) );
BUFx4f_ASAP7_75t_L g518 ( .A(n_519), .Y(n_518) );
INVx2_ASAP7_75t_L g549 ( .A(n_519), .Y(n_549) );
AND2x4_ASAP7_75t_L g519 ( .A(n_520), .B(n_521), .Y(n_519) );
BUFx3_ASAP7_75t_L g553 ( .A(n_520), .Y(n_553) );
INVx1_ASAP7_75t_L g557 ( .A(n_521), .Y(n_557) );
INVx4_ASAP7_75t_L g522 ( .A(n_523), .Y(n_522) );
INVx1_ASAP7_75t_L g537 ( .A(n_523), .Y(n_537) );
INVx5_ASAP7_75t_L g523 ( .A(n_524), .Y(n_523) );
AND2x4_ASAP7_75t_L g524 ( .A(n_525), .B(n_526), .Y(n_524) );
INVx1_ASAP7_75t_L g527 ( .A(n_528), .Y(n_527) );
INVx1_ASAP7_75t_L g531 ( .A(n_532), .Y(n_531) );
BUFx2_ASAP7_75t_L g532 ( .A(n_533), .Y(n_532) );
BUFx4_ASAP7_75t_L g538 ( .A(n_539), .Y(n_538) );
OR2x6_ASAP7_75t_L g541 ( .A(n_542), .B(n_544), .Y(n_541) );
INVx1_ASAP7_75t_L g550 ( .A(n_542), .Y(n_550) );
INVx1_ASAP7_75t_L g542 ( .A(n_543), .Y(n_542) );
AND2x2_ASAP7_75t_L g552 ( .A(n_543), .B(n_553), .Y(n_552) );
AND2x2_ASAP7_75t_L g555 ( .A(n_543), .B(n_556), .Y(n_555) );
BUFx6f_ASAP7_75t_L g544 ( .A(n_545), .Y(n_544) );
BUFx2_ASAP7_75t_L g546 ( .A(n_547), .Y(n_546) );
NAND2xp5_ASAP7_75t_L g547 ( .A(n_548), .B(n_550), .Y(n_547) );
INVx1_ASAP7_75t_L g548 ( .A(n_549), .Y(n_548) );
AOI22xp33_ASAP7_75t_SL g551 ( .A1(n_552), .A2(n_554), .B1(n_555), .B2(n_558), .Y(n_551) );
AOI22xp33_ASAP7_75t_L g645 ( .A1(n_554), .A2(n_646), .B1(n_651), .B2(n_655), .Y(n_645) );
INVx1_ASAP7_75t_L g556 ( .A(n_557), .Y(n_556) );
INVx1_ASAP7_75t_L g563 ( .A(n_564), .Y(n_563) );
INVx2_ASAP7_75t_L g564 ( .A(n_565), .Y(n_564) );
AND2x6_ASAP7_75t_L g570 ( .A(n_565), .B(n_571), .Y(n_570) );
INVx2_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
INVx1_ASAP7_75t_L g613 ( .A(n_566), .Y(n_613) );
OR2x2_ASAP7_75t_L g622 ( .A(n_566), .B(n_623), .Y(n_622) );
NOR3xp33_ASAP7_75t_L g567 ( .A(n_568), .B(n_631), .C(n_641), .Y(n_567) );
NAND2xp5_ASAP7_75t_SL g568 ( .A(n_569), .B(n_615), .Y(n_568) );
AOI33xp33_ASAP7_75t_L g569 ( .A1(n_570), .A2(n_576), .A3(n_592), .B1(n_602), .B2(n_606), .B3(n_610), .Y(n_569) );
AND2x2_ASAP7_75t_L g571 ( .A(n_572), .B(n_574), .Y(n_571) );
AND2x4_ASAP7_75t_L g614 ( .A(n_572), .B(n_575), .Y(n_614) );
BUFx2_ASAP7_75t_L g572 ( .A(n_573), .Y(n_572) );
OR2x6_ASAP7_75t_L g623 ( .A(n_573), .B(n_575), .Y(n_623) );
INVx1_ASAP7_75t_L g637 ( .A(n_573), .Y(n_637) );
INVx1_ASAP7_75t_L g574 ( .A(n_575), .Y(n_574) );
AND2x2_ASAP7_75t_L g636 ( .A(n_575), .B(n_637), .Y(n_636) );
OR2x2_ASAP7_75t_L g698 ( .A(n_575), .B(n_637), .Y(n_698) );
INVx2_ASAP7_75t_SL g577 ( .A(n_578), .Y(n_577) );
INVx1_ASAP7_75t_L g578 ( .A(n_579), .Y(n_578) );
BUFx12f_ASAP7_75t_L g579 ( .A(n_580), .Y(n_579) );
NAND2x1_ASAP7_75t_L g632 ( .A(n_580), .B(n_627), .Y(n_632) );
BUFx6f_ASAP7_75t_L g580 ( .A(n_581), .Y(n_580) );
AND2x2_ASAP7_75t_L g581 ( .A(n_582), .B(n_584), .Y(n_581) );
AND2x4_ASAP7_75t_L g601 ( .A(n_582), .B(n_591), .Y(n_601) );
INVx2_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
AND2x2_ASAP7_75t_L g595 ( .A(n_583), .B(n_584), .Y(n_595) );
INVx2_ASAP7_75t_L g591 ( .A(n_584), .Y(n_591) );
INVx2_ASAP7_75t_L g585 ( .A(n_586), .Y(n_585) );
INVx2_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
INVx3_ASAP7_75t_L g587 ( .A(n_588), .Y(n_587) );
INVx4_ASAP7_75t_L g588 ( .A(n_589), .Y(n_588) );
BUFx6f_ASAP7_75t_L g605 ( .A(n_589), .Y(n_605) );
BUFx3_ASAP7_75t_L g630 ( .A(n_589), .Y(n_630) );
AND2x4_ASAP7_75t_L g589 ( .A(n_590), .B(n_591), .Y(n_589) );
AND2x4_ASAP7_75t_L g620 ( .A(n_590), .B(n_621), .Y(n_620) );
INVx1_ASAP7_75t_L g654 ( .A(n_590), .Y(n_654) );
INVx3_ASAP7_75t_L g593 ( .A(n_594), .Y(n_593) );
INVx2_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
INVx1_ASAP7_75t_L g596 ( .A(n_597), .Y(n_596) );
INVx1_ASAP7_75t_L g597 ( .A(n_598), .Y(n_597) );
HB1xp67_ASAP7_75t_L g598 ( .A(n_599), .Y(n_598) );
BUFx6f_ASAP7_75t_SL g599 ( .A(n_600), .Y(n_599) );
BUFx6f_ASAP7_75t_L g609 ( .A(n_600), .Y(n_609) );
BUFx6f_ASAP7_75t_L g600 ( .A(n_601), .Y(n_600) );
BUFx6f_ASAP7_75t_L g640 ( .A(n_601), .Y(n_640) );
INVx2_ASAP7_75t_L g644 ( .A(n_601), .Y(n_644) );
INVx2_ASAP7_75t_L g603 ( .A(n_604), .Y(n_603) );
INVx2_ASAP7_75t_L g604 ( .A(n_605), .Y(n_604) );
INVx1_ASAP7_75t_L g607 ( .A(n_608), .Y(n_607) );
INVx1_ASAP7_75t_L g608 ( .A(n_609), .Y(n_608) );
CKINVDCx5p33_ASAP7_75t_R g610 ( .A(n_611), .Y(n_610) );
CKINVDCx8_ASAP7_75t_R g611 ( .A(n_612), .Y(n_611) );
AND2x6_ASAP7_75t_L g612 ( .A(n_613), .B(n_614), .Y(n_612) );
AND2x4_ASAP7_75t_L g635 ( .A(n_613), .B(n_636), .Y(n_635) );
AOI22xp33_ASAP7_75t_L g615 ( .A1(n_616), .A2(n_617), .B1(n_624), .B2(n_625), .Y(n_615) );
CKINVDCx5p33_ASAP7_75t_R g617 ( .A(n_618), .Y(n_617) );
OR2x6_ASAP7_75t_L g618 ( .A(n_619), .B(n_622), .Y(n_618) );
OR2x2_ASAP7_75t_L g633 ( .A(n_619), .B(n_634), .Y(n_633) );
INVx8_ASAP7_75t_L g619 ( .A(n_620), .Y(n_619) );
HB1xp67_ASAP7_75t_L g650 ( .A(n_621), .Y(n_650) );
INVx1_ASAP7_75t_L g696 ( .A(n_621), .Y(n_696) );
INVx2_ASAP7_75t_L g627 ( .A(n_622), .Y(n_627) );
BUFx2_ASAP7_75t_L g625 ( .A(n_626), .Y(n_625) );
AND2x4_ASAP7_75t_L g626 ( .A(n_627), .B(n_628), .Y(n_626) );
NAND2x1_ASAP7_75t_L g642 ( .A(n_627), .B(n_643), .Y(n_642) );
INVx1_ASAP7_75t_L g628 ( .A(n_629), .Y(n_628) );
INVx1_ASAP7_75t_L g629 ( .A(n_630), .Y(n_629) );
INVx2_ASAP7_75t_L g634 ( .A(n_635), .Y(n_634) );
AND2x4_ASAP7_75t_L g639 ( .A(n_635), .B(n_640), .Y(n_639) );
AND2x2_ASAP7_75t_L g648 ( .A(n_635), .B(n_649), .Y(n_648) );
AND2x4_ASAP7_75t_L g651 ( .A(n_635), .B(n_652), .Y(n_651) );
INVx1_ASAP7_75t_L g706 ( .A(n_636), .Y(n_706) );
CKINVDCx5p33_ASAP7_75t_R g638 ( .A(n_639), .Y(n_638) );
INVx4_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
INVx2_ASAP7_75t_L g646 ( .A(n_647), .Y(n_646) );
INVx2_ASAP7_75t_L g647 ( .A(n_648), .Y(n_647) );
INVx2_ASAP7_75t_L g649 ( .A(n_650), .Y(n_649) );
INVx1_ASAP7_75t_L g652 ( .A(n_653), .Y(n_652) );
INVx1_ASAP7_75t_L g653 ( .A(n_654), .Y(n_653) );
CKINVDCx20_ASAP7_75t_R g656 ( .A(n_657), .Y(n_656) );
CKINVDCx20_ASAP7_75t_R g657 ( .A(n_658), .Y(n_657) );
BUFx2_ASAP7_75t_L g658 ( .A(n_659), .Y(n_658) );
BUFx6f_ASAP7_75t_L g659 ( .A(n_660), .Y(n_659) );
NAND2xp5_ASAP7_75t_L g660 ( .A(n_661), .B(n_664), .Y(n_660) );
INVx1_ASAP7_75t_L g661 ( .A(n_662), .Y(n_661) );
BUFx2_ASAP7_75t_L g662 ( .A(n_663), .Y(n_662) );
INVx1_ASAP7_75t_L g691 ( .A(n_663), .Y(n_691) );
AND2x2_ASAP7_75t_L g723 ( .A(n_664), .B(n_724), .Y(n_723) );
INVx1_ASAP7_75t_L g664 ( .A(n_665), .Y(n_664) );
NAND2xp5_ASAP7_75t_L g690 ( .A(n_665), .B(n_691), .Y(n_690) );
AOI22xp33_ASAP7_75t_L g666 ( .A1(n_667), .A2(n_685), .B1(n_707), .B2(n_709), .Y(n_666) );
OAI22xp5_ASAP7_75t_L g716 ( .A1(n_667), .A2(n_707), .B1(n_717), .B2(n_719), .Y(n_716) );
XNOR2xp5_ASAP7_75t_L g667 ( .A(n_668), .B(n_676), .Y(n_667) );
INVx1_ASAP7_75t_L g670 ( .A(n_671), .Y(n_670) );
OAI22xp5_ASAP7_75t_L g671 ( .A1(n_672), .A2(n_673), .B1(n_674), .B2(n_675), .Y(n_671) );
INVx2_ASAP7_75t_L g672 ( .A(n_673), .Y(n_672) );
INVx1_ASAP7_75t_L g675 ( .A(n_674), .Y(n_675) );
AOI22xp5_ASAP7_75t_L g676 ( .A1(n_677), .A2(n_678), .B1(n_681), .B2(n_682), .Y(n_676) );
INVx1_ASAP7_75t_L g677 ( .A(n_678), .Y(n_677) );
INVx1_ASAP7_75t_L g681 ( .A(n_682), .Y(n_681) );
INVx1_ASAP7_75t_L g684 ( .A(n_683), .Y(n_684) );
INVx2_ASAP7_75t_L g685 ( .A(n_686), .Y(n_685) );
BUFx3_ASAP7_75t_L g686 ( .A(n_687), .Y(n_686) );
INVx1_ASAP7_75t_L g718 ( .A(n_687), .Y(n_718) );
INVx5_ASAP7_75t_L g687 ( .A(n_688), .Y(n_687) );
AND2x6_ASAP7_75t_L g688 ( .A(n_689), .B(n_699), .Y(n_688) );
NOR2xp33_ASAP7_75t_L g689 ( .A(n_690), .B(n_692), .Y(n_689) );
INVxp67_ASAP7_75t_L g713 ( .A(n_690), .Y(n_713) );
INVx1_ASAP7_75t_L g724 ( .A(n_691), .Y(n_724) );
INVxp67_ASAP7_75t_SL g692 ( .A(n_693), .Y(n_692) );
NAND2xp5_ASAP7_75t_L g714 ( .A(n_693), .B(n_703), .Y(n_714) );
NAND3xp33_ASAP7_75t_L g693 ( .A(n_694), .B(n_696), .C(n_697), .Y(n_693) );
INVx2_ASAP7_75t_L g694 ( .A(n_695), .Y(n_694) );
CKINVDCx11_ASAP7_75t_R g701 ( .A(n_695), .Y(n_701) );
AND2x4_ASAP7_75t_L g704 ( .A(n_696), .B(n_705), .Y(n_704) );
BUFx6f_ASAP7_75t_L g697 ( .A(n_698), .Y(n_697) );
NAND2xp5_ASAP7_75t_L g699 ( .A(n_700), .B(n_702), .Y(n_699) );
CKINVDCx5p33_ASAP7_75t_R g700 ( .A(n_701), .Y(n_700) );
INVx2_ASAP7_75t_SL g702 ( .A(n_703), .Y(n_702) );
INVx2_ASAP7_75t_SL g703 ( .A(n_704), .Y(n_703) );
INVx1_ASAP7_75t_L g705 ( .A(n_706), .Y(n_705) );
INVx1_ASAP7_75t_L g707 ( .A(n_708), .Y(n_707) );
INVx2_ASAP7_75t_L g709 ( .A(n_710), .Y(n_709) );
BUFx6f_ASAP7_75t_L g710 ( .A(n_711), .Y(n_710) );
BUFx6f_ASAP7_75t_L g719 ( .A(n_711), .Y(n_719) );
INVx4_ASAP7_75t_L g711 ( .A(n_712), .Y(n_711) );
AND2x2_ASAP7_75t_L g712 ( .A(n_713), .B(n_714), .Y(n_712) );
INVx1_ASAP7_75t_L g717 ( .A(n_718), .Y(n_717) );
CKINVDCx20_ASAP7_75t_R g720 ( .A(n_721), .Y(n_720) );
CKINVDCx20_ASAP7_75t_R g721 ( .A(n_722), .Y(n_721) );
endmodule