module real_aes_3763_n_360 (n_76, n_113, n_187, n_90, n_257, n_65, n_74, n_185, n_285, n_30, n_222, n_61, n_20, n_287, n_357, n_64, n_254, n_207, n_10, n_83, n_181, n_124, n_191, n_209, n_299, n_322, n_328, n_19, n_40, n_318, n_355, n_239, n_100, n_54, n_112, n_319, n_35, n_42, n_329, n_132, n_131, n_144, n_169, n_242, n_308, n_172, n_341, n_232, n_6, n_69, n_317, n_353, n_321, n_73, n_320, n_77, n_260, n_37, n_97, n_186, n_138, n_26, n_235, n_245, n_161, n_189, n_271, n_2, n_145, n_227, n_92, n_330, n_332, n_292, n_116, n_94, n_289, n_280, n_333, n_213, n_356, n_184, n_28, n_202, n_56, n_34, n_98, n_121, n_352, n_125, n_216, n_82, n_327, n_47, n_106, n_32, n_263, n_230, n_51, n_248, n_301, n_27, n_343, n_174, n_18, n_104, n_211, n_281, n_1210, n_173, n_234, n_284, n_153, n_316, n_75, n_178, n_298, n_49, n_43, n_297, n_9, n_119, n_310, n_164, n_231, n_44, n_102, n_122, n_141, n_128, n_111, n_167, n_80, n_179, n_12, n_68, n_129, n_345, n_304, n_311, n_324, n_25, n_278, n_236, n_267, n_218, n_48, n_204, n_339, n_89, n_277, n_331, n_93, n_182, n_323, n_199, n_350, n_142, n_223, n_67, n_250, n_85, n_45, n_5, n_244, n_118, n_139, n_87, n_171, n_78, n_146, n_17, n_226, n_255, n_286, n_120, n_261, n_238, n_58, n_165, n_246, n_176, n_163, n_29, n_52, n_251, n_220, n_197, n_296, n_3, n_41, n_256, n_71, n_302, n_351, n_126, n_200, n_115, n_96, n_110, n_150, n_147, n_288, n_23, n_334, n_274, n_160, n_303, n_95, n_188, n_269, n_201, n_306, n_158, n_4, n_346, n_193, n_293, n_162, n_358, n_275, n_214, n_46, n_109, n_59, n_203, n_81, n_133, n_273, n_114, n_276, n_295, n_265, n_354, n_154, n_127, n_326, n_24, n_217, n_55, n_62, n_291, n_148, n_88, n_159, n_11, n_108, n_60, n_233, n_290, n_155, n_243, n_268, n_136, n_157, n_282, n_101, n_309, n_344, n_229, n_107, n_33, n_53, n_36, n_149, n_190, n_262, n_134, n_349, n_336, n_195, n_300, n_252, n_283, n_314, n_249, n_221, n_156, n_359, n_57, n_66, n_21, n_31, n_8, n_312, n_183, n_266, n_205, n_335, n_177, n_313, n_22, n_140, n_219, n_180, n_212, n_210, n_325, n_338, n_103, n_166, n_224, n_151, n_130, n_253, n_99, n_15, n_72, n_152, n_198, n_7, n_228, n_272, n_196, n_347, n_315, n_123, n_279, n_79, n_270, n_305, n_117, n_208, n_215, n_135, n_70, n_50, n_170, n_86, n_340, n_13, n_168, n_175, n_241, n_105, n_84, n_294, n_258, n_206, n_307, n_342, n_348, n_14, n_194, n_137, n_225, n_16, n_39, n_337, n_247, n_240, n_38, n_259, n_143, n_192, n_0, n_264, n_63, n_1, n_237, n_91, n_360);
input n_76;
input n_113;
input n_187;
input n_90;
input n_257;
input n_65;
input n_74;
input n_185;
input n_285;
input n_30;
input n_222;
input n_61;
input n_20;
input n_287;
input n_357;
input n_64;
input n_254;
input n_207;
input n_10;
input n_83;
input n_181;
input n_124;
input n_191;
input n_209;
input n_299;
input n_322;
input n_328;
input n_19;
input n_40;
input n_318;
input n_355;
input n_239;
input n_100;
input n_54;
input n_112;
input n_319;
input n_35;
input n_42;
input n_329;
input n_132;
input n_131;
input n_144;
input n_169;
input n_242;
input n_308;
input n_172;
input n_341;
input n_232;
input n_6;
input n_69;
input n_317;
input n_353;
input n_321;
input n_73;
input n_320;
input n_77;
input n_260;
input n_37;
input n_97;
input n_186;
input n_138;
input n_26;
input n_235;
input n_245;
input n_161;
input n_189;
input n_271;
input n_2;
input n_145;
input n_227;
input n_92;
input n_330;
input n_332;
input n_292;
input n_116;
input n_94;
input n_289;
input n_280;
input n_333;
input n_213;
input n_356;
input n_184;
input n_28;
input n_202;
input n_56;
input n_34;
input n_98;
input n_121;
input n_352;
input n_125;
input n_216;
input n_82;
input n_327;
input n_47;
input n_106;
input n_32;
input n_263;
input n_230;
input n_51;
input n_248;
input n_301;
input n_27;
input n_343;
input n_174;
input n_18;
input n_104;
input n_211;
input n_281;
input n_1210;
input n_173;
input n_234;
input n_284;
input n_153;
input n_316;
input n_75;
input n_178;
input n_298;
input n_49;
input n_43;
input n_297;
input n_9;
input n_119;
input n_310;
input n_164;
input n_231;
input n_44;
input n_102;
input n_122;
input n_141;
input n_128;
input n_111;
input n_167;
input n_80;
input n_179;
input n_12;
input n_68;
input n_129;
input n_345;
input n_304;
input n_311;
input n_324;
input n_25;
input n_278;
input n_236;
input n_267;
input n_218;
input n_48;
input n_204;
input n_339;
input n_89;
input n_277;
input n_331;
input n_93;
input n_182;
input n_323;
input n_199;
input n_350;
input n_142;
input n_223;
input n_67;
input n_250;
input n_85;
input n_45;
input n_5;
input n_244;
input n_118;
input n_139;
input n_87;
input n_171;
input n_78;
input n_146;
input n_17;
input n_226;
input n_255;
input n_286;
input n_120;
input n_261;
input n_238;
input n_58;
input n_165;
input n_246;
input n_176;
input n_163;
input n_29;
input n_52;
input n_251;
input n_220;
input n_197;
input n_296;
input n_3;
input n_41;
input n_256;
input n_71;
input n_302;
input n_351;
input n_126;
input n_200;
input n_115;
input n_96;
input n_110;
input n_150;
input n_147;
input n_288;
input n_23;
input n_334;
input n_274;
input n_160;
input n_303;
input n_95;
input n_188;
input n_269;
input n_201;
input n_306;
input n_158;
input n_4;
input n_346;
input n_193;
input n_293;
input n_162;
input n_358;
input n_275;
input n_214;
input n_46;
input n_109;
input n_59;
input n_203;
input n_81;
input n_133;
input n_273;
input n_114;
input n_276;
input n_295;
input n_265;
input n_354;
input n_154;
input n_127;
input n_326;
input n_24;
input n_217;
input n_55;
input n_62;
input n_291;
input n_148;
input n_88;
input n_159;
input n_11;
input n_108;
input n_60;
input n_233;
input n_290;
input n_155;
input n_243;
input n_268;
input n_136;
input n_157;
input n_282;
input n_101;
input n_309;
input n_344;
input n_229;
input n_107;
input n_33;
input n_53;
input n_36;
input n_149;
input n_190;
input n_262;
input n_134;
input n_349;
input n_336;
input n_195;
input n_300;
input n_252;
input n_283;
input n_314;
input n_249;
input n_221;
input n_156;
input n_359;
input n_57;
input n_66;
input n_21;
input n_31;
input n_8;
input n_312;
input n_183;
input n_266;
input n_205;
input n_335;
input n_177;
input n_313;
input n_22;
input n_140;
input n_219;
input n_180;
input n_212;
input n_210;
input n_325;
input n_338;
input n_103;
input n_166;
input n_224;
input n_151;
input n_130;
input n_253;
input n_99;
input n_15;
input n_72;
input n_152;
input n_198;
input n_7;
input n_228;
input n_272;
input n_196;
input n_347;
input n_315;
input n_123;
input n_279;
input n_79;
input n_270;
input n_305;
input n_117;
input n_208;
input n_215;
input n_135;
input n_70;
input n_50;
input n_170;
input n_86;
input n_340;
input n_13;
input n_168;
input n_175;
input n_241;
input n_105;
input n_84;
input n_294;
input n_258;
input n_206;
input n_307;
input n_342;
input n_348;
input n_14;
input n_194;
input n_137;
input n_225;
input n_16;
input n_39;
input n_337;
input n_247;
input n_240;
input n_38;
input n_259;
input n_143;
input n_192;
input n_0;
input n_264;
input n_63;
input n_1;
input n_237;
input n_91;
output n_360;
wire n_480;
wire n_1177;
wire n_1073;
wire n_476;
wire n_758;
wire n_599;
wire n_436;
wire n_887;
wire n_684;
wire n_1066;
wire n_390;
wire n_1178;
wire n_1096;
wire n_821;
wire n_830;
wire n_624;
wire n_1018;
wire n_980;
wire n_800;
wire n_778;
wire n_618;
wire n_1175;
wire n_1106;
wire n_522;
wire n_1092;
wire n_838;
wire n_933;
wire n_1170;
wire n_485;
wire n_1205;
wire n_822;
wire n_846;
wire n_750;
wire n_631;
wire n_943;
wire n_977;
wire n_503;
wire n_792;
wire n_673;
wire n_386;
wire n_635;
wire n_518;
wire n_905;
wire n_1067;
wire n_878;
wire n_1192;
wire n_665;
wire n_667;
wire n_991;
wire n_1114;
wire n_580;
wire n_577;
wire n_1004;
wire n_469;
wire n_987;
wire n_362;
wire n_759;
wire n_979;
wire n_445;
wire n_1065;
wire n_596;
wire n_592;
wire n_540;
wire n_1064;
wire n_1075;
wire n_1197;
wire n_657;
wire n_900;
wire n_841;
wire n_718;
wire n_1129;
wire n_669;
wire n_1091;
wire n_423;
wire n_458;
wire n_1200;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_364;
wire n_421;
wire n_555;
wire n_766;
wire n_852;
wire n_1113;
wire n_974;
wire n_857;
wire n_919;
wire n_1089;
wire n_1122;
wire n_461;
wire n_1047;
wire n_1016;
wire n_908;
wire n_376;
wire n_571;
wire n_549;
wire n_694;
wire n_491;
wire n_894;
wire n_923;
wire n_1123;
wire n_1034;
wire n_952;
wire n_429;
wire n_1110;
wire n_752;
wire n_448;
wire n_545;
wire n_556;
wire n_1137;
wire n_593;
wire n_460;
wire n_937;
wire n_989;
wire n_773;
wire n_401;
wire n_538;
wire n_431;
wire n_1044;
wire n_963;
wire n_865;
wire n_537;
wire n_666;
wire n_551;
wire n_884;
wire n_560;
wire n_660;
wire n_1094;
wire n_814;
wire n_944;
wire n_886;
wire n_856;
wire n_594;
wire n_1146;
wire n_983;
wire n_767;
wire n_889;
wire n_696;
wire n_955;
wire n_1147;
wire n_975;
wire n_704;
wire n_941;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_932;
wire n_948;
wire n_399;
wire n_700;
wire n_1021;
wire n_677;
wire n_958;
wire n_1046;
wire n_378;
wire n_591;
wire n_775;
wire n_763;
wire n_1093;
wire n_1109;
wire n_870;
wire n_961;
wire n_489;
wire n_427;
wire n_678;
wire n_548;
wire n_415;
wire n_572;
wire n_564;
wire n_519;
wire n_638;
wire n_815;
wire n_1116;
wire n_573;
wire n_510;
wire n_1140;
wire n_1099;
wire n_709;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_816;
wire n_539;
wire n_400;
wire n_626;
wire n_625;
wire n_953;
wire n_462;
wire n_615;
wire n_1118;
wire n_990;
wire n_550;
wire n_966;
wire n_1160;
wire n_1108;
wire n_670;
wire n_818;
wire n_716;
wire n_883;
wire n_478;
wire n_918;
wire n_584;
wire n_896;
wire n_408;
wire n_553;
wire n_892;
wire n_578;
wire n_528;
wire n_372;
wire n_495;
wire n_994;
wire n_1078;
wire n_370;
wire n_1072;
wire n_744;
wire n_384;
wire n_938;
wire n_1128;
wire n_935;
wire n_824;
wire n_1098;
wire n_1199;
wire n_467;
wire n_875;
wire n_951;
wire n_774;
wire n_992;
wire n_813;
wire n_791;
wire n_981;
wire n_976;
wire n_466;
wire n_1182;
wire n_636;
wire n_559;
wire n_872;
wire n_906;
wire n_477;
wire n_515;
wire n_984;
wire n_1019;
wire n_680;
wire n_595;
wire n_1086;
wire n_369;
wire n_1189;
wire n_726;
wire n_1070;
wire n_1180;
wire n_517;
wire n_683;
wire n_780;
wire n_904;
wire n_840;
wire n_570;
wire n_675;
wire n_931;
wire n_920;
wire n_530;
wire n_835;
wire n_535;
wire n_732;
wire n_1117;
wire n_834;
wire n_882;
wire n_784;
wire n_962;
wire n_496;
wire n_693;
wire n_1082;
wire n_468;
wire n_746;
wire n_532;
wire n_656;
wire n_755;
wire n_1025;
wire n_1168;
wire n_1148;
wire n_409;
wire n_748;
wire n_781;
wire n_909;
wire n_523;
wire n_860;
wire n_996;
wire n_439;
wire n_1062;
wire n_576;
wire n_924;
wire n_956;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_1049;
wire n_874;
wire n_796;
wire n_1152;
wire n_801;
wire n_1126;
wire n_383;
wire n_529;
wire n_1115;
wire n_504;
wire n_455;
wire n_725;
wire n_973;
wire n_671;
wire n_960;
wire n_1081;
wire n_1084;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_903;
wire n_454;
wire n_1198;
wire n_817;
wire n_565;
wire n_443;
wire n_782;
wire n_760;
wire n_608;
wire n_812;
wire n_534;
wire n_925;
wire n_708;
wire n_1029;
wire n_1020;
wire n_457;
wire n_885;
wire n_1121;
wire n_1207;
wire n_1059;
wire n_950;
wire n_381;
wire n_993;
wire n_493;
wire n_664;
wire n_367;
wire n_819;
wire n_1196;
wire n_737;
wire n_1013;
wire n_1017;
wire n_581;
wire n_610;
wire n_936;
wire n_1035;
wire n_620;
wire n_582;
wire n_641;
wire n_1063;
wire n_1135;
wire n_828;
wire n_808;
wire n_770;
wire n_940;
wire n_745;
wire n_867;
wire n_722;
wire n_398;
wire n_1100;
wire n_1167;
wire n_1174;
wire n_688;
wire n_1193;
wire n_425;
wire n_609;
wire n_1042;
wire n_879;
wire n_417;
wire n_363;
wire n_449;
wire n_607;
wire n_754;
wire n_1006;
wire n_690;
wire n_629;
wire n_1053;
wire n_499;
wire n_508;
wire n_1142;
wire n_1141;
wire n_706;
wire n_901;
wire n_561;
wire n_970;
wire n_947;
wire n_876;
wire n_437;
wire n_1112;
wire n_428;
wire n_405;
wire n_1149;
wire n_621;
wire n_368;
wire n_783;
wire n_1107;
wire n_1012;
wire n_655;
wire n_654;
wire n_502;
wire n_505;
wire n_769;
wire n_527;
wire n_434;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_1054;
wire n_672;
wire n_567;
wire n_916;
wire n_406;
wire n_1050;
wire n_426;
wire n_1134;
wire n_733;
wire n_552;
wire n_602;
wire n_402;
wire n_617;
wire n_658;
wire n_676;
wire n_986;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_880;
wire n_1031;
wire n_1037;
wire n_1103;
wire n_1131;
wire n_1008;
wire n_807;
wire n_1011;
wire n_416;
wire n_790;
wire n_895;
wire n_832;
wire n_410;
wire n_799;
wire n_805;
wire n_751;
wire n_999;
wire n_490;
wire n_913;
wire n_619;
wire n_391;
wire n_1095;
wire n_1060;
wire n_859;
wire n_695;
wire n_1181;
wire n_685;
wire n_881;
wire n_1154;
wire n_1080;
wire n_361;
wire n_917;
wire n_632;
wire n_768;
wire n_412;
wire n_542;
wire n_645;
wire n_1145;
wire n_557;
wire n_714;
wire n_777;
wire n_985;
wire n_1077;
wire n_501;
wire n_488;
wire n_1041;
wire n_1111;
wire n_910;
wire n_642;
wire n_613;
wire n_869;
wire n_387;
wire n_1125;
wire n_957;
wire n_995;
wire n_1124;
wire n_702;
wire n_954;
wire n_969;
wire n_912;
wire n_1009;
wire n_1202;
wire n_1007;
wire n_464;
wire n_1163;
wire n_945;
wire n_604;
wire n_734;
wire n_898;
wire n_848;
wire n_392;
wire n_562;
wire n_1022;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_756;
wire n_1201;
wire n_1179;
wire n_569;
wire n_997;
wire n_785;
wire n_1203;
wire n_563;
wire n_1171;
wire n_891;
wire n_430;
wire n_568;
wire n_413;
wire n_471;
wire n_902;
wire n_1105;
wire n_1157;
wire n_1158;
wire n_1132;
wire n_853;
wire n_810;
wire n_843;
wire n_1079;
wire n_579;
wire n_1033;
wire n_699;
wire n_533;
wire n_1028;
wire n_1003;
wire n_1000;
wire n_1014;
wire n_1187;
wire n_366;
wire n_727;
wire n_1083;
wire n_649;
wire n_385;
wire n_397;
wire n_749;
wire n_663;
wire n_588;
wire n_536;
wire n_914;
wire n_707;
wire n_622;
wire n_470;
wire n_851;
wire n_915;
wire n_1002;
wire n_1155;
wire n_934;
wire n_1165;
wire n_494;
wire n_1001;
wire n_711;
wire n_864;
wire n_1027;
wire n_1169;
wire n_377;
wire n_1058;
wire n_1139;
wire n_927;
wire n_1038;
wire n_965;
wire n_723;
wire n_662;
wire n_1085;
wire n_382;
wire n_845;
wire n_850;
wire n_1043;
wire n_1136;
wire n_720;
wire n_972;
wire n_1127;
wire n_435;
wire n_968;
wire n_1026;
wire n_511;
wire n_484;
wire n_893;
wire n_492;
wire n_1068;
wire n_509;
wire n_407;
wire n_419;
wire n_730;
wire n_1023;
wire n_643;
wire n_747;
wire n_1204;
wire n_486;
wire n_930;
wire n_1057;
wire n_411;
wire n_697;
wire n_978;
wire n_847;
wire n_907;
wire n_779;
wire n_498;
wire n_481;
wire n_765;
wire n_691;
wire n_826;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_939;
wire n_1005;
wire n_487;
wire n_831;
wire n_653;
wire n_365;
wire n_526;
wire n_637;
wire n_899;
wire n_928;
wire n_692;
wire n_789;
wire n_544;
wire n_1087;
wire n_1051;
wire n_1194;
wire n_389;
wire n_738;
wire n_701;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_926;
wire n_922;
wire n_942;
wire n_1048;
wire n_472;
wire n_1120;
wire n_971;
wire n_866;
wire n_452;
wire n_787;
wire n_1071;
wire n_1052;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_1097;
wire n_715;
wire n_959;
wire n_1208;
wire n_946;
wire n_420;
wire n_612;
wire n_858;
wire n_873;
wire n_1130;
wire n_438;
wire n_764;
wire n_794;
wire n_741;
wire n_753;
wire n_1188;
wire n_623;
wire n_1032;
wire n_446;
wire n_721;
wire n_681;
wire n_1090;
wire n_456;
wire n_717;
wire n_982;
wire n_1133;
wire n_1164;
wire n_712;
wire n_1183;
wire n_433;
wire n_516;
wire n_627;
wire n_739;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_524;
wire n_861;
wire n_1162;
wire n_705;
wire n_1191;
wire n_1206;
wire n_1195;
wire n_575;
wire n_762;
wire n_479;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_541;
wire n_839;
wire n_546;
wire n_587;
wire n_639;
wire n_1186;
wire n_1010;
wire n_811;
wire n_1015;
wire n_459;
wire n_558;
wire n_1172;
wire n_863;
wire n_998;
wire n_724;
wire n_440;
wire n_525;
wire n_1074;
wire n_644;
wire n_674;
wire n_836;
wire n_888;
wire n_793;
wire n_1150;
wire n_1184;
wire n_1166;
wire n_1056;
wire n_583;
wire n_833;
wire n_414;
wire n_757;
wire n_1161;
wire n_929;
wire n_1143;
wire n_686;
wire n_776;
wire n_1190;
wire n_1138;
wire n_803;
wire n_890;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_949;
wire n_614;
wire n_586;
wire n_911;
wire n_772;
wire n_450;
wire n_788;
wire n_441;
wire n_585;
wire n_465;
wire n_719;
wire n_473;
wire n_566;
wire n_967;
wire n_837;
wire n_1045;
wire n_871;
wire n_474;
wire n_1159;
wire n_1156;
wire n_829;
wire n_1030;
wire n_988;
wire n_1088;
wire n_1055;
wire n_921;
wire n_375;
wire n_597;
wire n_640;
wire n_483;
wire n_611;
wire n_1176;
wire n_1151;
wire n_380;
wire n_1036;
wire n_394;
wire n_687;
wire n_729;
wire n_844;
wire n_646;
wire n_650;
wire n_710;
wire n_743;
wire n_823;
wire n_393;
wire n_652;
wire n_703;
wire n_1040;
wire n_500;
wire n_601;
wire n_1102;
wire n_661;
wire n_463;
wire n_1076;
wire n_396;
wire n_804;
wire n_1101;
wire n_447;
wire n_1185;
wire n_1173;
wire n_603;
wire n_403;
wire n_854;
wire n_424;
wire n_877;
wire n_802;
wire n_868;
wire n_1119;
wire n_1039;
wire n_574;
wire n_1069;
wire n_1024;
wire n_842;
wire n_1104;
wire n_1144;
wire n_849;
wire n_1061;
wire n_475;
wire n_554;
wire n_897;
wire n_1153;
wire n_855;
wire n_798;
wire n_797;
wire n_668;
wire n_862;
AOI22xp33_ASAP7_75t_L g836 ( .A1(n_0), .A2(n_102), .B1(n_582), .B2(n_733), .Y(n_836) );
AOI22x1_ASAP7_75t_L g774 ( .A1(n_1), .A2(n_216), .B1(n_429), .B2(n_731), .Y(n_774) );
AOI22xp33_ASAP7_75t_L g506 ( .A1(n_2), .A2(n_132), .B1(n_507), .B2(n_508), .Y(n_506) );
AOI22xp33_ASAP7_75t_L g885 ( .A1(n_3), .A2(n_221), .B1(n_501), .B2(n_502), .Y(n_885) );
AOI22xp33_ASAP7_75t_L g923 ( .A1(n_4), .A2(n_321), .B1(n_620), .B2(n_924), .Y(n_923) );
AOI22xp33_ASAP7_75t_L g544 ( .A1(n_5), .A2(n_273), .B1(n_545), .B2(n_546), .Y(n_544) );
AOI22xp33_ASAP7_75t_L g585 ( .A1(n_6), .A2(n_173), .B1(n_433), .B2(n_586), .Y(n_585) );
CKINVDCx5p33_ASAP7_75t_R g722 ( .A(n_7), .Y(n_722) );
INVx1_ASAP7_75t_L g865 ( .A(n_8), .Y(n_865) );
AOI221xp5_ASAP7_75t_L g651 ( .A1(n_9), .A2(n_285), .B1(n_619), .B2(n_652), .C(n_653), .Y(n_651) );
AOI22xp33_ASAP7_75t_L g513 ( .A1(n_10), .A2(n_301), .B1(n_486), .B2(n_488), .Y(n_513) );
AOI22xp5_ASAP7_75t_L g790 ( .A1(n_11), .A2(n_293), .B1(n_727), .B2(n_777), .Y(n_790) );
AOI22xp5_ASAP7_75t_L g920 ( .A1(n_12), .A2(n_82), .B1(n_867), .B2(n_921), .Y(n_920) );
AOI22xp33_ASAP7_75t_L g730 ( .A1(n_13), .A2(n_202), .B1(n_731), .B2(n_732), .Y(n_730) );
AOI22xp33_ASAP7_75t_L g500 ( .A1(n_14), .A2(n_186), .B1(n_501), .B2(n_502), .Y(n_500) );
NAND2xp5_ASAP7_75t_SL g399 ( .A(n_15), .B(n_388), .Y(n_399) );
AOI22xp5_ASAP7_75t_L g1200 ( .A1(n_16), .A2(n_1201), .B1(n_1202), .B2(n_1203), .Y(n_1200) );
CKINVDCx20_ASAP7_75t_R g1203 ( .A(n_16), .Y(n_1203) );
AOI22xp5_ASAP7_75t_L g961 ( .A1(n_17), .A2(n_334), .B1(n_962), .B2(n_966), .Y(n_961) );
AOI22xp33_ASAP7_75t_L g657 ( .A1(n_18), .A2(n_267), .B1(n_475), .B2(n_658), .Y(n_657) );
AOI22xp33_ASAP7_75t_L g432 ( .A1(n_19), .A2(n_93), .B1(n_433), .B2(n_437), .Y(n_432) );
AOI22xp33_ASAP7_75t_L g853 ( .A1(n_20), .A2(n_30), .B1(n_406), .B2(n_580), .Y(n_853) );
BUFx6f_ASAP7_75t_L g388 ( .A(n_21), .Y(n_388) );
AOI22xp5_ASAP7_75t_L g928 ( .A1(n_22), .A2(n_332), .B1(n_383), .B2(n_643), .Y(n_928) );
AOI22xp33_ASAP7_75t_L g693 ( .A1(n_23), .A2(n_32), .B1(n_504), .B2(n_507), .Y(n_693) );
INVx1_ASAP7_75t_L g944 ( .A(n_24), .Y(n_944) );
AOI22xp33_ASAP7_75t_L g522 ( .A1(n_25), .A2(n_71), .B1(n_505), .B2(n_508), .Y(n_522) );
AOI22xp33_ASAP7_75t_L g674 ( .A1(n_26), .A2(n_217), .B1(n_489), .B2(n_498), .Y(n_674) );
NAND2xp5_ASAP7_75t_L g696 ( .A(n_27), .B(n_552), .Y(n_696) );
AOI22xp5_ASAP7_75t_L g426 ( .A1(n_28), .A2(n_151), .B1(n_427), .B2(n_429), .Y(n_426) );
AOI22xp33_ASAP7_75t_L g648 ( .A1(n_29), .A2(n_168), .B1(n_437), .B2(n_649), .Y(n_648) );
AOI221xp5_ASAP7_75t_L g891 ( .A1(n_31), .A2(n_338), .B1(n_486), .B2(n_488), .C(n_892), .Y(n_891) );
AOI21xp33_ASAP7_75t_L g1187 ( .A1(n_33), .A2(n_552), .B(n_1188), .Y(n_1187) );
AOI21xp5_ASAP7_75t_L g622 ( .A1(n_34), .A2(n_623), .B(n_625), .Y(n_622) );
AOI22xp33_ASAP7_75t_L g795 ( .A1(n_35), .A2(n_180), .B1(n_591), .B2(n_658), .Y(n_795) );
INVx1_ASAP7_75t_L g495 ( .A(n_36), .Y(n_495) );
AOI22xp33_ASAP7_75t_L g937 ( .A1(n_37), .A2(n_103), .B1(n_580), .B2(n_678), .Y(n_937) );
AOI22xp33_ASAP7_75t_L g950 ( .A1(n_38), .A2(n_45), .B1(n_565), .B2(n_658), .Y(n_950) );
AOI22xp33_ASAP7_75t_L g845 ( .A1(n_39), .A2(n_201), .B1(n_658), .B2(n_846), .Y(n_845) );
AOI22xp33_ASAP7_75t_L g701 ( .A1(n_40), .A2(n_98), .B1(n_489), .B2(n_702), .Y(n_701) );
AOI22xp5_ASAP7_75t_L g1192 ( .A1(n_41), .A2(n_335), .B1(n_547), .B2(n_669), .Y(n_1192) );
AOI22xp33_ASAP7_75t_L g820 ( .A1(n_42), .A2(n_341), .B1(n_499), .B2(n_505), .Y(n_820) );
AOI22xp33_ASAP7_75t_L g382 ( .A1(n_43), .A2(n_128), .B1(n_383), .B2(n_406), .Y(n_382) );
AO22x1_ASAP7_75t_L g892 ( .A1(n_44), .A2(n_65), .B1(n_489), .B2(n_493), .Y(n_892) );
AOI22xp33_ASAP7_75t_L g813 ( .A1(n_46), .A2(n_289), .B1(n_488), .B2(n_489), .Y(n_813) );
NAND2xp5_ASAP7_75t_L g557 ( .A(n_47), .B(n_558), .Y(n_557) );
OA22x2_ASAP7_75t_L g393 ( .A1(n_48), .A2(n_140), .B1(n_388), .B2(n_392), .Y(n_393) );
INVx1_ASAP7_75t_L g412 ( .A(n_48), .Y(n_412) );
AOI22xp33_ASAP7_75t_L g581 ( .A1(n_49), .A2(n_117), .B1(n_429), .B2(n_582), .Y(n_581) );
AOI221xp5_ASAP7_75t_L g442 ( .A1(n_50), .A2(n_62), .B1(n_443), .B2(n_447), .C(n_450), .Y(n_442) );
AOI22xp33_ASAP7_75t_L g1092 ( .A1(n_51), .A2(n_192), .B1(n_989), .B2(n_1002), .Y(n_1092) );
AOI22xp33_ASAP7_75t_L g930 ( .A1(n_52), .A2(n_295), .B1(n_437), .B2(n_649), .Y(n_930) );
AOI221x1_ASAP7_75t_L g787 ( .A1(n_53), .A2(n_253), .B1(n_677), .B2(n_687), .C(n_788), .Y(n_787) );
INVxp67_ASAP7_75t_L g850 ( .A(n_54), .Y(n_850) );
AOI22xp33_ASAP7_75t_L g1011 ( .A1(n_54), .A2(n_171), .B1(n_969), .B2(n_972), .Y(n_1011) );
AOI22xp33_ASAP7_75t_L g857 ( .A1(n_55), .A2(n_131), .B1(n_433), .B2(n_586), .Y(n_857) );
AOI221xp5_ASAP7_75t_L g771 ( .A1(n_56), .A2(n_240), .B1(n_737), .B2(n_772), .C(n_773), .Y(n_771) );
AOI22xp33_ASAP7_75t_L g594 ( .A1(n_57), .A2(n_277), .B1(n_465), .B2(n_568), .Y(n_594) );
AOI22xp33_ASAP7_75t_L g854 ( .A1(n_58), .A2(n_353), .B1(n_383), .B2(n_427), .Y(n_854) );
AOI22xp33_ASAP7_75t_L g743 ( .A1(n_59), .A2(n_329), .B1(n_744), .B2(n_745), .Y(n_743) );
AOI22xp33_ASAP7_75t_L g487 ( .A1(n_60), .A2(n_323), .B1(n_488), .B2(n_489), .Y(n_487) );
NOR2xp33_ASAP7_75t_L g369 ( .A(n_61), .B(n_161), .Y(n_369) );
INVx1_ASAP7_75t_L g391 ( .A(n_61), .Y(n_391) );
OAI21xp33_ASAP7_75t_L g413 ( .A1(n_61), .A2(n_140), .B(n_414), .Y(n_413) );
INVx1_ASAP7_75t_L g809 ( .A(n_63), .Y(n_809) );
AO221x2_ASAP7_75t_L g987 ( .A1(n_63), .A2(n_336), .B1(n_969), .B2(n_976), .C(n_988), .Y(n_987) );
AOI22xp33_ASAP7_75t_L g901 ( .A1(n_64), .A2(n_166), .B1(n_462), .B2(n_902), .Y(n_901) );
AOI22xp33_ASAP7_75t_L g929 ( .A1(n_66), .A2(n_100), .B1(n_417), .B2(n_424), .Y(n_929) );
AOI22xp33_ASAP7_75t_L g560 ( .A1(n_67), .A2(n_153), .B1(n_561), .B2(n_562), .Y(n_560) );
INVx1_ASAP7_75t_L g608 ( .A(n_68), .Y(n_608) );
AOI22xp33_ASAP7_75t_L g886 ( .A1(n_69), .A2(n_197), .B1(n_485), .B2(n_504), .Y(n_886) );
AOI22xp33_ASAP7_75t_L g691 ( .A1(n_70), .A2(n_223), .B1(n_485), .B2(n_508), .Y(n_691) );
NOR3xp33_ASAP7_75t_L g784 ( .A(n_72), .B(n_785), .C(n_789), .Y(n_784) );
AOI22xp5_ASAP7_75t_L g805 ( .A1(n_72), .A2(n_789), .B1(n_794), .B2(n_1210), .Y(n_805) );
OAI21xp5_ASAP7_75t_L g806 ( .A1(n_72), .A2(n_785), .B(n_800), .Y(n_806) );
AOI22xp5_ASAP7_75t_L g982 ( .A1(n_72), .A2(n_326), .B1(n_972), .B2(n_983), .Y(n_982) );
AOI22xp33_ASAP7_75t_L g694 ( .A1(n_73), .A2(n_147), .B1(n_501), .B2(n_502), .Y(n_694) );
AOI21xp33_ASAP7_75t_L g698 ( .A1(n_74), .A2(n_498), .B(n_699), .Y(n_698) );
AOI22xp33_ASAP7_75t_L g936 ( .A1(n_75), .A2(n_78), .B1(n_427), .B2(n_539), .Y(n_936) );
AOI22xp33_ASAP7_75t_L g1001 ( .A1(n_76), .A2(n_339), .B1(n_962), .B2(n_1002), .Y(n_1001) );
AND2x4_ASAP7_75t_L g965 ( .A(n_77), .B(n_265), .Y(n_965) );
INVx1_ASAP7_75t_L g971 ( .A(n_77), .Y(n_971) );
AOI22xp33_ASAP7_75t_L g839 ( .A1(n_79), .A2(n_92), .B1(n_477), .B2(n_600), .Y(n_839) );
AOI22xp33_ASAP7_75t_L g692 ( .A1(n_80), .A2(n_86), .B1(n_499), .B2(n_505), .Y(n_692) );
AO22x1_ASAP7_75t_L g988 ( .A1(n_81), .A2(n_170), .B1(n_966), .B2(n_989), .Y(n_988) );
AOI22xp33_ASAP7_75t_L g618 ( .A1(n_83), .A2(n_224), .B1(n_619), .B2(n_620), .Y(n_618) );
AOI21xp33_ASAP7_75t_L g492 ( .A1(n_84), .A2(n_493), .B(n_494), .Y(n_492) );
AOI21xp5_ASAP7_75t_L g590 ( .A1(n_85), .A2(n_591), .B(n_592), .Y(n_590) );
XNOR2x2_ASAP7_75t_L g933 ( .A(n_87), .B(n_934), .Y(n_933) );
AOI211xp5_ASAP7_75t_L g762 ( .A1(n_88), .A2(n_763), .B(n_765), .C(n_769), .Y(n_762) );
AOI22xp5_ASAP7_75t_L g985 ( .A1(n_89), .A2(n_122), .B1(n_978), .B2(n_986), .Y(n_985) );
XNOR2x1_ASAP7_75t_L g510 ( .A(n_90), .B(n_511), .Y(n_510) );
AOI22xp33_ASAP7_75t_L g821 ( .A1(n_91), .A2(n_107), .B1(n_504), .B2(n_507), .Y(n_821) );
AOI22xp5_ASAP7_75t_L g766 ( .A1(n_94), .A2(n_176), .B1(n_443), .B2(n_477), .Y(n_766) );
AOI22xp33_ASAP7_75t_L g834 ( .A1(n_95), .A2(n_138), .B1(n_433), .B2(n_835), .Y(n_834) );
AOI22xp5_ASAP7_75t_L g672 ( .A1(n_96), .A2(n_142), .B1(n_488), .B2(n_673), .Y(n_672) );
AOI22xp33_ASAP7_75t_L g734 ( .A1(n_97), .A2(n_218), .B1(n_538), .B2(n_584), .Y(n_734) );
INVx1_ASAP7_75t_L g817 ( .A(n_99), .Y(n_817) );
AOI22xp5_ASAP7_75t_L g611 ( .A1(n_101), .A2(n_247), .B1(n_433), .B2(n_586), .Y(n_611) );
INVx1_ASAP7_75t_L g964 ( .A(n_104), .Y(n_964) );
AND2x4_ASAP7_75t_L g967 ( .A(n_104), .B(n_365), .Y(n_967) );
INVx1_ASAP7_75t_SL g984 ( .A(n_104), .Y(n_984) );
AOI22xp33_ASAP7_75t_L g686 ( .A1(n_105), .A2(n_350), .B1(n_437), .B2(n_687), .Y(n_686) );
AOI22xp33_ASAP7_75t_L g416 ( .A1(n_106), .A2(n_109), .B1(n_417), .B2(n_424), .Y(n_416) );
AOI22xp33_ASAP7_75t_L g524 ( .A1(n_108), .A2(n_264), .B1(n_499), .B2(n_507), .Y(n_524) );
AOI22xp33_ASAP7_75t_L g1010 ( .A1(n_110), .A2(n_137), .B1(n_962), .B2(n_966), .Y(n_1010) );
AOI22xp33_ASAP7_75t_L g720 ( .A1(n_111), .A2(n_258), .B1(n_558), .B2(n_658), .Y(n_720) );
XNOR2x1_ASAP7_75t_L g481 ( .A(n_112), .B(n_482), .Y(n_481) );
AOI22xp33_ASAP7_75t_L g697 ( .A1(n_113), .A2(n_291), .B1(n_486), .B2(n_488), .Y(n_697) );
NAND2xp5_ASAP7_75t_L g1184 ( .A(n_114), .B(n_619), .Y(n_1184) );
AOI22xp33_ASAP7_75t_L g668 ( .A1(n_115), .A2(n_219), .B1(n_669), .B2(n_670), .Y(n_668) );
AOI22xp5_ASAP7_75t_L g599 ( .A1(n_116), .A2(n_271), .B1(n_477), .B2(n_600), .Y(n_599) );
AOI22xp33_ASAP7_75t_L g503 ( .A1(n_118), .A2(n_152), .B1(n_504), .B2(n_505), .Y(n_503) );
AOI22xp33_ASAP7_75t_L g615 ( .A1(n_119), .A2(n_146), .B1(n_383), .B2(n_427), .Y(n_615) );
AOI22xp33_ASAP7_75t_L g617 ( .A1(n_120), .A2(n_302), .B1(n_475), .B2(n_568), .Y(n_617) );
AOI22xp33_ASAP7_75t_L g540 ( .A1(n_121), .A2(n_337), .B1(n_541), .B2(n_543), .Y(n_540) );
INVx1_ASAP7_75t_L g554 ( .A(n_123), .Y(n_554) );
NAND2xp5_ASAP7_75t_L g490 ( .A(n_124), .B(n_491), .Y(n_490) );
NAND2xp33_ASAP7_75t_L g786 ( .A(n_125), .B(n_678), .Y(n_786) );
AOI22xp33_ASAP7_75t_L g862 ( .A1(n_126), .A2(n_348), .B1(n_477), .B2(n_619), .Y(n_862) );
AOI22xp5_ASAP7_75t_L g583 ( .A1(n_127), .A2(n_345), .B1(n_383), .B2(n_584), .Y(n_583) );
AOI22xp5_ASAP7_75t_L g671 ( .A1(n_129), .A2(n_155), .B1(n_417), .B2(n_647), .Y(n_671) );
AOI22xp5_ASAP7_75t_L g530 ( .A1(n_130), .A2(n_215), .B1(n_531), .B2(n_534), .Y(n_530) );
INVx1_ASAP7_75t_L g700 ( .A(n_133), .Y(n_700) );
INVx1_ASAP7_75t_L g626 ( .A(n_134), .Y(n_626) );
AOI22xp33_ASAP7_75t_L g645 ( .A1(n_135), .A2(n_254), .B1(n_383), .B2(n_427), .Y(n_645) );
AO22x1_ASAP7_75t_L g779 ( .A1(n_136), .A2(n_214), .B1(n_584), .B2(n_780), .Y(n_779) );
INVx1_ASAP7_75t_L g405 ( .A(n_139), .Y(n_405) );
NAND2xp5_ASAP7_75t_L g460 ( .A(n_139), .B(n_410), .Y(n_460) );
NAND2xp5_ASAP7_75t_L g470 ( .A(n_139), .B(n_198), .Y(n_470) );
NOR2xp33_ASAP7_75t_L g368 ( .A(n_140), .B(n_281), .Y(n_368) );
AOI22xp33_ASAP7_75t_L g1089 ( .A1(n_141), .A2(n_208), .B1(n_999), .B2(n_1090), .Y(n_1089) );
AND2x2_ASAP7_75t_L g788 ( .A(n_143), .B(n_537), .Y(n_788) );
AOI22xp33_ASAP7_75t_SL g814 ( .A1(n_144), .A2(n_287), .B1(n_486), .B2(n_498), .Y(n_814) );
AOI22xp33_ASAP7_75t_L g461 ( .A1(n_145), .A2(n_150), .B1(n_462), .B2(n_465), .Y(n_461) );
AOI21xp33_ASAP7_75t_L g942 ( .A1(n_148), .A2(n_491), .B(n_943), .Y(n_942) );
XNOR2x1_ASAP7_75t_L g665 ( .A(n_149), .B(n_666), .Y(n_665) );
AOI22xp33_ASAP7_75t_L g840 ( .A1(n_154), .A2(n_268), .B1(n_462), .B2(n_841), .Y(n_840) );
NAND2xp5_ASAP7_75t_L g906 ( .A(n_156), .B(n_447), .Y(n_906) );
AO22x1_ASAP7_75t_L g769 ( .A1(n_157), .A2(n_299), .B1(n_580), .B2(n_770), .Y(n_769) );
AOI22xp33_ASAP7_75t_L g474 ( .A1(n_158), .A2(n_358), .B1(n_475), .B2(n_477), .Y(n_474) );
NAND2xp5_ASAP7_75t_L g629 ( .A(n_159), .B(n_558), .Y(n_629) );
AOI22xp5_ASAP7_75t_L g946 ( .A1(n_160), .A2(n_189), .B1(n_437), .B2(n_687), .Y(n_946) );
NAND2xp5_ASAP7_75t_L g397 ( .A(n_161), .B(n_398), .Y(n_397) );
AOI22xp33_ASAP7_75t_SL g1194 ( .A1(n_162), .A2(n_327), .B1(n_687), .B2(n_802), .Y(n_1194) );
AOI22xp5_ASAP7_75t_L g1193 ( .A1(n_163), .A2(n_331), .B1(n_677), .B2(n_948), .Y(n_1193) );
NAND2xp5_ASAP7_75t_L g595 ( .A(n_164), .B(n_596), .Y(n_595) );
AOI22xp5_ASAP7_75t_L g1191 ( .A1(n_165), .A2(n_297), .B1(n_539), .B2(n_678), .Y(n_1191) );
AOI22xp33_ASAP7_75t_L g855 ( .A1(n_167), .A2(n_190), .B1(n_582), .B2(n_856), .Y(n_855) );
INVx1_ASAP7_75t_L g939 ( .A(n_169), .Y(n_939) );
AOI22xp33_ASAP7_75t_L g676 ( .A1(n_172), .A2(n_262), .B1(n_677), .B2(n_678), .Y(n_676) );
AOI22xp33_ASAP7_75t_L g646 ( .A1(n_174), .A2(n_310), .B1(n_417), .B2(n_647), .Y(n_646) );
AOI22xp33_ASAP7_75t_L g925 ( .A1(n_175), .A2(n_250), .B1(n_902), .B2(n_926), .Y(n_925) );
AOI22xp33_ASAP7_75t_L g903 ( .A1(n_177), .A2(n_355), .B1(n_427), .B2(n_904), .Y(n_903) );
AOI22xp5_ASAP7_75t_L g910 ( .A1(n_178), .A2(n_229), .B1(n_516), .B2(n_911), .Y(n_910) );
INVx1_ASAP7_75t_L g703 ( .A(n_179), .Y(n_703) );
OA22x2_ASAP7_75t_L g881 ( .A1(n_181), .A2(n_882), .B1(n_893), .B2(n_894), .Y(n_881) );
INVx1_ASAP7_75t_L g894 ( .A(n_181), .Y(n_894) );
AOI221xp5_ASAP7_75t_L g775 ( .A1(n_182), .A2(n_191), .B1(n_776), .B2(n_778), .C(n_779), .Y(n_775) );
AOI21xp33_ASAP7_75t_SL g907 ( .A1(n_183), .A2(n_475), .B(n_908), .Y(n_907) );
AOI21xp5_ASAP7_75t_L g517 ( .A1(n_184), .A2(n_493), .B(n_518), .Y(n_517) );
AOI22xp33_ASAP7_75t_L g1185 ( .A1(n_185), .A2(n_356), .B1(n_902), .B2(n_926), .Y(n_1185) );
AOI22xp33_ASAP7_75t_L g535 ( .A1(n_187), .A2(n_245), .B1(n_536), .B2(n_538), .Y(n_535) );
AOI21xp33_ASAP7_75t_L g815 ( .A1(n_188), .A2(n_702), .B(n_816), .Y(n_815) );
INVx1_ASAP7_75t_L g917 ( .A(n_193), .Y(n_917) );
AOI22xp33_ASAP7_75t_L g525 ( .A1(n_194), .A2(n_342), .B1(n_501), .B2(n_502), .Y(n_525) );
AOI22xp5_ASAP7_75t_L g975 ( .A1(n_195), .A2(n_225), .B1(n_969), .B2(n_976), .Y(n_975) );
INVx1_ASAP7_75t_L g519 ( .A(n_196), .Y(n_519) );
INVx1_ASAP7_75t_L g389 ( .A(n_198), .Y(n_389) );
OAI22x1_ASAP7_75t_L g577 ( .A1(n_199), .A2(n_578), .B1(n_587), .B2(n_602), .Y(n_577) );
NAND5xp2_ASAP7_75t_SL g578 ( .A(n_199), .B(n_579), .C(n_581), .D(n_583), .E(n_585), .Y(n_578) );
INVx1_ASAP7_75t_L g717 ( .A(n_200), .Y(n_717) );
AOI22xp5_ASAP7_75t_L g884 ( .A1(n_203), .A2(n_357), .B1(n_499), .B2(n_505), .Y(n_884) );
AOI22xp33_ASAP7_75t_L g993 ( .A1(n_204), .A2(n_308), .B1(n_969), .B2(n_972), .Y(n_993) );
AOI22xp33_ASAP7_75t_L g1186 ( .A1(n_205), .A2(n_316), .B1(n_565), .B2(n_727), .Y(n_1186) );
AOI22xp33_ASAP7_75t_L g767 ( .A1(n_206), .A2(n_343), .B1(n_453), .B2(n_768), .Y(n_767) );
AOI22xp33_ASAP7_75t_L g833 ( .A1(n_207), .A2(n_346), .B1(n_383), .B2(n_584), .Y(n_833) );
INVx1_ASAP7_75t_L g724 ( .A(n_209), .Y(n_724) );
AOI22xp5_ASAP7_75t_L g968 ( .A1(n_210), .A2(n_255), .B1(n_969), .B2(n_972), .Y(n_968) );
AOI22xp33_ASAP7_75t_L g822 ( .A1(n_211), .A2(n_239), .B1(n_501), .B2(n_502), .Y(n_822) );
AOI22xp33_ASAP7_75t_L g579 ( .A1(n_212), .A2(n_252), .B1(n_406), .B2(n_580), .Y(n_579) );
AOI22xp33_ASAP7_75t_L g947 ( .A1(n_213), .A2(n_324), .B1(n_733), .B2(n_948), .Y(n_947) );
AOI22xp33_ASAP7_75t_L g819 ( .A1(n_220), .A2(n_347), .B1(n_485), .B2(n_508), .Y(n_819) );
AOI22xp5_ASAP7_75t_L g887 ( .A1(n_222), .A2(n_315), .B1(n_507), .B2(n_508), .Y(n_887) );
AOI222xp33_ASAP7_75t_L g1178 ( .A1(n_225), .A2(n_1179), .B1(n_1195), .B2(n_1199), .C1(n_1204), .C2(n_1206), .Y(n_1178) );
XNOR2x1_ASAP7_75t_L g1181 ( .A(n_225), .B(n_1182), .Y(n_1181) );
AOI22xp33_ASAP7_75t_L g898 ( .A1(n_226), .A2(n_227), .B1(n_433), .B2(n_586), .Y(n_898) );
AOI22xp33_ASAP7_75t_L g998 ( .A1(n_228), .A2(n_304), .B1(n_969), .B2(n_999), .Y(n_998) );
AOI22xp33_ASAP7_75t_L g992 ( .A1(n_230), .A2(n_300), .B1(n_966), .B2(n_989), .Y(n_992) );
INVx1_ASAP7_75t_L g451 ( .A(n_231), .Y(n_451) );
AOI22xp33_ASAP7_75t_L g484 ( .A1(n_232), .A2(n_244), .B1(n_485), .B2(n_486), .Y(n_484) );
AOI22xp5_ASAP7_75t_L g796 ( .A1(n_233), .A2(n_312), .B1(n_797), .B2(n_798), .Y(n_796) );
AOI22xp33_ASAP7_75t_L g736 ( .A1(n_234), .A2(n_349), .B1(n_737), .B2(n_739), .Y(n_736) );
AOI22xp5_ASAP7_75t_L g801 ( .A1(n_235), .A2(n_340), .B1(n_614), .B2(n_802), .Y(n_801) );
AOI22xp5_ASAP7_75t_L g899 ( .A1(n_236), .A2(n_269), .B1(n_580), .B2(n_770), .Y(n_899) );
AOI22xp33_ASAP7_75t_L g951 ( .A1(n_237), .A2(n_344), .B1(n_911), .B2(n_926), .Y(n_951) );
AOI22xp33_ASAP7_75t_L g523 ( .A1(n_238), .A2(n_325), .B1(n_485), .B2(n_504), .Y(n_523) );
AOI22xp5_ASAP7_75t_L g659 ( .A1(n_241), .A2(n_318), .B1(n_620), .B2(n_660), .Y(n_659) );
XNOR2xp5_ASAP7_75t_L g895 ( .A(n_242), .B(n_896), .Y(n_895) );
AOI22xp5_ASAP7_75t_L g977 ( .A1(n_243), .A2(n_333), .B1(n_962), .B2(n_978), .Y(n_977) );
AOI22xp33_ASAP7_75t_L g642 ( .A1(n_246), .A2(n_266), .B1(n_424), .B2(n_643), .Y(n_642) );
INVx1_ASAP7_75t_L g684 ( .A(n_248), .Y(n_684) );
NAND2xp5_ASAP7_75t_L g791 ( .A(n_249), .B(n_792), .Y(n_791) );
AOI221xp5_ASAP7_75t_SL g888 ( .A1(n_251), .A2(n_305), .B1(n_491), .B2(n_498), .C(n_889), .Y(n_888) );
INVx1_ASAP7_75t_L g828 ( .A(n_255), .Y(n_828) );
AOI22xp33_ASAP7_75t_L g514 ( .A1(n_256), .A2(n_298), .B1(n_489), .B2(n_498), .Y(n_514) );
AOI22xp5_ASAP7_75t_L g931 ( .A1(n_257), .A2(n_351), .B1(n_427), .B2(n_856), .Y(n_931) );
AOI22xp33_ASAP7_75t_L g612 ( .A1(n_259), .A2(n_278), .B1(n_406), .B2(n_580), .Y(n_612) );
INVx1_ASAP7_75t_L g748 ( .A(n_260), .Y(n_748) );
CKINVDCx5p33_ASAP7_75t_R g713 ( .A(n_261), .Y(n_713) );
AOI22xp33_ASAP7_75t_SL g563 ( .A1(n_263), .A2(n_290), .B1(n_564), .B2(n_566), .Y(n_563) );
HB1xp67_ASAP7_75t_L g370 ( .A(n_265), .Y(n_370) );
AND2x4_ASAP7_75t_L g970 ( .A(n_265), .B(n_971), .Y(n_970) );
AOI22xp5_ASAP7_75t_L g860 ( .A1(n_270), .A2(n_294), .B1(n_660), .B2(n_861), .Y(n_860) );
CKINVDCx5p33_ASAP7_75t_R g711 ( .A(n_272), .Y(n_711) );
AOI22xp33_ASAP7_75t_L g832 ( .A1(n_274), .A2(n_286), .B1(n_406), .B2(n_424), .Y(n_832) );
AOI22xp5_ASAP7_75t_L g803 ( .A1(n_275), .A2(n_319), .B1(n_417), .B2(n_670), .Y(n_803) );
NAND2xp5_ASAP7_75t_L g843 ( .A(n_276), .B(n_844), .Y(n_843) );
AOI22xp5_ASAP7_75t_L g912 ( .A1(n_279), .A2(n_306), .B1(n_417), .B2(n_614), .Y(n_912) );
INVx1_ASAP7_75t_L g654 ( .A(n_280), .Y(n_654) );
INVx1_ASAP7_75t_L g403 ( .A(n_281), .Y(n_403) );
INVxp67_ASAP7_75t_L g473 ( .A(n_281), .Y(n_473) );
AOI21xp33_ASAP7_75t_L g863 ( .A1(n_282), .A2(n_475), .B(n_864), .Y(n_863) );
INVx1_ASAP7_75t_L g909 ( .A(n_283), .Y(n_909) );
NAND2xp5_ASAP7_75t_L g922 ( .A(n_284), .B(n_443), .Y(n_922) );
INVx2_ASAP7_75t_L g365 ( .A(n_288), .Y(n_365) );
INVx1_ASAP7_75t_L g1189 ( .A(n_292), .Y(n_1189) );
AOI22xp33_ASAP7_75t_L g613 ( .A1(n_296), .A2(n_313), .B1(n_582), .B2(n_614), .Y(n_613) );
AOI221xp5_ASAP7_75t_L g679 ( .A1(n_303), .A2(n_328), .B1(n_680), .B2(n_681), .C(n_683), .Y(n_679) );
CKINVDCx5p33_ASAP7_75t_R g890 ( .A(n_307), .Y(n_890) );
CKINVDCx14_ASAP7_75t_R g760 ( .A(n_308), .Y(n_760) );
NAND2xp5_ASAP7_75t_L g859 ( .A(n_309), .B(n_719), .Y(n_859) );
NAND2xp5_ASAP7_75t_L g812 ( .A(n_311), .B(n_797), .Y(n_812) );
INVx1_ASAP7_75t_L g379 ( .A(n_314), .Y(n_379) );
AOI21xp33_ASAP7_75t_SL g549 ( .A1(n_317), .A2(n_550), .B(n_553), .Y(n_549) );
AOI22xp33_ASAP7_75t_L g497 ( .A1(n_320), .A2(n_352), .B1(n_498), .B2(n_499), .Y(n_497) );
INVx1_ASAP7_75t_L g593 ( .A(n_322), .Y(n_593) );
OAI22x1_ASAP7_75t_L g526 ( .A1(n_330), .A2(n_527), .B1(n_528), .B2(n_569), .Y(n_526) );
INVx1_ASAP7_75t_L g569 ( .A(n_330), .Y(n_569) );
AOI22x1_ASAP7_75t_L g571 ( .A1(n_330), .A2(n_527), .B1(n_528), .B2(n_569), .Y(n_571) );
NAND2xp5_ASAP7_75t_L g515 ( .A(n_354), .B(n_516), .Y(n_515) );
XNOR2x1_ASAP7_75t_L g639 ( .A(n_359), .B(n_640), .Y(n_639) );
AOI21xp5_ASAP7_75t_L g360 ( .A1(n_361), .A2(n_371), .B(n_954), .Y(n_360) );
INVx2_ASAP7_75t_SL g361 ( .A(n_362), .Y(n_361) );
NAND3xp33_ASAP7_75t_L g362 ( .A(n_363), .B(n_366), .C(n_370), .Y(n_362) );
AND2x2_ASAP7_75t_L g1196 ( .A(n_363), .B(n_1197), .Y(n_1196) );
AND2x2_ASAP7_75t_L g1205 ( .A(n_363), .B(n_1198), .Y(n_1205) );
INVx1_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
OA21x2_ASAP7_75t_L g1207 ( .A1(n_364), .A2(n_984), .B(n_1208), .Y(n_1207) );
HB1xp67_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
AND2x2_ASAP7_75t_L g963 ( .A(n_365), .B(n_964), .Y(n_963) );
AND3x4_ASAP7_75t_L g983 ( .A(n_365), .B(n_970), .C(n_984), .Y(n_983) );
NOR2xp33_ASAP7_75t_L g1197 ( .A(n_366), .B(n_1198), .Y(n_1197) );
HB1xp67_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
AO21x2_ASAP7_75t_L g456 ( .A1(n_367), .A2(n_457), .B(n_459), .Y(n_456) );
NAND2xp5_ASAP7_75t_L g367 ( .A(n_368), .B(n_369), .Y(n_367) );
INVx1_ASAP7_75t_L g1198 ( .A(n_370), .Y(n_1198) );
XNOR2xp5_ASAP7_75t_L g371 ( .A(n_372), .B(n_751), .Y(n_371) );
XNOR2xp5_ASAP7_75t_L g372 ( .A(n_373), .B(n_636), .Y(n_372) );
AOI22xp5_ASAP7_75t_L g373 ( .A1(n_374), .A2(n_375), .B1(n_572), .B2(n_573), .Y(n_373) );
INVx1_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
AO22x2_ASAP7_75t_L g375 ( .A1(n_376), .A2(n_526), .B1(n_570), .B2(n_571), .Y(n_375) );
INVx1_ASAP7_75t_L g570 ( .A(n_376), .Y(n_570) );
XNOR2xp5_ASAP7_75t_L g376 ( .A(n_377), .B(n_479), .Y(n_376) );
INVx2_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
XNOR2x1_ASAP7_75t_L g378 ( .A(n_379), .B(n_380), .Y(n_378) );
NOR2x1_ASAP7_75t_L g380 ( .A(n_381), .B(n_441), .Y(n_380) );
NAND4xp25_ASAP7_75t_L g381 ( .A(n_382), .B(n_416), .C(n_426), .D(n_432), .Y(n_381) );
BUFx6f_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
BUFx12f_ASAP7_75t_L g539 ( .A(n_384), .Y(n_539) );
BUFx6f_ASAP7_75t_L g670 ( .A(n_384), .Y(n_670) );
BUFx3_ASAP7_75t_L g780 ( .A(n_384), .Y(n_780) );
BUFx6f_ASAP7_75t_L g904 ( .A(n_384), .Y(n_904) );
AND2x4_ASAP7_75t_L g384 ( .A(n_385), .B(n_394), .Y(n_384) );
AND2x2_ASAP7_75t_L g428 ( .A(n_385), .B(n_422), .Y(n_428) );
AND2x2_ASAP7_75t_L g449 ( .A(n_385), .B(n_439), .Y(n_449) );
AND2x2_ASAP7_75t_L g464 ( .A(n_385), .B(n_435), .Y(n_464) );
AND2x4_ASAP7_75t_L g488 ( .A(n_385), .B(n_435), .Y(n_488) );
AND2x2_ASAP7_75t_L g493 ( .A(n_385), .B(n_439), .Y(n_493) );
AND2x4_ASAP7_75t_L g499 ( .A(n_385), .B(n_422), .Y(n_499) );
AND2x4_ASAP7_75t_L g505 ( .A(n_385), .B(n_415), .Y(n_505) );
AND2x2_ASAP7_75t_L g537 ( .A(n_385), .B(n_422), .Y(n_537) );
AND2x2_ASAP7_75t_L g385 ( .A(n_386), .B(n_393), .Y(n_385) );
INVx1_ASAP7_75t_L g420 ( .A(n_386), .Y(n_420) );
NAND2xp5_ASAP7_75t_L g386 ( .A(n_387), .B(n_390), .Y(n_386) );
NAND2xp33_ASAP7_75t_L g387 ( .A(n_388), .B(n_389), .Y(n_387) );
INVx2_ASAP7_75t_L g392 ( .A(n_388), .Y(n_392) );
INVx3_ASAP7_75t_L g398 ( .A(n_388), .Y(n_398) );
NAND2xp33_ASAP7_75t_L g404 ( .A(n_388), .B(n_405), .Y(n_404) );
INVx1_ASAP7_75t_L g414 ( .A(n_388), .Y(n_414) );
HB1xp67_ASAP7_75t_L g458 ( .A(n_388), .Y(n_458) );
NAND2xp5_ASAP7_75t_L g411 ( .A(n_389), .B(n_412), .Y(n_411) );
NAND2xp5_ASAP7_75t_L g390 ( .A(n_391), .B(n_392), .Y(n_390) );
OAI21xp5_ASAP7_75t_L g472 ( .A1(n_391), .A2(n_414), .B(n_473), .Y(n_472) );
INVx1_ASAP7_75t_L g421 ( .A(n_393), .Y(n_421) );
AND2x2_ASAP7_75t_L g446 ( .A(n_393), .B(n_420), .Y(n_446) );
AND2x2_ASAP7_75t_L g471 ( .A(n_393), .B(n_472), .Y(n_471) );
AND2x4_ASAP7_75t_L g485 ( .A(n_394), .B(n_419), .Y(n_485) );
INVx2_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
INVx2_ASAP7_75t_L g415 ( .A(n_395), .Y(n_415) );
OR2x2_ASAP7_75t_L g395 ( .A(n_396), .B(n_400), .Y(n_395) );
AND2x4_ASAP7_75t_L g422 ( .A(n_396), .B(n_423), .Y(n_422) );
AND2x4_ASAP7_75t_L g435 ( .A(n_396), .B(n_436), .Y(n_435) );
INVx2_ASAP7_75t_L g440 ( .A(n_396), .Y(n_440) );
AND2x2_ASAP7_75t_L g468 ( .A(n_396), .B(n_469), .Y(n_468) );
AND2x4_ASAP7_75t_L g396 ( .A(n_397), .B(n_399), .Y(n_396) );
NAND2xp5_ASAP7_75t_L g402 ( .A(n_398), .B(n_403), .Y(n_402) );
INVxp67_ASAP7_75t_L g410 ( .A(n_398), .Y(n_410) );
NAND3xp33_ASAP7_75t_L g459 ( .A(n_399), .B(n_409), .C(n_460), .Y(n_459) );
INVx1_ASAP7_75t_L g423 ( .A(n_400), .Y(n_423) );
INVx1_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
INVx1_ASAP7_75t_L g436 ( .A(n_401), .Y(n_436) );
AND2x2_ASAP7_75t_L g401 ( .A(n_402), .B(n_404), .Y(n_401) );
BUFx3_ASAP7_75t_L g534 ( .A(n_406), .Y(n_534) );
BUFx12f_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
INVx6_ASAP7_75t_L g644 ( .A(n_407), .Y(n_644) );
AND2x4_ASAP7_75t_L g407 ( .A(n_408), .B(n_415), .Y(n_407) );
AND2x4_ASAP7_75t_L g431 ( .A(n_408), .B(n_422), .Y(n_431) );
AND2x4_ASAP7_75t_L g478 ( .A(n_408), .B(n_439), .Y(n_478) );
AND2x4_ASAP7_75t_L g489 ( .A(n_408), .B(n_439), .Y(n_489) );
AND2x4_ASAP7_75t_L g507 ( .A(n_408), .B(n_422), .Y(n_507) );
AND2x4_ASAP7_75t_L g508 ( .A(n_408), .B(n_415), .Y(n_508) );
AND2x2_ASAP7_75t_L g408 ( .A(n_409), .B(n_413), .Y(n_408) );
NAND2xp5_ASAP7_75t_L g409 ( .A(n_410), .B(n_411), .Y(n_409) );
AND2x4_ASAP7_75t_L g425 ( .A(n_415), .B(n_419), .Y(n_425) );
BUFx6f_ASAP7_75t_L g545 ( .A(n_417), .Y(n_545) );
BUFx12f_ASAP7_75t_L g731 ( .A(n_417), .Y(n_731) );
BUFx12f_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
BUFx6f_ASAP7_75t_L g582 ( .A(n_418), .Y(n_582) );
BUFx6f_ASAP7_75t_L g948 ( .A(n_418), .Y(n_948) );
AND2x4_ASAP7_75t_L g418 ( .A(n_419), .B(n_422), .Y(n_418) );
AND2x4_ASAP7_75t_L g434 ( .A(n_419), .B(n_435), .Y(n_434) );
AND2x2_ASAP7_75t_L g438 ( .A(n_419), .B(n_439), .Y(n_438) );
AND2x4_ASAP7_75t_L g501 ( .A(n_419), .B(n_435), .Y(n_501) );
AND2x4_ASAP7_75t_L g502 ( .A(n_419), .B(n_439), .Y(n_502) );
AND2x4_ASAP7_75t_L g504 ( .A(n_419), .B(n_422), .Y(n_504) );
AND2x4_ASAP7_75t_L g419 ( .A(n_420), .B(n_421), .Y(n_419) );
BUFx6f_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
BUFx6f_ASAP7_75t_L g533 ( .A(n_425), .Y(n_533) );
BUFx6f_ASAP7_75t_L g580 ( .A(n_425), .Y(n_580) );
BUFx6f_ASAP7_75t_L g677 ( .A(n_425), .Y(n_677) );
BUFx6f_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
BUFx8_ASAP7_75t_L g584 ( .A(n_428), .Y(n_584) );
INVx4_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
INVx2_ASAP7_75t_L g547 ( .A(n_430), .Y(n_547) );
INVx4_ASAP7_75t_L g614 ( .A(n_430), .Y(n_614) );
INVx2_ASAP7_75t_SL g647 ( .A(n_430), .Y(n_647) );
INVx4_ASAP7_75t_L g733 ( .A(n_430), .Y(n_733) );
INVx2_ASAP7_75t_L g856 ( .A(n_430), .Y(n_856) );
INVx8_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
BUFx6f_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
INVx3_ASAP7_75t_L g542 ( .A(n_434), .Y(n_542) );
BUFx12f_ASAP7_75t_L g687 ( .A(n_434), .Y(n_687) );
AND2x4_ASAP7_75t_L g476 ( .A(n_435), .B(n_446), .Y(n_476) );
AND2x4_ASAP7_75t_L g498 ( .A(n_435), .B(n_446), .Y(n_498) );
AND2x4_ASAP7_75t_L g439 ( .A(n_436), .B(n_440), .Y(n_439) );
BUFx2_ASAP7_75t_SL g543 ( .A(n_437), .Y(n_543) );
BUFx6f_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
BUFx5_ASAP7_75t_L g586 ( .A(n_438), .Y(n_586) );
INVx1_ASAP7_75t_L g742 ( .A(n_438), .Y(n_742) );
BUFx3_ASAP7_75t_L g802 ( .A(n_438), .Y(n_802) );
AND2x4_ASAP7_75t_L g445 ( .A(n_439), .B(n_446), .Y(n_445) );
AND2x2_ASAP7_75t_L g702 ( .A(n_439), .B(n_446), .Y(n_702) );
NAND3xp33_ASAP7_75t_L g441 ( .A(n_442), .B(n_461), .C(n_474), .Y(n_441) );
INVx3_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
INVx2_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
BUFx6f_ASAP7_75t_L g491 ( .A(n_445), .Y(n_491) );
BUFx6f_ASAP7_75t_L g516 ( .A(n_445), .Y(n_516) );
INVx2_ASAP7_75t_L g601 ( .A(n_445), .Y(n_601) );
BUFx8_ASAP7_75t_SL g619 ( .A(n_445), .Y(n_619) );
BUFx3_ASAP7_75t_L g792 ( .A(n_445), .Y(n_792) );
INVx3_ASAP7_75t_SL g447 ( .A(n_448), .Y(n_447) );
INVx2_ASAP7_75t_L g652 ( .A(n_448), .Y(n_652) );
INVx2_ASAP7_75t_L g764 ( .A(n_448), .Y(n_764) );
INVx2_ASAP7_75t_L g921 ( .A(n_448), .Y(n_921) );
INVx3_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
BUFx3_ASAP7_75t_L g552 ( .A(n_449), .Y(n_552) );
INVx2_ASAP7_75t_L g598 ( .A(n_449), .Y(n_598) );
NOR2xp33_ASAP7_75t_L g450 ( .A(n_451), .B(n_452), .Y(n_450) );
INVx2_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
INVx4_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
NOR2xp33_ASAP7_75t_L g494 ( .A(n_454), .B(n_495), .Y(n_494) );
NOR2xp33_ASAP7_75t_L g592 ( .A(n_454), .B(n_593), .Y(n_592) );
NOR2xp33_ASAP7_75t_L g816 ( .A(n_454), .B(n_817), .Y(n_816) );
INVx4_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
INVx3_ASAP7_75t_L g559 ( .A(n_455), .Y(n_559) );
INVx3_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
BUFx6f_ASAP7_75t_L g520 ( .A(n_456), .Y(n_520) );
INVx1_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
NAND2xp5_ASAP7_75t_L g469 ( .A(n_458), .B(n_470), .Y(n_469) );
INVx1_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
BUFx6f_ASAP7_75t_L g661 ( .A(n_463), .Y(n_661) );
INVx2_ASAP7_75t_L g777 ( .A(n_463), .Y(n_777) );
INVx2_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
BUFx3_ASAP7_75t_L g568 ( .A(n_464), .Y(n_568) );
BUFx6f_ASAP7_75t_L g926 ( .A(n_464), .Y(n_926) );
INVx2_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
INVx4_ASAP7_75t_L g658 ( .A(n_466), .Y(n_658) );
INVx2_ASAP7_75t_L g673 ( .A(n_466), .Y(n_673) );
INVx3_ASAP7_75t_L g768 ( .A(n_466), .Y(n_768) );
INVx2_ASAP7_75t_L g861 ( .A(n_466), .Y(n_861) );
INVx5_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
BUFx4f_ASAP7_75t_L g556 ( .A(n_467), .Y(n_556) );
BUFx2_ASAP7_75t_L g902 ( .A(n_467), .Y(n_902) );
AND2x4_ASAP7_75t_L g467 ( .A(n_468), .B(n_471), .Y(n_467) );
AND2x2_ASAP7_75t_L g486 ( .A(n_468), .B(n_471), .Y(n_486) );
AND2x4_ASAP7_75t_L g628 ( .A(n_468), .B(n_471), .Y(n_628) );
INVx4_ASAP7_75t_L g712 ( .A(n_475), .Y(n_712) );
BUFx6f_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
BUFx3_ASAP7_75t_L g565 ( .A(n_476), .Y(n_565) );
BUFx3_ASAP7_75t_L g591 ( .A(n_476), .Y(n_591) );
INVx1_ASAP7_75t_L g842 ( .A(n_476), .Y(n_842) );
BUFx3_ASAP7_75t_L g562 ( .A(n_477), .Y(n_562) );
BUFx6f_ASAP7_75t_L g477 ( .A(n_478), .Y(n_477) );
INVx3_ASAP7_75t_L g621 ( .A(n_478), .Y(n_621) );
BUFx6f_ASAP7_75t_L g727 ( .A(n_478), .Y(n_727) );
OAI22xp5_ASAP7_75t_L g479 ( .A1(n_480), .A2(n_481), .B1(n_509), .B2(n_510), .Y(n_479) );
INVx1_ASAP7_75t_SL g480 ( .A(n_481), .Y(n_480) );
INVx1_ASAP7_75t_L g631 ( .A(n_481), .Y(n_631) );
NOR2x1_ASAP7_75t_L g482 ( .A(n_483), .B(n_496), .Y(n_482) );
NAND4xp25_ASAP7_75t_L g483 ( .A(n_484), .B(n_487), .C(n_490), .D(n_492), .Y(n_483) );
INVx2_ASAP7_75t_L g682 ( .A(n_493), .Y(n_682) );
NAND4xp25_ASAP7_75t_L g496 ( .A(n_497), .B(n_500), .C(n_503), .D(n_506), .Y(n_496) );
INVx2_ASAP7_75t_L g509 ( .A(n_510), .Y(n_509) );
OR2x2_ASAP7_75t_L g511 ( .A(n_512), .B(n_521), .Y(n_511) );
NAND4xp25_ASAP7_75t_L g512 ( .A(n_513), .B(n_514), .C(n_515), .D(n_517), .Y(n_512) );
BUFx3_ASAP7_75t_L g561 ( .A(n_516), .Y(n_561) );
NOR2xp33_ASAP7_75t_L g518 ( .A(n_519), .B(n_520), .Y(n_518) );
INVx2_ASAP7_75t_L g656 ( .A(n_520), .Y(n_656) );
BUFx6f_ASAP7_75t_L g685 ( .A(n_520), .Y(n_685) );
BUFx6f_ASAP7_75t_L g799 ( .A(n_520), .Y(n_799) );
INVx2_ASAP7_75t_SL g846 ( .A(n_520), .Y(n_846) );
INVx1_ASAP7_75t_L g867 ( .A(n_520), .Y(n_867) );
NOR2xp33_ASAP7_75t_L g889 ( .A(n_520), .B(n_890), .Y(n_889) );
NAND4xp25_ASAP7_75t_L g521 ( .A(n_522), .B(n_523), .C(n_524), .D(n_525), .Y(n_521) );
INVx2_ASAP7_75t_L g527 ( .A(n_528), .Y(n_527) );
OR2x2_ASAP7_75t_L g528 ( .A(n_529), .B(n_548), .Y(n_528) );
NAND4xp25_ASAP7_75t_SL g529 ( .A(n_530), .B(n_535), .C(n_540), .D(n_544), .Y(n_529) );
INVx1_ASAP7_75t_L g531 ( .A(n_532), .Y(n_531) );
INVx1_ASAP7_75t_L g532 ( .A(n_533), .Y(n_532) );
BUFx3_ASAP7_75t_L g744 ( .A(n_533), .Y(n_744) );
BUFx6f_ASAP7_75t_L g536 ( .A(n_537), .Y(n_536) );
BUFx4f_ASAP7_75t_L g669 ( .A(n_537), .Y(n_669) );
BUFx3_ASAP7_75t_L g538 ( .A(n_539), .Y(n_538) );
INVx1_ASAP7_75t_L g541 ( .A(n_542), .Y(n_541) );
INVx1_ASAP7_75t_L g649 ( .A(n_542), .Y(n_649) );
INVx2_ASAP7_75t_L g738 ( .A(n_542), .Y(n_738) );
BUFx2_ASAP7_75t_SL g546 ( .A(n_547), .Y(n_546) );
NAND3xp33_ASAP7_75t_L g548 ( .A(n_549), .B(n_560), .C(n_563), .Y(n_548) );
HB1xp67_ASAP7_75t_L g550 ( .A(n_551), .Y(n_550) );
BUFx3_ASAP7_75t_L g551 ( .A(n_552), .Y(n_551) );
INVx2_ASAP7_75t_L g624 ( .A(n_552), .Y(n_624) );
OAI21xp33_ASAP7_75t_L g553 ( .A1(n_554), .A2(n_555), .B(n_557), .Y(n_553) );
INVx2_ASAP7_75t_SL g555 ( .A(n_556), .Y(n_555) );
INVx4_ASAP7_75t_L g558 ( .A(n_559), .Y(n_558) );
NOR2xp33_ASAP7_75t_L g699 ( .A(n_559), .B(n_700), .Y(n_699) );
NOR2xp33_ASAP7_75t_L g908 ( .A(n_559), .B(n_909), .Y(n_908) );
INVx1_ASAP7_75t_L g723 ( .A(n_561), .Y(n_723) );
BUFx2_ASAP7_75t_L g564 ( .A(n_565), .Y(n_564) );
INVx2_ASAP7_75t_L g566 ( .A(n_567), .Y(n_566) );
INVx2_ASAP7_75t_L g567 ( .A(n_568), .Y(n_567) );
BUFx2_ASAP7_75t_L g715 ( .A(n_568), .Y(n_715) );
INVxp67_ASAP7_75t_L g572 ( .A(n_573), .Y(n_572) );
AOI22xp5_ASAP7_75t_L g573 ( .A1(n_574), .A2(n_606), .B1(n_633), .B2(n_635), .Y(n_573) );
INVx1_ASAP7_75t_L g574 ( .A(n_575), .Y(n_574) );
BUFx3_ASAP7_75t_L g575 ( .A(n_576), .Y(n_575) );
INVx2_ASAP7_75t_L g634 ( .A(n_576), .Y(n_634) );
BUFx3_ASAP7_75t_L g576 ( .A(n_577), .Y(n_576) );
NAND4xp25_ASAP7_75t_L g603 ( .A(n_579), .B(n_581), .C(n_585), .D(n_595), .Y(n_603) );
NAND2xp5_ASAP7_75t_L g605 ( .A(n_583), .B(n_599), .Y(n_605) );
NAND3xp33_ASAP7_75t_L g587 ( .A(n_588), .B(n_595), .C(n_599), .Y(n_587) );
INVxp67_ASAP7_75t_L g588 ( .A(n_589), .Y(n_588) );
OR2x2_ASAP7_75t_L g604 ( .A(n_589), .B(n_605), .Y(n_604) );
NAND2xp5_ASAP7_75t_L g589 ( .A(n_590), .B(n_594), .Y(n_589) );
HB1xp67_ASAP7_75t_L g778 ( .A(n_591), .Y(n_778) );
INVx2_ASAP7_75t_L g596 ( .A(n_597), .Y(n_596) );
INVx2_ASAP7_75t_L g719 ( .A(n_597), .Y(n_719) );
INVx2_ASAP7_75t_L g941 ( .A(n_597), .Y(n_941) );
BUFx6f_ASAP7_75t_L g597 ( .A(n_598), .Y(n_597) );
INVx2_ASAP7_75t_L g797 ( .A(n_598), .Y(n_797) );
INVx2_ASAP7_75t_SL g600 ( .A(n_601), .Y(n_600) );
INVx2_ASAP7_75t_SL g680 ( .A(n_601), .Y(n_680) );
NOR2x1_ASAP7_75t_L g602 ( .A(n_603), .B(n_604), .Y(n_602) );
INVx2_ASAP7_75t_L g635 ( .A(n_606), .Y(n_635) );
OA22x2_ASAP7_75t_L g606 ( .A1(n_607), .A2(n_630), .B1(n_631), .B2(n_632), .Y(n_606) );
INVx1_ASAP7_75t_L g632 ( .A(n_607), .Y(n_632) );
XNOR2x1_ASAP7_75t_L g607 ( .A(n_608), .B(n_609), .Y(n_607) );
NOR2x1_ASAP7_75t_L g609 ( .A(n_610), .B(n_616), .Y(n_609) );
NAND4xp25_ASAP7_75t_L g610 ( .A(n_611), .B(n_612), .C(n_613), .D(n_615), .Y(n_610) );
NAND3xp33_ASAP7_75t_L g616 ( .A(n_617), .B(n_618), .C(n_622), .Y(n_616) );
INVx3_ASAP7_75t_L g620 ( .A(n_621), .Y(n_620) );
INVx2_ASAP7_75t_L g911 ( .A(n_621), .Y(n_911) );
INVx2_ASAP7_75t_L g623 ( .A(n_624), .Y(n_623) );
OAI21xp5_ASAP7_75t_L g625 ( .A1(n_626), .A2(n_627), .B(n_629), .Y(n_625) );
INVx4_ASAP7_75t_L g627 ( .A(n_628), .Y(n_627) );
INVx1_ASAP7_75t_L g630 ( .A(n_631), .Y(n_630) );
INVx2_ASAP7_75t_L g633 ( .A(n_634), .Y(n_633) );
AOI22xp5_ASAP7_75t_L g636 ( .A1(n_637), .A2(n_662), .B1(n_749), .B2(n_750), .Y(n_636) );
INVxp67_ASAP7_75t_L g750 ( .A(n_637), .Y(n_750) );
INVx1_ASAP7_75t_L g637 ( .A(n_638), .Y(n_637) );
INVx2_ASAP7_75t_L g638 ( .A(n_639), .Y(n_638) );
NOR2x1_ASAP7_75t_L g640 ( .A(n_641), .B(n_650), .Y(n_640) );
NAND4xp25_ASAP7_75t_L g641 ( .A(n_642), .B(n_645), .C(n_646), .D(n_648), .Y(n_641) );
INVx3_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
INVx5_ASAP7_75t_L g678 ( .A(n_644), .Y(n_678) );
INVx2_ASAP7_75t_L g747 ( .A(n_644), .Y(n_747) );
INVx1_ASAP7_75t_L g770 ( .A(n_644), .Y(n_770) );
NAND3xp33_ASAP7_75t_L g650 ( .A(n_651), .B(n_657), .C(n_659), .Y(n_650) );
NOR2xp33_ASAP7_75t_L g653 ( .A(n_654), .B(n_655), .Y(n_653) );
NOR2xp33_ASAP7_75t_L g943 ( .A(n_655), .B(n_944), .Y(n_943) );
INVx3_ASAP7_75t_L g655 ( .A(n_656), .Y(n_655) );
INVx2_ASAP7_75t_L g660 ( .A(n_661), .Y(n_660) );
INVx2_ASAP7_75t_L g749 ( .A(n_662), .Y(n_749) );
OA22x2_ASAP7_75t_L g662 ( .A1(n_663), .A2(n_664), .B1(n_706), .B2(n_707), .Y(n_662) );
INVx2_ASAP7_75t_L g663 ( .A(n_664), .Y(n_663) );
OA22x2_ASAP7_75t_L g664 ( .A1(n_665), .A2(n_688), .B1(n_704), .B2(n_705), .Y(n_664) );
INVx1_ASAP7_75t_L g704 ( .A(n_665), .Y(n_704) );
NOR2x1_ASAP7_75t_L g666 ( .A(n_667), .B(n_675), .Y(n_666) );
NAND4xp25_ASAP7_75t_L g667 ( .A(n_668), .B(n_671), .C(n_672), .D(n_674), .Y(n_667) );
NAND3xp33_ASAP7_75t_L g675 ( .A(n_676), .B(n_679), .C(n_686), .Y(n_675) );
INVx2_ASAP7_75t_L g681 ( .A(n_682), .Y(n_681) );
NOR2xp33_ASAP7_75t_L g683 ( .A(n_684), .B(n_685), .Y(n_683) );
NOR2xp33_ASAP7_75t_L g1188 ( .A(n_685), .B(n_1189), .Y(n_1188) );
INVx2_ASAP7_75t_L g705 ( .A(n_688), .Y(n_705) );
XOR2x2_ASAP7_75t_L g688 ( .A(n_689), .B(n_703), .Y(n_688) );
NOR2xp67_ASAP7_75t_L g689 ( .A(n_690), .B(n_695), .Y(n_689) );
NAND4xp25_ASAP7_75t_L g690 ( .A(n_691), .B(n_692), .C(n_693), .D(n_694), .Y(n_690) );
NAND4xp25_ASAP7_75t_L g695 ( .A(n_696), .B(n_697), .C(n_698), .D(n_701), .Y(n_695) );
INVx2_ASAP7_75t_SL g706 ( .A(n_707), .Y(n_706) );
XOR2x2_ASAP7_75t_L g707 ( .A(n_708), .B(n_748), .Y(n_707) );
NAND2xp5_ASAP7_75t_L g708 ( .A(n_709), .B(n_728), .Y(n_708) );
NOR3xp33_ASAP7_75t_L g709 ( .A(n_710), .B(n_716), .C(n_721), .Y(n_709) );
OAI22xp5_ASAP7_75t_L g710 ( .A1(n_711), .A2(n_712), .B1(n_713), .B2(n_714), .Y(n_710) );
INVx1_ASAP7_75t_L g714 ( .A(n_715), .Y(n_714) );
OAI21xp33_ASAP7_75t_L g716 ( .A1(n_717), .A2(n_718), .B(n_720), .Y(n_716) );
INVx2_ASAP7_75t_L g718 ( .A(n_719), .Y(n_718) );
OAI22xp5_ASAP7_75t_L g721 ( .A1(n_722), .A2(n_723), .B1(n_724), .B2(n_725), .Y(n_721) );
INVx1_ASAP7_75t_L g725 ( .A(n_726), .Y(n_725) );
BUFx3_ASAP7_75t_L g726 ( .A(n_727), .Y(n_726) );
NOR2xp67_ASAP7_75t_L g728 ( .A(n_729), .B(n_735), .Y(n_728) );
NAND2xp5_ASAP7_75t_L g729 ( .A(n_730), .B(n_734), .Y(n_729) );
BUFx2_ASAP7_75t_L g732 ( .A(n_733), .Y(n_732) );
NAND2xp5_ASAP7_75t_L g735 ( .A(n_736), .B(n_743), .Y(n_735) );
BUFx4f_ASAP7_75t_L g737 ( .A(n_738), .Y(n_737) );
INVx1_ASAP7_75t_L g739 ( .A(n_740), .Y(n_739) );
INVx1_ASAP7_75t_L g835 ( .A(n_740), .Y(n_835) );
INVx1_ASAP7_75t_L g740 ( .A(n_741), .Y(n_740) );
BUFx6f_ASAP7_75t_L g772 ( .A(n_741), .Y(n_772) );
INVx2_ASAP7_75t_L g741 ( .A(n_742), .Y(n_741) );
INVx1_ASAP7_75t_L g745 ( .A(n_746), .Y(n_745) );
INVx1_ASAP7_75t_L g746 ( .A(n_747), .Y(n_746) );
OAI22xp5_ASAP7_75t_L g751 ( .A1(n_752), .A2(n_753), .B1(n_875), .B2(n_876), .Y(n_751) );
INVx1_ASAP7_75t_L g752 ( .A(n_753), .Y(n_752) );
AOI22xp5_ASAP7_75t_L g753 ( .A1(n_754), .A2(n_824), .B1(n_825), .B2(n_874), .Y(n_753) );
INVx1_ASAP7_75t_L g754 ( .A(n_755), .Y(n_754) );
INVx1_ASAP7_75t_L g755 ( .A(n_756), .Y(n_755) );
INVxp67_ASAP7_75t_SL g874 ( .A(n_756), .Y(n_874) );
INVx1_ASAP7_75t_L g756 ( .A(n_757), .Y(n_756) );
XNOR2x1_ASAP7_75t_L g757 ( .A(n_758), .B(n_781), .Y(n_757) );
INVx2_ASAP7_75t_L g758 ( .A(n_759), .Y(n_758) );
XNOR2x2_ASAP7_75t_L g759 ( .A(n_760), .B(n_761), .Y(n_759) );
NAND3xp33_ASAP7_75t_L g761 ( .A(n_762), .B(n_771), .C(n_775), .Y(n_761) );
HB1xp67_ASAP7_75t_L g763 ( .A(n_764), .Y(n_763) );
NAND2xp5_ASAP7_75t_L g765 ( .A(n_766), .B(n_767), .Y(n_765) );
INVx1_ASAP7_75t_L g773 ( .A(n_774), .Y(n_773) );
BUFx3_ASAP7_75t_L g776 ( .A(n_777), .Y(n_776) );
AO22x2_ASAP7_75t_L g781 ( .A1(n_782), .A2(n_783), .B1(n_807), .B2(n_808), .Y(n_781) );
INVx2_ASAP7_75t_SL g782 ( .A(n_783), .Y(n_782) );
XOR2x2_ASAP7_75t_L g848 ( .A(n_783), .B(n_849), .Y(n_848) );
AO21x2_ASAP7_75t_L g783 ( .A1(n_784), .A2(n_793), .B(n_804), .Y(n_783) );
NAND2xp5_ASAP7_75t_L g785 ( .A(n_786), .B(n_787), .Y(n_785) );
NAND2xp5_ASAP7_75t_SL g789 ( .A(n_790), .B(n_791), .Y(n_789) );
NOR2xp33_ASAP7_75t_L g793 ( .A(n_794), .B(n_800), .Y(n_793) );
NAND2xp5_ASAP7_75t_L g794 ( .A(n_795), .B(n_796), .Y(n_794) );
BUFx3_ASAP7_75t_L g844 ( .A(n_797), .Y(n_844) );
INVx2_ASAP7_75t_L g798 ( .A(n_799), .Y(n_798) );
NAND2x1_ASAP7_75t_SL g800 ( .A(n_801), .B(n_803), .Y(n_800) );
NAND2xp5_ASAP7_75t_L g804 ( .A(n_805), .B(n_806), .Y(n_804) );
INVx2_ASAP7_75t_L g807 ( .A(n_808), .Y(n_807) );
AO21x2_ASAP7_75t_L g808 ( .A1(n_809), .A2(n_810), .B(n_823), .Y(n_808) );
NOR3xp33_ASAP7_75t_SL g823 ( .A(n_809), .B(n_811), .C(n_818), .Y(n_823) );
OR2x2_ASAP7_75t_L g810 ( .A(n_811), .B(n_818), .Y(n_810) );
NAND4xp75_ASAP7_75t_L g811 ( .A(n_812), .B(n_813), .C(n_814), .D(n_815), .Y(n_811) );
NAND4xp25_ASAP7_75t_L g818 ( .A(n_819), .B(n_820), .C(n_821), .D(n_822), .Y(n_818) );
INVx1_ASAP7_75t_L g824 ( .A(n_825), .Y(n_824) );
XOR2x1_ASAP7_75t_L g825 ( .A(n_826), .B(n_848), .Y(n_825) );
INVx2_ASAP7_75t_L g826 ( .A(n_827), .Y(n_826) );
AO21x2_ASAP7_75t_L g827 ( .A1(n_828), .A2(n_829), .B(n_847), .Y(n_827) );
NOR3xp33_ASAP7_75t_SL g847 ( .A(n_828), .B(n_831), .C(n_838), .Y(n_847) );
NAND2xp5_ASAP7_75t_L g829 ( .A(n_830), .B(n_837), .Y(n_829) );
INVx1_ASAP7_75t_L g830 ( .A(n_831), .Y(n_830) );
NAND4xp25_ASAP7_75t_SL g831 ( .A(n_832), .B(n_833), .C(n_834), .D(n_836), .Y(n_831) );
INVx1_ASAP7_75t_L g837 ( .A(n_838), .Y(n_837) );
NAND4xp25_ASAP7_75t_L g838 ( .A(n_839), .B(n_840), .C(n_843), .D(n_845), .Y(n_838) );
INVx2_ASAP7_75t_L g841 ( .A(n_842), .Y(n_841) );
INVx2_ASAP7_75t_L g924 ( .A(n_842), .Y(n_924) );
OAI21xp5_ASAP7_75t_L g849 ( .A1(n_850), .A2(n_851), .B(n_868), .Y(n_849) );
NAND2xp5_ASAP7_75t_L g871 ( .A(n_850), .B(n_860), .Y(n_871) );
NOR2xp67_ASAP7_75t_L g851 ( .A(n_852), .B(n_858), .Y(n_851) );
INVx1_ASAP7_75t_L g869 ( .A(n_852), .Y(n_869) );
NAND4xp25_ASAP7_75t_L g852 ( .A(n_853), .B(n_854), .C(n_855), .D(n_857), .Y(n_852) );
NAND4xp25_ASAP7_75t_L g858 ( .A(n_859), .B(n_860), .C(n_862), .D(n_863), .Y(n_858) );
INVx1_ASAP7_75t_L g872 ( .A(n_859), .Y(n_872) );
NAND2xp5_ASAP7_75t_L g873 ( .A(n_862), .B(n_863), .Y(n_873) );
NOR2xp33_ASAP7_75t_L g864 ( .A(n_865), .B(n_866), .Y(n_864) );
INVx1_ASAP7_75t_L g866 ( .A(n_867), .Y(n_866) );
NAND2xp5_ASAP7_75t_L g868 ( .A(n_869), .B(n_870), .Y(n_868) );
NOR3xp33_ASAP7_75t_L g870 ( .A(n_871), .B(n_872), .C(n_873), .Y(n_870) );
INVx1_ASAP7_75t_L g875 ( .A(n_876), .Y(n_875) );
OAI22xp5_ASAP7_75t_L g876 ( .A1(n_877), .A2(n_932), .B1(n_952), .B2(n_953), .Y(n_876) );
INVx1_ASAP7_75t_L g877 ( .A(n_878), .Y(n_877) );
HB1xp67_ASAP7_75t_L g952 ( .A(n_878), .Y(n_952) );
XOR2x2_ASAP7_75t_L g878 ( .A(n_879), .B(n_914), .Y(n_878) );
OAI22xp5_ASAP7_75t_L g879 ( .A1(n_880), .A2(n_881), .B1(n_895), .B2(n_913), .Y(n_879) );
INVx2_ASAP7_75t_L g880 ( .A(n_881), .Y(n_880) );
INVx1_ASAP7_75t_L g893 ( .A(n_882), .Y(n_893) );
NAND3xp33_ASAP7_75t_L g882 ( .A(n_883), .B(n_888), .C(n_891), .Y(n_882) );
AND4x1_ASAP7_75t_L g883 ( .A(n_884), .B(n_885), .C(n_886), .D(n_887), .Y(n_883) );
INVx1_ASAP7_75t_L g913 ( .A(n_895), .Y(n_913) );
NOR3xp33_ASAP7_75t_L g896 ( .A(n_897), .B(n_900), .C(n_905), .Y(n_896) );
NAND2xp5_ASAP7_75t_L g897 ( .A(n_898), .B(n_899), .Y(n_897) );
NAND2xp5_ASAP7_75t_SL g900 ( .A(n_901), .B(n_903), .Y(n_900) );
NAND4xp25_ASAP7_75t_SL g905 ( .A(n_906), .B(n_907), .C(n_910), .D(n_912), .Y(n_905) );
INVx1_ASAP7_75t_L g914 ( .A(n_915), .Y(n_914) );
XNOR2xp5_ASAP7_75t_L g915 ( .A(n_916), .B(n_918), .Y(n_915) );
CKINVDCx5p33_ASAP7_75t_R g916 ( .A(n_917), .Y(n_916) );
NOR2x1_ASAP7_75t_L g918 ( .A(n_919), .B(n_927), .Y(n_918) );
NAND4xp25_ASAP7_75t_L g919 ( .A(n_920), .B(n_922), .C(n_923), .D(n_925), .Y(n_919) );
NAND4xp25_ASAP7_75t_L g927 ( .A(n_928), .B(n_929), .C(n_930), .D(n_931), .Y(n_927) );
HB1xp67_ASAP7_75t_L g932 ( .A(n_933), .Y(n_932) );
INVx2_ASAP7_75t_L g953 ( .A(n_933), .Y(n_953) );
NAND4xp75_ASAP7_75t_L g934 ( .A(n_935), .B(n_938), .C(n_945), .D(n_949), .Y(n_934) );
AND2x2_ASAP7_75t_L g935 ( .A(n_936), .B(n_937), .Y(n_935) );
OA21x2_ASAP7_75t_L g938 ( .A1(n_939), .A2(n_940), .B(n_942), .Y(n_938) );
INVx1_ASAP7_75t_L g940 ( .A(n_941), .Y(n_940) );
AND2x2_ASAP7_75t_L g945 ( .A(n_946), .B(n_947), .Y(n_945) );
AND2x2_ASAP7_75t_L g949 ( .A(n_950), .B(n_951), .Y(n_949) );
OAI21xp5_ASAP7_75t_SL g954 ( .A1(n_955), .A2(n_1175), .B(n_1178), .Y(n_954) );
AOI211xp5_ASAP7_75t_L g955 ( .A1(n_956), .A2(n_1086), .B(n_1093), .C(n_1142), .Y(n_955) );
NAND5xp2_ASAP7_75t_L g956 ( .A(n_957), .B(n_1031), .C(n_1056), .D(n_1068), .E(n_1073), .Y(n_956) );
AOI211xp5_ASAP7_75t_SL g957 ( .A1(n_958), .A2(n_990), .B(n_994), .C(n_1023), .Y(n_957) );
AND2x2_ASAP7_75t_L g958 ( .A(n_959), .B(n_973), .Y(n_958) );
NOR2xp33_ASAP7_75t_L g1025 ( .A(n_959), .B(n_1022), .Y(n_1025) );
NAND2xp5_ASAP7_75t_L g1072 ( .A(n_959), .B(n_1030), .Y(n_1072) );
AND2x2_ASAP7_75t_L g1074 ( .A(n_959), .B(n_1075), .Y(n_1074) );
NOR2xp33_ASAP7_75t_L g1126 ( .A(n_959), .B(n_1127), .Y(n_1126) );
NOR2xp33_ASAP7_75t_L g1159 ( .A(n_959), .B(n_1160), .Y(n_1159) );
INVx2_ASAP7_75t_L g959 ( .A(n_960), .Y(n_959) );
INVx3_ASAP7_75t_L g1017 ( .A(n_960), .Y(n_1017) );
AND2x2_ASAP7_75t_L g1055 ( .A(n_960), .B(n_1038), .Y(n_1055) );
NAND2xp5_ASAP7_75t_L g1063 ( .A(n_960), .B(n_996), .Y(n_1063) );
INVx2_ASAP7_75t_L g1096 ( .A(n_960), .Y(n_1096) );
NAND2xp5_ASAP7_75t_L g1105 ( .A(n_960), .B(n_1067), .Y(n_1105) );
NOR3xp33_ASAP7_75t_L g1152 ( .A(n_960), .B(n_1020), .C(n_1088), .Y(n_1152) );
NOR2xp33_ASAP7_75t_L g1174 ( .A(n_960), .B(n_1078), .Y(n_1174) );
AND2x2_ASAP7_75t_L g960 ( .A(n_961), .B(n_968), .Y(n_960) );
AND2x2_ASAP7_75t_L g962 ( .A(n_963), .B(n_965), .Y(n_962) );
AND2x4_ASAP7_75t_L g969 ( .A(n_963), .B(n_970), .Y(n_969) );
AND2x2_ASAP7_75t_L g986 ( .A(n_963), .B(n_965), .Y(n_986) );
AND2x4_ASAP7_75t_L g989 ( .A(n_963), .B(n_965), .Y(n_989) );
AND2x2_ASAP7_75t_L g966 ( .A(n_965), .B(n_967), .Y(n_966) );
AND2x2_ASAP7_75t_L g978 ( .A(n_965), .B(n_967), .Y(n_978) );
AND2x4_ASAP7_75t_L g1002 ( .A(n_965), .B(n_967), .Y(n_1002) );
AND2x4_ASAP7_75t_L g972 ( .A(n_967), .B(n_970), .Y(n_972) );
AND2x4_ASAP7_75t_L g976 ( .A(n_967), .B(n_970), .Y(n_976) );
NAND2xp5_ASAP7_75t_L g1177 ( .A(n_967), .B(n_970), .Y(n_1177) );
INVx3_ASAP7_75t_L g1091 ( .A(n_969), .Y(n_1091) );
CKINVDCx5p33_ASAP7_75t_R g1208 ( .A(n_970), .Y(n_1208) );
INVx2_ASAP7_75t_SL g1000 ( .A(n_972), .Y(n_1000) );
NAND2xp5_ASAP7_75t_L g1110 ( .A(n_973), .B(n_1028), .Y(n_1110) );
AND2x2_ASAP7_75t_L g973 ( .A(n_974), .B(n_979), .Y(n_973) );
AND2x2_ASAP7_75t_L g1015 ( .A(n_974), .B(n_1016), .Y(n_1015) );
AND2x2_ASAP7_75t_L g1030 ( .A(n_974), .B(n_1019), .Y(n_1030) );
AND2x2_ASAP7_75t_L g1032 ( .A(n_974), .B(n_1033), .Y(n_1032) );
CKINVDCx6p67_ASAP7_75t_R g1038 ( .A(n_974), .Y(n_1038) );
AOI32xp33_ASAP7_75t_L g1073 ( .A1(n_974), .A2(n_1074), .A3(n_1076), .B1(n_1079), .B2(n_1083), .Y(n_1073) );
NOR2xp33_ASAP7_75t_L g1085 ( .A(n_974), .B(n_980), .Y(n_1085) );
AND2x2_ASAP7_75t_L g1097 ( .A(n_974), .B(n_1013), .Y(n_1097) );
NAND2xp5_ASAP7_75t_L g1115 ( .A(n_974), .B(n_1020), .Y(n_1115) );
AND2x2_ASAP7_75t_L g1135 ( .A(n_974), .B(n_981), .Y(n_1135) );
AND2x2_ASAP7_75t_L g974 ( .A(n_975), .B(n_977), .Y(n_974) );
NAND2xp5_ASAP7_75t_L g1059 ( .A(n_979), .B(n_1015), .Y(n_1059) );
INVx1_ASAP7_75t_L g1078 ( .A(n_979), .Y(n_1078) );
AND2x2_ASAP7_75t_L g1101 ( .A(n_979), .B(n_1038), .Y(n_1101) );
AND2x2_ASAP7_75t_L g1109 ( .A(n_979), .B(n_1055), .Y(n_1109) );
AND2x2_ASAP7_75t_L g979 ( .A(n_980), .B(n_987), .Y(n_979) );
OAI221xp5_ASAP7_75t_L g1147 ( .A1(n_980), .A2(n_1028), .B1(n_1123), .B2(n_1148), .C(n_1149), .Y(n_1147) );
NAND2xp5_ASAP7_75t_L g1160 ( .A(n_980), .B(n_1038), .Y(n_1160) );
INVx1_ASAP7_75t_L g980 ( .A(n_981), .Y(n_980) );
OR2x2_ASAP7_75t_L g1014 ( .A(n_981), .B(n_987), .Y(n_1014) );
AND2x2_ASAP7_75t_L g1019 ( .A(n_981), .B(n_1020), .Y(n_1019) );
AND2x2_ASAP7_75t_L g1034 ( .A(n_981), .B(n_987), .Y(n_1034) );
AND2x2_ASAP7_75t_L g981 ( .A(n_982), .B(n_985), .Y(n_981) );
INVx1_ASAP7_75t_L g1020 ( .A(n_987), .Y(n_1020) );
NAND2xp5_ASAP7_75t_L g1044 ( .A(n_987), .B(n_1015), .Y(n_1044) );
AND2x2_ASAP7_75t_L g1132 ( .A(n_987), .B(n_1038), .Y(n_1132) );
INVxp67_ASAP7_75t_L g1003 ( .A(n_990), .Y(n_1003) );
OR2x2_ASAP7_75t_L g1043 ( .A(n_990), .B(n_1009), .Y(n_1043) );
OR2x2_ASAP7_75t_L g1048 ( .A(n_990), .B(n_1008), .Y(n_1048) );
AND2x2_ASAP7_75t_L g1067 ( .A(n_990), .B(n_1009), .Y(n_1067) );
INVx2_ASAP7_75t_L g1071 ( .A(n_990), .Y(n_1071) );
AND2x2_ASAP7_75t_L g1082 ( .A(n_990), .B(n_996), .Y(n_1082) );
INVx2_ASAP7_75t_L g990 ( .A(n_991), .Y(n_990) );
OR2x2_ASAP7_75t_L g1022 ( .A(n_991), .B(n_1009), .Y(n_1022) );
AND2x2_ASAP7_75t_L g1039 ( .A(n_991), .B(n_997), .Y(n_1039) );
NAND2xp5_ASAP7_75t_L g991 ( .A(n_992), .B(n_993), .Y(n_991) );
OAI21xp33_ASAP7_75t_L g994 ( .A1(n_995), .A2(n_1004), .B(n_1018), .Y(n_994) );
INVx1_ASAP7_75t_L g1130 ( .A(n_995), .Y(n_1130) );
AOI21xp33_ASAP7_75t_SL g1162 ( .A1(n_995), .A2(n_1145), .B(n_1163), .Y(n_1162) );
OR2x2_ASAP7_75t_L g995 ( .A(n_996), .B(n_1003), .Y(n_995) );
NOR2xp33_ASAP7_75t_L g1021 ( .A(n_996), .B(n_1022), .Y(n_1021) );
AND2x2_ASAP7_75t_L g1027 ( .A(n_996), .B(n_1028), .Y(n_1027) );
NAND2xp5_ASAP7_75t_L g1041 ( .A(n_996), .B(n_1042), .Y(n_1041) );
NAND2xp5_ASAP7_75t_L g1070 ( .A(n_996), .B(n_1071), .Y(n_1070) );
AOI32xp33_ASAP7_75t_L g1120 ( .A1(n_996), .A2(n_1074), .A3(n_1121), .B1(n_1122), .B2(n_1124), .Y(n_1120) );
INVx2_ASAP7_75t_L g1146 ( .A(n_996), .Y(n_1146) );
INVx4_ASAP7_75t_L g996 ( .A(n_997), .Y(n_996) );
NAND2xp5_ASAP7_75t_L g1061 ( .A(n_997), .B(n_1006), .Y(n_1061) );
NOR2xp33_ASAP7_75t_L g1141 ( .A(n_997), .B(n_1088), .Y(n_1141) );
AND2x2_ASAP7_75t_L g1153 ( .A(n_997), .B(n_1075), .Y(n_1153) );
NOR2xp33_ASAP7_75t_L g1155 ( .A(n_997), .B(n_1048), .Y(n_1155) );
AND2x2_ASAP7_75t_L g1161 ( .A(n_997), .B(n_1028), .Y(n_1161) );
AND2x2_ASAP7_75t_L g997 ( .A(n_998), .B(n_1001), .Y(n_997) );
INVx2_ASAP7_75t_L g999 ( .A(n_1000), .Y(n_999) );
INVx1_ASAP7_75t_L g1124 ( .A(n_1003), .Y(n_1124) );
NAND2xp5_ASAP7_75t_L g1004 ( .A(n_1005), .B(n_1012), .Y(n_1004) );
NOR2xp33_ASAP7_75t_L g1035 ( .A(n_1005), .B(n_1036), .Y(n_1035) );
INVx2_ASAP7_75t_L g1005 ( .A(n_1006), .Y(n_1005) );
INVx1_ASAP7_75t_L g1006 ( .A(n_1007), .Y(n_1006) );
INVx1_ASAP7_75t_L g1053 ( .A(n_1007), .Y(n_1053) );
INVx1_ASAP7_75t_L g1007 ( .A(n_1008), .Y(n_1007) );
INVx2_ASAP7_75t_L g1028 ( .A(n_1008), .Y(n_1028) );
INVx4_ASAP7_75t_L g1008 ( .A(n_1009), .Y(n_1008) );
NAND2xp5_ASAP7_75t_L g1165 ( .A(n_1009), .B(n_1096), .Y(n_1165) );
AND2x2_ASAP7_75t_L g1009 ( .A(n_1010), .B(n_1011), .Y(n_1009) );
NAND2xp5_ASAP7_75t_L g1118 ( .A(n_1012), .B(n_1119), .Y(n_1118) );
AND2x2_ASAP7_75t_L g1012 ( .A(n_1013), .B(n_1015), .Y(n_1012) );
AND2x2_ASAP7_75t_L g1037 ( .A(n_1013), .B(n_1038), .Y(n_1037) );
AND2x2_ASAP7_75t_L g1054 ( .A(n_1013), .B(n_1055), .Y(n_1054) );
INVx1_ASAP7_75t_L g1013 ( .A(n_1014), .Y(n_1013) );
NOR2x1_ASAP7_75t_L g1065 ( .A(n_1014), .B(n_1016), .Y(n_1065) );
NAND2xp5_ASAP7_75t_L g1123 ( .A(n_1015), .B(n_1034), .Y(n_1123) );
NOR2x1_ASAP7_75t_L g1057 ( .A(n_1016), .B(n_1047), .Y(n_1057) );
A2O1A1Ixp33_ASAP7_75t_L g1099 ( .A1(n_1016), .A2(n_1022), .B(n_1100), .C(n_1102), .Y(n_1099) );
AOI221xp5_ASAP7_75t_L g1106 ( .A1(n_1016), .A2(n_1082), .B1(n_1107), .B2(n_1112), .C(n_1117), .Y(n_1106) );
NAND2xp5_ASAP7_75t_L g1148 ( .A(n_1016), .B(n_1042), .Y(n_1148) );
INVx3_ASAP7_75t_L g1016 ( .A(n_1017), .Y(n_1016) );
AND2x2_ASAP7_75t_L g1033 ( .A(n_1017), .B(n_1034), .Y(n_1033) );
NAND2xp5_ASAP7_75t_L g1084 ( .A(n_1017), .B(n_1085), .Y(n_1084) );
AND2x2_ASAP7_75t_L g1136 ( .A(n_1017), .B(n_1042), .Y(n_1136) );
NAND2xp5_ASAP7_75t_L g1018 ( .A(n_1019), .B(n_1021), .Y(n_1018) );
NAND2xp5_ASAP7_75t_L g1047 ( .A(n_1019), .B(n_1038), .Y(n_1047) );
INVx1_ASAP7_75t_L g1077 ( .A(n_1019), .Y(n_1077) );
O2A1O1Ixp33_ASAP7_75t_L g1062 ( .A1(n_1020), .A2(n_1063), .B(n_1064), .C(n_1066), .Y(n_1062) );
NAND2xp5_ASAP7_75t_L g1104 ( .A(n_1020), .B(n_1038), .Y(n_1104) );
INVx1_ASAP7_75t_L g1150 ( .A(n_1022), .Y(n_1150) );
AOI21xp33_ASAP7_75t_SL g1171 ( .A1(n_1022), .A2(n_1172), .B(n_1173), .Y(n_1171) );
AOI21xp33_ASAP7_75t_L g1023 ( .A1(n_1024), .A2(n_1026), .B(n_1029), .Y(n_1023) );
INVx1_ASAP7_75t_L g1024 ( .A(n_1025), .Y(n_1024) );
INVx1_ASAP7_75t_L g1026 ( .A(n_1027), .Y(n_1026) );
AOI22xp5_ASAP7_75t_L g1154 ( .A1(n_1027), .A2(n_1046), .B1(n_1057), .B2(n_1155), .Y(n_1154) );
AOI32xp33_ASAP7_75t_L g1137 ( .A1(n_1028), .A2(n_1059), .A3(n_1100), .B1(n_1138), .B2(n_1139), .Y(n_1137) );
NAND2xp5_ASAP7_75t_L g1158 ( .A(n_1028), .B(n_1159), .Y(n_1158) );
NAND2xp5_ASAP7_75t_L g1114 ( .A(n_1029), .B(n_1100), .Y(n_1114) );
INVx1_ASAP7_75t_L g1029 ( .A(n_1030), .Y(n_1029) );
O2A1O1Ixp33_ASAP7_75t_L g1031 ( .A1(n_1032), .A2(n_1035), .B(n_1039), .C(n_1040), .Y(n_1031) );
INVx1_ASAP7_75t_L g1127 ( .A(n_1034), .Y(n_1127) );
NAND2xp5_ASAP7_75t_L g1170 ( .A(n_1034), .B(n_1055), .Y(n_1170) );
INVx1_ASAP7_75t_L g1036 ( .A(n_1037), .Y(n_1036) );
NAND2xp5_ASAP7_75t_L g1064 ( .A(n_1038), .B(n_1065), .Y(n_1064) );
A2O1A1Ixp33_ASAP7_75t_SL g1125 ( .A1(n_1039), .A2(n_1087), .B(n_1126), .C(n_1128), .Y(n_1125) );
OAI221xp5_ASAP7_75t_L g1040 ( .A1(n_1041), .A2(n_1044), .B1(n_1045), .B2(n_1048), .C(n_1049), .Y(n_1040) );
INVx1_ASAP7_75t_L g1042 ( .A(n_1043), .Y(n_1042) );
INVx2_ASAP7_75t_L g1045 ( .A(n_1046), .Y(n_1045) );
NAND2xp5_ASAP7_75t_L g1102 ( .A(n_1046), .B(n_1067), .Y(n_1102) );
INVx1_ASAP7_75t_L g1046 ( .A(n_1047), .Y(n_1046) );
INVx1_ASAP7_75t_L g1075 ( .A(n_1048), .Y(n_1075) );
OAI22xp5_ASAP7_75t_L g1112 ( .A1(n_1048), .A2(n_1113), .B1(n_1115), .B2(n_1116), .Y(n_1112) );
NAND2xp5_ASAP7_75t_L g1049 ( .A(n_1050), .B(n_1054), .Y(n_1049) );
HB1xp67_ASAP7_75t_L g1050 ( .A(n_1051), .Y(n_1050) );
NAND2xp5_ASAP7_75t_L g1108 ( .A(n_1051), .B(n_1109), .Y(n_1108) );
NOR2xp33_ASAP7_75t_L g1122 ( .A(n_1051), .B(n_1123), .Y(n_1122) );
HB1xp67_ASAP7_75t_L g1168 ( .A(n_1051), .Y(n_1168) );
INVx1_ASAP7_75t_L g1051 ( .A(n_1052), .Y(n_1051) );
INVx1_ASAP7_75t_L g1081 ( .A(n_1052), .Y(n_1081) );
INVx1_ASAP7_75t_L g1052 ( .A(n_1053), .Y(n_1052) );
HB1xp67_ASAP7_75t_L g1119 ( .A(n_1053), .Y(n_1119) );
INVx1_ASAP7_75t_L g1172 ( .A(n_1054), .Y(n_1172) );
O2A1O1Ixp33_ASAP7_75t_L g1056 ( .A1(n_1057), .A2(n_1058), .B(n_1060), .C(n_1062), .Y(n_1056) );
INVx1_ASAP7_75t_L g1058 ( .A(n_1059), .Y(n_1058) );
INVx1_ASAP7_75t_L g1060 ( .A(n_1061), .Y(n_1060) );
INVx1_ASAP7_75t_L g1138 ( .A(n_1065), .Y(n_1138) );
INVx1_ASAP7_75t_L g1066 ( .A(n_1067), .Y(n_1066) );
INVx1_ASAP7_75t_L g1068 ( .A(n_1069), .Y(n_1068) );
NOR2xp33_ASAP7_75t_L g1069 ( .A(n_1070), .B(n_1072), .Y(n_1069) );
INVx3_ASAP7_75t_SL g1098 ( .A(n_1071), .Y(n_1098) );
NAND2xp5_ASAP7_75t_L g1116 ( .A(n_1071), .B(n_1087), .Y(n_1116) );
AND2x2_ASAP7_75t_L g1076 ( .A(n_1077), .B(n_1078), .Y(n_1076) );
INVx1_ASAP7_75t_L g1079 ( .A(n_1080), .Y(n_1079) );
NAND2xp5_ASAP7_75t_L g1080 ( .A(n_1081), .B(n_1082), .Y(n_1080) );
HB1xp67_ASAP7_75t_L g1140 ( .A(n_1081), .Y(n_1140) );
INVxp33_ASAP7_75t_SL g1083 ( .A(n_1084), .Y(n_1083) );
OAI211xp5_ASAP7_75t_L g1093 ( .A1(n_1086), .A2(n_1094), .B(n_1106), .C(n_1133), .Y(n_1093) );
INVx2_ASAP7_75t_L g1086 ( .A(n_1087), .Y(n_1086) );
NAND2xp5_ASAP7_75t_L g1145 ( .A(n_1087), .B(n_1146), .Y(n_1145) );
CKINVDCx5p33_ASAP7_75t_R g1087 ( .A(n_1088), .Y(n_1087) );
AND2x2_ASAP7_75t_L g1088 ( .A(n_1089), .B(n_1092), .Y(n_1088) );
INVx1_ASAP7_75t_L g1090 ( .A(n_1091), .Y(n_1090) );
AOI211xp5_ASAP7_75t_L g1094 ( .A1(n_1095), .A2(n_1098), .B(n_1099), .C(n_1103), .Y(n_1094) );
INVx1_ASAP7_75t_L g1111 ( .A(n_1095), .Y(n_1111) );
AOI22xp33_ASAP7_75t_L g1143 ( .A1(n_1095), .A2(n_1144), .B1(n_1147), .B2(n_1150), .Y(n_1143) );
OAI31xp33_ASAP7_75t_L g1151 ( .A1(n_1095), .A2(n_1101), .A3(n_1152), .B(n_1153), .Y(n_1151) );
AND2x2_ASAP7_75t_L g1095 ( .A(n_1096), .B(n_1097), .Y(n_1095) );
AND2x2_ASAP7_75t_L g1131 ( .A(n_1096), .B(n_1132), .Y(n_1131) );
INVx1_ASAP7_75t_L g1149 ( .A(n_1097), .Y(n_1149) );
OAI211xp5_ASAP7_75t_SL g1117 ( .A1(n_1098), .A2(n_1118), .B(n_1120), .C(n_1125), .Y(n_1117) );
INVx1_ASAP7_75t_L g1100 ( .A(n_1101), .Y(n_1100) );
NOR2xp33_ASAP7_75t_L g1103 ( .A(n_1104), .B(n_1105), .Y(n_1103) );
INVx1_ASAP7_75t_L g1121 ( .A(n_1104), .Y(n_1121) );
NAND3xp33_ASAP7_75t_L g1107 ( .A(n_1108), .B(n_1110), .C(n_1111), .Y(n_1107) );
AOI221xp5_ASAP7_75t_L g1156 ( .A1(n_1109), .A2(n_1144), .B1(n_1157), .B2(n_1161), .C(n_1162), .Y(n_1156) );
INVx1_ASAP7_75t_L g1113 ( .A(n_1114), .Y(n_1113) );
INVxp67_ASAP7_75t_SL g1128 ( .A(n_1129), .Y(n_1128) );
NAND2xp5_ASAP7_75t_L g1129 ( .A(n_1130), .B(n_1131), .Y(n_1129) );
A2O1A1Ixp33_ASAP7_75t_SL g1133 ( .A1(n_1134), .A2(n_1136), .B(n_1137), .C(n_1141), .Y(n_1133) );
INVx1_ASAP7_75t_L g1134 ( .A(n_1135), .Y(n_1134) );
NAND2xp5_ASAP7_75t_L g1163 ( .A(n_1135), .B(n_1164), .Y(n_1163) );
HB1xp67_ASAP7_75t_L g1139 ( .A(n_1140), .Y(n_1139) );
NAND5xp2_ASAP7_75t_L g1142 ( .A(n_1143), .B(n_1151), .C(n_1154), .D(n_1156), .E(n_1166), .Y(n_1142) );
INVx1_ASAP7_75t_L g1144 ( .A(n_1145), .Y(n_1144) );
A2O1A1Ixp33_ASAP7_75t_L g1166 ( .A1(n_1146), .A2(n_1167), .B(n_1169), .C(n_1171), .Y(n_1166) );
INVxp67_ASAP7_75t_SL g1157 ( .A(n_1158), .Y(n_1157) );
INVx1_ASAP7_75t_L g1164 ( .A(n_1165), .Y(n_1164) );
HB1xp67_ASAP7_75t_L g1167 ( .A(n_1168), .Y(n_1167) );
INVx1_ASAP7_75t_L g1169 ( .A(n_1170), .Y(n_1169) );
INVx1_ASAP7_75t_L g1173 ( .A(n_1174), .Y(n_1173) );
BUFx2_ASAP7_75t_L g1175 ( .A(n_1176), .Y(n_1175) );
BUFx2_ASAP7_75t_L g1176 ( .A(n_1177), .Y(n_1176) );
INVx2_ASAP7_75t_L g1179 ( .A(n_1180), .Y(n_1179) );
INVx1_ASAP7_75t_SL g1180 ( .A(n_1181), .Y(n_1180) );
INVxp33_ASAP7_75t_SL g1202 ( .A(n_1182), .Y(n_1202) );
NOR2x1_ASAP7_75t_L g1182 ( .A(n_1183), .B(n_1190), .Y(n_1182) );
NAND4xp25_ASAP7_75t_L g1183 ( .A(n_1184), .B(n_1185), .C(n_1186), .D(n_1187), .Y(n_1183) );
NAND4xp25_ASAP7_75t_L g1190 ( .A(n_1191), .B(n_1192), .C(n_1193), .D(n_1194), .Y(n_1190) );
HB1xp67_ASAP7_75t_L g1195 ( .A(n_1196), .Y(n_1195) );
INVxp67_ASAP7_75t_L g1199 ( .A(n_1200), .Y(n_1199) );
INVx1_ASAP7_75t_L g1201 ( .A(n_1202), .Y(n_1201) );
BUFx2_ASAP7_75t_L g1204 ( .A(n_1205), .Y(n_1204) );
HB1xp67_ASAP7_75t_L g1206 ( .A(n_1207), .Y(n_1206) );
endmodule