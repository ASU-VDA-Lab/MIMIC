module fake_jpeg_346_n_430 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_430);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_430;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_15;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_256;
wire n_221;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_14),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_9),
.Y(n_16)
);

BUFx5_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_9),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_14),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

CKINVDCx16_ASAP7_75t_R g24 ( 
.A(n_7),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_9),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_0),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_1),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_14),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_2),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

BUFx12_ASAP7_75t_L g33 ( 
.A(n_11),
.Y(n_33)
);

BUFx24_ASAP7_75t_L g34 ( 
.A(n_1),
.Y(n_34)
);

BUFx12_ASAP7_75t_L g35 ( 
.A(n_9),
.Y(n_35)
);

BUFx12_ASAP7_75t_L g36 ( 
.A(n_0),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_11),
.Y(n_37)
);

BUFx10_ASAP7_75t_L g38 ( 
.A(n_1),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_11),
.Y(n_39)
);

BUFx16f_ASAP7_75t_L g40 ( 
.A(n_6),
.Y(n_40)
);

BUFx5_ASAP7_75t_L g41 ( 
.A(n_2),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_0),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_2),
.Y(n_43)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_10),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_12),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_8),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_5),
.Y(n_47)
);

BUFx12_ASAP7_75t_L g48 ( 
.A(n_40),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g104 ( 
.A(n_48),
.Y(n_104)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_22),
.Y(n_49)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_49),
.Y(n_101)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_17),
.Y(n_50)
);

INVx4_ASAP7_75t_L g119 ( 
.A(n_50),
.Y(n_119)
);

INVx8_ASAP7_75t_L g51 ( 
.A(n_40),
.Y(n_51)
);

INVx5_ASAP7_75t_L g111 ( 
.A(n_51),
.Y(n_111)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_17),
.Y(n_52)
);

INVx4_ASAP7_75t_L g125 ( 
.A(n_52),
.Y(n_125)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

BUFx2_ASAP7_75t_L g141 ( 
.A(n_53),
.Y(n_141)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_22),
.Y(n_54)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_54),
.Y(n_105)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_17),
.Y(n_55)
);

INVx4_ASAP7_75t_L g129 ( 
.A(n_55),
.Y(n_129)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_18),
.Y(n_56)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_56),
.Y(n_112)
);

INVx2_ASAP7_75t_SL g57 ( 
.A(n_34),
.Y(n_57)
);

INVx4_ASAP7_75t_L g153 ( 
.A(n_57),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_20),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_58),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_20),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_59),
.Y(n_108)
);

BUFx12_ASAP7_75t_L g60 ( 
.A(n_40),
.Y(n_60)
);

INVx6_ASAP7_75t_SL g150 ( 
.A(n_60),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_20),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_61),
.Y(n_109)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_18),
.Y(n_62)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_62),
.Y(n_116)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_23),
.Y(n_63)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_63),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_28),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_64),
.Y(n_121)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_41),
.Y(n_65)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_65),
.Y(n_120)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_18),
.Y(n_66)
);

INVx3_ASAP7_75t_L g139 ( 
.A(n_66),
.Y(n_139)
);

BUFx5_ASAP7_75t_L g67 ( 
.A(n_34),
.Y(n_67)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_67),
.Y(n_122)
);

INVx8_ASAP7_75t_L g68 ( 
.A(n_18),
.Y(n_68)
);

INVx6_ASAP7_75t_L g132 ( 
.A(n_68),
.Y(n_132)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_18),
.Y(n_69)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_69),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_28),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_70),
.Y(n_136)
);

INVx6_ASAP7_75t_L g71 ( 
.A(n_28),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g147 ( 
.A(n_71),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_15),
.B(n_13),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_72),
.B(n_98),
.Y(n_115)
);

CKINVDCx14_ASAP7_75t_R g73 ( 
.A(n_34),
.Y(n_73)
);

OR2x2_ASAP7_75t_L g135 ( 
.A(n_73),
.B(n_97),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_39),
.Y(n_74)
);

INVx6_ASAP7_75t_L g134 ( 
.A(n_74),
.Y(n_134)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_32),
.Y(n_75)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_75),
.Y(n_138)
);

INVx6_ASAP7_75t_L g76 ( 
.A(n_39),
.Y(n_76)
);

INVx8_ASAP7_75t_L g127 ( 
.A(n_76),
.Y(n_127)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_32),
.Y(n_77)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_77),
.Y(n_140)
);

BUFx3_ASAP7_75t_L g78 ( 
.A(n_39),
.Y(n_78)
);

INVx6_ASAP7_75t_L g151 ( 
.A(n_78),
.Y(n_151)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_32),
.Y(n_79)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_79),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_SL g80 ( 
.A(n_15),
.B(n_13),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_80),
.B(n_88),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_24),
.B(n_12),
.Y(n_81)
);

OAI21xp33_ASAP7_75t_L g118 ( 
.A1(n_81),
.A2(n_83),
.B(n_3),
.Y(n_118)
);

BUFx5_ASAP7_75t_L g82 ( 
.A(n_34),
.Y(n_82)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_82),
.Y(n_128)
);

NAND2x1_ASAP7_75t_L g83 ( 
.A(n_32),
.B(n_1),
.Y(n_83)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_32),
.Y(n_84)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_84),
.Y(n_131)
);

INVx8_ASAP7_75t_L g85 ( 
.A(n_47),
.Y(n_85)
);

AND2x2_ASAP7_75t_L g148 ( 
.A(n_85),
.B(n_89),
.Y(n_148)
);

INVx2_ASAP7_75t_SL g86 ( 
.A(n_34),
.Y(n_86)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_86),
.Y(n_137)
);

INVx13_ASAP7_75t_L g87 ( 
.A(n_24),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_87),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_SL g88 ( 
.A(n_30),
.B(n_12),
.Y(n_88)
);

INVx2_ASAP7_75t_SL g89 ( 
.A(n_41),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_47),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_90),
.Y(n_110)
);

BUFx3_ASAP7_75t_L g91 ( 
.A(n_47),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_91),
.B(n_93),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_23),
.B(n_2),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_92),
.B(n_95),
.Y(n_143)
);

BUFx12f_ASAP7_75t_L g93 ( 
.A(n_33),
.Y(n_93)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_19),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_94),
.B(n_96),
.Y(n_142)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_44),
.Y(n_95)
);

INVx5_ASAP7_75t_L g96 ( 
.A(n_44),
.Y(n_96)
);

INVx4_ASAP7_75t_SL g97 ( 
.A(n_41),
.Y(n_97)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_19),
.Y(n_98)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_44),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_99),
.B(n_100),
.Y(n_149)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_38),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g103 ( 
.A(n_81),
.B(n_30),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_103),
.B(n_118),
.Y(n_182)
);

AOI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_97),
.A2(n_45),
.B1(n_46),
.B2(n_42),
.Y(n_114)
);

OA22x2_ASAP7_75t_L g157 ( 
.A1(n_114),
.A2(n_152),
.B1(n_86),
.B2(n_73),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_92),
.A2(n_61),
.B1(n_90),
.B2(n_70),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_124),
.A2(n_126),
.B1(n_85),
.B2(n_53),
.Y(n_173)
);

AOI22xp33_ASAP7_75t_L g126 ( 
.A1(n_58),
.A2(n_46),
.B1(n_42),
.B2(n_37),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_83),
.B(n_45),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_130),
.B(n_4),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_89),
.B(n_25),
.C(n_37),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_133),
.B(n_31),
.C(n_27),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_59),
.Y(n_145)
);

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_145),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_64),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_146),
.B(n_154),
.Y(n_174)
);

AOI22xp33_ASAP7_75t_SL g152 ( 
.A1(n_57),
.A2(n_25),
.B1(n_43),
.B2(n_26),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_74),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_51),
.B(n_43),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_155),
.B(n_93),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_150),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_156),
.B(n_161),
.Y(n_203)
);

CKINVDCx16_ASAP7_75t_R g213 ( 
.A(n_157),
.Y(n_213)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_147),
.Y(n_159)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_159),
.Y(n_200)
);

BUFx3_ASAP7_75t_L g160 ( 
.A(n_111),
.Y(n_160)
);

BUFx3_ASAP7_75t_L g228 ( 
.A(n_160),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_142),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_141),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_162),
.B(n_172),
.Y(n_205)
);

AOI22xp33_ASAP7_75t_SL g163 ( 
.A1(n_148),
.A2(n_29),
.B1(n_16),
.B2(n_21),
.Y(n_163)
);

INVxp67_ASAP7_75t_SL g211 ( 
.A(n_163),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_143),
.A2(n_29),
.B1(n_16),
.B2(n_21),
.Y(n_164)
);

CKINVDCx16_ASAP7_75t_R g222 ( 
.A(n_164),
.Y(n_222)
);

AND2x2_ASAP7_75t_L g229 ( 
.A(n_165),
.B(n_173),
.Y(n_229)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_153),
.Y(n_166)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_166),
.Y(n_215)
);

AOI22xp33_ASAP7_75t_L g167 ( 
.A1(n_115),
.A2(n_31),
.B1(n_27),
.B2(n_26),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_167),
.A2(n_187),
.B1(n_152),
.B2(n_114),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_118),
.B(n_3),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_168),
.B(n_176),
.Y(n_201)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_153),
.Y(n_169)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_169),
.Y(n_220)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_147),
.Y(n_170)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_170),
.Y(n_202)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_137),
.Y(n_171)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_171),
.Y(n_223)
);

INVxp67_ASAP7_75t_L g172 ( 
.A(n_135),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_175),
.B(n_186),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_117),
.B(n_3),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_101),
.Y(n_177)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_177),
.Y(n_216)
);

INVx5_ASAP7_75t_L g178 ( 
.A(n_111),
.Y(n_178)
);

INVx4_ASAP7_75t_L g219 ( 
.A(n_178),
.Y(n_219)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_148),
.Y(n_179)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_179),
.Y(n_218)
);

INVx3_ASAP7_75t_SL g180 ( 
.A(n_127),
.Y(n_180)
);

INVx11_ASAP7_75t_L g217 ( 
.A(n_180),
.Y(n_217)
);

HB1xp67_ASAP7_75t_L g181 ( 
.A(n_139),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_181),
.Y(n_198)
);

AOI22xp33_ASAP7_75t_SL g183 ( 
.A1(n_110),
.A2(n_87),
.B1(n_38),
.B2(n_33),
.Y(n_183)
);

OAI22xp33_ASAP7_75t_L g206 ( 
.A1(n_183),
.A2(n_197),
.B1(n_180),
.B2(n_156),
.Y(n_206)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_134),
.Y(n_184)
);

INVx3_ASAP7_75t_L g208 ( 
.A(n_184),
.Y(n_208)
);

INVx5_ASAP7_75t_L g185 ( 
.A(n_104),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_185),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_126),
.A2(n_38),
.B1(n_48),
.B2(n_60),
.Y(n_187)
);

CKINVDCx16_ASAP7_75t_R g188 ( 
.A(n_135),
.Y(n_188)
);

INVx13_ASAP7_75t_L g207 ( 
.A(n_188),
.Y(n_207)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_131),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_189),
.B(n_191),
.Y(n_225)
);

INVx5_ASAP7_75t_L g190 ( 
.A(n_104),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_190),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_141),
.Y(n_191)
);

INVx8_ASAP7_75t_L g192 ( 
.A(n_104),
.Y(n_192)
);

BUFx12f_ASAP7_75t_L g221 ( 
.A(n_192),
.Y(n_221)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_149),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_193),
.B(n_194),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_105),
.B(n_4),
.Y(n_194)
);

INVx1_ASAP7_75t_SL g195 ( 
.A(n_128),
.Y(n_195)
);

INVx8_ASAP7_75t_L g212 ( 
.A(n_195),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_106),
.B(n_4),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_196),
.B(n_107),
.C(n_122),
.Y(n_199)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_134),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_199),
.B(n_195),
.Y(n_246)
);

AND2x2_ASAP7_75t_L g250 ( 
.A(n_204),
.B(n_158),
.Y(n_250)
);

INVx1_ASAP7_75t_SL g231 ( 
.A(n_206),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_164),
.A2(n_127),
.B1(n_136),
.B2(n_121),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_209),
.A2(n_187),
.B1(n_191),
.B2(n_162),
.Y(n_242)
);

AOI21xp5_ASAP7_75t_L g224 ( 
.A1(n_172),
.A2(n_157),
.B(n_168),
.Y(n_224)
);

INVxp67_ASAP7_75t_L g237 ( 
.A(n_224),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_213),
.A2(n_179),
.B1(n_173),
.B2(n_193),
.Y(n_230)
);

AO22x1_ASAP7_75t_SL g259 ( 
.A1(n_230),
.A2(n_232),
.B1(n_235),
.B2(n_204),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_213),
.A2(n_176),
.B1(n_182),
.B2(n_194),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_227),
.B(n_177),
.C(n_189),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_233),
.B(n_240),
.C(n_249),
.Y(n_255)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_216),
.Y(n_234)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_234),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_224),
.A2(n_157),
.B1(n_174),
.B2(n_136),
.Y(n_235)
);

AOI22xp33_ASAP7_75t_L g236 ( 
.A1(n_211),
.A2(n_180),
.B1(n_171),
.B2(n_157),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_L g258 ( 
.A1(n_236),
.A2(n_242),
.B1(n_217),
.B2(n_231),
.Y(n_258)
);

OR2x6_ASAP7_75t_L g238 ( 
.A(n_199),
.B(n_165),
.Y(n_238)
);

AOI21xp5_ASAP7_75t_SL g263 ( 
.A1(n_238),
.A2(n_207),
.B(n_113),
.Y(n_263)
);

OAI22x1_ASAP7_75t_L g239 ( 
.A1(n_229),
.A2(n_158),
.B1(n_190),
.B2(n_185),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_239),
.B(n_252),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_227),
.B(n_140),
.C(n_116),
.Y(n_240)
);

INVxp67_ASAP7_75t_L g241 ( 
.A(n_205),
.Y(n_241)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_241),
.Y(n_264)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_216),
.Y(n_243)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_243),
.Y(n_275)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_223),
.Y(n_244)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_244),
.Y(n_278)
);

INVx4_ASAP7_75t_L g245 ( 
.A(n_219),
.Y(n_245)
);

INVx3_ASAP7_75t_L g269 ( 
.A(n_245),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_SL g266 ( 
.A(n_246),
.B(n_254),
.Y(n_266)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_200),
.Y(n_247)
);

AND2x2_ASAP7_75t_L g270 ( 
.A(n_247),
.B(n_250),
.Y(n_270)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_223),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_SL g271 ( 
.A(n_248),
.B(n_253),
.Y(n_271)
);

MAJx2_ASAP7_75t_L g249 ( 
.A(n_229),
.B(n_169),
.C(n_166),
.Y(n_249)
);

INVxp67_ASAP7_75t_L g251 ( 
.A(n_225),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_251),
.Y(n_268)
);

INVxp33_ASAP7_75t_L g252 ( 
.A(n_225),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_215),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_203),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_237),
.A2(n_229),
.B1(n_222),
.B2(n_201),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_256),
.A2(n_265),
.B1(n_230),
.B2(n_235),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_258),
.A2(n_260),
.B1(n_261),
.B2(n_208),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_259),
.B(n_109),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_L g260 ( 
.A1(n_231),
.A2(n_222),
.B1(n_201),
.B2(n_218),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_L g261 ( 
.A1(n_241),
.A2(n_218),
.B1(n_209),
.B2(n_226),
.Y(n_261)
);

OAI21xp5_ASAP7_75t_SL g262 ( 
.A1(n_237),
.A2(n_207),
.B(n_198),
.Y(n_262)
);

AOI21xp5_ASAP7_75t_SL g288 ( 
.A1(n_262),
.A2(n_238),
.B(n_214),
.Y(n_288)
);

XOR2xp5_ASAP7_75t_L g283 ( 
.A(n_263),
.B(n_239),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_250),
.A2(n_206),
.B1(n_170),
.B2(n_159),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_249),
.B(n_220),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_272),
.B(n_273),
.C(n_276),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_233),
.B(n_198),
.C(n_220),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_251),
.B(n_215),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_274),
.B(n_252),
.Y(n_281)
);

XOR2xp5_ASAP7_75t_L g276 ( 
.A(n_240),
.B(n_144),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_238),
.B(n_112),
.C(n_138),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_277),
.B(n_250),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_L g320 ( 
.A1(n_279),
.A2(n_285),
.B1(n_290),
.B2(n_300),
.Y(n_320)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_278),
.Y(n_280)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_280),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_281),
.B(n_286),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_SL g282 ( 
.A(n_266),
.B(n_232),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_SL g315 ( 
.A(n_282),
.B(n_257),
.Y(n_315)
);

OR2x2_ASAP7_75t_L g319 ( 
.A(n_283),
.B(n_269),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_L g302 ( 
.A(n_284),
.B(n_276),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_268),
.A2(n_242),
.B1(n_238),
.B2(n_243),
.Y(n_285)
);

INVxp67_ASAP7_75t_L g286 ( 
.A(n_262),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_278),
.Y(n_287)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_287),
.Y(n_316)
);

AOI21xp5_ASAP7_75t_L g317 ( 
.A1(n_288),
.A2(n_275),
.B(n_257),
.Y(n_317)
);

OAI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_259),
.A2(n_238),
.B1(n_245),
.B2(n_214),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_289),
.A2(n_301),
.B1(n_267),
.B2(n_272),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_268),
.A2(n_210),
.B1(n_247),
.B2(n_219),
.Y(n_290)
);

INVxp67_ASAP7_75t_L g292 ( 
.A(n_270),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_292),
.B(n_293),
.Y(n_309)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_271),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_SL g294 ( 
.A1(n_259),
.A2(n_210),
.B1(n_184),
.B2(n_197),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_L g324 ( 
.A1(n_294),
.A2(n_121),
.B1(n_108),
.B2(n_109),
.Y(n_324)
);

A2O1A1O1Ixp25_ASAP7_75t_L g295 ( 
.A1(n_277),
.A2(n_123),
.B(n_202),
.C(n_200),
.D(n_212),
.Y(n_295)
);

FAx1_ASAP7_75t_SL g304 ( 
.A(n_295),
.B(n_273),
.CI(n_265),
.CON(n_304),
.SN(n_304)
);

XOR2xp5_ASAP7_75t_L g296 ( 
.A(n_255),
.B(n_202),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_296),
.B(n_139),
.C(n_120),
.Y(n_323)
);

CKINVDCx16_ASAP7_75t_R g297 ( 
.A(n_274),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_297),
.B(n_298),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g298 ( 
.A(n_270),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_264),
.B(n_208),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_299),
.B(n_269),
.Y(n_321)
);

XNOR2xp5_ASAP7_75t_SL g340 ( 
.A(n_302),
.B(n_318),
.Y(n_340)
);

AOI22xp5_ASAP7_75t_SL g303 ( 
.A1(n_286),
.A2(n_267),
.B1(n_270),
.B2(n_256),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_SL g346 ( 
.A1(n_303),
.A2(n_221),
.B1(n_151),
.B2(n_129),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_304),
.B(n_307),
.Y(n_328)
);

OAI22xp5_ASAP7_75t_L g336 ( 
.A1(n_305),
.A2(n_315),
.B1(n_324),
.B2(n_290),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_291),
.B(n_266),
.Y(n_307)
);

XOR2xp5_ASAP7_75t_L g308 ( 
.A(n_296),
.B(n_255),
.Y(n_308)
);

XOR2xp5_ASAP7_75t_L g331 ( 
.A(n_308),
.B(n_312),
.Y(n_331)
);

XNOR2xp5_ASAP7_75t_L g312 ( 
.A(n_291),
.B(n_263),
.Y(n_312)
);

HB1xp67_ASAP7_75t_L g313 ( 
.A(n_285),
.Y(n_313)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_313),
.Y(n_330)
);

XNOR2xp5_ASAP7_75t_L g314 ( 
.A(n_284),
.B(n_264),
.Y(n_314)
);

XOR2xp5_ASAP7_75t_L g337 ( 
.A(n_314),
.B(n_322),
.Y(n_337)
);

OAI21xp5_ASAP7_75t_L g335 ( 
.A1(n_317),
.A2(n_295),
.B(n_301),
.Y(n_335)
);

XNOR2xp5_ASAP7_75t_SL g318 ( 
.A(n_289),
.B(n_275),
.Y(n_318)
);

NAND2xp33_ASAP7_75t_SL g326 ( 
.A(n_319),
.B(n_294),
.Y(n_326)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_321),
.Y(n_332)
);

XOR2xp5_ASAP7_75t_L g322 ( 
.A(n_288),
.B(n_212),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_323),
.B(n_283),
.C(n_292),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g354 ( 
.A(n_325),
.B(n_329),
.C(n_341),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_326),
.B(n_346),
.Y(n_347)
);

XNOR2xp5_ASAP7_75t_L g327 ( 
.A(n_312),
.B(n_308),
.Y(n_327)
);

XOR2xp5_ASAP7_75t_L g352 ( 
.A(n_327),
.B(n_334),
.Y(n_352)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_302),
.B(n_279),
.C(n_281),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_309),
.B(n_299),
.Y(n_333)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_333),
.Y(n_348)
);

XNOR2xp5_ASAP7_75t_L g334 ( 
.A(n_314),
.B(n_300),
.Y(n_334)
);

AOI21xp5_ASAP7_75t_L g365 ( 
.A1(n_335),
.A2(n_132),
.B(n_38),
.Y(n_365)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_336),
.Y(n_349)
);

OAI22xp5_ASAP7_75t_L g338 ( 
.A1(n_320),
.A2(n_228),
.B1(n_217),
.B2(n_221),
.Y(n_338)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_338),
.Y(n_355)
);

AOI22xp5_ASAP7_75t_L g339 ( 
.A1(n_310),
.A2(n_228),
.B1(n_178),
.B2(n_108),
.Y(n_339)
);

INVxp67_ASAP7_75t_SL g358 ( 
.A(n_339),
.Y(n_358)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_323),
.B(n_160),
.C(n_120),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_311),
.B(n_221),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_SL g357 ( 
.A(n_342),
.B(n_316),
.Y(n_357)
);

XOR2xp5_ASAP7_75t_L g343 ( 
.A(n_303),
.B(n_192),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g356 ( 
.A(n_343),
.B(n_344),
.C(n_345),
.Y(n_356)
);

MAJIxp5_ASAP7_75t_L g344 ( 
.A(n_319),
.B(n_125),
.C(n_119),
.Y(n_344)
);

MAJIxp5_ASAP7_75t_L g345 ( 
.A(n_322),
.B(n_125),
.C(n_119),
.Y(n_345)
);

INVx2_ASAP7_75t_L g350 ( 
.A(n_332),
.Y(n_350)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_350),
.Y(n_376)
);

XNOR2x2_ASAP7_75t_L g351 ( 
.A(n_340),
.B(n_306),
.Y(n_351)
);

XNOR2xp5_ASAP7_75t_SL g373 ( 
.A(n_351),
.B(n_36),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_330),
.B(n_317),
.Y(n_353)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_353),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_357),
.Y(n_378)
);

CKINVDCx20_ASAP7_75t_R g359 ( 
.A(n_335),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_SL g379 ( 
.A(n_359),
.B(n_360),
.Y(n_379)
);

MAJIxp5_ASAP7_75t_L g360 ( 
.A(n_331),
.B(n_318),
.C(n_305),
.Y(n_360)
);

OAI22xp5_ASAP7_75t_SL g361 ( 
.A1(n_328),
.A2(n_304),
.B1(n_324),
.B2(n_221),
.Y(n_361)
);

AOI22xp5_ASAP7_75t_L g371 ( 
.A1(n_361),
.A2(n_362),
.B1(n_337),
.B2(n_36),
.Y(n_371)
);

OAI22xp5_ASAP7_75t_SL g362 ( 
.A1(n_334),
.A2(n_304),
.B1(n_102),
.B2(n_151),
.Y(n_362)
);

MAJIxp5_ASAP7_75t_L g363 ( 
.A(n_331),
.B(n_129),
.C(n_102),
.Y(n_363)
);

MAJIxp5_ASAP7_75t_L g367 ( 
.A(n_363),
.B(n_364),
.C(n_340),
.Y(n_367)
);

MAJIxp5_ASAP7_75t_L g364 ( 
.A(n_327),
.B(n_132),
.C(n_38),
.Y(n_364)
);

XOR2xp5_ASAP7_75t_L g372 ( 
.A(n_365),
.B(n_5),
.Y(n_372)
);

OAI22xp5_ASAP7_75t_L g366 ( 
.A1(n_348),
.A2(n_329),
.B1(n_343),
.B2(n_344),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_366),
.B(n_369),
.Y(n_382)
);

XOR2xp5_ASAP7_75t_L g390 ( 
.A(n_367),
.B(n_372),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_350),
.B(n_341),
.Y(n_368)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_368),
.Y(n_384)
);

OAI22xp5_ASAP7_75t_L g369 ( 
.A1(n_349),
.A2(n_345),
.B1(n_325),
.B2(n_337),
.Y(n_369)
);

HB1xp67_ASAP7_75t_L g370 ( 
.A(n_355),
.Y(n_370)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_370),
.Y(n_385)
);

HB1xp67_ASAP7_75t_L g389 ( 
.A(n_371),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_373),
.B(n_375),
.Y(n_391)
);

XOR2xp5_ASAP7_75t_L g374 ( 
.A(n_352),
.B(n_354),
.Y(n_374)
);

NOR2xp33_ASAP7_75t_L g394 ( 
.A(n_374),
.B(n_380),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_353),
.B(n_5),
.Y(n_375)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_358),
.Y(n_380)
);

MAJIxp5_ASAP7_75t_L g381 ( 
.A(n_354),
.B(n_352),
.C(n_360),
.Y(n_381)
);

MAJIxp5_ASAP7_75t_L g387 ( 
.A(n_381),
.B(n_356),
.C(n_364),
.Y(n_387)
);

AOI21xp5_ASAP7_75t_L g383 ( 
.A1(n_379),
.A2(n_361),
.B(n_363),
.Y(n_383)
);

AOI21xp5_ASAP7_75t_L g396 ( 
.A1(n_383),
.A2(n_386),
.B(n_393),
.Y(n_396)
);

AOI21xp5_ASAP7_75t_L g386 ( 
.A1(n_377),
.A2(n_356),
.B(n_362),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_387),
.B(n_388),
.Y(n_402)
);

MAJIxp5_ASAP7_75t_L g388 ( 
.A(n_374),
.B(n_351),
.C(n_347),
.Y(n_388)
);

AOI22xp5_ASAP7_75t_SL g392 ( 
.A1(n_368),
.A2(n_347),
.B1(n_365),
.B2(n_8),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_392),
.B(n_395),
.Y(n_405)
);

AOI21xp5_ASAP7_75t_SL g393 ( 
.A1(n_376),
.A2(n_6),
.B(n_7),
.Y(n_393)
);

MAJIxp5_ASAP7_75t_L g395 ( 
.A(n_381),
.B(n_33),
.C(n_35),
.Y(n_395)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_393),
.Y(n_397)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_397),
.Y(n_411)
);

NOR2x1_ASAP7_75t_SL g398 ( 
.A(n_388),
.B(n_378),
.Y(n_398)
);

AOI21xp5_ASAP7_75t_L g410 ( 
.A1(n_398),
.A2(n_7),
.B(n_8),
.Y(n_410)
);

OAI22xp5_ASAP7_75t_SL g399 ( 
.A1(n_389),
.A2(n_371),
.B1(n_373),
.B2(n_375),
.Y(n_399)
);

NOR2xp33_ASAP7_75t_L g413 ( 
.A(n_399),
.B(n_400),
.Y(n_413)
);

MAJIxp5_ASAP7_75t_L g400 ( 
.A(n_387),
.B(n_367),
.C(n_372),
.Y(n_400)
);

XOR2xp5_ASAP7_75t_L g401 ( 
.A(n_390),
.B(n_394),
.Y(n_401)
);

XNOR2xp5_ASAP7_75t_L g407 ( 
.A(n_401),
.B(n_403),
.Y(n_407)
);

XOR2xp5_ASAP7_75t_L g403 ( 
.A(n_390),
.B(n_33),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_385),
.Y(n_404)
);

NOR2xp33_ASAP7_75t_SL g412 ( 
.A(n_404),
.B(n_8),
.Y(n_412)
);

XOR2xp5_ASAP7_75t_L g406 ( 
.A(n_384),
.B(n_382),
.Y(n_406)
);

MAJIxp5_ASAP7_75t_L g408 ( 
.A(n_406),
.B(n_395),
.C(n_391),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_408),
.B(n_409),
.Y(n_416)
);

NOR2xp67_ASAP7_75t_L g409 ( 
.A(n_402),
.B(n_35),
.Y(n_409)
);

XNOR2xp5_ASAP7_75t_L g420 ( 
.A(n_410),
.B(n_403),
.Y(n_420)
);

NOR2xp33_ASAP7_75t_L g415 ( 
.A(n_412),
.B(n_10),
.Y(n_415)
);

NOR2xp33_ASAP7_75t_SL g414 ( 
.A(n_401),
.B(n_10),
.Y(n_414)
);

NOR2xp33_ASAP7_75t_SL g418 ( 
.A(n_414),
.B(n_399),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_415),
.B(n_417),
.Y(n_424)
);

NAND4xp25_ASAP7_75t_SL g417 ( 
.A(n_413),
.B(n_405),
.C(n_406),
.D(n_396),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_SL g421 ( 
.A(n_418),
.B(n_419),
.Y(n_421)
);

INVxp67_ASAP7_75t_L g419 ( 
.A(n_413),
.Y(n_419)
);

XOR2xp5_ASAP7_75t_L g422 ( 
.A(n_420),
.B(n_407),
.Y(n_422)
);

INVxp33_ASAP7_75t_SL g425 ( 
.A(n_422),
.Y(n_425)
);

AOI21xp5_ASAP7_75t_L g423 ( 
.A1(n_416),
.A2(n_411),
.B(n_400),
.Y(n_423)
);

AOI21xp5_ASAP7_75t_SL g426 ( 
.A1(n_423),
.A2(n_35),
.B(n_36),
.Y(n_426)
);

AOI22xp5_ASAP7_75t_L g427 ( 
.A1(n_426),
.A2(n_424),
.B1(n_421),
.B2(n_35),
.Y(n_427)
);

A2O1A1Ixp33_ASAP7_75t_SL g428 ( 
.A1(n_427),
.A2(n_425),
.B(n_11),
.C(n_10),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_428),
.Y(n_429)
);

XOR2xp5_ASAP7_75t_L g430 ( 
.A(n_429),
.B(n_36),
.Y(n_430)
);


endmodule