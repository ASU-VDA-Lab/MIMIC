module fake_jpeg_12544_n_173 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_173);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_173;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_96;

INVx2_ASAP7_75t_L g15 ( 
.A(n_4),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_1),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_5),
.B(n_8),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_4),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_0),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_0),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

INVx13_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_7),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_6),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_32),
.B(n_9),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_SL g69 ( 
.A(n_34),
.B(n_43),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_33),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_35),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_33),
.Y(n_36)
);

INVx5_ASAP7_75t_L g71 ( 
.A(n_36),
.Y(n_71)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_18),
.Y(n_37)
);

INVx1_ASAP7_75t_SL g57 ( 
.A(n_37),
.Y(n_57)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_19),
.Y(n_38)
);

INVx5_ASAP7_75t_L g64 ( 
.A(n_38),
.Y(n_64)
);

INVx5_ASAP7_75t_L g39 ( 
.A(n_33),
.Y(n_39)
);

BUFx2_ASAP7_75t_L g66 ( 
.A(n_39),
.Y(n_66)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_19),
.Y(n_40)
);

INVx5_ASAP7_75t_L g67 ( 
.A(n_40),
.Y(n_67)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_33),
.Y(n_41)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_41),
.Y(n_55)
);

BUFx5_ASAP7_75t_L g42 ( 
.A(n_19),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_42),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_SL g43 ( 
.A(n_21),
.B(n_9),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_32),
.B(n_13),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_44),
.B(n_47),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_26),
.Y(n_45)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_45),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_26),
.Y(n_46)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_46),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_17),
.B(n_1),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_47),
.B(n_15),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_49),
.B(n_28),
.Y(n_74)
);

OR2x2_ASAP7_75t_L g52 ( 
.A(n_43),
.B(n_31),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_52),
.B(n_53),
.Y(n_72)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_41),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_37),
.B(n_31),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_54),
.B(n_56),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_37),
.B(n_27),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_37),
.B(n_27),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_59),
.B(n_61),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g60 ( 
.A1(n_45),
.A2(n_15),
.B1(n_26),
.B2(n_16),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_60),
.A2(n_29),
.B1(n_20),
.B2(n_17),
.Y(n_94)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_38),
.Y(n_61)
);

INVxp67_ASAP7_75t_L g62 ( 
.A(n_40),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_62),
.B(n_70),
.Y(n_84)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_45),
.Y(n_65)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_65),
.Y(n_82)
);

INVx5_ASAP7_75t_SL g68 ( 
.A(n_39),
.Y(n_68)
);

OR2x2_ASAP7_75t_L g75 ( 
.A(n_68),
.B(n_36),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_35),
.B(n_23),
.Y(n_70)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_63),
.Y(n_73)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_73),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_74),
.B(n_85),
.Y(n_99)
);

INVx1_ASAP7_75t_SL g111 ( 
.A(n_75),
.Y(n_111)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_49),
.B(n_46),
.Y(n_77)
);

INVxp67_ASAP7_75t_SL g97 ( 
.A(n_77),
.Y(n_97)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_55),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_L g79 ( 
.A1(n_60),
.A2(n_46),
.B1(n_28),
.B2(n_25),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_79),
.A2(n_24),
.B1(n_67),
.B2(n_18),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_55),
.B(n_57),
.C(n_48),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_80),
.B(n_90),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_52),
.B(n_20),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_81),
.B(n_2),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_69),
.B(n_22),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_66),
.B(n_22),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_86),
.B(n_89),
.Y(n_104)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_50),
.Y(n_87)
);

HB1xp67_ASAP7_75t_L g98 ( 
.A(n_87),
.Y(n_98)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_50),
.Y(n_88)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_88),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_66),
.B(n_23),
.Y(n_89)
);

OR2x2_ASAP7_75t_L g90 ( 
.A(n_68),
.B(n_29),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_57),
.B(n_25),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_91),
.B(n_93),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_63),
.Y(n_92)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_92),
.Y(n_100)
);

NOR2x1_ASAP7_75t_L g93 ( 
.A(n_65),
.B(n_16),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_94),
.A2(n_24),
.B1(n_62),
.B2(n_64),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_64),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_95),
.B(n_67),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_101),
.A2(n_110),
.B1(n_113),
.B2(n_71),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_103),
.A2(n_114),
.B1(n_81),
.B2(n_95),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_105),
.B(n_109),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_90),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_106),
.B(n_112),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_94),
.A2(n_71),
.B1(n_58),
.B2(n_51),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_90),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_L g113 ( 
.A1(n_77),
.A2(n_58),
.B1(n_51),
.B2(n_30),
.Y(n_113)
);

OAI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_93),
.A2(n_75),
.B1(n_80),
.B2(n_74),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_SL g115 ( 
.A(n_99),
.B(n_72),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_115),
.B(n_120),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_97),
.B(n_77),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_117),
.B(n_123),
.Y(n_134)
);

AOI21xp5_ASAP7_75t_L g119 ( 
.A1(n_111),
.A2(n_75),
.B(n_93),
.Y(n_119)
);

AOI21xp5_ASAP7_75t_L g135 ( 
.A1(n_119),
.A2(n_107),
.B(n_110),
.Y(n_135)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_108),
.Y(n_120)
);

INVxp67_ASAP7_75t_L g136 ( 
.A(n_121),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_L g122 ( 
.A(n_96),
.B(n_76),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_122),
.B(n_129),
.C(n_82),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_96),
.B(n_83),
.Y(n_123)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_108),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_124),
.B(n_127),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_125),
.A2(n_112),
.B1(n_103),
.B2(n_101),
.Y(n_131)
);

AND2x2_ASAP7_75t_L g126 ( 
.A(n_111),
.B(n_84),
.Y(n_126)
);

XNOR2xp5_ASAP7_75t_L g132 ( 
.A(n_126),
.B(n_128),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_104),
.B(n_78),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_106),
.B(n_88),
.Y(n_128)
);

XOR2xp5_ASAP7_75t_L g129 ( 
.A(n_105),
.B(n_87),
.Y(n_129)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_98),
.Y(n_130)
);

CKINVDCx16_ASAP7_75t_R g138 ( 
.A(n_130),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_131),
.A2(n_139),
.B1(n_130),
.B2(n_102),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_128),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_133),
.B(n_92),
.Y(n_152)
);

NAND3xp33_ASAP7_75t_L g143 ( 
.A(n_135),
.B(n_119),
.C(n_116),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_L g137 ( 
.A(n_122),
.B(n_82),
.Y(n_137)
);

XOR2xp5_ASAP7_75t_L g148 ( 
.A(n_137),
.B(n_142),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_121),
.A2(n_102),
.B1(n_100),
.B2(n_73),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_L g156 ( 
.A(n_143),
.B(n_145),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_140),
.B(n_118),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_SL g154 ( 
.A(n_144),
.B(n_146),
.Y(n_154)
);

A2O1A1O1Ixp25_ASAP7_75t_L g145 ( 
.A1(n_134),
.A2(n_123),
.B(n_117),
.C(n_126),
.D(n_125),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_134),
.B(n_129),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_141),
.B(n_126),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_SL g155 ( 
.A(n_147),
.B(n_149),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_138),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_150),
.B(n_151),
.C(n_152),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_137),
.B(n_100),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_148),
.B(n_132),
.C(n_131),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_157),
.B(n_158),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_145),
.B(n_143),
.C(n_136),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_153),
.A2(n_136),
.B1(n_139),
.B2(n_42),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_159),
.A2(n_161),
.B1(n_3),
.B2(n_6),
.Y(n_165)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_155),
.Y(n_160)
);

AND2x2_ASAP7_75t_L g166 ( 
.A(n_160),
.B(n_162),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_156),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_154),
.A2(n_10),
.B1(n_12),
.B2(n_4),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_L g164 ( 
.A(n_163),
.B(n_2),
.Y(n_164)
);

AND2x2_ASAP7_75t_L g168 ( 
.A(n_164),
.B(n_166),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_165),
.A2(n_161),
.B1(n_162),
.B2(n_121),
.Y(n_167)
);

INVxp67_ASAP7_75t_L g169 ( 
.A(n_167),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_SL g170 ( 
.A(n_168),
.B(n_165),
.Y(n_170)
);

INVxp67_ASAP7_75t_L g171 ( 
.A(n_170),
.Y(n_171)
);

CKINVDCx16_ASAP7_75t_R g172 ( 
.A(n_171),
.Y(n_172)
);

XOR2xp5_ASAP7_75t_L g173 ( 
.A(n_172),
.B(n_169),
.Y(n_173)
);


endmodule