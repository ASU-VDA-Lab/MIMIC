module fake_jpeg_24756_n_337 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_337);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_337;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

INVxp67_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

INVx6_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_9),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_8),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_8),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_15),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_16),
.Y(n_29)
);

CKINVDCx16_ASAP7_75t_R g30 ( 
.A(n_5),
.Y(n_30)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

INVx11_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_10),
.Y(n_34)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_6),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_24),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_36),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_24),
.Y(n_37)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_37),
.Y(n_66)
);

INVx5_ASAP7_75t_L g38 ( 
.A(n_19),
.Y(n_38)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_38),
.A2(n_32),
.B1(n_19),
.B2(n_35),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_23),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_39),
.B(n_44),
.Y(n_48)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_31),
.Y(n_40)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_40),
.Y(n_68)
);

INVx2_ASAP7_75t_R g41 ( 
.A(n_24),
.Y(n_41)
);

OAI21xp33_ASAP7_75t_L g56 ( 
.A1(n_41),
.A2(n_32),
.B(n_36),
.Y(n_56)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_31),
.Y(n_42)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_42),
.Y(n_47)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_43),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_23),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_22),
.B(n_0),
.Y(n_45)
);

AND2x2_ASAP7_75t_L g62 ( 
.A(n_45),
.B(n_0),
.Y(n_62)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_24),
.Y(n_46)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_46),
.Y(n_60)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_45),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_50),
.B(n_64),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_45),
.B(n_22),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_51),
.B(n_62),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_L g52 ( 
.A1(n_38),
.A2(n_19),
.B1(n_31),
.B2(n_35),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_52),
.A2(n_65),
.B1(n_42),
.B2(n_40),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_36),
.Y(n_53)
);

BUFx2_ASAP7_75t_SL g89 ( 
.A(n_53),
.Y(n_89)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_36),
.Y(n_54)
);

INVx3_ASAP7_75t_SL g76 ( 
.A(n_54),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_55),
.A2(n_59),
.B1(n_61),
.B2(n_30),
.Y(n_95)
);

OAI21xp5_ASAP7_75t_SL g99 ( 
.A1(n_56),
.A2(n_40),
.B(n_28),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_39),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_SL g73 ( 
.A(n_57),
.B(n_63),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_L g58 ( 
.A1(n_38),
.A2(n_19),
.B1(n_31),
.B2(n_35),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_L g90 ( 
.A1(n_58),
.A2(n_43),
.B1(n_25),
.B2(n_68),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_41),
.A2(n_32),
.B1(n_35),
.B2(n_30),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_41),
.A2(n_30),
.B1(n_17),
.B2(n_27),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_39),
.B(n_17),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_44),
.B(n_17),
.Y(n_64)
);

OAI22xp33_ASAP7_75t_L g65 ( 
.A1(n_41),
.A2(n_25),
.B1(n_33),
.B2(n_34),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_44),
.B(n_22),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_67),
.B(n_26),
.Y(n_94)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_36),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_69),
.B(n_42),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_70),
.Y(n_74)
);

INVx4_ASAP7_75t_L g112 ( 
.A(n_74),
.Y(n_112)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_70),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_75),
.B(n_78),
.Y(n_103)
);

BUFx3_ASAP7_75t_L g77 ( 
.A(n_70),
.Y(n_77)
);

INVx4_ASAP7_75t_L g117 ( 
.A(n_77),
.Y(n_117)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_47),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_51),
.B(n_27),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_79),
.B(n_85),
.Y(n_104)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_67),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_80),
.B(n_84),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g81 ( 
.A(n_50),
.B(n_36),
.C(n_46),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_81),
.B(n_83),
.C(n_99),
.Y(n_115)
);

AOI21xp33_ASAP7_75t_L g82 ( 
.A1(n_62),
.A2(n_46),
.B(n_26),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_82),
.A2(n_88),
.B1(n_52),
.B2(n_47),
.Y(n_107)
);

OAI21xp5_ASAP7_75t_L g83 ( 
.A1(n_62),
.A2(n_18),
.B(n_46),
.Y(n_83)
);

INVx13_ASAP7_75t_L g84 ( 
.A(n_60),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_62),
.B(n_27),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_48),
.A2(n_18),
.B1(n_25),
.B2(n_46),
.Y(n_86)
);

INVxp67_ASAP7_75t_L g102 ( 
.A(n_86),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_66),
.Y(n_87)
);

INVx13_ASAP7_75t_L g106 ( 
.A(n_87),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_48),
.A2(n_25),
.B1(n_46),
.B2(n_43),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_90),
.A2(n_91),
.B1(n_97),
.B2(n_100),
.Y(n_109)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_63),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_92),
.B(n_98),
.Y(n_111)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_93),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_94),
.B(n_64),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_95),
.A2(n_29),
.B1(n_21),
.B2(n_60),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_66),
.Y(n_96)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_96),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_L g97 ( 
.A1(n_68),
.A2(n_28),
.B1(n_29),
.B2(n_21),
.Y(n_97)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_47),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_L g100 ( 
.A1(n_68),
.A2(n_21),
.B1(n_28),
.B2(n_29),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g155 ( 
.A(n_101),
.B(n_12),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_71),
.B(n_57),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_105),
.B(n_118),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_107),
.A2(n_120),
.B1(n_124),
.B2(n_126),
.Y(n_149)
);

AND2x6_ASAP7_75t_L g110 ( 
.A(n_99),
.B(n_16),
.Y(n_110)
);

XNOR2x1_ASAP7_75t_SL g139 ( 
.A(n_110),
.B(n_77),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_93),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_113),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_71),
.A2(n_49),
.B1(n_66),
.B2(n_60),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_116),
.A2(n_87),
.B1(n_96),
.B2(n_76),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_79),
.B(n_80),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_91),
.A2(n_49),
.B1(n_69),
.B2(n_54),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_94),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_121),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_73),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_122),
.Y(n_160)
);

INVxp67_ASAP7_75t_L g143 ( 
.A(n_123),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_82),
.A2(n_37),
.B1(n_26),
.B2(n_23),
.Y(n_124)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_72),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_125),
.B(n_127),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_81),
.A2(n_37),
.B1(n_20),
.B2(n_34),
.Y(n_126)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_72),
.Y(n_127)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_73),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_128),
.B(n_129),
.Y(n_145)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_88),
.Y(n_129)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_111),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_130),
.B(n_132),
.Y(n_166)
);

INVx2_ASAP7_75t_SL g131 ( 
.A(n_106),
.Y(n_131)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_131),
.Y(n_173)
);

CKINVDCx16_ASAP7_75t_R g132 ( 
.A(n_108),
.Y(n_132)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_111),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_133),
.B(n_140),
.Y(n_174)
);

AOI21xp5_ASAP7_75t_L g134 ( 
.A1(n_129),
.A2(n_83),
.B(n_98),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_SL g163 ( 
.A1(n_134),
.A2(n_139),
.B(n_150),
.Y(n_163)
);

OR2x2_ASAP7_75t_L g135 ( 
.A(n_122),
.B(n_85),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_135),
.B(n_137),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_105),
.B(n_92),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_102),
.A2(n_86),
.B1(n_78),
.B2(n_87),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_138),
.A2(n_152),
.B1(n_107),
.B2(n_126),
.Y(n_161)
);

CKINVDCx14_ASAP7_75t_R g140 ( 
.A(n_108),
.Y(n_140)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_103),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_142),
.B(n_148),
.Y(n_189)
);

AOI22xp33_ASAP7_75t_SL g144 ( 
.A1(n_106),
.A2(n_76),
.B1(n_84),
.B2(n_89),
.Y(n_144)
);

AOI21xp5_ASAP7_75t_L g171 ( 
.A1(n_144),
.A2(n_151),
.B(n_119),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_125),
.B(n_84),
.Y(n_146)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_146),
.Y(n_164)
);

INVx1_ASAP7_75t_SL g148 ( 
.A(n_106),
.Y(n_148)
);

AOI21xp5_ASAP7_75t_L g150 ( 
.A1(n_115),
.A2(n_75),
.B(n_89),
.Y(n_150)
);

AOI22xp33_ASAP7_75t_SL g151 ( 
.A1(n_112),
.A2(n_76),
.B1(n_77),
.B2(n_53),
.Y(n_151)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_103),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_153),
.B(n_155),
.Y(n_167)
);

CKINVDCx16_ASAP7_75t_R g154 ( 
.A(n_116),
.Y(n_154)
);

INVxp67_ASAP7_75t_SL g168 ( 
.A(n_154),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_121),
.B(n_53),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_156),
.B(n_158),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_124),
.B(n_37),
.Y(n_158)
);

AOI21xp5_ASAP7_75t_L g159 ( 
.A1(n_115),
.A2(n_110),
.B(n_113),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_SL g169 ( 
.A1(n_159),
.A2(n_104),
.B(n_127),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_L g200 ( 
.A1(n_161),
.A2(n_171),
.B1(n_151),
.B2(n_144),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_139),
.A2(n_110),
.B1(n_128),
.B2(n_118),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_165),
.A2(n_188),
.B1(n_112),
.B2(n_148),
.Y(n_217)
);

XOR2xp5_ASAP7_75t_L g202 ( 
.A(n_169),
.B(n_182),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g172 ( 
.A(n_150),
.B(n_104),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_172),
.B(n_177),
.C(n_180),
.Y(n_209)
);

OAI21xp5_ASAP7_75t_SL g175 ( 
.A1(n_134),
.A2(n_159),
.B(n_145),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_L g195 ( 
.A1(n_175),
.A2(n_176),
.B(n_143),
.Y(n_195)
);

AOI21xp5_ASAP7_75t_L g176 ( 
.A1(n_134),
.A2(n_114),
.B(n_101),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_136),
.B(n_114),
.C(n_120),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_136),
.B(n_109),
.Y(n_178)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_178),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_137),
.B(n_157),
.Y(n_179)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_179),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_149),
.B(n_119),
.C(n_109),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_156),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_181),
.B(n_193),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g182 ( 
.A(n_149),
.B(n_34),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_149),
.B(n_117),
.C(n_96),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_183),
.B(n_184),
.C(n_185),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_139),
.B(n_117),
.C(n_74),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_157),
.B(n_117),
.C(n_74),
.Y(n_185)
);

XOR2xp5_ASAP7_75t_L g186 ( 
.A(n_158),
.B(n_34),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_186),
.B(n_187),
.C(n_190),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g187 ( 
.A(n_145),
.B(n_33),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_154),
.A2(n_112),
.B1(n_20),
.B2(n_33),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_132),
.B(n_140),
.C(n_153),
.Y(n_190)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_131),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_191),
.B(n_131),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_SL g192 ( 
.A(n_138),
.B(n_33),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_192),
.B(n_20),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_141),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_SL g194 ( 
.A(n_165),
.B(n_141),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_194),
.B(n_206),
.C(n_214),
.Y(n_229)
);

AOI21xp5_ASAP7_75t_L g226 ( 
.A1(n_195),
.A2(n_198),
.B(n_170),
.Y(n_226)
);

INVxp33_ASAP7_75t_SL g196 ( 
.A(n_168),
.Y(n_196)
);

INVxp33_ASAP7_75t_SL g234 ( 
.A(n_196),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_179),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_197),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_L g198 ( 
.A1(n_176),
.A2(n_160),
.B(n_147),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_162),
.B(n_160),
.Y(n_199)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_199),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_L g241 ( 
.A1(n_200),
.A2(n_210),
.B1(n_217),
.B2(n_185),
.Y(n_241)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_203),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_SL g204 ( 
.A(n_174),
.B(n_146),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_204),
.B(n_207),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_SL g206 ( 
.A(n_172),
.B(n_138),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_191),
.B(n_147),
.Y(n_207)
);

OR2x2_ASAP7_75t_L g208 ( 
.A(n_166),
.B(n_135),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_208),
.B(n_162),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_L g210 ( 
.A1(n_161),
.A2(n_133),
.B1(n_130),
.B2(n_142),
.Y(n_210)
);

BUFx12f_ASAP7_75t_SL g211 ( 
.A(n_175),
.Y(n_211)
);

OAI21xp5_ASAP7_75t_SL g227 ( 
.A1(n_211),
.A2(n_171),
.B(n_184),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_163),
.B(n_152),
.C(n_135),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_215),
.B(n_192),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_SL g216 ( 
.A(n_167),
.B(n_155),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g243 ( 
.A(n_216),
.B(n_221),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_163),
.B(n_148),
.C(n_131),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_219),
.B(n_212),
.C(n_213),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_180),
.A2(n_20),
.B1(n_1),
.B2(n_2),
.Y(n_220)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_220),
.Y(n_235)
);

CKINVDCx14_ASAP7_75t_R g221 ( 
.A(n_189),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_164),
.B(n_16),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_222),
.B(n_167),
.Y(n_237)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_224),
.Y(n_252)
);

OAI21xp5_ASAP7_75t_SL g256 ( 
.A1(n_226),
.A2(n_248),
.B(n_224),
.Y(n_256)
);

AOI21xp5_ASAP7_75t_L g249 ( 
.A1(n_227),
.A2(n_247),
.B(n_219),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_228),
.B(n_244),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_230),
.B(n_239),
.Y(n_251)
);

HB1xp67_ASAP7_75t_L g231 ( 
.A(n_211),
.Y(n_231)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_231),
.Y(n_264)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_201),
.Y(n_232)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_232),
.Y(n_269)
);

CKINVDCx16_ASAP7_75t_R g236 ( 
.A(n_199),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g262 ( 
.A(n_236),
.B(n_237),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_206),
.B(n_169),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_209),
.B(n_177),
.C(n_183),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_240),
.B(n_244),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_241),
.A2(n_213),
.B1(n_218),
.B2(n_202),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_L g242 ( 
.A1(n_217),
.A2(n_178),
.B1(n_190),
.B2(n_170),
.Y(n_242)
);

CKINVDCx16_ASAP7_75t_R g267 ( 
.A(n_242),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_209),
.B(n_186),
.C(n_187),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_195),
.A2(n_182),
.B1(n_188),
.B2(n_173),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_245),
.A2(n_214),
.B1(n_205),
.B2(n_212),
.Y(n_259)
);

AOI21x1_ASAP7_75t_SL g246 ( 
.A1(n_198),
.A2(n_173),
.B(n_1),
.Y(n_246)
);

AOI21xp5_ASAP7_75t_SL g265 ( 
.A1(n_246),
.A2(n_0),
.B(n_2),
.Y(n_265)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_220),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_197),
.Y(n_248)
);

NAND4xp25_ASAP7_75t_L g279 ( 
.A(n_249),
.B(n_226),
.C(n_245),
.D(n_243),
.Y(n_279)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_250),
.B(n_253),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_229),
.B(n_202),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_SL g254 ( 
.A(n_239),
.B(n_194),
.Y(n_254)
);

XOR2xp5_ASAP7_75t_L g287 ( 
.A(n_254),
.B(n_270),
.Y(n_287)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_256),
.Y(n_276)
);

INVx8_ASAP7_75t_L g257 ( 
.A(n_234),
.Y(n_257)
);

AOI22xp33_ASAP7_75t_SL g272 ( 
.A1(n_257),
.A2(n_233),
.B1(n_247),
.B2(n_225),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_232),
.B(n_205),
.Y(n_258)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_258),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_259),
.A2(n_261),
.B1(n_263),
.B2(n_266),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_260),
.B(n_265),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_235),
.A2(n_218),
.B1(n_208),
.B2(n_216),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_235),
.A2(n_215),
.B1(n_1),
.B2(n_2),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_225),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_223),
.B(n_10),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_268),
.A2(n_233),
.B1(n_11),
.B2(n_12),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_229),
.B(n_10),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_L g292 ( 
.A1(n_272),
.A2(n_279),
.B1(n_262),
.B2(n_266),
.Y(n_292)
);

BUFx2_ASAP7_75t_L g274 ( 
.A(n_257),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_274),
.B(n_269),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_255),
.B(n_230),
.C(n_240),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_275),
.B(n_285),
.C(n_251),
.Y(n_293)
);

OR2x2_ASAP7_75t_L g277 ( 
.A(n_252),
.B(n_246),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_277),
.B(n_274),
.Y(n_298)
);

XNOR2x1_ASAP7_75t_L g278 ( 
.A(n_254),
.B(n_227),
.Y(n_278)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_278),
.B(n_281),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_250),
.B(n_228),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_260),
.B(n_238),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g296 ( 
.A(n_282),
.B(n_253),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_283),
.B(n_15),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_255),
.B(n_251),
.C(n_259),
.Y(n_285)
);

NAND4xp25_ASAP7_75t_L g286 ( 
.A(n_264),
.B(n_15),
.C(n_13),
.D(n_12),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_SL g289 ( 
.A(n_286),
.B(n_265),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_289),
.B(n_294),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_290),
.B(n_295),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_SL g291 ( 
.A1(n_276),
.A2(n_267),
.B1(n_261),
.B2(n_263),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_SL g310 ( 
.A1(n_291),
.A2(n_285),
.B1(n_287),
.B2(n_273),
.Y(n_310)
);

AOI21xp5_ASAP7_75t_L g313 ( 
.A1(n_292),
.A2(n_299),
.B(n_301),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_L g303 ( 
.A(n_293),
.B(n_296),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_SL g294 ( 
.A(n_283),
.B(n_270),
.Y(n_294)
);

OA21x2_ASAP7_75t_SL g297 ( 
.A1(n_278),
.A2(n_11),
.B(n_13),
.Y(n_297)
);

NOR2x1_ASAP7_75t_SL g312 ( 
.A(n_297),
.B(n_5),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_SL g304 ( 
.A1(n_298),
.A2(n_271),
.B1(n_302),
.B2(n_277),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_284),
.B(n_13),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_282),
.B(n_3),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_300),
.B(n_4),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_275),
.B(n_3),
.C(n_4),
.Y(n_301)
);

AOI21xp5_ASAP7_75t_L g302 ( 
.A1(n_280),
.A2(n_4),
.B(n_5),
.Y(n_302)
);

OAI21xp5_ASAP7_75t_L g314 ( 
.A1(n_302),
.A2(n_301),
.B(n_6),
.Y(n_314)
);

XOR2xp5_ASAP7_75t_L g316 ( 
.A(n_304),
.B(n_305),
.Y(n_316)
);

XNOR2xp5_ASAP7_75t_L g305 ( 
.A(n_296),
.B(n_281),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_SL g321 ( 
.A(n_307),
.B(n_308),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_291),
.B(n_287),
.Y(n_308)
);

HB1xp67_ASAP7_75t_L g309 ( 
.A(n_298),
.Y(n_309)
);

INVxp67_ASAP7_75t_L g319 ( 
.A(n_309),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_SL g322 ( 
.A(n_310),
.B(n_312),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_314),
.B(n_7),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_SL g315 ( 
.A(n_313),
.B(n_293),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_315),
.B(n_318),
.Y(n_328)
);

OAI22xp5_ASAP7_75t_L g317 ( 
.A1(n_311),
.A2(n_288),
.B1(n_273),
.B2(n_7),
.Y(n_317)
);

INVxp33_ASAP7_75t_L g326 ( 
.A(n_317),
.Y(n_326)
);

AOI21xp5_ASAP7_75t_SL g318 ( 
.A1(n_306),
.A2(n_288),
.B(n_6),
.Y(n_318)
);

BUFx24_ASAP7_75t_SL g320 ( 
.A(n_303),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_320),
.B(n_324),
.Y(n_329)
);

NOR4xp25_ASAP7_75t_L g330 ( 
.A(n_323),
.B(n_7),
.C(n_314),
.D(n_319),
.Y(n_330)
);

AOI21xp5_ASAP7_75t_SL g324 ( 
.A1(n_303),
.A2(n_5),
.B(n_6),
.Y(n_324)
);

XNOR2xp5_ASAP7_75t_L g325 ( 
.A(n_321),
.B(n_305),
.Y(n_325)
);

XOR2xp5_ASAP7_75t_L g332 ( 
.A(n_325),
.B(n_331),
.Y(n_332)
);

AND2x2_ASAP7_75t_L g327 ( 
.A(n_316),
.B(n_310),
.Y(n_327)
);

MAJx2_ASAP7_75t_L g333 ( 
.A(n_327),
.B(n_330),
.C(n_326),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_322),
.B(n_7),
.Y(n_331)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_333),
.Y(n_335)
);

INVxp67_ASAP7_75t_L g334 ( 
.A(n_328),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_335),
.B(n_332),
.C(n_329),
.Y(n_336)
);

XNOR2xp5_ASAP7_75t_L g337 ( 
.A(n_336),
.B(n_334),
.Y(n_337)
);


endmodule