module fake_jpeg_24878_n_206 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_206);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_206;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_125;
wire n_80;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_2),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_0),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_1),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_12),
.Y(n_16)
);

INVx13_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

INVx3_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_1),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_11),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_4),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_9),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_SL g26 ( 
.A(n_15),
.B(n_0),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_26),
.B(n_29),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

INVx5_ASAP7_75t_L g49 ( 
.A(n_27),
.Y(n_49)
);

INVx5_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

AOI22xp33_ASAP7_75t_SL g40 ( 
.A1(n_28),
.A2(n_31),
.B1(n_17),
.B2(n_18),
.Y(n_40)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_17),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_30),
.Y(n_46)
);

INVx11_ASAP7_75t_L g31 ( 
.A(n_17),
.Y(n_31)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_32),
.B(n_18),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_17),
.Y(n_33)
);

BUFx4f_ASAP7_75t_SL g36 ( 
.A(n_33),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_14),
.B(n_0),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_34),
.B(n_20),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_SL g35 ( 
.A(n_15),
.B(n_1),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_35),
.B(n_15),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g38 ( 
.A(n_26),
.B(n_24),
.Y(n_38)
);

OAI21xp33_ASAP7_75t_L g59 ( 
.A1(n_38),
.A2(n_42),
.B(n_48),
.Y(n_59)
);

AND2x2_ASAP7_75t_L g58 ( 
.A(n_39),
.B(n_33),
.Y(n_58)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_41),
.B(n_50),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_35),
.B(n_24),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_SL g43 ( 
.A1(n_28),
.A2(n_18),
.B1(n_24),
.B2(n_23),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_43),
.A2(n_28),
.B1(n_32),
.B2(n_31),
.Y(n_54)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_33),
.Y(n_44)
);

HB1xp67_ASAP7_75t_L g57 ( 
.A(n_44),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_L g45 ( 
.A1(n_28),
.A2(n_18),
.B1(n_23),
.B2(n_22),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_L g60 ( 
.A1(n_45),
.A2(n_29),
.B1(n_13),
.B2(n_25),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_34),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_47),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_34),
.B(n_16),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_31),
.B(n_16),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_51),
.B(n_32),
.Y(n_53)
);

CKINVDCx14_ASAP7_75t_R g70 ( 
.A(n_53),
.Y(n_70)
);

INVxp67_ASAP7_75t_L g81 ( 
.A(n_54),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_47),
.B(n_31),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_56),
.B(n_63),
.Y(n_75)
);

AND2x2_ASAP7_75t_L g71 ( 
.A(n_58),
.B(n_33),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_60),
.A2(n_64),
.B1(n_49),
.B2(n_29),
.Y(n_74)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_36),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_61),
.B(n_66),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_39),
.B(n_20),
.Y(n_63)
);

O2A1O1Ixp33_ASAP7_75t_SL g64 ( 
.A1(n_36),
.A2(n_33),
.B(n_30),
.C(n_27),
.Y(n_64)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_49),
.Y(n_65)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_65),
.Y(n_69)
);

INVx8_ASAP7_75t_L g66 ( 
.A(n_36),
.Y(n_66)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_49),
.Y(n_67)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_67),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_48),
.B(n_20),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_68),
.B(n_38),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_71),
.B(n_73),
.Y(n_96)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_57),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_72),
.B(n_74),
.Y(n_100)
);

XNOR2xp5_ASAP7_75t_L g73 ( 
.A(n_63),
.B(n_37),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_55),
.A2(n_30),
.B1(n_46),
.B2(n_51),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_76),
.A2(n_78),
.B1(n_64),
.B2(n_67),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_77),
.B(n_85),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_55),
.A2(n_46),
.B1(n_37),
.B2(n_29),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_57),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_79),
.B(n_84),
.Y(n_103)
);

AND2x2_ASAP7_75t_L g82 ( 
.A(n_56),
.B(n_33),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_82),
.B(n_58),
.Y(n_98)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_62),
.Y(n_84)
);

INVxp67_ASAP7_75t_SL g85 ( 
.A(n_65),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_62),
.B(n_42),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_86),
.B(n_41),
.Y(n_97)
);

OR2x2_ASAP7_75t_L g87 ( 
.A(n_70),
.B(n_52),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_87),
.B(n_101),
.Y(n_116)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_84),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_88),
.B(n_89),
.Y(n_118)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_83),
.Y(n_89)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_72),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_91),
.B(n_92),
.Y(n_108)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_75),
.Y(n_92)
);

OR2x2_ASAP7_75t_L g93 ( 
.A(n_78),
.B(n_52),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_93),
.B(n_94),
.Y(n_115)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_76),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_82),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_95),
.Y(n_107)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_97),
.Y(n_109)
);

OAI21xp5_ASAP7_75t_SL g110 ( 
.A1(n_98),
.A2(n_102),
.B(n_104),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_99),
.A2(n_40),
.B1(n_43),
.B2(n_53),
.Y(n_119)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_82),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_79),
.Y(n_102)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_74),
.Y(n_104)
);

INVxp67_ASAP7_75t_L g105 ( 
.A(n_103),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_105),
.B(n_117),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_96),
.B(n_71),
.C(n_73),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_106),
.B(n_113),
.C(n_92),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_104),
.A2(n_81),
.B1(n_71),
.B2(n_64),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_111),
.A2(n_112),
.B1(n_119),
.B2(n_46),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_94),
.A2(n_81),
.B1(n_58),
.B2(n_67),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_96),
.B(n_58),
.C(n_68),
.Y(n_113)
);

INVx1_ASAP7_75t_SL g114 ( 
.A(n_90),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_114),
.B(n_87),
.Y(n_128)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_88),
.Y(n_117)
);

XNOR2xp5_ASAP7_75t_L g120 ( 
.A(n_98),
.B(n_59),
.Y(n_120)
);

XNOR2xp5_ASAP7_75t_L g132 ( 
.A(n_120),
.B(n_50),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_SL g121 ( 
.A1(n_101),
.A2(n_95),
.B(n_100),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_L g127 ( 
.A1(n_121),
.A2(n_99),
.B(n_93),
.Y(n_127)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_118),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_122),
.B(n_138),
.Y(n_146)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_108),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_123),
.B(n_125),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_124),
.B(n_113),
.C(n_111),
.Y(n_145)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_110),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_115),
.B(n_87),
.Y(n_126)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_126),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_L g150 ( 
.A(n_127),
.B(n_132),
.Y(n_150)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_128),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_116),
.B(n_89),
.Y(n_129)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_129),
.Y(n_141)
);

HB1xp67_ASAP7_75t_L g130 ( 
.A(n_105),
.Y(n_130)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_130),
.Y(n_142)
);

OA21x2_ASAP7_75t_L g131 ( 
.A1(n_107),
.A2(n_102),
.B(n_36),
.Y(n_131)
);

OAI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_131),
.A2(n_133),
.B1(n_66),
.B2(n_61),
.Y(n_147)
);

OA21x2_ASAP7_75t_L g133 ( 
.A1(n_110),
.A2(n_36),
.B(n_65),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_L g135 ( 
.A1(n_116),
.A2(n_91),
.B(n_80),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_L g151 ( 
.A(n_135),
.B(n_137),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_114),
.B(n_69),
.Y(n_136)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_136),
.Y(n_143)
);

FAx1_ASAP7_75t_SL g138 ( 
.A(n_106),
.B(n_45),
.CI(n_44),
.CON(n_138),
.SN(n_138)
);

OAI21xp33_ASAP7_75t_L g144 ( 
.A1(n_126),
.A2(n_121),
.B(n_120),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_L g159 ( 
.A1(n_144),
.A2(n_153),
.B(n_146),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_L g154 ( 
.A(n_145),
.B(n_124),
.Y(n_154)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_147),
.Y(n_160)
);

XNOR2x1_ASAP7_75t_L g149 ( 
.A(n_133),
.B(n_112),
.Y(n_149)
);

OAI21x1_ASAP7_75t_SL g166 ( 
.A1(n_149),
.A2(n_20),
.B(n_19),
.Y(n_166)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_134),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_152),
.B(n_135),
.Y(n_158)
);

AND2x2_ASAP7_75t_L g153 ( 
.A(n_129),
.B(n_133),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_154),
.B(n_161),
.C(n_163),
.Y(n_174)
);

FAx1_ASAP7_75t_SL g155 ( 
.A(n_145),
.B(n_127),
.CI(n_150),
.CON(n_155),
.SN(n_155)
);

FAx1_ASAP7_75t_SL g171 ( 
.A(n_155),
.B(n_159),
.CI(n_19),
.CON(n_171),
.SN(n_171)
);

NOR2xp33_ASAP7_75t_SL g156 ( 
.A(n_143),
.B(n_109),
.Y(n_156)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_156),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_149),
.A2(n_122),
.B1(n_137),
.B2(n_131),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_157),
.A2(n_162),
.B1(n_166),
.B2(n_142),
.Y(n_169)
);

OAI211xp5_ASAP7_75t_L g167 ( 
.A1(n_158),
.A2(n_164),
.B(n_147),
.C(n_13),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_L g161 ( 
.A1(n_153),
.A2(n_131),
.B(n_138),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_148),
.A2(n_138),
.B1(n_132),
.B2(n_66),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_L g163 ( 
.A(n_151),
.B(n_61),
.Y(n_163)
);

OAI21x1_ASAP7_75t_L g164 ( 
.A1(n_144),
.A2(n_12),
.B(n_20),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_140),
.B(n_16),
.Y(n_165)
);

OR2x2_ASAP7_75t_L g168 ( 
.A(n_165),
.B(n_13),
.Y(n_168)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_167),
.Y(n_178)
);

AOI31xp67_ASAP7_75t_SL g179 ( 
.A1(n_168),
.A2(n_21),
.A3(n_3),
.B(n_4),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_169),
.A2(n_175),
.B1(n_2),
.B2(n_3),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_154),
.B(n_141),
.C(n_139),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_170),
.B(n_172),
.C(n_176),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_SL g180 ( 
.A(n_171),
.B(n_19),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_159),
.B(n_27),
.C(n_25),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_160),
.A2(n_25),
.B1(n_23),
.B2(n_22),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_161),
.B(n_155),
.C(n_163),
.Y(n_176)
);

A2O1A1Ixp33_ASAP7_75t_L g177 ( 
.A1(n_157),
.A2(n_22),
.B(n_21),
.C(n_19),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_177),
.B(n_21),
.Y(n_182)
);

OR2x2_ASAP7_75t_L g187 ( 
.A(n_179),
.B(n_168),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_180),
.B(n_186),
.C(n_5),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_L g181 ( 
.A(n_174),
.B(n_19),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_181),
.B(n_183),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_182),
.B(n_184),
.Y(n_192)
);

AND2x2_ASAP7_75t_L g183 ( 
.A(n_176),
.B(n_2),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_170),
.B(n_3),
.C(n_4),
.Y(n_186)
);

OR2x2_ASAP7_75t_L g195 ( 
.A(n_187),
.B(n_188),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_178),
.B(n_173),
.Y(n_188)
);

INVxp67_ASAP7_75t_L g189 ( 
.A(n_182),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_L g196 ( 
.A1(n_189),
.A2(n_193),
.B(n_5),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_185),
.A2(n_172),
.B1(n_171),
.B2(n_177),
.Y(n_191)
);

INVxp67_ASAP7_75t_L g198 ( 
.A(n_191),
.Y(n_198)
);

AOI21x1_ASAP7_75t_L g194 ( 
.A1(n_188),
.A2(n_183),
.B(n_6),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g201 ( 
.A(n_194),
.B(n_190),
.Y(n_201)
);

BUFx24_ASAP7_75t_SL g199 ( 
.A(n_196),
.Y(n_199)
);

A2O1A1Ixp33_ASAP7_75t_SL g197 ( 
.A1(n_192),
.A2(n_6),
.B(n_7),
.C(n_8),
.Y(n_197)
);

AOI21x1_ASAP7_75t_L g200 ( 
.A1(n_197),
.A2(n_6),
.B(n_7),
.Y(n_200)
);

O2A1O1Ixp33_ASAP7_75t_L g204 ( 
.A1(n_200),
.A2(n_201),
.B(n_195),
.C(n_10),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_198),
.B(n_27),
.C(n_9),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_202),
.B(n_8),
.C(n_9),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_203),
.B(n_204),
.C(n_199),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_L g206 ( 
.A(n_205),
.B(n_10),
.Y(n_206)
);


endmodule