module real_jpeg_22930_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_247;
wire n_146;
wire n_78;
wire n_83;
wire n_288;
wire n_166;
wire n_176;
wire n_215;
wire n_221;
wire n_249;
wire n_286;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_280;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_281;
wire n_271;
wire n_163;
wire n_276;
wire n_22;
wire n_287;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_105;
wire n_40;
wire n_243;
wire n_173;
wire n_255;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_275;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_120;
wire n_113;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_282;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_44;
wire n_28;
wire n_267;
wire n_208;
wire n_62;
wire n_239;
wire n_162;
wire n_290;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_211;
wire n_285;
wire n_45;
wire n_172;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_262;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_258;
wire n_205;
wire n_195;
wire n_110;
wire n_289;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_228;
wire n_150;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_278;
wire n_241;
wire n_103;
wire n_225;
wire n_259;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_284;
wire n_226;
wire n_277;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_191;
wire n_52;
wire n_58;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_279;
wire n_128;
wire n_244;
wire n_167;
wire n_179;
wire n_216;
wire n_202;
wire n_133;
wire n_213;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_206;
wire n_210;
wire n_127;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_181;
wire n_85;
wire n_283;
wire n_101;
wire n_256;
wire n_274;
wire n_182;
wire n_273;
wire n_96;
wire n_253;
wire n_269;
wire n_89;

INVx3_ASAP7_75t_L g62 ( 
.A(n_0),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_1),
.A2(n_67),
.B1(n_76),
.B2(n_166),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_1),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_1),
.A2(n_60),
.B1(n_61),
.B2(n_166),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_L g229 ( 
.A1(n_1),
.A2(n_42),
.B1(n_43),
.B2(n_166),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_1),
.A2(n_29),
.B1(n_31),
.B2(n_166),
.Y(n_254)
);

AOI22xp33_ASAP7_75t_SL g41 ( 
.A1(n_2),
.A2(n_42),
.B1(n_43),
.B2(n_44),
.Y(n_41)
);

CKINVDCx16_ASAP7_75t_R g44 ( 
.A(n_2),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_2),
.A2(n_44),
.B1(n_60),
.B2(n_61),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_2),
.A2(n_29),
.B1(n_31),
.B2(n_44),
.Y(n_182)
);

AOI21xp5_ASAP7_75t_L g160 ( 
.A1(n_3),
.A2(n_72),
.B(n_161),
.Y(n_160)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_3),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_3),
.B(n_59),
.Y(n_193)
);

OAI22xp33_ASAP7_75t_L g228 ( 
.A1(n_3),
.A2(n_42),
.B1(n_43),
.B2(n_163),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_3),
.B(n_29),
.C(n_47),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_3),
.B(n_80),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_3),
.A2(n_95),
.B1(n_247),
.B2(n_254),
.Y(n_256)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_4),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_6),
.A2(n_70),
.B1(n_71),
.B2(n_72),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_6),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g157 ( 
.A1(n_6),
.A2(n_60),
.B1(n_61),
.B2(n_70),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g211 ( 
.A1(n_6),
.A2(n_42),
.B1(n_43),
.B2(n_70),
.Y(n_211)
);

AOI22xp33_ASAP7_75t_L g239 ( 
.A1(n_6),
.A2(n_29),
.B1(n_31),
.B2(n_70),
.Y(n_239)
);

INVx8_ASAP7_75t_SL g65 ( 
.A(n_7),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_8),
.A2(n_76),
.B1(n_117),
.B2(n_118),
.Y(n_116)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_8),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_SL g156 ( 
.A1(n_8),
.A2(n_60),
.B1(n_61),
.B2(n_117),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g210 ( 
.A1(n_8),
.A2(n_42),
.B1(n_43),
.B2(n_117),
.Y(n_210)
);

AOI22xp33_ASAP7_75t_L g244 ( 
.A1(n_8),
.A2(n_29),
.B1(n_31),
.B2(n_117),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g52 ( 
.A1(n_9),
.A2(n_42),
.B1(n_43),
.B2(n_53),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_9),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_9),
.A2(n_29),
.B1(n_31),
.B2(n_53),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_9),
.A2(n_53),
.B1(n_60),
.B2(n_61),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g33 ( 
.A1(n_10),
.A2(n_29),
.B1(n_31),
.B2(n_34),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_10),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_10),
.A2(n_34),
.B1(n_60),
.B2(n_61),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_L g92 ( 
.A1(n_10),
.A2(n_34),
.B1(n_42),
.B2(n_43),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_L g137 ( 
.A1(n_10),
.A2(n_34),
.B1(n_67),
.B2(n_76),
.Y(n_137)
);

BUFx5_ASAP7_75t_L g81 ( 
.A(n_11),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g28 ( 
.A1(n_12),
.A2(n_29),
.B1(n_30),
.B2(n_31),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_12),
.Y(n_30)
);

AOI22xp33_ASAP7_75t_L g75 ( 
.A1(n_12),
.A2(n_30),
.B1(n_67),
.B2(n_76),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_12),
.A2(n_30),
.B1(n_60),
.B2(n_61),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_12),
.A2(n_30),
.B1(n_42),
.B2(n_43),
.Y(n_128)
);

INVx13_ASAP7_75t_L g67 ( 
.A(n_13),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_14),
.Y(n_43)
);

INVx6_ASAP7_75t_L g27 ( 
.A(n_15),
.Y(n_27)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_15),
.Y(n_37)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_15),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_146),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_144),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_120),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_SL g145 ( 
.A(n_19),
.B(n_120),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_88),
.C(n_99),
.Y(n_19)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_20),
.A2(n_21),
.B1(n_88),
.B2(n_289),
.Y(n_288)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

XNOR2xp5_ASAP7_75t_SL g21 ( 
.A(n_22),
.B(n_54),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_22),
.B(n_56),
.C(n_77),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_38),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_23),
.A2(n_24),
.B1(n_38),
.B2(n_39),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_24),
.Y(n_23)
);

AND2x2_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_32),
.Y(n_24)
);

OAI21xp5_ASAP7_75t_L g238 ( 
.A1(n_25),
.A2(n_95),
.B(n_239),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_28),
.Y(n_25)
);

INVx3_ASAP7_75t_SL g26 ( 
.A(n_27),
.Y(n_26)
);

INVx5_ASAP7_75t_L g105 ( 
.A(n_27),
.Y(n_105)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_28),
.Y(n_98)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_29),
.Y(n_31)
);

AOI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_29),
.A2(n_31),
.B1(n_47),
.B2(n_49),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_31),
.B(n_36),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_SL g257 ( 
.A(n_31),
.B(n_258),
.Y(n_257)
);

OAI21xp5_ASAP7_75t_L g190 ( 
.A1(n_32),
.A2(n_182),
.B(n_191),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_SL g32 ( 
.A(n_33),
.B(n_35),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_33),
.B(n_105),
.Y(n_104)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_35),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_35),
.A2(n_36),
.B1(n_103),
.B2(n_181),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_35),
.A2(n_243),
.B1(n_245),
.B2(n_246),
.Y(n_242)
);

INVx5_ASAP7_75t_L g191 ( 
.A(n_36),
.Y(n_191)
);

INVx5_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_37),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_39),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_L g39 ( 
.A1(n_40),
.A2(n_45),
.B1(n_51),
.B2(n_52),
.Y(n_39)
);

INVxp67_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

OAI21xp5_ASAP7_75t_L g106 ( 
.A1(n_41),
.A2(n_50),
.B(n_107),
.Y(n_106)
);

OAI22xp33_ASAP7_75t_L g46 ( 
.A1(n_42),
.A2(n_43),
.B1(n_47),
.B2(n_49),
.Y(n_46)
);

AO22x1_ASAP7_75t_L g80 ( 
.A1(n_42),
.A2(n_43),
.B1(n_81),
.B2(n_82),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_42),
.B(n_82),
.Y(n_206)
);

INVx1_ASAP7_75t_SL g42 ( 
.A(n_43),
.Y(n_42)
);

OAI32xp33_ASAP7_75t_L g204 ( 
.A1(n_43),
.A2(n_61),
.A3(n_81),
.B1(n_205),
.B2(n_206),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_43),
.B(n_231),
.Y(n_230)
);

AOI21xp5_ASAP7_75t_L g90 ( 
.A1(n_45),
.A2(n_52),
.B(n_91),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_45),
.B(n_108),
.Y(n_107)
);

AOI21xp5_ASAP7_75t_L g154 ( 
.A1(n_45),
.A2(n_91),
.B(n_128),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_45),
.A2(n_51),
.B1(n_210),
.B2(n_211),
.Y(n_209)
);

AOI21xp5_ASAP7_75t_L g221 ( 
.A1(n_45),
.A2(n_126),
.B(n_211),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_45),
.A2(n_51),
.B1(n_228),
.B2(n_229),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_45),
.A2(n_51),
.B1(n_210),
.B2(n_229),
.Y(n_236)
);

AND2x2_ASAP7_75t_L g45 ( 
.A(n_46),
.B(n_50),
.Y(n_45)
);

INVx13_ASAP7_75t_L g49 ( 
.A(n_47),
.Y(n_49)
);

BUFx24_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_50),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_50),
.B(n_92),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_50),
.B(n_127),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_SL g252 ( 
.A(n_50),
.B(n_163),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g54 ( 
.A1(n_55),
.A2(n_56),
.B1(n_77),
.B2(n_78),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

AOI21xp5_ASAP7_75t_L g56 ( 
.A1(n_57),
.A2(n_69),
.B(n_74),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_57),
.A2(n_59),
.B1(n_69),
.B2(n_116),
.Y(n_115)
);

AOI21xp5_ASAP7_75t_L g134 ( 
.A1(n_57),
.A2(n_135),
.B(n_136),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_57),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_57),
.A2(n_59),
.B1(n_116),
.B2(n_165),
.Y(n_172)
);

AND2x2_ASAP7_75t_SL g57 ( 
.A(n_58),
.B(n_66),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_58),
.B(n_75),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_58),
.B(n_137),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_58),
.A2(n_159),
.B1(n_160),
.B2(n_164),
.Y(n_158)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g59 ( 
.A1(n_60),
.A2(n_61),
.B1(n_63),
.B2(n_64),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_L g86 ( 
.A1(n_60),
.A2(n_61),
.B1(n_81),
.B2(n_82),
.Y(n_86)
);

A2O1A1Ixp33_ASAP7_75t_L g177 ( 
.A1(n_60),
.A2(n_64),
.B(n_162),
.C(n_178),
.Y(n_177)
);

HAxp5_ASAP7_75t_SL g205 ( 
.A(n_60),
.B(n_163),
.CON(n_205),
.SN(n_205)
);

INVx3_ASAP7_75t_SL g60 ( 
.A(n_61),
.Y(n_60)
);

NAND3xp33_ASAP7_75t_L g178 ( 
.A(n_61),
.B(n_63),
.C(n_119),
.Y(n_178)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

OAI22xp33_ASAP7_75t_L g66 ( 
.A1(n_63),
.A2(n_64),
.B1(n_67),
.B2(n_68),
.Y(n_66)
);

CKINVDCx5p33_ASAP7_75t_R g63 ( 
.A(n_64),
.Y(n_63)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx8_ASAP7_75t_L g68 ( 
.A(n_67),
.Y(n_68)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_67),
.Y(n_73)
);

INVx11_ASAP7_75t_L g76 ( 
.A(n_67),
.Y(n_76)
);

INVx8_ASAP7_75t_L g119 ( 
.A(n_67),
.Y(n_119)
);

INVx8_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx8_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_73),
.B(n_163),
.Y(n_162)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_75),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_78),
.Y(n_77)
);

OAI21xp5_ASAP7_75t_L g78 ( 
.A1(n_79),
.A2(n_83),
.B(n_84),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_79),
.A2(n_83),
.B1(n_113),
.B2(n_130),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_79),
.A2(n_113),
.B1(n_156),
.B2(n_157),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_79),
.A2(n_113),
.B1(n_156),
.B2(n_195),
.Y(n_194)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_80),
.B(n_86),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_80),
.B(n_87),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_80),
.B(n_112),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_80),
.A2(n_85),
.B1(n_196),
.B2(n_205),
.Y(n_208)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_81),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_85),
.B(n_87),
.Y(n_84)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_85),
.Y(n_113)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_88),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_89),
.A2(n_90),
.B1(n_93),
.B2(n_94),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_90),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_90),
.B(n_93),
.Y(n_139)
);

INVxp67_ASAP7_75t_L g108 ( 
.A(n_92),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_93),
.A2(n_94),
.B1(n_134),
.B2(n_138),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_94),
.Y(n_93)
);

AOI21xp5_ASAP7_75t_L g94 ( 
.A1(n_95),
.A2(n_96),
.B(n_98),
.Y(n_94)
);

OAI21xp5_ASAP7_75t_L g101 ( 
.A1(n_95),
.A2(n_102),
.B(n_104),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_L g207 ( 
.A1(n_95),
.A2(n_98),
.B(n_104),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_95),
.A2(n_96),
.B1(n_244),
.B2(n_254),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_96),
.B(n_163),
.Y(n_258)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_99),
.B(n_288),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_100),
.B(n_109),
.C(n_115),
.Y(n_99)
);

XNOR2xp5_ASAP7_75t_SL g279 ( 
.A(n_100),
.B(n_280),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_101),
.B(n_106),
.Y(n_100)
);

XOR2xp5_ASAP7_75t_L g151 ( 
.A(n_101),
.B(n_106),
.Y(n_151)
);

INVxp67_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_107),
.B(n_125),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_109),
.A2(n_110),
.B1(n_115),
.B2(n_281),
.Y(n_280)
);

CKINVDCx14_ASAP7_75t_R g109 ( 
.A(n_110),
.Y(n_109)
);

OAI21xp5_ASAP7_75t_L g110 ( 
.A1(n_111),
.A2(n_113),
.B(n_114),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

OAI21xp33_ASAP7_75t_L g174 ( 
.A1(n_113),
.A2(n_157),
.B(n_175),
.Y(n_174)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_115),
.Y(n_281)
);

INVx4_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_121),
.A2(n_122),
.B1(n_142),
.B2(n_143),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_123),
.A2(n_132),
.B1(n_140),
.B2(n_141),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_123),
.Y(n_140)
);

AOI21xp5_ASAP7_75t_L g123 ( 
.A1(n_124),
.A2(n_129),
.B(n_131),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_124),
.B(n_129),
.Y(n_131)
);

INVxp67_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_132),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_SL g132 ( 
.A(n_133),
.B(n_139),
.Y(n_132)
);

CKINVDCx16_ASAP7_75t_R g138 ( 
.A(n_134),
.Y(n_138)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_142),
.Y(n_143)
);

INVxp67_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_SL g146 ( 
.A1(n_147),
.A2(n_285),
.B(n_290),
.Y(n_146)
);

O2A1O1Ixp33_ASAP7_75t_SL g147 ( 
.A1(n_148),
.A2(n_197),
.B(n_273),
.C(n_284),
.Y(n_147)
);

AND2x2_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_183),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_149),
.B(n_183),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_169),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_151),
.A2(n_152),
.B1(n_167),
.B2(n_168),
.Y(n_150)
);

CKINVDCx16_ASAP7_75t_R g167 ( 
.A(n_151),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_151),
.B(n_168),
.C(n_169),
.Y(n_274)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_152),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_155),
.C(n_158),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_153),
.A2(n_154),
.B1(n_155),
.B2(n_186),
.Y(n_185)
);

CKINVDCx16_ASAP7_75t_R g153 ( 
.A(n_154),
.Y(n_153)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_155),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_SL g184 ( 
.A(n_158),
.B(n_185),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_162),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_165),
.Y(n_164)
);

XOR2xp5_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_176),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_171),
.A2(n_172),
.B1(n_173),
.B2(n_174),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_172),
.B(n_173),
.C(n_176),
.Y(n_282)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_177),
.B(n_179),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_177),
.A2(n_179),
.B1(n_180),
.B2(n_188),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_177),
.Y(n_188)
);

CKINVDCx16_ASAP7_75t_R g179 ( 
.A(n_180),
.Y(n_179)
);

INVxp67_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_187),
.C(n_189),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_184),
.B(n_271),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_187),
.B(n_189),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_190),
.B(n_192),
.C(n_194),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_190),
.A2(n_192),
.B1(n_193),
.B2(n_216),
.Y(n_215)
);

CKINVDCx14_ASAP7_75t_R g216 ( 
.A(n_190),
.Y(n_216)
);

CKINVDCx16_ASAP7_75t_R g192 ( 
.A(n_193),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g214 ( 
.A(n_194),
.B(n_215),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_196),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_199),
.Y(n_197)
);

AOI21xp5_ASAP7_75t_L g199 ( 
.A1(n_200),
.A2(n_268),
.B(n_272),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_L g200 ( 
.A1(n_201),
.A2(n_223),
.B(n_267),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_202),
.B(n_212),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g267 ( 
.A(n_202),
.B(n_212),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_203),
.B(n_208),
.C(n_209),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_203),
.B(n_265),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_SL g203 ( 
.A(n_204),
.B(n_207),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_204),
.B(n_207),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_208),
.B(n_209),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_213),
.A2(n_214),
.B1(n_217),
.B2(n_218),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_213),
.B(n_220),
.C(n_222),
.Y(n_269)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_219),
.A2(n_220),
.B1(n_221),
.B2(n_222),
.Y(n_218)
);

CKINVDCx16_ASAP7_75t_R g222 ( 
.A(n_219),
.Y(n_222)
);

CKINVDCx14_ASAP7_75t_R g220 ( 
.A(n_221),
.Y(n_220)
);

AOI21xp5_ASAP7_75t_L g223 ( 
.A1(n_224),
.A2(n_262),
.B(n_266),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_SL g224 ( 
.A1(n_225),
.A2(n_240),
.B(n_261),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_232),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_226),
.B(n_232),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_SL g226 ( 
.A(n_227),
.B(n_230),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_227),
.B(n_230),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_233),
.B(n_238),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_234),
.A2(n_235),
.B1(n_236),
.B2(n_237),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_234),
.B(n_237),
.C(n_238),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_235),
.Y(n_234)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_236),
.Y(n_237)
);

INVxp67_ASAP7_75t_L g245 ( 
.A(n_239),
.Y(n_245)
);

AOI21xp33_ASAP7_75t_L g240 ( 
.A1(n_241),
.A2(n_250),
.B(n_260),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_249),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_242),
.B(n_249),
.Y(n_260)
);

CKINVDCx16_ASAP7_75t_R g243 ( 
.A(n_244),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_247),
.Y(n_246)
);

BUFx2_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

OAI21xp5_ASAP7_75t_SL g250 ( 
.A1(n_251),
.A2(n_255),
.B(n_259),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_252),
.B(n_253),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_SL g259 ( 
.A(n_252),
.B(n_253),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_SL g255 ( 
.A(n_256),
.B(n_257),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_263),
.B(n_264),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_SL g266 ( 
.A(n_263),
.B(n_264),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_269),
.B(n_270),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_SL g272 ( 
.A(n_269),
.B(n_270),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_274),
.B(n_275),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_274),
.B(n_275),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_276),
.A2(n_277),
.B1(n_282),
.B2(n_283),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

XOR2xp5_ASAP7_75t_L g277 ( 
.A(n_278),
.B(n_279),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_278),
.B(n_279),
.C(n_283),
.Y(n_286)
);

CKINVDCx16_ASAP7_75t_R g283 ( 
.A(n_282),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_286),
.B(n_287),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_SL g290 ( 
.A(n_286),
.B(n_287),
.Y(n_290)
);


endmodule