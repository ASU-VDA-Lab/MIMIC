module fake_jpeg_9347_n_205 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_205);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_205;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx16f_ASAP7_75t_L g16 ( 
.A(n_15),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_9),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_13),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_6),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

BUFx8_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_13),
.Y(n_25)
);

INVx5_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_8),
.Y(n_27)
);

INVx11_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

INVx13_ASAP7_75t_L g31 ( 
.A(n_6),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

OR2x2_ASAP7_75t_L g33 ( 
.A(n_19),
.B(n_0),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_33),
.B(n_42),
.Y(n_49)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_16),
.Y(n_34)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_34),
.Y(n_57)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_28),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_35),
.B(n_38),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

CKINVDCx16_ASAP7_75t_R g45 ( 
.A(n_36),
.Y(n_45)
);

AOI21xp33_ASAP7_75t_SL g37 ( 
.A1(n_32),
.A2(n_16),
.B(n_20),
.Y(n_37)
);

OR2x2_ASAP7_75t_SL g46 ( 
.A(n_37),
.B(n_22),
.Y(n_46)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_28),
.Y(n_38)
);

INVx13_ASAP7_75t_L g39 ( 
.A(n_16),
.Y(n_39)
);

INVx5_ASAP7_75t_L g50 ( 
.A(n_39),
.Y(n_50)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_20),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_40),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_28),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_41),
.Y(n_62)
);

INVx5_ASAP7_75t_L g42 ( 
.A(n_22),
.Y(n_42)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_20),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_43),
.B(n_44),
.Y(n_53)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_21),
.Y(n_44)
);

AND2x2_ASAP7_75t_L g79 ( 
.A(n_46),
.B(n_54),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_40),
.A2(n_26),
.B1(n_23),
.B2(n_31),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g72 ( 
.A1(n_47),
.A2(n_58),
.B1(n_61),
.B2(n_64),
.Y(n_72)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_35),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_48),
.B(n_63),
.Y(n_67)
);

BUFx12_ASAP7_75t_L g52 ( 
.A(n_36),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_52),
.B(n_39),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_33),
.B(n_24),
.Y(n_54)
);

O2A1O1Ixp33_ASAP7_75t_L g55 ( 
.A1(n_37),
.A2(n_24),
.B(n_30),
.C(n_19),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_55),
.A2(n_27),
.B1(n_25),
.B2(n_42),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_33),
.B(n_18),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_SL g85 ( 
.A(n_56),
.B(n_59),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_L g58 ( 
.A1(n_40),
.A2(n_23),
.B1(n_26),
.B2(n_31),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_38),
.B(n_18),
.Y(n_59)
);

OAI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_44),
.A2(n_26),
.B1(n_31),
.B2(n_27),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_36),
.B(n_32),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_42),
.A2(n_30),
.B1(n_25),
.B2(n_17),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_41),
.B(n_17),
.Y(n_65)
);

AND2x2_ASAP7_75t_L g82 ( 
.A(n_65),
.B(n_0),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g66 ( 
.A1(n_46),
.A2(n_44),
.B1(n_43),
.B2(n_34),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_66),
.A2(n_80),
.B1(n_84),
.B2(n_57),
.Y(n_93)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_51),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_68),
.B(n_76),
.Y(n_89)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_50),
.Y(n_69)
);

INVx11_ASAP7_75t_L g95 ( 
.A(n_69),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_55),
.B(n_32),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_70),
.B(n_65),
.Y(n_100)
);

INVx11_ASAP7_75t_L g71 ( 
.A(n_62),
.Y(n_71)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_71),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g97 ( 
.A(n_73),
.Y(n_97)
);

XNOR2xp5_ASAP7_75t_L g87 ( 
.A(n_74),
.B(n_54),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g75 ( 
.A(n_53),
.Y(n_75)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_75),
.Y(n_98)
);

HB1xp67_ASAP7_75t_L g76 ( 
.A(n_52),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_57),
.A2(n_43),
.B1(n_34),
.B2(n_39),
.Y(n_77)
);

INVxp67_ASAP7_75t_L g105 ( 
.A(n_77),
.Y(n_105)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_50),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_78),
.B(n_81),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_60),
.A2(n_41),
.B1(n_21),
.B2(n_29),
.Y(n_80)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_62),
.Y(n_81)
);

OR2x2_ASAP7_75t_L g94 ( 
.A(n_82),
.B(n_0),
.Y(n_94)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_52),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_83),
.B(n_86),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_60),
.A2(n_21),
.B1(n_29),
.B2(n_32),
.Y(n_84)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_59),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_87),
.B(n_94),
.Y(n_114)
);

XNOR2xp5_ASAP7_75t_L g88 ( 
.A(n_70),
.B(n_49),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_88),
.B(n_96),
.C(n_86),
.Y(n_113)
);

A2O1A1Ixp33_ASAP7_75t_L g92 ( 
.A1(n_79),
.A2(n_49),
.B(n_56),
.C(n_63),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_92),
.B(n_106),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_93),
.A2(n_100),
.B1(n_68),
.B2(n_81),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_67),
.B(n_45),
.C(n_48),
.Y(n_96)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_67),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_99),
.B(n_101),
.Y(n_119)
);

HB1xp67_ASAP7_75t_L g101 ( 
.A(n_71),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_69),
.B(n_57),
.Y(n_103)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_103),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_78),
.B(n_52),
.Y(n_104)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_104),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_75),
.B(n_53),
.Y(n_106)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_80),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_107),
.B(n_108),
.Y(n_124)
);

OR2x2_ASAP7_75t_L g108 ( 
.A(n_85),
.B(n_1),
.Y(n_108)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_90),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_109),
.B(n_118),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_107),
.A2(n_100),
.B1(n_106),
.B2(n_74),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_110),
.A2(n_122),
.B1(n_98),
.B2(n_85),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_113),
.B(n_115),
.C(n_45),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_96),
.B(n_66),
.C(n_79),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_116),
.B(n_117),
.Y(n_136)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_89),
.Y(n_117)
);

INVxp67_ASAP7_75t_L g118 ( 
.A(n_91),
.Y(n_118)
);

INVx4_ASAP7_75t_L g120 ( 
.A(n_95),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_120),
.B(n_102),
.Y(n_129)
);

AOI21xp5_ASAP7_75t_L g121 ( 
.A1(n_105),
.A2(n_79),
.B(n_72),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_SL g141 ( 
.A1(n_121),
.A2(n_97),
.B(n_82),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_105),
.A2(n_92),
.B1(n_93),
.B2(n_98),
.Y(n_122)
);

BUFx24_ASAP7_75t_L g123 ( 
.A(n_102),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_123),
.B(n_126),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_99),
.B(n_88),
.Y(n_126)
);

A2O1A1Ixp33_ASAP7_75t_SL g127 ( 
.A1(n_87),
.A2(n_84),
.B(n_62),
.C(n_36),
.Y(n_127)
);

AO21x1_ASAP7_75t_L g142 ( 
.A1(n_127),
.A2(n_22),
.B(n_29),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_128),
.B(n_135),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_129),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_SL g130 ( 
.A(n_112),
.B(n_108),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_130),
.B(n_131),
.Y(n_147)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_119),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_SL g132 ( 
.A(n_121),
.B(n_94),
.C(n_82),
.Y(n_132)
);

NAND2xp33_ASAP7_75t_SL g149 ( 
.A(n_132),
.B(n_141),
.Y(n_149)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_123),
.Y(n_134)
);

INVxp67_ASAP7_75t_SL g159 ( 
.A(n_134),
.Y(n_159)
);

INVx5_ASAP7_75t_L g135 ( 
.A(n_123),
.Y(n_135)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_124),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_L g155 ( 
.A1(n_137),
.A2(n_139),
.B(n_111),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_138),
.B(n_140),
.C(n_144),
.Y(n_146)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_110),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_113),
.B(n_97),
.C(n_36),
.Y(n_140)
);

AO21x1_ASAP7_75t_L g151 ( 
.A1(n_141),
.A2(n_142),
.B(n_143),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_SL g143 ( 
.A1(n_125),
.A2(n_95),
.B(n_83),
.Y(n_143)
);

XOR2xp5_ASAP7_75t_L g144 ( 
.A(n_126),
.B(n_22),
.Y(n_144)
);

XOR2xp5_ASAP7_75t_L g148 ( 
.A(n_138),
.B(n_115),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_148),
.B(n_149),
.C(n_152),
.Y(n_164)
);

AOI22x1_ASAP7_75t_L g150 ( 
.A1(n_143),
.A2(n_125),
.B1(n_127),
.B2(n_118),
.Y(n_150)
);

AOI21xp5_ASAP7_75t_L g167 ( 
.A1(n_150),
.A2(n_136),
.B(n_120),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_140),
.B(n_114),
.C(n_109),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_155),
.B(n_158),
.Y(n_163)
);

HB1xp67_ASAP7_75t_L g156 ( 
.A(n_135),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_156),
.B(n_160),
.Y(n_170)
);

AOI221xp5_ASAP7_75t_L g157 ( 
.A1(n_128),
.A2(n_127),
.B1(n_10),
.B2(n_11),
.C(n_12),
.Y(n_157)
);

XOR2xp5_ASAP7_75t_L g171 ( 
.A(n_157),
.B(n_12),
.Y(n_171)
);

BUFx6f_ASAP7_75t_L g158 ( 
.A(n_134),
.Y(n_158)
);

A2O1A1O1Ixp25_ASAP7_75t_L g160 ( 
.A1(n_142),
.A2(n_127),
.B(n_2),
.C(n_3),
.D(n_4),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_147),
.Y(n_161)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_161),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_153),
.B(n_145),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_162),
.B(n_165),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_148),
.B(n_144),
.C(n_133),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_159),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_166),
.B(n_168),
.Y(n_176)
);

AOI21xp5_ASAP7_75t_SL g174 ( 
.A1(n_167),
.A2(n_151),
.B(n_146),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_150),
.B(n_1),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_159),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_SL g180 ( 
.A(n_169),
.B(n_171),
.Y(n_180)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_158),
.Y(n_172)
);

BUFx24_ASAP7_75t_SL g181 ( 
.A(n_172),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_154),
.B(n_160),
.Y(n_173)
);

OR2x2_ASAP7_75t_L g179 ( 
.A(n_173),
.B(n_170),
.Y(n_179)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_174),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_168),
.A2(n_151),
.B1(n_146),
.B2(n_11),
.Y(n_175)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_175),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_163),
.A2(n_10),
.B1(n_2),
.B2(n_3),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_177),
.B(n_179),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_182),
.B(n_164),
.C(n_165),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g190 ( 
.A(n_185),
.B(n_189),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_178),
.B(n_161),
.Y(n_186)
);

AOI21xp5_ASAP7_75t_L g191 ( 
.A1(n_186),
.A2(n_176),
.B(n_179),
.Y(n_191)
);

AOI21xp5_ASAP7_75t_L g187 ( 
.A1(n_180),
.A2(n_162),
.B(n_164),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_SL g195 ( 
.A1(n_187),
.A2(n_4),
.B(n_5),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_181),
.B(n_167),
.C(n_171),
.Y(n_189)
);

INVxp67_ASAP7_75t_L g199 ( 
.A(n_191),
.Y(n_199)
);

CKINVDCx16_ASAP7_75t_R g192 ( 
.A(n_188),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_192),
.B(n_193),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_184),
.B(n_174),
.Y(n_193)
);

AOI22xp33_ASAP7_75t_L g194 ( 
.A1(n_183),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_194)
);

AND2x2_ASAP7_75t_L g198 ( 
.A(n_194),
.B(n_195),
.Y(n_198)
);

NOR2xp67_ASAP7_75t_L g197 ( 
.A(n_190),
.B(n_186),
.Y(n_197)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_197),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_L g201 ( 
.A1(n_196),
.A2(n_194),
.B(n_4),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_201),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_199),
.B(n_198),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_202),
.B(n_200),
.Y(n_203)
);

XOR2xp5_ASAP7_75t_L g205 ( 
.A(n_203),
.B(n_204),
.Y(n_205)
);


endmodule