module fake_ariane_3345_n_46 (n_8, n_3, n_2, n_11, n_7, n_5, n_1, n_0, n_6, n_9, n_4, n_10, n_46);

input n_8;
input n_3;
input n_2;
input n_11;
input n_7;
input n_5;
input n_1;
input n_0;
input n_6;
input n_9;
input n_4;
input n_10;

output n_46;

wire n_24;
wire n_22;
wire n_43;
wire n_13;
wire n_20;
wire n_27;
wire n_29;
wire n_17;
wire n_41;
wire n_38;
wire n_18;
wire n_32;
wire n_28;
wire n_37;
wire n_45;
wire n_34;
wire n_26;
wire n_14;
wire n_36;
wire n_33;
wire n_44;
wire n_40;
wire n_30;
wire n_39;
wire n_19;
wire n_31;
wire n_42;
wire n_16;
wire n_12;
wire n_15;
wire n_21;
wire n_23;
wire n_35;
wire n_25;

INVx2_ASAP7_75t_SL g12 ( 
.A(n_3),
.Y(n_12)
);

INVx2_ASAP7_75t_L g13 ( 
.A(n_10),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_5),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_9),
.Y(n_15)
);

BUFx2_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_8),
.B(n_6),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_0),
.B(n_2),
.Y(n_22)
);

O2A1O1Ixp33_ASAP7_75t_L g23 ( 
.A1(n_22),
.A2(n_2),
.B(n_4),
.C(n_5),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_SL g24 ( 
.A(n_13),
.B(n_4),
.Y(n_24)
);

OAI22xp33_ASAP7_75t_L g25 ( 
.A1(n_16),
.A2(n_7),
.B1(n_12),
.B2(n_18),
.Y(n_25)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_18),
.Y(n_26)
);

OAI21xp5_ASAP7_75t_L g27 ( 
.A1(n_25),
.A2(n_13),
.B(n_21),
.Y(n_27)
);

OAI21x1_ASAP7_75t_L g28 ( 
.A1(n_24),
.A2(n_21),
.B(n_17),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_26),
.Y(n_29)
);

OAI21x1_ASAP7_75t_SL g30 ( 
.A1(n_23),
.A2(n_14),
.B(n_20),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_29),
.Y(n_31)
);

OAI21x1_ASAP7_75t_L g32 ( 
.A1(n_28),
.A2(n_26),
.B(n_15),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_29),
.Y(n_33)
);

CKINVDCx5p33_ASAP7_75t_R g34 ( 
.A(n_29),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_31),
.Y(n_35)
);

AND2x2_ASAP7_75t_L g36 ( 
.A(n_31),
.B(n_27),
.Y(n_36)
);

HB1xp67_ASAP7_75t_L g37 ( 
.A(n_36),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_37),
.Y(n_38)
);

AOI211xp5_ASAP7_75t_L g39 ( 
.A1(n_38),
.A2(n_28),
.B(n_36),
.C(n_29),
.Y(n_39)
);

AOI21xp5_ASAP7_75t_L g40 ( 
.A1(n_39),
.A2(n_35),
.B(n_32),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_L g41 ( 
.A1(n_40),
.A2(n_35),
.B1(n_34),
.B2(n_33),
.Y(n_41)
);

AOI222xp33_ASAP7_75t_L g42 ( 
.A1(n_40),
.A2(n_30),
.B1(n_29),
.B2(n_19),
.C1(n_15),
.C2(n_33),
.Y(n_42)
);

OAI211xp5_ASAP7_75t_SL g43 ( 
.A1(n_41),
.A2(n_32),
.B(n_15),
.C(n_19),
.Y(n_43)
);

OR2x6_ASAP7_75t_L g44 ( 
.A(n_42),
.B(n_32),
.Y(n_44)
);

OAI21xp5_ASAP7_75t_SL g45 ( 
.A1(n_43),
.A2(n_44),
.B(n_15),
.Y(n_45)
);

OR2x6_ASAP7_75t_L g46 ( 
.A(n_45),
.B(n_19),
.Y(n_46)
);


endmodule