module fake_jpeg_31668_n_88 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_88);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_88;

wire n_10;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_65;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_22;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;

INVx1_ASAP7_75t_L g10 ( 
.A(n_4),
.Y(n_10)
);

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_8),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_6),
.Y(n_12)
);

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_1),
.Y(n_13)
);

BUFx3_ASAP7_75t_L g14 ( 
.A(n_8),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_4),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_2),
.Y(n_17)
);

INVx8_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_SL g22 ( 
.A(n_11),
.B(n_3),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_22),
.B(n_25),
.Y(n_32)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_20),
.Y(n_23)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_23),
.Y(n_38)
);

INVx8_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

INVx13_ASAP7_75t_L g40 ( 
.A(n_24),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_12),
.B(n_5),
.Y(n_25)
);

INVx5_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

HB1xp67_ASAP7_75t_L g42 ( 
.A(n_26),
.Y(n_42)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_27),
.B(n_28),
.Y(n_34)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_21),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_20),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_29),
.B(n_31),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_17),
.B(n_5),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_30),
.Y(n_33)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_21),
.Y(n_31)
);

MAJIxp5_ASAP7_75t_L g35 ( 
.A(n_23),
.B(n_13),
.C(n_18),
.Y(n_35)
);

AND2x2_ASAP7_75t_L g48 ( 
.A(n_35),
.B(n_15),
.Y(n_48)
);

BUFx10_ASAP7_75t_L g37 ( 
.A(n_26),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_37),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_L g39 ( 
.A1(n_29),
.A2(n_24),
.B1(n_27),
.B2(n_28),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_39),
.B(n_41),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_L g41 ( 
.A1(n_31),
.A2(n_18),
.B1(n_19),
.B2(n_10),
.Y(n_41)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_40),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_43),
.B(n_47),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_33),
.B(n_22),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_SL g64 ( 
.A(n_45),
.B(n_49),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g47 ( 
.A(n_32),
.B(n_10),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_48),
.B(n_53),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_33),
.B(n_15),
.Y(n_49)
);

INVxp67_ASAP7_75t_L g50 ( 
.A(n_34),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_50),
.B(n_51),
.Y(n_63)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_32),
.B(n_16),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_52),
.Y(n_56)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_36),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_35),
.B(n_38),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_54),
.B(n_55),
.Y(n_58)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_38),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_51),
.A2(n_42),
.B1(n_19),
.B2(n_16),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_59),
.A2(n_60),
.B1(n_48),
.B2(n_46),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_53),
.A2(n_40),
.B1(n_37),
.B2(n_0),
.Y(n_60)
);

NOR3xp33_ASAP7_75t_L g61 ( 
.A(n_54),
.B(n_37),
.C(n_7),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_61),
.B(n_7),
.Y(n_68)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_59),
.Y(n_65)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_65),
.Y(n_75)
);

BUFx4f_ASAP7_75t_SL g66 ( 
.A(n_60),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_66),
.B(n_68),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_64),
.B(n_50),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_SL g74 ( 
.A(n_67),
.B(n_56),
.Y(n_74)
);

MAJx2_ASAP7_75t_L g69 ( 
.A(n_57),
.B(n_48),
.C(n_44),
.Y(n_69)
);

XOR2xp5_ASAP7_75t_L g73 ( 
.A(n_69),
.B(n_58),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_70),
.B(n_57),
.Y(n_72)
);

OAI32xp33_ASAP7_75t_L g76 ( 
.A1(n_72),
.A2(n_58),
.A3(n_63),
.B1(n_62),
.B2(n_69),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_73),
.B(n_66),
.C(n_55),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_74),
.Y(n_79)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_76),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_77),
.B(n_73),
.Y(n_80)
);

AOI21xp5_ASAP7_75t_L g78 ( 
.A1(n_71),
.A2(n_66),
.B(n_43),
.Y(n_78)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_78),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_80),
.B(n_37),
.C(n_40),
.Y(n_84)
);

NAND3xp33_ASAP7_75t_L g83 ( 
.A(n_81),
.B(n_79),
.C(n_75),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_83),
.B(n_84),
.Y(n_85)
);

AOI21x1_ASAP7_75t_L g86 ( 
.A1(n_85),
.A2(n_80),
.B(n_82),
.Y(n_86)
);

OAI21xp5_ASAP7_75t_SL g87 ( 
.A1(n_86),
.A2(n_9),
.B(n_0),
.Y(n_87)
);

NAND2xp33_ASAP7_75t_L g88 ( 
.A(n_87),
.B(n_0),
.Y(n_88)
);


endmodule