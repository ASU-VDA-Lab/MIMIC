module fake_netlist_5_993_n_1806 (n_137, n_168, n_164, n_91, n_82, n_122, n_142, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_165, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_60, n_155, n_152, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_125, n_35, n_167, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_156, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_157, n_29, n_79, n_131, n_151, n_47, n_25, n_53, n_160, n_8, n_158, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_85, n_159, n_163, n_95, n_119, n_59, n_26, n_133, n_55, n_99, n_2, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_12, n_67, n_121, n_36, n_76, n_87, n_150, n_162, n_27, n_64, n_77, n_102, n_106, n_161, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_134, n_32, n_41, n_104, n_103, n_56, n_51, n_63, n_97, n_141, n_166, n_11, n_153, n_7, n_15, n_145, n_48, n_50, n_52, n_88, n_110, n_1806);

input n_137;
input n_168;
input n_164;
input n_91;
input n_82;
input n_122;
input n_142;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_165;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_60;
input n_155;
input n_152;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_125;
input n_35;
input n_167;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_157;
input n_29;
input n_79;
input n_131;
input n_151;
input n_47;
input n_25;
input n_53;
input n_160;
input n_8;
input n_158;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_85;
input n_159;
input n_163;
input n_95;
input n_119;
input n_59;
input n_26;
input n_133;
input n_55;
input n_99;
input n_2;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_150;
input n_162;
input n_27;
input n_64;
input n_77;
input n_102;
input n_106;
input n_161;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_134;
input n_32;
input n_41;
input n_104;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_166;
input n_11;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_1806;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1729;
wire n_1166;
wire n_1751;
wire n_469;
wire n_1508;
wire n_785;
wire n_549;
wire n_532;
wire n_1161;
wire n_1677;
wire n_1150;
wire n_226;
wire n_1780;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_1501;
wire n_880;
wire n_544;
wire n_1007;
wire n_552;
wire n_1528;
wire n_1370;
wire n_1292;
wire n_1198;
wire n_1360;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1738;
wire n_1021;
wire n_551;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1695;
wire n_1353;
wire n_800;
wire n_1347;
wire n_1535;
wire n_1789;
wire n_1666;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_915;
wire n_1545;
wire n_864;
wire n_173;
wire n_859;
wire n_951;
wire n_1264;
wire n_447;
wire n_247;
wire n_1494;
wire n_292;
wire n_625;
wire n_854;
wire n_1462;
wire n_1799;
wire n_1580;
wire n_674;
wire n_417;
wire n_516;
wire n_933;
wire n_1152;
wire n_497;
wire n_1607;
wire n_1563;
wire n_606;
wire n_275;
wire n_877;
wire n_1696;
wire n_755;
wire n_1118;
wire n_1686;
wire n_947;
wire n_1285;
wire n_373;
wire n_307;
wire n_1359;
wire n_530;
wire n_1107;
wire n_1728;
wire n_556;
wire n_1230;
wire n_668;
wire n_375;
wire n_301;
wire n_929;
wire n_1124;
wire n_902;
wire n_1576;
wire n_191;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1705;
wire n_1257;
wire n_171;
wire n_1182;
wire n_579;
wire n_1698;
wire n_1261;
wire n_938;
wire n_1098;
wire n_320;
wire n_1154;
wire n_1242;
wire n_1135;
wire n_406;
wire n_519;
wire n_1016;
wire n_1243;
wire n_546;
wire n_1280;
wire n_281;
wire n_240;
wire n_291;
wire n_231;
wire n_257;
wire n_731;
wire n_371;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_317;
wire n_1236;
wire n_1633;
wire n_569;
wire n_1778;
wire n_227;
wire n_920;
wire n_1289;
wire n_1517;
wire n_335;
wire n_1669;
wire n_370;
wire n_976;
wire n_343;
wire n_1449;
wire n_308;
wire n_1566;
wire n_297;
wire n_1078;
wire n_1670;
wire n_775;
wire n_219;
wire n_600;
wire n_1484;
wire n_1374;
wire n_1328;
wire n_223;
wire n_264;
wire n_1598;
wire n_1723;
wire n_955;
wire n_339;
wire n_1146;
wire n_882;
wire n_183;
wire n_243;
wire n_1097;
wire n_1036;
wire n_1749;
wire n_347;
wire n_550;
wire n_696;
wire n_897;
wire n_215;
wire n_350;
wire n_196;
wire n_798;
wire n_646;
wire n_1428;
wire n_436;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_290;
wire n_580;
wire n_1040;
wire n_578;
wire n_926;
wire n_344;
wire n_1218;
wire n_422;
wire n_475;
wire n_777;
wire n_1070;
wire n_1547;
wire n_1030;
wire n_1755;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_1561;
wire n_496;
wire n_1801;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_1600;
wire n_521;
wire n_663;
wire n_845;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_1796;
wire n_680;
wire n_1473;
wire n_1587;
wire n_395;
wire n_553;
wire n_901;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_214;
wire n_1748;
wire n_1672;
wire n_675;
wire n_888;
wire n_1167;
wire n_1626;
wire n_637;
wire n_1384;
wire n_1556;
wire n_184;
wire n_446;
wire n_1064;
wire n_858;
wire n_923;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_1706;
wire n_468;
wire n_213;
wire n_342;
wire n_464;
wire n_363;
wire n_1582;
wire n_197;
wire n_1069;
wire n_1784;
wire n_1075;
wire n_1450;
wire n_1322;
wire n_1471;
wire n_1750;
wire n_1459;
wire n_460;
wire n_889;
wire n_973;
wire n_1700;
wire n_477;
wire n_571;
wire n_1585;
wire n_461;
wire n_1599;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_907;
wire n_1447;
wire n_1377;
wire n_190;
wire n_989;
wire n_1039;
wire n_228;
wire n_283;
wire n_1403;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_1002;
wire n_1463;
wire n_1581;
wire n_310;
wire n_593;
wire n_748;
wire n_586;
wire n_1058;
wire n_1667;
wire n_838;
wire n_332;
wire n_1053;
wire n_1224;
wire n_349;
wire n_1248;
wire n_230;
wire n_1331;
wire n_953;
wire n_279;
wire n_1014;
wire n_1241;
wire n_289;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_440;
wire n_793;
wire n_478;
wire n_476;
wire n_1527;
wire n_534;
wire n_884;
wire n_345;
wire n_944;
wire n_1754;
wire n_1623;
wire n_1565;
wire n_182;
wire n_647;
wire n_237;
wire n_407;
wire n_1072;
wire n_832;
wire n_857;
wire n_207;
wire n_561;
wire n_1319;
wire n_1712;
wire n_1387;
wire n_1532;
wire n_1027;
wire n_971;
wire n_1156;
wire n_794;
wire n_326;
wire n_404;
wire n_686;
wire n_847;
wire n_1393;
wire n_596;
wire n_1775;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_1709;
wire n_728;
wire n_266;
wire n_1162;
wire n_272;
wire n_1538;
wire n_1199;
wire n_1779;
wire n_352;
wire n_1038;
wire n_520;
wire n_1369;
wire n_409;
wire n_1660;
wire n_887;
wire n_300;
wire n_809;
wire n_931;
wire n_870;
wire n_599;
wire n_1711;
wire n_1662;
wire n_1481;
wire n_434;
wire n_1544;
wire n_868;
wire n_639;
wire n_914;
wire n_411;
wire n_414;
wire n_1629;
wire n_1293;
wire n_965;
wire n_1743;
wire n_935;
wire n_817;
wire n_1175;
wire n_360;
wire n_1479;
wire n_759;
wire n_806;
wire n_1766;
wire n_1477;
wire n_324;
wire n_1635;
wire n_1571;
wire n_187;
wire n_1189;
wire n_1259;
wire n_1690;
wire n_706;
wire n_746;
wire n_1649;
wire n_747;
wire n_784;
wire n_1733;
wire n_1244;
wire n_431;
wire n_1194;
wire n_615;
wire n_851;
wire n_1759;
wire n_843;
wire n_1788;
wire n_523;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_1679;
wire n_776;
wire n_1798;
wire n_1790;
wire n_1415;
wire n_367;
wire n_452;
wire n_525;
wire n_1260;
wire n_1746;
wire n_1647;
wire n_1464;
wire n_649;
wire n_547;
wire n_1444;
wire n_1191;
wire n_1674;
wire n_1710;
wire n_284;
wire n_1128;
wire n_1734;
wire n_744;
wire n_590;
wire n_629;
wire n_1308;
wire n_1767;
wire n_254;
wire n_1680;
wire n_1233;
wire n_1615;
wire n_1529;
wire n_526;
wire n_372;
wire n_293;
wire n_677;
wire n_244;
wire n_1333;
wire n_1121;
wire n_368;
wire n_433;
wire n_314;
wire n_604;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_1001;
wire n_1503;
wire n_498;
wire n_1468;
wire n_1559;
wire n_1765;
wire n_689;
wire n_738;
wire n_1624;
wire n_640;
wire n_1510;
wire n_252;
wire n_624;
wire n_1380;
wire n_1744;
wire n_1617;
wire n_295;
wire n_1010;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_1195;
wire n_610;
wire n_1760;
wire n_936;
wire n_568;
wire n_1500;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_259;
wire n_448;
wire n_758;
wire n_999;
wire n_1656;
wire n_1158;
wire n_1509;
wire n_563;
wire n_1145;
wire n_878;
wire n_524;
wire n_394;
wire n_204;
wire n_1678;
wire n_1049;
wire n_1153;
wire n_741;
wire n_1639;
wire n_1306;
wire n_1068;
wire n_331;
wire n_906;
wire n_1163;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_1781;
wire n_658;
wire n_1740;
wire n_1362;
wire n_1586;
wire n_456;
wire n_959;
wire n_535;
wire n_940;
wire n_1445;
wire n_1492;
wire n_1773;
wire n_592;
wire n_1169;
wire n_1596;
wire n_1692;
wire n_1017;
wire n_978;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_1095;
wire n_1614;
wire n_267;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_603;
wire n_1431;
wire n_484;
wire n_1593;
wire n_1033;
wire n_442;
wire n_636;
wire n_660;
wire n_1640;
wire n_1732;
wire n_1009;
wire n_1148;
wire n_742;
wire n_750;
wire n_995;
wire n_454;
wire n_1609;
wire n_374;
wire n_185;
wire n_396;
wire n_1383;
wire n_1073;
wire n_255;
wire n_662;
wire n_459;
wire n_218;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1065;
wire n_1592;
wire n_1336;
wire n_1721;
wire n_1758;
wire n_1574;
wire n_473;
wire n_1309;
wire n_1426;
wire n_1043;
wire n_355;
wire n_486;
wire n_1800;
wire n_1548;
wire n_614;
wire n_337;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_208;
wire n_743;
wire n_299;
wire n_303;
wire n_296;
wire n_613;
wire n_1119;
wire n_1240;
wire n_829;
wire n_1612;
wire n_1416;
wire n_1724;
wire n_361;
wire n_700;
wire n_1237;
wire n_573;
wire n_1420;
wire n_1132;
wire n_388;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_761;
wire n_1785;
wire n_1568;
wire n_1006;
wire n_329;
wire n_274;
wire n_1270;
wire n_1664;
wire n_1486;
wire n_582;
wire n_1332;
wire n_1390;
wire n_309;
wire n_512;
wire n_1591;
wire n_322;
wire n_1682;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1349;
wire n_1093;
wire n_288;
wire n_1031;
wire n_263;
wire n_609;
wire n_1041;
wire n_1265;
wire n_224;
wire n_1562;
wire n_383;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_239;
wire n_630;
wire n_504;
wire n_511;
wire n_874;
wire n_358;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_1304;
wire n_1324;
wire n_987;
wire n_261;
wire n_174;
wire n_1455;
wire n_767;
wire n_993;
wire n_1407;
wire n_1551;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_1805;
wire n_429;
wire n_948;
wire n_1217;
wire n_628;
wire n_365;
wire n_729;
wire n_1131;
wire n_1084;
wire n_970;
wire n_911;
wire n_1430;
wire n_513;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1534;
wire n_340;
wire n_1351;
wire n_1044;
wire n_1205;
wire n_346;
wire n_1209;
wire n_1552;
wire n_495;
wire n_602;
wire n_574;
wire n_1435;
wire n_879;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_1645;
wire n_490;
wire n_1327;
wire n_996;
wire n_921;
wire n_1684;
wire n_233;
wire n_1717;
wire n_572;
wire n_366;
wire n_815;
wire n_1795;
wire n_327;
wire n_1381;
wire n_1611;
wire n_1037;
wire n_1080;
wire n_1274;
wire n_1316;
wire n_1708;
wire n_426;
wire n_1438;
wire n_1082;
wire n_589;
wire n_716;
wire n_1630;
wire n_562;
wire n_1436;
wire n_1691;
wire n_952;
wire n_1229;
wire n_391;
wire n_701;
wire n_1437;
wire n_1023;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_238;
wire n_1776;
wire n_531;
wire n_1757;
wire n_890;
wire n_764;
wire n_1056;
wire n_1424;
wire n_960;
wire n_222;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_634;
wire n_199;
wire n_1252;
wire n_348;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_1311;
wire n_1519;
wire n_256;
wire n_950;
wire n_1553;
wire n_380;
wire n_419;
wire n_1346;
wire n_444;
wire n_1299;
wire n_1060;
wire n_1141;
wire n_316;
wire n_389;
wire n_418;
wire n_248;
wire n_912;
wire n_315;
wire n_968;
wire n_451;
wire n_619;
wire n_408;
wire n_1386;
wire n_1699;
wire n_376;
wire n_967;
wire n_1442;
wire n_1139;
wire n_515;
wire n_351;
wire n_885;
wire n_397;
wire n_1432;
wire n_1357;
wire n_483;
wire n_683;
wire n_1632;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_1608;
wire n_983;
wire n_280;
wire n_1305;
wire n_873;
wire n_378;
wire n_1112;
wire n_762;
wire n_1283;
wire n_1644;
wire n_690;
wire n_583;
wire n_302;
wire n_1343;
wire n_1203;
wire n_1631;
wire n_821;
wire n_1763;
wire n_1768;
wire n_321;
wire n_1179;
wire n_621;
wire n_753;
wire n_455;
wire n_1048;
wire n_1719;
wire n_1288;
wire n_385;
wire n_212;
wire n_507;
wire n_1560;
wire n_1605;
wire n_330;
wire n_1228;
wire n_972;
wire n_692;
wire n_820;
wire n_1200;
wire n_1301;
wire n_1363;
wire n_1668;
wire n_1185;
wire n_991;
wire n_828;
wire n_779;
wire n_576;
wire n_1143;
wire n_1579;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_537;
wire n_1688;
wire n_945;
wire n_492;
wire n_1504;
wire n_943;
wire n_341;
wire n_250;
wire n_992;
wire n_543;
wire n_260;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_286;
wire n_1643;
wire n_883;
wire n_470;
wire n_449;
wire n_325;
wire n_1594;
wire n_1214;
wire n_1342;
wire n_1400;
wire n_900;
wire n_856;
wire n_1793;
wire n_918;
wire n_942;
wire n_1804;
wire n_189;
wire n_1147;
wire n_1557;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_540;
wire n_618;
wire n_896;
wire n_323;
wire n_195;
wire n_356;
wire n_894;
wire n_1636;
wire n_1730;
wire n_831;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1470;
wire n_1096;
wire n_234;
wire n_1575;
wire n_1697;
wire n_1735;
wire n_833;
wire n_1646;
wire n_225;
wire n_1307;
wire n_988;
wire n_814;
wire n_192;
wire n_1549;
wire n_1201;
wire n_1114;
wire n_655;
wire n_1616;
wire n_1446;
wire n_669;
wire n_472;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_387;
wire n_1149;
wire n_398;
wire n_1671;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_211;
wire n_1219;
wire n_1204;
wire n_178;
wire n_1035;
wire n_287;
wire n_555;
wire n_783;
wire n_1188;
wire n_1722;
wire n_661;
wire n_1802;
wire n_849;
wire n_584;
wire n_681;
wire n_336;
wire n_1638;
wire n_1786;
wire n_430;
wire n_510;
wire n_216;
wire n_311;
wire n_830;
wire n_1296;
wire n_1413;
wire n_801;
wire n_241;
wire n_875;
wire n_357;
wire n_1110;
wire n_1655;
wire n_445;
wire n_749;
wire n_1134;
wire n_1358;
wire n_717;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_249;
wire n_304;
wire n_1338;
wire n_577;
wire n_1522;
wire n_1687;
wire n_1637;
wire n_1419;
wire n_338;
wire n_1653;
wire n_693;
wire n_1506;
wire n_836;
wire n_990;
wire n_1389;
wire n_975;
wire n_1256;
wire n_1702;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_306;
wire n_458;
wire n_770;
wire n_1375;
wire n_1102;
wire n_711;
wire n_1499;
wire n_1187;
wire n_1441;
wire n_1392;
wire n_1597;
wire n_1164;
wire n_1659;
wire n_489;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_1572;
wire n_876;
wire n_1516;
wire n_1190;
wire n_1736;
wire n_1685;
wire n_601;
wire n_917;
wire n_1714;
wire n_966;
wire n_253;
wire n_1116;
wire n_1661;
wire n_1212;
wire n_1541;
wire n_172;
wire n_206;
wire n_217;
wire n_726;
wire n_982;
wire n_1573;
wire n_1453;
wire n_1731;
wire n_818;
wire n_861;
wire n_1713;
wire n_1183;
wire n_1658;
wire n_899;
wire n_1253;
wire n_210;
wire n_1737;
wire n_774;
wire n_1628;
wire n_1335;
wire n_1514;
wire n_1777;
wire n_1059;
wire n_1345;
wire n_176;
wire n_1133;
wire n_1771;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_527;
wire n_1168;
wire n_707;
wire n_937;
wire n_1427;
wire n_393;
wire n_487;
wire n_1584;
wire n_665;
wire n_1726;
wire n_1440;
wire n_177;
wire n_421;
wire n_1356;
wire n_1787;
wire n_910;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1302;
wire n_1774;
wire n_1725;
wire n_205;
wire n_1136;
wire n_1313;
wire n_1491;
wire n_754;
wire n_1496;
wire n_179;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_735;
wire n_232;
wire n_1109;
wire n_895;
wire n_1310;
wire n_1803;
wire n_202;
wire n_427;
wire n_1399;
wire n_1543;
wire n_791;
wire n_732;
wire n_1533;
wire n_193;
wire n_808;
wire n_797;
wire n_1025;
wire n_500;
wire n_1067;
wire n_1720;
wire n_435;
wire n_766;
wire n_1457;
wire n_541;
wire n_538;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1742;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_594;
wire n_200;
wire n_1291;
wire n_1297;
wire n_1753;
wire n_1782;
wire n_1155;
wire n_1418;
wire n_1524;
wire n_1689;
wire n_1485;
wire n_1011;
wire n_1184;
wire n_985;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_1703;
wire n_1352;
wire n_626;
wire n_1650;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_1170;
wire n_305;
wire n_676;
wire n_294;
wire n_318;
wire n_653;
wire n_642;
wire n_1602;
wire n_194;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_268;
wire n_664;
wire n_503;
wire n_235;
wire n_1372;
wire n_605;
wire n_1273;
wire n_353;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_1282;
wire n_1318;
wire n_1783;
wire n_780;
wire n_998;
wire n_1454;
wire n_467;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_501;
wire n_823;
wire n_245;
wire n_725;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_672;
wire n_581;
wire n_382;
wire n_554;
wire n_1625;
wire n_898;
wire n_1762;
wire n_1013;
wire n_1452;
wire n_718;
wire n_265;
wire n_1120;
wire n_719;
wire n_443;
wire n_1791;
wire n_198;
wire n_1747;
wire n_714;
wire n_1683;
wire n_909;
wire n_1530;
wire n_1497;
wire n_997;
wire n_932;
wire n_612;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_508;
wire n_506;
wire n_1320;
wire n_1663;
wire n_737;
wire n_1718;
wire n_986;
wire n_509;
wire n_1317;
wire n_1715;
wire n_1518;
wire n_1281;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_209;
wire n_1792;
wire n_1564;
wire n_1613;
wire n_733;
wire n_1489;
wire n_1376;
wire n_941;
wire n_981;
wire n_1569;
wire n_867;
wire n_186;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_298;
wire n_518;
wire n_505;
wire n_1772;
wire n_282;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1620;
wire n_381;
wire n_220;
wire n_390;
wire n_1330;
wire n_481;
wire n_1675;
wire n_1727;
wire n_1554;
wire n_1745;
wire n_769;
wire n_1046;
wire n_271;
wire n_934;
wire n_1618;
wire n_826;
wire n_886;
wire n_1221;
wire n_654;
wire n_1172;
wire n_379;
wire n_428;
wire n_1341;
wire n_570;
wire n_1641;
wire n_1361;
wire n_1707;
wire n_853;
wire n_377;
wire n_751;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_392;
wire n_704;
wire n_787;
wire n_1770;
wire n_961;
wire n_1756;
wire n_771;
wire n_276;
wire n_1716;
wire n_1225;
wire n_1520;
wire n_169;
wire n_522;
wire n_1287;
wire n_1262;
wire n_400;
wire n_930;
wire n_181;
wire n_1411;
wire n_221;
wire n_622;
wire n_1577;
wire n_1087;
wire n_386;
wire n_994;
wire n_1701;
wire n_848;
wire n_1550;
wire n_1498;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1567;
wire n_1247;
wire n_922;
wire n_816;
wire n_1648;
wire n_591;
wire n_1536;
wire n_1344;
wire n_313;
wire n_631;
wire n_479;
wire n_1246;
wire n_1478;
wire n_1339;
wire n_1797;
wire n_432;
wire n_1769;
wire n_839;
wire n_1210;
wire n_1364;
wire n_328;
wire n_1250;
wire n_369;
wire n_871;
wire n_598;
wire n_685;
wire n_928;
wire n_608;
wire n_1367;
wire n_1460;
wire n_772;
wire n_1555;
wire n_499;
wire n_1589;
wire n_517;
wire n_413;
wire n_402;
wire n_1086;
wire n_796;
wire n_1619;
wire n_236;
wire n_1502;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_903;
wire n_1525;
wire n_1752;
wire n_740;
wire n_203;
wire n_384;
wire n_1404;
wire n_1794;
wire n_1315;
wire n_277;
wire n_1061;
wire n_333;
wire n_1298;
wire n_1652;
wire n_462;
wire n_1193;
wire n_1676;
wire n_1255;
wire n_258;
wire n_1113;
wire n_1226;
wire n_722;
wire n_1277;
wire n_188;
wire n_844;
wire n_201;
wire n_471;
wire n_852;
wire n_1487;
wire n_1028;
wire n_1601;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_1546;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_1627;
wire n_1245;
wire n_846;
wire n_1673;
wire n_465;
wire n_362;
wire n_1321;
wire n_170;
wire n_273;
wire n_585;
wire n_1739;
wire n_270;
wire n_616;
wire n_745;
wire n_1654;
wire n_1103;
wire n_648;
wire n_1379;
wire n_312;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_494;
wire n_1761;
wire n_641;
wire n_730;
wire n_1325;
wire n_1595;
wire n_354;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_695;
wire n_180;
wire n_656;
wire n_1606;
wire n_1220;
wire n_1694;
wire n_1540;
wire n_229;
wire n_437;
wire n_1642;
wire n_403;
wire n_453;
wire n_1130;
wire n_720;
wire n_1526;
wire n_863;
wire n_805;
wire n_1604;
wire n_1275;
wire n_1764;
wire n_712;
wire n_246;
wire n_1583;
wire n_1042;
wire n_1402;
wire n_269;
wire n_285;
wire n_412;
wire n_1493;
wire n_657;
wire n_644;
wire n_1741;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_1621;
wire n_251;
wire n_566;
wire n_565;
wire n_1448;
wire n_1507;
wire n_1398;
wire n_597;
wire n_1181;
wire n_1505;
wire n_1634;
wire n_1196;
wire n_651;
wire n_1340;
wire n_334;
wire n_811;
wire n_1558;
wire n_807;
wire n_835;
wire n_175;
wire n_666;
wire n_262;
wire n_1433;
wire n_1704;
wire n_1254;
wire n_1026;
wire n_1234;
wire n_319;
wire n_364;
wire n_1138;
wire n_927;
wire n_1089;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_242;
wire n_1681;
wire n_1018;
wire n_1693;
wire n_438;
wire n_713;
wire n_904;
wire n_1588;
wire n_1622;
wire n_1180;
wire n_1271;
wire n_533;
wire n_1542;
wire n_1251;
wire n_278;

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_3),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_72),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_68),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_51),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_163),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_26),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_37),
.Y(n_175)
);

BUFx3_ASAP7_75t_L g176 ( 
.A(n_118),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_101),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_162),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_37),
.Y(n_179)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_85),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_69),
.Y(n_181)
);

INVxp67_ASAP7_75t_L g182 ( 
.A(n_25),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_120),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_49),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_90),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_112),
.Y(n_186)
);

BUFx3_ASAP7_75t_L g187 ( 
.A(n_44),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_51),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_38),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_123),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_1),
.Y(n_191)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_61),
.Y(n_192)
);

INVx2_ASAP7_75t_SL g193 ( 
.A(n_17),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_148),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_57),
.Y(n_195)
);

CKINVDCx16_ASAP7_75t_R g196 ( 
.A(n_31),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_53),
.Y(n_197)
);

BUFx3_ASAP7_75t_L g198 ( 
.A(n_60),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_150),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_166),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_30),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_56),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_75),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_1),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_16),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_117),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_151),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_40),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_95),
.Y(n_209)
);

BUFx2_ASAP7_75t_L g210 ( 
.A(n_18),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_33),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_41),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_19),
.Y(n_213)
);

BUFx6f_ASAP7_75t_L g214 ( 
.A(n_92),
.Y(n_214)
);

CKINVDCx16_ASAP7_75t_R g215 ( 
.A(n_107),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_89),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_136),
.Y(n_217)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_88),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_44),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_70),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_141),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_87),
.Y(n_222)
);

INVx1_ASAP7_75t_SL g223 ( 
.A(n_64),
.Y(n_223)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_63),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_31),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_111),
.Y(n_226)
);

BUFx3_ASAP7_75t_L g227 ( 
.A(n_9),
.Y(n_227)
);

CKINVDCx14_ASAP7_75t_R g228 ( 
.A(n_99),
.Y(n_228)
);

BUFx2_ASAP7_75t_L g229 ( 
.A(n_114),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_158),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_5),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_130),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_7),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_124),
.Y(n_234)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_29),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_35),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_59),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_108),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_128),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_140),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_53),
.Y(n_241)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_155),
.Y(n_242)
);

BUFx10_ASAP7_75t_L g243 ( 
.A(n_160),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_125),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_131),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_122),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_45),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_49),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_137),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_25),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_115),
.Y(n_251)
);

BUFx2_ASAP7_75t_L g252 ( 
.A(n_10),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_50),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_23),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_109),
.Y(n_255)
);

BUFx5_ASAP7_75t_L g256 ( 
.A(n_152),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_116),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_134),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_98),
.Y(n_259)
);

BUFx3_ASAP7_75t_L g260 ( 
.A(n_67),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_26),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_119),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_102),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_43),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_146),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_22),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_127),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_82),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_74),
.Y(n_269)
);

INVxp67_ASAP7_75t_L g270 ( 
.A(n_100),
.Y(n_270)
);

INVx2_ASAP7_75t_SL g271 ( 
.A(n_41),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_103),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_161),
.Y(n_273)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_50),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_22),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_78),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_45),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_35),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_38),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_153),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_8),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_126),
.Y(n_282)
);

BUFx6f_ASAP7_75t_L g283 ( 
.A(n_4),
.Y(n_283)
);

INVx1_ASAP7_75t_SL g284 ( 
.A(n_65),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_19),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_28),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_33),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_157),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g289 ( 
.A(n_34),
.Y(n_289)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_86),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_39),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_13),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_139),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_52),
.Y(n_294)
);

BUFx5_ASAP7_75t_L g295 ( 
.A(n_28),
.Y(n_295)
);

INVx2_ASAP7_75t_L g296 ( 
.A(n_29),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_135),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_73),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_104),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_156),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_15),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_12),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_16),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_12),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_57),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g306 ( 
.A(n_143),
.Y(n_306)
);

INVx3_ASAP7_75t_L g307 ( 
.A(n_39),
.Y(n_307)
);

HB1xp67_ASAP7_75t_L g308 ( 
.A(n_10),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_154),
.Y(n_309)
);

CKINVDCx16_ASAP7_75t_R g310 ( 
.A(n_48),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_18),
.Y(n_311)
);

BUFx10_ASAP7_75t_L g312 ( 
.A(n_77),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_58),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_164),
.Y(n_314)
);

CKINVDCx20_ASAP7_75t_R g315 ( 
.A(n_80),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_54),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_9),
.Y(n_317)
);

INVx2_ASAP7_75t_L g318 ( 
.A(n_133),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_4),
.Y(n_319)
);

BUFx3_ASAP7_75t_L g320 ( 
.A(n_54),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_147),
.Y(n_321)
);

INVx2_ASAP7_75t_L g322 ( 
.A(n_20),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_13),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_129),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_159),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_34),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_81),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_83),
.Y(n_328)
);

CKINVDCx16_ASAP7_75t_R g329 ( 
.A(n_40),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_48),
.Y(n_330)
);

BUFx3_ASAP7_75t_L g331 ( 
.A(n_94),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_42),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_6),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g334 ( 
.A(n_24),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_23),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_46),
.Y(n_336)
);

INVx1_ASAP7_75t_SL g337 ( 
.A(n_17),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_8),
.Y(n_338)
);

CKINVDCx20_ASAP7_75t_R g339 ( 
.A(n_221),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_216),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_295),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_217),
.Y(n_342)
);

HB1xp67_ASAP7_75t_L g343 ( 
.A(n_196),
.Y(n_343)
);

INVxp33_ASAP7_75t_L g344 ( 
.A(n_308),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_220),
.Y(n_345)
);

NOR2xp33_ASAP7_75t_L g346 ( 
.A(n_229),
.B(n_0),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_295),
.Y(n_347)
);

INVxp67_ASAP7_75t_L g348 ( 
.A(n_210),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_295),
.Y(n_349)
);

INVx2_ASAP7_75t_L g350 ( 
.A(n_295),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_222),
.Y(n_351)
);

AND2x2_ASAP7_75t_L g352 ( 
.A(n_252),
.B(n_0),
.Y(n_352)
);

INVxp67_ASAP7_75t_SL g353 ( 
.A(n_307),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_295),
.Y(n_354)
);

INVx2_ASAP7_75t_L g355 ( 
.A(n_295),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_226),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_230),
.Y(n_357)
);

INVxp33_ASAP7_75t_L g358 ( 
.A(n_172),
.Y(n_358)
);

CKINVDCx20_ASAP7_75t_R g359 ( 
.A(n_238),
.Y(n_359)
);

CKINVDCx20_ASAP7_75t_R g360 ( 
.A(n_245),
.Y(n_360)
);

CKINVDCx20_ASAP7_75t_R g361 ( 
.A(n_306),
.Y(n_361)
);

CKINVDCx16_ASAP7_75t_R g362 ( 
.A(n_310),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_234),
.Y(n_363)
);

HB1xp67_ASAP7_75t_L g364 ( 
.A(n_329),
.Y(n_364)
);

CKINVDCx20_ASAP7_75t_R g365 ( 
.A(n_315),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_307),
.B(n_2),
.Y(n_366)
);

CKINVDCx20_ASAP7_75t_R g367 ( 
.A(n_215),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_239),
.Y(n_368)
);

HB1xp67_ASAP7_75t_L g369 ( 
.A(n_169),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_240),
.Y(n_370)
);

BUFx6f_ASAP7_75t_L g371 ( 
.A(n_214),
.Y(n_371)
);

NOR2xp67_ASAP7_75t_L g372 ( 
.A(n_307),
.B(n_2),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_295),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_295),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_283),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_283),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_246),
.Y(n_377)
);

INVx1_ASAP7_75t_SL g378 ( 
.A(n_337),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_283),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_283),
.Y(n_380)
);

CKINVDCx20_ASAP7_75t_R g381 ( 
.A(n_228),
.Y(n_381)
);

CKINVDCx20_ASAP7_75t_R g382 ( 
.A(n_249),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_251),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_259),
.Y(n_384)
);

INVxp67_ASAP7_75t_L g385 ( 
.A(n_193),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_283),
.Y(n_386)
);

INVxp67_ASAP7_75t_SL g387 ( 
.A(n_176),
.Y(n_387)
);

HB1xp67_ASAP7_75t_L g388 ( 
.A(n_169),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_235),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_235),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_265),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_274),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_274),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_268),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_296),
.Y(n_395)
);

INVxp67_ASAP7_75t_SL g396 ( 
.A(n_176),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_296),
.Y(n_397)
);

INVxp67_ASAP7_75t_L g398 ( 
.A(n_193),
.Y(n_398)
);

INVxp67_ASAP7_75t_SL g399 ( 
.A(n_198),
.Y(n_399)
);

CKINVDCx20_ASAP7_75t_R g400 ( 
.A(n_269),
.Y(n_400)
);

NOR2xp33_ASAP7_75t_L g401 ( 
.A(n_270),
.B(n_180),
.Y(n_401)
);

CKINVDCx20_ASAP7_75t_R g402 ( 
.A(n_273),
.Y(n_402)
);

INVx1_ASAP7_75t_SL g403 ( 
.A(n_231),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_322),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_322),
.Y(n_405)
);

CKINVDCx20_ASAP7_75t_R g406 ( 
.A(n_276),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_187),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_187),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_297),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_227),
.Y(n_410)
);

HB1xp67_ASAP7_75t_L g411 ( 
.A(n_174),
.Y(n_411)
);

HB1xp67_ASAP7_75t_L g412 ( 
.A(n_174),
.Y(n_412)
);

CKINVDCx14_ASAP7_75t_R g413 ( 
.A(n_243),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_227),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_320),
.Y(n_415)
);

INVxp67_ASAP7_75t_SL g416 ( 
.A(n_198),
.Y(n_416)
);

CKINVDCx20_ASAP7_75t_R g417 ( 
.A(n_298),
.Y(n_417)
);

NOR2xp67_ASAP7_75t_L g418 ( 
.A(n_271),
.B(n_3),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_320),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_225),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_175),
.Y(n_421)
);

AND2x2_ASAP7_75t_L g422 ( 
.A(n_353),
.B(n_260),
.Y(n_422)
);

INVx1_ASAP7_75t_SL g423 ( 
.A(n_378),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_375),
.Y(n_424)
);

AND2x2_ASAP7_75t_L g425 ( 
.A(n_387),
.B(n_260),
.Y(n_425)
);

AND2x2_ASAP7_75t_L g426 ( 
.A(n_396),
.B(n_331),
.Y(n_426)
);

AND2x2_ASAP7_75t_L g427 ( 
.A(n_399),
.B(n_331),
.Y(n_427)
);

INVx2_ASAP7_75t_L g428 ( 
.A(n_350),
.Y(n_428)
);

INVx2_ASAP7_75t_L g429 ( 
.A(n_350),
.Y(n_429)
);

INVx2_ASAP7_75t_L g430 ( 
.A(n_350),
.Y(n_430)
);

INVx3_ASAP7_75t_L g431 ( 
.A(n_371),
.Y(n_431)
);

OAI21x1_ASAP7_75t_L g432 ( 
.A1(n_355),
.A2(n_192),
.B(n_180),
.Y(n_432)
);

INVx2_ASAP7_75t_L g433 ( 
.A(n_355),
.Y(n_433)
);

INVx2_ASAP7_75t_L g434 ( 
.A(n_355),
.Y(n_434)
);

BUFx6f_ASAP7_75t_L g435 ( 
.A(n_371),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_L g436 ( 
.A(n_341),
.B(n_192),
.Y(n_436)
);

INVx2_ASAP7_75t_L g437 ( 
.A(n_371),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_375),
.Y(n_438)
);

BUFx6f_ASAP7_75t_L g439 ( 
.A(n_371),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_376),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_376),
.Y(n_441)
);

INVx2_ASAP7_75t_L g442 ( 
.A(n_371),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_379),
.Y(n_443)
);

INVx2_ASAP7_75t_L g444 ( 
.A(n_371),
.Y(n_444)
);

AND2x4_ASAP7_75t_L g445 ( 
.A(n_372),
.B(n_218),
.Y(n_445)
);

INVx2_ASAP7_75t_L g446 ( 
.A(n_341),
.Y(n_446)
);

INVxp67_ASAP7_75t_L g447 ( 
.A(n_378),
.Y(n_447)
);

OA21x2_ASAP7_75t_L g448 ( 
.A1(n_366),
.A2(n_184),
.B(n_179),
.Y(n_448)
);

OR2x6_ASAP7_75t_L g449 ( 
.A(n_366),
.B(n_372),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_401),
.B(n_170),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_379),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_416),
.B(n_170),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_380),
.Y(n_453)
);

HB1xp67_ASAP7_75t_L g454 ( 
.A(n_343),
.Y(n_454)
);

INVx2_ASAP7_75t_L g455 ( 
.A(n_347),
.Y(n_455)
);

HB1xp67_ASAP7_75t_L g456 ( 
.A(n_364),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_380),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_386),
.B(n_171),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_386),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_347),
.B(n_218),
.Y(n_460)
);

NOR2xp33_ASAP7_75t_L g461 ( 
.A(n_346),
.B(n_223),
.Y(n_461)
);

INVx3_ASAP7_75t_L g462 ( 
.A(n_349),
.Y(n_462)
);

INVx2_ASAP7_75t_L g463 ( 
.A(n_349),
.Y(n_463)
);

INVx3_ASAP7_75t_L g464 ( 
.A(n_354),
.Y(n_464)
);

INVx2_ASAP7_75t_L g465 ( 
.A(n_354),
.Y(n_465)
);

BUFx3_ASAP7_75t_L g466 ( 
.A(n_373),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_373),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_374),
.Y(n_468)
);

CKINVDCx5p33_ASAP7_75t_R g469 ( 
.A(n_382),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_374),
.Y(n_470)
);

INVx2_ASAP7_75t_L g471 ( 
.A(n_389),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_389),
.Y(n_472)
);

BUFx6f_ASAP7_75t_L g473 ( 
.A(n_390),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_407),
.B(n_171),
.Y(n_474)
);

INVx2_ASAP7_75t_L g475 ( 
.A(n_390),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_392),
.B(n_224),
.Y(n_476)
);

BUFx6f_ASAP7_75t_L g477 ( 
.A(n_392),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_393),
.Y(n_478)
);

INVx3_ASAP7_75t_L g479 ( 
.A(n_393),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_L g480 ( 
.A(n_407),
.B(n_178),
.Y(n_480)
);

OAI22xp5_ASAP7_75t_L g481 ( 
.A1(n_348),
.A2(n_289),
.B1(n_294),
.B2(n_233),
.Y(n_481)
);

AND2x4_ASAP7_75t_L g482 ( 
.A(n_418),
.B(n_224),
.Y(n_482)
);

INVx2_ASAP7_75t_L g483 ( 
.A(n_395),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_SL g484 ( 
.A(n_352),
.B(n_243),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_395),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_397),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_L g487 ( 
.A(n_397),
.B(n_242),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_404),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_404),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_405),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_L g491 ( 
.A(n_408),
.B(n_178),
.Y(n_491)
);

INVx2_ASAP7_75t_L g492 ( 
.A(n_405),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_421),
.Y(n_493)
);

INVx2_ASAP7_75t_L g494 ( 
.A(n_421),
.Y(n_494)
);

AND2x2_ASAP7_75t_L g495 ( 
.A(n_408),
.B(n_242),
.Y(n_495)
);

BUFx6f_ASAP7_75t_L g496 ( 
.A(n_410),
.Y(n_496)
);

AND2x2_ASAP7_75t_SL g497 ( 
.A(n_352),
.B(n_290),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_L g498 ( 
.A(n_497),
.B(n_340),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_L g499 ( 
.A(n_497),
.B(n_342),
.Y(n_499)
);

AND2x6_ASAP7_75t_L g500 ( 
.A(n_445),
.B(n_290),
.Y(n_500)
);

NAND2xp33_ASAP7_75t_L g501 ( 
.A(n_450),
.B(n_345),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_467),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_467),
.Y(n_503)
);

INVxp67_ASAP7_75t_SL g504 ( 
.A(n_447),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_L g505 ( 
.A(n_497),
.B(n_351),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_SL g506 ( 
.A(n_423),
.B(n_356),
.Y(n_506)
);

INVx2_ASAP7_75t_SL g507 ( 
.A(n_423),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_467),
.Y(n_508)
);

INVx2_ASAP7_75t_L g509 ( 
.A(n_428),
.Y(n_509)
);

BUFx3_ASAP7_75t_L g510 ( 
.A(n_466),
.Y(n_510)
);

INVx2_ASAP7_75t_L g511 ( 
.A(n_428),
.Y(n_511)
);

INVx4_ASAP7_75t_L g512 ( 
.A(n_449),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_L g513 ( 
.A(n_497),
.B(n_357),
.Y(n_513)
);

BUFx3_ASAP7_75t_L g514 ( 
.A(n_466),
.Y(n_514)
);

INVx2_ASAP7_75t_L g515 ( 
.A(n_428),
.Y(n_515)
);

INVx3_ASAP7_75t_L g516 ( 
.A(n_435),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_468),
.Y(n_517)
);

INVx2_ASAP7_75t_L g518 ( 
.A(n_428),
.Y(n_518)
);

INVx2_ASAP7_75t_L g519 ( 
.A(n_429),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_SL g520 ( 
.A(n_423),
.B(n_363),
.Y(n_520)
);

INVx2_ASAP7_75t_L g521 ( 
.A(n_429),
.Y(n_521)
);

BUFx3_ASAP7_75t_L g522 ( 
.A(n_466),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_L g523 ( 
.A(n_497),
.B(n_368),
.Y(n_523)
);

INVx4_ASAP7_75t_L g524 ( 
.A(n_449),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_468),
.Y(n_525)
);

NOR2xp33_ASAP7_75t_L g526 ( 
.A(n_461),
.B(n_370),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_468),
.Y(n_527)
);

INVx4_ASAP7_75t_SL g528 ( 
.A(n_449),
.Y(n_528)
);

INVx2_ASAP7_75t_L g529 ( 
.A(n_429),
.Y(n_529)
);

INVx2_ASAP7_75t_L g530 ( 
.A(n_429),
.Y(n_530)
);

NOR2xp33_ASAP7_75t_L g531 ( 
.A(n_461),
.B(n_377),
.Y(n_531)
);

CKINVDCx16_ASAP7_75t_R g532 ( 
.A(n_454),
.Y(n_532)
);

NOR2xp33_ASAP7_75t_L g533 ( 
.A(n_450),
.B(n_383),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_470),
.Y(n_534)
);

NOR2xp33_ASAP7_75t_L g535 ( 
.A(n_484),
.B(n_384),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_SL g536 ( 
.A(n_447),
.B(n_391),
.Y(n_536)
);

INVx2_ASAP7_75t_L g537 ( 
.A(n_430),
.Y(n_537)
);

INVx2_ASAP7_75t_L g538 ( 
.A(n_430),
.Y(n_538)
);

INVx2_ASAP7_75t_L g539 ( 
.A(n_430),
.Y(n_539)
);

NOR2xp33_ASAP7_75t_L g540 ( 
.A(n_484),
.B(n_394),
.Y(n_540)
);

INVx3_ASAP7_75t_L g541 ( 
.A(n_435),
.Y(n_541)
);

BUFx6f_ASAP7_75t_L g542 ( 
.A(n_435),
.Y(n_542)
);

BUFx2_ASAP7_75t_L g543 ( 
.A(n_454),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_470),
.Y(n_544)
);

INVx1_ASAP7_75t_SL g545 ( 
.A(n_469),
.Y(n_545)
);

INVx5_ASAP7_75t_L g546 ( 
.A(n_435),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_L g547 ( 
.A(n_466),
.B(n_409),
.Y(n_547)
);

INVx2_ASAP7_75t_L g548 ( 
.A(n_430),
.Y(n_548)
);

INVx4_ASAP7_75t_L g549 ( 
.A(n_449),
.Y(n_549)
);

NOR2xp33_ASAP7_75t_L g550 ( 
.A(n_452),
.B(n_420),
.Y(n_550)
);

AND2x2_ASAP7_75t_L g551 ( 
.A(n_425),
.B(n_410),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_470),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_462),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_462),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_462),
.Y(n_555)
);

INVx2_ASAP7_75t_L g556 ( 
.A(n_433),
.Y(n_556)
);

AND2x2_ASAP7_75t_L g557 ( 
.A(n_425),
.B(n_414),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_462),
.Y(n_558)
);

OAI22xp5_ASAP7_75t_L g559 ( 
.A1(n_449),
.A2(n_381),
.B1(n_400),
.B2(n_417),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_462),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_462),
.Y(n_561)
);

INVx2_ASAP7_75t_L g562 ( 
.A(n_433),
.Y(n_562)
);

INVx2_ASAP7_75t_L g563 ( 
.A(n_433),
.Y(n_563)
);

NAND2xp33_ASAP7_75t_SL g564 ( 
.A(n_456),
.B(n_367),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_L g565 ( 
.A(n_425),
.B(n_413),
.Y(n_565)
);

INVx2_ASAP7_75t_L g566 ( 
.A(n_433),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_L g567 ( 
.A(n_425),
.B(n_284),
.Y(n_567)
);

INVxp67_ASAP7_75t_SL g568 ( 
.A(n_464),
.Y(n_568)
);

AOI22xp33_ASAP7_75t_L g569 ( 
.A1(n_449),
.A2(n_418),
.B1(n_271),
.B2(n_344),
.Y(n_569)
);

AND2x4_ASAP7_75t_L g570 ( 
.A(n_445),
.B(n_318),
.Y(n_570)
);

BUFx3_ASAP7_75t_L g571 ( 
.A(n_448),
.Y(n_571)
);

NOR2xp33_ASAP7_75t_L g572 ( 
.A(n_452),
.B(n_402),
.Y(n_572)
);

INVx2_ASAP7_75t_L g573 ( 
.A(n_434),
.Y(n_573)
);

AOI22xp33_ASAP7_75t_L g574 ( 
.A1(n_449),
.A2(n_445),
.B1(n_482),
.B2(n_448),
.Y(n_574)
);

INVx2_ASAP7_75t_L g575 ( 
.A(n_434),
.Y(n_575)
);

INVx3_ASAP7_75t_L g576 ( 
.A(n_435),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_L g577 ( 
.A(n_426),
.B(n_173),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_L g578 ( 
.A(n_426),
.B(n_177),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_SL g579 ( 
.A(n_426),
.B(n_362),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_SL g580 ( 
.A(n_427),
.B(n_362),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_464),
.Y(n_581)
);

INVxp33_ASAP7_75t_SL g582 ( 
.A(n_469),
.Y(n_582)
);

OR2x2_ASAP7_75t_L g583 ( 
.A(n_456),
.B(n_403),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_L g584 ( 
.A(n_427),
.B(n_232),
.Y(n_584)
);

INVx3_ASAP7_75t_L g585 ( 
.A(n_435),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_L g586 ( 
.A(n_427),
.B(n_237),
.Y(n_586)
);

INVx3_ASAP7_75t_L g587 ( 
.A(n_435),
.Y(n_587)
);

INVx2_ASAP7_75t_SL g588 ( 
.A(n_427),
.Y(n_588)
);

AO21x2_ASAP7_75t_L g589 ( 
.A1(n_432),
.A2(n_255),
.B(n_244),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_L g590 ( 
.A(n_422),
.B(n_257),
.Y(n_590)
);

AND2x2_ASAP7_75t_L g591 ( 
.A(n_422),
.B(n_414),
.Y(n_591)
);

AOI22xp33_ASAP7_75t_L g592 ( 
.A1(n_449),
.A2(n_445),
.B1(n_482),
.B2(n_448),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_464),
.Y(n_593)
);

BUFx10_ASAP7_75t_L g594 ( 
.A(n_445),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_464),
.Y(n_595)
);

INVx2_ASAP7_75t_L g596 ( 
.A(n_434),
.Y(n_596)
);

INVx5_ASAP7_75t_L g597 ( 
.A(n_435),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_L g598 ( 
.A(n_422),
.B(n_258),
.Y(n_598)
);

INVx3_ASAP7_75t_L g599 ( 
.A(n_435),
.Y(n_599)
);

INVx2_ASAP7_75t_SL g600 ( 
.A(n_422),
.Y(n_600)
);

INVx2_ASAP7_75t_L g601 ( 
.A(n_434),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_464),
.Y(n_602)
);

BUFx4f_ASAP7_75t_L g603 ( 
.A(n_448),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_446),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_446),
.Y(n_605)
);

INVx3_ASAP7_75t_L g606 ( 
.A(n_439),
.Y(n_606)
);

AOI22xp33_ASAP7_75t_L g607 ( 
.A1(n_445),
.A2(n_236),
.B1(n_189),
.B2(n_205),
.Y(n_607)
);

INVx2_ASAP7_75t_L g608 ( 
.A(n_446),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_446),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_455),
.Y(n_610)
);

INVx3_ASAP7_75t_L g611 ( 
.A(n_439),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_455),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_455),
.Y(n_613)
);

INVx4_ASAP7_75t_L g614 ( 
.A(n_496),
.Y(n_614)
);

INVxp33_ASAP7_75t_SL g615 ( 
.A(n_481),
.Y(n_615)
);

INVx2_ASAP7_75t_L g616 ( 
.A(n_455),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_463),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_463),
.Y(n_618)
);

INVx2_ASAP7_75t_L g619 ( 
.A(n_463),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_L g620 ( 
.A(n_482),
.B(n_262),
.Y(n_620)
);

INVx2_ASAP7_75t_L g621 ( 
.A(n_463),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_465),
.Y(n_622)
);

NOR2xp33_ASAP7_75t_L g623 ( 
.A(n_474),
.B(n_406),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_SL g624 ( 
.A(n_474),
.B(n_243),
.Y(n_624)
);

INVx2_ASAP7_75t_SL g625 ( 
.A(n_448),
.Y(n_625)
);

INVx4_ASAP7_75t_SL g626 ( 
.A(n_439),
.Y(n_626)
);

INVx2_ASAP7_75t_L g627 ( 
.A(n_465),
.Y(n_627)
);

INVx6_ASAP7_75t_L g628 ( 
.A(n_482),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_465),
.Y(n_629)
);

OAI22xp5_ASAP7_75t_L g630 ( 
.A1(n_480),
.A2(n_182),
.B1(n_264),
.B2(n_286),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_SL g631 ( 
.A(n_480),
.B(n_312),
.Y(n_631)
);

INVx3_ASAP7_75t_L g632 ( 
.A(n_439),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_SL g633 ( 
.A(n_491),
.B(n_312),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_L g634 ( 
.A(n_482),
.B(n_458),
.Y(n_634)
);

INVx2_ASAP7_75t_SL g635 ( 
.A(n_448),
.Y(n_635)
);

INVx2_ASAP7_75t_SL g636 ( 
.A(n_448),
.Y(n_636)
);

INVx2_ASAP7_75t_L g637 ( 
.A(n_465),
.Y(n_637)
);

INVx6_ASAP7_75t_L g638 ( 
.A(n_482),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_424),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_L g640 ( 
.A(n_458),
.B(n_263),
.Y(n_640)
);

AOI22xp33_ASAP7_75t_L g641 ( 
.A1(n_495),
.A2(n_291),
.B1(n_213),
.B2(n_219),
.Y(n_641)
);

INVx3_ASAP7_75t_L g642 ( 
.A(n_439),
.Y(n_642)
);

INVx2_ASAP7_75t_L g643 ( 
.A(n_432),
.Y(n_643)
);

NOR3xp33_ASAP7_75t_L g644 ( 
.A(n_481),
.B(n_403),
.C(n_388),
.Y(n_644)
);

INVx2_ASAP7_75t_L g645 ( 
.A(n_432),
.Y(n_645)
);

INVxp67_ASAP7_75t_SL g646 ( 
.A(n_431),
.Y(n_646)
);

OAI22xp5_ASAP7_75t_L g647 ( 
.A1(n_491),
.A2(n_287),
.B1(n_241),
.B2(n_250),
.Y(n_647)
);

AOI22xp5_ASAP7_75t_L g648 ( 
.A1(n_481),
.A2(n_316),
.B1(n_333),
.B2(n_334),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_SL g649 ( 
.A(n_594),
.B(n_496),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_L g650 ( 
.A(n_533),
.B(n_496),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_L g651 ( 
.A(n_600),
.B(n_496),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_507),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_L g653 ( 
.A(n_600),
.B(n_496),
.Y(n_653)
);

INVx2_ASAP7_75t_L g654 ( 
.A(n_502),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_L g655 ( 
.A(n_588),
.B(n_550),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_507),
.Y(n_656)
);

INVx2_ASAP7_75t_L g657 ( 
.A(n_502),
.Y(n_657)
);

INVxp67_ASAP7_75t_L g658 ( 
.A(n_504),
.Y(n_658)
);

NOR2xp33_ASAP7_75t_L g659 ( 
.A(n_526),
.B(n_369),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_L g660 ( 
.A(n_588),
.B(n_496),
.Y(n_660)
);

OAI22xp5_ASAP7_75t_L g661 ( 
.A1(n_574),
.A2(n_365),
.B1(n_361),
.B2(n_360),
.Y(n_661)
);

OAI221xp5_ASAP7_75t_L g662 ( 
.A1(n_569),
.A2(n_278),
.B1(n_311),
.B2(n_303),
.C(n_301),
.Y(n_662)
);

INVx2_ASAP7_75t_L g663 ( 
.A(n_503),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_639),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_SL g665 ( 
.A(n_594),
.B(n_496),
.Y(n_665)
);

AOI22xp5_ASAP7_75t_L g666 ( 
.A1(n_498),
.A2(n_359),
.B1(n_339),
.B2(n_495),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_SL g667 ( 
.A(n_594),
.B(n_496),
.Y(n_667)
);

OAI22xp5_ASAP7_75t_L g668 ( 
.A1(n_592),
.A2(n_272),
.B1(n_267),
.B2(n_280),
.Y(n_668)
);

AO22x2_ASAP7_75t_L g669 ( 
.A1(n_644),
.A2(n_208),
.B1(n_248),
.B2(n_253),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_L g670 ( 
.A(n_531),
.B(n_496),
.Y(n_670)
);

CKINVDCx5p33_ASAP7_75t_R g671 ( 
.A(n_582),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_639),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_SL g673 ( 
.A(n_594),
.B(n_603),
.Y(n_673)
);

INVx2_ASAP7_75t_SL g674 ( 
.A(n_583),
.Y(n_674)
);

NOR2xp33_ASAP7_75t_L g675 ( 
.A(n_499),
.B(n_411),
.Y(n_675)
);

AO22x2_ASAP7_75t_L g676 ( 
.A1(n_625),
.A2(n_254),
.B1(n_281),
.B2(n_313),
.Y(n_676)
);

BUFx6f_ASAP7_75t_SL g677 ( 
.A(n_570),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_503),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_SL g679 ( 
.A(n_603),
.B(n_214),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_L g680 ( 
.A(n_634),
.B(n_436),
.Y(n_680)
);

INVx2_ASAP7_75t_L g681 ( 
.A(n_508),
.Y(n_681)
);

NOR2xp33_ASAP7_75t_L g682 ( 
.A(n_505),
.B(n_412),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_SL g683 ( 
.A(n_603),
.B(n_214),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_SL g684 ( 
.A(n_528),
.B(n_214),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_SL g685 ( 
.A(n_528),
.B(n_512),
.Y(n_685)
);

BUFx3_ASAP7_75t_L g686 ( 
.A(n_510),
.Y(n_686)
);

NOR2xp33_ASAP7_75t_L g687 ( 
.A(n_513),
.B(n_358),
.Y(n_687)
);

NOR2xp33_ASAP7_75t_L g688 ( 
.A(n_523),
.B(n_181),
.Y(n_688)
);

AOI22xp5_ASAP7_75t_L g689 ( 
.A1(n_535),
.A2(n_495),
.B1(n_200),
.B2(n_186),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_L g690 ( 
.A(n_568),
.B(n_436),
.Y(n_690)
);

OAI21xp5_ASAP7_75t_L g691 ( 
.A1(n_625),
.A2(n_432),
.B(n_460),
.Y(n_691)
);

INVx2_ASAP7_75t_L g692 ( 
.A(n_508),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_L g693 ( 
.A(n_591),
.B(n_460),
.Y(n_693)
);

NOR2xp33_ASAP7_75t_L g694 ( 
.A(n_567),
.B(n_181),
.Y(n_694)
);

CKINVDCx14_ASAP7_75t_R g695 ( 
.A(n_564),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_L g696 ( 
.A(n_591),
.B(n_495),
.Y(n_696)
);

INVx2_ASAP7_75t_L g697 ( 
.A(n_517),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_L g698 ( 
.A(n_628),
.B(n_479),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_L g699 ( 
.A(n_628),
.B(n_479),
.Y(n_699)
);

A2O1A1Ixp33_ASAP7_75t_L g700 ( 
.A1(n_571),
.A2(n_314),
.B(n_288),
.C(n_299),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_517),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_L g702 ( 
.A(n_628),
.B(n_479),
.Y(n_702)
);

BUFx6f_ASAP7_75t_L g703 ( 
.A(n_510),
.Y(n_703)
);

INVx3_ASAP7_75t_L g704 ( 
.A(n_628),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_L g705 ( 
.A(n_638),
.B(n_479),
.Y(n_705)
);

AOI22xp33_ASAP7_75t_L g706 ( 
.A1(n_571),
.A2(n_285),
.B1(n_493),
.B2(n_214),
.Y(n_706)
);

BUFx6f_ASAP7_75t_L g707 ( 
.A(n_510),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_525),
.Y(n_708)
);

BUFx3_ASAP7_75t_L g709 ( 
.A(n_514),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_L g710 ( 
.A(n_638),
.B(n_479),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_SL g711 ( 
.A(n_540),
.B(n_183),
.Y(n_711)
);

O2A1O1Ixp33_ASAP7_75t_L g712 ( 
.A1(n_635),
.A2(n_476),
.B(n_487),
.C(n_493),
.Y(n_712)
);

INVx2_ASAP7_75t_L g713 ( 
.A(n_525),
.Y(n_713)
);

NOR2xp33_ASAP7_75t_L g714 ( 
.A(n_623),
.B(n_183),
.Y(n_714)
);

NAND3xp33_ASAP7_75t_L g715 ( 
.A(n_579),
.B(n_261),
.C(n_247),
.Y(n_715)
);

INVx2_ASAP7_75t_SL g716 ( 
.A(n_583),
.Y(n_716)
);

INVx2_ASAP7_75t_L g717 ( 
.A(n_527),
.Y(n_717)
);

INVx2_ASAP7_75t_L g718 ( 
.A(n_527),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_L g719 ( 
.A(n_638),
.B(n_479),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_SL g720 ( 
.A(n_528),
.B(n_256),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_SL g721 ( 
.A(n_528),
.B(n_256),
.Y(n_721)
);

INVx3_ASAP7_75t_L g722 ( 
.A(n_638),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_L g723 ( 
.A(n_534),
.B(n_424),
.Y(n_723)
);

INVx2_ASAP7_75t_L g724 ( 
.A(n_534),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_L g725 ( 
.A(n_544),
.B(n_424),
.Y(n_725)
);

INVx2_ASAP7_75t_SL g726 ( 
.A(n_543),
.Y(n_726)
);

INVx2_ASAP7_75t_L g727 ( 
.A(n_544),
.Y(n_727)
);

INVx2_ASAP7_75t_L g728 ( 
.A(n_552),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_552),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_L g730 ( 
.A(n_551),
.B(n_557),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_551),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_557),
.Y(n_732)
);

INVx2_ASAP7_75t_SL g733 ( 
.A(n_543),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_L g734 ( 
.A(n_640),
.B(n_438),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_L g735 ( 
.A(n_547),
.B(n_438),
.Y(n_735)
);

INVx2_ASAP7_75t_L g736 ( 
.A(n_643),
.Y(n_736)
);

OAI22xp5_ASAP7_75t_L g737 ( 
.A1(n_512),
.A2(n_282),
.B1(n_293),
.B2(n_185),
.Y(n_737)
);

INVx2_ASAP7_75t_L g738 ( 
.A(n_643),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_L g739 ( 
.A(n_514),
.B(n_522),
.Y(n_739)
);

INVx2_ASAP7_75t_SL g740 ( 
.A(n_532),
.Y(n_740)
);

BUFx2_ASAP7_75t_L g741 ( 
.A(n_532),
.Y(n_741)
);

NOR2xp33_ASAP7_75t_L g742 ( 
.A(n_580),
.B(n_185),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_553),
.Y(n_743)
);

NOR2xp33_ASAP7_75t_L g744 ( 
.A(n_572),
.B(n_186),
.Y(n_744)
);

OAI22xp5_ASAP7_75t_L g745 ( 
.A1(n_512),
.A2(n_324),
.B1(n_194),
.B2(n_199),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_SL g746 ( 
.A(n_565),
.B(n_190),
.Y(n_746)
);

AOI22xp5_ASAP7_75t_L g747 ( 
.A1(n_501),
.A2(n_194),
.B1(n_328),
.B2(n_190),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_SL g748 ( 
.A(n_506),
.B(n_199),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_L g749 ( 
.A(n_514),
.B(n_438),
.Y(n_749)
);

INVx4_ASAP7_75t_L g750 ( 
.A(n_522),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_L g751 ( 
.A(n_522),
.B(n_440),
.Y(n_751)
);

OAI22xp5_ASAP7_75t_L g752 ( 
.A1(n_512),
.A2(n_325),
.B1(n_203),
.B2(n_206),
.Y(n_752)
);

AOI22xp5_ASAP7_75t_L g753 ( 
.A1(n_524),
.A2(n_200),
.B1(n_328),
.B2(n_203),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_SL g754 ( 
.A(n_520),
.B(n_206),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_553),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_554),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_SL g757 ( 
.A(n_536),
.B(n_207),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_L g758 ( 
.A(n_554),
.B(n_440),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_L g759 ( 
.A(n_555),
.B(n_440),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_L g760 ( 
.A(n_555),
.B(n_441),
.Y(n_760)
);

NAND3xp33_ASAP7_75t_L g761 ( 
.A(n_647),
.B(n_338),
.C(n_292),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_L g762 ( 
.A(n_558),
.B(n_441),
.Y(n_762)
);

INVx2_ASAP7_75t_SL g763 ( 
.A(n_577),
.Y(n_763)
);

INVx2_ASAP7_75t_L g764 ( 
.A(n_643),
.Y(n_764)
);

HB1xp67_ASAP7_75t_L g765 ( 
.A(n_578),
.Y(n_765)
);

O2A1O1Ixp33_ASAP7_75t_L g766 ( 
.A1(n_635),
.A2(n_476),
.B(n_487),
.C(n_493),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_L g767 ( 
.A(n_558),
.B(n_441),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_L g768 ( 
.A(n_560),
.B(n_443),
.Y(n_768)
);

NAND2xp33_ASAP7_75t_SL g769 ( 
.A(n_624),
.B(n_188),
.Y(n_769)
);

INVx2_ASAP7_75t_L g770 ( 
.A(n_645),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_L g771 ( 
.A(n_560),
.B(n_443),
.Y(n_771)
);

A2O1A1Ixp33_ASAP7_75t_L g772 ( 
.A1(n_571),
.A2(n_476),
.B(n_487),
.C(n_494),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_561),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_L g774 ( 
.A(n_561),
.B(n_443),
.Y(n_774)
);

OAI22xp5_ASAP7_75t_L g775 ( 
.A1(n_524),
.A2(n_207),
.B1(n_209),
.B2(n_300),
.Y(n_775)
);

NAND2xp33_ASAP7_75t_L g776 ( 
.A(n_500),
.B(n_256),
.Y(n_776)
);

OAI22xp5_ASAP7_75t_L g777 ( 
.A1(n_524),
.A2(n_321),
.B1(n_300),
.B2(n_309),
.Y(n_777)
);

NOR2xp33_ASAP7_75t_L g778 ( 
.A(n_590),
.B(n_598),
.Y(n_778)
);

NOR2xp33_ASAP7_75t_L g779 ( 
.A(n_584),
.B(n_209),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_L g780 ( 
.A(n_581),
.B(n_451),
.Y(n_780)
);

INVx2_ASAP7_75t_L g781 ( 
.A(n_645),
.Y(n_781)
);

INVx1_ASAP7_75t_L g782 ( 
.A(n_581),
.Y(n_782)
);

INVx2_ASAP7_75t_L g783 ( 
.A(n_645),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_L g784 ( 
.A(n_593),
.B(n_451),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_L g785 ( 
.A(n_593),
.B(n_451),
.Y(n_785)
);

NAND2xp33_ASAP7_75t_L g786 ( 
.A(n_500),
.B(n_636),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_L g787 ( 
.A(n_595),
.B(n_453),
.Y(n_787)
);

NAND2xp33_ASAP7_75t_L g788 ( 
.A(n_500),
.B(n_256),
.Y(n_788)
);

OAI22xp5_ASAP7_75t_L g789 ( 
.A1(n_524),
.A2(n_324),
.B1(n_321),
.B2(n_309),
.Y(n_789)
);

INVx1_ASAP7_75t_SL g790 ( 
.A(n_545),
.Y(n_790)
);

NOR2xp33_ASAP7_75t_L g791 ( 
.A(n_586),
.B(n_325),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_L g792 ( 
.A(n_595),
.B(n_453),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_L g793 ( 
.A(n_602),
.B(n_453),
.Y(n_793)
);

NAND2xp33_ASAP7_75t_L g794 ( 
.A(n_500),
.B(n_256),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_L g795 ( 
.A(n_602),
.B(n_570),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_L g796 ( 
.A(n_570),
.B(n_457),
.Y(n_796)
);

NOR2xp33_ASAP7_75t_L g797 ( 
.A(n_631),
.B(n_327),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_L g798 ( 
.A(n_570),
.B(n_646),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_620),
.Y(n_799)
);

AND2x2_ASAP7_75t_L g800 ( 
.A(n_559),
.B(n_385),
.Y(n_800)
);

BUFx6f_ASAP7_75t_L g801 ( 
.A(n_542),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_L g802 ( 
.A(n_516),
.B(n_457),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_L g803 ( 
.A(n_516),
.B(n_457),
.Y(n_803)
);

OR2x2_ASAP7_75t_L g804 ( 
.A(n_648),
.B(n_415),
.Y(n_804)
);

NAND2x1p5_ASAP7_75t_L g805 ( 
.A(n_549),
.B(n_494),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_604),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_604),
.Y(n_807)
);

AND2x2_ASAP7_75t_L g808 ( 
.A(n_633),
.B(n_385),
.Y(n_808)
);

AND2x2_ASAP7_75t_L g809 ( 
.A(n_648),
.B(n_398),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_605),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_L g811 ( 
.A(n_516),
.B(n_459),
.Y(n_811)
);

NAND3xp33_ASAP7_75t_L g812 ( 
.A(n_630),
.B(n_266),
.C(n_275),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_605),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_L g814 ( 
.A(n_516),
.B(n_459),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_SL g815 ( 
.A(n_528),
.B(n_256),
.Y(n_815)
);

BUFx12f_ASAP7_75t_L g816 ( 
.A(n_500),
.Y(n_816)
);

OAI22xp5_ASAP7_75t_L g817 ( 
.A1(n_655),
.A2(n_549),
.B1(n_615),
.B2(n_607),
.Y(n_817)
);

AOI21xp5_ASAP7_75t_L g818 ( 
.A1(n_680),
.A2(n_549),
.B(n_614),
.Y(n_818)
);

HB1xp67_ASAP7_75t_L g819 ( 
.A(n_726),
.Y(n_819)
);

O2A1O1Ixp5_ASAP7_75t_L g820 ( 
.A1(n_679),
.A2(n_608),
.B(n_616),
.C(n_619),
.Y(n_820)
);

A2O1A1Ixp33_ASAP7_75t_L g821 ( 
.A1(n_778),
.A2(n_641),
.B(n_613),
.C(n_618),
.Y(n_821)
);

HB1xp67_ASAP7_75t_L g822 ( 
.A(n_733),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_L g823 ( 
.A(n_778),
.B(n_500),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_L g824 ( 
.A(n_763),
.B(n_500),
.Y(n_824)
);

NOR3xp33_ASAP7_75t_L g825 ( 
.A(n_659),
.B(n_398),
.C(n_327),
.Y(n_825)
);

AOI21xp5_ASAP7_75t_L g826 ( 
.A1(n_690),
.A2(n_614),
.B(n_542),
.Y(n_826)
);

NOR2xp33_ASAP7_75t_L g827 ( 
.A(n_659),
.B(n_609),
.Y(n_827)
);

BUFx6f_ASAP7_75t_L g828 ( 
.A(n_801),
.Y(n_828)
);

INVx1_ASAP7_75t_SL g829 ( 
.A(n_790),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_SL g830 ( 
.A(n_693),
.B(n_542),
.Y(n_830)
);

OAI22xp5_ASAP7_75t_L g831 ( 
.A1(n_706),
.A2(n_612),
.B1(n_609),
.B2(n_610),
.Y(n_831)
);

NOR2xp33_ASAP7_75t_L g832 ( 
.A(n_744),
.B(n_610),
.Y(n_832)
);

AND2x2_ASAP7_75t_L g833 ( 
.A(n_674),
.B(n_415),
.Y(n_833)
);

AOI21xp5_ASAP7_75t_L g834 ( 
.A1(n_691),
.A2(n_542),
.B(n_546),
.Y(n_834)
);

OAI21xp33_ASAP7_75t_L g835 ( 
.A1(n_714),
.A2(n_191),
.B(n_188),
.Y(n_835)
);

A2O1A1Ixp33_ASAP7_75t_L g836 ( 
.A1(n_744),
.A2(n_622),
.B(n_617),
.C(n_612),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_L g837 ( 
.A(n_687),
.B(n_613),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_L g838 ( 
.A(n_687),
.B(n_617),
.Y(n_838)
);

HB1xp67_ASAP7_75t_SL g839 ( 
.A(n_671),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_L g840 ( 
.A(n_765),
.B(n_618),
.Y(n_840)
);

AOI21xp5_ASAP7_75t_L g841 ( 
.A1(n_786),
.A2(n_597),
.B(n_546),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_SL g842 ( 
.A(n_730),
.B(n_541),
.Y(n_842)
);

OAI21xp5_ASAP7_75t_L g843 ( 
.A1(n_772),
.A2(n_683),
.B(n_679),
.Y(n_843)
);

AOI21xp5_ASAP7_75t_L g844 ( 
.A1(n_798),
.A2(n_597),
.B(n_546),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_L g845 ( 
.A(n_714),
.B(n_622),
.Y(n_845)
);

A2O1A1Ixp33_ASAP7_75t_L g846 ( 
.A1(n_675),
.A2(n_629),
.B(n_616),
.C(n_608),
.Y(n_846)
);

INVx2_ASAP7_75t_L g847 ( 
.A(n_654),
.Y(n_847)
);

AND2x2_ASAP7_75t_L g848 ( 
.A(n_716),
.B(n_419),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_L g849 ( 
.A(n_694),
.B(n_629),
.Y(n_849)
);

AND2x2_ASAP7_75t_L g850 ( 
.A(n_809),
.B(n_419),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_L g851 ( 
.A(n_694),
.B(n_541),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_L g852 ( 
.A(n_779),
.B(n_541),
.Y(n_852)
);

NOR2xp33_ASAP7_75t_L g853 ( 
.A(n_652),
.B(n_621),
.Y(n_853)
);

OAI22xp5_ASAP7_75t_L g854 ( 
.A1(n_706),
.A2(n_642),
.B1(n_585),
.B2(n_632),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_657),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_L g856 ( 
.A(n_779),
.B(n_541),
.Y(n_856)
);

OAI21xp5_ASAP7_75t_L g857 ( 
.A1(n_683),
.A2(n_621),
.B(n_637),
.Y(n_857)
);

AOI21xp5_ASAP7_75t_L g858 ( 
.A1(n_739),
.A2(n_597),
.B(n_546),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_657),
.Y(n_859)
);

A2O1A1Ixp33_ASAP7_75t_L g860 ( 
.A1(n_675),
.A2(n_621),
.B(n_637),
.C(n_627),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_SL g861 ( 
.A(n_799),
.B(n_576),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_L g862 ( 
.A(n_791),
.B(n_576),
.Y(n_862)
);

A2O1A1Ixp33_ASAP7_75t_L g863 ( 
.A1(n_682),
.A2(n_627),
.B(n_637),
.C(n_632),
.Y(n_863)
);

NOR2xp33_ASAP7_75t_L g864 ( 
.A(n_656),
.B(n_627),
.Y(n_864)
);

O2A1O1Ixp33_ASAP7_75t_L g865 ( 
.A1(n_668),
.A2(n_562),
.B(n_548),
.C(n_556),
.Y(n_865)
);

BUFx12f_ASAP7_75t_L g866 ( 
.A(n_740),
.Y(n_866)
);

AOI21xp5_ASAP7_75t_L g867 ( 
.A1(n_650),
.A2(n_597),
.B(n_546),
.Y(n_867)
);

OR2x2_ASAP7_75t_L g868 ( 
.A(n_804),
.B(n_589),
.Y(n_868)
);

O2A1O1Ixp33_ASAP7_75t_L g869 ( 
.A1(n_731),
.A2(n_562),
.B(n_548),
.C(n_556),
.Y(n_869)
);

AOI21xp5_ASAP7_75t_L g870 ( 
.A1(n_649),
.A2(n_597),
.B(n_546),
.Y(n_870)
);

OAI21xp5_ASAP7_75t_L g871 ( 
.A1(n_712),
.A2(n_521),
.B(n_509),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_L g872 ( 
.A(n_791),
.B(n_642),
.Y(n_872)
);

BUFx3_ASAP7_75t_L g873 ( 
.A(n_741),
.Y(n_873)
);

AOI22xp5_ASAP7_75t_L g874 ( 
.A1(n_682),
.A2(n_589),
.B1(n_632),
.B2(n_576),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_L g875 ( 
.A(n_696),
.B(n_642),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_L g876 ( 
.A(n_688),
.B(n_642),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_L g877 ( 
.A(n_688),
.B(n_576),
.Y(n_877)
);

INVx2_ASAP7_75t_L g878 ( 
.A(n_663),
.Y(n_878)
);

BUFx6f_ASAP7_75t_L g879 ( 
.A(n_801),
.Y(n_879)
);

AND2x2_ASAP7_75t_L g880 ( 
.A(n_800),
.B(n_589),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_L g881 ( 
.A(n_735),
.B(n_585),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_L g882 ( 
.A(n_732),
.B(n_585),
.Y(n_882)
);

A2O1A1Ixp33_ASAP7_75t_L g883 ( 
.A1(n_742),
.A2(n_632),
.B(n_611),
.C(n_606),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_L g884 ( 
.A(n_664),
.B(n_672),
.Y(n_884)
);

AND2x4_ASAP7_75t_L g885 ( 
.A(n_686),
.B(n_472),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_SL g886 ( 
.A(n_658),
.B(n_312),
.Y(n_886)
);

NOR2xp33_ASAP7_75t_L g887 ( 
.A(n_666),
.B(n_742),
.Y(n_887)
);

AND2x4_ASAP7_75t_L g888 ( 
.A(n_686),
.B(n_709),
.Y(n_888)
);

NOR2xp67_ASAP7_75t_L g889 ( 
.A(n_715),
.B(n_472),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_SL g890 ( 
.A(n_670),
.B(n_585),
.Y(n_890)
);

BUFx6f_ASAP7_75t_L g891 ( 
.A(n_801),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_L g892 ( 
.A(n_678),
.B(n_587),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_SL g893 ( 
.A(n_704),
.B(n_587),
.Y(n_893)
);

AOI21xp5_ASAP7_75t_L g894 ( 
.A1(n_649),
.A2(n_597),
.B(n_611),
.Y(n_894)
);

INVx2_ASAP7_75t_L g895 ( 
.A(n_681),
.Y(n_895)
);

NAND2x1p5_ASAP7_75t_L g896 ( 
.A(n_685),
.B(n_587),
.Y(n_896)
);

INVx2_ASAP7_75t_L g897 ( 
.A(n_681),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_L g898 ( 
.A(n_701),
.B(n_587),
.Y(n_898)
);

O2A1O1Ixp33_ASAP7_75t_L g899 ( 
.A1(n_711),
.A2(n_662),
.B(n_737),
.C(n_766),
.Y(n_899)
);

INVx1_ASAP7_75t_L g900 ( 
.A(n_692),
.Y(n_900)
);

AOI21xp5_ASAP7_75t_L g901 ( 
.A1(n_665),
.A2(n_599),
.B(n_611),
.Y(n_901)
);

OR2x2_ASAP7_75t_L g902 ( 
.A(n_661),
.B(n_191),
.Y(n_902)
);

INVx1_ASAP7_75t_L g903 ( 
.A(n_692),
.Y(n_903)
);

INVx2_ASAP7_75t_L g904 ( 
.A(n_697),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_L g905 ( 
.A(n_708),
.B(n_729),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_697),
.Y(n_906)
);

BUFx4f_ASAP7_75t_L g907 ( 
.A(n_808),
.Y(n_907)
);

INVx3_ASAP7_75t_L g908 ( 
.A(n_703),
.Y(n_908)
);

AOI222xp33_ASAP7_75t_L g909 ( 
.A1(n_669),
.A2(n_335),
.B1(n_197),
.B2(n_201),
.C1(n_202),
.C2(n_204),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_L g910 ( 
.A(n_734),
.B(n_599),
.Y(n_910)
);

INVx4_ASAP7_75t_L g911 ( 
.A(n_703),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_L g912 ( 
.A(n_713),
.B(n_599),
.Y(n_912)
);

OAI22xp5_ASAP7_75t_L g913 ( 
.A1(n_685),
.A2(n_599),
.B1(n_611),
.B2(n_606),
.Y(n_913)
);

AOI21xp5_ASAP7_75t_L g914 ( 
.A1(n_665),
.A2(n_606),
.B(n_509),
.Y(n_914)
);

NOR2xp33_ASAP7_75t_L g915 ( 
.A(n_746),
.B(n_797),
.Y(n_915)
);

OAI21x1_ASAP7_75t_L g916 ( 
.A1(n_698),
.A2(n_606),
.B(n_548),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_L g917 ( 
.A(n_713),
.B(n_511),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_SL g918 ( 
.A(n_704),
.B(n_626),
.Y(n_918)
);

AOI21xp5_ASAP7_75t_L g919 ( 
.A1(n_667),
.A2(n_529),
.B(n_601),
.Y(n_919)
);

AOI21xp5_ASAP7_75t_L g920 ( 
.A1(n_667),
.A2(n_673),
.B(n_699),
.Y(n_920)
);

INVx1_ASAP7_75t_SL g921 ( 
.A(n_769),
.Y(n_921)
);

AND2x2_ASAP7_75t_L g922 ( 
.A(n_797),
.B(n_494),
.Y(n_922)
);

AOI21x1_ASAP7_75t_L g923 ( 
.A1(n_720),
.A2(n_515),
.B(n_601),
.Y(n_923)
);

BUFx12f_ASAP7_75t_L g924 ( 
.A(n_703),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_L g925 ( 
.A(n_717),
.B(n_511),
.Y(n_925)
);

HB1xp67_ASAP7_75t_L g926 ( 
.A(n_709),
.Y(n_926)
);

A2O1A1Ixp33_ASAP7_75t_L g927 ( 
.A1(n_795),
.A2(n_519),
.B(n_596),
.C(n_575),
.Y(n_927)
);

A2O1A1Ixp33_ASAP7_75t_L g928 ( 
.A1(n_689),
.A2(n_519),
.B(n_596),
.C(n_575),
.Y(n_928)
);

BUFx6f_ASAP7_75t_L g929 ( 
.A(n_801),
.Y(n_929)
);

NOR2xp33_ASAP7_75t_L g930 ( 
.A(n_748),
.B(n_277),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_717),
.Y(n_931)
);

INVx5_ASAP7_75t_L g932 ( 
.A(n_816),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_L g933 ( 
.A(n_718),
.B(n_518),
.Y(n_933)
);

AOI21xp5_ASAP7_75t_L g934 ( 
.A1(n_673),
.A2(n_521),
.B(n_529),
.Y(n_934)
);

OAI21xp33_ASAP7_75t_L g935 ( 
.A1(n_669),
.A2(n_197),
.B(n_201),
.Y(n_935)
);

AND2x2_ASAP7_75t_L g936 ( 
.A(n_669),
.B(n_494),
.Y(n_936)
);

NAND2xp5_ASAP7_75t_SL g937 ( 
.A(n_703),
.B(n_626),
.Y(n_937)
);

NAND2xp5_ASAP7_75t_L g938 ( 
.A(n_718),
.B(n_530),
.Y(n_938)
);

NOR2xp33_ASAP7_75t_R g939 ( 
.A(n_695),
.B(n_195),
.Y(n_939)
);

INVx1_ASAP7_75t_L g940 ( 
.A(n_724),
.Y(n_940)
);

INVx2_ASAP7_75t_L g941 ( 
.A(n_724),
.Y(n_941)
);

AOI21xp5_ASAP7_75t_L g942 ( 
.A1(n_702),
.A2(n_537),
.B(n_530),
.Y(n_942)
);

AOI21xp5_ASAP7_75t_L g943 ( 
.A1(n_705),
.A2(n_539),
.B(n_537),
.Y(n_943)
);

NOR2xp33_ASAP7_75t_L g944 ( 
.A(n_754),
.B(n_279),
.Y(n_944)
);

NOR2xp33_ASAP7_75t_SL g945 ( 
.A(n_677),
.B(n_195),
.Y(n_945)
);

OAI21xp5_ASAP7_75t_L g946 ( 
.A1(n_651),
.A2(n_538),
.B(n_539),
.Y(n_946)
);

O2A1O1Ixp33_ASAP7_75t_L g947 ( 
.A1(n_700),
.A2(n_573),
.B(n_566),
.C(n_563),
.Y(n_947)
);

INVx2_ASAP7_75t_L g948 ( 
.A(n_727),
.Y(n_948)
);

INVx2_ASAP7_75t_L g949 ( 
.A(n_727),
.Y(n_949)
);

OAI21xp5_ASAP7_75t_L g950 ( 
.A1(n_653),
.A2(n_538),
.B(n_573),
.Y(n_950)
);

INVx2_ASAP7_75t_L g951 ( 
.A(n_728),
.Y(n_951)
);

OR2x2_ASAP7_75t_L g952 ( 
.A(n_757),
.B(n_202),
.Y(n_952)
);

AOI22xp33_ASAP7_75t_L g953 ( 
.A1(n_676),
.A2(n_728),
.B1(n_783),
.B2(n_736),
.Y(n_953)
);

CKINVDCx5p33_ASAP7_75t_R g954 ( 
.A(n_747),
.Y(n_954)
);

AND2x2_ASAP7_75t_L g955 ( 
.A(n_812),
.B(n_204),
.Y(n_955)
);

AOI22xp5_ASAP7_75t_L g956 ( 
.A1(n_722),
.A2(n_573),
.B1(n_566),
.B2(n_563),
.Y(n_956)
);

AOI21x1_ASAP7_75t_L g957 ( 
.A1(n_720),
.A2(n_556),
.B(n_566),
.Y(n_957)
);

INVx1_ASAP7_75t_L g958 ( 
.A(n_743),
.Y(n_958)
);

A2O1A1Ixp33_ASAP7_75t_L g959 ( 
.A1(n_755),
.A2(n_562),
.B(n_563),
.C(n_486),
.Y(n_959)
);

AOI21xp33_ASAP7_75t_L g960 ( 
.A1(n_753),
.A2(n_211),
.B(n_212),
.Y(n_960)
);

INVxp33_ASAP7_75t_L g961 ( 
.A(n_761),
.Y(n_961)
);

O2A1O1Ixp5_ASAP7_75t_L g962 ( 
.A1(n_723),
.A2(n_459),
.B(n_492),
.C(n_471),
.Y(n_962)
);

NAND2xp5_ASAP7_75t_L g963 ( 
.A(n_736),
.B(n_626),
.Y(n_963)
);

NOR3xp33_ASAP7_75t_L g964 ( 
.A(n_745),
.B(n_330),
.C(n_212),
.Y(n_964)
);

BUFx6f_ASAP7_75t_L g965 ( 
.A(n_707),
.Y(n_965)
);

NAND2xp5_ASAP7_75t_L g966 ( 
.A(n_738),
.B(n_626),
.Y(n_966)
);

NAND2xp5_ASAP7_75t_SL g967 ( 
.A(n_722),
.B(n_626),
.Y(n_967)
);

AO21x1_ASAP7_75t_L g968 ( 
.A1(n_721),
.A2(n_478),
.B(n_490),
.Y(n_968)
);

CKINVDCx5p33_ASAP7_75t_R g969 ( 
.A(n_677),
.Y(n_969)
);

AO21x1_ASAP7_75t_L g970 ( 
.A1(n_721),
.A2(n_478),
.B(n_490),
.Y(n_970)
);

INVx3_ASAP7_75t_L g971 ( 
.A(n_707),
.Y(n_971)
);

O2A1O1Ixp33_ASAP7_75t_L g972 ( 
.A1(n_725),
.A2(n_485),
.B(n_490),
.C(n_489),
.Y(n_972)
);

AO21x1_ASAP7_75t_L g973 ( 
.A1(n_815),
.A2(n_478),
.B(n_489),
.Y(n_973)
);

AND2x2_ASAP7_75t_L g974 ( 
.A(n_752),
.B(n_211),
.Y(n_974)
);

NAND2xp5_ASAP7_75t_SL g975 ( 
.A(n_707),
.B(n_472),
.Y(n_975)
);

NAND2xp5_ASAP7_75t_L g976 ( 
.A(n_738),
.B(n_471),
.Y(n_976)
);

CKINVDCx5p33_ASAP7_75t_R g977 ( 
.A(n_775),
.Y(n_977)
);

AOI21xp5_ASAP7_75t_L g978 ( 
.A1(n_710),
.A2(n_439),
.B(n_431),
.Y(n_978)
);

AND2x2_ASAP7_75t_L g979 ( 
.A(n_777),
.B(n_302),
.Y(n_979)
);

OAI21xp5_ASAP7_75t_L g980 ( 
.A1(n_660),
.A2(n_437),
.B(n_442),
.Y(n_980)
);

AOI21xp5_ASAP7_75t_L g981 ( 
.A1(n_719),
.A2(n_439),
.B(n_431),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_L g982 ( 
.A(n_764),
.B(n_471),
.Y(n_982)
);

AND2x4_ASAP7_75t_L g983 ( 
.A(n_750),
.B(n_485),
.Y(n_983)
);

AOI21xp5_ASAP7_75t_L g984 ( 
.A1(n_796),
.A2(n_439),
.B(n_431),
.Y(n_984)
);

AOI21xp5_ASAP7_75t_L g985 ( 
.A1(n_749),
.A2(n_751),
.B(n_805),
.Y(n_985)
);

AOI21xp5_ASAP7_75t_L g986 ( 
.A1(n_805),
.A2(n_431),
.B(n_437),
.Y(n_986)
);

NAND2xp5_ASAP7_75t_L g987 ( 
.A(n_764),
.B(n_492),
.Y(n_987)
);

AND2x4_ASAP7_75t_L g988 ( 
.A(n_750),
.B(n_707),
.Y(n_988)
);

NAND2xp5_ASAP7_75t_L g989 ( 
.A(n_770),
.B(n_492),
.Y(n_989)
);

AOI21xp5_ASAP7_75t_L g990 ( 
.A1(n_776),
.A2(n_431),
.B(n_437),
.Y(n_990)
);

INVx1_ASAP7_75t_L g991 ( 
.A(n_756),
.Y(n_991)
);

AND2x2_ASAP7_75t_SL g992 ( 
.A(n_788),
.B(n_485),
.Y(n_992)
);

NAND2xp5_ASAP7_75t_L g993 ( 
.A(n_770),
.B(n_471),
.Y(n_993)
);

NAND2xp5_ASAP7_75t_L g994 ( 
.A(n_781),
.B(n_492),
.Y(n_994)
);

BUFx6f_ASAP7_75t_L g995 ( 
.A(n_816),
.Y(n_995)
);

A2O1A1Ixp33_ASAP7_75t_L g996 ( 
.A1(n_773),
.A2(n_489),
.B(n_488),
.C(n_486),
.Y(n_996)
);

NOR2xp33_ASAP7_75t_L g997 ( 
.A(n_789),
.B(n_302),
.Y(n_997)
);

NOR2xp33_ASAP7_75t_SL g998 ( 
.A(n_782),
.B(n_304),
.Y(n_998)
);

INVx1_ASAP7_75t_L g999 ( 
.A(n_806),
.Y(n_999)
);

NOR2xp33_ASAP7_75t_R g1000 ( 
.A(n_794),
.B(n_304),
.Y(n_1000)
);

AOI21xp5_ASAP7_75t_L g1001 ( 
.A1(n_823),
.A2(n_781),
.B(n_783),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_L g1002 ( 
.A(n_827),
.B(n_807),
.Y(n_1002)
);

NAND2xp5_ASAP7_75t_SL g1003 ( 
.A(n_907),
.B(n_810),
.Y(n_1003)
);

OR2x2_ASAP7_75t_L g1004 ( 
.A(n_829),
.B(n_815),
.Y(n_1004)
);

BUFx6f_ASAP7_75t_L g1005 ( 
.A(n_924),
.Y(n_1005)
);

NAND2xp5_ASAP7_75t_SL g1006 ( 
.A(n_907),
.B(n_813),
.Y(n_1006)
);

AND2x2_ASAP7_75t_L g1007 ( 
.A(n_850),
.B(n_676),
.Y(n_1007)
);

AOI22xp33_ASAP7_75t_L g1008 ( 
.A1(n_887),
.A2(n_676),
.B1(n_684),
.B2(n_758),
.Y(n_1008)
);

NAND2xp5_ASAP7_75t_L g1009 ( 
.A(n_827),
.B(n_832),
.Y(n_1009)
);

OR2x2_ASAP7_75t_L g1010 ( 
.A(n_902),
.B(n_759),
.Y(n_1010)
);

NOR2xp33_ASAP7_75t_R g1011 ( 
.A(n_839),
.B(n_760),
.Y(n_1011)
);

INVx1_ASAP7_75t_SL g1012 ( 
.A(n_873),
.Y(n_1012)
);

INVx4_ASAP7_75t_L g1013 ( 
.A(n_965),
.Y(n_1013)
);

AOI21xp5_ASAP7_75t_L g1014 ( 
.A1(n_818),
.A2(n_684),
.B(n_811),
.Y(n_1014)
);

NAND2xp5_ASAP7_75t_L g1015 ( 
.A(n_832),
.B(n_762),
.Y(n_1015)
);

INVxp67_ASAP7_75t_L g1016 ( 
.A(n_819),
.Y(n_1016)
);

BUFx6f_ASAP7_75t_L g1017 ( 
.A(n_995),
.Y(n_1017)
);

O2A1O1Ixp33_ASAP7_75t_L g1018 ( 
.A1(n_887),
.A2(n_825),
.B(n_915),
.C(n_997),
.Y(n_1018)
);

BUFx6f_ASAP7_75t_L g1019 ( 
.A(n_995),
.Y(n_1019)
);

OAI21xp5_ASAP7_75t_L g1020 ( 
.A1(n_843),
.A2(n_814),
.B(n_803),
.Y(n_1020)
);

O2A1O1Ixp33_ASAP7_75t_SL g1021 ( 
.A1(n_883),
.A2(n_768),
.B(n_793),
.C(n_792),
.Y(n_1021)
);

INVx4_ASAP7_75t_L g1022 ( 
.A(n_965),
.Y(n_1022)
);

NOR2xp33_ASAP7_75t_L g1023 ( 
.A(n_915),
.B(n_767),
.Y(n_1023)
);

NOR2xp33_ASAP7_75t_L g1024 ( 
.A(n_954),
.B(n_771),
.Y(n_1024)
);

A2O1A1Ixp33_ASAP7_75t_L g1025 ( 
.A1(n_899),
.A2(n_780),
.B(n_787),
.C(n_785),
.Y(n_1025)
);

O2A1O1Ixp33_ASAP7_75t_L g1026 ( 
.A1(n_825),
.A2(n_784),
.B(n_774),
.C(n_802),
.Y(n_1026)
);

NOR2xp33_ASAP7_75t_L g1027 ( 
.A(n_819),
.B(n_822),
.Y(n_1027)
);

NAND2xp5_ASAP7_75t_L g1028 ( 
.A(n_837),
.B(n_486),
.Y(n_1028)
);

OR2x6_ASAP7_75t_L g1029 ( 
.A(n_866),
.B(n_995),
.Y(n_1029)
);

INVx1_ASAP7_75t_L g1030 ( 
.A(n_855),
.Y(n_1030)
);

AOI21xp5_ASAP7_75t_L g1031 ( 
.A1(n_985),
.A2(n_444),
.B(n_442),
.Y(n_1031)
);

NOR3xp33_ASAP7_75t_SL g1032 ( 
.A(n_977),
.B(n_326),
.C(n_336),
.Y(n_1032)
);

NOR2xp33_ASAP7_75t_L g1033 ( 
.A(n_822),
.B(n_305),
.Y(n_1033)
);

INVx8_ASAP7_75t_L g1034 ( 
.A(n_888),
.Y(n_1034)
);

NOR3xp33_ASAP7_75t_SL g1035 ( 
.A(n_935),
.B(n_326),
.C(n_336),
.Y(n_1035)
);

A2O1A1Ixp33_ASAP7_75t_L g1036 ( 
.A1(n_930),
.A2(n_488),
.B(n_335),
.C(n_332),
.Y(n_1036)
);

NOR2xp33_ASAP7_75t_L g1037 ( 
.A(n_961),
.B(n_305),
.Y(n_1037)
);

A2O1A1Ixp33_ASAP7_75t_SL g1038 ( 
.A1(n_930),
.A2(n_483),
.B(n_475),
.C(n_444),
.Y(n_1038)
);

INVx1_ASAP7_75t_L g1039 ( 
.A(n_859),
.Y(n_1039)
);

HB1xp67_ASAP7_75t_L g1040 ( 
.A(n_926),
.Y(n_1040)
);

NAND2xp5_ASAP7_75t_L g1041 ( 
.A(n_838),
.B(n_483),
.Y(n_1041)
);

BUFx2_ASAP7_75t_L g1042 ( 
.A(n_939),
.Y(n_1042)
);

AOI21xp5_ASAP7_75t_L g1043 ( 
.A1(n_826),
.A2(n_444),
.B(n_442),
.Y(n_1043)
);

OAI22xp5_ASAP7_75t_L g1044 ( 
.A1(n_953),
.A2(n_332),
.B1(n_319),
.B2(n_323),
.Y(n_1044)
);

NAND2xp5_ASAP7_75t_L g1045 ( 
.A(n_840),
.B(n_483),
.Y(n_1045)
);

OAI22x1_ASAP7_75t_L g1046 ( 
.A1(n_997),
.A2(n_317),
.B1(n_319),
.B2(n_323),
.Y(n_1046)
);

OAI22x1_ASAP7_75t_L g1047 ( 
.A1(n_921),
.A2(n_317),
.B1(n_330),
.B2(n_7),
.Y(n_1047)
);

AOI221xp5_ASAP7_75t_L g1048 ( 
.A1(n_960),
.A2(n_475),
.B1(n_477),
.B2(n_473),
.C(n_14),
.Y(n_1048)
);

INVx3_ASAP7_75t_L g1049 ( 
.A(n_965),
.Y(n_1049)
);

AOI22xp5_ASAP7_75t_L g1050 ( 
.A1(n_817),
.A2(n_256),
.B1(n_475),
.B2(n_473),
.Y(n_1050)
);

A2O1A1Ixp33_ASAP7_75t_SL g1051 ( 
.A1(n_944),
.A2(n_256),
.B(n_79),
.C(n_168),
.Y(n_1051)
);

AOI21x1_ASAP7_75t_L g1052 ( 
.A1(n_834),
.A2(n_477),
.B(n_473),
.Y(n_1052)
);

AND2x2_ASAP7_75t_SL g1053 ( 
.A(n_964),
.B(n_5),
.Y(n_1053)
);

NAND2xp5_ASAP7_75t_L g1054 ( 
.A(n_880),
.B(n_477),
.Y(n_1054)
);

INVx4_ASAP7_75t_SL g1055 ( 
.A(n_828),
.Y(n_1055)
);

AOI22xp5_ASAP7_75t_L g1056 ( 
.A1(n_944),
.A2(n_473),
.B1(n_477),
.B2(n_76),
.Y(n_1056)
);

AOI21xp5_ASAP7_75t_L g1057 ( 
.A1(n_876),
.A2(n_477),
.B(n_473),
.Y(n_1057)
);

NOR2xp33_ASAP7_75t_L g1058 ( 
.A(n_998),
.B(n_6),
.Y(n_1058)
);

AOI21xp5_ASAP7_75t_L g1059 ( 
.A1(n_877),
.A2(n_477),
.B(n_473),
.Y(n_1059)
);

OAI21x1_ASAP7_75t_L g1060 ( 
.A1(n_957),
.A2(n_84),
.B(n_167),
.Y(n_1060)
);

OR2x2_ASAP7_75t_L g1061 ( 
.A(n_833),
.B(n_477),
.Y(n_1061)
);

AND2x2_ASAP7_75t_L g1062 ( 
.A(n_848),
.B(n_477),
.Y(n_1062)
);

NOR2xp33_ASAP7_75t_L g1063 ( 
.A(n_835),
.B(n_955),
.Y(n_1063)
);

AOI21xp5_ASAP7_75t_L g1064 ( 
.A1(n_852),
.A2(n_473),
.B(n_71),
.Y(n_1064)
);

NAND2xp5_ASAP7_75t_L g1065 ( 
.A(n_922),
.B(n_473),
.Y(n_1065)
);

O2A1O1Ixp33_ASAP7_75t_L g1066 ( 
.A1(n_964),
.A2(n_11),
.B(n_14),
.C(n_15),
.Y(n_1066)
);

AND3x1_ASAP7_75t_SL g1067 ( 
.A(n_909),
.B(n_939),
.C(n_958),
.Y(n_1067)
);

AOI22xp33_ASAP7_75t_L g1068 ( 
.A1(n_868),
.A2(n_11),
.B1(n_20),
.B2(n_21),
.Y(n_1068)
);

NAND2xp5_ASAP7_75t_L g1069 ( 
.A(n_884),
.B(n_21),
.Y(n_1069)
);

OAI22xp5_ASAP7_75t_L g1070 ( 
.A1(n_953),
.A2(n_24),
.B1(n_27),
.B2(n_30),
.Y(n_1070)
);

BUFx3_ASAP7_75t_L g1071 ( 
.A(n_969),
.Y(n_1071)
);

NOR2xp33_ASAP7_75t_L g1072 ( 
.A(n_926),
.B(n_27),
.Y(n_1072)
);

AOI21xp5_ASAP7_75t_L g1073 ( 
.A1(n_856),
.A2(n_97),
.B(n_149),
.Y(n_1073)
);

NAND2xp5_ASAP7_75t_L g1074 ( 
.A(n_905),
.B(n_32),
.Y(n_1074)
);

INVx1_ASAP7_75t_L g1075 ( 
.A(n_900),
.Y(n_1075)
);

NAND2xp5_ASAP7_75t_L g1076 ( 
.A(n_845),
.B(n_32),
.Y(n_1076)
);

AOI22xp5_ASAP7_75t_L g1077 ( 
.A1(n_889),
.A2(n_96),
.B1(n_145),
.B2(n_144),
.Y(n_1077)
);

A2O1A1Ixp33_ASAP7_75t_L g1078 ( 
.A1(n_920),
.A2(n_36),
.B(n_42),
.C(n_43),
.Y(n_1078)
);

OAI21x1_ASAP7_75t_L g1079 ( 
.A1(n_923),
.A2(n_916),
.B(n_934),
.Y(n_1079)
);

NOR2xp33_ASAP7_75t_L g1080 ( 
.A(n_886),
.B(n_36),
.Y(n_1080)
);

BUFx3_ASAP7_75t_L g1081 ( 
.A(n_995),
.Y(n_1081)
);

BUFx8_ASAP7_75t_L g1082 ( 
.A(n_936),
.Y(n_1082)
);

NAND3xp33_ASAP7_75t_SL g1083 ( 
.A(n_945),
.B(n_46),
.C(n_47),
.Y(n_1083)
);

BUFx2_ASAP7_75t_L g1084 ( 
.A(n_1000),
.Y(n_1084)
);

INVx1_ASAP7_75t_L g1085 ( 
.A(n_903),
.Y(n_1085)
);

NOR2xp33_ASAP7_75t_L g1086 ( 
.A(n_974),
.B(n_47),
.Y(n_1086)
);

NAND2xp5_ASAP7_75t_L g1087 ( 
.A(n_849),
.B(n_52),
.Y(n_1087)
);

AOI22xp5_ASAP7_75t_L g1088 ( 
.A1(n_885),
.A2(n_106),
.B1(n_142),
.B2(n_138),
.Y(n_1088)
);

AOI21xp5_ASAP7_75t_L g1089 ( 
.A1(n_862),
.A2(n_93),
.B(n_132),
.Y(n_1089)
);

AOI21xp5_ASAP7_75t_L g1090 ( 
.A1(n_872),
.A2(n_91),
.B(n_121),
.Y(n_1090)
);

OAI22xp5_ASAP7_75t_L g1091 ( 
.A1(n_992),
.A2(n_821),
.B1(n_999),
.B2(n_991),
.Y(n_1091)
);

INVx2_ASAP7_75t_L g1092 ( 
.A(n_847),
.Y(n_1092)
);

OAI22xp5_ASAP7_75t_L g1093 ( 
.A1(n_992),
.A2(n_55),
.B1(n_56),
.B2(n_58),
.Y(n_1093)
);

OAI22xp5_ASAP7_75t_L g1094 ( 
.A1(n_874),
.A2(n_55),
.B1(n_62),
.B2(n_66),
.Y(n_1094)
);

NOR2xp33_ASAP7_75t_L g1095 ( 
.A(n_979),
.B(n_952),
.Y(n_1095)
);

NAND2xp5_ASAP7_75t_L g1096 ( 
.A(n_885),
.B(n_853),
.Y(n_1096)
);

NAND2xp5_ASAP7_75t_L g1097 ( 
.A(n_906),
.B(n_105),
.Y(n_1097)
);

NAND2xp5_ASAP7_75t_L g1098 ( 
.A(n_853),
.B(n_110),
.Y(n_1098)
);

AOI21xp5_ASAP7_75t_L g1099 ( 
.A1(n_875),
.A2(n_113),
.B(n_165),
.Y(n_1099)
);

NAND2xp5_ASAP7_75t_L g1100 ( 
.A(n_864),
.B(n_931),
.Y(n_1100)
);

AND2x4_ASAP7_75t_L g1101 ( 
.A(n_988),
.B(n_932),
.Y(n_1101)
);

INVx8_ASAP7_75t_L g1102 ( 
.A(n_988),
.Y(n_1102)
);

AO32x2_ASAP7_75t_L g1103 ( 
.A1(n_831),
.A2(n_854),
.A3(n_913),
.B1(n_911),
.B2(n_962),
.Y(n_1103)
);

NAND3xp33_ASAP7_75t_SL g1104 ( 
.A(n_1000),
.B(n_824),
.C(n_851),
.Y(n_1104)
);

OAI321xp33_ASAP7_75t_L g1105 ( 
.A1(n_940),
.A2(n_864),
.A3(n_910),
.B1(n_881),
.B2(n_882),
.C(n_871),
.Y(n_1105)
);

INVx8_ASAP7_75t_L g1106 ( 
.A(n_932),
.Y(n_1106)
);

NOR2xp33_ASAP7_75t_L g1107 ( 
.A(n_839),
.B(n_878),
.Y(n_1107)
);

INVx2_ASAP7_75t_L g1108 ( 
.A(n_895),
.Y(n_1108)
);

INVx1_ASAP7_75t_L g1109 ( 
.A(n_897),
.Y(n_1109)
);

O2A1O1Ixp33_ASAP7_75t_L g1110 ( 
.A1(n_996),
.A2(n_863),
.B(n_836),
.C(n_846),
.Y(n_1110)
);

AOI221xp5_ASAP7_75t_L g1111 ( 
.A1(n_972),
.A2(n_842),
.B1(n_861),
.B2(n_904),
.C(n_948),
.Y(n_1111)
);

INVx3_ASAP7_75t_L g1112 ( 
.A(n_911),
.Y(n_1112)
);

OAI22xp5_ASAP7_75t_L g1113 ( 
.A1(n_896),
.A2(n_949),
.B1(n_951),
.B2(n_941),
.Y(n_1113)
);

AOI21xp5_ASAP7_75t_L g1114 ( 
.A1(n_890),
.A2(n_830),
.B(n_842),
.Y(n_1114)
);

AOI22xp5_ASAP7_75t_L g1115 ( 
.A1(n_983),
.A2(n_975),
.B1(n_861),
.B2(n_893),
.Y(n_1115)
);

BUFx2_ASAP7_75t_SL g1116 ( 
.A(n_828),
.Y(n_1116)
);

NAND2xp5_ASAP7_75t_L g1117 ( 
.A(n_983),
.B(n_908),
.Y(n_1117)
);

AOI21xp5_ASAP7_75t_L g1118 ( 
.A1(n_912),
.A2(n_841),
.B(n_963),
.Y(n_1118)
);

INVx2_ASAP7_75t_L g1119 ( 
.A(n_917),
.Y(n_1119)
);

NAND2xp5_ASAP7_75t_L g1120 ( 
.A(n_908),
.B(n_971),
.Y(n_1120)
);

INVx4_ASAP7_75t_L g1121 ( 
.A(n_828),
.Y(n_1121)
);

INVx3_ASAP7_75t_SL g1122 ( 
.A(n_828),
.Y(n_1122)
);

CKINVDCx5p33_ASAP7_75t_R g1123 ( 
.A(n_879),
.Y(n_1123)
);

OAI21xp33_ASAP7_75t_SL g1124 ( 
.A1(n_892),
.A2(n_898),
.B(n_857),
.Y(n_1124)
);

AOI21xp5_ASAP7_75t_L g1125 ( 
.A1(n_966),
.A2(n_844),
.B(n_858),
.Y(n_1125)
);

OAI22xp5_ASAP7_75t_L g1126 ( 
.A1(n_896),
.A2(n_860),
.B1(n_929),
.B2(n_891),
.Y(n_1126)
);

OAI21xp33_ASAP7_75t_L g1127 ( 
.A1(n_925),
.A2(n_938),
.B(n_933),
.Y(n_1127)
);

AOI21xp5_ASAP7_75t_L g1128 ( 
.A1(n_867),
.A2(n_980),
.B(n_950),
.Y(n_1128)
);

NOR2xp33_ASAP7_75t_L g1129 ( 
.A(n_918),
.B(n_967),
.Y(n_1129)
);

AOI221xp5_ASAP7_75t_L g1130 ( 
.A1(n_869),
.A2(n_962),
.B1(n_865),
.B2(n_928),
.C(n_968),
.Y(n_1130)
);

O2A1O1Ixp33_ASAP7_75t_SL g1131 ( 
.A1(n_918),
.A2(n_967),
.B(n_959),
.C(n_927),
.Y(n_1131)
);

NAND2xp5_ASAP7_75t_L g1132 ( 
.A(n_976),
.B(n_994),
.Y(n_1132)
);

HB1xp67_ASAP7_75t_L g1133 ( 
.A(n_879),
.Y(n_1133)
);

CKINVDCx5p33_ASAP7_75t_R g1134 ( 
.A(n_879),
.Y(n_1134)
);

NOR2xp33_ASAP7_75t_L g1135 ( 
.A(n_970),
.B(n_973),
.Y(n_1135)
);

BUFx12f_ASAP7_75t_L g1136 ( 
.A(n_879),
.Y(n_1136)
);

NAND2xp5_ASAP7_75t_SL g1137 ( 
.A(n_891),
.B(n_929),
.Y(n_1137)
);

INVx2_ASAP7_75t_L g1138 ( 
.A(n_982),
.Y(n_1138)
);

INVxp67_ASAP7_75t_L g1139 ( 
.A(n_891),
.Y(n_1139)
);

AOI21xp5_ASAP7_75t_L g1140 ( 
.A1(n_901),
.A2(n_946),
.B(n_894),
.Y(n_1140)
);

BUFx2_ASAP7_75t_L g1141 ( 
.A(n_891),
.Y(n_1141)
);

AOI21xp5_ASAP7_75t_L g1142 ( 
.A1(n_987),
.A2(n_993),
.B(n_989),
.Y(n_1142)
);

AOI21xp5_ASAP7_75t_L g1143 ( 
.A1(n_820),
.A2(n_914),
.B(n_937),
.Y(n_1143)
);

INVx2_ASAP7_75t_L g1144 ( 
.A(n_929),
.Y(n_1144)
);

AOI21xp5_ASAP7_75t_L g1145 ( 
.A1(n_820),
.A2(n_870),
.B(n_929),
.Y(n_1145)
);

OAI21x1_ASAP7_75t_L g1146 ( 
.A1(n_1079),
.A2(n_919),
.B(n_942),
.Y(n_1146)
);

AO22x2_ASAP7_75t_L g1147 ( 
.A1(n_1094),
.A2(n_943),
.B1(n_981),
.B2(n_978),
.Y(n_1147)
);

NAND2xp5_ASAP7_75t_L g1148 ( 
.A(n_1009),
.B(n_984),
.Y(n_1148)
);

NOR2xp33_ASAP7_75t_L g1149 ( 
.A(n_1024),
.B(n_956),
.Y(n_1149)
);

BUFx6f_ASAP7_75t_L g1150 ( 
.A(n_1017),
.Y(n_1150)
);

OAI22xp5_ASAP7_75t_L g1151 ( 
.A1(n_1002),
.A2(n_990),
.B1(n_986),
.B2(n_947),
.Y(n_1151)
);

OAI21x1_ASAP7_75t_L g1152 ( 
.A1(n_1118),
.A2(n_1001),
.B(n_1031),
.Y(n_1152)
);

HB1xp67_ASAP7_75t_L g1153 ( 
.A(n_1040),
.Y(n_1153)
);

AO22x2_ASAP7_75t_L g1154 ( 
.A1(n_1094),
.A2(n_1093),
.B1(n_1070),
.B2(n_1083),
.Y(n_1154)
);

BUFx3_ASAP7_75t_L g1155 ( 
.A(n_1005),
.Y(n_1155)
);

NAND2xp5_ASAP7_75t_L g1156 ( 
.A(n_1023),
.B(n_1015),
.Y(n_1156)
);

INVx1_ASAP7_75t_L g1157 ( 
.A(n_1030),
.Y(n_1157)
);

INVx1_ASAP7_75t_L g1158 ( 
.A(n_1039),
.Y(n_1158)
);

AOI21xp5_ASAP7_75t_L g1159 ( 
.A1(n_1128),
.A2(n_1140),
.B(n_1025),
.Y(n_1159)
);

AOI21xp5_ASAP7_75t_L g1160 ( 
.A1(n_1014),
.A2(n_1021),
.B(n_1065),
.Y(n_1160)
);

AOI21xp5_ASAP7_75t_L g1161 ( 
.A1(n_1020),
.A2(n_1098),
.B(n_1041),
.Y(n_1161)
);

INVx5_ASAP7_75t_L g1162 ( 
.A(n_1106),
.Y(n_1162)
);

OA22x2_ASAP7_75t_L g1163 ( 
.A1(n_1046),
.A2(n_1047),
.B1(n_1093),
.B2(n_1070),
.Y(n_1163)
);

INVx1_ASAP7_75t_L g1164 ( 
.A(n_1075),
.Y(n_1164)
);

INVx1_ASAP7_75t_L g1165 ( 
.A(n_1085),
.Y(n_1165)
);

AOI21x1_ASAP7_75t_L g1166 ( 
.A1(n_1114),
.A2(n_1143),
.B(n_1126),
.Y(n_1166)
);

O2A1O1Ixp33_ASAP7_75t_SL g1167 ( 
.A1(n_1018),
.A2(n_1078),
.B(n_1051),
.C(n_1097),
.Y(n_1167)
);

NAND2xp5_ASAP7_75t_L g1168 ( 
.A(n_1010),
.B(n_1095),
.Y(n_1168)
);

AOI21xp5_ASAP7_75t_L g1169 ( 
.A1(n_1020),
.A2(n_1105),
.B(n_1054),
.Y(n_1169)
);

AOI22xp5_ASAP7_75t_L g1170 ( 
.A1(n_1086),
.A2(n_1053),
.B1(n_1058),
.B2(n_1063),
.Y(n_1170)
);

O2A1O1Ixp33_ASAP7_75t_L g1171 ( 
.A1(n_1036),
.A2(n_1080),
.B(n_1066),
.C(n_1037),
.Y(n_1171)
);

INVx1_ASAP7_75t_L g1172 ( 
.A(n_1109),
.Y(n_1172)
);

OR2x2_ASAP7_75t_L g1173 ( 
.A(n_1012),
.B(n_1004),
.Y(n_1173)
);

OAI21xp5_ASAP7_75t_L g1174 ( 
.A1(n_1026),
.A2(n_1135),
.B(n_1008),
.Y(n_1174)
);

A2O1A1Ixp33_ASAP7_75t_L g1175 ( 
.A1(n_1048),
.A2(n_1076),
.B(n_1087),
.C(n_1056),
.Y(n_1175)
);

OAI21xp5_ASAP7_75t_L g1176 ( 
.A1(n_1096),
.A2(n_1104),
.B(n_1091),
.Y(n_1176)
);

CKINVDCx20_ASAP7_75t_R g1177 ( 
.A(n_1071),
.Y(n_1177)
);

BUFx6f_ASAP7_75t_L g1178 ( 
.A(n_1017),
.Y(n_1178)
);

A2O1A1Ixp33_ASAP7_75t_L g1179 ( 
.A1(n_1069),
.A2(n_1074),
.B(n_1035),
.C(n_1091),
.Y(n_1179)
);

NOR2xp33_ASAP7_75t_SL g1180 ( 
.A(n_1106),
.B(n_1102),
.Y(n_1180)
);

OAI21xp5_ASAP7_75t_L g1181 ( 
.A1(n_1124),
.A2(n_1105),
.B(n_1115),
.Y(n_1181)
);

AOI21xp5_ASAP7_75t_L g1182 ( 
.A1(n_1100),
.A2(n_1132),
.B(n_1142),
.Y(n_1182)
);

AOI21xp5_ASAP7_75t_L g1183 ( 
.A1(n_1110),
.A2(n_1127),
.B(n_1028),
.Y(n_1183)
);

AO31x2_ASAP7_75t_L g1184 ( 
.A1(n_1126),
.A2(n_1113),
.A3(n_1064),
.B(n_1059),
.Y(n_1184)
);

AOI21xp5_ASAP7_75t_L g1185 ( 
.A1(n_1130),
.A2(n_1045),
.B(n_1131),
.Y(n_1185)
);

NAND3xp33_ASAP7_75t_L g1186 ( 
.A(n_1068),
.B(n_1033),
.C(n_1027),
.Y(n_1186)
);

A2O1A1Ixp33_ASAP7_75t_L g1187 ( 
.A1(n_1007),
.A2(n_1111),
.B(n_1073),
.C(n_1089),
.Y(n_1187)
);

AOI21xp5_ASAP7_75t_L g1188 ( 
.A1(n_1119),
.A2(n_1113),
.B(n_1138),
.Y(n_1188)
);

OAI21x1_ASAP7_75t_L g1189 ( 
.A1(n_1043),
.A2(n_1060),
.B(n_1057),
.Y(n_1189)
);

OR2x2_ASAP7_75t_L g1190 ( 
.A(n_1012),
.B(n_1016),
.Y(n_1190)
);

BUFx4_ASAP7_75t_SL g1191 ( 
.A(n_1029),
.Y(n_1191)
);

CKINVDCx5p33_ASAP7_75t_R g1192 ( 
.A(n_1042),
.Y(n_1192)
);

HB1xp67_ASAP7_75t_L g1193 ( 
.A(n_1123),
.Y(n_1193)
);

O2A1O1Ixp33_ASAP7_75t_SL g1194 ( 
.A1(n_1097),
.A2(n_1003),
.B(n_1006),
.C(n_1038),
.Y(n_1194)
);

NAND2xp5_ASAP7_75t_L g1195 ( 
.A(n_1107),
.B(n_1062),
.Y(n_1195)
);

OAI22xp5_ASAP7_75t_L g1196 ( 
.A1(n_1117),
.A2(n_1134),
.B1(n_1102),
.B2(n_1061),
.Y(n_1196)
);

AOI21xp5_ASAP7_75t_L g1197 ( 
.A1(n_1090),
.A2(n_1137),
.B(n_1102),
.Y(n_1197)
);

AO31x2_ASAP7_75t_L g1198 ( 
.A1(n_1129),
.A2(n_1099),
.A3(n_1120),
.B(n_1072),
.Y(n_1198)
);

AO31x2_ASAP7_75t_L g1199 ( 
.A1(n_1092),
.A2(n_1108),
.A3(n_1044),
.B(n_1103),
.Y(n_1199)
);

INVx1_ASAP7_75t_SL g1200 ( 
.A(n_1122),
.Y(n_1200)
);

NOR2xp33_ASAP7_75t_L g1201 ( 
.A(n_1084),
.B(n_1005),
.Y(n_1201)
);

OAI22x1_ASAP7_75t_L g1202 ( 
.A1(n_1067),
.A2(n_1088),
.B1(n_1050),
.B2(n_1077),
.Y(n_1202)
);

AO31x2_ASAP7_75t_L g1203 ( 
.A1(n_1044),
.A2(n_1103),
.A3(n_1144),
.B(n_1013),
.Y(n_1203)
);

INVx1_ASAP7_75t_L g1204 ( 
.A(n_1133),
.Y(n_1204)
);

INVx1_ASAP7_75t_L g1205 ( 
.A(n_1141),
.Y(n_1205)
);

NOR2xp33_ASAP7_75t_L g1206 ( 
.A(n_1005),
.B(n_1034),
.Y(n_1206)
);

NAND2xp5_ASAP7_75t_L g1207 ( 
.A(n_1034),
.B(n_1011),
.Y(n_1207)
);

INVx1_ASAP7_75t_L g1208 ( 
.A(n_1055),
.Y(n_1208)
);

INVx2_ASAP7_75t_L g1209 ( 
.A(n_1112),
.Y(n_1209)
);

OR2x6_ASAP7_75t_L g1210 ( 
.A(n_1106),
.B(n_1034),
.Y(n_1210)
);

INVx1_ASAP7_75t_L g1211 ( 
.A(n_1055),
.Y(n_1211)
);

OAI21x1_ASAP7_75t_L g1212 ( 
.A1(n_1049),
.A2(n_1103),
.B(n_1055),
.Y(n_1212)
);

OAI21xp5_ASAP7_75t_L g1213 ( 
.A1(n_1139),
.A2(n_1049),
.B(n_1032),
.Y(n_1213)
);

A2O1A1Ixp33_ASAP7_75t_L g1214 ( 
.A1(n_1101),
.A2(n_1081),
.B(n_1019),
.C(n_1017),
.Y(n_1214)
);

AOI221x1_ASAP7_75t_L g1215 ( 
.A1(n_1022),
.A2(n_1121),
.B1(n_1116),
.B2(n_1019),
.C(n_1082),
.Y(n_1215)
);

AO31x2_ASAP7_75t_L g1216 ( 
.A1(n_1121),
.A2(n_1082),
.A3(n_1136),
.B(n_1019),
.Y(n_1216)
);

AND2x4_ASAP7_75t_L g1217 ( 
.A(n_1029),
.B(n_1101),
.Y(n_1217)
);

AND2x4_ASAP7_75t_L g1218 ( 
.A(n_1029),
.B(n_1101),
.Y(n_1218)
);

AO31x2_ASAP7_75t_L g1219 ( 
.A1(n_1135),
.A2(n_1128),
.A3(n_1091),
.B(n_1126),
.Y(n_1219)
);

INVxp67_ASAP7_75t_L g1220 ( 
.A(n_1027),
.Y(n_1220)
);

AND2x4_ASAP7_75t_L g1221 ( 
.A(n_1101),
.B(n_1081),
.Y(n_1221)
);

NOR2x1_ASAP7_75t_L g1222 ( 
.A(n_1009),
.B(n_1002),
.Y(n_1222)
);

AOI21xp5_ASAP7_75t_L g1223 ( 
.A1(n_1128),
.A2(n_680),
.B(n_786),
.Y(n_1223)
);

A2O1A1Ixp33_ASAP7_75t_L g1224 ( 
.A1(n_1018),
.A2(n_887),
.B(n_915),
.C(n_1009),
.Y(n_1224)
);

AOI22xp33_ASAP7_75t_L g1225 ( 
.A1(n_1086),
.A2(n_887),
.B1(n_615),
.B2(n_744),
.Y(n_1225)
);

AO21x1_ASAP7_75t_L g1226 ( 
.A1(n_1009),
.A2(n_1018),
.B(n_1094),
.Y(n_1226)
);

INVx3_ASAP7_75t_L g1227 ( 
.A(n_1101),
.Y(n_1227)
);

NAND2xp5_ASAP7_75t_L g1228 ( 
.A(n_1009),
.B(n_1023),
.Y(n_1228)
);

A2O1A1Ixp33_ASAP7_75t_L g1229 ( 
.A1(n_1018),
.A2(n_887),
.B(n_915),
.C(n_1009),
.Y(n_1229)
);

NOR2xp33_ASAP7_75t_L g1230 ( 
.A(n_1024),
.B(n_659),
.Y(n_1230)
);

NAND2xp5_ASAP7_75t_L g1231 ( 
.A(n_1009),
.B(n_1023),
.Y(n_1231)
);

AO31x2_ASAP7_75t_L g1232 ( 
.A1(n_1135),
.A2(n_1128),
.A3(n_1091),
.B(n_1126),
.Y(n_1232)
);

OA21x2_ASAP7_75t_L g1233 ( 
.A1(n_1128),
.A2(n_1130),
.B(n_843),
.Y(n_1233)
);

INVx1_ASAP7_75t_L g1234 ( 
.A(n_1030),
.Y(n_1234)
);

OR2x2_ASAP7_75t_L g1235 ( 
.A(n_1010),
.B(n_507),
.Y(n_1235)
);

NOR2xp33_ASAP7_75t_L g1236 ( 
.A(n_1024),
.B(n_659),
.Y(n_1236)
);

NOR4xp25_ASAP7_75t_L g1237 ( 
.A(n_1018),
.B(n_1066),
.C(n_1093),
.D(n_1009),
.Y(n_1237)
);

A2O1A1Ixp33_ASAP7_75t_L g1238 ( 
.A1(n_1018),
.A2(n_887),
.B(n_915),
.C(n_1009),
.Y(n_1238)
);

INVx1_ASAP7_75t_SL g1239 ( 
.A(n_1012),
.Y(n_1239)
);

AOI21xp5_ASAP7_75t_L g1240 ( 
.A1(n_1128),
.A2(n_680),
.B(n_786),
.Y(n_1240)
);

NOR2xp33_ASAP7_75t_L g1241 ( 
.A(n_1024),
.B(n_659),
.Y(n_1241)
);

OAI21xp5_ASAP7_75t_L g1242 ( 
.A1(n_1009),
.A2(n_1018),
.B(n_887),
.Y(n_1242)
);

BUFx2_ASAP7_75t_L g1243 ( 
.A(n_1012),
.Y(n_1243)
);

OAI21xp5_ASAP7_75t_L g1244 ( 
.A1(n_1018),
.A2(n_843),
.B(n_1009),
.Y(n_1244)
);

NAND2xp5_ASAP7_75t_L g1245 ( 
.A(n_1009),
.B(n_1023),
.Y(n_1245)
);

AOI21x1_ASAP7_75t_L g1246 ( 
.A1(n_1052),
.A2(n_1145),
.B(n_1128),
.Y(n_1246)
);

OA21x2_ASAP7_75t_L g1247 ( 
.A1(n_1128),
.A2(n_1130),
.B(n_843),
.Y(n_1247)
);

AOI22xp5_ASAP7_75t_L g1248 ( 
.A1(n_1009),
.A2(n_887),
.B1(n_659),
.B2(n_1086),
.Y(n_1248)
);

NAND2xp5_ASAP7_75t_L g1249 ( 
.A(n_1009),
.B(n_1023),
.Y(n_1249)
);

AO31x2_ASAP7_75t_L g1250 ( 
.A1(n_1135),
.A2(n_1128),
.A3(n_1091),
.B(n_1126),
.Y(n_1250)
);

NAND2xp5_ASAP7_75t_L g1251 ( 
.A(n_1009),
.B(n_1023),
.Y(n_1251)
);

INVx1_ASAP7_75t_L g1252 ( 
.A(n_1030),
.Y(n_1252)
);

AOI21xp5_ASAP7_75t_L g1253 ( 
.A1(n_1128),
.A2(n_680),
.B(n_786),
.Y(n_1253)
);

AOI21xp5_ASAP7_75t_L g1254 ( 
.A1(n_1128),
.A2(n_680),
.B(n_786),
.Y(n_1254)
);

AOI21xp5_ASAP7_75t_L g1255 ( 
.A1(n_1128),
.A2(n_680),
.B(n_786),
.Y(n_1255)
);

OAI21x1_ASAP7_75t_L g1256 ( 
.A1(n_1079),
.A2(n_916),
.B(n_1145),
.Y(n_1256)
);

NOR2xp33_ASAP7_75t_L g1257 ( 
.A(n_1024),
.B(n_659),
.Y(n_1257)
);

AND2x4_ASAP7_75t_L g1258 ( 
.A(n_1101),
.B(n_1081),
.Y(n_1258)
);

CKINVDCx5p33_ASAP7_75t_R g1259 ( 
.A(n_1071),
.Y(n_1259)
);

INVx3_ASAP7_75t_L g1260 ( 
.A(n_1101),
.Y(n_1260)
);

AOI21xp5_ASAP7_75t_L g1261 ( 
.A1(n_1128),
.A2(n_680),
.B(n_786),
.Y(n_1261)
);

BUFx2_ASAP7_75t_R g1262 ( 
.A(n_1071),
.Y(n_1262)
);

NOR3xp33_ASAP7_75t_L g1263 ( 
.A(n_1018),
.B(n_887),
.C(n_659),
.Y(n_1263)
);

AOI21xp5_ASAP7_75t_L g1264 ( 
.A1(n_1128),
.A2(n_680),
.B(n_786),
.Y(n_1264)
);

AOI21xp5_ASAP7_75t_L g1265 ( 
.A1(n_1128),
.A2(n_680),
.B(n_786),
.Y(n_1265)
);

AOI221x1_ASAP7_75t_L g1266 ( 
.A1(n_1094),
.A2(n_1009),
.B1(n_887),
.B2(n_825),
.C(n_1078),
.Y(n_1266)
);

AND2x2_ASAP7_75t_L g1267 ( 
.A(n_1024),
.B(n_507),
.Y(n_1267)
);

AOI221xp5_ASAP7_75t_SL g1268 ( 
.A1(n_1018),
.A2(n_1009),
.B1(n_1070),
.B2(n_1093),
.C(n_1086),
.Y(n_1268)
);

INVx4_ASAP7_75t_L g1269 ( 
.A(n_1106),
.Y(n_1269)
);

OAI22xp5_ASAP7_75t_L g1270 ( 
.A1(n_1009),
.A2(n_1024),
.B1(n_887),
.B2(n_1002),
.Y(n_1270)
);

AOI21xp5_ASAP7_75t_L g1271 ( 
.A1(n_1128),
.A2(n_680),
.B(n_786),
.Y(n_1271)
);

BUFx3_ASAP7_75t_L g1272 ( 
.A(n_1005),
.Y(n_1272)
);

AND2x4_ASAP7_75t_L g1273 ( 
.A(n_1101),
.B(n_1081),
.Y(n_1273)
);

BUFx4_ASAP7_75t_SL g1274 ( 
.A(n_1029),
.Y(n_1274)
);

INVx1_ASAP7_75t_L g1275 ( 
.A(n_1030),
.Y(n_1275)
);

CKINVDCx5p33_ASAP7_75t_R g1276 ( 
.A(n_1071),
.Y(n_1276)
);

AO32x2_ASAP7_75t_L g1277 ( 
.A1(n_1091),
.A2(n_1094),
.A3(n_1093),
.B1(n_1070),
.B2(n_1126),
.Y(n_1277)
);

INVx2_ASAP7_75t_SL g1278 ( 
.A(n_1005),
.Y(n_1278)
);

AOI21xp5_ASAP7_75t_L g1279 ( 
.A1(n_1128),
.A2(n_680),
.B(n_786),
.Y(n_1279)
);

OAI21xp5_ASAP7_75t_SL g1280 ( 
.A1(n_1018),
.A2(n_887),
.B(n_659),
.Y(n_1280)
);

AOI22x1_ASAP7_75t_L g1281 ( 
.A1(n_1064),
.A2(n_922),
.B1(n_1125),
.B2(n_1114),
.Y(n_1281)
);

NOR3xp33_ASAP7_75t_L g1282 ( 
.A(n_1018),
.B(n_887),
.C(n_659),
.Y(n_1282)
);

O2A1O1Ixp33_ASAP7_75t_SL g1283 ( 
.A1(n_1009),
.A2(n_1018),
.B(n_1078),
.C(n_1051),
.Y(n_1283)
);

AOI22xp5_ASAP7_75t_L g1284 ( 
.A1(n_1009),
.A2(n_887),
.B1(n_659),
.B2(n_1086),
.Y(n_1284)
);

AOI21xp5_ASAP7_75t_L g1285 ( 
.A1(n_1128),
.A2(n_680),
.B(n_786),
.Y(n_1285)
);

INVx3_ASAP7_75t_SL g1286 ( 
.A(n_1029),
.Y(n_1286)
);

NAND2xp5_ASAP7_75t_L g1287 ( 
.A(n_1009),
.B(n_1023),
.Y(n_1287)
);

CKINVDCx20_ASAP7_75t_R g1288 ( 
.A(n_1071),
.Y(n_1288)
);

AOI21xp5_ASAP7_75t_L g1289 ( 
.A1(n_1128),
.A2(n_680),
.B(n_786),
.Y(n_1289)
);

CKINVDCx6p67_ASAP7_75t_R g1290 ( 
.A(n_1286),
.Y(n_1290)
);

CKINVDCx20_ASAP7_75t_R g1291 ( 
.A(n_1177),
.Y(n_1291)
);

BUFx3_ASAP7_75t_L g1292 ( 
.A(n_1288),
.Y(n_1292)
);

BUFx6f_ASAP7_75t_L g1293 ( 
.A(n_1150),
.Y(n_1293)
);

INVx1_ASAP7_75t_SL g1294 ( 
.A(n_1239),
.Y(n_1294)
);

BUFx2_ASAP7_75t_SL g1295 ( 
.A(n_1155),
.Y(n_1295)
);

BUFx6f_ASAP7_75t_L g1296 ( 
.A(n_1150),
.Y(n_1296)
);

INVx3_ASAP7_75t_SL g1297 ( 
.A(n_1192),
.Y(n_1297)
);

INVx4_ASAP7_75t_SL g1298 ( 
.A(n_1216),
.Y(n_1298)
);

INVx6_ASAP7_75t_L g1299 ( 
.A(n_1162),
.Y(n_1299)
);

INVx3_ASAP7_75t_L g1300 ( 
.A(n_1269),
.Y(n_1300)
);

INVx1_ASAP7_75t_L g1301 ( 
.A(n_1157),
.Y(n_1301)
);

AOI22xp33_ASAP7_75t_L g1302 ( 
.A1(n_1263),
.A2(n_1282),
.B1(n_1241),
.B2(n_1236),
.Y(n_1302)
);

CKINVDCx5p33_ASAP7_75t_R g1303 ( 
.A(n_1259),
.Y(n_1303)
);

AOI22xp33_ASAP7_75t_L g1304 ( 
.A1(n_1230),
.A2(n_1257),
.B1(n_1225),
.B2(n_1284),
.Y(n_1304)
);

OAI22xp5_ASAP7_75t_L g1305 ( 
.A1(n_1248),
.A2(n_1284),
.B1(n_1170),
.B2(n_1251),
.Y(n_1305)
);

AOI22xp33_ASAP7_75t_SL g1306 ( 
.A1(n_1163),
.A2(n_1270),
.B1(n_1154),
.B2(n_1186),
.Y(n_1306)
);

AOI22xp33_ASAP7_75t_L g1307 ( 
.A1(n_1248),
.A2(n_1242),
.B1(n_1170),
.B2(n_1154),
.Y(n_1307)
);

NAND2xp5_ASAP7_75t_L g1308 ( 
.A(n_1228),
.B(n_1231),
.Y(n_1308)
);

OAI22xp5_ASAP7_75t_L g1309 ( 
.A1(n_1245),
.A2(n_1249),
.B1(n_1287),
.B2(n_1156),
.Y(n_1309)
);

OAI21xp5_ASAP7_75t_SL g1310 ( 
.A1(n_1280),
.A2(n_1171),
.B(n_1186),
.Y(n_1310)
);

INVx1_ASAP7_75t_L g1311 ( 
.A(n_1158),
.Y(n_1311)
);

INVx6_ASAP7_75t_L g1312 ( 
.A(n_1162),
.Y(n_1312)
);

BUFx2_ASAP7_75t_L g1313 ( 
.A(n_1243),
.Y(n_1313)
);

CKINVDCx6p67_ASAP7_75t_R g1314 ( 
.A(n_1272),
.Y(n_1314)
);

CKINVDCx11_ASAP7_75t_R g1315 ( 
.A(n_1239),
.Y(n_1315)
);

INVx1_ASAP7_75t_L g1316 ( 
.A(n_1164),
.Y(n_1316)
);

BUFx3_ASAP7_75t_L g1317 ( 
.A(n_1276),
.Y(n_1317)
);

BUFx4_ASAP7_75t_SL g1318 ( 
.A(n_1210),
.Y(n_1318)
);

INVx1_ASAP7_75t_L g1319 ( 
.A(n_1165),
.Y(n_1319)
);

INVx6_ASAP7_75t_L g1320 ( 
.A(n_1269),
.Y(n_1320)
);

CKINVDCx11_ASAP7_75t_R g1321 ( 
.A(n_1200),
.Y(n_1321)
);

AOI22xp33_ASAP7_75t_L g1322 ( 
.A1(n_1226),
.A2(n_1244),
.B1(n_1174),
.B2(n_1202),
.Y(n_1322)
);

INVx4_ASAP7_75t_L g1323 ( 
.A(n_1150),
.Y(n_1323)
);

INVx1_ASAP7_75t_L g1324 ( 
.A(n_1234),
.Y(n_1324)
);

BUFx2_ASAP7_75t_L g1325 ( 
.A(n_1193),
.Y(n_1325)
);

OAI22xp33_ASAP7_75t_R g1326 ( 
.A1(n_1173),
.A2(n_1190),
.B1(n_1235),
.B2(n_1201),
.Y(n_1326)
);

AOI22xp33_ASAP7_75t_SL g1327 ( 
.A1(n_1267),
.A2(n_1168),
.B1(n_1244),
.B2(n_1149),
.Y(n_1327)
);

AOI22xp33_ASAP7_75t_L g1328 ( 
.A1(n_1222),
.A2(n_1176),
.B1(n_1280),
.B2(n_1181),
.Y(n_1328)
);

AOI22xp33_ASAP7_75t_L g1329 ( 
.A1(n_1222),
.A2(n_1233),
.B1(n_1247),
.B2(n_1183),
.Y(n_1329)
);

INVx3_ASAP7_75t_L g1330 ( 
.A(n_1227),
.Y(n_1330)
);

CKINVDCx6p67_ASAP7_75t_R g1331 ( 
.A(n_1200),
.Y(n_1331)
);

AOI22xp33_ASAP7_75t_L g1332 ( 
.A1(n_1233),
.A2(n_1247),
.B1(n_1195),
.B2(n_1185),
.Y(n_1332)
);

CKINVDCx5p33_ASAP7_75t_R g1333 ( 
.A(n_1191),
.Y(n_1333)
);

INVx3_ASAP7_75t_L g1334 ( 
.A(n_1227),
.Y(n_1334)
);

INVx1_ASAP7_75t_SL g1335 ( 
.A(n_1262),
.Y(n_1335)
);

AOI22xp33_ASAP7_75t_L g1336 ( 
.A1(n_1268),
.A2(n_1169),
.B1(n_1148),
.B2(n_1229),
.Y(n_1336)
);

CKINVDCx20_ASAP7_75t_R g1337 ( 
.A(n_1207),
.Y(n_1337)
);

CKINVDCx5p33_ASAP7_75t_R g1338 ( 
.A(n_1274),
.Y(n_1338)
);

BUFx4f_ASAP7_75t_SL g1339 ( 
.A(n_1178),
.Y(n_1339)
);

INVx2_ASAP7_75t_SL g1340 ( 
.A(n_1278),
.Y(n_1340)
);

INVxp67_ASAP7_75t_SL g1341 ( 
.A(n_1212),
.Y(n_1341)
);

AOI22xp33_ASAP7_75t_L g1342 ( 
.A1(n_1268),
.A2(n_1224),
.B1(n_1238),
.B2(n_1172),
.Y(n_1342)
);

INVx1_ASAP7_75t_L g1343 ( 
.A(n_1252),
.Y(n_1343)
);

BUFx8_ASAP7_75t_SL g1344 ( 
.A(n_1217),
.Y(n_1344)
);

CKINVDCx6p67_ASAP7_75t_R g1345 ( 
.A(n_1178),
.Y(n_1345)
);

INVx3_ASAP7_75t_L g1346 ( 
.A(n_1260),
.Y(n_1346)
);

BUFx12f_ASAP7_75t_L g1347 ( 
.A(n_1217),
.Y(n_1347)
);

INVx5_ASAP7_75t_SL g1348 ( 
.A(n_1210),
.Y(n_1348)
);

AOI22xp33_ASAP7_75t_SL g1349 ( 
.A1(n_1277),
.A2(n_1237),
.B1(n_1266),
.B2(n_1180),
.Y(n_1349)
);

INVx1_ASAP7_75t_L g1350 ( 
.A(n_1275),
.Y(n_1350)
);

CKINVDCx20_ASAP7_75t_R g1351 ( 
.A(n_1206),
.Y(n_1351)
);

AOI22xp5_ASAP7_75t_L g1352 ( 
.A1(n_1237),
.A2(n_1218),
.B1(n_1196),
.B2(n_1220),
.Y(n_1352)
);

BUFx2_ASAP7_75t_L g1353 ( 
.A(n_1153),
.Y(n_1353)
);

INVx1_ASAP7_75t_SL g1354 ( 
.A(n_1205),
.Y(n_1354)
);

AND2x2_ASAP7_75t_L g1355 ( 
.A(n_1221),
.B(n_1258),
.Y(n_1355)
);

AOI21xp5_ASAP7_75t_L g1356 ( 
.A1(n_1159),
.A2(n_1182),
.B(n_1223),
.Y(n_1356)
);

BUFx6f_ASAP7_75t_L g1357 ( 
.A(n_1178),
.Y(n_1357)
);

CKINVDCx5p33_ASAP7_75t_R g1358 ( 
.A(n_1258),
.Y(n_1358)
);

INVx6_ASAP7_75t_L g1359 ( 
.A(n_1273),
.Y(n_1359)
);

INVx2_ASAP7_75t_L g1360 ( 
.A(n_1209),
.Y(n_1360)
);

INVx6_ASAP7_75t_L g1361 ( 
.A(n_1273),
.Y(n_1361)
);

INVx2_ASAP7_75t_L g1362 ( 
.A(n_1204),
.Y(n_1362)
);

OAI22xp33_ASAP7_75t_L g1363 ( 
.A1(n_1180),
.A2(n_1215),
.B1(n_1277),
.B2(n_1188),
.Y(n_1363)
);

AOI22xp33_ASAP7_75t_L g1364 ( 
.A1(n_1161),
.A2(n_1213),
.B1(n_1281),
.B2(n_1277),
.Y(n_1364)
);

INVx6_ASAP7_75t_L g1365 ( 
.A(n_1210),
.Y(n_1365)
);

CKINVDCx6p67_ASAP7_75t_R g1366 ( 
.A(n_1208),
.Y(n_1366)
);

NAND3xp33_ASAP7_75t_L g1367 ( 
.A(n_1179),
.B(n_1175),
.C(n_1283),
.Y(n_1367)
);

CKINVDCx11_ASAP7_75t_R g1368 ( 
.A(n_1211),
.Y(n_1368)
);

INVx2_ASAP7_75t_SL g1369 ( 
.A(n_1216),
.Y(n_1369)
);

AOI22xp33_ASAP7_75t_L g1370 ( 
.A1(n_1147),
.A2(n_1289),
.B1(n_1253),
.B2(n_1254),
.Y(n_1370)
);

INVx1_ASAP7_75t_L g1371 ( 
.A(n_1199),
.Y(n_1371)
);

HB1xp67_ASAP7_75t_L g1372 ( 
.A(n_1203),
.Y(n_1372)
);

AOI22xp5_ASAP7_75t_L g1373 ( 
.A1(n_1167),
.A2(n_1187),
.B1(n_1214),
.B2(n_1197),
.Y(n_1373)
);

AOI22xp33_ASAP7_75t_SL g1374 ( 
.A1(n_1147),
.A2(n_1285),
.B1(n_1240),
.B2(n_1279),
.Y(n_1374)
);

INVx1_ASAP7_75t_L g1375 ( 
.A(n_1199),
.Y(n_1375)
);

CKINVDCx6p67_ASAP7_75t_R g1376 ( 
.A(n_1194),
.Y(n_1376)
);

INVx2_ASAP7_75t_L g1377 ( 
.A(n_1203),
.Y(n_1377)
);

CKINVDCx11_ASAP7_75t_R g1378 ( 
.A(n_1151),
.Y(n_1378)
);

AOI22xp33_ASAP7_75t_L g1379 ( 
.A1(n_1255),
.A2(n_1265),
.B1(n_1261),
.B2(n_1264),
.Y(n_1379)
);

OAI22xp5_ASAP7_75t_L g1380 ( 
.A1(n_1271),
.A2(n_1160),
.B1(n_1166),
.B2(n_1246),
.Y(n_1380)
);

INVx1_ASAP7_75t_L g1381 ( 
.A(n_1219),
.Y(n_1381)
);

BUFx2_ASAP7_75t_L g1382 ( 
.A(n_1198),
.Y(n_1382)
);

AOI22xp33_ASAP7_75t_L g1383 ( 
.A1(n_1152),
.A2(n_1232),
.B1(n_1250),
.B2(n_1219),
.Y(n_1383)
);

INVx1_ASAP7_75t_L g1384 ( 
.A(n_1219),
.Y(n_1384)
);

BUFx2_ASAP7_75t_L g1385 ( 
.A(n_1198),
.Y(n_1385)
);

OAI22xp33_ASAP7_75t_L g1386 ( 
.A1(n_1232),
.A2(n_1250),
.B1(n_1184),
.B2(n_1189),
.Y(n_1386)
);

AOI22xp33_ASAP7_75t_L g1387 ( 
.A1(n_1232),
.A2(n_1250),
.B1(n_1256),
.B2(n_1146),
.Y(n_1387)
);

INVx2_ASAP7_75t_R g1388 ( 
.A(n_1184),
.Y(n_1388)
);

BUFx10_ASAP7_75t_L g1389 ( 
.A(n_1201),
.Y(n_1389)
);

CKINVDCx11_ASAP7_75t_R g1390 ( 
.A(n_1177),
.Y(n_1390)
);

AOI22xp33_ASAP7_75t_L g1391 ( 
.A1(n_1263),
.A2(n_1282),
.B1(n_1241),
.B2(n_1230),
.Y(n_1391)
);

NAND2xp5_ASAP7_75t_L g1392 ( 
.A(n_1230),
.B(n_1236),
.Y(n_1392)
);

INVx6_ASAP7_75t_L g1393 ( 
.A(n_1162),
.Y(n_1393)
);

CKINVDCx5p33_ASAP7_75t_R g1394 ( 
.A(n_1259),
.Y(n_1394)
);

AOI22xp33_ASAP7_75t_L g1395 ( 
.A1(n_1263),
.A2(n_1282),
.B1(n_1241),
.B2(n_1230),
.Y(n_1395)
);

AOI22xp33_ASAP7_75t_L g1396 ( 
.A1(n_1263),
.A2(n_1282),
.B1(n_1241),
.B2(n_1230),
.Y(n_1396)
);

BUFx4f_ASAP7_75t_L g1397 ( 
.A(n_1286),
.Y(n_1397)
);

BUFx8_ASAP7_75t_SL g1398 ( 
.A(n_1177),
.Y(n_1398)
);

OAI22x1_ASAP7_75t_SL g1399 ( 
.A1(n_1259),
.A2(n_615),
.B1(n_469),
.B2(n_582),
.Y(n_1399)
);

BUFx6f_ASAP7_75t_L g1400 ( 
.A(n_1150),
.Y(n_1400)
);

INVx6_ASAP7_75t_L g1401 ( 
.A(n_1162),
.Y(n_1401)
);

BUFx6f_ASAP7_75t_L g1402 ( 
.A(n_1150),
.Y(n_1402)
);

INVx6_ASAP7_75t_L g1403 ( 
.A(n_1162),
.Y(n_1403)
);

AOI22xp5_ASAP7_75t_L g1404 ( 
.A1(n_1230),
.A2(n_1241),
.B1(n_1257),
.B2(n_1236),
.Y(n_1404)
);

AOI22xp33_ASAP7_75t_SL g1405 ( 
.A1(n_1230),
.A2(n_1236),
.B1(n_1257),
.B2(n_1241),
.Y(n_1405)
);

AOI22xp33_ASAP7_75t_SL g1406 ( 
.A1(n_1230),
.A2(n_1236),
.B1(n_1257),
.B2(n_1241),
.Y(n_1406)
);

INVx1_ASAP7_75t_L g1407 ( 
.A(n_1157),
.Y(n_1407)
);

INVxp67_ASAP7_75t_L g1408 ( 
.A(n_1153),
.Y(n_1408)
);

BUFx4f_ASAP7_75t_SL g1409 ( 
.A(n_1177),
.Y(n_1409)
);

NAND2xp5_ASAP7_75t_L g1410 ( 
.A(n_1230),
.B(n_1236),
.Y(n_1410)
);

BUFx12f_ASAP7_75t_L g1411 ( 
.A(n_1390),
.Y(n_1411)
);

INVx1_ASAP7_75t_L g1412 ( 
.A(n_1371),
.Y(n_1412)
);

INVx1_ASAP7_75t_L g1413 ( 
.A(n_1375),
.Y(n_1413)
);

OR2x2_ASAP7_75t_L g1414 ( 
.A(n_1381),
.B(n_1384),
.Y(n_1414)
);

BUFx3_ASAP7_75t_L g1415 ( 
.A(n_1344),
.Y(n_1415)
);

INVx1_ASAP7_75t_L g1416 ( 
.A(n_1377),
.Y(n_1416)
);

OAI22xp5_ASAP7_75t_L g1417 ( 
.A1(n_1405),
.A2(n_1406),
.B1(n_1404),
.B2(n_1304),
.Y(n_1417)
);

BUFx3_ASAP7_75t_L g1418 ( 
.A(n_1347),
.Y(n_1418)
);

AND2x4_ASAP7_75t_L g1419 ( 
.A(n_1298),
.B(n_1369),
.Y(n_1419)
);

INVx1_ASAP7_75t_L g1420 ( 
.A(n_1372),
.Y(n_1420)
);

INVx2_ASAP7_75t_L g1421 ( 
.A(n_1301),
.Y(n_1421)
);

AOI21x1_ASAP7_75t_L g1422 ( 
.A1(n_1380),
.A2(n_1356),
.B(n_1382),
.Y(n_1422)
);

INVx2_ASAP7_75t_SL g1423 ( 
.A(n_1365),
.Y(n_1423)
);

CKINVDCx16_ASAP7_75t_R g1424 ( 
.A(n_1351),
.Y(n_1424)
);

NOR2xp33_ASAP7_75t_L g1425 ( 
.A(n_1392),
.B(n_1410),
.Y(n_1425)
);

INVx2_ASAP7_75t_L g1426 ( 
.A(n_1311),
.Y(n_1426)
);

INVxp67_ASAP7_75t_L g1427 ( 
.A(n_1353),
.Y(n_1427)
);

NAND2x1p5_ASAP7_75t_L g1428 ( 
.A(n_1373),
.B(n_1385),
.Y(n_1428)
);

AO21x2_ASAP7_75t_L g1429 ( 
.A1(n_1386),
.A2(n_1363),
.B(n_1310),
.Y(n_1429)
);

INVx2_ASAP7_75t_L g1430 ( 
.A(n_1316),
.Y(n_1430)
);

OA21x2_ASAP7_75t_L g1431 ( 
.A1(n_1370),
.A2(n_1364),
.B(n_1379),
.Y(n_1431)
);

INVx1_ASAP7_75t_L g1432 ( 
.A(n_1372),
.Y(n_1432)
);

AND2x2_ASAP7_75t_L g1433 ( 
.A(n_1349),
.B(n_1307),
.Y(n_1433)
);

OR2x2_ASAP7_75t_L g1434 ( 
.A(n_1383),
.B(n_1307),
.Y(n_1434)
);

INVx1_ASAP7_75t_L g1435 ( 
.A(n_1341),
.Y(n_1435)
);

AOI221xp5_ASAP7_75t_L g1436 ( 
.A1(n_1304),
.A2(n_1395),
.B1(n_1396),
.B2(n_1302),
.C(n_1391),
.Y(n_1436)
);

BUFx4f_ASAP7_75t_L g1437 ( 
.A(n_1365),
.Y(n_1437)
);

INVx2_ASAP7_75t_L g1438 ( 
.A(n_1319),
.Y(n_1438)
);

INVx2_ASAP7_75t_L g1439 ( 
.A(n_1324),
.Y(n_1439)
);

INVx2_ASAP7_75t_L g1440 ( 
.A(n_1343),
.Y(n_1440)
);

INVx2_ASAP7_75t_L g1441 ( 
.A(n_1350),
.Y(n_1441)
);

AND2x2_ASAP7_75t_L g1442 ( 
.A(n_1349),
.B(n_1322),
.Y(n_1442)
);

OR2x2_ASAP7_75t_L g1443 ( 
.A(n_1383),
.B(n_1322),
.Y(n_1443)
);

HB1xp67_ASAP7_75t_L g1444 ( 
.A(n_1294),
.Y(n_1444)
);

HB1xp67_ASAP7_75t_L g1445 ( 
.A(n_1313),
.Y(n_1445)
);

INVx1_ASAP7_75t_L g1446 ( 
.A(n_1407),
.Y(n_1446)
);

INVx1_ASAP7_75t_L g1447 ( 
.A(n_1386),
.Y(n_1447)
);

AND2x2_ASAP7_75t_L g1448 ( 
.A(n_1306),
.B(n_1328),
.Y(n_1448)
);

INVx1_ASAP7_75t_L g1449 ( 
.A(n_1329),
.Y(n_1449)
);

AND2x2_ASAP7_75t_L g1450 ( 
.A(n_1306),
.B(n_1328),
.Y(n_1450)
);

INVx1_ASAP7_75t_L g1451 ( 
.A(n_1329),
.Y(n_1451)
);

INVx2_ASAP7_75t_SL g1452 ( 
.A(n_1299),
.Y(n_1452)
);

INVx1_ASAP7_75t_L g1453 ( 
.A(n_1388),
.Y(n_1453)
);

CKINVDCx20_ASAP7_75t_R g1454 ( 
.A(n_1398),
.Y(n_1454)
);

INVx1_ASAP7_75t_L g1455 ( 
.A(n_1388),
.Y(n_1455)
);

INVx1_ASAP7_75t_L g1456 ( 
.A(n_1387),
.Y(n_1456)
);

INVx1_ASAP7_75t_L g1457 ( 
.A(n_1387),
.Y(n_1457)
);

INVx1_ASAP7_75t_L g1458 ( 
.A(n_1367),
.Y(n_1458)
);

BUFx2_ASAP7_75t_L g1459 ( 
.A(n_1352),
.Y(n_1459)
);

BUFx6f_ASAP7_75t_L g1460 ( 
.A(n_1299),
.Y(n_1460)
);

AND2x2_ASAP7_75t_L g1461 ( 
.A(n_1327),
.B(n_1336),
.Y(n_1461)
);

INVx1_ASAP7_75t_L g1462 ( 
.A(n_1332),
.Y(n_1462)
);

OAI21x1_ASAP7_75t_L g1463 ( 
.A1(n_1379),
.A2(n_1370),
.B(n_1364),
.Y(n_1463)
);

INVx1_ASAP7_75t_L g1464 ( 
.A(n_1332),
.Y(n_1464)
);

AND2x2_ASAP7_75t_L g1465 ( 
.A(n_1327),
.B(n_1336),
.Y(n_1465)
);

INVx2_ASAP7_75t_SL g1466 ( 
.A(n_1312),
.Y(n_1466)
);

NAND2xp5_ASAP7_75t_L g1467 ( 
.A(n_1309),
.B(n_1302),
.Y(n_1467)
);

INVx1_ASAP7_75t_SL g1468 ( 
.A(n_1315),
.Y(n_1468)
);

INVx1_ASAP7_75t_L g1469 ( 
.A(n_1363),
.Y(n_1469)
);

AND2x2_ASAP7_75t_L g1470 ( 
.A(n_1391),
.B(n_1395),
.Y(n_1470)
);

INVx1_ASAP7_75t_L g1471 ( 
.A(n_1342),
.Y(n_1471)
);

OA21x2_ASAP7_75t_L g1472 ( 
.A1(n_1342),
.A2(n_1396),
.B(n_1305),
.Y(n_1472)
);

BUFx2_ASAP7_75t_L g1473 ( 
.A(n_1298),
.Y(n_1473)
);

OR2x6_ASAP7_75t_L g1474 ( 
.A(n_1312),
.B(n_1393),
.Y(n_1474)
);

NAND2xp5_ASAP7_75t_L g1475 ( 
.A(n_1405),
.B(n_1406),
.Y(n_1475)
);

INVx1_ASAP7_75t_L g1476 ( 
.A(n_1376),
.Y(n_1476)
);

OAI21xp5_ASAP7_75t_L g1477 ( 
.A1(n_1308),
.A2(n_1374),
.B(n_1408),
.Y(n_1477)
);

AND2x2_ASAP7_75t_L g1478 ( 
.A(n_1360),
.B(n_1362),
.Y(n_1478)
);

INVx1_ASAP7_75t_L g1479 ( 
.A(n_1374),
.Y(n_1479)
);

AOI22xp33_ASAP7_75t_L g1480 ( 
.A1(n_1378),
.A2(n_1326),
.B1(n_1325),
.B2(n_1337),
.Y(n_1480)
);

AND2x2_ASAP7_75t_L g1481 ( 
.A(n_1330),
.B(n_1334),
.Y(n_1481)
);

BUFx2_ASAP7_75t_L g1482 ( 
.A(n_1408),
.Y(n_1482)
);

INVx1_ASAP7_75t_L g1483 ( 
.A(n_1346),
.Y(n_1483)
);

OR2x2_ASAP7_75t_L g1484 ( 
.A(n_1354),
.B(n_1348),
.Y(n_1484)
);

A2O1A1Ixp33_ASAP7_75t_SL g1485 ( 
.A1(n_1300),
.A2(n_1355),
.B(n_1399),
.C(n_1318),
.Y(n_1485)
);

NAND2x1_ASAP7_75t_L g1486 ( 
.A(n_1401),
.B(n_1403),
.Y(n_1486)
);

BUFx2_ASAP7_75t_SL g1487 ( 
.A(n_1389),
.Y(n_1487)
);

NAND2x1p5_ASAP7_75t_L g1488 ( 
.A(n_1300),
.B(n_1397),
.Y(n_1488)
);

CKINVDCx5p33_ASAP7_75t_R g1489 ( 
.A(n_1321),
.Y(n_1489)
);

OAI21xp5_ASAP7_75t_L g1490 ( 
.A1(n_1436),
.A2(n_1397),
.B(n_1335),
.Y(n_1490)
);

OA21x2_ASAP7_75t_L g1491 ( 
.A1(n_1463),
.A2(n_1340),
.B(n_1358),
.Y(n_1491)
);

A2O1A1Ixp33_ASAP7_75t_L g1492 ( 
.A1(n_1417),
.A2(n_1318),
.B(n_1295),
.C(n_1317),
.Y(n_1492)
);

AND2x2_ASAP7_75t_L g1493 ( 
.A(n_1459),
.B(n_1292),
.Y(n_1493)
);

NOR2xp33_ASAP7_75t_SL g1494 ( 
.A(n_1411),
.B(n_1409),
.Y(n_1494)
);

AND2x2_ASAP7_75t_L g1495 ( 
.A(n_1459),
.B(n_1445),
.Y(n_1495)
);

OAI211xp5_ASAP7_75t_L g1496 ( 
.A1(n_1475),
.A2(n_1368),
.B(n_1394),
.C(n_1303),
.Y(n_1496)
);

OR2x2_ASAP7_75t_L g1497 ( 
.A(n_1421),
.B(n_1331),
.Y(n_1497)
);

NAND4xp25_ASAP7_75t_L g1498 ( 
.A(n_1425),
.B(n_1323),
.C(n_1290),
.D(n_1314),
.Y(n_1498)
);

NAND2xp33_ASAP7_75t_L g1499 ( 
.A(n_1467),
.B(n_1470),
.Y(n_1499)
);

INVxp67_ASAP7_75t_L g1500 ( 
.A(n_1444),
.Y(n_1500)
);

AOI221xp5_ASAP7_75t_L g1501 ( 
.A1(n_1470),
.A2(n_1338),
.B1(n_1333),
.B2(n_1297),
.C(n_1291),
.Y(n_1501)
);

OR2x2_ASAP7_75t_L g1502 ( 
.A(n_1421),
.B(n_1297),
.Y(n_1502)
);

O2A1O1Ixp33_ASAP7_75t_L g1503 ( 
.A1(n_1485),
.A2(n_1458),
.B(n_1477),
.C(n_1450),
.Y(n_1503)
);

NOR2xp33_ASAP7_75t_L g1504 ( 
.A(n_1458),
.B(n_1361),
.Y(n_1504)
);

OR2x2_ASAP7_75t_L g1505 ( 
.A(n_1426),
.B(n_1366),
.Y(n_1505)
);

INVx4_ASAP7_75t_L g1506 ( 
.A(n_1474),
.Y(n_1506)
);

AND2x2_ASAP7_75t_L g1507 ( 
.A(n_1429),
.B(n_1479),
.Y(n_1507)
);

INVx2_ASAP7_75t_L g1508 ( 
.A(n_1426),
.Y(n_1508)
);

AND2x2_ASAP7_75t_L g1509 ( 
.A(n_1429),
.B(n_1402),
.Y(n_1509)
);

O2A1O1Ixp33_ASAP7_75t_SL g1510 ( 
.A1(n_1476),
.A2(n_1403),
.B(n_1401),
.C(n_1320),
.Y(n_1510)
);

OAI21xp5_ASAP7_75t_L g1511 ( 
.A1(n_1472),
.A2(n_1323),
.B(n_1409),
.Y(n_1511)
);

A2O1A1Ixp33_ASAP7_75t_L g1512 ( 
.A1(n_1448),
.A2(n_1402),
.B(n_1296),
.C(n_1357),
.Y(n_1512)
);

NAND2xp5_ASAP7_75t_L g1513 ( 
.A(n_1482),
.B(n_1478),
.Y(n_1513)
);

AND2x2_ASAP7_75t_L g1514 ( 
.A(n_1479),
.B(n_1400),
.Y(n_1514)
);

OR2x6_ASAP7_75t_L g1515 ( 
.A(n_1428),
.B(n_1320),
.Y(n_1515)
);

INVx4_ASAP7_75t_L g1516 ( 
.A(n_1474),
.Y(n_1516)
);

BUFx2_ASAP7_75t_L g1517 ( 
.A(n_1484),
.Y(n_1517)
);

AOI21xp5_ASAP7_75t_L g1518 ( 
.A1(n_1437),
.A2(n_1293),
.B(n_1296),
.Y(n_1518)
);

AOI22xp5_ASAP7_75t_L g1519 ( 
.A1(n_1450),
.A2(n_1359),
.B1(n_1320),
.B2(n_1339),
.Y(n_1519)
);

A2O1A1Ixp33_ASAP7_75t_L g1520 ( 
.A1(n_1461),
.A2(n_1293),
.B(n_1296),
.C(n_1357),
.Y(n_1520)
);

OAI21xp5_ASAP7_75t_L g1521 ( 
.A1(n_1472),
.A2(n_1359),
.B(n_1345),
.Y(n_1521)
);

AOI21xp5_ASAP7_75t_L g1522 ( 
.A1(n_1437),
.A2(n_1357),
.B(n_1339),
.Y(n_1522)
);

AO32x2_ASAP7_75t_L g1523 ( 
.A1(n_1423),
.A2(n_1466),
.A3(n_1452),
.B1(n_1469),
.B2(n_1432),
.Y(n_1523)
);

HB1xp67_ASAP7_75t_L g1524 ( 
.A(n_1483),
.Y(n_1524)
);

AND2x2_ASAP7_75t_L g1525 ( 
.A(n_1456),
.B(n_1457),
.Y(n_1525)
);

CKINVDCx5p33_ASAP7_75t_R g1526 ( 
.A(n_1454),
.Y(n_1526)
);

NAND2xp5_ASAP7_75t_L g1527 ( 
.A(n_1427),
.B(n_1461),
.Y(n_1527)
);

INVx2_ASAP7_75t_L g1528 ( 
.A(n_1430),
.Y(n_1528)
);

OR2x2_ASAP7_75t_L g1529 ( 
.A(n_1430),
.B(n_1438),
.Y(n_1529)
);

AND2x4_ASAP7_75t_L g1530 ( 
.A(n_1419),
.B(n_1473),
.Y(n_1530)
);

OAI21x1_ASAP7_75t_SL g1531 ( 
.A1(n_1471),
.A2(n_1472),
.B(n_1423),
.Y(n_1531)
);

AND2x2_ASAP7_75t_SL g1532 ( 
.A(n_1431),
.B(n_1442),
.Y(n_1532)
);

AO32x2_ASAP7_75t_L g1533 ( 
.A1(n_1452),
.A2(n_1466),
.A3(n_1469),
.B1(n_1420),
.B2(n_1432),
.Y(n_1533)
);

AOI22xp5_ASAP7_75t_L g1534 ( 
.A1(n_1472),
.A2(n_1465),
.B1(n_1480),
.B2(n_1442),
.Y(n_1534)
);

AND2x2_ASAP7_75t_L g1535 ( 
.A(n_1481),
.B(n_1438),
.Y(n_1535)
);

A2O1A1Ixp33_ASAP7_75t_L g1536 ( 
.A1(n_1465),
.A2(n_1463),
.B(n_1433),
.C(n_1471),
.Y(n_1536)
);

AND2x2_ASAP7_75t_L g1537 ( 
.A(n_1439),
.B(n_1440),
.Y(n_1537)
);

AND2x2_ASAP7_75t_L g1538 ( 
.A(n_1449),
.B(n_1451),
.Y(n_1538)
);

AOI221xp5_ASAP7_75t_L g1539 ( 
.A1(n_1447),
.A2(n_1451),
.B1(n_1464),
.B2(n_1462),
.C(n_1443),
.Y(n_1539)
);

OR2x2_ASAP7_75t_L g1540 ( 
.A(n_1440),
.B(n_1441),
.Y(n_1540)
);

BUFx10_ASAP7_75t_L g1541 ( 
.A(n_1476),
.Y(n_1541)
);

OR2x2_ASAP7_75t_L g1542 ( 
.A(n_1507),
.B(n_1435),
.Y(n_1542)
);

AND2x2_ASAP7_75t_L g1543 ( 
.A(n_1507),
.B(n_1453),
.Y(n_1543)
);

INVx2_ASAP7_75t_L g1544 ( 
.A(n_1508),
.Y(n_1544)
);

NOR2xp33_ASAP7_75t_L g1545 ( 
.A(n_1496),
.B(n_1424),
.Y(n_1545)
);

CKINVDCx20_ASAP7_75t_R g1546 ( 
.A(n_1526),
.Y(n_1546)
);

AND2x2_ASAP7_75t_L g1547 ( 
.A(n_1532),
.B(n_1453),
.Y(n_1547)
);

INVxp67_ASAP7_75t_SL g1548 ( 
.A(n_1524),
.Y(n_1548)
);

INVx4_ASAP7_75t_L g1549 ( 
.A(n_1515),
.Y(n_1549)
);

AND2x2_ASAP7_75t_L g1550 ( 
.A(n_1532),
.B(n_1455),
.Y(n_1550)
);

NAND2xp5_ASAP7_75t_L g1551 ( 
.A(n_1538),
.B(n_1462),
.Y(n_1551)
);

AND2x2_ASAP7_75t_L g1552 ( 
.A(n_1533),
.B(n_1455),
.Y(n_1552)
);

AND2x2_ASAP7_75t_L g1553 ( 
.A(n_1533),
.B(n_1422),
.Y(n_1553)
);

AND2x2_ASAP7_75t_SL g1554 ( 
.A(n_1499),
.B(n_1431),
.Y(n_1554)
);

OAI21xp33_ASAP7_75t_L g1555 ( 
.A1(n_1499),
.A2(n_1443),
.B(n_1434),
.Y(n_1555)
);

AOI22xp33_ASAP7_75t_SL g1556 ( 
.A1(n_1490),
.A2(n_1431),
.B1(n_1428),
.B2(n_1434),
.Y(n_1556)
);

NAND2xp5_ASAP7_75t_SL g1557 ( 
.A(n_1492),
.B(n_1437),
.Y(n_1557)
);

HB1xp67_ASAP7_75t_L g1558 ( 
.A(n_1528),
.Y(n_1558)
);

INVx2_ASAP7_75t_SL g1559 ( 
.A(n_1530),
.Y(n_1559)
);

AND2x2_ASAP7_75t_L g1560 ( 
.A(n_1533),
.B(n_1431),
.Y(n_1560)
);

AND2x2_ASAP7_75t_L g1561 ( 
.A(n_1523),
.B(n_1412),
.Y(n_1561)
);

AND2x2_ASAP7_75t_L g1562 ( 
.A(n_1523),
.B(n_1413),
.Y(n_1562)
);

INVx1_ASAP7_75t_L g1563 ( 
.A(n_1529),
.Y(n_1563)
);

OAI22xp33_ASAP7_75t_L g1564 ( 
.A1(n_1534),
.A2(n_1428),
.B1(n_1424),
.B2(n_1484),
.Y(n_1564)
);

OR2x2_ASAP7_75t_L g1565 ( 
.A(n_1525),
.B(n_1414),
.Y(n_1565)
);

AND2x2_ASAP7_75t_L g1566 ( 
.A(n_1523),
.B(n_1416),
.Y(n_1566)
);

INVx1_ASAP7_75t_SL g1567 ( 
.A(n_1502),
.Y(n_1567)
);

NOR2xp33_ASAP7_75t_L g1568 ( 
.A(n_1498),
.B(n_1468),
.Y(n_1568)
);

NAND2xp5_ASAP7_75t_L g1569 ( 
.A(n_1539),
.B(n_1446),
.Y(n_1569)
);

AOI22xp33_ASAP7_75t_SL g1570 ( 
.A1(n_1511),
.A2(n_1411),
.B1(n_1489),
.B2(n_1487),
.Y(n_1570)
);

AND2x2_ASAP7_75t_L g1571 ( 
.A(n_1547),
.B(n_1517),
.Y(n_1571)
);

NAND2xp5_ASAP7_75t_L g1572 ( 
.A(n_1563),
.B(n_1537),
.Y(n_1572)
);

NAND2xp5_ASAP7_75t_L g1573 ( 
.A(n_1563),
.B(n_1536),
.Y(n_1573)
);

INVx1_ASAP7_75t_L g1574 ( 
.A(n_1558),
.Y(n_1574)
);

INVx1_ASAP7_75t_L g1575 ( 
.A(n_1558),
.Y(n_1575)
);

INVx2_ASAP7_75t_L g1576 ( 
.A(n_1566),
.Y(n_1576)
);

OAI22xp5_ASAP7_75t_L g1577 ( 
.A1(n_1556),
.A2(n_1555),
.B1(n_1492),
.B2(n_1536),
.Y(n_1577)
);

AND2x2_ASAP7_75t_L g1578 ( 
.A(n_1547),
.B(n_1509),
.Y(n_1578)
);

INVx1_ASAP7_75t_L g1579 ( 
.A(n_1544),
.Y(n_1579)
);

AND2x2_ASAP7_75t_L g1580 ( 
.A(n_1550),
.B(n_1509),
.Y(n_1580)
);

AND2x2_ASAP7_75t_L g1581 ( 
.A(n_1550),
.B(n_1495),
.Y(n_1581)
);

BUFx2_ASAP7_75t_L g1582 ( 
.A(n_1548),
.Y(n_1582)
);

OR2x2_ASAP7_75t_L g1583 ( 
.A(n_1565),
.B(n_1513),
.Y(n_1583)
);

NOR2xp33_ASAP7_75t_SL g1584 ( 
.A(n_1555),
.B(n_1506),
.Y(n_1584)
);

INVx2_ASAP7_75t_L g1585 ( 
.A(n_1566),
.Y(n_1585)
);

AOI22xp33_ASAP7_75t_L g1586 ( 
.A1(n_1556),
.A2(n_1493),
.B1(n_1506),
.B2(n_1516),
.Y(n_1586)
);

AND2x2_ASAP7_75t_L g1587 ( 
.A(n_1550),
.B(n_1491),
.Y(n_1587)
);

AND3x1_ASAP7_75t_L g1588 ( 
.A(n_1545),
.B(n_1494),
.C(n_1501),
.Y(n_1588)
);

INVx2_ASAP7_75t_L g1589 ( 
.A(n_1566),
.Y(n_1589)
);

HB1xp67_ASAP7_75t_L g1590 ( 
.A(n_1542),
.Y(n_1590)
);

NOR2xp33_ASAP7_75t_L g1591 ( 
.A(n_1568),
.B(n_1500),
.Y(n_1591)
);

BUFx6f_ASAP7_75t_L g1592 ( 
.A(n_1554),
.Y(n_1592)
);

AND2x2_ASAP7_75t_L g1593 ( 
.A(n_1567),
.B(n_1491),
.Y(n_1593)
);

AND2x4_ASAP7_75t_L g1594 ( 
.A(n_1549),
.B(n_1530),
.Y(n_1594)
);

NAND2xp5_ASAP7_75t_L g1595 ( 
.A(n_1551),
.B(n_1535),
.Y(n_1595)
);

NOR2x1_ASAP7_75t_L g1596 ( 
.A(n_1549),
.B(n_1515),
.Y(n_1596)
);

OAI222xp33_ASAP7_75t_L g1597 ( 
.A1(n_1570),
.A2(n_1503),
.B1(n_1519),
.B2(n_1527),
.C1(n_1515),
.C2(n_1497),
.Y(n_1597)
);

NAND3xp33_ASAP7_75t_SL g1598 ( 
.A(n_1570),
.B(n_1521),
.C(n_1520),
.Y(n_1598)
);

NAND2xp5_ASAP7_75t_L g1599 ( 
.A(n_1551),
.B(n_1540),
.Y(n_1599)
);

AOI221xp5_ASAP7_75t_L g1600 ( 
.A1(n_1564),
.A2(n_1504),
.B1(n_1531),
.B2(n_1514),
.C(n_1510),
.Y(n_1600)
);

AOI22xp33_ASAP7_75t_L g1601 ( 
.A1(n_1564),
.A2(n_1516),
.B1(n_1506),
.B2(n_1515),
.Y(n_1601)
);

INVxp67_ASAP7_75t_L g1602 ( 
.A(n_1573),
.Y(n_1602)
);

INVx1_ASAP7_75t_L g1603 ( 
.A(n_1590),
.Y(n_1603)
);

NAND2xp5_ASAP7_75t_L g1604 ( 
.A(n_1573),
.B(n_1552),
.Y(n_1604)
);

HB1xp67_ASAP7_75t_L g1605 ( 
.A(n_1582),
.Y(n_1605)
);

NAND2xp5_ASAP7_75t_L g1606 ( 
.A(n_1582),
.B(n_1552),
.Y(n_1606)
);

INVx2_ASAP7_75t_L g1607 ( 
.A(n_1576),
.Y(n_1607)
);

INVxp67_ASAP7_75t_L g1608 ( 
.A(n_1591),
.Y(n_1608)
);

INVx1_ASAP7_75t_L g1609 ( 
.A(n_1574),
.Y(n_1609)
);

INVx2_ASAP7_75t_L g1610 ( 
.A(n_1576),
.Y(n_1610)
);

INVx1_ASAP7_75t_L g1611 ( 
.A(n_1574),
.Y(n_1611)
);

INVx1_ASAP7_75t_L g1612 ( 
.A(n_1575),
.Y(n_1612)
);

BUFx2_ASAP7_75t_L g1613 ( 
.A(n_1596),
.Y(n_1613)
);

AND2x2_ASAP7_75t_L g1614 ( 
.A(n_1578),
.B(n_1559),
.Y(n_1614)
);

AND2x4_ASAP7_75t_SL g1615 ( 
.A(n_1571),
.B(n_1541),
.Y(n_1615)
);

INVx1_ASAP7_75t_L g1616 ( 
.A(n_1575),
.Y(n_1616)
);

INVx2_ASAP7_75t_L g1617 ( 
.A(n_1576),
.Y(n_1617)
);

AND2x2_ASAP7_75t_L g1618 ( 
.A(n_1578),
.B(n_1567),
.Y(n_1618)
);

AND2x2_ASAP7_75t_L g1619 ( 
.A(n_1580),
.B(n_1543),
.Y(n_1619)
);

NAND2xp5_ASAP7_75t_L g1620 ( 
.A(n_1593),
.B(n_1552),
.Y(n_1620)
);

AND2x4_ASAP7_75t_L g1621 ( 
.A(n_1596),
.B(n_1549),
.Y(n_1621)
);

OAI211xp5_ASAP7_75t_SL g1622 ( 
.A1(n_1577),
.A2(n_1569),
.B(n_1557),
.C(n_1505),
.Y(n_1622)
);

NAND2xp5_ASAP7_75t_L g1623 ( 
.A(n_1593),
.B(n_1561),
.Y(n_1623)
);

INVx1_ASAP7_75t_SL g1624 ( 
.A(n_1571),
.Y(n_1624)
);

AND2x4_ASAP7_75t_L g1625 ( 
.A(n_1592),
.B(n_1561),
.Y(n_1625)
);

AND2x4_ASAP7_75t_L g1626 ( 
.A(n_1592),
.B(n_1562),
.Y(n_1626)
);

NAND2xp5_ASAP7_75t_L g1627 ( 
.A(n_1595),
.B(n_1562),
.Y(n_1627)
);

AND2x2_ASAP7_75t_L g1628 ( 
.A(n_1592),
.B(n_1554),
.Y(n_1628)
);

AND2x2_ASAP7_75t_L g1629 ( 
.A(n_1592),
.B(n_1554),
.Y(n_1629)
);

INVx1_ASAP7_75t_L g1630 ( 
.A(n_1609),
.Y(n_1630)
);

OR2x2_ASAP7_75t_L g1631 ( 
.A(n_1602),
.B(n_1583),
.Y(n_1631)
);

INVxp67_ASAP7_75t_L g1632 ( 
.A(n_1605),
.Y(n_1632)
);

AND2x2_ASAP7_75t_L g1633 ( 
.A(n_1628),
.B(n_1592),
.Y(n_1633)
);

INVx1_ASAP7_75t_L g1634 ( 
.A(n_1609),
.Y(n_1634)
);

AND2x2_ASAP7_75t_L g1635 ( 
.A(n_1628),
.B(n_1587),
.Y(n_1635)
);

AND2x2_ASAP7_75t_L g1636 ( 
.A(n_1625),
.B(n_1585),
.Y(n_1636)
);

NOR2xp33_ASAP7_75t_SL g1637 ( 
.A(n_1613),
.B(n_1597),
.Y(n_1637)
);

INVx2_ASAP7_75t_SL g1638 ( 
.A(n_1615),
.Y(n_1638)
);

AND2x2_ASAP7_75t_L g1639 ( 
.A(n_1625),
.B(n_1585),
.Y(n_1639)
);

AND2x2_ASAP7_75t_L g1640 ( 
.A(n_1629),
.B(n_1587),
.Y(n_1640)
);

INVx2_ASAP7_75t_L g1641 ( 
.A(n_1607),
.Y(n_1641)
);

INVx2_ASAP7_75t_L g1642 ( 
.A(n_1607),
.Y(n_1642)
);

OAI21xp5_ASAP7_75t_L g1643 ( 
.A1(n_1622),
.A2(n_1577),
.B(n_1588),
.Y(n_1643)
);

AND2x2_ASAP7_75t_L g1644 ( 
.A(n_1629),
.B(n_1589),
.Y(n_1644)
);

NAND2x1p5_ASAP7_75t_L g1645 ( 
.A(n_1613),
.B(n_1621),
.Y(n_1645)
);

INVx1_ASAP7_75t_L g1646 ( 
.A(n_1611),
.Y(n_1646)
);

NAND2xp5_ASAP7_75t_L g1647 ( 
.A(n_1602),
.B(n_1599),
.Y(n_1647)
);

AND2x2_ASAP7_75t_L g1648 ( 
.A(n_1625),
.B(n_1594),
.Y(n_1648)
);

AND2x2_ASAP7_75t_L g1649 ( 
.A(n_1625),
.B(n_1560),
.Y(n_1649)
);

AOI21xp5_ASAP7_75t_L g1650 ( 
.A1(n_1622),
.A2(n_1598),
.B(n_1584),
.Y(n_1650)
);

INVx1_ASAP7_75t_L g1651 ( 
.A(n_1611),
.Y(n_1651)
);

INVx1_ASAP7_75t_L g1652 ( 
.A(n_1612),
.Y(n_1652)
);

AND2x2_ASAP7_75t_L g1653 ( 
.A(n_1626),
.B(n_1560),
.Y(n_1653)
);

INVx1_ASAP7_75t_L g1654 ( 
.A(n_1612),
.Y(n_1654)
);

NAND2xp5_ASAP7_75t_L g1655 ( 
.A(n_1604),
.B(n_1599),
.Y(n_1655)
);

INVx1_ASAP7_75t_L g1656 ( 
.A(n_1616),
.Y(n_1656)
);

OR2x2_ASAP7_75t_L g1657 ( 
.A(n_1604),
.B(n_1583),
.Y(n_1657)
);

INVx1_ASAP7_75t_L g1658 ( 
.A(n_1616),
.Y(n_1658)
);

NAND2xp5_ASAP7_75t_L g1659 ( 
.A(n_1603),
.B(n_1581),
.Y(n_1659)
);

AOI21xp33_ASAP7_75t_SL g1660 ( 
.A1(n_1608),
.A2(n_1489),
.B(n_1526),
.Y(n_1660)
);

OR2x2_ASAP7_75t_L g1661 ( 
.A(n_1603),
.B(n_1572),
.Y(n_1661)
);

NAND2xp5_ASAP7_75t_L g1662 ( 
.A(n_1608),
.B(n_1581),
.Y(n_1662)
);

INVx2_ASAP7_75t_L g1663 ( 
.A(n_1607),
.Y(n_1663)
);

NAND2xp5_ASAP7_75t_L g1664 ( 
.A(n_1627),
.B(n_1579),
.Y(n_1664)
);

NOR2xp33_ASAP7_75t_SL g1665 ( 
.A(n_1621),
.B(n_1584),
.Y(n_1665)
);

INVx2_ASAP7_75t_L g1666 ( 
.A(n_1610),
.Y(n_1666)
);

INVx2_ASAP7_75t_L g1667 ( 
.A(n_1610),
.Y(n_1667)
);

AND2x4_ASAP7_75t_L g1668 ( 
.A(n_1621),
.B(n_1594),
.Y(n_1668)
);

AND2x2_ASAP7_75t_L g1669 ( 
.A(n_1626),
.B(n_1594),
.Y(n_1669)
);

NAND3xp33_ASAP7_75t_L g1670 ( 
.A(n_1606),
.B(n_1588),
.C(n_1600),
.Y(n_1670)
);

OR2x2_ASAP7_75t_L g1671 ( 
.A(n_1631),
.B(n_1620),
.Y(n_1671)
);

INVx2_ASAP7_75t_L g1672 ( 
.A(n_1636),
.Y(n_1672)
);

AND2x2_ASAP7_75t_L g1673 ( 
.A(n_1633),
.B(n_1626),
.Y(n_1673)
);

INVx2_ASAP7_75t_L g1674 ( 
.A(n_1636),
.Y(n_1674)
);

INVx1_ASAP7_75t_L g1675 ( 
.A(n_1630),
.Y(n_1675)
);

NAND2xp5_ASAP7_75t_L g1676 ( 
.A(n_1643),
.B(n_1624),
.Y(n_1676)
);

INVx2_ASAP7_75t_L g1677 ( 
.A(n_1636),
.Y(n_1677)
);

OR2x2_ASAP7_75t_L g1678 ( 
.A(n_1631),
.B(n_1620),
.Y(n_1678)
);

NAND2xp5_ASAP7_75t_L g1679 ( 
.A(n_1643),
.B(n_1624),
.Y(n_1679)
);

INVx1_ASAP7_75t_L g1680 ( 
.A(n_1630),
.Y(n_1680)
);

NAND2xp5_ASAP7_75t_L g1681 ( 
.A(n_1662),
.B(n_1618),
.Y(n_1681)
);

INVx1_ASAP7_75t_L g1682 ( 
.A(n_1634),
.Y(n_1682)
);

AOI21xp5_ASAP7_75t_L g1683 ( 
.A1(n_1637),
.A2(n_1621),
.B(n_1510),
.Y(n_1683)
);

OR2x2_ASAP7_75t_L g1684 ( 
.A(n_1657),
.B(n_1623),
.Y(n_1684)
);

AND2x2_ASAP7_75t_SL g1685 ( 
.A(n_1637),
.B(n_1586),
.Y(n_1685)
);

OR2x2_ASAP7_75t_L g1686 ( 
.A(n_1657),
.B(n_1662),
.Y(n_1686)
);

INVxp67_ASAP7_75t_L g1687 ( 
.A(n_1650),
.Y(n_1687)
);

AND2x2_ASAP7_75t_L g1688 ( 
.A(n_1633),
.B(n_1626),
.Y(n_1688)
);

INVx1_ASAP7_75t_L g1689 ( 
.A(n_1634),
.Y(n_1689)
);

INVx1_ASAP7_75t_L g1690 ( 
.A(n_1646),
.Y(n_1690)
);

AND2x2_ASAP7_75t_L g1691 ( 
.A(n_1648),
.B(n_1615),
.Y(n_1691)
);

INVx1_ASAP7_75t_SL g1692 ( 
.A(n_1638),
.Y(n_1692)
);

AOI21xp33_ASAP7_75t_L g1693 ( 
.A1(n_1670),
.A2(n_1601),
.B(n_1569),
.Y(n_1693)
);

INVxp67_ASAP7_75t_L g1694 ( 
.A(n_1650),
.Y(n_1694)
);

AND2x2_ASAP7_75t_L g1695 ( 
.A(n_1648),
.B(n_1615),
.Y(n_1695)
);

OAI22x1_ASAP7_75t_L g1696 ( 
.A1(n_1670),
.A2(n_1606),
.B1(n_1618),
.B2(n_1614),
.Y(n_1696)
);

OR2x2_ASAP7_75t_L g1697 ( 
.A(n_1647),
.B(n_1623),
.Y(n_1697)
);

INVx2_ASAP7_75t_L g1698 ( 
.A(n_1639),
.Y(n_1698)
);

AND2x2_ASAP7_75t_L g1699 ( 
.A(n_1669),
.B(n_1619),
.Y(n_1699)
);

NOR2xp33_ASAP7_75t_L g1700 ( 
.A(n_1660),
.B(n_1546),
.Y(n_1700)
);

INVx1_ASAP7_75t_L g1701 ( 
.A(n_1646),
.Y(n_1701)
);

INVx1_ASAP7_75t_L g1702 ( 
.A(n_1651),
.Y(n_1702)
);

INVx2_ASAP7_75t_L g1703 ( 
.A(n_1639),
.Y(n_1703)
);

INVx1_ASAP7_75t_L g1704 ( 
.A(n_1651),
.Y(n_1704)
);

OAI21xp5_ASAP7_75t_L g1705 ( 
.A1(n_1665),
.A2(n_1512),
.B(n_1553),
.Y(n_1705)
);

NAND2xp5_ASAP7_75t_L g1706 ( 
.A(n_1647),
.B(n_1619),
.Y(n_1706)
);

INVx1_ASAP7_75t_L g1707 ( 
.A(n_1675),
.Y(n_1707)
);

INVx1_ASAP7_75t_L g1708 ( 
.A(n_1675),
.Y(n_1708)
);

NAND2xp5_ASAP7_75t_L g1709 ( 
.A(n_1687),
.B(n_1632),
.Y(n_1709)
);

INVx1_ASAP7_75t_L g1710 ( 
.A(n_1680),
.Y(n_1710)
);

INVx1_ASAP7_75t_SL g1711 ( 
.A(n_1692),
.Y(n_1711)
);

INVx2_ASAP7_75t_SL g1712 ( 
.A(n_1673),
.Y(n_1712)
);

AOI21xp5_ASAP7_75t_L g1713 ( 
.A1(n_1685),
.A2(n_1665),
.B(n_1660),
.Y(n_1713)
);

NOR2xp33_ASAP7_75t_L g1714 ( 
.A(n_1700),
.B(n_1415),
.Y(n_1714)
);

NAND2xp33_ASAP7_75t_SL g1715 ( 
.A(n_1676),
.B(n_1679),
.Y(n_1715)
);

NOR2xp33_ASAP7_75t_SL g1716 ( 
.A(n_1694),
.B(n_1638),
.Y(n_1716)
);

NAND2xp5_ASAP7_75t_L g1717 ( 
.A(n_1693),
.B(n_1632),
.Y(n_1717)
);

INVx1_ASAP7_75t_L g1718 ( 
.A(n_1680),
.Y(n_1718)
);

INVx1_ASAP7_75t_L g1719 ( 
.A(n_1682),
.Y(n_1719)
);

INVx1_ASAP7_75t_L g1720 ( 
.A(n_1682),
.Y(n_1720)
);

NOR3xp33_ASAP7_75t_L g1721 ( 
.A(n_1683),
.B(n_1638),
.C(n_1415),
.Y(n_1721)
);

NAND2xp5_ASAP7_75t_L g1722 ( 
.A(n_1685),
.B(n_1655),
.Y(n_1722)
);

NOR2xp33_ASAP7_75t_L g1723 ( 
.A(n_1685),
.B(n_1655),
.Y(n_1723)
);

INVx1_ASAP7_75t_L g1724 ( 
.A(n_1689),
.Y(n_1724)
);

AOI221xp5_ASAP7_75t_L g1725 ( 
.A1(n_1696),
.A2(n_1645),
.B1(n_1656),
.B2(n_1658),
.C(n_1654),
.Y(n_1725)
);

AND2x2_ASAP7_75t_L g1726 ( 
.A(n_1673),
.B(n_1669),
.Y(n_1726)
);

OAI22xp33_ASAP7_75t_SL g1727 ( 
.A1(n_1686),
.A2(n_1645),
.B1(n_1668),
.B2(n_1659),
.Y(n_1727)
);

AOI21xp33_ASAP7_75t_SL g1728 ( 
.A1(n_1696),
.A2(n_1645),
.B(n_1668),
.Y(n_1728)
);

OAI321xp33_ASAP7_75t_L g1729 ( 
.A1(n_1705),
.A2(n_1645),
.A3(n_1659),
.B1(n_1658),
.B2(n_1652),
.C(n_1654),
.Y(n_1729)
);

AOI21xp5_ASAP7_75t_L g1730 ( 
.A1(n_1681),
.A2(n_1656),
.B(n_1652),
.Y(n_1730)
);

OAI21xp5_ASAP7_75t_SL g1731 ( 
.A1(n_1688),
.A2(n_1668),
.B(n_1640),
.Y(n_1731)
);

NAND2xp5_ASAP7_75t_SL g1732 ( 
.A(n_1688),
.B(n_1668),
.Y(n_1732)
);

NOR2xp33_ASAP7_75t_L g1733 ( 
.A(n_1686),
.B(n_1706),
.Y(n_1733)
);

AOI222xp33_ASAP7_75t_L g1734 ( 
.A1(n_1715),
.A2(n_1698),
.B1(n_1703),
.B2(n_1677),
.C1(n_1674),
.C2(n_1672),
.Y(n_1734)
);

INVx1_ASAP7_75t_SL g1735 ( 
.A(n_1711),
.Y(n_1735)
);

INVxp67_ASAP7_75t_SL g1736 ( 
.A(n_1723),
.Y(n_1736)
);

OAI22xp33_ASAP7_75t_L g1737 ( 
.A1(n_1722),
.A2(n_1697),
.B1(n_1678),
.B2(n_1671),
.Y(n_1737)
);

OAI211xp5_ASAP7_75t_L g1738 ( 
.A1(n_1725),
.A2(n_1704),
.B(n_1689),
.C(n_1702),
.Y(n_1738)
);

A2O1A1Ixp33_ASAP7_75t_L g1739 ( 
.A1(n_1713),
.A2(n_1697),
.B(n_1671),
.C(n_1678),
.Y(n_1739)
);

AND2x2_ASAP7_75t_L g1740 ( 
.A(n_1726),
.B(n_1691),
.Y(n_1740)
);

INVx1_ASAP7_75t_L g1741 ( 
.A(n_1707),
.Y(n_1741)
);

AO22x1_ASAP7_75t_L g1742 ( 
.A1(n_1723),
.A2(n_1695),
.B1(n_1691),
.B2(n_1702),
.Y(n_1742)
);

INVx1_ASAP7_75t_L g1743 ( 
.A(n_1708),
.Y(n_1743)
);

OAI21xp33_ASAP7_75t_L g1744 ( 
.A1(n_1717),
.A2(n_1684),
.B(n_1695),
.Y(n_1744)
);

AOI22xp5_ASAP7_75t_L g1745 ( 
.A1(n_1716),
.A2(n_1672),
.B1(n_1703),
.B2(n_1674),
.Y(n_1745)
);

INVx2_ASAP7_75t_SL g1746 ( 
.A(n_1712),
.Y(n_1746)
);

NAND2xp5_ASAP7_75t_L g1747 ( 
.A(n_1733),
.B(n_1699),
.Y(n_1747)
);

NAND3xp33_ASAP7_75t_L g1748 ( 
.A(n_1728),
.B(n_1704),
.C(n_1701),
.Y(n_1748)
);

INVx1_ASAP7_75t_L g1749 ( 
.A(n_1710),
.Y(n_1749)
);

NAND2xp5_ASAP7_75t_L g1750 ( 
.A(n_1733),
.B(n_1699),
.Y(n_1750)
);

INVx1_ASAP7_75t_SL g1751 ( 
.A(n_1709),
.Y(n_1751)
);

AOI22x1_ASAP7_75t_L g1752 ( 
.A1(n_1730),
.A2(n_1701),
.B1(n_1690),
.B2(n_1684),
.Y(n_1752)
);

OAI21xp33_ASAP7_75t_L g1753 ( 
.A1(n_1727),
.A2(n_1698),
.B(n_1677),
.Y(n_1753)
);

AOI21xp33_ASAP7_75t_L g1754 ( 
.A1(n_1736),
.A2(n_1729),
.B(n_1714),
.Y(n_1754)
);

INVx1_ASAP7_75t_L g1755 ( 
.A(n_1741),
.Y(n_1755)
);

OAI22xp33_ASAP7_75t_L g1756 ( 
.A1(n_1745),
.A2(n_1731),
.B1(n_1732),
.B2(n_1661),
.Y(n_1756)
);

NAND2xp5_ASAP7_75t_SL g1757 ( 
.A(n_1735),
.B(n_1721),
.Y(n_1757)
);

NAND2xp5_ASAP7_75t_SL g1758 ( 
.A(n_1737),
.B(n_1721),
.Y(n_1758)
);

OAI22xp5_ASAP7_75t_L g1759 ( 
.A1(n_1736),
.A2(n_1661),
.B1(n_1649),
.B2(n_1653),
.Y(n_1759)
);

NAND2xp5_ASAP7_75t_L g1760 ( 
.A(n_1746),
.B(n_1744),
.Y(n_1760)
);

INVx1_ASAP7_75t_L g1761 ( 
.A(n_1743),
.Y(n_1761)
);

OAI22xp33_ASAP7_75t_SL g1762 ( 
.A1(n_1752),
.A2(n_1724),
.B1(n_1720),
.B2(n_1719),
.Y(n_1762)
);

OR2x2_ASAP7_75t_L g1763 ( 
.A(n_1747),
.B(n_1718),
.Y(n_1763)
);

AOI22xp5_ASAP7_75t_L g1764 ( 
.A1(n_1740),
.A2(n_1690),
.B1(n_1635),
.B2(n_1640),
.Y(n_1764)
);

INVx2_ASAP7_75t_L g1765 ( 
.A(n_1763),
.Y(n_1765)
);

O2A1O1Ixp5_ASAP7_75t_L g1766 ( 
.A1(n_1758),
.A2(n_1742),
.B(n_1738),
.C(n_1748),
.Y(n_1766)
);

NAND3xp33_ASAP7_75t_L g1767 ( 
.A(n_1754),
.B(n_1734),
.C(n_1739),
.Y(n_1767)
);

INVx2_ASAP7_75t_SL g1768 ( 
.A(n_1757),
.Y(n_1768)
);

NAND2xp33_ASAP7_75t_SL g1769 ( 
.A(n_1760),
.B(n_1750),
.Y(n_1769)
);

NAND2xp5_ASAP7_75t_L g1770 ( 
.A(n_1756),
.B(n_1751),
.Y(n_1770)
);

NOR3xp33_ASAP7_75t_L g1771 ( 
.A(n_1762),
.B(n_1761),
.C(n_1755),
.Y(n_1771)
);

INVx2_ASAP7_75t_SL g1772 ( 
.A(n_1764),
.Y(n_1772)
);

NAND2xp5_ASAP7_75t_L g1773 ( 
.A(n_1759),
.B(n_1749),
.Y(n_1773)
);

NAND3xp33_ASAP7_75t_L g1774 ( 
.A(n_1754),
.B(n_1738),
.C(n_1753),
.Y(n_1774)
);

NAND4xp25_ASAP7_75t_L g1775 ( 
.A(n_1766),
.B(n_1418),
.C(n_1635),
.D(n_1522),
.Y(n_1775)
);

O2A1O1Ixp33_ASAP7_75t_L g1776 ( 
.A1(n_1774),
.A2(n_1667),
.B(n_1666),
.C(n_1641),
.Y(n_1776)
);

OAI211xp5_ASAP7_75t_SL g1777 ( 
.A1(n_1767),
.A2(n_1667),
.B(n_1666),
.C(n_1663),
.Y(n_1777)
);

AOI22x1_ASAP7_75t_L g1778 ( 
.A1(n_1768),
.A2(n_1487),
.B1(n_1666),
.B2(n_1663),
.Y(n_1778)
);

OAI211xp5_ASAP7_75t_L g1779 ( 
.A1(n_1770),
.A2(n_1418),
.B(n_1639),
.C(n_1649),
.Y(n_1779)
);

AOI221x1_ASAP7_75t_SL g1780 ( 
.A1(n_1775),
.A2(n_1773),
.B1(n_1765),
.B2(n_1771),
.C(n_1769),
.Y(n_1780)
);

INVx1_ASAP7_75t_L g1781 ( 
.A(n_1777),
.Y(n_1781)
);

INVxp33_ASAP7_75t_SL g1782 ( 
.A(n_1778),
.Y(n_1782)
);

INVx1_ASAP7_75t_L g1783 ( 
.A(n_1779),
.Y(n_1783)
);

NAND2x1_ASAP7_75t_L g1784 ( 
.A(n_1776),
.B(n_1772),
.Y(n_1784)
);

INVxp67_ASAP7_75t_SL g1785 ( 
.A(n_1775),
.Y(n_1785)
);

NAND2xp5_ASAP7_75t_L g1786 ( 
.A(n_1780),
.B(n_1644),
.Y(n_1786)
);

INVx1_ASAP7_75t_L g1787 ( 
.A(n_1784),
.Y(n_1787)
);

INVx2_ASAP7_75t_L g1788 ( 
.A(n_1783),
.Y(n_1788)
);

NAND2x1p5_ASAP7_75t_L g1789 ( 
.A(n_1781),
.B(n_1486),
.Y(n_1789)
);

INVxp67_ASAP7_75t_L g1790 ( 
.A(n_1785),
.Y(n_1790)
);

XNOR2xp5_ASAP7_75t_L g1791 ( 
.A(n_1787),
.B(n_1782),
.Y(n_1791)
);

AOI221xp5_ASAP7_75t_L g1792 ( 
.A1(n_1790),
.A2(n_1782),
.B1(n_1667),
.B2(n_1663),
.C(n_1641),
.Y(n_1792)
);

AND2x4_ASAP7_75t_L g1793 ( 
.A(n_1788),
.B(n_1644),
.Y(n_1793)
);

NAND2xp5_ASAP7_75t_L g1794 ( 
.A(n_1793),
.B(n_1786),
.Y(n_1794)
);

NOR4xp25_ASAP7_75t_L g1795 ( 
.A(n_1794),
.B(n_1792),
.C(n_1791),
.D(n_1789),
.Y(n_1795)
);

XNOR2x1_ASAP7_75t_L g1796 ( 
.A(n_1795),
.B(n_1488),
.Y(n_1796)
);

XNOR2xp5_ASAP7_75t_L g1797 ( 
.A(n_1795),
.B(n_1488),
.Y(n_1797)
);

INVxp67_ASAP7_75t_L g1798 ( 
.A(n_1796),
.Y(n_1798)
);

NOR2x1p5_ASAP7_75t_L g1799 ( 
.A(n_1797),
.B(n_1486),
.Y(n_1799)
);

INVx1_ASAP7_75t_L g1800 ( 
.A(n_1798),
.Y(n_1800)
);

NAND2xp5_ASAP7_75t_L g1801 ( 
.A(n_1799),
.B(n_1641),
.Y(n_1801)
);

NAND2xp5_ASAP7_75t_L g1802 ( 
.A(n_1800),
.B(n_1642),
.Y(n_1802)
);

NAND2xp5_ASAP7_75t_L g1803 ( 
.A(n_1802),
.B(n_1801),
.Y(n_1803)
);

OAI22xp33_ASAP7_75t_L g1804 ( 
.A1(n_1803),
.A2(n_1642),
.B1(n_1664),
.B2(n_1617),
.Y(n_1804)
);

OAI221xp5_ASAP7_75t_R g1805 ( 
.A1(n_1804),
.A2(n_1642),
.B1(n_1653),
.B2(n_1649),
.C(n_1541),
.Y(n_1805)
);

AOI211xp5_ASAP7_75t_L g1806 ( 
.A1(n_1805),
.A2(n_1518),
.B(n_1653),
.C(n_1460),
.Y(n_1806)
);


endmodule