module real_jpeg_27174_n_21 (n_17, n_108, n_8, n_0, n_111, n_2, n_10, n_114, n_9, n_12, n_107, n_6, n_106, n_11, n_14, n_110, n_112, n_7, n_18, n_3, n_5, n_4, n_105, n_109, n_1, n_20, n_19, n_16, n_15, n_13, n_113, n_21);

input n_17;
input n_108;
input n_8;
input n_0;
input n_111;
input n_2;
input n_10;
input n_114;
input n_9;
input n_12;
input n_107;
input n_6;
input n_106;
input n_11;
input n_14;
input n_110;
input n_112;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_105;
input n_109;
input n_1;
input n_20;
input n_19;
input n_16;
input n_15;
input n_13;
input n_113;

output n_21;

wire n_54;
wire n_37;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_68;
wire n_83;
wire n_78;
wire n_64;
wire n_47;
wire n_22;
wire n_87;
wire n_40;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_93;
wire n_95;
wire n_65;
wire n_33;
wire n_76;
wire n_67;
wire n_79;
wire n_66;
wire n_28;
wire n_44;
wire n_62;
wire n_45;
wire n_42;
wire n_77;
wire n_39;
wire n_94;
wire n_26;
wire n_50;
wire n_69;
wire n_31;
wire n_72;
wire n_100;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_30;
wire n_103;
wire n_43;
wire n_57;
wire n_84;
wire n_82;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_24;
wire n_92;
wire n_97;
wire n_75;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_25;
wire n_53;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_101;
wire n_96;
wire n_89;

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_0),
.B(n_71),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_0),
.B(n_71),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_1),
.B(n_58),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_1),
.B(n_58),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_2),
.B(n_61),
.Y(n_60)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

BUFx12_ASAP7_75t_L g41 ( 
.A(n_3),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_SL g58 ( 
.A(n_3),
.B(n_59),
.Y(n_58)
);

BUFx12_ASAP7_75t_L g62 ( 
.A(n_3),
.Y(n_62)
);

OR2x2_ASAP7_75t_L g67 ( 
.A(n_3),
.B(n_68),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_4),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g35 ( 
.A(n_5),
.B(n_36),
.C(n_100),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_6),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_7),
.B(n_46),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_7),
.B(n_46),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_8),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_9),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_10),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g39 ( 
.A(n_11),
.B(n_40),
.Y(n_39)
);

OR2x2_ASAP7_75t_L g86 ( 
.A(n_11),
.B(n_40),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_12),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_13),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_14),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_SL g32 ( 
.A(n_15),
.B(n_33),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_15),
.B(n_33),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_16),
.B(n_88),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_16),
.B(n_88),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_17),
.B(n_97),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_17),
.B(n_97),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_18),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_19),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_20),
.B(n_51),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_20),
.B(n_51),
.Y(n_79)
);

XOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_31),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_30),
.Y(n_22)
);

INVxp67_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_26),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_SL g30 ( 
.A(n_25),
.B(n_26),
.Y(n_30)
);

OR2x2_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_28),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_28),
.B(n_34),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_SL g46 ( 
.A(n_28),
.B(n_47),
.Y(n_46)
);

OR2x2_ASAP7_75t_L g82 ( 
.A(n_28),
.B(n_83),
.Y(n_82)
);

OR2x2_ASAP7_75t_L g92 ( 
.A(n_28),
.B(n_93),
.Y(n_92)
);

INVx11_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_29),
.Y(n_102)
);

OAI21xp5_ASAP7_75t_L g31 ( 
.A1(n_32),
.A2(n_35),
.B(n_103),
.Y(n_31)
);

OAI21xp5_ASAP7_75t_SL g36 ( 
.A1(n_37),
.A2(n_96),
.B(n_99),
.Y(n_36)
);

AOI21xp5_ASAP7_75t_SL g37 ( 
.A1(n_38),
.A2(n_91),
.B(n_95),
.Y(n_37)
);

A2O1A1Ixp33_ASAP7_75t_SL g38 ( 
.A1(n_39),
.A2(n_43),
.B(n_87),
.C(n_90),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_SL g40 ( 
.A(n_41),
.B(n_42),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_SL g51 ( 
.A(n_41),
.B(n_52),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_SL g88 ( 
.A(n_41),
.B(n_89),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_41),
.B(n_98),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g43 ( 
.A(n_44),
.B(n_86),
.Y(n_43)
);

OAI21xp5_ASAP7_75t_L g44 ( 
.A1(n_45),
.A2(n_48),
.B(n_85),
.Y(n_44)
);

AOI21xp5_ASAP7_75t_L g48 ( 
.A1(n_49),
.A2(n_80),
.B(n_84),
.Y(n_48)
);

OAI21xp5_ASAP7_75t_L g49 ( 
.A1(n_50),
.A2(n_53),
.B(n_79),
.Y(n_49)
);

AOI21xp5_ASAP7_75t_L g53 ( 
.A1(n_54),
.A2(n_74),
.B(n_78),
.Y(n_53)
);

OAI21xp5_ASAP7_75t_SL g54 ( 
.A1(n_55),
.A2(n_70),
.B(n_73),
.Y(n_54)
);

AOI21xp5_ASAP7_75t_L g55 ( 
.A1(n_56),
.A2(n_65),
.B(n_69),
.Y(n_55)
);

OAI21xp5_ASAP7_75t_SL g56 ( 
.A1(n_57),
.A2(n_60),
.B(n_64),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_SL g61 ( 
.A(n_62),
.B(n_63),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_SL g71 ( 
.A(n_62),
.B(n_72),
.Y(n_71)
);

OR2x2_ASAP7_75t_L g76 ( 
.A(n_62),
.B(n_77),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_66),
.B(n_67),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_66),
.B(n_67),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_75),
.B(n_76),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g78 ( 
.A(n_75),
.B(n_76),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_81),
.B(n_82),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_81),
.B(n_82),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_92),
.B(n_94),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_92),
.B(n_94),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_101),
.B(n_102),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_105),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_106),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_107),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_108),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_109),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_110),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_111),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_112),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_113),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_114),
.Y(n_89)
);


endmodule