module fake_jpeg_11544_n_138 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_138);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_138;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_124;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_6),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_30),
.Y(n_40)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_37),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_33),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_36),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_6),
.Y(n_44)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_29),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_25),
.Y(n_46)
);

INVx6_ASAP7_75t_SL g47 ( 
.A(n_17),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_35),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_26),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_5),
.Y(n_50)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_19),
.Y(n_51)
);

BUFx5_ASAP7_75t_L g52 ( 
.A(n_0),
.Y(n_52)
);

BUFx5_ASAP7_75t_L g53 ( 
.A(n_38),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_20),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_7),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_42),
.Y(n_56)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_56),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_47),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_57),
.B(n_59),
.Y(n_66)
);

INVx5_ASAP7_75t_L g58 ( 
.A(n_46),
.Y(n_58)
);

INVx5_ASAP7_75t_L g71 ( 
.A(n_58),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_40),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_50),
.B(n_0),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_60),
.B(n_1),
.Y(n_70)
);

INVx4_ASAP7_75t_SL g61 ( 
.A(n_39),
.Y(n_61)
);

INVx5_ASAP7_75t_L g75 ( 
.A(n_61),
.Y(n_75)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_43),
.Y(n_62)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_62),
.Y(n_69)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_44),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_63),
.B(n_48),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_41),
.Y(n_64)
);

INVx5_ASAP7_75t_L g78 ( 
.A(n_64),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_SL g65 ( 
.A(n_56),
.B(n_55),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g79 ( 
.A(n_65),
.B(n_72),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_68),
.B(n_46),
.Y(n_80)
);

AND2x2_ASAP7_75t_L g92 ( 
.A(n_70),
.B(n_2),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_62),
.B(n_54),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_58),
.B(n_49),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_73),
.B(n_74),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_64),
.B(n_45),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_61),
.B(n_45),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_76),
.B(n_77),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_60),
.B(n_51),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_80),
.B(n_8),
.Y(n_97)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_67),
.Y(n_81)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_81),
.Y(n_100)
);

HB1xp67_ASAP7_75t_L g82 ( 
.A(n_71),
.Y(n_82)
);

HB1xp67_ASAP7_75t_L g111 ( 
.A(n_82),
.Y(n_111)
);

OA22x2_ASAP7_75t_L g84 ( 
.A1(n_69),
.A2(n_39),
.B1(n_51),
.B2(n_46),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_84),
.A2(n_95),
.B1(n_16),
.B2(n_18),
.Y(n_110)
);

BUFx2_ASAP7_75t_L g85 ( 
.A(n_71),
.Y(n_85)
);

INVx1_ASAP7_75t_SL g104 ( 
.A(n_85),
.Y(n_104)
);

NAND2xp33_ASAP7_75t_SL g87 ( 
.A(n_67),
.B(n_52),
.Y(n_87)
);

AOI21xp5_ASAP7_75t_L g108 ( 
.A1(n_87),
.A2(n_94),
.B(n_14),
.Y(n_108)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_78),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_88),
.B(n_91),
.Y(n_99)
);

OAI21xp33_ASAP7_75t_SL g89 ( 
.A1(n_75),
.A2(n_53),
.B(n_52),
.Y(n_89)
);

NAND2xp33_ASAP7_75t_SL g109 ( 
.A(n_89),
.B(n_15),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_66),
.B(n_41),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_SL g102 ( 
.A(n_90),
.B(n_92),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_75),
.B(n_1),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_78),
.B(n_2),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_93),
.B(n_13),
.Y(n_107)
);

AOI21xp5_ASAP7_75t_L g94 ( 
.A1(n_76),
.A2(n_53),
.B(n_4),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_74),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_83),
.A2(n_3),
.B1(n_7),
.B2(n_8),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_96),
.A2(n_110),
.B1(n_89),
.B2(n_22),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_SL g112 ( 
.A(n_97),
.B(n_98),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_79),
.B(n_9),
.Y(n_98)
);

AOI21xp5_ASAP7_75t_SL g101 ( 
.A1(n_86),
.A2(n_9),
.B(n_10),
.Y(n_101)
);

AND2x2_ASAP7_75t_L g122 ( 
.A(n_101),
.B(n_107),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_92),
.B(n_82),
.Y(n_103)
);

XNOR2xp5_ASAP7_75t_L g119 ( 
.A(n_103),
.B(n_105),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_84),
.B(n_11),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_SL g106 ( 
.A(n_84),
.B(n_12),
.Y(n_106)
);

CKINVDCx14_ASAP7_75t_R g118 ( 
.A(n_106),
.Y(n_118)
);

AOI21xp5_ASAP7_75t_L g117 ( 
.A1(n_108),
.A2(n_109),
.B(n_23),
.Y(n_117)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_100),
.Y(n_113)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_113),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_114),
.B(n_115),
.Y(n_124)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_111),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_99),
.B(n_21),
.Y(n_116)
);

A2O1A1O1Ixp25_ASAP7_75t_L g126 ( 
.A1(n_116),
.A2(n_121),
.B(n_101),
.C(n_27),
.D(n_28),
.Y(n_126)
);

XOR2xp5_ASAP7_75t_L g127 ( 
.A(n_117),
.B(n_120),
.Y(n_127)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_104),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_104),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_118),
.A2(n_110),
.B1(n_102),
.B2(n_109),
.Y(n_125)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_125),
.Y(n_130)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_126),
.Y(n_129)
);

XOR2xp5_ASAP7_75t_L g128 ( 
.A(n_127),
.B(n_119),
.Y(n_128)
);

AND2x2_ASAP7_75t_L g132 ( 
.A(n_128),
.B(n_124),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_L g131 ( 
.A1(n_130),
.A2(n_124),
.B(n_116),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_L g133 ( 
.A(n_131),
.B(n_132),
.Y(n_133)
);

OAI31xp33_ASAP7_75t_L g134 ( 
.A1(n_133),
.A2(n_129),
.A3(n_123),
.B(n_128),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_134),
.B(n_122),
.C(n_112),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_L g136 ( 
.A1(n_135),
.A2(n_122),
.B(n_31),
.Y(n_136)
);

OAI21xp33_ASAP7_75t_SL g137 ( 
.A1(n_136),
.A2(n_24),
.B(n_32),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_L g138 ( 
.A(n_137),
.B(n_34),
.Y(n_138)
);


endmodule