module real_aes_9016_n_105 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_104, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_103, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_105);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_104;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_103;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_105;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_555;
wire n_421;
wire n_766;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_666;
wire n_551;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_578;
wire n_528;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_774;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_535;
wire n_732;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_755;
wire n_656;
wire n_178;
wire n_409;
wire n_748;
wire n_781;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_455;
wire n_119;
wire n_504;
wire n_310;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_782;
wire n_443;
wire n_565;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_770;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_527;
wire n_769;
wire n_434;
wire n_505;
wire n_502;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_768;
wire n_176;
wire n_412;
wire n_542;
wire n_163;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_288;
wire n_147;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_749;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_419;
wire n_217;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_148;
wire n_498;
wire n_481;
wire n_765;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_679;
wire n_520;
wire n_633;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_456;
wire n_156;
wire n_359;
wire n_717;
wire n_312;
wire n_266;
wire n_183;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_521;
wire n_140;
wire n_418;
wire n_422;
wire n_771;
wire n_524;
wire n_219;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_639;
wire n_587;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_554;
wire n_475;
wire n_264;
wire n_237;
wire n_668;
A2O1A1Ixp33_ASAP7_75t_SL g523 ( .A1(n_0), .A2(n_169), .B(n_524), .C(n_527), .Y(n_523) );
NAND2xp5_ASAP7_75t_L g528 ( .A(n_1), .B(n_519), .Y(n_528) );
NAND3xp33_ASAP7_75t_SL g113 ( .A(n_2), .B(n_114), .C(n_115), .Y(n_113) );
INVx1_ASAP7_75t_L g467 ( .A(n_2), .Y(n_467) );
INVx1_ASAP7_75t_L g167 ( .A(n_3), .Y(n_167) );
NAND2xp5_ASAP7_75t_SL g592 ( .A(n_4), .B(n_170), .Y(n_592) );
AOI21xp5_ASAP7_75t_L g562 ( .A1(n_5), .A2(n_488), .B(n_563), .Y(n_562) );
OAI22xp5_ASAP7_75t_SL g770 ( .A1(n_6), .A2(n_771), .B1(n_774), .B2(n_775), .Y(n_770) );
CKINVDCx20_ASAP7_75t_R g775 ( .A(n_6), .Y(n_775) );
AO21x2_ASAP7_75t_L g541 ( .A1(n_7), .A2(n_177), .B(n_542), .Y(n_541) );
AOI22xp33_ASAP7_75t_L g223 ( .A1(n_8), .A2(n_37), .B1(n_157), .B2(n_205), .Y(n_223) );
NAND2xp5_ASAP7_75t_L g185 ( .A(n_9), .B(n_177), .Y(n_185) );
AND2x6_ASAP7_75t_L g172 ( .A(n_10), .B(n_173), .Y(n_172) );
A2O1A1Ixp33_ASAP7_75t_L g535 ( .A1(n_11), .A2(n_172), .B(n_493), .C(n_536), .Y(n_535) );
OAI22xp5_ASAP7_75t_L g771 ( .A1(n_12), .A2(n_41), .B1(n_772), .B2(n_773), .Y(n_771) );
CKINVDCx20_ASAP7_75t_R g772 ( .A(n_12), .Y(n_772) );
INVx1_ASAP7_75t_L g111 ( .A(n_13), .Y(n_111) );
NOR2xp33_ASAP7_75t_L g468 ( .A(n_13), .B(n_38), .Y(n_468) );
INVx1_ASAP7_75t_L g151 ( .A(n_14), .Y(n_151) );
INVx1_ASAP7_75t_L g148 ( .A(n_15), .Y(n_148) );
NAND2xp5_ASAP7_75t_L g214 ( .A(n_16), .B(n_153), .Y(n_214) );
NAND2xp5_ASAP7_75t_SL g547 ( .A(n_17), .B(n_170), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g251 ( .A(n_18), .B(n_144), .Y(n_251) );
AO32x2_ASAP7_75t_L g221 ( .A1(n_19), .A2(n_143), .A3(n_177), .B1(n_196), .B2(n_222), .Y(n_221) );
NAND2xp5_ASAP7_75t_SL g218 ( .A(n_20), .B(n_157), .Y(n_218) );
NAND2xp5_ASAP7_75t_L g174 ( .A(n_21), .B(n_144), .Y(n_174) );
AOI22xp33_ASAP7_75t_L g224 ( .A1(n_22), .A2(n_57), .B1(n_157), .B2(n_205), .Y(n_224) );
AOI22xp33_ASAP7_75t_SL g207 ( .A1(n_23), .A2(n_85), .B1(n_153), .B2(n_157), .Y(n_207) );
NAND2xp5_ASAP7_75t_SL g237 ( .A(n_24), .B(n_157), .Y(n_237) );
A2O1A1Ixp33_ASAP7_75t_L g510 ( .A1(n_25), .A2(n_196), .B(n_493), .C(n_511), .Y(n_510) );
A2O1A1Ixp33_ASAP7_75t_L g544 ( .A1(n_26), .A2(n_196), .B(n_493), .C(n_545), .Y(n_544) );
BUFx6f_ASAP7_75t_L g162 ( .A(n_27), .Y(n_162) );
NAND2xp5_ASAP7_75t_L g197 ( .A(n_28), .B(n_198), .Y(n_197) );
AOI22xp5_ASAP7_75t_L g767 ( .A1(n_29), .A2(n_768), .B1(n_769), .B2(n_770), .Y(n_767) );
CKINVDCx20_ASAP7_75t_R g768 ( .A(n_29), .Y(n_768) );
AOI21xp5_ASAP7_75t_L g520 ( .A1(n_30), .A2(n_488), .B(n_521), .Y(n_520) );
NAND2xp5_ASAP7_75t_L g239 ( .A(n_31), .B(n_198), .Y(n_239) );
INVx2_ASAP7_75t_L g155 ( .A(n_32), .Y(n_155) );
A2O1A1Ixp33_ASAP7_75t_L g490 ( .A1(n_33), .A2(n_491), .B(n_495), .C(n_501), .Y(n_490) );
NAND2xp5_ASAP7_75t_SL g189 ( .A(n_34), .B(n_157), .Y(n_189) );
NAND2xp5_ASAP7_75t_L g220 ( .A(n_35), .B(n_198), .Y(n_220) );
NAND2xp5_ASAP7_75t_L g546 ( .A(n_36), .B(n_216), .Y(n_546) );
NAND2xp5_ASAP7_75t_L g110 ( .A(n_38), .B(n_111), .Y(n_110) );
NAND2xp5_ASAP7_75t_L g508 ( .A(n_39), .B(n_509), .Y(n_508) );
CKINVDCx20_ASAP7_75t_R g540 ( .A(n_40), .Y(n_540) );
INVx1_ASAP7_75t_L g773 ( .A(n_41), .Y(n_773) );
NAND2xp5_ASAP7_75t_L g557 ( .A(n_42), .B(n_170), .Y(n_557) );
OAI22xp5_ASAP7_75t_SL g454 ( .A1(n_43), .A2(n_455), .B1(n_458), .B2(n_459), .Y(n_454) );
CKINVDCx20_ASAP7_75t_R g458 ( .A(n_43), .Y(n_458) );
NAND2xp5_ASAP7_75t_L g543 ( .A(n_44), .B(n_488), .Y(n_543) );
OAI22xp5_ASAP7_75t_SL g455 ( .A1(n_45), .A2(n_47), .B1(n_456), .B2(n_457), .Y(n_455) );
INVx1_ASAP7_75t_L g457 ( .A(n_45), .Y(n_457) );
OAI22xp5_ASAP7_75t_SL g475 ( .A1(n_45), .A2(n_131), .B1(n_132), .B2(n_457), .Y(n_475) );
A2O1A1Ixp33_ASAP7_75t_L g554 ( .A1(n_46), .A2(n_491), .B(n_501), .C(n_555), .Y(n_554) );
CKINVDCx20_ASAP7_75t_R g456 ( .A(n_47), .Y(n_456) );
NAND2xp5_ASAP7_75t_SL g180 ( .A(n_48), .B(n_157), .Y(n_180) );
INVx1_ASAP7_75t_L g525 ( .A(n_49), .Y(n_525) );
AOI22xp33_ASAP7_75t_L g204 ( .A1(n_50), .A2(n_94), .B1(n_205), .B2(n_206), .Y(n_204) );
NAND2xp5_ASAP7_75t_L g469 ( .A(n_51), .B(n_470), .Y(n_469) );
NAND2xp5_ASAP7_75t_SL g183 ( .A(n_52), .B(n_157), .Y(n_183) );
NAND2xp5_ASAP7_75t_L g156 ( .A(n_53), .B(n_157), .Y(n_156) );
INVx1_ASAP7_75t_L g556 ( .A(n_54), .Y(n_556) );
NAND2xp5_ASAP7_75t_L g553 ( .A(n_55), .B(n_488), .Y(n_553) );
NAND2xp5_ASAP7_75t_L g184 ( .A(n_56), .B(n_165), .Y(n_184) );
AOI22xp33_ASAP7_75t_SL g249 ( .A1(n_58), .A2(n_62), .B1(n_153), .B2(n_157), .Y(n_249) );
OAI22xp5_ASAP7_75t_SL g126 ( .A1(n_59), .A2(n_70), .B1(n_127), .B2(n_128), .Y(n_126) );
CKINVDCx20_ASAP7_75t_R g127 ( .A(n_59), .Y(n_127) );
NAND2xp5_ASAP7_75t_SL g193 ( .A(n_60), .B(n_157), .Y(n_193) );
NAND2xp5_ASAP7_75t_SL g213 ( .A(n_61), .B(n_157), .Y(n_213) );
INVx1_ASAP7_75t_L g173 ( .A(n_63), .Y(n_173) );
NAND2xp5_ASAP7_75t_L g594 ( .A(n_64), .B(n_488), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g568 ( .A(n_65), .B(n_519), .Y(n_568) );
A2O1A1Ixp33_ASAP7_75t_L g565 ( .A1(n_66), .A2(n_159), .B(n_165), .C(n_566), .Y(n_565) );
AOI22xp33_ASAP7_75t_L g105 ( .A1(n_67), .A2(n_106), .B1(n_118), .B2(n_785), .Y(n_105) );
NAND2xp5_ASAP7_75t_L g168 ( .A(n_68), .B(n_157), .Y(n_168) );
INVx1_ASAP7_75t_L g147 ( .A(n_69), .Y(n_147) );
CKINVDCx20_ASAP7_75t_R g128 ( .A(n_70), .Y(n_128) );
CKINVDCx20_ASAP7_75t_R g123 ( .A(n_71), .Y(n_123) );
NAND2xp5_ASAP7_75t_SL g499 ( .A(n_72), .B(n_170), .Y(n_499) );
AO32x2_ASAP7_75t_L g202 ( .A1(n_73), .A2(n_177), .A3(n_196), .B1(n_203), .B2(n_208), .Y(n_202) );
NAND2xp5_ASAP7_75t_L g537 ( .A(n_74), .B(n_171), .Y(n_537) );
INVx1_ASAP7_75t_L g192 ( .A(n_75), .Y(n_192) );
INVx1_ASAP7_75t_L g234 ( .A(n_76), .Y(n_234) );
CKINVDCx16_ASAP7_75t_R g522 ( .A(n_77), .Y(n_522) );
NAND2xp5_ASAP7_75t_L g512 ( .A(n_78), .B(n_498), .Y(n_512) );
A2O1A1Ixp33_ASAP7_75t_L g589 ( .A1(n_79), .A2(n_493), .B(n_501), .C(n_590), .Y(n_589) );
AOI222xp33_ASAP7_75t_L g473 ( .A1(n_80), .A2(n_474), .B1(n_766), .B2(n_767), .C1(n_776), .C2(n_780), .Y(n_473) );
NAND2xp5_ASAP7_75t_SL g235 ( .A(n_81), .B(n_153), .Y(n_235) );
CKINVDCx16_ASAP7_75t_R g564 ( .A(n_82), .Y(n_564) );
INVx1_ASAP7_75t_L g117 ( .A(n_83), .Y(n_117) );
NAND2xp5_ASAP7_75t_SL g513 ( .A(n_84), .B(n_497), .Y(n_513) );
NAND2xp5_ASAP7_75t_L g219 ( .A(n_86), .B(n_205), .Y(n_219) );
CKINVDCx20_ASAP7_75t_R g504 ( .A(n_87), .Y(n_504) );
NAND2xp5_ASAP7_75t_SL g238 ( .A(n_88), .B(n_153), .Y(n_238) );
INVx2_ASAP7_75t_L g145 ( .A(n_89), .Y(n_145) );
CKINVDCx20_ASAP7_75t_R g596 ( .A(n_90), .Y(n_596) );
NAND2xp5_ASAP7_75t_SL g538 ( .A(n_91), .B(n_195), .Y(n_538) );
NAND2xp5_ASAP7_75t_L g181 ( .A(n_92), .B(n_153), .Y(n_181) );
INVx2_ASAP7_75t_L g114 ( .A(n_93), .Y(n_114) );
OR2x2_ASAP7_75t_L g464 ( .A(n_93), .B(n_465), .Y(n_464) );
OR2x2_ASAP7_75t_L g478 ( .A(n_93), .B(n_466), .Y(n_478) );
AOI22xp33_ASAP7_75t_L g248 ( .A1(n_95), .A2(n_104), .B1(n_153), .B2(n_154), .Y(n_248) );
NAND2xp5_ASAP7_75t_L g487 ( .A(n_96), .B(n_488), .Y(n_487) );
INVx1_ASAP7_75t_L g496 ( .A(n_97), .Y(n_496) );
INVxp67_ASAP7_75t_L g567 ( .A(n_98), .Y(n_567) );
NAND2xp5_ASAP7_75t_L g190 ( .A(n_99), .B(n_153), .Y(n_190) );
NAND2xp5_ASAP7_75t_L g116 ( .A(n_100), .B(n_117), .Y(n_116) );
INVx1_ASAP7_75t_L g533 ( .A(n_101), .Y(n_533) );
INVx1_ASAP7_75t_L g591 ( .A(n_102), .Y(n_591) );
AND2x2_ASAP7_75t_L g558 ( .A(n_103), .B(n_198), .Y(n_558) );
INVx1_ASAP7_75t_L g106 ( .A(n_107), .Y(n_106) );
INVx2_ASAP7_75t_L g107 ( .A(n_108), .Y(n_107) );
INVx2_ASAP7_75t_SL g785 ( .A(n_108), .Y(n_785) );
AND2x2_ASAP7_75t_L g108 ( .A(n_109), .B(n_112), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_110), .Y(n_109) );
INVx1_ASAP7_75t_L g112 ( .A(n_113), .Y(n_112) );
OR2x2_ASAP7_75t_L g765 ( .A(n_114), .B(n_466), .Y(n_765) );
NOR2x2_ASAP7_75t_L g782 ( .A(n_114), .B(n_465), .Y(n_782) );
INVx1_ASAP7_75t_SL g115 ( .A(n_116), .Y(n_115) );
OA21x2_ASAP7_75t_L g118 ( .A1(n_119), .A2(n_124), .B(n_472), .Y(n_118) );
BUFx2_ASAP7_75t_SL g119 ( .A(n_120), .Y(n_119) );
CKINVDCx20_ASAP7_75t_R g120 ( .A(n_121), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
INVx1_ASAP7_75t_SL g784 ( .A(n_122), .Y(n_784) );
INVx2_ASAP7_75t_L g122 ( .A(n_123), .Y(n_122) );
OAI21xp5_ASAP7_75t_SL g124 ( .A1(n_125), .A2(n_461), .B(n_469), .Y(n_124) );
AOI22xp33_ASAP7_75t_L g125 ( .A1(n_126), .A2(n_129), .B1(n_130), .B2(n_460), .Y(n_125) );
CKINVDCx20_ASAP7_75t_R g460 ( .A(n_126), .Y(n_460) );
NOR2xp33_ASAP7_75t_L g515 ( .A(n_127), .B(n_516), .Y(n_515) );
INVx1_ASAP7_75t_L g129 ( .A(n_130), .Y(n_129) );
OAI22xp5_ASAP7_75t_SL g130 ( .A1(n_131), .A2(n_132), .B1(n_453), .B2(n_454), .Y(n_130) );
INVx1_ASAP7_75t_L g131 ( .A(n_132), .Y(n_131) );
AND2x2_ASAP7_75t_SL g132 ( .A(n_133), .B(n_419), .Y(n_132) );
NOR3xp33_ASAP7_75t_L g133 ( .A(n_134), .B(n_323), .C(n_407), .Y(n_133) );
NAND4xp25_ASAP7_75t_L g134 ( .A(n_135), .B(n_266), .C(n_288), .D(n_304), .Y(n_134) );
AOI221xp5_ASAP7_75t_L g135 ( .A1(n_136), .A2(n_199), .B1(n_225), .B2(n_244), .C(n_252), .Y(n_135) );
INVx1_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
NAND2xp5_ASAP7_75t_L g137 ( .A(n_138), .B(n_175), .Y(n_137) );
NAND2xp5_ASAP7_75t_SL g278 ( .A(n_138), .B(n_244), .Y(n_278) );
NAND4xp25_ASAP7_75t_L g318 ( .A(n_138), .B(n_306), .C(n_319), .D(n_321), .Y(n_318) );
INVxp67_ASAP7_75t_L g435 ( .A(n_138), .Y(n_435) );
INVx3_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
OR2x2_ASAP7_75t_L g317 ( .A(n_139), .B(n_255), .Y(n_317) );
AND2x2_ASAP7_75t_L g341 ( .A(n_139), .B(n_175), .Y(n_341) );
INVx2_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
AND2x2_ASAP7_75t_L g308 ( .A(n_140), .B(n_243), .Y(n_308) );
AND2x2_ASAP7_75t_L g348 ( .A(n_140), .B(n_329), .Y(n_348) );
AND2x2_ASAP7_75t_L g365 ( .A(n_140), .B(n_366), .Y(n_365) );
NAND2xp5_ASAP7_75t_L g389 ( .A(n_140), .B(n_176), .Y(n_389) );
INVx2_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
AND2x2_ASAP7_75t_L g242 ( .A(n_141), .B(n_243), .Y(n_242) );
AND2x2_ASAP7_75t_L g260 ( .A(n_141), .B(n_261), .Y(n_260) );
AND2x2_ASAP7_75t_L g272 ( .A(n_141), .B(n_176), .Y(n_272) );
NAND2xp5_ASAP7_75t_L g294 ( .A(n_141), .B(n_186), .Y(n_294) );
OA21x2_ASAP7_75t_L g141 ( .A1(n_142), .A2(n_149), .B(n_174), .Y(n_141) );
OA21x2_ASAP7_75t_L g186 ( .A1(n_142), .A2(n_187), .B(n_197), .Y(n_186) );
INVx2_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
NOR2xp33_ASAP7_75t_L g539 ( .A(n_143), .B(n_540), .Y(n_539) );
INVx1_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
BUFx6f_ASAP7_75t_L g177 ( .A(n_144), .Y(n_177) );
AND2x2_ASAP7_75t_L g144 ( .A(n_145), .B(n_146), .Y(n_144) );
AND2x2_ASAP7_75t_SL g198 ( .A(n_145), .B(n_146), .Y(n_198) );
NAND2xp5_ASAP7_75t_L g146 ( .A(n_147), .B(n_148), .Y(n_146) );
OAI21xp5_ASAP7_75t_L g149 ( .A1(n_150), .A2(n_163), .B(n_172), .Y(n_149) );
O2A1O1Ixp33_ASAP7_75t_L g150 ( .A1(n_151), .A2(n_152), .B(n_156), .C(n_159), .Y(n_150) );
AOI21xp5_ASAP7_75t_L g536 ( .A1(n_152), .A2(n_537), .B(n_538), .Y(n_536) );
AOI21xp5_ASAP7_75t_L g545 ( .A1(n_152), .A2(n_546), .B(n_547), .Y(n_545) );
INVx2_ASAP7_75t_L g152 ( .A(n_153), .Y(n_152) );
INVx3_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
INVx1_ASAP7_75t_L g154 ( .A(n_155), .Y(n_154) );
INVx2_ASAP7_75t_L g158 ( .A(n_155), .Y(n_158) );
INVx1_ASAP7_75t_L g166 ( .A(n_155), .Y(n_166) );
INVx3_ASAP7_75t_L g233 ( .A(n_157), .Y(n_233) );
HB1xp67_ASAP7_75t_L g593 ( .A(n_157), .Y(n_593) );
BUFx6f_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
INVx1_ASAP7_75t_L g205 ( .A(n_158), .Y(n_205) );
BUFx3_ASAP7_75t_L g206 ( .A(n_158), .Y(n_206) );
AND2x6_ASAP7_75t_L g493 ( .A(n_158), .B(n_494), .Y(n_493) );
O2A1O1Ixp33_ASAP7_75t_L g590 ( .A1(n_159), .A2(n_591), .B(n_592), .C(n_593), .Y(n_590) );
INVx1_ASAP7_75t_L g159 ( .A(n_160), .Y(n_159) );
AOI21xp5_ASAP7_75t_L g236 ( .A1(n_160), .A2(n_237), .B(n_238), .Y(n_236) );
INVx4_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
INVx2_ASAP7_75t_L g498 ( .A(n_161), .Y(n_498) );
BUFx6f_ASAP7_75t_L g161 ( .A(n_162), .Y(n_161) );
INVx3_ASAP7_75t_L g171 ( .A(n_162), .Y(n_171) );
BUFx6f_ASAP7_75t_L g195 ( .A(n_162), .Y(n_195) );
INVx1_ASAP7_75t_L g216 ( .A(n_162), .Y(n_216) );
AND2x2_ASAP7_75t_L g489 ( .A(n_162), .B(n_166), .Y(n_489) );
INVx1_ASAP7_75t_L g494 ( .A(n_162), .Y(n_494) );
O2A1O1Ixp33_ASAP7_75t_L g163 ( .A1(n_164), .A2(n_167), .B(n_168), .C(n_169), .Y(n_163) );
O2A1O1Ixp5_ASAP7_75t_L g191 ( .A1(n_164), .A2(n_192), .B(n_193), .C(n_194), .Y(n_191) );
AOI21xp5_ASAP7_75t_L g511 ( .A1(n_164), .A2(n_512), .B(n_513), .Y(n_511) );
INVx2_ASAP7_75t_L g164 ( .A(n_165), .Y(n_164) );
INVx1_ASAP7_75t_L g165 ( .A(n_166), .Y(n_165) );
AOI21xp5_ASAP7_75t_L g182 ( .A1(n_169), .A2(n_183), .B(n_184), .Y(n_182) );
OAI22xp5_ASAP7_75t_L g222 ( .A1(n_169), .A2(n_195), .B1(n_223), .B2(n_224), .Y(n_222) );
OAI22xp5_ASAP7_75t_L g247 ( .A1(n_169), .A2(n_195), .B1(n_248), .B2(n_249), .Y(n_247) );
INVx2_ASAP7_75t_L g169 ( .A(n_170), .Y(n_169) );
AOI21xp5_ASAP7_75t_L g179 ( .A1(n_170), .A2(n_180), .B(n_181), .Y(n_179) );
AOI21xp5_ASAP7_75t_L g188 ( .A1(n_170), .A2(n_189), .B(n_190), .Y(n_188) );
O2A1O1Ixp5_ASAP7_75t_SL g232 ( .A1(n_170), .A2(n_233), .B(n_234), .C(n_235), .Y(n_232) );
NOR2xp33_ASAP7_75t_L g566 ( .A(n_170), .B(n_567), .Y(n_566) );
INVx5_ASAP7_75t_L g170 ( .A(n_171), .Y(n_170) );
OAI22xp5_ASAP7_75t_SL g203 ( .A1(n_171), .A2(n_195), .B1(n_204), .B2(n_207), .Y(n_203) );
OAI21xp5_ASAP7_75t_L g178 ( .A1(n_172), .A2(n_179), .B(n_182), .Y(n_178) );
BUFx3_ASAP7_75t_L g196 ( .A(n_172), .Y(n_196) );
OAI21xp5_ASAP7_75t_L g211 ( .A1(n_172), .A2(n_212), .B(n_217), .Y(n_211) );
OAI21xp5_ASAP7_75t_L g231 ( .A1(n_172), .A2(n_232), .B(n_236), .Y(n_231) );
AND2x4_ASAP7_75t_L g488 ( .A(n_172), .B(n_489), .Y(n_488) );
INVx4_ASAP7_75t_SL g502 ( .A(n_172), .Y(n_502) );
NAND2x1p5_ASAP7_75t_L g534 ( .A(n_172), .B(n_489), .Y(n_534) );
AND2x2_ASAP7_75t_L g275 ( .A(n_175), .B(n_276), .Y(n_275) );
AOI221xp5_ASAP7_75t_L g324 ( .A1(n_175), .A2(n_325), .B1(n_328), .B2(n_330), .C(n_334), .Y(n_324) );
AND2x2_ASAP7_75t_L g383 ( .A(n_175), .B(n_348), .Y(n_383) );
NAND2xp5_ASAP7_75t_L g417 ( .A(n_175), .B(n_365), .Y(n_417) );
AND2x2_ASAP7_75t_L g175 ( .A(n_176), .B(n_186), .Y(n_175) );
INVx3_ASAP7_75t_L g243 ( .A(n_176), .Y(n_243) );
AND2x2_ASAP7_75t_L g292 ( .A(n_176), .B(n_293), .Y(n_292) );
AND2x2_ASAP7_75t_L g346 ( .A(n_176), .B(n_261), .Y(n_346) );
AND2x2_ASAP7_75t_L g404 ( .A(n_176), .B(n_405), .Y(n_404) );
OA21x2_ASAP7_75t_L g176 ( .A1(n_177), .A2(n_178), .B(n_185), .Y(n_176) );
INVx4_ASAP7_75t_L g246 ( .A(n_177), .Y(n_246) );
AOI21xp5_ASAP7_75t_L g542 ( .A1(n_177), .A2(n_543), .B(n_544), .Y(n_542) );
HB1xp67_ASAP7_75t_L g561 ( .A(n_177), .Y(n_561) );
AND2x2_ASAP7_75t_L g244 ( .A(n_186), .B(n_245), .Y(n_244) );
INVx2_ASAP7_75t_L g261 ( .A(n_186), .Y(n_261) );
INVx1_ASAP7_75t_L g316 ( .A(n_186), .Y(n_316) );
HB1xp67_ASAP7_75t_L g322 ( .A(n_186), .Y(n_322) );
AND2x2_ASAP7_75t_L g367 ( .A(n_186), .B(n_243), .Y(n_367) );
OR2x2_ASAP7_75t_L g406 ( .A(n_186), .B(n_245), .Y(n_406) );
OAI21xp5_ASAP7_75t_L g187 ( .A1(n_188), .A2(n_191), .B(n_196), .Y(n_187) );
AOI21xp5_ASAP7_75t_L g217 ( .A1(n_194), .A2(n_218), .B(n_219), .Y(n_217) );
INVx2_ASAP7_75t_L g194 ( .A(n_195), .Y(n_194) );
INVx4_ASAP7_75t_L g526 ( .A(n_195), .Y(n_526) );
NAND3xp33_ASAP7_75t_L g265 ( .A(n_196), .B(n_246), .C(n_247), .Y(n_265) );
INVx2_ASAP7_75t_L g208 ( .A(n_198), .Y(n_208) );
OA21x2_ASAP7_75t_L g210 ( .A1(n_198), .A2(n_211), .B(n_220), .Y(n_210) );
OA21x2_ASAP7_75t_L g230 ( .A1(n_198), .A2(n_231), .B(n_239), .Y(n_230) );
AOI21xp5_ASAP7_75t_L g486 ( .A1(n_198), .A2(n_487), .B(n_490), .Y(n_486) );
INVx1_ASAP7_75t_L g516 ( .A(n_198), .Y(n_516) );
AOI21xp5_ASAP7_75t_L g552 ( .A1(n_198), .A2(n_553), .B(n_554), .Y(n_552) );
NAND2xp5_ASAP7_75t_L g285 ( .A(n_199), .B(n_286), .Y(n_285) );
AND2x2_ASAP7_75t_L g199 ( .A(n_200), .B(n_209), .Y(n_199) );
AND2x2_ASAP7_75t_L g402 ( .A(n_200), .B(n_399), .Y(n_402) );
NAND2xp5_ASAP7_75t_L g434 ( .A(n_200), .B(n_384), .Y(n_434) );
BUFx2_ASAP7_75t_L g200 ( .A(n_201), .Y(n_200) );
AND2x2_ASAP7_75t_L g333 ( .A(n_201), .B(n_257), .Y(n_333) );
AND2x2_ASAP7_75t_L g382 ( .A(n_201), .B(n_228), .Y(n_382) );
INVx1_ASAP7_75t_L g428 ( .A(n_201), .Y(n_428) );
INVx1_ASAP7_75t_L g201 ( .A(n_202), .Y(n_201) );
BUFx6f_ASAP7_75t_L g241 ( .A(n_202), .Y(n_241) );
AND2x2_ASAP7_75t_L g283 ( .A(n_202), .B(n_257), .Y(n_283) );
INVx1_ASAP7_75t_L g300 ( .A(n_202), .Y(n_300) );
AND2x2_ASAP7_75t_L g306 ( .A(n_202), .B(n_221), .Y(n_306) );
HB1xp67_ASAP7_75t_L g500 ( .A(n_206), .Y(n_500) );
INVx2_ASAP7_75t_L g527 ( .A(n_206), .Y(n_527) );
INVx1_ASAP7_75t_L g514 ( .A(n_208), .Y(n_514) );
AND2x2_ASAP7_75t_L g374 ( .A(n_209), .B(n_282), .Y(n_374) );
INVx2_ASAP7_75t_L g439 ( .A(n_209), .Y(n_439) );
AND2x2_ASAP7_75t_L g209 ( .A(n_210), .B(n_221), .Y(n_209) );
AND2x2_ASAP7_75t_L g256 ( .A(n_210), .B(n_257), .Y(n_256) );
OR2x2_ASAP7_75t_L g269 ( .A(n_210), .B(n_229), .Y(n_269) );
NAND2xp5_ASAP7_75t_L g297 ( .A(n_210), .B(n_228), .Y(n_297) );
INVx1_ASAP7_75t_L g303 ( .A(n_210), .Y(n_303) );
INVx1_ASAP7_75t_L g320 ( .A(n_210), .Y(n_320) );
HB1xp67_ASAP7_75t_L g332 ( .A(n_210), .Y(n_332) );
INVx2_ASAP7_75t_L g400 ( .A(n_210), .Y(n_400) );
AOI21xp5_ASAP7_75t_L g212 ( .A1(n_213), .A2(n_214), .B(n_215), .Y(n_212) );
INVx1_ASAP7_75t_L g215 ( .A(n_216), .Y(n_215) );
INVx2_ASAP7_75t_L g257 ( .A(n_221), .Y(n_257) );
BUFx2_ASAP7_75t_L g354 ( .A(n_221), .Y(n_354) );
AND2x2_ASAP7_75t_L g399 ( .A(n_221), .B(n_400), .Y(n_399) );
INVx1_ASAP7_75t_L g225 ( .A(n_226), .Y(n_225) );
NAND2xp5_ASAP7_75t_L g226 ( .A(n_227), .B(n_240), .Y(n_226) );
NAND2xp5_ASAP7_75t_L g335 ( .A(n_227), .B(n_336), .Y(n_335) );
AOI21xp5_ASAP7_75t_L g422 ( .A1(n_227), .A2(n_398), .B(n_412), .Y(n_422) );
AND2x2_ASAP7_75t_L g447 ( .A(n_227), .B(n_333), .Y(n_447) );
BUFx2_ASAP7_75t_L g227 ( .A(n_228), .Y(n_227) );
INVx2_ASAP7_75t_L g228 ( .A(n_229), .Y(n_228) );
INVx1_ASAP7_75t_L g369 ( .A(n_229), .Y(n_369) );
AND2x2_ASAP7_75t_L g398 ( .A(n_229), .B(n_399), .Y(n_398) );
INVx2_ASAP7_75t_L g229 ( .A(n_230), .Y(n_229) );
HB1xp67_ASAP7_75t_L g282 ( .A(n_230), .Y(n_282) );
INVx2_ASAP7_75t_L g301 ( .A(n_230), .Y(n_301) );
OR2x2_ASAP7_75t_L g302 ( .A(n_230), .B(n_303), .Y(n_302) );
AND2x2_ASAP7_75t_L g240 ( .A(n_241), .B(n_242), .Y(n_240) );
INVx2_ASAP7_75t_L g255 ( .A(n_241), .Y(n_255) );
OR2x2_ASAP7_75t_L g268 ( .A(n_241), .B(n_269), .Y(n_268) );
AND2x2_ASAP7_75t_L g336 ( .A(n_241), .B(n_332), .Y(n_336) );
NAND2xp5_ASAP7_75t_L g431 ( .A(n_241), .B(n_432), .Y(n_431) );
OR2x2_ASAP7_75t_L g437 ( .A(n_241), .B(n_438), .Y(n_437) );
NAND2xp5_ASAP7_75t_L g449 ( .A(n_241), .B(n_374), .Y(n_449) );
AND2x2_ASAP7_75t_L g328 ( .A(n_242), .B(n_329), .Y(n_328) );
AND2x2_ASAP7_75t_L g351 ( .A(n_242), .B(n_244), .Y(n_351) );
INVx2_ASAP7_75t_L g263 ( .A(n_243), .Y(n_263) );
AND2x2_ASAP7_75t_L g291 ( .A(n_243), .B(n_264), .Y(n_291) );
NAND2xp5_ASAP7_75t_L g372 ( .A(n_243), .B(n_316), .Y(n_372) );
AND2x2_ASAP7_75t_L g286 ( .A(n_244), .B(n_287), .Y(n_286) );
INVx1_ASAP7_75t_L g433 ( .A(n_244), .Y(n_433) );
AND2x2_ASAP7_75t_L g445 ( .A(n_244), .B(n_308), .Y(n_445) );
AND2x2_ASAP7_75t_L g271 ( .A(n_245), .B(n_261), .Y(n_271) );
INVx1_ASAP7_75t_L g366 ( .A(n_245), .Y(n_366) );
AO21x1_ASAP7_75t_L g245 ( .A1(n_246), .A2(n_247), .B(n_250), .Y(n_245) );
NOR2xp33_ASAP7_75t_L g503 ( .A(n_246), .B(n_504), .Y(n_503) );
INVx3_ASAP7_75t_L g519 ( .A(n_246), .Y(n_519) );
AO21x2_ASAP7_75t_L g531 ( .A1(n_246), .A2(n_532), .B(n_539), .Y(n_531) );
AO21x2_ASAP7_75t_L g587 ( .A1(n_246), .A2(n_588), .B(n_595), .Y(n_587) );
NOR2xp33_ASAP7_75t_L g595 ( .A(n_246), .B(n_596), .Y(n_595) );
INVx1_ASAP7_75t_L g250 ( .A(n_251), .Y(n_250) );
AND2x4_ASAP7_75t_L g264 ( .A(n_251), .B(n_265), .Y(n_264) );
INVxp67_ASAP7_75t_L g252 ( .A(n_253), .Y(n_252) );
NAND2xp5_ASAP7_75t_L g253 ( .A(n_254), .B(n_258), .Y(n_253) );
AND2x2_ASAP7_75t_L g254 ( .A(n_255), .B(n_256), .Y(n_254) );
NOR2xp33_ASAP7_75t_L g311 ( .A(n_255), .B(n_302), .Y(n_311) );
OR2x2_ASAP7_75t_L g443 ( .A(n_255), .B(n_444), .Y(n_443) );
AND2x2_ASAP7_75t_L g360 ( .A(n_256), .B(n_301), .Y(n_360) );
AND2x2_ASAP7_75t_L g368 ( .A(n_256), .B(n_369), .Y(n_368) );
AND2x2_ASAP7_75t_L g427 ( .A(n_256), .B(n_428), .Y(n_427) );
AND2x2_ASAP7_75t_L g451 ( .A(n_256), .B(n_298), .Y(n_451) );
NOR2xp67_ASAP7_75t_L g409 ( .A(n_257), .B(n_410), .Y(n_409) );
OR2x2_ASAP7_75t_L g438 ( .A(n_257), .B(n_301), .Y(n_438) );
INVx1_ASAP7_75t_L g258 ( .A(n_259), .Y(n_258) );
NAND2x1p5_ASAP7_75t_L g259 ( .A(n_260), .B(n_262), .Y(n_259) );
AND2x2_ASAP7_75t_L g290 ( .A(n_260), .B(n_291), .Y(n_290) );
INVxp67_ASAP7_75t_L g452 ( .A(n_260), .Y(n_452) );
NOR2x1_ASAP7_75t_L g262 ( .A(n_263), .B(n_264), .Y(n_262) );
INVx1_ASAP7_75t_L g287 ( .A(n_263), .Y(n_287) );
AND2x2_ASAP7_75t_L g338 ( .A(n_263), .B(n_271), .Y(n_338) );
NOR2xp33_ASAP7_75t_L g432 ( .A(n_263), .B(n_406), .Y(n_432) );
INVx2_ASAP7_75t_L g277 ( .A(n_264), .Y(n_277) );
INVx3_ASAP7_75t_L g329 ( .A(n_264), .Y(n_329) );
OR2x2_ASAP7_75t_L g357 ( .A(n_264), .B(n_358), .Y(n_357) );
AOI311xp33_ASAP7_75t_L g266 ( .A1(n_267), .A2(n_270), .A3(n_272), .B(n_273), .C(n_284), .Y(n_266) );
O2A1O1Ixp33_ASAP7_75t_L g304 ( .A1(n_267), .A2(n_305), .B(n_307), .C(n_309), .Y(n_304) );
INVx2_ASAP7_75t_L g267 ( .A(n_268), .Y(n_267) );
INVx2_ASAP7_75t_SL g289 ( .A(n_269), .Y(n_289) );
INVx2_ASAP7_75t_L g270 ( .A(n_271), .Y(n_270) );
AND2x2_ASAP7_75t_L g307 ( .A(n_271), .B(n_308), .Y(n_307) );
NAND2xp5_ASAP7_75t_L g392 ( .A(n_271), .B(n_287), .Y(n_392) );
NAND2xp5_ASAP7_75t_L g440 ( .A(n_271), .B(n_272), .Y(n_440) );
AND2x2_ASAP7_75t_L g362 ( .A(n_272), .B(n_276), .Y(n_362) );
AOI21xp33_ASAP7_75t_L g273 ( .A1(n_274), .A2(n_278), .B(n_279), .Y(n_273) );
INVx1_ASAP7_75t_L g274 ( .A(n_275), .Y(n_274) );
AND2x2_ASAP7_75t_L g420 ( .A(n_276), .B(n_308), .Y(n_420) );
INVx2_ASAP7_75t_L g276 ( .A(n_277), .Y(n_276) );
NOR2xp33_ASAP7_75t_L g293 ( .A(n_277), .B(n_294), .Y(n_293) );
INVx1_ASAP7_75t_L g314 ( .A(n_277), .Y(n_314) );
INVx1_ASAP7_75t_L g279 ( .A(n_280), .Y(n_279) );
AND2x2_ASAP7_75t_L g280 ( .A(n_281), .B(n_283), .Y(n_280) );
AND2x2_ASAP7_75t_L g305 ( .A(n_281), .B(n_306), .Y(n_305) );
INVx1_ASAP7_75t_L g281 ( .A(n_282), .Y(n_281) );
INVx1_ASAP7_75t_L g350 ( .A(n_283), .Y(n_350) );
AND2x4_ASAP7_75t_L g412 ( .A(n_283), .B(n_381), .Y(n_412) );
INVx1_ASAP7_75t_L g284 ( .A(n_285), .Y(n_284) );
AOI222xp33_ASAP7_75t_L g363 ( .A1(n_286), .A2(n_352), .B1(n_364), .B2(n_368), .C1(n_370), .C2(n_374), .Y(n_363) );
A2O1A1Ixp33_ASAP7_75t_L g288 ( .A1(n_289), .A2(n_290), .B(n_292), .C(n_295), .Y(n_288) );
NAND2xp5_ASAP7_75t_L g356 ( .A(n_289), .B(n_333), .Y(n_356) );
INVx1_ASAP7_75t_L g378 ( .A(n_291), .Y(n_378) );
INVx1_ASAP7_75t_L g312 ( .A(n_293), .Y(n_312) );
OR2x2_ASAP7_75t_L g377 ( .A(n_294), .B(n_378), .Y(n_377) );
OAI21xp33_ASAP7_75t_SL g295 ( .A1(n_296), .A2(n_298), .B(n_302), .Y(n_295) );
NAND3xp33_ASAP7_75t_L g313 ( .A(n_296), .B(n_314), .C(n_315), .Y(n_313) );
AOI21xp5_ASAP7_75t_L g411 ( .A1(n_296), .A2(n_333), .B(n_412), .Y(n_411) );
INVx1_ASAP7_75t_L g296 ( .A(n_297), .Y(n_296) );
INVx1_ASAP7_75t_SL g298 ( .A(n_299), .Y(n_298) );
NAND2xp5_ASAP7_75t_L g299 ( .A(n_300), .B(n_301), .Y(n_299) );
HB1xp67_ASAP7_75t_L g353 ( .A(n_300), .Y(n_353) );
AND2x2_ASAP7_75t_SL g319 ( .A(n_301), .B(n_320), .Y(n_319) );
INVx1_ASAP7_75t_L g410 ( .A(n_301), .Y(n_410) );
HB1xp67_ASAP7_75t_L g426 ( .A(n_301), .Y(n_426) );
INVx2_ASAP7_75t_L g384 ( .A(n_302), .Y(n_384) );
NAND2xp5_ASAP7_75t_L g326 ( .A(n_306), .B(n_327), .Y(n_326) );
INVx2_ASAP7_75t_L g358 ( .A(n_308), .Y(n_358) );
OAI221xp5_ASAP7_75t_L g309 ( .A1(n_310), .A2(n_312), .B1(n_313), .B2(n_317), .C(n_318), .Y(n_309) );
INVx1_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
NAND2xp5_ASAP7_75t_SL g391 ( .A(n_312), .B(n_392), .Y(n_391) );
INVx1_ASAP7_75t_SL g446 ( .A(n_312), .Y(n_446) );
INVx1_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
INVx2_ASAP7_75t_L g327 ( .A(n_319), .Y(n_327) );
NOR2xp33_ASAP7_75t_L g349 ( .A(n_319), .B(n_350), .Y(n_349) );
AND2x2_ASAP7_75t_L g385 ( .A(n_319), .B(n_333), .Y(n_385) );
NAND2xp5_ASAP7_75t_L g394 ( .A(n_319), .B(n_395), .Y(n_394) );
AND2x2_ASAP7_75t_L g418 ( .A(n_319), .B(n_353), .Y(n_418) );
BUFx3_ASAP7_75t_L g381 ( .A(n_320), .Y(n_381) );
INVx1_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
NAND5xp2_ASAP7_75t_L g323 ( .A(n_324), .B(n_342), .C(n_363), .D(n_375), .E(n_390), .Y(n_323) );
INVx1_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
AOI32xp33_ASAP7_75t_L g415 ( .A1(n_327), .A2(n_354), .A3(n_370), .B1(n_416), .B2(n_418), .Y(n_415) );
NAND2xp5_ASAP7_75t_L g387 ( .A(n_329), .B(n_388), .Y(n_387) );
AND2x2_ASAP7_75t_L g330 ( .A(n_331), .B(n_333), .Y(n_330) );
INVx1_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
INVx1_ASAP7_75t_SL g339 ( .A(n_333), .Y(n_339) );
OAI22xp5_ASAP7_75t_L g334 ( .A1(n_335), .A2(n_337), .B1(n_339), .B2(n_340), .Y(n_334) );
INVx1_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
INVx1_ASAP7_75t_SL g340 ( .A(n_341), .Y(n_340) );
AOI221xp5_ASAP7_75t_L g342 ( .A1(n_343), .A2(n_349), .B1(n_351), .B2(n_352), .C(n_355), .Y(n_342) );
INVx2_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
OR2x2_ASAP7_75t_L g344 ( .A(n_345), .B(n_347), .Y(n_344) );
INVx1_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
AND2x2_ASAP7_75t_L g414 ( .A(n_346), .B(n_365), .Y(n_414) );
INVx1_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
AOI221xp5_ASAP7_75t_L g429 ( .A1(n_351), .A2(n_412), .B1(n_430), .B2(n_435), .C(n_436), .Y(n_429) );
AND2x2_ASAP7_75t_L g352 ( .A(n_353), .B(n_354), .Y(n_352) );
INVx2_ASAP7_75t_L g395 ( .A(n_354), .Y(n_395) );
OAI22xp5_ASAP7_75t_L g355 ( .A1(n_356), .A2(n_357), .B1(n_359), .B2(n_361), .Y(n_355) );
INVx1_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
INVx1_ASAP7_75t_SL g361 ( .A(n_362), .Y(n_361) );
AND2x2_ASAP7_75t_L g364 ( .A(n_365), .B(n_367), .Y(n_364) );
INVx1_ASAP7_75t_L g373 ( .A(n_365), .Y(n_373) );
INVx1_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
OR2x2_ASAP7_75t_L g371 ( .A(n_372), .B(n_373), .Y(n_371) );
AOI222xp33_ASAP7_75t_L g375 ( .A1(n_376), .A2(n_379), .B1(n_383), .B2(n_384), .C1(n_385), .C2(n_386), .Y(n_375) );
INVx1_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
AND2x2_ASAP7_75t_L g379 ( .A(n_380), .B(n_382), .Y(n_379) );
INVxp67_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
OAI22xp33_ASAP7_75t_L g430 ( .A1(n_384), .A2(n_431), .B1(n_433), .B2(n_434), .Y(n_430) );
INVx1_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
INVx1_ASAP7_75t_SL g388 ( .A(n_389), .Y(n_388) );
AOI21xp5_ASAP7_75t_L g390 ( .A1(n_391), .A2(n_393), .B(n_396), .Y(n_390) );
INVx1_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
AOI21xp33_ASAP7_75t_L g396 ( .A1(n_397), .A2(n_401), .B(n_403), .Y(n_396) );
INVx2_ASAP7_75t_SL g397 ( .A(n_398), .Y(n_397) );
INVx1_ASAP7_75t_L g444 ( .A(n_399), .Y(n_444) );
INVx1_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
INVx1_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
INVx1_ASAP7_75t_SL g405 ( .A(n_406), .Y(n_405) );
A2O1A1Ixp33_ASAP7_75t_L g407 ( .A1(n_408), .A2(n_411), .B(n_413), .C(n_415), .Y(n_407) );
INVx1_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
INVx1_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
INVx1_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
AOI211xp5_ASAP7_75t_L g419 ( .A1(n_420), .A2(n_421), .B(n_423), .C(n_448), .Y(n_419) );
CKINVDCx16_ASAP7_75t_R g424 ( .A(n_420), .Y(n_424) );
INVxp67_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
OAI211xp5_ASAP7_75t_L g423 ( .A1(n_424), .A2(n_425), .B(n_429), .C(n_441), .Y(n_423) );
NAND2xp5_ASAP7_75t_L g425 ( .A(n_426), .B(n_427), .Y(n_425) );
AOI21xp33_ASAP7_75t_L g436 ( .A1(n_437), .A2(n_439), .B(n_440), .Y(n_436) );
AOI22xp5_ASAP7_75t_L g441 ( .A1(n_442), .A2(n_445), .B1(n_446), .B2(n_447), .Y(n_441) );
INVx1_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
AOI21xp33_ASAP7_75t_L g448 ( .A1(n_449), .A2(n_450), .B(n_452), .Y(n_448) );
INVx1_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
INVx1_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
CKINVDCx20_ASAP7_75t_R g459 ( .A(n_455), .Y(n_459) );
INVx1_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
INVx1_ASAP7_75t_SL g462 ( .A(n_463), .Y(n_462) );
INVx1_ASAP7_75t_SL g463 ( .A(n_464), .Y(n_463) );
HB1xp67_ASAP7_75t_L g471 ( .A(n_464), .Y(n_471) );
INVx2_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
AND2x2_ASAP7_75t_L g466 ( .A(n_467), .B(n_468), .Y(n_466) );
NAND3xp33_ASAP7_75t_L g472 ( .A(n_469), .B(n_473), .C(n_783), .Y(n_472) );
INVx1_ASAP7_75t_L g470 ( .A(n_471), .Y(n_470) );
OAI22xp5_ASAP7_75t_SL g474 ( .A1(n_475), .A2(n_476), .B1(n_479), .B2(n_765), .Y(n_474) );
INVx1_ASAP7_75t_L g777 ( .A(n_475), .Y(n_777) );
OAI22x1_ASAP7_75t_SL g776 ( .A1(n_476), .A2(n_480), .B1(n_777), .B2(n_778), .Y(n_776) );
INVx2_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
INVx1_ASAP7_75t_L g477 ( .A(n_478), .Y(n_477) );
INVx2_ASAP7_75t_L g479 ( .A(n_480), .Y(n_479) );
OR3x2_ASAP7_75t_L g480 ( .A(n_481), .B(n_679), .C(n_722), .Y(n_480) );
NAND5xp2_ASAP7_75t_L g481 ( .A(n_482), .B(n_606), .C(n_636), .D(n_653), .E(n_668), .Y(n_481) );
AOI221xp5_ASAP7_75t_SL g482 ( .A1(n_483), .A2(n_529), .B1(n_569), .B2(n_575), .C(n_579), .Y(n_482) );
AND2x2_ASAP7_75t_L g483 ( .A(n_484), .B(n_505), .Y(n_483) );
OR2x2_ASAP7_75t_L g584 ( .A(n_484), .B(n_585), .Y(n_584) );
AND2x2_ASAP7_75t_L g623 ( .A(n_484), .B(n_624), .Y(n_623) );
AND2x2_ASAP7_75t_L g641 ( .A(n_484), .B(n_642), .Y(n_641) );
NAND2xp5_ASAP7_75t_L g658 ( .A(n_484), .B(n_577), .Y(n_658) );
OR2x2_ASAP7_75t_L g670 ( .A(n_484), .B(n_671), .Y(n_670) );
NAND2xp5_ASAP7_75t_L g684 ( .A(n_484), .B(n_629), .Y(n_684) );
NAND2xp5_ASAP7_75t_L g702 ( .A(n_484), .B(n_703), .Y(n_702) );
NAND2xp5_ASAP7_75t_L g712 ( .A(n_484), .B(n_607), .Y(n_712) );
NAND2xp5_ASAP7_75t_L g721 ( .A(n_484), .B(n_615), .Y(n_721) );
AND2x2_ASAP7_75t_L g753 ( .A(n_484), .B(n_517), .Y(n_753) );
HB1xp67_ASAP7_75t_L g761 ( .A(n_484), .Y(n_761) );
INVx5_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
NAND2xp5_ASAP7_75t_L g576 ( .A(n_485), .B(n_577), .Y(n_576) );
AND2x2_ASAP7_75t_L g581 ( .A(n_485), .B(n_559), .Y(n_581) );
BUFx2_ASAP7_75t_L g603 ( .A(n_485), .Y(n_603) );
AND2x2_ASAP7_75t_L g632 ( .A(n_485), .B(n_506), .Y(n_632) );
AND2x2_ASAP7_75t_L g687 ( .A(n_485), .B(n_585), .Y(n_687) );
OR2x6_ASAP7_75t_L g485 ( .A(n_486), .B(n_503), .Y(n_485) );
BUFx2_ASAP7_75t_L g509 ( .A(n_488), .Y(n_509) );
INVx2_ASAP7_75t_L g491 ( .A(n_492), .Y(n_491) );
O2A1O1Ixp33_ASAP7_75t_SL g521 ( .A1(n_492), .A2(n_502), .B(n_522), .C(n_523), .Y(n_521) );
O2A1O1Ixp33_ASAP7_75t_L g563 ( .A1(n_492), .A2(n_502), .B(n_564), .C(n_565), .Y(n_563) );
INVx5_ASAP7_75t_L g492 ( .A(n_493), .Y(n_492) );
O2A1O1Ixp33_ASAP7_75t_L g495 ( .A1(n_496), .A2(n_497), .B(n_499), .C(n_500), .Y(n_495) );
O2A1O1Ixp33_ASAP7_75t_L g555 ( .A1(n_497), .A2(n_500), .B(n_556), .C(n_557), .Y(n_555) );
INVx2_ASAP7_75t_L g497 ( .A(n_498), .Y(n_497) );
INVx1_ASAP7_75t_L g501 ( .A(n_502), .Y(n_501) );
NAND2xp5_ASAP7_75t_L g650 ( .A(n_505), .B(n_641), .Y(n_650) );
OAI32xp33_ASAP7_75t_L g664 ( .A1(n_505), .A2(n_600), .A3(n_665), .B1(n_666), .B2(n_667), .Y(n_664) );
NAND2xp5_ASAP7_75t_L g696 ( .A(n_505), .B(n_666), .Y(n_696) );
NOR2xp33_ASAP7_75t_L g707 ( .A(n_505), .B(n_584), .Y(n_707) );
INVx1_ASAP7_75t_SL g736 ( .A(n_505), .Y(n_736) );
NAND4xp25_ASAP7_75t_L g745 ( .A(n_505), .B(n_531), .C(n_687), .D(n_746), .Y(n_745) );
AND2x4_ASAP7_75t_L g505 ( .A(n_506), .B(n_517), .Y(n_505) );
INVx5_ASAP7_75t_L g578 ( .A(n_506), .Y(n_578) );
AND2x2_ASAP7_75t_L g607 ( .A(n_506), .B(n_518), .Y(n_607) );
HB1xp67_ASAP7_75t_L g686 ( .A(n_506), .Y(n_686) );
AND2x2_ASAP7_75t_L g756 ( .A(n_506), .B(n_703), .Y(n_756) );
OR2x6_ASAP7_75t_L g506 ( .A(n_507), .B(n_515), .Y(n_506) );
AOI21xp5_ASAP7_75t_SL g507 ( .A1(n_508), .A2(n_510), .B(n_514), .Y(n_507) );
AND2x4_ASAP7_75t_L g629 ( .A(n_517), .B(n_578), .Y(n_629) );
NAND2xp5_ASAP7_75t_L g638 ( .A(n_517), .B(n_639), .Y(n_638) );
AND2x2_ASAP7_75t_L g663 ( .A(n_517), .B(n_585), .Y(n_663) );
INVx2_ASAP7_75t_L g517 ( .A(n_518), .Y(n_517) );
AND2x2_ASAP7_75t_L g577 ( .A(n_518), .B(n_578), .Y(n_577) );
AND2x2_ASAP7_75t_L g615 ( .A(n_518), .B(n_587), .Y(n_615) );
AND2x2_ASAP7_75t_L g624 ( .A(n_518), .B(n_586), .Y(n_624) );
OA21x2_ASAP7_75t_L g518 ( .A1(n_519), .A2(n_520), .B(n_528), .Y(n_518) );
NOR2xp33_ASAP7_75t_L g524 ( .A(n_525), .B(n_526), .Y(n_524) );
AOI222xp33_ASAP7_75t_L g692 ( .A1(n_529), .A2(n_693), .B1(n_695), .B2(n_697), .C1(n_700), .C2(n_701), .Y(n_692) );
AND2x4_ASAP7_75t_L g529 ( .A(n_530), .B(n_548), .Y(n_529) );
AND2x2_ASAP7_75t_L g625 ( .A(n_530), .B(n_626), .Y(n_625) );
NAND3xp33_ASAP7_75t_L g742 ( .A(n_530), .B(n_603), .C(n_743), .Y(n_742) );
AND2x2_ASAP7_75t_L g530 ( .A(n_531), .B(n_541), .Y(n_530) );
INVx5_ASAP7_75t_SL g574 ( .A(n_531), .Y(n_574) );
OAI322xp33_ASAP7_75t_L g579 ( .A1(n_531), .A2(n_580), .A3(n_582), .B1(n_583), .B2(n_597), .C1(n_600), .C2(n_602), .Y(n_579) );
NAND2xp5_ASAP7_75t_SL g645 ( .A(n_531), .B(n_572), .Y(n_645) );
NAND2xp5_ASAP7_75t_L g751 ( .A(n_531), .B(n_560), .Y(n_751) );
OAI21xp5_ASAP7_75t_L g532 ( .A1(n_533), .A2(n_534), .B(n_535), .Y(n_532) );
INVx2_ASAP7_75t_L g572 ( .A(n_541), .Y(n_572) );
NAND2xp5_ASAP7_75t_L g656 ( .A(n_541), .B(n_550), .Y(n_656) );
NAND2xp5_ASAP7_75t_L g665 ( .A(n_548), .B(n_610), .Y(n_665) );
INVx2_ASAP7_75t_L g548 ( .A(n_549), .Y(n_548) );
OR2x2_ASAP7_75t_L g644 ( .A(n_549), .B(n_645), .Y(n_644) );
NAND2xp5_ASAP7_75t_L g549 ( .A(n_550), .B(n_559), .Y(n_549) );
OR2x2_ASAP7_75t_L g573 ( .A(n_550), .B(n_574), .Y(n_573) );
NAND2xp5_ASAP7_75t_L g580 ( .A(n_550), .B(n_581), .Y(n_580) );
OR2x2_ASAP7_75t_L g612 ( .A(n_550), .B(n_560), .Y(n_612) );
AND2x2_ASAP7_75t_L g635 ( .A(n_550), .B(n_572), .Y(n_635) );
NOR2xp33_ASAP7_75t_L g646 ( .A(n_550), .B(n_647), .Y(n_646) );
AND2x2_ASAP7_75t_L g651 ( .A(n_550), .B(n_610), .Y(n_651) );
AND2x2_ASAP7_75t_L g659 ( .A(n_550), .B(n_660), .Y(n_659) );
NAND2xp5_ASAP7_75t_L g709 ( .A(n_550), .B(n_619), .Y(n_709) );
INVx5_ASAP7_75t_SL g550 ( .A(n_551), .Y(n_550) );
AND2x2_ASAP7_75t_L g599 ( .A(n_551), .B(n_574), .Y(n_599) );
OR2x2_ASAP7_75t_L g600 ( .A(n_551), .B(n_601), .Y(n_600) );
AND2x2_ASAP7_75t_L g626 ( .A(n_551), .B(n_560), .Y(n_626) );
NAND2xp5_ASAP7_75t_L g714 ( .A(n_551), .B(n_673), .Y(n_714) );
OR2x2_ASAP7_75t_L g730 ( .A(n_551), .B(n_674), .Y(n_730) );
AND2x2_ASAP7_75t_SL g737 ( .A(n_551), .B(n_691), .Y(n_737) );
HB1xp67_ASAP7_75t_L g744 ( .A(n_551), .Y(n_744) );
OR2x6_ASAP7_75t_L g551 ( .A(n_552), .B(n_558), .Y(n_551) );
AND2x2_ASAP7_75t_L g598 ( .A(n_559), .B(n_599), .Y(n_598) );
AND2x2_ASAP7_75t_L g648 ( .A(n_559), .B(n_572), .Y(n_648) );
NAND2xp5_ASAP7_75t_L g699 ( .A(n_559), .B(n_574), .Y(n_699) );
NAND2xp5_ASAP7_75t_L g732 ( .A(n_559), .B(n_610), .Y(n_732) );
INVx3_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
NAND2xp5_ASAP7_75t_L g601 ( .A(n_560), .B(n_574), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g620 ( .A(n_560), .B(n_572), .Y(n_620) );
OR2x2_ASAP7_75t_L g674 ( .A(n_560), .B(n_572), .Y(n_674) );
AND2x2_ASAP7_75t_L g691 ( .A(n_560), .B(n_571), .Y(n_691) );
INVxp67_ASAP7_75t_L g713 ( .A(n_560), .Y(n_713) );
AND2x2_ASAP7_75t_L g740 ( .A(n_560), .B(n_610), .Y(n_740) );
HB1xp67_ASAP7_75t_L g747 ( .A(n_560), .Y(n_747) );
OA21x2_ASAP7_75t_L g560 ( .A1(n_561), .A2(n_562), .B(n_568), .Y(n_560) );
INVx1_ASAP7_75t_L g569 ( .A(n_570), .Y(n_569) );
OR2x2_ASAP7_75t_L g570 ( .A(n_571), .B(n_573), .Y(n_570) );
NAND2xp5_ASAP7_75t_L g694 ( .A(n_571), .B(n_621), .Y(n_694) );
INVx1_ASAP7_75t_SL g571 ( .A(n_572), .Y(n_571) );
AND2x2_ASAP7_75t_L g610 ( .A(n_572), .B(n_574), .Y(n_610) );
OR2x2_ASAP7_75t_L g677 ( .A(n_572), .B(n_678), .Y(n_677) );
INVx2_ASAP7_75t_L g621 ( .A(n_573), .Y(n_621) );
OR2x2_ASAP7_75t_L g682 ( .A(n_573), .B(n_674), .Y(n_682) );
INVx1_ASAP7_75t_L g575 ( .A(n_576), .Y(n_575) );
INVx1_ASAP7_75t_L g582 ( .A(n_577), .Y(n_582) );
NAND2xp5_ASAP7_75t_L g640 ( .A(n_577), .B(n_641), .Y(n_640) );
OR2x2_ASAP7_75t_L g583 ( .A(n_578), .B(n_584), .Y(n_583) );
NAND2xp5_ASAP7_75t_L g604 ( .A(n_578), .B(n_605), .Y(n_604) );
NAND2xp5_ASAP7_75t_L g617 ( .A(n_578), .B(n_585), .Y(n_617) );
INVx2_ASAP7_75t_L g662 ( .A(n_578), .Y(n_662) );
AND2x2_ASAP7_75t_L g675 ( .A(n_578), .B(n_615), .Y(n_675) );
AND2x2_ASAP7_75t_L g700 ( .A(n_578), .B(n_624), .Y(n_700) );
INVx1_ASAP7_75t_L g652 ( .A(n_583), .Y(n_652) );
INVx2_ASAP7_75t_SL g639 ( .A(n_584), .Y(n_639) );
INVx1_ASAP7_75t_L g642 ( .A(n_585), .Y(n_642) );
INVx2_ASAP7_75t_L g585 ( .A(n_586), .Y(n_585) );
HB1xp67_ASAP7_75t_L g605 ( .A(n_586), .Y(n_605) );
INVx2_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
BUFx2_ASAP7_75t_L g703 ( .A(n_587), .Y(n_703) );
NAND2xp5_ASAP7_75t_L g588 ( .A(n_589), .B(n_594), .Y(n_588) );
INVx1_ASAP7_75t_L g597 ( .A(n_598), .Y(n_597) );
AND2x2_ASAP7_75t_L g672 ( .A(n_599), .B(n_673), .Y(n_672) );
INVx1_ASAP7_75t_L g678 ( .A(n_599), .Y(n_678) );
AOI22xp5_ASAP7_75t_L g680 ( .A1(n_599), .A2(n_681), .B1(n_683), .B2(n_688), .Y(n_680) );
NAND2xp5_ASAP7_75t_L g718 ( .A(n_599), .B(n_691), .Y(n_718) );
NAND2xp5_ASAP7_75t_L g693 ( .A(n_600), .B(n_694), .Y(n_693) );
INVx1_ASAP7_75t_SL g634 ( .A(n_601), .Y(n_634) );
OR2x2_ASAP7_75t_L g602 ( .A(n_603), .B(n_604), .Y(n_602) );
OR2x2_ASAP7_75t_L g616 ( .A(n_603), .B(n_617), .Y(n_616) );
NAND2xp5_ASAP7_75t_L g667 ( .A(n_603), .B(n_607), .Y(n_667) );
AND2x2_ASAP7_75t_L g690 ( .A(n_603), .B(n_691), .Y(n_690) );
BUFx2_ASAP7_75t_L g666 ( .A(n_605), .Y(n_666) );
AOI211xp5_ASAP7_75t_L g606 ( .A1(n_607), .A2(n_608), .B(n_613), .C(n_627), .Y(n_606) );
INVx1_ASAP7_75t_L g630 ( .A(n_607), .Y(n_630) );
OAI221xp5_ASAP7_75t_SL g738 ( .A1(n_607), .A2(n_739), .B1(n_741), .B2(n_742), .C(n_745), .Y(n_738) );
INVx1_ASAP7_75t_L g608 ( .A(n_609), .Y(n_608) );
NAND2xp5_ASAP7_75t_L g609 ( .A(n_610), .B(n_611), .Y(n_609) );
INVx1_ASAP7_75t_L g757 ( .A(n_610), .Y(n_757) );
INVx1_ASAP7_75t_L g611 ( .A(n_612), .Y(n_611) );
OR2x2_ASAP7_75t_L g706 ( .A(n_612), .B(n_645), .Y(n_706) );
A2O1A1Ixp33_ASAP7_75t_L g613 ( .A1(n_614), .A2(n_616), .B(n_618), .C(n_622), .Y(n_613) );
INVx1_ASAP7_75t_L g614 ( .A(n_615), .Y(n_614) );
NAND2xp5_ASAP7_75t_L g618 ( .A(n_619), .B(n_621), .Y(n_618) );
INVx1_ASAP7_75t_SL g619 ( .A(n_620), .Y(n_619) );
OAI32xp33_ASAP7_75t_L g731 ( .A1(n_620), .A2(n_621), .A3(n_684), .B1(n_721), .B2(n_732), .Y(n_731) );
NAND2xp5_ASAP7_75t_L g622 ( .A(n_623), .B(n_625), .Y(n_622) );
AND2x2_ASAP7_75t_L g763 ( .A(n_623), .B(n_662), .Y(n_763) );
AND2x2_ASAP7_75t_L g710 ( .A(n_624), .B(n_662), .Y(n_710) );
NAND2xp5_ASAP7_75t_L g728 ( .A(n_624), .B(n_632), .Y(n_728) );
AOI31xp33_ASAP7_75t_SL g627 ( .A1(n_628), .A2(n_630), .A3(n_631), .B(n_633), .Y(n_627) );
INVxp67_ASAP7_75t_L g628 ( .A(n_629), .Y(n_628) );
NAND2xp5_ASAP7_75t_L g715 ( .A(n_629), .B(n_641), .Y(n_715) );
NAND2xp5_ASAP7_75t_L g726 ( .A(n_629), .B(n_639), .Y(n_726) );
AOI221xp5_ASAP7_75t_L g748 ( .A1(n_629), .A2(n_659), .B1(n_749), .B2(n_752), .C(n_754), .Y(n_748) );
CKINVDCx16_ASAP7_75t_R g631 ( .A(n_632), .Y(n_631) );
NAND2xp5_ASAP7_75t_L g633 ( .A(n_634), .B(n_635), .Y(n_633) );
AND2x2_ASAP7_75t_L g654 ( .A(n_634), .B(n_655), .Y(n_654) );
AOI222xp33_ASAP7_75t_L g636 ( .A1(n_637), .A2(n_643), .B1(n_646), .B2(n_649), .C1(n_651), .C2(n_652), .Y(n_636) );
NAND2xp5_ASAP7_75t_SL g637 ( .A(n_638), .B(n_640), .Y(n_637) );
INVx1_ASAP7_75t_L g719 ( .A(n_638), .Y(n_719) );
INVx1_ASAP7_75t_L g741 ( .A(n_641), .Y(n_741) );
INVx2_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
OAI22xp5_ASAP7_75t_L g754 ( .A1(n_644), .A2(n_755), .B1(n_757), .B2(n_758), .Y(n_754) );
INVx1_ASAP7_75t_L g660 ( .A(n_645), .Y(n_660) );
INVx1_ASAP7_75t_SL g647 ( .A(n_648), .Y(n_647) );
INVx1_ASAP7_75t_L g649 ( .A(n_650), .Y(n_649) );
AOI221xp5_ASAP7_75t_L g653 ( .A1(n_654), .A2(n_657), .B1(n_659), .B2(n_661), .C(n_664), .Y(n_653) );
INVx1_ASAP7_75t_SL g655 ( .A(n_656), .Y(n_655) );
OR2x2_ASAP7_75t_L g698 ( .A(n_656), .B(n_699), .Y(n_698) );
OR2x2_ASAP7_75t_L g750 ( .A(n_656), .B(n_751), .Y(n_750) );
INVx1_ASAP7_75t_L g657 ( .A(n_658), .Y(n_657) );
INVx1_ASAP7_75t_L g725 ( .A(n_661), .Y(n_725) );
AND2x2_ASAP7_75t_L g661 ( .A(n_662), .B(n_663), .Y(n_661) );
INVx1_ASAP7_75t_L g689 ( .A(n_662), .Y(n_689) );
INVx1_ASAP7_75t_L g671 ( .A(n_663), .Y(n_671) );
NAND2xp5_ASAP7_75t_L g758 ( .A(n_666), .B(n_753), .Y(n_758) );
AOI22xp33_ASAP7_75t_L g668 ( .A1(n_669), .A2(n_672), .B1(n_675), .B2(n_676), .Y(n_668) );
INVx1_ASAP7_75t_L g669 ( .A(n_670), .Y(n_669) );
INVx1_ASAP7_75t_SL g673 ( .A(n_674), .Y(n_673) );
INVx1_ASAP7_75t_SL g762 ( .A(n_675), .Y(n_762) );
INVxp33_ASAP7_75t_L g676 ( .A(n_677), .Y(n_676) );
NOR2xp33_ASAP7_75t_L g720 ( .A(n_677), .B(n_721), .Y(n_720) );
OAI32xp33_ASAP7_75t_L g711 ( .A1(n_678), .A2(n_712), .A3(n_713), .B1(n_714), .B2(n_715), .Y(n_711) );
NAND4xp25_ASAP7_75t_L g679 ( .A(n_680), .B(n_692), .C(n_704), .D(n_716), .Y(n_679) );
INVx1_ASAP7_75t_SL g681 ( .A(n_682), .Y(n_681) );
NAND2xp33_ASAP7_75t_SL g683 ( .A(n_684), .B(n_685), .Y(n_683) );
NAND2xp5_ASAP7_75t_L g685 ( .A(n_686), .B(n_687), .Y(n_685) );
NAND2xp5_ASAP7_75t_L g735 ( .A(n_687), .B(n_736), .Y(n_735) );
AND2x2_ASAP7_75t_L g688 ( .A(n_689), .B(n_690), .Y(n_688) );
INVx1_ASAP7_75t_L g695 ( .A(n_696), .Y(n_695) );
CKINVDCx16_ASAP7_75t_R g697 ( .A(n_698), .Y(n_697) );
AOI221xp5_ASAP7_75t_L g733 ( .A1(n_701), .A2(n_717), .B1(n_734), .B2(n_737), .C(n_738), .Y(n_733) );
INVx1_ASAP7_75t_L g701 ( .A(n_702), .Y(n_701) );
AND2x2_ASAP7_75t_L g752 ( .A(n_703), .B(n_753), .Y(n_752) );
AOI221xp5_ASAP7_75t_L g704 ( .A1(n_705), .A2(n_707), .B1(n_708), .B2(n_710), .C(n_711), .Y(n_704) );
INVx1_ASAP7_75t_SL g705 ( .A(n_706), .Y(n_705) );
INVx1_ASAP7_75t_L g708 ( .A(n_709), .Y(n_708) );
NOR2xp33_ASAP7_75t_L g743 ( .A(n_713), .B(n_744), .Y(n_743) );
AOI21xp5_ASAP7_75t_L g716 ( .A1(n_717), .A2(n_719), .B(n_720), .Y(n_716) );
INVx1_ASAP7_75t_L g717 ( .A(n_718), .Y(n_717) );
NAND4xp25_ASAP7_75t_L g722 ( .A(n_723), .B(n_733), .C(n_748), .D(n_759), .Y(n_722) );
O2A1O1Ixp33_ASAP7_75t_L g723 ( .A1(n_724), .A2(n_727), .B(n_729), .C(n_731), .Y(n_723) );
NAND2xp5_ASAP7_75t_SL g724 ( .A(n_725), .B(n_726), .Y(n_724) );
INVx1_ASAP7_75t_L g727 ( .A(n_728), .Y(n_727) );
INVx1_ASAP7_75t_L g729 ( .A(n_730), .Y(n_729) );
INVxp67_ASAP7_75t_L g734 ( .A(n_735), .Y(n_734) );
INVx1_ASAP7_75t_SL g739 ( .A(n_740), .Y(n_739) );
INVx1_ASAP7_75t_L g746 ( .A(n_747), .Y(n_746) );
INVx1_ASAP7_75t_L g749 ( .A(n_750), .Y(n_749) );
INVx1_ASAP7_75t_L g764 ( .A(n_751), .Y(n_764) );
INVx2_ASAP7_75t_L g755 ( .A(n_756), .Y(n_755) );
OAI21xp5_ASAP7_75t_L g759 ( .A1(n_760), .A2(n_763), .B(n_764), .Y(n_759) );
NOR2xp33_ASAP7_75t_L g760 ( .A(n_761), .B(n_762), .Y(n_760) );
INVx1_ASAP7_75t_L g779 ( .A(n_765), .Y(n_779) );
INVx1_ASAP7_75t_L g766 ( .A(n_767), .Y(n_766) );
INVx1_ASAP7_75t_L g769 ( .A(n_770), .Y(n_769) );
CKINVDCx14_ASAP7_75t_R g774 ( .A(n_771), .Y(n_774) );
INVx2_ASAP7_75t_L g778 ( .A(n_779), .Y(n_778) );
INVx2_ASAP7_75t_L g780 ( .A(n_781), .Y(n_780) );
INVx2_ASAP7_75t_L g781 ( .A(n_782), .Y(n_781) );
INVx1_ASAP7_75t_SL g783 ( .A(n_784), .Y(n_783) );
endmodule