module real_aes_8272_n_350 (n_76, n_113, n_187, n_90, n_257, n_65, n_74, n_185, n_285, n_30, n_222, n_61, n_20, n_287, n_64, n_254, n_207, n_10, n_83, n_181, n_124, n_191, n_209, n_299, n_322, n_328, n_19, n_40, n_318, n_239, n_100, n_54, n_112, n_319, n_35, n_42, n_329, n_132, n_131, n_144, n_169, n_242, n_308, n_172, n_341, n_232, n_6, n_69, n_317, n_321, n_73, n_320, n_77, n_260, n_37, n_97, n_186, n_138, n_26, n_235, n_245, n_161, n_189, n_271, n_2, n_145, n_227, n_92, n_330, n_332, n_292, n_116, n_94, n_289, n_280, n_333, n_213, n_184, n_28, n_202, n_56, n_34, n_98, n_121, n_125, n_216, n_82, n_327, n_47, n_106, n_32, n_263, n_230, n_51, n_248, n_301, n_27, n_343, n_174, n_18, n_104, n_211, n_281, n_173, n_234, n_284, n_153, n_316, n_75, n_178, n_298, n_49, n_43, n_297, n_9, n_119, n_310, n_164, n_231, n_44, n_102, n_122, n_141, n_128, n_111, n_167, n_80, n_179, n_12, n_68, n_129, n_345, n_304, n_311, n_324, n_25, n_278, n_236, n_267, n_218, n_48, n_204, n_339, n_89, n_277, n_331, n_93, n_182, n_323, n_199, n_142, n_223, n_67, n_250, n_85, n_45, n_5, n_244, n_118, n_139, n_87, n_171, n_78, n_146, n_17, n_226, n_255, n_286, n_120, n_261, n_238, n_58, n_165, n_246, n_176, n_163, n_29, n_52, n_251, n_220, n_197, n_296, n_3, n_41, n_256, n_71, n_302, n_126, n_200, n_115, n_96, n_110, n_150, n_147, n_288, n_23, n_334, n_274, n_160, n_303, n_95, n_188, n_269, n_201, n_306, n_158, n_4, n_346, n_193, n_293, n_162, n_275, n_214, n_46, n_109, n_59, n_203, n_81, n_133, n_273, n_114, n_276, n_295, n_265, n_154, n_127, n_326, n_24, n_217, n_55, n_62, n_291, n_148, n_88, n_159, n_11, n_108, n_60, n_233, n_290, n_155, n_243, n_268, n_136, n_157, n_282, n_101, n_309, n_344, n_229, n_107, n_33, n_53, n_36, n_149, n_190, n_262, n_134, n_349, n_336, n_195, n_300, n_252, n_283, n_314, n_249, n_221, n_156, n_57, n_66, n_21, n_31, n_8, n_312, n_183, n_266, n_205, n_335, n_177, n_313, n_22, n_140, n_219, n_180, n_212, n_210, n_325, n_338, n_103, n_166, n_224, n_151, n_130, n_253, n_99, n_15, n_72, n_152, n_198, n_7, n_228, n_272, n_196, n_347, n_315, n_123, n_279, n_79, n_270, n_305, n_117, n_208, n_215, n_135, n_70, n_50, n_170, n_86, n_340, n_13, n_168, n_175, n_241, n_105, n_84, n_294, n_258, n_206, n_307, n_342, n_348, n_14, n_194, n_137, n_225, n_16, n_39, n_337, n_247, n_240, n_38, n_259, n_143, n_192, n_0, n_264, n_63, n_1, n_237, n_91, n_350);
input n_76;
input n_113;
input n_187;
input n_90;
input n_257;
input n_65;
input n_74;
input n_185;
input n_285;
input n_30;
input n_222;
input n_61;
input n_20;
input n_287;
input n_64;
input n_254;
input n_207;
input n_10;
input n_83;
input n_181;
input n_124;
input n_191;
input n_209;
input n_299;
input n_322;
input n_328;
input n_19;
input n_40;
input n_318;
input n_239;
input n_100;
input n_54;
input n_112;
input n_319;
input n_35;
input n_42;
input n_329;
input n_132;
input n_131;
input n_144;
input n_169;
input n_242;
input n_308;
input n_172;
input n_341;
input n_232;
input n_6;
input n_69;
input n_317;
input n_321;
input n_73;
input n_320;
input n_77;
input n_260;
input n_37;
input n_97;
input n_186;
input n_138;
input n_26;
input n_235;
input n_245;
input n_161;
input n_189;
input n_271;
input n_2;
input n_145;
input n_227;
input n_92;
input n_330;
input n_332;
input n_292;
input n_116;
input n_94;
input n_289;
input n_280;
input n_333;
input n_213;
input n_184;
input n_28;
input n_202;
input n_56;
input n_34;
input n_98;
input n_121;
input n_125;
input n_216;
input n_82;
input n_327;
input n_47;
input n_106;
input n_32;
input n_263;
input n_230;
input n_51;
input n_248;
input n_301;
input n_27;
input n_343;
input n_174;
input n_18;
input n_104;
input n_211;
input n_281;
input n_173;
input n_234;
input n_284;
input n_153;
input n_316;
input n_75;
input n_178;
input n_298;
input n_49;
input n_43;
input n_297;
input n_9;
input n_119;
input n_310;
input n_164;
input n_231;
input n_44;
input n_102;
input n_122;
input n_141;
input n_128;
input n_111;
input n_167;
input n_80;
input n_179;
input n_12;
input n_68;
input n_129;
input n_345;
input n_304;
input n_311;
input n_324;
input n_25;
input n_278;
input n_236;
input n_267;
input n_218;
input n_48;
input n_204;
input n_339;
input n_89;
input n_277;
input n_331;
input n_93;
input n_182;
input n_323;
input n_199;
input n_142;
input n_223;
input n_67;
input n_250;
input n_85;
input n_45;
input n_5;
input n_244;
input n_118;
input n_139;
input n_87;
input n_171;
input n_78;
input n_146;
input n_17;
input n_226;
input n_255;
input n_286;
input n_120;
input n_261;
input n_238;
input n_58;
input n_165;
input n_246;
input n_176;
input n_163;
input n_29;
input n_52;
input n_251;
input n_220;
input n_197;
input n_296;
input n_3;
input n_41;
input n_256;
input n_71;
input n_302;
input n_126;
input n_200;
input n_115;
input n_96;
input n_110;
input n_150;
input n_147;
input n_288;
input n_23;
input n_334;
input n_274;
input n_160;
input n_303;
input n_95;
input n_188;
input n_269;
input n_201;
input n_306;
input n_158;
input n_4;
input n_346;
input n_193;
input n_293;
input n_162;
input n_275;
input n_214;
input n_46;
input n_109;
input n_59;
input n_203;
input n_81;
input n_133;
input n_273;
input n_114;
input n_276;
input n_295;
input n_265;
input n_154;
input n_127;
input n_326;
input n_24;
input n_217;
input n_55;
input n_62;
input n_291;
input n_148;
input n_88;
input n_159;
input n_11;
input n_108;
input n_60;
input n_233;
input n_290;
input n_155;
input n_243;
input n_268;
input n_136;
input n_157;
input n_282;
input n_101;
input n_309;
input n_344;
input n_229;
input n_107;
input n_33;
input n_53;
input n_36;
input n_149;
input n_190;
input n_262;
input n_134;
input n_349;
input n_336;
input n_195;
input n_300;
input n_252;
input n_283;
input n_314;
input n_249;
input n_221;
input n_156;
input n_57;
input n_66;
input n_21;
input n_31;
input n_8;
input n_312;
input n_183;
input n_266;
input n_205;
input n_335;
input n_177;
input n_313;
input n_22;
input n_140;
input n_219;
input n_180;
input n_212;
input n_210;
input n_325;
input n_338;
input n_103;
input n_166;
input n_224;
input n_151;
input n_130;
input n_253;
input n_99;
input n_15;
input n_72;
input n_152;
input n_198;
input n_7;
input n_228;
input n_272;
input n_196;
input n_347;
input n_315;
input n_123;
input n_279;
input n_79;
input n_270;
input n_305;
input n_117;
input n_208;
input n_215;
input n_135;
input n_70;
input n_50;
input n_170;
input n_86;
input n_340;
input n_13;
input n_168;
input n_175;
input n_241;
input n_105;
input n_84;
input n_294;
input n_258;
input n_206;
input n_307;
input n_342;
input n_348;
input n_14;
input n_194;
input n_137;
input n_225;
input n_16;
input n_39;
input n_337;
input n_247;
input n_240;
input n_38;
input n_259;
input n_143;
input n_192;
input n_0;
input n_264;
input n_63;
input n_1;
input n_237;
input n_91;
output n_350;
wire n_480;
wire n_476;
wire n_758;
wire n_887;
wire n_436;
wire n_599;
wire n_684;
wire n_390;
wire n_821;
wire n_830;
wire n_624;
wire n_1018;
wire n_980;
wire n_800;
wire n_618;
wire n_778;
wire n_522;
wire n_838;
wire n_933;
wire n_485;
wire n_822;
wire n_846;
wire n_750;
wire n_631;
wire n_943;
wire n_977;
wire n_357;
wire n_503;
wire n_792;
wire n_386;
wire n_673;
wire n_635;
wire n_518;
wire n_905;
wire n_878;
wire n_665;
wire n_667;
wire n_991;
wire n_1004;
wire n_577;
wire n_580;
wire n_469;
wire n_987;
wire n_362;
wire n_979;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_657;
wire n_900;
wire n_718;
wire n_841;
wire n_355;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_364;
wire n_555;
wire n_421;
wire n_766;
wire n_852;
wire n_974;
wire n_919;
wire n_857;
wire n_461;
wire n_1016;
wire n_908;
wire n_376;
wire n_571;
wire n_549;
wire n_694;
wire n_491;
wire n_894;
wire n_923;
wire n_1034;
wire n_952;
wire n_429;
wire n_752;
wire n_448;
wire n_556;
wire n_545;
wire n_593;
wire n_460;
wire n_937;
wire n_773;
wire n_989;
wire n_401;
wire n_538;
wire n_353;
wire n_431;
wire n_1044;
wire n_963;
wire n_865;
wire n_537;
wire n_551;
wire n_666;
wire n_884;
wire n_560;
wire n_660;
wire n_814;
wire n_944;
wire n_886;
wire n_856;
wire n_594;
wire n_983;
wire n_767;
wire n_696;
wire n_889;
wire n_955;
wire n_975;
wire n_704;
wire n_941;
wire n_379;
wire n_374;
wire n_453;
wire n_932;
wire n_647;
wire n_399;
wire n_948;
wire n_700;
wire n_1021;
wire n_958;
wire n_677;
wire n_378;
wire n_591;
wire n_775;
wire n_763;
wire n_870;
wire n_961;
wire n_489;
wire n_427;
wire n_678;
wire n_548;
wire n_1040;
wire n_415;
wire n_572;
wire n_564;
wire n_815;
wire n_519;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_626;
wire n_539;
wire n_400;
wire n_816;
wire n_625;
wire n_953;
wire n_462;
wire n_615;
wire n_990;
wire n_550;
wire n_966;
wire n_670;
wire n_818;
wire n_716;
wire n_883;
wire n_356;
wire n_478;
wire n_918;
wire n_584;
wire n_896;
wire n_408;
wire n_553;
wire n_892;
wire n_372;
wire n_528;
wire n_578;
wire n_495;
wire n_994;
wire n_370;
wire n_384;
wire n_744;
wire n_938;
wire n_352;
wire n_935;
wire n_824;
wire n_467;
wire n_875;
wire n_951;
wire n_774;
wire n_992;
wire n_813;
wire n_981;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_872;
wire n_976;
wire n_906;
wire n_477;
wire n_515;
wire n_984;
wire n_1019;
wire n_680;
wire n_595;
wire n_726;
wire n_369;
wire n_517;
wire n_931;
wire n_780;
wire n_683;
wire n_840;
wire n_570;
wire n_675;
wire n_904;
wire n_920;
wire n_530;
wire n_835;
wire n_535;
wire n_732;
wire n_834;
wire n_882;
wire n_784;
wire n_496;
wire n_962;
wire n_693;
wire n_468;
wire n_746;
wire n_532;
wire n_1025;
wire n_656;
wire n_755;
wire n_409;
wire n_748;
wire n_781;
wire n_909;
wire n_996;
wire n_523;
wire n_860;
wire n_439;
wire n_576;
wire n_924;
wire n_956;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_874;
wire n_796;
wire n_801;
wire n_383;
wire n_529;
wire n_455;
wire n_504;
wire n_725;
wire n_960;
wire n_671;
wire n_973;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_903;
wire n_454;
wire n_812;
wire n_782;
wire n_443;
wire n_565;
wire n_817;
wire n_760;
wire n_608;
wire n_925;
wire n_534;
wire n_708;
wire n_1029;
wire n_1020;
wire n_457;
wire n_885;
wire n_950;
wire n_381;
wire n_993;
wire n_493;
wire n_664;
wire n_367;
wire n_819;
wire n_737;
wire n_1013;
wire n_1017;
wire n_581;
wire n_610;
wire n_936;
wire n_1035;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_940;
wire n_745;
wire n_722;
wire n_867;
wire n_398;
wire n_688;
wire n_425;
wire n_609;
wire n_1042;
wire n_879;
wire n_417;
wire n_363;
wire n_449;
wire n_607;
wire n_754;
wire n_1006;
wire n_690;
wire n_629;
wire n_499;
wire n_508;
wire n_706;
wire n_901;
wire n_561;
wire n_970;
wire n_947;
wire n_876;
wire n_437;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_1012;
wire n_655;
wire n_654;
wire n_527;
wire n_505;
wire n_434;
wire n_502;
wire n_769;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_672;
wire n_567;
wire n_916;
wire n_406;
wire n_426;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_658;
wire n_676;
wire n_986;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_880;
wire n_1031;
wire n_1037;
wire n_1008;
wire n_807;
wire n_1011;
wire n_416;
wire n_790;
wire n_895;
wire n_832;
wire n_410;
wire n_799;
wire n_805;
wire n_751;
wire n_999;
wire n_490;
wire n_913;
wire n_619;
wire n_391;
wire n_360;
wire n_859;
wire n_695;
wire n_685;
wire n_881;
wire n_361;
wire n_917;
wire n_632;
wire n_768;
wire n_412;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_985;
wire n_488;
wire n_1041;
wire n_501;
wire n_910;
wire n_642;
wire n_613;
wire n_869;
wire n_387;
wire n_957;
wire n_995;
wire n_702;
wire n_954;
wire n_969;
wire n_912;
wire n_1009;
wire n_1007;
wire n_464;
wire n_351;
wire n_945;
wire n_604;
wire n_734;
wire n_898;
wire n_848;
wire n_392;
wire n_562;
wire n_1022;
wire n_404;
wire n_598;
wire n_713;
wire n_735;
wire n_728;
wire n_756;
wire n_569;
wire n_997;
wire n_563;
wire n_785;
wire n_891;
wire n_430;
wire n_568;
wire n_413;
wire n_471;
wire n_902;
wire n_853;
wire n_810;
wire n_843;
wire n_579;
wire n_1033;
wire n_699;
wire n_533;
wire n_1000;
wire n_1003;
wire n_1028;
wire n_366;
wire n_727;
wire n_1014;
wire n_649;
wire n_358;
wire n_385;
wire n_397;
wire n_663;
wire n_749;
wire n_588;
wire n_536;
wire n_914;
wire n_707;
wire n_622;
wire n_470;
wire n_851;
wire n_915;
wire n_1002;
wire n_934;
wire n_494;
wire n_1001;
wire n_711;
wire n_864;
wire n_1027;
wire n_377;
wire n_927;
wire n_1038;
wire n_965;
wire n_723;
wire n_662;
wire n_382;
wire n_845;
wire n_850;
wire n_1043;
wire n_354;
wire n_720;
wire n_972;
wire n_435;
wire n_1026;
wire n_511;
wire n_484;
wire n_893;
wire n_492;
wire n_509;
wire n_407;
wire n_419;
wire n_730;
wire n_1023;
wire n_643;
wire n_747;
wire n_486;
wire n_930;
wire n_411;
wire n_697;
wire n_978;
wire n_907;
wire n_847;
wire n_779;
wire n_498;
wire n_481;
wire n_765;
wire n_691;
wire n_826;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_939;
wire n_1005;
wire n_487;
wire n_831;
wire n_365;
wire n_899;
wire n_637;
wire n_928;
wire n_526;
wire n_653;
wire n_692;
wire n_544;
wire n_789;
wire n_389;
wire n_738;
wire n_701;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_922;
wire n_926;
wire n_942;
wire n_472;
wire n_971;
wire n_866;
wire n_452;
wire n_787;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_959;
wire n_715;
wire n_946;
wire n_420;
wire n_612;
wire n_858;
wire n_873;
wire n_438;
wire n_764;
wire n_794;
wire n_753;
wire n_741;
wire n_623;
wire n_1032;
wire n_446;
wire n_721;
wire n_681;
wire n_982;
wire n_359;
wire n_456;
wire n_717;
wire n_712;
wire n_433;
wire n_516;
wire n_627;
wire n_739;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_524;
wire n_861;
wire n_705;
wire n_575;
wire n_762;
wire n_479;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_541;
wire n_839;
wire n_546;
wire n_587;
wire n_639;
wire n_1010;
wire n_811;
wire n_1015;
wire n_459;
wire n_558;
wire n_863;
wire n_998;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_836;
wire n_888;
wire n_793;
wire n_583;
wire n_833;
wire n_414;
wire n_757;
wire n_929;
wire n_686;
wire n_776;
wire n_803;
wire n_890;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_949;
wire n_614;
wire n_586;
wire n_911;
wire n_772;
wire n_450;
wire n_788;
wire n_441;
wire n_585;
wire n_465;
wire n_719;
wire n_473;
wire n_967;
wire n_566;
wire n_837;
wire n_1045;
wire n_871;
wire n_474;
wire n_829;
wire n_1030;
wire n_988;
wire n_921;
wire n_375;
wire n_597;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_1036;
wire n_394;
wire n_687;
wire n_729;
wire n_844;
wire n_968;
wire n_650;
wire n_646;
wire n_743;
wire n_710;
wire n_393;
wire n_652;
wire n_703;
wire n_823;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_603;
wire n_403;
wire n_854;
wire n_424;
wire n_877;
wire n_802;
wire n_868;
wire n_1039;
wire n_574;
wire n_1024;
wire n_842;
wire n_849;
wire n_554;
wire n_475;
wire n_897;
wire n_855;
wire n_798;
wire n_668;
wire n_797;
wire n_862;
AOI22xp33_ASAP7_75t_L g966 ( .A1(n_0), .A2(n_175), .B1(n_967), .B2(n_968), .Y(n_966) );
INVx1_ASAP7_75t_L g825 ( .A(n_1), .Y(n_825) );
AOI22xp33_ASAP7_75t_SL g536 ( .A1(n_2), .A2(n_222), .B1(n_472), .B2(n_537), .Y(n_536) );
AOI222xp33_ASAP7_75t_L g767 ( .A1(n_3), .A2(n_167), .B1(n_307), .B2(n_442), .C1(n_550), .C2(n_649), .Y(n_767) );
AOI22xp33_ASAP7_75t_L g616 ( .A1(n_4), .A2(n_235), .B1(n_369), .B2(n_386), .Y(n_616) );
AOI211xp5_ASAP7_75t_L g350 ( .A1(n_5), .A2(n_351), .B(n_360), .C(n_996), .Y(n_350) );
AOI22xp33_ASAP7_75t_L g1002 ( .A1(n_6), .A2(n_101), .B1(n_402), .B2(n_887), .Y(n_1002) );
AOI221xp5_ASAP7_75t_L g401 ( .A1(n_7), .A2(n_302), .B1(n_402), .B2(n_406), .C(n_411), .Y(n_401) );
AOI22xp33_ASAP7_75t_SL g744 ( .A1(n_8), .A2(n_148), .B1(n_745), .B2(n_746), .Y(n_744) );
AOI22xp5_ASAP7_75t_L g699 ( .A1(n_9), .A2(n_92), .B1(n_470), .B2(n_700), .Y(n_699) );
AOI22xp33_ASAP7_75t_L g607 ( .A1(n_10), .A2(n_77), .B1(n_550), .B2(n_586), .Y(n_607) );
NAND2xp5_ASAP7_75t_SL g738 ( .A(n_11), .B(n_739), .Y(n_738) );
AO22x2_ASAP7_75t_L g383 ( .A1(n_12), .A2(n_208), .B1(n_375), .B2(n_380), .Y(n_383) );
INVx1_ASAP7_75t_L g994 ( .A(n_12), .Y(n_994) );
AOI22xp33_ASAP7_75t_L g761 ( .A1(n_13), .A2(n_159), .B1(n_542), .B2(n_562), .Y(n_761) );
AOI22xp33_ASAP7_75t_SL g866 ( .A1(n_14), .A2(n_331), .B1(n_446), .B2(n_555), .Y(n_866) );
AOI22xp5_ASAP7_75t_L g915 ( .A1(n_15), .A2(n_145), .B1(n_407), .B2(n_750), .Y(n_915) );
CKINVDCx20_ASAP7_75t_R g935 ( .A(n_16), .Y(n_935) );
CKINVDCx20_ASAP7_75t_R g946 ( .A(n_17), .Y(n_946) );
AOI22xp33_ASAP7_75t_L g558 ( .A1(n_18), .A2(n_181), .B1(n_423), .B2(n_426), .Y(n_558) );
AOI22xp33_ASAP7_75t_L g859 ( .A1(n_19), .A2(n_231), .B1(n_407), .B2(n_722), .Y(n_859) );
AOI22xp33_ASAP7_75t_L g1006 ( .A1(n_20), .A2(n_297), .B1(n_698), .B2(n_892), .Y(n_1006) );
AOI222xp33_ASAP7_75t_L g725 ( .A1(n_21), .A2(n_63), .B1(n_259), .B2(n_446), .C1(n_726), .C2(n_727), .Y(n_725) );
AOI22xp33_ASAP7_75t_SL g894 ( .A1(n_22), .A2(n_286), .B1(n_393), .B2(n_895), .Y(n_894) );
AOI22xp5_ASAP7_75t_SL g855 ( .A1(n_23), .A2(n_227), .B1(n_750), .B2(n_856), .Y(n_855) );
CKINVDCx20_ASAP7_75t_R g902 ( .A(n_24), .Y(n_902) );
AOI221xp5_ASAP7_75t_L g421 ( .A1(n_25), .A2(n_36), .B1(n_422), .B2(n_426), .C(n_428), .Y(n_421) );
AOI22xp33_ASAP7_75t_SL g886 ( .A1(n_26), .A2(n_284), .B1(n_787), .B2(n_887), .Y(n_886) );
AOI22xp33_ASAP7_75t_L g541 ( .A1(n_27), .A2(n_233), .B1(n_369), .B2(n_542), .Y(n_541) );
AOI22xp33_ASAP7_75t_L g916 ( .A1(n_28), .A2(n_335), .B1(n_724), .B2(n_746), .Y(n_916) );
CKINVDCx20_ASAP7_75t_R g929 ( .A(n_29), .Y(n_929) );
AOI22xp33_ASAP7_75t_L g561 ( .A1(n_30), .A2(n_225), .B1(n_470), .B2(n_562), .Y(n_561) );
CKINVDCx20_ASAP7_75t_R g1033 ( .A(n_31), .Y(n_1033) );
AO22x2_ASAP7_75t_L g385 ( .A1(n_32), .A2(n_115), .B1(n_375), .B2(n_376), .Y(n_385) );
AOI22xp33_ASAP7_75t_L g568 ( .A1(n_33), .A2(n_163), .B1(n_394), .B2(n_418), .Y(n_568) );
CKINVDCx20_ASAP7_75t_R g729 ( .A(n_34), .Y(n_729) );
AOI22xp5_ASAP7_75t_L g952 ( .A1(n_35), .A2(n_953), .B1(n_974), .B2(n_975), .Y(n_952) );
INVx1_ASAP7_75t_L g975 ( .A(n_35), .Y(n_975) );
AOI22xp33_ASAP7_75t_SL g566 ( .A1(n_37), .A2(n_59), .B1(n_542), .B2(n_567), .Y(n_566) );
CKINVDCx20_ASAP7_75t_R g690 ( .A(n_38), .Y(n_690) );
INVx1_ASAP7_75t_L g803 ( .A(n_39), .Y(n_803) );
AOI22xp5_ASAP7_75t_L g549 ( .A1(n_40), .A2(n_270), .B1(n_550), .B2(n_551), .Y(n_549) );
AOI22xp5_ASAP7_75t_L g464 ( .A1(n_41), .A2(n_60), .B1(n_404), .B2(n_465), .Y(n_464) );
AOI22xp33_ASAP7_75t_L g783 ( .A1(n_42), .A2(n_152), .B1(n_562), .B2(n_666), .Y(n_783) );
INVx1_ASAP7_75t_L g415 ( .A(n_43), .Y(n_415) );
AOI22xp33_ASAP7_75t_L g972 ( .A1(n_44), .A2(n_281), .B1(n_402), .B2(n_472), .Y(n_972) );
INVx1_ASAP7_75t_L g779 ( .A(n_45), .Y(n_779) );
AOI22xp5_ASAP7_75t_L g801 ( .A1(n_46), .A2(n_197), .B1(n_452), .B2(n_491), .Y(n_801) );
AOI222xp33_ASAP7_75t_L g441 ( .A1(n_47), .A2(n_130), .B1(n_137), .B2(n_442), .C1(n_444), .C2(n_450), .Y(n_441) );
AOI22xp5_ASAP7_75t_SL g854 ( .A1(n_48), .A2(n_293), .B1(n_386), .B2(n_461), .Y(n_854) );
AOI222xp33_ASAP7_75t_L g1011 ( .A1(n_49), .A2(n_278), .B1(n_296), .B2(n_554), .C1(n_907), .C2(n_959), .Y(n_1011) );
CKINVDCx20_ASAP7_75t_R g768 ( .A(n_50), .Y(n_768) );
AOI22xp5_ASAP7_75t_SL g460 ( .A1(n_51), .A2(n_206), .B1(n_407), .B2(n_461), .Y(n_460) );
AOI22xp33_ASAP7_75t_SL g878 ( .A1(n_52), .A2(n_71), .B1(n_444), .B2(n_489), .Y(n_878) );
CKINVDCx20_ASAP7_75t_R g933 ( .A(n_53), .Y(n_933) );
AOI22xp33_ASAP7_75t_L g660 ( .A1(n_54), .A2(n_165), .B1(n_417), .B2(n_661), .Y(n_660) );
AOI22xp33_ASAP7_75t_L g717 ( .A1(n_55), .A2(n_303), .B1(n_718), .B2(n_719), .Y(n_717) );
CKINVDCx16_ASAP7_75t_R g925 ( .A(n_56), .Y(n_925) );
AOI22xp33_ASAP7_75t_L g642 ( .A1(n_57), .A2(n_280), .B1(n_643), .B2(n_645), .Y(n_642) );
CKINVDCx20_ASAP7_75t_R g682 ( .A(n_58), .Y(n_682) );
CKINVDCx20_ASAP7_75t_R g569 ( .A(n_61), .Y(n_569) );
AOI22xp33_ASAP7_75t_SL g847 ( .A1(n_62), .A2(n_226), .B1(n_531), .B2(n_848), .Y(n_847) );
AOI22xp5_ASAP7_75t_L g780 ( .A1(n_64), .A2(n_91), .B1(n_550), .B2(n_719), .Y(n_780) );
AOI22xp33_ASAP7_75t_SL g742 ( .A1(n_65), .A2(n_123), .B1(n_564), .B2(n_743), .Y(n_742) );
INVx1_ASAP7_75t_L g822 ( .A(n_66), .Y(n_822) );
NAND2xp5_ASAP7_75t_SL g812 ( .A(n_67), .B(n_473), .Y(n_812) );
CKINVDCx20_ASAP7_75t_R g956 ( .A(n_68), .Y(n_956) );
AOI22xp33_ASAP7_75t_SL g530 ( .A1(n_69), .A2(n_191), .B1(n_531), .B2(n_534), .Y(n_530) );
AOI22xp33_ASAP7_75t_L g1037 ( .A1(n_70), .A2(n_103), .B1(n_531), .B2(n_1038), .Y(n_1037) );
AOI22xp33_ASAP7_75t_L g615 ( .A1(n_72), .A2(n_90), .B1(n_527), .B2(n_529), .Y(n_615) );
AOI22xp33_ASAP7_75t_L g867 ( .A1(n_73), .A2(n_204), .B1(n_423), .B2(n_427), .Y(n_867) );
CKINVDCx20_ASAP7_75t_R g913 ( .A(n_74), .Y(n_913) );
AOI22xp33_ASAP7_75t_L g693 ( .A1(n_75), .A2(n_213), .B1(n_657), .B2(n_658), .Y(n_693) );
INVx1_ASAP7_75t_L g518 ( .A(n_76), .Y(n_518) );
AOI22xp33_ASAP7_75t_SL g850 ( .A1(n_78), .A2(n_211), .B1(n_469), .B2(n_589), .Y(n_850) );
AOI22xp5_ASAP7_75t_SL g468 ( .A1(n_79), .A2(n_96), .B1(n_469), .B2(n_470), .Y(n_468) );
AOI22xp33_ASAP7_75t_L g663 ( .A1(n_80), .A2(n_139), .B1(n_664), .B2(n_667), .Y(n_663) );
AO22x2_ASAP7_75t_L g379 ( .A1(n_81), .A2(n_238), .B1(n_375), .B2(n_380), .Y(n_379) );
INVx1_ASAP7_75t_L g991 ( .A(n_81), .Y(n_991) );
AOI22xp33_ASAP7_75t_SL g526 ( .A1(n_82), .A2(n_83), .B1(n_527), .B2(n_529), .Y(n_526) );
AOI22xp33_ASAP7_75t_L g723 ( .A1(n_84), .A2(n_248), .B1(n_418), .B2(n_724), .Y(n_723) );
AOI22xp33_ASAP7_75t_L g908 ( .A1(n_85), .A2(n_326), .B1(n_727), .B2(n_909), .Y(n_908) );
AOI22xp33_ASAP7_75t_L g918 ( .A1(n_86), .A2(n_323), .B1(n_666), .B2(n_712), .Y(n_918) );
AOI22xp33_ASAP7_75t_L g961 ( .A1(n_87), .A2(n_274), .B1(n_716), .B2(n_962), .Y(n_961) );
AOI22xp5_ASAP7_75t_L g957 ( .A1(n_88), .A2(n_201), .B1(n_958), .B2(n_959), .Y(n_957) );
CKINVDCx20_ASAP7_75t_R g877 ( .A(n_89), .Y(n_877) );
AOI22xp5_ASAP7_75t_L g997 ( .A1(n_93), .A2(n_998), .B1(n_999), .B2(n_1012), .Y(n_997) );
CKINVDCx20_ASAP7_75t_R g1012 ( .A(n_93), .Y(n_1012) );
AOI22xp33_ASAP7_75t_L g694 ( .A1(n_94), .A2(n_268), .B1(n_417), .B2(n_695), .Y(n_694) );
AOI22xp33_ASAP7_75t_L g917 ( .A1(n_95), .A2(n_288), .B1(n_465), .B2(n_743), .Y(n_917) );
AOI22xp33_ASAP7_75t_SL g471 ( .A1(n_97), .A2(n_193), .B1(n_472), .B2(n_473), .Y(n_471) );
AOI22xp5_ASAP7_75t_L g784 ( .A1(n_98), .A2(n_112), .B1(n_470), .B2(n_564), .Y(n_784) );
AOI22xp33_ASAP7_75t_SL g553 ( .A1(n_99), .A2(n_105), .B1(n_554), .B2(n_555), .Y(n_553) );
INVx1_ASAP7_75t_L g457 ( .A(n_100), .Y(n_457) );
AOI22xp33_ASAP7_75t_L g969 ( .A1(n_102), .A2(n_122), .B1(n_702), .B2(n_970), .Y(n_969) );
AOI22xp33_ASAP7_75t_SL g838 ( .A1(n_104), .A2(n_147), .B1(n_645), .B2(n_839), .Y(n_838) );
CKINVDCx20_ASAP7_75t_R g684 ( .A(n_106), .Y(n_684) );
CKINVDCx20_ASAP7_75t_R g862 ( .A(n_107), .Y(n_862) );
CKINVDCx20_ASAP7_75t_R g811 ( .A(n_108), .Y(n_811) );
NAND2xp5_ASAP7_75t_L g774 ( .A(n_109), .B(n_775), .Y(n_774) );
CKINVDCx20_ASAP7_75t_R g804 ( .A(n_110), .Y(n_804) );
CKINVDCx20_ASAP7_75t_R g641 ( .A(n_111), .Y(n_641) );
AOI22xp5_ASAP7_75t_L g588 ( .A1(n_113), .A2(n_258), .B1(n_461), .B2(n_589), .Y(n_588) );
INVx1_ASAP7_75t_L g584 ( .A(n_114), .Y(n_584) );
INVx1_ASAP7_75t_L g995 ( .A(n_115), .Y(n_995) );
AOI22xp33_ASAP7_75t_SL g889 ( .A1(n_116), .A2(n_136), .B1(n_417), .B2(n_890), .Y(n_889) );
CKINVDCx20_ASAP7_75t_R g734 ( .A(n_117), .Y(n_734) );
AOI22xp5_ASAP7_75t_L g581 ( .A1(n_118), .A2(n_189), .B1(n_556), .B2(n_582), .Y(n_581) );
AOI22xp33_ASAP7_75t_L g788 ( .A1(n_119), .A2(n_126), .B1(n_472), .B2(n_591), .Y(n_788) );
OAI22xp5_ASAP7_75t_L g504 ( .A1(n_120), .A2(n_505), .B1(n_506), .B2(n_507), .Y(n_504) );
INVx1_ASAP7_75t_L g505 ( .A(n_120), .Y(n_505) );
CKINVDCx20_ASAP7_75t_R g651 ( .A(n_121), .Y(n_651) );
AOI22xp33_ASAP7_75t_L g656 ( .A1(n_124), .A2(n_192), .B1(n_657), .B2(n_658), .Y(n_656) );
CKINVDCx20_ASAP7_75t_R g479 ( .A(n_125), .Y(n_479) );
AOI211xp5_ASAP7_75t_L g927 ( .A1(n_127), .A2(n_907), .B(n_928), .C(n_932), .Y(n_927) );
INVx1_ASAP7_75t_L g595 ( .A(n_128), .Y(n_595) );
CKINVDCx20_ASAP7_75t_R g808 ( .A(n_129), .Y(n_808) );
CKINVDCx20_ASAP7_75t_R g638 ( .A(n_131), .Y(n_638) );
INVx1_ASAP7_75t_L g789 ( .A(n_132), .Y(n_789) );
AOI22xp5_ASAP7_75t_L g563 ( .A1(n_133), .A2(n_162), .B1(n_539), .B2(n_564), .Y(n_563) );
AOI22xp33_ASAP7_75t_L g1007 ( .A1(n_134), .A2(n_310), .B1(n_594), .B2(n_620), .Y(n_1007) );
AOI22xp5_ASAP7_75t_L g488 ( .A1(n_135), .A2(n_237), .B1(n_489), .B2(n_490), .Y(n_488) );
AOI22xp33_ASAP7_75t_L g777 ( .A1(n_138), .A2(n_333), .B1(n_446), .B2(n_555), .Y(n_777) );
AOI22xp33_ASAP7_75t_L g697 ( .A1(n_140), .A2(n_244), .B1(n_667), .B2(n_698), .Y(n_697) );
AOI22xp33_ASAP7_75t_L g759 ( .A1(n_141), .A2(n_172), .B1(n_418), .B2(n_567), .Y(n_759) );
AOI22xp33_ASAP7_75t_L g931 ( .A1(n_142), .A2(n_332), .B1(n_645), .B2(n_839), .Y(n_931) );
AOI22xp33_ASAP7_75t_L g1010 ( .A1(n_143), .A2(n_252), .B1(n_491), .B2(n_839), .Y(n_1010) );
AOI22xp33_ASAP7_75t_L g973 ( .A1(n_144), .A2(n_217), .B1(n_695), .B2(n_848), .Y(n_973) );
AND2x6_ASAP7_75t_L g355 ( .A(n_146), .B(n_356), .Y(n_355) );
HB1xp67_ASAP7_75t_L g988 ( .A(n_146), .Y(n_988) );
CKINVDCx20_ASAP7_75t_R g806 ( .A(n_149), .Y(n_806) );
CKINVDCx20_ASAP7_75t_R g494 ( .A(n_150), .Y(n_494) );
CKINVDCx20_ASAP7_75t_R g689 ( .A(n_151), .Y(n_689) );
AOI22xp33_ASAP7_75t_SL g786 ( .A1(n_153), .A2(n_328), .B1(n_567), .B2(n_787), .Y(n_786) );
AOI22xp5_ASAP7_75t_L g864 ( .A1(n_154), .A2(n_221), .B1(n_491), .B2(n_550), .Y(n_864) );
CKINVDCx20_ASAP7_75t_R g1025 ( .A(n_155), .Y(n_1025) );
AO22x1_ASAP7_75t_L g391 ( .A1(n_156), .A2(n_168), .B1(n_392), .B2(n_396), .Y(n_391) );
AOI22xp33_ASAP7_75t_SL g748 ( .A1(n_157), .A2(n_340), .B1(n_470), .B2(n_562), .Y(n_748) );
CKINVDCx20_ASAP7_75t_R g751 ( .A(n_158), .Y(n_751) );
AOI221xp5_ASAP7_75t_L g368 ( .A1(n_160), .A2(n_309), .B1(n_369), .B2(n_386), .C(n_391), .Y(n_368) );
AOI22xp33_ASAP7_75t_L g1003 ( .A1(n_161), .A2(n_247), .B1(n_890), .B2(n_1004), .Y(n_1003) );
AOI22xp5_ASAP7_75t_L g585 ( .A1(n_164), .A2(n_346), .B1(n_451), .B2(n_586), .Y(n_585) );
INVx1_ASAP7_75t_L g522 ( .A(n_166), .Y(n_522) );
AOI22xp33_ASAP7_75t_SL g590 ( .A1(n_169), .A2(n_173), .B1(n_393), .B2(n_591), .Y(n_590) );
AOI22xp33_ASAP7_75t_SL g891 ( .A1(n_170), .A2(n_246), .B1(n_892), .B2(n_893), .Y(n_891) );
AO22x2_ASAP7_75t_L g374 ( .A1(n_171), .A2(n_228), .B1(n_375), .B2(n_376), .Y(n_374) );
NOR2xp33_ASAP7_75t_L g992 ( .A(n_171), .B(n_993), .Y(n_992) );
CKINVDCx20_ASAP7_75t_R g903 ( .A(n_174), .Y(n_903) );
AOI22xp33_ASAP7_75t_SL g749 ( .A1(n_176), .A2(n_245), .B1(n_386), .B2(n_750), .Y(n_749) );
AOI22xp33_ASAP7_75t_L g758 ( .A1(n_177), .A2(n_232), .B1(n_465), .B2(n_539), .Y(n_758) );
AOI22xp33_ASAP7_75t_L g835 ( .A1(n_178), .A2(n_285), .B1(n_489), .B2(n_836), .Y(n_835) );
AOI22xp33_ASAP7_75t_SL g592 ( .A1(n_179), .A2(n_318), .B1(n_407), .B2(n_539), .Y(n_592) );
CKINVDCx20_ASAP7_75t_R g687 ( .A(n_180), .Y(n_687) );
CKINVDCx20_ASAP7_75t_R g1026 ( .A(n_182), .Y(n_1026) );
CKINVDCx20_ASAP7_75t_R g1028 ( .A(n_183), .Y(n_1028) );
AOI22xp33_ASAP7_75t_L g519 ( .A1(n_184), .A2(n_349), .B1(n_446), .B2(n_489), .Y(n_519) );
INVx1_ASAP7_75t_L g510 ( .A(n_185), .Y(n_510) );
INVx1_ASAP7_75t_L g521 ( .A(n_186), .Y(n_521) );
AOI22xp5_ASAP7_75t_SL g858 ( .A1(n_187), .A2(n_254), .B1(n_473), .B2(n_846), .Y(n_858) );
CKINVDCx20_ASAP7_75t_R g609 ( .A(n_188), .Y(n_609) );
AOI22xp33_ASAP7_75t_L g711 ( .A1(n_190), .A2(n_220), .B1(n_562), .B2(n_712), .Y(n_711) );
AOI22xp5_ASAP7_75t_L g619 ( .A1(n_194), .A2(n_315), .B1(n_418), .B2(n_620), .Y(n_619) );
CKINVDCx20_ASAP7_75t_R g622 ( .A(n_195), .Y(n_622) );
NAND2xp5_ASAP7_75t_L g765 ( .A(n_196), .B(n_579), .Y(n_765) );
AOI22xp33_ASAP7_75t_SL g884 ( .A1(n_198), .A2(n_229), .B1(n_645), .B2(n_839), .Y(n_884) );
AOI22xp33_ASAP7_75t_L g1030 ( .A1(n_199), .A2(n_207), .B1(n_451), .B2(n_836), .Y(n_1030) );
AOI22xp33_ASAP7_75t_SL g618 ( .A1(n_200), .A2(n_341), .B1(n_402), .B2(n_461), .Y(n_618) );
CKINVDCx20_ASAP7_75t_R g942 ( .A(n_202), .Y(n_942) );
AOI22xp5_ASAP7_75t_L g364 ( .A1(n_203), .A2(n_365), .B1(n_366), .B2(n_454), .Y(n_364) );
INVx1_ASAP7_75t_L g454 ( .A(n_203), .Y(n_454) );
CKINVDCx20_ASAP7_75t_R g905 ( .A(n_205), .Y(n_905) );
AOI22xp5_ASAP7_75t_L g677 ( .A1(n_209), .A2(n_678), .B1(n_703), .B2(n_704), .Y(n_677) );
INVx1_ASAP7_75t_L g703 ( .A(n_209), .Y(n_703) );
AOI22xp33_ASAP7_75t_L g939 ( .A1(n_210), .A2(n_329), .B1(n_594), .B2(n_620), .Y(n_939) );
NAND2xp5_ASAP7_75t_L g580 ( .A(n_212), .B(n_426), .Y(n_580) );
AOI22xp33_ASAP7_75t_L g963 ( .A1(n_214), .A2(n_276), .B1(n_643), .B2(n_645), .Y(n_963) );
AOI22xp33_ASAP7_75t_L g762 ( .A1(n_215), .A2(n_337), .B1(n_393), .B2(n_712), .Y(n_762) );
CKINVDCx20_ASAP7_75t_R g868 ( .A(n_216), .Y(n_868) );
XNOR2xp5_ASAP7_75t_L g873 ( .A(n_218), .B(n_874), .Y(n_873) );
AOI22xp33_ASAP7_75t_SL g844 ( .A1(n_219), .A2(n_249), .B1(n_845), .B2(n_846), .Y(n_844) );
INVx2_ASAP7_75t_L g359 ( .A(n_223), .Y(n_359) );
AOI22xp33_ASAP7_75t_SL g735 ( .A1(n_224), .A2(n_301), .B1(n_446), .B2(n_452), .Y(n_735) );
AOI22xp5_ASAP7_75t_L g1040 ( .A1(n_230), .A2(n_240), .B1(n_698), .B2(n_1041), .Y(n_1040) );
AOI22xp33_ASAP7_75t_L g713 ( .A1(n_234), .A2(n_243), .B1(n_386), .B2(n_589), .Y(n_713) );
AOI22xp33_ASAP7_75t_L g721 ( .A1(n_236), .A2(n_291), .B1(n_564), .B2(n_722), .Y(n_721) );
AOI22xp33_ASAP7_75t_L g940 ( .A1(n_239), .A2(n_290), .B1(n_745), .B2(n_848), .Y(n_940) );
INVx1_ASAP7_75t_L g800 ( .A(n_241), .Y(n_800) );
CKINVDCx20_ASAP7_75t_R g834 ( .A(n_242), .Y(n_834) );
AOI22xp33_ASAP7_75t_L g1036 ( .A1(n_250), .A2(n_343), .B1(n_856), .B2(n_968), .Y(n_1036) );
AOI22xp33_ASAP7_75t_L g1009 ( .A1(n_251), .A2(n_295), .B1(n_422), .B2(n_962), .Y(n_1009) );
NAND2xp5_ASAP7_75t_SL g737 ( .A(n_253), .B(n_426), .Y(n_737) );
CKINVDCx20_ASAP7_75t_R g820 ( .A(n_255), .Y(n_820) );
AOI22xp33_ASAP7_75t_L g668 ( .A1(n_256), .A2(n_305), .B1(n_669), .B2(n_671), .Y(n_668) );
AOI22xp33_ASAP7_75t_L g715 ( .A1(n_257), .A2(n_336), .B1(n_426), .B2(n_716), .Y(n_715) );
AOI22xp33_ASAP7_75t_SL g851 ( .A1(n_260), .A2(n_348), .B1(n_369), .B2(n_527), .Y(n_851) );
CKINVDCx20_ASAP7_75t_R g482 ( .A(n_261), .Y(n_482) );
INVx1_ASAP7_75t_L g375 ( .A(n_262), .Y(n_375) );
INVx1_ASAP7_75t_L g377 ( .A(n_262), .Y(n_377) );
AOI22xp33_ASAP7_75t_L g840 ( .A1(n_263), .A2(n_269), .B1(n_422), .B2(n_841), .Y(n_840) );
AOI22xp33_ASAP7_75t_L g1042 ( .A1(n_264), .A2(n_339), .B1(n_407), .B2(n_750), .Y(n_1042) );
INVx1_ASAP7_75t_L g513 ( .A(n_265), .Y(n_513) );
INVx1_ASAP7_75t_L g604 ( .A(n_266), .Y(n_604) );
AOI22xp5_ASAP7_75t_L g633 ( .A1(n_267), .A2(n_634), .B1(n_672), .B2(n_673), .Y(n_633) );
CKINVDCx20_ASAP7_75t_R g672 ( .A(n_267), .Y(n_672) );
CKINVDCx20_ASAP7_75t_R g814 ( .A(n_271), .Y(n_814) );
CKINVDCx20_ASAP7_75t_R g818 ( .A(n_272), .Y(n_818) );
CKINVDCx20_ASAP7_75t_R g429 ( .A(n_273), .Y(n_429) );
AOI22xp5_ASAP7_75t_L g593 ( .A1(n_275), .A2(n_313), .B1(n_564), .B2(n_594), .Y(n_593) );
INVx1_ASAP7_75t_L g602 ( .A(n_277), .Y(n_602) );
CKINVDCx20_ASAP7_75t_R g496 ( .A(n_279), .Y(n_496) );
AOI22xp33_ASAP7_75t_SL g740 ( .A1(n_282), .A2(n_321), .B1(n_556), .B2(n_719), .Y(n_740) );
CKINVDCx20_ASAP7_75t_R g650 ( .A(n_283), .Y(n_650) );
CKINVDCx20_ASAP7_75t_R g911 ( .A(n_287), .Y(n_911) );
AOI22xp33_ASAP7_75t_L g766 ( .A1(n_289), .A2(n_314), .B1(n_490), .B2(n_555), .Y(n_766) );
NAND2xp5_ASAP7_75t_SL g883 ( .A(n_292), .B(n_423), .Y(n_883) );
AO22x2_ASAP7_75t_L g898 ( .A1(n_294), .A2(n_899), .B1(n_919), .B2(n_920), .Y(n_898) );
CKINVDCx20_ASAP7_75t_R g920 ( .A(n_294), .Y(n_920) );
CKINVDCx20_ASAP7_75t_R g829 ( .A(n_298), .Y(n_829) );
INVx1_ASAP7_75t_L g358 ( .A(n_299), .Y(n_358) );
INVx1_ASAP7_75t_L g356 ( .A(n_300), .Y(n_356) );
NAND2xp5_ASAP7_75t_L g776 ( .A(n_304), .B(n_579), .Y(n_776) );
NAND2xp5_ASAP7_75t_L g880 ( .A(n_306), .B(n_881), .Y(n_880) );
INVx1_ASAP7_75t_L g826 ( .A(n_308), .Y(n_826) );
CKINVDCx20_ASAP7_75t_R g685 ( .A(n_311), .Y(n_685) );
NAND2xp5_ASAP7_75t_L g930 ( .A(n_312), .B(n_716), .Y(n_930) );
CKINVDCx20_ASAP7_75t_R g815 ( .A(n_316), .Y(n_815) );
CKINVDCx20_ASAP7_75t_R g487 ( .A(n_317), .Y(n_487) );
CKINVDCx20_ASAP7_75t_R g681 ( .A(n_319), .Y(n_681) );
CKINVDCx20_ASAP7_75t_R g764 ( .A(n_320), .Y(n_764) );
INVx1_ASAP7_75t_L g1020 ( .A(n_322), .Y(n_1020) );
CKINVDCx20_ASAP7_75t_R g611 ( .A(n_324), .Y(n_611) );
CKINVDCx20_ASAP7_75t_R g1032 ( .A(n_325), .Y(n_1032) );
INVx1_ASAP7_75t_L g948 ( .A(n_327), .Y(n_948) );
NAND2xp5_ASAP7_75t_L g578 ( .A(n_330), .B(n_579), .Y(n_578) );
CKINVDCx20_ASAP7_75t_R g944 ( .A(n_334), .Y(n_944) );
INVx1_ASAP7_75t_L g412 ( .A(n_338), .Y(n_412) );
CKINVDCx20_ASAP7_75t_R g653 ( .A(n_342), .Y(n_653) );
CKINVDCx20_ASAP7_75t_R g606 ( .A(n_344), .Y(n_606) );
CKINVDCx20_ASAP7_75t_R g433 ( .A(n_345), .Y(n_433) );
CKINVDCx20_ASAP7_75t_R g547 ( .A(n_347), .Y(n_547) );
CKINVDCx20_ASAP7_75t_R g351 ( .A(n_352), .Y(n_351) );
CKINVDCx20_ASAP7_75t_R g352 ( .A(n_353), .Y(n_352) );
HB1xp67_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
AND2x4_ASAP7_75t_L g354 ( .A(n_355), .B(n_357), .Y(n_354) );
HB1xp67_ASAP7_75t_L g987 ( .A(n_356), .Y(n_987) );
OAI21xp5_ASAP7_75t_L g1018 ( .A1(n_357), .A2(n_986), .B(n_1019), .Y(n_1018) );
AND2x2_ASAP7_75t_L g357 ( .A(n_358), .B(n_359), .Y(n_357) );
AOI221xp5_ASAP7_75t_L g360 ( .A1(n_361), .A2(n_627), .B1(n_981), .B2(n_982), .C(n_983), .Y(n_360) );
INVx1_ASAP7_75t_L g982 ( .A(n_361), .Y(n_982) );
AOI22xp5_ASAP7_75t_L g361 ( .A1(n_362), .A2(n_499), .B1(n_625), .B2(n_626), .Y(n_361) );
INVx1_ASAP7_75t_L g625 ( .A(n_362), .Y(n_625) );
OAI22xp5_ASAP7_75t_L g362 ( .A1(n_363), .A2(n_455), .B1(n_497), .B2(n_498), .Y(n_362) );
INVx1_ASAP7_75t_L g497 ( .A(n_363), .Y(n_497) );
INVx1_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
INVx2_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
INVx1_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
AND4x1_ASAP7_75t_L g367 ( .A(n_368), .B(n_401), .C(n_421), .D(n_441), .Y(n_367) );
INVx1_ASAP7_75t_SL g947 ( .A(n_369), .Y(n_947) );
BUFx6f_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
BUFx3_ASAP7_75t_L g657 ( .A(n_370), .Y(n_657) );
BUFx3_ASAP7_75t_L g892 ( .A(n_370), .Y(n_892) );
BUFx6f_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
INVx2_ASAP7_75t_L g466 ( .A(n_371), .Y(n_466) );
BUFx2_ASAP7_75t_SL g856 ( .A(n_371), .Y(n_856) );
BUFx2_ASAP7_75t_SL g970 ( .A(n_371), .Y(n_970) );
AND2x2_ASAP7_75t_L g371 ( .A(n_372), .B(n_381), .Y(n_371) );
AND2x6_ASAP7_75t_L g388 ( .A(n_372), .B(n_389), .Y(n_388) );
AND2x4_ASAP7_75t_L g404 ( .A(n_372), .B(n_405), .Y(n_404) );
AND2x6_ASAP7_75t_L g443 ( .A(n_372), .B(n_438), .Y(n_443) );
AND2x2_ASAP7_75t_L g372 ( .A(n_373), .B(n_378), .Y(n_372) );
AND2x2_ASAP7_75t_L g395 ( .A(n_373), .B(n_379), .Y(n_395) );
INVx2_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
NAND2xp5_ASAP7_75t_L g400 ( .A(n_374), .B(n_379), .Y(n_400) );
AND2x2_ASAP7_75t_L g409 ( .A(n_374), .B(n_410), .Y(n_409) );
AND2x2_ASAP7_75t_L g431 ( .A(n_374), .B(n_383), .Y(n_431) );
INVx1_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
INVx1_ASAP7_75t_L g380 ( .A(n_377), .Y(n_380) );
INVx1_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
INVx1_ASAP7_75t_L g410 ( .A(n_379), .Y(n_410) );
INVx1_ASAP7_75t_L g449 ( .A(n_379), .Y(n_449) );
AND2x4_ASAP7_75t_L g394 ( .A(n_381), .B(n_395), .Y(n_394) );
AND2x4_ASAP7_75t_L g398 ( .A(n_381), .B(n_399), .Y(n_398) );
AND2x2_ASAP7_75t_L g408 ( .A(n_381), .B(n_409), .Y(n_408) );
NAND2xp5_ASAP7_75t_L g823 ( .A(n_381), .B(n_409), .Y(n_823) );
AND2x2_ASAP7_75t_L g381 ( .A(n_382), .B(n_384), .Y(n_381) );
OR2x2_ASAP7_75t_L g390 ( .A(n_382), .B(n_385), .Y(n_390) );
AND2x2_ASAP7_75t_L g405 ( .A(n_382), .B(n_385), .Y(n_405) );
INVx2_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
AND2x2_ASAP7_75t_L g438 ( .A(n_383), .B(n_385), .Y(n_438) );
INVx1_ASAP7_75t_L g432 ( .A(n_384), .Y(n_432) );
AND2x2_ASAP7_75t_L g448 ( .A(n_384), .B(n_449), .Y(n_448) );
INVx2_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
INVx1_ASAP7_75t_L g420 ( .A(n_385), .Y(n_420) );
INVx1_ASAP7_75t_L g943 ( .A(n_386), .Y(n_943) );
INVx3_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
INVx4_ASAP7_75t_L g469 ( .A(n_387), .Y(n_469) );
INVx2_ASAP7_75t_SL g698 ( .A(n_387), .Y(n_698) );
INVx11_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
INVx11_ASAP7_75t_L g540 ( .A(n_388), .Y(n_540) );
AND2x4_ASAP7_75t_L g425 ( .A(n_389), .B(n_395), .Y(n_425) );
INVx2_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
OR2x2_ASAP7_75t_L g485 ( .A(n_390), .B(n_486), .Y(n_485) );
BUFx2_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
BUFx3_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
BUFx6f_ASAP7_75t_L g472 ( .A(n_394), .Y(n_472) );
INVx2_ASAP7_75t_L g659 ( .A(n_394), .Y(n_659) );
BUFx3_ASAP7_75t_L g722 ( .A(n_394), .Y(n_722) );
BUFx3_ASAP7_75t_L g743 ( .A(n_394), .Y(n_743) );
AND2x6_ASAP7_75t_L g427 ( .A(n_395), .B(n_405), .Y(n_427) );
NAND2x1p5_ASAP7_75t_L g478 ( .A(n_395), .B(n_405), .Y(n_478) );
INVx1_ASAP7_75t_L g486 ( .A(n_395), .Y(n_486) );
HB1xp67_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
INVx2_ASAP7_75t_L g896 ( .A(n_397), .Y(n_896) );
BUFx3_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
BUFx3_ASAP7_75t_L g470 ( .A(n_398), .Y(n_470) );
BUFx2_ASAP7_75t_SL g529 ( .A(n_398), .Y(n_529) );
BUFx2_ASAP7_75t_L g594 ( .A(n_398), .Y(n_594) );
BUFx3_ASAP7_75t_L g712 ( .A(n_398), .Y(n_712) );
INVx1_ASAP7_75t_L g819 ( .A(n_398), .Y(n_819) );
BUFx3_ASAP7_75t_L g846 ( .A(n_398), .Y(n_846) );
BUFx2_ASAP7_75t_SL g968 ( .A(n_398), .Y(n_968) );
AND2x2_ASAP7_75t_L g473 ( .A(n_399), .B(n_432), .Y(n_473) );
INVx1_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
OR2x6_ASAP7_75t_L g419 ( .A(n_400), .B(n_420), .Y(n_419) );
INVx2_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
INVx3_ASAP7_75t_L g542 ( .A(n_403), .Y(n_542) );
INVx2_ASAP7_75t_L g589 ( .A(n_403), .Y(n_589) );
INVx2_ASAP7_75t_L g667 ( .A(n_403), .Y(n_667) );
OAI22xp5_ASAP7_75t_SL g813 ( .A1(n_403), .A2(n_466), .B1(n_814), .B2(n_815), .Y(n_813) );
OAI22xp5_ASAP7_75t_L g941 ( .A1(n_403), .A2(n_942), .B1(n_943), .B2(n_944), .Y(n_941) );
INVx6_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
BUFx3_ASAP7_75t_L g750 ( .A(n_404), .Y(n_750) );
BUFx3_ASAP7_75t_L g787 ( .A(n_404), .Y(n_787) );
NAND2xp5_ASAP7_75t_SL g414 ( .A(n_405), .B(n_409), .Y(n_414) );
AND2x2_ASAP7_75t_L g463 ( .A(n_405), .B(n_409), .Y(n_463) );
BUFx2_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
INVx1_ASAP7_75t_L g888 ( .A(n_407), .Y(n_888) );
BUFx3_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
BUFx3_ASAP7_75t_L g528 ( .A(n_408), .Y(n_528) );
BUFx3_ASAP7_75t_L g562 ( .A(n_408), .Y(n_562) );
BUFx3_ASAP7_75t_L g702 ( .A(n_408), .Y(n_702) );
INVx1_ASAP7_75t_L g440 ( .A(n_410), .Y(n_440) );
OAI22xp5_ASAP7_75t_L g411 ( .A1(n_412), .A2(n_413), .B1(n_415), .B2(n_416), .Y(n_411) );
BUFx2_ASAP7_75t_R g413 ( .A(n_414), .Y(n_413) );
OAI22xp5_ASAP7_75t_L g817 ( .A1(n_414), .A2(n_818), .B1(n_819), .B2(n_820), .Y(n_817) );
CKINVDCx20_ASAP7_75t_R g416 ( .A(n_417), .Y(n_416) );
BUFx4f_ASAP7_75t_SL g417 ( .A(n_418), .Y(n_417) );
BUFx2_ASAP7_75t_L g534 ( .A(n_418), .Y(n_534) );
BUFx2_ASAP7_75t_L g746 ( .A(n_418), .Y(n_746) );
BUFx2_ASAP7_75t_L g1004 ( .A(n_418), .Y(n_1004) );
INVx6_ASAP7_75t_SL g418 ( .A(n_419), .Y(n_418) );
INVx1_ASAP7_75t_SL g591 ( .A(n_419), .Y(n_591) );
INVx1_ASAP7_75t_SL g848 ( .A(n_419), .Y(n_848) );
INVx1_ASAP7_75t_L g1038 ( .A(n_419), .Y(n_1038) );
INVx1_ASAP7_75t_L g557 ( .A(n_420), .Y(n_557) );
BUFx6f_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
INVx5_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
INVx2_ASAP7_75t_L g579 ( .A(n_424), .Y(n_579) );
INVx2_ASAP7_75t_L g716 ( .A(n_424), .Y(n_716) );
INVx2_ASAP7_75t_L g739 ( .A(n_424), .Y(n_739) );
INVx4_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
INVx1_ASAP7_75t_L g882 ( .A(n_426), .Y(n_882) );
BUFx4f_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
BUFx2_ASAP7_75t_L g775 ( .A(n_427), .Y(n_775) );
INVx1_ASAP7_75t_SL g842 ( .A(n_427), .Y(n_842) );
BUFx2_ASAP7_75t_L g962 ( .A(n_427), .Y(n_962) );
OAI22xp5_ASAP7_75t_L g428 ( .A1(n_429), .A2(n_430), .B1(n_433), .B2(n_434), .Y(n_428) );
INVx4_ASAP7_75t_L g481 ( .A(n_430), .Y(n_481) );
OAI22xp5_ASAP7_75t_L g520 ( .A1(n_430), .A2(n_521), .B1(n_522), .B2(n_523), .Y(n_520) );
HB1xp67_ASAP7_75t_L g612 ( .A(n_430), .Y(n_612) );
OAI22xp5_ASAP7_75t_L g802 ( .A1(n_430), .A2(n_515), .B1(n_803), .B2(n_804), .Y(n_802) );
NAND2x1p5_ASAP7_75t_L g430 ( .A(n_431), .B(n_432), .Y(n_430) );
AND2x4_ASAP7_75t_L g447 ( .A(n_431), .B(n_448), .Y(n_447) );
AND2x4_ASAP7_75t_L g452 ( .A(n_431), .B(n_453), .Y(n_452) );
AND2x4_ASAP7_75t_L g556 ( .A(n_431), .B(n_557), .Y(n_556) );
OAI22xp5_ASAP7_75t_L g688 ( .A1(n_434), .A2(n_612), .B1(n_689), .B2(n_690), .Y(n_688) );
OAI22xp5_ASAP7_75t_L g1031 ( .A1(n_434), .A2(n_480), .B1(n_1032), .B2(n_1033), .Y(n_1031) );
INVx2_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
CKINVDCx16_ASAP7_75t_R g435 ( .A(n_436), .Y(n_435) );
BUFx2_ASAP7_75t_L g523 ( .A(n_436), .Y(n_523) );
OAI22xp5_ASAP7_75t_L g910 ( .A1(n_436), .A2(n_911), .B1(n_912), .B2(n_913), .Y(n_910) );
OR2x6_ASAP7_75t_L g436 ( .A(n_437), .B(n_439), .Y(n_436) );
INVx1_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
AND2x4_ASAP7_75t_L g491 ( .A(n_438), .B(n_440), .Y(n_491) );
INVx1_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
INVx2_ASAP7_75t_SL g517 ( .A(n_442), .Y(n_517) );
INVx2_ASAP7_75t_L g833 ( .A(n_442), .Y(n_833) );
BUFx6f_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
INVx4_ASAP7_75t_L g493 ( .A(n_443), .Y(n_493) );
INVx2_ASAP7_75t_L g548 ( .A(n_443), .Y(n_548) );
INVx2_ASAP7_75t_SL g807 ( .A(n_443), .Y(n_807) );
INVx2_ASAP7_75t_L g863 ( .A(n_443), .Y(n_863) );
BUFx3_ASAP7_75t_L g907 ( .A(n_443), .Y(n_907) );
INVx3_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
OAI222xp33_ASAP7_75t_L g683 ( .A1(n_445), .A2(n_517), .B1(n_684), .B2(n_685), .C1(n_686), .C2(n_687), .Y(n_683) );
OAI22xp5_ASAP7_75t_L g805 ( .A1(n_445), .A2(n_806), .B1(n_807), .B2(n_808), .Y(n_805) );
INVx4_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
INVx2_ASAP7_75t_L g495 ( .A(n_446), .Y(n_495) );
BUFx2_ASAP7_75t_L g836 ( .A(n_446), .Y(n_836) );
BUFx6f_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
BUFx4f_ASAP7_75t_SL g554 ( .A(n_447), .Y(n_554) );
BUFx6f_ASAP7_75t_L g582 ( .A(n_447), .Y(n_582) );
BUFx6f_ASAP7_75t_L g649 ( .A(n_447), .Y(n_649) );
BUFx2_ASAP7_75t_L g909 ( .A(n_447), .Y(n_909) );
INVx1_ASAP7_75t_L g453 ( .A(n_449), .Y(n_453) );
INVx2_ASAP7_75t_L g652 ( .A(n_450), .Y(n_652) );
BUFx3_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
INVx2_ASAP7_75t_L g686 ( .A(n_451), .Y(n_686) );
BUFx6f_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
BUFx6f_ASAP7_75t_L g489 ( .A(n_452), .Y(n_489) );
BUFx12f_ASAP7_75t_L g550 ( .A(n_452), .Y(n_550) );
INVx1_ASAP7_75t_SL g498 ( .A(n_455), .Y(n_498) );
HB1xp67_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
XNOR2xp5_ASAP7_75t_L g456 ( .A(n_457), .B(n_458), .Y(n_456) );
NAND3x1_ASAP7_75t_SL g458 ( .A(n_459), .B(n_467), .C(n_474), .Y(n_458) );
AND2x2_ASAP7_75t_L g459 ( .A(n_460), .B(n_464), .Y(n_459) );
INVx3_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
INVx4_ASAP7_75t_L g533 ( .A(n_462), .Y(n_533) );
INVx5_ASAP7_75t_L g567 ( .A(n_462), .Y(n_567) );
INVx2_ASAP7_75t_L g724 ( .A(n_462), .Y(n_724) );
INVx1_ASAP7_75t_L g745 ( .A(n_462), .Y(n_745) );
INVx8_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
INVx3_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
INVx3_ASAP7_75t_L g564 ( .A(n_466), .Y(n_564) );
AND2x2_ASAP7_75t_L g467 ( .A(n_468), .B(n_471), .Y(n_467) );
BUFx2_ASAP7_75t_L g671 ( .A(n_470), .Y(n_671) );
INVx4_ASAP7_75t_L g621 ( .A(n_472), .Y(n_621) );
NOR3xp33_ASAP7_75t_L g474 ( .A(n_475), .B(n_483), .C(n_492), .Y(n_474) );
OAI22xp5_ASAP7_75t_SL g475 ( .A1(n_476), .A2(n_479), .B1(n_480), .B2(n_482), .Y(n_475) );
OAI22xp5_ASAP7_75t_L g901 ( .A1(n_476), .A2(n_637), .B1(n_902), .B2(n_903), .Y(n_901) );
INVx2_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
INVx1_ASAP7_75t_L g477 ( .A(n_478), .Y(n_477) );
BUFx3_ASAP7_75t_L g515 ( .A(n_478), .Y(n_515) );
INVx3_ASAP7_75t_SL g480 ( .A(n_481), .Y(n_480) );
INVx2_ASAP7_75t_L g912 ( .A(n_481), .Y(n_912) );
OAI21xp5_ASAP7_75t_SL g483 ( .A1(n_484), .A2(n_487), .B(n_488), .Y(n_483) );
BUFx6f_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
INVx2_ASAP7_75t_L g512 ( .A(n_485), .Y(n_512) );
OAI21xp5_ASAP7_75t_L g799 ( .A1(n_485), .A2(n_800), .B(n_801), .Y(n_799) );
INVx1_ASAP7_75t_SL g646 ( .A(n_490), .Y(n_646) );
BUFx6f_ASAP7_75t_L g490 ( .A(n_491), .Y(n_490) );
BUFx2_ASAP7_75t_SL g551 ( .A(n_491), .Y(n_551) );
BUFx2_ASAP7_75t_SL g586 ( .A(n_491), .Y(n_586) );
BUFx3_ASAP7_75t_L g719 ( .A(n_491), .Y(n_719) );
OAI22xp5_ASAP7_75t_SL g492 ( .A1(n_493), .A2(n_494), .B1(n_495), .B2(n_496), .Y(n_492) );
INVx4_ASAP7_75t_L g726 ( .A(n_493), .Y(n_726) );
BUFx2_ASAP7_75t_L g1029 ( .A(n_493), .Y(n_1029) );
INVx1_ASAP7_75t_L g626 ( .A(n_499), .Y(n_626) );
AOI22xp5_ASAP7_75t_L g499 ( .A1(n_500), .A2(n_501), .B1(n_571), .B2(n_624), .Y(n_499) );
INVx1_ASAP7_75t_L g500 ( .A(n_501), .Y(n_500) );
BUFx2_ASAP7_75t_L g501 ( .A(n_502), .Y(n_501) );
AO22x1_ASAP7_75t_L g502 ( .A1(n_503), .A2(n_504), .B1(n_543), .B2(n_570), .Y(n_502) );
INVx1_ASAP7_75t_L g503 ( .A(n_504), .Y(n_503) );
INVx1_ASAP7_75t_SL g506 ( .A(n_507), .Y(n_506) );
AND2x2_ASAP7_75t_L g507 ( .A(n_508), .B(n_524), .Y(n_507) );
NOR3xp33_ASAP7_75t_L g508 ( .A(n_509), .B(n_516), .C(n_520), .Y(n_508) );
OAI22xp5_ASAP7_75t_L g509 ( .A1(n_510), .A2(n_511), .B1(n_513), .B2(n_514), .Y(n_509) );
INVx2_ASAP7_75t_L g511 ( .A(n_512), .Y(n_511) );
INVx1_ASAP7_75t_SL g603 ( .A(n_512), .Y(n_603) );
INVx2_ASAP7_75t_L g637 ( .A(n_512), .Y(n_637) );
BUFx3_ASAP7_75t_L g514 ( .A(n_515), .Y(n_514) );
OAI22xp5_ASAP7_75t_L g601 ( .A1(n_515), .A2(n_602), .B1(n_603), .B2(n_604), .Y(n_601) );
INVx2_ASAP7_75t_L g640 ( .A(n_515), .Y(n_640) );
OAI22xp5_ASAP7_75t_L g680 ( .A1(n_515), .A2(n_637), .B1(n_681), .B2(n_682), .Y(n_680) );
OA211x2_ASAP7_75t_L g763 ( .A1(n_515), .A2(n_764), .B(n_765), .C(n_766), .Y(n_763) );
OAI21xp33_ASAP7_75t_SL g516 ( .A1(n_517), .A2(n_518), .B(n_519), .Y(n_516) );
OAI21xp33_ASAP7_75t_L g605 ( .A1(n_517), .A2(n_606), .B(n_607), .Y(n_605) );
NOR2xp33_ASAP7_75t_L g524 ( .A(n_525), .B(n_535), .Y(n_524) );
NAND2xp5_ASAP7_75t_L g525 ( .A(n_526), .B(n_530), .Y(n_525) );
BUFx4f_ASAP7_75t_SL g527 ( .A(n_528), .Y(n_527) );
INVx1_ASAP7_75t_L g670 ( .A(n_528), .Y(n_670) );
INVx3_ASAP7_75t_L g531 ( .A(n_532), .Y(n_531) );
INVx2_ASAP7_75t_L g532 ( .A(n_533), .Y(n_532) );
BUFx2_ASAP7_75t_L g890 ( .A(n_533), .Y(n_890) );
NAND2xp5_ASAP7_75t_L g535 ( .A(n_536), .B(n_541), .Y(n_535) );
INVx2_ASAP7_75t_L g537 ( .A(n_538), .Y(n_537) );
INVx1_ASAP7_75t_L g538 ( .A(n_539), .Y(n_538) );
INVx5_ASAP7_75t_SL g539 ( .A(n_540), .Y(n_539) );
INVx2_ASAP7_75t_SL g666 ( .A(n_540), .Y(n_666) );
NOR2xp33_ASAP7_75t_L g824 ( .A(n_540), .B(n_825), .Y(n_824) );
INVx4_ASAP7_75t_L g893 ( .A(n_540), .Y(n_893) );
INVx2_ASAP7_75t_L g967 ( .A(n_540), .Y(n_967) );
INVx3_ASAP7_75t_SL g570 ( .A(n_543), .Y(n_570) );
OAI22xp5_ASAP7_75t_L g596 ( .A1(n_543), .A2(n_570), .B1(n_597), .B2(n_598), .Y(n_596) );
XOR2x2_ASAP7_75t_L g543 ( .A(n_544), .B(n_569), .Y(n_543) );
NAND2xp5_ASAP7_75t_SL g544 ( .A(n_545), .B(n_559), .Y(n_544) );
NOR2xp33_ASAP7_75t_L g545 ( .A(n_546), .B(n_552), .Y(n_545) );
OAI21xp5_ASAP7_75t_L g546 ( .A1(n_547), .A2(n_548), .B(n_549), .Y(n_546) );
OAI21xp5_ASAP7_75t_L g583 ( .A1(n_548), .A2(n_584), .B(n_585), .Y(n_583) );
OAI222xp33_ASAP7_75t_L g647 ( .A1(n_548), .A2(n_648), .B1(n_650), .B2(n_651), .C1(n_652), .C2(n_653), .Y(n_647) );
OAI21xp5_ASAP7_75t_SL g733 ( .A1(n_548), .A2(n_734), .B(n_735), .Y(n_733) );
OAI21xp5_ASAP7_75t_SL g778 ( .A1(n_548), .A2(n_779), .B(n_780), .Y(n_778) );
OAI21xp5_ASAP7_75t_SL g955 ( .A1(n_548), .A2(n_956), .B(n_957), .Y(n_955) );
INVx2_ASAP7_75t_L g728 ( .A(n_550), .Y(n_728) );
BUFx4f_ASAP7_75t_SL g959 ( .A(n_550), .Y(n_959) );
NAND2xp5_ASAP7_75t_L g552 ( .A(n_553), .B(n_558), .Y(n_552) );
INVx1_ASAP7_75t_L g610 ( .A(n_554), .Y(n_610) );
BUFx3_ASAP7_75t_L g555 ( .A(n_556), .Y(n_555) );
INVx1_ASAP7_75t_L g644 ( .A(n_556), .Y(n_644) );
BUFx2_ASAP7_75t_L g718 ( .A(n_556), .Y(n_718) );
BUFx2_ASAP7_75t_L g839 ( .A(n_556), .Y(n_839) );
NOR2xp33_ASAP7_75t_L g559 ( .A(n_560), .B(n_565), .Y(n_559) );
NAND2xp5_ASAP7_75t_L g560 ( .A(n_561), .B(n_563), .Y(n_560) );
NAND2xp5_ASAP7_75t_L g565 ( .A(n_566), .B(n_568), .Y(n_565) );
BUFx2_ASAP7_75t_L g661 ( .A(n_567), .Y(n_661) );
BUFx6f_ASAP7_75t_L g695 ( .A(n_567), .Y(n_695) );
INVx2_ASAP7_75t_L g624 ( .A(n_571), .Y(n_624) );
HB1xp67_ASAP7_75t_L g571 ( .A(n_572), .Y(n_571) );
OA22x2_ASAP7_75t_L g572 ( .A1(n_573), .A2(n_574), .B1(n_596), .B2(n_623), .Y(n_572) );
INVx1_ASAP7_75t_L g573 ( .A(n_574), .Y(n_573) );
XOR2x2_ASAP7_75t_L g574 ( .A(n_575), .B(n_595), .Y(n_574) );
NAND4xp75_ASAP7_75t_SL g575 ( .A(n_576), .B(n_587), .C(n_592), .D(n_593), .Y(n_575) );
NOR2xp67_ASAP7_75t_SL g576 ( .A(n_577), .B(n_583), .Y(n_576) );
NAND3xp33_ASAP7_75t_L g577 ( .A(n_578), .B(n_580), .C(n_581), .Y(n_577) );
INVx1_ASAP7_75t_L g934 ( .A(n_582), .Y(n_934) );
BUFx6f_ASAP7_75t_L g958 ( .A(n_582), .Y(n_958) );
AND2x2_ASAP7_75t_L g587 ( .A(n_588), .B(n_590), .Y(n_587) );
INVx1_ASAP7_75t_L g623 ( .A(n_596), .Y(n_623) );
INVx1_ASAP7_75t_SL g597 ( .A(n_598), .Y(n_597) );
XNOR2x1_ASAP7_75t_L g598 ( .A(n_599), .B(n_622), .Y(n_598) );
AND2x2_ASAP7_75t_L g599 ( .A(n_600), .B(n_613), .Y(n_599) );
NOR3xp33_ASAP7_75t_L g600 ( .A(n_601), .B(n_605), .C(n_608), .Y(n_600) );
OAI22xp5_ASAP7_75t_L g1024 ( .A1(n_603), .A2(n_639), .B1(n_1025), .B2(n_1026), .Y(n_1024) );
OAI22xp5_ASAP7_75t_L g608 ( .A1(n_609), .A2(n_610), .B1(n_611), .B2(n_612), .Y(n_608) );
NOR2xp33_ASAP7_75t_L g613 ( .A(n_614), .B(n_617), .Y(n_613) );
NAND2xp5_ASAP7_75t_L g614 ( .A(n_615), .B(n_616), .Y(n_614) );
NAND2xp5_ASAP7_75t_L g617 ( .A(n_618), .B(n_619), .Y(n_617) );
INVx3_ASAP7_75t_L g620 ( .A(n_621), .Y(n_620) );
INVx4_ASAP7_75t_L g1041 ( .A(n_621), .Y(n_1041) );
INVx1_ASAP7_75t_L g981 ( .A(n_627), .Y(n_981) );
AOI22xp5_ASAP7_75t_L g627 ( .A1(n_628), .A2(n_792), .B1(n_979), .B2(n_980), .Y(n_627) );
INVx1_ASAP7_75t_L g980 ( .A(n_628), .Y(n_980) );
OAI22xp5_ASAP7_75t_SL g628 ( .A1(n_629), .A2(n_630), .B1(n_753), .B2(n_754), .Y(n_628) );
INVx1_ASAP7_75t_L g629 ( .A(n_630), .Y(n_629) );
XNOR2x1_ASAP7_75t_L g630 ( .A(n_631), .B(n_674), .Y(n_630) );
INVx1_ASAP7_75t_L g631 ( .A(n_632), .Y(n_631) );
INVx1_ASAP7_75t_L g632 ( .A(n_633), .Y(n_632) );
INVx1_ASAP7_75t_SL g673 ( .A(n_634), .Y(n_673) );
AND2x2_ASAP7_75t_L g634 ( .A(n_635), .B(n_654), .Y(n_634) );
NOR2xp33_ASAP7_75t_SL g635 ( .A(n_636), .B(n_647), .Y(n_635) );
OAI221xp5_ASAP7_75t_L g636 ( .A1(n_637), .A2(n_638), .B1(n_639), .B2(n_641), .C(n_642), .Y(n_636) );
OAI211xp5_ASAP7_75t_L g928 ( .A1(n_639), .A2(n_929), .B(n_930), .C(n_931), .Y(n_928) );
INVx2_ASAP7_75t_L g639 ( .A(n_640), .Y(n_639) );
INVx1_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
INVx2_ASAP7_75t_L g645 ( .A(n_646), .Y(n_645) );
CKINVDCx20_ASAP7_75t_R g648 ( .A(n_649), .Y(n_648) );
NOR2xp33_ASAP7_75t_L g654 ( .A(n_655), .B(n_662), .Y(n_654) );
NAND2xp5_ASAP7_75t_L g655 ( .A(n_656), .B(n_660), .Y(n_655) );
INVx1_ASAP7_75t_L g658 ( .A(n_659), .Y(n_658) );
OAI21xp5_ASAP7_75t_SL g810 ( .A1(n_659), .A2(n_811), .B(n_812), .Y(n_810) );
INVx2_ASAP7_75t_L g845 ( .A(n_659), .Y(n_845) );
NAND2xp5_ASAP7_75t_SL g662 ( .A(n_663), .B(n_668), .Y(n_662) );
INVx1_ASAP7_75t_L g664 ( .A(n_665), .Y(n_664) );
INVx1_ASAP7_75t_L g665 ( .A(n_666), .Y(n_665) );
INVx1_ASAP7_75t_L g669 ( .A(n_670), .Y(n_669) );
BUFx3_ASAP7_75t_L g674 ( .A(n_675), .Y(n_674) );
AOI22xp5_ASAP7_75t_L g675 ( .A1(n_676), .A2(n_677), .B1(n_705), .B2(n_706), .Y(n_675) );
INVx1_ASAP7_75t_L g676 ( .A(n_677), .Y(n_676) );
INVx1_ASAP7_75t_L g704 ( .A(n_678), .Y(n_704) );
AND2x2_ASAP7_75t_L g678 ( .A(n_679), .B(n_691), .Y(n_678) );
NOR3xp33_ASAP7_75t_L g679 ( .A(n_680), .B(n_683), .C(n_688), .Y(n_679) );
NOR2xp33_ASAP7_75t_L g691 ( .A(n_692), .B(n_696), .Y(n_691) );
NAND2xp5_ASAP7_75t_L g692 ( .A(n_693), .B(n_694), .Y(n_692) );
NAND2xp5_ASAP7_75t_SL g696 ( .A(n_697), .B(n_699), .Y(n_696) );
INVx1_ASAP7_75t_L g700 ( .A(n_701), .Y(n_700) );
INVx1_ASAP7_75t_L g701 ( .A(n_702), .Y(n_701) );
INVx1_ASAP7_75t_L g705 ( .A(n_706), .Y(n_705) );
AO22x2_ASAP7_75t_L g706 ( .A1(n_707), .A2(n_708), .B1(n_730), .B2(n_752), .Y(n_706) );
INVx2_ASAP7_75t_SL g707 ( .A(n_708), .Y(n_707) );
XOR2x2_ASAP7_75t_L g708 ( .A(n_709), .B(n_729), .Y(n_708) );
NAND4xp75_ASAP7_75t_L g709 ( .A(n_710), .B(n_714), .C(n_720), .D(n_725), .Y(n_709) );
AND2x2_ASAP7_75t_L g710 ( .A(n_711), .B(n_713), .Y(n_710) );
AND2x2_ASAP7_75t_SL g714 ( .A(n_715), .B(n_717), .Y(n_714) );
AND2x2_ASAP7_75t_L g720 ( .A(n_721), .B(n_723), .Y(n_720) );
INVx1_ASAP7_75t_L g936 ( .A(n_727), .Y(n_936) );
INVx3_ASAP7_75t_L g727 ( .A(n_728), .Y(n_727) );
INVx4_ASAP7_75t_SL g752 ( .A(n_730), .Y(n_752) );
XOR2x2_ASAP7_75t_L g730 ( .A(n_731), .B(n_751), .Y(n_730) );
NAND3x1_ASAP7_75t_L g731 ( .A(n_732), .B(n_741), .C(n_747), .Y(n_731) );
NOR2xp33_ASAP7_75t_L g732 ( .A(n_733), .B(n_736), .Y(n_732) );
NAND3xp33_ASAP7_75t_L g736 ( .A(n_737), .B(n_738), .C(n_740), .Y(n_736) );
AND2x2_ASAP7_75t_L g741 ( .A(n_742), .B(n_744), .Y(n_741) );
AND2x2_ASAP7_75t_L g747 ( .A(n_748), .B(n_749), .Y(n_747) );
INVx1_ASAP7_75t_L g753 ( .A(n_754), .Y(n_753) );
OAI22xp5_ASAP7_75t_SL g754 ( .A1(n_755), .A2(n_769), .B1(n_790), .B2(n_791), .Y(n_754) );
INVx2_ASAP7_75t_SL g790 ( .A(n_755), .Y(n_790) );
XOR2x2_ASAP7_75t_L g755 ( .A(n_756), .B(n_768), .Y(n_755) );
NAND4xp75_ASAP7_75t_L g756 ( .A(n_757), .B(n_760), .C(n_763), .D(n_767), .Y(n_756) );
AND2x2_ASAP7_75t_L g757 ( .A(n_758), .B(n_759), .Y(n_757) );
AND2x2_ASAP7_75t_L g760 ( .A(n_761), .B(n_762), .Y(n_760) );
INVx1_ASAP7_75t_SL g791 ( .A(n_769), .Y(n_791) );
INVx1_ASAP7_75t_L g769 ( .A(n_770), .Y(n_769) );
XOR2x2_ASAP7_75t_SL g770 ( .A(n_771), .B(n_789), .Y(n_770) );
NAND2x1p5_ASAP7_75t_L g771 ( .A(n_772), .B(n_781), .Y(n_771) );
NOR2xp33_ASAP7_75t_L g772 ( .A(n_773), .B(n_778), .Y(n_772) );
NAND3xp33_ASAP7_75t_L g773 ( .A(n_774), .B(n_776), .C(n_777), .Y(n_773) );
NOR2x1_ASAP7_75t_L g781 ( .A(n_782), .B(n_785), .Y(n_781) );
NAND2xp5_ASAP7_75t_L g782 ( .A(n_783), .B(n_784), .Y(n_782) );
NAND2xp5_ASAP7_75t_L g785 ( .A(n_786), .B(n_788), .Y(n_785) );
INVx1_ASAP7_75t_L g979 ( .A(n_792), .Y(n_979) );
XOR2xp5_ASAP7_75t_L g792 ( .A(n_793), .B(n_869), .Y(n_792) );
INVx1_ASAP7_75t_L g793 ( .A(n_794), .Y(n_793) );
XNOR2xp5_ASAP7_75t_L g794 ( .A(n_795), .B(n_827), .Y(n_794) );
BUFx2_ASAP7_75t_L g795 ( .A(n_796), .Y(n_795) );
XNOR2x1_ASAP7_75t_L g796 ( .A(n_797), .B(n_826), .Y(n_796) );
AND3x2_ASAP7_75t_L g797 ( .A(n_798), .B(n_809), .C(n_816), .Y(n_797) );
NOR3xp33_ASAP7_75t_L g798 ( .A(n_799), .B(n_802), .C(n_805), .Y(n_798) );
NOR2xp33_ASAP7_75t_L g809 ( .A(n_810), .B(n_813), .Y(n_809) );
NOR3xp33_ASAP7_75t_L g816 ( .A(n_817), .B(n_821), .C(n_824), .Y(n_816) );
NOR2xp33_ASAP7_75t_L g821 ( .A(n_822), .B(n_823), .Y(n_821) );
INVx1_ASAP7_75t_L g950 ( .A(n_823), .Y(n_950) );
XOR2x2_ASAP7_75t_L g827 ( .A(n_828), .B(n_852), .Y(n_827) );
XNOR2xp5_ASAP7_75t_L g828 ( .A(n_829), .B(n_830), .Y(n_828) );
NAND3xp33_ASAP7_75t_L g830 ( .A(n_831), .B(n_843), .C(n_849), .Y(n_830) );
NOR2xp33_ASAP7_75t_L g831 ( .A(n_832), .B(n_837), .Y(n_831) );
OAI21xp5_ASAP7_75t_SL g832 ( .A1(n_833), .A2(n_834), .B(n_835), .Y(n_832) );
OAI21xp5_ASAP7_75t_SL g876 ( .A1(n_833), .A2(n_877), .B(n_878), .Y(n_876) );
NAND2xp5_ASAP7_75t_L g837 ( .A(n_838), .B(n_840), .Y(n_837) );
INVx1_ASAP7_75t_SL g841 ( .A(n_842), .Y(n_841) );
AND2x2_ASAP7_75t_L g843 ( .A(n_844), .B(n_847), .Y(n_843) );
AND2x2_ASAP7_75t_L g849 ( .A(n_850), .B(n_851), .Y(n_849) );
XOR2x2_ASAP7_75t_L g852 ( .A(n_853), .B(n_868), .Y(n_852) );
NAND4xp75_ASAP7_75t_SL g853 ( .A(n_854), .B(n_855), .C(n_857), .D(n_860), .Y(n_853) );
AND2x2_ASAP7_75t_L g857 ( .A(n_858), .B(n_859), .Y(n_857) );
NOR2xp33_ASAP7_75t_L g860 ( .A(n_861), .B(n_865), .Y(n_860) );
OAI21xp5_ASAP7_75t_L g861 ( .A1(n_862), .A2(n_863), .B(n_864), .Y(n_861) );
NAND2xp5_ASAP7_75t_L g865 ( .A(n_866), .B(n_867), .Y(n_865) );
AOI22xp33_ASAP7_75t_L g869 ( .A1(n_870), .A2(n_921), .B1(n_977), .B2(n_978), .Y(n_869) );
INVx1_ASAP7_75t_L g977 ( .A(n_870), .Y(n_977) );
INVx2_ASAP7_75t_L g870 ( .A(n_871), .Y(n_870) );
AO22x1_ASAP7_75t_L g871 ( .A1(n_872), .A2(n_873), .B1(n_897), .B2(n_898), .Y(n_871) );
INVx1_ASAP7_75t_L g872 ( .A(n_873), .Y(n_872) );
NAND4xp75_ASAP7_75t_SL g874 ( .A(n_875), .B(n_885), .C(n_891), .D(n_894), .Y(n_874) );
NOR2xp67_ASAP7_75t_L g875 ( .A(n_876), .B(n_879), .Y(n_875) );
NAND3xp33_ASAP7_75t_L g879 ( .A(n_880), .B(n_883), .C(n_884), .Y(n_879) );
INVx1_ASAP7_75t_L g881 ( .A(n_882), .Y(n_881) );
AND2x2_ASAP7_75t_L g885 ( .A(n_886), .B(n_889), .Y(n_885) );
INVx2_ASAP7_75t_L g887 ( .A(n_888), .Y(n_887) );
INVx2_ASAP7_75t_L g895 ( .A(n_896), .Y(n_895) );
INVx2_ASAP7_75t_L g897 ( .A(n_898), .Y(n_897) );
XNOR2x2_ASAP7_75t_L g951 ( .A(n_898), .B(n_952), .Y(n_951) );
INVx1_ASAP7_75t_SL g919 ( .A(n_899), .Y(n_919) );
AND2x2_ASAP7_75t_SL g899 ( .A(n_900), .B(n_914), .Y(n_899) );
NOR3xp33_ASAP7_75t_L g900 ( .A(n_901), .B(n_904), .C(n_910), .Y(n_900) );
OAI21xp33_ASAP7_75t_L g904 ( .A1(n_905), .A2(n_906), .B(n_908), .Y(n_904) );
INVx3_ASAP7_75t_L g906 ( .A(n_907), .Y(n_906) );
AND4x1_ASAP7_75t_L g914 ( .A(n_915), .B(n_916), .C(n_917), .D(n_918), .Y(n_914) );
INVx2_ASAP7_75t_SL g978 ( .A(n_921), .Y(n_978) );
AOI22xp5_ASAP7_75t_L g921 ( .A1(n_922), .A2(n_923), .B1(n_951), .B2(n_976), .Y(n_921) );
INVx1_ASAP7_75t_L g922 ( .A(n_923), .Y(n_922) );
INVx2_ASAP7_75t_L g923 ( .A(n_924), .Y(n_923) );
XNOR2xp5_ASAP7_75t_L g924 ( .A(n_925), .B(n_926), .Y(n_924) );
AND2x2_ASAP7_75t_L g926 ( .A(n_927), .B(n_937), .Y(n_926) );
OAI22xp5_ASAP7_75t_L g932 ( .A1(n_933), .A2(n_934), .B1(n_935), .B2(n_936), .Y(n_932) );
NOR3xp33_ASAP7_75t_L g937 ( .A(n_938), .B(n_941), .C(n_945), .Y(n_937) );
NAND2xp5_ASAP7_75t_L g938 ( .A(n_939), .B(n_940), .Y(n_938) );
OAI22xp5_ASAP7_75t_L g945 ( .A1(n_946), .A2(n_947), .B1(n_948), .B2(n_949), .Y(n_945) );
INVx1_ASAP7_75t_L g949 ( .A(n_950), .Y(n_949) );
INVx2_ASAP7_75t_L g976 ( .A(n_951), .Y(n_976) );
INVx2_ASAP7_75t_SL g974 ( .A(n_953), .Y(n_974) );
AND2x2_ASAP7_75t_L g953 ( .A(n_954), .B(n_964), .Y(n_953) );
NOR2xp33_ASAP7_75t_L g954 ( .A(n_955), .B(n_960), .Y(n_954) );
NAND2xp5_ASAP7_75t_SL g960 ( .A(n_961), .B(n_963), .Y(n_960) );
NOR2xp33_ASAP7_75t_L g964 ( .A(n_965), .B(n_971), .Y(n_964) );
NAND2xp5_ASAP7_75t_L g965 ( .A(n_966), .B(n_969), .Y(n_965) );
NAND2xp5_ASAP7_75t_L g971 ( .A(n_972), .B(n_973), .Y(n_971) );
INVx1_ASAP7_75t_SL g983 ( .A(n_984), .Y(n_983) );
NOR2x1_ASAP7_75t_L g984 ( .A(n_985), .B(n_989), .Y(n_984) );
OR2x2_ASAP7_75t_SL g1045 ( .A(n_985), .B(n_990), .Y(n_1045) );
NAND2xp5_ASAP7_75t_L g985 ( .A(n_986), .B(n_988), .Y(n_985) );
INVx1_ASAP7_75t_L g986 ( .A(n_987), .Y(n_986) );
HB1xp67_ASAP7_75t_L g1013 ( .A(n_987), .Y(n_1013) );
NAND2xp5_ASAP7_75t_L g1019 ( .A(n_987), .B(n_1016), .Y(n_1019) );
CKINVDCx16_ASAP7_75t_R g1016 ( .A(n_988), .Y(n_1016) );
CKINVDCx20_ASAP7_75t_R g989 ( .A(n_990), .Y(n_989) );
NAND2xp5_ASAP7_75t_L g990 ( .A(n_991), .B(n_992), .Y(n_990) );
NAND2xp5_ASAP7_75t_L g993 ( .A(n_994), .B(n_995), .Y(n_993) );
OAI322xp33_ASAP7_75t_L g996 ( .A1(n_997), .A2(n_1013), .A3(n_1014), .B1(n_1017), .B2(n_1020), .C1(n_1021), .C2(n_1043), .Y(n_996) );
CKINVDCx20_ASAP7_75t_R g998 ( .A(n_999), .Y(n_998) );
HB1xp67_ASAP7_75t_L g999 ( .A(n_1000), .Y(n_999) );
NAND4xp75_ASAP7_75t_L g1000 ( .A(n_1001), .B(n_1005), .C(n_1008), .D(n_1011), .Y(n_1000) );
AND2x2_ASAP7_75t_L g1001 ( .A(n_1002), .B(n_1003), .Y(n_1001) );
AND2x2_ASAP7_75t_L g1005 ( .A(n_1006), .B(n_1007), .Y(n_1005) );
AND2x2_ASAP7_75t_SL g1008 ( .A(n_1009), .B(n_1010), .Y(n_1008) );
HB1xp67_ASAP7_75t_L g1014 ( .A(n_1015), .Y(n_1014) );
INVx1_ASAP7_75t_L g1015 ( .A(n_1016), .Y(n_1015) );
CKINVDCx16_ASAP7_75t_R g1017 ( .A(n_1018), .Y(n_1017) );
XOR2x2_ASAP7_75t_L g1021 ( .A(n_1020), .B(n_1022), .Y(n_1021) );
NAND2xp5_ASAP7_75t_L g1022 ( .A(n_1023), .B(n_1034), .Y(n_1022) );
NOR3xp33_ASAP7_75t_L g1023 ( .A(n_1024), .B(n_1027), .C(n_1031), .Y(n_1023) );
OAI21xp33_ASAP7_75t_L g1027 ( .A1(n_1028), .A2(n_1029), .B(n_1030), .Y(n_1027) );
NOR2xp33_ASAP7_75t_L g1034 ( .A(n_1035), .B(n_1039), .Y(n_1034) );
NAND2xp5_ASAP7_75t_L g1035 ( .A(n_1036), .B(n_1037), .Y(n_1035) );
NAND2xp5_ASAP7_75t_L g1039 ( .A(n_1040), .B(n_1042), .Y(n_1039) );
CKINVDCx20_ASAP7_75t_R g1043 ( .A(n_1044), .Y(n_1043) );
CKINVDCx20_ASAP7_75t_R g1044 ( .A(n_1045), .Y(n_1044) );
endmodule