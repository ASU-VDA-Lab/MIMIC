module fake_jpeg_1706_n_207 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_51, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_52, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_207);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_51;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_52;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_207;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_143;
wire n_202;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_94;
wire n_206;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g53 ( 
.A(n_24),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_10),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_30),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_15),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_52),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_11),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_6),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_36),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_0),
.Y(n_61)
);

INVx11_ASAP7_75t_SL g62 ( 
.A(n_32),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_27),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_44),
.Y(n_64)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_41),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_50),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_42),
.Y(n_67)
);

HB1xp67_ASAP7_75t_L g68 ( 
.A(n_8),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_2),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_26),
.Y(n_70)
);

BUFx10_ASAP7_75t_L g71 ( 
.A(n_45),
.Y(n_71)
);

INVx8_ASAP7_75t_L g72 ( 
.A(n_10),
.Y(n_72)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_48),
.Y(n_73)
);

INVx11_ASAP7_75t_L g74 ( 
.A(n_40),
.Y(n_74)
);

BUFx5_ASAP7_75t_L g75 ( 
.A(n_7),
.Y(n_75)
);

BUFx12_ASAP7_75t_L g76 ( 
.A(n_34),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_1),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_16),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_7),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_54),
.B(n_0),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_80),
.B(n_86),
.Y(n_89)
);

BUFx12f_ASAP7_75t_L g81 ( 
.A(n_62),
.Y(n_81)
);

BUFx3_ASAP7_75t_L g96 ( 
.A(n_81),
.Y(n_96)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_62),
.Y(n_82)
);

BUFx2_ASAP7_75t_L g99 ( 
.A(n_82),
.Y(n_99)
);

INVx11_ASAP7_75t_L g83 ( 
.A(n_71),
.Y(n_83)
);

INVx6_ASAP7_75t_L g93 ( 
.A(n_83),
.Y(n_93)
);

INVx5_ASAP7_75t_L g84 ( 
.A(n_72),
.Y(n_84)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_84),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_55),
.Y(n_85)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_85),
.Y(n_90)
);

BUFx12f_ASAP7_75t_L g86 ( 
.A(n_76),
.Y(n_86)
);

INVx6_ASAP7_75t_L g87 ( 
.A(n_55),
.Y(n_87)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_87),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_58),
.B(n_1),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_88),
.B(n_69),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_91),
.B(n_95),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_85),
.A2(n_65),
.B1(n_56),
.B2(n_61),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_94),
.A2(n_97),
.B1(n_102),
.B2(n_81),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_88),
.B(n_78),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_85),
.A2(n_65),
.B1(n_56),
.B2(n_61),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_86),
.B(n_78),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_98),
.B(n_81),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_87),
.B(n_53),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_100),
.B(n_70),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_83),
.A2(n_68),
.B1(n_72),
.B2(n_77),
.Y(n_102)
);

O2A1O1Ixp33_ASAP7_75t_SL g103 ( 
.A1(n_101),
.A2(n_90),
.B(n_89),
.C(n_97),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_103),
.A2(n_106),
.B1(n_86),
.B2(n_75),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_94),
.A2(n_84),
.B1(n_79),
.B2(n_73),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_104),
.A2(n_105),
.B1(n_120),
.B2(n_76),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_100),
.A2(n_79),
.B1(n_73),
.B2(n_67),
.Y(n_105)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_101),
.Y(n_108)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_108),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_109),
.B(n_2),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_99),
.B(n_67),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_110),
.B(n_111),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_99),
.B(n_77),
.Y(n_111)
);

A2O1A1Ixp33_ASAP7_75t_L g112 ( 
.A1(n_92),
.A2(n_59),
.B(n_57),
.C(n_64),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_112),
.B(n_115),
.Y(n_140)
);

AND2x2_ASAP7_75t_L g113 ( 
.A(n_92),
.B(n_90),
.Y(n_113)
);

CKINVDCx14_ASAP7_75t_R g139 ( 
.A(n_113),
.Y(n_139)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_96),
.Y(n_114)
);

INVx3_ASAP7_75t_L g125 ( 
.A(n_114),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_93),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_116),
.B(n_117),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_96),
.B(n_66),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_93),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_118),
.B(n_23),
.Y(n_136)
);

A2O1A1Ixp33_ASAP7_75t_L g119 ( 
.A1(n_89),
.A2(n_63),
.B(n_60),
.C(n_71),
.Y(n_119)
);

AND2x2_ASAP7_75t_L g141 ( 
.A(n_119),
.B(n_5),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_L g120 ( 
.A1(n_90),
.A2(n_82),
.B1(n_74),
.B2(n_81),
.Y(n_120)
);

HB1xp67_ASAP7_75t_L g121 ( 
.A(n_92),
.Y(n_121)
);

BUFx2_ASAP7_75t_SL g146 ( 
.A(n_121),
.Y(n_146)
);

O2A1O1Ixp33_ASAP7_75t_L g122 ( 
.A1(n_92),
.A2(n_86),
.B(n_71),
.C(n_74),
.Y(n_122)
);

INVxp67_ASAP7_75t_L g144 ( 
.A(n_122),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_124),
.A2(n_126),
.B1(n_135),
.B2(n_143),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_106),
.A2(n_75),
.B1(n_76),
.B2(n_4),
.Y(n_126)
);

AND2x2_ASAP7_75t_L g162 ( 
.A(n_128),
.B(n_141),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_116),
.B(n_21),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_129),
.B(n_132),
.Y(n_148)
);

INVxp67_ASAP7_75t_L g153 ( 
.A(n_130),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_107),
.B(n_3),
.Y(n_132)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_108),
.Y(n_133)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_133),
.Y(n_154)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_113),
.Y(n_134)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_134),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_104),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_136),
.B(n_145),
.Y(n_150)
);

INVx8_ASAP7_75t_L g137 ( 
.A(n_122),
.Y(n_137)
);

INVx4_ASAP7_75t_L g157 ( 
.A(n_137),
.Y(n_157)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_113),
.Y(n_138)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_138),
.Y(n_169)
);

AND2x2_ASAP7_75t_L g142 ( 
.A(n_119),
.B(n_6),
.Y(n_142)
);

AND2x2_ASAP7_75t_L g168 ( 
.A(n_142),
.B(n_25),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_105),
.A2(n_8),
.B1(n_9),
.B2(n_11),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_112),
.B(n_9),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_L g147 ( 
.A1(n_144),
.A2(n_103),
.B1(n_114),
.B2(n_14),
.Y(n_147)
);

INVxp67_ASAP7_75t_L g179 ( 
.A(n_147),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_123),
.B(n_12),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_149),
.B(n_156),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_124),
.A2(n_12),
.B1(n_13),
.B2(n_14),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_139),
.B(n_31),
.C(n_49),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_152),
.B(n_143),
.C(n_33),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_144),
.A2(n_29),
.B1(n_47),
.B2(n_46),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_131),
.B(n_142),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_SL g158 ( 
.A1(n_140),
.A2(n_13),
.B(n_15),
.Y(n_158)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_158),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_129),
.B(n_17),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_159),
.B(n_160),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_141),
.B(n_127),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_137),
.A2(n_18),
.B1(n_19),
.B2(n_20),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_125),
.B(n_19),
.Y(n_163)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_163),
.Y(n_175)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_146),
.Y(n_165)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_165),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_125),
.B(n_22),
.Y(n_166)
);

CKINVDCx16_ASAP7_75t_R g180 ( 
.A(n_166),
.Y(n_180)
);

CKINVDCx16_ASAP7_75t_R g181 ( 
.A(n_168),
.Y(n_181)
);

OAI322xp33_ASAP7_75t_L g188 ( 
.A1(n_170),
.A2(n_168),
.A3(n_148),
.B1(n_43),
.B2(n_39),
.C1(n_37),
.C2(n_153),
.Y(n_188)
);

BUFx6f_ASAP7_75t_L g171 ( 
.A(n_154),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_171),
.A2(n_182),
.B1(n_157),
.B2(n_162),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_164),
.B(n_28),
.C(n_35),
.Y(n_172)
);

XOR2xp5_ASAP7_75t_L g183 ( 
.A(n_172),
.B(n_152),
.Y(n_183)
);

AOI21xp5_ASAP7_75t_L g174 ( 
.A1(n_157),
.A2(n_51),
.B(n_38),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_L g185 ( 
.A1(n_174),
.A2(n_155),
.B(n_172),
.Y(n_185)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_169),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g192 ( 
.A(n_183),
.B(n_186),
.Y(n_192)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_184),
.Y(n_195)
);

HB1xp67_ASAP7_75t_L g194 ( 
.A(n_185),
.Y(n_194)
);

AOI22xp33_ASAP7_75t_L g186 ( 
.A1(n_179),
.A2(n_167),
.B1(n_147),
.B2(n_162),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_179),
.A2(n_161),
.B1(n_151),
.B2(n_150),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_187),
.B(n_188),
.C(n_189),
.Y(n_191)
);

XOR2xp5_ASAP7_75t_L g189 ( 
.A(n_176),
.B(n_153),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_SL g190 ( 
.A1(n_173),
.A2(n_174),
.B(n_176),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_190),
.B(n_181),
.C(n_177),
.Y(n_193)
);

XOR2xp5_ASAP7_75t_L g198 ( 
.A(n_193),
.B(n_183),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_SL g196 ( 
.A(n_191),
.B(n_189),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_R g199 ( 
.A(n_196),
.B(n_194),
.Y(n_199)
);

INVx2_ASAP7_75t_SL g197 ( 
.A(n_195),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_197),
.B(n_198),
.Y(n_200)
);

CKINVDCx16_ASAP7_75t_R g201 ( 
.A(n_199),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_201),
.B(n_200),
.C(n_192),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_202),
.Y(n_203)
);

AO21x2_ASAP7_75t_L g204 ( 
.A1(n_203),
.A2(n_175),
.B(n_197),
.Y(n_204)
);

CKINVDCx16_ASAP7_75t_R g205 ( 
.A(n_204),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_L g206 ( 
.A1(n_205),
.A2(n_180),
.B(n_186),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_206),
.B(n_178),
.Y(n_207)
);


endmodule