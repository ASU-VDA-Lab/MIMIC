module fake_jpeg_28467_n_146 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_146);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_146;

wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVxp67_ASAP7_75t_L g13 ( 
.A(n_10),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_12),
.Y(n_14)
);

INVx6_ASAP7_75t_L g15 ( 
.A(n_3),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_2),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_11),
.Y(n_18)
);

INVx4_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_7),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_5),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_11),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_10),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_19),
.Y(n_30)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_30),
.Y(n_47)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_19),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_31),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_32),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_33),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_15),
.Y(n_34)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_34),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_13),
.B(n_20),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_35),
.B(n_38),
.Y(n_48)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_19),
.Y(n_36)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

INVx11_ASAP7_75t_L g37 ( 
.A(n_22),
.Y(n_37)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_37),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_14),
.B(n_9),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_22),
.Y(n_39)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_39),
.Y(n_52)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_22),
.Y(n_40)
);

CKINVDCx16_ASAP7_75t_R g56 ( 
.A(n_40),
.Y(n_56)
);

AND2x2_ASAP7_75t_L g41 ( 
.A(n_23),
.B(n_29),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_41),
.B(n_29),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_SL g45 ( 
.A(n_30),
.B(n_20),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_45),
.B(n_50),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_L g49 ( 
.A1(n_39),
.A2(n_28),
.B1(n_26),
.B2(n_17),
.Y(n_49)
);

OAI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_49),
.A2(n_33),
.B1(n_34),
.B2(n_18),
.Y(n_76)
);

A2O1A1Ixp33_ASAP7_75t_L g50 ( 
.A1(n_41),
.A2(n_21),
.B(n_16),
.C(n_24),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_41),
.B(n_24),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_53),
.B(n_27),
.Y(n_68)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_36),
.Y(n_55)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_55),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_40),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_57),
.B(n_60),
.Y(n_66)
);

AND2x2_ASAP7_75t_L g69 ( 
.A(n_58),
.B(n_23),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g59 ( 
.A1(n_39),
.A2(n_28),
.B1(n_26),
.B2(n_23),
.Y(n_59)
);

OA22x2_ASAP7_75t_L g61 ( 
.A1(n_59),
.A2(n_37),
.B1(n_21),
.B2(n_16),
.Y(n_61)
);

CKINVDCx16_ASAP7_75t_R g60 ( 
.A(n_31),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_61),
.A2(n_54),
.B1(n_1),
.B2(n_2),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_48),
.B(n_18),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_63),
.B(n_68),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_50),
.A2(n_17),
.B1(n_27),
.B2(n_25),
.Y(n_65)
);

OAI21xp5_ASAP7_75t_SL g86 ( 
.A1(n_65),
.A2(n_71),
.B(n_74),
.Y(n_86)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_47),
.Y(n_67)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_67),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_69),
.B(n_78),
.Y(n_84)
);

HB1xp67_ASAP7_75t_L g70 ( 
.A(n_51),
.Y(n_70)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_70),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_55),
.A2(n_40),
.B1(n_28),
.B2(n_26),
.Y(n_71)
);

HB1xp67_ASAP7_75t_L g72 ( 
.A(n_51),
.Y(n_72)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_72),
.Y(n_91)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_47),
.Y(n_73)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_73),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_52),
.A2(n_40),
.B1(n_32),
.B2(n_33),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_53),
.B(n_25),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_75),
.B(n_77),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_76),
.A2(n_46),
.B1(n_43),
.B2(n_42),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_57),
.B(n_14),
.Y(n_77)
);

INVxp67_ASAP7_75t_L g78 ( 
.A(n_52),
.Y(n_78)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_44),
.Y(n_79)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_79),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_56),
.B(n_9),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_80),
.B(n_81),
.Y(n_94)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_59),
.B(n_34),
.Y(n_81)
);

OAI32xp33_ASAP7_75t_L g87 ( 
.A1(n_64),
.A2(n_43),
.A3(n_44),
.B1(n_46),
.B2(n_42),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_87),
.B(n_61),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_77),
.B(n_0),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_88),
.B(n_90),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_89),
.A2(n_93),
.B1(n_81),
.B2(n_61),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_75),
.B(n_0),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_80),
.B(n_0),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_97),
.B(n_68),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_83),
.B(n_64),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_99),
.B(n_100),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_94),
.B(n_66),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_94),
.B(n_66),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_101),
.B(n_102),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_84),
.B(n_69),
.C(n_83),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_103),
.B(n_86),
.C(n_91),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_104),
.Y(n_112)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_105),
.Y(n_114)
);

BUFx2_ASAP7_75t_L g106 ( 
.A(n_92),
.Y(n_106)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_106),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_82),
.B(n_65),
.Y(n_107)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_107),
.Y(n_120)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_95),
.Y(n_108)
);

HB1xp67_ASAP7_75t_L g119 ( 
.A(n_108),
.Y(n_119)
);

NAND2xp33_ASAP7_75t_SL g109 ( 
.A(n_87),
.B(n_62),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_109),
.A2(n_86),
.B1(n_92),
.B2(n_95),
.Y(n_111)
);

A2O1A1O1Ixp25_ASAP7_75t_L g110 ( 
.A1(n_93),
.A2(n_69),
.B(n_62),
.C(n_61),
.D(n_73),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_110),
.B(n_81),
.C(n_89),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_111),
.A2(n_109),
.B1(n_110),
.B2(n_102),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_113),
.B(n_96),
.C(n_78),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_L g122 ( 
.A(n_115),
.B(n_103),
.Y(n_122)
);

NOR3xp33_ASAP7_75t_L g121 ( 
.A(n_120),
.B(n_101),
.C(n_100),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_121),
.A2(n_124),
.B1(n_125),
.B2(n_126),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_122),
.B(n_123),
.C(n_127),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_L g123 ( 
.A(n_113),
.B(n_98),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_112),
.B(n_106),
.Y(n_125)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_119),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_112),
.B(n_91),
.C(n_96),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_128),
.A2(n_117),
.B1(n_114),
.B2(n_116),
.Y(n_130)
);

XOR2xp5_ASAP7_75t_L g136 ( 
.A(n_130),
.B(n_131),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_121),
.A2(n_114),
.B1(n_118),
.B2(n_85),
.Y(n_131)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_131),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_128),
.A2(n_85),
.B1(n_79),
.B2(n_67),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_132),
.B(n_133),
.Y(n_134)
);

OAI221xp5_ASAP7_75t_L g138 ( 
.A1(n_134),
.A2(n_132),
.B1(n_130),
.B2(n_129),
.C(n_5),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_SL g139 ( 
.A(n_136),
.B(n_137),
.Y(n_139)
);

XOR2xp5_ASAP7_75t_L g137 ( 
.A(n_129),
.B(n_54),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_138),
.A2(n_140),
.B1(n_1),
.B2(n_3),
.Y(n_142)
);

NOR2xp67_ASAP7_75t_L g140 ( 
.A(n_136),
.B(n_1),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_139),
.B(n_135),
.C(n_2),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_141),
.B(n_142),
.Y(n_143)
);

AOI21xp5_ASAP7_75t_SL g144 ( 
.A1(n_143),
.A2(n_3),
.B(n_5),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_144),
.B(n_6),
.Y(n_145)
);

XOR2xp5_ASAP7_75t_L g146 ( 
.A(n_145),
.B(n_6),
.Y(n_146)
);


endmodule