module fake_jpeg_29815_n_140 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_140);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_140;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

INVx1_ASAP7_75t_L g12 ( 
.A(n_4),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_6),
.Y(n_13)
);

INVx8_ASAP7_75t_L g14 ( 
.A(n_0),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_9),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

INVx11_ASAP7_75t_SL g17 ( 
.A(n_11),
.Y(n_17)
);

BUFx10_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_4),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_4),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_10),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_1),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_7),
.Y(n_25)
);

BUFx12_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

INVx2_ASAP7_75t_SL g27 ( 
.A(n_17),
.Y(n_27)
);

BUFx8_ASAP7_75t_L g47 ( 
.A(n_27),
.Y(n_47)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_28),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_16),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_29),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_16),
.Y(n_30)
);

INVx5_ASAP7_75t_L g52 ( 
.A(n_30),
.Y(n_52)
);

CKINVDCx14_ASAP7_75t_R g31 ( 
.A(n_19),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_31),
.B(n_37),
.Y(n_46)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_19),
.Y(n_32)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_32),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_33),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_34),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_16),
.Y(n_35)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_35),
.Y(n_57)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_18),
.Y(n_36)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_36),
.Y(n_60)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_12),
.Y(n_37)
);

INVx5_ASAP7_75t_L g38 ( 
.A(n_18),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_38),
.B(n_39),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_18),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_20),
.B(n_0),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_40),
.B(n_21),
.Y(n_58)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_18),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_41),
.B(n_42),
.Y(n_54)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_26),
.Y(n_42)
);

INVxp67_ASAP7_75t_L g43 ( 
.A(n_27),
.Y(n_43)
);

INVx13_ASAP7_75t_L g73 ( 
.A(n_43),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_L g50 ( 
.A1(n_29),
.A2(n_30),
.B1(n_35),
.B2(n_39),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g68 ( 
.A1(n_50),
.A2(n_51),
.B1(n_56),
.B2(n_38),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_36),
.A2(n_12),
.B1(n_20),
.B2(n_24),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_42),
.B(n_22),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_55),
.B(n_26),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_41),
.A2(n_24),
.B1(n_21),
.B2(n_13),
.Y(n_56)
);

OR2x2_ASAP7_75t_L g75 ( 
.A(n_58),
.B(n_15),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_46),
.B(n_25),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_61),
.B(n_64),
.Y(n_89)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_44),
.Y(n_62)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_62),
.Y(n_88)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_48),
.Y(n_63)
);

BUFx2_ASAP7_75t_L g80 ( 
.A(n_63),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_44),
.B(n_25),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_57),
.B(n_13),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_65),
.B(n_70),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_66),
.B(n_74),
.Y(n_84)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_59),
.Y(n_67)
);

INVxp67_ASAP7_75t_L g91 ( 
.A(n_67),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_68),
.A2(n_52),
.B1(n_49),
.B2(n_33),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_47),
.B(n_22),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g93 ( 
.A(n_69),
.B(n_72),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_57),
.B(n_23),
.Y(n_70)
);

XOR2x2_ASAP7_75t_L g71 ( 
.A(n_54),
.B(n_26),
.Y(n_71)
);

XNOR2xp5_ASAP7_75t_L g86 ( 
.A(n_71),
.B(n_76),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_SL g72 ( 
.A(n_47),
.B(n_23),
.Y(n_72)
);

INVxp67_ASAP7_75t_L g74 ( 
.A(n_47),
.Y(n_74)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_75),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_45),
.B(n_15),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_60),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_77),
.A2(n_78),
.B1(n_1),
.B2(n_2),
.Y(n_92)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_48),
.Y(n_78)
);

AND2x2_ASAP7_75t_L g79 ( 
.A(n_53),
.B(n_34),
.Y(n_79)
);

AO22x1_ASAP7_75t_L g87 ( 
.A1(n_79),
.A2(n_43),
.B1(n_26),
.B2(n_3),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_71),
.A2(n_49),
.B1(n_45),
.B2(n_52),
.Y(n_82)
);

INVxp67_ASAP7_75t_L g102 ( 
.A(n_82),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_83),
.B(n_79),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_L g85 ( 
.A1(n_62),
.A2(n_60),
.B1(n_59),
.B2(n_47),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_85),
.B(n_73),
.Y(n_96)
);

OAI21xp5_ASAP7_75t_SL g94 ( 
.A1(n_87),
.A2(n_92),
.B(n_74),
.Y(n_94)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_94),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_95),
.A2(n_87),
.B1(n_89),
.B2(n_70),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_96),
.A2(n_77),
.B1(n_91),
.B2(n_78),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_93),
.B(n_72),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_97),
.B(n_99),
.Y(n_107)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_88),
.Y(n_98)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_98),
.Y(n_106)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_80),
.Y(n_99)
);

XNOR2xp5_ASAP7_75t_L g100 ( 
.A(n_86),
.B(n_79),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_100),
.B(n_76),
.C(n_64),
.Y(n_109)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_80),
.Y(n_101)
);

NOR3xp33_ASAP7_75t_L g110 ( 
.A(n_101),
.B(n_103),
.C(n_104),
.Y(n_110)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_84),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_89),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_102),
.A2(n_82),
.B1(n_86),
.B2(n_81),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_105),
.A2(n_111),
.B1(n_91),
.B2(n_99),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_108),
.B(n_98),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_109),
.B(n_65),
.C(n_61),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_102),
.A2(n_87),
.B1(n_83),
.B2(n_90),
.Y(n_111)
);

OR2x2_ASAP7_75t_L g120 ( 
.A(n_113),
.B(n_63),
.Y(n_120)
);

NOR2xp67_ASAP7_75t_L g114 ( 
.A(n_110),
.B(n_100),
.Y(n_114)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_114),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_SL g124 ( 
.A1(n_115),
.A2(n_117),
.B(n_73),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_116),
.A2(n_120),
.B1(n_1),
.B2(n_2),
.Y(n_127)
);

AOI21xp33_ASAP7_75t_L g117 ( 
.A1(n_107),
.A2(n_94),
.B(n_75),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_SL g118 ( 
.A1(n_112),
.A2(n_105),
.B(n_111),
.Y(n_118)
);

AOI21xp5_ASAP7_75t_L g123 ( 
.A1(n_118),
.A2(n_112),
.B(n_67),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_106),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_119),
.Y(n_125)
);

AND2x2_ASAP7_75t_L g122 ( 
.A(n_121),
.B(n_109),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_122),
.B(n_115),
.Y(n_130)
);

AOI21xp5_ASAP7_75t_L g129 ( 
.A1(n_123),
.A2(n_127),
.B(n_120),
.Y(n_129)
);

MAJx2_ASAP7_75t_L g128 ( 
.A(n_124),
.B(n_118),
.C(n_116),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_128),
.B(n_130),
.C(n_122),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_129),
.B(n_125),
.Y(n_133)
);

NOR2xp67_ASAP7_75t_SL g131 ( 
.A(n_126),
.B(n_5),
.Y(n_131)
);

NAND4xp25_ASAP7_75t_L g134 ( 
.A(n_131),
.B(n_5),
.C(n_6),
.D(n_8),
.Y(n_134)
);

INVxp67_ASAP7_75t_L g136 ( 
.A(n_132),
.Y(n_136)
);

A2O1A1Ixp33_ASAP7_75t_SL g135 ( 
.A1(n_133),
.A2(n_134),
.B(n_11),
.C(n_8),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_135),
.B(n_3),
.Y(n_137)
);

INVxp67_ASAP7_75t_L g138 ( 
.A(n_137),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_138),
.B(n_136),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_L g140 ( 
.A(n_139),
.B(n_3),
.Y(n_140)
);


endmodule