module fake_jpeg_14813_n_245 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_245);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_245;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_233;
wire n_102;
wire n_121;
wire n_130;
wire n_99;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_145;
wire n_18;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_11),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

BUFx10_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_5),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_2),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_0),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_8),
.Y(n_30)
);

INVx2_ASAP7_75t_R g31 ( 
.A(n_4),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_13),
.Y(n_32)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_28),
.Y(n_33)
);

INVx5_ASAP7_75t_L g52 ( 
.A(n_33),
.Y(n_52)
);

INVx11_ASAP7_75t_L g34 ( 
.A(n_31),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_34),
.Y(n_57)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_28),
.Y(n_35)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_35),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_28),
.Y(n_36)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_36),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_25),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_37),
.B(n_38),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_20),
.B(n_0),
.Y(n_38)
);

INVx11_ASAP7_75t_L g39 ( 
.A(n_31),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_39),
.B(n_40),
.Y(n_46)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_25),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_20),
.B(n_0),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_41),
.B(n_16),
.Y(n_53)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_35),
.Y(n_42)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_42),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_38),
.B(n_24),
.Y(n_47)
);

AND2x2_ASAP7_75t_L g60 ( 
.A(n_47),
.B(n_50),
.Y(n_60)
);

OA22x2_ASAP7_75t_L g48 ( 
.A1(n_35),
.A2(n_31),
.B1(n_19),
.B2(n_30),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_48),
.A2(n_51),
.B1(n_55),
.B2(n_39),
.Y(n_72)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_49),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_38),
.B(n_24),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g51 ( 
.A1(n_41),
.A2(n_24),
.B1(n_31),
.B2(n_30),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_53),
.B(n_21),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_41),
.B(n_16),
.Y(n_54)
);

AND2x2_ASAP7_75t_L g80 ( 
.A(n_54),
.B(n_29),
.Y(n_80)
);

OAI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_34),
.A2(n_39),
.B1(n_29),
.B2(n_26),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_34),
.B(n_17),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_SL g81 ( 
.A(n_56),
.B(n_25),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_54),
.B(n_22),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_58),
.B(n_62),
.Y(n_102)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_44),
.Y(n_59)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_59),
.Y(n_88)
);

INVx1_ASAP7_75t_SL g61 ( 
.A(n_57),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_61),
.B(n_63),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_43),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_53),
.B(n_32),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_64),
.B(n_65),
.Y(n_98)
);

CKINVDCx16_ASAP7_75t_R g65 ( 
.A(n_46),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_56),
.B(n_32),
.Y(n_67)
);

CKINVDCx16_ASAP7_75t_R g96 ( 
.A(n_67),
.Y(n_96)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_44),
.Y(n_69)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_69),
.Y(n_90)
);

A2O1A1Ixp33_ASAP7_75t_L g70 ( 
.A1(n_45),
.A2(n_34),
.B(n_39),
.C(n_26),
.Y(n_70)
);

MAJIxp5_ASAP7_75t_SL g104 ( 
.A(n_70),
.B(n_72),
.C(n_80),
.Y(n_104)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_43),
.Y(n_71)
);

CKINVDCx16_ASAP7_75t_R g100 ( 
.A(n_71),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g73 ( 
.A(n_46),
.Y(n_73)
);

CKINVDCx16_ASAP7_75t_R g110 ( 
.A(n_73),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_52),
.A2(n_33),
.B1(n_40),
.B2(n_23),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_74),
.A2(n_83),
.B1(n_27),
.B2(n_36),
.Y(n_109)
);

AO22x2_ASAP7_75t_SL g75 ( 
.A1(n_48),
.A2(n_36),
.B1(n_40),
.B2(n_33),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_75),
.A2(n_33),
.B1(n_36),
.B2(n_37),
.Y(n_107)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_52),
.Y(n_76)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_76),
.Y(n_91)
);

INVx4_ASAP7_75t_SL g77 ( 
.A(n_57),
.Y(n_77)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_77),
.Y(n_92)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_57),
.Y(n_78)
);

INVxp67_ASAP7_75t_L g99 ( 
.A(n_78),
.Y(n_99)
);

INVxp67_ASAP7_75t_L g79 ( 
.A(n_48),
.Y(n_79)
);

INVxp67_ASAP7_75t_L g106 ( 
.A(n_79),
.Y(n_106)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_81),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_48),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_82),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_42),
.A2(n_33),
.B1(n_40),
.B2(n_17),
.Y(n_83)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_47),
.B(n_21),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g93 ( 
.A(n_84),
.B(n_86),
.Y(n_93)
);

INVx8_ASAP7_75t_L g85 ( 
.A(n_49),
.Y(n_85)
);

INVx8_ASAP7_75t_L g89 ( 
.A(n_85),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_50),
.B(n_23),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_45),
.B(n_22),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_87),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_60),
.B(n_36),
.C(n_51),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_94),
.B(n_72),
.C(n_73),
.Y(n_118)
);

NOR2x1_ASAP7_75t_L g97 ( 
.A(n_75),
.B(n_48),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g130 ( 
.A(n_97),
.B(n_37),
.Y(n_130)
);

AND2x2_ASAP7_75t_L g101 ( 
.A(n_75),
.B(n_36),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_SL g139 ( 
.A1(n_101),
.A2(n_77),
.B(n_78),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_107),
.A2(n_109),
.B1(n_111),
.B2(n_61),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_60),
.B(n_84),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_108),
.B(n_60),
.Y(n_115)
);

OAI22xp33_ASAP7_75t_L g111 ( 
.A1(n_79),
.A2(n_19),
.B1(n_36),
.B2(n_27),
.Y(n_111)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_69),
.Y(n_113)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_113),
.Y(n_119)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_95),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_114),
.B(n_117),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_L g158 ( 
.A(n_115),
.B(n_102),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_116),
.A2(n_101),
.B1(n_97),
.B2(n_106),
.Y(n_143)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_98),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_118),
.B(n_124),
.C(n_136),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_88),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_120),
.B(n_122),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_96),
.B(n_71),
.Y(n_121)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_121),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_88),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_108),
.B(n_84),
.Y(n_123)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_123),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_94),
.B(n_37),
.C(n_70),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_103),
.B(n_80),
.Y(n_125)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_125),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_90),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_126),
.B(n_129),
.Y(n_157)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_90),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_127),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_93),
.B(n_80),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_L g142 ( 
.A1(n_128),
.A2(n_130),
.B(n_131),
.Y(n_142)
);

CKINVDCx16_ASAP7_75t_R g129 ( 
.A(n_92),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_93),
.B(n_68),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_113),
.Y(n_132)
);

INVxp67_ASAP7_75t_SL g155 ( 
.A(n_132),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_91),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_SL g156 ( 
.A(n_133),
.B(n_134),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_105),
.B(n_66),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_105),
.B(n_66),
.Y(n_135)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_135),
.Y(n_145)
);

XOR2xp5_ASAP7_75t_L g136 ( 
.A(n_104),
.B(n_28),
.Y(n_136)
);

CKINVDCx14_ASAP7_75t_R g137 ( 
.A(n_107),
.Y(n_137)
);

INVx1_ASAP7_75t_SL g153 ( 
.A(n_137),
.Y(n_153)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_91),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_138),
.A2(n_110),
.B1(n_100),
.B2(n_68),
.Y(n_148)
);

AOI21xp5_ASAP7_75t_L g152 ( 
.A1(n_139),
.A2(n_106),
.B(n_101),
.Y(n_152)
);

XOR2xp5_ASAP7_75t_L g140 ( 
.A(n_118),
.B(n_104),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_140),
.B(n_141),
.C(n_158),
.Y(n_180)
);

XOR2xp5_ASAP7_75t_L g141 ( 
.A(n_136),
.B(n_93),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_143),
.A2(n_152),
.B1(n_85),
.B2(n_127),
.Y(n_169)
);

AND2x2_ASAP7_75t_L g176 ( 
.A(n_148),
.B(n_99),
.Y(n_176)
);

INVxp67_ASAP7_75t_L g150 ( 
.A(n_134),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_150),
.B(n_162),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_115),
.B(n_124),
.C(n_131),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_159),
.B(n_164),
.Y(n_182)
);

AOI21xp5_ASAP7_75t_L g161 ( 
.A1(n_130),
.A2(n_112),
.B(n_111),
.Y(n_161)
);

NOR3xp33_ASAP7_75t_L g170 ( 
.A(n_161),
.B(n_132),
.C(n_119),
.Y(n_170)
);

INVxp67_ASAP7_75t_L g162 ( 
.A(n_135),
.Y(n_162)
);

AOI211xp5_ASAP7_75t_L g163 ( 
.A1(n_128),
.A2(n_112),
.B(n_92),
.C(n_99),
.Y(n_163)
);

AOI21xp33_ASAP7_75t_L g165 ( 
.A1(n_163),
.A2(n_125),
.B(n_139),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_123),
.B(n_76),
.C(n_89),
.Y(n_164)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_165),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_153),
.A2(n_116),
.B1(n_133),
.B2(n_126),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_166),
.A2(n_167),
.B1(n_168),
.B2(n_175),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_153),
.A2(n_120),
.B1(n_122),
.B2(n_89),
.Y(n_167)
);

AOI21xp5_ASAP7_75t_L g168 ( 
.A1(n_142),
.A2(n_129),
.B(n_138),
.Y(n_168)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_169),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_170),
.B(n_176),
.Y(n_196)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_147),
.Y(n_171)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_171),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_SL g172 ( 
.A(n_144),
.B(n_119),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_SL g188 ( 
.A(n_172),
.B(n_173),
.Y(n_188)
);

AOI322xp5_ASAP7_75t_SL g173 ( 
.A1(n_163),
.A2(n_15),
.A3(n_14),
.B1(n_12),
.B2(n_4),
.C1(n_5),
.C2(n_6),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_157),
.Y(n_174)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_174),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_154),
.A2(n_159),
.B1(n_162),
.B2(n_145),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_145),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_177),
.A2(n_181),
.B1(n_183),
.B2(n_148),
.Y(n_198)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_156),
.Y(n_178)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_178),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_143),
.A2(n_19),
.B1(n_28),
.B2(n_18),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_160),
.A2(n_18),
.B1(n_25),
.B2(n_15),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_149),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_184),
.B(n_150),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_180),
.B(n_151),
.C(n_140),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g212 ( 
.A(n_186),
.B(n_191),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_L g206 ( 
.A1(n_187),
.A2(n_200),
.B(n_1),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_180),
.B(n_151),
.C(n_141),
.Y(n_191)
);

FAx1_ASAP7_75t_SL g192 ( 
.A(n_175),
.B(n_142),
.CI(n_158),
.CON(n_192),
.SN(n_192)
);

XNOR2xp5_ASAP7_75t_L g210 ( 
.A(n_192),
.B(n_194),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_182),
.B(n_164),
.C(n_146),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_L g209 ( 
.A1(n_198),
.A2(n_2),
.B1(n_5),
.B2(n_6),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_168),
.B(n_155),
.C(n_25),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_199),
.B(n_6),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_179),
.B(n_18),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_185),
.A2(n_176),
.B1(n_174),
.B2(n_181),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_201),
.B(n_189),
.Y(n_214)
);

XOR2x2_ASAP7_75t_L g202 ( 
.A(n_192),
.B(n_166),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_L g219 ( 
.A1(n_202),
.A2(n_204),
.B1(n_205),
.B2(n_209),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_SL g203 ( 
.A(n_192),
.B(n_193),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_203),
.B(n_207),
.C(n_208),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_190),
.A2(n_176),
.B1(n_167),
.B2(n_183),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_196),
.A2(n_177),
.B1(n_12),
.B2(n_3),
.Y(n_205)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_206),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g207 ( 
.A(n_186),
.B(n_191),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_193),
.B(n_1),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_211),
.B(n_188),
.Y(n_222)
);

OAI21xp5_ASAP7_75t_L g224 ( 
.A1(n_214),
.A2(n_194),
.B(n_195),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_208),
.B(n_189),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_215),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_210),
.B(n_197),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_216),
.B(n_217),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_SL g217 ( 
.A(n_202),
.B(n_195),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_203),
.B(n_187),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_218),
.B(n_212),
.Y(n_228)
);

OR2x2_ASAP7_75t_L g221 ( 
.A(n_207),
.B(n_200),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_221),
.B(n_222),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_SL g232 ( 
.A(n_224),
.B(n_221),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_213),
.B(n_199),
.Y(n_226)
);

OR2x2_ASAP7_75t_L g234 ( 
.A(n_226),
.B(n_220),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_219),
.B(n_198),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_227),
.B(n_228),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_229),
.B(n_218),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_231),
.B(n_232),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_223),
.B(n_220),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_233),
.B(n_234),
.Y(n_238)
);

NAND2xp33_ASAP7_75t_R g235 ( 
.A(n_231),
.B(n_225),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_235),
.B(n_9),
.C(n_10),
.Y(n_240)
);

AOI21xp5_ASAP7_75t_L g236 ( 
.A1(n_230),
.A2(n_228),
.B(n_9),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_236),
.B(n_9),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g239 ( 
.A(n_237),
.B(n_7),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_239),
.B(n_238),
.C(n_10),
.Y(n_243)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_240),
.B(n_241),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_243),
.B(n_239),
.Y(n_244)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_244),
.B(n_242),
.Y(n_245)
);


endmodule