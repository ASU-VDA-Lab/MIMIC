module fake_netlist_5_882_n_1693 (n_137, n_164, n_91, n_82, n_122, n_142, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_165, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_60, n_155, n_152, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_125, n_35, n_167, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_156, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_157, n_29, n_79, n_131, n_151, n_47, n_25, n_53, n_160, n_8, n_158, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_85, n_159, n_163, n_95, n_119, n_59, n_26, n_133, n_55, n_99, n_2, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_12, n_67, n_121, n_36, n_76, n_87, n_150, n_162, n_27, n_64, n_77, n_102, n_106, n_161, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_134, n_32, n_41, n_104, n_103, n_56, n_51, n_63, n_97, n_141, n_166, n_11, n_153, n_7, n_15, n_145, n_48, n_50, n_52, n_88, n_110, n_1693);

input n_137;
input n_164;
input n_91;
input n_82;
input n_122;
input n_142;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_165;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_60;
input n_155;
input n_152;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_125;
input n_35;
input n_167;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_157;
input n_29;
input n_79;
input n_131;
input n_151;
input n_47;
input n_25;
input n_53;
input n_160;
input n_8;
input n_158;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_85;
input n_159;
input n_163;
input n_95;
input n_119;
input n_59;
input n_26;
input n_133;
input n_55;
input n_99;
input n_2;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_150;
input n_162;
input n_27;
input n_64;
input n_77;
input n_102;
input n_106;
input n_161;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_134;
input n_32;
input n_41;
input n_104;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_166;
input n_11;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_1693;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1166;
wire n_469;
wire n_1508;
wire n_785;
wire n_549;
wire n_532;
wire n_1161;
wire n_1677;
wire n_1150;
wire n_226;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_1501;
wire n_880;
wire n_544;
wire n_1007;
wire n_552;
wire n_1528;
wire n_1370;
wire n_1292;
wire n_1198;
wire n_1360;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1021;
wire n_551;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1353;
wire n_800;
wire n_1347;
wire n_1535;
wire n_1666;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_915;
wire n_1545;
wire n_864;
wire n_173;
wire n_859;
wire n_951;
wire n_1264;
wire n_447;
wire n_247;
wire n_1494;
wire n_292;
wire n_625;
wire n_854;
wire n_1462;
wire n_1580;
wire n_674;
wire n_417;
wire n_516;
wire n_933;
wire n_1152;
wire n_497;
wire n_1607;
wire n_1563;
wire n_606;
wire n_275;
wire n_877;
wire n_755;
wire n_1118;
wire n_1686;
wire n_947;
wire n_1285;
wire n_373;
wire n_307;
wire n_1359;
wire n_530;
wire n_1107;
wire n_556;
wire n_1230;
wire n_668;
wire n_375;
wire n_301;
wire n_929;
wire n_1124;
wire n_902;
wire n_1576;
wire n_191;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1257;
wire n_171;
wire n_1182;
wire n_579;
wire n_1261;
wire n_938;
wire n_1098;
wire n_320;
wire n_1154;
wire n_1242;
wire n_1135;
wire n_406;
wire n_519;
wire n_1016;
wire n_1243;
wire n_546;
wire n_1280;
wire n_281;
wire n_240;
wire n_291;
wire n_231;
wire n_257;
wire n_731;
wire n_371;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_317;
wire n_1236;
wire n_1633;
wire n_569;
wire n_227;
wire n_920;
wire n_1289;
wire n_1517;
wire n_335;
wire n_1669;
wire n_370;
wire n_976;
wire n_343;
wire n_1449;
wire n_308;
wire n_1566;
wire n_297;
wire n_1078;
wire n_1670;
wire n_775;
wire n_219;
wire n_600;
wire n_1484;
wire n_1374;
wire n_1328;
wire n_223;
wire n_264;
wire n_1598;
wire n_955;
wire n_339;
wire n_1146;
wire n_882;
wire n_183;
wire n_243;
wire n_1097;
wire n_1036;
wire n_347;
wire n_550;
wire n_696;
wire n_897;
wire n_215;
wire n_350;
wire n_196;
wire n_798;
wire n_646;
wire n_1428;
wire n_436;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_580;
wire n_290;
wire n_1040;
wire n_578;
wire n_926;
wire n_344;
wire n_1218;
wire n_422;
wire n_475;
wire n_777;
wire n_1070;
wire n_1547;
wire n_1030;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_1561;
wire n_496;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_1600;
wire n_521;
wire n_663;
wire n_845;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_680;
wire n_1473;
wire n_1587;
wire n_395;
wire n_553;
wire n_901;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_214;
wire n_1672;
wire n_675;
wire n_888;
wire n_1167;
wire n_1626;
wire n_637;
wire n_1384;
wire n_1556;
wire n_184;
wire n_446;
wire n_1064;
wire n_858;
wire n_923;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_468;
wire n_213;
wire n_342;
wire n_464;
wire n_363;
wire n_1582;
wire n_197;
wire n_1069;
wire n_1075;
wire n_1450;
wire n_1322;
wire n_1471;
wire n_1459;
wire n_460;
wire n_889;
wire n_973;
wire n_477;
wire n_571;
wire n_1585;
wire n_461;
wire n_1599;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_907;
wire n_1447;
wire n_1377;
wire n_190;
wire n_989;
wire n_1039;
wire n_228;
wire n_283;
wire n_1403;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_1002;
wire n_1463;
wire n_1581;
wire n_310;
wire n_593;
wire n_748;
wire n_586;
wire n_1058;
wire n_1667;
wire n_838;
wire n_332;
wire n_1053;
wire n_1224;
wire n_349;
wire n_1248;
wire n_230;
wire n_1331;
wire n_953;
wire n_279;
wire n_1014;
wire n_1241;
wire n_289;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_440;
wire n_793;
wire n_478;
wire n_476;
wire n_1527;
wire n_534;
wire n_884;
wire n_345;
wire n_944;
wire n_1623;
wire n_1565;
wire n_182;
wire n_647;
wire n_237;
wire n_407;
wire n_1072;
wire n_857;
wire n_832;
wire n_207;
wire n_561;
wire n_1319;
wire n_1387;
wire n_1532;
wire n_1027;
wire n_971;
wire n_1156;
wire n_326;
wire n_794;
wire n_404;
wire n_686;
wire n_847;
wire n_1393;
wire n_596;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_728;
wire n_266;
wire n_1162;
wire n_272;
wire n_1538;
wire n_1199;
wire n_352;
wire n_1038;
wire n_520;
wire n_1369;
wire n_409;
wire n_1660;
wire n_887;
wire n_300;
wire n_809;
wire n_870;
wire n_931;
wire n_599;
wire n_1662;
wire n_1481;
wire n_434;
wire n_1544;
wire n_868;
wire n_639;
wire n_914;
wire n_411;
wire n_414;
wire n_1629;
wire n_1293;
wire n_965;
wire n_935;
wire n_1175;
wire n_817;
wire n_360;
wire n_1479;
wire n_759;
wire n_806;
wire n_1477;
wire n_324;
wire n_1635;
wire n_1571;
wire n_187;
wire n_1189;
wire n_1259;
wire n_1690;
wire n_706;
wire n_746;
wire n_1649;
wire n_747;
wire n_784;
wire n_1244;
wire n_431;
wire n_1194;
wire n_615;
wire n_851;
wire n_843;
wire n_523;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_1679;
wire n_776;
wire n_1415;
wire n_367;
wire n_452;
wire n_525;
wire n_1260;
wire n_1647;
wire n_1464;
wire n_649;
wire n_547;
wire n_1444;
wire n_1191;
wire n_1674;
wire n_284;
wire n_1128;
wire n_744;
wire n_590;
wire n_629;
wire n_1308;
wire n_254;
wire n_1680;
wire n_1233;
wire n_1615;
wire n_1529;
wire n_526;
wire n_372;
wire n_293;
wire n_677;
wire n_244;
wire n_1333;
wire n_1121;
wire n_368;
wire n_433;
wire n_314;
wire n_604;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_1001;
wire n_1503;
wire n_498;
wire n_1468;
wire n_1559;
wire n_689;
wire n_738;
wire n_1624;
wire n_640;
wire n_1510;
wire n_252;
wire n_624;
wire n_1380;
wire n_1617;
wire n_295;
wire n_1010;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_1195;
wire n_610;
wire n_936;
wire n_568;
wire n_1500;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_259;
wire n_448;
wire n_758;
wire n_999;
wire n_1656;
wire n_1158;
wire n_1509;
wire n_563;
wire n_1145;
wire n_878;
wire n_524;
wire n_394;
wire n_204;
wire n_1678;
wire n_1049;
wire n_1153;
wire n_741;
wire n_1639;
wire n_1306;
wire n_1068;
wire n_331;
wire n_906;
wire n_1163;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_658;
wire n_1362;
wire n_1586;
wire n_456;
wire n_959;
wire n_535;
wire n_940;
wire n_1445;
wire n_1492;
wire n_592;
wire n_1169;
wire n_1596;
wire n_1692;
wire n_1017;
wire n_978;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_1095;
wire n_1614;
wire n_267;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_603;
wire n_1431;
wire n_484;
wire n_1593;
wire n_1033;
wire n_442;
wire n_636;
wire n_660;
wire n_1640;
wire n_1009;
wire n_1148;
wire n_750;
wire n_742;
wire n_995;
wire n_454;
wire n_1609;
wire n_374;
wire n_185;
wire n_396;
wire n_1383;
wire n_1073;
wire n_255;
wire n_662;
wire n_459;
wire n_218;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1065;
wire n_1592;
wire n_1336;
wire n_1574;
wire n_473;
wire n_1309;
wire n_1426;
wire n_1043;
wire n_355;
wire n_486;
wire n_1548;
wire n_614;
wire n_337;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_168;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_208;
wire n_743;
wire n_299;
wire n_303;
wire n_296;
wire n_613;
wire n_1119;
wire n_1240;
wire n_829;
wire n_1612;
wire n_1416;
wire n_361;
wire n_700;
wire n_1237;
wire n_573;
wire n_1420;
wire n_1132;
wire n_388;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_761;
wire n_1568;
wire n_1006;
wire n_329;
wire n_274;
wire n_1270;
wire n_1664;
wire n_1486;
wire n_582;
wire n_1332;
wire n_1390;
wire n_309;
wire n_512;
wire n_1591;
wire n_322;
wire n_1682;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1349;
wire n_1093;
wire n_288;
wire n_1031;
wire n_263;
wire n_609;
wire n_1041;
wire n_1265;
wire n_224;
wire n_1562;
wire n_383;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_239;
wire n_630;
wire n_504;
wire n_511;
wire n_874;
wire n_358;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_1304;
wire n_1324;
wire n_987;
wire n_261;
wire n_174;
wire n_1455;
wire n_767;
wire n_993;
wire n_1407;
wire n_1551;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_429;
wire n_948;
wire n_1217;
wire n_628;
wire n_365;
wire n_729;
wire n_1131;
wire n_1084;
wire n_970;
wire n_911;
wire n_1430;
wire n_513;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1534;
wire n_340;
wire n_1351;
wire n_1044;
wire n_1205;
wire n_346;
wire n_1209;
wire n_1552;
wire n_495;
wire n_602;
wire n_574;
wire n_1435;
wire n_879;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_1645;
wire n_490;
wire n_1327;
wire n_996;
wire n_921;
wire n_1684;
wire n_233;
wire n_572;
wire n_366;
wire n_815;
wire n_327;
wire n_1381;
wire n_1611;
wire n_1037;
wire n_1080;
wire n_1274;
wire n_1316;
wire n_426;
wire n_1438;
wire n_1082;
wire n_589;
wire n_716;
wire n_1630;
wire n_562;
wire n_1436;
wire n_1691;
wire n_952;
wire n_1229;
wire n_391;
wire n_701;
wire n_1437;
wire n_1023;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_238;
wire n_531;
wire n_890;
wire n_764;
wire n_1056;
wire n_1424;
wire n_960;
wire n_222;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_634;
wire n_199;
wire n_1252;
wire n_348;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_1311;
wire n_1519;
wire n_256;
wire n_950;
wire n_1553;
wire n_380;
wire n_419;
wire n_1346;
wire n_444;
wire n_1299;
wire n_1060;
wire n_1141;
wire n_316;
wire n_389;
wire n_418;
wire n_248;
wire n_912;
wire n_315;
wire n_968;
wire n_451;
wire n_619;
wire n_408;
wire n_1386;
wire n_376;
wire n_967;
wire n_1442;
wire n_1139;
wire n_515;
wire n_351;
wire n_885;
wire n_397;
wire n_1432;
wire n_1357;
wire n_483;
wire n_683;
wire n_1632;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_1608;
wire n_983;
wire n_280;
wire n_1305;
wire n_873;
wire n_378;
wire n_1112;
wire n_762;
wire n_1283;
wire n_1644;
wire n_690;
wire n_583;
wire n_302;
wire n_1343;
wire n_1203;
wire n_1631;
wire n_821;
wire n_321;
wire n_1179;
wire n_621;
wire n_753;
wire n_455;
wire n_1048;
wire n_1288;
wire n_212;
wire n_385;
wire n_507;
wire n_1560;
wire n_1605;
wire n_330;
wire n_1228;
wire n_972;
wire n_692;
wire n_820;
wire n_1200;
wire n_1301;
wire n_1363;
wire n_1668;
wire n_1185;
wire n_991;
wire n_828;
wire n_779;
wire n_576;
wire n_1143;
wire n_1579;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_537;
wire n_1688;
wire n_945;
wire n_492;
wire n_1504;
wire n_943;
wire n_341;
wire n_250;
wire n_992;
wire n_543;
wire n_260;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_286;
wire n_1643;
wire n_883;
wire n_470;
wire n_325;
wire n_449;
wire n_1594;
wire n_1214;
wire n_1342;
wire n_1400;
wire n_900;
wire n_856;
wire n_918;
wire n_942;
wire n_189;
wire n_1147;
wire n_1557;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_540;
wire n_618;
wire n_896;
wire n_323;
wire n_195;
wire n_356;
wire n_894;
wire n_1636;
wire n_831;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1470;
wire n_1096;
wire n_234;
wire n_1575;
wire n_833;
wire n_1646;
wire n_225;
wire n_1307;
wire n_988;
wire n_814;
wire n_192;
wire n_1549;
wire n_1201;
wire n_1114;
wire n_655;
wire n_1616;
wire n_1446;
wire n_669;
wire n_472;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_387;
wire n_1149;
wire n_398;
wire n_1671;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_211;
wire n_1219;
wire n_1204;
wire n_178;
wire n_1035;
wire n_287;
wire n_555;
wire n_783;
wire n_1188;
wire n_661;
wire n_849;
wire n_336;
wire n_584;
wire n_681;
wire n_1638;
wire n_430;
wire n_510;
wire n_216;
wire n_311;
wire n_830;
wire n_1296;
wire n_1413;
wire n_801;
wire n_241;
wire n_875;
wire n_357;
wire n_1110;
wire n_1655;
wire n_445;
wire n_749;
wire n_1134;
wire n_1358;
wire n_717;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_249;
wire n_304;
wire n_1338;
wire n_577;
wire n_1522;
wire n_1687;
wire n_1637;
wire n_1419;
wire n_338;
wire n_1653;
wire n_693;
wire n_1506;
wire n_836;
wire n_990;
wire n_1389;
wire n_975;
wire n_1256;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_306;
wire n_458;
wire n_770;
wire n_1375;
wire n_1102;
wire n_711;
wire n_1499;
wire n_1187;
wire n_1441;
wire n_1392;
wire n_1597;
wire n_1164;
wire n_1659;
wire n_489;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_1572;
wire n_876;
wire n_1516;
wire n_1190;
wire n_1685;
wire n_601;
wire n_917;
wire n_966;
wire n_253;
wire n_1116;
wire n_1661;
wire n_1212;
wire n_1541;
wire n_206;
wire n_172;
wire n_217;
wire n_726;
wire n_982;
wire n_1573;
wire n_1453;
wire n_818;
wire n_861;
wire n_1183;
wire n_1658;
wire n_899;
wire n_1253;
wire n_210;
wire n_774;
wire n_1628;
wire n_1335;
wire n_1514;
wire n_1059;
wire n_1345;
wire n_176;
wire n_1133;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_527;
wire n_1168;
wire n_707;
wire n_937;
wire n_1427;
wire n_393;
wire n_487;
wire n_1584;
wire n_665;
wire n_1440;
wire n_177;
wire n_421;
wire n_1356;
wire n_910;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1302;
wire n_205;
wire n_1136;
wire n_1313;
wire n_1491;
wire n_754;
wire n_1496;
wire n_179;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_735;
wire n_232;
wire n_1109;
wire n_895;
wire n_1310;
wire n_202;
wire n_427;
wire n_1399;
wire n_1543;
wire n_791;
wire n_732;
wire n_1533;
wire n_193;
wire n_808;
wire n_797;
wire n_1025;
wire n_500;
wire n_1067;
wire n_435;
wire n_766;
wire n_1457;
wire n_541;
wire n_538;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_594;
wire n_200;
wire n_1291;
wire n_1297;
wire n_1155;
wire n_1418;
wire n_1524;
wire n_1689;
wire n_1485;
wire n_1011;
wire n_1184;
wire n_985;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_1352;
wire n_626;
wire n_1650;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_1170;
wire n_305;
wire n_676;
wire n_294;
wire n_318;
wire n_653;
wire n_642;
wire n_1602;
wire n_194;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_268;
wire n_664;
wire n_503;
wire n_235;
wire n_1372;
wire n_605;
wire n_1273;
wire n_353;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_1282;
wire n_1318;
wire n_780;
wire n_998;
wire n_1454;
wire n_467;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_501;
wire n_823;
wire n_245;
wire n_725;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_672;
wire n_581;
wire n_382;
wire n_554;
wire n_1625;
wire n_898;
wire n_1013;
wire n_1452;
wire n_718;
wire n_265;
wire n_1120;
wire n_719;
wire n_443;
wire n_198;
wire n_714;
wire n_1683;
wire n_909;
wire n_1530;
wire n_1497;
wire n_997;
wire n_932;
wire n_612;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_508;
wire n_506;
wire n_1320;
wire n_1663;
wire n_737;
wire n_986;
wire n_509;
wire n_1317;
wire n_1518;
wire n_1281;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_209;
wire n_1564;
wire n_1613;
wire n_733;
wire n_1489;
wire n_1376;
wire n_941;
wire n_981;
wire n_1569;
wire n_867;
wire n_186;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_298;
wire n_518;
wire n_505;
wire n_282;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1620;
wire n_381;
wire n_220;
wire n_390;
wire n_1330;
wire n_481;
wire n_1675;
wire n_1554;
wire n_769;
wire n_1046;
wire n_271;
wire n_934;
wire n_1618;
wire n_826;
wire n_886;
wire n_1221;
wire n_654;
wire n_1172;
wire n_379;
wire n_428;
wire n_1341;
wire n_570;
wire n_1641;
wire n_1361;
wire n_853;
wire n_377;
wire n_751;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_392;
wire n_704;
wire n_787;
wire n_961;
wire n_771;
wire n_276;
wire n_1225;
wire n_1520;
wire n_169;
wire n_522;
wire n_1287;
wire n_1262;
wire n_400;
wire n_930;
wire n_181;
wire n_1411;
wire n_221;
wire n_622;
wire n_1577;
wire n_1087;
wire n_386;
wire n_994;
wire n_848;
wire n_1550;
wire n_1498;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1567;
wire n_1247;
wire n_922;
wire n_816;
wire n_1648;
wire n_591;
wire n_1536;
wire n_1344;
wire n_313;
wire n_631;
wire n_479;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_432;
wire n_839;
wire n_1210;
wire n_1364;
wire n_328;
wire n_1250;
wire n_369;
wire n_871;
wire n_598;
wire n_685;
wire n_928;
wire n_608;
wire n_1367;
wire n_1460;
wire n_772;
wire n_1555;
wire n_499;
wire n_1589;
wire n_517;
wire n_413;
wire n_402;
wire n_1086;
wire n_796;
wire n_1619;
wire n_236;
wire n_1502;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_903;
wire n_1525;
wire n_740;
wire n_203;
wire n_384;
wire n_1404;
wire n_1315;
wire n_277;
wire n_1061;
wire n_333;
wire n_1298;
wire n_1652;
wire n_462;
wire n_1193;
wire n_1676;
wire n_1255;
wire n_258;
wire n_1113;
wire n_1226;
wire n_722;
wire n_1277;
wire n_188;
wire n_844;
wire n_201;
wire n_471;
wire n_852;
wire n_1487;
wire n_1028;
wire n_1601;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_1546;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_1627;
wire n_1245;
wire n_846;
wire n_1673;
wire n_465;
wire n_362;
wire n_1321;
wire n_170;
wire n_273;
wire n_585;
wire n_270;
wire n_616;
wire n_745;
wire n_1654;
wire n_1103;
wire n_648;
wire n_1379;
wire n_312;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_494;
wire n_641;
wire n_730;
wire n_1325;
wire n_1595;
wire n_354;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_695;
wire n_180;
wire n_656;
wire n_1606;
wire n_1220;
wire n_1540;
wire n_229;
wire n_437;
wire n_1642;
wire n_403;
wire n_453;
wire n_1130;
wire n_720;
wire n_1526;
wire n_863;
wire n_805;
wire n_1604;
wire n_1275;
wire n_712;
wire n_246;
wire n_1583;
wire n_1042;
wire n_1402;
wire n_269;
wire n_285;
wire n_412;
wire n_1493;
wire n_657;
wire n_644;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_1621;
wire n_251;
wire n_566;
wire n_565;
wire n_1448;
wire n_1507;
wire n_1398;
wire n_597;
wire n_1181;
wire n_1505;
wire n_1634;
wire n_1196;
wire n_651;
wire n_1340;
wire n_334;
wire n_811;
wire n_1558;
wire n_807;
wire n_835;
wire n_175;
wire n_666;
wire n_262;
wire n_1433;
wire n_1254;
wire n_1026;
wire n_1234;
wire n_319;
wire n_364;
wire n_1138;
wire n_927;
wire n_1089;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_242;
wire n_1681;
wire n_1018;
wire n_438;
wire n_713;
wire n_904;
wire n_1588;
wire n_1622;
wire n_1180;
wire n_1271;
wire n_533;
wire n_1542;
wire n_1251;
wire n_278;

INVx1_ASAP7_75t_L g168 ( 
.A(n_128),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_108),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_84),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_75),
.Y(n_171)
);

CKINVDCx16_ASAP7_75t_R g172 ( 
.A(n_73),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_11),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_60),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_9),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_18),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_92),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_79),
.Y(n_178)
);

BUFx3_ASAP7_75t_L g179 ( 
.A(n_150),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_20),
.Y(n_180)
);

BUFx6f_ASAP7_75t_L g181 ( 
.A(n_143),
.Y(n_181)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_20),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_24),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_103),
.Y(n_184)
);

BUFx10_ASAP7_75t_L g185 ( 
.A(n_124),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_107),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_17),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_30),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_89),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_114),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_105),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_134),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_130),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_87),
.Y(n_194)
);

BUFx2_ASAP7_75t_L g195 ( 
.A(n_110),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_122),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_167),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_47),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_93),
.Y(n_199)
);

CKINVDCx16_ASAP7_75t_R g200 ( 
.A(n_19),
.Y(n_200)
);

INVx1_ASAP7_75t_SL g201 ( 
.A(n_5),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_163),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_60),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_7),
.Y(n_204)
);

BUFx6f_ASAP7_75t_L g205 ( 
.A(n_29),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_99),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_145),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_44),
.Y(n_208)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_152),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_141),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_11),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_151),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_142),
.Y(n_213)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_136),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_3),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_50),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_32),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_54),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_61),
.Y(n_219)
);

BUFx2_ASAP7_75t_L g220 ( 
.A(n_80),
.Y(n_220)
);

BUFx10_ASAP7_75t_L g221 ( 
.A(n_147),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_12),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_48),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_12),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_121),
.Y(n_225)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_81),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_86),
.Y(n_227)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_3),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_159),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_71),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_111),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_120),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_33),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_18),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_115),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_9),
.Y(n_236)
);

BUFx3_ASAP7_75t_L g237 ( 
.A(n_35),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_102),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_45),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_39),
.Y(n_240)
);

INVx2_ASAP7_75t_SL g241 ( 
.A(n_54),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_138),
.Y(n_242)
);

HB1xp67_ASAP7_75t_L g243 ( 
.A(n_94),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_135),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_41),
.Y(n_245)
);

INVxp67_ASAP7_75t_SL g246 ( 
.A(n_1),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_66),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_117),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_10),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_52),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_95),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_65),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_32),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_4),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_56),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_63),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_6),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_83),
.Y(n_258)
);

BUFx3_ASAP7_75t_L g259 ( 
.A(n_56),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_17),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_100),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_15),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_34),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_25),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_36),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_68),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_165),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_47),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_43),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_161),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_13),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_162),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_125),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_90),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_19),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_156),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_67),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_50),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_118),
.Y(n_279)
);

INVx1_ASAP7_75t_SL g280 ( 
.A(n_144),
.Y(n_280)
);

BUFx2_ASAP7_75t_L g281 ( 
.A(n_97),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_57),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_149),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_98),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_85),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_146),
.Y(n_286)
);

INVx1_ASAP7_75t_SL g287 ( 
.A(n_129),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_123),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_72),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_21),
.Y(n_290)
);

BUFx8_ASAP7_75t_SL g291 ( 
.A(n_30),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_43),
.Y(n_292)
);

BUFx10_ASAP7_75t_L g293 ( 
.A(n_27),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_8),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_116),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_158),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_119),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_160),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_77),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_137),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g301 ( 
.A(n_133),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_88),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_78),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_139),
.Y(n_304)
);

CKINVDCx20_ASAP7_75t_R g305 ( 
.A(n_37),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_155),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_53),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_2),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_132),
.Y(n_309)
);

HB1xp67_ASAP7_75t_L g310 ( 
.A(n_59),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_49),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_53),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_157),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_96),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_23),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_42),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_14),
.Y(n_317)
);

BUFx10_ASAP7_75t_L g318 ( 
.A(n_164),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_0),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_16),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_39),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_51),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_104),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g324 ( 
.A(n_21),
.Y(n_324)
);

CKINVDCx16_ASAP7_75t_R g325 ( 
.A(n_42),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_13),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g327 ( 
.A(n_74),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_33),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_52),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_15),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_109),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_131),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_57),
.Y(n_333)
);

INVx1_ASAP7_75t_SL g334 ( 
.A(n_10),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_35),
.Y(n_335)
);

INVx2_ASAP7_75t_L g336 ( 
.A(n_148),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_291),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_205),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_169),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_205),
.Y(n_340)
);

CKINVDCx20_ASAP7_75t_R g341 ( 
.A(n_202),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_170),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_205),
.Y(n_343)
);

INVxp67_ASAP7_75t_L g344 ( 
.A(n_310),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_171),
.Y(n_345)
);

INVxp33_ASAP7_75t_L g346 ( 
.A(n_180),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_177),
.Y(n_347)
);

CKINVDCx20_ASAP7_75t_R g348 ( 
.A(n_247),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_186),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_205),
.Y(n_350)
);

CKINVDCx20_ASAP7_75t_R g351 ( 
.A(n_279),
.Y(n_351)
);

INVxp33_ASAP7_75t_SL g352 ( 
.A(n_173),
.Y(n_352)
);

CKINVDCx16_ASAP7_75t_R g353 ( 
.A(n_200),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_205),
.Y(n_354)
);

CKINVDCx20_ASAP7_75t_R g355 ( 
.A(n_301),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_205),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_182),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_182),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_228),
.Y(n_359)
);

OR2x2_ASAP7_75t_L g360 ( 
.A(n_180),
.B(n_0),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_189),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_190),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_228),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_259),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_191),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_259),
.Y(n_366)
);

CKINVDCx20_ASAP7_75t_R g367 ( 
.A(n_327),
.Y(n_367)
);

NOR2xp33_ASAP7_75t_L g368 ( 
.A(n_195),
.B(n_1),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_192),
.Y(n_369)
);

CKINVDCx20_ASAP7_75t_R g370 ( 
.A(n_172),
.Y(n_370)
);

BUFx2_ASAP7_75t_L g371 ( 
.A(n_259),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_203),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_196),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_203),
.Y(n_374)
);

INVxp67_ASAP7_75t_SL g375 ( 
.A(n_243),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_215),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_197),
.Y(n_377)
);

INVxp67_ASAP7_75t_SL g378 ( 
.A(n_195),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_215),
.Y(n_379)
);

CKINVDCx20_ASAP7_75t_R g380 ( 
.A(n_172),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_220),
.B(n_281),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_217),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_217),
.Y(n_383)
);

NOR2xp33_ASAP7_75t_L g384 ( 
.A(n_220),
.B(n_2),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_206),
.Y(n_385)
);

HB1xp67_ASAP7_75t_L g386 ( 
.A(n_200),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_222),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_222),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_210),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_281),
.B(n_5),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_223),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_223),
.Y(n_392)
);

AND2x2_ASAP7_75t_L g393 ( 
.A(n_237),
.B(n_325),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_233),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_233),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_212),
.Y(n_396)
);

INVxp67_ASAP7_75t_L g397 ( 
.A(n_236),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_213),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_236),
.Y(n_399)
);

INVxp67_ASAP7_75t_L g400 ( 
.A(n_249),
.Y(n_400)
);

INVx1_ASAP7_75t_SL g401 ( 
.A(n_305),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_225),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_249),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_227),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_250),
.Y(n_405)
);

INVxp33_ASAP7_75t_SL g406 ( 
.A(n_174),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_250),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_229),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_260),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_260),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_231),
.Y(n_411)
);

NOR2xp33_ASAP7_75t_L g412 ( 
.A(n_168),
.B(n_6),
.Y(n_412)
);

CKINVDCx20_ASAP7_75t_R g413 ( 
.A(n_232),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_235),
.Y(n_414)
);

CKINVDCx20_ASAP7_75t_R g415 ( 
.A(n_244),
.Y(n_415)
);

INVxp67_ASAP7_75t_SL g416 ( 
.A(n_179),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_262),
.Y(n_417)
);

NOR2xp33_ASAP7_75t_L g418 ( 
.A(n_168),
.B(n_8),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_262),
.Y(n_419)
);

CKINVDCx20_ASAP7_75t_R g420 ( 
.A(n_248),
.Y(n_420)
);

INVxp67_ASAP7_75t_SL g421 ( 
.A(n_179),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_252),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_256),
.Y(n_423)
);

INVxp67_ASAP7_75t_L g424 ( 
.A(n_263),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_263),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_258),
.Y(n_426)
);

HB1xp67_ASAP7_75t_L g427 ( 
.A(n_325),
.Y(n_427)
);

BUFx3_ASAP7_75t_L g428 ( 
.A(n_364),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_338),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_338),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_340),
.Y(n_431)
);

INVx3_ASAP7_75t_L g432 ( 
.A(n_340),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_339),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_343),
.Y(n_434)
);

AND2x4_ASAP7_75t_L g435 ( 
.A(n_343),
.B(n_179),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_350),
.Y(n_436)
);

CKINVDCx20_ASAP7_75t_R g437 ( 
.A(n_341),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_350),
.Y(n_438)
);

INVx2_ASAP7_75t_L g439 ( 
.A(n_354),
.Y(n_439)
);

AND2x2_ASAP7_75t_L g440 ( 
.A(n_416),
.B(n_237),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_354),
.Y(n_441)
);

BUFx2_ASAP7_75t_L g442 ( 
.A(n_370),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_356),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_356),
.Y(n_444)
);

CKINVDCx5p33_ASAP7_75t_R g445 ( 
.A(n_342),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_372),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_372),
.Y(n_447)
);

CKINVDCx5p33_ASAP7_75t_R g448 ( 
.A(n_345),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_374),
.Y(n_449)
);

BUFx6f_ASAP7_75t_L g450 ( 
.A(n_357),
.Y(n_450)
);

CKINVDCx5p33_ASAP7_75t_R g451 ( 
.A(n_347),
.Y(n_451)
);

INVxp67_ASAP7_75t_L g452 ( 
.A(n_386),
.Y(n_452)
);

INVx2_ASAP7_75t_L g453 ( 
.A(n_357),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_374),
.Y(n_454)
);

CKINVDCx5p33_ASAP7_75t_R g455 ( 
.A(n_349),
.Y(n_455)
);

INVx3_ASAP7_75t_L g456 ( 
.A(n_358),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_376),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_376),
.Y(n_458)
);

BUFx6f_ASAP7_75t_L g459 ( 
.A(n_358),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_379),
.Y(n_460)
);

NOR2xp33_ASAP7_75t_SL g461 ( 
.A(n_368),
.B(n_293),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_361),
.B(n_362),
.Y(n_462)
);

BUFx3_ASAP7_75t_L g463 ( 
.A(n_364),
.Y(n_463)
);

CKINVDCx5p33_ASAP7_75t_R g464 ( 
.A(n_365),
.Y(n_464)
);

CKINVDCx5p33_ASAP7_75t_R g465 ( 
.A(n_369),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_379),
.Y(n_466)
);

HB1xp67_ASAP7_75t_L g467 ( 
.A(n_427),
.Y(n_467)
);

INVx2_ASAP7_75t_L g468 ( 
.A(n_359),
.Y(n_468)
);

NAND3xp33_ASAP7_75t_L g469 ( 
.A(n_381),
.B(n_275),
.C(n_271),
.Y(n_469)
);

INVxp67_ASAP7_75t_L g470 ( 
.A(n_393),
.Y(n_470)
);

HB1xp67_ASAP7_75t_L g471 ( 
.A(n_401),
.Y(n_471)
);

INVx2_ASAP7_75t_L g472 ( 
.A(n_363),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_382),
.Y(n_473)
);

CKINVDCx5p33_ASAP7_75t_R g474 ( 
.A(n_373),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_SL g475 ( 
.A(n_353),
.B(n_185),
.Y(n_475)
);

HB1xp67_ASAP7_75t_L g476 ( 
.A(n_377),
.Y(n_476)
);

CKINVDCx5p33_ASAP7_75t_R g477 ( 
.A(n_385),
.Y(n_477)
);

CKINVDCx8_ASAP7_75t_R g478 ( 
.A(n_337),
.Y(n_478)
);

CKINVDCx5p33_ASAP7_75t_R g479 ( 
.A(n_389),
.Y(n_479)
);

BUFx6f_ASAP7_75t_L g480 ( 
.A(n_363),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_L g481 ( 
.A(n_396),
.B(n_209),
.Y(n_481)
);

CKINVDCx5p33_ASAP7_75t_R g482 ( 
.A(n_398),
.Y(n_482)
);

NOR2xp33_ASAP7_75t_R g483 ( 
.A(n_413),
.B(n_261),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_L g484 ( 
.A(n_421),
.B(n_266),
.Y(n_484)
);

INVxp67_ASAP7_75t_L g485 ( 
.A(n_393),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_382),
.Y(n_486)
);

INVx2_ASAP7_75t_L g487 ( 
.A(n_383),
.Y(n_487)
);

BUFx6f_ASAP7_75t_L g488 ( 
.A(n_387),
.Y(n_488)
);

INVx2_ASAP7_75t_L g489 ( 
.A(n_387),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_L g490 ( 
.A(n_366),
.B(n_270),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_388),
.Y(n_491)
);

CKINVDCx5p33_ASAP7_75t_R g492 ( 
.A(n_402),
.Y(n_492)
);

INVx1_ASAP7_75t_SL g493 ( 
.A(n_380),
.Y(n_493)
);

AND2x4_ASAP7_75t_L g494 ( 
.A(n_366),
.B(n_209),
.Y(n_494)
);

INVx2_ASAP7_75t_L g495 ( 
.A(n_388),
.Y(n_495)
);

CKINVDCx5p33_ASAP7_75t_R g496 ( 
.A(n_404),
.Y(n_496)
);

AND2x2_ASAP7_75t_SL g497 ( 
.A(n_384),
.B(n_181),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_391),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_391),
.Y(n_499)
);

INVx2_ASAP7_75t_L g500 ( 
.A(n_392),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_392),
.Y(n_501)
);

INVxp67_ASAP7_75t_L g502 ( 
.A(n_371),
.Y(n_502)
);

CKINVDCx5p33_ASAP7_75t_R g503 ( 
.A(n_408),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_394),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_L g505 ( 
.A(n_484),
.B(n_411),
.Y(n_505)
);

INVx2_ASAP7_75t_L g506 ( 
.A(n_439),
.Y(n_506)
);

INVx3_ASAP7_75t_L g507 ( 
.A(n_432),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_428),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_428),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_L g510 ( 
.A(n_484),
.B(n_414),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_L g511 ( 
.A(n_481),
.B(n_422),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_L g512 ( 
.A(n_490),
.B(n_423),
.Y(n_512)
);

INVx5_ASAP7_75t_L g513 ( 
.A(n_432),
.Y(n_513)
);

NOR2xp33_ASAP7_75t_L g514 ( 
.A(n_461),
.B(n_352),
.Y(n_514)
);

INVx4_ASAP7_75t_SL g515 ( 
.A(n_435),
.Y(n_515)
);

INVx2_ASAP7_75t_L g516 ( 
.A(n_439),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_L g517 ( 
.A(n_490),
.B(n_426),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_463),
.Y(n_518)
);

INVx2_ASAP7_75t_L g519 ( 
.A(n_429),
.Y(n_519)
);

INVx2_ASAP7_75t_L g520 ( 
.A(n_429),
.Y(n_520)
);

AND2x4_ASAP7_75t_L g521 ( 
.A(n_435),
.B(n_178),
.Y(n_521)
);

AND2x2_ASAP7_75t_L g522 ( 
.A(n_440),
.B(n_378),
.Y(n_522)
);

NOR2xp33_ASAP7_75t_L g523 ( 
.A(n_461),
.B(n_406),
.Y(n_523)
);

AOI22xp33_ASAP7_75t_L g524 ( 
.A1(n_497),
.A2(n_390),
.B1(n_418),
.B2(n_412),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_463),
.Y(n_525)
);

AND2x4_ASAP7_75t_L g526 ( 
.A(n_435),
.B(n_178),
.Y(n_526)
);

CKINVDCx20_ASAP7_75t_R g527 ( 
.A(n_437),
.Y(n_527)
);

AND2x6_ASAP7_75t_L g528 ( 
.A(n_440),
.B(n_181),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_L g529 ( 
.A(n_497),
.B(n_375),
.Y(n_529)
);

INVx1_ASAP7_75t_SL g530 ( 
.A(n_471),
.Y(n_530)
);

BUFx10_ASAP7_75t_L g531 ( 
.A(n_433),
.Y(n_531)
);

BUFx4f_ASAP7_75t_L g532 ( 
.A(n_497),
.Y(n_532)
);

INVx5_ASAP7_75t_L g533 ( 
.A(n_432),
.Y(n_533)
);

NOR2xp33_ASAP7_75t_L g534 ( 
.A(n_462),
.B(n_415),
.Y(n_534)
);

INVx2_ASAP7_75t_L g535 ( 
.A(n_430),
.Y(n_535)
);

AO22x2_ASAP7_75t_L g536 ( 
.A1(n_469),
.A2(n_360),
.B1(n_241),
.B2(n_275),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_L g537 ( 
.A(n_463),
.B(n_280),
.Y(n_537)
);

INVx6_ASAP7_75t_L g538 ( 
.A(n_494),
.Y(n_538)
);

INVx2_ASAP7_75t_L g539 ( 
.A(n_430),
.Y(n_539)
);

BUFx2_ASAP7_75t_L g540 ( 
.A(n_502),
.Y(n_540)
);

BUFx3_ASAP7_75t_L g541 ( 
.A(n_494),
.Y(n_541)
);

AOI22xp33_ASAP7_75t_L g542 ( 
.A1(n_469),
.A2(n_360),
.B1(n_241),
.B2(n_344),
.Y(n_542)
);

NOR2xp33_ASAP7_75t_L g543 ( 
.A(n_470),
.B(n_420),
.Y(n_543)
);

BUFx2_ASAP7_75t_L g544 ( 
.A(n_467),
.Y(n_544)
);

INVx2_ASAP7_75t_L g545 ( 
.A(n_431),
.Y(n_545)
);

CKINVDCx20_ASAP7_75t_R g546 ( 
.A(n_442),
.Y(n_546)
);

INVx5_ASAP7_75t_L g547 ( 
.A(n_432),
.Y(n_547)
);

INVx3_ASAP7_75t_L g548 ( 
.A(n_488),
.Y(n_548)
);

BUFx3_ASAP7_75t_L g549 ( 
.A(n_494),
.Y(n_549)
);

NOR2xp33_ASAP7_75t_L g550 ( 
.A(n_485),
.B(n_371),
.Y(n_550)
);

AOI21x1_ASAP7_75t_L g551 ( 
.A1(n_431),
.A2(n_193),
.B(n_184),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_L g552 ( 
.A(n_434),
.B(n_287),
.Y(n_552)
);

NOR2xp33_ASAP7_75t_L g553 ( 
.A(n_445),
.B(n_346),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_488),
.Y(n_554)
);

INVx2_ASAP7_75t_L g555 ( 
.A(n_434),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_SL g556 ( 
.A(n_448),
.B(n_185),
.Y(n_556)
);

CKINVDCx5p33_ASAP7_75t_R g557 ( 
.A(n_483),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_488),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_SL g559 ( 
.A(n_451),
.B(n_185),
.Y(n_559)
);

INVx2_ASAP7_75t_L g560 ( 
.A(n_436),
.Y(n_560)
);

INVx2_ASAP7_75t_L g561 ( 
.A(n_436),
.Y(n_561)
);

NAND3xp33_ASAP7_75t_L g562 ( 
.A(n_452),
.B(n_400),
.C(n_397),
.Y(n_562)
);

INVx2_ASAP7_75t_L g563 ( 
.A(n_438),
.Y(n_563)
);

AND2x2_ASAP7_75t_SL g564 ( 
.A(n_494),
.B(n_214),
.Y(n_564)
);

INVx6_ASAP7_75t_L g565 ( 
.A(n_488),
.Y(n_565)
);

BUFx3_ASAP7_75t_L g566 ( 
.A(n_441),
.Y(n_566)
);

BUFx4f_ASAP7_75t_L g567 ( 
.A(n_450),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_L g568 ( 
.A(n_441),
.B(n_272),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_SL g569 ( 
.A(n_455),
.B(n_185),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_443),
.Y(n_570)
);

BUFx8_ASAP7_75t_SL g571 ( 
.A(n_442),
.Y(n_571)
);

AND2x2_ASAP7_75t_L g572 ( 
.A(n_446),
.B(n_394),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_L g573 ( 
.A(n_443),
.B(n_273),
.Y(n_573)
);

INVx2_ASAP7_75t_L g574 ( 
.A(n_444),
.Y(n_574)
);

BUFx6f_ASAP7_75t_L g575 ( 
.A(n_450),
.Y(n_575)
);

AND2x2_ASAP7_75t_L g576 ( 
.A(n_446),
.B(n_395),
.Y(n_576)
);

AND3x2_ASAP7_75t_L g577 ( 
.A(n_476),
.B(n_226),
.C(n_214),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_444),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_L g579 ( 
.A(n_447),
.B(n_274),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_447),
.Y(n_580)
);

OR2x6_ASAP7_75t_L g581 ( 
.A(n_475),
.B(n_424),
.Y(n_581)
);

BUFx2_ASAP7_75t_L g582 ( 
.A(n_493),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_449),
.Y(n_583)
);

INVx2_ASAP7_75t_L g584 ( 
.A(n_450),
.Y(n_584)
);

INVx2_ASAP7_75t_L g585 ( 
.A(n_450),
.Y(n_585)
);

INVx3_ASAP7_75t_L g586 ( 
.A(n_459),
.Y(n_586)
);

INVx3_ASAP7_75t_L g587 ( 
.A(n_459),
.Y(n_587)
);

INVx2_ASAP7_75t_L g588 ( 
.A(n_459),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_L g589 ( 
.A(n_454),
.B(n_277),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_454),
.Y(n_590)
);

AOI22xp33_ASAP7_75t_L g591 ( 
.A1(n_457),
.A2(n_320),
.B1(n_292),
.B2(n_271),
.Y(n_591)
);

INVx2_ASAP7_75t_L g592 ( 
.A(n_459),
.Y(n_592)
);

INVx2_ASAP7_75t_L g593 ( 
.A(n_459),
.Y(n_593)
);

INVx1_ASAP7_75t_SL g594 ( 
.A(n_493),
.Y(n_594)
);

BUFx10_ASAP7_75t_L g595 ( 
.A(n_464),
.Y(n_595)
);

OR2x2_ASAP7_75t_L g596 ( 
.A(n_458),
.B(n_201),
.Y(n_596)
);

INVx4_ASAP7_75t_SL g597 ( 
.A(n_480),
.Y(n_597)
);

BUFx3_ASAP7_75t_L g598 ( 
.A(n_460),
.Y(n_598)
);

AND2x2_ASAP7_75t_L g599 ( 
.A(n_466),
.B(n_395),
.Y(n_599)
);

AND2x2_ASAP7_75t_L g600 ( 
.A(n_466),
.B(n_399),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_L g601 ( 
.A(n_473),
.B(n_486),
.Y(n_601)
);

BUFx3_ASAP7_75t_L g602 ( 
.A(n_473),
.Y(n_602)
);

AO21x2_ASAP7_75t_L g603 ( 
.A1(n_486),
.A2(n_193),
.B(n_184),
.Y(n_603)
);

BUFx2_ASAP7_75t_L g604 ( 
.A(n_465),
.Y(n_604)
);

INVx4_ASAP7_75t_SL g605 ( 
.A(n_480),
.Y(n_605)
);

BUFx2_ASAP7_75t_L g606 ( 
.A(n_474),
.Y(n_606)
);

INVx5_ASAP7_75t_L g607 ( 
.A(n_480),
.Y(n_607)
);

OR2x2_ASAP7_75t_L g608 ( 
.A(n_491),
.B(n_334),
.Y(n_608)
);

BUFx10_ASAP7_75t_L g609 ( 
.A(n_477),
.Y(n_609)
);

NOR2xp33_ASAP7_75t_L g610 ( 
.A(n_479),
.B(n_348),
.Y(n_610)
);

AND2x6_ASAP7_75t_L g611 ( 
.A(n_491),
.B(n_181),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_L g612 ( 
.A(n_498),
.B(n_499),
.Y(n_612)
);

INVxp67_ASAP7_75t_L g613 ( 
.A(n_498),
.Y(n_613)
);

BUFx6f_ASAP7_75t_L g614 ( 
.A(n_487),
.Y(n_614)
);

CKINVDCx5p33_ASAP7_75t_R g615 ( 
.A(n_482),
.Y(n_615)
);

INVxp67_ASAP7_75t_L g616 ( 
.A(n_499),
.Y(n_616)
);

INVx2_ASAP7_75t_L g617 ( 
.A(n_456),
.Y(n_617)
);

NOR2xp33_ASAP7_75t_L g618 ( 
.A(n_492),
.B(n_351),
.Y(n_618)
);

INVx2_ASAP7_75t_L g619 ( 
.A(n_456),
.Y(n_619)
);

HAxp5_ASAP7_75t_SL g620 ( 
.A(n_501),
.B(n_282),
.CON(n_620),
.SN(n_620)
);

CKINVDCx5p33_ASAP7_75t_R g621 ( 
.A(n_496),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_L g622 ( 
.A(n_504),
.B(n_284),
.Y(n_622)
);

BUFx3_ASAP7_75t_L g623 ( 
.A(n_504),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_487),
.Y(n_624)
);

CKINVDCx5p33_ASAP7_75t_R g625 ( 
.A(n_503),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_487),
.Y(n_626)
);

BUFx3_ASAP7_75t_L g627 ( 
.A(n_489),
.Y(n_627)
);

NAND2xp33_ASAP7_75t_SL g628 ( 
.A(n_489),
.B(n_311),
.Y(n_628)
);

BUFx10_ASAP7_75t_L g629 ( 
.A(n_478),
.Y(n_629)
);

BUFx2_ASAP7_75t_L g630 ( 
.A(n_489),
.Y(n_630)
);

INVx2_ASAP7_75t_L g631 ( 
.A(n_456),
.Y(n_631)
);

INVx5_ASAP7_75t_L g632 ( 
.A(n_495),
.Y(n_632)
);

AND2x4_ASAP7_75t_L g633 ( 
.A(n_495),
.B(n_194),
.Y(n_633)
);

BUFx2_ASAP7_75t_L g634 ( 
.A(n_500),
.Y(n_634)
);

AOI22xp33_ASAP7_75t_L g635 ( 
.A1(n_500),
.A2(n_320),
.B1(n_292),
.B2(n_282),
.Y(n_635)
);

NOR2xp33_ASAP7_75t_SL g636 ( 
.A(n_478),
.B(n_355),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_SL g637 ( 
.A(n_532),
.B(n_181),
.Y(n_637)
);

INVx2_ASAP7_75t_L g638 ( 
.A(n_627),
.Y(n_638)
);

NOR2xp33_ASAP7_75t_L g639 ( 
.A(n_512),
.B(n_175),
.Y(n_639)
);

AOI22xp5_ASAP7_75t_L g640 ( 
.A1(n_529),
.A2(n_367),
.B1(n_286),
.B2(n_288),
.Y(n_640)
);

INVxp67_ASAP7_75t_L g641 ( 
.A(n_530),
.Y(n_641)
);

AOI22xp5_ASAP7_75t_L g642 ( 
.A1(n_514),
.A2(n_297),
.B1(n_289),
.B2(n_332),
.Y(n_642)
);

INVx8_ASAP7_75t_L g643 ( 
.A(n_581),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_L g644 ( 
.A(n_564),
.B(n_194),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_L g645 ( 
.A(n_564),
.B(n_199),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_L g646 ( 
.A(n_564),
.B(n_199),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_541),
.Y(n_647)
);

NOR2xp33_ASAP7_75t_L g648 ( 
.A(n_517),
.B(n_176),
.Y(n_648)
);

INVx2_ASAP7_75t_L g649 ( 
.A(n_506),
.Y(n_649)
);

NOR2xp67_ASAP7_75t_L g650 ( 
.A(n_557),
.B(n_296),
.Y(n_650)
);

INVxp67_ASAP7_75t_SL g651 ( 
.A(n_630),
.Y(n_651)
);

OR2x2_ASAP7_75t_L g652 ( 
.A(n_596),
.B(n_246),
.Y(n_652)
);

AOI22xp5_ASAP7_75t_L g653 ( 
.A1(n_523),
.A2(n_304),
.B1(n_298),
.B2(n_299),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_SL g654 ( 
.A(n_532),
.B(n_181),
.Y(n_654)
);

AO221x1_ASAP7_75t_L g655 ( 
.A1(n_536),
.A2(n_181),
.B1(n_307),
.B2(n_317),
.C(n_329),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_L g656 ( 
.A(n_634),
.B(n_207),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_SL g657 ( 
.A(n_553),
.B(n_303),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_549),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_549),
.Y(n_659)
);

AOI22xp5_ASAP7_75t_L g660 ( 
.A1(n_532),
.A2(n_309),
.B1(n_314),
.B2(n_331),
.Y(n_660)
);

NAND2x1p5_ASAP7_75t_L g661 ( 
.A(n_634),
.B(n_230),
.Y(n_661)
);

OR2x6_ASAP7_75t_L g662 ( 
.A(n_582),
.B(n_307),
.Y(n_662)
);

NOR2xp67_ASAP7_75t_SL g663 ( 
.A(n_538),
.B(n_230),
.Y(n_663)
);

NAND2xp33_ASAP7_75t_L g664 ( 
.A(n_524),
.B(n_226),
.Y(n_664)
);

OAI22xp33_ASAP7_75t_L g665 ( 
.A1(n_581),
.A2(n_317),
.B1(n_329),
.B2(n_324),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_508),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_L g667 ( 
.A(n_508),
.B(n_238),
.Y(n_667)
);

INVx2_ASAP7_75t_SL g668 ( 
.A(n_596),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_L g669 ( 
.A(n_509),
.B(n_238),
.Y(n_669)
);

INVx2_ASAP7_75t_SL g670 ( 
.A(n_608),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_L g671 ( 
.A(n_509),
.B(n_242),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_L g672 ( 
.A(n_518),
.B(n_242),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_L g673 ( 
.A(n_518),
.B(n_251),
.Y(n_673)
);

BUFx6f_ASAP7_75t_L g674 ( 
.A(n_598),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_L g675 ( 
.A(n_525),
.B(n_251),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_SL g676 ( 
.A(n_522),
.B(n_221),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_525),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_L g678 ( 
.A(n_505),
.B(n_510),
.Y(n_678)
);

AND2x2_ASAP7_75t_SL g679 ( 
.A(n_521),
.B(n_336),
.Y(n_679)
);

INVx2_ASAP7_75t_L g680 ( 
.A(n_516),
.Y(n_680)
);

AND2x6_ASAP7_75t_SL g681 ( 
.A(n_610),
.B(n_399),
.Y(n_681)
);

OR2x2_ASAP7_75t_L g682 ( 
.A(n_608),
.B(n_403),
.Y(n_682)
);

AOI22xp33_ASAP7_75t_L g683 ( 
.A1(n_536),
.A2(n_276),
.B1(n_306),
.B2(n_302),
.Y(n_683)
);

BUFx6f_ASAP7_75t_L g684 ( 
.A(n_598),
.Y(n_684)
);

AOI22xp33_ASAP7_75t_L g685 ( 
.A1(n_536),
.A2(n_276),
.B1(n_306),
.B2(n_302),
.Y(n_685)
);

BUFx2_ASAP7_75t_L g686 ( 
.A(n_582),
.Y(n_686)
);

OR2x2_ASAP7_75t_L g687 ( 
.A(n_544),
.B(n_403),
.Y(n_687)
);

NOR2xp33_ASAP7_75t_L g688 ( 
.A(n_550),
.B(n_183),
.Y(n_688)
);

NOR2xp33_ASAP7_75t_L g689 ( 
.A(n_522),
.B(n_187),
.Y(n_689)
);

OAI22xp5_ASAP7_75t_L g690 ( 
.A1(n_511),
.A2(n_336),
.B1(n_267),
.B2(n_283),
.Y(n_690)
);

AND2x2_ASAP7_75t_L g691 ( 
.A(n_540),
.B(n_293),
.Y(n_691)
);

AOI221xp5_ASAP7_75t_L g692 ( 
.A1(n_542),
.A2(n_218),
.B1(n_211),
.B2(n_208),
.C(n_204),
.Y(n_692)
);

INVxp67_ASAP7_75t_SL g693 ( 
.A(n_601),
.Y(n_693)
);

INVx2_ASAP7_75t_SL g694 ( 
.A(n_544),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_572),
.Y(n_695)
);

INVx3_ASAP7_75t_L g696 ( 
.A(n_538),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_L g697 ( 
.A(n_566),
.B(n_267),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_L g698 ( 
.A(n_580),
.B(n_285),
.Y(n_698)
);

BUFx6f_ASAP7_75t_L g699 ( 
.A(n_602),
.Y(n_699)
);

OAI221xp5_ASAP7_75t_L g700 ( 
.A1(n_591),
.A2(n_635),
.B1(n_613),
.B2(n_616),
.C(n_612),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_L g701 ( 
.A(n_583),
.B(n_285),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_L g702 ( 
.A(n_583),
.B(n_295),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_576),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_SL g704 ( 
.A(n_557),
.B(n_221),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_L g705 ( 
.A(n_590),
.B(n_295),
.Y(n_705)
);

AOI22xp33_ASAP7_75t_L g706 ( 
.A1(n_536),
.A2(n_323),
.B1(n_313),
.B2(n_300),
.Y(n_706)
);

INVx2_ASAP7_75t_L g707 ( 
.A(n_614),
.Y(n_707)
);

NOR2xp33_ASAP7_75t_L g708 ( 
.A(n_537),
.B(n_188),
.Y(n_708)
);

NOR2xp33_ASAP7_75t_L g709 ( 
.A(n_602),
.B(n_198),
.Y(n_709)
);

AOI22xp33_ASAP7_75t_L g710 ( 
.A1(n_603),
.A2(n_300),
.B1(n_313),
.B2(n_323),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_L g711 ( 
.A(n_590),
.B(n_453),
.Y(n_711)
);

NOR2xp33_ASAP7_75t_L g712 ( 
.A(n_623),
.B(n_216),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_599),
.Y(n_713)
);

OR2x6_ASAP7_75t_L g714 ( 
.A(n_604),
.B(n_606),
.Y(n_714)
);

INVx2_ASAP7_75t_L g715 ( 
.A(n_614),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_SL g716 ( 
.A(n_540),
.B(n_221),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_SL g717 ( 
.A(n_534),
.B(n_552),
.Y(n_717)
);

OR2x2_ASAP7_75t_L g718 ( 
.A(n_594),
.B(n_405),
.Y(n_718)
);

AOI21xp5_ASAP7_75t_L g719 ( 
.A1(n_567),
.A2(n_472),
.B(n_468),
.Y(n_719)
);

AOI22xp33_ASAP7_75t_L g720 ( 
.A1(n_603),
.A2(n_293),
.B1(n_417),
.B2(n_425),
.Y(n_720)
);

AND2x2_ASAP7_75t_L g721 ( 
.A(n_604),
.B(n_293),
.Y(n_721)
);

CKINVDCx5p33_ASAP7_75t_R g722 ( 
.A(n_615),
.Y(n_722)
);

NOR2xp33_ASAP7_75t_L g723 ( 
.A(n_623),
.B(n_219),
.Y(n_723)
);

OAI22xp33_ASAP7_75t_L g724 ( 
.A1(n_581),
.A2(n_308),
.B1(n_234),
.B2(n_239),
.Y(n_724)
);

BUFx2_ASAP7_75t_L g725 ( 
.A(n_546),
.Y(n_725)
);

INVx2_ASAP7_75t_L g726 ( 
.A(n_614),
.Y(n_726)
);

BUFx8_ASAP7_75t_L g727 ( 
.A(n_606),
.Y(n_727)
);

O2A1O1Ixp33_ASAP7_75t_L g728 ( 
.A1(n_600),
.A2(n_410),
.B(n_425),
.C(n_419),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_600),
.Y(n_729)
);

NOR2xp33_ASAP7_75t_L g730 ( 
.A(n_579),
.B(n_224),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_L g731 ( 
.A(n_521),
.B(n_472),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_L g732 ( 
.A(n_526),
.B(n_472),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_L g733 ( 
.A(n_526),
.B(n_407),
.Y(n_733)
);

HB1xp67_ASAP7_75t_L g734 ( 
.A(n_603),
.Y(n_734)
);

AOI22xp5_ASAP7_75t_L g735 ( 
.A1(n_538),
.A2(n_318),
.B1(n_240),
.B2(n_290),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_570),
.Y(n_736)
);

INVx2_ASAP7_75t_L g737 ( 
.A(n_614),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_L g738 ( 
.A(n_570),
.B(n_407),
.Y(n_738)
);

NOR2xp33_ASAP7_75t_L g739 ( 
.A(n_589),
.B(n_245),
.Y(n_739)
);

BUFx6f_ASAP7_75t_SL g740 ( 
.A(n_629),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_L g741 ( 
.A(n_578),
.B(n_409),
.Y(n_741)
);

INVx3_ASAP7_75t_L g742 ( 
.A(n_507),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_L g743 ( 
.A(n_578),
.B(n_409),
.Y(n_743)
);

NAND3xp33_ASAP7_75t_L g744 ( 
.A(n_620),
.B(n_294),
.C(n_253),
.Y(n_744)
);

HB1xp67_ASAP7_75t_L g745 ( 
.A(n_581),
.Y(n_745)
);

AOI221xp5_ASAP7_75t_L g746 ( 
.A1(n_628),
.A2(n_312),
.B1(n_255),
.B2(n_257),
.C(n_335),
.Y(n_746)
);

BUFx8_ASAP7_75t_L g747 ( 
.A(n_571),
.Y(n_747)
);

INVx2_ASAP7_75t_L g748 ( 
.A(n_617),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_SL g749 ( 
.A(n_622),
.B(n_254),
.Y(n_749)
);

NOR2xp33_ASAP7_75t_L g750 ( 
.A(n_556),
.B(n_264),
.Y(n_750)
);

INVx4_ASAP7_75t_L g751 ( 
.A(n_515),
.Y(n_751)
);

CKINVDCx5p33_ASAP7_75t_R g752 ( 
.A(n_615),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_507),
.Y(n_753)
);

INVx8_ASAP7_75t_L g754 ( 
.A(n_621),
.Y(n_754)
);

INVx2_ASAP7_75t_SL g755 ( 
.A(n_577),
.Y(n_755)
);

CKINVDCx5p33_ASAP7_75t_R g756 ( 
.A(n_621),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_617),
.Y(n_757)
);

OR2x2_ASAP7_75t_L g758 ( 
.A(n_562),
.B(n_419),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_SL g759 ( 
.A(n_543),
.B(n_265),
.Y(n_759)
);

AOI22xp33_ASAP7_75t_SL g760 ( 
.A1(n_636),
.A2(n_333),
.B1(n_330),
.B2(n_328),
.Y(n_760)
);

NOR2x1p5_ASAP7_75t_L g761 ( 
.A(n_625),
.B(n_268),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_619),
.Y(n_762)
);

CKINVDCx11_ASAP7_75t_R g763 ( 
.A(n_629),
.Y(n_763)
);

NOR2xp33_ASAP7_75t_L g764 ( 
.A(n_559),
.B(n_269),
.Y(n_764)
);

BUFx8_ASAP7_75t_L g765 ( 
.A(n_629),
.Y(n_765)
);

NOR2xp33_ASAP7_75t_L g766 ( 
.A(n_569),
.B(n_278),
.Y(n_766)
);

NOR3xp33_ASAP7_75t_L g767 ( 
.A(n_568),
.B(n_326),
.C(n_322),
.Y(n_767)
);

AOI22xp5_ASAP7_75t_L g768 ( 
.A1(n_573),
.A2(n_321),
.B1(n_319),
.B2(n_316),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_L g769 ( 
.A(n_519),
.B(n_315),
.Y(n_769)
);

AOI22xp33_ASAP7_75t_L g770 ( 
.A1(n_633),
.A2(n_14),
.B1(n_16),
.B2(n_22),
.Y(n_770)
);

AND2x2_ASAP7_75t_L g771 ( 
.A(n_531),
.B(n_22),
.Y(n_771)
);

NAND3xp33_ASAP7_75t_L g772 ( 
.A(n_620),
.B(n_23),
.C(n_24),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_631),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_L g774 ( 
.A(n_693),
.B(n_520),
.Y(n_774)
);

O2A1O1Ixp5_ASAP7_75t_L g775 ( 
.A1(n_637),
.A2(n_551),
.B(n_633),
.C(n_520),
.Y(n_775)
);

INVx2_ASAP7_75t_L g776 ( 
.A(n_638),
.Y(n_776)
);

BUFx2_ASAP7_75t_L g777 ( 
.A(n_686),
.Y(n_777)
);

O2A1O1Ixp33_ASAP7_75t_L g778 ( 
.A1(n_664),
.A2(n_644),
.B(n_646),
.C(n_645),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_666),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_L g780 ( 
.A(n_678),
.B(n_535),
.Y(n_780)
);

OAI21xp5_ASAP7_75t_L g781 ( 
.A1(n_637),
.A2(n_554),
.B(n_558),
.Y(n_781)
);

OAI21xp5_ASAP7_75t_L g782 ( 
.A1(n_654),
.A2(n_554),
.B(n_558),
.Y(n_782)
);

CKINVDCx14_ASAP7_75t_R g783 ( 
.A(n_763),
.Y(n_783)
);

CKINVDCx10_ASAP7_75t_R g784 ( 
.A(n_740),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_L g785 ( 
.A(n_651),
.B(n_535),
.Y(n_785)
);

AND2x2_ASAP7_75t_L g786 ( 
.A(n_668),
.B(n_531),
.Y(n_786)
);

BUFx4f_ASAP7_75t_L g787 ( 
.A(n_754),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_L g788 ( 
.A(n_651),
.B(n_539),
.Y(n_788)
);

NAND3xp33_ASAP7_75t_SL g789 ( 
.A(n_746),
.B(n_546),
.C(n_527),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_L g790 ( 
.A(n_639),
.B(n_648),
.Y(n_790)
);

NOR2xp33_ASAP7_75t_L g791 ( 
.A(n_641),
.B(n_618),
.Y(n_791)
);

INVx4_ASAP7_75t_L g792 ( 
.A(n_674),
.Y(n_792)
);

NOR2xp33_ASAP7_75t_L g793 ( 
.A(n_641),
.B(n_531),
.Y(n_793)
);

BUFx2_ASAP7_75t_L g794 ( 
.A(n_694),
.Y(n_794)
);

NOR2xp33_ASAP7_75t_L g795 ( 
.A(n_717),
.B(n_595),
.Y(n_795)
);

A2O1A1Ixp33_ASAP7_75t_L g796 ( 
.A1(n_648),
.A2(n_633),
.B(n_545),
.C(n_574),
.Y(n_796)
);

OAI21xp5_ASAP7_75t_L g797 ( 
.A1(n_734),
.A2(n_624),
.B(n_626),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_L g798 ( 
.A(n_708),
.B(n_545),
.Y(n_798)
);

OAI21xp5_ASAP7_75t_L g799 ( 
.A1(n_734),
.A2(n_561),
.B(n_563),
.Y(n_799)
);

AOI21xp5_ASAP7_75t_L g800 ( 
.A1(n_731),
.A2(n_588),
.B(n_592),
.Y(n_800)
);

AOI22xp5_ASAP7_75t_L g801 ( 
.A1(n_679),
.A2(n_528),
.B1(n_555),
.B2(n_560),
.Y(n_801)
);

BUFx6f_ASAP7_75t_L g802 ( 
.A(n_674),
.Y(n_802)
);

AOI21xp5_ASAP7_75t_L g803 ( 
.A1(n_732),
.A2(n_593),
.B(n_584),
.Y(n_803)
);

INVx3_ASAP7_75t_SL g804 ( 
.A(n_722),
.Y(n_804)
);

AOI21x1_ASAP7_75t_L g805 ( 
.A1(n_711),
.A2(n_584),
.B(n_593),
.Y(n_805)
);

INVx2_ASAP7_75t_L g806 ( 
.A(n_748),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_L g807 ( 
.A(n_730),
.B(n_528),
.Y(n_807)
);

OR2x6_ASAP7_75t_L g808 ( 
.A(n_754),
.B(n_595),
.Y(n_808)
);

CKINVDCx20_ASAP7_75t_R g809 ( 
.A(n_752),
.Y(n_809)
);

AOI21xp5_ASAP7_75t_L g810 ( 
.A1(n_679),
.A2(n_592),
.B(n_585),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_677),
.Y(n_811)
);

NOR2xp33_ASAP7_75t_L g812 ( 
.A(n_670),
.B(n_595),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_L g813 ( 
.A(n_730),
.B(n_739),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_L g814 ( 
.A(n_739),
.B(n_528),
.Y(n_814)
);

CKINVDCx6p67_ASAP7_75t_R g815 ( 
.A(n_740),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_736),
.Y(n_816)
);

AND2x2_ASAP7_75t_L g817 ( 
.A(n_718),
.B(n_609),
.Y(n_817)
);

AND2x4_ASAP7_75t_L g818 ( 
.A(n_695),
.B(n_515),
.Y(n_818)
);

OAI21xp5_ASAP7_75t_L g819 ( 
.A1(n_753),
.A2(n_528),
.B(n_548),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_L g820 ( 
.A(n_688),
.B(n_548),
.Y(n_820)
);

INVx1_ASAP7_75t_L g821 ( 
.A(n_757),
.Y(n_821)
);

NOR2xp33_ASAP7_75t_L g822 ( 
.A(n_759),
.B(n_609),
.Y(n_822)
);

AOI21xp33_ASAP7_75t_L g823 ( 
.A1(n_750),
.A2(n_527),
.B(n_609),
.Y(n_823)
);

BUFx2_ASAP7_75t_L g824 ( 
.A(n_725),
.Y(n_824)
);

OAI21xp33_ASAP7_75t_L g825 ( 
.A1(n_689),
.A2(n_551),
.B(n_586),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_L g826 ( 
.A(n_703),
.B(n_587),
.Y(n_826)
);

NOR3xp33_ASAP7_75t_L g827 ( 
.A(n_764),
.B(n_766),
.C(n_704),
.Y(n_827)
);

HB1xp67_ASAP7_75t_L g828 ( 
.A(n_662),
.Y(n_828)
);

INVx2_ASAP7_75t_L g829 ( 
.A(n_742),
.Y(n_829)
);

INVx3_ASAP7_75t_L g830 ( 
.A(n_742),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_L g831 ( 
.A(n_713),
.B(n_515),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_762),
.Y(n_832)
);

AOI33xp33_ASAP7_75t_L g833 ( 
.A1(n_665),
.A2(n_770),
.A3(n_724),
.B1(n_760),
.B2(n_683),
.B3(n_685),
.Y(n_833)
);

AOI22xp5_ASAP7_75t_L g834 ( 
.A1(n_647),
.A2(n_565),
.B1(n_575),
.B2(n_611),
.Y(n_834)
);

INVx2_ASAP7_75t_L g835 ( 
.A(n_773),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_658),
.Y(n_836)
);

HB1xp67_ASAP7_75t_L g837 ( 
.A(n_662),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_659),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_L g839 ( 
.A(n_729),
.B(n_733),
.Y(n_839)
);

NOR2x1p5_ASAP7_75t_SL g840 ( 
.A(n_707),
.B(n_597),
.Y(n_840)
);

A2O1A1Ixp33_ASAP7_75t_L g841 ( 
.A1(n_764),
.A2(n_547),
.B(n_533),
.C(n_513),
.Y(n_841)
);

INVx2_ASAP7_75t_L g842 ( 
.A(n_649),
.Y(n_842)
);

AOI21xp5_ASAP7_75t_L g843 ( 
.A1(n_656),
.A2(n_607),
.B(n_632),
.Y(n_843)
);

O2A1O1Ixp33_ASAP7_75t_L g844 ( 
.A1(n_700),
.A2(n_25),
.B(n_26),
.C(n_27),
.Y(n_844)
);

AOI21xp5_ASAP7_75t_L g845 ( 
.A1(n_769),
.A2(n_607),
.B(n_632),
.Y(n_845)
);

AOI21xp5_ASAP7_75t_L g846 ( 
.A1(n_697),
.A2(n_607),
.B(n_632),
.Y(n_846)
);

HB1xp67_ASAP7_75t_L g847 ( 
.A(n_662),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_SL g848 ( 
.A(n_684),
.B(n_513),
.Y(n_848)
);

AND2x2_ASAP7_75t_L g849 ( 
.A(n_691),
.B(n_597),
.Y(n_849)
);

AOI21xp5_ASAP7_75t_L g850 ( 
.A1(n_667),
.A2(n_607),
.B(n_632),
.Y(n_850)
);

XNOR2xp5_ASAP7_75t_L g851 ( 
.A(n_756),
.B(n_76),
.Y(n_851)
);

AOI21xp5_ASAP7_75t_L g852 ( 
.A1(n_669),
.A2(n_632),
.B(n_547),
.Y(n_852)
);

NAND2x1p5_ASAP7_75t_L g853 ( 
.A(n_696),
.B(n_699),
.Y(n_853)
);

NOR3xp33_ASAP7_75t_L g854 ( 
.A(n_766),
.B(n_26),
.C(n_28),
.Y(n_854)
);

AOI21xp5_ASAP7_75t_L g855 ( 
.A1(n_671),
.A2(n_547),
.B(n_533),
.Y(n_855)
);

NOR2xp33_ASAP7_75t_SL g856 ( 
.A(n_754),
.B(n_611),
.Y(n_856)
);

AOI21xp5_ASAP7_75t_L g857 ( 
.A1(n_672),
.A2(n_675),
.B(n_673),
.Y(n_857)
);

OAI21xp33_ASAP7_75t_L g858 ( 
.A1(n_682),
.A2(n_28),
.B(n_29),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_738),
.Y(n_859)
);

INVx1_ASAP7_75t_L g860 ( 
.A(n_741),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_L g861 ( 
.A(n_709),
.B(n_712),
.Y(n_861)
);

BUFx6f_ASAP7_75t_L g862 ( 
.A(n_696),
.Y(n_862)
);

AOI21xp5_ASAP7_75t_L g863 ( 
.A1(n_715),
.A2(n_533),
.B(n_605),
.Y(n_863)
);

INVx2_ASAP7_75t_L g864 ( 
.A(n_680),
.Y(n_864)
);

NOR2xp33_ASAP7_75t_L g865 ( 
.A(n_652),
.B(n_533),
.Y(n_865)
);

INVx4_ASAP7_75t_L g866 ( 
.A(n_714),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_743),
.Y(n_867)
);

NOR2xp33_ASAP7_75t_L g868 ( 
.A(n_640),
.B(n_31),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_698),
.Y(n_869)
);

HB1xp67_ASAP7_75t_L g870 ( 
.A(n_687),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_L g871 ( 
.A(n_712),
.B(n_605),
.Y(n_871)
);

INVx3_ASAP7_75t_L g872 ( 
.A(n_726),
.Y(n_872)
);

BUFx6f_ASAP7_75t_L g873 ( 
.A(n_737),
.Y(n_873)
);

AND2x6_ASAP7_75t_L g874 ( 
.A(n_771),
.B(n_605),
.Y(n_874)
);

NOR3xp33_ASAP7_75t_L g875 ( 
.A(n_744),
.B(n_31),
.C(n_34),
.Y(n_875)
);

INVx2_ASAP7_75t_L g876 ( 
.A(n_661),
.Y(n_876)
);

INVx2_ASAP7_75t_L g877 ( 
.A(n_661),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_701),
.Y(n_878)
);

AOI21xp5_ASAP7_75t_L g879 ( 
.A1(n_719),
.A2(n_597),
.B(n_611),
.Y(n_879)
);

CKINVDCx8_ASAP7_75t_R g880 ( 
.A(n_681),
.Y(n_880)
);

INVx1_ASAP7_75t_L g881 ( 
.A(n_702),
.Y(n_881)
);

O2A1O1Ixp33_ASAP7_75t_L g882 ( 
.A1(n_690),
.A2(n_36),
.B(n_38),
.C(n_40),
.Y(n_882)
);

NOR2xp33_ASAP7_75t_L g883 ( 
.A(n_657),
.B(n_721),
.Y(n_883)
);

AOI21xp5_ASAP7_75t_L g884 ( 
.A1(n_705),
.A2(n_710),
.B(n_676),
.Y(n_884)
);

INVx3_ASAP7_75t_L g885 ( 
.A(n_758),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_L g886 ( 
.A(n_723),
.B(n_611),
.Y(n_886)
);

OAI21xp33_ASAP7_75t_L g887 ( 
.A1(n_692),
.A2(n_38),
.B(n_41),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_L g888 ( 
.A(n_723),
.B(n_44),
.Y(n_888)
);

AND2x2_ASAP7_75t_L g889 ( 
.A(n_714),
.B(n_45),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_SL g890 ( 
.A(n_767),
.B(n_91),
.Y(n_890)
);

OAI21xp5_ASAP7_75t_L g891 ( 
.A1(n_710),
.A2(n_660),
.B(n_749),
.Y(n_891)
);

BUFx4f_ASAP7_75t_L g892 ( 
.A(n_714),
.Y(n_892)
);

INVxp67_ASAP7_75t_L g893 ( 
.A(n_716),
.Y(n_893)
);

NOR2xp33_ASAP7_75t_L g894 ( 
.A(n_665),
.B(n_46),
.Y(n_894)
);

OR2x4_ASAP7_75t_L g895 ( 
.A(n_761),
.B(n_643),
.Y(n_895)
);

INVx1_ASAP7_75t_SL g896 ( 
.A(n_745),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_SL g897 ( 
.A(n_650),
.B(n_101),
.Y(n_897)
);

INVx1_ASAP7_75t_L g898 ( 
.A(n_728),
.Y(n_898)
);

OAI22xp5_ASAP7_75t_L g899 ( 
.A1(n_683),
.A2(n_82),
.B1(n_154),
.B2(n_153),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_SL g900 ( 
.A(n_642),
.B(n_70),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_L g901 ( 
.A(n_685),
.B(n_706),
.Y(n_901)
);

OAI22xp5_ASAP7_75t_L g902 ( 
.A1(n_706),
.A2(n_69),
.B1(n_140),
.B2(n_127),
.Y(n_902)
);

AOI21x1_ASAP7_75t_L g903 ( 
.A1(n_663),
.A2(n_64),
.B(n_126),
.Y(n_903)
);

A2O1A1Ixp33_ASAP7_75t_L g904 ( 
.A1(n_720),
.A2(n_49),
.B(n_51),
.C(n_55),
.Y(n_904)
);

BUFx6f_ASAP7_75t_L g905 ( 
.A(n_755),
.Y(n_905)
);

AOI21xp5_ASAP7_75t_L g906 ( 
.A1(n_720),
.A2(n_106),
.B(n_113),
.Y(n_906)
);

BUFx2_ASAP7_75t_L g907 ( 
.A(n_745),
.Y(n_907)
);

OAI21xp5_ASAP7_75t_L g908 ( 
.A1(n_653),
.A2(n_768),
.B(n_735),
.Y(n_908)
);

INVx1_ASAP7_75t_L g909 ( 
.A(n_655),
.Y(n_909)
);

NAND2x1p5_ASAP7_75t_L g910 ( 
.A(n_643),
.B(n_770),
.Y(n_910)
);

NAND2xp5_ASAP7_75t_SL g911 ( 
.A(n_643),
.B(n_62),
.Y(n_911)
);

HB1xp67_ASAP7_75t_L g912 ( 
.A(n_727),
.Y(n_912)
);

CKINVDCx5p33_ASAP7_75t_R g913 ( 
.A(n_809),
.Y(n_913)
);

NOR2x1_ASAP7_75t_L g914 ( 
.A(n_808),
.B(n_772),
.Y(n_914)
);

BUFx6f_ASAP7_75t_L g915 ( 
.A(n_802),
.Y(n_915)
);

NOR2xp33_ASAP7_75t_L g916 ( 
.A(n_813),
.B(n_727),
.Y(n_916)
);

OAI21x1_ASAP7_75t_L g917 ( 
.A1(n_800),
.A2(n_112),
.B(n_166),
.Y(n_917)
);

OAI21xp5_ASAP7_75t_L g918 ( 
.A1(n_778),
.A2(n_765),
.B(n_59),
.Y(n_918)
);

AOI21xp5_ASAP7_75t_L g919 ( 
.A1(n_774),
.A2(n_765),
.B(n_61),
.Y(n_919)
);

OAI21x1_ASAP7_75t_L g920 ( 
.A1(n_800),
.A2(n_58),
.B(n_747),
.Y(n_920)
);

A2O1A1Ixp33_ASAP7_75t_L g921 ( 
.A1(n_790),
.A2(n_861),
.B(n_827),
.C(n_891),
.Y(n_921)
);

BUFx2_ASAP7_75t_L g922 ( 
.A(n_777),
.Y(n_922)
);

AND2x4_ASAP7_75t_L g923 ( 
.A(n_885),
.B(n_866),
.Y(n_923)
);

INVx1_ASAP7_75t_L g924 ( 
.A(n_816),
.Y(n_924)
);

NOR2xp33_ASAP7_75t_SL g925 ( 
.A(n_910),
.B(n_787),
.Y(n_925)
);

INVx1_ASAP7_75t_SL g926 ( 
.A(n_870),
.Y(n_926)
);

OAI21xp5_ASAP7_75t_L g927 ( 
.A1(n_775),
.A2(n_884),
.B(n_909),
.Y(n_927)
);

OAI21xp5_ASAP7_75t_L g928 ( 
.A1(n_884),
.A2(n_796),
.B(n_857),
.Y(n_928)
);

NAND2xp5_ASAP7_75t_L g929 ( 
.A(n_780),
.B(n_859),
.Y(n_929)
);

INVx1_ASAP7_75t_L g930 ( 
.A(n_779),
.Y(n_930)
);

NAND2xp5_ASAP7_75t_L g931 ( 
.A(n_860),
.B(n_867),
.Y(n_931)
);

OAI22x1_ASAP7_75t_L g932 ( 
.A1(n_894),
.A2(n_868),
.B1(n_910),
.B2(n_791),
.Y(n_932)
);

OAI21xp5_ASAP7_75t_L g933 ( 
.A1(n_810),
.A2(n_799),
.B(n_825),
.Y(n_933)
);

NAND2xp5_ASAP7_75t_L g934 ( 
.A(n_869),
.B(n_878),
.Y(n_934)
);

NAND2xp5_ASAP7_75t_L g935 ( 
.A(n_881),
.B(n_839),
.Y(n_935)
);

INVx1_ASAP7_75t_SL g936 ( 
.A(n_794),
.Y(n_936)
);

NAND2xp5_ASAP7_75t_L g937 ( 
.A(n_785),
.B(n_788),
.Y(n_937)
);

BUFx2_ASAP7_75t_L g938 ( 
.A(n_824),
.Y(n_938)
);

AOI221x1_ASAP7_75t_L g939 ( 
.A1(n_888),
.A2(n_854),
.B1(n_906),
.B2(n_875),
.C(n_807),
.Y(n_939)
);

AOI21xp5_ASAP7_75t_L g940 ( 
.A1(n_820),
.A2(n_814),
.B(n_797),
.Y(n_940)
);

AOI221x1_ASAP7_75t_L g941 ( 
.A1(n_906),
.A2(n_781),
.B1(n_782),
.B2(n_887),
.C(n_908),
.Y(n_941)
);

AND2x2_ASAP7_75t_L g942 ( 
.A(n_817),
.B(n_885),
.Y(n_942)
);

OR2x6_ASAP7_75t_L g943 ( 
.A(n_808),
.B(n_866),
.Y(n_943)
);

AOI21x1_ASAP7_75t_SL g944 ( 
.A1(n_871),
.A2(n_886),
.B(n_831),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_L g945 ( 
.A(n_883),
.B(n_798),
.Y(n_945)
);

AND3x4_ASAP7_75t_L g946 ( 
.A(n_880),
.B(n_876),
.C(n_877),
.Y(n_946)
);

OAI21xp5_ASAP7_75t_L g947 ( 
.A1(n_801),
.A2(n_901),
.B(n_819),
.Y(n_947)
);

AOI22xp5_ASAP7_75t_L g948 ( 
.A1(n_789),
.A2(n_795),
.B1(n_822),
.B2(n_893),
.Y(n_948)
);

NOR2xp33_ASAP7_75t_L g949 ( 
.A(n_793),
.B(n_823),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_L g950 ( 
.A(n_811),
.B(n_833),
.Y(n_950)
);

AO21x1_ASAP7_75t_L g951 ( 
.A1(n_900),
.A2(n_890),
.B(n_844),
.Y(n_951)
);

BUFx6f_ASAP7_75t_L g952 ( 
.A(n_802),
.Y(n_952)
);

CKINVDCx5p33_ASAP7_75t_R g953 ( 
.A(n_804),
.Y(n_953)
);

BUFx2_ASAP7_75t_L g954 ( 
.A(n_907),
.Y(n_954)
);

AOI21xp5_ASAP7_75t_L g955 ( 
.A1(n_830),
.A2(n_849),
.B(n_848),
.Y(n_955)
);

NOR3xp33_ASAP7_75t_L g956 ( 
.A(n_812),
.B(n_786),
.C(n_911),
.Y(n_956)
);

AOI21xp33_ASAP7_75t_L g957 ( 
.A1(n_898),
.A2(n_858),
.B(n_882),
.Y(n_957)
);

NAND2xp5_ASAP7_75t_SL g958 ( 
.A(n_802),
.B(n_787),
.Y(n_958)
);

BUFx2_ASAP7_75t_SL g959 ( 
.A(n_905),
.Y(n_959)
);

NAND2xp5_ASAP7_75t_L g960 ( 
.A(n_829),
.B(n_865),
.Y(n_960)
);

OAI22xp5_ASAP7_75t_L g961 ( 
.A1(n_904),
.A2(n_899),
.B1(n_902),
.B2(n_838),
.Y(n_961)
);

AND2x2_ASAP7_75t_L g962 ( 
.A(n_828),
.B(n_847),
.Y(n_962)
);

AND2x2_ASAP7_75t_L g963 ( 
.A(n_837),
.B(n_889),
.Y(n_963)
);

XOR2xp5_ASAP7_75t_L g964 ( 
.A(n_783),
.B(n_851),
.Y(n_964)
);

OR2x2_ASAP7_75t_L g965 ( 
.A(n_896),
.B(n_836),
.Y(n_965)
);

NAND2xp5_ASAP7_75t_L g966 ( 
.A(n_821),
.B(n_832),
.Y(n_966)
);

NAND2xp5_ASAP7_75t_L g967 ( 
.A(n_826),
.B(n_835),
.Y(n_967)
);

AND2x2_ASAP7_75t_L g968 ( 
.A(n_905),
.B(n_808),
.Y(n_968)
);

NOR2xp33_ASAP7_75t_L g969 ( 
.A(n_905),
.B(n_776),
.Y(n_969)
);

OAI21x1_ASAP7_75t_L g970 ( 
.A1(n_863),
.A2(n_845),
.B(n_879),
.Y(n_970)
);

INVx2_ASAP7_75t_SL g971 ( 
.A(n_892),
.Y(n_971)
);

OR2x6_ASAP7_75t_L g972 ( 
.A(n_912),
.B(n_792),
.Y(n_972)
);

OAI21x1_ASAP7_75t_L g973 ( 
.A1(n_863),
.A2(n_843),
.B(n_846),
.Y(n_973)
);

INVxp67_ASAP7_75t_L g974 ( 
.A(n_892),
.Y(n_974)
);

AOI22xp5_ASAP7_75t_L g975 ( 
.A1(n_818),
.A2(n_895),
.B1(n_862),
.B2(n_897),
.Y(n_975)
);

INVx3_ASAP7_75t_SL g976 ( 
.A(n_815),
.Y(n_976)
);

OR2x6_ASAP7_75t_L g977 ( 
.A(n_792),
.B(n_853),
.Y(n_977)
);

INVx1_ASAP7_75t_L g978 ( 
.A(n_842),
.Y(n_978)
);

NAND2xp5_ASAP7_75t_SL g979 ( 
.A(n_862),
.B(n_856),
.Y(n_979)
);

OAI21xp5_ASAP7_75t_L g980 ( 
.A1(n_855),
.A2(n_852),
.B(n_850),
.Y(n_980)
);

NAND2x1p5_ASAP7_75t_L g981 ( 
.A(n_862),
.B(n_873),
.Y(n_981)
);

INVx2_ASAP7_75t_SL g982 ( 
.A(n_895),
.Y(n_982)
);

BUFx3_ASAP7_75t_L g983 ( 
.A(n_873),
.Y(n_983)
);

OAI21x1_ASAP7_75t_L g984 ( 
.A1(n_872),
.A2(n_903),
.B(n_806),
.Y(n_984)
);

INVxp67_ASAP7_75t_L g985 ( 
.A(n_864),
.Y(n_985)
);

AOI21xp5_ASAP7_75t_L g986 ( 
.A1(n_872),
.A2(n_873),
.B(n_834),
.Y(n_986)
);

OAI21x1_ASAP7_75t_L g987 ( 
.A1(n_840),
.A2(n_874),
.B(n_784),
.Y(n_987)
);

NAND2xp5_ASAP7_75t_L g988 ( 
.A(n_874),
.B(n_813),
.Y(n_988)
);

AO21x1_ASAP7_75t_L g989 ( 
.A1(n_874),
.A2(n_790),
.B(n_813),
.Y(n_989)
);

A2O1A1Ixp33_ASAP7_75t_L g990 ( 
.A1(n_874),
.A2(n_790),
.B(n_813),
.C(n_532),
.Y(n_990)
);

INVx1_ASAP7_75t_L g991 ( 
.A(n_874),
.Y(n_991)
);

A2O1A1Ixp33_ASAP7_75t_L g992 ( 
.A1(n_790),
.A2(n_813),
.B(n_532),
.C(n_861),
.Y(n_992)
);

NAND2xp5_ASAP7_75t_L g993 ( 
.A(n_813),
.B(n_790),
.Y(n_993)
);

NAND2xp5_ASAP7_75t_L g994 ( 
.A(n_813),
.B(n_790),
.Y(n_994)
);

INVx3_ASAP7_75t_L g995 ( 
.A(n_818),
.Y(n_995)
);

A2O1A1Ixp33_ASAP7_75t_L g996 ( 
.A1(n_790),
.A2(n_813),
.B(n_532),
.C(n_861),
.Y(n_996)
);

HB1xp67_ASAP7_75t_L g997 ( 
.A(n_777),
.Y(n_997)
);

NAND2xp5_ASAP7_75t_L g998 ( 
.A(n_790),
.B(n_813),
.Y(n_998)
);

NAND2xp5_ASAP7_75t_L g999 ( 
.A(n_790),
.B(n_813),
.Y(n_999)
);

A2O1A1Ixp33_ASAP7_75t_L g1000 ( 
.A1(n_790),
.A2(n_813),
.B(n_532),
.C(n_861),
.Y(n_1000)
);

A2O1A1Ixp33_ASAP7_75t_L g1001 ( 
.A1(n_790),
.A2(n_813),
.B(n_532),
.C(n_861),
.Y(n_1001)
);

BUFx10_ASAP7_75t_L g1002 ( 
.A(n_793),
.Y(n_1002)
);

A2O1A1Ixp33_ASAP7_75t_L g1003 ( 
.A1(n_790),
.A2(n_813),
.B(n_532),
.C(n_861),
.Y(n_1003)
);

OAI21xp33_ASAP7_75t_SL g1004 ( 
.A1(n_901),
.A2(n_790),
.B(n_833),
.Y(n_1004)
);

AND2x2_ASAP7_75t_L g1005 ( 
.A(n_817),
.B(n_668),
.Y(n_1005)
);

A2O1A1Ixp33_ASAP7_75t_L g1006 ( 
.A1(n_790),
.A2(n_813),
.B(n_532),
.C(n_861),
.Y(n_1006)
);

NAND3xp33_ASAP7_75t_L g1007 ( 
.A(n_813),
.B(n_790),
.C(n_523),
.Y(n_1007)
);

OAI21xp5_ASAP7_75t_L g1008 ( 
.A1(n_778),
.A2(n_532),
.B(n_790),
.Y(n_1008)
);

HB1xp67_ASAP7_75t_L g1009 ( 
.A(n_777),
.Y(n_1009)
);

NOR2xp33_ASAP7_75t_L g1010 ( 
.A(n_813),
.B(n_790),
.Y(n_1010)
);

NAND2xp5_ASAP7_75t_L g1011 ( 
.A(n_790),
.B(n_813),
.Y(n_1011)
);

OAI21x1_ASAP7_75t_L g1012 ( 
.A1(n_800),
.A2(n_803),
.B(n_805),
.Y(n_1012)
);

OAI21xp5_ASAP7_75t_L g1013 ( 
.A1(n_778),
.A2(n_532),
.B(n_790),
.Y(n_1013)
);

BUFx2_ASAP7_75t_L g1014 ( 
.A(n_777),
.Y(n_1014)
);

AO31x2_ASAP7_75t_L g1015 ( 
.A1(n_796),
.A2(n_841),
.A3(n_909),
.B(n_884),
.Y(n_1015)
);

NAND2x1p5_ASAP7_75t_L g1016 ( 
.A(n_792),
.B(n_802),
.Y(n_1016)
);

OAI21x1_ASAP7_75t_L g1017 ( 
.A1(n_800),
.A2(n_803),
.B(n_805),
.Y(n_1017)
);

NAND2xp5_ASAP7_75t_L g1018 ( 
.A(n_813),
.B(n_790),
.Y(n_1018)
);

NAND2xp5_ASAP7_75t_L g1019 ( 
.A(n_790),
.B(n_813),
.Y(n_1019)
);

INVx3_ASAP7_75t_L g1020 ( 
.A(n_818),
.Y(n_1020)
);

OAI21xp5_ASAP7_75t_L g1021 ( 
.A1(n_778),
.A2(n_532),
.B(n_790),
.Y(n_1021)
);

NAND2x1_ASAP7_75t_L g1022 ( 
.A(n_792),
.B(n_751),
.Y(n_1022)
);

BUFx2_ASAP7_75t_L g1023 ( 
.A(n_777),
.Y(n_1023)
);

OAI21x1_ASAP7_75t_L g1024 ( 
.A1(n_800),
.A2(n_803),
.B(n_805),
.Y(n_1024)
);

OAI21xp33_ASAP7_75t_L g1025 ( 
.A1(n_813),
.A2(n_523),
.B(n_514),
.Y(n_1025)
);

OR2x2_ASAP7_75t_L g1026 ( 
.A(n_870),
.B(n_530),
.Y(n_1026)
);

INVx1_ASAP7_75t_L g1027 ( 
.A(n_816),
.Y(n_1027)
);

OAI21xp5_ASAP7_75t_L g1028 ( 
.A1(n_778),
.A2(n_532),
.B(n_790),
.Y(n_1028)
);

AOI21xp33_ASAP7_75t_L g1029 ( 
.A1(n_790),
.A2(n_813),
.B(n_861),
.Y(n_1029)
);

AO31x2_ASAP7_75t_L g1030 ( 
.A1(n_796),
.A2(n_841),
.A3(n_909),
.B(n_884),
.Y(n_1030)
);

BUFx3_ASAP7_75t_L g1031 ( 
.A(n_777),
.Y(n_1031)
);

AOI21xp33_ASAP7_75t_L g1032 ( 
.A1(n_790),
.A2(n_813),
.B(n_861),
.Y(n_1032)
);

AND2x4_ASAP7_75t_L g1033 ( 
.A(n_982),
.B(n_923),
.Y(n_1033)
);

INVx1_ASAP7_75t_L g1034 ( 
.A(n_924),
.Y(n_1034)
);

NAND2xp5_ASAP7_75t_L g1035 ( 
.A(n_1010),
.B(n_998),
.Y(n_1035)
);

AND2x2_ASAP7_75t_L g1036 ( 
.A(n_1005),
.B(n_963),
.Y(n_1036)
);

INVx4_ASAP7_75t_L g1037 ( 
.A(n_915),
.Y(n_1037)
);

INVx2_ASAP7_75t_L g1038 ( 
.A(n_930),
.Y(n_1038)
);

O2A1O1Ixp33_ASAP7_75t_L g1039 ( 
.A1(n_1025),
.A2(n_921),
.B(n_999),
.C(n_998),
.Y(n_1039)
);

AND2x4_ASAP7_75t_L g1040 ( 
.A(n_923),
.B(n_968),
.Y(n_1040)
);

INVx2_ASAP7_75t_L g1041 ( 
.A(n_1027),
.Y(n_1041)
);

AND2x4_ASAP7_75t_L g1042 ( 
.A(n_971),
.B(n_943),
.Y(n_1042)
);

NAND2xp5_ASAP7_75t_SL g1043 ( 
.A(n_948),
.B(n_949),
.Y(n_1043)
);

INVxp67_ASAP7_75t_L g1044 ( 
.A(n_1026),
.Y(n_1044)
);

INVx1_ASAP7_75t_SL g1045 ( 
.A(n_936),
.Y(n_1045)
);

INVx4_ASAP7_75t_L g1046 ( 
.A(n_915),
.Y(n_1046)
);

AOI22xp5_ASAP7_75t_L g1047 ( 
.A1(n_932),
.A2(n_916),
.B1(n_1007),
.B2(n_956),
.Y(n_1047)
);

INVx1_ASAP7_75t_L g1048 ( 
.A(n_966),
.Y(n_1048)
);

AOI22xp33_ASAP7_75t_L g1049 ( 
.A1(n_1029),
.A2(n_1032),
.B1(n_951),
.B2(n_918),
.Y(n_1049)
);

OAI21xp5_ASAP7_75t_L g1050 ( 
.A1(n_992),
.A2(n_1000),
.B(n_996),
.Y(n_1050)
);

AOI22xp33_ASAP7_75t_L g1051 ( 
.A1(n_1029),
.A2(n_1032),
.B1(n_918),
.B2(n_994),
.Y(n_1051)
);

OAI22xp5_ASAP7_75t_SL g1052 ( 
.A1(n_946),
.A2(n_964),
.B1(n_974),
.B2(n_913),
.Y(n_1052)
);

OAI22xp5_ASAP7_75t_L g1053 ( 
.A1(n_999),
.A2(n_1019),
.B1(n_1011),
.B2(n_993),
.Y(n_1053)
);

NAND2xp5_ASAP7_75t_L g1054 ( 
.A(n_1011),
.B(n_1019),
.Y(n_1054)
);

NAND2xp5_ASAP7_75t_L g1055 ( 
.A(n_1018),
.B(n_929),
.Y(n_1055)
);

BUFx3_ASAP7_75t_L g1056 ( 
.A(n_1031),
.Y(n_1056)
);

NAND2xp5_ASAP7_75t_L g1057 ( 
.A(n_929),
.B(n_945),
.Y(n_1057)
);

AND2x4_ASAP7_75t_L g1058 ( 
.A(n_943),
.B(n_942),
.Y(n_1058)
);

BUFx3_ASAP7_75t_L g1059 ( 
.A(n_922),
.Y(n_1059)
);

OAI22xp5_ASAP7_75t_L g1060 ( 
.A1(n_931),
.A2(n_935),
.B1(n_934),
.B2(n_950),
.Y(n_1060)
);

NAND2xp5_ASAP7_75t_L g1061 ( 
.A(n_931),
.B(n_934),
.Y(n_1061)
);

BUFx12f_ASAP7_75t_L g1062 ( 
.A(n_953),
.Y(n_1062)
);

OR2x2_ASAP7_75t_L g1063 ( 
.A(n_926),
.B(n_1014),
.Y(n_1063)
);

OAI22xp5_ASAP7_75t_L g1064 ( 
.A1(n_1001),
.A2(n_1003),
.B1(n_1006),
.B2(n_937),
.Y(n_1064)
);

OAI22xp5_ASAP7_75t_L g1065 ( 
.A1(n_961),
.A2(n_947),
.B1(n_990),
.B2(n_1021),
.Y(n_1065)
);

NOR2xp33_ASAP7_75t_L g1066 ( 
.A(n_926),
.B(n_936),
.Y(n_1066)
);

OAI221xp5_ASAP7_75t_L g1067 ( 
.A1(n_1004),
.A2(n_957),
.B1(n_961),
.B2(n_919),
.C(n_914),
.Y(n_1067)
);

OR2x6_ASAP7_75t_L g1068 ( 
.A(n_959),
.B(n_943),
.Y(n_1068)
);

OAI22xp5_ASAP7_75t_L g1069 ( 
.A1(n_947),
.A2(n_1028),
.B1(n_1021),
.B2(n_1013),
.Y(n_1069)
);

A2O1A1Ixp33_ASAP7_75t_L g1070 ( 
.A1(n_957),
.A2(n_1008),
.B(n_1028),
.C(n_1013),
.Y(n_1070)
);

AND2x4_ASAP7_75t_L g1071 ( 
.A(n_995),
.B(n_1020),
.Y(n_1071)
);

NOR2xp33_ASAP7_75t_L g1072 ( 
.A(n_997),
.B(n_1009),
.Y(n_1072)
);

OAI22xp5_ASAP7_75t_L g1073 ( 
.A1(n_1008),
.A2(n_988),
.B1(n_967),
.B2(n_933),
.Y(n_1073)
);

INVx2_ASAP7_75t_L g1074 ( 
.A(n_978),
.Y(n_1074)
);

INVx1_ASAP7_75t_L g1075 ( 
.A(n_985),
.Y(n_1075)
);

INVx1_ASAP7_75t_L g1076 ( 
.A(n_965),
.Y(n_1076)
);

NOR2xp33_ASAP7_75t_L g1077 ( 
.A(n_1023),
.B(n_938),
.Y(n_1077)
);

HB1xp67_ASAP7_75t_L g1078 ( 
.A(n_954),
.Y(n_1078)
);

INVx3_ASAP7_75t_SL g1079 ( 
.A(n_976),
.Y(n_1079)
);

AND2x2_ASAP7_75t_L g1080 ( 
.A(n_962),
.B(n_1002),
.Y(n_1080)
);

OAI22xp5_ASAP7_75t_L g1081 ( 
.A1(n_933),
.A2(n_927),
.B1(n_975),
.B2(n_928),
.Y(n_1081)
);

OAI22xp33_ASAP7_75t_SL g1082 ( 
.A1(n_925),
.A2(n_960),
.B1(n_972),
.B2(n_958),
.Y(n_1082)
);

INVx1_ASAP7_75t_L g1083 ( 
.A(n_969),
.Y(n_1083)
);

INVx1_ASAP7_75t_SL g1084 ( 
.A(n_1002),
.Y(n_1084)
);

AND2x4_ASAP7_75t_L g1085 ( 
.A(n_995),
.B(n_1020),
.Y(n_1085)
);

OAI22xp5_ASAP7_75t_L g1086 ( 
.A1(n_927),
.A2(n_928),
.B1(n_960),
.B2(n_979),
.Y(n_1086)
);

NOR2xp67_ASAP7_75t_L g1087 ( 
.A(n_983),
.B(n_955),
.Y(n_1087)
);

OR2x6_ASAP7_75t_L g1088 ( 
.A(n_972),
.B(n_977),
.Y(n_1088)
);

NAND2xp5_ASAP7_75t_L g1089 ( 
.A(n_939),
.B(n_941),
.Y(n_1089)
);

INVxp67_ASAP7_75t_L g1090 ( 
.A(n_972),
.Y(n_1090)
);

AND2x4_ASAP7_75t_L g1091 ( 
.A(n_987),
.B(n_977),
.Y(n_1091)
);

INVx2_ASAP7_75t_L g1092 ( 
.A(n_981),
.Y(n_1092)
);

BUFx3_ASAP7_75t_L g1093 ( 
.A(n_915),
.Y(n_1093)
);

INVx2_ASAP7_75t_L g1094 ( 
.A(n_1016),
.Y(n_1094)
);

INVx1_ASAP7_75t_L g1095 ( 
.A(n_952),
.Y(n_1095)
);

INVx2_ASAP7_75t_L g1096 ( 
.A(n_1016),
.Y(n_1096)
);

NAND2xp5_ASAP7_75t_L g1097 ( 
.A(n_925),
.B(n_986),
.Y(n_1097)
);

NAND2x1_ASAP7_75t_L g1098 ( 
.A(n_977),
.B(n_952),
.Y(n_1098)
);

AOI22xp33_ASAP7_75t_L g1099 ( 
.A1(n_989),
.A2(n_991),
.B1(n_920),
.B2(n_980),
.Y(n_1099)
);

AND2x2_ASAP7_75t_L g1100 ( 
.A(n_1015),
.B(n_1030),
.Y(n_1100)
);

AND2x2_ASAP7_75t_L g1101 ( 
.A(n_1015),
.B(n_1030),
.Y(n_1101)
);

BUFx3_ASAP7_75t_L g1102 ( 
.A(n_1022),
.Y(n_1102)
);

HB1xp67_ASAP7_75t_L g1103 ( 
.A(n_917),
.Y(n_1103)
);

NOR2xp33_ASAP7_75t_L g1104 ( 
.A(n_970),
.B(n_973),
.Y(n_1104)
);

AND2x2_ASAP7_75t_SL g1105 ( 
.A(n_944),
.B(n_984),
.Y(n_1105)
);

CKINVDCx5p33_ASAP7_75t_R g1106 ( 
.A(n_1012),
.Y(n_1106)
);

INVx5_ASAP7_75t_L g1107 ( 
.A(n_1017),
.Y(n_1107)
);

BUFx3_ASAP7_75t_L g1108 ( 
.A(n_1024),
.Y(n_1108)
);

INVx4_ASAP7_75t_L g1109 ( 
.A(n_915),
.Y(n_1109)
);

OA21x2_ASAP7_75t_L g1110 ( 
.A1(n_927),
.A2(n_928),
.B(n_933),
.Y(n_1110)
);

INVx1_ASAP7_75t_SL g1111 ( 
.A(n_936),
.Y(n_1111)
);

AND2x4_ASAP7_75t_L g1112 ( 
.A(n_982),
.B(n_923),
.Y(n_1112)
);

AOI22xp33_ASAP7_75t_L g1113 ( 
.A1(n_1025),
.A2(n_790),
.B1(n_813),
.B2(n_868),
.Y(n_1113)
);

INVx5_ASAP7_75t_L g1114 ( 
.A(n_915),
.Y(n_1114)
);

NAND2xp33_ASAP7_75t_L g1115 ( 
.A(n_1025),
.B(n_827),
.Y(n_1115)
);

NOR2xp33_ASAP7_75t_L g1116 ( 
.A(n_1010),
.B(n_813),
.Y(n_1116)
);

INVx3_ASAP7_75t_L g1117 ( 
.A(n_981),
.Y(n_1117)
);

INVx3_ASAP7_75t_L g1118 ( 
.A(n_981),
.Y(n_1118)
);

NAND2xp5_ASAP7_75t_L g1119 ( 
.A(n_1010),
.B(n_998),
.Y(n_1119)
);

AND2x2_ASAP7_75t_L g1120 ( 
.A(n_1005),
.B(n_817),
.Y(n_1120)
);

NAND2xp5_ASAP7_75t_L g1121 ( 
.A(n_1010),
.B(n_998),
.Y(n_1121)
);

BUFx8_ASAP7_75t_SL g1122 ( 
.A(n_913),
.Y(n_1122)
);

NAND3xp33_ASAP7_75t_L g1123 ( 
.A(n_1010),
.B(n_813),
.C(n_790),
.Y(n_1123)
);

A2O1A1Ixp33_ASAP7_75t_L g1124 ( 
.A1(n_1010),
.A2(n_813),
.B(n_790),
.C(n_1025),
.Y(n_1124)
);

NAND2x1p5_ASAP7_75t_L g1125 ( 
.A(n_958),
.B(n_792),
.Y(n_1125)
);

AND2x4_ASAP7_75t_L g1126 ( 
.A(n_982),
.B(n_923),
.Y(n_1126)
);

AND2x4_ASAP7_75t_L g1127 ( 
.A(n_982),
.B(n_923),
.Y(n_1127)
);

OAI22xp5_ASAP7_75t_L g1128 ( 
.A1(n_1010),
.A2(n_532),
.B1(n_999),
.B2(n_998),
.Y(n_1128)
);

O2A1O1Ixp5_ASAP7_75t_SL g1129 ( 
.A1(n_918),
.A2(n_1032),
.B(n_1029),
.C(n_980),
.Y(n_1129)
);

OAI22xp5_ASAP7_75t_L g1130 ( 
.A1(n_1010),
.A2(n_532),
.B1(n_999),
.B2(n_998),
.Y(n_1130)
);

AOI21xp33_ASAP7_75t_SL g1131 ( 
.A1(n_946),
.A2(n_523),
.B(n_514),
.Y(n_1131)
);

HB1xp67_ASAP7_75t_L g1132 ( 
.A(n_997),
.Y(n_1132)
);

NAND2xp5_ASAP7_75t_L g1133 ( 
.A(n_1010),
.B(n_998),
.Y(n_1133)
);

AOI21xp33_ASAP7_75t_SL g1134 ( 
.A1(n_946),
.A2(n_523),
.B(n_514),
.Y(n_1134)
);

NAND2xp5_ASAP7_75t_SL g1135 ( 
.A(n_948),
.B(n_791),
.Y(n_1135)
);

INVx1_ASAP7_75t_SL g1136 ( 
.A(n_936),
.Y(n_1136)
);

AND2x2_ASAP7_75t_L g1137 ( 
.A(n_1005),
.B(n_817),
.Y(n_1137)
);

CKINVDCx5p33_ASAP7_75t_R g1138 ( 
.A(n_913),
.Y(n_1138)
);

NAND2xp5_ASAP7_75t_SL g1139 ( 
.A(n_948),
.B(n_791),
.Y(n_1139)
);

AOI21xp5_ASAP7_75t_L g1140 ( 
.A1(n_940),
.A2(n_532),
.B(n_790),
.Y(n_1140)
);

INVx1_ASAP7_75t_L g1141 ( 
.A(n_924),
.Y(n_1141)
);

AND2x2_ASAP7_75t_L g1142 ( 
.A(n_1005),
.B(n_817),
.Y(n_1142)
);

HB1xp67_ASAP7_75t_L g1143 ( 
.A(n_997),
.Y(n_1143)
);

HB1xp67_ASAP7_75t_L g1144 ( 
.A(n_997),
.Y(n_1144)
);

AOI21xp5_ASAP7_75t_L g1145 ( 
.A1(n_940),
.A2(n_532),
.B(n_790),
.Y(n_1145)
);

AOI21xp5_ASAP7_75t_L g1146 ( 
.A1(n_940),
.A2(n_532),
.B(n_790),
.Y(n_1146)
);

AOI21xp5_ASAP7_75t_L g1147 ( 
.A1(n_940),
.A2(n_532),
.B(n_790),
.Y(n_1147)
);

OAI21xp5_ASAP7_75t_L g1148 ( 
.A1(n_921),
.A2(n_790),
.B(n_992),
.Y(n_1148)
);

A2O1A1Ixp33_ASAP7_75t_L g1149 ( 
.A1(n_1010),
.A2(n_813),
.B(n_790),
.C(n_1025),
.Y(n_1149)
);

INVx2_ASAP7_75t_L g1150 ( 
.A(n_924),
.Y(n_1150)
);

NOR2xp33_ASAP7_75t_L g1151 ( 
.A(n_1010),
.B(n_813),
.Y(n_1151)
);

INVx1_ASAP7_75t_L g1152 ( 
.A(n_924),
.Y(n_1152)
);

BUFx3_ASAP7_75t_L g1153 ( 
.A(n_1031),
.Y(n_1153)
);

NAND2xp5_ASAP7_75t_L g1154 ( 
.A(n_1010),
.B(n_998),
.Y(n_1154)
);

NAND2xp5_ASAP7_75t_L g1155 ( 
.A(n_1010),
.B(n_998),
.Y(n_1155)
);

OAI22xp5_ASAP7_75t_L g1156 ( 
.A1(n_1010),
.A2(n_532),
.B1(n_999),
.B2(n_998),
.Y(n_1156)
);

INVx1_ASAP7_75t_SL g1157 ( 
.A(n_936),
.Y(n_1157)
);

BUFx8_ASAP7_75t_L g1158 ( 
.A(n_922),
.Y(n_1158)
);

NAND2xp5_ASAP7_75t_L g1159 ( 
.A(n_1010),
.B(n_998),
.Y(n_1159)
);

OAI22xp5_ASAP7_75t_L g1160 ( 
.A1(n_1010),
.A2(n_532),
.B1(n_999),
.B2(n_998),
.Y(n_1160)
);

OAI21xp5_ASAP7_75t_L g1161 ( 
.A1(n_921),
.A2(n_790),
.B(n_992),
.Y(n_1161)
);

INVxp67_ASAP7_75t_L g1162 ( 
.A(n_1066),
.Y(n_1162)
);

AO21x1_ASAP7_75t_L g1163 ( 
.A1(n_1065),
.A2(n_1069),
.B(n_1148),
.Y(n_1163)
);

BUFx6f_ASAP7_75t_L g1164 ( 
.A(n_1114),
.Y(n_1164)
);

BUFx2_ASAP7_75t_L g1165 ( 
.A(n_1063),
.Y(n_1165)
);

INVxp67_ASAP7_75t_L g1166 ( 
.A(n_1072),
.Y(n_1166)
);

AOI22xp33_ASAP7_75t_L g1167 ( 
.A1(n_1043),
.A2(n_1139),
.B1(n_1135),
.B2(n_1151),
.Y(n_1167)
);

AOI22xp33_ASAP7_75t_SL g1168 ( 
.A1(n_1116),
.A2(n_1115),
.B1(n_1123),
.B2(n_1067),
.Y(n_1168)
);

AOI22xp33_ASAP7_75t_SL g1169 ( 
.A1(n_1065),
.A2(n_1069),
.B1(n_1035),
.B2(n_1119),
.Y(n_1169)
);

AOI22xp33_ASAP7_75t_SL g1170 ( 
.A1(n_1119),
.A2(n_1159),
.B1(n_1154),
.B2(n_1155),
.Y(n_1170)
);

INVx1_ASAP7_75t_L g1171 ( 
.A(n_1100),
.Y(n_1171)
);

INVx1_ASAP7_75t_L g1172 ( 
.A(n_1041),
.Y(n_1172)
);

HB1xp67_ASAP7_75t_L g1173 ( 
.A(n_1045),
.Y(n_1173)
);

INVx1_ASAP7_75t_L g1174 ( 
.A(n_1150),
.Y(n_1174)
);

INVx3_ASAP7_75t_L g1175 ( 
.A(n_1091),
.Y(n_1175)
);

INVx1_ASAP7_75t_L g1176 ( 
.A(n_1034),
.Y(n_1176)
);

INVx3_ASAP7_75t_L g1177 ( 
.A(n_1091),
.Y(n_1177)
);

INVx6_ASAP7_75t_L g1178 ( 
.A(n_1114),
.Y(n_1178)
);

AOI22xp33_ASAP7_75t_L g1179 ( 
.A1(n_1113),
.A2(n_1120),
.B1(n_1137),
.B2(n_1142),
.Y(n_1179)
);

CKINVDCx5p33_ASAP7_75t_R g1180 ( 
.A(n_1122),
.Y(n_1180)
);

OAI22xp5_ASAP7_75t_L g1181 ( 
.A1(n_1121),
.A2(n_1155),
.B1(n_1154),
.B2(n_1133),
.Y(n_1181)
);

BUFx2_ASAP7_75t_L g1182 ( 
.A(n_1097),
.Y(n_1182)
);

AND2x2_ASAP7_75t_L g1183 ( 
.A(n_1054),
.B(n_1053),
.Y(n_1183)
);

BUFx2_ASAP7_75t_L g1184 ( 
.A(n_1097),
.Y(n_1184)
);

INVx2_ASAP7_75t_SL g1185 ( 
.A(n_1114),
.Y(n_1185)
);

AND2x2_ASAP7_75t_L g1186 ( 
.A(n_1054),
.B(n_1053),
.Y(n_1186)
);

BUFx3_ASAP7_75t_L g1187 ( 
.A(n_1056),
.Y(n_1187)
);

INVx2_ASAP7_75t_SL g1188 ( 
.A(n_1114),
.Y(n_1188)
);

AND2x4_ASAP7_75t_L g1189 ( 
.A(n_1058),
.B(n_1040),
.Y(n_1189)
);

AOI22xp5_ASAP7_75t_SL g1190 ( 
.A1(n_1058),
.A2(n_1133),
.B1(n_1159),
.B2(n_1121),
.Y(n_1190)
);

BUFx12f_ASAP7_75t_L g1191 ( 
.A(n_1138),
.Y(n_1191)
);

HB1xp67_ASAP7_75t_L g1192 ( 
.A(n_1111),
.Y(n_1192)
);

INVx1_ASAP7_75t_L g1193 ( 
.A(n_1141),
.Y(n_1193)
);

AND2x4_ASAP7_75t_L g1194 ( 
.A(n_1040),
.B(n_1042),
.Y(n_1194)
);

AOI22xp33_ASAP7_75t_L g1195 ( 
.A1(n_1047),
.A2(n_1051),
.B1(n_1049),
.B2(n_1060),
.Y(n_1195)
);

INVx1_ASAP7_75t_L g1196 ( 
.A(n_1152),
.Y(n_1196)
);

CKINVDCx6p67_ASAP7_75t_R g1197 ( 
.A(n_1079),
.Y(n_1197)
);

INVx1_ASAP7_75t_L g1198 ( 
.A(n_1101),
.Y(n_1198)
);

OAI22xp5_ASAP7_75t_L g1199 ( 
.A1(n_1055),
.A2(n_1061),
.B1(n_1057),
.B2(n_1131),
.Y(n_1199)
);

BUFx8_ASAP7_75t_SL g1200 ( 
.A(n_1062),
.Y(n_1200)
);

OR2x2_ASAP7_75t_L g1201 ( 
.A(n_1110),
.B(n_1081),
.Y(n_1201)
);

BUFx3_ASAP7_75t_L g1202 ( 
.A(n_1153),
.Y(n_1202)
);

INVx1_ASAP7_75t_L g1203 ( 
.A(n_1074),
.Y(n_1203)
);

OAI22xp5_ASAP7_75t_L g1204 ( 
.A1(n_1055),
.A2(n_1061),
.B1(n_1057),
.B2(n_1134),
.Y(n_1204)
);

OAI22xp5_ASAP7_75t_L g1205 ( 
.A1(n_1048),
.A2(n_1149),
.B1(n_1124),
.B2(n_1083),
.Y(n_1205)
);

AND2x2_ASAP7_75t_L g1206 ( 
.A(n_1060),
.B(n_1128),
.Y(n_1206)
);

BUFx3_ASAP7_75t_L g1207 ( 
.A(n_1158),
.Y(n_1207)
);

INVx3_ASAP7_75t_L g1208 ( 
.A(n_1108),
.Y(n_1208)
);

BUFx12f_ASAP7_75t_L g1209 ( 
.A(n_1158),
.Y(n_1209)
);

HB1xp67_ASAP7_75t_L g1210 ( 
.A(n_1136),
.Y(n_1210)
);

INVx1_ASAP7_75t_L g1211 ( 
.A(n_1076),
.Y(n_1211)
);

NOR2xp33_ASAP7_75t_L g1212 ( 
.A(n_1077),
.B(n_1044),
.Y(n_1212)
);

INVx1_ASAP7_75t_L g1213 ( 
.A(n_1095),
.Y(n_1213)
);

BUFx6f_ASAP7_75t_L g1214 ( 
.A(n_1088),
.Y(n_1214)
);

HB1xp67_ASAP7_75t_L g1215 ( 
.A(n_1157),
.Y(n_1215)
);

NAND2x1p5_ASAP7_75t_L g1216 ( 
.A(n_1110),
.B(n_1107),
.Y(n_1216)
);

INVx1_ASAP7_75t_L g1217 ( 
.A(n_1092),
.Y(n_1217)
);

CKINVDCx20_ASAP7_75t_R g1218 ( 
.A(n_1052),
.Y(n_1218)
);

BUFx2_ASAP7_75t_L g1219 ( 
.A(n_1088),
.Y(n_1219)
);

OAI22xp5_ASAP7_75t_L g1220 ( 
.A1(n_1084),
.A2(n_1088),
.B1(n_1130),
.B2(n_1160),
.Y(n_1220)
);

HB1xp67_ASAP7_75t_L g1221 ( 
.A(n_1132),
.Y(n_1221)
);

INVx2_ASAP7_75t_SL g1222 ( 
.A(n_1059),
.Y(n_1222)
);

BUFx2_ASAP7_75t_L g1223 ( 
.A(n_1143),
.Y(n_1223)
);

BUFx2_ASAP7_75t_L g1224 ( 
.A(n_1144),
.Y(n_1224)
);

BUFx3_ASAP7_75t_L g1225 ( 
.A(n_1093),
.Y(n_1225)
);

BUFx2_ASAP7_75t_L g1226 ( 
.A(n_1078),
.Y(n_1226)
);

AOI22xp33_ASAP7_75t_SL g1227 ( 
.A1(n_1082),
.A2(n_1161),
.B1(n_1156),
.B2(n_1080),
.Y(n_1227)
);

NAND2x1p5_ASAP7_75t_L g1228 ( 
.A(n_1107),
.B(n_1105),
.Y(n_1228)
);

INVx1_ASAP7_75t_L g1229 ( 
.A(n_1094),
.Y(n_1229)
);

INVx1_ASAP7_75t_L g1230 ( 
.A(n_1096),
.Y(n_1230)
);

INVxp33_ASAP7_75t_L g1231 ( 
.A(n_1036),
.Y(n_1231)
);

AOI22xp33_ASAP7_75t_SL g1232 ( 
.A1(n_1086),
.A2(n_1050),
.B1(n_1042),
.B2(n_1064),
.Y(n_1232)
);

INVx3_ASAP7_75t_L g1233 ( 
.A(n_1117),
.Y(n_1233)
);

INVx2_ASAP7_75t_L g1234 ( 
.A(n_1107),
.Y(n_1234)
);

BUFx3_ASAP7_75t_L g1235 ( 
.A(n_1033),
.Y(n_1235)
);

AND2x2_ASAP7_75t_L g1236 ( 
.A(n_1039),
.B(n_1086),
.Y(n_1236)
);

AO21x1_ASAP7_75t_SL g1237 ( 
.A1(n_1099),
.A2(n_1089),
.B(n_1103),
.Y(n_1237)
);

OAI22xp33_ASAP7_75t_L g1238 ( 
.A1(n_1068),
.A2(n_1075),
.B1(n_1090),
.B2(n_1106),
.Y(n_1238)
);

CKINVDCx5p33_ASAP7_75t_R g1239 ( 
.A(n_1068),
.Y(n_1239)
);

AOI22xp33_ASAP7_75t_SL g1240 ( 
.A1(n_1064),
.A2(n_1089),
.B1(n_1068),
.B2(n_1073),
.Y(n_1240)
);

OAI22xp5_ASAP7_75t_L g1241 ( 
.A1(n_1070),
.A2(n_1125),
.B1(n_1112),
.B2(n_1126),
.Y(n_1241)
);

INVx1_ASAP7_75t_L g1242 ( 
.A(n_1073),
.Y(n_1242)
);

BUFx6f_ASAP7_75t_L g1243 ( 
.A(n_1098),
.Y(n_1243)
);

BUFx2_ASAP7_75t_SL g1244 ( 
.A(n_1037),
.Y(n_1244)
);

AND2x2_ASAP7_75t_L g1245 ( 
.A(n_1129),
.B(n_1118),
.Y(n_1245)
);

INVx1_ASAP7_75t_L g1246 ( 
.A(n_1125),
.Y(n_1246)
);

AOI22xp33_ASAP7_75t_L g1247 ( 
.A1(n_1071),
.A2(n_1085),
.B1(n_1112),
.B2(n_1127),
.Y(n_1247)
);

AOI22xp33_ASAP7_75t_L g1248 ( 
.A1(n_1033),
.A2(n_1127),
.B1(n_1126),
.B2(n_1147),
.Y(n_1248)
);

BUFx2_ASAP7_75t_L g1249 ( 
.A(n_1037),
.Y(n_1249)
);

NAND2xp5_ASAP7_75t_L g1250 ( 
.A(n_1146),
.B(n_1145),
.Y(n_1250)
);

BUFx2_ASAP7_75t_L g1251 ( 
.A(n_1046),
.Y(n_1251)
);

INVx1_ASAP7_75t_L g1252 ( 
.A(n_1087),
.Y(n_1252)
);

INVx2_ASAP7_75t_L g1253 ( 
.A(n_1104),
.Y(n_1253)
);

AOI22xp33_ASAP7_75t_SL g1254 ( 
.A1(n_1140),
.A2(n_1102),
.B1(n_1046),
.B2(n_1109),
.Y(n_1254)
);

INVxp67_ASAP7_75t_L g1255 ( 
.A(n_1066),
.Y(n_1255)
);

INVx4_ASAP7_75t_L g1256 ( 
.A(n_1114),
.Y(n_1256)
);

NAND2xp5_ASAP7_75t_L g1257 ( 
.A(n_1116),
.B(n_1151),
.Y(n_1257)
);

AOI22xp33_ASAP7_75t_SL g1258 ( 
.A1(n_1116),
.A2(n_813),
.B1(n_790),
.B2(n_949),
.Y(n_1258)
);

AND2x2_ASAP7_75t_L g1259 ( 
.A(n_1054),
.B(n_1053),
.Y(n_1259)
);

AND2x2_ASAP7_75t_L g1260 ( 
.A(n_1054),
.B(n_1053),
.Y(n_1260)
);

INVx1_ASAP7_75t_L g1261 ( 
.A(n_1038),
.Y(n_1261)
);

BUFx10_ASAP7_75t_L g1262 ( 
.A(n_1066),
.Y(n_1262)
);

INVx1_ASAP7_75t_L g1263 ( 
.A(n_1038),
.Y(n_1263)
);

INVx1_ASAP7_75t_L g1264 ( 
.A(n_1038),
.Y(n_1264)
);

INVx1_ASAP7_75t_L g1265 ( 
.A(n_1038),
.Y(n_1265)
);

CKINVDCx5p33_ASAP7_75t_R g1266 ( 
.A(n_1122),
.Y(n_1266)
);

CKINVDCx6p67_ASAP7_75t_R g1267 ( 
.A(n_1079),
.Y(n_1267)
);

BUFx8_ASAP7_75t_L g1268 ( 
.A(n_1062),
.Y(n_1268)
);

AND2x2_ASAP7_75t_L g1269 ( 
.A(n_1054),
.B(n_1053),
.Y(n_1269)
);

AND2x2_ASAP7_75t_L g1270 ( 
.A(n_1054),
.B(n_1053),
.Y(n_1270)
);

BUFx2_ASAP7_75t_L g1271 ( 
.A(n_1063),
.Y(n_1271)
);

AOI22xp33_ASAP7_75t_SL g1272 ( 
.A1(n_1116),
.A2(n_813),
.B1(n_790),
.B2(n_949),
.Y(n_1272)
);

INVx3_ASAP7_75t_L g1273 ( 
.A(n_1091),
.Y(n_1273)
);

NAND2xp5_ASAP7_75t_L g1274 ( 
.A(n_1116),
.B(n_1151),
.Y(n_1274)
);

HB1xp67_ASAP7_75t_L g1275 ( 
.A(n_1223),
.Y(n_1275)
);

OR2x6_ASAP7_75t_L g1276 ( 
.A(n_1250),
.B(n_1163),
.Y(n_1276)
);

INVx1_ASAP7_75t_L g1277 ( 
.A(n_1171),
.Y(n_1277)
);

OAI21xp33_ASAP7_75t_SL g1278 ( 
.A1(n_1236),
.A2(n_1186),
.B(n_1183),
.Y(n_1278)
);

AND2x2_ASAP7_75t_L g1279 ( 
.A(n_1198),
.B(n_1182),
.Y(n_1279)
);

INVx3_ASAP7_75t_L g1280 ( 
.A(n_1216),
.Y(n_1280)
);

BUFx3_ASAP7_75t_L g1281 ( 
.A(n_1214),
.Y(n_1281)
);

INVx3_ASAP7_75t_L g1282 ( 
.A(n_1216),
.Y(n_1282)
);

AND2x2_ASAP7_75t_L g1283 ( 
.A(n_1182),
.B(n_1184),
.Y(n_1283)
);

INVx3_ASAP7_75t_L g1284 ( 
.A(n_1216),
.Y(n_1284)
);

AND2x4_ASAP7_75t_L g1285 ( 
.A(n_1175),
.B(n_1177),
.Y(n_1285)
);

INVx1_ASAP7_75t_L g1286 ( 
.A(n_1184),
.Y(n_1286)
);

OA21x2_ASAP7_75t_L g1287 ( 
.A1(n_1206),
.A2(n_1242),
.B(n_1245),
.Y(n_1287)
);

INVx2_ASAP7_75t_L g1288 ( 
.A(n_1201),
.Y(n_1288)
);

AND2x4_ASAP7_75t_L g1289 ( 
.A(n_1175),
.B(n_1177),
.Y(n_1289)
);

HB1xp67_ASAP7_75t_L g1290 ( 
.A(n_1224),
.Y(n_1290)
);

INVx2_ASAP7_75t_L g1291 ( 
.A(n_1201),
.Y(n_1291)
);

AND2x2_ASAP7_75t_L g1292 ( 
.A(n_1183),
.B(n_1186),
.Y(n_1292)
);

INVx1_ASAP7_75t_L g1293 ( 
.A(n_1253),
.Y(n_1293)
);

BUFx2_ASAP7_75t_SL g1294 ( 
.A(n_1243),
.Y(n_1294)
);

BUFx8_ASAP7_75t_SL g1295 ( 
.A(n_1180),
.Y(n_1295)
);

AO21x2_ASAP7_75t_L g1296 ( 
.A1(n_1245),
.A2(n_1220),
.B(n_1236),
.Y(n_1296)
);

AND2x4_ASAP7_75t_L g1297 ( 
.A(n_1175),
.B(n_1177),
.Y(n_1297)
);

AOI22xp5_ASAP7_75t_L g1298 ( 
.A1(n_1167),
.A2(n_1272),
.B1(n_1258),
.B2(n_1168),
.Y(n_1298)
);

INVx1_ASAP7_75t_L g1299 ( 
.A(n_1206),
.Y(n_1299)
);

AOI21x1_ASAP7_75t_L g1300 ( 
.A1(n_1205),
.A2(n_1234),
.B(n_1241),
.Y(n_1300)
);

AOI22xp33_ASAP7_75t_SL g1301 ( 
.A1(n_1190),
.A2(n_1274),
.B1(n_1257),
.B2(n_1259),
.Y(n_1301)
);

INVx2_ASAP7_75t_SL g1302 ( 
.A(n_1228),
.Y(n_1302)
);

NAND2xp5_ASAP7_75t_L g1303 ( 
.A(n_1259),
.B(n_1260),
.Y(n_1303)
);

OAI21xp5_ASAP7_75t_L g1304 ( 
.A1(n_1195),
.A2(n_1169),
.B(n_1199),
.Y(n_1304)
);

INVx1_ASAP7_75t_L g1305 ( 
.A(n_1260),
.Y(n_1305)
);

OR2x2_ASAP7_75t_L g1306 ( 
.A(n_1269),
.B(n_1270),
.Y(n_1306)
);

NOR2x1_ASAP7_75t_L g1307 ( 
.A(n_1204),
.B(n_1252),
.Y(n_1307)
);

INVx1_ASAP7_75t_L g1308 ( 
.A(n_1269),
.Y(n_1308)
);

AND2x2_ASAP7_75t_L g1309 ( 
.A(n_1270),
.B(n_1232),
.Y(n_1309)
);

HB1xp67_ASAP7_75t_L g1310 ( 
.A(n_1224),
.Y(n_1310)
);

AND2x2_ASAP7_75t_L g1311 ( 
.A(n_1240),
.B(n_1273),
.Y(n_1311)
);

OR2x2_ASAP7_75t_L g1312 ( 
.A(n_1165),
.B(n_1271),
.Y(n_1312)
);

INVx4_ASAP7_75t_L g1313 ( 
.A(n_1164),
.Y(n_1313)
);

HB1xp67_ASAP7_75t_L g1314 ( 
.A(n_1165),
.Y(n_1314)
);

INVx1_ASAP7_75t_L g1315 ( 
.A(n_1176),
.Y(n_1315)
);

BUFx2_ASAP7_75t_L g1316 ( 
.A(n_1219),
.Y(n_1316)
);

INVx2_ASAP7_75t_L g1317 ( 
.A(n_1193),
.Y(n_1317)
);

INVx2_ASAP7_75t_L g1318 ( 
.A(n_1196),
.Y(n_1318)
);

AND2x4_ASAP7_75t_L g1319 ( 
.A(n_1214),
.B(n_1208),
.Y(n_1319)
);

BUFx6f_ASAP7_75t_L g1320 ( 
.A(n_1214),
.Y(n_1320)
);

HB1xp67_ASAP7_75t_L g1321 ( 
.A(n_1271),
.Y(n_1321)
);

OAI22xp33_ASAP7_75t_L g1322 ( 
.A1(n_1231),
.A2(n_1162),
.B1(n_1255),
.B2(n_1239),
.Y(n_1322)
);

HB1xp67_ASAP7_75t_SL g1323 ( 
.A(n_1268),
.Y(n_1323)
);

HB1xp67_ASAP7_75t_L g1324 ( 
.A(n_1226),
.Y(n_1324)
);

INVx1_ASAP7_75t_L g1325 ( 
.A(n_1172),
.Y(n_1325)
);

NAND2xp5_ASAP7_75t_L g1326 ( 
.A(n_1170),
.B(n_1181),
.Y(n_1326)
);

AND2x4_ASAP7_75t_L g1327 ( 
.A(n_1214),
.B(n_1219),
.Y(n_1327)
);

HB1xp67_ASAP7_75t_L g1328 ( 
.A(n_1226),
.Y(n_1328)
);

OAI21x1_ASAP7_75t_L g1329 ( 
.A1(n_1248),
.A2(n_1246),
.B(n_1233),
.Y(n_1329)
);

OR2x2_ASAP7_75t_L g1330 ( 
.A(n_1179),
.B(n_1221),
.Y(n_1330)
);

INVx1_ASAP7_75t_L g1331 ( 
.A(n_1174),
.Y(n_1331)
);

OAI21xp5_ASAP7_75t_L g1332 ( 
.A1(n_1227),
.A2(n_1254),
.B(n_1231),
.Y(n_1332)
);

BUFx2_ASAP7_75t_L g1333 ( 
.A(n_1239),
.Y(n_1333)
);

AND2x2_ASAP7_75t_L g1334 ( 
.A(n_1237),
.B(n_1265),
.Y(n_1334)
);

AND2x2_ASAP7_75t_L g1335 ( 
.A(n_1237),
.B(n_1263),
.Y(n_1335)
);

BUFx8_ASAP7_75t_SL g1336 ( 
.A(n_1180),
.Y(n_1336)
);

INVx2_ASAP7_75t_L g1337 ( 
.A(n_1261),
.Y(n_1337)
);

INVx1_ASAP7_75t_L g1338 ( 
.A(n_1264),
.Y(n_1338)
);

NAND2xp5_ASAP7_75t_L g1339 ( 
.A(n_1238),
.B(n_1211),
.Y(n_1339)
);

HB1xp67_ASAP7_75t_SL g1340 ( 
.A(n_1268),
.Y(n_1340)
);

INVx1_ASAP7_75t_L g1341 ( 
.A(n_1203),
.Y(n_1341)
);

INVx1_ASAP7_75t_L g1342 ( 
.A(n_1213),
.Y(n_1342)
);

NAND2xp5_ASAP7_75t_L g1343 ( 
.A(n_1292),
.B(n_1262),
.Y(n_1343)
);

OAI21xp33_ASAP7_75t_L g1344 ( 
.A1(n_1298),
.A2(n_1212),
.B(n_1166),
.Y(n_1344)
);

NAND2xp5_ASAP7_75t_L g1345 ( 
.A(n_1303),
.B(n_1305),
.Y(n_1345)
);

AND2x4_ASAP7_75t_L g1346 ( 
.A(n_1280),
.B(n_1243),
.Y(n_1346)
);

OR2x2_ASAP7_75t_L g1347 ( 
.A(n_1288),
.B(n_1291),
.Y(n_1347)
);

AND2x2_ASAP7_75t_L g1348 ( 
.A(n_1306),
.B(n_1217),
.Y(n_1348)
);

INVx1_ASAP7_75t_L g1349 ( 
.A(n_1277),
.Y(n_1349)
);

INVx5_ASAP7_75t_L g1350 ( 
.A(n_1276),
.Y(n_1350)
);

BUFx3_ASAP7_75t_L g1351 ( 
.A(n_1319),
.Y(n_1351)
);

BUFx3_ASAP7_75t_L g1352 ( 
.A(n_1319),
.Y(n_1352)
);

AND2x2_ASAP7_75t_L g1353 ( 
.A(n_1306),
.B(n_1229),
.Y(n_1353)
);

BUFx3_ASAP7_75t_L g1354 ( 
.A(n_1319),
.Y(n_1354)
);

AND2x2_ASAP7_75t_L g1355 ( 
.A(n_1303),
.B(n_1230),
.Y(n_1355)
);

AND2x2_ASAP7_75t_L g1356 ( 
.A(n_1305),
.B(n_1262),
.Y(n_1356)
);

NOR2xp33_ASAP7_75t_R g1357 ( 
.A(n_1323),
.B(n_1266),
.Y(n_1357)
);

AOI221xp5_ASAP7_75t_L g1358 ( 
.A1(n_1304),
.A2(n_1215),
.B1(n_1173),
.B2(n_1210),
.C(n_1192),
.Y(n_1358)
);

AND2x2_ASAP7_75t_L g1359 ( 
.A(n_1308),
.B(n_1296),
.Y(n_1359)
);

AND2x2_ASAP7_75t_L g1360 ( 
.A(n_1308),
.B(n_1262),
.Y(n_1360)
);

HB1xp67_ASAP7_75t_L g1361 ( 
.A(n_1314),
.Y(n_1361)
);

HB1xp67_ASAP7_75t_L g1362 ( 
.A(n_1321),
.Y(n_1362)
);

AND2x2_ASAP7_75t_L g1363 ( 
.A(n_1296),
.B(n_1194),
.Y(n_1363)
);

INVx1_ASAP7_75t_SL g1364 ( 
.A(n_1312),
.Y(n_1364)
);

OAI22xp33_ASAP7_75t_L g1365 ( 
.A1(n_1298),
.A2(n_1235),
.B1(n_1218),
.B2(n_1243),
.Y(n_1365)
);

AOI22xp33_ASAP7_75t_SL g1366 ( 
.A1(n_1304),
.A2(n_1218),
.B1(n_1209),
.B2(n_1207),
.Y(n_1366)
);

AND2x2_ASAP7_75t_L g1367 ( 
.A(n_1296),
.B(n_1194),
.Y(n_1367)
);

OR2x2_ASAP7_75t_L g1368 ( 
.A(n_1288),
.B(n_1222),
.Y(n_1368)
);

INVx5_ASAP7_75t_L g1369 ( 
.A(n_1276),
.Y(n_1369)
);

AND2x2_ASAP7_75t_L g1370 ( 
.A(n_1296),
.B(n_1194),
.Y(n_1370)
);

BUFx3_ASAP7_75t_L g1371 ( 
.A(n_1319),
.Y(n_1371)
);

OAI211xp5_ASAP7_75t_SL g1372 ( 
.A1(n_1301),
.A2(n_1247),
.B(n_1222),
.C(n_1185),
.Y(n_1372)
);

OAI22xp33_ASAP7_75t_L g1373 ( 
.A1(n_1326),
.A2(n_1235),
.B1(n_1197),
.B2(n_1267),
.Y(n_1373)
);

AOI22xp33_ASAP7_75t_L g1374 ( 
.A1(n_1301),
.A2(n_1189),
.B1(n_1209),
.B2(n_1207),
.Y(n_1374)
);

AND2x2_ASAP7_75t_L g1375 ( 
.A(n_1279),
.B(n_1249),
.Y(n_1375)
);

INVxp67_ASAP7_75t_L g1376 ( 
.A(n_1307),
.Y(n_1376)
);

AOI22xp5_ASAP7_75t_L g1377 ( 
.A1(n_1326),
.A2(n_1267),
.B1(n_1197),
.B2(n_1191),
.Y(n_1377)
);

HB1xp67_ASAP7_75t_L g1378 ( 
.A(n_1324),
.Y(n_1378)
);

AND2x2_ASAP7_75t_L g1379 ( 
.A(n_1283),
.B(n_1251),
.Y(n_1379)
);

OAI221xp5_ASAP7_75t_L g1380 ( 
.A1(n_1332),
.A2(n_1187),
.B1(n_1202),
.B2(n_1225),
.C(n_1188),
.Y(n_1380)
);

AND2x2_ASAP7_75t_L g1381 ( 
.A(n_1283),
.B(n_1225),
.Y(n_1381)
);

OR2x2_ASAP7_75t_L g1382 ( 
.A(n_1291),
.B(n_1202),
.Y(n_1382)
);

INVxp67_ASAP7_75t_L g1383 ( 
.A(n_1307),
.Y(n_1383)
);

AOI221xp5_ASAP7_75t_L g1384 ( 
.A1(n_1332),
.A2(n_1187),
.B1(n_1266),
.B2(n_1244),
.C(n_1164),
.Y(n_1384)
);

INVxp67_ASAP7_75t_L g1385 ( 
.A(n_1328),
.Y(n_1385)
);

AND2x2_ASAP7_75t_L g1386 ( 
.A(n_1291),
.B(n_1276),
.Y(n_1386)
);

NAND2xp5_ASAP7_75t_L g1387 ( 
.A(n_1364),
.B(n_1312),
.Y(n_1387)
);

OAI22xp33_ASAP7_75t_L g1388 ( 
.A1(n_1380),
.A2(n_1339),
.B1(n_1330),
.B2(n_1276),
.Y(n_1388)
);

NAND2xp5_ASAP7_75t_L g1389 ( 
.A(n_1364),
.B(n_1275),
.Y(n_1389)
);

AND2x2_ASAP7_75t_L g1390 ( 
.A(n_1363),
.B(n_1287),
.Y(n_1390)
);

NOR2xp33_ASAP7_75t_L g1391 ( 
.A(n_1344),
.B(n_1322),
.Y(n_1391)
);

AND2x2_ASAP7_75t_L g1392 ( 
.A(n_1363),
.B(n_1287),
.Y(n_1392)
);

NAND3xp33_ASAP7_75t_L g1393 ( 
.A(n_1358),
.B(n_1339),
.C(n_1276),
.Y(n_1393)
);

OAI221xp5_ASAP7_75t_SL g1394 ( 
.A1(n_1344),
.A2(n_1278),
.B1(n_1309),
.B2(n_1330),
.C(n_1311),
.Y(n_1394)
);

AND2x2_ASAP7_75t_L g1395 ( 
.A(n_1367),
.B(n_1287),
.Y(n_1395)
);

NAND4xp25_ASAP7_75t_L g1396 ( 
.A(n_1358),
.B(n_1316),
.C(n_1309),
.D(n_1315),
.Y(n_1396)
);

OAI22xp5_ASAP7_75t_L g1397 ( 
.A1(n_1366),
.A2(n_1323),
.B1(n_1340),
.B2(n_1333),
.Y(n_1397)
);

AND2x2_ASAP7_75t_L g1398 ( 
.A(n_1367),
.B(n_1287),
.Y(n_1398)
);

AND2x2_ASAP7_75t_L g1399 ( 
.A(n_1370),
.B(n_1280),
.Y(n_1399)
);

NAND2xp5_ASAP7_75t_L g1400 ( 
.A(n_1355),
.B(n_1290),
.Y(n_1400)
);

NAND2xp5_ASAP7_75t_L g1401 ( 
.A(n_1343),
.B(n_1361),
.Y(n_1401)
);

OAI22xp5_ASAP7_75t_L g1402 ( 
.A1(n_1366),
.A2(n_1374),
.B1(n_1365),
.B2(n_1384),
.Y(n_1402)
);

NAND2xp5_ASAP7_75t_L g1403 ( 
.A(n_1343),
.B(n_1310),
.Y(n_1403)
);

OAI31xp33_ASAP7_75t_SL g1404 ( 
.A1(n_1372),
.A2(n_1311),
.A3(n_1327),
.B(n_1334),
.Y(n_1404)
);

AND2x2_ASAP7_75t_L g1405 ( 
.A(n_1370),
.B(n_1359),
.Y(n_1405)
);

NAND2xp5_ASAP7_75t_L g1406 ( 
.A(n_1362),
.B(n_1286),
.Y(n_1406)
);

NAND2xp5_ASAP7_75t_L g1407 ( 
.A(n_1378),
.B(n_1316),
.Y(n_1407)
);

NOR3xp33_ASAP7_75t_L g1408 ( 
.A(n_1373),
.B(n_1300),
.C(n_1278),
.Y(n_1408)
);

NAND3xp33_ASAP7_75t_SL g1409 ( 
.A(n_1384),
.B(n_1333),
.C(n_1334),
.Y(n_1409)
);

NAND3xp33_ASAP7_75t_L g1410 ( 
.A(n_1380),
.B(n_1341),
.C(n_1325),
.Y(n_1410)
);

AOI21xp33_ASAP7_75t_L g1411 ( 
.A1(n_1376),
.A2(n_1335),
.B(n_1302),
.Y(n_1411)
);

OAI21xp5_ASAP7_75t_L g1412 ( 
.A1(n_1376),
.A2(n_1329),
.B(n_1335),
.Y(n_1412)
);

NAND2xp5_ASAP7_75t_L g1413 ( 
.A(n_1348),
.B(n_1317),
.Y(n_1413)
);

NAND3xp33_ASAP7_75t_L g1414 ( 
.A(n_1383),
.B(n_1341),
.C(n_1325),
.Y(n_1414)
);

NAND3xp33_ASAP7_75t_L g1415 ( 
.A(n_1383),
.B(n_1331),
.C(n_1338),
.Y(n_1415)
);

NAND2xp5_ASAP7_75t_L g1416 ( 
.A(n_1353),
.B(n_1317),
.Y(n_1416)
);

AND2x2_ASAP7_75t_L g1417 ( 
.A(n_1386),
.B(n_1282),
.Y(n_1417)
);

NAND2xp5_ASAP7_75t_L g1418 ( 
.A(n_1353),
.B(n_1318),
.Y(n_1418)
);

AOI21xp5_ASAP7_75t_SL g1419 ( 
.A1(n_1377),
.A2(n_1164),
.B(n_1320),
.Y(n_1419)
);

INVx1_ASAP7_75t_L g1420 ( 
.A(n_1349),
.Y(n_1420)
);

NAND2xp5_ASAP7_75t_L g1421 ( 
.A(n_1385),
.B(n_1318),
.Y(n_1421)
);

NOR3xp33_ASAP7_75t_L g1422 ( 
.A(n_1372),
.B(n_1300),
.C(n_1313),
.Y(n_1422)
);

AND2x2_ASAP7_75t_L g1423 ( 
.A(n_1386),
.B(n_1282),
.Y(n_1423)
);

NAND3xp33_ASAP7_75t_L g1424 ( 
.A(n_1377),
.B(n_1331),
.C(n_1338),
.Y(n_1424)
);

NAND2xp5_ASAP7_75t_L g1425 ( 
.A(n_1385),
.B(n_1318),
.Y(n_1425)
);

OAI21xp5_ASAP7_75t_SL g1426 ( 
.A1(n_1356),
.A2(n_1340),
.B(n_1327),
.Y(n_1426)
);

NOR2xp33_ASAP7_75t_L g1427 ( 
.A(n_1381),
.B(n_1382),
.Y(n_1427)
);

AND2x2_ASAP7_75t_L g1428 ( 
.A(n_1351),
.B(n_1284),
.Y(n_1428)
);

OAI22xp5_ASAP7_75t_L g1429 ( 
.A1(n_1350),
.A2(n_1369),
.B1(n_1299),
.B2(n_1327),
.Y(n_1429)
);

AND2x2_ASAP7_75t_L g1430 ( 
.A(n_1351),
.B(n_1284),
.Y(n_1430)
);

INVxp67_ASAP7_75t_L g1431 ( 
.A(n_1368),
.Y(n_1431)
);

AND2x2_ASAP7_75t_L g1432 ( 
.A(n_1352),
.B(n_1354),
.Y(n_1432)
);

NAND2xp5_ASAP7_75t_L g1433 ( 
.A(n_1345),
.B(n_1315),
.Y(n_1433)
);

AOI22xp33_ASAP7_75t_L g1434 ( 
.A1(n_1356),
.A2(n_1327),
.B1(n_1289),
.B2(n_1285),
.Y(n_1434)
);

AOI22xp33_ASAP7_75t_L g1435 ( 
.A1(n_1360),
.A2(n_1289),
.B1(n_1285),
.B2(n_1297),
.Y(n_1435)
);

NAND2xp5_ASAP7_75t_L g1436 ( 
.A(n_1345),
.B(n_1337),
.Y(n_1436)
);

OAI22xp5_ASAP7_75t_L g1437 ( 
.A1(n_1350),
.A2(n_1294),
.B1(n_1281),
.B2(n_1178),
.Y(n_1437)
);

NAND3xp33_ASAP7_75t_L g1438 ( 
.A(n_1350),
.B(n_1342),
.C(n_1293),
.Y(n_1438)
);

OAI22xp5_ASAP7_75t_L g1439 ( 
.A1(n_1350),
.A2(n_1294),
.B1(n_1281),
.B2(n_1178),
.Y(n_1439)
);

OAI22xp5_ASAP7_75t_L g1440 ( 
.A1(n_1350),
.A2(n_1281),
.B1(n_1178),
.B2(n_1320),
.Y(n_1440)
);

OR2x2_ASAP7_75t_L g1441 ( 
.A(n_1390),
.B(n_1347),
.Y(n_1441)
);

NAND2xp5_ASAP7_75t_SL g1442 ( 
.A(n_1397),
.B(n_1357),
.Y(n_1442)
);

BUFx3_ASAP7_75t_L g1443 ( 
.A(n_1407),
.Y(n_1443)
);

NOR2x1_ASAP7_75t_L g1444 ( 
.A(n_1419),
.B(n_1368),
.Y(n_1444)
);

AND2x4_ASAP7_75t_L g1445 ( 
.A(n_1438),
.B(n_1350),
.Y(n_1445)
);

NAND2xp5_ASAP7_75t_L g1446 ( 
.A(n_1401),
.B(n_1379),
.Y(n_1446)
);

AND2x2_ASAP7_75t_L g1447 ( 
.A(n_1405),
.B(n_1350),
.Y(n_1447)
);

INVx1_ASAP7_75t_L g1448 ( 
.A(n_1420),
.Y(n_1448)
);

INVx1_ASAP7_75t_L g1449 ( 
.A(n_1420),
.Y(n_1449)
);

AND2x2_ASAP7_75t_L g1450 ( 
.A(n_1405),
.B(n_1369),
.Y(n_1450)
);

NAND2xp5_ASAP7_75t_L g1451 ( 
.A(n_1403),
.B(n_1379),
.Y(n_1451)
);

AND2x4_ASAP7_75t_L g1452 ( 
.A(n_1438),
.B(n_1369),
.Y(n_1452)
);

INVx1_ASAP7_75t_L g1453 ( 
.A(n_1421),
.Y(n_1453)
);

INVx1_ASAP7_75t_L g1454 ( 
.A(n_1425),
.Y(n_1454)
);

INVx1_ASAP7_75t_L g1455 ( 
.A(n_1414),
.Y(n_1455)
);

INVx1_ASAP7_75t_L g1456 ( 
.A(n_1414),
.Y(n_1456)
);

INVx1_ASAP7_75t_L g1457 ( 
.A(n_1415),
.Y(n_1457)
);

AND2x4_ASAP7_75t_SL g1458 ( 
.A(n_1408),
.B(n_1346),
.Y(n_1458)
);

INVx6_ASAP7_75t_L g1459 ( 
.A(n_1432),
.Y(n_1459)
);

AND2x2_ASAP7_75t_L g1460 ( 
.A(n_1390),
.B(n_1369),
.Y(n_1460)
);

INVxp67_ASAP7_75t_SL g1461 ( 
.A(n_1415),
.Y(n_1461)
);

NAND2xp5_ASAP7_75t_SL g1462 ( 
.A(n_1424),
.B(n_1346),
.Y(n_1462)
);

AND2x2_ASAP7_75t_L g1463 ( 
.A(n_1392),
.B(n_1369),
.Y(n_1463)
);

INVx1_ASAP7_75t_L g1464 ( 
.A(n_1392),
.Y(n_1464)
);

AND2x2_ASAP7_75t_L g1465 ( 
.A(n_1395),
.B(n_1369),
.Y(n_1465)
);

NAND2xp5_ASAP7_75t_L g1466 ( 
.A(n_1387),
.B(n_1360),
.Y(n_1466)
);

NAND2xp5_ASAP7_75t_L g1467 ( 
.A(n_1389),
.B(n_1375),
.Y(n_1467)
);

INVx1_ASAP7_75t_L g1468 ( 
.A(n_1395),
.Y(n_1468)
);

BUFx2_ASAP7_75t_SL g1469 ( 
.A(n_1428),
.Y(n_1469)
);

BUFx2_ASAP7_75t_L g1470 ( 
.A(n_1399),
.Y(n_1470)
);

INVx1_ASAP7_75t_L g1471 ( 
.A(n_1398),
.Y(n_1471)
);

INVx2_ASAP7_75t_L g1472 ( 
.A(n_1398),
.Y(n_1472)
);

INVx5_ASAP7_75t_L g1473 ( 
.A(n_1430),
.Y(n_1473)
);

INVx1_ASAP7_75t_L g1474 ( 
.A(n_1431),
.Y(n_1474)
);

NAND2xp5_ASAP7_75t_L g1475 ( 
.A(n_1400),
.B(n_1375),
.Y(n_1475)
);

AOI22xp33_ASAP7_75t_L g1476 ( 
.A1(n_1391),
.A2(n_1369),
.B1(n_1371),
.B2(n_1289),
.Y(n_1476)
);

INVx1_ASAP7_75t_L g1477 ( 
.A(n_1406),
.Y(n_1477)
);

INVx1_ASAP7_75t_L g1478 ( 
.A(n_1448),
.Y(n_1478)
);

OR2x2_ASAP7_75t_L g1479 ( 
.A(n_1461),
.B(n_1413),
.Y(n_1479)
);

INVx1_ASAP7_75t_L g1480 ( 
.A(n_1448),
.Y(n_1480)
);

INVx2_ASAP7_75t_L g1481 ( 
.A(n_1449),
.Y(n_1481)
);

INVx1_ASAP7_75t_L g1482 ( 
.A(n_1449),
.Y(n_1482)
);

INVx2_ASAP7_75t_L g1483 ( 
.A(n_1472),
.Y(n_1483)
);

AND2x2_ASAP7_75t_L g1484 ( 
.A(n_1469),
.B(n_1432),
.Y(n_1484)
);

INVx2_ASAP7_75t_L g1485 ( 
.A(n_1472),
.Y(n_1485)
);

NAND2xp5_ASAP7_75t_L g1486 ( 
.A(n_1455),
.B(n_1433),
.Y(n_1486)
);

AND2x4_ASAP7_75t_L g1487 ( 
.A(n_1473),
.B(n_1412),
.Y(n_1487)
);

AND2x2_ASAP7_75t_L g1488 ( 
.A(n_1469),
.B(n_1417),
.Y(n_1488)
);

INVx1_ASAP7_75t_L g1489 ( 
.A(n_1441),
.Y(n_1489)
);

AND2x2_ASAP7_75t_L g1490 ( 
.A(n_1473),
.B(n_1423),
.Y(n_1490)
);

INVx2_ASAP7_75t_L g1491 ( 
.A(n_1464),
.Y(n_1491)
);

OAI21xp33_ASAP7_75t_L g1492 ( 
.A1(n_1455),
.A2(n_1396),
.B(n_1393),
.Y(n_1492)
);

NAND2xp5_ASAP7_75t_L g1493 ( 
.A(n_1456),
.B(n_1436),
.Y(n_1493)
);

INVx1_ASAP7_75t_L g1494 ( 
.A(n_1441),
.Y(n_1494)
);

INVx1_ASAP7_75t_L g1495 ( 
.A(n_1474),
.Y(n_1495)
);

NAND2xp5_ASAP7_75t_L g1496 ( 
.A(n_1456),
.B(n_1416),
.Y(n_1496)
);

INVx2_ASAP7_75t_L g1497 ( 
.A(n_1468),
.Y(n_1497)
);

NAND2xp5_ASAP7_75t_L g1498 ( 
.A(n_1457),
.B(n_1418),
.Y(n_1498)
);

AND2x2_ASAP7_75t_L g1499 ( 
.A(n_1473),
.B(n_1423),
.Y(n_1499)
);

AND2x2_ASAP7_75t_L g1500 ( 
.A(n_1473),
.B(n_1427),
.Y(n_1500)
);

NOR3xp33_ASAP7_75t_L g1501 ( 
.A(n_1442),
.B(n_1402),
.C(n_1393),
.Y(n_1501)
);

INVx2_ASAP7_75t_L g1502 ( 
.A(n_1468),
.Y(n_1502)
);

OR2x2_ASAP7_75t_L g1503 ( 
.A(n_1471),
.B(n_1457),
.Y(n_1503)
);

OAI21xp33_ASAP7_75t_L g1504 ( 
.A1(n_1462),
.A2(n_1394),
.B(n_1409),
.Y(n_1504)
);

INVx1_ASAP7_75t_L g1505 ( 
.A(n_1474),
.Y(n_1505)
);

OAI21xp33_ASAP7_75t_SL g1506 ( 
.A1(n_1444),
.A2(n_1419),
.B(n_1404),
.Y(n_1506)
);

OR2x6_ASAP7_75t_L g1507 ( 
.A(n_1445),
.B(n_1410),
.Y(n_1507)
);

INVx2_ASAP7_75t_L g1508 ( 
.A(n_1470),
.Y(n_1508)
);

INVx2_ASAP7_75t_L g1509 ( 
.A(n_1470),
.Y(n_1509)
);

AND2x2_ASAP7_75t_L g1510 ( 
.A(n_1473),
.B(n_1371),
.Y(n_1510)
);

AND2x2_ASAP7_75t_L g1511 ( 
.A(n_1473),
.B(n_1447),
.Y(n_1511)
);

AND2x2_ASAP7_75t_L g1512 ( 
.A(n_1447),
.B(n_1429),
.Y(n_1512)
);

OR2x2_ASAP7_75t_L g1513 ( 
.A(n_1453),
.B(n_1454),
.Y(n_1513)
);

NAND2xp5_ASAP7_75t_L g1514 ( 
.A(n_1504),
.B(n_1492),
.Y(n_1514)
);

NOR2xp67_ASAP7_75t_L g1515 ( 
.A(n_1506),
.B(n_1445),
.Y(n_1515)
);

INVx1_ASAP7_75t_L g1516 ( 
.A(n_1478),
.Y(n_1516)
);

INVx1_ASAP7_75t_L g1517 ( 
.A(n_1478),
.Y(n_1517)
);

NAND2x1p5_ASAP7_75t_L g1518 ( 
.A(n_1487),
.B(n_1445),
.Y(n_1518)
);

INVx1_ASAP7_75t_L g1519 ( 
.A(n_1480),
.Y(n_1519)
);

INVxp67_ASAP7_75t_SL g1520 ( 
.A(n_1486),
.Y(n_1520)
);

AND2x2_ASAP7_75t_L g1521 ( 
.A(n_1511),
.B(n_1512),
.Y(n_1521)
);

INVx2_ASAP7_75t_L g1522 ( 
.A(n_1481),
.Y(n_1522)
);

AND2x2_ASAP7_75t_L g1523 ( 
.A(n_1511),
.B(n_1460),
.Y(n_1523)
);

NAND2xp5_ASAP7_75t_L g1524 ( 
.A(n_1504),
.B(n_1477),
.Y(n_1524)
);

INVx1_ASAP7_75t_L g1525 ( 
.A(n_1480),
.Y(n_1525)
);

AND2x2_ASAP7_75t_L g1526 ( 
.A(n_1512),
.B(n_1460),
.Y(n_1526)
);

INVx1_ASAP7_75t_L g1527 ( 
.A(n_1482),
.Y(n_1527)
);

AND2x2_ASAP7_75t_L g1528 ( 
.A(n_1500),
.B(n_1463),
.Y(n_1528)
);

NOR2x1_ASAP7_75t_L g1529 ( 
.A(n_1507),
.B(n_1410),
.Y(n_1529)
);

NOR2xp67_ASAP7_75t_L g1530 ( 
.A(n_1506),
.B(n_1445),
.Y(n_1530)
);

INVx3_ASAP7_75t_L g1531 ( 
.A(n_1487),
.Y(n_1531)
);

AND2x2_ASAP7_75t_L g1532 ( 
.A(n_1500),
.B(n_1463),
.Y(n_1532)
);

INVx1_ASAP7_75t_L g1533 ( 
.A(n_1482),
.Y(n_1533)
);

OR2x2_ASAP7_75t_L g1534 ( 
.A(n_1503),
.B(n_1453),
.Y(n_1534)
);

A2O1A1Ixp33_ASAP7_75t_L g1535 ( 
.A1(n_1501),
.A2(n_1458),
.B(n_1424),
.C(n_1452),
.Y(n_1535)
);

OR2x2_ASAP7_75t_L g1536 ( 
.A(n_1503),
.B(n_1454),
.Y(n_1536)
);

OR2x2_ASAP7_75t_L g1537 ( 
.A(n_1479),
.B(n_1489),
.Y(n_1537)
);

INVxp67_ASAP7_75t_L g1538 ( 
.A(n_1486),
.Y(n_1538)
);

AND2x2_ASAP7_75t_L g1539 ( 
.A(n_1487),
.B(n_1465),
.Y(n_1539)
);

AOI32xp33_ASAP7_75t_SL g1540 ( 
.A1(n_1501),
.A2(n_1477),
.A3(n_1466),
.B1(n_1467),
.B2(n_1451),
.Y(n_1540)
);

AND2x2_ASAP7_75t_L g1541 ( 
.A(n_1487),
.B(n_1465),
.Y(n_1541)
);

NAND2xp5_ASAP7_75t_SL g1542 ( 
.A(n_1492),
.B(n_1452),
.Y(n_1542)
);

NOR3xp33_ASAP7_75t_L g1543 ( 
.A(n_1493),
.B(n_1388),
.C(n_1496),
.Y(n_1543)
);

INVx1_ASAP7_75t_L g1544 ( 
.A(n_1495),
.Y(n_1544)
);

AOI211xp5_ASAP7_75t_SL g1545 ( 
.A1(n_1493),
.A2(n_1437),
.B(n_1439),
.C(n_1440),
.Y(n_1545)
);

NAND2xp5_ASAP7_75t_L g1546 ( 
.A(n_1496),
.B(n_1443),
.Y(n_1546)
);

OR2x2_ASAP7_75t_L g1547 ( 
.A(n_1479),
.B(n_1446),
.Y(n_1547)
);

AND2x2_ASAP7_75t_L g1548 ( 
.A(n_1484),
.B(n_1450),
.Y(n_1548)
);

AND2x2_ASAP7_75t_L g1549 ( 
.A(n_1484),
.B(n_1450),
.Y(n_1549)
);

INVx1_ASAP7_75t_L g1550 ( 
.A(n_1495),
.Y(n_1550)
);

INVx1_ASAP7_75t_L g1551 ( 
.A(n_1505),
.Y(n_1551)
);

OR2x2_ASAP7_75t_L g1552 ( 
.A(n_1489),
.B(n_1494),
.Y(n_1552)
);

OR2x2_ASAP7_75t_L g1553 ( 
.A(n_1494),
.B(n_1475),
.Y(n_1553)
);

AOI22xp5_ASAP7_75t_L g1554 ( 
.A1(n_1507),
.A2(n_1458),
.B1(n_1426),
.B2(n_1422),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_1505),
.Y(n_1555)
);

INVx2_ASAP7_75t_SL g1556 ( 
.A(n_1508),
.Y(n_1556)
);

INVx1_ASAP7_75t_SL g1557 ( 
.A(n_1521),
.Y(n_1557)
);

NAND2xp5_ASAP7_75t_L g1558 ( 
.A(n_1514),
.B(n_1524),
.Y(n_1558)
);

AND2x2_ASAP7_75t_L g1559 ( 
.A(n_1515),
.B(n_1507),
.Y(n_1559)
);

INVx1_ASAP7_75t_L g1560 ( 
.A(n_1516),
.Y(n_1560)
);

INVx1_ASAP7_75t_L g1561 ( 
.A(n_1517),
.Y(n_1561)
);

INVx1_ASAP7_75t_SL g1562 ( 
.A(n_1521),
.Y(n_1562)
);

AND2x2_ASAP7_75t_L g1563 ( 
.A(n_1530),
.B(n_1507),
.Y(n_1563)
);

INVx1_ASAP7_75t_L g1564 ( 
.A(n_1544),
.Y(n_1564)
);

INVx2_ASAP7_75t_L g1565 ( 
.A(n_1556),
.Y(n_1565)
);

OA21x2_ASAP7_75t_L g1566 ( 
.A1(n_1542),
.A2(n_1481),
.B(n_1508),
.Y(n_1566)
);

INVx1_ASAP7_75t_L g1567 ( 
.A(n_1519),
.Y(n_1567)
);

NAND2xp5_ASAP7_75t_L g1568 ( 
.A(n_1543),
.B(n_1498),
.Y(n_1568)
);

OA21x2_ASAP7_75t_L g1569 ( 
.A1(n_1542),
.A2(n_1481),
.B(n_1508),
.Y(n_1569)
);

BUFx3_ASAP7_75t_L g1570 ( 
.A(n_1556),
.Y(n_1570)
);

AOI22xp5_ASAP7_75t_L g1571 ( 
.A1(n_1529),
.A2(n_1507),
.B1(n_1452),
.B2(n_1498),
.Y(n_1571)
);

INVx1_ASAP7_75t_L g1572 ( 
.A(n_1525),
.Y(n_1572)
);

INVx1_ASAP7_75t_L g1573 ( 
.A(n_1527),
.Y(n_1573)
);

INVx4_ASAP7_75t_L g1574 ( 
.A(n_1531),
.Y(n_1574)
);

INVx1_ASAP7_75t_L g1575 ( 
.A(n_1533),
.Y(n_1575)
);

INVx1_ASAP7_75t_L g1576 ( 
.A(n_1550),
.Y(n_1576)
);

AND2x2_ASAP7_75t_L g1577 ( 
.A(n_1526),
.B(n_1509),
.Y(n_1577)
);

INVx1_ASAP7_75t_L g1578 ( 
.A(n_1551),
.Y(n_1578)
);

OR2x2_ASAP7_75t_L g1579 ( 
.A(n_1537),
.B(n_1513),
.Y(n_1579)
);

AND2x2_ASAP7_75t_L g1580 ( 
.A(n_1526),
.B(n_1509),
.Y(n_1580)
);

AND2x2_ASAP7_75t_L g1581 ( 
.A(n_1523),
.B(n_1509),
.Y(n_1581)
);

INVx1_ASAP7_75t_L g1582 ( 
.A(n_1555),
.Y(n_1582)
);

INVx1_ASAP7_75t_L g1583 ( 
.A(n_1552),
.Y(n_1583)
);

OR2x2_ASAP7_75t_L g1584 ( 
.A(n_1537),
.B(n_1513),
.Y(n_1584)
);

AND2x2_ASAP7_75t_L g1585 ( 
.A(n_1523),
.B(n_1528),
.Y(n_1585)
);

OR2x2_ASAP7_75t_L g1586 ( 
.A(n_1552),
.B(n_1491),
.Y(n_1586)
);

CKINVDCx16_ASAP7_75t_R g1587 ( 
.A(n_1554),
.Y(n_1587)
);

AND2x2_ASAP7_75t_L g1588 ( 
.A(n_1528),
.B(n_1490),
.Y(n_1588)
);

AOI21xp5_ASAP7_75t_L g1589 ( 
.A1(n_1535),
.A2(n_1452),
.B(n_1510),
.Y(n_1589)
);

INVx1_ASAP7_75t_L g1590 ( 
.A(n_1534),
.Y(n_1590)
);

INVx1_ASAP7_75t_L g1591 ( 
.A(n_1534),
.Y(n_1591)
);

INVx1_ASAP7_75t_L g1592 ( 
.A(n_1536),
.Y(n_1592)
);

AOI22xp5_ASAP7_75t_L g1593 ( 
.A1(n_1587),
.A2(n_1535),
.B1(n_1538),
.B2(n_1520),
.Y(n_1593)
);

OAI21xp33_ASAP7_75t_SL g1594 ( 
.A1(n_1571),
.A2(n_1541),
.B(n_1539),
.Y(n_1594)
);

OAI21xp5_ASAP7_75t_L g1595 ( 
.A1(n_1558),
.A2(n_1545),
.B(n_1540),
.Y(n_1595)
);

XOR2x2_ASAP7_75t_L g1596 ( 
.A(n_1568),
.B(n_1518),
.Y(n_1596)
);

O2A1O1Ixp33_ASAP7_75t_L g1597 ( 
.A1(n_1589),
.A2(n_1531),
.B(n_1518),
.C(n_1546),
.Y(n_1597)
);

AND2x2_ASAP7_75t_L g1598 ( 
.A(n_1585),
.B(n_1548),
.Y(n_1598)
);

OAI22xp5_ASAP7_75t_L g1599 ( 
.A1(n_1566),
.A2(n_1531),
.B1(n_1547),
.B2(n_1476),
.Y(n_1599)
);

INVx1_ASAP7_75t_L g1600 ( 
.A(n_1560),
.Y(n_1600)
);

NAND2xp5_ASAP7_75t_L g1601 ( 
.A(n_1557),
.B(n_1548),
.Y(n_1601)
);

AOI22xp5_ASAP7_75t_L g1602 ( 
.A1(n_1562),
.A2(n_1539),
.B1(n_1541),
.B2(n_1532),
.Y(n_1602)
);

INVx1_ASAP7_75t_L g1603 ( 
.A(n_1560),
.Y(n_1603)
);

INVx1_ASAP7_75t_L g1604 ( 
.A(n_1561),
.Y(n_1604)
);

INVx2_ASAP7_75t_SL g1605 ( 
.A(n_1570),
.Y(n_1605)
);

NAND2xp5_ASAP7_75t_L g1606 ( 
.A(n_1585),
.B(n_1549),
.Y(n_1606)
);

INVx2_ASAP7_75t_SL g1607 ( 
.A(n_1570),
.Y(n_1607)
);

AND2x2_ASAP7_75t_L g1608 ( 
.A(n_1581),
.B(n_1549),
.Y(n_1608)
);

AOI211xp5_ASAP7_75t_SL g1609 ( 
.A1(n_1559),
.A2(n_1200),
.B(n_1532),
.C(n_1336),
.Y(n_1609)
);

INVx2_ASAP7_75t_L g1610 ( 
.A(n_1574),
.Y(n_1610)
);

NAND2xp5_ASAP7_75t_L g1611 ( 
.A(n_1583),
.B(n_1547),
.Y(n_1611)
);

INVxp67_ASAP7_75t_L g1612 ( 
.A(n_1559),
.Y(n_1612)
);

INVx1_ASAP7_75t_L g1613 ( 
.A(n_1561),
.Y(n_1613)
);

O2A1O1Ixp33_ASAP7_75t_L g1614 ( 
.A1(n_1563),
.A2(n_1536),
.B(n_1522),
.C(n_1553),
.Y(n_1614)
);

AOI22xp5_ASAP7_75t_L g1615 ( 
.A1(n_1563),
.A2(n_1510),
.B1(n_1459),
.B2(n_1553),
.Y(n_1615)
);

NAND3xp33_ASAP7_75t_L g1616 ( 
.A(n_1566),
.B(n_1522),
.C(n_1411),
.Y(n_1616)
);

NOR3xp33_ASAP7_75t_L g1617 ( 
.A(n_1574),
.B(n_1499),
.C(n_1490),
.Y(n_1617)
);

OAI22xp5_ASAP7_75t_L g1618 ( 
.A1(n_1566),
.A2(n_1459),
.B1(n_1443),
.B2(n_1499),
.Y(n_1618)
);

INVx1_ASAP7_75t_SL g1619 ( 
.A(n_1596),
.Y(n_1619)
);

NOR2xp33_ASAP7_75t_L g1620 ( 
.A(n_1612),
.B(n_1295),
.Y(n_1620)
);

NAND2xp5_ASAP7_75t_L g1621 ( 
.A(n_1605),
.B(n_1581),
.Y(n_1621)
);

INVx1_ASAP7_75t_L g1622 ( 
.A(n_1600),
.Y(n_1622)
);

INVxp67_ASAP7_75t_SL g1623 ( 
.A(n_1607),
.Y(n_1623)
);

NOR2xp33_ASAP7_75t_L g1624 ( 
.A(n_1595),
.B(n_1574),
.Y(n_1624)
);

INVx1_ASAP7_75t_L g1625 ( 
.A(n_1603),
.Y(n_1625)
);

NOR2xp33_ASAP7_75t_L g1626 ( 
.A(n_1595),
.B(n_1590),
.Y(n_1626)
);

AND2x2_ASAP7_75t_L g1627 ( 
.A(n_1609),
.B(n_1588),
.Y(n_1627)
);

NOR2xp33_ASAP7_75t_L g1628 ( 
.A(n_1594),
.B(n_1200),
.Y(n_1628)
);

INVx1_ASAP7_75t_L g1629 ( 
.A(n_1604),
.Y(n_1629)
);

NAND3xp33_ASAP7_75t_SL g1630 ( 
.A(n_1593),
.B(n_1565),
.C(n_1579),
.Y(n_1630)
);

NAND2xp5_ASAP7_75t_L g1631 ( 
.A(n_1598),
.B(n_1577),
.Y(n_1631)
);

OAI222xp33_ASAP7_75t_L g1632 ( 
.A1(n_1597),
.A2(n_1584),
.B1(n_1579),
.B2(n_1588),
.C1(n_1577),
.C2(n_1580),
.Y(n_1632)
);

BUFx2_ASAP7_75t_L g1633 ( 
.A(n_1610),
.Y(n_1633)
);

NAND2x1_ASAP7_75t_SL g1634 ( 
.A(n_1602),
.B(n_1566),
.Y(n_1634)
);

OR2x2_ASAP7_75t_L g1635 ( 
.A(n_1601),
.B(n_1584),
.Y(n_1635)
);

CKINVDCx20_ASAP7_75t_R g1636 ( 
.A(n_1615),
.Y(n_1636)
);

INVx1_ASAP7_75t_L g1637 ( 
.A(n_1613),
.Y(n_1637)
);

NOR2xp33_ASAP7_75t_R g1638 ( 
.A(n_1611),
.B(n_1268),
.Y(n_1638)
);

AOI221x1_ASAP7_75t_L g1639 ( 
.A1(n_1630),
.A2(n_1617),
.B1(n_1618),
.B2(n_1565),
.C(n_1599),
.Y(n_1639)
);

AOI221xp5_ASAP7_75t_L g1640 ( 
.A1(n_1626),
.A2(n_1599),
.B1(n_1618),
.B2(n_1614),
.C(n_1616),
.Y(n_1640)
);

NAND2xp5_ASAP7_75t_L g1641 ( 
.A(n_1623),
.B(n_1608),
.Y(n_1641)
);

OR2x2_ASAP7_75t_L g1642 ( 
.A(n_1631),
.B(n_1606),
.Y(n_1642)
);

NAND2xp5_ASAP7_75t_L g1643 ( 
.A(n_1633),
.B(n_1609),
.Y(n_1643)
);

NAND2xp5_ASAP7_75t_L g1644 ( 
.A(n_1626),
.B(n_1580),
.Y(n_1644)
);

O2A1O1Ixp33_ASAP7_75t_L g1645 ( 
.A1(n_1624),
.A2(n_1569),
.B(n_1582),
.C(n_1564),
.Y(n_1645)
);

AOI21xp5_ASAP7_75t_L g1646 ( 
.A1(n_1624),
.A2(n_1619),
.B(n_1632),
.Y(n_1646)
);

OAI21xp33_ASAP7_75t_L g1647 ( 
.A1(n_1634),
.A2(n_1591),
.B(n_1590),
.Y(n_1647)
);

NAND2xp5_ASAP7_75t_L g1648 ( 
.A(n_1627),
.B(n_1591),
.Y(n_1648)
);

AOI221xp5_ASAP7_75t_L g1649 ( 
.A1(n_1621),
.A2(n_1592),
.B1(n_1567),
.B2(n_1578),
.C(n_1576),
.Y(n_1649)
);

NAND2xp5_ASAP7_75t_L g1650 ( 
.A(n_1620),
.B(n_1592),
.Y(n_1650)
);

NOR2x1p5_ASAP7_75t_L g1651 ( 
.A(n_1643),
.B(n_1635),
.Y(n_1651)
);

NOR4xp75_ASAP7_75t_L g1652 ( 
.A(n_1641),
.B(n_1636),
.C(n_1638),
.D(n_1628),
.Y(n_1652)
);

OA22x2_ASAP7_75t_L g1653 ( 
.A1(n_1639),
.A2(n_1629),
.B1(n_1625),
.B2(n_1622),
.Y(n_1653)
);

NAND2xp5_ASAP7_75t_L g1654 ( 
.A(n_1646),
.B(n_1620),
.Y(n_1654)
);

NOR2x1p5_ASAP7_75t_L g1655 ( 
.A(n_1648),
.B(n_1637),
.Y(n_1655)
);

INVx1_ASAP7_75t_L g1656 ( 
.A(n_1642),
.Y(n_1656)
);

NOR3xp33_ASAP7_75t_L g1657 ( 
.A(n_1650),
.B(n_1572),
.C(n_1567),
.Y(n_1657)
);

NOR2xp33_ASAP7_75t_L g1658 ( 
.A(n_1644),
.B(n_1191),
.Y(n_1658)
);

NOR2xp33_ASAP7_75t_L g1659 ( 
.A(n_1647),
.B(n_1572),
.Y(n_1659)
);

NOR3xp33_ASAP7_75t_L g1660 ( 
.A(n_1640),
.B(n_1575),
.C(n_1573),
.Y(n_1660)
);

NAND2x1_ASAP7_75t_SL g1661 ( 
.A(n_1645),
.B(n_1569),
.Y(n_1661)
);

NAND4xp25_ASAP7_75t_L g1662 ( 
.A(n_1654),
.B(n_1649),
.C(n_1576),
.D(n_1578),
.Y(n_1662)
);

NOR3xp33_ASAP7_75t_L g1663 ( 
.A(n_1656),
.B(n_1575),
.C(n_1573),
.Y(n_1663)
);

AOI21xp5_ASAP7_75t_L g1664 ( 
.A1(n_1653),
.A2(n_1659),
.B(n_1660),
.Y(n_1664)
);

O2A1O1Ixp5_ASAP7_75t_L g1665 ( 
.A1(n_1658),
.A2(n_1586),
.B(n_1569),
.C(n_1491),
.Y(n_1665)
);

NOR2x1_ASAP7_75t_L g1666 ( 
.A(n_1651),
.B(n_1569),
.Y(n_1666)
);

NAND5xp2_ASAP7_75t_L g1667 ( 
.A(n_1657),
.B(n_1434),
.C(n_1435),
.D(n_1488),
.E(n_1381),
.Y(n_1667)
);

INVx1_ASAP7_75t_L g1668 ( 
.A(n_1666),
.Y(n_1668)
);

HB1xp67_ASAP7_75t_L g1669 ( 
.A(n_1662),
.Y(n_1669)
);

INVx1_ASAP7_75t_L g1670 ( 
.A(n_1663),
.Y(n_1670)
);

INVx2_ASAP7_75t_L g1671 ( 
.A(n_1665),
.Y(n_1671)
);

AND2x2_ASAP7_75t_L g1672 ( 
.A(n_1664),
.B(n_1655),
.Y(n_1672)
);

INVx1_ASAP7_75t_L g1673 ( 
.A(n_1667),
.Y(n_1673)
);

NOR2xp67_ASAP7_75t_L g1674 ( 
.A(n_1668),
.B(n_1586),
.Y(n_1674)
);

INVx2_ASAP7_75t_L g1675 ( 
.A(n_1670),
.Y(n_1675)
);

NOR2xp67_ASAP7_75t_L g1676 ( 
.A(n_1671),
.B(n_1652),
.Y(n_1676)
);

NAND2x1p5_ASAP7_75t_L g1677 ( 
.A(n_1672),
.B(n_1256),
.Y(n_1677)
);

NOR2x1_ASAP7_75t_L g1678 ( 
.A(n_1671),
.B(n_1661),
.Y(n_1678)
);

INVx1_ASAP7_75t_L g1679 ( 
.A(n_1674),
.Y(n_1679)
);

NAND3x1_ASAP7_75t_L g1680 ( 
.A(n_1678),
.B(n_1673),
.C(n_1669),
.Y(n_1680)
);

NAND2xp5_ASAP7_75t_L g1681 ( 
.A(n_1676),
.B(n_1669),
.Y(n_1681)
);

INVx1_ASAP7_75t_L g1682 ( 
.A(n_1679),
.Y(n_1682)
);

NAND3xp33_ASAP7_75t_SL g1683 ( 
.A(n_1682),
.B(n_1681),
.C(n_1677),
.Y(n_1683)
);

INVx2_ASAP7_75t_SL g1684 ( 
.A(n_1683),
.Y(n_1684)
);

AOI21xp5_ASAP7_75t_L g1685 ( 
.A1(n_1683),
.A2(n_1675),
.B(n_1680),
.Y(n_1685)
);

AOI22xp5_ASAP7_75t_L g1686 ( 
.A1(n_1684),
.A2(n_1459),
.B1(n_1502),
.B2(n_1497),
.Y(n_1686)
);

NOR2xp33_ASAP7_75t_L g1687 ( 
.A(n_1685),
.B(n_1459),
.Y(n_1687)
);

INVx1_ASAP7_75t_L g1688 ( 
.A(n_1687),
.Y(n_1688)
);

XNOR2xp5_ASAP7_75t_L g1689 ( 
.A(n_1686),
.B(n_1244),
.Y(n_1689)
);

XNOR2xp5_ASAP7_75t_L g1690 ( 
.A(n_1688),
.B(n_1488),
.Y(n_1690)
);

AOI322xp5_ASAP7_75t_L g1691 ( 
.A1(n_1690),
.A2(n_1689),
.A3(n_1502),
.B1(n_1497),
.B2(n_1491),
.C1(n_1485),
.C2(n_1483),
.Y(n_1691)
);

AOI221xp5_ASAP7_75t_L g1692 ( 
.A1(n_1691),
.A2(n_1502),
.B1(n_1497),
.B2(n_1485),
.C(n_1483),
.Y(n_1692)
);

AOI211xp5_ASAP7_75t_L g1693 ( 
.A1(n_1692),
.A2(n_1164),
.B(n_1485),
.C(n_1483),
.Y(n_1693)
);


endmodule