module real_jpeg_27627_n_18 (n_17, n_8, n_0, n_2, n_10, n_9, n_298, n_12, n_6, n_11, n_14, n_7, n_3, n_5, n_4, n_1, n_16, n_15, n_13, n_18);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_298;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;

output n_18;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_78;
wire n_83;
wire n_286;
wire n_166;
wire n_176;
wire n_288;
wire n_292;
wire n_215;
wire n_221;
wire n_249;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_280;
wire n_64;
wire n_177;
wire n_291;
wire n_236;
wire n_47;
wire n_131;
wire n_271;
wire n_281;
wire n_163;
wire n_276;
wire n_22;
wire n_287;
wire n_174;
wire n_237;
wire n_87;
wire n_255;
wire n_40;
wire n_105;
wire n_173;
wire n_197;
wire n_243;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_293;
wire n_200;
wire n_275;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_282;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_44;
wire n_28;
wire n_267;
wire n_208;
wire n_62;
wire n_239;
wire n_162;
wire n_290;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_172;
wire n_160;
wire n_211;
wire n_45;
wire n_285;
wire n_112;
wire n_42;
wire n_268;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_222;
wire n_148;
wire n_262;
wire n_118;
wire n_220;
wire n_294;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_198;
wire n_192;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_205;
wire n_258;
wire n_289;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_228;
wire n_150;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_278;
wire n_241;
wire n_103;
wire n_225;
wire n_259;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_284;
wire n_226;
wire n_277;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_230;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_279;
wire n_59;
wire n_169;
wire n_128;
wire n_167;
wire n_213;
wire n_179;
wire n_202;
wire n_244;
wire n_133;
wire n_216;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_210;
wire n_206;
wire n_224;
wire n_119;
wire n_36;
wire n_102;
wire n_81;
wire n_85;
wire n_181;
wire n_283;
wire n_101;
wire n_274;
wire n_256;
wire n_182;
wire n_269;
wire n_96;
wire n_253;
wire n_273;
wire n_89;

OAI22xp5_ASAP7_75t_L g41 ( 
.A1(n_0),
.A2(n_42),
.B1(n_43),
.B2(n_44),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_0),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_L g136 ( 
.A1(n_0),
.A2(n_42),
.B1(n_50),
.B2(n_51),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_SL g176 ( 
.A1(n_0),
.A2(n_42),
.B1(n_63),
.B2(n_64),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_0),
.A2(n_29),
.B1(n_36),
.B2(n_42),
.Y(n_223)
);

HB1xp67_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

INVx11_ASAP7_75t_L g34 ( 
.A(n_1),
.Y(n_34)
);

INVx5_ASAP7_75t_L g239 ( 
.A(n_1),
.Y(n_239)
);

AOI22xp33_ASAP7_75t_L g62 ( 
.A1(n_2),
.A2(n_63),
.B1(n_64),
.B2(n_65),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_2),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_2),
.A2(n_50),
.B1(n_51),
.B2(n_65),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_2),
.A2(n_29),
.B1(n_36),
.B2(n_65),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_3),
.Y(n_145)
);

AOI21xp33_ASAP7_75t_SL g146 ( 
.A1(n_3),
.A2(n_47),
.B(n_51),
.Y(n_146)
);

OAI22xp33_ASAP7_75t_SL g178 ( 
.A1(n_3),
.A2(n_43),
.B1(n_44),
.B2(n_145),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_3),
.B(n_49),
.Y(n_187)
);

AOI21xp5_ASAP7_75t_L g207 ( 
.A1(n_3),
.A2(n_63),
.B(n_208),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_3),
.B(n_63),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_3),
.B(n_95),
.Y(n_217)
);

OAI22xp33_ASAP7_75t_SL g238 ( 
.A1(n_3),
.A2(n_27),
.B1(n_235),
.B2(n_239),
.Y(n_238)
);

AOI21xp5_ASAP7_75t_L g250 ( 
.A1(n_3),
.A2(n_50),
.B(n_251),
.Y(n_250)
);

BUFx12_ASAP7_75t_L g47 ( 
.A(n_4),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_5),
.A2(n_43),
.B1(n_44),
.B2(n_141),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_5),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_L g184 ( 
.A1(n_5),
.A2(n_50),
.B1(n_51),
.B2(n_141),
.Y(n_184)
);

AOI22xp33_ASAP7_75t_SL g209 ( 
.A1(n_5),
.A2(n_63),
.B1(n_64),
.B2(n_141),
.Y(n_209)
);

AOI22xp33_ASAP7_75t_SL g235 ( 
.A1(n_5),
.A2(n_29),
.B1(n_36),
.B2(n_141),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_6),
.A2(n_50),
.B1(n_51),
.B2(n_85),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_6),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_L g100 ( 
.A1(n_6),
.A2(n_63),
.B1(n_64),
.B2(n_85),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_6),
.A2(n_43),
.B1(n_44),
.B2(n_85),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_6),
.A2(n_29),
.B1(n_36),
.B2(n_85),
.Y(n_148)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_7),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g35 ( 
.A1(n_8),
.A2(n_29),
.B1(n_36),
.B2(n_37),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_8),
.Y(n_37)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_8),
.A2(n_37),
.B1(n_63),
.B2(n_64),
.Y(n_88)
);

BUFx10_ASAP7_75t_L g43 ( 
.A(n_9),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_10),
.A2(n_43),
.B1(n_44),
.B2(n_55),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_10),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_10),
.A2(n_50),
.B1(n_51),
.B2(n_55),
.Y(n_93)
);

OAI22xp33_ASAP7_75t_L g130 ( 
.A1(n_10),
.A2(n_55),
.B1(n_63),
.B2(n_64),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_10),
.A2(n_29),
.B1(n_36),
.B2(n_55),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g68 ( 
.A1(n_11),
.A2(n_29),
.B1(n_36),
.B2(n_69),
.Y(n_68)
);

INVx11_ASAP7_75t_L g69 ( 
.A(n_11),
.Y(n_69)
);

OAI22xp33_ASAP7_75t_L g70 ( 
.A1(n_11),
.A2(n_63),
.B1(n_64),
.B2(n_69),
.Y(n_70)
);

OAI32xp33_ASAP7_75t_L g211 ( 
.A1(n_11),
.A2(n_36),
.A3(n_63),
.B1(n_212),
.B2(n_213),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_12),
.A2(n_43),
.B1(n_44),
.B2(n_103),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_12),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g151 ( 
.A1(n_12),
.A2(n_50),
.B1(n_51),
.B2(n_103),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_L g222 ( 
.A1(n_12),
.A2(n_29),
.B1(n_36),
.B2(n_103),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_12),
.A2(n_63),
.B1(n_64),
.B2(n_103),
.Y(n_255)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_13),
.Y(n_52)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_14),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_14),
.B(n_50),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_14),
.A2(n_63),
.B1(n_64),
.B2(n_80),
.Y(n_82)
);

INVx4_ASAP7_75t_L g261 ( 
.A(n_14),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_15),
.A2(n_63),
.B1(n_64),
.B2(n_73),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_15),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_L g98 ( 
.A1(n_15),
.A2(n_29),
.B1(n_36),
.B2(n_73),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_15),
.A2(n_50),
.B1(n_51),
.B2(n_73),
.Y(n_112)
);

INVx11_ASAP7_75t_SL g30 ( 
.A(n_16),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_17),
.A2(n_43),
.B1(n_44),
.B2(n_134),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_17),
.Y(n_134)
);

OAI22xp33_ASAP7_75t_L g172 ( 
.A1(n_17),
.A2(n_50),
.B1(n_51),
.B2(n_134),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_SL g220 ( 
.A1(n_17),
.A2(n_63),
.B1(n_64),
.B2(n_134),
.Y(n_220)
);

AOI22xp33_ASAP7_75t_SL g229 ( 
.A1(n_17),
.A2(n_29),
.B1(n_36),
.B2(n_134),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_119),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_118),
.Y(n_19)
);

INVxp67_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_104),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_22),
.B(n_104),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_76),
.C(n_90),
.Y(n_22)
);

XOR2xp5_ASAP7_75t_L g163 ( 
.A(n_23),
.B(n_76),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_57),
.B1(n_58),
.B2(n_75),
.Y(n_23)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_24),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_26),
.B1(n_38),
.B2(n_39),
.Y(n_24)
);

OAI21xp5_ASAP7_75t_L g117 ( 
.A1(n_25),
.A2(n_39),
.B(n_57),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_25),
.A2(n_26),
.B1(n_59),
.B2(n_60),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_26),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_26),
.B(n_59),
.Y(n_58)
);

AOI21xp5_ASAP7_75t_L g26 ( 
.A1(n_27),
.A2(n_32),
.B(n_35),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_27),
.A2(n_34),
.B1(n_35),
.B2(n_98),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_27),
.A2(n_32),
.B1(n_98),
.B2(n_126),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_27),
.A2(n_222),
.B1(n_223),
.B2(n_224),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_27),
.A2(n_34),
.B1(n_229),
.B2(n_235),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_L g264 ( 
.A1(n_27),
.A2(n_223),
.B1(n_224),
.B2(n_265),
.Y(n_264)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_28),
.A2(n_127),
.B1(n_148),
.B2(n_149),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_28),
.A2(n_33),
.B1(n_148),
.B2(n_186),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_28),
.A2(n_33),
.B1(n_228),
.B2(n_230),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_31),
.Y(n_28)
);

INVx11_ASAP7_75t_L g36 ( 
.A(n_29),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_SL g213 ( 
.A(n_29),
.B(n_69),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_SL g240 ( 
.A(n_29),
.B(n_241),
.Y(n_240)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_32),
.Y(n_149)
);

INVx11_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx5_ASAP7_75t_SL g224 ( 
.A(n_33),
.Y(n_224)
);

INVx11_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_L g39 ( 
.A1(n_40),
.A2(n_45),
.B1(n_54),
.B2(n_56),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_41),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_41),
.A2(n_46),
.B1(n_49),
.B2(n_102),
.Y(n_101)
);

INVx13_ASAP7_75t_L g44 ( 
.A(n_43),
.Y(n_44)
);

A2O1A1Ixp33_ASAP7_75t_L g144 ( 
.A1(n_43),
.A2(n_53),
.B(n_145),
.C(n_146),
.Y(n_144)
);

O2A1O1Ixp33_ASAP7_75t_L g46 ( 
.A1(n_44),
.A2(n_47),
.B(n_48),
.C(n_49),
.Y(n_46)
);

NAND2xp33_ASAP7_75t_SL g48 ( 
.A(n_44),
.B(n_47),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_45),
.A2(n_54),
.B1(n_56),
.B2(n_108),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_45),
.A2(n_56),
.B1(n_139),
.B2(n_142),
.Y(n_138)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_46),
.A2(n_49),
.B1(n_102),
.B2(n_133),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_46),
.A2(n_49),
.B1(n_140),
.B2(n_178),
.Y(n_177)
);

AO22x1_ASAP7_75t_L g49 ( 
.A1(n_47),
.A2(n_50),
.B1(n_51),
.B2(n_53),
.Y(n_49)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_47),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_49),
.Y(n_56)
);

A2O1A1Ixp33_ASAP7_75t_L g78 ( 
.A1(n_50),
.A2(n_79),
.B(n_81),
.C(n_82),
.Y(n_78)
);

OAI32xp33_ASAP7_75t_L g259 ( 
.A1(n_50),
.A2(n_64),
.A3(n_252),
.B1(n_260),
.B2(n_262),
.Y(n_259)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_51),
.B(n_145),
.Y(n_252)
);

INVx11_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g60 ( 
.A1(n_61),
.A2(n_66),
.B1(n_71),
.B2(n_74),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_62),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_62),
.A2(n_67),
.B1(n_68),
.B2(n_100),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_SL g262 ( 
.A(n_63),
.B(n_263),
.Y(n_262)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_66),
.A2(n_74),
.B1(n_130),
.B2(n_175),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_66),
.A2(n_74),
.B1(n_254),
.B2(n_255),
.Y(n_253)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_67),
.A2(n_68),
.B1(n_72),
.B2(n_88),
.Y(n_87)
);

AOI21xp5_ASAP7_75t_L g113 ( 
.A1(n_67),
.A2(n_68),
.B(n_88),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_67),
.A2(n_68),
.B1(n_100),
.B2(n_129),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g206 ( 
.A1(n_67),
.A2(n_68),
.B1(n_207),
.B2(n_209),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_67),
.A2(n_68),
.B1(n_209),
.B2(n_220),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_67),
.A2(n_68),
.B1(n_176),
.B2(n_279),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_68),
.B(n_70),
.Y(n_67)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_68),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g236 ( 
.A(n_68),
.B(n_145),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_72),
.Y(n_71)
);

AOI21xp5_ASAP7_75t_L g76 ( 
.A1(n_77),
.A2(n_87),
.B(n_89),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_77),
.B(n_87),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_78),
.A2(n_82),
.B1(n_83),
.B2(n_86),
.Y(n_77)
);

CKINVDCx16_ASAP7_75t_R g94 ( 
.A(n_78),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_78),
.A2(n_82),
.B1(n_151),
.B2(n_152),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_78),
.A2(n_82),
.B1(n_151),
.B2(n_171),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g249 ( 
.A1(n_78),
.A2(n_82),
.B1(n_184),
.B2(n_250),
.Y(n_249)
);

INVx1_ASAP7_75t_SL g79 ( 
.A(n_80),
.Y(n_79)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_82),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_84),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_84),
.A2(n_93),
.B1(n_94),
.B2(n_95),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_86),
.Y(n_111)
);

FAx1_ASAP7_75t_SL g104 ( 
.A(n_89),
.B(n_105),
.CI(n_117),
.CON(n_104),
.SN(n_104)
);

AOI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_90),
.A2(n_91),
.B1(n_162),
.B2(n_163),
.Y(n_161)
);

CKINVDCx16_ASAP7_75t_R g90 ( 
.A(n_91),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_92),
.B(n_96),
.C(n_101),
.Y(n_91)
);

FAx1_ASAP7_75t_SL g157 ( 
.A(n_92),
.B(n_96),
.CI(n_101),
.CON(n_157),
.SN(n_157)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_93),
.A2(n_94),
.B1(n_95),
.B2(n_136),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_94),
.A2(n_95),
.B1(n_111),
.B2(n_112),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_94),
.A2(n_95),
.B1(n_172),
.B2(n_183),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_99),
.Y(n_96)
);

XNOR2xp5_ASAP7_75t_L g153 ( 
.A(n_97),
.B(n_99),
.Y(n_153)
);

BUFx24_ASAP7_75t_SL g296 ( 
.A(n_104),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_106),
.A2(n_107),
.B1(n_109),
.B2(n_116),
.Y(n_105)
);

CKINVDCx14_ASAP7_75t_R g106 ( 
.A(n_107),
.Y(n_106)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_109),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_L g109 ( 
.A1(n_110),
.A2(n_113),
.B1(n_114),
.B2(n_115),
.Y(n_109)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_110),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_113),
.Y(n_115)
);

AOI321xp33_ASAP7_75t_L g119 ( 
.A1(n_120),
.A2(n_159),
.A3(n_164),
.B1(n_289),
.B2(n_294),
.C(n_298),
.Y(n_119)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_SL g289 ( 
.A1(n_121),
.A2(n_290),
.B(n_293),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_122),
.B(n_154),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g293 ( 
.A(n_122),
.B(n_154),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_123),
.B(n_137),
.C(n_153),
.Y(n_122)
);

XNOR2xp5_ASAP7_75t_L g198 ( 
.A(n_123),
.B(n_153),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_SL g123 ( 
.A(n_124),
.B(n_131),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_124),
.B(n_132),
.C(n_135),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_125),
.B(n_128),
.Y(n_124)
);

XOR2xp5_ASAP7_75t_L g190 ( 
.A(n_125),
.B(n_128),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_127),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_130),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_L g131 ( 
.A(n_132),
.B(n_135),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_133),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_136),
.Y(n_152)
);

XNOR2xp5_ASAP7_75t_L g197 ( 
.A(n_137),
.B(n_198),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_143),
.C(n_150),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_138),
.B(n_150),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_140),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_SL g192 ( 
.A(n_143),
.B(n_193),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_147),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_144),
.B(n_147),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_145),
.B(n_239),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_158),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_157),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_156),
.B(n_157),
.C(n_158),
.Y(n_160)
);

BUFx24_ASAP7_75t_SL g297 ( 
.A(n_157),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_161),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_160),
.B(n_161),
.Y(n_294)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

NOR3xp33_ASAP7_75t_SL g164 ( 
.A(n_165),
.B(n_194),
.C(n_199),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_188),
.Y(n_165)
);

AND2x2_ASAP7_75t_L g291 ( 
.A(n_166),
.B(n_188),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_167),
.B(n_179),
.C(n_180),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g285 ( 
.A(n_167),
.B(n_286),
.Y(n_285)
);

XOR2xp5_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_177),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_169),
.A2(n_170),
.B1(n_173),
.B2(n_174),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_169),
.B(n_174),
.C(n_177),
.Y(n_191)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_172),
.Y(n_171)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_176),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_L g286 ( 
.A1(n_179),
.A2(n_180),
.B1(n_181),
.B2(n_287),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_179),
.Y(n_287)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_182),
.B(n_185),
.C(n_187),
.Y(n_181)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_182),
.B(n_274),
.Y(n_273)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_185),
.B(n_187),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_186),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g188 ( 
.A(n_189),
.B(n_192),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_L g189 ( 
.A(n_190),
.B(n_191),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_190),
.B(n_191),
.C(n_192),
.Y(n_196)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

AOI21xp33_ASAP7_75t_L g290 ( 
.A1(n_195),
.A2(n_291),
.B(n_292),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_197),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_SL g292 ( 
.A(n_196),
.B(n_197),
.Y(n_292)
);

AOI21xp5_ASAP7_75t_L g199 ( 
.A1(n_200),
.A2(n_283),
.B(n_288),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_SL g200 ( 
.A1(n_201),
.A2(n_269),
.B(n_282),
.Y(n_200)
);

AOI21xp5_ASAP7_75t_L g201 ( 
.A1(n_202),
.A2(n_245),
.B(n_268),
.Y(n_201)
);

OAI21xp5_ASAP7_75t_SL g202 ( 
.A1(n_203),
.A2(n_225),
.B(n_244),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_204),
.B(n_214),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g244 ( 
.A(n_204),
.B(n_214),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_SL g204 ( 
.A(n_205),
.B(n_210),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_205),
.A2(n_206),
.B1(n_210),
.B2(n_211),
.Y(n_231)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

CKINVDCx16_ASAP7_75t_R g212 ( 
.A(n_208),
.Y(n_212)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_L g214 ( 
.A(n_215),
.B(n_221),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_216),
.A2(n_217),
.B1(n_218),
.B2(n_219),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_216),
.B(n_219),
.C(n_221),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_217),
.Y(n_216)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_220),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_222),
.Y(n_230)
);

AOI21xp5_ASAP7_75t_L g225 ( 
.A1(n_226),
.A2(n_232),
.B(n_243),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_227),
.B(n_231),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_SL g243 ( 
.A(n_227),
.B(n_231),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_229),
.Y(n_228)
);

OAI21xp5_ASAP7_75t_SL g232 ( 
.A1(n_233),
.A2(n_237),
.B(n_242),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_234),
.B(n_236),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_SL g242 ( 
.A(n_234),
.B(n_236),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_238),
.B(n_240),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_246),
.B(n_247),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_SL g268 ( 
.A(n_246),
.B(n_247),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_248),
.A2(n_258),
.B1(n_266),
.B2(n_267),
.Y(n_247)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_248),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_249),
.A2(n_253),
.B1(n_256),
.B2(n_257),
.Y(n_248)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_249),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_252),
.Y(n_251)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_253),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_253),
.B(n_257),
.C(n_267),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_255),
.Y(n_279)
);

CKINVDCx16_ASAP7_75t_R g267 ( 
.A(n_258),
.Y(n_267)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_259),
.B(n_264),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_259),
.B(n_264),
.Y(n_277)
);

INVx6_ASAP7_75t_L g263 ( 
.A(n_260),
.Y(n_263)
);

INVx8_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_270),
.B(n_271),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_SL g282 ( 
.A(n_270),
.B(n_271),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_272),
.A2(n_273),
.B1(n_275),
.B2(n_276),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_272),
.B(n_278),
.C(n_280),
.Y(n_284)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_277),
.A2(n_278),
.B1(n_280),
.B2(n_281),
.Y(n_276)
);

CKINVDCx16_ASAP7_75t_R g280 ( 
.A(n_277),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_278),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_284),
.B(n_285),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_SL g288 ( 
.A(n_284),
.B(n_285),
.Y(n_288)
);


endmodule