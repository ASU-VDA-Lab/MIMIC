module fake_netlist_6_4959_n_1868 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_161, n_68, n_166, n_28, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_167, n_144, n_127, n_125, n_153, n_168, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_165, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_173, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_171, n_31, n_57, n_169, n_53, n_51, n_44, n_56, n_1868);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_161;
input n_68;
input n_166;
input n_28;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_167;
input n_144;
input n_127;
input n_125;
input n_153;
input n_168;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_165;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_173;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_171;
input n_31;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1868;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_1853;
wire n_783;
wire n_1738;
wire n_798;
wire n_188;
wire n_1575;
wire n_1854;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1691;
wire n_1688;
wire n_1009;
wire n_1743;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_1844;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_1786;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_200;
wire n_447;
wire n_1803;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1867;
wire n_1704;
wire n_1078;
wire n_250;
wire n_544;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_658;
wire n_616;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1842;
wire n_1620;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1798;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_1820;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_1815;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1644;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_577;
wire n_1843;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1762;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1697;
wire n_243;
wire n_979;
wire n_905;
wire n_1866;
wire n_1680;
wire n_175;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1865;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_530;
wire n_1563;
wire n_277;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_1760;
wire n_210;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_178;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_429;
wire n_1747;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1802;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_1801;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_1813;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_1709;
wire n_1825;
wire n_1757;
wire n_1796;
wire n_1792;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_462;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_595;
wire n_627;
wire n_297;
wire n_1767;
wire n_1779;
wire n_524;
wire n_1465;
wire n_342;
wire n_1858;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_1839;
wire n_685;
wire n_1765;
wire n_353;
wire n_605;
wire n_1514;
wire n_1863;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_1808;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_1788;
wire n_622;
wire n_1469;
wire n_1838;
wire n_1835;
wire n_1766;
wire n_1776;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_1771;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_899;
wire n_189;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_1577;
wire n_1181;
wire n_1822;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_1817;
wire n_927;
wire n_1849;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_184;
wire n_552;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_216;
wire n_912;
wire n_1857;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_755;
wire n_931;
wire n_1021;
wire n_527;
wire n_683;
wire n_811;
wire n_474;
wire n_1207;
wire n_312;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_1837;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_211;
wire n_1483;
wire n_1834;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_1787;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1769;
wire n_1220;
wire n_556;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1775;
wire n_1773;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_1745;
wire n_914;
wire n_759;
wire n_1831;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1580;
wire n_1425;
wire n_1281;
wire n_1267;
wire n_1806;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_177;
wire n_1855;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_1832;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1594;
wire n_664;
wire n_1764;
wire n_1429;
wire n_1610;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_186;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_1859;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1852;
wire n_1024;
wire n_1768;
wire n_198;
wire n_1847;
wire n_179;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1841;
wire n_1639;
wire n_1623;
wire n_183;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1818;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1686;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1262;
wire n_218;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1827;
wire n_1361;
wire n_1864;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_370;
wire n_1695;
wire n_1828;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_1823;
wire n_227;
wire n_1720;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_1795;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1845;
wire n_1489;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_1846;
wire n_533;
wire n_806;
wire n_959;
wire n_879;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_1782;
wire n_282;
wire n_1676;
wire n_833;
wire n_1830;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_1086;
wire n_1066;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1484;
wire n_1321;
wire n_1241;
wire n_1672;
wire n_569;
wire n_1758;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1794;
wire n_1236;
wire n_1559;
wire n_1725;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1746;
wire n_1325;
wire n_1002;
wire n_1741;
wire n_545;
wire n_489;
wire n_1804;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1860;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_187;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1800;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_1826;
wire n_566;
wire n_1023;
wire n_1076;
wire n_1118;
wire n_194;
wire n_1007;
wire n_1807;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1814;
wire n_1631;
wire n_591;
wire n_1377;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1824;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_180;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_181;
wire n_1810;
wire n_182;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_1729;
wire n_669;
wire n_176;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1785;
wire n_763;
wire n_1147;
wire n_1848;
wire n_360;
wire n_1754;
wire n_1506;
wire n_1652;
wire n_1812;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_174;
wire n_1173;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1821;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_185;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1525;
wire n_455;
wire n_1585;
wire n_1851;
wire n_363;
wire n_1799;
wire n_1090;
wire n_592;
wire n_1816;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_1829;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_1789;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_271;
wire n_404;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1819;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_1861;
wire n_373;
wire n_1632;
wire n_1805;
wire n_257;
wire n_1557;
wire n_1833;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_1850;
wire n_207;
wire n_1089;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_1836;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_1856;
wire n_1862;
wire n_339;
wire n_784;
wire n_434;
wire n_315;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_1259;
wire n_192;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

INVx1_ASAP7_75t_L g174 ( 
.A(n_16),
.Y(n_174)
);

CKINVDCx16_ASAP7_75t_R g175 ( 
.A(n_74),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_122),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_168),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_108),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_78),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_148),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_62),
.Y(n_181)
);

CKINVDCx16_ASAP7_75t_R g182 ( 
.A(n_130),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_8),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_29),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_50),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_35),
.Y(n_186)
);

BUFx6f_ASAP7_75t_L g187 ( 
.A(n_77),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_32),
.Y(n_188)
);

BUFx8_ASAP7_75t_SL g189 ( 
.A(n_22),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_123),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_56),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_88),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_91),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_112),
.Y(n_194)
);

BUFx10_ASAP7_75t_L g195 ( 
.A(n_65),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_99),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_55),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_142),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_155),
.Y(n_199)
);

BUFx2_ASAP7_75t_L g200 ( 
.A(n_73),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_58),
.Y(n_201)
);

INVx2_ASAP7_75t_SL g202 ( 
.A(n_154),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_21),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_125),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_103),
.Y(n_205)
);

INVxp33_ASAP7_75t_R g206 ( 
.A(n_70),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_63),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_162),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_46),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_61),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_43),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_102),
.Y(n_212)
);

BUFx10_ASAP7_75t_L g213 ( 
.A(n_172),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_65),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_13),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_115),
.Y(n_216)
);

BUFx3_ASAP7_75t_L g217 ( 
.A(n_32),
.Y(n_217)
);

BUFx6f_ASAP7_75t_L g218 ( 
.A(n_76),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_151),
.Y(n_219)
);

BUFx3_ASAP7_75t_L g220 ( 
.A(n_82),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_38),
.Y(n_221)
);

INVx1_ASAP7_75t_SL g222 ( 
.A(n_93),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_48),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_106),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_121),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_48),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_45),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_21),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_43),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_38),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_64),
.Y(n_231)
);

BUFx6f_ASAP7_75t_L g232 ( 
.A(n_57),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_169),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_79),
.Y(n_234)
);

BUFx2_ASAP7_75t_L g235 ( 
.A(n_46),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_33),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_19),
.Y(n_237)
);

HB1xp67_ASAP7_75t_L g238 ( 
.A(n_2),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_13),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_57),
.Y(n_240)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_158),
.Y(n_241)
);

BUFx6f_ASAP7_75t_L g242 ( 
.A(n_161),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_118),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_80),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_66),
.Y(n_245)
);

BUFx6f_ASAP7_75t_L g246 ( 
.A(n_28),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_85),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_146),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_109),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_89),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_72),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_136),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_64),
.Y(n_253)
);

INVx1_ASAP7_75t_SL g254 ( 
.A(n_127),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_105),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_39),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_14),
.Y(n_257)
);

INVx2_ASAP7_75t_SL g258 ( 
.A(n_101),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_92),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_137),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_152),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_3),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_150),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_149),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_8),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_143),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_55),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_11),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_52),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_173),
.Y(n_270)
);

INVx3_ASAP7_75t_L g271 ( 
.A(n_45),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_94),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_14),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_25),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_16),
.Y(n_275)
);

INVx1_ASAP7_75t_SL g276 ( 
.A(n_170),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_166),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_10),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_163),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_12),
.Y(n_280)
);

CKINVDCx16_ASAP7_75t_R g281 ( 
.A(n_128),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_114),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_7),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_51),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_134),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_6),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_36),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_18),
.Y(n_288)
);

BUFx8_ASAP7_75t_SL g289 ( 
.A(n_5),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_54),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_34),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_60),
.Y(n_292)
);

INVx1_ASAP7_75t_SL g293 ( 
.A(n_37),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_31),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_147),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_138),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_20),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_5),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_83),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g300 ( 
.A(n_84),
.Y(n_300)
);

INVx3_ASAP7_75t_L g301 ( 
.A(n_34),
.Y(n_301)
);

INVxp67_ASAP7_75t_L g302 ( 
.A(n_69),
.Y(n_302)
);

INVx2_ASAP7_75t_L g303 ( 
.A(n_11),
.Y(n_303)
);

INVx2_ASAP7_75t_L g304 ( 
.A(n_54),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_59),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_139),
.Y(n_306)
);

BUFx3_ASAP7_75t_L g307 ( 
.A(n_61),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_126),
.Y(n_308)
);

INVx1_ASAP7_75t_SL g309 ( 
.A(n_171),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_10),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_29),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_81),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_87),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_22),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_2),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_86),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_23),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_7),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_124),
.Y(n_319)
);

INVx1_ASAP7_75t_SL g320 ( 
.A(n_52),
.Y(n_320)
);

BUFx3_ASAP7_75t_L g321 ( 
.A(n_30),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_110),
.Y(n_322)
);

INVxp67_ASAP7_75t_L g323 ( 
.A(n_67),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_40),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_159),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_119),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_165),
.Y(n_327)
);

CKINVDCx16_ASAP7_75t_R g328 ( 
.A(n_42),
.Y(n_328)
);

CKINVDCx14_ASAP7_75t_R g329 ( 
.A(n_96),
.Y(n_329)
);

BUFx2_ASAP7_75t_SL g330 ( 
.A(n_9),
.Y(n_330)
);

HB1xp67_ASAP7_75t_L g331 ( 
.A(n_28),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_153),
.Y(n_332)
);

INVx2_ASAP7_75t_L g333 ( 
.A(n_135),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_17),
.Y(n_334)
);

BUFx3_ASAP7_75t_L g335 ( 
.A(n_24),
.Y(n_335)
);

BUFx3_ASAP7_75t_L g336 ( 
.A(n_33),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_95),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_31),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_132),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_140),
.Y(n_340)
);

CKINVDCx16_ASAP7_75t_R g341 ( 
.A(n_59),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_3),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_117),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_40),
.Y(n_344)
);

BUFx2_ASAP7_75t_SL g345 ( 
.A(n_68),
.Y(n_345)
);

CKINVDCx20_ASAP7_75t_R g346 ( 
.A(n_12),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_113),
.Y(n_347)
);

CKINVDCx16_ASAP7_75t_R g348 ( 
.A(n_41),
.Y(n_348)
);

HB1xp67_ASAP7_75t_L g349 ( 
.A(n_24),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_232),
.Y(n_350)
);

INVxp67_ASAP7_75t_L g351 ( 
.A(n_235),
.Y(n_351)
);

INVx2_ASAP7_75t_SL g352 ( 
.A(n_195),
.Y(n_352)
);

CKINVDCx20_ASAP7_75t_R g353 ( 
.A(n_192),
.Y(n_353)
);

HB1xp67_ASAP7_75t_L g354 ( 
.A(n_235),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_189),
.Y(n_355)
);

CKINVDCx20_ASAP7_75t_R g356 ( 
.A(n_205),
.Y(n_356)
);

AND2x2_ASAP7_75t_L g357 ( 
.A(n_217),
.B(n_0),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_232),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_289),
.Y(n_359)
);

INVxp33_ASAP7_75t_L g360 ( 
.A(n_238),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_232),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_232),
.Y(n_362)
);

NOR2xp67_ASAP7_75t_L g363 ( 
.A(n_271),
.B(n_0),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_176),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_177),
.Y(n_365)
);

CKINVDCx20_ASAP7_75t_R g366 ( 
.A(n_248),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_232),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_178),
.Y(n_368)
);

CKINVDCx20_ASAP7_75t_R g369 ( 
.A(n_266),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_232),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_246),
.Y(n_371)
);

INVx2_ASAP7_75t_L g372 ( 
.A(n_242),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_179),
.Y(n_373)
);

INVxp67_ASAP7_75t_SL g374 ( 
.A(n_200),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_180),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_190),
.Y(n_376)
);

INVxp33_ASAP7_75t_SL g377 ( 
.A(n_331),
.Y(n_377)
);

CKINVDCx20_ASAP7_75t_R g378 ( 
.A(n_300),
.Y(n_378)
);

CKINVDCx20_ASAP7_75t_R g379 ( 
.A(n_175),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_246),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_193),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_196),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_246),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_246),
.Y(n_384)
);

NOR2xp67_ASAP7_75t_L g385 ( 
.A(n_271),
.B(n_1),
.Y(n_385)
);

CKINVDCx20_ASAP7_75t_R g386 ( 
.A(n_175),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_198),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_246),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_271),
.Y(n_389)
);

CKINVDCx20_ASAP7_75t_R g390 ( 
.A(n_182),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_271),
.Y(n_391)
);

AND2x2_ASAP7_75t_L g392 ( 
.A(n_217),
.B(n_1),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_301),
.B(n_4),
.Y(n_393)
);

HB1xp67_ASAP7_75t_L g394 ( 
.A(n_328),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_301),
.Y(n_395)
);

INVxp33_ASAP7_75t_SL g396 ( 
.A(n_349),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_301),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_301),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_303),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_303),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_212),
.Y(n_401)
);

BUFx3_ASAP7_75t_L g402 ( 
.A(n_220),
.Y(n_402)
);

INVxp33_ASAP7_75t_SL g403 ( 
.A(n_181),
.Y(n_403)
);

CKINVDCx20_ASAP7_75t_R g404 ( 
.A(n_182),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_304),
.Y(n_405)
);

CKINVDCx20_ASAP7_75t_R g406 ( 
.A(n_281),
.Y(n_406)
);

HB1xp67_ASAP7_75t_L g407 ( 
.A(n_328),
.Y(n_407)
);

CKINVDCx20_ASAP7_75t_R g408 ( 
.A(n_281),
.Y(n_408)
);

INVx2_ASAP7_75t_L g409 ( 
.A(n_242),
.Y(n_409)
);

CKINVDCx20_ASAP7_75t_R g410 ( 
.A(n_329),
.Y(n_410)
);

CKINVDCx20_ASAP7_75t_R g411 ( 
.A(n_216),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_219),
.Y(n_412)
);

HB1xp67_ASAP7_75t_L g413 ( 
.A(n_341),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_304),
.Y(n_414)
);

CKINVDCx20_ASAP7_75t_R g415 ( 
.A(n_224),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_174),
.Y(n_416)
);

NOR2xp33_ASAP7_75t_L g417 ( 
.A(n_200),
.B(n_4),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_L g418 ( 
.A(n_202),
.B(n_6),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_174),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_185),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_225),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_185),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_233),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_186),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_243),
.Y(n_425)
);

BUFx2_ASAP7_75t_SL g426 ( 
.A(n_202),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_186),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_191),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_191),
.Y(n_429)
);

CKINVDCx20_ASAP7_75t_R g430 ( 
.A(n_245),
.Y(n_430)
);

INVxp67_ASAP7_75t_SL g431 ( 
.A(n_220),
.Y(n_431)
);

INVxp33_ASAP7_75t_SL g432 ( 
.A(n_183),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_209),
.Y(n_433)
);

CKINVDCx20_ASAP7_75t_R g434 ( 
.A(n_250),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_209),
.Y(n_435)
);

INVx2_ASAP7_75t_L g436 ( 
.A(n_242),
.Y(n_436)
);

INVxp67_ASAP7_75t_SL g437 ( 
.A(n_214),
.Y(n_437)
);

INVx2_ASAP7_75t_L g438 ( 
.A(n_372),
.Y(n_438)
);

INVx2_ASAP7_75t_L g439 ( 
.A(n_372),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_350),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_L g441 ( 
.A(n_431),
.B(n_258),
.Y(n_441)
);

INVx3_ASAP7_75t_L g442 ( 
.A(n_372),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_371),
.B(n_258),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g444 ( 
.A(n_371),
.B(n_380),
.Y(n_444)
);

HB1xp67_ASAP7_75t_L g445 ( 
.A(n_394),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_L g446 ( 
.A(n_380),
.B(n_252),
.Y(n_446)
);

INVx3_ASAP7_75t_L g447 ( 
.A(n_409),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_SL g448 ( 
.A(n_417),
.B(n_341),
.Y(n_448)
);

AND2x2_ASAP7_75t_L g449 ( 
.A(n_357),
.B(n_307),
.Y(n_449)
);

INVx3_ASAP7_75t_L g450 ( 
.A(n_409),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_350),
.Y(n_451)
);

INVx2_ASAP7_75t_L g452 ( 
.A(n_409),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_358),
.Y(n_453)
);

HB1xp67_ASAP7_75t_L g454 ( 
.A(n_407),
.Y(n_454)
);

BUFx2_ASAP7_75t_L g455 ( 
.A(n_379),
.Y(n_455)
);

BUFx6f_ASAP7_75t_L g456 ( 
.A(n_436),
.Y(n_456)
);

BUFx6f_ASAP7_75t_L g457 ( 
.A(n_436),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_383),
.B(n_259),
.Y(n_458)
);

HB1xp67_ASAP7_75t_L g459 ( 
.A(n_413),
.Y(n_459)
);

AND2x2_ASAP7_75t_L g460 ( 
.A(n_357),
.B(n_307),
.Y(n_460)
);

NOR2x1_ASAP7_75t_L g461 ( 
.A(n_393),
.B(n_241),
.Y(n_461)
);

BUFx8_ASAP7_75t_L g462 ( 
.A(n_392),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_383),
.B(n_260),
.Y(n_463)
);

AND2x2_ASAP7_75t_L g464 ( 
.A(n_392),
.B(n_194),
.Y(n_464)
);

AND2x2_ASAP7_75t_L g465 ( 
.A(n_389),
.B(n_321),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_358),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_361),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_L g468 ( 
.A(n_384),
.B(n_261),
.Y(n_468)
);

INVx3_ASAP7_75t_L g469 ( 
.A(n_436),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_L g470 ( 
.A(n_384),
.B(n_263),
.Y(n_470)
);

AND2x4_ASAP7_75t_L g471 ( 
.A(n_363),
.B(n_385),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_361),
.Y(n_472)
);

BUFx6f_ASAP7_75t_L g473 ( 
.A(n_362),
.Y(n_473)
);

BUFx6f_ASAP7_75t_L g474 ( 
.A(n_362),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_367),
.Y(n_475)
);

NOR2xp33_ASAP7_75t_L g476 ( 
.A(n_426),
.B(n_348),
.Y(n_476)
);

AND2x4_ASAP7_75t_L g477 ( 
.A(n_363),
.B(n_241),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_367),
.Y(n_478)
);

BUFx6f_ASAP7_75t_L g479 ( 
.A(n_370),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_L g480 ( 
.A(n_388),
.B(n_264),
.Y(n_480)
);

INVx2_ASAP7_75t_L g481 ( 
.A(n_370),
.Y(n_481)
);

AND2x4_ASAP7_75t_L g482 ( 
.A(n_385),
.B(n_389),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_L g483 ( 
.A(n_388),
.B(n_270),
.Y(n_483)
);

BUFx6f_ASAP7_75t_L g484 ( 
.A(n_391),
.Y(n_484)
);

INVx5_ASAP7_75t_L g485 ( 
.A(n_402),
.Y(n_485)
);

BUFx6f_ASAP7_75t_L g486 ( 
.A(n_391),
.Y(n_486)
);

INVx2_ASAP7_75t_L g487 ( 
.A(n_395),
.Y(n_487)
);

INVx2_ASAP7_75t_L g488 ( 
.A(n_395),
.Y(n_488)
);

AND2x2_ASAP7_75t_L g489 ( 
.A(n_397),
.B(n_321),
.Y(n_489)
);

INVx3_ASAP7_75t_L g490 ( 
.A(n_397),
.Y(n_490)
);

INVx3_ASAP7_75t_L g491 ( 
.A(n_398),
.Y(n_491)
);

BUFx6f_ASAP7_75t_L g492 ( 
.A(n_398),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_399),
.Y(n_493)
);

OA21x2_ASAP7_75t_L g494 ( 
.A1(n_393),
.A2(n_215),
.B(n_214),
.Y(n_494)
);

INVx2_ASAP7_75t_L g495 ( 
.A(n_399),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_400),
.Y(n_496)
);

INVx6_ASAP7_75t_L g497 ( 
.A(n_402),
.Y(n_497)
);

INVx2_ASAP7_75t_L g498 ( 
.A(n_400),
.Y(n_498)
);

AND2x2_ASAP7_75t_L g499 ( 
.A(n_402),
.B(n_194),
.Y(n_499)
);

CKINVDCx8_ASAP7_75t_R g500 ( 
.A(n_355),
.Y(n_500)
);

INVx2_ASAP7_75t_L g501 ( 
.A(n_405),
.Y(n_501)
);

OR2x2_ASAP7_75t_L g502 ( 
.A(n_418),
.B(n_348),
.Y(n_502)
);

INVx2_ASAP7_75t_L g503 ( 
.A(n_405),
.Y(n_503)
);

INVx2_ASAP7_75t_L g504 ( 
.A(n_414),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_414),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_L g506 ( 
.A(n_426),
.B(n_272),
.Y(n_506)
);

BUFx2_ASAP7_75t_L g507 ( 
.A(n_386),
.Y(n_507)
);

HB1xp67_ASAP7_75t_L g508 ( 
.A(n_354),
.Y(n_508)
);

INVx6_ASAP7_75t_L g509 ( 
.A(n_437),
.Y(n_509)
);

INVx2_ASAP7_75t_L g510 ( 
.A(n_416),
.Y(n_510)
);

BUFx6f_ASAP7_75t_L g511 ( 
.A(n_416),
.Y(n_511)
);

CKINVDCx5p33_ASAP7_75t_R g512 ( 
.A(n_411),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_419),
.Y(n_513)
);

INVx3_ASAP7_75t_L g514 ( 
.A(n_419),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_509),
.B(n_364),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_513),
.Y(n_516)
);

INVx3_ASAP7_75t_L g517 ( 
.A(n_456),
.Y(n_517)
);

AOI22xp5_ASAP7_75t_L g518 ( 
.A1(n_448),
.A2(n_374),
.B1(n_396),
.B2(n_377),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_L g519 ( 
.A(n_509),
.B(n_365),
.Y(n_519)
);

AOI22xp33_ASAP7_75t_L g520 ( 
.A1(n_461),
.A2(n_418),
.B1(n_351),
.B2(n_437),
.Y(n_520)
);

INVx2_ASAP7_75t_L g521 ( 
.A(n_481),
.Y(n_521)
);

INVx2_ASAP7_75t_L g522 ( 
.A(n_481),
.Y(n_522)
);

AND2x6_ASAP7_75t_L g523 ( 
.A(n_461),
.B(n_187),
.Y(n_523)
);

AND2x6_ASAP7_75t_L g524 ( 
.A(n_461),
.B(n_187),
.Y(n_524)
);

INVx3_ASAP7_75t_L g525 ( 
.A(n_456),
.Y(n_525)
);

INVx3_ASAP7_75t_L g526 ( 
.A(n_456),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_513),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_513),
.Y(n_528)
);

BUFx3_ASAP7_75t_L g529 ( 
.A(n_497),
.Y(n_529)
);

OR2x6_ASAP7_75t_L g530 ( 
.A(n_509),
.B(n_345),
.Y(n_530)
);

INVx2_ASAP7_75t_L g531 ( 
.A(n_481),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_L g532 ( 
.A(n_509),
.B(n_471),
.Y(n_532)
);

BUFx3_ASAP7_75t_L g533 ( 
.A(n_497),
.Y(n_533)
);

CKINVDCx5p33_ASAP7_75t_R g534 ( 
.A(n_512),
.Y(n_534)
);

AOI22xp33_ASAP7_75t_L g535 ( 
.A1(n_509),
.A2(n_351),
.B1(n_336),
.B2(n_335),
.Y(n_535)
);

AND2x2_ASAP7_75t_L g536 ( 
.A(n_509),
.B(n_352),
.Y(n_536)
);

NOR2xp33_ASAP7_75t_L g537 ( 
.A(n_509),
.B(n_403),
.Y(n_537)
);

BUFx6f_ASAP7_75t_L g538 ( 
.A(n_511),
.Y(n_538)
);

INVx2_ASAP7_75t_L g539 ( 
.A(n_481),
.Y(n_539)
);

INVx2_ASAP7_75t_L g540 ( 
.A(n_440),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_444),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_SL g542 ( 
.A(n_476),
.B(n_368),
.Y(n_542)
);

INVx8_ASAP7_75t_L g543 ( 
.A(n_471),
.Y(n_543)
);

AND2x2_ASAP7_75t_L g544 ( 
.A(n_499),
.B(n_352),
.Y(n_544)
);

INVx2_ASAP7_75t_L g545 ( 
.A(n_440),
.Y(n_545)
);

NOR2xp33_ASAP7_75t_SL g546 ( 
.A(n_500),
.B(n_359),
.Y(n_546)
);

NOR2xp33_ASAP7_75t_L g547 ( 
.A(n_506),
.B(n_432),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_444),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_440),
.Y(n_549)
);

INVx6_ASAP7_75t_L g550 ( 
.A(n_485),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_451),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_451),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_L g553 ( 
.A(n_471),
.B(n_373),
.Y(n_553)
);

INVx2_ASAP7_75t_L g554 ( 
.A(n_451),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_453),
.Y(n_555)
);

AOI22xp33_ASAP7_75t_L g556 ( 
.A1(n_464),
.A2(n_336),
.B1(n_335),
.B2(n_360),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_SL g557 ( 
.A(n_476),
.B(n_375),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_453),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_453),
.Y(n_559)
);

OAI21xp33_ASAP7_75t_SL g560 ( 
.A1(n_448),
.A2(n_230),
.B(n_215),
.Y(n_560)
);

AOI22xp5_ASAP7_75t_L g561 ( 
.A1(n_502),
.A2(n_227),
.B1(n_211),
.B2(n_310),
.Y(n_561)
);

CKINVDCx5p33_ASAP7_75t_R g562 ( 
.A(n_512),
.Y(n_562)
);

INVx2_ASAP7_75t_L g563 ( 
.A(n_466),
.Y(n_563)
);

INVx4_ASAP7_75t_L g564 ( 
.A(n_485),
.Y(n_564)
);

INVx2_ASAP7_75t_L g565 ( 
.A(n_466),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_466),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_SL g567 ( 
.A(n_506),
.B(n_376),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_467),
.Y(n_568)
);

INVx2_ASAP7_75t_L g569 ( 
.A(n_467),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_467),
.Y(n_570)
);

INVx2_ASAP7_75t_SL g571 ( 
.A(n_471),
.Y(n_571)
);

INVx2_ASAP7_75t_L g572 ( 
.A(n_472),
.Y(n_572)
);

INVx2_ASAP7_75t_L g573 ( 
.A(n_472),
.Y(n_573)
);

NAND3xp33_ASAP7_75t_L g574 ( 
.A(n_494),
.B(n_204),
.C(n_199),
.Y(n_574)
);

INVx2_ASAP7_75t_L g575 ( 
.A(n_472),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_L g576 ( 
.A(n_471),
.B(n_381),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_475),
.Y(n_577)
);

INVx2_ASAP7_75t_L g578 ( 
.A(n_475),
.Y(n_578)
);

CKINVDCx5p33_ASAP7_75t_R g579 ( 
.A(n_500),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_475),
.Y(n_580)
);

INVx2_ASAP7_75t_L g581 ( 
.A(n_438),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_SL g582 ( 
.A(n_502),
.B(n_382),
.Y(n_582)
);

OR2x6_ASAP7_75t_L g583 ( 
.A(n_502),
.B(n_345),
.Y(n_583)
);

AND2x2_ASAP7_75t_L g584 ( 
.A(n_499),
.B(n_420),
.Y(n_584)
);

INVx2_ASAP7_75t_L g585 ( 
.A(n_478),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_478),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_478),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_514),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_SL g589 ( 
.A(n_471),
.B(n_387),
.Y(n_589)
);

CKINVDCx6p67_ASAP7_75t_R g590 ( 
.A(n_455),
.Y(n_590)
);

INVx4_ASAP7_75t_L g591 ( 
.A(n_485),
.Y(n_591)
);

NOR2xp33_ASAP7_75t_L g592 ( 
.A(n_441),
.B(n_401),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_514),
.Y(n_593)
);

INVx3_ASAP7_75t_L g594 ( 
.A(n_456),
.Y(n_594)
);

NOR2xp33_ASAP7_75t_L g595 ( 
.A(n_441),
.B(n_412),
.Y(n_595)
);

INVx2_ASAP7_75t_SL g596 ( 
.A(n_497),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_514),
.Y(n_597)
);

BUFx6f_ASAP7_75t_L g598 ( 
.A(n_511),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_514),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_514),
.Y(n_600)
);

INVx2_ASAP7_75t_L g601 ( 
.A(n_495),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_L g602 ( 
.A(n_446),
.B(n_421),
.Y(n_602)
);

INVx2_ASAP7_75t_L g603 ( 
.A(n_495),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_514),
.Y(n_604)
);

INVx2_ASAP7_75t_L g605 ( 
.A(n_495),
.Y(n_605)
);

INVxp67_ASAP7_75t_L g606 ( 
.A(n_508),
.Y(n_606)
);

INVx3_ASAP7_75t_L g607 ( 
.A(n_456),
.Y(n_607)
);

INVx3_ASAP7_75t_L g608 ( 
.A(n_456),
.Y(n_608)
);

INVx2_ASAP7_75t_SL g609 ( 
.A(n_497),
.Y(n_609)
);

BUFx6f_ASAP7_75t_SL g610 ( 
.A(n_477),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_L g611 ( 
.A(n_446),
.B(n_458),
.Y(n_611)
);

HB1xp67_ASAP7_75t_L g612 ( 
.A(n_445),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_L g613 ( 
.A(n_458),
.B(n_423),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_490),
.Y(n_614)
);

AND2x2_ASAP7_75t_L g615 ( 
.A(n_499),
.B(n_420),
.Y(n_615)
);

INVx4_ASAP7_75t_L g616 ( 
.A(n_485),
.Y(n_616)
);

NAND2xp33_ASAP7_75t_L g617 ( 
.A(n_463),
.B(n_425),
.Y(n_617)
);

AND3x2_ASAP7_75t_L g618 ( 
.A(n_445),
.B(n_323),
.C(n_302),
.Y(n_618)
);

NOR2x1p5_ASAP7_75t_L g619 ( 
.A(n_449),
.B(n_230),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_490),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_490),
.Y(n_621)
);

INVx2_ASAP7_75t_L g622 ( 
.A(n_495),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_L g623 ( 
.A(n_463),
.B(n_222),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_SL g624 ( 
.A(n_462),
.B(n_410),
.Y(n_624)
);

INVx4_ASAP7_75t_L g625 ( 
.A(n_485),
.Y(n_625)
);

BUFx3_ASAP7_75t_L g626 ( 
.A(n_497),
.Y(n_626)
);

BUFx10_ASAP7_75t_L g627 ( 
.A(n_497),
.Y(n_627)
);

BUFx6f_ASAP7_75t_SL g628 ( 
.A(n_477),
.Y(n_628)
);

AOI22xp33_ASAP7_75t_SL g629 ( 
.A1(n_462),
.A2(n_406),
.B1(n_390),
.B2(n_408),
.Y(n_629)
);

NOR2xp33_ASAP7_75t_L g630 ( 
.A(n_468),
.B(n_415),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_490),
.Y(n_631)
);

BUFx4f_ASAP7_75t_L g632 ( 
.A(n_494),
.Y(n_632)
);

INVx2_ASAP7_75t_L g633 ( 
.A(n_498),
.Y(n_633)
);

INVx2_ASAP7_75t_L g634 ( 
.A(n_498),
.Y(n_634)
);

INVx3_ASAP7_75t_L g635 ( 
.A(n_456),
.Y(n_635)
);

INVx3_ASAP7_75t_L g636 ( 
.A(n_456),
.Y(n_636)
);

INVx2_ASAP7_75t_L g637 ( 
.A(n_498),
.Y(n_637)
);

INVx2_ASAP7_75t_L g638 ( 
.A(n_498),
.Y(n_638)
);

INVx2_ASAP7_75t_L g639 ( 
.A(n_501),
.Y(n_639)
);

INVx5_ASAP7_75t_L g640 ( 
.A(n_456),
.Y(n_640)
);

INVx5_ASAP7_75t_L g641 ( 
.A(n_457),
.Y(n_641)
);

NOR2xp33_ASAP7_75t_L g642 ( 
.A(n_468),
.B(n_430),
.Y(n_642)
);

INVx2_ASAP7_75t_L g643 ( 
.A(n_501),
.Y(n_643)
);

INVx2_ASAP7_75t_L g644 ( 
.A(n_501),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_490),
.Y(n_645)
);

INVx2_ASAP7_75t_SL g646 ( 
.A(n_497),
.Y(n_646)
);

OR2x2_ASAP7_75t_L g647 ( 
.A(n_508),
.B(n_454),
.Y(n_647)
);

INVx2_ASAP7_75t_L g648 ( 
.A(n_501),
.Y(n_648)
);

AND2x4_ASAP7_75t_L g649 ( 
.A(n_482),
.B(n_199),
.Y(n_649)
);

NOR2x1p5_ASAP7_75t_L g650 ( 
.A(n_449),
.B(n_231),
.Y(n_650)
);

BUFx3_ASAP7_75t_L g651 ( 
.A(n_494),
.Y(n_651)
);

OAI22xp33_ASAP7_75t_L g652 ( 
.A1(n_454),
.A2(n_293),
.B1(n_320),
.B2(n_228),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_490),
.Y(n_653)
);

INVx2_ASAP7_75t_L g654 ( 
.A(n_503),
.Y(n_654)
);

INVx5_ASAP7_75t_L g655 ( 
.A(n_457),
.Y(n_655)
);

INVx3_ASAP7_75t_L g656 ( 
.A(n_457),
.Y(n_656)
);

AND2x2_ASAP7_75t_L g657 ( 
.A(n_499),
.B(n_422),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_491),
.Y(n_658)
);

BUFx3_ASAP7_75t_L g659 ( 
.A(n_494),
.Y(n_659)
);

INVx4_ASAP7_75t_L g660 ( 
.A(n_485),
.Y(n_660)
);

NOR2xp33_ASAP7_75t_L g661 ( 
.A(n_470),
.B(n_434),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_491),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_SL g663 ( 
.A(n_462),
.B(n_404),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_491),
.Y(n_664)
);

NOR2xp33_ASAP7_75t_L g665 ( 
.A(n_470),
.B(n_353),
.Y(n_665)
);

INVx2_ASAP7_75t_L g666 ( 
.A(n_438),
.Y(n_666)
);

INVx2_ASAP7_75t_L g667 ( 
.A(n_438),
.Y(n_667)
);

INVx2_ASAP7_75t_SL g668 ( 
.A(n_619),
.Y(n_668)
);

INVx2_ASAP7_75t_L g669 ( 
.A(n_516),
.Y(n_669)
);

AND2x4_ASAP7_75t_SL g670 ( 
.A(n_590),
.B(n_612),
.Y(n_670)
);

NAND2xp33_ASAP7_75t_SL g671 ( 
.A(n_579),
.B(n_356),
.Y(n_671)
);

O2A1O1Ixp33_ASAP7_75t_L g672 ( 
.A1(n_541),
.A2(n_443),
.B(n_494),
.C(n_483),
.Y(n_672)
);

BUFx3_ASAP7_75t_L g673 ( 
.A(n_536),
.Y(n_673)
);

INVxp33_ASAP7_75t_SL g674 ( 
.A(n_534),
.Y(n_674)
);

NOR2xp33_ASAP7_75t_L g675 ( 
.A(n_611),
.B(n_459),
.Y(n_675)
);

NOR2xp33_ASAP7_75t_L g676 ( 
.A(n_592),
.B(n_459),
.Y(n_676)
);

NAND2xp33_ASAP7_75t_L g677 ( 
.A(n_523),
.B(n_277),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_L g678 ( 
.A(n_541),
.B(n_462),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_516),
.Y(n_679)
);

AOI22xp5_ASAP7_75t_SL g680 ( 
.A1(n_547),
.A2(n_369),
.B1(n_378),
.B2(n_366),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_527),
.Y(n_681)
);

NOR2xp33_ASAP7_75t_L g682 ( 
.A(n_595),
.B(n_480),
.Y(n_682)
);

INVx2_ASAP7_75t_L g683 ( 
.A(n_527),
.Y(n_683)
);

AND2x6_ASAP7_75t_L g684 ( 
.A(n_651),
.B(n_464),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_528),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_528),
.Y(n_686)
);

A2O1A1Ixp33_ASAP7_75t_L g687 ( 
.A1(n_632),
.A2(n_464),
.B(n_477),
.C(n_482),
.Y(n_687)
);

OR2x2_ASAP7_75t_L g688 ( 
.A(n_647),
.B(n_606),
.Y(n_688)
);

INVx2_ASAP7_75t_L g689 ( 
.A(n_540),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_584),
.Y(n_690)
);

INVx2_ASAP7_75t_L g691 ( 
.A(n_540),
.Y(n_691)
);

INVx2_ASAP7_75t_L g692 ( 
.A(n_545),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_L g693 ( 
.A(n_548),
.B(n_462),
.Y(n_693)
);

OAI21xp5_ASAP7_75t_L g694 ( 
.A1(n_632),
.A2(n_464),
.B(n_494),
.Y(n_694)
);

INVx2_ASAP7_75t_L g695 ( 
.A(n_545),
.Y(n_695)
);

AOI221xp5_ASAP7_75t_L g696 ( 
.A1(n_652),
.A2(n_346),
.B1(n_286),
.B2(n_290),
.C(n_291),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_SL g697 ( 
.A(n_537),
.B(n_462),
.Y(n_697)
);

NAND2xp33_ASAP7_75t_L g698 ( 
.A(n_523),
.B(n_524),
.Y(n_698)
);

AOI22xp33_ASAP7_75t_L g699 ( 
.A1(n_651),
.A2(n_477),
.B1(n_482),
.B2(n_236),
.Y(n_699)
);

INVx3_ASAP7_75t_L g700 ( 
.A(n_610),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_L g701 ( 
.A(n_548),
.B(n_482),
.Y(n_701)
);

INVx2_ASAP7_75t_L g702 ( 
.A(n_554),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_L g703 ( 
.A(n_536),
.B(n_482),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_584),
.Y(n_704)
);

INVxp67_ASAP7_75t_L g705 ( 
.A(n_647),
.Y(n_705)
);

HB1xp67_ASAP7_75t_L g706 ( 
.A(n_583),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_SL g707 ( 
.A(n_632),
.B(n_482),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_L g708 ( 
.A(n_623),
.B(n_477),
.Y(n_708)
);

BUFx5_ASAP7_75t_L g709 ( 
.A(n_651),
.Y(n_709)
);

INVxp67_ASAP7_75t_L g710 ( 
.A(n_582),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_L g711 ( 
.A(n_571),
.B(n_477),
.Y(n_711)
);

INVx2_ASAP7_75t_L g712 ( 
.A(n_554),
.Y(n_712)
);

INVx2_ASAP7_75t_L g713 ( 
.A(n_563),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_615),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_L g715 ( 
.A(n_571),
.B(n_480),
.Y(n_715)
);

NAND3xp33_ASAP7_75t_L g716 ( 
.A(n_520),
.B(n_483),
.C(n_460),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_615),
.Y(n_717)
);

INVxp67_ASAP7_75t_SL g718 ( 
.A(n_532),
.Y(n_718)
);

BUFx6f_ASAP7_75t_L g719 ( 
.A(n_543),
.Y(n_719)
);

INVx2_ASAP7_75t_L g720 ( 
.A(n_563),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_657),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_L g722 ( 
.A(n_515),
.B(n_449),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_657),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_L g724 ( 
.A(n_519),
.B(n_460),
.Y(n_724)
);

INVxp67_ASAP7_75t_L g725 ( 
.A(n_518),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_SL g726 ( 
.A(n_630),
.B(n_500),
.Y(n_726)
);

NOR2xp67_ASAP7_75t_L g727 ( 
.A(n_642),
.B(n_485),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_L g728 ( 
.A(n_602),
.B(n_460),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_549),
.Y(n_729)
);

AOI22xp5_ASAP7_75t_L g730 ( 
.A1(n_661),
.A2(n_309),
.B1(n_254),
.B2(n_276),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_L g731 ( 
.A(n_613),
.B(n_485),
.Y(n_731)
);

NAND3xp33_ASAP7_75t_SL g732 ( 
.A(n_518),
.B(n_507),
.C(n_455),
.Y(n_732)
);

OAI22xp33_ASAP7_75t_L g733 ( 
.A1(n_583),
.A2(n_312),
.B1(n_279),
.B2(n_204),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_L g734 ( 
.A(n_544),
.B(n_485),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_549),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_551),
.Y(n_736)
);

AOI22xp5_ASAP7_75t_L g737 ( 
.A1(n_665),
.A2(n_282),
.B1(n_295),
.B2(n_296),
.Y(n_737)
);

BUFx2_ASAP7_75t_L g738 ( 
.A(n_590),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_SL g739 ( 
.A(n_544),
.B(n_500),
.Y(n_739)
);

INVx8_ASAP7_75t_L g740 ( 
.A(n_583),
.Y(n_740)
);

NOR3xp33_ASAP7_75t_L g741 ( 
.A(n_542),
.B(n_507),
.C(n_455),
.Y(n_741)
);

NOR3xp33_ASAP7_75t_L g742 ( 
.A(n_557),
.B(n_507),
.C(n_489),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_552),
.Y(n_743)
);

AOI22xp33_ASAP7_75t_L g744 ( 
.A1(n_659),
.A2(n_315),
.B1(n_231),
.B2(n_236),
.Y(n_744)
);

INVx2_ASAP7_75t_L g745 ( 
.A(n_565),
.Y(n_745)
);

NOR3xp33_ASAP7_75t_L g746 ( 
.A(n_560),
.B(n_489),
.C(n_465),
.Y(n_746)
);

INVx2_ASAP7_75t_L g747 ( 
.A(n_565),
.Y(n_747)
);

NOR2xp33_ASAP7_75t_L g748 ( 
.A(n_553),
.B(n_206),
.Y(n_748)
);

INVx2_ASAP7_75t_L g749 ( 
.A(n_569),
.Y(n_749)
);

INVx2_ASAP7_75t_L g750 ( 
.A(n_569),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_L g751 ( 
.A(n_576),
.B(n_485),
.Y(n_751)
);

INVx2_ASAP7_75t_L g752 ( 
.A(n_572),
.Y(n_752)
);

AOI22xp5_ASAP7_75t_L g753 ( 
.A1(n_583),
.A2(n_617),
.B1(n_560),
.B2(n_619),
.Y(n_753)
);

NOR2xp33_ASAP7_75t_L g754 ( 
.A(n_567),
.B(n_184),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_SL g755 ( 
.A(n_589),
.B(n_299),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_552),
.Y(n_756)
);

NOR2xp33_ASAP7_75t_L g757 ( 
.A(n_659),
.B(n_649),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_L g758 ( 
.A(n_649),
.B(n_491),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_SL g759 ( 
.A(n_546),
.B(n_306),
.Y(n_759)
);

OAI22xp5_ASAP7_75t_L g760 ( 
.A1(n_530),
.A2(n_333),
.B1(n_208),
.B2(n_251),
.Y(n_760)
);

BUFx6f_ASAP7_75t_SL g761 ( 
.A(n_649),
.Y(n_761)
);

AOI22xp33_ASAP7_75t_L g762 ( 
.A1(n_659),
.A2(n_317),
.B1(n_237),
.B2(n_239),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_555),
.Y(n_763)
);

INVx2_ASAP7_75t_L g764 ( 
.A(n_572),
.Y(n_764)
);

AND2x2_ASAP7_75t_L g765 ( 
.A(n_556),
.B(n_535),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_L g766 ( 
.A(n_649),
.B(n_491),
.Y(n_766)
);

INVx2_ASAP7_75t_L g767 ( 
.A(n_573),
.Y(n_767)
);

INVx8_ASAP7_75t_L g768 ( 
.A(n_610),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_SL g769 ( 
.A(n_629),
.B(n_308),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_555),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_L g771 ( 
.A(n_588),
.B(n_491),
.Y(n_771)
);

NOR2xp33_ASAP7_75t_L g772 ( 
.A(n_558),
.B(n_188),
.Y(n_772)
);

A2O1A1Ixp33_ASAP7_75t_L g773 ( 
.A1(n_574),
.A2(n_333),
.B(n_339),
.C(n_247),
.Y(n_773)
);

INVx3_ASAP7_75t_L g774 ( 
.A(n_610),
.Y(n_774)
);

INVx6_ASAP7_75t_L g775 ( 
.A(n_650),
.Y(n_775)
);

NOR2xp33_ASAP7_75t_L g776 ( 
.A(n_558),
.B(n_197),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_SL g777 ( 
.A(n_624),
.B(n_313),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_L g778 ( 
.A(n_588),
.B(n_511),
.Y(n_778)
);

AND2x6_ASAP7_75t_SL g779 ( 
.A(n_562),
.B(n_237),
.Y(n_779)
);

NOR2xp33_ASAP7_75t_R g780 ( 
.A(n_610),
.B(n_316),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_L g781 ( 
.A(n_593),
.B(n_511),
.Y(n_781)
);

INVxp33_ASAP7_75t_SL g782 ( 
.A(n_561),
.Y(n_782)
);

AND2x2_ASAP7_75t_L g783 ( 
.A(n_650),
.B(n_465),
.Y(n_783)
);

INVx1_ASAP7_75t_L g784 ( 
.A(n_559),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_SL g785 ( 
.A(n_543),
.B(n_319),
.Y(n_785)
);

NOR2xp33_ASAP7_75t_L g786 ( 
.A(n_559),
.B(n_201),
.Y(n_786)
);

BUFx6f_ASAP7_75t_L g787 ( 
.A(n_543),
.Y(n_787)
);

INVx2_ASAP7_75t_L g788 ( 
.A(n_573),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_SL g789 ( 
.A(n_543),
.B(n_322),
.Y(n_789)
);

OAI22xp5_ASAP7_75t_L g790 ( 
.A1(n_530),
.A2(n_249),
.B1(n_208),
.B2(n_234),
.Y(n_790)
);

AOI22xp5_ASAP7_75t_L g791 ( 
.A1(n_628),
.A2(n_332),
.B1(n_325),
.B2(n_326),
.Y(n_791)
);

NAND2xp33_ASAP7_75t_L g792 ( 
.A(n_523),
.B(n_327),
.Y(n_792)
);

NOR2xp33_ASAP7_75t_SL g793 ( 
.A(n_628),
.B(n_213),
.Y(n_793)
);

AOI22xp33_ASAP7_75t_L g794 ( 
.A1(n_574),
.A2(n_317),
.B1(n_292),
.B2(n_239),
.Y(n_794)
);

AOI21xp5_ASAP7_75t_L g795 ( 
.A1(n_530),
.A2(n_443),
.B(n_465),
.Y(n_795)
);

NAND2xp33_ASAP7_75t_L g796 ( 
.A(n_523),
.B(n_340),
.Y(n_796)
);

OAI21xp5_ASAP7_75t_L g797 ( 
.A1(n_593),
.A2(n_488),
.B(n_487),
.Y(n_797)
);

NOR2xp33_ASAP7_75t_L g798 ( 
.A(n_566),
.B(n_203),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_L g799 ( 
.A(n_597),
.B(n_511),
.Y(n_799)
);

OR2x2_ASAP7_75t_L g800 ( 
.A(n_561),
.B(n_489),
.Y(n_800)
);

BUFx3_ASAP7_75t_L g801 ( 
.A(n_543),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_L g802 ( 
.A(n_597),
.B(n_599),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_566),
.Y(n_803)
);

CKINVDCx20_ASAP7_75t_R g804 ( 
.A(n_663),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_SL g805 ( 
.A(n_568),
.B(n_343),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_SL g806 ( 
.A(n_570),
.B(n_213),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_L g807 ( 
.A(n_599),
.B(n_511),
.Y(n_807)
);

NOR2xp67_ASAP7_75t_SL g808 ( 
.A(n_538),
.B(n_187),
.Y(n_808)
);

INVx2_ASAP7_75t_L g809 ( 
.A(n_575),
.Y(n_809)
);

NOR2x1p5_ASAP7_75t_L g810 ( 
.A(n_618),
.B(n_207),
.Y(n_810)
);

AOI22xp33_ASAP7_75t_L g811 ( 
.A1(n_523),
.A2(n_292),
.B1(n_257),
.B2(n_267),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_570),
.Y(n_812)
);

BUFx6f_ASAP7_75t_L g813 ( 
.A(n_529),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_L g814 ( 
.A(n_600),
.B(n_511),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_SL g815 ( 
.A(n_577),
.B(n_213),
.Y(n_815)
);

NOR2xp33_ASAP7_75t_SL g816 ( 
.A(n_628),
.B(n_213),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_L g817 ( 
.A(n_600),
.B(n_511),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_SL g818 ( 
.A(n_577),
.B(n_242),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_580),
.Y(n_819)
);

INVx8_ASAP7_75t_L g820 ( 
.A(n_628),
.Y(n_820)
);

NAND2xp33_ASAP7_75t_L g821 ( 
.A(n_523),
.B(n_187),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_L g822 ( 
.A(n_604),
.B(n_511),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_580),
.Y(n_823)
);

INVx2_ASAP7_75t_L g824 ( 
.A(n_575),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_586),
.Y(n_825)
);

NOR2xp33_ASAP7_75t_L g826 ( 
.A(n_586),
.B(n_210),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_SL g827 ( 
.A(n_604),
.B(n_187),
.Y(n_827)
);

INVx3_ASAP7_75t_L g828 ( 
.A(n_578),
.Y(n_828)
);

NOR2xp33_ASAP7_75t_L g829 ( 
.A(n_587),
.B(n_221),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_SL g830 ( 
.A(n_614),
.B(n_187),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_SL g831 ( 
.A(n_614),
.B(n_218),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_L g832 ( 
.A(n_587),
.B(n_510),
.Y(n_832)
);

BUFx3_ASAP7_75t_L g833 ( 
.A(n_620),
.Y(n_833)
);

NAND2xp33_ASAP7_75t_L g834 ( 
.A(n_523),
.B(n_524),
.Y(n_834)
);

AOI22xp5_ASAP7_75t_L g835 ( 
.A1(n_530),
.A2(n_339),
.B1(n_234),
.B2(n_244),
.Y(n_835)
);

OAI21xp5_ASAP7_75t_L g836 ( 
.A1(n_694),
.A2(n_687),
.B(n_707),
.Y(n_836)
);

AOI21xp5_ASAP7_75t_L g837 ( 
.A1(n_718),
.A2(n_609),
.B(n_596),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_L g838 ( 
.A(n_682),
.B(n_524),
.Y(n_838)
);

OAI21xp5_ASAP7_75t_L g839 ( 
.A1(n_707),
.A2(n_621),
.B(n_620),
.Y(n_839)
);

A2O1A1Ixp33_ASAP7_75t_L g840 ( 
.A1(n_682),
.A2(n_344),
.B(n_334),
.C(n_257),
.Y(n_840)
);

AND2x2_ASAP7_75t_SL g841 ( 
.A(n_744),
.B(n_244),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_L g842 ( 
.A(n_728),
.B(n_524),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_L g843 ( 
.A(n_722),
.B(n_524),
.Y(n_843)
);

AOI21xp5_ASAP7_75t_L g844 ( 
.A1(n_711),
.A2(n_609),
.B(n_596),
.Y(n_844)
);

NOR2xp67_ASAP7_75t_L g845 ( 
.A(n_710),
.B(n_621),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_L g846 ( 
.A(n_724),
.B(n_524),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_L g847 ( 
.A(n_708),
.B(n_524),
.Y(n_847)
);

INVx11_ASAP7_75t_L g848 ( 
.A(n_684),
.Y(n_848)
);

OAI21xp5_ASAP7_75t_L g849 ( 
.A1(n_757),
.A2(n_645),
.B(n_631),
.Y(n_849)
);

AND2x2_ASAP7_75t_L g850 ( 
.A(n_675),
.B(n_195),
.Y(n_850)
);

NAND3xp33_ASAP7_75t_SL g851 ( 
.A(n_696),
.B(n_226),
.C(n_223),
.Y(n_851)
);

AOI21xp5_ASAP7_75t_L g852 ( 
.A1(n_703),
.A2(n_646),
.B(n_533),
.Y(n_852)
);

NOR2x1p5_ASAP7_75t_SL g853 ( 
.A(n_709),
.B(n_631),
.Y(n_853)
);

AOI21xp5_ASAP7_75t_L g854 ( 
.A1(n_715),
.A2(n_646),
.B(n_533),
.Y(n_854)
);

AOI22xp5_ASAP7_75t_L g855 ( 
.A1(n_757),
.A2(n_684),
.B1(n_748),
.B2(n_693),
.Y(n_855)
);

AND2x2_ASAP7_75t_L g856 ( 
.A(n_675),
.B(n_195),
.Y(n_856)
);

AOI21xp5_ASAP7_75t_L g857 ( 
.A1(n_701),
.A2(n_734),
.B(n_698),
.Y(n_857)
);

AND2x2_ASAP7_75t_L g858 ( 
.A(n_676),
.B(n_195),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_SL g859 ( 
.A(n_709),
.B(n_645),
.Y(n_859)
);

INVx1_ASAP7_75t_L g860 ( 
.A(n_669),
.Y(n_860)
);

AOI21xp5_ASAP7_75t_L g861 ( 
.A1(n_834),
.A2(n_533),
.B(n_529),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_L g862 ( 
.A(n_676),
.B(n_653),
.Y(n_862)
);

AOI21xp5_ASAP7_75t_L g863 ( 
.A1(n_751),
.A2(n_626),
.B(n_529),
.Y(n_863)
);

BUFx3_ASAP7_75t_L g864 ( 
.A(n_674),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_L g865 ( 
.A(n_699),
.B(n_653),
.Y(n_865)
);

NOR2xp33_ASAP7_75t_SL g866 ( 
.A(n_738),
.B(n_229),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_L g867 ( 
.A(n_699),
.B(n_658),
.Y(n_867)
);

NOR2xp33_ASAP7_75t_L g868 ( 
.A(n_725),
.B(n_658),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_L g869 ( 
.A(n_765),
.B(n_662),
.Y(n_869)
);

NAND2xp5_ASAP7_75t_L g870 ( 
.A(n_783),
.B(n_662),
.Y(n_870)
);

NOR2xp33_ASAP7_75t_L g871 ( 
.A(n_705),
.B(n_664),
.Y(n_871)
);

AOI21xp5_ASAP7_75t_L g872 ( 
.A1(n_758),
.A2(n_626),
.B(n_627),
.Y(n_872)
);

AOI21x1_ASAP7_75t_L g873 ( 
.A1(n_832),
.A2(n_585),
.B(n_578),
.Y(n_873)
);

NOR2xp33_ASAP7_75t_L g874 ( 
.A(n_726),
.B(n_240),
.Y(n_874)
);

INVx2_ASAP7_75t_L g875 ( 
.A(n_683),
.Y(n_875)
);

A2O1A1Ixp33_ASAP7_75t_L g876 ( 
.A1(n_744),
.A2(n_344),
.B(n_291),
.C(n_290),
.Y(n_876)
);

AND2x4_ASAP7_75t_L g877 ( 
.A(n_690),
.B(n_626),
.Y(n_877)
);

INVx4_ASAP7_75t_L g878 ( 
.A(n_719),
.Y(n_878)
);

AOI22xp5_ASAP7_75t_L g879 ( 
.A1(n_684),
.A2(n_517),
.B1(n_525),
.B2(n_656),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_SL g880 ( 
.A(n_709),
.B(n_538),
.Y(n_880)
);

HB1xp67_ASAP7_75t_L g881 ( 
.A(n_673),
.Y(n_881)
);

NOR2xp33_ASAP7_75t_L g882 ( 
.A(n_688),
.B(n_253),
.Y(n_882)
);

AOI21xp5_ASAP7_75t_L g883 ( 
.A1(n_766),
.A2(n_627),
.B(n_591),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_SL g884 ( 
.A(n_709),
.B(n_538),
.Y(n_884)
);

AND2x4_ASAP7_75t_L g885 ( 
.A(n_704),
.B(n_422),
.Y(n_885)
);

AND2x4_ASAP7_75t_L g886 ( 
.A(n_714),
.B(n_424),
.Y(n_886)
);

OAI21xp33_ASAP7_75t_L g887 ( 
.A1(n_730),
.A2(n_262),
.B(n_256),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_L g888 ( 
.A(n_679),
.B(n_517),
.Y(n_888)
);

NOR2xp33_ASAP7_75t_L g889 ( 
.A(n_748),
.B(n_265),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_L g890 ( 
.A(n_681),
.B(n_517),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_L g891 ( 
.A(n_685),
.B(n_686),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_SL g892 ( 
.A(n_709),
.B(n_538),
.Y(n_892)
);

AOI21x1_ASAP7_75t_L g893 ( 
.A1(n_795),
.A2(n_522),
.B(n_521),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_L g894 ( 
.A(n_729),
.B(n_517),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_L g895 ( 
.A(n_735),
.B(n_525),
.Y(n_895)
);

AOI21xp5_ASAP7_75t_L g896 ( 
.A1(n_731),
.A2(n_627),
.B(n_591),
.Y(n_896)
);

INVx1_ASAP7_75t_L g897 ( 
.A(n_833),
.Y(n_897)
);

AOI21xp5_ASAP7_75t_L g898 ( 
.A1(n_797),
.A2(n_627),
.B(n_591),
.Y(n_898)
);

OAI21xp5_ASAP7_75t_L g899 ( 
.A1(n_672),
.A2(n_603),
.B(n_601),
.Y(n_899)
);

NOR2x1_ASAP7_75t_L g900 ( 
.A(n_678),
.B(n_247),
.Y(n_900)
);

NOR2x1p5_ASAP7_75t_L g901 ( 
.A(n_732),
.B(n_268),
.Y(n_901)
);

AOI21xp5_ASAP7_75t_L g902 ( 
.A1(n_697),
.A2(n_591),
.B(n_564),
.Y(n_902)
);

NOR2x1_ASAP7_75t_R g903 ( 
.A(n_775),
.B(n_330),
.Y(n_903)
);

NOR3xp33_ASAP7_75t_L g904 ( 
.A(n_739),
.B(n_251),
.C(n_249),
.Y(n_904)
);

AND2x2_ASAP7_75t_L g905 ( 
.A(n_717),
.B(n_424),
.Y(n_905)
);

NOR2xp33_ASAP7_75t_L g906 ( 
.A(n_782),
.B(n_273),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_SL g907 ( 
.A(n_709),
.B(n_538),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_L g908 ( 
.A(n_736),
.B(n_525),
.Y(n_908)
);

AOI21xp5_ASAP7_75t_L g909 ( 
.A1(n_821),
.A2(n_616),
.B(n_564),
.Y(n_909)
);

NOR2xp67_ASAP7_75t_SL g910 ( 
.A(n_719),
.B(n_330),
.Y(n_910)
);

NOR2x1_ASAP7_75t_L g911 ( 
.A(n_716),
.B(n_255),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_L g912 ( 
.A(n_743),
.B(n_526),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_L g913 ( 
.A(n_756),
.B(n_526),
.Y(n_913)
);

OAI22xp5_ASAP7_75t_L g914 ( 
.A1(n_762),
.A2(n_312),
.B1(n_347),
.B2(n_337),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_L g915 ( 
.A(n_763),
.B(n_526),
.Y(n_915)
);

AOI21xp5_ASAP7_75t_L g916 ( 
.A1(n_802),
.A2(n_616),
.B(n_564),
.Y(n_916)
);

O2A1O1Ixp5_ASAP7_75t_L g917 ( 
.A1(n_805),
.A2(n_526),
.B(n_594),
.C(n_656),
.Y(n_917)
);

OAI21xp5_ASAP7_75t_L g918 ( 
.A1(n_771),
.A2(n_603),
.B(n_601),
.Y(n_918)
);

NAND2xp5_ASAP7_75t_SL g919 ( 
.A(n_753),
.B(n_538),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_L g920 ( 
.A(n_770),
.B(n_594),
.Y(n_920)
);

O2A1O1Ixp5_ASAP7_75t_L g921 ( 
.A1(n_784),
.A2(n_594),
.B(n_607),
.C(n_608),
.Y(n_921)
);

INVx1_ASAP7_75t_L g922 ( 
.A(n_803),
.Y(n_922)
);

NAND2xp5_ASAP7_75t_SL g923 ( 
.A(n_673),
.B(n_719),
.Y(n_923)
);

BUFx6f_ASAP7_75t_L g924 ( 
.A(n_719),
.Y(n_924)
);

AO21x1_ASAP7_75t_L g925 ( 
.A1(n_733),
.A2(n_279),
.B(n_255),
.Y(n_925)
);

OAI22xp5_ASAP7_75t_L g926 ( 
.A1(n_762),
.A2(n_337),
.B1(n_347),
.B2(n_285),
.Y(n_926)
);

AOI21x1_ASAP7_75t_L g927 ( 
.A1(n_778),
.A2(n_522),
.B(n_521),
.Y(n_927)
);

AOI21xp5_ASAP7_75t_L g928 ( 
.A1(n_813),
.A2(n_616),
.B(n_564),
.Y(n_928)
);

AND2x2_ASAP7_75t_L g929 ( 
.A(n_721),
.B(n_427),
.Y(n_929)
);

NOR2xp33_ASAP7_75t_L g930 ( 
.A(n_800),
.B(n_274),
.Y(n_930)
);

OR2x2_ASAP7_75t_L g931 ( 
.A(n_671),
.B(n_427),
.Y(n_931)
);

AOI21xp5_ASAP7_75t_L g932 ( 
.A1(n_813),
.A2(n_625),
.B(n_616),
.Y(n_932)
);

O2A1O1Ixp33_ASAP7_75t_L g933 ( 
.A1(n_723),
.A2(n_285),
.B(n_639),
.C(n_638),
.Y(n_933)
);

AO21x1_ASAP7_75t_L g934 ( 
.A1(n_760),
.A2(n_269),
.B(n_267),
.Y(n_934)
);

NAND2xp5_ASAP7_75t_L g935 ( 
.A(n_812),
.B(n_594),
.Y(n_935)
);

NAND2xp5_ASAP7_75t_SL g936 ( 
.A(n_787),
.B(n_598),
.Y(n_936)
);

CKINVDCx11_ASAP7_75t_R g937 ( 
.A(n_779),
.Y(n_937)
);

NAND2xp5_ASAP7_75t_L g938 ( 
.A(n_819),
.B(n_607),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_L g939 ( 
.A(n_823),
.B(n_607),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_L g940 ( 
.A(n_825),
.B(n_607),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_L g941 ( 
.A(n_746),
.B(n_608),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_L g942 ( 
.A(n_772),
.B(n_608),
.Y(n_942)
);

INVx2_ASAP7_75t_L g943 ( 
.A(n_689),
.Y(n_943)
);

NAND2xp5_ASAP7_75t_SL g944 ( 
.A(n_787),
.B(n_598),
.Y(n_944)
);

INVx2_ASAP7_75t_L g945 ( 
.A(n_689),
.Y(n_945)
);

NAND2xp5_ASAP7_75t_L g946 ( 
.A(n_772),
.B(n_635),
.Y(n_946)
);

BUFx4f_ASAP7_75t_L g947 ( 
.A(n_670),
.Y(n_947)
);

NOR2xp33_ASAP7_75t_L g948 ( 
.A(n_775),
.B(n_275),
.Y(n_948)
);

OAI22xp5_ASAP7_75t_L g949 ( 
.A1(n_668),
.A2(n_636),
.B1(n_656),
.B2(n_635),
.Y(n_949)
);

A2O1A1Ixp33_ASAP7_75t_L g950 ( 
.A1(n_754),
.A2(n_269),
.B(n_278),
.C(n_283),
.Y(n_950)
);

OAI22x1_ASAP7_75t_L g951 ( 
.A1(n_769),
.A2(n_297),
.B1(n_280),
.B2(n_287),
.Y(n_951)
);

AOI21xp5_ASAP7_75t_L g952 ( 
.A1(n_813),
.A2(n_727),
.B(n_785),
.Y(n_952)
);

NAND3xp33_ASAP7_75t_L g953 ( 
.A(n_754),
.B(n_298),
.C(n_342),
.Y(n_953)
);

OAI21xp5_ASAP7_75t_L g954 ( 
.A1(n_684),
.A2(n_634),
.B(n_637),
.Y(n_954)
);

BUFx2_ASAP7_75t_L g955 ( 
.A(n_804),
.Y(n_955)
);

AOI21xp5_ASAP7_75t_L g956 ( 
.A1(n_813),
.A2(n_625),
.B(n_660),
.Y(n_956)
);

O2A1O1Ixp5_ASAP7_75t_L g957 ( 
.A1(n_776),
.A2(n_636),
.B(n_635),
.C(n_622),
.Y(n_957)
);

OAI21xp5_ASAP7_75t_L g958 ( 
.A1(n_684),
.A2(n_638),
.B(n_605),
.Y(n_958)
);

AOI22xp5_ASAP7_75t_L g959 ( 
.A1(n_775),
.A2(n_742),
.B1(n_761),
.B2(n_706),
.Y(n_959)
);

A2O1A1Ixp33_ASAP7_75t_L g960 ( 
.A1(n_794),
.A2(n_278),
.B(n_283),
.C(n_284),
.Y(n_960)
);

O2A1O1Ixp33_ASAP7_75t_L g961 ( 
.A1(n_773),
.A2(n_633),
.B(n_622),
.C(n_654),
.Y(n_961)
);

INVx2_ASAP7_75t_SL g962 ( 
.A(n_670),
.Y(n_962)
);

AOI21xp5_ASAP7_75t_L g963 ( 
.A1(n_789),
.A2(n_625),
.B(n_660),
.Y(n_963)
);

NAND2xp5_ASAP7_75t_L g964 ( 
.A(n_776),
.B(n_636),
.Y(n_964)
);

O2A1O1Ixp33_ASAP7_75t_L g965 ( 
.A1(n_790),
.A2(n_634),
.B(n_633),
.C(n_654),
.Y(n_965)
);

AOI21xp5_ASAP7_75t_L g966 ( 
.A1(n_677),
.A2(n_796),
.B(n_792),
.Y(n_966)
);

BUFx3_ASAP7_75t_L g967 ( 
.A(n_740),
.Y(n_967)
);

NAND2xp5_ASAP7_75t_L g968 ( 
.A(n_786),
.B(n_636),
.Y(n_968)
);

OAI22xp5_ASAP7_75t_L g969 ( 
.A1(n_801),
.A2(n_637),
.B1(n_605),
.B2(n_648),
.Y(n_969)
);

NOR2xp33_ASAP7_75t_L g970 ( 
.A(n_786),
.B(n_288),
.Y(n_970)
);

AND2x2_ASAP7_75t_L g971 ( 
.A(n_680),
.B(n_428),
.Y(n_971)
);

AOI21xp5_ASAP7_75t_L g972 ( 
.A1(n_781),
.A2(n_625),
.B(n_660),
.Y(n_972)
);

BUFx6f_ASAP7_75t_L g973 ( 
.A(n_787),
.Y(n_973)
);

NAND2xp5_ASAP7_75t_L g974 ( 
.A(n_798),
.B(n_639),
.Y(n_974)
);

OAI321xp33_ASAP7_75t_L g975 ( 
.A1(n_794),
.A2(n_314),
.A3(n_338),
.B1(n_334),
.B2(n_315),
.C(n_284),
.Y(n_975)
);

NAND2xp5_ASAP7_75t_L g976 ( 
.A(n_798),
.B(n_643),
.Y(n_976)
);

NAND2xp5_ASAP7_75t_L g977 ( 
.A(n_826),
.B(n_829),
.Y(n_977)
);

INVx3_ASAP7_75t_L g978 ( 
.A(n_828),
.Y(n_978)
);

INVx1_ASAP7_75t_L g979 ( 
.A(n_691),
.Y(n_979)
);

AND2x2_ASAP7_75t_L g980 ( 
.A(n_826),
.B(n_428),
.Y(n_980)
);

INVx1_ASAP7_75t_L g981 ( 
.A(n_691),
.Y(n_981)
);

INVx2_ASAP7_75t_L g982 ( 
.A(n_692),
.Y(n_982)
);

AOI21xp5_ASAP7_75t_L g983 ( 
.A1(n_799),
.A2(n_660),
.B(n_598),
.Y(n_983)
);

INVx11_ASAP7_75t_L g984 ( 
.A(n_810),
.Y(n_984)
);

NAND3xp33_ASAP7_75t_L g985 ( 
.A(n_737),
.B(n_311),
.C(n_294),
.Y(n_985)
);

INVx1_ASAP7_75t_L g986 ( 
.A(n_692),
.Y(n_986)
);

A2O1A1Ixp33_ASAP7_75t_L g987 ( 
.A1(n_811),
.A2(n_338),
.B(n_314),
.C(n_429),
.Y(n_987)
);

OAI22xp5_ASAP7_75t_L g988 ( 
.A1(n_801),
.A2(n_644),
.B1(n_643),
.B2(n_648),
.Y(n_988)
);

NAND2xp5_ASAP7_75t_L g989 ( 
.A(n_829),
.B(n_828),
.Y(n_989)
);

O2A1O1Ixp33_ASAP7_75t_L g990 ( 
.A1(n_777),
.A2(n_644),
.B(n_539),
.C(n_531),
.Y(n_990)
);

AOI21xp5_ASAP7_75t_L g991 ( 
.A1(n_807),
.A2(n_598),
.B(n_655),
.Y(n_991)
);

OAI21xp5_ASAP7_75t_L g992 ( 
.A1(n_695),
.A2(n_712),
.B(n_702),
.Y(n_992)
);

NOR2xp33_ASAP7_75t_L g993 ( 
.A(n_759),
.B(n_305),
.Y(n_993)
);

NAND2xp5_ASAP7_75t_L g994 ( 
.A(n_695),
.B(n_531),
.Y(n_994)
);

INVx3_ASAP7_75t_L g995 ( 
.A(n_702),
.Y(n_995)
);

NAND2xp5_ASAP7_75t_L g996 ( 
.A(n_712),
.B(n_539),
.Y(n_996)
);

NAND3x1_ASAP7_75t_L g997 ( 
.A(n_741),
.B(n_435),
.C(n_433),
.Y(n_997)
);

INVx3_ASAP7_75t_L g998 ( 
.A(n_713),
.Y(n_998)
);

O2A1O1Ixp33_ASAP7_75t_L g999 ( 
.A1(n_827),
.A2(n_510),
.B(n_487),
.C(n_488),
.Y(n_999)
);

AO21x1_ASAP7_75t_L g1000 ( 
.A1(n_827),
.A2(n_488),
.B(n_487),
.Y(n_1000)
);

HB1xp67_ASAP7_75t_L g1001 ( 
.A(n_761),
.Y(n_1001)
);

OAI21xp5_ASAP7_75t_L g1002 ( 
.A1(n_713),
.A2(n_667),
.B(n_666),
.Y(n_1002)
);

A2O1A1Ixp33_ASAP7_75t_L g1003 ( 
.A1(n_811),
.A2(n_435),
.B(n_429),
.C(n_433),
.Y(n_1003)
);

AOI21xp5_ASAP7_75t_L g1004 ( 
.A1(n_814),
.A2(n_598),
.B(n_655),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_L g1005 ( 
.A(n_720),
.B(n_598),
.Y(n_1005)
);

NAND2xp5_ASAP7_75t_L g1006 ( 
.A(n_720),
.B(n_510),
.Y(n_1006)
);

AOI21xp5_ASAP7_75t_L g1007 ( 
.A1(n_817),
.A2(n_822),
.B(n_787),
.Y(n_1007)
);

AOI21xp5_ASAP7_75t_L g1008 ( 
.A1(n_700),
.A2(n_774),
.B(n_788),
.Y(n_1008)
);

NAND2xp5_ASAP7_75t_L g1009 ( 
.A(n_745),
.B(n_747),
.Y(n_1009)
);

HB1xp67_ASAP7_75t_L g1010 ( 
.A(n_745),
.Y(n_1010)
);

AOI21xp5_ASAP7_75t_L g1011 ( 
.A1(n_700),
.A2(n_655),
.B(n_641),
.Y(n_1011)
);

AOI21xp5_ASAP7_75t_L g1012 ( 
.A1(n_774),
.A2(n_655),
.B(n_641),
.Y(n_1012)
);

OAI21xp33_ASAP7_75t_L g1013 ( 
.A1(n_793),
.A2(n_324),
.B(n_318),
.Y(n_1013)
);

AOI21xp5_ASAP7_75t_L g1014 ( 
.A1(n_747),
.A2(n_655),
.B(n_641),
.Y(n_1014)
);

NAND2xp5_ASAP7_75t_L g1015 ( 
.A(n_749),
.B(n_750),
.Y(n_1015)
);

NOR3xp33_ASAP7_75t_L g1016 ( 
.A(n_755),
.B(n_493),
.C(n_496),
.Y(n_1016)
);

NAND2xp5_ASAP7_75t_L g1017 ( 
.A(n_749),
.B(n_581),
.Y(n_1017)
);

INVx2_ASAP7_75t_L g1018 ( 
.A(n_750),
.Y(n_1018)
);

AOI21xp5_ASAP7_75t_L g1019 ( 
.A1(n_752),
.A2(n_655),
.B(n_641),
.Y(n_1019)
);

NOR2xp33_ASAP7_75t_SL g1020 ( 
.A(n_816),
.B(n_218),
.Y(n_1020)
);

OAI21xp33_ASAP7_75t_L g1021 ( 
.A1(n_806),
.A2(n_493),
.B(n_505),
.Y(n_1021)
);

OAI21xp33_ASAP7_75t_L g1022 ( 
.A1(n_815),
.A2(n_493),
.B(n_505),
.Y(n_1022)
);

OAI21xp33_ASAP7_75t_L g1023 ( 
.A1(n_970),
.A2(n_791),
.B(n_835),
.Y(n_1023)
);

AOI22xp5_ASAP7_75t_L g1024 ( 
.A1(n_970),
.A2(n_740),
.B1(n_768),
.B2(n_820),
.Y(n_1024)
);

NOR2xp33_ASAP7_75t_L g1025 ( 
.A(n_977),
.B(n_740),
.Y(n_1025)
);

AOI21xp5_ASAP7_75t_L g1026 ( 
.A1(n_836),
.A2(n_788),
.B(n_767),
.Y(n_1026)
);

OAI22xp5_ASAP7_75t_SL g1027 ( 
.A1(n_906),
.A2(n_218),
.B1(n_242),
.B2(n_752),
.Y(n_1027)
);

AND2x2_ASAP7_75t_L g1028 ( 
.A(n_850),
.B(n_780),
.Y(n_1028)
);

A2O1A1Ixp33_ASAP7_75t_SL g1029 ( 
.A1(n_889),
.A2(n_808),
.B(n_767),
.C(n_824),
.Y(n_1029)
);

AOI21xp5_ASAP7_75t_L g1030 ( 
.A1(n_966),
.A2(n_809),
.B(n_764),
.Y(n_1030)
);

INVx1_ASAP7_75t_L g1031 ( 
.A(n_1010),
.Y(n_1031)
);

OAI22xp5_ASAP7_75t_L g1032 ( 
.A1(n_855),
.A2(n_820),
.B1(n_768),
.B2(n_831),
.Y(n_1032)
);

CKINVDCx16_ASAP7_75t_R g1033 ( 
.A(n_864),
.Y(n_1033)
);

INVx1_ASAP7_75t_L g1034 ( 
.A(n_1010),
.Y(n_1034)
);

NAND2xp5_ASAP7_75t_SL g1035 ( 
.A(n_980),
.B(n_768),
.Y(n_1035)
);

NOR2xp33_ASAP7_75t_L g1036 ( 
.A(n_906),
.B(n_820),
.Y(n_1036)
);

O2A1O1Ixp33_ASAP7_75t_L g1037 ( 
.A1(n_950),
.A2(n_818),
.B(n_831),
.C(n_830),
.Y(n_1037)
);

NOR2xp33_ASAP7_75t_L g1038 ( 
.A(n_930),
.B(n_830),
.Y(n_1038)
);

O2A1O1Ixp33_ASAP7_75t_L g1039 ( 
.A1(n_950),
.A2(n_487),
.B(n_496),
.C(n_505),
.Y(n_1039)
);

INVxp67_ASAP7_75t_SL g1040 ( 
.A(n_881),
.Y(n_1040)
);

OR2x2_ASAP7_75t_L g1041 ( 
.A(n_955),
.B(n_496),
.Y(n_1041)
);

NAND2xp5_ASAP7_75t_L g1042 ( 
.A(n_868),
.B(n_484),
.Y(n_1042)
);

INVx4_ASAP7_75t_L g1043 ( 
.A(n_924),
.Y(n_1043)
);

NOR2xp33_ASAP7_75t_SL g1044 ( 
.A(n_864),
.B(n_218),
.Y(n_1044)
);

A2O1A1Ixp33_ASAP7_75t_L g1045 ( 
.A1(n_874),
.A2(n_930),
.B(n_993),
.C(n_868),
.Y(n_1045)
);

O2A1O1Ixp33_ASAP7_75t_L g1046 ( 
.A1(n_851),
.A2(n_504),
.B(n_503),
.C(n_581),
.Y(n_1046)
);

NAND2xp5_ASAP7_75t_SL g1047 ( 
.A(n_881),
.B(n_218),
.Y(n_1047)
);

A2O1A1Ixp33_ASAP7_75t_L g1048 ( 
.A1(n_874),
.A2(n_218),
.B(n_503),
.C(n_504),
.Y(n_1048)
);

NAND2xp5_ASAP7_75t_L g1049 ( 
.A(n_862),
.B(n_484),
.Y(n_1049)
);

BUFx6f_ASAP7_75t_L g1050 ( 
.A(n_924),
.Y(n_1050)
);

AND2x2_ASAP7_75t_L g1051 ( 
.A(n_856),
.B(n_882),
.Y(n_1051)
);

NAND2x1_ASAP7_75t_L g1052 ( 
.A(n_878),
.B(n_550),
.Y(n_1052)
);

BUFx6f_ASAP7_75t_L g1053 ( 
.A(n_924),
.Y(n_1053)
);

AOI21xp5_ASAP7_75t_L g1054 ( 
.A1(n_847),
.A2(n_667),
.B(n_666),
.Y(n_1054)
);

INVx2_ASAP7_75t_L g1055 ( 
.A(n_995),
.Y(n_1055)
);

NAND2xp5_ASAP7_75t_SL g1056 ( 
.A(n_845),
.B(n_931),
.Y(n_1056)
);

OAI22xp5_ASAP7_75t_L g1057 ( 
.A1(n_838),
.A2(n_484),
.B1(n_486),
.B2(n_492),
.Y(n_1057)
);

OAI22xp5_ASAP7_75t_SL g1058 ( 
.A1(n_841),
.A2(n_9),
.B1(n_15),
.B2(n_17),
.Y(n_1058)
);

NOR3xp33_ASAP7_75t_L g1059 ( 
.A(n_993),
.B(n_503),
.C(n_504),
.Y(n_1059)
);

O2A1O1Ixp33_ASAP7_75t_L g1060 ( 
.A1(n_840),
.A2(n_504),
.B(n_666),
.C(n_581),
.Y(n_1060)
);

OAI22xp5_ASAP7_75t_L g1061 ( 
.A1(n_865),
.A2(n_486),
.B1(n_484),
.B2(n_492),
.Y(n_1061)
);

BUFx6f_ASAP7_75t_SL g1062 ( 
.A(n_962),
.Y(n_1062)
);

A2O1A1Ixp33_ASAP7_75t_L g1063 ( 
.A1(n_953),
.A2(n_667),
.B(n_486),
.C(n_492),
.Y(n_1063)
);

BUFx6f_ASAP7_75t_L g1064 ( 
.A(n_924),
.Y(n_1064)
);

OAI21xp33_ASAP7_75t_L g1065 ( 
.A1(n_882),
.A2(n_492),
.B(n_486),
.Y(n_1065)
);

INVx3_ASAP7_75t_L g1066 ( 
.A(n_973),
.Y(n_1066)
);

AOI21xp5_ASAP7_75t_L g1067 ( 
.A1(n_857),
.A2(n_641),
.B(n_640),
.Y(n_1067)
);

OAI22xp5_ASAP7_75t_L g1068 ( 
.A1(n_867),
.A2(n_484),
.B1(n_486),
.B2(n_492),
.Y(n_1068)
);

AO22x1_ASAP7_75t_L g1069 ( 
.A1(n_971),
.A2(n_15),
.B1(n_18),
.B2(n_19),
.Y(n_1069)
);

BUFx6f_ASAP7_75t_L g1070 ( 
.A(n_973),
.Y(n_1070)
);

O2A1O1Ixp33_ASAP7_75t_L g1071 ( 
.A1(n_840),
.A2(n_438),
.B(n_439),
.C(n_452),
.Y(n_1071)
);

AOI21xp5_ASAP7_75t_L g1072 ( 
.A1(n_919),
.A2(n_641),
.B(n_640),
.Y(n_1072)
);

INVx3_ASAP7_75t_L g1073 ( 
.A(n_973),
.Y(n_1073)
);

AOI21xp5_ASAP7_75t_L g1074 ( 
.A1(n_919),
.A2(n_946),
.B(n_942),
.Y(n_1074)
);

NAND2xp5_ASAP7_75t_SL g1075 ( 
.A(n_1020),
.B(n_492),
.Y(n_1075)
);

INVx2_ASAP7_75t_SL g1076 ( 
.A(n_901),
.Y(n_1076)
);

INVx1_ASAP7_75t_SL g1077 ( 
.A(n_1001),
.Y(n_1077)
);

AND2x4_ASAP7_75t_L g1078 ( 
.A(n_967),
.B(n_885),
.Y(n_1078)
);

CKINVDCx16_ASAP7_75t_R g1079 ( 
.A(n_866),
.Y(n_1079)
);

OAI21xp5_ASAP7_75t_L g1080 ( 
.A1(n_842),
.A2(n_439),
.B(n_452),
.Y(n_1080)
);

BUFx3_ASAP7_75t_L g1081 ( 
.A(n_947),
.Y(n_1081)
);

OAI21xp33_ASAP7_75t_L g1082 ( 
.A1(n_887),
.A2(n_948),
.B(n_1013),
.Y(n_1082)
);

O2A1O1Ixp33_ASAP7_75t_L g1083 ( 
.A1(n_914),
.A2(n_439),
.B(n_452),
.C(n_447),
.Y(n_1083)
);

NAND2xp5_ASAP7_75t_SL g1084 ( 
.A(n_897),
.B(n_492),
.Y(n_1084)
);

INVx1_ASAP7_75t_L g1085 ( 
.A(n_860),
.Y(n_1085)
);

NAND3xp33_ASAP7_75t_L g1086 ( 
.A(n_985),
.B(n_492),
.C(n_486),
.Y(n_1086)
);

NOR2x1_ASAP7_75t_SL g1087 ( 
.A(n_973),
.B(n_492),
.Y(n_1087)
);

AOI21x1_ASAP7_75t_L g1088 ( 
.A1(n_893),
.A2(n_439),
.B(n_452),
.Y(n_1088)
);

NOR3xp33_ASAP7_75t_SL g1089 ( 
.A(n_948),
.B(n_20),
.C(n_23),
.Y(n_1089)
);

INVx2_ASAP7_75t_SL g1090 ( 
.A(n_947),
.Y(n_1090)
);

AOI21xp5_ASAP7_75t_L g1091 ( 
.A1(n_964),
.A2(n_640),
.B(n_442),
.Y(n_1091)
);

AOI21x1_ASAP7_75t_L g1092 ( 
.A1(n_936),
.A2(n_640),
.B(n_457),
.Y(n_1092)
);

OAI22xp5_ASAP7_75t_L g1093 ( 
.A1(n_989),
.A2(n_486),
.B1(n_484),
.B2(n_550),
.Y(n_1093)
);

BUFx2_ASAP7_75t_L g1094 ( 
.A(n_1001),
.Y(n_1094)
);

AOI21xp5_ASAP7_75t_L g1095 ( 
.A1(n_968),
.A2(n_640),
.B(n_442),
.Y(n_1095)
);

INVx2_ASAP7_75t_SL g1096 ( 
.A(n_885),
.Y(n_1096)
);

AND2x2_ASAP7_75t_L g1097 ( 
.A(n_905),
.B(n_484),
.Y(n_1097)
);

INVx3_ASAP7_75t_L g1098 ( 
.A(n_878),
.Y(n_1098)
);

INVx1_ASAP7_75t_L g1099 ( 
.A(n_875),
.Y(n_1099)
);

NOR2xp67_ASAP7_75t_L g1100 ( 
.A(n_959),
.B(n_107),
.Y(n_1100)
);

NAND2xp5_ASAP7_75t_L g1101 ( 
.A(n_841),
.B(n_486),
.Y(n_1101)
);

AO22x1_ASAP7_75t_L g1102 ( 
.A1(n_904),
.A2(n_25),
.B1(n_26),
.B2(n_27),
.Y(n_1102)
);

NAND2x1p5_ASAP7_75t_L g1103 ( 
.A(n_967),
.B(n_640),
.Y(n_1103)
);

AOI21xp5_ASAP7_75t_L g1104 ( 
.A1(n_1007),
.A2(n_442),
.B(n_447),
.Y(n_1104)
);

AOI21xp5_ASAP7_75t_L g1105 ( 
.A1(n_843),
.A2(n_442),
.B(n_447),
.Y(n_1105)
);

O2A1O1Ixp33_ASAP7_75t_L g1106 ( 
.A1(n_926),
.A2(n_442),
.B(n_447),
.C(n_450),
.Y(n_1106)
);

INVx1_ASAP7_75t_L g1107 ( 
.A(n_922),
.Y(n_1107)
);

OAI22xp5_ASAP7_75t_L g1108 ( 
.A1(n_848),
.A2(n_486),
.B1(n_484),
.B2(n_550),
.Y(n_1108)
);

OR2x2_ASAP7_75t_L g1109 ( 
.A(n_886),
.B(n_484),
.Y(n_1109)
);

NAND2xp5_ASAP7_75t_L g1110 ( 
.A(n_871),
.B(n_447),
.Y(n_1110)
);

O2A1O1Ixp5_ASAP7_75t_L g1111 ( 
.A1(n_899),
.A2(n_447),
.B(n_469),
.C(n_450),
.Y(n_1111)
);

A2O1A1Ixp33_ASAP7_75t_SL g1112 ( 
.A1(n_910),
.A2(n_450),
.B(n_469),
.C(n_98),
.Y(n_1112)
);

NAND2xp5_ASAP7_75t_L g1113 ( 
.A(n_871),
.B(n_450),
.Y(n_1113)
);

AOI21xp5_ASAP7_75t_L g1114 ( 
.A1(n_846),
.A2(n_469),
.B(n_450),
.Y(n_1114)
);

AOI22xp33_ASAP7_75t_L g1115 ( 
.A1(n_911),
.A2(n_479),
.B1(n_474),
.B2(n_473),
.Y(n_1115)
);

A2O1A1Ixp33_ASAP7_75t_L g1116 ( 
.A1(n_1021),
.A2(n_469),
.B(n_457),
.C(n_473),
.Y(n_1116)
);

O2A1O1Ixp33_ASAP7_75t_L g1117 ( 
.A1(n_891),
.A2(n_469),
.B(n_30),
.C(n_35),
.Y(n_1117)
);

BUFx2_ASAP7_75t_L g1118 ( 
.A(n_903),
.Y(n_1118)
);

INVx1_ASAP7_75t_L g1119 ( 
.A(n_979),
.Y(n_1119)
);

BUFx12f_ASAP7_75t_L g1120 ( 
.A(n_937),
.Y(n_1120)
);

NAND2xp5_ASAP7_75t_L g1121 ( 
.A(n_869),
.B(n_473),
.Y(n_1121)
);

NOR2xp33_ASAP7_75t_L g1122 ( 
.A(n_870),
.B(n_27),
.Y(n_1122)
);

NAND2xp5_ASAP7_75t_L g1123 ( 
.A(n_929),
.B(n_473),
.Y(n_1123)
);

INVx2_ASAP7_75t_L g1124 ( 
.A(n_998),
.Y(n_1124)
);

OAI22xp5_ASAP7_75t_L g1125 ( 
.A1(n_974),
.A2(n_550),
.B1(n_457),
.B2(n_474),
.Y(n_1125)
);

NAND2xp5_ASAP7_75t_L g1126 ( 
.A(n_976),
.B(n_479),
.Y(n_1126)
);

OAI22xp5_ASAP7_75t_L g1127 ( 
.A1(n_941),
.A2(n_457),
.B1(n_474),
.B2(n_473),
.Y(n_1127)
);

INVx1_ASAP7_75t_L g1128 ( 
.A(n_981),
.Y(n_1128)
);

NAND2xp5_ASAP7_75t_L g1129 ( 
.A(n_877),
.B(n_479),
.Y(n_1129)
);

O2A1O1Ixp33_ASAP7_75t_L g1130 ( 
.A1(n_876),
.A2(n_36),
.B(n_37),
.C(n_39),
.Y(n_1130)
);

BUFx6f_ASAP7_75t_L g1131 ( 
.A(n_877),
.Y(n_1131)
);

O2A1O1Ixp33_ASAP7_75t_L g1132 ( 
.A1(n_960),
.A2(n_41),
.B(n_42),
.C(n_44),
.Y(n_1132)
);

INVx1_ASAP7_75t_L g1133 ( 
.A(n_986),
.Y(n_1133)
);

HB1xp67_ASAP7_75t_L g1134 ( 
.A(n_978),
.Y(n_1134)
);

NAND2xp5_ASAP7_75t_L g1135 ( 
.A(n_978),
.B(n_943),
.Y(n_1135)
);

O2A1O1Ixp33_ASAP7_75t_L g1136 ( 
.A1(n_960),
.A2(n_44),
.B(n_47),
.C(n_49),
.Y(n_1136)
);

HB1xp67_ASAP7_75t_L g1137 ( 
.A(n_951),
.Y(n_1137)
);

NOR2xp33_ASAP7_75t_L g1138 ( 
.A(n_1022),
.B(n_47),
.Y(n_1138)
);

NOR2xp33_ASAP7_75t_L g1139 ( 
.A(n_923),
.B(n_49),
.Y(n_1139)
);

NAND2xp5_ASAP7_75t_SL g1140 ( 
.A(n_900),
.B(n_975),
.Y(n_1140)
);

NAND2xp5_ASAP7_75t_L g1141 ( 
.A(n_943),
.B(n_479),
.Y(n_1141)
);

INVx1_ASAP7_75t_L g1142 ( 
.A(n_1018),
.Y(n_1142)
);

INVx2_ASAP7_75t_L g1143 ( 
.A(n_998),
.Y(n_1143)
);

NAND2xp5_ASAP7_75t_L g1144 ( 
.A(n_1018),
.B(n_479),
.Y(n_1144)
);

AND2x2_ASAP7_75t_L g1145 ( 
.A(n_945),
.B(n_982),
.Y(n_1145)
);

OAI22xp5_ASAP7_75t_SL g1146 ( 
.A1(n_984),
.A2(n_50),
.B1(n_51),
.B2(n_53),
.Y(n_1146)
);

NAND2xp5_ASAP7_75t_SL g1147 ( 
.A(n_923),
.B(n_479),
.Y(n_1147)
);

O2A1O1Ixp33_ASAP7_75t_SL g1148 ( 
.A1(n_936),
.A2(n_944),
.B(n_987),
.C(n_859),
.Y(n_1148)
);

O2A1O1Ixp33_ASAP7_75t_L g1149 ( 
.A1(n_949),
.A2(n_53),
.B(n_56),
.C(n_58),
.Y(n_1149)
);

AOI22xp33_ASAP7_75t_L g1150 ( 
.A1(n_1016),
.A2(n_479),
.B1(n_474),
.B2(n_473),
.Y(n_1150)
);

NAND2xp5_ASAP7_75t_SL g1151 ( 
.A(n_849),
.B(n_879),
.Y(n_1151)
);

AOI22x1_ASAP7_75t_L g1152 ( 
.A1(n_1008),
.A2(n_457),
.B1(n_474),
.B2(n_473),
.Y(n_1152)
);

INVx4_ASAP7_75t_L g1153 ( 
.A(n_853),
.Y(n_1153)
);

BUFx2_ASAP7_75t_L g1154 ( 
.A(n_997),
.Y(n_1154)
);

NOR2xp33_ASAP7_75t_L g1155 ( 
.A(n_859),
.B(n_60),
.Y(n_1155)
);

NAND2xp5_ASAP7_75t_L g1156 ( 
.A(n_1009),
.B(n_479),
.Y(n_1156)
);

A2O1A1Ixp33_ASAP7_75t_L g1157 ( 
.A1(n_839),
.A2(n_457),
.B(n_474),
.C(n_473),
.Y(n_1157)
);

NAND2x1p5_ASAP7_75t_L g1158 ( 
.A(n_944),
.B(n_479),
.Y(n_1158)
);

AOI21xp5_ASAP7_75t_L g1159 ( 
.A1(n_952),
.A2(n_474),
.B(n_131),
.Y(n_1159)
);

OAI21x1_ASAP7_75t_SL g1160 ( 
.A1(n_934),
.A2(n_129),
.B(n_167),
.Y(n_1160)
);

AOI21xp5_ASAP7_75t_L g1161 ( 
.A1(n_852),
.A2(n_474),
.B(n_120),
.Y(n_1161)
);

BUFx2_ASAP7_75t_L g1162 ( 
.A(n_925),
.Y(n_1162)
);

NOR2xp33_ASAP7_75t_L g1163 ( 
.A(n_880),
.B(n_71),
.Y(n_1163)
);

NOR2xp33_ASAP7_75t_L g1164 ( 
.A(n_880),
.B(n_75),
.Y(n_1164)
);

AOI22xp33_ASAP7_75t_L g1165 ( 
.A1(n_888),
.A2(n_474),
.B1(n_90),
.B2(n_97),
.Y(n_1165)
);

OAI22x1_ASAP7_75t_L g1166 ( 
.A1(n_884),
.A2(n_100),
.B1(n_104),
.B2(n_111),
.Y(n_1166)
);

AOI21xp5_ASAP7_75t_L g1167 ( 
.A1(n_898),
.A2(n_116),
.B(n_133),
.Y(n_1167)
);

AOI21xp5_ASAP7_75t_L g1168 ( 
.A1(n_854),
.A2(n_141),
.B(n_144),
.Y(n_1168)
);

INVx2_ASAP7_75t_L g1169 ( 
.A(n_1015),
.Y(n_1169)
);

NAND2xp5_ASAP7_75t_SL g1170 ( 
.A(n_954),
.B(n_145),
.Y(n_1170)
);

CKINVDCx5p33_ASAP7_75t_R g1171 ( 
.A(n_890),
.Y(n_1171)
);

BUFx8_ASAP7_75t_L g1172 ( 
.A(n_1003),
.Y(n_1172)
);

OR2x2_ASAP7_75t_L g1173 ( 
.A(n_1041),
.B(n_1031),
.Y(n_1173)
);

O2A1O1Ixp33_ASAP7_75t_L g1174 ( 
.A1(n_1045),
.A2(n_933),
.B(n_1003),
.C(n_988),
.Y(n_1174)
);

OA21x2_ASAP7_75t_L g1175 ( 
.A1(n_1074),
.A2(n_957),
.B(n_921),
.Y(n_1175)
);

NOR2xp67_ASAP7_75t_L g1176 ( 
.A(n_1090),
.B(n_908),
.Y(n_1176)
);

INVxp67_ASAP7_75t_L g1177 ( 
.A(n_1094),
.Y(n_1177)
);

BUFx2_ASAP7_75t_L g1178 ( 
.A(n_1033),
.Y(n_1178)
);

AOI22xp5_ASAP7_75t_L g1179 ( 
.A1(n_1051),
.A2(n_907),
.B1(n_892),
.B2(n_884),
.Y(n_1179)
);

O2A1O1Ixp33_ASAP7_75t_L g1180 ( 
.A1(n_1023),
.A2(n_969),
.B(n_990),
.C(n_920),
.Y(n_1180)
);

NAND2x1p5_ASAP7_75t_L g1181 ( 
.A(n_1098),
.B(n_892),
.Y(n_1181)
);

BUFx3_ASAP7_75t_L g1182 ( 
.A(n_1081),
.Y(n_1182)
);

NAND3xp33_ASAP7_75t_L g1183 ( 
.A(n_1089),
.B(n_917),
.C(n_844),
.Y(n_1183)
);

AO31x2_ASAP7_75t_L g1184 ( 
.A1(n_1157),
.A2(n_1000),
.A3(n_863),
.B(n_1004),
.Y(n_1184)
);

O2A1O1Ixp33_ASAP7_75t_SL g1185 ( 
.A1(n_1140),
.A2(n_907),
.B(n_895),
.C(n_938),
.Y(n_1185)
);

AO31x2_ASAP7_75t_L g1186 ( 
.A1(n_1074),
.A2(n_991),
.A3(n_939),
.B(n_935),
.Y(n_1186)
);

A2O1A1Ixp33_ASAP7_75t_L g1187 ( 
.A1(n_1038),
.A2(n_965),
.B(n_837),
.C(n_961),
.Y(n_1187)
);

INVx5_ASAP7_75t_L g1188 ( 
.A(n_1050),
.Y(n_1188)
);

NAND2xp5_ASAP7_75t_L g1189 ( 
.A(n_1171),
.B(n_913),
.Y(n_1189)
);

OAI21x1_ASAP7_75t_L g1190 ( 
.A1(n_1088),
.A2(n_927),
.B(n_873),
.Y(n_1190)
);

AO31x2_ASAP7_75t_L g1191 ( 
.A1(n_1048),
.A2(n_940),
.A3(n_915),
.B(n_912),
.Y(n_1191)
);

CKINVDCx5p33_ASAP7_75t_R g1192 ( 
.A(n_1079),
.Y(n_1192)
);

AOI21xp5_ASAP7_75t_L g1193 ( 
.A1(n_1151),
.A2(n_1030),
.B(n_1025),
.Y(n_1193)
);

BUFx2_ASAP7_75t_L g1194 ( 
.A(n_1040),
.Y(n_1194)
);

CKINVDCx20_ASAP7_75t_R g1195 ( 
.A(n_1120),
.Y(n_1195)
);

INVx3_ASAP7_75t_SL g1196 ( 
.A(n_1076),
.Y(n_1196)
);

INVx1_ASAP7_75t_L g1197 ( 
.A(n_1142),
.Y(n_1197)
);

BUFx3_ASAP7_75t_L g1198 ( 
.A(n_1077),
.Y(n_1198)
);

AND2x4_ASAP7_75t_L g1199 ( 
.A(n_1078),
.B(n_1096),
.Y(n_1199)
);

HB1xp67_ASAP7_75t_L g1200 ( 
.A(n_1034),
.Y(n_1200)
);

AO32x2_ASAP7_75t_L g1201 ( 
.A1(n_1058),
.A2(n_992),
.A3(n_918),
.B1(n_1006),
.B2(n_958),
.Y(n_1201)
);

AO32x2_ASAP7_75t_L g1202 ( 
.A1(n_1027),
.A2(n_1032),
.A3(n_1068),
.B1(n_1061),
.B2(n_1127),
.Y(n_1202)
);

INVx1_ASAP7_75t_L g1203 ( 
.A(n_1107),
.Y(n_1203)
);

A2O1A1Ixp33_ASAP7_75t_L g1204 ( 
.A1(n_1082),
.A2(n_861),
.B(n_872),
.C(n_894),
.Y(n_1204)
);

AOI22xp5_ASAP7_75t_L g1205 ( 
.A1(n_1028),
.A2(n_1005),
.B1(n_996),
.B2(n_994),
.Y(n_1205)
);

INVx2_ASAP7_75t_SL g1206 ( 
.A(n_1078),
.Y(n_1206)
);

AO32x2_ASAP7_75t_L g1207 ( 
.A1(n_1153),
.A2(n_999),
.A3(n_1002),
.B1(n_1017),
.B2(n_1019),
.Y(n_1207)
);

BUFx6f_ASAP7_75t_L g1208 ( 
.A(n_1050),
.Y(n_1208)
);

OAI21x1_ASAP7_75t_L g1209 ( 
.A1(n_1030),
.A2(n_1067),
.B(n_1026),
.Y(n_1209)
);

INVx2_ASAP7_75t_L g1210 ( 
.A(n_1145),
.Y(n_1210)
);

AO31x2_ASAP7_75t_L g1211 ( 
.A1(n_1063),
.A2(n_1014),
.A3(n_902),
.B(n_983),
.Y(n_1211)
);

AOI22xp5_ASAP7_75t_L g1212 ( 
.A1(n_1036),
.A2(n_883),
.B1(n_916),
.B2(n_963),
.Y(n_1212)
);

INVx4_ASAP7_75t_L g1213 ( 
.A(n_1050),
.Y(n_1213)
);

A2O1A1Ixp33_ASAP7_75t_L g1214 ( 
.A1(n_1122),
.A2(n_896),
.B(n_972),
.C(n_1011),
.Y(n_1214)
);

AOI22xp5_ASAP7_75t_L g1215 ( 
.A1(n_1100),
.A2(n_909),
.B1(n_956),
.B2(n_932),
.Y(n_1215)
);

AND2x4_ASAP7_75t_L g1216 ( 
.A(n_1131),
.B(n_1012),
.Y(n_1216)
);

NAND3xp33_ASAP7_75t_SL g1217 ( 
.A(n_1154),
.B(n_928),
.C(n_157),
.Y(n_1217)
);

O2A1O1Ixp33_ASAP7_75t_L g1218 ( 
.A1(n_1137),
.A2(n_156),
.B(n_160),
.C(n_164),
.Y(n_1218)
);

A2O1A1Ixp33_ASAP7_75t_L g1219 ( 
.A1(n_1155),
.A2(n_1138),
.B(n_1164),
.C(n_1163),
.Y(n_1219)
);

HB1xp67_ASAP7_75t_L g1220 ( 
.A(n_1134),
.Y(n_1220)
);

NAND2xp5_ASAP7_75t_L g1221 ( 
.A(n_1169),
.B(n_1056),
.Y(n_1221)
);

BUFx2_ASAP7_75t_L g1222 ( 
.A(n_1131),
.Y(n_1222)
);

NAND2xp5_ASAP7_75t_L g1223 ( 
.A(n_1131),
.B(n_1139),
.Y(n_1223)
);

NAND2xp5_ASAP7_75t_L g1224 ( 
.A(n_1097),
.B(n_1085),
.Y(n_1224)
);

OAI21x1_ASAP7_75t_L g1225 ( 
.A1(n_1067),
.A2(n_1054),
.B(n_1092),
.Y(n_1225)
);

A2O1A1Ixp33_ASAP7_75t_L g1226 ( 
.A1(n_1065),
.A2(n_1149),
.B(n_1167),
.C(n_1037),
.Y(n_1226)
);

A2O1A1Ixp33_ASAP7_75t_L g1227 ( 
.A1(n_1167),
.A2(n_1037),
.B(n_1170),
.C(n_1086),
.Y(n_1227)
);

NOR2xp33_ASAP7_75t_L g1228 ( 
.A(n_1118),
.B(n_1044),
.Y(n_1228)
);

INVx1_ASAP7_75t_L g1229 ( 
.A(n_1135),
.Y(n_1229)
);

AOI21xp5_ASAP7_75t_L g1230 ( 
.A1(n_1049),
.A2(n_1126),
.B(n_1121),
.Y(n_1230)
);

NAND2xp5_ASAP7_75t_L g1231 ( 
.A(n_1099),
.B(n_1119),
.Y(n_1231)
);

AOI21xp5_ASAP7_75t_L g1232 ( 
.A1(n_1042),
.A2(n_1148),
.B(n_1123),
.Y(n_1232)
);

AND2x4_ASAP7_75t_L g1233 ( 
.A(n_1035),
.B(n_1098),
.Y(n_1233)
);

AOI21xp5_ASAP7_75t_SL g1234 ( 
.A1(n_1024),
.A2(n_1087),
.B(n_1101),
.Y(n_1234)
);

AOI21xp5_ASAP7_75t_L g1235 ( 
.A1(n_1159),
.A2(n_1029),
.B(n_1156),
.Y(n_1235)
);

O2A1O1Ixp33_ASAP7_75t_SL g1236 ( 
.A1(n_1112),
.A2(n_1147),
.B(n_1047),
.C(n_1075),
.Y(n_1236)
);

OR2x2_ASAP7_75t_L g1237 ( 
.A(n_1109),
.B(n_1128),
.Y(n_1237)
);

OAI21x1_ASAP7_75t_L g1238 ( 
.A1(n_1054),
.A2(n_1104),
.B(n_1072),
.Y(n_1238)
);

O2A1O1Ixp33_ASAP7_75t_SL g1239 ( 
.A1(n_1132),
.A2(n_1136),
.B(n_1129),
.C(n_1130),
.Y(n_1239)
);

AOI21xp5_ASAP7_75t_L g1240 ( 
.A1(n_1159),
.A2(n_1161),
.B(n_1110),
.Y(n_1240)
);

AOI21xp5_ASAP7_75t_L g1241 ( 
.A1(n_1113),
.A2(n_1080),
.B(n_1072),
.Y(n_1241)
);

HB1xp67_ASAP7_75t_L g1242 ( 
.A(n_1053),
.Y(n_1242)
);

NOR2x1_ASAP7_75t_SL g1243 ( 
.A(n_1053),
.B(n_1070),
.Y(n_1243)
);

CKINVDCx5p33_ASAP7_75t_R g1244 ( 
.A(n_1062),
.Y(n_1244)
);

O2A1O1Ixp33_ASAP7_75t_SL g1245 ( 
.A1(n_1132),
.A2(n_1136),
.B(n_1116),
.C(n_1084),
.Y(n_1245)
);

NOR2xp33_ASAP7_75t_L g1246 ( 
.A(n_1055),
.B(n_1143),
.Y(n_1246)
);

OA21x2_ASAP7_75t_L g1247 ( 
.A1(n_1091),
.A2(n_1095),
.B(n_1111),
.Y(n_1247)
);

NAND2xp5_ASAP7_75t_L g1248 ( 
.A(n_1133),
.B(n_1162),
.Y(n_1248)
);

NOR2xp33_ASAP7_75t_L g1249 ( 
.A(n_1124),
.B(n_1153),
.Y(n_1249)
);

CKINVDCx5p33_ASAP7_75t_R g1250 ( 
.A(n_1062),
.Y(n_1250)
);

AND2x2_ASAP7_75t_L g1251 ( 
.A(n_1069),
.B(n_1059),
.Y(n_1251)
);

OAI21x1_ASAP7_75t_L g1252 ( 
.A1(n_1104),
.A2(n_1114),
.B(n_1105),
.Y(n_1252)
);

AOI21x1_ASAP7_75t_L g1253 ( 
.A1(n_1091),
.A2(n_1095),
.B(n_1105),
.Y(n_1253)
);

AOI221x1_ASAP7_75t_L g1254 ( 
.A1(n_1166),
.A2(n_1160),
.B1(n_1168),
.B2(n_1146),
.C(n_1114),
.Y(n_1254)
);

BUFx8_ASAP7_75t_L g1255 ( 
.A(n_1053),
.Y(n_1255)
);

INVx1_ASAP7_75t_L g1256 ( 
.A(n_1060),
.Y(n_1256)
);

BUFx10_ASAP7_75t_L g1257 ( 
.A(n_1064),
.Y(n_1257)
);

AO31x2_ASAP7_75t_L g1258 ( 
.A1(n_1057),
.A2(n_1168),
.A3(n_1093),
.B(n_1125),
.Y(n_1258)
);

OAI21x1_ASAP7_75t_L g1259 ( 
.A1(n_1152),
.A2(n_1141),
.B(n_1144),
.Y(n_1259)
);

INVx5_ASAP7_75t_SL g1260 ( 
.A(n_1064),
.Y(n_1260)
);

AOI21xp5_ASAP7_75t_L g1261 ( 
.A1(n_1165),
.A2(n_1108),
.B(n_1158),
.Y(n_1261)
);

OAI21x1_ASAP7_75t_L g1262 ( 
.A1(n_1158),
.A2(n_1046),
.B(n_1071),
.Y(n_1262)
);

BUFx2_ASAP7_75t_L g1263 ( 
.A(n_1064),
.Y(n_1263)
);

AOI21xp5_ASAP7_75t_L g1264 ( 
.A1(n_1052),
.A2(n_1043),
.B(n_1066),
.Y(n_1264)
);

INVx1_ASAP7_75t_L g1265 ( 
.A(n_1039),
.Y(n_1265)
);

AO31x2_ASAP7_75t_L g1266 ( 
.A1(n_1039),
.A2(n_1117),
.A3(n_1172),
.B(n_1102),
.Y(n_1266)
);

INVx2_ASAP7_75t_L g1267 ( 
.A(n_1066),
.Y(n_1267)
);

INVx5_ASAP7_75t_L g1268 ( 
.A(n_1070),
.Y(n_1268)
);

NAND2xp5_ASAP7_75t_L g1269 ( 
.A(n_1073),
.B(n_1070),
.Y(n_1269)
);

AO21x1_ASAP7_75t_L g1270 ( 
.A1(n_1103),
.A2(n_1083),
.B(n_1106),
.Y(n_1270)
);

NOR2xp33_ASAP7_75t_L g1271 ( 
.A(n_1073),
.B(n_1103),
.Y(n_1271)
);

NAND2xp5_ASAP7_75t_L g1272 ( 
.A(n_1150),
.B(n_1115),
.Y(n_1272)
);

INVx1_ASAP7_75t_L g1273 ( 
.A(n_1083),
.Y(n_1273)
);

O2A1O1Ixp33_ASAP7_75t_L g1274 ( 
.A1(n_1106),
.A2(n_1045),
.B(n_977),
.C(n_970),
.Y(n_1274)
);

NOR2xp33_ASAP7_75t_L g1275 ( 
.A(n_1051),
.B(n_353),
.Y(n_1275)
);

AO31x2_ASAP7_75t_L g1276 ( 
.A1(n_1157),
.A2(n_1074),
.A3(n_1045),
.B(n_1048),
.Y(n_1276)
);

AND2x2_ASAP7_75t_L g1277 ( 
.A(n_1051),
.B(n_858),
.Y(n_1277)
);

AO31x2_ASAP7_75t_L g1278 ( 
.A1(n_1157),
.A2(n_1074),
.A3(n_1045),
.B(n_1048),
.Y(n_1278)
);

AOI221x1_ASAP7_75t_L g1279 ( 
.A1(n_1045),
.A2(n_977),
.B1(n_970),
.B2(n_1023),
.C(n_1074),
.Y(n_1279)
);

AOI22xp33_ASAP7_75t_L g1280 ( 
.A1(n_1023),
.A2(n_782),
.B1(n_851),
.B2(n_970),
.Y(n_1280)
);

NAND2xp5_ASAP7_75t_L g1281 ( 
.A(n_1051),
.B(n_980),
.Y(n_1281)
);

CKINVDCx5p33_ASAP7_75t_R g1282 ( 
.A(n_1033),
.Y(n_1282)
);

NOR2xp33_ASAP7_75t_L g1283 ( 
.A(n_1051),
.B(n_353),
.Y(n_1283)
);

AOI21xp5_ASAP7_75t_L g1284 ( 
.A1(n_1074),
.A2(n_543),
.B(n_966),
.Y(n_1284)
);

AO31x2_ASAP7_75t_L g1285 ( 
.A1(n_1157),
.A2(n_1074),
.A3(n_1045),
.B(n_1048),
.Y(n_1285)
);

AO31x2_ASAP7_75t_L g1286 ( 
.A1(n_1157),
.A2(n_1074),
.A3(n_1045),
.B(n_1048),
.Y(n_1286)
);

NAND2xp5_ASAP7_75t_L g1287 ( 
.A(n_1051),
.B(n_980),
.Y(n_1287)
);

NAND2xp5_ASAP7_75t_L g1288 ( 
.A(n_1051),
.B(n_980),
.Y(n_1288)
);

AO31x2_ASAP7_75t_L g1289 ( 
.A1(n_1157),
.A2(n_1074),
.A3(n_1045),
.B(n_1048),
.Y(n_1289)
);

NAND2xp5_ASAP7_75t_L g1290 ( 
.A(n_1051),
.B(n_980),
.Y(n_1290)
);

AOI21xp5_ASAP7_75t_L g1291 ( 
.A1(n_1074),
.A2(n_543),
.B(n_966),
.Y(n_1291)
);

A2O1A1Ixp33_ASAP7_75t_L g1292 ( 
.A1(n_1045),
.A2(n_977),
.B(n_1038),
.C(n_1023),
.Y(n_1292)
);

INVx1_ASAP7_75t_SL g1293 ( 
.A(n_1077),
.Y(n_1293)
);

O2A1O1Ixp5_ASAP7_75t_L g1294 ( 
.A1(n_1045),
.A2(n_977),
.B(n_970),
.C(n_697),
.Y(n_1294)
);

BUFx6f_ASAP7_75t_L g1295 ( 
.A(n_1050),
.Y(n_1295)
);

INVxp67_ASAP7_75t_SL g1296 ( 
.A(n_1040),
.Y(n_1296)
);

OAI21x1_ASAP7_75t_L g1297 ( 
.A1(n_1088),
.A2(n_1030),
.B(n_893),
.Y(n_1297)
);

BUFx2_ASAP7_75t_R g1298 ( 
.A(n_1081),
.Y(n_1298)
);

NOR2xp33_ASAP7_75t_L g1299 ( 
.A(n_1051),
.B(n_353),
.Y(n_1299)
);

AOI21xp5_ASAP7_75t_L g1300 ( 
.A1(n_1074),
.A2(n_543),
.B(n_966),
.Y(n_1300)
);

OAI21xp5_ASAP7_75t_L g1301 ( 
.A1(n_1045),
.A2(n_977),
.B(n_1038),
.Y(n_1301)
);

NAND2x2_ASAP7_75t_L g1302 ( 
.A(n_1081),
.B(n_864),
.Y(n_1302)
);

AOI21xp5_ASAP7_75t_L g1303 ( 
.A1(n_1074),
.A2(n_543),
.B(n_966),
.Y(n_1303)
);

OAI21x1_ASAP7_75t_L g1304 ( 
.A1(n_1088),
.A2(n_1030),
.B(n_893),
.Y(n_1304)
);

AOI21xp5_ASAP7_75t_L g1305 ( 
.A1(n_1074),
.A2(n_543),
.B(n_966),
.Y(n_1305)
);

AOI21xp5_ASAP7_75t_L g1306 ( 
.A1(n_1074),
.A2(n_543),
.B(n_966),
.Y(n_1306)
);

INVxp67_ASAP7_75t_SL g1307 ( 
.A(n_1040),
.Y(n_1307)
);

AOI22xp33_ASAP7_75t_L g1308 ( 
.A1(n_1023),
.A2(n_782),
.B1(n_851),
.B2(n_970),
.Y(n_1308)
);

NAND2xp5_ASAP7_75t_L g1309 ( 
.A(n_1051),
.B(n_980),
.Y(n_1309)
);

OAI21x1_ASAP7_75t_L g1310 ( 
.A1(n_1088),
.A2(n_1030),
.B(n_893),
.Y(n_1310)
);

A2O1A1Ixp33_ASAP7_75t_L g1311 ( 
.A1(n_1045),
.A2(n_977),
.B(n_1038),
.C(n_1023),
.Y(n_1311)
);

HB1xp67_ASAP7_75t_L g1312 ( 
.A(n_1031),
.Y(n_1312)
);

INVx1_ASAP7_75t_L g1313 ( 
.A(n_1142),
.Y(n_1313)
);

CKINVDCx20_ASAP7_75t_R g1314 ( 
.A(n_1033),
.Y(n_1314)
);

AOI221xp5_ASAP7_75t_SL g1315 ( 
.A1(n_1045),
.A2(n_725),
.B1(n_448),
.B2(n_696),
.C(n_970),
.Y(n_1315)
);

OAI21x1_ASAP7_75t_L g1316 ( 
.A1(n_1088),
.A2(n_1030),
.B(n_893),
.Y(n_1316)
);

OR2x2_ASAP7_75t_L g1317 ( 
.A(n_1041),
.B(n_688),
.Y(n_1317)
);

AO31x2_ASAP7_75t_L g1318 ( 
.A1(n_1157),
.A2(n_1074),
.A3(n_1045),
.B(n_1048),
.Y(n_1318)
);

NOR2xp33_ASAP7_75t_L g1319 ( 
.A(n_1051),
.B(n_353),
.Y(n_1319)
);

AO31x2_ASAP7_75t_L g1320 ( 
.A1(n_1157),
.A2(n_1074),
.A3(n_1045),
.B(n_1048),
.Y(n_1320)
);

AOI22xp5_ASAP7_75t_L g1321 ( 
.A1(n_1045),
.A2(n_970),
.B1(n_671),
.B2(n_906),
.Y(n_1321)
);

OAI21x1_ASAP7_75t_L g1322 ( 
.A1(n_1088),
.A2(n_1030),
.B(n_893),
.Y(n_1322)
);

HB1xp67_ASAP7_75t_L g1323 ( 
.A(n_1031),
.Y(n_1323)
);

AOI222xp33_ASAP7_75t_L g1324 ( 
.A1(n_1058),
.A2(n_696),
.B1(n_782),
.B2(n_725),
.C1(n_732),
.C2(n_851),
.Y(n_1324)
);

BUFx6f_ASAP7_75t_L g1325 ( 
.A(n_1050),
.Y(n_1325)
);

BUFx8_ASAP7_75t_SL g1326 ( 
.A(n_1195),
.Y(n_1326)
);

BUFx2_ASAP7_75t_SL g1327 ( 
.A(n_1314),
.Y(n_1327)
);

OAI22xp5_ASAP7_75t_L g1328 ( 
.A1(n_1219),
.A2(n_1311),
.B1(n_1292),
.B2(n_1301),
.Y(n_1328)
);

NAND2xp5_ASAP7_75t_L g1329 ( 
.A(n_1321),
.B(n_1315),
.Y(n_1329)
);

INVx1_ASAP7_75t_L g1330 ( 
.A(n_1203),
.Y(n_1330)
);

INVx6_ASAP7_75t_L g1331 ( 
.A(n_1255),
.Y(n_1331)
);

BUFx6f_ASAP7_75t_L g1332 ( 
.A(n_1188),
.Y(n_1332)
);

BUFx12f_ASAP7_75t_L g1333 ( 
.A(n_1282),
.Y(n_1333)
);

AOI22xp33_ASAP7_75t_L g1334 ( 
.A1(n_1280),
.A2(n_1308),
.B1(n_1324),
.B2(n_1277),
.Y(n_1334)
);

OAI21xp5_ASAP7_75t_L g1335 ( 
.A1(n_1294),
.A2(n_1279),
.B(n_1274),
.Y(n_1335)
);

AND2x2_ASAP7_75t_L g1336 ( 
.A(n_1275),
.B(n_1283),
.Y(n_1336)
);

INVx1_ASAP7_75t_L g1337 ( 
.A(n_1231),
.Y(n_1337)
);

BUFx8_ASAP7_75t_SL g1338 ( 
.A(n_1178),
.Y(n_1338)
);

BUFx2_ASAP7_75t_L g1339 ( 
.A(n_1198),
.Y(n_1339)
);

INVx1_ASAP7_75t_L g1340 ( 
.A(n_1197),
.Y(n_1340)
);

AOI22xp33_ASAP7_75t_SL g1341 ( 
.A1(n_1299),
.A2(n_1319),
.B1(n_1251),
.B2(n_1287),
.Y(n_1341)
);

CKINVDCx11_ASAP7_75t_R g1342 ( 
.A(n_1196),
.Y(n_1342)
);

AOI22xp33_ASAP7_75t_L g1343 ( 
.A1(n_1281),
.A2(n_1309),
.B1(n_1290),
.B2(n_1288),
.Y(n_1343)
);

CKINVDCx11_ASAP7_75t_R g1344 ( 
.A(n_1302),
.Y(n_1344)
);

AOI22xp33_ASAP7_75t_SL g1345 ( 
.A1(n_1189),
.A2(n_1228),
.B1(n_1192),
.B2(n_1223),
.Y(n_1345)
);

CKINVDCx20_ASAP7_75t_R g1346 ( 
.A(n_1182),
.Y(n_1346)
);

OAI22xp33_ASAP7_75t_L g1347 ( 
.A1(n_1317),
.A2(n_1173),
.B1(n_1293),
.B2(n_1221),
.Y(n_1347)
);

INVxp67_ASAP7_75t_L g1348 ( 
.A(n_1200),
.Y(n_1348)
);

BUFx6f_ASAP7_75t_L g1349 ( 
.A(n_1188),
.Y(n_1349)
);

BUFx3_ASAP7_75t_L g1350 ( 
.A(n_1255),
.Y(n_1350)
);

CKINVDCx6p67_ASAP7_75t_R g1351 ( 
.A(n_1188),
.Y(n_1351)
);

OAI22xp5_ASAP7_75t_L g1352 ( 
.A1(n_1248),
.A2(n_1226),
.B1(n_1296),
.B2(n_1307),
.Y(n_1352)
);

INVx11_ASAP7_75t_L g1353 ( 
.A(n_1260),
.Y(n_1353)
);

AOI22xp5_ASAP7_75t_L g1354 ( 
.A1(n_1199),
.A2(n_1233),
.B1(n_1206),
.B2(n_1176),
.Y(n_1354)
);

CKINVDCx20_ASAP7_75t_R g1355 ( 
.A(n_1244),
.Y(n_1355)
);

OAI22xp5_ASAP7_75t_L g1356 ( 
.A1(n_1194),
.A2(n_1224),
.B1(n_1237),
.B2(n_1210),
.Y(n_1356)
);

OAI22xp33_ASAP7_75t_SL g1357 ( 
.A1(n_1177),
.A2(n_1229),
.B1(n_1323),
.B2(n_1312),
.Y(n_1357)
);

INVx6_ASAP7_75t_L g1358 ( 
.A(n_1257),
.Y(n_1358)
);

AOI22xp33_ASAP7_75t_SL g1359 ( 
.A1(n_1261),
.A2(n_1233),
.B1(n_1250),
.B2(n_1220),
.Y(n_1359)
);

INVx1_ASAP7_75t_SL g1360 ( 
.A(n_1263),
.Y(n_1360)
);

NAND2x1p5_ASAP7_75t_L g1361 ( 
.A(n_1268),
.B(n_1229),
.Y(n_1361)
);

OAI22xp5_ASAP7_75t_L g1362 ( 
.A1(n_1272),
.A2(n_1265),
.B1(n_1313),
.B2(n_1227),
.Y(n_1362)
);

AOI22xp33_ASAP7_75t_SL g1363 ( 
.A1(n_1249),
.A2(n_1183),
.B1(n_1222),
.B2(n_1193),
.Y(n_1363)
);

INVx1_ASAP7_75t_SL g1364 ( 
.A(n_1298),
.Y(n_1364)
);

BUFx2_ASAP7_75t_L g1365 ( 
.A(n_1242),
.Y(n_1365)
);

CKINVDCx11_ASAP7_75t_R g1366 ( 
.A(n_1257),
.Y(n_1366)
);

OAI21xp33_ASAP7_75t_SL g1367 ( 
.A1(n_1179),
.A2(n_1256),
.B(n_1205),
.Y(n_1367)
);

CKINVDCx6p67_ASAP7_75t_R g1368 ( 
.A(n_1268),
.Y(n_1368)
);

AOI22xp33_ASAP7_75t_L g1369 ( 
.A1(n_1217),
.A2(n_1273),
.B1(n_1270),
.B2(n_1216),
.Y(n_1369)
);

AOI22xp33_ASAP7_75t_L g1370 ( 
.A1(n_1273),
.A2(n_1216),
.B1(n_1256),
.B2(n_1246),
.Y(n_1370)
);

NAND2xp5_ASAP7_75t_L g1371 ( 
.A(n_1239),
.B(n_1232),
.Y(n_1371)
);

OAI22xp5_ASAP7_75t_L g1372 ( 
.A1(n_1187),
.A2(n_1268),
.B1(n_1260),
.B2(n_1174),
.Y(n_1372)
);

AOI22xp33_ASAP7_75t_L g1373 ( 
.A1(n_1267),
.A2(n_1240),
.B1(n_1271),
.B2(n_1235),
.Y(n_1373)
);

OAI22xp33_ASAP7_75t_L g1374 ( 
.A1(n_1254),
.A2(n_1215),
.B1(n_1212),
.B2(n_1181),
.Y(n_1374)
);

CKINVDCx11_ASAP7_75t_R g1375 ( 
.A(n_1208),
.Y(n_1375)
);

OAI21xp5_ASAP7_75t_SL g1376 ( 
.A1(n_1218),
.A2(n_1180),
.B(n_1291),
.Y(n_1376)
);

INVx1_ASAP7_75t_L g1377 ( 
.A(n_1269),
.Y(n_1377)
);

CKINVDCx11_ASAP7_75t_R g1378 ( 
.A(n_1208),
.Y(n_1378)
);

INVx1_ASAP7_75t_L g1379 ( 
.A(n_1243),
.Y(n_1379)
);

INVx6_ASAP7_75t_L g1380 ( 
.A(n_1208),
.Y(n_1380)
);

CKINVDCx8_ASAP7_75t_R g1381 ( 
.A(n_1325),
.Y(n_1381)
);

AOI22xp33_ASAP7_75t_SL g1382 ( 
.A1(n_1284),
.A2(n_1306),
.B1(n_1305),
.B2(n_1303),
.Y(n_1382)
);

BUFx6f_ASAP7_75t_L g1383 ( 
.A(n_1295),
.Y(n_1383)
);

OAI22xp5_ASAP7_75t_L g1384 ( 
.A1(n_1234),
.A2(n_1204),
.B1(n_1201),
.B2(n_1230),
.Y(n_1384)
);

INVx6_ASAP7_75t_L g1385 ( 
.A(n_1295),
.Y(n_1385)
);

INVx3_ASAP7_75t_L g1386 ( 
.A(n_1213),
.Y(n_1386)
);

AOI22xp33_ASAP7_75t_SL g1387 ( 
.A1(n_1300),
.A2(n_1201),
.B1(n_1266),
.B2(n_1262),
.Y(n_1387)
);

BUFx12f_ASAP7_75t_L g1388 ( 
.A(n_1264),
.Y(n_1388)
);

CKINVDCx20_ASAP7_75t_R g1389 ( 
.A(n_1247),
.Y(n_1389)
);

INVx1_ASAP7_75t_L g1390 ( 
.A(n_1253),
.Y(n_1390)
);

OAI22xp5_ASAP7_75t_L g1391 ( 
.A1(n_1201),
.A2(n_1241),
.B1(n_1214),
.B2(n_1245),
.Y(n_1391)
);

AOI22xp33_ASAP7_75t_L g1392 ( 
.A1(n_1247),
.A2(n_1252),
.B1(n_1175),
.B2(n_1238),
.Y(n_1392)
);

INVx6_ASAP7_75t_L g1393 ( 
.A(n_1185),
.Y(n_1393)
);

AND2x4_ASAP7_75t_L g1394 ( 
.A(n_1266),
.B(n_1289),
.Y(n_1394)
);

AOI22xp33_ASAP7_75t_SL g1395 ( 
.A1(n_1266),
.A2(n_1202),
.B1(n_1175),
.B2(n_1209),
.Y(n_1395)
);

BUFx2_ASAP7_75t_L g1396 ( 
.A(n_1276),
.Y(n_1396)
);

BUFx10_ASAP7_75t_L g1397 ( 
.A(n_1236),
.Y(n_1397)
);

AOI22xp33_ASAP7_75t_SL g1398 ( 
.A1(n_1202),
.A2(n_1278),
.B1(n_1320),
.B2(n_1318),
.Y(n_1398)
);

BUFx12f_ASAP7_75t_L g1399 ( 
.A(n_1191),
.Y(n_1399)
);

AOI22xp33_ASAP7_75t_L g1400 ( 
.A1(n_1225),
.A2(n_1190),
.B1(n_1316),
.B2(n_1322),
.Y(n_1400)
);

OAI22xp5_ASAP7_75t_L g1401 ( 
.A1(n_1276),
.A2(n_1278),
.B1(n_1318),
.B2(n_1289),
.Y(n_1401)
);

AOI22xp5_ASAP7_75t_L g1402 ( 
.A1(n_1297),
.A2(n_1310),
.B1(n_1304),
.B2(n_1259),
.Y(n_1402)
);

BUFx12f_ASAP7_75t_L g1403 ( 
.A(n_1191),
.Y(n_1403)
);

OAI22xp5_ASAP7_75t_L g1404 ( 
.A1(n_1285),
.A2(n_1318),
.B1(n_1289),
.B2(n_1286),
.Y(n_1404)
);

OAI22xp5_ASAP7_75t_L g1405 ( 
.A1(n_1285),
.A2(n_1286),
.B1(n_1320),
.B2(n_1207),
.Y(n_1405)
);

CKINVDCx20_ASAP7_75t_R g1406 ( 
.A(n_1285),
.Y(n_1406)
);

AOI22xp33_ASAP7_75t_SL g1407 ( 
.A1(n_1258),
.A2(n_1191),
.B1(n_1207),
.B2(n_1186),
.Y(n_1407)
);

CKINVDCx11_ASAP7_75t_R g1408 ( 
.A(n_1186),
.Y(n_1408)
);

AOI22xp33_ASAP7_75t_L g1409 ( 
.A1(n_1258),
.A2(n_1186),
.B1(n_1211),
.B2(n_1184),
.Y(n_1409)
);

CKINVDCx5p33_ASAP7_75t_R g1410 ( 
.A(n_1184),
.Y(n_1410)
);

INVx5_ASAP7_75t_L g1411 ( 
.A(n_1211),
.Y(n_1411)
);

BUFx8_ASAP7_75t_L g1412 ( 
.A(n_1258),
.Y(n_1412)
);

BUFx4_ASAP7_75t_SL g1413 ( 
.A(n_1195),
.Y(n_1413)
);

BUFx6f_ASAP7_75t_L g1414 ( 
.A(n_1188),
.Y(n_1414)
);

INVx1_ASAP7_75t_SL g1415 ( 
.A(n_1173),
.Y(n_1415)
);

INVx1_ASAP7_75t_L g1416 ( 
.A(n_1203),
.Y(n_1416)
);

CKINVDCx20_ASAP7_75t_R g1417 ( 
.A(n_1314),
.Y(n_1417)
);

BUFx6f_ASAP7_75t_L g1418 ( 
.A(n_1188),
.Y(n_1418)
);

AOI22xp33_ASAP7_75t_L g1419 ( 
.A1(n_1280),
.A2(n_1308),
.B1(n_1324),
.B2(n_906),
.Y(n_1419)
);

AOI22xp33_ASAP7_75t_L g1420 ( 
.A1(n_1280),
.A2(n_1308),
.B1(n_1324),
.B2(n_906),
.Y(n_1420)
);

INVx3_ASAP7_75t_L g1421 ( 
.A(n_1257),
.Y(n_1421)
);

AOI22xp33_ASAP7_75t_L g1422 ( 
.A1(n_1280),
.A2(n_1308),
.B1(n_1324),
.B2(n_906),
.Y(n_1422)
);

OAI21xp33_ASAP7_75t_L g1423 ( 
.A1(n_1280),
.A2(n_970),
.B(n_676),
.Y(n_1423)
);

INVx1_ASAP7_75t_SL g1424 ( 
.A(n_1173),
.Y(n_1424)
);

CKINVDCx5p33_ASAP7_75t_R g1425 ( 
.A(n_1192),
.Y(n_1425)
);

NAND2x1p5_ASAP7_75t_L g1426 ( 
.A(n_1188),
.B(n_1268),
.Y(n_1426)
);

AOI22xp33_ASAP7_75t_L g1427 ( 
.A1(n_1280),
.A2(n_1308),
.B1(n_1324),
.B2(n_906),
.Y(n_1427)
);

INVx6_ASAP7_75t_L g1428 ( 
.A(n_1255),
.Y(n_1428)
);

AOI22xp33_ASAP7_75t_SL g1429 ( 
.A1(n_1301),
.A2(n_782),
.B1(n_680),
.B2(n_676),
.Y(n_1429)
);

INVx6_ASAP7_75t_L g1430 ( 
.A(n_1255),
.Y(n_1430)
);

CKINVDCx11_ASAP7_75t_R g1431 ( 
.A(n_1195),
.Y(n_1431)
);

CKINVDCx11_ASAP7_75t_R g1432 ( 
.A(n_1195),
.Y(n_1432)
);

INVx1_ASAP7_75t_L g1433 ( 
.A(n_1203),
.Y(n_1433)
);

INVx1_ASAP7_75t_L g1434 ( 
.A(n_1203),
.Y(n_1434)
);

OAI22xp5_ASAP7_75t_L g1435 ( 
.A1(n_1219),
.A2(n_841),
.B1(n_1045),
.B2(n_1292),
.Y(n_1435)
);

BUFx8_ASAP7_75t_L g1436 ( 
.A(n_1178),
.Y(n_1436)
);

CKINVDCx11_ASAP7_75t_R g1437 ( 
.A(n_1195),
.Y(n_1437)
);

NAND2xp5_ASAP7_75t_L g1438 ( 
.A(n_1301),
.B(n_1045),
.Y(n_1438)
);

AOI22xp33_ASAP7_75t_SL g1439 ( 
.A1(n_1301),
.A2(n_782),
.B1(n_680),
.B2(n_676),
.Y(n_1439)
);

NAND2xp5_ASAP7_75t_L g1440 ( 
.A(n_1281),
.B(n_1287),
.Y(n_1440)
);

CKINVDCx11_ASAP7_75t_R g1441 ( 
.A(n_1195),
.Y(n_1441)
);

OAI22xp5_ASAP7_75t_L g1442 ( 
.A1(n_1219),
.A2(n_841),
.B1(n_1045),
.B2(n_1292),
.Y(n_1442)
);

OAI21xp5_ASAP7_75t_L g1443 ( 
.A1(n_1292),
.A2(n_1311),
.B(n_1301),
.Y(n_1443)
);

AOI22xp33_ASAP7_75t_L g1444 ( 
.A1(n_1280),
.A2(n_1308),
.B1(n_1324),
.B2(n_906),
.Y(n_1444)
);

BUFx10_ASAP7_75t_L g1445 ( 
.A(n_1282),
.Y(n_1445)
);

INVx4_ASAP7_75t_L g1446 ( 
.A(n_1188),
.Y(n_1446)
);

CKINVDCx16_ASAP7_75t_R g1447 ( 
.A(n_1314),
.Y(n_1447)
);

INVx2_ASAP7_75t_L g1448 ( 
.A(n_1340),
.Y(n_1448)
);

HB1xp67_ASAP7_75t_L g1449 ( 
.A(n_1415),
.Y(n_1449)
);

AND2x2_ASAP7_75t_L g1450 ( 
.A(n_1396),
.B(n_1406),
.Y(n_1450)
);

AO21x2_ASAP7_75t_L g1451 ( 
.A1(n_1335),
.A2(n_1374),
.B(n_1402),
.Y(n_1451)
);

HB1xp67_ASAP7_75t_L g1452 ( 
.A(n_1415),
.Y(n_1452)
);

OAI21x1_ASAP7_75t_L g1453 ( 
.A1(n_1392),
.A2(n_1400),
.B(n_1390),
.Y(n_1453)
);

BUFx3_ASAP7_75t_L g1454 ( 
.A(n_1361),
.Y(n_1454)
);

INVx1_ASAP7_75t_L g1455 ( 
.A(n_1410),
.Y(n_1455)
);

INVx6_ASAP7_75t_L g1456 ( 
.A(n_1332),
.Y(n_1456)
);

AND2x2_ASAP7_75t_L g1457 ( 
.A(n_1394),
.B(n_1398),
.Y(n_1457)
);

INVx2_ASAP7_75t_SL g1458 ( 
.A(n_1330),
.Y(n_1458)
);

OR2x2_ASAP7_75t_L g1459 ( 
.A(n_1401),
.B(n_1404),
.Y(n_1459)
);

BUFx6f_ASAP7_75t_L g1460 ( 
.A(n_1408),
.Y(n_1460)
);

CKINVDCx11_ASAP7_75t_R g1461 ( 
.A(n_1431),
.Y(n_1461)
);

NAND2xp5_ASAP7_75t_L g1462 ( 
.A(n_1440),
.B(n_1343),
.Y(n_1462)
);

HB1xp67_ASAP7_75t_L g1463 ( 
.A(n_1424),
.Y(n_1463)
);

CKINVDCx12_ASAP7_75t_R g1464 ( 
.A(n_1413),
.Y(n_1464)
);

OA21x2_ASAP7_75t_L g1465 ( 
.A1(n_1335),
.A2(n_1376),
.B(n_1409),
.Y(n_1465)
);

INVx1_ASAP7_75t_L g1466 ( 
.A(n_1371),
.Y(n_1466)
);

INVx1_ASAP7_75t_L g1467 ( 
.A(n_1371),
.Y(n_1467)
);

INVx1_ASAP7_75t_L g1468 ( 
.A(n_1401),
.Y(n_1468)
);

INVx2_ASAP7_75t_L g1469 ( 
.A(n_1416),
.Y(n_1469)
);

INVx2_ASAP7_75t_L g1470 ( 
.A(n_1433),
.Y(n_1470)
);

AND2x2_ASAP7_75t_L g1471 ( 
.A(n_1438),
.B(n_1329),
.Y(n_1471)
);

INVx1_ASAP7_75t_L g1472 ( 
.A(n_1405),
.Y(n_1472)
);

NOR2xp33_ASAP7_75t_L g1473 ( 
.A(n_1336),
.B(n_1339),
.Y(n_1473)
);

INVx1_ASAP7_75t_L g1474 ( 
.A(n_1362),
.Y(n_1474)
);

AND2x2_ASAP7_75t_L g1475 ( 
.A(n_1438),
.B(n_1329),
.Y(n_1475)
);

INVx1_ASAP7_75t_L g1476 ( 
.A(n_1362),
.Y(n_1476)
);

INVx1_ASAP7_75t_L g1477 ( 
.A(n_1399),
.Y(n_1477)
);

AND2x2_ASAP7_75t_L g1478 ( 
.A(n_1443),
.B(n_1377),
.Y(n_1478)
);

INVx1_ASAP7_75t_L g1479 ( 
.A(n_1403),
.Y(n_1479)
);

OR2x6_ASAP7_75t_L g1480 ( 
.A(n_1443),
.B(n_1376),
.Y(n_1480)
);

INVx2_ASAP7_75t_SL g1481 ( 
.A(n_1434),
.Y(n_1481)
);

NOR2xp33_ASAP7_75t_L g1482 ( 
.A(n_1447),
.B(n_1345),
.Y(n_1482)
);

AND2x4_ASAP7_75t_L g1483 ( 
.A(n_1411),
.B(n_1373),
.Y(n_1483)
);

INVx1_ASAP7_75t_L g1484 ( 
.A(n_1389),
.Y(n_1484)
);

INVx1_ASAP7_75t_L g1485 ( 
.A(n_1412),
.Y(n_1485)
);

INVx1_ASAP7_75t_L g1486 ( 
.A(n_1412),
.Y(n_1486)
);

HB1xp67_ASAP7_75t_L g1487 ( 
.A(n_1424),
.Y(n_1487)
);

INVx1_ASAP7_75t_L g1488 ( 
.A(n_1391),
.Y(n_1488)
);

INVx1_ASAP7_75t_L g1489 ( 
.A(n_1395),
.Y(n_1489)
);

INVx1_ASAP7_75t_L g1490 ( 
.A(n_1407),
.Y(n_1490)
);

BUFx2_ASAP7_75t_L g1491 ( 
.A(n_1367),
.Y(n_1491)
);

INVx1_ASAP7_75t_L g1492 ( 
.A(n_1328),
.Y(n_1492)
);

INVx1_ASAP7_75t_L g1493 ( 
.A(n_1328),
.Y(n_1493)
);

INVx1_ASAP7_75t_L g1494 ( 
.A(n_1384),
.Y(n_1494)
);

INVx1_ASAP7_75t_L g1495 ( 
.A(n_1384),
.Y(n_1495)
);

OR2x6_ASAP7_75t_L g1496 ( 
.A(n_1435),
.B(n_1442),
.Y(n_1496)
);

OAI22xp5_ASAP7_75t_SL g1497 ( 
.A1(n_1429),
.A2(n_1439),
.B1(n_1419),
.B2(n_1427),
.Y(n_1497)
);

INVx2_ASAP7_75t_SL g1498 ( 
.A(n_1332),
.Y(n_1498)
);

HB1xp67_ASAP7_75t_L g1499 ( 
.A(n_1348),
.Y(n_1499)
);

AOI21x1_ASAP7_75t_L g1500 ( 
.A1(n_1435),
.A2(n_1442),
.B(n_1372),
.Y(n_1500)
);

INVx4_ASAP7_75t_L g1501 ( 
.A(n_1388),
.Y(n_1501)
);

AOI21x1_ASAP7_75t_L g1502 ( 
.A1(n_1372),
.A2(n_1352),
.B(n_1356),
.Y(n_1502)
);

NOR2x1_ASAP7_75t_SL g1503 ( 
.A(n_1352),
.B(n_1356),
.Y(n_1503)
);

BUFx3_ASAP7_75t_L g1504 ( 
.A(n_1436),
.Y(n_1504)
);

BUFx12f_ASAP7_75t_L g1505 ( 
.A(n_1432),
.Y(n_1505)
);

INVx2_ASAP7_75t_SL g1506 ( 
.A(n_1332),
.Y(n_1506)
);

BUFx3_ASAP7_75t_L g1507 ( 
.A(n_1436),
.Y(n_1507)
);

INVxp67_ASAP7_75t_L g1508 ( 
.A(n_1365),
.Y(n_1508)
);

CKINVDCx5p33_ASAP7_75t_R g1509 ( 
.A(n_1326),
.Y(n_1509)
);

OR2x6_ASAP7_75t_L g1510 ( 
.A(n_1393),
.B(n_1426),
.Y(n_1510)
);

AND2x2_ASAP7_75t_L g1511 ( 
.A(n_1387),
.B(n_1337),
.Y(n_1511)
);

INVx1_ASAP7_75t_L g1512 ( 
.A(n_1393),
.Y(n_1512)
);

HB1xp67_ASAP7_75t_L g1513 ( 
.A(n_1360),
.Y(n_1513)
);

NAND2xp5_ASAP7_75t_L g1514 ( 
.A(n_1347),
.B(n_1341),
.Y(n_1514)
);

INVx2_ASAP7_75t_SL g1515 ( 
.A(n_1349),
.Y(n_1515)
);

INVx1_ASAP7_75t_L g1516 ( 
.A(n_1397),
.Y(n_1516)
);

INVx2_ASAP7_75t_L g1517 ( 
.A(n_1397),
.Y(n_1517)
);

INVx2_ASAP7_75t_L g1518 ( 
.A(n_1379),
.Y(n_1518)
);

INVx1_ASAP7_75t_L g1519 ( 
.A(n_1357),
.Y(n_1519)
);

INVx2_ASAP7_75t_SL g1520 ( 
.A(n_1349),
.Y(n_1520)
);

INVx1_ASAP7_75t_L g1521 ( 
.A(n_1382),
.Y(n_1521)
);

BUFx6f_ASAP7_75t_L g1522 ( 
.A(n_1349),
.Y(n_1522)
);

HB1xp67_ASAP7_75t_L g1523 ( 
.A(n_1360),
.Y(n_1523)
);

INVx1_ASAP7_75t_L g1524 ( 
.A(n_1363),
.Y(n_1524)
);

INVxp67_ASAP7_75t_SL g1525 ( 
.A(n_1370),
.Y(n_1525)
);

INVx1_ASAP7_75t_L g1526 ( 
.A(n_1369),
.Y(n_1526)
);

INVx1_ASAP7_75t_L g1527 ( 
.A(n_1359),
.Y(n_1527)
);

BUFx3_ASAP7_75t_L g1528 ( 
.A(n_1354),
.Y(n_1528)
);

INVx4_ASAP7_75t_L g1529 ( 
.A(n_1414),
.Y(n_1529)
);

NAND2x1_ASAP7_75t_L g1530 ( 
.A(n_1446),
.B(n_1386),
.Y(n_1530)
);

INVxp67_ASAP7_75t_L g1531 ( 
.A(n_1338),
.Y(n_1531)
);

BUFx3_ASAP7_75t_L g1532 ( 
.A(n_1331),
.Y(n_1532)
);

INVx1_ASAP7_75t_L g1533 ( 
.A(n_1446),
.Y(n_1533)
);

AOI21xp5_ASAP7_75t_L g1534 ( 
.A1(n_1480),
.A2(n_1423),
.B(n_1444),
.Y(n_1534)
);

INVx1_ASAP7_75t_SL g1535 ( 
.A(n_1449),
.Y(n_1535)
);

NAND2xp5_ASAP7_75t_L g1536 ( 
.A(n_1471),
.B(n_1475),
.Y(n_1536)
);

NAND2xp5_ASAP7_75t_L g1537 ( 
.A(n_1471),
.B(n_1422),
.Y(n_1537)
);

O2A1O1Ixp33_ASAP7_75t_SL g1538 ( 
.A1(n_1516),
.A2(n_1364),
.B(n_1355),
.C(n_1417),
.Y(n_1538)
);

AND2x2_ASAP7_75t_SL g1539 ( 
.A(n_1491),
.B(n_1420),
.Y(n_1539)
);

AND2x2_ASAP7_75t_L g1540 ( 
.A(n_1484),
.B(n_1327),
.Y(n_1540)
);

CKINVDCx20_ASAP7_75t_R g1541 ( 
.A(n_1461),
.Y(n_1541)
);

OR2x2_ASAP7_75t_L g1542 ( 
.A(n_1455),
.B(n_1364),
.Y(n_1542)
);

AND2x4_ASAP7_75t_L g1543 ( 
.A(n_1477),
.B(n_1350),
.Y(n_1543)
);

NAND2xp5_ASAP7_75t_L g1544 ( 
.A(n_1475),
.B(n_1334),
.Y(n_1544)
);

NOR2x1_ASAP7_75t_L g1545 ( 
.A(n_1501),
.B(n_1421),
.Y(n_1545)
);

O2A1O1Ixp33_ASAP7_75t_SL g1546 ( 
.A1(n_1516),
.A2(n_1346),
.B(n_1351),
.C(n_1368),
.Y(n_1546)
);

NOR2xp33_ASAP7_75t_L g1547 ( 
.A(n_1462),
.B(n_1331),
.Y(n_1547)
);

OR2x2_ASAP7_75t_L g1548 ( 
.A(n_1455),
.B(n_1425),
.Y(n_1548)
);

OA21x2_ASAP7_75t_L g1549 ( 
.A1(n_1453),
.A2(n_1381),
.B(n_1385),
.Y(n_1549)
);

AOI22xp5_ASAP7_75t_L g1550 ( 
.A1(n_1497),
.A2(n_1344),
.B1(n_1430),
.B2(n_1428),
.Y(n_1550)
);

OAI211xp5_ASAP7_75t_L g1551 ( 
.A1(n_1514),
.A2(n_1342),
.B(n_1366),
.C(n_1437),
.Y(n_1551)
);

AND2x2_ASAP7_75t_L g1552 ( 
.A(n_1450),
.B(n_1445),
.Y(n_1552)
);

AND2x4_ASAP7_75t_L g1553 ( 
.A(n_1477),
.B(n_1383),
.Y(n_1553)
);

O2A1O1Ixp33_ASAP7_75t_SL g1554 ( 
.A1(n_1512),
.A2(n_1428),
.B(n_1430),
.C(n_1441),
.Y(n_1554)
);

BUFx3_ASAP7_75t_L g1555 ( 
.A(n_1532),
.Y(n_1555)
);

OA21x2_ASAP7_75t_L g1556 ( 
.A1(n_1453),
.A2(n_1380),
.B(n_1385),
.Y(n_1556)
);

AO32x2_ASAP7_75t_L g1557 ( 
.A1(n_1458),
.A2(n_1378),
.A3(n_1375),
.B1(n_1445),
.B2(n_1380),
.Y(n_1557)
);

AOI21xp5_ASAP7_75t_L g1558 ( 
.A1(n_1480),
.A2(n_1414),
.B(n_1418),
.Y(n_1558)
);

OR2x2_ASAP7_75t_L g1559 ( 
.A(n_1452),
.B(n_1383),
.Y(n_1559)
);

AND2x2_ASAP7_75t_L g1560 ( 
.A(n_1519),
.B(n_1383),
.Y(n_1560)
);

OR2x6_ASAP7_75t_L g1561 ( 
.A(n_1480),
.B(n_1414),
.Y(n_1561)
);

INVx1_ASAP7_75t_L g1562 ( 
.A(n_1448),
.Y(n_1562)
);

AND2x4_ASAP7_75t_L g1563 ( 
.A(n_1479),
.B(n_1353),
.Y(n_1563)
);

O2A1O1Ixp33_ASAP7_75t_SL g1564 ( 
.A1(n_1512),
.A2(n_1333),
.B(n_1358),
.C(n_1517),
.Y(n_1564)
);

AND2x2_ASAP7_75t_L g1565 ( 
.A(n_1519),
.B(n_1358),
.Y(n_1565)
);

AND2x2_ASAP7_75t_L g1566 ( 
.A(n_1478),
.B(n_1460),
.Y(n_1566)
);

O2A1O1Ixp33_ASAP7_75t_SL g1567 ( 
.A1(n_1517),
.A2(n_1531),
.B(n_1486),
.C(n_1485),
.Y(n_1567)
);

NOR2xp33_ASAP7_75t_L g1568 ( 
.A(n_1524),
.B(n_1491),
.Y(n_1568)
);

AO32x2_ASAP7_75t_L g1569 ( 
.A1(n_1458),
.A2(n_1481),
.A3(n_1497),
.B1(n_1501),
.B2(n_1498),
.Y(n_1569)
);

OAI21xp5_ASAP7_75t_L g1570 ( 
.A1(n_1500),
.A2(n_1496),
.B(n_1521),
.Y(n_1570)
);

BUFx3_ASAP7_75t_L g1571 ( 
.A(n_1532),
.Y(n_1571)
);

O2A1O1Ixp33_ASAP7_75t_SL g1572 ( 
.A1(n_1485),
.A2(n_1486),
.B(n_1524),
.C(n_1526),
.Y(n_1572)
);

A2O1A1Ixp33_ASAP7_75t_L g1573 ( 
.A1(n_1482),
.A2(n_1526),
.B(n_1521),
.C(n_1525),
.Y(n_1573)
);

A2O1A1Ixp33_ASAP7_75t_L g1574 ( 
.A1(n_1527),
.A2(n_1528),
.B(n_1495),
.C(n_1494),
.Y(n_1574)
);

OAI22xp5_ASAP7_75t_L g1575 ( 
.A1(n_1496),
.A2(n_1492),
.B1(n_1493),
.B2(n_1487),
.Y(n_1575)
);

OAI22xp5_ASAP7_75t_L g1576 ( 
.A1(n_1496),
.A2(n_1493),
.B1(n_1492),
.B2(n_1463),
.Y(n_1576)
);

AO21x1_ASAP7_75t_L g1577 ( 
.A1(n_1527),
.A2(n_1466),
.B(n_1467),
.Y(n_1577)
);

AND2x2_ASAP7_75t_L g1578 ( 
.A(n_1478),
.B(n_1460),
.Y(n_1578)
);

CKINVDCx20_ASAP7_75t_R g1579 ( 
.A(n_1464),
.Y(n_1579)
);

O2A1O1Ixp33_ASAP7_75t_SL g1580 ( 
.A1(n_1530),
.A2(n_1513),
.B(n_1523),
.C(n_1515),
.Y(n_1580)
);

OAI21xp5_ASAP7_75t_L g1581 ( 
.A1(n_1496),
.A2(n_1502),
.B(n_1476),
.Y(n_1581)
);

OAI211xp5_ASAP7_75t_L g1582 ( 
.A1(n_1474),
.A2(n_1499),
.B(n_1465),
.C(n_1528),
.Y(n_1582)
);

NOR2x1_ASAP7_75t_SL g1583 ( 
.A(n_1510),
.B(n_1460),
.Y(n_1583)
);

AND2x2_ASAP7_75t_L g1584 ( 
.A(n_1460),
.B(n_1511),
.Y(n_1584)
);

AND2x2_ASAP7_75t_L g1585 ( 
.A(n_1460),
.B(n_1511),
.Y(n_1585)
);

AO32x2_ASAP7_75t_L g1586 ( 
.A1(n_1481),
.A2(n_1501),
.A3(n_1498),
.B1(n_1506),
.B2(n_1515),
.Y(n_1586)
);

BUFx12f_ASAP7_75t_L g1587 ( 
.A(n_1505),
.Y(n_1587)
);

NOR2xp33_ASAP7_75t_L g1588 ( 
.A(n_1528),
.B(n_1501),
.Y(n_1588)
);

NOR2x1_ASAP7_75t_L g1589 ( 
.A(n_1510),
.B(n_1533),
.Y(n_1589)
);

NAND2x1_ASAP7_75t_L g1590 ( 
.A(n_1510),
.B(n_1466),
.Y(n_1590)
);

NOR2x1_ASAP7_75t_SL g1591 ( 
.A(n_1510),
.B(n_1496),
.Y(n_1591)
);

AOI211xp5_ASAP7_75t_L g1592 ( 
.A1(n_1473),
.A2(n_1489),
.B(n_1508),
.C(n_1490),
.Y(n_1592)
);

BUFx3_ASAP7_75t_L g1593 ( 
.A(n_1532),
.Y(n_1593)
);

OR2x6_ASAP7_75t_L g1594 ( 
.A(n_1483),
.B(n_1510),
.Y(n_1594)
);

AND2x2_ASAP7_75t_L g1595 ( 
.A(n_1566),
.B(n_1457),
.Y(n_1595)
);

INVxp67_ASAP7_75t_SL g1596 ( 
.A(n_1577),
.Y(n_1596)
);

AND2x2_ASAP7_75t_L g1597 ( 
.A(n_1578),
.B(n_1457),
.Y(n_1597)
);

AND2x2_ASAP7_75t_L g1598 ( 
.A(n_1594),
.B(n_1489),
.Y(n_1598)
);

OAI22xp5_ASAP7_75t_L g1599 ( 
.A1(n_1550),
.A2(n_1507),
.B1(n_1504),
.B2(n_1454),
.Y(n_1599)
);

INVx1_ASAP7_75t_SL g1600 ( 
.A(n_1548),
.Y(n_1600)
);

OR2x6_ASAP7_75t_SL g1601 ( 
.A(n_1575),
.B(n_1509),
.Y(n_1601)
);

NOR2x1_ASAP7_75t_L g1602 ( 
.A(n_1589),
.B(n_1454),
.Y(n_1602)
);

INVx1_ASAP7_75t_L g1603 ( 
.A(n_1562),
.Y(n_1603)
);

OR2x2_ASAP7_75t_L g1604 ( 
.A(n_1536),
.B(n_1535),
.Y(n_1604)
);

BUFx2_ASAP7_75t_L g1605 ( 
.A(n_1586),
.Y(n_1605)
);

INVx4_ASAP7_75t_L g1606 ( 
.A(n_1561),
.Y(n_1606)
);

AOI22xp33_ASAP7_75t_L g1607 ( 
.A1(n_1534),
.A2(n_1451),
.B1(n_1483),
.B2(n_1490),
.Y(n_1607)
);

NAND2xp5_ASAP7_75t_L g1608 ( 
.A(n_1536),
.B(n_1469),
.Y(n_1608)
);

NOR2x1p5_ASAP7_75t_L g1609 ( 
.A(n_1587),
.B(n_1505),
.Y(n_1609)
);

OR2x2_ASAP7_75t_L g1610 ( 
.A(n_1581),
.B(n_1459),
.Y(n_1610)
);

NAND2xp5_ASAP7_75t_SL g1611 ( 
.A(n_1588),
.B(n_1454),
.Y(n_1611)
);

NAND2xp5_ASAP7_75t_L g1612 ( 
.A(n_1568),
.B(n_1470),
.Y(n_1612)
);

NOR2x1_ASAP7_75t_L g1613 ( 
.A(n_1588),
.B(n_1507),
.Y(n_1613)
);

AOI22xp33_ASAP7_75t_L g1614 ( 
.A1(n_1534),
.A2(n_1451),
.B1(n_1483),
.B2(n_1465),
.Y(n_1614)
);

INVx1_ASAP7_75t_L g1615 ( 
.A(n_1586),
.Y(n_1615)
);

INVx1_ASAP7_75t_L g1616 ( 
.A(n_1586),
.Y(n_1616)
);

INVx1_ASAP7_75t_L g1617 ( 
.A(n_1556),
.Y(n_1617)
);

NAND2xp5_ASAP7_75t_L g1618 ( 
.A(n_1568),
.B(n_1470),
.Y(n_1618)
);

INVx2_ASAP7_75t_L g1619 ( 
.A(n_1590),
.Y(n_1619)
);

AND2x2_ASAP7_75t_L g1620 ( 
.A(n_1584),
.B(n_1451),
.Y(n_1620)
);

NAND2xp5_ASAP7_75t_SL g1621 ( 
.A(n_1539),
.B(n_1573),
.Y(n_1621)
);

OAI21xp33_ASAP7_75t_L g1622 ( 
.A1(n_1539),
.A2(n_1518),
.B(n_1488),
.Y(n_1622)
);

INVx1_ASAP7_75t_L g1623 ( 
.A(n_1575),
.Y(n_1623)
);

INVx1_ASAP7_75t_L g1624 ( 
.A(n_1576),
.Y(n_1624)
);

OR2x2_ASAP7_75t_L g1625 ( 
.A(n_1581),
.B(n_1459),
.Y(n_1625)
);

AND2x4_ASAP7_75t_L g1626 ( 
.A(n_1617),
.B(n_1591),
.Y(n_1626)
);

INVx3_ASAP7_75t_L g1627 ( 
.A(n_1617),
.Y(n_1627)
);

NAND3xp33_ASAP7_75t_L g1628 ( 
.A(n_1621),
.B(n_1592),
.C(n_1582),
.Y(n_1628)
);

AOI22xp5_ASAP7_75t_L g1629 ( 
.A1(n_1622),
.A2(n_1544),
.B1(n_1537),
.B2(n_1547),
.Y(n_1629)
);

AND2x2_ASAP7_75t_L g1630 ( 
.A(n_1605),
.B(n_1549),
.Y(n_1630)
);

INVx2_ASAP7_75t_L g1631 ( 
.A(n_1615),
.Y(n_1631)
);

OAI211xp5_ASAP7_75t_L g1632 ( 
.A1(n_1596),
.A2(n_1582),
.B(n_1574),
.C(n_1570),
.Y(n_1632)
);

AOI32xp33_ASAP7_75t_L g1633 ( 
.A1(n_1607),
.A2(n_1576),
.A3(n_1585),
.B1(n_1544),
.B2(n_1537),
.Y(n_1633)
);

NAND3xp33_ASAP7_75t_L g1634 ( 
.A(n_1614),
.B(n_1570),
.C(n_1547),
.Y(n_1634)
);

HB1xp67_ASAP7_75t_L g1635 ( 
.A(n_1615),
.Y(n_1635)
);

OR2x2_ASAP7_75t_L g1636 ( 
.A(n_1605),
.B(n_1472),
.Y(n_1636)
);

AND2x2_ASAP7_75t_L g1637 ( 
.A(n_1616),
.B(n_1549),
.Y(n_1637)
);

AND2x2_ASAP7_75t_L g1638 ( 
.A(n_1616),
.B(n_1620),
.Y(n_1638)
);

NOR2xp33_ASAP7_75t_L g1639 ( 
.A(n_1600),
.B(n_1565),
.Y(n_1639)
);

AND2x2_ASAP7_75t_L g1640 ( 
.A(n_1620),
.B(n_1569),
.Y(n_1640)
);

BUFx3_ASAP7_75t_L g1641 ( 
.A(n_1601),
.Y(n_1641)
);

AND2x2_ASAP7_75t_L g1642 ( 
.A(n_1595),
.B(n_1569),
.Y(n_1642)
);

AND2x2_ASAP7_75t_L g1643 ( 
.A(n_1595),
.B(n_1569),
.Y(n_1643)
);

INVx2_ASAP7_75t_L g1644 ( 
.A(n_1603),
.Y(n_1644)
);

AND2x2_ASAP7_75t_L g1645 ( 
.A(n_1597),
.B(n_1472),
.Y(n_1645)
);

AOI31xp33_ASAP7_75t_L g1646 ( 
.A1(n_1599),
.A2(n_1564),
.A3(n_1546),
.B(n_1554),
.Y(n_1646)
);

NAND2xp5_ASAP7_75t_L g1647 ( 
.A(n_1604),
.B(n_1468),
.Y(n_1647)
);

INVx2_ASAP7_75t_SL g1648 ( 
.A(n_1619),
.Y(n_1648)
);

A2O1A1Ixp33_ASAP7_75t_SL g1649 ( 
.A1(n_1623),
.A2(n_1551),
.B(n_1533),
.C(n_1558),
.Y(n_1649)
);

NAND3xp33_ASAP7_75t_L g1650 ( 
.A(n_1610),
.B(n_1572),
.C(n_1560),
.Y(n_1650)
);

INVxp67_ASAP7_75t_SL g1651 ( 
.A(n_1612),
.Y(n_1651)
);

INVxp67_ASAP7_75t_SL g1652 ( 
.A(n_1618),
.Y(n_1652)
);

AND2x4_ASAP7_75t_L g1653 ( 
.A(n_1606),
.B(n_1583),
.Y(n_1653)
);

AND2x4_ASAP7_75t_L g1654 ( 
.A(n_1626),
.B(n_1606),
.Y(n_1654)
);

INVx1_ASAP7_75t_SL g1655 ( 
.A(n_1637),
.Y(n_1655)
);

INVx1_ASAP7_75t_SL g1656 ( 
.A(n_1637),
.Y(n_1656)
);

INVx2_ASAP7_75t_L g1657 ( 
.A(n_1627),
.Y(n_1657)
);

AND2x2_ASAP7_75t_L g1658 ( 
.A(n_1630),
.B(n_1597),
.Y(n_1658)
);

AND2x2_ASAP7_75t_L g1659 ( 
.A(n_1630),
.B(n_1598),
.Y(n_1659)
);

NOR2x1_ASAP7_75t_L g1660 ( 
.A(n_1628),
.B(n_1613),
.Y(n_1660)
);

AND2x2_ASAP7_75t_L g1661 ( 
.A(n_1630),
.B(n_1598),
.Y(n_1661)
);

INVx1_ASAP7_75t_L g1662 ( 
.A(n_1644),
.Y(n_1662)
);

AND2x2_ASAP7_75t_L g1663 ( 
.A(n_1631),
.B(n_1638),
.Y(n_1663)
);

AND2x2_ASAP7_75t_L g1664 ( 
.A(n_1631),
.B(n_1623),
.Y(n_1664)
);

INVx1_ASAP7_75t_L g1665 ( 
.A(n_1644),
.Y(n_1665)
);

AND2x2_ASAP7_75t_L g1666 ( 
.A(n_1631),
.B(n_1624),
.Y(n_1666)
);

INVx2_ASAP7_75t_L g1667 ( 
.A(n_1627),
.Y(n_1667)
);

AND2x4_ASAP7_75t_L g1668 ( 
.A(n_1626),
.B(n_1606),
.Y(n_1668)
);

OR2x2_ASAP7_75t_L g1669 ( 
.A(n_1631),
.B(n_1604),
.Y(n_1669)
);

NOR2xp33_ASAP7_75t_L g1670 ( 
.A(n_1628),
.B(n_1552),
.Y(n_1670)
);

INVx2_ASAP7_75t_L g1671 ( 
.A(n_1627),
.Y(n_1671)
);

AND2x2_ASAP7_75t_L g1672 ( 
.A(n_1638),
.B(n_1640),
.Y(n_1672)
);

BUFx2_ASAP7_75t_L g1673 ( 
.A(n_1626),
.Y(n_1673)
);

AND2x2_ASAP7_75t_L g1674 ( 
.A(n_1640),
.B(n_1624),
.Y(n_1674)
);

BUFx2_ASAP7_75t_L g1675 ( 
.A(n_1626),
.Y(n_1675)
);

AND2x4_ASAP7_75t_L g1676 ( 
.A(n_1626),
.B(n_1619),
.Y(n_1676)
);

AND2x2_ASAP7_75t_L g1677 ( 
.A(n_1640),
.B(n_1642),
.Y(n_1677)
);

BUFx2_ASAP7_75t_L g1678 ( 
.A(n_1641),
.Y(n_1678)
);

AND2x2_ASAP7_75t_SL g1679 ( 
.A(n_1653),
.B(n_1610),
.Y(n_1679)
);

AND2x2_ASAP7_75t_L g1680 ( 
.A(n_1642),
.B(n_1643),
.Y(n_1680)
);

NAND2xp5_ASAP7_75t_L g1681 ( 
.A(n_1651),
.B(n_1608),
.Y(n_1681)
);

NOR2xp33_ASAP7_75t_L g1682 ( 
.A(n_1639),
.B(n_1551),
.Y(n_1682)
);

AND2x2_ASAP7_75t_L g1683 ( 
.A(n_1642),
.B(n_1643),
.Y(n_1683)
);

BUFx2_ASAP7_75t_L g1684 ( 
.A(n_1641),
.Y(n_1684)
);

INVx2_ASAP7_75t_L g1685 ( 
.A(n_1627),
.Y(n_1685)
);

INVx1_ASAP7_75t_L g1686 ( 
.A(n_1664),
.Y(n_1686)
);

INVx1_ASAP7_75t_L g1687 ( 
.A(n_1664),
.Y(n_1687)
);

INVx3_ASAP7_75t_L g1688 ( 
.A(n_1654),
.Y(n_1688)
);

OR2x2_ASAP7_75t_L g1689 ( 
.A(n_1669),
.B(n_1636),
.Y(n_1689)
);

HB1xp67_ASAP7_75t_L g1690 ( 
.A(n_1678),
.Y(n_1690)
);

NAND2xp5_ASAP7_75t_L g1691 ( 
.A(n_1670),
.B(n_1651),
.Y(n_1691)
);

INVx2_ASAP7_75t_SL g1692 ( 
.A(n_1678),
.Y(n_1692)
);

INVx1_ASAP7_75t_L g1693 ( 
.A(n_1664),
.Y(n_1693)
);

AND2x2_ASAP7_75t_L g1694 ( 
.A(n_1680),
.B(n_1643),
.Y(n_1694)
);

INVx1_ASAP7_75t_L g1695 ( 
.A(n_1664),
.Y(n_1695)
);

INVx1_ASAP7_75t_L g1696 ( 
.A(n_1666),
.Y(n_1696)
);

HB1xp67_ASAP7_75t_L g1697 ( 
.A(n_1678),
.Y(n_1697)
);

NOR2xp33_ASAP7_75t_L g1698 ( 
.A(n_1670),
.B(n_1541),
.Y(n_1698)
);

INVx1_ASAP7_75t_L g1699 ( 
.A(n_1666),
.Y(n_1699)
);

INVx1_ASAP7_75t_L g1700 ( 
.A(n_1666),
.Y(n_1700)
);

NAND2xp5_ASAP7_75t_L g1701 ( 
.A(n_1660),
.B(n_1652),
.Y(n_1701)
);

INVx2_ASAP7_75t_L g1702 ( 
.A(n_1663),
.Y(n_1702)
);

AND2x2_ASAP7_75t_L g1703 ( 
.A(n_1680),
.B(n_1641),
.Y(n_1703)
);

AND2x2_ASAP7_75t_L g1704 ( 
.A(n_1680),
.B(n_1641),
.Y(n_1704)
);

AND2x2_ASAP7_75t_L g1705 ( 
.A(n_1683),
.B(n_1652),
.Y(n_1705)
);

AOI22xp5_ASAP7_75t_L g1706 ( 
.A1(n_1660),
.A2(n_1632),
.B1(n_1634),
.B2(n_1629),
.Y(n_1706)
);

NOR2xp33_ASAP7_75t_SL g1707 ( 
.A(n_1660),
.B(n_1650),
.Y(n_1707)
);

INVx2_ASAP7_75t_L g1708 ( 
.A(n_1663),
.Y(n_1708)
);

INVx1_ASAP7_75t_L g1709 ( 
.A(n_1666),
.Y(n_1709)
);

AOI22xp5_ASAP7_75t_L g1710 ( 
.A1(n_1682),
.A2(n_1632),
.B1(n_1634),
.B2(n_1629),
.Y(n_1710)
);

INVx3_ASAP7_75t_SL g1711 ( 
.A(n_1679),
.Y(n_1711)
);

NAND2xp5_ASAP7_75t_L g1712 ( 
.A(n_1684),
.B(n_1633),
.Y(n_1712)
);

OAI22xp33_ASAP7_75t_L g1713 ( 
.A1(n_1684),
.A2(n_1650),
.B1(n_1625),
.B2(n_1646),
.Y(n_1713)
);

INVx6_ASAP7_75t_L g1714 ( 
.A(n_1679),
.Y(n_1714)
);

AND2x2_ASAP7_75t_L g1715 ( 
.A(n_1683),
.B(n_1635),
.Y(n_1715)
);

AND2x4_ASAP7_75t_L g1716 ( 
.A(n_1684),
.B(n_1654),
.Y(n_1716)
);

INVx1_ASAP7_75t_L g1717 ( 
.A(n_1662),
.Y(n_1717)
);

INVx1_ASAP7_75t_L g1718 ( 
.A(n_1662),
.Y(n_1718)
);

NAND2xp5_ASAP7_75t_L g1719 ( 
.A(n_1681),
.B(n_1633),
.Y(n_1719)
);

OR2x2_ASAP7_75t_L g1720 ( 
.A(n_1669),
.B(n_1636),
.Y(n_1720)
);

AND2x2_ASAP7_75t_L g1721 ( 
.A(n_1683),
.B(n_1635),
.Y(n_1721)
);

INVx1_ASAP7_75t_L g1722 ( 
.A(n_1662),
.Y(n_1722)
);

AND2x2_ASAP7_75t_L g1723 ( 
.A(n_1679),
.B(n_1645),
.Y(n_1723)
);

INVx1_ASAP7_75t_SL g1724 ( 
.A(n_1679),
.Y(n_1724)
);

AND2x2_ASAP7_75t_L g1725 ( 
.A(n_1677),
.B(n_1645),
.Y(n_1725)
);

INVx1_ASAP7_75t_L g1726 ( 
.A(n_1665),
.Y(n_1726)
);

AND2x2_ASAP7_75t_L g1727 ( 
.A(n_1677),
.B(n_1645),
.Y(n_1727)
);

NAND2xp5_ASAP7_75t_L g1728 ( 
.A(n_1681),
.B(n_1647),
.Y(n_1728)
);

INVxp67_ASAP7_75t_L g1729 ( 
.A(n_1707),
.Y(n_1729)
);

NAND2xp5_ASAP7_75t_L g1730 ( 
.A(n_1710),
.B(n_1659),
.Y(n_1730)
);

INVx1_ASAP7_75t_SL g1731 ( 
.A(n_1711),
.Y(n_1731)
);

AND2x2_ASAP7_75t_L g1732 ( 
.A(n_1711),
.B(n_1677),
.Y(n_1732)
);

OR2x2_ASAP7_75t_L g1733 ( 
.A(n_1728),
.B(n_1701),
.Y(n_1733)
);

NAND2xp5_ASAP7_75t_L g1734 ( 
.A(n_1710),
.B(n_1659),
.Y(n_1734)
);

INVx1_ASAP7_75t_L g1735 ( 
.A(n_1690),
.Y(n_1735)
);

INVx1_ASAP7_75t_L g1736 ( 
.A(n_1697),
.Y(n_1736)
);

OR2x2_ASAP7_75t_L g1737 ( 
.A(n_1689),
.B(n_1669),
.Y(n_1737)
);

AND2x4_ASAP7_75t_L g1738 ( 
.A(n_1703),
.B(n_1654),
.Y(n_1738)
);

INVx1_ASAP7_75t_L g1739 ( 
.A(n_1717),
.Y(n_1739)
);

NAND2xp5_ASAP7_75t_L g1740 ( 
.A(n_1706),
.B(n_1659),
.Y(n_1740)
);

INVx1_ASAP7_75t_L g1741 ( 
.A(n_1692),
.Y(n_1741)
);

NOR2xp33_ASAP7_75t_L g1742 ( 
.A(n_1698),
.B(n_1682),
.Y(n_1742)
);

INVxp67_ASAP7_75t_L g1743 ( 
.A(n_1703),
.Y(n_1743)
);

NAND2xp5_ASAP7_75t_L g1744 ( 
.A(n_1719),
.B(n_1659),
.Y(n_1744)
);

INVx2_ASAP7_75t_SL g1745 ( 
.A(n_1692),
.Y(n_1745)
);

INVxp67_ASAP7_75t_L g1746 ( 
.A(n_1704),
.Y(n_1746)
);

HB1xp67_ASAP7_75t_L g1747 ( 
.A(n_1704),
.Y(n_1747)
);

NAND2xp5_ASAP7_75t_L g1748 ( 
.A(n_1712),
.B(n_1661),
.Y(n_1748)
);

NAND2xp5_ASAP7_75t_L g1749 ( 
.A(n_1691),
.B(n_1661),
.Y(n_1749)
);

HB1xp67_ASAP7_75t_L g1750 ( 
.A(n_1715),
.Y(n_1750)
);

AND2x2_ASAP7_75t_L g1751 ( 
.A(n_1711),
.B(n_1677),
.Y(n_1751)
);

INVx1_ASAP7_75t_L g1752 ( 
.A(n_1725),
.Y(n_1752)
);

HB1xp67_ASAP7_75t_L g1753 ( 
.A(n_1715),
.Y(n_1753)
);

INVx1_ASAP7_75t_L g1754 ( 
.A(n_1717),
.Y(n_1754)
);

NAND2xp5_ASAP7_75t_L g1755 ( 
.A(n_1713),
.B(n_1661),
.Y(n_1755)
);

NAND2xp5_ASAP7_75t_L g1756 ( 
.A(n_1705),
.B(n_1661),
.Y(n_1756)
);

INVx1_ASAP7_75t_L g1757 ( 
.A(n_1725),
.Y(n_1757)
);

NAND2xp5_ASAP7_75t_L g1758 ( 
.A(n_1705),
.B(n_1658),
.Y(n_1758)
);

AOI22xp33_ASAP7_75t_L g1759 ( 
.A1(n_1714),
.A2(n_1668),
.B1(n_1654),
.B2(n_1625),
.Y(n_1759)
);

NAND2xp5_ASAP7_75t_L g1760 ( 
.A(n_1723),
.B(n_1658),
.Y(n_1760)
);

OR2x2_ASAP7_75t_L g1761 ( 
.A(n_1689),
.B(n_1655),
.Y(n_1761)
);

AND2x2_ASAP7_75t_L g1762 ( 
.A(n_1694),
.B(n_1672),
.Y(n_1762)
);

INVx1_ASAP7_75t_L g1763 ( 
.A(n_1727),
.Y(n_1763)
);

INVx1_ASAP7_75t_L g1764 ( 
.A(n_1718),
.Y(n_1764)
);

OR2x2_ASAP7_75t_L g1765 ( 
.A(n_1720),
.B(n_1655),
.Y(n_1765)
);

OAI22xp5_ASAP7_75t_L g1766 ( 
.A1(n_1729),
.A2(n_1714),
.B1(n_1724),
.B2(n_1601),
.Y(n_1766)
);

AOI21xp33_ASAP7_75t_L g1767 ( 
.A1(n_1731),
.A2(n_1649),
.B(n_1716),
.Y(n_1767)
);

OAI22xp33_ASAP7_75t_L g1768 ( 
.A1(n_1730),
.A2(n_1646),
.B1(n_1714),
.B2(n_1656),
.Y(n_1768)
);

AOI22xp5_ASAP7_75t_L g1769 ( 
.A1(n_1742),
.A2(n_1714),
.B1(n_1716),
.B2(n_1668),
.Y(n_1769)
);

NAND2xp5_ASAP7_75t_L g1770 ( 
.A(n_1743),
.B(n_1723),
.Y(n_1770)
);

NAND2xp5_ASAP7_75t_L g1771 ( 
.A(n_1746),
.B(n_1716),
.Y(n_1771)
);

NAND3xp33_ASAP7_75t_L g1772 ( 
.A(n_1734),
.B(n_1649),
.C(n_1716),
.Y(n_1772)
);

NAND2xp5_ASAP7_75t_L g1773 ( 
.A(n_1747),
.B(n_1694),
.Y(n_1773)
);

OAI22xp33_ASAP7_75t_SL g1774 ( 
.A1(n_1755),
.A2(n_1688),
.B1(n_1656),
.B2(n_1720),
.Y(n_1774)
);

INVx1_ASAP7_75t_L g1775 ( 
.A(n_1739),
.Y(n_1775)
);

OAI21xp5_ASAP7_75t_L g1776 ( 
.A1(n_1740),
.A2(n_1668),
.B(n_1654),
.Y(n_1776)
);

OAI21xp33_ASAP7_75t_L g1777 ( 
.A1(n_1744),
.A2(n_1748),
.B(n_1732),
.Y(n_1777)
);

OAI22xp33_ASAP7_75t_L g1778 ( 
.A1(n_1760),
.A2(n_1756),
.B1(n_1750),
.B2(n_1753),
.Y(n_1778)
);

AOI22xp5_ASAP7_75t_L g1779 ( 
.A1(n_1732),
.A2(n_1668),
.B1(n_1654),
.B2(n_1653),
.Y(n_1779)
);

OAI22xp5_ASAP7_75t_L g1780 ( 
.A1(n_1759),
.A2(n_1688),
.B1(n_1668),
.B2(n_1727),
.Y(n_1780)
);

NOR2xp33_ASAP7_75t_L g1781 ( 
.A(n_1733),
.B(n_1579),
.Y(n_1781)
);

INVx1_ASAP7_75t_L g1782 ( 
.A(n_1739),
.Y(n_1782)
);

INVx2_ASAP7_75t_L g1783 ( 
.A(n_1738),
.Y(n_1783)
);

INVx1_ASAP7_75t_L g1784 ( 
.A(n_1754),
.Y(n_1784)
);

OAI21xp33_ASAP7_75t_L g1785 ( 
.A1(n_1751),
.A2(n_1721),
.B(n_1708),
.Y(n_1785)
);

OAI21xp5_ASAP7_75t_L g1786 ( 
.A1(n_1751),
.A2(n_1668),
.B(n_1688),
.Y(n_1786)
);

AOI222xp33_ASAP7_75t_L g1787 ( 
.A1(n_1735),
.A2(n_1721),
.B1(n_1503),
.B2(n_1637),
.C1(n_1675),
.C2(n_1673),
.Y(n_1787)
);

INVxp67_ASAP7_75t_L g1788 ( 
.A(n_1745),
.Y(n_1788)
);

NAND2xp5_ASAP7_75t_L g1789 ( 
.A(n_1736),
.B(n_1658),
.Y(n_1789)
);

AOI221x1_ASAP7_75t_L g1790 ( 
.A1(n_1736),
.A2(n_1687),
.B1(n_1695),
.B2(n_1696),
.C(n_1709),
.Y(n_1790)
);

AOI221xp5_ASAP7_75t_L g1791 ( 
.A1(n_1741),
.A2(n_1693),
.B1(n_1686),
.B2(n_1687),
.C(n_1709),
.Y(n_1791)
);

OAI31xp33_ASAP7_75t_L g1792 ( 
.A1(n_1768),
.A2(n_1733),
.A3(n_1745),
.B(n_1738),
.Y(n_1792)
);

AOI21xp33_ASAP7_75t_L g1793 ( 
.A1(n_1768),
.A2(n_1778),
.B(n_1774),
.Y(n_1793)
);

OAI21xp5_ASAP7_75t_L g1794 ( 
.A1(n_1772),
.A2(n_1738),
.B(n_1749),
.Y(n_1794)
);

OAI21xp5_ASAP7_75t_L g1795 ( 
.A1(n_1766),
.A2(n_1769),
.B(n_1790),
.Y(n_1795)
);

INVxp67_ASAP7_75t_SL g1796 ( 
.A(n_1788),
.Y(n_1796)
);

AOI21xp33_ASAP7_75t_L g1797 ( 
.A1(n_1781),
.A2(n_1765),
.B(n_1761),
.Y(n_1797)
);

NAND3xp33_ASAP7_75t_L g1798 ( 
.A(n_1767),
.B(n_1765),
.C(n_1761),
.Y(n_1798)
);

INVx1_ASAP7_75t_L g1799 ( 
.A(n_1775),
.Y(n_1799)
);

OAI21xp5_ASAP7_75t_L g1800 ( 
.A1(n_1788),
.A2(n_1758),
.B(n_1757),
.Y(n_1800)
);

AOI22xp5_ASAP7_75t_L g1801 ( 
.A1(n_1777),
.A2(n_1752),
.B1(n_1763),
.B2(n_1762),
.Y(n_1801)
);

INVxp67_ASAP7_75t_L g1802 ( 
.A(n_1771),
.Y(n_1802)
);

NAND2xp5_ASAP7_75t_L g1803 ( 
.A(n_1783),
.B(n_1762),
.Y(n_1803)
);

AND2x4_ASAP7_75t_L g1804 ( 
.A(n_1786),
.B(n_1609),
.Y(n_1804)
);

AND2x2_ASAP7_75t_L g1805 ( 
.A(n_1776),
.B(n_1658),
.Y(n_1805)
);

NAND2xp5_ASAP7_75t_SL g1806 ( 
.A(n_1787),
.B(n_1737),
.Y(n_1806)
);

INVx2_ASAP7_75t_L g1807 ( 
.A(n_1773),
.Y(n_1807)
);

NAND4xp25_ASAP7_75t_SL g1808 ( 
.A(n_1779),
.B(n_1737),
.C(n_1708),
.D(n_1702),
.Y(n_1808)
);

NAND4xp25_ASAP7_75t_L g1809 ( 
.A(n_1770),
.B(n_1780),
.C(n_1785),
.D(n_1791),
.Y(n_1809)
);

NAND2xp5_ASAP7_75t_L g1810 ( 
.A(n_1782),
.B(n_1674),
.Y(n_1810)
);

HB1xp67_ASAP7_75t_L g1811 ( 
.A(n_1784),
.Y(n_1811)
);

OAI221xp5_ASAP7_75t_L g1812 ( 
.A1(n_1795),
.A2(n_1789),
.B1(n_1673),
.B2(n_1675),
.C(n_1764),
.Y(n_1812)
);

NAND2xp5_ASAP7_75t_L g1813 ( 
.A(n_1796),
.B(n_1672),
.Y(n_1813)
);

OAI21xp5_ASAP7_75t_SL g1814 ( 
.A1(n_1793),
.A2(n_1653),
.B(n_1563),
.Y(n_1814)
);

INVx1_ASAP7_75t_L g1815 ( 
.A(n_1796),
.Y(n_1815)
);

OR2x2_ASAP7_75t_L g1816 ( 
.A(n_1803),
.B(n_1702),
.Y(n_1816)
);

AOI22xp33_ASAP7_75t_L g1817 ( 
.A1(n_1792),
.A2(n_1764),
.B1(n_1754),
.B2(n_1540),
.Y(n_1817)
);

INVx1_ASAP7_75t_SL g1818 ( 
.A(n_1804),
.Y(n_1818)
);

INVx1_ASAP7_75t_SL g1819 ( 
.A(n_1804),
.Y(n_1819)
);

NAND2xp5_ASAP7_75t_L g1820 ( 
.A(n_1802),
.B(n_1672),
.Y(n_1820)
);

INVx1_ASAP7_75t_L g1821 ( 
.A(n_1811),
.Y(n_1821)
);

NAND3xp33_ASAP7_75t_SL g1822 ( 
.A(n_1794),
.B(n_1675),
.C(n_1673),
.Y(n_1822)
);

NAND2xp5_ASAP7_75t_SL g1823 ( 
.A(n_1797),
.B(n_1653),
.Y(n_1823)
);

NOR5xp2_ASAP7_75t_L g1824 ( 
.A(n_1812),
.B(n_1811),
.C(n_1798),
.D(n_1802),
.E(n_1809),
.Y(n_1824)
);

O2A1O1Ixp5_ASAP7_75t_L g1825 ( 
.A1(n_1815),
.A2(n_1806),
.B(n_1800),
.C(n_1807),
.Y(n_1825)
);

O2A1O1Ixp5_ASAP7_75t_SL g1826 ( 
.A1(n_1821),
.A2(n_1799),
.B(n_1810),
.C(n_1722),
.Y(n_1826)
);

NAND3xp33_ASAP7_75t_L g1827 ( 
.A(n_1817),
.B(n_1801),
.C(n_1805),
.Y(n_1827)
);

NOR2xp33_ASAP7_75t_L g1828 ( 
.A(n_1818),
.B(n_1808),
.Y(n_1828)
);

NAND2xp5_ASAP7_75t_L g1829 ( 
.A(n_1819),
.B(n_1674),
.Y(n_1829)
);

OAI211xp5_ASAP7_75t_SL g1830 ( 
.A1(n_1814),
.A2(n_1538),
.B(n_1542),
.C(n_1686),
.Y(n_1830)
);

NAND2xp5_ASAP7_75t_L g1831 ( 
.A(n_1817),
.B(n_1674),
.Y(n_1831)
);

NAND3xp33_ASAP7_75t_L g1832 ( 
.A(n_1813),
.B(n_1722),
.C(n_1718),
.Y(n_1832)
);

AND2x2_ASAP7_75t_SL g1833 ( 
.A(n_1820),
.B(n_1464),
.Y(n_1833)
);

AOI21xp5_ASAP7_75t_L g1834 ( 
.A1(n_1825),
.A2(n_1827),
.B(n_1822),
.Y(n_1834)
);

O2A1O1Ixp5_ASAP7_75t_L g1835 ( 
.A1(n_1828),
.A2(n_1823),
.B(n_1816),
.C(n_1726),
.Y(n_1835)
);

AOI21xp5_ASAP7_75t_L g1836 ( 
.A1(n_1833),
.A2(n_1507),
.B(n_1504),
.Y(n_1836)
);

OAI32xp33_ASAP7_75t_L g1837 ( 
.A1(n_1824),
.A2(n_1700),
.A3(n_1699),
.B1(n_1693),
.B2(n_1696),
.Y(n_1837)
);

NOR3x1_ASAP7_75t_L g1838 ( 
.A(n_1829),
.B(n_1699),
.C(n_1695),
.Y(n_1838)
);

NAND4xp25_ASAP7_75t_L g1839 ( 
.A(n_1830),
.B(n_1504),
.C(n_1543),
.D(n_1563),
.Y(n_1839)
);

NAND2xp5_ASAP7_75t_L g1840 ( 
.A(n_1831),
.B(n_1700),
.Y(n_1840)
);

OAI21xp33_ASAP7_75t_L g1841 ( 
.A1(n_1839),
.A2(n_1826),
.B(n_1832),
.Y(n_1841)
);

OAI21xp33_ASAP7_75t_L g1842 ( 
.A1(n_1834),
.A2(n_1726),
.B(n_1593),
.Y(n_1842)
);

OAI221xp5_ASAP7_75t_L g1843 ( 
.A1(n_1835),
.A2(n_1545),
.B1(n_1567),
.B2(n_1639),
.C(n_1555),
.Y(n_1843)
);

AOI21xp5_ASAP7_75t_L g1844 ( 
.A1(n_1837),
.A2(n_1543),
.B(n_1685),
.Y(n_1844)
);

OAI211xp5_ASAP7_75t_SL g1845 ( 
.A1(n_1836),
.A2(n_1840),
.B(n_1838),
.C(n_1558),
.Y(n_1845)
);

AOI22xp33_ASAP7_75t_L g1846 ( 
.A1(n_1834),
.A2(n_1653),
.B1(n_1561),
.B2(n_1571),
.Y(n_1846)
);

OAI211xp5_ASAP7_75t_SL g1847 ( 
.A1(n_1834),
.A2(n_1611),
.B(n_1602),
.C(n_1657),
.Y(n_1847)
);

NOR3xp33_ASAP7_75t_L g1848 ( 
.A(n_1842),
.B(n_1841),
.C(n_1845),
.Y(n_1848)
);

INVx2_ASAP7_75t_SL g1849 ( 
.A(n_1847),
.Y(n_1849)
);

NOR2x1_ASAP7_75t_L g1850 ( 
.A(n_1843),
.B(n_1657),
.Y(n_1850)
);

INVx1_ASAP7_75t_L g1851 ( 
.A(n_1846),
.Y(n_1851)
);

AO22x2_ASAP7_75t_L g1852 ( 
.A1(n_1844),
.A2(n_1685),
.B1(n_1671),
.B2(n_1667),
.Y(n_1852)
);

OAI211xp5_ASAP7_75t_SL g1853 ( 
.A1(n_1851),
.A2(n_1559),
.B(n_1685),
.C(n_1657),
.Y(n_1853)
);

NOR2x1p5_ASAP7_75t_L g1854 ( 
.A(n_1848),
.B(n_1529),
.Y(n_1854)
);

OAI21xp5_ASAP7_75t_L g1855 ( 
.A1(n_1849),
.A2(n_1676),
.B(n_1674),
.Y(n_1855)
);

INVx1_ASAP7_75t_L g1856 ( 
.A(n_1854),
.Y(n_1856)
);

INVx1_ASAP7_75t_L g1857 ( 
.A(n_1856),
.Y(n_1857)
);

OAI22xp5_ASAP7_75t_L g1858 ( 
.A1(n_1857),
.A2(n_1850),
.B1(n_1855),
.B2(n_1852),
.Y(n_1858)
);

OAI22xp5_ASAP7_75t_SL g1859 ( 
.A1(n_1857),
.A2(n_1853),
.B1(n_1456),
.B2(n_1529),
.Y(n_1859)
);

INVx1_ASAP7_75t_L g1860 ( 
.A(n_1858),
.Y(n_1860)
);

AND2x4_ASAP7_75t_L g1861 ( 
.A(n_1859),
.B(n_1676),
.Y(n_1861)
);

INVx2_ASAP7_75t_L g1862 ( 
.A(n_1861),
.Y(n_1862)
);

INVx1_ASAP7_75t_L g1863 ( 
.A(n_1860),
.Y(n_1863)
);

INVx1_ASAP7_75t_L g1864 ( 
.A(n_1863),
.Y(n_1864)
);

OAI21xp5_ASAP7_75t_SL g1865 ( 
.A1(n_1864),
.A2(n_1862),
.B(n_1553),
.Y(n_1865)
);

OAI222xp33_ASAP7_75t_L g1866 ( 
.A1(n_1865),
.A2(n_1685),
.B1(n_1657),
.B2(n_1667),
.C1(n_1671),
.C2(n_1648),
.Y(n_1866)
);

OAI221xp5_ASAP7_75t_R g1867 ( 
.A1(n_1866),
.A2(n_1557),
.B1(n_1667),
.B2(n_1671),
.C(n_1648),
.Y(n_1867)
);

AOI211xp5_ASAP7_75t_L g1868 ( 
.A1(n_1867),
.A2(n_1522),
.B(n_1580),
.C(n_1520),
.Y(n_1868)
);


endmodule