module fake_jpeg_21504_n_152 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_152);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_152;

wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_51;
wire n_147;
wire n_73;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_150;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_138;
wire n_101;
wire n_149;
wire n_87;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_135;
wire n_62;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_39),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_24),
.Y(n_50)
);

CKINVDCx14_ASAP7_75t_R g51 ( 
.A(n_19),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_28),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_32),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_25),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_15),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_0),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_33),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_48),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_37),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_1),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_44),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_41),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_11),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_20),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_34),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_12),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_30),
.Y(n_67)
);

BUFx16f_ASAP7_75t_L g68 ( 
.A(n_14),
.Y(n_68)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_40),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_6),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_38),
.Y(n_71)
);

BUFx10_ASAP7_75t_L g72 ( 
.A(n_18),
.Y(n_72)
);

BUFx2_ASAP7_75t_L g73 ( 
.A(n_0),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_2),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_17),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_27),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_50),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_77),
.B(n_79),
.Y(n_93)
);

BUFx12f_ASAP7_75t_L g78 ( 
.A(n_63),
.Y(n_78)
);

BUFx2_ASAP7_75t_L g94 ( 
.A(n_78),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_52),
.Y(n_79)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_69),
.Y(n_80)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_80),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_55),
.Y(n_81)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_81),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_55),
.Y(n_82)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_82),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_76),
.Y(n_83)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_83),
.Y(n_91)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_73),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_84),
.A2(n_72),
.B1(n_68),
.B2(n_75),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_L g85 ( 
.A1(n_80),
.A2(n_51),
.B1(n_73),
.B2(n_65),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_85),
.A2(n_89),
.B1(n_90),
.B2(n_92),
.Y(n_108)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_88),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_81),
.A2(n_72),
.B1(n_54),
.B2(n_57),
.Y(n_89)
);

OAI22xp33_ASAP7_75t_L g90 ( 
.A1(n_82),
.A2(n_51),
.B1(n_72),
.B2(n_75),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_78),
.A2(n_62),
.B1(n_71),
.B2(n_59),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_91),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_96),
.B(n_101),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_93),
.B(n_74),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_97),
.B(n_103),
.Y(n_122)
);

BUFx3_ASAP7_75t_L g99 ( 
.A(n_94),
.Y(n_99)
);

O2A1O1Ixp33_ASAP7_75t_L g100 ( 
.A1(n_87),
.A2(n_78),
.B(n_49),
.C(n_61),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_100),
.A2(n_102),
.B1(n_106),
.B2(n_3),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_89),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_88),
.A2(n_53),
.B1(n_64),
.B2(n_66),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_86),
.B(n_56),
.Y(n_103)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_95),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_104),
.B(n_3),
.Y(n_116)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_94),
.Y(n_105)
);

INVx6_ASAP7_75t_L g109 ( 
.A(n_105),
.Y(n_109)
);

OAI22xp33_ASAP7_75t_L g106 ( 
.A1(n_95),
.A2(n_65),
.B1(n_58),
.B2(n_68),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_92),
.B(n_60),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_SL g113 ( 
.A(n_107),
.B(n_1),
.Y(n_113)
);

CKINVDCx12_ASAP7_75t_R g111 ( 
.A(n_99),
.Y(n_111)
);

INVxp67_ASAP7_75t_L g128 ( 
.A(n_111),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_98),
.A2(n_70),
.B1(n_58),
.B2(n_67),
.Y(n_112)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_112),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_113),
.B(n_114),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_108),
.B(n_22),
.C(n_46),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_104),
.B(n_2),
.Y(n_115)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_115),
.Y(n_127)
);

CKINVDCx16_ASAP7_75t_R g131 ( 
.A(n_116),
.Y(n_131)
);

AND2x6_ASAP7_75t_L g117 ( 
.A(n_100),
.B(n_21),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_117),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_106),
.B(n_23),
.C(n_45),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_118),
.A2(n_4),
.B1(n_5),
.B2(n_7),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_96),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_119),
.Y(n_124)
);

XOR2xp5_ASAP7_75t_L g120 ( 
.A(n_108),
.B(n_16),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_120),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_121),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_126),
.A2(n_109),
.B1(n_8),
.B2(n_9),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_111),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_132),
.B(n_133),
.Y(n_139)
);

XOR2xp5_ASAP7_75t_L g134 ( 
.A(n_130),
.B(n_110),
.Y(n_134)
);

XNOR2xp5_ASAP7_75t_L g141 ( 
.A(n_134),
.B(n_136),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_124),
.B(n_110),
.Y(n_135)
);

INVxp67_ASAP7_75t_L g140 ( 
.A(n_135),
.Y(n_140)
);

AOI21xp5_ASAP7_75t_SL g136 ( 
.A1(n_127),
.A2(n_115),
.B(n_122),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_128),
.Y(n_137)
);

AOI21xp5_ASAP7_75t_L g142 ( 
.A1(n_140),
.A2(n_135),
.B(n_137),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_142),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_143),
.B(n_131),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_144),
.B(n_139),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_SL g146 ( 
.A1(n_145),
.A2(n_123),
.B(n_128),
.Y(n_146)
);

HB1xp67_ASAP7_75t_L g147 ( 
.A(n_146),
.Y(n_147)
);

AOI322xp5_ASAP7_75t_L g148 ( 
.A1(n_147),
.A2(n_141),
.A3(n_129),
.B1(n_126),
.B2(n_138),
.C1(n_13),
.C2(n_26),
.Y(n_148)
);

AOI322xp5_ASAP7_75t_L g149 ( 
.A1(n_148),
.A2(n_129),
.A3(n_36),
.B1(n_42),
.B2(n_10),
.C1(n_29),
.C2(n_31),
.Y(n_149)
);

AOI21xp5_ASAP7_75t_L g150 ( 
.A1(n_149),
.A2(n_43),
.B(n_47),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_150),
.B(n_35),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_L g152 ( 
.A(n_151),
.B(n_125),
.Y(n_152)
);


endmodule