module fake_jpeg_2925_n_497 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_497);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_497;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_490;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_12),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_16),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_3),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

BUFx24_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_17),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_17),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_15),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_16),
.Y(n_33)
);

BUFx6f_ASAP7_75t_SL g34 ( 
.A(n_3),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_15),
.Y(n_35)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

BUFx10_ASAP7_75t_L g37 ( 
.A(n_1),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_13),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_17),
.Y(n_39)
);

BUFx5_ASAP7_75t_L g40 ( 
.A(n_4),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_8),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_3),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_SL g43 ( 
.A(n_5),
.B(n_10),
.Y(n_43)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_8),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_8),
.Y(n_45)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_14),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_8),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_2),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_12),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_7),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_12),
.Y(n_51)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_2),
.Y(n_52)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_10),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_5),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_5),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_7),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_43),
.B(n_18),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_57),
.B(n_69),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g58 ( 
.A(n_18),
.B(n_14),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_58),
.B(n_66),
.Y(n_122)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_52),
.Y(n_59)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_59),
.Y(n_127)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_27),
.Y(n_60)
);

BUFx2_ASAP7_75t_L g175 ( 
.A(n_60),
.Y(n_175)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_24),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g142 ( 
.A(n_61),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_24),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g148 ( 
.A(n_62),
.Y(n_148)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_26),
.Y(n_63)
);

INVx5_ASAP7_75t_L g138 ( 
.A(n_63),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_24),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g152 ( 
.A(n_64),
.Y(n_152)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_52),
.Y(n_65)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_65),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_SL g66 ( 
.A(n_32),
.B(n_13),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_41),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g156 ( 
.A(n_67),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_41),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g157 ( 
.A(n_68),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_43),
.B(n_0),
.Y(n_69)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_53),
.Y(n_70)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_70),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_41),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g171 ( 
.A(n_71),
.Y(n_171)
);

INVx11_ASAP7_75t_L g72 ( 
.A(n_23),
.Y(n_72)
);

INVx11_ASAP7_75t_L g143 ( 
.A(n_72),
.Y(n_143)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_53),
.Y(n_73)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_73),
.Y(n_176)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_46),
.Y(n_74)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_74),
.Y(n_182)
);

INVx5_ASAP7_75t_L g75 ( 
.A(n_44),
.Y(n_75)
);

BUFx2_ASAP7_75t_L g190 ( 
.A(n_75),
.Y(n_190)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_55),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g180 ( 
.A(n_76),
.Y(n_180)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_55),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g183 ( 
.A(n_77),
.Y(n_183)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_55),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g187 ( 
.A(n_78),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_32),
.B(n_0),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_79),
.B(n_93),
.Y(n_167)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_26),
.Y(n_80)
);

INVx2_ASAP7_75t_SL g174 ( 
.A(n_80),
.Y(n_174)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_28),
.Y(n_81)
);

INVx6_ASAP7_75t_L g132 ( 
.A(n_81),
.Y(n_132)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_46),
.Y(n_82)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_82),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_28),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_83),
.B(n_99),
.Y(n_124)
);

BUFx3_ASAP7_75t_L g84 ( 
.A(n_27),
.Y(n_84)
);

INVx4_ASAP7_75t_L g135 ( 
.A(n_84),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_28),
.Y(n_85)
);

INVx6_ASAP7_75t_L g145 ( 
.A(n_85),
.Y(n_145)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_22),
.Y(n_86)
);

INVx3_ASAP7_75t_L g194 ( 
.A(n_86),
.Y(n_194)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_20),
.Y(n_87)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_87),
.Y(n_121)
);

BUFx5_ASAP7_75t_L g88 ( 
.A(n_23),
.Y(n_88)
);

INVx4_ASAP7_75t_L g149 ( 
.A(n_88),
.Y(n_149)
);

INVx5_ASAP7_75t_L g89 ( 
.A(n_44),
.Y(n_89)
);

INVx4_ASAP7_75t_L g168 ( 
.A(n_89),
.Y(n_168)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_26),
.Y(n_90)
);

INVx1_ASAP7_75t_SL g139 ( 
.A(n_90),
.Y(n_139)
);

INVx11_ASAP7_75t_L g91 ( 
.A(n_23),
.Y(n_91)
);

CKINVDCx16_ASAP7_75t_R g153 ( 
.A(n_91),
.Y(n_153)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_19),
.Y(n_92)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_92),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_35),
.B(n_0),
.Y(n_93)
);

AND2x2_ASAP7_75t_SL g94 ( 
.A(n_26),
.B(n_0),
.Y(n_94)
);

AND2x2_ASAP7_75t_L g126 ( 
.A(n_94),
.B(n_114),
.Y(n_126)
);

BUFx12f_ASAP7_75t_L g95 ( 
.A(n_44),
.Y(n_95)
);

INVx8_ASAP7_75t_L g146 ( 
.A(n_95),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_35),
.B(n_1),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_96),
.B(n_98),
.Y(n_177)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_29),
.Y(n_97)
);

BUFx12f_ASAP7_75t_L g154 ( 
.A(n_97),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_39),
.B(n_1),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g99 ( 
.A(n_39),
.B(n_1),
.Y(n_99)
);

INVx5_ASAP7_75t_L g100 ( 
.A(n_36),
.Y(n_100)
);

INVx3_ASAP7_75t_L g125 ( 
.A(n_100),
.Y(n_125)
);

BUFx5_ASAP7_75t_L g101 ( 
.A(n_23),
.Y(n_101)
);

BUFx12f_ASAP7_75t_L g155 ( 
.A(n_101),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_29),
.Y(n_102)
);

BUFx12f_ASAP7_75t_L g161 ( 
.A(n_102),
.Y(n_161)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_27),
.Y(n_103)
);

HB1xp67_ASAP7_75t_L g185 ( 
.A(n_103),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_29),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_104),
.B(n_117),
.Y(n_131)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_42),
.Y(n_105)
);

HB1xp67_ASAP7_75t_L g186 ( 
.A(n_105),
.Y(n_186)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_42),
.Y(n_106)
);

INVx3_ASAP7_75t_L g178 ( 
.A(n_106),
.Y(n_178)
);

INVx8_ASAP7_75t_L g107 ( 
.A(n_30),
.Y(n_107)
);

INVx3_ASAP7_75t_L g193 ( 
.A(n_107),
.Y(n_193)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_22),
.Y(n_108)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_108),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_30),
.Y(n_109)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_109),
.Y(n_147)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_20),
.Y(n_110)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_110),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_30),
.Y(n_111)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_111),
.Y(n_165)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_25),
.Y(n_112)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_112),
.Y(n_184)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_33),
.Y(n_113)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_113),
.Y(n_195)
);

INVx5_ASAP7_75t_L g114 ( 
.A(n_42),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_33),
.Y(n_115)
);

AND2x2_ASAP7_75t_L g170 ( 
.A(n_115),
.B(n_118),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_49),
.B(n_2),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_SL g140 ( 
.A(n_116),
.B(n_50),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_SL g117 ( 
.A(n_49),
.B(n_2),
.Y(n_117)
);

INVx8_ASAP7_75t_L g118 ( 
.A(n_33),
.Y(n_118)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_25),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_119),
.B(n_19),
.Y(n_144)
);

INVx4_ASAP7_75t_L g120 ( 
.A(n_40),
.Y(n_120)
);

AND2x2_ASAP7_75t_L g189 ( 
.A(n_120),
.B(n_75),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_94),
.A2(n_36),
.B1(n_51),
.B2(n_38),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_123),
.A2(n_197),
.B1(n_153),
.B2(n_125),
.Y(n_240)
);

AOI22xp33_ASAP7_75t_L g129 ( 
.A1(n_61),
.A2(n_34),
.B1(n_45),
.B2(n_31),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g249 ( 
.A1(n_129),
.A2(n_137),
.B1(n_158),
.B2(n_173),
.Y(n_249)
);

AOI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_86),
.A2(n_34),
.B1(n_56),
.B2(n_36),
.Y(n_130)
);

OA22x2_ASAP7_75t_L g241 ( 
.A1(n_130),
.A2(n_151),
.B1(n_181),
.B2(n_149),
.Y(n_241)
);

AOI21xp33_ASAP7_75t_SL g134 ( 
.A1(n_60),
.A2(n_56),
.B(n_38),
.Y(n_134)
);

OAI21xp33_ASAP7_75t_L g257 ( 
.A1(n_134),
.A2(n_156),
.B(n_157),
.Y(n_257)
);

OR2x2_ASAP7_75t_L g136 ( 
.A(n_108),
.B(n_51),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_136),
.B(n_140),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_81),
.A2(n_56),
.B1(n_31),
.B2(n_45),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_85),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_SL g226 ( 
.A(n_141),
.B(n_159),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_144),
.B(n_172),
.Y(n_200)
);

OA22x2_ASAP7_75t_L g151 ( 
.A1(n_120),
.A2(n_37),
.B1(n_40),
.B2(n_54),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g158 ( 
.A1(n_97),
.A2(n_54),
.B1(n_50),
.B2(n_48),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_63),
.B(n_48),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_102),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_SL g227 ( 
.A(n_162),
.B(n_164),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_84),
.B(n_47),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_114),
.B(n_47),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_SL g239 ( 
.A(n_166),
.B(n_169),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_109),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_L g172 ( 
.A1(n_107),
.A2(n_21),
.B(n_37),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_L g173 ( 
.A1(n_62),
.A2(n_21),
.B1(n_37),
.B2(n_6),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_95),
.B(n_4),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_179),
.B(n_188),
.Y(n_211)
);

AOI22xp33_ASAP7_75t_SL g181 ( 
.A1(n_72),
.A2(n_37),
.B1(n_5),
.B2(n_6),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_95),
.B(n_4),
.Y(n_188)
);

INVxp67_ASAP7_75t_L g221 ( 
.A(n_189),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_111),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_196),
.B(n_170),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_113),
.A2(n_37),
.B1(n_7),
.B2(n_9),
.Y(n_197)
);

AOI22xp33_ASAP7_75t_SL g198 ( 
.A1(n_189),
.A2(n_91),
.B1(n_89),
.B2(n_118),
.Y(n_198)
);

INVxp67_ASAP7_75t_L g303 ( 
.A(n_198),
.Y(n_303)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_147),
.Y(n_199)
);

INVx2_ASAP7_75t_L g281 ( 
.A(n_199),
.Y(n_281)
);

AOI22xp33_ASAP7_75t_SL g201 ( 
.A1(n_126),
.A2(n_67),
.B1(n_78),
.B2(n_77),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_L g263 ( 
.A1(n_201),
.A2(n_230),
.B1(n_232),
.B2(n_236),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_185),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g265 ( 
.A(n_202),
.B(n_204),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_126),
.A2(n_64),
.B1(n_76),
.B2(n_71),
.Y(n_203)
);

CKINVDCx16_ASAP7_75t_R g270 ( 
.A(n_203),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_186),
.Y(n_204)
);

INVx3_ASAP7_75t_L g205 ( 
.A(n_138),
.Y(n_205)
);

INVx4_ASAP7_75t_L g299 ( 
.A(n_205),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_175),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g300 ( 
.A(n_206),
.B(n_214),
.Y(n_300)
);

FAx1_ASAP7_75t_SL g207 ( 
.A(n_167),
.B(n_6),
.CI(n_7),
.CON(n_207),
.SN(n_207)
);

XNOR2xp5_ASAP7_75t_L g301 ( 
.A(n_207),
.B(n_217),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_124),
.B(n_68),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_208),
.B(n_213),
.Y(n_268)
);

BUFx3_ASAP7_75t_L g209 ( 
.A(n_138),
.Y(n_209)
);

INVx3_ASAP7_75t_L g276 ( 
.A(n_209),
.Y(n_276)
);

BUFx6f_ASAP7_75t_L g210 ( 
.A(n_142),
.Y(n_210)
);

INVx2_ASAP7_75t_SL g297 ( 
.A(n_210),
.Y(n_297)
);

INVx3_ASAP7_75t_L g212 ( 
.A(n_146),
.Y(n_212)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_212),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_131),
.B(n_115),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_175),
.Y(n_214)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_192),
.Y(n_216)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_216),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_177),
.A2(n_6),
.B1(n_9),
.B2(n_10),
.Y(n_217)
);

OAI22xp33_ASAP7_75t_SL g264 ( 
.A1(n_217),
.A2(n_225),
.B1(n_254),
.B2(n_180),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_190),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_SL g309 ( 
.A(n_218),
.B(n_224),
.Y(n_309)
);

BUFx3_ASAP7_75t_L g219 ( 
.A(n_146),
.Y(n_219)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_219),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_121),
.B(n_10),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_220),
.B(n_234),
.Y(n_277)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_165),
.Y(n_222)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_222),
.Y(n_274)
);

INVx3_ASAP7_75t_SL g223 ( 
.A(n_135),
.Y(n_223)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_223),
.Y(n_284)
);

A2O1A1Ixp33_ASAP7_75t_L g224 ( 
.A1(n_128),
.A2(n_11),
.B(n_122),
.C(n_136),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_151),
.A2(n_11),
.B1(n_170),
.B2(n_130),
.Y(n_225)
);

CKINVDCx14_ASAP7_75t_R g282 ( 
.A(n_228),
.Y(n_282)
);

INVx4_ASAP7_75t_L g229 ( 
.A(n_168),
.Y(n_229)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_229),
.Y(n_307)
);

AOI22xp33_ASAP7_75t_SL g230 ( 
.A1(n_151),
.A2(n_194),
.B1(n_133),
.B2(n_178),
.Y(n_230)
);

INVxp67_ASAP7_75t_L g231 ( 
.A(n_178),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_231),
.B(n_244),
.Y(n_285)
);

AOI22xp33_ASAP7_75t_SL g232 ( 
.A1(n_125),
.A2(n_139),
.B1(n_190),
.B2(n_149),
.Y(n_232)
);

AND2x2_ASAP7_75t_SL g233 ( 
.A(n_127),
.B(n_160),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_233),
.B(n_247),
.C(n_262),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_163),
.B(n_184),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_195),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_235),
.B(n_237),
.Y(n_280)
);

AOI22xp33_ASAP7_75t_L g236 ( 
.A1(n_129),
.A2(n_173),
.B1(n_150),
.B2(n_176),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_193),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_182),
.B(n_191),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_238),
.B(n_242),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_240),
.A2(n_249),
.B1(n_221),
.B2(n_242),
.Y(n_272)
);

A2O1A1Ixp33_ASAP7_75t_SL g286 ( 
.A1(n_241),
.A2(n_257),
.B(n_245),
.C(n_256),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_193),
.B(n_135),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_168),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_243),
.B(n_251),
.Y(n_294)
);

INVx3_ASAP7_75t_L g244 ( 
.A(n_139),
.Y(n_244)
);

O2A1O1Ixp33_ASAP7_75t_L g245 ( 
.A1(n_181),
.A2(n_143),
.B(n_155),
.C(n_174),
.Y(n_245)
);

AOI21xp5_ASAP7_75t_L g306 ( 
.A1(n_245),
.A2(n_205),
.B(n_241),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_132),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_246),
.B(n_248),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_SL g247 ( 
.A(n_174),
.B(n_155),
.Y(n_247)
);

INVx3_ASAP7_75t_L g248 ( 
.A(n_154),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_154),
.B(n_161),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_250),
.B(n_253),
.Y(n_293)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_132),
.Y(n_251)
);

AOI22xp33_ASAP7_75t_SL g252 ( 
.A1(n_155),
.A2(n_143),
.B1(n_161),
.B2(n_154),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_252),
.A2(n_218),
.B1(n_214),
.B2(n_206),
.Y(n_289)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_145),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_142),
.A2(n_187),
.B1(n_148),
.B2(n_152),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_161),
.B(n_145),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_255),
.B(n_256),
.Y(n_296)
);

NOR2x1_ASAP7_75t_L g256 ( 
.A(n_148),
.B(n_152),
.Y(n_256)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_156),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_258),
.B(n_260),
.Y(n_298)
);

BUFx3_ASAP7_75t_L g259 ( 
.A(n_187),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_259),
.B(n_248),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_157),
.B(n_183),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_183),
.B(n_171),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_261),
.B(n_254),
.Y(n_310)
);

XOR2xp5_ASAP7_75t_L g262 ( 
.A(n_171),
.B(n_180),
.Y(n_262)
);

INVxp67_ASAP7_75t_L g314 ( 
.A(n_264),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_247),
.B(n_234),
.C(n_200),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_271),
.B(n_287),
.C(n_292),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_L g312 ( 
.A1(n_272),
.A2(n_279),
.B1(n_258),
.B2(n_207),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_240),
.A2(n_262),
.B1(n_261),
.B2(n_260),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_L g317 ( 
.A1(n_275),
.A2(n_283),
.B1(n_295),
.B2(n_304),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_226),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_278),
.B(n_288),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_225),
.A2(n_203),
.B1(n_208),
.B2(n_213),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_220),
.A2(n_238),
.B1(n_221),
.B2(n_211),
.Y(n_283)
);

OAI21xp5_ASAP7_75t_L g316 ( 
.A1(n_286),
.A2(n_223),
.B(n_209),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_233),
.B(n_216),
.C(n_237),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_227),
.Y(n_288)
);

CKINVDCx16_ASAP7_75t_R g323 ( 
.A(n_289),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_233),
.B(n_243),
.C(n_231),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_241),
.A2(n_239),
.B1(n_224),
.B2(n_251),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_301),
.B(n_305),
.Y(n_326)
);

INVxp33_ASAP7_75t_L g320 ( 
.A(n_302),
.Y(n_320)
);

AOI22xp33_ASAP7_75t_L g304 ( 
.A1(n_222),
.A2(n_235),
.B1(n_241),
.B2(n_199),
.Y(n_304)
);

CKINVDCx20_ASAP7_75t_R g305 ( 
.A(n_210),
.Y(n_305)
);

CKINVDCx16_ASAP7_75t_R g329 ( 
.A(n_306),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_215),
.B(n_244),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_308),
.B(n_278),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_SL g341 ( 
.A(n_310),
.B(n_271),
.Y(n_341)
);

XOR2xp5_ASAP7_75t_L g311 ( 
.A(n_207),
.B(n_253),
.Y(n_311)
);

XOR2xp5_ASAP7_75t_L g346 ( 
.A(n_311),
.B(n_291),
.Y(n_346)
);

OAI22xp5_ASAP7_75t_SL g370 ( 
.A1(n_312),
.A2(n_341),
.B1(n_326),
.B2(n_340),
.Y(n_370)
);

AOI21xp5_ASAP7_75t_L g313 ( 
.A1(n_306),
.A2(n_212),
.B(n_229),
.Y(n_313)
);

OA21x2_ASAP7_75t_L g351 ( 
.A1(n_313),
.A2(n_316),
.B(n_331),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_290),
.B(n_259),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_318),
.B(n_322),
.Y(n_355)
);

CKINVDCx20_ASAP7_75t_R g319 ( 
.A(n_280),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g367 ( 
.A(n_319),
.B(n_324),
.Y(n_367)
);

OAI22xp5_ASAP7_75t_SL g322 ( 
.A1(n_272),
.A2(n_219),
.B1(n_275),
.B2(n_295),
.Y(n_322)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_280),
.Y(n_324)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_324),
.Y(n_352)
);

INVx2_ASAP7_75t_L g325 ( 
.A(n_284),
.Y(n_325)
);

INVx2_ASAP7_75t_L g377 ( 
.A(n_325),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_SL g366 ( 
.A(n_327),
.B(n_341),
.Y(n_366)
);

INVx3_ASAP7_75t_L g328 ( 
.A(n_299),
.Y(n_328)
);

INVx4_ASAP7_75t_L g360 ( 
.A(n_328),
.Y(n_360)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_294),
.Y(n_330)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_330),
.Y(n_356)
);

AOI21xp5_ASAP7_75t_L g331 ( 
.A1(n_303),
.A2(n_286),
.B(n_269),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_294),
.Y(n_332)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_332),
.Y(n_357)
);

OAI22xp5_ASAP7_75t_L g333 ( 
.A1(n_310),
.A2(n_283),
.B1(n_290),
.B2(n_268),
.Y(n_333)
);

OAI22xp5_ASAP7_75t_L g353 ( 
.A1(n_333),
.A2(n_334),
.B1(n_342),
.B2(n_349),
.Y(n_353)
);

AOI22xp5_ASAP7_75t_L g334 ( 
.A1(n_279),
.A2(n_270),
.B1(n_298),
.B2(n_268),
.Y(n_334)
);

INVx2_ASAP7_75t_L g335 ( 
.A(n_284),
.Y(n_335)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_335),
.Y(n_358)
);

AOI22xp33_ASAP7_75t_L g336 ( 
.A1(n_263),
.A2(n_296),
.B1(n_286),
.B2(n_303),
.Y(n_336)
);

AOI22xp33_ASAP7_75t_L g362 ( 
.A1(n_336),
.A2(n_297),
.B1(n_273),
.B2(n_276),
.Y(n_362)
);

OAI22xp5_ASAP7_75t_SL g337 ( 
.A1(n_277),
.A2(n_298),
.B1(n_286),
.B2(n_309),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_337),
.B(n_338),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_L g338 ( 
.A(n_282),
.B(n_265),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_277),
.B(n_269),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_339),
.B(n_340),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_311),
.B(n_287),
.Y(n_340)
);

AOI22xp5_ASAP7_75t_L g342 ( 
.A1(n_286),
.A2(n_292),
.B1(n_301),
.B2(n_293),
.Y(n_342)
);

OAI21xp5_ASAP7_75t_L g343 ( 
.A1(n_300),
.A2(n_289),
.B(n_274),
.Y(n_343)
);

XNOR2xp5_ASAP7_75t_SL g376 ( 
.A(n_343),
.B(n_346),
.Y(n_376)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_274),
.Y(n_344)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_344),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_285),
.B(n_267),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_SL g369 ( 
.A(n_345),
.B(n_348),
.Y(n_369)
);

NAND2x1p5_ASAP7_75t_L g347 ( 
.A(n_267),
.B(n_266),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_L g354 ( 
.A(n_347),
.B(n_307),
.C(n_273),
.Y(n_354)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_281),
.Y(n_348)
);

OAI22xp5_ASAP7_75t_SL g349 ( 
.A1(n_297),
.A2(n_266),
.B1(n_299),
.B2(n_281),
.Y(n_349)
);

XOR2x2_ASAP7_75t_L g350 ( 
.A(n_346),
.B(n_276),
.Y(n_350)
);

XOR2xp5_ASAP7_75t_L g381 ( 
.A(n_350),
.B(n_315),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_SL g394 ( 
.A(n_354),
.B(n_370),
.Y(n_394)
);

OAI22xp5_ASAP7_75t_L g359 ( 
.A1(n_334),
.A2(n_333),
.B1(n_317),
.B2(n_319),
.Y(n_359)
);

OAI22xp5_ASAP7_75t_L g398 ( 
.A1(n_359),
.A2(n_362),
.B1(n_363),
.B2(n_373),
.Y(n_398)
);

INVx3_ASAP7_75t_L g361 ( 
.A(n_328),
.Y(n_361)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_361),
.Y(n_380)
);

AOI22xp33_ASAP7_75t_L g363 ( 
.A1(n_314),
.A2(n_297),
.B1(n_307),
.B2(n_323),
.Y(n_363)
);

CKINVDCx12_ASAP7_75t_R g365 ( 
.A(n_320),
.Y(n_365)
);

CKINVDCx20_ASAP7_75t_R g391 ( 
.A(n_365),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_367),
.B(n_374),
.Y(n_393)
);

AND2x6_ASAP7_75t_L g368 ( 
.A(n_331),
.B(n_342),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_368),
.B(n_353),
.Y(n_404)
);

NOR2xp33_ASAP7_75t_L g372 ( 
.A(n_338),
.B(n_327),
.Y(n_372)
);

NOR2xp33_ASAP7_75t_L g397 ( 
.A(n_372),
.B(n_378),
.Y(n_397)
);

OAI22xp5_ASAP7_75t_L g373 ( 
.A1(n_317),
.A2(n_330),
.B1(n_332),
.B2(n_329),
.Y(n_373)
);

OAI22xp5_ASAP7_75t_SL g374 ( 
.A1(n_312),
.A2(n_329),
.B1(n_323),
.B2(n_313),
.Y(n_374)
);

AND2x6_ASAP7_75t_L g375 ( 
.A(n_339),
.B(n_337),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_375),
.B(n_349),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_SL g378 ( 
.A(n_321),
.B(n_345),
.Y(n_378)
);

XOR2xp5_ASAP7_75t_L g410 ( 
.A(n_381),
.B(n_385),
.Y(n_410)
);

AOI21xp5_ASAP7_75t_L g382 ( 
.A1(n_351),
.A2(n_316),
.B(n_343),
.Y(n_382)
);

OAI21xp5_ASAP7_75t_SL g407 ( 
.A1(n_382),
.A2(n_383),
.B(n_389),
.Y(n_407)
);

AOI21xp5_ASAP7_75t_L g383 ( 
.A1(n_351),
.A2(n_322),
.B(n_347),
.Y(n_383)
);

XOR2xp5_ASAP7_75t_L g384 ( 
.A(n_379),
.B(n_315),
.Y(n_384)
);

MAJIxp5_ASAP7_75t_L g419 ( 
.A(n_384),
.B(n_392),
.C(n_396),
.Y(n_419)
);

XNOR2xp5_ASAP7_75t_L g385 ( 
.A(n_379),
.B(n_326),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_371),
.Y(n_386)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_386),
.Y(n_417)
);

OAI32xp33_ASAP7_75t_L g387 ( 
.A1(n_364),
.A2(n_318),
.A3(n_321),
.B1(n_344),
.B2(n_335),
.Y(n_387)
);

INVxp67_ASAP7_75t_L g421 ( 
.A(n_387),
.Y(n_421)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_371),
.Y(n_388)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_388),
.Y(n_424)
);

AOI21xp5_ASAP7_75t_L g389 ( 
.A1(n_351),
.A2(n_347),
.B(n_325),
.Y(n_389)
);

OAI21xp5_ASAP7_75t_L g390 ( 
.A1(n_374),
.A2(n_364),
.B(n_355),
.Y(n_390)
);

AND2x2_ASAP7_75t_L g405 ( 
.A(n_390),
.B(n_373),
.Y(n_405)
);

XNOR2xp5_ASAP7_75t_SL g392 ( 
.A(n_370),
.B(n_347),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_395),
.B(n_399),
.Y(n_412)
);

XNOR2xp5_ASAP7_75t_SL g396 ( 
.A(n_376),
.B(n_348),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g399 ( 
.A(n_369),
.B(n_352),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_358),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_400),
.B(n_358),
.Y(n_413)
);

CKINVDCx16_ASAP7_75t_R g401 ( 
.A(n_354),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_SL g425 ( 
.A(n_401),
.B(n_381),
.Y(n_425)
);

MAJIxp5_ASAP7_75t_L g402 ( 
.A(n_350),
.B(n_376),
.C(n_366),
.Y(n_402)
);

MAJIxp5_ASAP7_75t_L g426 ( 
.A(n_402),
.B(n_403),
.C(n_401),
.Y(n_426)
);

XNOR2xp5_ASAP7_75t_L g403 ( 
.A(n_359),
.B(n_353),
.Y(n_403)
);

OAI22xp5_ASAP7_75t_L g420 ( 
.A1(n_404),
.A2(n_360),
.B1(n_383),
.B2(n_395),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_SL g437 ( 
.A(n_405),
.B(n_407),
.Y(n_437)
);

AOI22xp5_ASAP7_75t_L g406 ( 
.A1(n_403),
.A2(n_355),
.B1(n_352),
.B2(n_356),
.Y(n_406)
);

OAI22xp5_ASAP7_75t_SL g430 ( 
.A1(n_406),
.A2(n_416),
.B1(n_418),
.B2(n_405),
.Y(n_430)
);

XNOR2xp5_ASAP7_75t_L g408 ( 
.A(n_384),
.B(n_356),
.Y(n_408)
);

XOR2xp5_ASAP7_75t_L g433 ( 
.A(n_408),
.B(n_426),
.Y(n_433)
);

NOR2xp33_ASAP7_75t_L g409 ( 
.A(n_391),
.B(n_357),
.Y(n_409)
);

INVxp67_ASAP7_75t_SL g429 ( 
.A(n_409),
.Y(n_429)
);

CKINVDCx14_ASAP7_75t_R g411 ( 
.A(n_397),
.Y(n_411)
);

CKINVDCx20_ASAP7_75t_R g428 ( 
.A(n_411),
.Y(n_428)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_413),
.Y(n_439)
);

CKINVDCx16_ASAP7_75t_R g414 ( 
.A(n_393),
.Y(n_414)
);

NOR2xp33_ASAP7_75t_L g435 ( 
.A(n_414),
.B(n_423),
.Y(n_435)
);

AND2x2_ASAP7_75t_L g415 ( 
.A(n_389),
.B(n_357),
.Y(n_415)
);

CKINVDCx16_ASAP7_75t_R g442 ( 
.A(n_415),
.Y(n_442)
);

AOI22xp5_ASAP7_75t_L g416 ( 
.A1(n_390),
.A2(n_375),
.B1(n_368),
.B2(n_377),
.Y(n_416)
);

AOI22xp5_ASAP7_75t_L g418 ( 
.A1(n_398),
.A2(n_377),
.B1(n_361),
.B2(n_360),
.Y(n_418)
);

OAI21xp5_ASAP7_75t_SL g431 ( 
.A1(n_420),
.A2(n_393),
.B(n_404),
.Y(n_431)
);

AND2x2_ASAP7_75t_L g422 ( 
.A(n_382),
.B(n_398),
.Y(n_422)
);

CKINVDCx14_ASAP7_75t_R g443 ( 
.A(n_422),
.Y(n_443)
);

CKINVDCx20_ASAP7_75t_R g423 ( 
.A(n_399),
.Y(n_423)
);

XNOR2xp5_ASAP7_75t_L g441 ( 
.A(n_425),
.B(n_380),
.Y(n_441)
);

MAJIxp5_ASAP7_75t_L g427 ( 
.A(n_410),
.B(n_394),
.C(n_402),
.Y(n_427)
);

MAJIxp5_ASAP7_75t_L g447 ( 
.A(n_427),
.B(n_438),
.C(n_440),
.Y(n_447)
);

AOI22xp5_ASAP7_75t_L g449 ( 
.A1(n_430),
.A2(n_432),
.B1(n_436),
.B2(n_405),
.Y(n_449)
);

INVxp67_ASAP7_75t_L g457 ( 
.A(n_431),
.Y(n_457)
);

OAI22xp5_ASAP7_75t_SL g432 ( 
.A1(n_421),
.A2(n_394),
.B1(n_392),
.B2(n_387),
.Y(n_432)
);

XOR2xp5_ASAP7_75t_L g434 ( 
.A(n_410),
.B(n_396),
.Y(n_434)
);

XOR2xp5_ASAP7_75t_L g448 ( 
.A(n_434),
.B(n_441),
.Y(n_448)
);

AOI22xp5_ASAP7_75t_L g436 ( 
.A1(n_421),
.A2(n_385),
.B1(n_397),
.B2(n_386),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_437),
.B(n_407),
.Y(n_451)
);

MAJIxp5_ASAP7_75t_L g438 ( 
.A(n_426),
.B(n_408),
.C(n_419),
.Y(n_438)
);

MAJIxp5_ASAP7_75t_L g440 ( 
.A(n_419),
.B(n_400),
.C(n_388),
.Y(n_440)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_413),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_444),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_SL g446 ( 
.A(n_428),
.B(n_391),
.Y(n_446)
);

NOR2xp33_ASAP7_75t_L g459 ( 
.A(n_446),
.B(n_449),
.Y(n_459)
);

XNOR2xp5_ASAP7_75t_L g450 ( 
.A(n_440),
.B(n_416),
.Y(n_450)
);

NOR2xp33_ASAP7_75t_L g467 ( 
.A(n_450),
.B(n_454),
.Y(n_467)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_451),
.Y(n_460)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_435),
.Y(n_452)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_452),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_428),
.B(n_406),
.Y(n_453)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_453),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_429),
.B(n_380),
.Y(n_454)
);

AOI21xp5_ASAP7_75t_L g455 ( 
.A1(n_437),
.A2(n_415),
.B(n_422),
.Y(n_455)
);

OAI21xp5_ASAP7_75t_SL g463 ( 
.A1(n_455),
.A2(n_422),
.B(n_415),
.Y(n_463)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_439),
.Y(n_456)
);

NOR2xp33_ASAP7_75t_L g468 ( 
.A(n_456),
.B(n_417),
.Y(n_468)
);

BUFx6f_ASAP7_75t_L g458 ( 
.A(n_445),
.Y(n_458)
);

NOR2xp33_ASAP7_75t_L g474 ( 
.A(n_458),
.B(n_468),
.Y(n_474)
);

AOI21xp5_ASAP7_75t_L g461 ( 
.A1(n_451),
.A2(n_455),
.B(n_457),
.Y(n_461)
);

AND2x2_ASAP7_75t_L g475 ( 
.A(n_461),
.B(n_453),
.Y(n_475)
);

XOR2xp5_ASAP7_75t_L g473 ( 
.A(n_463),
.B(n_461),
.Y(n_473)
);

MAJIxp5_ASAP7_75t_L g464 ( 
.A(n_447),
.B(n_433),
.C(n_438),
.Y(n_464)
);

NOR2xp67_ASAP7_75t_SL g471 ( 
.A(n_464),
.B(n_465),
.Y(n_471)
);

MAJIxp5_ASAP7_75t_L g465 ( 
.A(n_447),
.B(n_433),
.C(n_427),
.Y(n_465)
);

NOR2xp33_ASAP7_75t_SL g469 ( 
.A(n_466),
.B(n_436),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_L g481 ( 
.A(n_469),
.B(n_477),
.Y(n_481)
);

OAI22xp5_ASAP7_75t_SL g470 ( 
.A1(n_459),
.A2(n_449),
.B1(n_457),
.B2(n_412),
.Y(n_470)
);

AOI22xp5_ASAP7_75t_L g482 ( 
.A1(n_470),
.A2(n_475),
.B1(n_462),
.B2(n_412),
.Y(n_482)
);

MAJIxp5_ASAP7_75t_L g472 ( 
.A(n_464),
.B(n_450),
.C(n_441),
.Y(n_472)
);

OR2x2_ASAP7_75t_L g479 ( 
.A(n_472),
.B(n_476),
.Y(n_479)
);

XNOR2xp5_ASAP7_75t_L g484 ( 
.A(n_473),
.B(n_448),
.Y(n_484)
);

AOI22xp5_ASAP7_75t_SL g476 ( 
.A1(n_460),
.A2(n_430),
.B1(n_443),
.B2(n_432),
.Y(n_476)
);

XNOR2xp5_ASAP7_75t_L g477 ( 
.A(n_465),
.B(n_448),
.Y(n_477)
);

MAJIxp5_ASAP7_75t_L g478 ( 
.A(n_471),
.B(n_467),
.C(n_460),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_L g489 ( 
.A(n_478),
.B(n_474),
.Y(n_489)
);

AOI221xp5_ASAP7_75t_L g480 ( 
.A1(n_475),
.A2(n_462),
.B1(n_439),
.B2(n_444),
.C(n_442),
.Y(n_480)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_480),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_L g488 ( 
.A(n_482),
.B(n_483),
.Y(n_488)
);

AOI322xp5_ASAP7_75t_L g483 ( 
.A1(n_476),
.A2(n_431),
.A3(n_463),
.B1(n_458),
.B2(n_442),
.C1(n_417),
.C2(n_424),
.Y(n_483)
);

AND2x2_ASAP7_75t_L g485 ( 
.A(n_484),
.B(n_472),
.Y(n_485)
);

XOR2xp5_ASAP7_75t_L g490 ( 
.A(n_485),
.B(n_488),
.Y(n_490)
);

XOR2xp5_ASAP7_75t_L g486 ( 
.A(n_481),
.B(n_473),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_L g492 ( 
.A(n_486),
.B(n_489),
.Y(n_492)
);

AOI21xp5_ASAP7_75t_SL g494 ( 
.A1(n_490),
.A2(n_491),
.B(n_487),
.Y(n_494)
);

OAI21xp5_ASAP7_75t_SL g491 ( 
.A1(n_485),
.A2(n_479),
.B(n_480),
.Y(n_491)
);

BUFx24_ASAP7_75t_SL g493 ( 
.A(n_492),
.Y(n_493)
);

OAI22xp5_ASAP7_75t_L g495 ( 
.A1(n_493),
.A2(n_494),
.B1(n_424),
.B2(n_418),
.Y(n_495)
);

OAI21xp5_ASAP7_75t_L g496 ( 
.A1(n_495),
.A2(n_483),
.B(n_434),
.Y(n_496)
);

BUFx24_ASAP7_75t_SL g497 ( 
.A(n_496),
.Y(n_497)
);


endmodule