module fake_jpeg_28813_n_540 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_540);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_540;

wire n_529;
wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_17),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_4),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_5),
.Y(n_22)
);

INVx6_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_17),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_9),
.Y(n_25)
);

BUFx12_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_0),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_2),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_0),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_17),
.Y(n_33)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_12),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_10),
.Y(n_35)
);

INVxp67_ASAP7_75t_L g36 ( 
.A(n_13),
.Y(n_36)
);

BUFx5_ASAP7_75t_L g37 ( 
.A(n_7),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_10),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_11),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_0),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_2),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_8),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_0),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_4),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_2),
.Y(n_45)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_15),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_5),
.Y(n_47)
);

INVx1_ASAP7_75t_SL g48 ( 
.A(n_8),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_4),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_12),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_16),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_10),
.Y(n_52)
);

BUFx5_ASAP7_75t_L g53 ( 
.A(n_6),
.Y(n_53)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_6),
.Y(n_54)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_27),
.Y(n_55)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_55),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_35),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_56),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_35),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_57),
.Y(n_131)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_35),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_58),
.Y(n_135)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_27),
.Y(n_59)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_59),
.Y(n_112)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_37),
.Y(n_60)
);

INVx5_ASAP7_75t_L g141 ( 
.A(n_60),
.Y(n_141)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_34),
.Y(n_61)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_61),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_36),
.B(n_15),
.Y(n_62)
);

AND2x2_ASAP7_75t_L g144 ( 
.A(n_62),
.B(n_85),
.Y(n_144)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_35),
.Y(n_63)
);

INVx3_ASAP7_75t_L g158 ( 
.A(n_63),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_31),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g148 ( 
.A(n_64),
.Y(n_148)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_33),
.Y(n_65)
);

INVx3_ASAP7_75t_L g165 ( 
.A(n_65),
.Y(n_165)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_31),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g151 ( 
.A(n_66),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_31),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g154 ( 
.A(n_67),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_24),
.B(n_16),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_68),
.B(n_103),
.Y(n_152)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_34),
.Y(n_69)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_69),
.Y(n_123)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_37),
.Y(n_70)
);

INVx8_ASAP7_75t_L g119 ( 
.A(n_70),
.Y(n_119)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_33),
.Y(n_71)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_71),
.Y(n_127)
);

INVx11_ASAP7_75t_L g72 ( 
.A(n_54),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g172 ( 
.A(n_72),
.Y(n_172)
);

BUFx3_ASAP7_75t_L g73 ( 
.A(n_37),
.Y(n_73)
);

INVx5_ASAP7_75t_L g143 ( 
.A(n_73),
.Y(n_143)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_34),
.Y(n_74)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_74),
.Y(n_129)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_33),
.Y(n_75)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_75),
.Y(n_136)
);

INVx6_ASAP7_75t_L g76 ( 
.A(n_39),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g173 ( 
.A(n_76),
.Y(n_173)
);

INVx11_ASAP7_75t_L g77 ( 
.A(n_54),
.Y(n_77)
);

INVx5_ASAP7_75t_L g149 ( 
.A(n_77),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_39),
.Y(n_78)
);

INVx6_ASAP7_75t_L g164 ( 
.A(n_78),
.Y(n_164)
);

INVx5_ASAP7_75t_L g79 ( 
.A(n_53),
.Y(n_79)
);

INVx5_ASAP7_75t_L g155 ( 
.A(n_79),
.Y(n_155)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_46),
.Y(n_80)
);

INVx4_ASAP7_75t_L g121 ( 
.A(n_80),
.Y(n_121)
);

INVx8_ASAP7_75t_L g81 ( 
.A(n_53),
.Y(n_81)
);

INVx8_ASAP7_75t_L g163 ( 
.A(n_81),
.Y(n_163)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_46),
.Y(n_82)
);

INVx4_ASAP7_75t_L g122 ( 
.A(n_82),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_39),
.Y(n_83)
);

INVx6_ASAP7_75t_L g170 ( 
.A(n_83),
.Y(n_170)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_46),
.Y(n_84)
);

INVx4_ASAP7_75t_L g146 ( 
.A(n_84),
.Y(n_146)
);

AND2x2_ASAP7_75t_SL g85 ( 
.A(n_19),
.B(n_1),
.Y(n_85)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_48),
.B(n_16),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_86),
.B(n_87),
.Y(n_115)
);

INVx1_ASAP7_75t_SL g87 ( 
.A(n_18),
.Y(n_87)
);

INVx13_ASAP7_75t_L g88 ( 
.A(n_54),
.Y(n_88)
);

BUFx12f_ASAP7_75t_L g114 ( 
.A(n_88),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_42),
.Y(n_89)
);

INVx6_ASAP7_75t_L g171 ( 
.A(n_89),
.Y(n_171)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_23),
.Y(n_90)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_90),
.Y(n_138)
);

BUFx3_ASAP7_75t_L g91 ( 
.A(n_53),
.Y(n_91)
);

BUFx3_ASAP7_75t_L g140 ( 
.A(n_91),
.Y(n_140)
);

AOI21xp33_ASAP7_75t_L g92 ( 
.A1(n_18),
.A2(n_15),
.B(n_14),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g153 ( 
.A(n_92),
.B(n_106),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_42),
.Y(n_93)
);

INVx3_ASAP7_75t_SL g120 ( 
.A(n_93),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_42),
.Y(n_94)
);

BUFx2_ASAP7_75t_L g126 ( 
.A(n_94),
.Y(n_126)
);

INVx8_ASAP7_75t_L g95 ( 
.A(n_49),
.Y(n_95)
);

INVx4_ASAP7_75t_L g159 ( 
.A(n_95),
.Y(n_159)
);

BUFx3_ASAP7_75t_L g96 ( 
.A(n_44),
.Y(n_96)
);

INVx4_ASAP7_75t_L g162 ( 
.A(n_96),
.Y(n_162)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_48),
.B(n_14),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_97),
.B(n_48),
.Y(n_130)
);

BUFx3_ASAP7_75t_L g98 ( 
.A(n_44),
.Y(n_98)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_98),
.Y(n_167)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_23),
.Y(n_99)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_99),
.Y(n_168)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_23),
.Y(n_100)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_100),
.Y(n_145)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_44),
.Y(n_101)
);

INVx13_ASAP7_75t_L g124 ( 
.A(n_101),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_49),
.Y(n_102)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_102),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_49),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_50),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_104),
.B(n_105),
.Y(n_161)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_50),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_24),
.B(n_51),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_50),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_107),
.A2(n_108),
.B1(n_110),
.B2(n_32),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_19),
.Y(n_108)
);

BUFx5_ASAP7_75t_L g109 ( 
.A(n_32),
.Y(n_109)
);

INVx13_ASAP7_75t_L g132 ( 
.A(n_109),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_19),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_106),
.B(n_51),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_117),
.B(n_142),
.Y(n_226)
);

INVxp67_ASAP7_75t_L g220 ( 
.A(n_118),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_62),
.A2(n_25),
.B1(n_20),
.B2(n_47),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g188 ( 
.A1(n_125),
.A2(n_133),
.B1(n_139),
.B2(n_30),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g128 ( 
.A(n_88),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_128),
.B(n_157),
.Y(n_183)
);

AND2x2_ASAP7_75t_L g215 ( 
.A(n_130),
.B(n_146),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_85),
.A2(n_22),
.B1(n_47),
.B2(n_45),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_86),
.B(n_22),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_SL g194 ( 
.A(n_134),
.B(n_137),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_97),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_SL g139 ( 
.A1(n_95),
.A2(n_32),
.B1(n_52),
.B2(n_21),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_70),
.B(n_45),
.Y(n_142)
);

AOI21xp33_ASAP7_75t_L g147 ( 
.A1(n_81),
.A2(n_21),
.B(n_43),
.Y(n_147)
);

AOI21xp33_ASAP7_75t_L g178 ( 
.A1(n_147),
.A2(n_41),
.B(n_40),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_SL g156 ( 
.A(n_63),
.B(n_20),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_156),
.B(n_28),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_63),
.B(n_25),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_108),
.B(n_38),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_160),
.B(n_169),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_110),
.B(n_38),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_166),
.B(n_29),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_SL g169 ( 
.A(n_66),
.B(n_30),
.Y(n_169)
);

BUFx3_ASAP7_75t_L g174 ( 
.A(n_140),
.Y(n_174)
);

CKINVDCx14_ASAP7_75t_R g244 ( 
.A(n_174),
.Y(n_244)
);

BUFx2_ASAP7_75t_L g175 ( 
.A(n_167),
.Y(n_175)
);

INVx3_ASAP7_75t_L g231 ( 
.A(n_175),
.Y(n_231)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_127),
.Y(n_176)
);

CKINVDCx16_ASAP7_75t_R g248 ( 
.A(n_176),
.Y(n_248)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_111),
.Y(n_177)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_177),
.Y(n_230)
);

AO21x1_ASAP7_75t_L g241 ( 
.A1(n_178),
.A2(n_202),
.B(n_215),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_126),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g243 ( 
.A(n_179),
.B(n_212),
.Y(n_243)
);

AND2x4_ASAP7_75t_L g180 ( 
.A(n_152),
.B(n_32),
.Y(n_180)
);

AND2x2_ASAP7_75t_L g232 ( 
.A(n_180),
.B(n_188),
.Y(n_232)
);

INVx3_ASAP7_75t_L g181 ( 
.A(n_114),
.Y(n_181)
);

INVx3_ASAP7_75t_L g235 ( 
.A(n_181),
.Y(n_235)
);

AOI22xp33_ASAP7_75t_L g182 ( 
.A1(n_164),
.A2(n_76),
.B1(n_107),
.B2(n_103),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g250 ( 
.A1(n_182),
.A2(n_189),
.B1(n_192),
.B2(n_193),
.Y(n_250)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_145),
.Y(n_184)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_184),
.Y(n_238)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_113),
.Y(n_185)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_185),
.Y(n_239)
);

INVx4_ASAP7_75t_L g186 ( 
.A(n_158),
.Y(n_186)
);

INVx3_ASAP7_75t_L g237 ( 
.A(n_186),
.Y(n_237)
);

AOI21xp5_ASAP7_75t_L g187 ( 
.A1(n_153),
.A2(n_14),
.B(n_58),
.Y(n_187)
);

INVxp67_ASAP7_75t_L g247 ( 
.A(n_187),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_144),
.A2(n_78),
.B1(n_102),
.B2(n_94),
.Y(n_189)
);

INVx3_ASAP7_75t_L g190 ( 
.A(n_114),
.Y(n_190)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_190),
.Y(n_251)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_123),
.Y(n_191)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_191),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_144),
.A2(n_104),
.B1(n_93),
.B2(n_89),
.Y(n_192)
);

AOI22xp33_ASAP7_75t_L g193 ( 
.A1(n_164),
.A2(n_67),
.B1(n_64),
.B2(n_83),
.Y(n_193)
);

INVx6_ASAP7_75t_L g195 ( 
.A(n_116),
.Y(n_195)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_195),
.Y(n_254)
);

INVx6_ASAP7_75t_L g196 ( 
.A(n_116),
.Y(n_196)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_196),
.Y(n_272)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_112),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_197),
.B(n_198),
.Y(n_242)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_129),
.Y(n_198)
);

INVx3_ASAP7_75t_L g199 ( 
.A(n_114),
.Y(n_199)
);

INVx11_ASAP7_75t_L g265 ( 
.A(n_199),
.Y(n_265)
);

AOI21xp5_ASAP7_75t_L g200 ( 
.A1(n_115),
.A2(n_43),
.B(n_41),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_200),
.B(n_201),
.Y(n_245)
);

AND2x2_ASAP7_75t_SL g201 ( 
.A(n_161),
.B(n_136),
.Y(n_201)
);

OAI21xp33_ASAP7_75t_L g202 ( 
.A1(n_120),
.A2(n_52),
.B(n_40),
.Y(n_202)
);

OAI22xp33_ASAP7_75t_SL g203 ( 
.A1(n_150),
.A2(n_57),
.B1(n_56),
.B2(n_32),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_L g269 ( 
.A1(n_203),
.A2(n_154),
.B1(n_148),
.B2(n_131),
.Y(n_269)
);

CKINVDCx16_ASAP7_75t_R g204 ( 
.A(n_139),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_204),
.B(n_205),
.Y(n_255)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_138),
.Y(n_205)
);

BUFx3_ASAP7_75t_L g206 ( 
.A(n_140),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_206),
.Y(n_233)
);

INVx5_ASAP7_75t_L g207 ( 
.A(n_132),
.Y(n_207)
);

BUFx12f_ASAP7_75t_L g273 ( 
.A(n_207),
.Y(n_273)
);

INVx6_ASAP7_75t_L g208 ( 
.A(n_131),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_208),
.B(n_209),
.Y(n_259)
);

INVx3_ASAP7_75t_L g209 ( 
.A(n_149),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_168),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_210),
.B(n_213),
.Y(n_260)
);

INVx5_ASAP7_75t_L g211 ( 
.A(n_132),
.Y(n_211)
);

BUFx12_ASAP7_75t_L g249 ( 
.A(n_211),
.Y(n_249)
);

CKINVDCx14_ASAP7_75t_R g212 ( 
.A(n_124),
.Y(n_212)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_151),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_126),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_SL g253 ( 
.A(n_214),
.B(n_228),
.Y(n_253)
);

HB1xp67_ASAP7_75t_L g216 ( 
.A(n_165),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_216),
.B(n_218),
.Y(n_263)
);

INVx2_ASAP7_75t_SL g217 ( 
.A(n_170),
.Y(n_217)
);

BUFx24_ASAP7_75t_L g268 ( 
.A(n_217),
.Y(n_268)
);

INVx4_ASAP7_75t_L g218 ( 
.A(n_162),
.Y(n_218)
);

AOI22xp33_ASAP7_75t_SL g219 ( 
.A1(n_141),
.A2(n_29),
.B1(n_28),
.B2(n_5),
.Y(n_219)
);

AOI22xp33_ASAP7_75t_SL g257 ( 
.A1(n_219),
.A2(n_221),
.B1(n_171),
.B2(n_170),
.Y(n_257)
);

BUFx6f_ASAP7_75t_L g221 ( 
.A(n_148),
.Y(n_221)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_173),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_222),
.B(n_223),
.Y(n_264)
);

INVx3_ASAP7_75t_L g223 ( 
.A(n_172),
.Y(n_223)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_173),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_225),
.B(n_227),
.Y(n_271)
);

HB1xp67_ASAP7_75t_L g227 ( 
.A(n_121),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_SL g270 ( 
.A(n_229),
.B(n_146),
.Y(n_270)
);

AO22x1_ASAP7_75t_SL g234 ( 
.A1(n_180),
.A2(n_120),
.B1(n_151),
.B2(n_135),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_234),
.B(n_240),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_175),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g291 ( 
.A(n_236),
.B(n_252),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_180),
.B(n_171),
.Y(n_240)
);

MAJx2_ASAP7_75t_L g246 ( 
.A(n_215),
.B(n_118),
.C(n_124),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_246),
.B(n_262),
.C(n_202),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_201),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_183),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_SL g292 ( 
.A(n_256),
.B(n_258),
.Y(n_292)
);

INVxp67_ASAP7_75t_L g288 ( 
.A(n_257),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_SL g258 ( 
.A(n_224),
.B(n_122),
.Y(n_258)
);

AOI22xp33_ASAP7_75t_SL g261 ( 
.A1(n_220),
.A2(n_143),
.B1(n_119),
.B2(n_163),
.Y(n_261)
);

INVxp67_ASAP7_75t_L g305 ( 
.A(n_261),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_226),
.B(n_121),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_174),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_SL g293 ( 
.A(n_267),
.B(n_190),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_269),
.A2(n_203),
.B1(n_154),
.B2(n_208),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_SL g274 ( 
.A(n_270),
.B(n_253),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_274),
.B(n_287),
.Y(n_339)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_239),
.Y(n_275)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_275),
.Y(n_310)
);

HB1xp67_ASAP7_75t_L g276 ( 
.A(n_235),
.Y(n_276)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_276),
.Y(n_315)
);

AOI21xp5_ASAP7_75t_L g277 ( 
.A1(n_255),
.A2(n_220),
.B(n_207),
.Y(n_277)
);

AOI21xp5_ASAP7_75t_L g320 ( 
.A1(n_277),
.A2(n_241),
.B(n_259),
.Y(n_320)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_239),
.Y(n_279)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_279),
.Y(n_326)
);

BUFx6f_ASAP7_75t_L g280 ( 
.A(n_254),
.Y(n_280)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_280),
.Y(n_338)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_266),
.Y(n_281)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_281),
.Y(n_340)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_266),
.Y(n_282)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_282),
.Y(n_342)
);

INVx11_ASAP7_75t_L g283 ( 
.A(n_273),
.Y(n_283)
);

INVx2_ASAP7_75t_SL g332 ( 
.A(n_283),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_252),
.B(n_218),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_284),
.B(n_285),
.Y(n_317)
);

BUFx8_ASAP7_75t_L g286 ( 
.A(n_273),
.Y(n_286)
);

CKINVDCx14_ASAP7_75t_R g333 ( 
.A(n_286),
.Y(n_333)
);

INVx5_ASAP7_75t_L g287 ( 
.A(n_235),
.Y(n_287)
);

AOI22xp33_ASAP7_75t_SL g289 ( 
.A1(n_256),
.A2(n_211),
.B1(n_206),
.B2(n_119),
.Y(n_289)
);

AOI22xp33_ASAP7_75t_SL g328 ( 
.A1(n_289),
.A2(n_299),
.B1(n_273),
.B2(n_199),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_262),
.B(n_194),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_290),
.B(n_298),
.Y(n_330)
);

CKINVDCx14_ASAP7_75t_R g337 ( 
.A(n_293),
.Y(n_337)
);

OAI22xp5_ASAP7_75t_L g323 ( 
.A1(n_294),
.A2(n_300),
.B1(n_304),
.B2(n_278),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_242),
.Y(n_295)
);

OR2x2_ASAP7_75t_L g329 ( 
.A(n_295),
.B(n_264),
.Y(n_329)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_238),
.Y(n_296)
);

CKINVDCx16_ASAP7_75t_R g316 ( 
.A(n_296),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_SL g297 ( 
.A1(n_247),
.A2(n_182),
.B1(n_193),
.B2(n_219),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_L g312 ( 
.A1(n_297),
.A2(n_250),
.B1(n_269),
.B2(n_247),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_232),
.B(n_217),
.Y(n_298)
);

INVx2_ASAP7_75t_L g299 ( 
.A(n_230),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g300 ( 
.A1(n_232),
.A2(n_135),
.B1(n_159),
.B2(n_196),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_SL g325 ( 
.A1(n_300),
.A2(n_304),
.B1(n_236),
.B2(n_231),
.Y(n_325)
);

BUFx24_ASAP7_75t_SL g301 ( 
.A(n_258),
.Y(n_301)
);

INVxp67_ASAP7_75t_L g318 ( 
.A(n_301),
.Y(n_318)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_238),
.Y(n_302)
);

CKINVDCx16_ASAP7_75t_R g327 ( 
.A(n_302),
.Y(n_327)
);

XOR2xp5_ASAP7_75t_L g303 ( 
.A(n_245),
.B(n_122),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_SL g311 ( 
.A(n_303),
.B(n_306),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_232),
.A2(n_159),
.B1(n_195),
.B2(n_221),
.Y(n_304)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_260),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_SL g307 ( 
.A(n_245),
.B(n_162),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_SL g314 ( 
.A(n_307),
.B(n_308),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_240),
.B(n_209),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_243),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_SL g321 ( 
.A(n_309),
.B(n_248),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_SL g349 ( 
.A1(n_312),
.A2(n_313),
.B1(n_341),
.B2(n_305),
.Y(n_349)
);

AOI22xp33_ASAP7_75t_L g313 ( 
.A1(n_297),
.A2(n_250),
.B1(n_246),
.B2(n_234),
.Y(n_313)
);

OAI21xp33_ASAP7_75t_SL g319 ( 
.A1(n_278),
.A2(n_241),
.B(n_234),
.Y(n_319)
);

OAI21xp33_ASAP7_75t_SL g347 ( 
.A1(n_319),
.A2(n_320),
.B(n_277),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_SL g373 ( 
.A(n_321),
.B(n_329),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_SL g322 ( 
.A(n_295),
.B(n_271),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_322),
.B(n_324),
.Y(n_344)
);

AOI22xp5_ASAP7_75t_SL g371 ( 
.A1(n_323),
.A2(n_325),
.B1(n_268),
.B2(n_251),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_SL g324 ( 
.A(n_292),
.B(n_263),
.Y(n_324)
);

INVxp67_ASAP7_75t_L g343 ( 
.A(n_328),
.Y(n_343)
);

OAI22xp5_ASAP7_75t_SL g331 ( 
.A1(n_298),
.A2(n_254),
.B1(n_272),
.B2(n_223),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_331),
.B(n_334),
.Y(n_348)
);

OAI22xp5_ASAP7_75t_SL g334 ( 
.A1(n_285),
.A2(n_272),
.B1(n_233),
.B2(n_267),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_SL g335 ( 
.A(n_308),
.B(n_230),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_335),
.B(n_284),
.Y(n_353)
);

AOI22xp5_ASAP7_75t_SL g336 ( 
.A1(n_288),
.A2(n_233),
.B1(n_244),
.B2(n_237),
.Y(n_336)
);

AND2x2_ASAP7_75t_L g361 ( 
.A(n_336),
.B(n_287),
.Y(n_361)
);

AOI22xp5_ASAP7_75t_L g341 ( 
.A1(n_288),
.A2(n_231),
.B1(n_237),
.B2(n_163),
.Y(n_341)
);

CKINVDCx20_ASAP7_75t_R g345 ( 
.A(n_329),
.Y(n_345)
);

INVx11_ASAP7_75t_L g403 ( 
.A(n_345),
.Y(n_403)
);

XNOR2xp5_ASAP7_75t_SL g346 ( 
.A(n_314),
.B(n_311),
.Y(n_346)
);

XOR2xp5_ASAP7_75t_L g383 ( 
.A(n_346),
.B(n_331),
.Y(n_383)
);

AOI21xp5_ASAP7_75t_L g400 ( 
.A1(n_347),
.A2(n_361),
.B(n_332),
.Y(n_400)
);

AOI22xp5_ASAP7_75t_L g390 ( 
.A1(n_349),
.A2(n_358),
.B1(n_362),
.B2(n_366),
.Y(n_390)
);

MAJIxp5_ASAP7_75t_L g350 ( 
.A(n_311),
.B(n_307),
.C(n_303),
.Y(n_350)
);

MAJIxp5_ASAP7_75t_L g380 ( 
.A(n_350),
.B(n_352),
.C(n_356),
.Y(n_380)
);

NOR2xp33_ASAP7_75t_SL g351 ( 
.A(n_339),
.B(n_321),
.Y(n_351)
);

CKINVDCx14_ASAP7_75t_R g392 ( 
.A(n_351),
.Y(n_392)
);

MAJIxp5_ASAP7_75t_L g352 ( 
.A(n_314),
.B(n_290),
.C(n_291),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_353),
.B(n_360),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_L g354 ( 
.A(n_329),
.B(n_306),
.Y(n_354)
);

CKINVDCx16_ASAP7_75t_R g385 ( 
.A(n_354),
.Y(n_385)
);

NOR2xp33_ASAP7_75t_L g355 ( 
.A(n_339),
.B(n_265),
.Y(n_355)
);

NOR2xp33_ASAP7_75t_SL g376 ( 
.A(n_355),
.B(n_363),
.Y(n_376)
);

XNOR2xp5_ASAP7_75t_L g356 ( 
.A(n_317),
.B(n_302),
.Y(n_356)
);

OAI21xp5_ASAP7_75t_L g357 ( 
.A1(n_320),
.A2(n_305),
.B(n_296),
.Y(n_357)
);

OAI21xp5_ASAP7_75t_L g386 ( 
.A1(n_357),
.A2(n_342),
.B(n_340),
.Y(n_386)
);

OAI22xp5_ASAP7_75t_SL g358 ( 
.A1(n_313),
.A2(n_294),
.B1(n_275),
.B2(n_279),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_310),
.Y(n_359)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_359),
.Y(n_381)
);

CKINVDCx20_ASAP7_75t_R g360 ( 
.A(n_322),
.Y(n_360)
);

OAI22xp5_ASAP7_75t_SL g362 ( 
.A1(n_312),
.A2(n_319),
.B1(n_317),
.B2(n_330),
.Y(n_362)
);

NOR2xp33_ASAP7_75t_L g363 ( 
.A(n_324),
.B(n_330),
.Y(n_363)
);

CKINVDCx20_ASAP7_75t_R g364 ( 
.A(n_335),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_364),
.B(n_368),
.Y(n_378)
);

HB1xp67_ASAP7_75t_L g365 ( 
.A(n_315),
.Y(n_365)
);

INVxp67_ASAP7_75t_L g377 ( 
.A(n_365),
.Y(n_377)
);

OAI22xp5_ASAP7_75t_SL g366 ( 
.A1(n_337),
.A2(n_282),
.B1(n_281),
.B2(n_280),
.Y(n_366)
);

AND2x2_ASAP7_75t_L g367 ( 
.A(n_336),
.B(n_286),
.Y(n_367)
);

INVxp67_ASAP7_75t_L g388 ( 
.A(n_367),
.Y(n_388)
);

CKINVDCx20_ASAP7_75t_R g368 ( 
.A(n_316),
.Y(n_368)
);

OAI22xp5_ASAP7_75t_SL g369 ( 
.A1(n_337),
.A2(n_299),
.B1(n_283),
.B2(n_251),
.Y(n_369)
);

AOI22xp5_ASAP7_75t_L g394 ( 
.A1(n_369),
.A2(n_332),
.B1(n_333),
.B2(n_338),
.Y(n_394)
);

AOI32xp33_ASAP7_75t_L g370 ( 
.A1(n_334),
.A2(n_181),
.A3(n_186),
.B1(n_268),
.B2(n_273),
.Y(n_370)
);

NOR2xp33_ASAP7_75t_SL g391 ( 
.A(n_370),
.B(n_357),
.Y(n_391)
);

OAI22xp5_ASAP7_75t_SL g382 ( 
.A1(n_371),
.A2(n_341),
.B1(n_325),
.B2(n_323),
.Y(n_382)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_310),
.Y(n_372)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_372),
.Y(n_396)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_326),
.Y(n_374)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_374),
.Y(n_399)
);

HB1xp67_ASAP7_75t_L g379 ( 
.A(n_348),
.Y(n_379)
);

NOR2xp33_ASAP7_75t_L g422 ( 
.A(n_379),
.B(n_368),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_382),
.B(n_358),
.Y(n_408)
);

XOR2xp5_ASAP7_75t_L g425 ( 
.A(n_383),
.B(n_384),
.Y(n_425)
);

XOR2xp5_ASAP7_75t_L g384 ( 
.A(n_350),
.B(n_342),
.Y(n_384)
);

AOI21xp5_ASAP7_75t_L g416 ( 
.A1(n_386),
.A2(n_400),
.B(n_404),
.Y(n_416)
);

OAI22xp5_ASAP7_75t_SL g387 ( 
.A1(n_371),
.A2(n_316),
.B1(n_327),
.B2(n_326),
.Y(n_387)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_387),
.Y(n_411)
);

AOI22xp5_ASAP7_75t_SL g389 ( 
.A1(n_349),
.A2(n_343),
.B1(n_361),
.B2(n_367),
.Y(n_389)
);

OAI22xp5_ASAP7_75t_L g424 ( 
.A1(n_389),
.A2(n_394),
.B1(n_348),
.B2(n_374),
.Y(n_424)
);

CKINVDCx14_ASAP7_75t_R g410 ( 
.A(n_391),
.Y(n_410)
);

MAJIxp5_ASAP7_75t_L g393 ( 
.A(n_356),
.B(n_327),
.C(n_315),
.Y(n_393)
);

MAJIxp5_ASAP7_75t_L g423 ( 
.A(n_393),
.B(n_398),
.C(n_402),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_345),
.B(n_360),
.Y(n_395)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_395),
.Y(n_415)
);

OAI21xp33_ASAP7_75t_L g397 ( 
.A1(n_373),
.A2(n_333),
.B(n_340),
.Y(n_397)
);

BUFx12_ASAP7_75t_L g414 ( 
.A(n_397),
.Y(n_414)
);

MAJIxp5_ASAP7_75t_L g398 ( 
.A(n_346),
.B(n_338),
.C(n_332),
.Y(n_398)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_359),
.Y(n_401)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_401),
.Y(n_417)
);

MAJIxp5_ASAP7_75t_L g402 ( 
.A(n_352),
.B(n_318),
.C(n_268),
.Y(n_402)
);

AOI21xp5_ASAP7_75t_L g404 ( 
.A1(n_367),
.A2(n_286),
.B(n_155),
.Y(n_404)
);

MAJIxp5_ASAP7_75t_L g405 ( 
.A(n_362),
.B(n_268),
.C(n_172),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_SL g429 ( 
.A(n_405),
.B(n_398),
.Y(n_429)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_372),
.Y(n_406)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_406),
.Y(n_419)
);

XNOR2xp5_ASAP7_75t_L g407 ( 
.A(n_384),
.B(n_344),
.Y(n_407)
);

MAJIxp5_ASAP7_75t_L g441 ( 
.A(n_407),
.B(n_423),
.C(n_380),
.Y(n_441)
);

OAI22xp5_ASAP7_75t_SL g455 ( 
.A1(n_408),
.A2(n_265),
.B1(n_249),
.B2(n_26),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_395),
.B(n_344),
.Y(n_409)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_409),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_SL g412 ( 
.A(n_392),
.B(n_364),
.Y(n_412)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_412),
.Y(n_440)
);

INVxp67_ASAP7_75t_SL g413 ( 
.A(n_378),
.Y(n_413)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_413),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_L g418 ( 
.A(n_378),
.B(n_353),
.Y(n_418)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_418),
.Y(n_456)
);

AOI21xp5_ASAP7_75t_L g420 ( 
.A1(n_388),
.A2(n_361),
.B(n_343),
.Y(n_420)
);

CKINVDCx20_ASAP7_75t_R g453 ( 
.A(n_420),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_375),
.B(n_366),
.Y(n_421)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_421),
.Y(n_457)
);

OAI22xp5_ASAP7_75t_L g442 ( 
.A1(n_422),
.A2(n_431),
.B1(n_434),
.B2(n_435),
.Y(n_442)
);

AOI22xp5_ASAP7_75t_L g436 ( 
.A1(n_424),
.A2(n_382),
.B1(n_387),
.B2(n_383),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_375),
.B(n_369),
.Y(n_426)
);

XOR2xp5_ASAP7_75t_L g443 ( 
.A(n_426),
.B(n_427),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_377),
.B(n_286),
.Y(n_427)
);

INVxp33_ASAP7_75t_L g428 ( 
.A(n_376),
.Y(n_428)
);

INVx2_ASAP7_75t_SL g454 ( 
.A(n_428),
.Y(n_454)
);

XOR2xp5_ASAP7_75t_L g445 ( 
.A(n_429),
.B(n_430),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_377),
.B(n_1),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_403),
.Y(n_431)
);

XOR2xp5_ASAP7_75t_L g432 ( 
.A(n_380),
.B(n_249),
.Y(n_432)
);

XOR2xp5_ASAP7_75t_L g449 ( 
.A(n_432),
.B(n_433),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_385),
.B(n_1),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_SL g434 ( 
.A(n_386),
.B(n_3),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_403),
.Y(n_435)
);

XOR2xp5_ASAP7_75t_L g468 ( 
.A(n_436),
.B(n_408),
.Y(n_468)
);

AOI22xp5_ASAP7_75t_L g438 ( 
.A1(n_424),
.A2(n_400),
.B1(n_388),
.B2(n_390),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_438),
.B(n_439),
.Y(n_469)
);

AOI22xp5_ASAP7_75t_L g439 ( 
.A1(n_411),
.A2(n_390),
.B1(n_405),
.B2(n_389),
.Y(n_439)
);

XNOR2xp5_ASAP7_75t_L g459 ( 
.A(n_441),
.B(n_409),
.Y(n_459)
);

NAND3xp33_ASAP7_75t_L g444 ( 
.A(n_410),
.B(n_406),
.C(n_381),
.Y(n_444)
);

CKINVDCx14_ASAP7_75t_R g463 ( 
.A(n_444),
.Y(n_463)
);

MAJIxp5_ASAP7_75t_L g447 ( 
.A(n_423),
.B(n_393),
.C(n_402),
.Y(n_447)
);

MAJIxp5_ASAP7_75t_L g461 ( 
.A(n_447),
.B(n_451),
.C(n_452),
.Y(n_461)
);

AOI22xp5_ASAP7_75t_L g448 ( 
.A1(n_411),
.A2(n_404),
.B1(n_401),
.B2(n_399),
.Y(n_448)
);

NOR2xp33_ASAP7_75t_L g467 ( 
.A(n_448),
.B(n_450),
.Y(n_467)
);

AOI22xp5_ASAP7_75t_L g450 ( 
.A1(n_415),
.A2(n_399),
.B1(n_396),
.B2(n_381),
.Y(n_450)
);

MAJIxp5_ASAP7_75t_L g451 ( 
.A(n_432),
.B(n_394),
.C(n_396),
.Y(n_451)
);

MAJIxp5_ASAP7_75t_L g452 ( 
.A(n_425),
.B(n_407),
.C(n_415),
.Y(n_452)
);

AOI22xp5_ASAP7_75t_L g460 ( 
.A1(n_455),
.A2(n_435),
.B1(n_431),
.B2(n_419),
.Y(n_460)
);

MAJIxp5_ASAP7_75t_L g458 ( 
.A(n_425),
.B(n_249),
.C(n_26),
.Y(n_458)
);

MAJIxp5_ASAP7_75t_L g464 ( 
.A(n_458),
.B(n_427),
.C(n_416),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_L g490 ( 
.A(n_459),
.B(n_464),
.Y(n_490)
);

OAI22xp5_ASAP7_75t_SL g484 ( 
.A1(n_460),
.A2(n_475),
.B1(n_419),
.B2(n_417),
.Y(n_484)
);

XNOR2x1_ASAP7_75t_L g462 ( 
.A(n_451),
.B(n_421),
.Y(n_462)
);

XNOR2xp5_ASAP7_75t_SL g479 ( 
.A(n_462),
.B(n_474),
.Y(n_479)
);

HB1xp67_ASAP7_75t_L g465 ( 
.A(n_440),
.Y(n_465)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_465),
.Y(n_485)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_450),
.Y(n_466)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_466),
.Y(n_489)
);

XOR2xp5_ASAP7_75t_L g483 ( 
.A(n_468),
.B(n_476),
.Y(n_483)
);

NOR2xp33_ASAP7_75t_SL g470 ( 
.A(n_454),
.B(n_412),
.Y(n_470)
);

CKINVDCx16_ASAP7_75t_R g492 ( 
.A(n_470),
.Y(n_492)
);

AOI21xp33_ASAP7_75t_L g471 ( 
.A1(n_446),
.A2(n_418),
.B(n_414),
.Y(n_471)
);

AOI21xp5_ASAP7_75t_L g493 ( 
.A1(n_471),
.A2(n_477),
.B(n_434),
.Y(n_493)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_442),
.Y(n_472)
);

HB1xp67_ASAP7_75t_L g491 ( 
.A(n_472),
.Y(n_491)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_437),
.Y(n_473)
);

CKINVDCx14_ASAP7_75t_R g481 ( 
.A(n_473),
.Y(n_481)
);

XOR2x2_ASAP7_75t_L g474 ( 
.A(n_443),
.B(n_416),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_456),
.Y(n_475)
);

XNOR2xp5_ASAP7_75t_SL g476 ( 
.A(n_449),
.B(n_452),
.Y(n_476)
);

OAI21xp5_ASAP7_75t_SL g477 ( 
.A1(n_454),
.A2(n_420),
.B(n_426),
.Y(n_477)
);

AOI22xp5_ASAP7_75t_L g478 ( 
.A1(n_468),
.A2(n_457),
.B1(n_453),
.B2(n_443),
.Y(n_478)
);

OAI22xp5_ASAP7_75t_SL g495 ( 
.A1(n_478),
.A2(n_482),
.B1(n_464),
.B2(n_474),
.Y(n_495)
);

BUFx24_ASAP7_75t_SL g480 ( 
.A(n_463),
.Y(n_480)
);

NOR2xp33_ASAP7_75t_SL g502 ( 
.A(n_480),
.B(n_494),
.Y(n_502)
);

AOI22xp5_ASAP7_75t_L g482 ( 
.A1(n_467),
.A2(n_445),
.B1(n_439),
.B2(n_436),
.Y(n_482)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_484),
.Y(n_499)
);

MAJx2_ASAP7_75t_L g486 ( 
.A(n_461),
.B(n_447),
.C(n_441),
.Y(n_486)
);

XNOR2xp5_ASAP7_75t_SL g496 ( 
.A(n_486),
.B(n_493),
.Y(n_496)
);

MAJIxp5_ASAP7_75t_L g487 ( 
.A(n_459),
.B(n_445),
.C(n_449),
.Y(n_487)
);

MAJIxp5_ASAP7_75t_L g508 ( 
.A(n_487),
.B(n_26),
.C(n_6),
.Y(n_508)
);

OAI22xp5_ASAP7_75t_SL g488 ( 
.A1(n_469),
.A2(n_438),
.B1(n_460),
.B2(n_448),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_SL g507 ( 
.A(n_488),
.B(n_3),
.Y(n_507)
);

FAx1_ASAP7_75t_SL g494 ( 
.A(n_469),
.B(n_414),
.CI(n_433),
.CON(n_494),
.SN(n_494)
);

NAND2xp5_ASAP7_75t_L g511 ( 
.A(n_495),
.B(n_497),
.Y(n_511)
);

NOR2xp33_ASAP7_75t_L g497 ( 
.A(n_492),
.B(n_414),
.Y(n_497)
);

XOR2xp5_ASAP7_75t_L g498 ( 
.A(n_483),
.B(n_462),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_L g512 ( 
.A(n_498),
.B(n_500),
.Y(n_512)
);

XOR2xp5_ASAP7_75t_L g500 ( 
.A(n_483),
.B(n_461),
.Y(n_500)
);

MAJx2_ASAP7_75t_L g501 ( 
.A(n_487),
.B(n_477),
.C(n_476),
.Y(n_501)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_501),
.Y(n_515)
);

OAI22xp5_ASAP7_75t_SL g503 ( 
.A1(n_482),
.A2(n_417),
.B1(n_414),
.B2(n_430),
.Y(n_503)
);

AOI22xp5_ASAP7_75t_SL g513 ( 
.A1(n_503),
.A2(n_481),
.B1(n_489),
.B2(n_491),
.Y(n_513)
);

NOR2xp67_ASAP7_75t_SL g504 ( 
.A(n_479),
.B(n_458),
.Y(n_504)
);

AOI21xp5_ASAP7_75t_L g519 ( 
.A1(n_504),
.A2(n_506),
.B(n_3),
.Y(n_519)
);

XNOR2xp5_ASAP7_75t_L g505 ( 
.A(n_486),
.B(n_455),
.Y(n_505)
);

NOR2xp33_ASAP7_75t_L g510 ( 
.A(n_505),
.B(n_509),
.Y(n_510)
);

MAJIxp5_ASAP7_75t_L g506 ( 
.A(n_490),
.B(n_249),
.C(n_26),
.Y(n_506)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_507),
.Y(n_516)
);

MAJx2_ASAP7_75t_L g518 ( 
.A(n_508),
.B(n_494),
.C(n_479),
.Y(n_518)
);

NOR2xp33_ASAP7_75t_L g509 ( 
.A(n_494),
.B(n_3),
.Y(n_509)
);

XNOR2xp5_ASAP7_75t_L g521 ( 
.A(n_513),
.B(n_518),
.Y(n_521)
);

BUFx6f_ASAP7_75t_L g514 ( 
.A(n_496),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_SL g524 ( 
.A(n_514),
.B(n_498),
.Y(n_524)
);

OAI22xp5_ASAP7_75t_L g517 ( 
.A1(n_502),
.A2(n_499),
.B1(n_478),
.B2(n_485),
.Y(n_517)
);

AOI22xp5_ASAP7_75t_L g525 ( 
.A1(n_517),
.A2(n_520),
.B1(n_7),
.B2(n_8),
.Y(n_525)
);

XNOR2xp5_ASAP7_75t_L g526 ( 
.A(n_519),
.B(n_7),
.Y(n_526)
);

INVxp33_ASAP7_75t_L g520 ( 
.A(n_496),
.Y(n_520)
);

XOR2xp5_ASAP7_75t_L g522 ( 
.A(n_512),
.B(n_501),
.Y(n_522)
);

MAJIxp5_ASAP7_75t_L g528 ( 
.A(n_522),
.B(n_523),
.C(n_525),
.Y(n_528)
);

OAI21xp5_ASAP7_75t_SL g523 ( 
.A1(n_515),
.A2(n_500),
.B(n_508),
.Y(n_523)
);

OAI21xp5_ASAP7_75t_L g529 ( 
.A1(n_524),
.A2(n_526),
.B(n_527),
.Y(n_529)
);

XNOR2xp5_ASAP7_75t_L g527 ( 
.A(n_511),
.B(n_26),
.Y(n_527)
);

OAI21xp5_ASAP7_75t_SL g530 ( 
.A1(n_522),
.A2(n_510),
.B(n_514),
.Y(n_530)
);

O2A1O1Ixp33_ASAP7_75t_SL g533 ( 
.A1(n_530),
.A2(n_528),
.B(n_529),
.C(n_9),
.Y(n_533)
);

OAI21xp5_ASAP7_75t_L g531 ( 
.A1(n_521),
.A2(n_510),
.B(n_516),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_L g532 ( 
.A(n_531),
.B(n_521),
.Y(n_532)
);

OAI21x1_ASAP7_75t_L g535 ( 
.A1(n_532),
.A2(n_533),
.B(n_534),
.Y(n_535)
);

INVxp67_ASAP7_75t_L g534 ( 
.A(n_531),
.Y(n_534)
);

AOI22xp5_ASAP7_75t_L g536 ( 
.A1(n_535),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_L g537 ( 
.A(n_536),
.B(n_9),
.Y(n_537)
);

OAI221xp5_ASAP7_75t_L g538 ( 
.A1(n_537),
.A2(n_10),
.B1(n_11),
.B2(n_13),
.C(n_536),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_L g539 ( 
.A(n_538),
.B(n_11),
.Y(n_539)
);

XOR2xp5_ASAP7_75t_L g540 ( 
.A(n_539),
.B(n_11),
.Y(n_540)
);


endmodule