module fake_jpeg_24923_n_64 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_7, n_64);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;
input n_7;

output n_64;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_55;
wire n_22;
wire n_51;
wire n_47;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_59;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_62;
wire n_17;
wire n_25;
wire n_31;
wire n_56;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_8;
wire n_15;

BUFx6f_ASAP7_75t_L g8 ( 
.A(n_0),
.Y(n_8)
);

CKINVDCx20_ASAP7_75t_R g9 ( 
.A(n_1),
.Y(n_9)
);

INVx3_ASAP7_75t_L g10 ( 
.A(n_4),
.Y(n_10)
);

BUFx6f_ASAP7_75t_L g11 ( 
.A(n_6),
.Y(n_11)
);

INVx6_ASAP7_75t_L g12 ( 
.A(n_4),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_2),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_5),
.Y(n_14)
);

INVx11_ASAP7_75t_L g15 ( 
.A(n_0),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

INVx11_ASAP7_75t_L g17 ( 
.A(n_15),
.Y(n_17)
);

AOI22xp33_ASAP7_75t_SL g25 ( 
.A1(n_17),
.A2(n_19),
.B1(n_12),
.B2(n_15),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_18),
.Y(n_26)
);

AOI22xp33_ASAP7_75t_SL g19 ( 
.A1(n_12),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_10),
.B(n_3),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_20),
.B(n_16),
.Y(n_23)
);

A2O1A1Ixp33_ASAP7_75t_L g21 ( 
.A1(n_11),
.A2(n_3),
.B(n_5),
.C(n_6),
.Y(n_21)
);

NOR2x1_ASAP7_75t_L g24 ( 
.A(n_21),
.B(n_10),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_20),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_SL g27 ( 
.A(n_22),
.B(n_23),
.Y(n_27)
);

INVx2_ASAP7_75t_R g30 ( 
.A(n_24),
.Y(n_30)
);

OAI22xp33_ASAP7_75t_SL g34 ( 
.A1(n_25),
.A2(n_15),
.B1(n_17),
.B2(n_11),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_22),
.B(n_21),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_SL g43 ( 
.A(n_28),
.B(n_31),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_SL g29 ( 
.A1(n_24),
.A2(n_17),
.B1(n_12),
.B2(n_10),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_SL g37 ( 
.A1(n_29),
.A2(n_34),
.B1(n_16),
.B2(n_9),
.Y(n_37)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_23),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_26),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_32),
.B(n_33),
.Y(n_36)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_26),
.Y(n_33)
);

CKINVDCx16_ASAP7_75t_R g35 ( 
.A(n_26),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_35),
.B(n_9),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_SL g46 ( 
.A1(n_37),
.A2(n_14),
.B1(n_32),
.B2(n_8),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_38),
.Y(n_47)
);

OR2x2_ASAP7_75t_L g39 ( 
.A(n_30),
.B(n_13),
.Y(n_39)
);

AND2x2_ASAP7_75t_SL g48 ( 
.A(n_39),
.B(n_7),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_31),
.B(n_13),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_SL g45 ( 
.A(n_40),
.B(n_41),
.Y(n_45)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_33),
.Y(n_41)
);

MAJIxp5_ASAP7_75t_L g42 ( 
.A(n_29),
.B(n_18),
.C(n_14),
.Y(n_42)
);

MAJIxp5_ASAP7_75t_L g44 ( 
.A(n_42),
.B(n_30),
.C(n_27),
.Y(n_44)
);

MAJIxp5_ASAP7_75t_L g52 ( 
.A(n_44),
.B(n_48),
.C(n_49),
.Y(n_52)
);

XOR2xp5_ASAP7_75t_L g54 ( 
.A(n_46),
.B(n_37),
.Y(n_54)
);

MAJIxp5_ASAP7_75t_L g49 ( 
.A(n_43),
.B(n_18),
.C(n_8),
.Y(n_49)
);

BUFx2_ASAP7_75t_L g50 ( 
.A(n_45),
.Y(n_50)
);

CKINVDCx16_ASAP7_75t_R g56 ( 
.A(n_50),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_45),
.Y(n_51)
);

CKINVDCx16_ASAP7_75t_R g57 ( 
.A(n_51),
.Y(n_57)
);

AOI21xp5_ASAP7_75t_L g53 ( 
.A1(n_47),
.A2(n_42),
.B(n_39),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_53),
.A2(n_54),
.B1(n_48),
.B2(n_36),
.Y(n_55)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_55),
.Y(n_58)
);

AOI21xp5_ASAP7_75t_L g59 ( 
.A1(n_56),
.A2(n_50),
.B(n_52),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_59),
.B(n_57),
.Y(n_60)
);

INVxp67_ASAP7_75t_L g62 ( 
.A(n_60),
.Y(n_62)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_58),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_62),
.B(n_61),
.Y(n_63)
);

XNOR2xp5_ASAP7_75t_L g64 ( 
.A(n_63),
.B(n_41),
.Y(n_64)
);


endmodule