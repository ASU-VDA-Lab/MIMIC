module real_jpeg_24070_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_78;
wire n_83;
wire n_249;
wire n_166;
wire n_176;
wire n_215;
wire n_300;
wire n_292;
wire n_221;
wire n_286;
wire n_288;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_301;
wire n_280;
wire n_64;
wire n_177;
wire n_291;
wire n_236;
wire n_131;
wire n_47;
wire n_271;
wire n_281;
wire n_163;
wire n_276;
wire n_22;
wire n_287;
wire n_174;
wire n_237;
wire n_87;
wire n_255;
wire n_105;
wire n_40;
wire n_243;
wire n_173;
wire n_197;
wire n_115;
wire n_299;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_293;
wire n_275;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_242;
wire n_141;
wire n_139;
wire n_33;
wire n_65;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_282;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_290;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_285;
wire n_268;
wire n_42;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_148;
wire n_19;
wire n_222;
wire n_262;
wire n_118;
wire n_220;
wire n_294;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_298;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_296;
wire n_134;
wire n_270;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_192;
wire n_203;
wire n_100;
wire n_198;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_205;
wire n_258;
wire n_289;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_228;
wire n_150;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_278;
wire n_241;
wire n_103;
wire n_225;
wire n_259;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_284;
wire n_226;
wire n_277;
wire n_125;
wire n_185;
wire n_297;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_240;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_169;
wire n_88;
wire n_59;
wire n_279;
wire n_128;
wire n_244;
wire n_167;
wire n_179;
wire n_202;
wire n_213;
wire n_133;
wire n_216;
wire n_295;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_210;
wire n_127;
wire n_206;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_283;
wire n_101;
wire n_256;
wire n_274;
wire n_182;
wire n_273;
wire n_96;
wire n_253;
wire n_269;
wire n_89;

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_0),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g35 ( 
.A1(n_1),
.A2(n_28),
.B1(n_30),
.B2(n_36),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_1),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_1),
.A2(n_36),
.B1(n_74),
.B2(n_75),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_1),
.A2(n_36),
.B1(n_61),
.B2(n_62),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_1),
.A2(n_36),
.B1(n_41),
.B2(n_42),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g52 ( 
.A1(n_2),
.A2(n_41),
.B1(n_42),
.B2(n_53),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_2),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_2),
.A2(n_28),
.B1(n_30),
.B2(n_53),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_2),
.A2(n_53),
.B1(n_61),
.B2(n_62),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_3),
.A2(n_68),
.B1(n_174),
.B2(n_175),
.Y(n_173)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_3),
.Y(n_175)
);

AOI22xp33_ASAP7_75t_L g210 ( 
.A1(n_3),
.A2(n_61),
.B1(n_62),
.B2(n_175),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_L g226 ( 
.A1(n_3),
.A2(n_41),
.B1(n_42),
.B2(n_175),
.Y(n_226)
);

AOI22xp33_ASAP7_75t_L g251 ( 
.A1(n_3),
.A2(n_28),
.B1(n_30),
.B2(n_175),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_4),
.A2(n_66),
.B1(n_69),
.B2(n_71),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_4),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_4),
.A2(n_61),
.B1(n_62),
.B2(n_71),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_4),
.A2(n_28),
.B1(n_30),
.B2(n_71),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_L g268 ( 
.A1(n_4),
.A2(n_41),
.B1(n_42),
.B2(n_71),
.Y(n_268)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_5),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_6),
.A2(n_114),
.B1(n_115),
.B2(n_116),
.Y(n_113)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_6),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_6),
.A2(n_61),
.B1(n_62),
.B2(n_116),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_L g234 ( 
.A1(n_6),
.A2(n_41),
.B1(n_42),
.B2(n_116),
.Y(n_234)
);

AOI22xp33_ASAP7_75t_L g242 ( 
.A1(n_6),
.A2(n_28),
.B1(n_30),
.B2(n_116),
.Y(n_242)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

INVx8_ASAP7_75t_SL g60 ( 
.A(n_8),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_SL g26 ( 
.A1(n_9),
.A2(n_27),
.B1(n_28),
.B2(n_30),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_9),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_9),
.A2(n_27),
.B1(n_61),
.B2(n_62),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_9),
.A2(n_27),
.B1(n_41),
.B2(n_42),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_9),
.A2(n_27),
.B1(n_66),
.B2(n_115),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_SL g40 ( 
.A1(n_10),
.A2(n_41),
.B1(n_42),
.B2(n_44),
.Y(n_40)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_10),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_10),
.A2(n_44),
.B1(n_61),
.B2(n_62),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_L g170 ( 
.A1(n_10),
.A2(n_28),
.B1(n_30),
.B2(n_44),
.Y(n_170)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_11),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_11),
.B(n_76),
.Y(n_211)
);

AOI22xp33_ASAP7_75t_L g224 ( 
.A1(n_11),
.A2(n_41),
.B1(n_42),
.B2(n_165),
.Y(n_224)
);

AOI21xp5_ASAP7_75t_L g228 ( 
.A1(n_11),
.A2(n_28),
.B(n_48),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_11),
.B(n_121),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_11),
.A2(n_89),
.B1(n_90),
.B2(n_251),
.Y(n_253)
);

AOI21xp5_ASAP7_75t_L g264 ( 
.A1(n_11),
.A2(n_61),
.B(n_265),
.Y(n_264)
);

BUFx12f_ASAP7_75t_L g79 ( 
.A(n_12),
.Y(n_79)
);

INVx13_ASAP7_75t_L g68 ( 
.A(n_13),
.Y(n_68)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_14),
.Y(n_43)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_15),
.Y(n_38)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_15),
.Y(n_90)
);

INVx6_ASAP7_75t_L g108 ( 
.A(n_15),
.Y(n_108)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_148),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_SL g17 ( 
.A(n_18),
.B(n_146),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_122),
.Y(n_19)
);

AND2x2_ASAP7_75t_L g147 ( 
.A(n_20),
.B(n_122),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_87),
.C(n_98),
.Y(n_20)
);

FAx1_ASAP7_75t_SL g178 ( 
.A(n_21),
.B(n_87),
.CI(n_98),
.CON(n_178),
.SN(n_178)
);

AOI22xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_23),
.B1(n_54),
.B2(n_86),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_22),
.B(n_55),
.C(n_77),
.Y(n_145)
);

CKINVDCx14_ASAP7_75t_R g22 ( 
.A(n_23),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_39),
.Y(n_23)
);

XOR2xp5_ASAP7_75t_L g156 ( 
.A(n_24),
.B(n_39),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_34),
.Y(n_24)
);

OAI21xp5_ASAP7_75t_L g213 ( 
.A1(n_25),
.A2(n_108),
.B(n_170),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_SL g25 ( 
.A(n_26),
.B(n_31),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_26),
.B(n_105),
.Y(n_104)
);

INVx5_ASAP7_75t_L g30 ( 
.A(n_28),
.Y(n_30)
);

AOI22xp5_ASAP7_75t_L g51 ( 
.A1(n_28),
.A2(n_30),
.B1(n_48),
.B2(n_50),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_30),
.B(n_32),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_SL g254 ( 
.A(n_30),
.B(n_255),
.Y(n_254)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_31),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_31),
.A2(n_103),
.B1(n_169),
.B2(n_171),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_31),
.A2(n_241),
.B1(n_243),
.B2(n_244),
.Y(n_240)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

OAI21xp5_ASAP7_75t_L g236 ( 
.A1(n_34),
.A2(n_89),
.B(n_237),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g34 ( 
.A(n_35),
.B(n_37),
.Y(n_34)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_35),
.Y(n_91)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_38),
.A2(n_89),
.B1(n_242),
.B2(n_251),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_L g39 ( 
.A1(n_40),
.A2(n_45),
.B1(n_51),
.B2(n_52),
.Y(n_39)
);

OAI21xp5_ASAP7_75t_L g109 ( 
.A1(n_40),
.A2(n_51),
.B(n_110),
.Y(n_109)
);

OAI22xp33_ASAP7_75t_L g47 ( 
.A1(n_41),
.A2(n_42),
.B1(n_48),
.B2(n_50),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_41),
.A2(n_42),
.B1(n_79),
.B2(n_80),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_SL g273 ( 
.A(n_41),
.B(n_80),
.Y(n_273)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

A2O1A1Ixp33_ASAP7_75t_SL g227 ( 
.A1(n_42),
.A2(n_50),
.B(n_165),
.C(n_228),
.Y(n_227)
);

OAI32xp33_ASAP7_75t_L g272 ( 
.A1(n_42),
.A2(n_61),
.A3(n_79),
.B1(n_266),
.B2(n_273),
.Y(n_272)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

OAI21xp5_ASAP7_75t_SL g93 ( 
.A1(n_45),
.A2(n_52),
.B(n_94),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g223 ( 
.A1(n_45),
.A2(n_51),
.B1(n_224),
.B2(n_225),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_SL g288 ( 
.A1(n_45),
.A2(n_129),
.B(n_289),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_46),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_46),
.B(n_111),
.Y(n_110)
);

AOI21xp5_ASAP7_75t_L g188 ( 
.A1(n_46),
.A2(n_95),
.B(n_130),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_46),
.A2(n_131),
.B1(n_226),
.B2(n_234),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_46),
.A2(n_131),
.B1(n_234),
.B2(n_268),
.Y(n_267)
);

AND2x2_ASAP7_75t_L g46 ( 
.A(n_47),
.B(n_51),
.Y(n_46)
);

INVx13_ASAP7_75t_L g50 ( 
.A(n_48),
.Y(n_50)
);

BUFx24_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_51),
.B(n_96),
.Y(n_95)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_51),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_SL g249 ( 
.A(n_51),
.B(n_165),
.Y(n_249)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_54),
.Y(n_86)
);

XNOR2xp5_ASAP7_75t_SL g54 ( 
.A(n_55),
.B(n_77),
.Y(n_54)
);

OAI21xp5_ASAP7_75t_SL g55 ( 
.A1(n_56),
.A2(n_70),
.B(n_72),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_56),
.A2(n_57),
.B1(n_70),
.B2(n_113),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_SL g138 ( 
.A1(n_56),
.A2(n_139),
.B(n_140),
.Y(n_138)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_56),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g56 ( 
.A(n_57),
.B(n_65),
.Y(n_56)
);

CKINVDCx16_ASAP7_75t_R g76 ( 
.A(n_57),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g57 ( 
.A1(n_58),
.A2(n_59),
.B1(n_61),
.B2(n_62),
.Y(n_57)
);

OAI22xp33_ASAP7_75t_L g65 ( 
.A1(n_58),
.A2(n_59),
.B1(n_66),
.B2(n_69),
.Y(n_65)
);

OAI32xp33_ASAP7_75t_L g163 ( 
.A1(n_58),
.A2(n_62),
.A3(n_68),
.B1(n_164),
.B2(n_166),
.Y(n_163)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_59),
.B(n_61),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_61),
.A2(n_62),
.B1(n_79),
.B2(n_80),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_62),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_62),
.B(n_165),
.Y(n_266)
);

BUFx12f_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx8_ASAP7_75t_L g174 ( 
.A(n_66),
.Y(n_174)
);

INVx8_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx8_ASAP7_75t_L g69 ( 
.A(n_68),
.Y(n_69)
);

INVx11_ASAP7_75t_L g74 ( 
.A(n_68),
.Y(n_74)
);

INVx8_ASAP7_75t_L g115 ( 
.A(n_68),
.Y(n_115)
);

OAI21xp33_ASAP7_75t_L g190 ( 
.A1(n_69),
.A2(n_164),
.B(n_165),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_73),
.B(n_76),
.Y(n_72)
);

CKINVDCx16_ASAP7_75t_R g139 ( 
.A(n_73),
.Y(n_139)
);

INVx8_ASAP7_75t_L g75 ( 
.A(n_74),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_74),
.B(n_165),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_76),
.B(n_141),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_76),
.A2(n_173),
.B1(n_176),
.B2(n_177),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_76),
.A2(n_173),
.B1(n_176),
.B2(n_190),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_L g77 ( 
.A1(n_78),
.A2(n_81),
.B(n_82),
.Y(n_77)
);

AND2x2_ASAP7_75t_L g83 ( 
.A(n_78),
.B(n_84),
.Y(n_83)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_78),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_78),
.B(n_119),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g263 ( 
.A1(n_78),
.A2(n_118),
.B1(n_210),
.B2(n_264),
.Y(n_263)
);

INVx5_ASAP7_75t_L g80 ( 
.A(n_79),
.Y(n_80)
);

CKINVDCx14_ASAP7_75t_R g126 ( 
.A(n_81),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_83),
.B(n_85),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_83),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_83),
.A2(n_121),
.B1(n_126),
.B2(n_127),
.Y(n_125)
);

AOI21xp5_ASAP7_75t_L g159 ( 
.A1(n_83),
.A2(n_160),
.B(n_161),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_83),
.A2(n_121),
.B1(n_160),
.B2(n_192),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_83),
.A2(n_121),
.B1(n_192),
.B2(n_209),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_85),
.B(n_121),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_88),
.A2(n_92),
.B1(n_93),
.B2(n_97),
.Y(n_87)
);

CKINVDCx16_ASAP7_75t_R g97 ( 
.A(n_88),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_88),
.B(n_93),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_88),
.A2(n_97),
.B1(n_137),
.B2(n_138),
.Y(n_136)
);

AOI21xp5_ASAP7_75t_L g88 ( 
.A1(n_89),
.A2(n_90),
.B(n_91),
.Y(n_88)
);

OAI21xp5_ASAP7_75t_L g101 ( 
.A1(n_89),
.A2(n_102),
.B(n_104),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_L g274 ( 
.A1(n_89),
.A2(n_91),
.B(n_104),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_90),
.B(n_165),
.Y(n_255)
);

INVxp67_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVxp67_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_96),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_112),
.C(n_117),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_99),
.A2(n_100),
.B1(n_153),
.B2(n_154),
.Y(n_152)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_101),
.B(n_109),
.Y(n_100)
);

XOR2xp5_ASAP7_75t_L g193 ( 
.A(n_101),
.B(n_109),
.Y(n_193)
);

INVxp67_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx5_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

INVx8_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx5_ASAP7_75t_L g171 ( 
.A(n_108),
.Y(n_171)
);

INVx3_ASAP7_75t_SL g244 ( 
.A(n_108),
.Y(n_244)
);

AND2x2_ASAP7_75t_L g128 ( 
.A(n_110),
.B(n_129),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_SL g154 ( 
.A(n_112),
.B(n_117),
.Y(n_154)
);

CKINVDCx16_ASAP7_75t_R g177 ( 
.A(n_113),
.Y(n_177)
);

INVx4_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_SL g117 ( 
.A1(n_118),
.A2(n_119),
.B(n_120),
.Y(n_117)
);

XOR2xp5_ASAP7_75t_L g122 ( 
.A(n_123),
.B(n_145),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_124),
.A2(n_133),
.B1(n_143),
.B2(n_144),
.Y(n_123)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_124),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_L g124 ( 
.A1(n_125),
.A2(n_128),
.B(n_132),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_125),
.B(n_128),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_130),
.B(n_131),
.Y(n_129)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_133),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_134),
.A2(n_135),
.B1(n_136),
.B2(n_142),
.Y(n_133)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_136),
.Y(n_142)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

CKINVDCx16_ASAP7_75t_R g146 ( 
.A(n_147),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_L g148 ( 
.A1(n_149),
.A2(n_179),
.B(n_301),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_178),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g301 ( 
.A(n_150),
.B(n_178),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_155),
.C(n_157),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_151),
.A2(n_152),
.B1(n_155),
.B2(n_156),
.Y(n_195)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_157),
.A2(n_158),
.B1(n_195),
.B2(n_196),
.Y(n_194)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_162),
.C(n_172),
.Y(n_158)
);

XOR2xp5_ASAP7_75t_L g186 ( 
.A(n_159),
.B(n_172),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g185 ( 
.A(n_162),
.B(n_186),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_167),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_163),
.A2(n_167),
.B1(n_168),
.B2(n_205),
.Y(n_204)
);

CKINVDCx14_ASAP7_75t_R g205 ( 
.A(n_163),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_168),
.Y(n_167)
);

INVxp67_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

BUFx24_ASAP7_75t_SL g302 ( 
.A(n_178),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_215),
.Y(n_179)
);

INVxp33_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

AOI21xp33_ASAP7_75t_L g181 ( 
.A1(n_182),
.A2(n_197),
.B(n_214),
.Y(n_181)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_182),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_194),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_SL g214 ( 
.A(n_183),
.B(n_194),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_187),
.C(n_193),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_L g198 ( 
.A1(n_184),
.A2(n_185),
.B1(n_199),
.B2(n_200),
.Y(n_198)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_SL g200 ( 
.A(n_187),
.B(n_193),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_188),
.B(n_189),
.C(n_191),
.Y(n_187)
);

XOR2xp5_ASAP7_75t_L g203 ( 
.A(n_188),
.B(n_191),
.Y(n_203)
);

XOR2xp5_ASAP7_75t_L g202 ( 
.A(n_189),
.B(n_203),
.Y(n_202)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_195),
.Y(n_196)
);

AND2x2_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_201),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_198),
.B(n_201),
.Y(n_300)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_202),
.B(n_204),
.C(n_206),
.Y(n_201)
);

XOR2xp5_ASAP7_75t_L g295 ( 
.A(n_202),
.B(n_296),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_L g296 ( 
.A1(n_204),
.A2(n_206),
.B1(n_207),
.B2(n_297),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_204),
.Y(n_297)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_211),
.C(n_212),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_SL g282 ( 
.A(n_208),
.B(n_283),
.Y(n_282)
);

CKINVDCx14_ASAP7_75t_R g209 ( 
.A(n_210),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_211),
.A2(n_212),
.B1(n_213),
.B2(n_284),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_211),
.Y(n_284)
);

CKINVDCx16_ASAP7_75t_R g212 ( 
.A(n_213),
.Y(n_212)
);

NOR3xp33_ASAP7_75t_L g215 ( 
.A(n_216),
.B(n_299),
.C(n_300),
.Y(n_215)
);

AOI21xp5_ASAP7_75t_L g216 ( 
.A1(n_217),
.A2(n_293),
.B(n_298),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_SL g217 ( 
.A1(n_218),
.A2(n_278),
.B(n_292),
.Y(n_217)
);

AOI21xp5_ASAP7_75t_L g218 ( 
.A1(n_219),
.A2(n_259),
.B(n_277),
.Y(n_218)
);

OAI21xp5_ASAP7_75t_SL g219 ( 
.A1(n_220),
.A2(n_238),
.B(n_258),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_221),
.B(n_229),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_SL g258 ( 
.A(n_221),
.B(n_229),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_SL g221 ( 
.A(n_222),
.B(n_227),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_222),
.A2(n_223),
.B1(n_227),
.B2(n_246),
.Y(n_245)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

CKINVDCx16_ASAP7_75t_R g225 ( 
.A(n_226),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_227),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_230),
.B(n_236),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_231),
.A2(n_232),
.B1(n_233),
.B2(n_235),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_231),
.B(n_235),
.C(n_236),
.Y(n_260)
);

CKINVDCx14_ASAP7_75t_R g231 ( 
.A(n_232),
.Y(n_231)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_233),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_237),
.Y(n_243)
);

AOI21xp5_ASAP7_75t_L g238 ( 
.A1(n_239),
.A2(n_247),
.B(n_257),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_240),
.B(n_245),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_SL g257 ( 
.A(n_240),
.B(n_245),
.Y(n_257)
);

CKINVDCx16_ASAP7_75t_R g241 ( 
.A(n_242),
.Y(n_241)
);

OAI21xp5_ASAP7_75t_SL g247 ( 
.A1(n_248),
.A2(n_252),
.B(n_256),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_249),
.B(n_250),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_SL g256 ( 
.A(n_249),
.B(n_250),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_253),
.B(n_254),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_260),
.B(n_261),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_SL g277 ( 
.A(n_260),
.B(n_261),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_262),
.A2(n_271),
.B1(n_275),
.B2(n_276),
.Y(n_261)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_262),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_263),
.A2(n_267),
.B1(n_269),
.B2(n_270),
.Y(n_262)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_263),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_266),
.Y(n_265)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_267),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_267),
.B(n_270),
.C(n_275),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g289 ( 
.A(n_268),
.Y(n_289)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_271),
.Y(n_275)
);

XOR2xp5_ASAP7_75t_L g271 ( 
.A(n_272),
.B(n_274),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_272),
.B(n_274),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_279),
.B(n_280),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_SL g292 ( 
.A(n_279),
.B(n_280),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_281),
.A2(n_282),
.B1(n_285),
.B2(n_286),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_281),
.B(n_288),
.C(n_290),
.Y(n_294)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_SL g286 ( 
.A1(n_287),
.A2(n_288),
.B1(n_290),
.B2(n_291),
.Y(n_286)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_287),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_288),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_294),
.B(n_295),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_SL g298 ( 
.A(n_294),
.B(n_295),
.Y(n_298)
);


endmodule