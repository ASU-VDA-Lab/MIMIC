module real_jpeg_6267_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_384;
wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_50;
wire n_409;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_393;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_387;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_402;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_404;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_364;

INVx8_ASAP7_75t_L g45 ( 
.A(n_0),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_1),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_1),
.Y(n_111)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_1),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g156 ( 
.A(n_1),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g204 ( 
.A(n_1),
.Y(n_204)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_2),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_3),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_3),
.B(n_230),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_3),
.B(n_275),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_3),
.B(n_285),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_SL g295 ( 
.A(n_3),
.B(n_296),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_3),
.B(n_81),
.Y(n_311)
);

INVx6_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

INVx8_ASAP7_75t_L g105 ( 
.A(n_5),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g294 ( 
.A(n_5),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_6),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_6),
.B(n_113),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_6),
.B(n_118),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_6),
.B(n_148),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_6),
.B(n_221),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_6),
.B(n_251),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_6),
.B(n_269),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_6),
.B(n_292),
.Y(n_291)
);

AND2x2_ASAP7_75t_L g110 ( 
.A(n_7),
.B(n_111),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_7),
.B(n_136),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_7),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_7),
.B(n_325),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g362 ( 
.A(n_7),
.B(n_363),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_8),
.B(n_42),
.Y(n_41)
);

AND2x2_ASAP7_75t_SL g94 ( 
.A(n_8),
.B(n_95),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_8),
.B(n_140),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_8),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_8),
.B(n_184),
.Y(n_183)
);

BUFx5_ASAP7_75t_L g54 ( 
.A(n_9),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g153 ( 
.A(n_9),
.Y(n_153)
);

INVx3_ASAP7_75t_L g231 ( 
.A(n_9),
.Y(n_231)
);

INVx8_ASAP7_75t_L g76 ( 
.A(n_10),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_11),
.B(n_39),
.Y(n_38)
);

AND2x2_ASAP7_75t_L g80 ( 
.A(n_11),
.B(n_81),
.Y(n_80)
);

AND2x2_ASAP7_75t_SL g90 ( 
.A(n_11),
.B(n_91),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_11),
.B(n_134),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_11),
.B(n_172),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_11),
.B(n_227),
.Y(n_226)
);

AND2x2_ASAP7_75t_L g108 ( 
.A(n_12),
.B(n_109),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_12),
.B(n_152),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_12),
.B(n_256),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_12),
.B(n_39),
.Y(n_267)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_12),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_12),
.B(n_313),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_12),
.B(n_261),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_12),
.B(n_367),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_13),
.B(n_27),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_SL g29 ( 
.A(n_13),
.B(n_30),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_13),
.B(n_35),
.Y(n_34)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_13),
.B(n_78),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_13),
.B(n_102),
.Y(n_101)
);

AND2x2_ASAP7_75t_L g121 ( 
.A(n_13),
.B(n_122),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_13),
.B(n_190),
.Y(n_189)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_14),
.Y(n_36)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_14),
.Y(n_83)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_14),
.Y(n_177)
);

INVx1_ASAP7_75t_SL g24 ( 
.A(n_15),
.Y(n_24)
);

AND2x2_ASAP7_75t_L g51 ( 
.A(n_15),
.B(n_52),
.Y(n_51)
);

AND2x2_ASAP7_75t_L g57 ( 
.A(n_15),
.B(n_58),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_15),
.B(n_144),
.Y(n_143)
);

AND2x2_ASAP7_75t_L g203 ( 
.A(n_15),
.B(n_204),
.Y(n_203)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_207),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_206),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_166),
.Y(n_18)
);

OR2x2_ASAP7_75t_L g206 ( 
.A(n_19),
.B(n_166),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_19),
.B(n_210),
.Y(n_209)
);

OR2x2_ASAP7_75t_L g414 ( 
.A(n_19),
.B(n_210),
.Y(n_414)
);

FAx1_ASAP7_75t_SL g19 ( 
.A(n_20),
.B(n_63),
.CI(n_128),
.CON(n_19),
.SN(n_19)
);

XNOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_49),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_32),
.B1(n_47),
.B2(n_48),
.Y(n_21)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_22),
.Y(n_47)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_22),
.B(n_48),
.C(n_49),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_26),
.C(n_29),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_L g55 ( 
.A1(n_23),
.A2(n_56),
.B1(n_57),
.B2(n_61),
.Y(n_55)
);

CKINVDCx16_ASAP7_75t_R g61 ( 
.A(n_23),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g67 ( 
.A1(n_23),
.A2(n_29),
.B1(n_61),
.B2(n_68),
.Y(n_67)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_23),
.B(n_51),
.C(n_57),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g298 ( 
.A1(n_23),
.A2(n_61),
.B1(n_273),
.B2(n_274),
.Y(n_298)
);

OR2x2_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_25),
.Y(n_23)
);

OR2x2_ASAP7_75t_SL g86 ( 
.A(n_24),
.B(n_87),
.Y(n_86)
);

OR2x2_ASAP7_75t_SL g106 ( 
.A(n_24),
.B(n_107),
.Y(n_106)
);

OR2x2_ASAP7_75t_L g175 ( 
.A(n_24),
.B(n_176),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_26),
.A2(n_66),
.B1(n_67),
.B2(n_69),
.Y(n_65)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_26),
.Y(n_69)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_28),
.Y(n_40)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_28),
.Y(n_148)
);

INVx3_ASAP7_75t_L g186 ( 
.A(n_28),
.Y(n_186)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_29),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_29),
.B(n_175),
.C(n_220),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g348 ( 
.A1(n_29),
.A2(n_68),
.B1(n_174),
.B2(n_175),
.Y(n_348)
);

BUFx2_ASAP7_75t_L g134 ( 
.A(n_30),
.Y(n_134)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

BUFx8_ASAP7_75t_L g253 ( 
.A(n_31),
.Y(n_253)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_32),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g32 ( 
.A1(n_33),
.A2(n_34),
.B1(n_37),
.B2(n_46),
.Y(n_32)
);

AOI22xp5_ASAP7_75t_L g382 ( 
.A1(n_33),
.A2(n_34),
.B1(n_147),
.B2(n_383),
.Y(n_382)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_34),
.B(n_143),
.C(n_147),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_34),
.B(n_38),
.C(n_41),
.Y(n_179)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_37),
.Y(n_46)
);

XNOR2xp5_ASAP7_75t_SL g37 ( 
.A(n_38),
.B(n_41),
.Y(n_37)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_39),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx4_ASAP7_75t_SL g42 ( 
.A(n_43),
.Y(n_42)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_44),
.Y(n_79)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_45),
.Y(n_93)
);

INVx11_ASAP7_75t_L g146 ( 
.A(n_45),
.Y(n_146)
);

BUFx3_ASAP7_75t_L g222 ( 
.A(n_45),
.Y(n_222)
);

BUFx5_ASAP7_75t_L g297 ( 
.A(n_45),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_L g49 ( 
.A1(n_50),
.A2(n_51),
.B1(n_55),
.B2(n_62),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_53),
.B(n_163),
.Y(n_162)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx6_ASAP7_75t_L g114 ( 
.A(n_54),
.Y(n_114)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_55),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_56),
.A2(n_57),
.B1(n_174),
.B2(n_175),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_56),
.A2(n_57),
.B1(n_264),
.B2(n_265),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_57),
.Y(n_56)
);

MAJIxp5_ASAP7_75t_L g350 ( 
.A(n_57),
.B(n_266),
.C(n_270),
.Y(n_350)
);

BUFx6f_ASAP7_75t_L g161 ( 
.A(n_58),
.Y(n_161)
);

INVx3_ASAP7_75t_L g327 ( 
.A(n_58),
.Y(n_327)
);

INVx5_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g304 ( 
.A(n_59),
.Y(n_304)
);

INVx2_ASAP7_75t_L g315 ( 
.A(n_59),
.Y(n_315)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g272 ( 
.A(n_61),
.B(n_273),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_SL g63 ( 
.A(n_64),
.B(n_97),
.Y(n_63)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_64),
.B(n_98),
.C(n_115),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g64 ( 
.A(n_65),
.B(n_70),
.C(n_84),
.Y(n_64)
);

XOR2xp5_ASAP7_75t_L g214 ( 
.A(n_65),
.B(n_215),
.Y(n_214)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_70),
.B(n_84),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g70 ( 
.A(n_71),
.B(n_77),
.C(n_80),
.Y(n_70)
);

XNOR2xp5_ASAP7_75t_SL g130 ( 
.A(n_71),
.B(n_131),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_72),
.B(n_73),
.Y(n_71)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

BUFx12f_ASAP7_75t_L g172 ( 
.A(n_74),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_75),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_75),
.Y(n_122)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_75),
.Y(n_286)
);

INVx6_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g138 ( 
.A(n_76),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_L g131 ( 
.A(n_77),
.B(n_80),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_77),
.A2(n_183),
.B1(n_187),
.B2(n_188),
.Y(n_182)
);

INVx1_ASAP7_75t_SL g188 ( 
.A(n_77),
.Y(n_188)
);

INVx5_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_83),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_85),
.A2(n_86),
.B1(n_89),
.B2(n_96),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_86),
.B(n_126),
.C(n_127),
.Y(n_125)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx5_ASAP7_75t_L g368 ( 
.A(n_88),
.Y(n_368)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_89),
.Y(n_96)
);

XNOR2xp5_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_94),
.Y(n_89)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_90),
.Y(n_126)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_94),
.Y(n_127)
);

XNOR2xp5_ASAP7_75t_L g97 ( 
.A(n_98),
.B(n_115),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_110),
.C(n_112),
.Y(n_98)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

XNOR2xp5_ASAP7_75t_L g164 ( 
.A(n_100),
.B(n_165),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_101),
.B(n_106),
.C(n_108),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_101),
.A2(n_108),
.B1(n_236),
.B2(n_237),
.Y(n_235)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_101),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_101),
.A2(n_237),
.B1(n_283),
.B2(n_284),
.Y(n_282)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g141 ( 
.A(n_105),
.Y(n_141)
);

INVx4_ASAP7_75t_L g227 ( 
.A(n_105),
.Y(n_227)
);

INVx2_ASAP7_75t_L g308 ( 
.A(n_105),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_106),
.A2(n_233),
.B1(n_234),
.B2(n_235),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_106),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_108),
.Y(n_236)
);

XOR2xp5_ASAP7_75t_L g165 ( 
.A(n_110),
.B(n_112),
.Y(n_165)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

XNOR2xp5_ASAP7_75t_L g115 ( 
.A(n_116),
.B(n_125),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_117),
.A2(n_121),
.B1(n_123),
.B2(n_124),
.Y(n_116)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_117),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_121),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_121),
.B(n_123),
.C(n_198),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_121),
.A2(n_124),
.B1(n_202),
.B2(n_203),
.Y(n_201)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_125),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_129),
.B(n_149),
.C(n_164),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_SL g212 ( 
.A(n_129),
.B(n_213),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_132),
.C(n_142),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_L g403 ( 
.A(n_130),
.B(n_142),
.Y(n_403)
);

XNOR2xp5_ASAP7_75t_L g402 ( 
.A(n_132),
.B(n_403),
.Y(n_402)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_133),
.B(n_135),
.C(n_139),
.Y(n_132)
);

FAx1_ASAP7_75t_SL g218 ( 
.A(n_133),
.B(n_135),
.CI(n_139),
.CON(n_218),
.SN(n_218)
);

INVx5_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

INVx8_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g380 ( 
.A1(n_143),
.A2(n_381),
.B1(n_382),
.B2(n_384),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_143),
.Y(n_381)
);

INVx6_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

INVx6_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g258 ( 
.A(n_146),
.Y(n_258)
);

INVx5_ASAP7_75t_L g281 ( 
.A(n_146),
.Y(n_281)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_147),
.Y(n_383)
);

XNOR2xp5_ASAP7_75t_L g213 ( 
.A(n_149),
.B(n_164),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_158),
.C(n_162),
.Y(n_149)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_150),
.B(n_239),
.Y(n_238)
);

OAI21xp5_ASAP7_75t_L g379 ( 
.A1(n_150),
.A2(n_151),
.B(n_154),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_154),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

INVx4_ASAP7_75t_L g191 ( 
.A(n_153),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_SL g154 ( 
.A(n_155),
.B(n_157),
.Y(n_154)
);

INVx8_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_157),
.B(n_304),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_158),
.B(n_162),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_160),
.Y(n_158)
);

INVx3_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_163),
.B(n_260),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_163),
.B(n_278),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_163),
.B(n_318),
.Y(n_317)
);

XNOR2xp5_ASAP7_75t_L g166 ( 
.A(n_167),
.B(n_168),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_193),
.Y(n_168)
);

XOR2xp5_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_178),
.Y(n_169)
);

XOR2xp5_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_173),
.Y(n_170)
);

CKINVDCx16_ASAP7_75t_R g174 ( 
.A(n_175),
.Y(n_174)
);

BUFx5_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g262 ( 
.A(n_177),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_180),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_181),
.A2(n_182),
.B1(n_189),
.B2(n_192),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_183),
.Y(n_187)
);

INVx6_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

INVx8_ASAP7_75t_L g275 ( 
.A(n_185),
.Y(n_275)
);

INVx4_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

BUFx6f_ASAP7_75t_L g365 ( 
.A(n_186),
.Y(n_365)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_189),
.Y(n_192)
);

INVx6_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_194),
.A2(n_195),
.B1(n_196),
.B2(n_205),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_196),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_SL g196 ( 
.A(n_197),
.B(n_199),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g199 ( 
.A(n_200),
.B(n_201),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_203),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_L g207 ( 
.A1(n_208),
.A2(n_240),
.B(n_414),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_211),
.B(n_214),
.C(n_216),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g408 ( 
.A1(n_211),
.A2(n_212),
.B1(n_214),
.B2(n_409),
.Y(n_408)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_214),
.Y(n_409)
);

XOR2xp5_ASAP7_75t_L g407 ( 
.A(n_216),
.B(n_408),
.Y(n_407)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_217),
.B(n_232),
.C(n_238),
.Y(n_216)
);

XOR2xp5_ASAP7_75t_L g398 ( 
.A(n_217),
.B(n_399),
.Y(n_398)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_219),
.C(n_223),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g389 ( 
.A(n_218),
.B(n_390),
.Y(n_389)
);

BUFx24_ASAP7_75t_SL g415 ( 
.A(n_218),
.Y(n_415)
);

AOI22xp5_ASAP7_75t_L g390 ( 
.A1(n_219),
.A2(n_223),
.B1(n_224),
.B2(n_391),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_219),
.Y(n_391)
);

XNOR2xp5_ASAP7_75t_SL g347 ( 
.A(n_220),
.B(n_348),
.Y(n_347)
);

INVx3_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_225),
.B(n_228),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g351 ( 
.A1(n_225),
.A2(n_226),
.B1(n_228),
.B2(n_229),
.Y(n_351)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

INVx3_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g399 ( 
.A(n_232),
.B(n_238),
.Y(n_399)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_237),
.B(n_283),
.Y(n_358)
);

AOI21xp5_ASAP7_75t_L g240 ( 
.A1(n_241),
.A2(n_394),
.B(n_410),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

AOI21xp5_ASAP7_75t_L g242 ( 
.A1(n_243),
.A2(n_372),
.B(n_393),
.Y(n_242)
);

OAI21xp5_ASAP7_75t_SL g243 ( 
.A1(n_244),
.A2(n_342),
.B(n_371),
.Y(n_243)
);

AOI21xp5_ASAP7_75t_L g244 ( 
.A1(n_245),
.A2(n_299),
.B(n_341),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_SL g245 ( 
.A(n_246),
.B(n_287),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g341 ( 
.A(n_246),
.B(n_287),
.Y(n_341)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_247),
.B(n_271),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_248),
.B(n_263),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g343 ( 
.A(n_248),
.B(n_263),
.C(n_271),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_249),
.B(n_254),
.C(n_259),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_249),
.A2(n_250),
.B1(n_254),
.B2(n_255),
.Y(n_289)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

INVx8_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

INVx3_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_SL g288 ( 
.A(n_259),
.B(n_289),
.Y(n_288)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

INVx3_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

INVx3_ASAP7_75t_L g269 ( 
.A(n_262),
.Y(n_269)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_L g265 ( 
.A1(n_266),
.A2(n_267),
.B1(n_268),
.B2(n_270),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_268),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_SL g271 ( 
.A(n_272),
.B(n_276),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g354 ( 
.A(n_272),
.B(n_355),
.C(n_356),
.Y(n_354)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_277),
.B(n_282),
.Y(n_276)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_277),
.Y(n_355)
);

INVx1_ASAP7_75t_SL g278 ( 
.A(n_279),
.Y(n_278)
);

BUFx3_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

INVx5_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_282),
.Y(n_356)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_288),
.B(n_290),
.C(n_298),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_L g337 ( 
.A(n_288),
.B(n_338),
.Y(n_337)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_290),
.Y(n_333)
);

AOI22xp5_ASAP7_75t_L g338 ( 
.A1(n_290),
.A2(n_298),
.B1(n_333),
.B2(n_339),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_SL g290 ( 
.A(n_291),
.B(n_295),
.Y(n_290)
);

INVxp67_ASAP7_75t_L g331 ( 
.A(n_291),
.Y(n_331)
);

INVx2_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

INVx3_ASAP7_75t_L g318 ( 
.A(n_294),
.Y(n_318)
);

INVxp67_ASAP7_75t_L g332 ( 
.A(n_295),
.Y(n_332)
);

INVx5_ASAP7_75t_L g296 ( 
.A(n_297),
.Y(n_296)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_298),
.Y(n_339)
);

OAI21xp5_ASAP7_75t_L g299 ( 
.A1(n_300),
.A2(n_335),
.B(n_340),
.Y(n_299)
);

AOI21xp5_ASAP7_75t_L g300 ( 
.A1(n_301),
.A2(n_320),
.B(n_334),
.Y(n_300)
);

OAI21xp5_ASAP7_75t_L g301 ( 
.A1(n_302),
.A2(n_309),
.B(n_319),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_303),
.B(n_305),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_306),
.B(n_307),
.Y(n_305)
);

INVx4_ASAP7_75t_L g307 ( 
.A(n_308),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_SL g309 ( 
.A(n_310),
.B(n_317),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_310),
.B(n_317),
.Y(n_319)
);

AOI21xp5_ASAP7_75t_L g310 ( 
.A1(n_311),
.A2(n_312),
.B(n_316),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_311),
.B(n_312),
.Y(n_316)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_314),
.Y(n_313)
);

INVx4_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_L g321 ( 
.A1(n_316),
.A2(n_322),
.B1(n_328),
.B2(n_329),
.Y(n_321)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_316),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_SL g320 ( 
.A(n_321),
.B(n_330),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_321),
.B(n_330),
.Y(n_334)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_322),
.Y(n_329)
);

XNOR2xp5_ASAP7_75t_SL g322 ( 
.A(n_323),
.B(n_324),
.Y(n_322)
);

OAI21xp5_ASAP7_75t_SL g336 ( 
.A1(n_323),
.A2(n_324),
.B(n_328),
.Y(n_336)
);

INVx2_ASAP7_75t_L g325 ( 
.A(n_326),
.Y(n_325)
);

HB1xp67_ASAP7_75t_L g326 ( 
.A(n_327),
.Y(n_326)
);

OAI21xp5_ASAP7_75t_SL g330 ( 
.A1(n_331),
.A2(n_332),
.B(n_333),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_336),
.B(n_337),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_336),
.B(n_337),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_L g342 ( 
.A(n_343),
.B(n_344),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_343),
.B(n_344),
.Y(n_371)
);

OAI22xp5_ASAP7_75t_L g344 ( 
.A1(n_345),
.A2(n_346),
.B1(n_352),
.B2(n_353),
.Y(n_344)
);

MAJIxp5_ASAP7_75t_L g373 ( 
.A(n_345),
.B(n_354),
.C(n_357),
.Y(n_373)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_346),
.Y(n_345)
);

XOR2xp5_ASAP7_75t_L g346 ( 
.A(n_347),
.B(n_349),
.Y(n_346)
);

MAJIxp5_ASAP7_75t_L g388 ( 
.A(n_347),
.B(n_350),
.C(n_351),
.Y(n_388)
);

XOR2xp5_ASAP7_75t_L g349 ( 
.A(n_350),
.B(n_351),
.Y(n_349)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_353),
.Y(n_352)
);

XOR2xp5_ASAP7_75t_L g353 ( 
.A(n_354),
.B(n_357),
.Y(n_353)
);

OAI22xp5_ASAP7_75t_L g357 ( 
.A1(n_358),
.A2(n_359),
.B1(n_360),
.B2(n_370),
.Y(n_357)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_358),
.Y(n_370)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_360),
.Y(n_359)
);

AOI22xp5_ASAP7_75t_L g360 ( 
.A1(n_361),
.A2(n_362),
.B1(n_366),
.B2(n_369),
.Y(n_360)
);

MAJIxp5_ASAP7_75t_L g377 ( 
.A(n_361),
.B(n_369),
.C(n_370),
.Y(n_377)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_362),
.Y(n_361)
);

INVx5_ASAP7_75t_L g363 ( 
.A(n_364),
.Y(n_363)
);

INVx5_ASAP7_75t_L g364 ( 
.A(n_365),
.Y(n_364)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_366),
.Y(n_369)
);

INVx4_ASAP7_75t_SL g367 ( 
.A(n_368),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_373),
.B(n_374),
.Y(n_372)
);

NOR2xp33_ASAP7_75t_L g393 ( 
.A(n_373),
.B(n_374),
.Y(n_393)
);

AOI22xp5_ASAP7_75t_L g374 ( 
.A1(n_375),
.A2(n_376),
.B1(n_387),
.B2(n_392),
.Y(n_374)
);

MAJIxp5_ASAP7_75t_L g404 ( 
.A(n_375),
.B(n_388),
.C(n_389),
.Y(n_404)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_376),
.Y(n_375)
);

XNOR2xp5_ASAP7_75t_SL g376 ( 
.A(n_377),
.B(n_378),
.Y(n_376)
);

MAJIxp5_ASAP7_75t_L g401 ( 
.A(n_377),
.B(n_380),
.C(n_385),
.Y(n_401)
);

AOI22xp5_ASAP7_75t_L g378 ( 
.A1(n_379),
.A2(n_380),
.B1(n_385),
.B2(n_386),
.Y(n_378)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_379),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_380),
.Y(n_386)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_382),
.Y(n_384)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_387),
.Y(n_392)
);

XNOR2xp5_ASAP7_75t_SL g387 ( 
.A(n_388),
.B(n_389),
.Y(n_387)
);

INVxp67_ASAP7_75t_L g394 ( 
.A(n_395),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_396),
.B(n_405),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_SL g396 ( 
.A(n_397),
.B(n_404),
.Y(n_396)
);

NOR2xp33_ASAP7_75t_L g412 ( 
.A(n_397),
.B(n_404),
.Y(n_412)
);

XOR2xp5_ASAP7_75t_L g397 ( 
.A(n_398),
.B(n_400),
.Y(n_397)
);

MAJIxp5_ASAP7_75t_L g406 ( 
.A(n_398),
.B(n_401),
.C(n_402),
.Y(n_406)
);

XNOR2xp5_ASAP7_75t_L g400 ( 
.A(n_401),
.B(n_402),
.Y(n_400)
);

AOI21xp5_ASAP7_75t_L g411 ( 
.A1(n_405),
.A2(n_412),
.B(n_413),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_406),
.B(n_407),
.Y(n_405)
);

NOR2xp33_ASAP7_75t_L g413 ( 
.A(n_406),
.B(n_407),
.Y(n_413)
);

INVxp67_ASAP7_75t_L g410 ( 
.A(n_411),
.Y(n_410)
);


endmodule