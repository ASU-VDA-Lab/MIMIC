module fake_jpeg_23407_n_345 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_345);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_345;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx13_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

INVx6_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

BUFx4f_ASAP7_75t_SL g18 ( 
.A(n_10),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_11),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_5),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_14),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_2),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_7),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

INVx5_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_1),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_4),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_2),
.Y(n_34)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_5),
.Y(n_35)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_21),
.Y(n_36)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_36),
.A2(n_16),
.B1(n_31),
.B2(n_35),
.Y(n_54)
);

CKINVDCx5p33_ASAP7_75t_R g37 ( 
.A(n_18),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_37),
.B(n_46),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_16),
.B(n_0),
.Y(n_38)
);

A2O1A1Ixp33_ASAP7_75t_L g64 ( 
.A1(n_38),
.A2(n_41),
.B(n_27),
.C(n_24),
.Y(n_64)
);

BUFx5_ASAP7_75t_L g39 ( 
.A(n_18),
.Y(n_39)
);

INVxp67_ASAP7_75t_SL g53 ( 
.A(n_39),
.Y(n_53)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_18),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_40),
.B(n_43),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_19),
.B(n_15),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_18),
.Y(n_42)
);

BUFx10_ASAP7_75t_L g76 ( 
.A(n_42),
.Y(n_76)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_18),
.Y(n_43)
);

INVx11_ASAP7_75t_L g44 ( 
.A(n_16),
.Y(n_44)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_44),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g45 ( 
.A(n_17),
.B(n_0),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_45),
.B(n_47),
.Y(n_58)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_18),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g47 ( 
.A(n_17),
.B(n_0),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_23),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_48),
.B(n_34),
.Y(n_73)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_33),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_49),
.B(n_35),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_33),
.Y(n_50)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_50),
.Y(n_61)
);

INVx11_ASAP7_75t_L g51 ( 
.A(n_16),
.Y(n_51)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_51),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_54),
.A2(n_59),
.B1(n_65),
.B2(n_36),
.Y(n_110)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

CKINVDCx14_ASAP7_75t_R g106 ( 
.A(n_55),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_36),
.A2(n_31),
.B1(n_35),
.B2(n_17),
.Y(n_59)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_39),
.Y(n_60)
);

INVx11_ASAP7_75t_L g117 ( 
.A(n_60),
.Y(n_117)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_38),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_63),
.B(n_64),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_36),
.A2(n_31),
.B1(n_35),
.B2(n_17),
.Y(n_65)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_39),
.Y(n_66)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_66),
.Y(n_91)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_50),
.Y(n_67)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_67),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_41),
.B(n_20),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_68),
.B(n_73),
.Y(n_96)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_69),
.Y(n_100)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_44),
.Y(n_70)
);

INVx8_ASAP7_75t_L g88 ( 
.A(n_70),
.Y(n_88)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_50),
.Y(n_71)
);

HB1xp67_ASAP7_75t_L g94 ( 
.A(n_71),
.Y(n_94)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_50),
.Y(n_72)
);

HB1xp67_ASAP7_75t_L g101 ( 
.A(n_72),
.Y(n_101)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_50),
.Y(n_74)
);

INVx1_ASAP7_75t_SL g114 ( 
.A(n_74),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_48),
.B(n_19),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_75),
.B(n_79),
.Y(n_98)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_49),
.Y(n_77)
);

INVx1_ASAP7_75t_SL g115 ( 
.A(n_77),
.Y(n_115)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_49),
.Y(n_78)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_78),
.Y(n_102)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_44),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_45),
.A2(n_33),
.B1(n_34),
.B2(n_32),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_80),
.A2(n_20),
.B1(n_22),
.B2(n_25),
.Y(n_120)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_37),
.Y(n_81)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_81),
.Y(n_104)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_53),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_82),
.B(n_83),
.Y(n_135)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_55),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_57),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_SL g128 ( 
.A(n_84),
.B(n_103),
.Y(n_128)
);

O2A1O1Ixp33_ASAP7_75t_L g85 ( 
.A1(n_80),
.A2(n_47),
.B(n_45),
.C(n_38),
.Y(n_85)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_85),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_55),
.Y(n_86)
);

INVxp67_ASAP7_75t_SL g149 ( 
.A(n_86),
.Y(n_149)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_61),
.Y(n_87)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_87),
.Y(n_140)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_61),
.Y(n_89)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_89),
.Y(n_151)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_77),
.Y(n_90)
);

HB1xp67_ASAP7_75t_L g143 ( 
.A(n_90),
.Y(n_143)
);

BUFx12f_ASAP7_75t_L g92 ( 
.A(n_60),
.Y(n_92)
);

INVx5_ASAP7_75t_L g141 ( 
.A(n_92),
.Y(n_141)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_78),
.Y(n_93)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_93),
.Y(n_147)
);

AOI32xp33_ASAP7_75t_L g95 ( 
.A1(n_52),
.A2(n_51),
.A3(n_44),
.B1(n_33),
.B2(n_37),
.Y(n_95)
);

AOI32xp33_ASAP7_75t_L g142 ( 
.A1(n_95),
.A2(n_90),
.A3(n_118),
.B1(n_117),
.B2(n_101),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_67),
.Y(n_97)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_97),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_58),
.B(n_48),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_62),
.B(n_47),
.Y(n_105)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_105),
.Y(n_126)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_62),
.Y(n_107)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_107),
.Y(n_148)
);

A2O1A1Ixp33_ASAP7_75t_L g109 ( 
.A1(n_64),
.A2(n_51),
.B(n_42),
.C(n_22),
.Y(n_109)
);

XNOR2xp5_ASAP7_75t_SL g132 ( 
.A(n_109),
.B(n_120),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_SL g138 ( 
.A1(n_110),
.A2(n_113),
.B1(n_118),
.B2(n_56),
.Y(n_138)
);

INVx2_ASAP7_75t_SL g111 ( 
.A(n_70),
.Y(n_111)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_111),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_79),
.B(n_19),
.Y(n_112)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_112),
.Y(n_145)
);

INVx2_ASAP7_75t_SL g113 ( 
.A(n_71),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_76),
.B(n_20),
.Y(n_116)
);

AND2x2_ASAP7_75t_L g125 ( 
.A(n_116),
.B(n_25),
.Y(n_125)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_72),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_74),
.Y(n_119)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_119),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_98),
.B(n_37),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_123),
.B(n_127),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_125),
.B(n_129),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_85),
.B(n_21),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_108),
.B(n_21),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_120),
.B(n_21),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_130),
.B(n_131),
.Y(n_177)
);

OAI32xp33_ASAP7_75t_L g131 ( 
.A1(n_109),
.A2(n_40),
.A3(n_43),
.B1(n_81),
.B2(n_46),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_96),
.A2(n_51),
.B1(n_66),
.B2(n_56),
.Y(n_134)
);

INVxp67_ASAP7_75t_L g160 ( 
.A(n_134),
.Y(n_160)
);

O2A1O1Ixp33_ASAP7_75t_SL g136 ( 
.A1(n_94),
.A2(n_43),
.B(n_40),
.C(n_42),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_136),
.A2(n_142),
.B1(n_150),
.B2(n_111),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_L g137 ( 
.A1(n_100),
.A2(n_23),
.B(n_26),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_L g152 ( 
.A1(n_137),
.A2(n_32),
.B(n_28),
.Y(n_152)
);

INVxp67_ASAP7_75t_L g161 ( 
.A(n_138),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_L g139 ( 
.A1(n_88),
.A2(n_22),
.B1(n_25),
.B2(n_24),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_139),
.A2(n_88),
.B1(n_107),
.B2(n_87),
.Y(n_154)
);

AND2x2_ASAP7_75t_L g144 ( 
.A(n_106),
.B(n_1),
.Y(n_144)
);

AND2x2_ASAP7_75t_L g170 ( 
.A(n_144),
.B(n_15),
.Y(n_170)
);

OAI32xp33_ASAP7_75t_L g146 ( 
.A1(n_104),
.A2(n_46),
.A3(n_42),
.B1(n_27),
.B2(n_24),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_146),
.B(n_76),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_99),
.A2(n_23),
.B1(n_26),
.B2(n_34),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_L g187 ( 
.A1(n_152),
.A2(n_169),
.B(n_137),
.Y(n_187)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_143),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_153),
.B(n_156),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_154),
.A2(n_158),
.B1(n_124),
.B2(n_133),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_L g204 ( 
.A1(n_155),
.A2(n_157),
.B1(n_159),
.B2(n_181),
.Y(n_204)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_135),
.Y(n_156)
);

AOI22xp33_ASAP7_75t_SL g157 ( 
.A1(n_122),
.A2(n_82),
.B1(n_113),
.B2(n_89),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_121),
.A2(n_93),
.B1(n_102),
.B2(n_91),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_121),
.A2(n_115),
.B1(n_114),
.B2(n_117),
.Y(n_159)
);

HB1xp67_ASAP7_75t_L g162 ( 
.A(n_149),
.Y(n_162)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_162),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_SL g164 ( 
.A(n_128),
.B(n_83),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_164),
.B(n_167),
.Y(n_211)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_148),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_165),
.B(n_175),
.Y(n_203)
);

BUFx24_ASAP7_75t_L g166 ( 
.A(n_141),
.Y(n_166)
);

INVx1_ASAP7_75t_SL g189 ( 
.A(n_166),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_145),
.B(n_115),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_L g168 ( 
.A(n_132),
.B(n_92),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_L g192 ( 
.A(n_168),
.B(n_183),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_L g169 ( 
.A1(n_129),
.A2(n_28),
.B(n_26),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_170),
.B(n_172),
.Y(n_212)
);

OAI32xp33_ASAP7_75t_L g171 ( 
.A1(n_127),
.A2(n_92),
.A3(n_42),
.B1(n_24),
.B2(n_27),
.Y(n_171)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_171),
.B(n_182),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_SL g172 ( 
.A(n_145),
.B(n_32),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_133),
.B(n_114),
.Y(n_173)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_173),
.Y(n_194)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_148),
.Y(n_175)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_122),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_176),
.B(n_124),
.Y(n_205)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_136),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_178),
.B(n_184),
.Y(n_197)
);

AND2x2_ASAP7_75t_L g179 ( 
.A(n_123),
.B(n_1),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_SL g195 ( 
.A1(n_179),
.A2(n_180),
.B(n_144),
.Y(n_195)
);

OA21x2_ASAP7_75t_L g180 ( 
.A1(n_131),
.A2(n_28),
.B(n_76),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_126),
.B(n_76),
.C(n_86),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_132),
.B(n_27),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_136),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_150),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_185),
.B(n_144),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_126),
.B(n_119),
.C(n_97),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_186),
.B(n_30),
.Y(n_217)
);

FAx1_ASAP7_75t_SL g232 ( 
.A(n_187),
.B(n_180),
.CI(n_171),
.CON(n_232),
.SN(n_232)
);

AOI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_160),
.A2(n_130),
.B1(n_134),
.B2(n_146),
.Y(n_188)
);

OAI21xp33_ASAP7_75t_SL g236 ( 
.A1(n_188),
.A2(n_195),
.B(n_200),
.Y(n_236)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_166),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_193),
.B(n_198),
.Y(n_222)
);

OR2x6_ASAP7_75t_L g196 ( 
.A(n_170),
.B(n_125),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_SL g228 ( 
.A1(n_196),
.A2(n_161),
.B(n_179),
.Y(n_228)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_158),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_L g199 ( 
.A(n_168),
.B(n_125),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_199),
.B(n_207),
.Y(n_224)
);

OAI21xp33_ASAP7_75t_L g225 ( 
.A1(n_201),
.A2(n_196),
.B(n_211),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_152),
.B(n_151),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_202),
.B(n_206),
.Y(n_229)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_205),
.Y(n_234)
);

INVxp67_ASAP7_75t_L g206 ( 
.A(n_166),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_183),
.B(n_141),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_160),
.A2(n_140),
.B1(n_147),
.B2(n_30),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_L g235 ( 
.A1(n_208),
.A2(n_210),
.B1(n_176),
.B2(n_175),
.Y(n_235)
);

CKINVDCx14_ASAP7_75t_R g209 ( 
.A(n_186),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_209),
.B(n_213),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_177),
.A2(n_147),
.B1(n_30),
.B2(n_29),
.Y(n_210)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_159),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_155),
.A2(n_30),
.B1(n_29),
.B2(n_4),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_214),
.A2(n_219),
.B1(n_154),
.B2(n_196),
.Y(n_226)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_182),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_215),
.B(n_15),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_217),
.B(n_216),
.C(n_208),
.Y(n_230)
);

OAI21xp5_ASAP7_75t_L g218 ( 
.A1(n_174),
.A2(n_29),
.B(n_3),
.Y(n_218)
);

OAI21xp5_ASAP7_75t_L g233 ( 
.A1(n_218),
.A2(n_197),
.B(n_212),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_174),
.A2(n_29),
.B1(n_3),
.B2(n_4),
.Y(n_219)
);

OAI32xp33_ASAP7_75t_L g220 ( 
.A1(n_180),
.A2(n_2),
.A3(n_3),
.B1(n_5),
.B2(n_6),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_220),
.B(n_169),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_SL g221 ( 
.A(n_196),
.B(n_163),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_221),
.B(n_225),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_223),
.B(n_226),
.Y(n_258)
);

NAND3xp33_ASAP7_75t_L g227 ( 
.A(n_196),
.B(n_170),
.C(n_179),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_227),
.Y(n_262)
);

AOI21xp5_ASAP7_75t_L g269 ( 
.A1(n_228),
.A2(n_237),
.B(n_243),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_230),
.B(n_239),
.C(n_217),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_SL g249 ( 
.A(n_232),
.B(n_226),
.Y(n_249)
);

AOI21xp5_ASAP7_75t_SL g256 ( 
.A1(n_233),
.A2(n_214),
.B(n_204),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_235),
.A2(n_189),
.B1(n_194),
.B2(n_200),
.Y(n_259)
);

XOR2x2_ASAP7_75t_L g237 ( 
.A(n_192),
.B(n_161),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_220),
.A2(n_165),
.B1(n_10),
.B2(n_12),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_238),
.A2(n_246),
.B1(n_206),
.B2(n_188),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_192),
.B(n_2),
.C(n_3),
.Y(n_239)
);

INVxp67_ASAP7_75t_L g240 ( 
.A(n_203),
.Y(n_240)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_240),
.Y(n_253)
);

INVxp67_ASAP7_75t_L g264 ( 
.A(n_241),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_191),
.B(n_6),
.Y(n_242)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_242),
.Y(n_266)
);

OAI21xp5_ASAP7_75t_L g243 ( 
.A1(n_187),
.A2(n_6),
.B(n_7),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_189),
.B(n_6),
.Y(n_244)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_244),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_218),
.B(n_7),
.Y(n_245)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_245),
.Y(n_260)
);

AOI21xp5_ASAP7_75t_L g246 ( 
.A1(n_195),
.A2(n_7),
.B(n_8),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_190),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_247),
.Y(n_263)
);

HB1xp67_ASAP7_75t_L g248 ( 
.A(n_193),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_248),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_SL g277 ( 
.A(n_249),
.B(n_231),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_250),
.A2(n_235),
.B1(n_229),
.B2(n_228),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_251),
.B(n_252),
.C(n_230),
.Y(n_276)
);

XOR2xp5_ASAP7_75t_L g252 ( 
.A(n_224),
.B(n_207),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_221),
.B(n_219),
.Y(n_255)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_255),
.Y(n_281)
);

OAI21xp5_ASAP7_75t_L g282 ( 
.A1(n_256),
.A2(n_246),
.B(n_223),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_224),
.B(n_199),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g290 ( 
.A(n_257),
.B(n_265),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_259),
.A2(n_261),
.B1(n_238),
.B2(n_222),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_236),
.A2(n_216),
.B1(n_210),
.B2(n_9),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g265 ( 
.A(n_237),
.B(n_13),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_245),
.B(n_8),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_267),
.Y(n_274)
);

BUFx6f_ASAP7_75t_L g271 ( 
.A(n_248),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_271),
.B(n_268),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_263),
.B(n_244),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_SL g297 ( 
.A(n_272),
.B(n_287),
.Y(n_297)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_273),
.Y(n_301)
);

AND2x2_ASAP7_75t_L g275 ( 
.A(n_262),
.B(n_237),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_275),
.B(n_254),
.Y(n_291)
);

XOR2xp5_ASAP7_75t_L g294 ( 
.A(n_276),
.B(n_277),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_SL g278 ( 
.A(n_258),
.B(n_231),
.Y(n_278)
);

XOR2xp5_ASAP7_75t_L g296 ( 
.A(n_278),
.B(n_282),
.Y(n_296)
);

INVx2_ASAP7_75t_L g279 ( 
.A(n_271),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_279),
.B(n_285),
.Y(n_295)
);

HB1xp67_ASAP7_75t_L g280 ( 
.A(n_253),
.Y(n_280)
);

INVx13_ASAP7_75t_L g303 ( 
.A(n_280),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_SL g283 ( 
.A(n_261),
.B(n_229),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_283),
.B(n_289),
.C(n_269),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_SL g299 ( 
.A1(n_284),
.A2(n_260),
.B1(n_256),
.B2(n_267),
.Y(n_299)
);

INVxp67_ASAP7_75t_SL g286 ( 
.A(n_259),
.Y(n_286)
);

INVxp33_ASAP7_75t_L g304 ( 
.A(n_286),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_264),
.B(n_234),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_250),
.A2(n_222),
.B1(n_234),
.B2(n_241),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_L g302 ( 
.A1(n_288),
.A2(n_264),
.B1(n_232),
.B2(n_247),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_SL g289 ( 
.A(n_249),
.B(n_233),
.Y(n_289)
);

AOI21xp5_ASAP7_75t_L g315 ( 
.A1(n_291),
.A2(n_298),
.B(n_300),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_286),
.A2(n_255),
.B1(n_260),
.B2(n_269),
.Y(n_292)
);

XOR2xp5_ASAP7_75t_L g313 ( 
.A(n_292),
.B(n_293),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_SL g298 ( 
.A(n_281),
.B(n_270),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_L g316 ( 
.A1(n_299),
.A2(n_302),
.B1(n_232),
.B2(n_290),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_274),
.B(n_266),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_282),
.B(n_242),
.Y(n_305)
);

OAI21xp5_ASAP7_75t_SL g310 ( 
.A1(n_305),
.A2(n_239),
.B(n_283),
.Y(n_310)
);

OAI21xp5_ASAP7_75t_L g306 ( 
.A1(n_291),
.A2(n_276),
.B(n_251),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_306),
.B(n_307),
.C(n_308),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_294),
.B(n_252),
.C(n_278),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_L g308 ( 
.A(n_296),
.B(n_277),
.Y(n_308)
);

INVxp33_ASAP7_75t_SL g309 ( 
.A(n_304),
.Y(n_309)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_309),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_310),
.B(n_314),
.Y(n_319)
);

OAI221xp5_ASAP7_75t_L g311 ( 
.A1(n_300),
.A2(n_243),
.B1(n_275),
.B2(n_289),
.C(n_265),
.Y(n_311)
);

AOI31xp33_ASAP7_75t_L g320 ( 
.A1(n_311),
.A2(n_302),
.A3(n_309),
.B(n_292),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_294),
.B(n_290),
.C(n_257),
.Y(n_312)
);

OAI21xp5_ASAP7_75t_SL g325 ( 
.A1(n_312),
.A2(n_318),
.B(n_297),
.Y(n_325)
);

INVxp67_ASAP7_75t_SL g314 ( 
.A(n_303),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_316),
.B(n_317),
.Y(n_324)
);

OAI21xp5_ASAP7_75t_L g317 ( 
.A1(n_301),
.A2(n_13),
.B(n_14),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_301),
.B(n_296),
.C(n_293),
.Y(n_318)
);

AOI21xp5_ASAP7_75t_L g334 ( 
.A1(n_320),
.A2(n_323),
.B(n_325),
.Y(n_334)
);

AOI22xp5_ASAP7_75t_L g322 ( 
.A1(n_318),
.A2(n_295),
.B1(n_299),
.B2(n_298),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_322),
.B(n_327),
.Y(n_328)
);

AND2x2_ASAP7_75t_L g323 ( 
.A(n_313),
.B(n_303),
.Y(n_323)
);

HB1xp67_ASAP7_75t_L g327 ( 
.A(n_315),
.Y(n_327)
);

NOR2xp67_ASAP7_75t_SL g329 ( 
.A(n_323),
.B(n_313),
.Y(n_329)
);

AOI21xp5_ASAP7_75t_L g335 ( 
.A1(n_329),
.A2(n_330),
.B(n_331),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_324),
.B(n_308),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_324),
.B(n_307),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_321),
.B(n_312),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_332),
.B(n_333),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_326),
.B(n_8),
.C(n_9),
.Y(n_333)
);

INVxp67_ASAP7_75t_L g336 ( 
.A(n_328),
.Y(n_336)
);

CKINVDCx20_ASAP7_75t_R g340 ( 
.A(n_336),
.Y(n_340)
);

XNOR2xp5_ASAP7_75t_L g338 ( 
.A(n_333),
.B(n_319),
.Y(n_338)
);

INVxp67_ASAP7_75t_L g339 ( 
.A(n_338),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_L g341 ( 
.A(n_340),
.B(n_335),
.Y(n_341)
);

AOI22xp33_ASAP7_75t_L g342 ( 
.A1(n_341),
.A2(n_334),
.B1(n_337),
.B2(n_339),
.Y(n_342)
);

OAI21xp5_ASAP7_75t_SL g343 ( 
.A1(n_342),
.A2(n_14),
.B(n_8),
.Y(n_343)
);

XOR2xp5_ASAP7_75t_L g344 ( 
.A(n_343),
.B(n_9),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_344),
.B(n_9),
.Y(n_345)
);


endmodule