module fake_jpeg_2786_n_541 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_541);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_541;

wire n_529;
wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_393;
wire n_349;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_341;
wire n_151;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx3_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_2),
.B(n_4),
.Y(n_20)
);

INVx11_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_15),
.Y(n_24)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_14),
.Y(n_26)
);

BUFx10_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_3),
.Y(n_30)
);

BUFx10_ASAP7_75t_L g31 ( 
.A(n_15),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_5),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_5),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_6),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_0),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_10),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_8),
.Y(n_38)
);

CKINVDCx16_ASAP7_75t_R g39 ( 
.A(n_0),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_1),
.Y(n_40)
);

INVx11_ASAP7_75t_L g41 ( 
.A(n_5),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_3),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_2),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_3),
.Y(n_44)
);

CKINVDCx12_ASAP7_75t_R g45 ( 
.A(n_2),
.Y(n_45)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_4),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_5),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_7),
.Y(n_48)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_24),
.Y(n_49)
);

INVx2_ASAP7_75t_SL g145 ( 
.A(n_49),
.Y(n_145)
);

INVx11_ASAP7_75t_L g50 ( 
.A(n_33),
.Y(n_50)
);

INVx11_ASAP7_75t_L g135 ( 
.A(n_50),
.Y(n_135)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_28),
.Y(n_51)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_51),
.Y(n_109)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_24),
.Y(n_52)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_52),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_20),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_53),
.B(n_57),
.Y(n_106)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_17),
.Y(n_54)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_54),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_20),
.B(n_0),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_55),
.B(n_59),
.Y(n_102)
);

INVx11_ASAP7_75t_L g56 ( 
.A(n_33),
.Y(n_56)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_56),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_44),
.Y(n_57)
);

INVx3_ASAP7_75t_SL g58 ( 
.A(n_24),
.Y(n_58)
);

HB1xp67_ASAP7_75t_L g143 ( 
.A(n_58),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_17),
.B(n_9),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_18),
.Y(n_60)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_60),
.Y(n_146)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_18),
.Y(n_61)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_61),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_44),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_62),
.Y(n_121)
);

INVx5_ASAP7_75t_L g63 ( 
.A(n_16),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g149 ( 
.A(n_63),
.Y(n_149)
);

BUFx5_ASAP7_75t_L g64 ( 
.A(n_45),
.Y(n_64)
);

INVx4_ASAP7_75t_L g116 ( 
.A(n_64),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g65 ( 
.A1(n_28),
.A2(n_10),
.B1(n_14),
.B2(n_3),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_65),
.B(n_70),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_44),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_66),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_44),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_67),
.B(n_75),
.Y(n_108)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_22),
.Y(n_68)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_68),
.Y(n_122)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_22),
.Y(n_69)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_69),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_23),
.B(n_10),
.Y(n_70)
);

INVx6_ASAP7_75t_L g71 ( 
.A(n_48),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_71),
.Y(n_134)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_23),
.Y(n_72)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_72),
.Y(n_138)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_29),
.Y(n_73)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_73),
.Y(n_142)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_25),
.Y(n_74)
);

INVx3_ASAP7_75t_L g148 ( 
.A(n_74),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_SL g75 ( 
.A1(n_29),
.A2(n_10),
.B(n_14),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_32),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_76),
.B(n_77),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_48),
.Y(n_77)
);

INVx5_ASAP7_75t_L g78 ( 
.A(n_16),
.Y(n_78)
);

INVx4_ASAP7_75t_L g123 ( 
.A(n_78),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_48),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_79),
.B(n_83),
.Y(n_137)
);

BUFx8_ASAP7_75t_L g80 ( 
.A(n_45),
.Y(n_80)
);

INVx13_ASAP7_75t_L g141 ( 
.A(n_80),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_48),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g151 ( 
.A(n_81),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_19),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g155 ( 
.A(n_82),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_19),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_19),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g162 ( 
.A(n_84),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_27),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_85),
.B(n_87),
.Y(n_154)
);

BUFx5_ASAP7_75t_L g86 ( 
.A(n_46),
.Y(n_86)
);

INVx4_ASAP7_75t_L g128 ( 
.A(n_86),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_27),
.Y(n_87)
);

BUFx5_ASAP7_75t_L g88 ( 
.A(n_46),
.Y(n_88)
);

BUFx12f_ASAP7_75t_L g107 ( 
.A(n_88),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_32),
.B(n_8),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_89),
.B(n_39),
.Y(n_139)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_25),
.Y(n_90)
);

INVx3_ASAP7_75t_L g152 ( 
.A(n_90),
.Y(n_152)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_25),
.Y(n_91)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_91),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_16),
.Y(n_92)
);

INVx6_ASAP7_75t_L g131 ( 
.A(n_92),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_47),
.Y(n_93)
);

INVx8_ASAP7_75t_L g130 ( 
.A(n_93),
.Y(n_130)
);

BUFx3_ASAP7_75t_L g94 ( 
.A(n_42),
.Y(n_94)
);

INVx5_ASAP7_75t_L g132 ( 
.A(n_94),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_47),
.Y(n_95)
);

INVx8_ASAP7_75t_L g156 ( 
.A(n_95),
.Y(n_156)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_21),
.Y(n_96)
);

INVx3_ASAP7_75t_L g153 ( 
.A(n_96),
.Y(n_153)
);

INVx1_ASAP7_75t_SL g97 ( 
.A(n_33),
.Y(n_97)
);

AND2x2_ASAP7_75t_L g113 ( 
.A(n_97),
.B(n_39),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_47),
.Y(n_98)
);

INVx5_ASAP7_75t_L g133 ( 
.A(n_98),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_42),
.Y(n_99)
);

INVx5_ASAP7_75t_L g159 ( 
.A(n_99),
.Y(n_159)
);

INVx6_ASAP7_75t_L g100 ( 
.A(n_33),
.Y(n_100)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_100),
.Y(n_158)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_42),
.Y(n_101)
);

BUFx12f_ASAP7_75t_L g140 ( 
.A(n_101),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_SL g103 ( 
.A(n_55),
.B(n_30),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_SL g194 ( 
.A(n_103),
.B(n_111),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_91),
.A2(n_30),
.B1(n_37),
.B2(n_34),
.Y(n_105)
);

OA22x2_ASAP7_75t_L g179 ( 
.A1(n_105),
.A2(n_114),
.B1(n_96),
.B2(n_63),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_80),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_80),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_112),
.B(n_118),
.Y(n_181)
);

INVx1_ASAP7_75t_SL g190 ( 
.A(n_113),
.Y(n_190)
);

AOI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_97),
.A2(n_41),
.B1(n_21),
.B2(n_33),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_54),
.B(n_34),
.Y(n_118)
);

AND2x2_ASAP7_75t_L g120 ( 
.A(n_58),
.B(n_35),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_120),
.B(n_127),
.Y(n_189)
);

CKINVDCx14_ASAP7_75t_R g124 ( 
.A(n_64),
.Y(n_124)
);

INVx2_ASAP7_75t_R g175 ( 
.A(n_124),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_SL g127 ( 
.A(n_60),
.B(n_26),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_100),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_136),
.B(n_157),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_139),
.B(n_163),
.Y(n_172)
);

BUFx12f_ASAP7_75t_L g147 ( 
.A(n_101),
.Y(n_147)
);

INVx4_ASAP7_75t_SL g166 ( 
.A(n_147),
.Y(n_166)
);

BUFx16f_ASAP7_75t_L g150 ( 
.A(n_50),
.Y(n_150)
);

BUFx12f_ASAP7_75t_L g187 ( 
.A(n_150),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_71),
.Y(n_157)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_51),
.Y(n_160)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_160),
.Y(n_168)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_73),
.Y(n_161)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_161),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_61),
.B(n_43),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_62),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_164),
.B(n_99),
.Y(n_196)
);

INVx11_ASAP7_75t_L g165 ( 
.A(n_150),
.Y(n_165)
);

INVx4_ASAP7_75t_L g216 ( 
.A(n_165),
.Y(n_216)
);

NAND2xp33_ASAP7_75t_SL g167 ( 
.A(n_113),
.B(n_75),
.Y(n_167)
);

INVx1_ASAP7_75t_SL g233 ( 
.A(n_167),
.Y(n_233)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_154),
.Y(n_169)
);

INVx1_ASAP7_75t_SL g240 ( 
.A(n_169),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_L g170 ( 
.A1(n_115),
.A2(n_65),
.B1(n_84),
.B2(n_82),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_170),
.A2(n_183),
.B1(n_207),
.B2(n_210),
.Y(n_232)
);

AOI22xp33_ASAP7_75t_SL g171 ( 
.A1(n_108),
.A2(n_41),
.B1(n_21),
.B2(n_38),
.Y(n_171)
);

INVxp67_ASAP7_75t_L g248 ( 
.A(n_171),
.Y(n_248)
);

INVx6_ASAP7_75t_L g173 ( 
.A(n_155),
.Y(n_173)
);

BUFx6f_ASAP7_75t_L g219 ( 
.A(n_173),
.Y(n_219)
);

INVx4_ASAP7_75t_L g174 ( 
.A(n_123),
.Y(n_174)
);

BUFx2_ASAP7_75t_L g250 ( 
.A(n_174),
.Y(n_250)
);

INVx4_ASAP7_75t_L g176 ( 
.A(n_123),
.Y(n_176)
);

INVx3_ASAP7_75t_L g236 ( 
.A(n_176),
.Y(n_236)
);

INVx3_ASAP7_75t_L g177 ( 
.A(n_132),
.Y(n_177)
);

BUFx3_ASAP7_75t_L g242 ( 
.A(n_177),
.Y(n_242)
);

AOI22xp33_ASAP7_75t_L g178 ( 
.A1(n_110),
.A2(n_40),
.B1(n_36),
.B2(n_68),
.Y(n_178)
);

AOI22xp33_ASAP7_75t_SL g220 ( 
.A1(n_178),
.A2(n_203),
.B1(n_209),
.B2(n_213),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_179),
.A2(n_78),
.B1(n_94),
.B2(n_133),
.Y(n_235)
);

INVx3_ASAP7_75t_SL g182 ( 
.A(n_130),
.Y(n_182)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_182),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_102),
.A2(n_81),
.B1(n_66),
.B2(n_69),
.Y(n_183)
);

BUFx3_ASAP7_75t_L g184 ( 
.A(n_132),
.Y(n_184)
);

INVx5_ASAP7_75t_L g224 ( 
.A(n_184),
.Y(n_224)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_117),
.Y(n_185)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_185),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_137),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_SL g251 ( 
.A(n_186),
.B(n_192),
.Y(n_251)
);

INVx3_ASAP7_75t_L g188 ( 
.A(n_149),
.Y(n_188)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_188),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_143),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_146),
.Y(n_193)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_193),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_106),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_195),
.B(n_205),
.Y(n_243)
);

CKINVDCx14_ASAP7_75t_R g215 ( 
.A(n_196),
.Y(n_215)
);

INVx3_ASAP7_75t_L g197 ( 
.A(n_149),
.Y(n_197)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_197),
.Y(n_237)
);

INVx1_ASAP7_75t_SL g198 ( 
.A(n_141),
.Y(n_198)
);

AND2x2_ASAP7_75t_L g245 ( 
.A(n_198),
.B(n_212),
.Y(n_245)
);

HB1xp67_ASAP7_75t_L g199 ( 
.A(n_145),
.Y(n_199)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_199),
.Y(n_244)
);

INVx4_ASAP7_75t_L g200 ( 
.A(n_135),
.Y(n_200)
);

BUFx6f_ASAP7_75t_L g223 ( 
.A(n_200),
.Y(n_223)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_158),
.Y(n_201)
);

BUFx6f_ASAP7_75t_L g229 ( 
.A(n_201),
.Y(n_229)
);

BUFx12f_ASAP7_75t_L g202 ( 
.A(n_141),
.Y(n_202)
);

INVx11_ASAP7_75t_L g218 ( 
.A(n_202),
.Y(n_218)
);

INVx8_ASAP7_75t_L g203 ( 
.A(n_140),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_119),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_204),
.B(n_206),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_122),
.B(n_72),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_125),
.B(n_43),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_109),
.A2(n_98),
.B1(n_95),
.B2(n_92),
.Y(n_207)
);

BUFx12f_ASAP7_75t_L g208 ( 
.A(n_130),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_208),
.B(n_211),
.Y(n_246)
);

AOI22xp33_ASAP7_75t_L g209 ( 
.A1(n_138),
.A2(n_36),
.B1(n_40),
.B2(n_37),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_142),
.A2(n_90),
.B1(n_49),
.B2(n_52),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_131),
.Y(n_211)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_145),
.Y(n_212)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_129),
.Y(n_213)
);

INVx4_ASAP7_75t_L g214 ( 
.A(n_135),
.Y(n_214)
);

OR2x2_ASAP7_75t_L g225 ( 
.A(n_214),
.B(n_116),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_167),
.B(n_144),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_217),
.B(n_222),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_191),
.B(n_120),
.Y(n_222)
);

CKINVDCx16_ASAP7_75t_R g265 ( 
.A(n_225),
.Y(n_265)
);

OR2x2_ASAP7_75t_L g227 ( 
.A(n_190),
.B(n_116),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_227),
.B(n_241),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_172),
.B(n_129),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_230),
.B(n_231),
.Y(n_260)
);

AO22x1_ASAP7_75t_SL g231 ( 
.A1(n_190),
.A2(n_148),
.B1(n_152),
.B2(n_74),
.Y(n_231)
);

OAI22xp33_ASAP7_75t_L g234 ( 
.A1(n_183),
.A2(n_114),
.B1(n_131),
.B2(n_159),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_234),
.A2(n_232),
.B1(n_207),
.B2(n_217),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_L g271 ( 
.A1(n_235),
.A2(n_179),
.B1(n_107),
.B2(n_128),
.Y(n_271)
);

OR2x2_ASAP7_75t_L g241 ( 
.A(n_194),
.B(n_152),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_189),
.B(n_93),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_247),
.B(n_249),
.C(n_198),
.Y(n_261)
);

OAI21xp5_ASAP7_75t_SL g249 ( 
.A1(n_181),
.A2(n_148),
.B(n_153),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_L g291 ( 
.A1(n_252),
.A2(n_255),
.B1(n_269),
.B2(n_277),
.Y(n_291)
);

INVxp67_ASAP7_75t_L g253 ( 
.A(n_245),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_253),
.B(n_261),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_232),
.A2(n_179),
.B1(n_210),
.B2(n_134),
.Y(n_255)
);

INVx13_ASAP7_75t_L g256 ( 
.A(n_218),
.Y(n_256)
);

INVx1_ASAP7_75t_SL g300 ( 
.A(n_256),
.Y(n_300)
);

INVx13_ASAP7_75t_L g257 ( 
.A(n_218),
.Y(n_257)
);

INVxp67_ASAP7_75t_L g311 ( 
.A(n_257),
.Y(n_311)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_229),
.Y(n_258)
);

INVx2_ASAP7_75t_L g303 ( 
.A(n_258),
.Y(n_303)
);

CKINVDCx10_ASAP7_75t_R g259 ( 
.A(n_216),
.Y(n_259)
);

CKINVDCx16_ASAP7_75t_R g314 ( 
.A(n_259),
.Y(n_314)
);

BUFx6f_ASAP7_75t_L g262 ( 
.A(n_219),
.Y(n_262)
);

INVx4_ASAP7_75t_L g294 ( 
.A(n_262),
.Y(n_294)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_245),
.Y(n_263)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_263),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_SL g264 ( 
.A(n_233),
.B(n_175),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g284 ( 
.A(n_264),
.B(n_247),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_251),
.B(n_240),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_SL g285 ( 
.A(n_266),
.B(n_281),
.Y(n_285)
);

BUFx6f_ASAP7_75t_L g267 ( 
.A(n_219),
.Y(n_267)
);

INVx4_ASAP7_75t_L g308 ( 
.A(n_267),
.Y(n_308)
);

INVx4_ASAP7_75t_L g268 ( 
.A(n_221),
.Y(n_268)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_268),
.Y(n_299)
);

AOI22xp33_ASAP7_75t_SL g269 ( 
.A1(n_248),
.A2(n_177),
.B1(n_184),
.B2(n_197),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_271),
.A2(n_276),
.B1(n_166),
.B2(n_182),
.Y(n_304)
);

INVx13_ASAP7_75t_L g272 ( 
.A(n_216),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_272),
.Y(n_288)
);

CKINVDCx16_ASAP7_75t_R g273 ( 
.A(n_245),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_273),
.B(n_274),
.Y(n_287)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_229),
.Y(n_274)
);

CKINVDCx10_ASAP7_75t_R g275 ( 
.A(n_225),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_275),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_233),
.A2(n_179),
.B1(n_134),
.B2(n_155),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_L g277 ( 
.A1(n_235),
.A2(n_248),
.B1(n_230),
.B2(n_215),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_239),
.B(n_180),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_278),
.B(n_279),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_243),
.B(n_180),
.Y(n_279)
);

A2O1A1Ixp33_ASAP7_75t_L g280 ( 
.A1(n_222),
.A2(n_175),
.B(n_168),
.C(n_212),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_280),
.B(n_202),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_240),
.B(n_202),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_228),
.B(n_168),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_SL g306 ( 
.A(n_282),
.B(n_221),
.Y(n_306)
);

INVx13_ASAP7_75t_L g283 ( 
.A(n_224),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_283),
.Y(n_310)
);

XOR2xp5_ASAP7_75t_L g319 ( 
.A(n_284),
.B(n_312),
.Y(n_319)
);

MAJx2_ASAP7_75t_L g286 ( 
.A(n_264),
.B(n_241),
.C(n_227),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_286),
.B(n_290),
.C(n_297),
.Y(n_329)
);

XOR2xp5_ASAP7_75t_SL g289 ( 
.A(n_254),
.B(n_249),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_SL g324 ( 
.A(n_289),
.B(n_259),
.C(n_282),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_254),
.B(n_238),
.C(n_246),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_L g292 ( 
.A1(n_252),
.A2(n_220),
.B1(n_234),
.B2(n_231),
.Y(n_292)
);

AND2x2_ASAP7_75t_L g339 ( 
.A(n_292),
.B(n_208),
.Y(n_339)
);

OAI21xp5_ASAP7_75t_L g296 ( 
.A1(n_270),
.A2(n_244),
.B(n_231),
.Y(n_296)
);

OAI21xp5_ASAP7_75t_SL g317 ( 
.A1(n_296),
.A2(n_309),
.B(n_313),
.Y(n_317)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_261),
.B(n_244),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_255),
.A2(n_173),
.B1(n_162),
.B2(n_121),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_301),
.B(n_307),
.Y(n_326)
);

AOI21xp5_ASAP7_75t_L g302 ( 
.A1(n_275),
.A2(n_226),
.B(n_237),
.Y(n_302)
);

AOI21xp5_ASAP7_75t_L g333 ( 
.A1(n_302),
.A2(n_257),
.B(n_256),
.Y(n_333)
);

OAI22xp5_ASAP7_75t_L g318 ( 
.A1(n_304),
.A2(n_271),
.B1(n_260),
.B2(n_265),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_306),
.B(n_268),
.Y(n_325)
);

AO22x1_ASAP7_75t_L g307 ( 
.A1(n_277),
.A2(n_237),
.B1(n_226),
.B2(n_201),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_273),
.B(n_263),
.C(n_279),
.Y(n_312)
);

AOI21xp5_ASAP7_75t_SL g313 ( 
.A1(n_270),
.A2(n_250),
.B(n_38),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_SL g315 ( 
.A1(n_260),
.A2(n_162),
.B1(n_121),
.B2(n_126),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_315),
.B(n_301),
.Y(n_343)
);

BUFx24_ASAP7_75t_SL g316 ( 
.A(n_285),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_SL g362 ( 
.A(n_316),
.B(n_335),
.Y(n_362)
);

OAI22xp5_ASAP7_75t_L g361 ( 
.A1(n_318),
.A2(n_339),
.B1(n_313),
.B2(n_310),
.Y(n_361)
);

OAI22xp5_ASAP7_75t_SL g320 ( 
.A1(n_304),
.A2(n_265),
.B1(n_276),
.B2(n_278),
.Y(n_320)
);

AOI22xp5_ASAP7_75t_L g377 ( 
.A1(n_320),
.A2(n_328),
.B1(n_315),
.B2(n_310),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_SL g321 ( 
.A(n_298),
.B(n_280),
.Y(n_321)
);

CKINVDCx14_ASAP7_75t_R g380 ( 
.A(n_321),
.Y(n_380)
);

INVxp67_ASAP7_75t_L g322 ( 
.A(n_309),
.Y(n_322)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_322),
.Y(n_353)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_298),
.Y(n_323)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_323),
.Y(n_368)
);

XNOR2xp5_ASAP7_75t_L g350 ( 
.A(n_324),
.B(n_286),
.Y(n_350)
);

OAI21xp33_ASAP7_75t_SL g357 ( 
.A1(n_325),
.A2(n_332),
.B(n_340),
.Y(n_357)
);

INVx13_ASAP7_75t_L g327 ( 
.A(n_300),
.Y(n_327)
);

INVx1_ASAP7_75t_SL g360 ( 
.A(n_327),
.Y(n_360)
);

OAI22xp5_ASAP7_75t_SL g328 ( 
.A1(n_293),
.A2(n_267),
.B1(n_262),
.B2(n_258),
.Y(n_328)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_287),
.Y(n_330)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_330),
.Y(n_370)
);

OAI32xp33_ASAP7_75t_L g331 ( 
.A1(n_293),
.A2(n_274),
.A3(n_213),
.B1(n_272),
.B2(n_256),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_331),
.B(n_336),
.Y(n_366)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_290),
.B(n_242),
.Y(n_332)
);

NAND2xp33_ASAP7_75t_SL g372 ( 
.A(n_333),
.B(n_334),
.Y(n_372)
);

NAND2x1p5_ASAP7_75t_L g334 ( 
.A(n_287),
.B(n_236),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_SL g335 ( 
.A(n_295),
.B(n_242),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g336 ( 
.A(n_302),
.Y(n_336)
);

CKINVDCx20_ASAP7_75t_R g337 ( 
.A(n_311),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_337),
.B(n_345),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_SL g338 ( 
.A(n_312),
.B(n_289),
.Y(n_338)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_338),
.Y(n_371)
);

AOI21xp5_ASAP7_75t_L g340 ( 
.A1(n_295),
.A2(n_257),
.B(n_272),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_303),
.Y(n_341)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_341),
.Y(n_374)
);

INVx13_ASAP7_75t_L g342 ( 
.A(n_300),
.Y(n_342)
);

INVx4_ASAP7_75t_L g363 ( 
.A(n_342),
.Y(n_363)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_343),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_296),
.B(n_267),
.Y(n_344)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_344),
.Y(n_356)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_299),
.B(n_236),
.Y(n_345)
);

CKINVDCx20_ASAP7_75t_R g346 ( 
.A(n_311),
.Y(n_346)
);

NOR2xp33_ASAP7_75t_L g354 ( 
.A(n_346),
.B(n_314),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_307),
.B(n_262),
.Y(n_347)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_347),
.Y(n_365)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_303),
.Y(n_348)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_348),
.Y(n_379)
);

XNOR2x2_ASAP7_75t_SL g397 ( 
.A(n_350),
.B(n_334),
.Y(n_397)
);

MAJIxp5_ASAP7_75t_L g351 ( 
.A(n_319),
.B(n_329),
.C(n_297),
.Y(n_351)
);

MAJIxp5_ASAP7_75t_L g394 ( 
.A(n_351),
.B(n_352),
.C(n_364),
.Y(n_394)
);

MAJIxp5_ASAP7_75t_L g352 ( 
.A(n_319),
.B(n_329),
.C(n_338),
.Y(n_352)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_354),
.Y(n_386)
);

OAI22xp5_ASAP7_75t_SL g355 ( 
.A1(n_330),
.A2(n_336),
.B1(n_339),
.B2(n_321),
.Y(n_355)
);

AOI22xp5_ASAP7_75t_SL g400 ( 
.A1(n_355),
.A2(n_358),
.B1(n_361),
.B2(n_331),
.Y(n_400)
);

OAI22xp5_ASAP7_75t_SL g358 ( 
.A1(n_339),
.A2(n_291),
.B1(n_305),
.B2(n_307),
.Y(n_358)
);

XNOR2x2_ASAP7_75t_SL g359 ( 
.A(n_324),
.B(n_284),
.Y(n_359)
);

XNOR2xp5_ASAP7_75t_L g383 ( 
.A(n_359),
.B(n_317),
.Y(n_383)
);

MAJIxp5_ASAP7_75t_L g364 ( 
.A(n_332),
.B(n_323),
.C(n_318),
.Y(n_364)
);

AND2x2_ASAP7_75t_L g367 ( 
.A(n_337),
.B(n_288),
.Y(n_367)
);

CKINVDCx20_ASAP7_75t_R g385 ( 
.A(n_367),
.Y(n_385)
);

CKINVDCx16_ASAP7_75t_R g369 ( 
.A(n_345),
.Y(n_369)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_369),
.Y(n_387)
);

CKINVDCx20_ASAP7_75t_R g375 ( 
.A(n_335),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_SL g408 ( 
.A(n_375),
.B(n_283),
.Y(n_408)
);

OAI22xp5_ASAP7_75t_L g376 ( 
.A1(n_343),
.A2(n_326),
.B1(n_347),
.B2(n_344),
.Y(n_376)
);

OAI22xp5_ASAP7_75t_L g391 ( 
.A1(n_376),
.A2(n_377),
.B1(n_381),
.B2(n_346),
.Y(n_391)
);

MAJIxp5_ASAP7_75t_L g378 ( 
.A(n_334),
.B(n_299),
.C(n_188),
.Y(n_378)
);

MAJIxp5_ASAP7_75t_L g398 ( 
.A(n_378),
.B(n_334),
.C(n_342),
.Y(n_398)
);

OAI22xp5_ASAP7_75t_L g381 ( 
.A1(n_326),
.A2(n_288),
.B1(n_294),
.B2(n_308),
.Y(n_381)
);

AOI22xp5_ASAP7_75t_L g382 ( 
.A1(n_320),
.A2(n_308),
.B1(n_294),
.B2(n_224),
.Y(n_382)
);

OAI22xp5_ASAP7_75t_SL g396 ( 
.A1(n_382),
.A2(n_341),
.B1(n_342),
.B2(n_327),
.Y(n_396)
);

XNOR2xp5_ASAP7_75t_SL g429 ( 
.A(n_383),
.B(n_388),
.Y(n_429)
);

INVx2_ASAP7_75t_SL g384 ( 
.A(n_367),
.Y(n_384)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_384),
.Y(n_416)
);

XNOR2xp5_ASAP7_75t_SL g388 ( 
.A(n_350),
.B(n_317),
.Y(n_388)
);

OAI21xp5_ASAP7_75t_SL g389 ( 
.A1(n_371),
.A2(n_333),
.B(n_340),
.Y(n_389)
);

CKINVDCx14_ASAP7_75t_R g420 ( 
.A(n_389),
.Y(n_420)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_373),
.Y(n_390)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_390),
.Y(n_418)
);

OAI22xp5_ASAP7_75t_L g415 ( 
.A1(n_391),
.A2(n_406),
.B1(n_408),
.B2(n_387),
.Y(n_415)
);

MAJIxp5_ASAP7_75t_SL g392 ( 
.A(n_352),
.B(n_328),
.C(n_348),
.Y(n_392)
);

OAI22xp5_ASAP7_75t_SL g427 ( 
.A1(n_392),
.A2(n_360),
.B1(n_363),
.B2(n_379),
.Y(n_427)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_373),
.Y(n_393)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_393),
.Y(n_423)
);

XNOR2xp5_ASAP7_75t_L g395 ( 
.A(n_351),
.B(n_325),
.Y(n_395)
);

XNOR2xp5_ASAP7_75t_L g430 ( 
.A(n_395),
.B(n_397),
.Y(n_430)
);

HB1xp67_ASAP7_75t_L g414 ( 
.A(n_396),
.Y(n_414)
);

XNOR2xp5_ASAP7_75t_L g436 ( 
.A(n_398),
.B(n_403),
.Y(n_436)
);

XNOR2xp5_ASAP7_75t_L g399 ( 
.A(n_359),
.B(n_250),
.Y(n_399)
);

HB1xp67_ASAP7_75t_L g425 ( 
.A(n_399),
.Y(n_425)
);

OAI22xp5_ASAP7_75t_SL g424 ( 
.A1(n_400),
.A2(n_349),
.B1(n_382),
.B2(n_377),
.Y(n_424)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_367),
.Y(n_401)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_401),
.Y(n_431)
);

XNOR2xp5_ASAP7_75t_L g402 ( 
.A(n_364),
.B(n_223),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_SL g421 ( 
.A(n_402),
.B(n_374),
.Y(n_421)
);

XNOR2xp5_ASAP7_75t_L g403 ( 
.A(n_353),
.B(n_223),
.Y(n_403)
);

HB1xp67_ASAP7_75t_L g404 ( 
.A(n_366),
.Y(n_404)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_404),
.Y(n_434)
);

XOR2xp5_ASAP7_75t_L g405 ( 
.A(n_355),
.B(n_370),
.Y(n_405)
);

XOR2xp5_ASAP7_75t_L g417 ( 
.A(n_405),
.B(n_409),
.Y(n_417)
);

OAI22xp5_ASAP7_75t_L g406 ( 
.A1(n_380),
.A2(n_327),
.B1(n_26),
.B2(n_208),
.Y(n_406)
);

MAJIxp5_ASAP7_75t_L g407 ( 
.A(n_358),
.B(n_174),
.C(n_176),
.Y(n_407)
);

MAJIxp5_ASAP7_75t_L g428 ( 
.A(n_407),
.B(n_410),
.C(n_411),
.Y(n_428)
);

XOR2xp5_ASAP7_75t_L g409 ( 
.A(n_357),
.B(n_283),
.Y(n_409)
);

MAJIxp5_ASAP7_75t_L g410 ( 
.A(n_356),
.B(n_166),
.C(n_214),
.Y(n_410)
);

MAJIxp5_ASAP7_75t_L g411 ( 
.A(n_356),
.B(n_200),
.C(n_128),
.Y(n_411)
);

XOR2xp5_ASAP7_75t_L g412 ( 
.A(n_366),
.B(n_203),
.Y(n_412)
);

XOR2xp5_ASAP7_75t_L g426 ( 
.A(n_412),
.B(n_372),
.Y(n_426)
);

MAJIxp5_ASAP7_75t_L g413 ( 
.A(n_378),
.B(n_104),
.C(n_153),
.Y(n_413)
);

MAJIxp5_ASAP7_75t_L g432 ( 
.A(n_413),
.B(n_360),
.C(n_379),
.Y(n_432)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_415),
.Y(n_441)
);

XNOR2x1_ASAP7_75t_L g419 ( 
.A(n_405),
.B(n_365),
.Y(n_419)
);

XOR2xp5_ASAP7_75t_L g442 ( 
.A(n_419),
.B(n_412),
.Y(n_442)
);

XNOR2xp5_ASAP7_75t_L g449 ( 
.A(n_421),
.B(n_426),
.Y(n_449)
);

A2O1A1Ixp33_ASAP7_75t_L g422 ( 
.A1(n_385),
.A2(n_372),
.B(n_365),
.C(n_349),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_422),
.B(n_435),
.Y(n_448)
);

AOI22xp5_ASAP7_75t_L g447 ( 
.A1(n_424),
.A2(n_440),
.B1(n_407),
.B2(n_409),
.Y(n_447)
);

NOR2xp33_ASAP7_75t_L g450 ( 
.A(n_427),
.B(n_398),
.Y(n_450)
);

XNOR2xp5_ASAP7_75t_L g463 ( 
.A(n_432),
.B(n_147),
.Y(n_463)
);

MAJIxp5_ASAP7_75t_L g433 ( 
.A(n_394),
.B(n_368),
.C(n_363),
.Y(n_433)
);

MAJIxp5_ASAP7_75t_L g458 ( 
.A(n_433),
.B(n_187),
.C(n_165),
.Y(n_458)
);

CKINVDCx14_ASAP7_75t_R g435 ( 
.A(n_410),
.Y(n_435)
);

INVxp67_ASAP7_75t_L g437 ( 
.A(n_403),
.Y(n_437)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_437),
.Y(n_453)
);

OAI22xp5_ASAP7_75t_SL g438 ( 
.A1(n_400),
.A2(n_362),
.B1(n_151),
.B2(n_126),
.Y(n_438)
);

INVxp67_ASAP7_75t_L g445 ( 
.A(n_438),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_SL g439 ( 
.A(n_386),
.B(n_187),
.Y(n_439)
);

NOR2xp33_ASAP7_75t_SL g461 ( 
.A(n_439),
.B(n_11),
.Y(n_461)
);

OAI22xp5_ASAP7_75t_SL g440 ( 
.A1(n_384),
.A2(n_151),
.B1(n_159),
.B2(n_133),
.Y(n_440)
);

XOR2xp5_ASAP7_75t_L g465 ( 
.A(n_442),
.B(n_417),
.Y(n_465)
);

CKINVDCx20_ASAP7_75t_R g443 ( 
.A(n_420),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_SL g469 ( 
.A(n_443),
.B(n_456),
.Y(n_469)
);

XOR2xp5_ASAP7_75t_L g444 ( 
.A(n_436),
.B(n_395),
.Y(n_444)
);

XNOR2xp5_ASAP7_75t_L g483 ( 
.A(n_444),
.B(n_463),
.Y(n_483)
);

INVx2_ASAP7_75t_L g446 ( 
.A(n_416),
.Y(n_446)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_446),
.Y(n_470)
);

OAI22xp5_ASAP7_75t_SL g467 ( 
.A1(n_447),
.A2(n_457),
.B1(n_437),
.B2(n_440),
.Y(n_467)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_450),
.Y(n_472)
);

AOI221xp5_ASAP7_75t_L g451 ( 
.A1(n_418),
.A2(n_394),
.B1(n_397),
.B2(n_388),
.C(n_411),
.Y(n_451)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_451),
.Y(n_477)
);

AOI21xp5_ASAP7_75t_L g452 ( 
.A1(n_422),
.A2(n_413),
.B(n_104),
.Y(n_452)
);

OAI21xp5_ASAP7_75t_L g468 ( 
.A1(n_452),
.A2(n_459),
.B(n_457),
.Y(n_468)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_431),
.Y(n_454)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_454),
.Y(n_479)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_434),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g473 ( 
.A(n_455),
.B(n_462),
.Y(n_473)
);

CKINVDCx20_ASAP7_75t_R g456 ( 
.A(n_414),
.Y(n_456)
);

AOI22xp5_ASAP7_75t_L g457 ( 
.A1(n_424),
.A2(n_156),
.B1(n_140),
.B2(n_147),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_SL g476 ( 
.A(n_458),
.B(n_460),
.Y(n_476)
);

OAI21xp5_ASAP7_75t_SL g459 ( 
.A1(n_423),
.A2(n_187),
.B(n_156),
.Y(n_459)
);

AO221x1_ASAP7_75t_L g460 ( 
.A1(n_433),
.A2(n_27),
.B1(n_31),
.B2(n_107),
.C(n_41),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_SL g481 ( 
.A(n_461),
.B(n_12),
.Y(n_481)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_432),
.Y(n_462)
);

AOI211xp5_ASAP7_75t_L g464 ( 
.A1(n_448),
.A2(n_419),
.B(n_425),
.C(n_426),
.Y(n_464)
);

AOI22xp5_ASAP7_75t_L g495 ( 
.A1(n_464),
.A2(n_466),
.B1(n_13),
.B2(n_15),
.Y(n_495)
);

XOR2xp5_ASAP7_75t_L g497 ( 
.A(n_465),
.B(n_467),
.Y(n_497)
);

INVxp67_ASAP7_75t_SL g466 ( 
.A(n_441),
.Y(n_466)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_468),
.Y(n_489)
);

MAJIxp5_ASAP7_75t_L g471 ( 
.A(n_444),
.B(n_436),
.C(n_428),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_471),
.B(n_474),
.Y(n_494)
);

MAJIxp5_ASAP7_75t_L g474 ( 
.A(n_463),
.B(n_428),
.C(n_430),
.Y(n_474)
);

MAJIxp5_ASAP7_75t_L g475 ( 
.A(n_453),
.B(n_430),
.C(n_417),
.Y(n_475)
);

MAJIxp5_ASAP7_75t_L g492 ( 
.A(n_475),
.B(n_445),
.C(n_140),
.Y(n_492)
);

XOR2xp5_ASAP7_75t_L g478 ( 
.A(n_449),
.B(n_429),
.Y(n_478)
);

AND2x2_ASAP7_75t_L g490 ( 
.A(n_478),
.B(n_458),
.Y(n_490)
);

CKINVDCx20_ASAP7_75t_R g480 ( 
.A(n_448),
.Y(n_480)
);

NOR2xp33_ASAP7_75t_SL g484 ( 
.A(n_480),
.B(n_481),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_L g482 ( 
.A(n_446),
.B(n_429),
.Y(n_482)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_482),
.Y(n_496)
);

XNOR2xp5_ASAP7_75t_L g485 ( 
.A(n_471),
.B(n_449),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_L g513 ( 
.A(n_485),
.B(n_488),
.Y(n_513)
);

OAI21xp5_ASAP7_75t_L g486 ( 
.A1(n_482),
.A2(n_442),
.B(n_452),
.Y(n_486)
);

AOI21xp5_ASAP7_75t_L g511 ( 
.A1(n_486),
.A2(n_500),
.B(n_464),
.Y(n_511)
);

AOI21xp33_ASAP7_75t_L g487 ( 
.A1(n_473),
.A2(n_447),
.B(n_459),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_L g504 ( 
.A(n_487),
.B(n_491),
.Y(n_504)
);

XNOR2xp5_ASAP7_75t_L g488 ( 
.A(n_472),
.B(n_483),
.Y(n_488)
);

XOR2xp5_ASAP7_75t_L g512 ( 
.A(n_490),
.B(n_31),
.Y(n_512)
);

XNOR2xp5_ASAP7_75t_L g491 ( 
.A(n_483),
.B(n_445),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_SL g503 ( 
.A(n_492),
.B(n_498),
.Y(n_503)
);

OAI22xp5_ASAP7_75t_SL g493 ( 
.A1(n_477),
.A2(n_107),
.B1(n_35),
.B2(n_56),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_L g507 ( 
.A(n_493),
.B(n_499),
.Y(n_507)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_495),
.Y(n_505)
);

NOR2xp33_ASAP7_75t_SL g498 ( 
.A(n_469),
.B(n_13),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_470),
.Y(n_499)
);

AOI21xp5_ASAP7_75t_L g500 ( 
.A1(n_473),
.A2(n_88),
.B(n_86),
.Y(n_500)
);

OAI22xp5_ASAP7_75t_L g501 ( 
.A1(n_489),
.A2(n_468),
.B1(n_479),
.B2(n_474),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_501),
.B(n_502),
.Y(n_515)
);

MAJIxp5_ASAP7_75t_L g502 ( 
.A(n_494),
.B(n_475),
.C(n_465),
.Y(n_502)
);

NOR2xp33_ASAP7_75t_SL g506 ( 
.A(n_488),
.B(n_478),
.Y(n_506)
);

CKINVDCx20_ASAP7_75t_R g517 ( 
.A(n_506),
.Y(n_517)
);

CKINVDCx20_ASAP7_75t_R g508 ( 
.A(n_484),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_L g522 ( 
.A(n_508),
.B(n_509),
.Y(n_522)
);

NOR2xp33_ASAP7_75t_L g509 ( 
.A(n_485),
.B(n_467),
.Y(n_509)
);

NOR2xp33_ASAP7_75t_L g510 ( 
.A(n_491),
.B(n_476),
.Y(n_510)
);

AOI21xp5_ASAP7_75t_L g519 ( 
.A1(n_510),
.A2(n_514),
.B(n_486),
.Y(n_519)
);

XNOR2xp5_ASAP7_75t_L g520 ( 
.A(n_511),
.B(n_512),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_SL g514 ( 
.A(n_497),
.B(n_35),
.Y(n_514)
);

MAJIxp5_ASAP7_75t_L g516 ( 
.A(n_513),
.B(n_497),
.C(n_490),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_SL g531 ( 
.A(n_516),
.B(n_518),
.Y(n_531)
);

OAI21xp33_ASAP7_75t_L g518 ( 
.A1(n_504),
.A2(n_496),
.B(n_492),
.Y(n_518)
);

NOR2xp33_ASAP7_75t_L g526 ( 
.A(n_519),
.B(n_521),
.Y(n_526)
);

NOR2xp33_ASAP7_75t_L g521 ( 
.A(n_513),
.B(n_35),
.Y(n_521)
);

XNOR2xp5_ASAP7_75t_L g523 ( 
.A(n_502),
.B(n_31),
.Y(n_523)
);

MAJIxp5_ASAP7_75t_L g525 ( 
.A(n_523),
.B(n_524),
.C(n_522),
.Y(n_525)
);

AOI322xp5_ASAP7_75t_L g524 ( 
.A1(n_507),
.A2(n_31),
.A3(n_27),
.B1(n_35),
.B2(n_6),
.C1(n_8),
.C2(n_11),
.Y(n_524)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_525),
.Y(n_534)
);

MAJIxp5_ASAP7_75t_L g527 ( 
.A(n_517),
.B(n_511),
.C(n_505),
.Y(n_527)
);

OAI21xp5_ASAP7_75t_L g535 ( 
.A1(n_527),
.A2(n_529),
.B(n_530),
.Y(n_535)
);

A2O1A1O1Ixp25_ASAP7_75t_SL g528 ( 
.A1(n_518),
.A2(n_512),
.B(n_503),
.C(n_4),
.D(n_6),
.Y(n_528)
);

AOI322xp5_ASAP7_75t_L g532 ( 
.A1(n_528),
.A2(n_520),
.A3(n_11),
.B1(n_6),
.B2(n_8),
.C1(n_12),
.C2(n_13),
.Y(n_532)
);

MAJIxp5_ASAP7_75t_L g529 ( 
.A(n_515),
.B(n_31),
.C(n_27),
.Y(n_529)
);

OAI21xp5_ASAP7_75t_SL g530 ( 
.A1(n_516),
.A2(n_31),
.B(n_27),
.Y(n_530)
);

AO21x1_ASAP7_75t_L g536 ( 
.A1(n_532),
.A2(n_526),
.B(n_0),
.Y(n_536)
);

OAI22xp5_ASAP7_75t_L g533 ( 
.A1(n_531),
.A2(n_11),
.B1(n_15),
.B2(n_0),
.Y(n_533)
);

MAJIxp5_ASAP7_75t_L g537 ( 
.A(n_533),
.B(n_526),
.C(n_1),
.Y(n_537)
);

MAJIxp5_ASAP7_75t_L g538 ( 
.A(n_536),
.B(n_537),
.C(n_535),
.Y(n_538)
);

OAI21xp5_ASAP7_75t_SL g539 ( 
.A1(n_538),
.A2(n_534),
.B(n_1),
.Y(n_539)
);

XOR2xp5_ASAP7_75t_L g540 ( 
.A(n_539),
.B(n_1),
.Y(n_540)
);

NOR2xp33_ASAP7_75t_L g541 ( 
.A(n_540),
.B(n_1),
.Y(n_541)
);


endmodule