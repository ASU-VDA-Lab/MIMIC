module fake_jpeg_3358_n_644 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_644);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_644;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_620;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_635;
wire n_517;
wire n_629;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_643;
wire n_170;
wire n_602;
wire n_313;
wire n_574;
wire n_542;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_641;
wire n_48;
wire n_465;
wire n_638;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_623;
wire n_579;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_637;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_624;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_634;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_639;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_622;
wire n_463;
wire n_92;
wire n_332;
wire n_640;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_626;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_642;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_615;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_631;
wire n_433;
wire n_636;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_599;
wire n_239;
wire n_243;
wire n_481;
wire n_628;
wire n_619;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_625;
wire n_147;
wire n_449;
wire n_627;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_613;
wire n_630;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_633;
wire n_112;
wire n_632;
wire n_616;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_621;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_2),
.Y(n_20)
);

BUFx6f_ASAP7_75t_SL g21 ( 
.A(n_1),
.Y(n_21)
);

INVx4_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_0),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_17),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_14),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_13),
.Y(n_29)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

INVx13_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_16),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_2),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_4),
.Y(n_34)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_13),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_16),
.Y(n_36)
);

INVx13_ASAP7_75t_L g37 ( 
.A(n_11),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_9),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_1),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_11),
.Y(n_40)
);

CKINVDCx14_ASAP7_75t_R g41 ( 
.A(n_14),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_16),
.Y(n_42)
);

INVx2_ASAP7_75t_R g43 ( 
.A(n_11),
.Y(n_43)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_9),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_18),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_0),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_10),
.Y(n_47)
);

BUFx24_ASAP7_75t_L g48 ( 
.A(n_10),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_9),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_5),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_7),
.Y(n_51)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_14),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_14),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_8),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_16),
.Y(n_55)
);

INVx13_ASAP7_75t_L g56 ( 
.A(n_6),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_4),
.Y(n_57)
);

BUFx5_ASAP7_75t_L g58 ( 
.A(n_48),
.Y(n_58)
);

INVx4_ASAP7_75t_L g137 ( 
.A(n_58),
.Y(n_137)
);

BUFx5_ASAP7_75t_L g59 ( 
.A(n_48),
.Y(n_59)
);

INVx4_ASAP7_75t_L g142 ( 
.A(n_59),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_23),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_60),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_23),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g157 ( 
.A(n_61),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_52),
.B(n_19),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_62),
.B(n_74),
.Y(n_153)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_44),
.Y(n_63)
);

INVx4_ASAP7_75t_SL g191 ( 
.A(n_63),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_23),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_64),
.B(n_69),
.Y(n_131)
);

INVx4_ASAP7_75t_SL g65 ( 
.A(n_32),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g202 ( 
.A(n_65),
.Y(n_202)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_23),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g171 ( 
.A(n_66),
.Y(n_171)
);

INVx5_ASAP7_75t_L g67 ( 
.A(n_44),
.Y(n_67)
);

BUFx2_ASAP7_75t_L g208 ( 
.A(n_67),
.Y(n_208)
);

INVx8_ASAP7_75t_L g68 ( 
.A(n_57),
.Y(n_68)
);

INVx5_ASAP7_75t_L g160 ( 
.A(n_68),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_57),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_39),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g180 ( 
.A(n_70),
.Y(n_180)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_39),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g196 ( 
.A(n_71),
.Y(n_196)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_52),
.Y(n_72)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_72),
.Y(n_144)
);

BUFx3_ASAP7_75t_L g73 ( 
.A(n_55),
.Y(n_73)
);

INVx5_ASAP7_75t_L g163 ( 
.A(n_73),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_20),
.B(n_19),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_57),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_75),
.B(n_78),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_39),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g205 ( 
.A(n_76),
.Y(n_205)
);

BUFx3_ASAP7_75t_L g77 ( 
.A(n_55),
.Y(n_77)
);

INVx5_ASAP7_75t_L g170 ( 
.A(n_77),
.Y(n_170)
);

CKINVDCx16_ASAP7_75t_R g78 ( 
.A(n_39),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_46),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g213 ( 
.A(n_79),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_46),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_80),
.B(n_88),
.Y(n_138)
);

BUFx3_ASAP7_75t_L g81 ( 
.A(n_55),
.Y(n_81)
);

INVx4_ASAP7_75t_L g150 ( 
.A(n_81),
.Y(n_150)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_52),
.Y(n_82)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_82),
.Y(n_133)
);

BUFx12f_ASAP7_75t_L g83 ( 
.A(n_44),
.Y(n_83)
);

INVx8_ASAP7_75t_L g135 ( 
.A(n_83),
.Y(n_135)
);

INVx2_ASAP7_75t_SL g84 ( 
.A(n_48),
.Y(n_84)
);

INVx4_ASAP7_75t_L g152 ( 
.A(n_84),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_20),
.B(n_19),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_85),
.B(n_96),
.Y(n_156)
);

BUFx12f_ASAP7_75t_L g86 ( 
.A(n_44),
.Y(n_86)
);

INVx8_ASAP7_75t_L g154 ( 
.A(n_86),
.Y(n_154)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_32),
.Y(n_87)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_87),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_46),
.Y(n_88)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_22),
.Y(n_89)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_89),
.Y(n_167)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_32),
.Y(n_90)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_90),
.Y(n_136)
);

INVx8_ASAP7_75t_L g91 ( 
.A(n_57),
.Y(n_91)
);

INVx3_ASAP7_75t_L g181 ( 
.A(n_91),
.Y(n_181)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_35),
.Y(n_92)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_92),
.Y(n_151)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_22),
.Y(n_93)
);

INVx3_ASAP7_75t_L g143 ( 
.A(n_93),
.Y(n_143)
);

BUFx2_ASAP7_75t_L g94 ( 
.A(n_35),
.Y(n_94)
);

CKINVDCx16_ASAP7_75t_R g221 ( 
.A(n_94),
.Y(n_221)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_46),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g228 ( 
.A(n_95),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_24),
.B(n_0),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_47),
.Y(n_97)
);

INVx6_ASAP7_75t_L g141 ( 
.A(n_97),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_47),
.Y(n_98)
);

INVx6_ASAP7_75t_L g192 ( 
.A(n_98),
.Y(n_192)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_22),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_99),
.B(n_100),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_47),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_47),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_101),
.B(n_108),
.Y(n_176)
);

BUFx24_ASAP7_75t_L g102 ( 
.A(n_48),
.Y(n_102)
);

INVx11_ASAP7_75t_L g175 ( 
.A(n_102),
.Y(n_175)
);

INVx11_ASAP7_75t_L g103 ( 
.A(n_48),
.Y(n_103)
);

INVx4_ASAP7_75t_L g201 ( 
.A(n_103),
.Y(n_201)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_30),
.Y(n_104)
);

INVx6_ASAP7_75t_L g198 ( 
.A(n_104),
.Y(n_198)
);

BUFx4f_ASAP7_75t_SL g105 ( 
.A(n_35),
.Y(n_105)
);

INVx8_ASAP7_75t_L g209 ( 
.A(n_105),
.Y(n_209)
);

INVx8_ASAP7_75t_L g106 ( 
.A(n_48),
.Y(n_106)
);

INVx3_ASAP7_75t_L g207 ( 
.A(n_106),
.Y(n_207)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_30),
.Y(n_107)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_107),
.Y(n_159)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_30),
.Y(n_108)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_25),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_109),
.B(n_112),
.Y(n_177)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_25),
.Y(n_110)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_110),
.Y(n_161)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_25),
.Y(n_111)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_111),
.Y(n_162)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_26),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_26),
.Y(n_113)
);

INVx6_ASAP7_75t_L g219 ( 
.A(n_113),
.Y(n_219)
);

CKINVDCx14_ASAP7_75t_R g114 ( 
.A(n_43),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_114),
.B(n_118),
.Y(n_184)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_26),
.Y(n_115)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_115),
.Y(n_172)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_27),
.Y(n_116)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_116),
.Y(n_187)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_27),
.Y(n_117)
);

INVx3_ASAP7_75t_L g224 ( 
.A(n_117),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_41),
.Y(n_118)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_27),
.Y(n_119)
);

INVx3_ASAP7_75t_L g147 ( 
.A(n_119),
.Y(n_147)
);

INVx8_ASAP7_75t_L g120 ( 
.A(n_31),
.Y(n_120)
);

INVx4_ASAP7_75t_L g214 ( 
.A(n_120),
.Y(n_214)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_34),
.Y(n_121)
);

INVx3_ASAP7_75t_L g149 ( 
.A(n_121),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_24),
.B(n_0),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_122),
.B(n_1),
.Y(n_190)
);

BUFx12f_ASAP7_75t_L g123 ( 
.A(n_31),
.Y(n_123)
);

INVx4_ASAP7_75t_L g218 ( 
.A(n_123),
.Y(n_218)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_34),
.Y(n_124)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_124),
.Y(n_204)
);

BUFx3_ASAP7_75t_L g125 ( 
.A(n_34),
.Y(n_125)
);

INVx3_ASAP7_75t_L g183 ( 
.A(n_125),
.Y(n_183)
);

INVx4_ASAP7_75t_SL g126 ( 
.A(n_43),
.Y(n_126)
);

OR2x2_ASAP7_75t_L g188 ( 
.A(n_126),
.B(n_130),
.Y(n_188)
);

INVx8_ASAP7_75t_L g127 ( 
.A(n_31),
.Y(n_127)
);

INVx3_ASAP7_75t_L g195 ( 
.A(n_127),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_41),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_128),
.B(n_2),
.Y(n_194)
);

INVx5_ASAP7_75t_L g129 ( 
.A(n_21),
.Y(n_129)
);

INVx3_ASAP7_75t_L g211 ( 
.A(n_129),
.Y(n_211)
);

HAxp5_ASAP7_75t_SL g130 ( 
.A(n_43),
.B(n_1),
.CON(n_130),
.SN(n_130)
);

AOI22xp33_ASAP7_75t_L g139 ( 
.A1(n_126),
.A2(n_21),
.B1(n_54),
.B2(n_53),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g232 ( 
.A1(n_139),
.A2(n_148),
.B1(n_155),
.B2(n_164),
.Y(n_232)
);

OAI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_82),
.A2(n_66),
.B1(n_61),
.B2(n_70),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_140),
.A2(n_215),
.B1(n_15),
.B2(n_17),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_60),
.A2(n_29),
.B1(n_36),
.B2(n_38),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_71),
.A2(n_29),
.B1(n_36),
.B2(n_38),
.Y(n_155)
);

AO22x1_ASAP7_75t_SL g158 ( 
.A1(n_93),
.A2(n_43),
.B1(n_54),
.B2(n_53),
.Y(n_158)
);

AO22x1_ASAP7_75t_SL g279 ( 
.A1(n_158),
.A2(n_137),
.B1(n_150),
.B2(n_214),
.Y(n_279)
);

AOI22xp33_ASAP7_75t_L g164 ( 
.A1(n_76),
.A2(n_21),
.B1(n_54),
.B2(n_53),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_129),
.A2(n_28),
.B1(n_33),
.B2(n_40),
.Y(n_165)
);

XNOR2x1_ASAP7_75t_L g292 ( 
.A(n_165),
.B(n_210),
.Y(n_292)
);

AOI22xp33_ASAP7_75t_L g166 ( 
.A1(n_79),
.A2(n_42),
.B1(n_51),
.B2(n_50),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g245 ( 
.A1(n_166),
.A2(n_168),
.B1(n_169),
.B2(n_173),
.Y(n_245)
);

AOI22xp33_ASAP7_75t_L g168 ( 
.A1(n_95),
.A2(n_98),
.B1(n_97),
.B2(n_116),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_94),
.A2(n_28),
.B1(n_33),
.B2(n_40),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_SL g173 ( 
.A1(n_84),
.A2(n_45),
.B1(n_51),
.B2(n_50),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_105),
.B(n_49),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_SL g235 ( 
.A(n_174),
.B(n_186),
.Y(n_235)
);

AOI22xp33_ASAP7_75t_SL g178 ( 
.A1(n_65),
.A2(n_45),
.B1(n_51),
.B2(n_50),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_L g249 ( 
.A1(n_178),
.A2(n_185),
.B1(n_189),
.B2(n_200),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_SL g179 ( 
.A(n_73),
.B(n_49),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g265 ( 
.A(n_179),
.B(n_199),
.Y(n_265)
);

HB1xp67_ASAP7_75t_L g182 ( 
.A(n_119),
.Y(n_182)
);

INVxp67_ASAP7_75t_L g281 ( 
.A(n_182),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_L g185 ( 
.A1(n_68),
.A2(n_45),
.B1(n_42),
.B2(n_56),
.Y(n_185)
);

AND2x2_ASAP7_75t_L g186 ( 
.A(n_121),
.B(n_42),
.Y(n_186)
);

AOI22xp33_ASAP7_75t_L g189 ( 
.A1(n_110),
.A2(n_56),
.B1(n_37),
.B2(n_31),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_SL g260 ( 
.A(n_190),
.B(n_212),
.Y(n_260)
);

AND2x2_ASAP7_75t_SL g193 ( 
.A(n_130),
.B(n_56),
.Y(n_193)
);

NAND2x1_ASAP7_75t_SL g257 ( 
.A(n_193),
.B(n_15),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_194),
.B(n_197),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_105),
.B(n_2),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_SL g199 ( 
.A(n_77),
.B(n_3),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_111),
.A2(n_56),
.B1(n_37),
.B2(n_5),
.Y(n_200)
);

AOI22xp33_ASAP7_75t_L g203 ( 
.A1(n_113),
.A2(n_37),
.B1(n_4),
.B2(n_5),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_203),
.A2(n_225),
.B1(n_227),
.B2(n_102),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_81),
.B(n_37),
.C(n_4),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_206),
.B(n_17),
.C(n_18),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_67),
.A2(n_3),
.B1(n_5),
.B2(n_6),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_125),
.B(n_3),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_L g215 ( 
.A1(n_91),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_117),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_216),
.B(n_223),
.Y(n_253)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_124),
.Y(n_217)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_217),
.Y(n_234)
);

HB1xp67_ASAP7_75t_L g220 ( 
.A(n_123),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_220),
.Y(n_233)
);

AOI22xp33_ASAP7_75t_SL g222 ( 
.A1(n_106),
.A2(n_103),
.B1(n_123),
.B2(n_63),
.Y(n_222)
);

AOI22xp33_ASAP7_75t_SL g246 ( 
.A1(n_222),
.A2(n_86),
.B1(n_58),
.B2(n_59),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_104),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_63),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_225)
);

INVx3_ASAP7_75t_L g226 ( 
.A(n_120),
.Y(n_226)
);

INVx4_ASAP7_75t_SL g295 ( 
.A(n_226),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_83),
.A2(n_7),
.B1(n_10),
.B2(n_11),
.Y(n_227)
);

AND2x2_ASAP7_75t_L g229 ( 
.A(n_188),
.B(n_127),
.Y(n_229)
);

CKINVDCx16_ASAP7_75t_R g350 ( 
.A(n_229),
.Y(n_350)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_152),
.Y(n_230)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_230),
.Y(n_314)
);

INVx5_ASAP7_75t_L g236 ( 
.A(n_209),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g339 ( 
.A1(n_237),
.A2(n_239),
.B1(n_254),
.B2(n_274),
.Y(n_339)
);

AOI22xp33_ASAP7_75t_L g238 ( 
.A1(n_140),
.A2(n_102),
.B1(n_86),
.B2(n_83),
.Y(n_238)
);

OAI22xp33_ASAP7_75t_SL g359 ( 
.A1(n_238),
.A2(n_270),
.B1(n_278),
.B2(n_283),
.Y(n_359)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_168),
.A2(n_188),
.B1(n_164),
.B2(n_193),
.Y(n_239)
);

CKINVDCx16_ASAP7_75t_R g240 ( 
.A(n_184),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_240),
.B(n_264),
.Y(n_333)
);

BUFx6f_ASAP7_75t_L g241 ( 
.A(n_145),
.Y(n_241)
);

INVx3_ASAP7_75t_L g242 ( 
.A(n_218),
.Y(n_242)
);

INVx2_ASAP7_75t_SL g351 ( 
.A(n_242),
.Y(n_351)
);

INVx3_ASAP7_75t_L g243 ( 
.A(n_218),
.Y(n_243)
);

HB1xp67_ASAP7_75t_L g356 ( 
.A(n_243),
.Y(n_356)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_152),
.Y(n_244)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_244),
.Y(n_318)
);

AOI22xp33_ASAP7_75t_SL g317 ( 
.A1(n_246),
.A2(n_272),
.B1(n_275),
.B2(n_294),
.Y(n_317)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_153),
.B(n_12),
.Y(n_247)
);

AND2x2_ASAP7_75t_L g344 ( 
.A(n_247),
.B(n_257),
.Y(n_344)
);

OAI21xp5_ASAP7_75t_L g248 ( 
.A1(n_186),
.A2(n_12),
.B(n_15),
.Y(n_248)
);

OAI21xp5_ASAP7_75t_L g328 ( 
.A1(n_248),
.A2(n_259),
.B(n_269),
.Y(n_328)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_161),
.Y(n_250)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_250),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_177),
.B(n_12),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_251),
.B(n_252),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_158),
.B(n_12),
.Y(n_252)
);

INVx4_ASAP7_75t_L g255 ( 
.A(n_214),
.Y(n_255)
);

AND2x2_ASAP7_75t_L g256 ( 
.A(n_147),
.B(n_15),
.Y(n_256)
);

CKINVDCx14_ASAP7_75t_R g319 ( 
.A(n_256),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_SL g363 ( 
.A(n_258),
.B(n_280),
.Y(n_363)
);

AOI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_156),
.A2(n_172),
.B1(n_162),
.B2(n_187),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_146),
.B(n_17),
.Y(n_261)
);

INVxp67_ASAP7_75t_L g323 ( 
.A(n_261),
.Y(n_323)
);

INVx8_ASAP7_75t_L g262 ( 
.A(n_198),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_204),
.Y(n_263)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_263),
.Y(n_353)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_176),
.Y(n_264)
);

AND2x2_ASAP7_75t_L g266 ( 
.A(n_149),
.B(n_18),
.Y(n_266)
);

INVxp67_ASAP7_75t_L g364 ( 
.A(n_266),
.Y(n_364)
);

INVx5_ASAP7_75t_L g267 ( 
.A(n_209),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_144),
.B(n_18),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_268),
.B(n_276),
.Y(n_330)
);

AOI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_224),
.A2(n_163),
.B1(n_170),
.B2(n_183),
.Y(n_269)
);

AOI22xp33_ASAP7_75t_L g270 ( 
.A1(n_224),
.A2(n_136),
.B1(n_151),
.B2(n_134),
.Y(n_270)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_133),
.Y(n_271)
);

AOI22xp33_ASAP7_75t_SL g272 ( 
.A1(n_175),
.A2(n_202),
.B1(n_207),
.B2(n_142),
.Y(n_272)
);

OR2x2_ASAP7_75t_SL g273 ( 
.A(n_167),
.B(n_150),
.Y(n_273)
);

AOI21xp33_ASAP7_75t_L g347 ( 
.A1(n_273),
.A2(n_297),
.B(n_309),
.Y(n_347)
);

OAI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_203),
.A2(n_166),
.B1(n_139),
.B2(n_189),
.Y(n_274)
);

AOI22xp33_ASAP7_75t_SL g275 ( 
.A1(n_175),
.A2(n_202),
.B1(n_207),
.B2(n_142),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_132),
.B(n_131),
.Y(n_276)
);

BUFx12f_ASAP7_75t_L g277 ( 
.A(n_135),
.Y(n_277)
);

AOI22xp33_ASAP7_75t_L g278 ( 
.A1(n_138),
.A2(n_159),
.B1(n_213),
.B2(n_205),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_279),
.B(n_298),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_143),
.B(n_221),
.Y(n_280)
);

INVx8_ASAP7_75t_L g282 ( 
.A(n_198),
.Y(n_282)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_282),
.Y(n_355)
);

AOI22xp33_ASAP7_75t_L g283 ( 
.A1(n_145),
.A2(n_228),
.B1(n_213),
.B2(n_205),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_219),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g358 ( 
.A(n_284),
.B(n_285),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_SL g285 ( 
.A(n_208),
.B(n_181),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_191),
.B(n_170),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_286),
.B(n_293),
.Y(n_325)
);

OAI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_219),
.A2(n_178),
.B1(n_141),
.B2(n_192),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g341 ( 
.A1(n_287),
.A2(n_307),
.B1(n_274),
.B2(n_237),
.Y(n_341)
);

INVx2_ASAP7_75t_L g288 ( 
.A(n_141),
.Y(n_288)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_288),
.Y(n_361)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_228),
.A2(n_196),
.B1(n_180),
.B2(n_171),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_L g324 ( 
.A1(n_289),
.A2(n_312),
.B1(n_245),
.B2(n_232),
.Y(n_324)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_181),
.Y(n_290)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_290),
.Y(n_362)
);

NOR2xp33_ASAP7_75t_SL g291 ( 
.A(n_195),
.B(n_163),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g367 ( 
.A(n_291),
.B(n_301),
.Y(n_367)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_191),
.B(n_135),
.Y(n_293)
);

AOI22xp33_ASAP7_75t_SL g294 ( 
.A1(n_137),
.A2(n_208),
.B1(n_211),
.B2(n_160),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_154),
.B(n_160),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_296),
.B(n_306),
.Y(n_332)
);

AOI22xp33_ASAP7_75t_SL g297 ( 
.A1(n_201),
.A2(n_154),
.B1(n_173),
.B2(n_222),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_192),
.B(n_157),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_L g299 ( 
.A(n_157),
.B(n_171),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_SL g329 ( 
.A(n_299),
.B(n_302),
.Y(n_329)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_201),
.Y(n_300)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_300),
.Y(n_365)
);

BUFx3_ASAP7_75t_L g301 ( 
.A(n_180),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_SL g302 ( 
.A(n_196),
.B(n_153),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_SL g303 ( 
.A(n_153),
.B(n_184),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_SL g331 ( 
.A(n_303),
.B(n_304),
.Y(n_331)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_152),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_152),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_SL g352 ( 
.A(n_305),
.B(n_308),
.Y(n_352)
);

CKINVDCx16_ASAP7_75t_R g306 ( 
.A(n_220),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_SL g307 ( 
.A1(n_168),
.A2(n_188),
.B1(n_164),
.B2(n_212),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_152),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_SL g309 ( 
.A(n_153),
.B(n_156),
.Y(n_309)
);

O2A1O1Ixp33_ASAP7_75t_SL g310 ( 
.A1(n_188),
.A2(n_193),
.B(n_189),
.C(n_139),
.Y(n_310)
);

O2A1O1Ixp33_ASAP7_75t_L g349 ( 
.A1(n_310),
.A2(n_235),
.B(n_248),
.C(n_279),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_193),
.B(n_177),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_311),
.B(n_257),
.Y(n_338)
);

AOI22xp5_ASAP7_75t_L g312 ( 
.A1(n_140),
.A2(n_188),
.B1(n_212),
.B2(n_215),
.Y(n_312)
);

INVx6_ASAP7_75t_L g313 ( 
.A(n_145),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_313),
.Y(n_320)
);

OAI22xp5_ASAP7_75t_SL g315 ( 
.A1(n_312),
.A2(n_252),
.B1(n_254),
.B2(n_310),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_L g375 ( 
.A1(n_315),
.A2(n_324),
.B1(n_341),
.B2(n_346),
.Y(n_375)
);

AND2x4_ASAP7_75t_L g316 ( 
.A(n_229),
.B(n_239),
.Y(n_316)
);

CKINVDCx16_ASAP7_75t_R g395 ( 
.A(n_316),
.Y(n_395)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_253),
.Y(n_321)
);

CKINVDCx14_ASAP7_75t_R g391 ( 
.A(n_321),
.Y(n_391)
);

CKINVDCx20_ASAP7_75t_R g322 ( 
.A(n_236),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g381 ( 
.A(n_322),
.B(n_336),
.Y(n_381)
);

AOI21xp5_ASAP7_75t_L g334 ( 
.A1(n_229),
.A2(n_310),
.B(n_249),
.Y(n_334)
);

AOI21xp5_ASAP7_75t_L g409 ( 
.A1(n_334),
.A2(n_366),
.B(n_255),
.Y(n_409)
);

CKINVDCx20_ASAP7_75t_R g336 ( 
.A(n_267),
.Y(n_336)
);

AOI32xp33_ASAP7_75t_L g337 ( 
.A1(n_311),
.A2(n_231),
.A3(n_292),
.B1(n_302),
.B2(n_257),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_L g385 ( 
.A(n_337),
.B(n_345),
.Y(n_385)
);

XNOR2xp5_ASAP7_75t_SL g390 ( 
.A(n_338),
.B(n_258),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_268),
.B(n_299),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_340),
.B(n_343),
.Y(n_384)
);

CKINVDCx20_ASAP7_75t_R g342 ( 
.A(n_281),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_L g415 ( 
.A(n_342),
.B(n_354),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_247),
.B(n_260),
.Y(n_343)
);

CKINVDCx20_ASAP7_75t_R g345 ( 
.A(n_281),
.Y(n_345)
);

OAI22xp5_ASAP7_75t_L g346 ( 
.A1(n_235),
.A2(n_307),
.B1(n_259),
.B2(n_298),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_260),
.B(n_256),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_348),
.B(n_244),
.Y(n_402)
);

INVxp67_ASAP7_75t_L g405 ( 
.A(n_349),
.Y(n_405)
);

CKINVDCx20_ASAP7_75t_R g354 ( 
.A(n_291),
.Y(n_354)
);

CKINVDCx20_ASAP7_75t_R g357 ( 
.A(n_256),
.Y(n_357)
);

NOR2xp33_ASAP7_75t_L g393 ( 
.A(n_357),
.B(n_360),
.Y(n_393)
);

NOR2xp33_ASAP7_75t_L g360 ( 
.A(n_264),
.B(n_276),
.Y(n_360)
);

AOI21xp5_ASAP7_75t_L g366 ( 
.A1(n_279),
.A2(n_292),
.B(n_287),
.Y(n_366)
);

AOI32xp33_ASAP7_75t_L g368 ( 
.A1(n_337),
.A2(n_251),
.A3(n_273),
.B1(n_265),
.B2(n_284),
.Y(n_368)
);

NOR2xp33_ASAP7_75t_L g443 ( 
.A(n_368),
.B(n_376),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_SL g369 ( 
.A(n_340),
.B(n_303),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_SL g419 ( 
.A(n_369),
.B(n_400),
.Y(n_419)
);

OAI22xp5_ASAP7_75t_SL g370 ( 
.A1(n_341),
.A2(n_289),
.B1(n_269),
.B2(n_266),
.Y(n_370)
);

AOI22xp5_ASAP7_75t_L g450 ( 
.A1(n_370),
.A2(n_404),
.B1(n_359),
.B2(n_320),
.Y(n_450)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_352),
.Y(n_371)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_371),
.Y(n_432)
);

INVx2_ASAP7_75t_L g372 ( 
.A(n_362),
.Y(n_372)
);

INVxp67_ASAP7_75t_L g430 ( 
.A(n_372),
.Y(n_430)
);

AND2x2_ASAP7_75t_L g373 ( 
.A(n_316),
.B(n_266),
.Y(n_373)
);

AND2x2_ASAP7_75t_L g449 ( 
.A(n_373),
.B(n_379),
.Y(n_449)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_352),
.Y(n_374)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_374),
.Y(n_442)
);

CKINVDCx20_ASAP7_75t_R g376 ( 
.A(n_356),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_327),
.Y(n_377)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_377),
.Y(n_451)
);

OR2x2_ASAP7_75t_L g378 ( 
.A(n_334),
.B(n_230),
.Y(n_378)
);

OAI21xp5_ASAP7_75t_L g420 ( 
.A1(n_378),
.A2(n_349),
.B(n_335),
.Y(n_420)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_327),
.Y(n_379)
);

AND2x2_ASAP7_75t_SL g380 ( 
.A(n_329),
.B(n_316),
.Y(n_380)
);

INVxp67_ASAP7_75t_L g455 ( 
.A(n_380),
.Y(n_455)
);

INVx2_ASAP7_75t_L g382 ( 
.A(n_362),
.Y(n_382)
);

HB1xp67_ASAP7_75t_L g424 ( 
.A(n_382),
.Y(n_424)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_353),
.Y(n_383)
);

HB1xp67_ASAP7_75t_L g447 ( 
.A(n_383),
.Y(n_447)
);

INVx2_ASAP7_75t_L g386 ( 
.A(n_361),
.Y(n_386)
);

AOI22xp33_ASAP7_75t_SL g437 ( 
.A1(n_386),
.A2(n_388),
.B1(n_389),
.B2(n_351),
.Y(n_437)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_353),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_SL g436 ( 
.A(n_387),
.B(n_406),
.Y(n_436)
);

AOI22xp33_ASAP7_75t_SL g388 ( 
.A1(n_316),
.A2(n_295),
.B1(n_304),
.B2(n_308),
.Y(n_388)
);

INVx2_ASAP7_75t_L g389 ( 
.A(n_361),
.Y(n_389)
);

XNOR2xp5_ASAP7_75t_SL g453 ( 
.A(n_390),
.B(n_402),
.Y(n_453)
);

AND2x2_ASAP7_75t_L g392 ( 
.A(n_316),
.B(n_234),
.Y(n_392)
);

CKINVDCx16_ASAP7_75t_R g452 ( 
.A(n_392),
.Y(n_452)
);

XOR2xp5_ASAP7_75t_L g394 ( 
.A(n_329),
.B(n_250),
.Y(n_394)
);

MAJIxp5_ASAP7_75t_L g435 ( 
.A(n_394),
.B(n_398),
.C(n_408),
.Y(n_435)
);

CKINVDCx20_ASAP7_75t_R g396 ( 
.A(n_358),
.Y(n_396)
);

NOR2xp33_ASAP7_75t_L g454 ( 
.A(n_396),
.B(n_407),
.Y(n_454)
);

AND2x2_ASAP7_75t_L g397 ( 
.A(n_350),
.B(n_234),
.Y(n_397)
);

OAI21xp5_ASAP7_75t_SL g421 ( 
.A1(n_397),
.A2(n_399),
.B(n_409),
.Y(n_421)
);

MAJIxp5_ASAP7_75t_L g398 ( 
.A(n_350),
.B(n_233),
.C(n_271),
.Y(n_398)
);

AND2x2_ASAP7_75t_L g399 ( 
.A(n_346),
.B(n_263),
.Y(n_399)
);

FAx1_ASAP7_75t_SL g400 ( 
.A(n_315),
.B(n_233),
.CI(n_305),
.CON(n_400),
.SN(n_400)
);

NAND2xp5_ASAP7_75t_SL g401 ( 
.A(n_330),
.B(n_290),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g418 ( 
.A(n_401),
.B(n_411),
.Y(n_418)
);

AOI22xp5_ASAP7_75t_L g403 ( 
.A1(n_324),
.A2(n_288),
.B1(n_282),
.B2(n_262),
.Y(n_403)
);

OAI22xp5_ASAP7_75t_L g428 ( 
.A1(n_403),
.A2(n_413),
.B1(n_336),
.B2(n_322),
.Y(n_428)
);

OAI22xp33_ASAP7_75t_L g404 ( 
.A1(n_339),
.A2(n_295),
.B1(n_313),
.B2(n_241),
.Y(n_404)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_365),
.Y(n_406)
);

CKINVDCx16_ASAP7_75t_R g407 ( 
.A(n_325),
.Y(n_407)
);

MAJIxp5_ASAP7_75t_L g408 ( 
.A(n_343),
.B(n_242),
.C(n_243),
.Y(n_408)
);

AOI21xp5_ASAP7_75t_L g410 ( 
.A1(n_366),
.A2(n_300),
.B(n_277),
.Y(n_410)
);

AOI21xp5_ASAP7_75t_L g426 ( 
.A1(n_410),
.A2(n_328),
.B(n_317),
.Y(n_426)
);

CKINVDCx20_ASAP7_75t_R g411 ( 
.A(n_358),
.Y(n_411)
);

XOR2xp5_ASAP7_75t_L g412 ( 
.A(n_344),
.B(n_277),
.Y(n_412)
);

MAJIxp5_ASAP7_75t_L g444 ( 
.A(n_412),
.B(n_367),
.C(n_344),
.Y(n_444)
);

AOI22xp5_ASAP7_75t_L g413 ( 
.A1(n_339),
.A2(n_277),
.B1(n_301),
.B2(n_335),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_365),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_414),
.B(n_314),
.Y(n_422)
);

CKINVDCx20_ASAP7_75t_R g416 ( 
.A(n_391),
.Y(n_416)
);

NOR2xp33_ASAP7_75t_L g480 ( 
.A(n_416),
.B(n_417),
.Y(n_480)
);

CKINVDCx20_ASAP7_75t_R g417 ( 
.A(n_381),
.Y(n_417)
);

INVx1_ASAP7_75t_SL g487 ( 
.A(n_420),
.Y(n_487)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_422),
.Y(n_457)
);

OAI22xp5_ASAP7_75t_SL g423 ( 
.A1(n_375),
.A2(n_354),
.B1(n_357),
.B2(n_326),
.Y(n_423)
);

AOI22xp5_ASAP7_75t_L g459 ( 
.A1(n_423),
.A2(n_428),
.B1(n_429),
.B2(n_433),
.Y(n_459)
);

OAI21xp5_ASAP7_75t_L g425 ( 
.A1(n_395),
.A2(n_347),
.B(n_328),
.Y(n_425)
);

OAI21xp5_ASAP7_75t_SL g470 ( 
.A1(n_425),
.A2(n_426),
.B(n_441),
.Y(n_470)
);

AOI22x1_ASAP7_75t_L g427 ( 
.A1(n_405),
.A2(n_399),
.B1(n_370),
.B2(n_409),
.Y(n_427)
);

OAI22xp5_ASAP7_75t_L g486 ( 
.A1(n_427),
.A2(n_397),
.B1(n_406),
.B2(n_414),
.Y(n_486)
);

OAI22xp5_ASAP7_75t_SL g429 ( 
.A1(n_375),
.A2(n_326),
.B1(n_319),
.B2(n_330),
.Y(n_429)
);

XOR2xp5_ASAP7_75t_L g431 ( 
.A(n_384),
.B(n_363),
.Y(n_431)
);

MAJIxp5_ASAP7_75t_L g467 ( 
.A(n_431),
.B(n_444),
.C(n_445),
.Y(n_467)
);

OAI22xp5_ASAP7_75t_SL g433 ( 
.A1(n_378),
.A2(n_331),
.B1(n_348),
.B2(n_364),
.Y(n_433)
);

INVx5_ASAP7_75t_L g434 ( 
.A(n_376),
.Y(n_434)
);

INVx2_ASAP7_75t_L g461 ( 
.A(n_434),
.Y(n_461)
);

INVxp67_ASAP7_75t_L g460 ( 
.A(n_437),
.Y(n_460)
);

INVx5_ASAP7_75t_L g438 ( 
.A(n_413),
.Y(n_438)
);

NOR2xp33_ASAP7_75t_L g482 ( 
.A(n_438),
.B(n_345),
.Y(n_482)
);

AOI21xp5_ASAP7_75t_L g439 ( 
.A1(n_405),
.A2(n_367),
.B(n_332),
.Y(n_439)
);

AOI21xp5_ASAP7_75t_L g488 ( 
.A1(n_439),
.A2(n_333),
.B(n_377),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_396),
.B(n_331),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_440),
.B(n_446),
.Y(n_471)
);

AOI22xp5_ASAP7_75t_SL g441 ( 
.A1(n_411),
.A2(n_415),
.B1(n_399),
.B2(n_395),
.Y(n_441)
);

XOR2xp5_ASAP7_75t_L g445 ( 
.A(n_384),
.B(n_363),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_L g446 ( 
.A(n_401),
.B(n_344),
.Y(n_446)
);

OAI32xp33_ASAP7_75t_L g448 ( 
.A1(n_385),
.A2(n_333),
.A3(n_338),
.B1(n_323),
.B2(n_314),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_L g477 ( 
.A(n_448),
.B(n_450),
.Y(n_477)
);

AOI22xp5_ASAP7_75t_L g456 ( 
.A1(n_403),
.A2(n_320),
.B1(n_321),
.B2(n_355),
.Y(n_456)
);

OAI22xp5_ASAP7_75t_SL g465 ( 
.A1(n_456),
.A2(n_371),
.B1(n_378),
.B2(n_392),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_SL g458 ( 
.A(n_440),
.B(n_374),
.Y(n_458)
);

CKINVDCx14_ASAP7_75t_R g504 ( 
.A(n_458),
.Y(n_504)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_422),
.Y(n_462)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_462),
.Y(n_497)
);

NOR2xp33_ASAP7_75t_SL g463 ( 
.A(n_454),
.B(n_393),
.Y(n_463)
);

NOR2xp33_ASAP7_75t_SL g518 ( 
.A(n_463),
.B(n_473),
.Y(n_518)
);

INVxp67_ASAP7_75t_L g464 ( 
.A(n_449),
.Y(n_464)
);

NOR2xp33_ASAP7_75t_L g496 ( 
.A(n_464),
.B(n_466),
.Y(n_496)
);

AOI22xp5_ASAP7_75t_L g524 ( 
.A1(n_465),
.A2(n_469),
.B1(n_474),
.B2(n_452),
.Y(n_524)
);

CKINVDCx14_ASAP7_75t_R g466 ( 
.A(n_418),
.Y(n_466)
);

OR2x2_ASAP7_75t_L g468 ( 
.A(n_420),
.B(n_400),
.Y(n_468)
);

CKINVDCx20_ASAP7_75t_R g499 ( 
.A(n_468),
.Y(n_499)
);

OAI22xp5_ASAP7_75t_SL g469 ( 
.A1(n_441),
.A2(n_410),
.B1(n_380),
.B2(n_373),
.Y(n_469)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_436),
.Y(n_472)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_472),
.Y(n_498)
);

NOR2xp33_ASAP7_75t_SL g473 ( 
.A(n_416),
.B(n_369),
.Y(n_473)
);

OAI22xp5_ASAP7_75t_SL g474 ( 
.A1(n_426),
.A2(n_380),
.B1(n_373),
.B2(n_400),
.Y(n_474)
);

AOI22xp5_ASAP7_75t_SL g475 ( 
.A1(n_433),
.A2(n_392),
.B1(n_407),
.B2(n_368),
.Y(n_475)
);

OAI21xp5_ASAP7_75t_SL g503 ( 
.A1(n_475),
.A2(n_483),
.B(n_485),
.Y(n_503)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_436),
.Y(n_476)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_476),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_L g478 ( 
.A(n_418),
.B(n_402),
.Y(n_478)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_478),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_L g479 ( 
.A(n_432),
.B(n_408),
.Y(n_479)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_479),
.Y(n_507)
);

CKINVDCx20_ASAP7_75t_R g481 ( 
.A(n_447),
.Y(n_481)
);

NOR2xp33_ASAP7_75t_L g523 ( 
.A(n_481),
.B(n_491),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_L g495 ( 
.A(n_482),
.B(n_494),
.Y(n_495)
);

OAI21xp5_ASAP7_75t_L g483 ( 
.A1(n_425),
.A2(n_421),
.B(n_455),
.Y(n_483)
);

MAJIxp5_ASAP7_75t_L g484 ( 
.A(n_435),
.B(n_394),
.C(n_412),
.Y(n_484)
);

MAJIxp5_ASAP7_75t_L g513 ( 
.A(n_484),
.B(n_490),
.C(n_453),
.Y(n_513)
);

OAI21xp5_ASAP7_75t_L g485 ( 
.A1(n_421),
.A2(n_398),
.B(n_397),
.Y(n_485)
);

OA21x2_ASAP7_75t_L g502 ( 
.A1(n_486),
.A2(n_428),
.B(n_450),
.Y(n_502)
);

HB1xp67_ASAP7_75t_L g517 ( 
.A(n_488),
.Y(n_517)
);

XNOR2xp5_ASAP7_75t_L g489 ( 
.A(n_431),
.B(n_390),
.Y(n_489)
);

XOR2xp5_ASAP7_75t_L g508 ( 
.A(n_489),
.B(n_493),
.Y(n_508)
);

XOR2xp5_ASAP7_75t_L g490 ( 
.A(n_445),
.B(n_387),
.Y(n_490)
);

CKINVDCx16_ASAP7_75t_R g491 ( 
.A(n_424),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_451),
.Y(n_492)
);

XNOR2xp5_ASAP7_75t_L g493 ( 
.A(n_453),
.B(n_383),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_451),
.Y(n_494)
);

OAI22xp5_ASAP7_75t_SL g500 ( 
.A1(n_459),
.A2(n_477),
.B1(n_475),
.B2(n_487),
.Y(n_500)
);

AOI22xp5_ASAP7_75t_L g532 ( 
.A1(n_500),
.A2(n_511),
.B1(n_527),
.B2(n_486),
.Y(n_532)
);

OAI22xp5_ASAP7_75t_L g548 ( 
.A1(n_502),
.A2(n_519),
.B1(n_494),
.B2(n_372),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_L g505 ( 
.A(n_480),
.B(n_442),
.Y(n_505)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_505),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_L g509 ( 
.A(n_480),
.B(n_442),
.Y(n_509)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_509),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_L g510 ( 
.A(n_472),
.B(n_432),
.Y(n_510)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_510),
.Y(n_547)
);

OAI22xp5_ASAP7_75t_SL g511 ( 
.A1(n_459),
.A2(n_443),
.B1(n_438),
.B2(n_455),
.Y(n_511)
);

XOR2xp5_ASAP7_75t_L g512 ( 
.A(n_467),
.B(n_489),
.Y(n_512)
);

XOR2xp5_ASAP7_75t_L g529 ( 
.A(n_512),
.B(n_513),
.Y(n_529)
);

AOI21xp5_ASAP7_75t_L g514 ( 
.A1(n_470),
.A2(n_427),
.B(n_439),
.Y(n_514)
);

AOI21xp5_ASAP7_75t_L g556 ( 
.A1(n_514),
.A2(n_521),
.B(n_522),
.Y(n_556)
);

CKINVDCx20_ASAP7_75t_R g515 ( 
.A(n_463),
.Y(n_515)
);

AOI22xp33_ASAP7_75t_L g538 ( 
.A1(n_515),
.A2(n_462),
.B1(n_471),
.B2(n_478),
.Y(n_538)
);

XOR2x1_ASAP7_75t_L g516 ( 
.A(n_474),
.B(n_427),
.Y(n_516)
);

XNOR2x1_ASAP7_75t_L g550 ( 
.A(n_516),
.B(n_524),
.Y(n_550)
);

OAI22xp5_ASAP7_75t_L g519 ( 
.A1(n_457),
.A2(n_456),
.B1(n_419),
.B2(n_417),
.Y(n_519)
);

MAJIxp5_ASAP7_75t_L g520 ( 
.A(n_484),
.B(n_435),
.C(n_444),
.Y(n_520)
);

MAJIxp5_ASAP7_75t_L g536 ( 
.A(n_520),
.B(n_528),
.C(n_479),
.Y(n_536)
);

AOI211xp5_ASAP7_75t_SL g521 ( 
.A1(n_468),
.A2(n_419),
.B(n_448),
.C(n_423),
.Y(n_521)
);

AOI21xp5_ASAP7_75t_L g522 ( 
.A1(n_470),
.A2(n_449),
.B(n_429),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_476),
.B(n_434),
.Y(n_525)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_525),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_L g526 ( 
.A(n_458),
.B(n_430),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_L g540 ( 
.A(n_526),
.B(n_481),
.Y(n_540)
);

OAI22xp5_ASAP7_75t_SL g527 ( 
.A1(n_477),
.A2(n_452),
.B1(n_446),
.B2(n_449),
.Y(n_527)
);

MAJIxp5_ASAP7_75t_L g528 ( 
.A(n_467),
.B(n_379),
.C(n_430),
.Y(n_528)
);

XNOR2xp5_ASAP7_75t_L g530 ( 
.A(n_528),
.B(n_490),
.Y(n_530)
);

XOR2xp5_ASAP7_75t_L g559 ( 
.A(n_530),
.B(n_533),
.Y(n_559)
);

OAI22xp5_ASAP7_75t_L g567 ( 
.A1(n_532),
.A2(n_538),
.B1(n_543),
.B2(n_502),
.Y(n_567)
);

XNOR2xp5_ASAP7_75t_L g533 ( 
.A(n_512),
.B(n_493),
.Y(n_533)
);

XNOR2xp5_ASAP7_75t_SL g534 ( 
.A(n_508),
.B(n_487),
.Y(n_534)
);

XOR2xp5_ASAP7_75t_L g573 ( 
.A(n_534),
.B(n_537),
.Y(n_573)
);

OAI22xp5_ASAP7_75t_SL g535 ( 
.A1(n_524),
.A2(n_468),
.B1(n_471),
.B2(n_457),
.Y(n_535)
);

AOI22xp5_ASAP7_75t_L g562 ( 
.A1(n_535),
.A2(n_548),
.B1(n_502),
.B2(n_501),
.Y(n_562)
);

MAJIxp5_ASAP7_75t_L g561 ( 
.A(n_536),
.B(n_544),
.C(n_545),
.Y(n_561)
);

XOR2xp5_ASAP7_75t_L g537 ( 
.A(n_513),
.B(n_483),
.Y(n_537)
);

XOR2x2_ASAP7_75t_SL g539 ( 
.A(n_527),
.B(n_469),
.Y(n_539)
);

FAx1_ASAP7_75t_SL g564 ( 
.A(n_539),
.B(n_511),
.CI(n_516),
.CON(n_564),
.SN(n_564)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_540),
.Y(n_568)
);

XNOR2xp5_ASAP7_75t_SL g542 ( 
.A(n_508),
.B(n_485),
.Y(n_542)
);

AOI22xp5_ASAP7_75t_L g543 ( 
.A1(n_502),
.A2(n_465),
.B1(n_460),
.B2(n_488),
.Y(n_543)
);

MAJIxp5_ASAP7_75t_L g544 ( 
.A(n_520),
.B(n_491),
.C(n_461),
.Y(n_544)
);

MAJIxp5_ASAP7_75t_L g545 ( 
.A(n_507),
.B(n_461),
.C(n_492),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_L g546 ( 
.A(n_515),
.B(n_473),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_SL g565 ( 
.A(n_546),
.B(n_552),
.Y(n_565)
);

XNOR2xp5_ASAP7_75t_L g549 ( 
.A(n_507),
.B(n_382),
.Y(n_549)
);

HB1xp67_ASAP7_75t_L g570 ( 
.A(n_549),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_L g552 ( 
.A(n_523),
.B(n_342),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_SL g553 ( 
.A(n_518),
.B(n_318),
.Y(n_553)
);

NOR2xp33_ASAP7_75t_SL g563 ( 
.A(n_553),
.B(n_557),
.Y(n_563)
);

XOR2xp5_ASAP7_75t_L g554 ( 
.A(n_503),
.B(n_389),
.Y(n_554)
);

MAJIxp5_ASAP7_75t_L g578 ( 
.A(n_554),
.B(n_517),
.C(n_516),
.Y(n_578)
);

INVx2_ASAP7_75t_SL g555 ( 
.A(n_525),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_L g558 ( 
.A(n_555),
.B(n_526),
.Y(n_558)
);

NOR2xp33_ASAP7_75t_L g557 ( 
.A(n_518),
.B(n_318),
.Y(n_557)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_558),
.Y(n_586)
);

NOR2xp33_ASAP7_75t_L g560 ( 
.A(n_544),
.B(n_500),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_L g594 ( 
.A(n_560),
.B(n_564),
.Y(n_594)
);

AOI22xp5_ASAP7_75t_L g581 ( 
.A1(n_562),
.A2(n_567),
.B1(n_569),
.B2(n_574),
.Y(n_581)
);

BUFx2_ASAP7_75t_L g566 ( 
.A(n_531),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_L g595 ( 
.A(n_566),
.B(n_571),
.Y(n_595)
);

OAI321xp33_ASAP7_75t_L g569 ( 
.A1(n_556),
.A2(n_499),
.A3(n_514),
.B1(n_521),
.B2(n_522),
.C(n_506),
.Y(n_569)
);

CKINVDCx20_ASAP7_75t_R g571 ( 
.A(n_555),
.Y(n_571)
);

NOR2xp33_ASAP7_75t_L g572 ( 
.A(n_536),
.B(n_519),
.Y(n_572)
);

XNOR2xp5_ASAP7_75t_L g596 ( 
.A(n_572),
.B(n_575),
.Y(n_596)
);

OAI22xp5_ASAP7_75t_L g574 ( 
.A1(n_532),
.A2(n_504),
.B1(n_543),
.B2(n_547),
.Y(n_574)
);

NOR2xp33_ASAP7_75t_L g575 ( 
.A(n_545),
.B(n_506),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_L g576 ( 
.A(n_549),
.B(n_523),
.Y(n_576)
);

OAI21xp5_ASAP7_75t_L g597 ( 
.A1(n_576),
.A2(n_495),
.B(n_505),
.Y(n_597)
);

CKINVDCx20_ASAP7_75t_R g577 ( 
.A(n_556),
.Y(n_577)
);

NOR2xp33_ASAP7_75t_L g585 ( 
.A(n_577),
.B(n_579),
.Y(n_585)
);

XOR2xp5_ASAP7_75t_L g580 ( 
.A(n_578),
.B(n_539),
.Y(n_580)
);

INVxp67_ASAP7_75t_L g579 ( 
.A(n_554),
.Y(n_579)
);

XNOR2xp5_ASAP7_75t_L g601 ( 
.A(n_580),
.B(n_582),
.Y(n_601)
);

XOR2xp5_ASAP7_75t_L g582 ( 
.A(n_573),
.B(n_533),
.Y(n_582)
);

MAJIxp5_ASAP7_75t_L g583 ( 
.A(n_561),
.B(n_529),
.C(n_530),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_L g599 ( 
.A(n_583),
.B(n_584),
.Y(n_599)
);

NAND2x1p5_ASAP7_75t_L g584 ( 
.A(n_558),
.B(n_535),
.Y(n_584)
);

XOR2xp5_ASAP7_75t_L g587 ( 
.A(n_573),
.B(n_537),
.Y(n_587)
);

XNOR2xp5_ASAP7_75t_L g613 ( 
.A(n_587),
.B(n_588),
.Y(n_613)
);

XOR2xp5_ASAP7_75t_L g588 ( 
.A(n_559),
.B(n_529),
.Y(n_588)
);

MAJIxp5_ASAP7_75t_L g589 ( 
.A(n_561),
.B(n_542),
.C(n_550),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_L g602 ( 
.A(n_589),
.B(n_591),
.Y(n_602)
);

BUFx24_ASAP7_75t_SL g590 ( 
.A(n_565),
.Y(n_590)
);

NOR2xp33_ASAP7_75t_SL g612 ( 
.A(n_590),
.B(n_598),
.Y(n_612)
);

MAJIxp5_ASAP7_75t_L g591 ( 
.A(n_559),
.B(n_550),
.C(n_534),
.Y(n_591)
);

XNOR2xp5_ASAP7_75t_L g592 ( 
.A(n_578),
.B(n_503),
.Y(n_592)
);

HB1xp67_ASAP7_75t_L g610 ( 
.A(n_592),
.Y(n_610)
);

AOI22xp5_ASAP7_75t_L g593 ( 
.A1(n_568),
.A2(n_541),
.B1(n_551),
.B2(n_495),
.Y(n_593)
);

HB1xp67_ASAP7_75t_L g614 ( 
.A(n_593),
.Y(n_614)
);

XOR2xp5_ASAP7_75t_L g607 ( 
.A(n_597),
.B(n_576),
.Y(n_607)
);

FAx1_ASAP7_75t_SL g598 ( 
.A(n_569),
.B(n_499),
.CI(n_496),
.CON(n_598),
.SN(n_598)
);

NOR2xp33_ASAP7_75t_L g600 ( 
.A(n_596),
.B(n_563),
.Y(n_600)
);

OR2x2_ASAP7_75t_L g616 ( 
.A(n_600),
.B(n_606),
.Y(n_616)
);

AOI21xp5_ASAP7_75t_SL g603 ( 
.A1(n_585),
.A2(n_568),
.B(n_496),
.Y(n_603)
);

AOI21xp5_ASAP7_75t_L g623 ( 
.A1(n_603),
.A2(n_510),
.B(n_498),
.Y(n_623)
);

CKINVDCx20_ASAP7_75t_R g604 ( 
.A(n_595),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_L g621 ( 
.A(n_604),
.B(n_605),
.Y(n_621)
);

OAI22xp5_ASAP7_75t_SL g605 ( 
.A1(n_581),
.A2(n_562),
.B1(n_577),
.B2(n_571),
.Y(n_605)
);

NOR2xp33_ASAP7_75t_L g606 ( 
.A(n_594),
.B(n_563),
.Y(n_606)
);

AND2x2_ASAP7_75t_L g615 ( 
.A(n_607),
.B(n_584),
.Y(n_615)
);

NOR2xp33_ASAP7_75t_L g608 ( 
.A(n_583),
.B(n_566),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_L g625 ( 
.A(n_608),
.B(n_609),
.Y(n_625)
);

OAI22xp5_ASAP7_75t_SL g609 ( 
.A1(n_598),
.A2(n_564),
.B1(n_497),
.B2(n_579),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_SL g611 ( 
.A(n_589),
.B(n_509),
.Y(n_611)
);

NOR2xp33_ASAP7_75t_SL g619 ( 
.A(n_611),
.B(n_592),
.Y(n_619)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_615),
.Y(n_627)
);

NOR2xp33_ASAP7_75t_L g617 ( 
.A(n_612),
.B(n_586),
.Y(n_617)
);

NOR2xp33_ASAP7_75t_SL g631 ( 
.A(n_617),
.B(n_618),
.Y(n_631)
);

MAJIxp5_ASAP7_75t_L g618 ( 
.A(n_602),
.B(n_588),
.C(n_580),
.Y(n_618)
);

NOR2xp33_ASAP7_75t_L g626 ( 
.A(n_619),
.B(n_601),
.Y(n_626)
);

NOR2xp33_ASAP7_75t_L g620 ( 
.A(n_614),
.B(n_501),
.Y(n_620)
);

AND2x2_ASAP7_75t_L g629 ( 
.A(n_620),
.B(n_623),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_SL g622 ( 
.A(n_599),
.B(n_498),
.Y(n_622)
);

XNOR2xp5_ASAP7_75t_L g632 ( 
.A(n_622),
.B(n_624),
.Y(n_632)
);

MAJIxp5_ASAP7_75t_L g624 ( 
.A(n_610),
.B(n_570),
.C(n_582),
.Y(n_624)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_626),
.Y(n_636)
);

NOR2xp33_ASAP7_75t_L g628 ( 
.A(n_616),
.B(n_609),
.Y(n_628)
);

AOI21xp5_ASAP7_75t_L g638 ( 
.A1(n_628),
.A2(n_630),
.B(n_613),
.Y(n_638)
);

MAJIxp5_ASAP7_75t_L g630 ( 
.A(n_625),
.B(n_601),
.C(n_613),
.Y(n_630)
);

XNOR2xp5_ASAP7_75t_L g633 ( 
.A(n_615),
.B(n_607),
.Y(n_633)
);

MAJIxp5_ASAP7_75t_L g635 ( 
.A(n_633),
.B(n_621),
.C(n_603),
.Y(n_635)
);

INVxp67_ASAP7_75t_L g634 ( 
.A(n_630),
.Y(n_634)
);

OAI21xp5_ASAP7_75t_L g639 ( 
.A1(n_634),
.A2(n_635),
.B(n_638),
.Y(n_639)
);

OAI22xp5_ASAP7_75t_L g637 ( 
.A1(n_627),
.A2(n_617),
.B1(n_620),
.B2(n_497),
.Y(n_637)
);

NAND2xp33_ASAP7_75t_L g640 ( 
.A(n_637),
.B(n_632),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_L g641 ( 
.A(n_640),
.B(n_636),
.Y(n_641)
);

OAI21xp5_ASAP7_75t_L g642 ( 
.A1(n_641),
.A2(n_639),
.B(n_631),
.Y(n_642)
);

AOI31xp33_ASAP7_75t_SL g643 ( 
.A1(n_642),
.A2(n_629),
.A3(n_633),
.B(n_591),
.Y(n_643)
);

OAI311xp33_ASAP7_75t_L g644 ( 
.A1(n_643),
.A2(n_629),
.A3(n_605),
.B1(n_564),
.C1(n_587),
.Y(n_644)
);


endmodule