module real_aes_6025_n_77 (n_17, n_28, n_76, n_56, n_34, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_43, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_44, n_7, n_4, n_6, n_12, n_68, n_69, n_46, n_59, n_25, n_73, n_48, n_37, n_70, n_50, n_26, n_13, n_24, n_2, n_55, n_62, n_67, n_33, n_14, n_11, n_16, n_39, n_5, n_45, n_60, n_38, n_0, n_63, n_1, n_53, n_36, n_77);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_43;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_44;
input n_7;
input n_4;
input n_6;
input n_12;
input n_68;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_48;
input n_37;
input n_70;
input n_50;
input n_26;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_67;
input n_33;
input n_14;
input n_11;
input n_16;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_0;
input n_63;
input n_1;
input n_53;
input n_36;
output n_77;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_90;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_503;
wire n_635;
wire n_287;
wire n_357;
wire n_386;
wire n_518;
wire n_254;
wire n_207;
wire n_580;
wire n_577;
wire n_469;
wire n_83;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_322;
wire n_328;
wire n_318;
wire n_355;
wire n_239;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_364;
wire n_319;
wire n_555;
wire n_421;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_571;
wire n_376;
wire n_549;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_551;
wire n_320;
wire n_560;
wire n_260;
wire n_594;
wire n_97;
wire n_186;
wire n_138;
wire n_379;
wire n_374;
wire n_453;
wire n_235;
wire n_399;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_92;
wire n_519;
wire n_564;
wire n_573;
wire n_510;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_94;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_578;
wire n_528;
wire n_202;
wire n_495;
wire n_370;
wire n_98;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_82;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_517;
wire n_174;
wire n_570;
wire n_530;
wire n_104;
wire n_535;
wire n_211;
wire n_281;
wire n_496;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_178;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_297;
wire n_383;
wire n_529;
wire n_455;
wire n_119;
wire n_310;
wire n_504;
wire n_164;
wire n_231;
wire n_547;
wire n_102;
wire n_634;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_80;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_367;
wire n_267;
wire n_218;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_339;
wire n_398;
wire n_89;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_93;
wire n_182;
wire n_449;
wire n_417;
wire n_363;
wire n_607;
wire n_323;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_600;
wire n_250;
wire n_605;
wire n_85;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_87;
wire n_171;
wire n_78;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_557;
wire n_488;
wire n_501;
wire n_251;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_96;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_95;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_533;
wire n_366;
wire n_346;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_622;
wire n_470;
wire n_81;
wire n_133;
wire n_494;
wire n_377;
wire n_273;
wire n_114;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_486;
wire n_411;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_88;
wire n_159;
wire n_108;
wire n_373;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_526;
wire n_155;
wire n_243;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_633;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_249;
wire n_623;
wire n_446;
wire n_221;
wire n_156;
wire n_359;
wire n_456;
wire n_312;
wire n_183;
wire n_266;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_524;
wire n_219;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_371;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_99;
wire n_440;
wire n_525;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_79;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_566;
wire n_474;
wire n_170;
wire n_86;
wire n_375;
wire n_597;
wire n_340;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_241;
wire n_175;
wire n_105;
wire n_84;
wire n_393;
wire n_294;
wire n_258;
wire n_206;
wire n_307;
wire n_500;
wire n_601;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_554;
wire n_475;
wire n_264;
wire n_237;
wire n_91;
INVx1_ASAP7_75t_L g266 ( .A(n_0), .Y(n_266) );
AOI22xp5_ASAP7_75t_L g237 ( .A1(n_1), .A2(n_14), .B1(n_84), .B2(n_217), .Y(n_237) );
AOI22xp33_ASAP7_75t_L g590 ( .A1(n_2), .A2(n_37), .B1(n_591), .B2(n_592), .Y(n_590) );
INVx2_ASAP7_75t_L g127 ( .A(n_3), .Y(n_127) );
INVx1_ASAP7_75t_SL g186 ( .A(n_4), .Y(n_186) );
HB1xp67_ASAP7_75t_L g597 ( .A(n_5), .Y(n_597) );
NAND2xp5_ASAP7_75t_L g256 ( .A(n_6), .B(n_257), .Y(n_256) );
NAND2xp5_ASAP7_75t_L g168 ( .A(n_7), .B(n_169), .Y(n_168) );
INVx1_ASAP7_75t_L g529 ( .A(n_8), .Y(n_529) );
NOR2xp33_ASAP7_75t_L g565 ( .A(n_8), .B(n_59), .Y(n_565) );
INVxp67_ASAP7_75t_L g578 ( .A(n_8), .Y(n_578) );
AOI22xp33_ASAP7_75t_L g162 ( .A1(n_9), .A2(n_46), .B1(n_163), .B2(n_164), .Y(n_162) );
INVx1_ASAP7_75t_L g636 ( .A(n_9), .Y(n_636) );
AOI221xp5_ASAP7_75t_L g553 ( .A1(n_10), .A2(n_25), .B1(n_554), .B2(n_555), .C(n_557), .Y(n_553) );
OAI22xp33_ASAP7_75t_SL g628 ( .A1(n_11), .A2(n_502), .B1(n_503), .B2(n_629), .Y(n_628) );
CKINVDCx5p33_ASAP7_75t_R g629 ( .A(n_11), .Y(n_629) );
OA21x2_ASAP7_75t_L g108 ( .A1(n_12), .A2(n_57), .B(n_109), .Y(n_108) );
OA21x2_ASAP7_75t_L g157 ( .A1(n_12), .A2(n_57), .B(n_109), .Y(n_157) );
NAND2xp5_ASAP7_75t_SL g525 ( .A(n_13), .B(n_514), .Y(n_525) );
NOR2xp33_ASAP7_75t_L g227 ( .A(n_15), .B(n_123), .Y(n_227) );
AOI22xp5_ASAP7_75t_L g111 ( .A1(n_16), .A2(n_63), .B1(n_112), .B2(n_115), .Y(n_111) );
INVx2_ASAP7_75t_L g221 ( .A(n_17), .Y(n_221) );
AOI22xp33_ASAP7_75t_L g506 ( .A1(n_18), .A2(n_55), .B1(n_507), .B2(n_532), .Y(n_506) );
AOI22xp5_ASAP7_75t_L g238 ( .A1(n_19), .A2(n_24), .B1(n_147), .B2(n_185), .Y(n_238) );
BUFx3_ASAP7_75t_L g610 ( .A(n_20), .Y(n_610) );
O2A1O1Ixp5_ASAP7_75t_L g214 ( .A1(n_21), .A2(n_88), .B(n_215), .C(n_216), .Y(n_214) );
AOI22xp33_ASAP7_75t_L g119 ( .A1(n_22), .A2(n_51), .B1(n_120), .B2(n_122), .Y(n_119) );
HB1xp67_ASAP7_75t_L g501 ( .A(n_23), .Y(n_501) );
CKINVDCx5p33_ASAP7_75t_R g149 ( .A(n_26), .Y(n_149) );
AOI22xp5_ASAP7_75t_L g583 ( .A1(n_27), .A2(n_50), .B1(n_584), .B2(n_588), .Y(n_583) );
BUFx6f_ASAP7_75t_L g514 ( .A(n_28), .Y(n_514) );
AOI22xp33_ASAP7_75t_L g579 ( .A1(n_29), .A2(n_56), .B1(n_580), .B2(n_581), .Y(n_579) );
AOI22xp33_ASAP7_75t_L g570 ( .A1(n_30), .A2(n_54), .B1(n_571), .B2(n_572), .Y(n_570) );
AOI22xp5_ASAP7_75t_L g536 ( .A1(n_31), .A2(n_74), .B1(n_537), .B2(n_542), .Y(n_536) );
AOI22xp5_ASAP7_75t_L g171 ( .A1(n_32), .A2(n_65), .B1(n_172), .B2(n_174), .Y(n_171) );
INVx1_ASAP7_75t_L g210 ( .A(n_33), .Y(n_210) );
INVx1_ASAP7_75t_L g515 ( .A(n_34), .Y(n_515) );
NAND2xp5_ASAP7_75t_L g575 ( .A(n_34), .B(n_58), .Y(n_575) );
HB1xp67_ASAP7_75t_L g600 ( .A(n_35), .Y(n_600) );
INVx1_ASAP7_75t_L g558 ( .A(n_36), .Y(n_558) );
NAND2xp5_ASAP7_75t_L g261 ( .A(n_38), .B(n_206), .Y(n_261) );
INVx2_ASAP7_75t_L g218 ( .A(n_39), .Y(n_218) );
CKINVDCx5p33_ASAP7_75t_R g151 ( .A(n_40), .Y(n_151) );
INVx2_ASAP7_75t_L g226 ( .A(n_41), .Y(n_226) );
NAND2xp5_ASAP7_75t_L g258 ( .A(n_42), .B(n_259), .Y(n_258) );
INVx1_ASAP7_75t_SL g190 ( .A(n_43), .Y(n_190) );
INVx1_ASAP7_75t_L g143 ( .A(n_44), .Y(n_143) );
HB1xp67_ASAP7_75t_L g601 ( .A(n_44), .Y(n_601) );
INVx1_ASAP7_75t_L g109 ( .A(n_45), .Y(n_109) );
AND2x4_ASAP7_75t_L g91 ( .A(n_47), .B(n_92), .Y(n_91) );
AND2x4_ASAP7_75t_L g138 ( .A(n_47), .B(n_92), .Y(n_138) );
HB1xp67_ASAP7_75t_L g620 ( .A(n_47), .Y(n_620) );
INVx1_ASAP7_75t_L g195 ( .A(n_48), .Y(n_195) );
BUFx6f_ASAP7_75t_L g89 ( .A(n_49), .Y(n_89) );
NOR2xp33_ASAP7_75t_L g230 ( .A(n_52), .B(n_188), .Y(n_230) );
OA22x2_ASAP7_75t_L g520 ( .A1(n_53), .A2(n_59), .B1(n_514), .B2(n_518), .Y(n_520) );
INVx1_ASAP7_75t_L g549 ( .A(n_53), .Y(n_549) );
INVx1_ASAP7_75t_L g531 ( .A(n_58), .Y(n_531) );
NAND2xp5_ASAP7_75t_L g568 ( .A(n_58), .B(n_547), .Y(n_568) );
HB1xp67_ASAP7_75t_L g613 ( .A(n_58), .Y(n_613) );
OAI21xp33_ASAP7_75t_L g550 ( .A1(n_59), .A2(n_64), .B(n_551), .Y(n_550) );
CKINVDCx5p33_ASAP7_75t_R g134 ( .A(n_60), .Y(n_134) );
CKINVDCx5p33_ASAP7_75t_R g208 ( .A(n_61), .Y(n_208) );
NOR2xp33_ASAP7_75t_L g192 ( .A(n_62), .B(n_116), .Y(n_192) );
INVx1_ASAP7_75t_L g517 ( .A(n_64), .Y(n_517) );
NOR2xp33_ASAP7_75t_L g566 ( .A(n_64), .B(n_75), .Y(n_566) );
INVx1_ASAP7_75t_L g624 ( .A(n_65), .Y(n_624) );
HB1xp67_ASAP7_75t_L g595 ( .A(n_66), .Y(n_595) );
BUFx6f_ASAP7_75t_L g85 ( .A(n_67), .Y(n_85) );
INVx1_ASAP7_75t_L g114 ( .A(n_67), .Y(n_114) );
BUFx5_ASAP7_75t_L g148 ( .A(n_67), .Y(n_148) );
NOR2xp33_ASAP7_75t_L g187 ( .A(n_68), .B(n_188), .Y(n_187) );
INVx2_ASAP7_75t_L g229 ( .A(n_69), .Y(n_229) );
INVx1_ASAP7_75t_L g233 ( .A(n_70), .Y(n_233) );
INVx2_ASAP7_75t_L g155 ( .A(n_71), .Y(n_155) );
INVx2_ASAP7_75t_SL g92 ( .A(n_72), .Y(n_92) );
NAND2xp5_ASAP7_75t_SL g252 ( .A(n_73), .B(n_253), .Y(n_252) );
NAND2xp5_ASAP7_75t_L g523 ( .A(n_75), .B(n_524), .Y(n_523) );
AO32x2_ASAP7_75t_L g235 ( .A1(n_76), .A2(n_90), .A3(n_219), .B1(n_236), .B2(n_240), .Y(n_235) );
AO22x2_ASAP7_75t_L g271 ( .A1(n_76), .A2(n_236), .B1(n_272), .B2(n_274), .Y(n_271) );
AOI221xp5_ASAP7_75t_L g77 ( .A1(n_78), .A2(n_93), .B1(n_499), .B2(n_605), .C(n_621), .Y(n_77) );
BUFx2_ASAP7_75t_L g78 ( .A(n_79), .Y(n_78) );
AND2x2_ASAP7_75t_L g79 ( .A(n_80), .B(n_90), .Y(n_79) );
OA21x2_ASAP7_75t_L g633 ( .A1(n_80), .A2(n_634), .B(n_635), .Y(n_633) );
NOR2xp33_ASAP7_75t_L g80 ( .A(n_81), .B(n_86), .Y(n_80) );
CKINVDCx16_ASAP7_75t_R g81 ( .A(n_82), .Y(n_81) );
HB1xp67_ASAP7_75t_L g82 ( .A(n_83), .Y(n_82) );
INVx1_ASAP7_75t_L g83 ( .A(n_84), .Y(n_83) );
INVxp67_ASAP7_75t_SL g174 ( .A(n_84), .Y(n_174) );
INVx2_ASAP7_75t_L g212 ( .A(n_84), .Y(n_212) );
INVx2_ASAP7_75t_L g84 ( .A(n_85), .Y(n_84) );
INVx3_ASAP7_75t_L g116 ( .A(n_85), .Y(n_116) );
INVx6_ASAP7_75t_L g123 ( .A(n_85), .Y(n_123) );
INVx2_ASAP7_75t_L g141 ( .A(n_85), .Y(n_141) );
HB1xp67_ASAP7_75t_L g86 ( .A(n_87), .Y(n_86) );
NOR2xp33_ASAP7_75t_L g145 ( .A(n_87), .B(n_137), .Y(n_145) );
INVx4_ASAP7_75t_L g87 ( .A(n_88), .Y(n_87) );
OAI22xp5_ASAP7_75t_L g236 ( .A1(n_88), .A2(n_237), .B1(n_238), .B2(n_239), .Y(n_236) );
AOI21xp5_ASAP7_75t_L g255 ( .A1(n_88), .A2(n_256), .B(n_258), .Y(n_255) );
BUFx6f_ASAP7_75t_L g88 ( .A(n_89), .Y(n_88) );
BUFx6f_ASAP7_75t_L g118 ( .A(n_89), .Y(n_118) );
INVx3_ASAP7_75t_L g125 ( .A(n_89), .Y(n_125) );
INVx1_ASAP7_75t_L g176 ( .A(n_89), .Y(n_176) );
INVx4_ASAP7_75t_L g207 ( .A(n_89), .Y(n_207) );
BUFx6f_ASAP7_75t_L g90 ( .A(n_91), .Y(n_90) );
AND2x2_ASAP7_75t_L g104 ( .A(n_91), .B(n_105), .Y(n_104) );
INVx3_ASAP7_75t_L g167 ( .A(n_91), .Y(n_167) );
AND2x2_ASAP7_75t_L g272 ( .A(n_91), .B(n_273), .Y(n_272) );
HB1xp67_ASAP7_75t_L g618 ( .A(n_92), .Y(n_618) );
INVx1_ASAP7_75t_L g93 ( .A(n_94), .Y(n_93) );
BUFx3_ASAP7_75t_L g94 ( .A(n_95), .Y(n_94) );
AND2x4_ASAP7_75t_L g95 ( .A(n_96), .B(n_423), .Y(n_95) );
NOR2xp67_ASAP7_75t_L g96 ( .A(n_97), .B(n_345), .Y(n_96) );
NAND3xp33_ASAP7_75t_L g97 ( .A(n_98), .B(n_287), .C(n_324), .Y(n_97) );
AOI21xp5_ASAP7_75t_L g98 ( .A1(n_99), .A2(n_196), .B(n_241), .Y(n_98) );
OAI31xp33_ASAP7_75t_L g99 ( .A1(n_100), .A2(n_129), .A3(n_158), .B(n_177), .Y(n_99) );
INVx1_ASAP7_75t_L g482 ( .A(n_100), .Y(n_482) );
BUFx3_ASAP7_75t_L g100 ( .A(n_101), .Y(n_100) );
OR2x2_ASAP7_75t_L g319 ( .A(n_101), .B(n_320), .Y(n_319) );
AND2x2_ASAP7_75t_L g351 ( .A(n_101), .B(n_352), .Y(n_351) );
NAND2xp5_ASAP7_75t_L g365 ( .A(n_101), .B(n_278), .Y(n_365) );
AND2x2_ASAP7_75t_L g469 ( .A(n_101), .B(n_455), .Y(n_469) );
INVx2_ASAP7_75t_L g101 ( .A(n_102), .Y(n_101) );
AND2x2_ASAP7_75t_L g343 ( .A(n_102), .B(n_299), .Y(n_343) );
AND2x2_ASAP7_75t_L g382 ( .A(n_102), .B(n_279), .Y(n_382) );
HB1xp67_ASAP7_75t_L g416 ( .A(n_102), .Y(n_416) );
INVx1_ASAP7_75t_L g102 ( .A(n_103), .Y(n_102) );
INVx1_ASAP7_75t_L g296 ( .A(n_103), .Y(n_296) );
INVx1_ASAP7_75t_L g315 ( .A(n_103), .Y(n_315) );
AOI21x1_ASAP7_75t_L g103 ( .A1(n_104), .A2(n_110), .B(n_126), .Y(n_103) );
INVx2_ASAP7_75t_L g105 ( .A(n_106), .Y(n_105) );
NOR2xp33_ASAP7_75t_L g182 ( .A(n_106), .B(n_167), .Y(n_182) );
INVx2_ASAP7_75t_L g106 ( .A(n_107), .Y(n_106) );
INVx4_ASAP7_75t_L g107 ( .A(n_108), .Y(n_107) );
INVx2_ASAP7_75t_L g128 ( .A(n_108), .Y(n_128) );
BUFx3_ASAP7_75t_L g153 ( .A(n_108), .Y(n_153) );
OAI22xp5_ASAP7_75t_L g110 ( .A1(n_111), .A2(n_117), .B1(n_119), .B2(n_124), .Y(n_110) );
INVx2_ASAP7_75t_L g112 ( .A(n_113), .Y(n_112) );
INVx2_ASAP7_75t_L g135 ( .A(n_113), .Y(n_135) );
INVx2_ASAP7_75t_L g113 ( .A(n_114), .Y(n_113) );
INVx2_ASAP7_75t_L g121 ( .A(n_114), .Y(n_121) );
INVx2_ASAP7_75t_L g115 ( .A(n_116), .Y(n_115) );
INVx1_ASAP7_75t_L g164 ( .A(n_116), .Y(n_164) );
INVx2_ASAP7_75t_L g185 ( .A(n_116), .Y(n_185) );
INVx1_ASAP7_75t_L g257 ( .A(n_116), .Y(n_257) );
INVx1_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
NAND2xp5_ASAP7_75t_SL g165 ( .A(n_118), .B(n_166), .Y(n_165) );
A2O1A1Ixp33_ASAP7_75t_L g183 ( .A1(n_118), .A2(n_184), .B(n_186), .C(n_187), .Y(n_183) );
A2O1A1Ixp33_ASAP7_75t_L g228 ( .A1(n_118), .A2(n_135), .B(n_229), .C(n_230), .Y(n_228) );
INVx1_ASAP7_75t_L g239 ( .A(n_118), .Y(n_239) );
INVx3_ASAP7_75t_L g215 ( .A(n_120), .Y(n_215) );
INVx2_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
INVx1_ASAP7_75t_L g188 ( .A(n_121), .Y(n_188) );
INVx1_ASAP7_75t_L g225 ( .A(n_122), .Y(n_225) );
INVx1_ASAP7_75t_L g122 ( .A(n_123), .Y(n_122) );
INVx2_ASAP7_75t_L g150 ( .A(n_123), .Y(n_150) );
INVx2_ASAP7_75t_L g204 ( .A(n_123), .Y(n_204) );
INVx2_ASAP7_75t_SL g217 ( .A(n_123), .Y(n_217) );
NOR2xp33_ASAP7_75t_L g136 ( .A(n_124), .B(n_137), .Y(n_136) );
NOR3xp33_ASAP7_75t_L g142 ( .A(n_124), .B(n_137), .C(n_143), .Y(n_142) );
INVx3_ASAP7_75t_L g124 ( .A(n_125), .Y(n_124) );
A2O1A1Ixp33_ASAP7_75t_L g189 ( .A1(n_125), .A2(n_190), .B(n_191), .C(n_192), .Y(n_189) );
A2O1A1Ixp33_ASAP7_75t_L g224 ( .A1(n_125), .A2(n_225), .B(n_226), .C(n_227), .Y(n_224) );
NOR2xp33_ASAP7_75t_L g126 ( .A(n_127), .B(n_128), .Y(n_126) );
BUFx3_ASAP7_75t_L g219 ( .A(n_128), .Y(n_219) );
NOR2xp33_ASAP7_75t_L g220 ( .A(n_128), .B(n_221), .Y(n_220) );
INVx3_ASAP7_75t_L g253 ( .A(n_128), .Y(n_253) );
INVx2_ASAP7_75t_L g306 ( .A(n_129), .Y(n_306) );
NAND2xp5_ASAP7_75t_L g399 ( .A(n_129), .B(n_307), .Y(n_399) );
BUFx2_ASAP7_75t_L g129 ( .A(n_130), .Y(n_129) );
OR2x2_ASAP7_75t_L g180 ( .A(n_130), .B(n_181), .Y(n_180) );
INVx2_ASAP7_75t_L g284 ( .A(n_130), .Y(n_284) );
AND2x2_ASAP7_75t_L g417 ( .A(n_130), .B(n_320), .Y(n_417) );
AO21x2_ASAP7_75t_L g130 ( .A1(n_131), .A2(n_152), .B(n_154), .Y(n_130) );
AO21x2_ASAP7_75t_L g247 ( .A1(n_131), .A2(n_154), .B(n_248), .Y(n_247) );
NAND2xp5_ASAP7_75t_L g131 ( .A(n_132), .B(n_144), .Y(n_131) );
AOI22xp5_ASAP7_75t_L g132 ( .A1(n_133), .A2(n_136), .B1(n_139), .B2(n_142), .Y(n_132) );
NOR2xp67_ASAP7_75t_L g133 ( .A(n_134), .B(n_135), .Y(n_133) );
AOI221x1_ASAP7_75t_L g201 ( .A1(n_137), .A2(n_202), .B1(n_205), .B2(n_209), .C(n_211), .Y(n_201) );
INVx4_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
INVx1_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
INVx1_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
INVx2_ASAP7_75t_L g173 ( .A(n_141), .Y(n_173) );
NAND2xp5_ASAP7_75t_L g144 ( .A(n_145), .B(n_146), .Y(n_144) );
OAI22xp33_ASAP7_75t_L g146 ( .A1(n_147), .A2(n_149), .B1(n_150), .B2(n_151), .Y(n_146) );
INVx2_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
INVx2_ASAP7_75t_L g163 ( .A(n_148), .Y(n_163) );
INVx2_ASAP7_75t_L g191 ( .A(n_148), .Y(n_191) );
INVx2_ASAP7_75t_L g259 ( .A(n_148), .Y(n_259) );
INVx1_ASAP7_75t_L g263 ( .A(n_148), .Y(n_263) );
NAND2xp5_ASAP7_75t_L g264 ( .A(n_150), .B(n_265), .Y(n_264) );
INVx3_ASAP7_75t_L g152 ( .A(n_153), .Y(n_152) );
NOR2xp33_ASAP7_75t_L g154 ( .A(n_155), .B(n_156), .Y(n_154) );
INVx1_ASAP7_75t_L g240 ( .A(n_156), .Y(n_240) );
INVx1_ASAP7_75t_L g156 ( .A(n_157), .Y(n_156) );
NOR2xp67_ASAP7_75t_L g166 ( .A(n_157), .B(n_167), .Y(n_166) );
BUFx3_ASAP7_75t_L g169 ( .A(n_157), .Y(n_169) );
INVx1_ASAP7_75t_L g194 ( .A(n_157), .Y(n_194) );
NOR2xp33_ASAP7_75t_L g231 ( .A(n_157), .B(n_167), .Y(n_231) );
NOR2xp33_ASAP7_75t_L g267 ( .A(n_157), .B(n_167), .Y(n_267) );
INVx1_ASAP7_75t_L g273 ( .A(n_157), .Y(n_273) );
BUFx3_ASAP7_75t_L g158 ( .A(n_159), .Y(n_158) );
AND2x2_ASAP7_75t_L g447 ( .A(n_159), .B(n_358), .Y(n_447) );
INVx1_ASAP7_75t_L g159 ( .A(n_160), .Y(n_159) );
INVx1_ASAP7_75t_L g179 ( .A(n_160), .Y(n_179) );
INVx2_ASAP7_75t_L g283 ( .A(n_160), .Y(n_283) );
AND2x2_ASAP7_75t_L g302 ( .A(n_160), .B(n_251), .Y(n_302) );
AND2x2_ASAP7_75t_L g307 ( .A(n_160), .B(n_308), .Y(n_307) );
NAND2x1p5_ASAP7_75t_L g160 ( .A(n_161), .B(n_170), .Y(n_160) );
AND2x2_ASAP7_75t_SL g246 ( .A(n_161), .B(n_170), .Y(n_246) );
OA21x2_ASAP7_75t_L g161 ( .A1(n_162), .A2(n_165), .B(n_168), .Y(n_161) );
NAND2xp5_ASAP7_75t_L g175 ( .A(n_166), .B(n_176), .Y(n_175) );
OR2x2_ASAP7_75t_L g170 ( .A(n_171), .B(n_175), .Y(n_170) );
INVx1_ASAP7_75t_L g172 ( .A(n_173), .Y(n_172) );
INVx2_ASAP7_75t_L g461 ( .A(n_177), .Y(n_461) );
OR2x2_ASAP7_75t_L g177 ( .A(n_178), .B(n_180), .Y(n_177) );
AND2x4_ASAP7_75t_L g386 ( .A(n_178), .B(n_387), .Y(n_386) );
INVx2_ASAP7_75t_L g178 ( .A(n_179), .Y(n_178) );
AND2x2_ASAP7_75t_L g401 ( .A(n_179), .B(n_285), .Y(n_401) );
INVx2_ASAP7_75t_L g363 ( .A(n_180), .Y(n_363) );
INVx1_ASAP7_75t_L g268 ( .A(n_181), .Y(n_268) );
INVx2_ASAP7_75t_L g286 ( .A(n_181), .Y(n_286) );
HB1xp67_ASAP7_75t_L g301 ( .A(n_181), .Y(n_301) );
INVx2_ASAP7_75t_L g320 ( .A(n_181), .Y(n_320) );
AND2x2_ASAP7_75t_L g334 ( .A(n_181), .B(n_247), .Y(n_334) );
INVx1_ASAP7_75t_L g359 ( .A(n_181), .Y(n_359) );
AO31x2_ASAP7_75t_L g181 ( .A1(n_182), .A2(n_183), .A3(n_189), .B(n_193), .Y(n_181) );
INVx1_ASAP7_75t_L g184 ( .A(n_185), .Y(n_184) );
NOR2xp33_ASAP7_75t_SL g193 ( .A(n_194), .B(n_195), .Y(n_193) );
NOR2xp33_ASAP7_75t_L g232 ( .A(n_194), .B(n_233), .Y(n_232) );
INVx1_ASAP7_75t_L g196 ( .A(n_197), .Y(n_196) );
INVx1_ASAP7_75t_L g197 ( .A(n_198), .Y(n_197) );
NAND2xp5_ASAP7_75t_L g435 ( .A(n_198), .B(n_436), .Y(n_435) );
AND2x2_ASAP7_75t_L g198 ( .A(n_199), .B(n_234), .Y(n_198) );
AND2x2_ASAP7_75t_L g290 ( .A(n_199), .B(n_291), .Y(n_290) );
INVx2_ASAP7_75t_L g318 ( .A(n_199), .Y(n_318) );
INVx2_ASAP7_75t_L g376 ( .A(n_199), .Y(n_376) );
AND2x2_ASAP7_75t_L g199 ( .A(n_200), .B(n_222), .Y(n_199) );
INVx2_ASAP7_75t_L g279 ( .A(n_200), .Y(n_279) );
NAND2xp5_ASAP7_75t_L g295 ( .A(n_200), .B(n_296), .Y(n_295) );
OR2x2_ASAP7_75t_L g350 ( .A(n_200), .B(n_296), .Y(n_350) );
INVx1_ASAP7_75t_L g391 ( .A(n_200), .Y(n_391) );
AND2x2_ASAP7_75t_L g455 ( .A(n_200), .B(n_299), .Y(n_455) );
AO31x2_ASAP7_75t_L g200 ( .A1(n_201), .A2(n_213), .A3(n_219), .B(n_220), .Y(n_200) );
INVx1_ASAP7_75t_L g202 ( .A(n_203), .Y(n_202) );
INVx1_ASAP7_75t_L g203 ( .A(n_204), .Y(n_203) );
AND2x2_ASAP7_75t_L g205 ( .A(n_206), .B(n_208), .Y(n_205) );
AND2x2_ASAP7_75t_L g209 ( .A(n_206), .B(n_210), .Y(n_209) );
INVx2_ASAP7_75t_L g206 ( .A(n_207), .Y(n_206) );
NOR2xp33_ASAP7_75t_L g265 ( .A(n_207), .B(n_266), .Y(n_265) );
INVx1_ASAP7_75t_L g211 ( .A(n_212), .Y(n_211) );
INVx1_ASAP7_75t_L g213 ( .A(n_214), .Y(n_213) );
NAND2xp5_ASAP7_75t_L g216 ( .A(n_217), .B(n_218), .Y(n_216) );
INVx2_ASAP7_75t_L g274 ( .A(n_219), .Y(n_274) );
BUFx3_ASAP7_75t_L g275 ( .A(n_222), .Y(n_275) );
INVx2_ASAP7_75t_L g299 ( .A(n_222), .Y(n_299) );
AND2x4_ASAP7_75t_L g311 ( .A(n_222), .B(n_312), .Y(n_311) );
INVx1_ASAP7_75t_L g353 ( .A(n_222), .Y(n_353) );
AND2x4_ASAP7_75t_L g390 ( .A(n_222), .B(n_391), .Y(n_390) );
INVx3_ASAP7_75t_L g222 ( .A(n_223), .Y(n_222) );
AO31x2_ASAP7_75t_L g223 ( .A1(n_224), .A2(n_228), .A3(n_231), .B(n_232), .Y(n_223) );
INVx1_ASAP7_75t_L g366 ( .A(n_234), .Y(n_366) );
INVx2_ASAP7_75t_L g368 ( .A(n_234), .Y(n_368) );
AND2x4_ASAP7_75t_L g397 ( .A(n_234), .B(n_382), .Y(n_397) );
AND2x2_ASAP7_75t_L g463 ( .A(n_234), .B(n_464), .Y(n_463) );
BUFx8_ASAP7_75t_L g234 ( .A(n_235), .Y(n_234) );
INVx2_ASAP7_75t_L g312 ( .A(n_235), .Y(n_312) );
AND2x2_ASAP7_75t_L g327 ( .A(n_235), .B(n_328), .Y(n_327) );
INVxp67_ASAP7_75t_L g248 ( .A(n_240), .Y(n_248) );
OAI22xp5_ASAP7_75t_L g241 ( .A1(n_242), .A2(n_269), .B1(n_276), .B2(n_280), .Y(n_241) );
NAND2xp5_ASAP7_75t_L g392 ( .A(n_242), .B(n_393), .Y(n_392) );
INVx2_ASAP7_75t_L g242 ( .A(n_243), .Y(n_242) );
AOI211xp5_ASAP7_75t_L g442 ( .A1(n_243), .A2(n_325), .B(n_443), .C(n_449), .Y(n_442) );
AND2x4_ASAP7_75t_L g243 ( .A(n_244), .B(n_249), .Y(n_243) );
AND2x2_ASAP7_75t_L g244 ( .A(n_245), .B(n_247), .Y(n_244) );
NOR2xp67_ASAP7_75t_SL g436 ( .A(n_245), .B(n_338), .Y(n_436) );
INVx2_ASAP7_75t_L g245 ( .A(n_246), .Y(n_245) );
AND2x2_ASAP7_75t_L g371 ( .A(n_246), .B(n_372), .Y(n_371) );
AND2x2_ASAP7_75t_L g378 ( .A(n_246), .B(n_372), .Y(n_378) );
INVx1_ASAP7_75t_L g484 ( .A(n_246), .Y(n_484) );
OR2x2_ASAP7_75t_L g323 ( .A(n_247), .B(n_308), .Y(n_323) );
AND2x2_ASAP7_75t_L g330 ( .A(n_247), .B(n_283), .Y(n_330) );
AND2x2_ASAP7_75t_L g448 ( .A(n_247), .B(n_250), .Y(n_448) );
AND2x2_ASAP7_75t_L g407 ( .A(n_249), .B(n_330), .Y(n_407) );
AND2x2_ASAP7_75t_L g249 ( .A(n_250), .B(n_268), .Y(n_249) );
OR2x2_ASAP7_75t_L g338 ( .A(n_250), .B(n_284), .Y(n_338) );
INVx1_ASAP7_75t_L g432 ( .A(n_250), .Y(n_432) );
INVx1_ASAP7_75t_L g250 ( .A(n_251), .Y(n_250) );
AND2x2_ASAP7_75t_L g285 ( .A(n_251), .B(n_286), .Y(n_285) );
INVx2_ASAP7_75t_L g308 ( .A(n_251), .Y(n_308) );
HB1xp67_ASAP7_75t_L g360 ( .A(n_251), .Y(n_360) );
INVx1_ASAP7_75t_L g372 ( .A(n_251), .Y(n_372) );
AND2x4_ASAP7_75t_L g251 ( .A(n_252), .B(n_254), .Y(n_251) );
OAI21xp5_ASAP7_75t_L g254 ( .A1(n_255), .A2(n_260), .B(n_267), .Y(n_254) );
OAI21xp5_ASAP7_75t_L g260 ( .A1(n_261), .A2(n_262), .B(n_264), .Y(n_260) );
INVx1_ASAP7_75t_L g262 ( .A(n_263), .Y(n_262) );
INVxp67_ASAP7_75t_L g344 ( .A(n_268), .Y(n_344) );
NAND2xp5_ASAP7_75t_L g470 ( .A(n_268), .B(n_458), .Y(n_470) );
A2O1A1Ixp33_ASAP7_75t_L g496 ( .A1(n_269), .A2(n_364), .B(n_497), .C(n_498), .Y(n_496) );
INVx2_ASAP7_75t_L g269 ( .A(n_270), .Y(n_269) );
AND2x4_ASAP7_75t_L g270 ( .A(n_271), .B(n_275), .Y(n_270) );
INVx1_ASAP7_75t_L g291 ( .A(n_271), .Y(n_291) );
AND2x4_ASAP7_75t_L g298 ( .A(n_271), .B(n_299), .Y(n_298) );
INVx1_ASAP7_75t_L g354 ( .A(n_271), .Y(n_354) );
AND2x2_ASAP7_75t_L g472 ( .A(n_271), .B(n_296), .Y(n_472) );
INVx2_ASAP7_75t_SL g348 ( .A(n_275), .Y(n_348) );
INVxp67_ASAP7_75t_SL g276 ( .A(n_277), .Y(n_276) );
NAND2xp5_ASAP7_75t_L g420 ( .A(n_277), .B(n_348), .Y(n_420) );
INVx1_ASAP7_75t_L g277 ( .A(n_278), .Y(n_277) );
AND2x2_ASAP7_75t_L g339 ( .A(n_278), .B(n_312), .Y(n_339) );
INVx2_ASAP7_75t_SL g278 ( .A(n_279), .Y(n_278) );
INVx1_ASAP7_75t_L g326 ( .A(n_279), .Y(n_326) );
NAND2xp5_ASAP7_75t_L g341 ( .A(n_279), .B(n_312), .Y(n_341) );
BUFx3_ASAP7_75t_L g439 ( .A(n_279), .Y(n_439) );
INVx1_ASAP7_75t_L g280 ( .A(n_281), .Y(n_280) );
AND2x2_ASAP7_75t_L g281 ( .A(n_282), .B(n_285), .Y(n_281) );
AOI22xp33_ASAP7_75t_SL g336 ( .A1(n_282), .A2(n_337), .B1(n_339), .B2(n_340), .Y(n_336) );
AND2x2_ASAP7_75t_L g282 ( .A(n_283), .B(n_284), .Y(n_282) );
HB1xp67_ASAP7_75t_L g411 ( .A(n_283), .Y(n_411) );
BUFx2_ASAP7_75t_L g458 ( .A(n_283), .Y(n_458) );
AND2x4_ASAP7_75t_L g395 ( .A(n_284), .B(n_396), .Y(n_395) );
AND2x2_ASAP7_75t_L g329 ( .A(n_285), .B(n_330), .Y(n_329) );
INVx1_ASAP7_75t_L g396 ( .A(n_286), .Y(n_396) );
AOI21xp5_ASAP7_75t_L g287 ( .A1(n_288), .A2(n_300), .B(n_303), .Y(n_287) );
NAND2xp5_ASAP7_75t_L g288 ( .A(n_289), .B(n_292), .Y(n_288) );
INVx2_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
NAND2xp5_ASAP7_75t_L g487 ( .A(n_290), .B(n_482), .Y(n_487) );
INVx1_ASAP7_75t_L g292 ( .A(n_293), .Y(n_292) );
AND2x2_ASAP7_75t_L g293 ( .A(n_294), .B(n_297), .Y(n_293) );
OAI21xp33_ASAP7_75t_SL g331 ( .A1(n_294), .A2(n_297), .B(n_332), .Y(n_331) );
INVx2_ASAP7_75t_L g427 ( .A(n_294), .Y(n_427) );
INVx1_ASAP7_75t_L g294 ( .A(n_295), .Y(n_294) );
INVx1_ASAP7_75t_L g464 ( .A(n_295), .Y(n_464) );
HB1xp67_ASAP7_75t_L g495 ( .A(n_296), .Y(n_495) );
INVx4_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
NAND2xp5_ASAP7_75t_L g381 ( .A(n_298), .B(n_382), .Y(n_381) );
AND2x2_ASAP7_75t_L g300 ( .A(n_301), .B(n_302), .Y(n_300) );
AND2x2_ASAP7_75t_L g333 ( .A(n_302), .B(n_334), .Y(n_333) );
INVx1_ASAP7_75t_L g414 ( .A(n_302), .Y(n_414) );
AND2x2_ASAP7_75t_L g462 ( .A(n_302), .B(n_417), .Y(n_462) );
OAI22xp5_ASAP7_75t_L g303 ( .A1(n_304), .A2(n_309), .B1(n_316), .B2(n_321), .Y(n_303) );
INVx1_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
AND2x2_ASAP7_75t_L g305 ( .A(n_306), .B(n_307), .Y(n_305) );
NOR2xp33_ASAP7_75t_L g488 ( .A(n_306), .B(n_489), .Y(n_488) );
NAND2xp67_ASAP7_75t_L g362 ( .A(n_307), .B(n_363), .Y(n_362) );
BUFx3_ASAP7_75t_L g384 ( .A(n_307), .Y(n_384) );
AND2x2_ASAP7_75t_L g492 ( .A(n_307), .B(n_395), .Y(n_492) );
AND2x2_ASAP7_75t_L g498 ( .A(n_307), .B(n_334), .Y(n_498) );
INVx1_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
AND2x2_ASAP7_75t_L g310 ( .A(n_311), .B(n_313), .Y(n_310) );
NAND2xp5_ASAP7_75t_L g332 ( .A(n_311), .B(n_314), .Y(n_332) );
INVx2_ASAP7_75t_L g444 ( .A(n_311), .Y(n_444) );
NAND2xp5_ASAP7_75t_L g406 ( .A(n_312), .B(n_328), .Y(n_406) );
INVx2_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
HB1xp67_ASAP7_75t_SL g379 ( .A(n_314), .Y(n_379) );
AND2x2_ASAP7_75t_L g480 ( .A(n_314), .B(n_390), .Y(n_480) );
BUFx3_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
INVx1_ASAP7_75t_L g328 ( .A(n_315), .Y(n_328) );
INVxp67_ASAP7_75t_SL g316 ( .A(n_317), .Y(n_316) );
NOR2xp67_ASAP7_75t_L g317 ( .A(n_318), .B(n_319), .Y(n_317) );
INVxp67_ASAP7_75t_SL g422 ( .A(n_320), .Y(n_422) );
INVx1_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
AND2x2_ASAP7_75t_L g467 ( .A(n_322), .B(n_447), .Y(n_467) );
INVx1_ASAP7_75t_L g322 ( .A(n_323), .Y(n_322) );
INVxp67_ASAP7_75t_L g387 ( .A(n_323), .Y(n_387) );
OR2x6_ASAP7_75t_L g421 ( .A(n_323), .B(n_422), .Y(n_421) );
INVxp67_ASAP7_75t_SL g441 ( .A(n_323), .Y(n_441) );
AOI221xp5_ASAP7_75t_L g324 ( .A1(n_325), .A2(n_329), .B1(n_331), .B2(n_333), .C(n_335), .Y(n_324) );
AND2x4_ASAP7_75t_SL g325 ( .A(n_326), .B(n_327), .Y(n_325) );
INVx1_ASAP7_75t_L g451 ( .A(n_327), .Y(n_451) );
AND2x4_ASAP7_75t_L g356 ( .A(n_330), .B(n_357), .Y(n_356) );
NOR3xp33_ASAP7_75t_L g335 ( .A(n_336), .B(n_342), .C(n_344), .Y(n_335) );
INVx1_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
INVxp67_ASAP7_75t_SL g340 ( .A(n_341), .Y(n_340) );
OR2x2_ASAP7_75t_L g494 ( .A(n_341), .B(n_495), .Y(n_494) );
INVx1_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
AND2x2_ASAP7_75t_L g438 ( .A(n_343), .B(n_439), .Y(n_438) );
NAND4xp25_ASAP7_75t_L g345 ( .A(n_346), .B(n_373), .C(n_389), .D(n_402), .Y(n_345) );
O2A1O1Ixp5_ASAP7_75t_L g346 ( .A1(n_347), .A2(n_351), .B(n_355), .C(n_361), .Y(n_346) );
AND2x2_ASAP7_75t_L g347 ( .A(n_348), .B(n_349), .Y(n_347) );
INVx1_ASAP7_75t_L g413 ( .A(n_348), .Y(n_413) );
OAI32xp33_ASAP7_75t_L g481 ( .A1(n_348), .A2(n_369), .A3(n_450), .B1(n_482), .B2(n_483), .Y(n_481) );
INVx2_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
OR2x2_ASAP7_75t_L g367 ( .A(n_350), .B(n_368), .Y(n_367) );
INVx2_ASAP7_75t_L g476 ( .A(n_350), .Y(n_476) );
INVx1_ASAP7_75t_L g412 ( .A(n_352), .Y(n_412) );
NAND2xp5_ASAP7_75t_L g475 ( .A(n_352), .B(n_476), .Y(n_475) );
AND2x2_ASAP7_75t_L g497 ( .A(n_352), .B(n_439), .Y(n_497) );
AND2x4_ASAP7_75t_SL g352 ( .A(n_353), .B(n_354), .Y(n_352) );
HB1xp67_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
AND2x2_ASAP7_75t_L g357 ( .A(n_358), .B(n_360), .Y(n_357) );
HB1xp67_ASAP7_75t_L g370 ( .A(n_358), .Y(n_370) );
INVx2_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
OAI32xp33_ASAP7_75t_L g361 ( .A1(n_362), .A2(n_364), .A3(n_366), .B1(n_367), .B2(n_369), .Y(n_361) );
AND2x2_ASAP7_75t_L g377 ( .A(n_363), .B(n_378), .Y(n_377) );
INVx2_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
INVx2_ASAP7_75t_L g428 ( .A(n_367), .Y(n_428) );
AND2x2_ASAP7_75t_L g454 ( .A(n_368), .B(n_455), .Y(n_454) );
NAND2xp5_ASAP7_75t_L g369 ( .A(n_370), .B(n_371), .Y(n_369) );
INVx1_ASAP7_75t_L g489 ( .A(n_371), .Y(n_489) );
AOI21xp5_ASAP7_75t_L g373 ( .A1(n_374), .A2(n_379), .B(n_380), .Y(n_373) );
AND2x2_ASAP7_75t_L g374 ( .A(n_375), .B(n_377), .Y(n_374) );
INVx1_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
HB1xp67_ASAP7_75t_L g388 ( .A(n_376), .Y(n_388) );
NAND2xp5_ASAP7_75t_L g404 ( .A(n_376), .B(n_405), .Y(n_404) );
AND2x2_ASAP7_75t_L g394 ( .A(n_378), .B(n_395), .Y(n_394) );
OAI22xp5_ASAP7_75t_L g380 ( .A1(n_381), .A2(n_383), .B1(n_385), .B2(n_388), .Y(n_380) );
NOR2xp33_ASAP7_75t_SL g419 ( .A(n_382), .B(n_405), .Y(n_419) );
INVx1_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
INVx3_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
AOI21xp33_ASAP7_75t_L g443 ( .A1(n_388), .A2(n_444), .B(n_445), .Y(n_443) );
AOI22xp33_ASAP7_75t_L g389 ( .A1(n_390), .A2(n_392), .B1(n_397), .B2(n_398), .Y(n_389) );
INVx2_ASAP7_75t_L g452 ( .A(n_390), .Y(n_452) );
NAND2xp5_ASAP7_75t_L g471 ( .A(n_390), .B(n_472), .Y(n_471) );
INVx2_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
AND2x4_ASAP7_75t_L g431 ( .A(n_395), .B(n_432), .Y(n_431) );
AND2x2_ASAP7_75t_L g457 ( .A(n_395), .B(n_458), .Y(n_457) );
NAND2xp5_ASAP7_75t_L g398 ( .A(n_399), .B(n_400), .Y(n_398) );
INVx1_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
AOI221xp5_ASAP7_75t_SL g402 ( .A1(n_403), .A2(n_407), .B1(n_408), .B2(n_415), .C(n_418), .Y(n_402) );
INVxp67_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
INVx1_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
OAI22xp5_ASAP7_75t_L g408 ( .A1(n_409), .A2(n_412), .B1(n_413), .B2(n_414), .Y(n_408) );
INVxp67_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
NAND2xp5_ASAP7_75t_L g430 ( .A(n_410), .B(n_431), .Y(n_430) );
INVx1_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
AND2x4_ASAP7_75t_L g440 ( .A(n_411), .B(n_441), .Y(n_440) );
AND2x4_ASAP7_75t_L g415 ( .A(n_416), .B(n_417), .Y(n_415) );
INVx2_ASAP7_75t_L g479 ( .A(n_417), .Y(n_479) );
NAND2x1p5_ASAP7_75t_L g483 ( .A(n_417), .B(n_484), .Y(n_483) );
AOI21xp5_ASAP7_75t_L g418 ( .A1(n_419), .A2(n_420), .B(n_421), .Y(n_418) );
NOR2x1_ASAP7_75t_L g423 ( .A(n_424), .B(n_459), .Y(n_423) );
NAND3xp33_ASAP7_75t_L g424 ( .A(n_425), .B(n_433), .C(n_442), .Y(n_424) );
OAI21xp33_ASAP7_75t_L g425 ( .A1(n_426), .A2(n_428), .B(n_429), .Y(n_425) );
CKINVDCx5p33_ASAP7_75t_R g426 ( .A(n_427), .Y(n_426) );
INVx1_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
INVxp67_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
NAND2xp5_ASAP7_75t_L g434 ( .A(n_435), .B(n_437), .Y(n_434) );
AOI221xp5_ASAP7_75t_L g473 ( .A1(n_436), .A2(n_474), .B1(n_477), .B2(n_480), .C(n_481), .Y(n_473) );
NAND2xp5_ASAP7_75t_L g437 ( .A(n_438), .B(n_440), .Y(n_437) );
INVx2_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
AND2x4_ASAP7_75t_L g446 ( .A(n_447), .B(n_448), .Y(n_446) );
AOI21xp5_ASAP7_75t_L g449 ( .A1(n_450), .A2(n_453), .B(n_456), .Y(n_449) );
OR2x2_ASAP7_75t_L g450 ( .A(n_451), .B(n_452), .Y(n_450) );
INVx2_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
INVx1_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
INVx1_ASAP7_75t_L g478 ( .A(n_458), .Y(n_478) );
NAND3xp33_ASAP7_75t_SL g459 ( .A(n_460), .B(n_473), .C(n_485), .Y(n_459) );
O2A1O1Ixp33_ASAP7_75t_L g460 ( .A1(n_461), .A2(n_462), .B(n_463), .C(n_465), .Y(n_460) );
OAI22xp5_ASAP7_75t_L g465 ( .A1(n_466), .A2(n_468), .B1(n_470), .B2(n_471), .Y(n_465) );
INVx1_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
INVx1_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
INVx1_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
NOR2x1p5_ASAP7_75t_L g477 ( .A(n_478), .B(n_479), .Y(n_477) );
AOI21xp5_ASAP7_75t_L g485 ( .A1(n_486), .A2(n_488), .B(n_490), .Y(n_485) );
INVx1_ASAP7_75t_L g486 ( .A(n_487), .Y(n_486) );
OAI21xp5_ASAP7_75t_L g490 ( .A1(n_491), .A2(n_493), .B(n_496), .Y(n_490) );
INVx2_ASAP7_75t_L g491 ( .A(n_492), .Y(n_491) );
HB1xp67_ASAP7_75t_L g493 ( .A(n_494), .Y(n_493) );
XOR2xp5_ASAP7_75t_L g499 ( .A(n_500), .B(n_594), .Y(n_499) );
OAI22xp33_ASAP7_75t_SL g500 ( .A1(n_501), .A2(n_502), .B1(n_503), .B2(n_593), .Y(n_500) );
CKINVDCx5p33_ASAP7_75t_R g593 ( .A(n_501), .Y(n_593) );
OAI22xp33_ASAP7_75t_L g622 ( .A1(n_502), .A2(n_503), .B1(n_623), .B2(n_624), .Y(n_622) );
INVx1_ASAP7_75t_L g502 ( .A(n_503), .Y(n_502) );
HB1xp67_ASAP7_75t_L g503 ( .A(n_504), .Y(n_503) );
AND3x1_ASAP7_75t_L g504 ( .A(n_505), .B(n_552), .C(n_582), .Y(n_504) );
AND2x2_ASAP7_75t_L g505 ( .A(n_506), .B(n_536), .Y(n_505) );
INVx1_ASAP7_75t_L g507 ( .A(n_508), .Y(n_507) );
INVx3_ASAP7_75t_L g508 ( .A(n_509), .Y(n_508) );
AND2x4_ASAP7_75t_L g509 ( .A(n_510), .B(n_521), .Y(n_509) );
AND2x2_ASAP7_75t_L g533 ( .A(n_510), .B(n_534), .Y(n_533) );
AND2x4_ASAP7_75t_L g585 ( .A(n_510), .B(n_586), .Y(n_585) );
AND2x4_ASAP7_75t_L g589 ( .A(n_510), .B(n_539), .Y(n_589) );
AND2x4_ASAP7_75t_L g510 ( .A(n_511), .B(n_519), .Y(n_510) );
AND2x2_ASAP7_75t_L g556 ( .A(n_511), .B(n_520), .Y(n_556) );
INVx1_ASAP7_75t_L g511 ( .A(n_512), .Y(n_511) );
AND2x2_ASAP7_75t_L g538 ( .A(n_512), .B(n_520), .Y(n_538) );
NAND2xp5_ASAP7_75t_L g512 ( .A(n_513), .B(n_516), .Y(n_512) );
NAND2xp33_ASAP7_75t_L g513 ( .A(n_514), .B(n_515), .Y(n_513) );
INVx2_ASAP7_75t_L g518 ( .A(n_514), .Y(n_518) );
INVx3_ASAP7_75t_L g524 ( .A(n_514), .Y(n_524) );
NAND2xp33_ASAP7_75t_L g530 ( .A(n_514), .B(n_531), .Y(n_530) );
INVx1_ASAP7_75t_L g551 ( .A(n_514), .Y(n_551) );
HB1xp67_ASAP7_75t_L g563 ( .A(n_514), .Y(n_563) );
NAND2xp5_ASAP7_75t_L g548 ( .A(n_515), .B(n_549), .Y(n_548) );
INVxp67_ASAP7_75t_L g614 ( .A(n_515), .Y(n_614) );
NAND2xp5_ASAP7_75t_L g516 ( .A(n_517), .B(n_518), .Y(n_516) );
OAI21xp5_ASAP7_75t_L g577 ( .A1(n_517), .A2(n_551), .B(n_578), .Y(n_577) );
INVx1_ASAP7_75t_L g519 ( .A(n_520), .Y(n_519) );
AND2x2_ASAP7_75t_L g576 ( .A(n_520), .B(n_577), .Y(n_576) );
AND2x4_ASAP7_75t_L g571 ( .A(n_521), .B(n_538), .Y(n_571) );
AND2x4_ASAP7_75t_L g580 ( .A(n_521), .B(n_556), .Y(n_580) );
AND2x4_ASAP7_75t_L g521 ( .A(n_522), .B(n_526), .Y(n_521) );
INVx2_ASAP7_75t_L g535 ( .A(n_522), .Y(n_535) );
OR2x2_ASAP7_75t_L g540 ( .A(n_522), .B(n_541), .Y(n_540) );
AND2x2_ASAP7_75t_L g573 ( .A(n_522), .B(n_574), .Y(n_573) );
AND2x4_ASAP7_75t_L g586 ( .A(n_522), .B(n_587), .Y(n_586) );
AND2x4_ASAP7_75t_L g522 ( .A(n_523), .B(n_525), .Y(n_522) );
NAND2xp5_ASAP7_75t_L g528 ( .A(n_524), .B(n_529), .Y(n_528) );
INVxp67_ASAP7_75t_L g547 ( .A(n_524), .Y(n_547) );
NAND3xp33_ASAP7_75t_L g567 ( .A(n_525), .B(n_546), .C(n_568), .Y(n_567) );
AND2x4_ASAP7_75t_L g534 ( .A(n_526), .B(n_535), .Y(n_534) );
INVx1_ASAP7_75t_L g526 ( .A(n_527), .Y(n_526) );
INVx1_ASAP7_75t_L g541 ( .A(n_527), .Y(n_541) );
AND2x2_ASAP7_75t_L g527 ( .A(n_528), .B(n_530), .Y(n_527) );
BUFx3_ASAP7_75t_L g532 ( .A(n_533), .Y(n_532) );
AND2x2_ASAP7_75t_L g554 ( .A(n_534), .B(n_538), .Y(n_554) );
AND2x2_ASAP7_75t_L g555 ( .A(n_534), .B(n_556), .Y(n_555) );
AND2x4_ASAP7_75t_L g581 ( .A(n_534), .B(n_545), .Y(n_581) );
AND2x4_ASAP7_75t_L g537 ( .A(n_538), .B(n_539), .Y(n_537) );
AND2x4_ASAP7_75t_L g591 ( .A(n_538), .B(n_586), .Y(n_591) );
AND2x4_ASAP7_75t_L g544 ( .A(n_539), .B(n_545), .Y(n_544) );
INVx2_ASAP7_75t_L g539 ( .A(n_540), .Y(n_539) );
INVx1_ASAP7_75t_L g587 ( .A(n_541), .Y(n_587) );
INVx3_ASAP7_75t_L g542 ( .A(n_543), .Y(n_542) );
INVx6_ASAP7_75t_L g543 ( .A(n_544), .Y(n_543) );
AND2x4_ASAP7_75t_L g592 ( .A(n_545), .B(n_586), .Y(n_592) );
AND2x2_ASAP7_75t_L g545 ( .A(n_546), .B(n_550), .Y(n_545) );
NAND2xp5_ASAP7_75t_L g546 ( .A(n_547), .B(n_548), .Y(n_546) );
HB1xp67_ASAP7_75t_L g615 ( .A(n_549), .Y(n_615) );
AND2x2_ASAP7_75t_L g552 ( .A(n_553), .B(n_569), .Y(n_552) );
NOR2xp33_ASAP7_75t_L g557 ( .A(n_558), .B(n_559), .Y(n_557) );
INVx3_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
INVx3_ASAP7_75t_L g560 ( .A(n_561), .Y(n_560) );
AO21x2_ASAP7_75t_L g561 ( .A1(n_562), .A2(n_564), .B(n_567), .Y(n_561) );
INVx1_ASAP7_75t_L g562 ( .A(n_563), .Y(n_562) );
NAND2xp5_ASAP7_75t_L g574 ( .A(n_563), .B(n_575), .Y(n_574) );
NAND2xp5_ASAP7_75t_L g564 ( .A(n_565), .B(n_566), .Y(n_564) );
AND2x2_ASAP7_75t_L g569 ( .A(n_570), .B(n_579), .Y(n_569) );
AND2x4_ASAP7_75t_L g572 ( .A(n_573), .B(n_576), .Y(n_572) );
HB1xp67_ASAP7_75t_L g611 ( .A(n_575), .Y(n_611) );
AND2x2_ASAP7_75t_L g582 ( .A(n_583), .B(n_590), .Y(n_582) );
BUFx12f_ASAP7_75t_L g584 ( .A(n_585), .Y(n_584) );
BUFx6f_ASAP7_75t_L g588 ( .A(n_589), .Y(n_588) );
AOI22xp5_ASAP7_75t_L g594 ( .A1(n_595), .A2(n_596), .B1(n_603), .B2(n_604), .Y(n_594) );
CKINVDCx5p33_ASAP7_75t_R g603 ( .A(n_595), .Y(n_603) );
CKINVDCx20_ASAP7_75t_R g604 ( .A(n_596), .Y(n_604) );
AOI22xp5_ASAP7_75t_L g596 ( .A1(n_597), .A2(n_598), .B1(n_599), .B2(n_602), .Y(n_596) );
CKINVDCx5p33_ASAP7_75t_R g602 ( .A(n_597), .Y(n_602) );
INVx1_ASAP7_75t_L g598 ( .A(n_599), .Y(n_598) );
XOR2xp5_ASAP7_75t_L g599 ( .A(n_600), .B(n_601), .Y(n_599) );
BUFx3_ASAP7_75t_L g605 ( .A(n_606), .Y(n_605) );
CKINVDCx5p33_ASAP7_75t_R g606 ( .A(n_607), .Y(n_606) );
NAND2xp5_ASAP7_75t_L g607 ( .A(n_608), .B(n_616), .Y(n_607) );
INVxp67_ASAP7_75t_SL g608 ( .A(n_609), .Y(n_608) );
AND2x2_ASAP7_75t_L g626 ( .A(n_609), .B(n_616), .Y(n_626) );
AOI211xp5_ASAP7_75t_L g609 ( .A1(n_610), .A2(n_611), .B(n_612), .C(n_615), .Y(n_609) );
NOR2xp33_ASAP7_75t_L g612 ( .A(n_613), .B(n_614), .Y(n_612) );
NOR2xp33_ASAP7_75t_L g616 ( .A(n_617), .B(n_619), .Y(n_616) );
OR2x2_ASAP7_75t_L g631 ( .A(n_617), .B(n_620), .Y(n_631) );
INVx1_ASAP7_75t_L g634 ( .A(n_617), .Y(n_634) );
NAND2xp5_ASAP7_75t_L g635 ( .A(n_617), .B(n_619), .Y(n_635) );
HB1xp67_ASAP7_75t_L g617 ( .A(n_618), .Y(n_617) );
INVx1_ASAP7_75t_L g619 ( .A(n_620), .Y(n_619) );
OAI222xp33_ASAP7_75t_L g621 ( .A1(n_622), .A2(n_625), .B1(n_627), .B2(n_630), .C1(n_632), .C2(n_636), .Y(n_621) );
CKINVDCx20_ASAP7_75t_R g623 ( .A(n_624), .Y(n_623) );
INVx1_ASAP7_75t_SL g625 ( .A(n_626), .Y(n_625) );
INVx1_ASAP7_75t_L g627 ( .A(n_628), .Y(n_627) );
HB1xp67_ASAP7_75t_L g630 ( .A(n_631), .Y(n_630) );
BUFx3_ASAP7_75t_L g632 ( .A(n_633), .Y(n_632) );
endmodule