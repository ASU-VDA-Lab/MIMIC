module fake_ariane_2166_n_1828 (n_83, n_8, n_56, n_60, n_170, n_160, n_64, n_119, n_124, n_167, n_90, n_38, n_47, n_110, n_153, n_18, n_86, n_75, n_89, n_67, n_176, n_149, n_34, n_158, n_172, n_69, n_95, n_175, n_92, n_143, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_152, n_120, n_169, n_106, n_12, n_53, n_173, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_156, n_49, n_20, n_174, n_100, n_17, n_50, n_132, n_62, n_147, n_51, n_166, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_159, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_148, n_164, n_52, n_157, n_135, n_73, n_77, n_171, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_151, n_136, n_28, n_80, n_146, n_97, n_154, n_142, n_161, n_14, n_163, n_88, n_141, n_68, n_116, n_104, n_145, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_1828);

input n_83;
input n_8;
input n_56;
input n_60;
input n_170;
input n_160;
input n_64;
input n_119;
input n_124;
input n_167;
input n_90;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_176;
input n_149;
input n_34;
input n_158;
input n_172;
input n_69;
input n_95;
input n_175;
input n_92;
input n_143;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_152;
input n_120;
input n_169;
input n_106;
input n_12;
input n_53;
input n_173;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_156;
input n_49;
input n_20;
input n_174;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_147;
input n_51;
input n_166;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_159;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_164;
input n_52;
input n_157;
input n_135;
input n_73;
input n_77;
input n_171;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_151;
input n_136;
input n_28;
input n_80;
input n_146;
input n_97;
input n_154;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_1828;

wire n_913;
wire n_1681;
wire n_1507;
wire n_1486;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_1250;
wire n_1169;
wire n_789;
wire n_850;
wire n_610;
wire n_245;
wire n_1713;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_187;
wire n_1463;
wire n_1238;
wire n_1515;
wire n_817;
wire n_924;
wire n_781;
wire n_1566;
wire n_189;
wire n_717;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_1706;
wire n_524;
wire n_1214;
wire n_634;
wire n_1246;
wire n_1138;
wire n_214;
wire n_764;
wire n_1503;
wire n_462;
wire n_1196;
wire n_1181;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1745;
wire n_1366;
wire n_232;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1457;
wire n_377;
wire n_1682;
wire n_520;
wire n_870;
wire n_1453;
wire n_279;
wire n_958;
wire n_945;
wire n_813;
wire n_419;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1184;
wire n_202;
wire n_1535;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_1277;
wire n_1746;
wire n_829;
wire n_1761;
wire n_1062;
wire n_339;
wire n_738;
wire n_1690;
wire n_672;
wire n_740;
wire n_1283;
wire n_1736;
wire n_1018;
wire n_259;
wire n_953;
wire n_1364;
wire n_1224;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_1688;
wire n_989;
wire n_645;
wire n_242;
wire n_331;
wire n_559;
wire n_495;
wire n_267;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_200;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_1522;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_1404;
wire n_868;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_1676;
wire n_1085;
wire n_277;
wire n_1636;
wire n_432;
wire n_293;
wire n_823;
wire n_620;
wire n_1074;
wire n_859;
wire n_1765;
wire n_587;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_352;
wire n_206;
wire n_899;
wire n_1703;
wire n_611;
wire n_1295;
wire n_238;
wire n_365;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_334;
wire n_192;
wire n_661;
wire n_1751;
wire n_300;
wire n_533;
wire n_438;
wire n_1654;
wire n_1560;
wire n_1548;
wire n_1811;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_376;
wire n_512;
wire n_1597;
wire n_1771;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1354;
wire n_1790;
wire n_1213;
wire n_237;
wire n_780;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_209;
wire n_490;
wire n_1461;
wire n_1391;
wire n_225;
wire n_1599;
wire n_1006;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_1594;
wire n_680;
wire n_287;
wire n_1716;
wire n_302;
wire n_380;
wire n_1585;
wire n_1432;
wire n_249;
wire n_1108;
wire n_355;
wire n_212;
wire n_444;
wire n_851;
wire n_1590;
wire n_1351;
wire n_1274;
wire n_257;
wire n_652;
wire n_1819;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_182;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_407;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_460;
wire n_1555;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_992;
wire n_966;
wire n_955;
wire n_1182;
wire n_794;
wire n_1692;
wire n_1562;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_288;
wire n_179;
wire n_1292;
wire n_1178;
wire n_1435;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_306;
wire n_203;
wire n_436;
wire n_324;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_437;
wire n_337;
wire n_274;
wire n_967;
wire n_1083;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1787;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_1717;
wire n_1812;
wire n_824;
wire n_428;
wire n_892;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_990;
wire n_1623;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_1780;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1825;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1680;
wire n_964;
wire n_1627;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_1731;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_934;
wire n_1447;
wire n_1220;
wire n_356;
wire n_698;
wire n_1674;
wire n_307;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_1633;
wire n_404;
wire n_1058;
wire n_347;
wire n_1042;
wire n_183;
wire n_1234;
wire n_479;
wire n_1578;
wire n_1455;
wire n_299;
wire n_836;
wire n_1279;
wire n_564;
wire n_205;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_1689;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_1728;
wire n_370;
wire n_706;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_1817;
wire n_552;
wire n_348;
wire n_670;
wire n_1826;
wire n_379;
wire n_264;
wire n_441;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_1618;
wire n_1743;
wire n_905;
wire n_207;
wire n_720;
wire n_926;
wire n_194;
wire n_1802;
wire n_1163;
wire n_186;
wire n_1795;
wire n_1384;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1648;
wire n_1413;
wire n_855;
wire n_808;
wire n_1365;
wire n_553;
wire n_1439;
wire n_814;
wire n_578;
wire n_1665;
wire n_1287;
wire n_405;
wire n_1611;
wire n_320;
wire n_1414;
wire n_1134;
wire n_1484;
wire n_647;
wire n_1423;
wire n_481;
wire n_600;
wire n_1053;
wire n_1609;
wire n_529;
wire n_502;
wire n_218;
wire n_1467;
wire n_247;
wire n_1798;
wire n_1304;
wire n_1608;
wire n_1744;
wire n_1105;
wire n_547;
wire n_439;
wire n_604;
wire n_677;
wire n_478;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_1278;
wire n_707;
wire n_983;
wire n_590;
wire n_699;
wire n_727;
wire n_301;
wire n_1726;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_325;
wire n_1740;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_729;
wire n_887;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_1693;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1823;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_233;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_321;
wire n_221;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1763;
wire n_1666;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_281;
wire n_262;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_1667;
wire n_845;
wire n_888;
wire n_1649;
wire n_1677;
wire n_1297;
wire n_178;
wire n_551;
wire n_417;
wire n_1708;
wire n_343;
wire n_1222;
wire n_582;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_534;
wire n_1791;
wire n_1460;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_451;
wire n_745;
wire n_1741;
wire n_1572;
wire n_1793;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_769;
wire n_1797;
wire n_1753;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_982;
wire n_1800;
wire n_915;
wire n_215;
wire n_1075;
wire n_454;
wire n_298;
wire n_1331;
wire n_1529;
wire n_1227;
wire n_655;
wire n_1734;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_1700;
wire n_659;
wire n_1332;
wire n_509;
wire n_666;
wire n_1747;
wire n_430;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1766;
wire n_1338;
wire n_1342;
wire n_456;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_521;
wire n_873;
wire n_1301;
wire n_1748;
wire n_1243;
wire n_1400;
wire n_342;
wire n_1466;
wire n_1513;
wire n_1527;
wire n_358;
wire n_1783;
wire n_608;
wire n_1538;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1668;
wire n_1605;
wire n_1078;
wire n_266;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_687;
wire n_797;
wire n_1786;
wire n_480;
wire n_1327;
wire n_1475;
wire n_211;
wire n_642;
wire n_1804;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_1757;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_393;
wire n_1632;
wire n_1769;
wire n_474;
wire n_805;
wire n_295;
wire n_1658;
wire n_190;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_180;
wire n_730;
wire n_386;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1137;
wire n_1258;
wire n_640;
wire n_197;
wire n_463;
wire n_1476;
wire n_1524;
wire n_1733;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_1807;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_1784;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_283;
wire n_806;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_1824;
wire n_643;
wire n_1492;
wire n_226;
wire n_1441;
wire n_1822;
wire n_682;
wire n_1616;
wire n_819;
wire n_586;
wire n_1324;
wire n_1429;
wire n_1778;
wire n_1776;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1759;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_1815;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_198;
wire n_1208;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1577;
wire n_1448;
wire n_1009;
wire n_230;
wire n_1133;
wire n_883;
wire n_473;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_594;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_1201;
wire n_1288;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_426;
wire n_433;
wire n_398;
wire n_210;
wire n_1090;
wire n_1367;
wire n_253;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_224;
wire n_894;
wire n_1380;
wire n_1624;
wire n_1801;
wire n_420;
wire n_1291;
wire n_562;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1023;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_467;
wire n_1511;
wire n_1422;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_1641;
wire n_538;
wire n_1517;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_1307;
wire n_1128;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1773;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_810;
wire n_1290;
wire n_181;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_628;
wire n_1300;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_414;
wire n_571;
wire n_1521;
wire n_1694;
wire n_284;
wire n_593;
wire n_1695;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_1774;
wire n_409;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_526;
wire n_1767;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1444;
wire n_1803;
wire n_820;
wire n_1749;
wire n_872;
wire n_1653;
wire n_254;
wire n_1157;
wire n_1584;
wire n_234;
wire n_848;
wire n_1664;
wire n_280;
wire n_629;
wire n_1739;
wire n_1814;
wire n_532;
wire n_1789;
wire n_763;
wire n_540;
wire n_216;
wire n_692;
wire n_984;
wire n_1687;
wire n_223;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_1816;
wire n_1756;
wire n_1606;
wire n_395;
wire n_621;
wire n_1587;
wire n_213;
wire n_1772;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_493;
wire n_1311;
wire n_1589;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_697;
wire n_622;
wire n_1626;
wire n_1335;
wire n_1715;
wire n_296;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_1785;
wire n_792;
wire n_1262;
wire n_580;
wire n_1579;
wire n_494;
wire n_434;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1183;
wire n_1326;
wire n_1805;
wire n_981;
wire n_1110;
wire n_1758;
wire n_243;
wire n_1407;
wire n_185;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_184;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_1054;
wire n_508;
wire n_1679;
wire n_353;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_191;
wire n_1011;
wire n_978;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_1721;
wire n_653;
wire n_1445;
wire n_1317;
wire n_783;
wire n_556;
wire n_1127;
wire n_1536;
wire n_1471;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_541;
wire n_499;
wire n_1775;
wire n_788;
wire n_908;
wire n_1036;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_1663;
wire n_1625;
wire n_318;
wire n_1458;
wire n_679;
wire n_244;
wire n_1630;
wire n_220;
wire n_663;
wire n_1720;
wire n_443;
wire n_1412;
wire n_1738;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_1735;
wire n_1788;
wire n_391;
wire n_940;
wire n_1537;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_765;
wire n_1809;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_1530;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_857;
wire n_898;
wire n_363;
wire n_968;
wire n_1067;
wire n_1323;
wire n_1235;
wire n_1462;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_1755;
wire n_1285;
wire n_193;
wire n_733;
wire n_761;
wire n_731;
wire n_336;
wire n_1813;
wire n_315;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_1106;
wire n_648;
wire n_784;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_1348;
wire n_753;
wire n_1770;
wire n_701;
wire n_1003;
wire n_1125;
wire n_1710;
wire n_309;
wire n_1344;
wire n_1390;
wire n_401;
wire n_485;
wire n_1792;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_291;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1510;
wire n_1099;
wire n_839;
wire n_1754;
wire n_759;
wire n_567;
wire n_240;
wire n_369;
wire n_1727;
wire n_1575;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_188;
wire n_323;
wire n_550;
wire n_1315;
wire n_1660;
wire n_997;
wire n_635;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_248;
wire n_1152;
wire n_921;
wire n_1615;
wire n_1236;
wire n_228;
wire n_1265;
wire n_1576;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1806;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1684;
wire n_1673;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_1696;
wire n_498;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1497;
wire n_459;
wire n_1136;
wire n_1782;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_383;
wire n_838;
wire n_1558;
wire n_1316;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_1781;
wire n_709;
wire n_809;
wire n_1686;
wire n_235;
wire n_881;
wire n_1019;
wire n_1477;
wire n_1777;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_199;
wire n_217;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_708;
wire n_308;
wire n_1223;
wire n_201;
wire n_1768;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1041;
wire n_993;
wire n_948;
wire n_922;
wire n_1004;
wire n_1810;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_1764;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_196;
wire n_1337;
wire n_774;
wire n_933;
wire n_1779;
wire n_596;
wire n_954;
wire n_1168;
wire n_1821;
wire n_219;
wire n_1310;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_252;
wire n_664;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_1732;
wire n_415;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1724;
wire n_1670;
wire n_1707;
wire n_1799;
wire n_1126;
wire n_195;
wire n_938;
wire n_1328;
wire n_895;
wire n_304;
wire n_1639;
wire n_583;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_946;
wire n_757;
wire n_375;
wire n_1655;
wire n_1818;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_472;
wire n_937;
wire n_1474;
wire n_265;
wire n_1583;
wire n_1604;
wire n_208;
wire n_1631;
wire n_1702;
wire n_275;
wire n_1794;
wire n_1375;
wire n_204;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_496;
wire n_1827;
wire n_866;
wire n_246;
wire n_925;
wire n_1752;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_1129;
wire n_1252;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_329;
wire n_718;
wire n_1434;
wire n_340;
wire n_1569;
wire n_289;
wire n_548;
wire n_523;
wire n_1662;
wire n_457;
wire n_1299;
wire n_177;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1228;
wire n_1244;
wire n_1796;
wire n_411;
wire n_484;
wire n_849;
wire n_1820;
wire n_357;
wire n_412;
wire n_1251;
wire n_447;
wire n_1421;
wire n_1762;
wire n_1233;
wire n_1808;
wire n_1574;
wire n_1672;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_1487;
wire n_675;

INVx1_ASAP7_75t_L g177 ( 
.A(n_163),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_108),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_106),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_114),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_59),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_156),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_127),
.Y(n_183)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_85),
.Y(n_184)
);

BUFx2_ASAP7_75t_SL g185 ( 
.A(n_0),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_59),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_81),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_19),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_111),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_137),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_98),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_43),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_27),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_153),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_1),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_145),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_155),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_58),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_4),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_138),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_54),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_84),
.Y(n_202)
);

INVx2_ASAP7_75t_SL g203 ( 
.A(n_44),
.Y(n_203)
);

BUFx3_ASAP7_75t_L g204 ( 
.A(n_1),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_41),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_113),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_40),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_105),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_40),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_101),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_42),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_73),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_52),
.Y(n_213)
);

BUFx10_ASAP7_75t_L g214 ( 
.A(n_117),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_169),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_71),
.Y(n_216)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_164),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_165),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_32),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_82),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_132),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_86),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_97),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_118),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_94),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_62),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_66),
.Y(n_227)
);

CKINVDCx16_ASAP7_75t_R g228 ( 
.A(n_151),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_142),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_95),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_173),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_90),
.Y(n_232)
);

INVx2_ASAP7_75t_SL g233 ( 
.A(n_53),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_15),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_103),
.Y(n_235)
);

INVx1_ASAP7_75t_SL g236 ( 
.A(n_121),
.Y(n_236)
);

INVxp67_ASAP7_75t_L g237 ( 
.A(n_63),
.Y(n_237)
);

CKINVDCx16_ASAP7_75t_R g238 ( 
.A(n_150),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_55),
.Y(n_239)
);

BUFx8_ASAP7_75t_SL g240 ( 
.A(n_12),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_5),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_76),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_58),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_126),
.Y(n_244)
);

INVx1_ASAP7_75t_SL g245 ( 
.A(n_19),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_36),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_93),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_4),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_99),
.Y(n_249)
);

BUFx5_ASAP7_75t_L g250 ( 
.A(n_0),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_161),
.Y(n_251)
);

BUFx3_ASAP7_75t_L g252 ( 
.A(n_141),
.Y(n_252)
);

INVx1_ASAP7_75t_SL g253 ( 
.A(n_77),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_74),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_140),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_7),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_162),
.Y(n_257)
);

INVx2_ASAP7_75t_SL g258 ( 
.A(n_26),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_61),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_158),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_147),
.Y(n_261)
);

INVx2_ASAP7_75t_SL g262 ( 
.A(n_32),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_91),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_122),
.Y(n_264)
);

CKINVDCx16_ASAP7_75t_R g265 ( 
.A(n_78),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_130),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_107),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_75),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_143),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_67),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_55),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_2),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_56),
.Y(n_273)
);

BUFx6f_ASAP7_75t_L g274 ( 
.A(n_87),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_115),
.Y(n_275)
);

BUFx2_ASAP7_75t_L g276 ( 
.A(n_120),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_174),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_15),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_134),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_27),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_17),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_53),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_135),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_50),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_109),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_149),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_13),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_44),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_52),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_20),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_57),
.Y(n_291)
);

INVx2_ASAP7_75t_L g292 ( 
.A(n_176),
.Y(n_292)
);

BUFx10_ASAP7_75t_L g293 ( 
.A(n_37),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_29),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_175),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_28),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_92),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_131),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_139),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_61),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_170),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_129),
.Y(n_302)
);

INVx2_ASAP7_75t_L g303 ( 
.A(n_8),
.Y(n_303)
);

BUFx8_ASAP7_75t_SL g304 ( 
.A(n_6),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_166),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_51),
.Y(n_306)
);

HB1xp67_ASAP7_75t_L g307 ( 
.A(n_5),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_18),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_16),
.Y(n_309)
);

BUFx6f_ASAP7_75t_L g310 ( 
.A(n_157),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_146),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_47),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_37),
.Y(n_313)
);

BUFx8_ASAP7_75t_SL g314 ( 
.A(n_172),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_128),
.Y(n_315)
);

INVx2_ASAP7_75t_L g316 ( 
.A(n_18),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_50),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_38),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_112),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_100),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_144),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_148),
.Y(n_322)
);

BUFx3_ASAP7_75t_L g323 ( 
.A(n_20),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_11),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_42),
.Y(n_325)
);

INVx2_ASAP7_75t_SL g326 ( 
.A(n_124),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_64),
.Y(n_327)
);

BUFx2_ASAP7_75t_L g328 ( 
.A(n_38),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_49),
.Y(n_329)
);

CKINVDCx20_ASAP7_75t_R g330 ( 
.A(n_70),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_51),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_30),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_24),
.Y(n_333)
);

CKINVDCx16_ASAP7_75t_R g334 ( 
.A(n_36),
.Y(n_334)
);

BUFx2_ASAP7_75t_L g335 ( 
.A(n_23),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g336 ( 
.A(n_96),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_8),
.Y(n_337)
);

BUFx2_ASAP7_75t_L g338 ( 
.A(n_25),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_159),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_83),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_34),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_72),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_30),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_41),
.Y(n_344)
);

CKINVDCx16_ASAP7_75t_R g345 ( 
.A(n_60),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_7),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_14),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_16),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_125),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_33),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_31),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_79),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_250),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_240),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_250),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_304),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_314),
.Y(n_357)
);

NAND2xp33_ASAP7_75t_R g358 ( 
.A(n_276),
.B(n_179),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_250),
.Y(n_359)
);

NOR2xp67_ASAP7_75t_L g360 ( 
.A(n_203),
.B(n_2),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_250),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_250),
.Y(n_362)
);

HB1xp67_ASAP7_75t_L g363 ( 
.A(n_328),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_250),
.Y(n_364)
);

CKINVDCx20_ASAP7_75t_R g365 ( 
.A(n_178),
.Y(n_365)
);

CKINVDCx20_ASAP7_75t_R g366 ( 
.A(n_191),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_334),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_250),
.Y(n_368)
);

CKINVDCx20_ASAP7_75t_R g369 ( 
.A(n_218),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_250),
.Y(n_370)
);

INVxp67_ASAP7_75t_SL g371 ( 
.A(n_204),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_345),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_251),
.Y(n_373)
);

NOR2xp33_ASAP7_75t_L g374 ( 
.A(n_276),
.B(n_3),
.Y(n_374)
);

CKINVDCx20_ASAP7_75t_R g375 ( 
.A(n_261),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_250),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_275),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_321),
.Y(n_378)
);

BUFx3_ASAP7_75t_L g379 ( 
.A(n_252),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_177),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_177),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_180),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_330),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_336),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_180),
.Y(n_385)
);

INVxp67_ASAP7_75t_L g386 ( 
.A(n_328),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_181),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_189),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_189),
.Y(n_389)
);

INVx2_ASAP7_75t_L g390 ( 
.A(n_200),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_200),
.Y(n_391)
);

CKINVDCx20_ASAP7_75t_R g392 ( 
.A(n_281),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_188),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_202),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_202),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_193),
.Y(n_396)
);

INVx1_ASAP7_75t_SL g397 ( 
.A(n_245),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_208),
.Y(n_398)
);

INVxp67_ASAP7_75t_SL g399 ( 
.A(n_204),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_208),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_195),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_210),
.Y(n_402)
);

CKINVDCx20_ASAP7_75t_R g403 ( 
.A(n_228),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_199),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_210),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_205),
.Y(n_406)
);

CKINVDCx20_ASAP7_75t_R g407 ( 
.A(n_238),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_215),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_215),
.Y(n_409)
);

OR2x2_ASAP7_75t_L g410 ( 
.A(n_335),
.B(n_3),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_207),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_219),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_226),
.Y(n_413)
);

CKINVDCx20_ASAP7_75t_R g414 ( 
.A(n_265),
.Y(n_414)
);

CKINVDCx20_ASAP7_75t_R g415 ( 
.A(n_214),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_216),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_216),
.Y(n_417)
);

CKINVDCx20_ASAP7_75t_R g418 ( 
.A(n_214),
.Y(n_418)
);

BUFx2_ASAP7_75t_SL g419 ( 
.A(n_214),
.Y(n_419)
);

INVxp33_ASAP7_75t_L g420 ( 
.A(n_307),
.Y(n_420)
);

INVx2_ASAP7_75t_L g421 ( 
.A(n_220),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_220),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_232),
.Y(n_423)
);

INVxp67_ASAP7_75t_SL g424 ( 
.A(n_323),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_234),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_232),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_235),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_241),
.Y(n_428)
);

INVxp67_ASAP7_75t_SL g429 ( 
.A(n_323),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_246),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_235),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_247),
.Y(n_432)
);

NOR2xp67_ASAP7_75t_L g433 ( 
.A(n_203),
.B(n_6),
.Y(n_433)
);

CKINVDCx20_ASAP7_75t_R g434 ( 
.A(n_252),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_248),
.Y(n_435)
);

BUFx2_ASAP7_75t_L g436 ( 
.A(n_335),
.Y(n_436)
);

INVxp67_ASAP7_75t_SL g437 ( 
.A(n_186),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_259),
.Y(n_438)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_273),
.Y(n_439)
);

CKINVDCx5p33_ASAP7_75t_R g440 ( 
.A(n_280),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_L g441 ( 
.A(n_380),
.B(n_247),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_353),
.Y(n_442)
);

BUFx6f_ASAP7_75t_L g443 ( 
.A(n_353),
.Y(n_443)
);

NAND3xp33_ASAP7_75t_L g444 ( 
.A(n_374),
.B(n_192),
.C(n_186),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_355),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_355),
.Y(n_446)
);

BUFx6f_ASAP7_75t_L g447 ( 
.A(n_359),
.Y(n_447)
);

BUFx6f_ASAP7_75t_L g448 ( 
.A(n_359),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_361),
.Y(n_449)
);

INVx2_ASAP7_75t_L g450 ( 
.A(n_361),
.Y(n_450)
);

BUFx3_ASAP7_75t_L g451 ( 
.A(n_379),
.Y(n_451)
);

INVx3_ASAP7_75t_L g452 ( 
.A(n_390),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_380),
.B(n_260),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_362),
.Y(n_454)
);

INVx2_ASAP7_75t_L g455 ( 
.A(n_362),
.Y(n_455)
);

INVx2_ASAP7_75t_L g456 ( 
.A(n_364),
.Y(n_456)
);

HB1xp67_ASAP7_75t_L g457 ( 
.A(n_397),
.Y(n_457)
);

CKINVDCx5p33_ASAP7_75t_R g458 ( 
.A(n_373),
.Y(n_458)
);

CKINVDCx5p33_ASAP7_75t_R g459 ( 
.A(n_377),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_364),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_368),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_368),
.Y(n_462)
);

NAND2xp33_ASAP7_75t_L g463 ( 
.A(n_387),
.B(n_233),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_370),
.Y(n_464)
);

AND2x2_ASAP7_75t_L g465 ( 
.A(n_381),
.B(n_338),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_370),
.Y(n_466)
);

BUFx6f_ASAP7_75t_L g467 ( 
.A(n_376),
.Y(n_467)
);

AND2x4_ASAP7_75t_L g468 ( 
.A(n_379),
.B(n_233),
.Y(n_468)
);

AND3x2_ASAP7_75t_L g469 ( 
.A(n_436),
.B(n_338),
.C(n_237),
.Y(n_469)
);

AND2x2_ASAP7_75t_L g470 ( 
.A(n_381),
.B(n_303),
.Y(n_470)
);

AND2x4_ASAP7_75t_L g471 ( 
.A(n_382),
.B(n_258),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_376),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_390),
.Y(n_473)
);

BUFx6f_ASAP7_75t_L g474 ( 
.A(n_421),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_421),
.Y(n_475)
);

INVx3_ASAP7_75t_L g476 ( 
.A(n_382),
.Y(n_476)
);

BUFx6f_ASAP7_75t_L g477 ( 
.A(n_385),
.Y(n_477)
);

BUFx6f_ASAP7_75t_L g478 ( 
.A(n_385),
.Y(n_478)
);

INVx2_ASAP7_75t_L g479 ( 
.A(n_388),
.Y(n_479)
);

BUFx6f_ASAP7_75t_L g480 ( 
.A(n_388),
.Y(n_480)
);

INVx2_ASAP7_75t_L g481 ( 
.A(n_389),
.Y(n_481)
);

NAND2x1_ASAP7_75t_L g482 ( 
.A(n_389),
.B(n_326),
.Y(n_482)
);

AND2x2_ASAP7_75t_L g483 ( 
.A(n_391),
.B(n_303),
.Y(n_483)
);

AND2x4_ASAP7_75t_L g484 ( 
.A(n_391),
.B(n_258),
.Y(n_484)
);

AND2x4_ASAP7_75t_L g485 ( 
.A(n_394),
.B(n_262),
.Y(n_485)
);

INVx2_ASAP7_75t_L g486 ( 
.A(n_394),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_395),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_395),
.Y(n_488)
);

OAI22xp5_ASAP7_75t_L g489 ( 
.A1(n_410),
.A2(n_386),
.B1(n_420),
.B2(n_436),
.Y(n_489)
);

BUFx6f_ASAP7_75t_L g490 ( 
.A(n_398),
.Y(n_490)
);

BUFx6f_ASAP7_75t_L g491 ( 
.A(n_398),
.Y(n_491)
);

BUFx6f_ASAP7_75t_L g492 ( 
.A(n_400),
.Y(n_492)
);

INVx2_ASAP7_75t_L g493 ( 
.A(n_400),
.Y(n_493)
);

CKINVDCx5p33_ASAP7_75t_R g494 ( 
.A(n_378),
.Y(n_494)
);

BUFx6f_ASAP7_75t_L g495 ( 
.A(n_402),
.Y(n_495)
);

BUFx6f_ASAP7_75t_L g496 ( 
.A(n_402),
.Y(n_496)
);

HB1xp67_ASAP7_75t_L g497 ( 
.A(n_363),
.Y(n_497)
);

OAI21x1_ASAP7_75t_L g498 ( 
.A1(n_405),
.A2(n_263),
.B(n_260),
.Y(n_498)
);

INVx2_ASAP7_75t_L g499 ( 
.A(n_405),
.Y(n_499)
);

INVx2_ASAP7_75t_L g500 ( 
.A(n_408),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_408),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_409),
.Y(n_502)
);

INVx2_ASAP7_75t_L g503 ( 
.A(n_409),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_416),
.Y(n_504)
);

INVx2_ASAP7_75t_L g505 ( 
.A(n_416),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_L g506 ( 
.A(n_417),
.B(n_422),
.Y(n_506)
);

BUFx6f_ASAP7_75t_L g507 ( 
.A(n_417),
.Y(n_507)
);

AOI22xp5_ASAP7_75t_L g508 ( 
.A1(n_358),
.A2(n_262),
.B1(n_351),
.B2(n_308),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_422),
.Y(n_509)
);

CKINVDCx8_ASAP7_75t_R g510 ( 
.A(n_357),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_423),
.Y(n_511)
);

AND2x4_ASAP7_75t_L g512 ( 
.A(n_423),
.B(n_316),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_426),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_426),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_427),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_427),
.Y(n_516)
);

BUFx6f_ASAP7_75t_L g517 ( 
.A(n_431),
.Y(n_517)
);

INVx2_ASAP7_75t_L g518 ( 
.A(n_450),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_L g519 ( 
.A(n_476),
.B(n_419),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_L g520 ( 
.A(n_476),
.B(n_419),
.Y(n_520)
);

AND2x2_ASAP7_75t_L g521 ( 
.A(n_470),
.B(n_371),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_507),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_L g523 ( 
.A(n_476),
.B(n_431),
.Y(n_523)
);

INVxp67_ASAP7_75t_SL g524 ( 
.A(n_457),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_507),
.Y(n_525)
);

NOR2xp33_ASAP7_75t_L g526 ( 
.A(n_451),
.B(n_393),
.Y(n_526)
);

BUFx6f_ASAP7_75t_SL g527 ( 
.A(n_468),
.Y(n_527)
);

INVx2_ASAP7_75t_L g528 ( 
.A(n_450),
.Y(n_528)
);

NOR2xp33_ASAP7_75t_L g529 ( 
.A(n_451),
.B(n_396),
.Y(n_529)
);

INVx3_ASAP7_75t_L g530 ( 
.A(n_477),
.Y(n_530)
);

OR2x6_ASAP7_75t_L g531 ( 
.A(n_482),
.B(n_410),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_L g532 ( 
.A(n_476),
.B(n_432),
.Y(n_532)
);

NOR2xp33_ASAP7_75t_L g533 ( 
.A(n_463),
.B(n_401),
.Y(n_533)
);

INVx2_ASAP7_75t_L g534 ( 
.A(n_450),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_L g535 ( 
.A(n_487),
.B(n_404),
.Y(n_535)
);

INVx2_ASAP7_75t_L g536 ( 
.A(n_455),
.Y(n_536)
);

INVx2_ASAP7_75t_L g537 ( 
.A(n_455),
.Y(n_537)
);

INVx2_ASAP7_75t_SL g538 ( 
.A(n_457),
.Y(n_538)
);

NOR2xp33_ASAP7_75t_L g539 ( 
.A(n_508),
.B(n_406),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_L g540 ( 
.A(n_487),
.B(n_411),
.Y(n_540)
);

BUFx6f_ASAP7_75t_L g541 ( 
.A(n_474),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_SL g542 ( 
.A(n_508),
.B(n_412),
.Y(n_542)
);

AOI22xp33_ASAP7_75t_L g543 ( 
.A1(n_444),
.A2(n_360),
.B1(n_433),
.B2(n_434),
.Y(n_543)
);

AND3x2_ASAP7_75t_L g544 ( 
.A(n_497),
.B(n_198),
.C(n_192),
.Y(n_544)
);

INVx2_ASAP7_75t_SL g545 ( 
.A(n_471),
.Y(n_545)
);

INVx3_ASAP7_75t_L g546 ( 
.A(n_477),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_507),
.Y(n_547)
);

AOI22xp33_ASAP7_75t_L g548 ( 
.A1(n_444),
.A2(n_360),
.B1(n_433),
.B2(n_316),
.Y(n_548)
);

BUFx3_ASAP7_75t_L g549 ( 
.A(n_442),
.Y(n_549)
);

INVx2_ASAP7_75t_L g550 ( 
.A(n_455),
.Y(n_550)
);

OAI22xp33_ASAP7_75t_L g551 ( 
.A1(n_489),
.A2(n_372),
.B1(n_367),
.B2(n_438),
.Y(n_551)
);

BUFx4f_ASAP7_75t_L g552 ( 
.A(n_477),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_507),
.Y(n_553)
);

AND2x2_ASAP7_75t_L g554 ( 
.A(n_470),
.B(n_399),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_507),
.Y(n_555)
);

AOI22xp33_ASAP7_75t_L g556 ( 
.A1(n_489),
.A2(n_437),
.B1(n_209),
.B2(n_313),
.Y(n_556)
);

INVx2_ASAP7_75t_L g557 ( 
.A(n_456),
.Y(n_557)
);

AND2x2_ASAP7_75t_L g558 ( 
.A(n_470),
.B(n_424),
.Y(n_558)
);

NAND3xp33_ASAP7_75t_L g559 ( 
.A(n_477),
.B(n_266),
.C(n_263),
.Y(n_559)
);

INVx2_ASAP7_75t_L g560 ( 
.A(n_456),
.Y(n_560)
);

AND2x2_ASAP7_75t_SL g561 ( 
.A(n_471),
.B(n_184),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_507),
.Y(n_562)
);

INVx2_ASAP7_75t_L g563 ( 
.A(n_456),
.Y(n_563)
);

INVx2_ASAP7_75t_L g564 ( 
.A(n_443),
.Y(n_564)
);

INVx2_ASAP7_75t_L g565 ( 
.A(n_443),
.Y(n_565)
);

OR2x2_ASAP7_75t_L g566 ( 
.A(n_497),
.B(n_383),
.Y(n_566)
);

NOR2xp33_ASAP7_75t_L g567 ( 
.A(n_488),
.B(n_413),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_507),
.Y(n_568)
);

BUFx6f_ASAP7_75t_L g569 ( 
.A(n_474),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_L g570 ( 
.A(n_488),
.B(n_425),
.Y(n_570)
);

NAND3xp33_ASAP7_75t_L g571 ( 
.A(n_477),
.B(n_268),
.C(n_266),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_517),
.Y(n_572)
);

NOR2xp33_ASAP7_75t_L g573 ( 
.A(n_501),
.B(n_428),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_517),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_517),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_517),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_517),
.Y(n_577)
);

INVx2_ASAP7_75t_L g578 ( 
.A(n_443),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_517),
.Y(n_579)
);

INVx3_ASAP7_75t_L g580 ( 
.A(n_477),
.Y(n_580)
);

INVx2_ASAP7_75t_L g581 ( 
.A(n_443),
.Y(n_581)
);

INVx2_ASAP7_75t_L g582 ( 
.A(n_443),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_517),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_478),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_478),
.Y(n_585)
);

INVx2_ASAP7_75t_L g586 ( 
.A(n_443),
.Y(n_586)
);

INVx2_ASAP7_75t_L g587 ( 
.A(n_447),
.Y(n_587)
);

CKINVDCx5p33_ASAP7_75t_R g588 ( 
.A(n_458),
.Y(n_588)
);

BUFx3_ASAP7_75t_L g589 ( 
.A(n_442),
.Y(n_589)
);

AOI22xp5_ASAP7_75t_L g590 ( 
.A1(n_465),
.A2(n_300),
.B1(n_284),
.B2(n_287),
.Y(n_590)
);

BUFx6f_ASAP7_75t_L g591 ( 
.A(n_474),
.Y(n_591)
);

INVx3_ASAP7_75t_L g592 ( 
.A(n_478),
.Y(n_592)
);

INVxp67_ASAP7_75t_L g593 ( 
.A(n_459),
.Y(n_593)
);

INVx1_ASAP7_75t_SL g594 ( 
.A(n_494),
.Y(n_594)
);

BUFx10_ASAP7_75t_L g595 ( 
.A(n_468),
.Y(n_595)
);

BUFx3_ASAP7_75t_L g596 ( 
.A(n_445),
.Y(n_596)
);

INVxp67_ASAP7_75t_SL g597 ( 
.A(n_506),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_478),
.Y(n_598)
);

INVx3_ASAP7_75t_L g599 ( 
.A(n_478),
.Y(n_599)
);

BUFx6f_ASAP7_75t_L g600 ( 
.A(n_474),
.Y(n_600)
);

BUFx3_ASAP7_75t_L g601 ( 
.A(n_445),
.Y(n_601)
);

INVx2_ASAP7_75t_SL g602 ( 
.A(n_471),
.Y(n_602)
);

INVx4_ASAP7_75t_L g603 ( 
.A(n_478),
.Y(n_603)
);

INVx1_ASAP7_75t_SL g604 ( 
.A(n_465),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_480),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_L g606 ( 
.A(n_501),
.B(n_430),
.Y(n_606)
);

INVx2_ASAP7_75t_L g607 ( 
.A(n_447),
.Y(n_607)
);

NOR2xp33_ASAP7_75t_L g608 ( 
.A(n_502),
.B(n_435),
.Y(n_608)
);

AND2x4_ASAP7_75t_L g609 ( 
.A(n_471),
.B(n_429),
.Y(n_609)
);

AOI22xp33_ASAP7_75t_L g610 ( 
.A1(n_484),
.A2(n_288),
.B1(n_198),
.B2(n_256),
.Y(n_610)
);

BUFx3_ASAP7_75t_L g611 ( 
.A(n_446),
.Y(n_611)
);

INVx2_ASAP7_75t_L g612 ( 
.A(n_447),
.Y(n_612)
);

AOI22xp5_ASAP7_75t_L g613 ( 
.A1(n_465),
.A2(n_485),
.B1(n_484),
.B2(n_290),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_SL g614 ( 
.A(n_468),
.B(n_439),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_480),
.Y(n_615)
);

CKINVDCx5p33_ASAP7_75t_R g616 ( 
.A(n_510),
.Y(n_616)
);

OAI22xp33_ASAP7_75t_L g617 ( 
.A1(n_441),
.A2(n_440),
.B1(n_403),
.B2(n_407),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_480),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_L g619 ( 
.A(n_502),
.B(n_236),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_SL g620 ( 
.A(n_468),
.B(n_484),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_L g621 ( 
.A(n_504),
.B(n_253),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_SL g622 ( 
.A(n_484),
.B(n_384),
.Y(n_622)
);

BUFx10_ASAP7_75t_L g623 ( 
.A(n_469),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_480),
.Y(n_624)
);

OAI22xp33_ASAP7_75t_L g625 ( 
.A1(n_441),
.A2(n_414),
.B1(n_289),
.B2(n_318),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_480),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_480),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_490),
.Y(n_628)
);

INVx2_ASAP7_75t_L g629 ( 
.A(n_447),
.Y(n_629)
);

INVx2_ASAP7_75t_L g630 ( 
.A(n_447),
.Y(n_630)
);

INVx2_ASAP7_75t_L g631 ( 
.A(n_447),
.Y(n_631)
);

NOR2xp33_ASAP7_75t_L g632 ( 
.A(n_504),
.B(n_415),
.Y(n_632)
);

NOR2xp33_ASAP7_75t_L g633 ( 
.A(n_509),
.B(n_418),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_SL g634 ( 
.A(n_485),
.B(n_291),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_490),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_490),
.Y(n_636)
);

NOR2xp33_ASAP7_75t_L g637 ( 
.A(n_509),
.B(n_511),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_SL g638 ( 
.A(n_485),
.B(n_296),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_490),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_490),
.Y(n_640)
);

NAND3xp33_ASAP7_75t_L g641 ( 
.A(n_490),
.B(n_285),
.C(n_268),
.Y(n_641)
);

INVx2_ASAP7_75t_L g642 ( 
.A(n_448),
.Y(n_642)
);

INVx3_ASAP7_75t_L g643 ( 
.A(n_491),
.Y(n_643)
);

INVx2_ASAP7_75t_L g644 ( 
.A(n_448),
.Y(n_644)
);

INVx3_ASAP7_75t_L g645 ( 
.A(n_491),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_491),
.Y(n_646)
);

AND2x6_ASAP7_75t_L g647 ( 
.A(n_479),
.B(n_285),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_L g648 ( 
.A(n_511),
.B(n_295),
.Y(n_648)
);

NOR2xp33_ASAP7_75t_L g649 ( 
.A(n_513),
.B(n_365),
.Y(n_649)
);

AND2x6_ASAP7_75t_L g650 ( 
.A(n_479),
.B(n_295),
.Y(n_650)
);

NOR2xp33_ASAP7_75t_L g651 ( 
.A(n_513),
.B(n_366),
.Y(n_651)
);

BUFx6f_ASAP7_75t_L g652 ( 
.A(n_474),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_SL g653 ( 
.A(n_485),
.B(n_306),
.Y(n_653)
);

INVx5_ASAP7_75t_L g654 ( 
.A(n_448),
.Y(n_654)
);

HB1xp67_ASAP7_75t_L g655 ( 
.A(n_483),
.Y(n_655)
);

NAND2xp33_ASAP7_75t_L g656 ( 
.A(n_491),
.B(n_182),
.Y(n_656)
);

INVx2_ASAP7_75t_L g657 ( 
.A(n_448),
.Y(n_657)
);

INVx2_ASAP7_75t_L g658 ( 
.A(n_448),
.Y(n_658)
);

INVx3_ASAP7_75t_L g659 ( 
.A(n_491),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_SL g660 ( 
.A(n_510),
.B(n_309),
.Y(n_660)
);

OR2x2_ASAP7_75t_L g661 ( 
.A(n_506),
.B(n_354),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_SL g662 ( 
.A(n_510),
.B(n_312),
.Y(n_662)
);

INVx2_ASAP7_75t_L g663 ( 
.A(n_448),
.Y(n_663)
);

INVx5_ASAP7_75t_L g664 ( 
.A(n_467),
.Y(n_664)
);

INVxp67_ASAP7_75t_SL g665 ( 
.A(n_491),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_L g666 ( 
.A(n_514),
.B(n_297),
.Y(n_666)
);

INVx2_ASAP7_75t_L g667 ( 
.A(n_467),
.Y(n_667)
);

INVx1_ASAP7_75t_SL g668 ( 
.A(n_469),
.Y(n_668)
);

INVx2_ASAP7_75t_SL g669 ( 
.A(n_482),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_L g670 ( 
.A(n_597),
.B(n_514),
.Y(n_670)
);

OR2x2_ASAP7_75t_L g671 ( 
.A(n_538),
.B(n_356),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_L g672 ( 
.A(n_545),
.B(n_515),
.Y(n_672)
);

NOR2xp33_ASAP7_75t_R g673 ( 
.A(n_616),
.B(n_369),
.Y(n_673)
);

NOR2xp67_ASAP7_75t_SL g674 ( 
.A(n_545),
.B(n_185),
.Y(n_674)
);

AND2x2_ASAP7_75t_L g675 ( 
.A(n_538),
.B(n_483),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_SL g676 ( 
.A(n_561),
.B(n_446),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_SL g677 ( 
.A(n_561),
.B(n_449),
.Y(n_677)
);

INVx2_ASAP7_75t_SL g678 ( 
.A(n_566),
.Y(n_678)
);

AND2x4_ASAP7_75t_L g679 ( 
.A(n_521),
.B(n_554),
.Y(n_679)
);

A2O1A1Ixp33_ASAP7_75t_L g680 ( 
.A1(n_539),
.A2(n_498),
.B(n_453),
.C(n_505),
.Y(n_680)
);

AND2x6_ASAP7_75t_SL g681 ( 
.A(n_533),
.B(n_201),
.Y(n_681)
);

NAND3xp33_ASAP7_75t_L g682 ( 
.A(n_567),
.B(n_495),
.C(n_492),
.Y(n_682)
);

AND2x2_ASAP7_75t_L g683 ( 
.A(n_524),
.B(n_483),
.Y(n_683)
);

INVxp67_ASAP7_75t_L g684 ( 
.A(n_632),
.Y(n_684)
);

INVx2_ASAP7_75t_L g685 ( 
.A(n_518),
.Y(n_685)
);

AOI22xp33_ASAP7_75t_L g686 ( 
.A1(n_561),
.A2(n_475),
.B1(n_473),
.B2(n_512),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_L g687 ( 
.A(n_602),
.B(n_516),
.Y(n_687)
);

INVxp67_ASAP7_75t_SL g688 ( 
.A(n_549),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_L g689 ( 
.A(n_573),
.B(n_516),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_L g690 ( 
.A(n_608),
.B(n_609),
.Y(n_690)
);

AND2x4_ASAP7_75t_L g691 ( 
.A(n_531),
.B(n_512),
.Y(n_691)
);

OAI22xp5_ASAP7_75t_SL g692 ( 
.A1(n_616),
.A2(n_392),
.B1(n_375),
.B2(n_317),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_549),
.Y(n_693)
);

NOR2x1_ASAP7_75t_L g694 ( 
.A(n_661),
.B(n_453),
.Y(n_694)
);

NAND2xp33_ASAP7_75t_L g695 ( 
.A(n_519),
.B(n_492),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_L g696 ( 
.A(n_609),
.B(n_492),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_589),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_589),
.Y(n_698)
);

NOR2xp33_ASAP7_75t_L g699 ( 
.A(n_535),
.B(n_449),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_SL g700 ( 
.A(n_669),
.B(n_454),
.Y(n_700)
);

INVx8_ASAP7_75t_L g701 ( 
.A(n_527),
.Y(n_701)
);

INVx2_ASAP7_75t_L g702 ( 
.A(n_518),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_SL g703 ( 
.A(n_669),
.B(n_454),
.Y(n_703)
);

OAI22xp5_ASAP7_75t_L g704 ( 
.A1(n_520),
.A2(n_479),
.B1(n_505),
.B2(n_503),
.Y(n_704)
);

OR2x2_ASAP7_75t_L g705 ( 
.A(n_566),
.B(n_512),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_596),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_L g707 ( 
.A(n_609),
.B(n_526),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_L g708 ( 
.A(n_529),
.B(n_492),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_596),
.Y(n_709)
);

INVx2_ASAP7_75t_SL g710 ( 
.A(n_661),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_601),
.Y(n_711)
);

AND2x4_ASAP7_75t_L g712 ( 
.A(n_521),
.B(n_512),
.Y(n_712)
);

INVx2_ASAP7_75t_L g713 ( 
.A(n_528),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_SL g714 ( 
.A(n_601),
.B(n_460),
.Y(n_714)
);

INVx2_ASAP7_75t_L g715 ( 
.A(n_528),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_L g716 ( 
.A(n_540),
.B(n_492),
.Y(n_716)
);

AND2x4_ASAP7_75t_L g717 ( 
.A(n_554),
.B(n_481),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_SL g718 ( 
.A(n_611),
.B(n_460),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_SL g719 ( 
.A(n_611),
.B(n_461),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_L g720 ( 
.A(n_570),
.B(n_495),
.Y(n_720)
);

A2O1A1Ixp33_ASAP7_75t_L g721 ( 
.A1(n_637),
.A2(n_498),
.B(n_503),
.C(n_500),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_L g722 ( 
.A(n_606),
.B(n_495),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_L g723 ( 
.A(n_619),
.B(n_495),
.Y(n_723)
);

INVxp67_ASAP7_75t_SL g724 ( 
.A(n_541),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_SL g725 ( 
.A(n_595),
.B(n_461),
.Y(n_725)
);

AOI22xp5_ASAP7_75t_L g726 ( 
.A1(n_531),
.A2(n_505),
.B1(n_503),
.B2(n_500),
.Y(n_726)
);

NAND3xp33_ASAP7_75t_L g727 ( 
.A(n_633),
.B(n_496),
.C(n_495),
.Y(n_727)
);

NAND2x1p5_ASAP7_75t_L g728 ( 
.A(n_558),
.B(n_452),
.Y(n_728)
);

NOR2xp33_ASAP7_75t_L g729 ( 
.A(n_542),
.B(n_462),
.Y(n_729)
);

AND2x2_ASAP7_75t_L g730 ( 
.A(n_604),
.B(n_594),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_L g731 ( 
.A(n_621),
.B(n_495),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_SL g732 ( 
.A(n_595),
.B(n_462),
.Y(n_732)
);

A2O1A1Ixp33_ASAP7_75t_L g733 ( 
.A1(n_556),
.A2(n_498),
.B(n_499),
.C(n_500),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_L g734 ( 
.A(n_558),
.B(n_496),
.Y(n_734)
);

INVx3_ASAP7_75t_L g735 ( 
.A(n_530),
.Y(n_735)
);

INVx2_ASAP7_75t_L g736 ( 
.A(n_534),
.Y(n_736)
);

INVxp67_ASAP7_75t_L g737 ( 
.A(n_649),
.Y(n_737)
);

NOR2xp33_ASAP7_75t_L g738 ( 
.A(n_655),
.B(n_464),
.Y(n_738)
);

A2O1A1Ixp33_ASAP7_75t_L g739 ( 
.A1(n_613),
.A2(n_499),
.B(n_493),
.C(n_486),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_523),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_L g741 ( 
.A(n_620),
.B(n_496),
.Y(n_741)
);

NOR2xp33_ASAP7_75t_L g742 ( 
.A(n_614),
.B(n_464),
.Y(n_742)
);

OR2x2_ASAP7_75t_L g743 ( 
.A(n_588),
.B(n_452),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_L g744 ( 
.A(n_532),
.B(n_496),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_L g745 ( 
.A(n_613),
.B(n_496),
.Y(n_745)
);

A2O1A1Ixp33_ASAP7_75t_L g746 ( 
.A1(n_590),
.A2(n_651),
.B(n_481),
.C(n_493),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_L g747 ( 
.A(n_548),
.B(n_481),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_L g748 ( 
.A(n_543),
.B(n_595),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_534),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_SL g750 ( 
.A(n_595),
.B(n_552),
.Y(n_750)
);

NOR2x1p5_ASAP7_75t_L g751 ( 
.A(n_588),
.B(n_324),
.Y(n_751)
);

NAND3xp33_ASAP7_75t_L g752 ( 
.A(n_590),
.B(n_472),
.C(n_466),
.Y(n_752)
);

INVx2_ASAP7_75t_L g753 ( 
.A(n_536),
.Y(n_753)
);

OAI21xp5_ASAP7_75t_L g754 ( 
.A1(n_536),
.A2(n_472),
.B(n_466),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_L g755 ( 
.A(n_537),
.B(n_550),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_L g756 ( 
.A(n_537),
.B(n_486),
.Y(n_756)
);

O2A1O1Ixp33_ASAP7_75t_L g757 ( 
.A1(n_648),
.A2(n_666),
.B(n_638),
.C(n_653),
.Y(n_757)
);

OR2x6_ASAP7_75t_L g758 ( 
.A(n_593),
.B(n_185),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_557),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_SL g760 ( 
.A(n_552),
.B(n_467),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_557),
.Y(n_761)
);

AOI22xp33_ASAP7_75t_L g762 ( 
.A1(n_647),
.A2(n_475),
.B1(n_473),
.B2(n_474),
.Y(n_762)
);

AOI21xp5_ASAP7_75t_L g763 ( 
.A1(n_665),
.A2(n_467),
.B(n_486),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_L g764 ( 
.A(n_560),
.B(n_493),
.Y(n_764)
);

AND2x2_ASAP7_75t_L g765 ( 
.A(n_668),
.B(n_623),
.Y(n_765)
);

INVx2_ASAP7_75t_L g766 ( 
.A(n_560),
.Y(n_766)
);

CKINVDCx5p33_ASAP7_75t_R g767 ( 
.A(n_623),
.Y(n_767)
);

NOR2xp33_ASAP7_75t_L g768 ( 
.A(n_634),
.B(n_499),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_SL g769 ( 
.A(n_552),
.B(n_467),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_563),
.Y(n_770)
);

AND2x2_ASAP7_75t_L g771 ( 
.A(n_623),
.B(n_452),
.Y(n_771)
);

AOI22xp5_ASAP7_75t_L g772 ( 
.A1(n_531),
.A2(n_452),
.B1(n_297),
.B2(n_352),
.Y(n_772)
);

AND2x4_ASAP7_75t_L g773 ( 
.A(n_531),
.B(n_201),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_L g774 ( 
.A(n_531),
.B(n_301),
.Y(n_774)
);

BUFx3_ASAP7_75t_L g775 ( 
.A(n_530),
.Y(n_775)
);

AOI22xp5_ASAP7_75t_L g776 ( 
.A1(n_527),
.A2(n_622),
.B1(n_551),
.B2(n_625),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_SL g777 ( 
.A(n_603),
.B(n_301),
.Y(n_777)
);

NAND3xp33_ASAP7_75t_L g778 ( 
.A(n_610),
.B(n_329),
.C(n_325),
.Y(n_778)
);

AND2x2_ASAP7_75t_L g779 ( 
.A(n_623),
.B(n_293),
.Y(n_779)
);

NOR2xp33_ASAP7_75t_L g780 ( 
.A(n_527),
.B(n_331),
.Y(n_780)
);

NOR2x1p5_ASAP7_75t_L g781 ( 
.A(n_617),
.B(n_332),
.Y(n_781)
);

INVx2_ASAP7_75t_L g782 ( 
.A(n_564),
.Y(n_782)
);

INVx2_ASAP7_75t_SL g783 ( 
.A(n_544),
.Y(n_783)
);

INVx1_ASAP7_75t_L g784 ( 
.A(n_584),
.Y(n_784)
);

AND2x2_ASAP7_75t_L g785 ( 
.A(n_660),
.B(n_293),
.Y(n_785)
);

INVxp67_ASAP7_75t_L g786 ( 
.A(n_662),
.Y(n_786)
);

INVx2_ASAP7_75t_L g787 ( 
.A(n_564),
.Y(n_787)
);

NAND2x1p5_ASAP7_75t_L g788 ( 
.A(n_603),
.B(n_311),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_L g789 ( 
.A(n_530),
.B(n_311),
.Y(n_789)
);

AND2x4_ASAP7_75t_L g790 ( 
.A(n_603),
.B(n_209),
.Y(n_790)
);

INVx2_ASAP7_75t_SL g791 ( 
.A(n_546),
.Y(n_791)
);

BUFx3_ASAP7_75t_L g792 ( 
.A(n_546),
.Y(n_792)
);

NAND3xp33_ASAP7_75t_L g793 ( 
.A(n_584),
.B(n_346),
.C(n_337),
.Y(n_793)
);

INVx2_ASAP7_75t_SL g794 ( 
.A(n_546),
.Y(n_794)
);

INVx2_ASAP7_75t_L g795 ( 
.A(n_565),
.Y(n_795)
);

INVxp67_ASAP7_75t_L g796 ( 
.A(n_647),
.Y(n_796)
);

INVx2_ASAP7_75t_L g797 ( 
.A(n_565),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_SL g798 ( 
.A(n_654),
.B(n_322),
.Y(n_798)
);

NAND2xp33_ASAP7_75t_L g799 ( 
.A(n_522),
.B(n_343),
.Y(n_799)
);

INVx2_ASAP7_75t_L g800 ( 
.A(n_578),
.Y(n_800)
);

INVx3_ASAP7_75t_L g801 ( 
.A(n_580),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_585),
.Y(n_802)
);

AOI22xp5_ASAP7_75t_L g803 ( 
.A1(n_585),
.A2(n_352),
.B1(n_339),
.B2(n_322),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_SL g804 ( 
.A(n_654),
.B(n_664),
.Y(n_804)
);

AND2x2_ASAP7_75t_L g805 ( 
.A(n_580),
.B(n_293),
.Y(n_805)
);

CKINVDCx5p33_ASAP7_75t_R g806 ( 
.A(n_647),
.Y(n_806)
);

INVx2_ASAP7_75t_L g807 ( 
.A(n_578),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_L g808 ( 
.A(n_580),
.B(n_339),
.Y(n_808)
);

AOI22xp5_ASAP7_75t_L g809 ( 
.A1(n_598),
.A2(n_206),
.B1(n_349),
.B2(n_183),
.Y(n_809)
);

INVx2_ASAP7_75t_L g810 ( 
.A(n_581),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_L g811 ( 
.A(n_592),
.B(n_211),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_L g812 ( 
.A(n_592),
.B(n_211),
.Y(n_812)
);

NOR2xp33_ASAP7_75t_SL g813 ( 
.A(n_559),
.B(n_344),
.Y(n_813)
);

INVx3_ASAP7_75t_L g814 ( 
.A(n_592),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_L g815 ( 
.A(n_599),
.B(n_213),
.Y(n_815)
);

INVx2_ASAP7_75t_L g816 ( 
.A(n_582),
.Y(n_816)
);

INVx2_ASAP7_75t_L g817 ( 
.A(n_582),
.Y(n_817)
);

INVx2_ASAP7_75t_SL g818 ( 
.A(n_599),
.Y(n_818)
);

A2O1A1Ixp33_ASAP7_75t_L g819 ( 
.A1(n_571),
.A2(n_350),
.B(n_348),
.C(n_213),
.Y(n_819)
);

CKINVDCx5p33_ASAP7_75t_R g820 ( 
.A(n_647),
.Y(n_820)
);

INVx1_ASAP7_75t_L g821 ( 
.A(n_598),
.Y(n_821)
);

AND2x4_ASAP7_75t_L g822 ( 
.A(n_599),
.B(n_643),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_SL g823 ( 
.A(n_654),
.B(n_184),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_L g824 ( 
.A(n_643),
.B(n_256),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_L g825 ( 
.A(n_643),
.B(n_271),
.Y(n_825)
);

INVx2_ASAP7_75t_L g826 ( 
.A(n_586),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_L g827 ( 
.A(n_645),
.B(n_659),
.Y(n_827)
);

NOR3xp33_ASAP7_75t_L g828 ( 
.A(n_645),
.B(n_239),
.C(n_243),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_L g829 ( 
.A(n_645),
.B(n_271),
.Y(n_829)
);

INVx3_ASAP7_75t_L g830 ( 
.A(n_659),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_SL g831 ( 
.A(n_654),
.B(n_217),
.Y(n_831)
);

NAND2xp33_ASAP7_75t_L g832 ( 
.A(n_522),
.B(n_347),
.Y(n_832)
);

NAND2xp33_ASAP7_75t_L g833 ( 
.A(n_525),
.B(n_272),
.Y(n_833)
);

INVx2_ASAP7_75t_L g834 ( 
.A(n_586),
.Y(n_834)
);

OR2x6_ASAP7_75t_L g835 ( 
.A(n_701),
.B(n_571),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_696),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_L g837 ( 
.A(n_690),
.B(n_605),
.Y(n_837)
);

INVxp67_ASAP7_75t_L g838 ( 
.A(n_730),
.Y(n_838)
);

AO21x1_ASAP7_75t_L g839 ( 
.A1(n_708),
.A2(n_547),
.B(n_525),
.Y(n_839)
);

INVx2_ASAP7_75t_L g840 ( 
.A(n_685),
.Y(n_840)
);

AOI21x1_ASAP7_75t_L g841 ( 
.A1(n_760),
.A2(n_615),
.B(n_605),
.Y(n_841)
);

NOR2xp33_ASAP7_75t_L g842 ( 
.A(n_737),
.B(n_587),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_L g843 ( 
.A(n_689),
.B(n_615),
.Y(n_843)
);

OAI21xp5_ASAP7_75t_L g844 ( 
.A1(n_733),
.A2(n_553),
.B(n_547),
.Y(n_844)
);

NOR2xp33_ASAP7_75t_L g845 ( 
.A(n_684),
.B(n_587),
.Y(n_845)
);

O2A1O1Ixp33_ASAP7_75t_SL g846 ( 
.A1(n_680),
.A2(n_577),
.B(n_553),
.C(n_555),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_L g847 ( 
.A(n_707),
.B(n_618),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_L g848 ( 
.A(n_694),
.B(n_618),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_L g849 ( 
.A(n_699),
.B(n_624),
.Y(n_849)
);

BUFx6f_ASAP7_75t_L g850 ( 
.A(n_701),
.Y(n_850)
);

AOI21xp5_ASAP7_75t_L g851 ( 
.A1(n_716),
.A2(n_612),
.B(n_607),
.Y(n_851)
);

AOI21x1_ASAP7_75t_L g852 ( 
.A1(n_760),
.A2(n_626),
.B(n_624),
.Y(n_852)
);

OAI22xp5_ASAP7_75t_L g853 ( 
.A1(n_699),
.A2(n_577),
.B1(n_555),
.B2(n_562),
.Y(n_853)
);

AOI21xp5_ASAP7_75t_L g854 ( 
.A1(n_720),
.A2(n_612),
.B(n_607),
.Y(n_854)
);

A2O1A1Ixp33_ASAP7_75t_L g855 ( 
.A1(n_729),
.A2(n_640),
.B(n_626),
.C(n_627),
.Y(n_855)
);

NOR3xp33_ASAP7_75t_L g856 ( 
.A(n_710),
.B(n_282),
.C(n_278),
.Y(n_856)
);

OAI21xp5_ASAP7_75t_L g857 ( 
.A1(n_733),
.A2(n_568),
.B(n_562),
.Y(n_857)
);

HB1xp67_ASAP7_75t_L g858 ( 
.A(n_679),
.Y(n_858)
);

INVx6_ASAP7_75t_L g859 ( 
.A(n_701),
.Y(n_859)
);

AOI21xp5_ASAP7_75t_L g860 ( 
.A1(n_722),
.A2(n_630),
.B(n_629),
.Y(n_860)
);

INVx4_ASAP7_75t_L g861 ( 
.A(n_691),
.Y(n_861)
);

OAI22xp5_ASAP7_75t_L g862 ( 
.A1(n_670),
.A2(n_568),
.B1(n_572),
.B2(n_574),
.Y(n_862)
);

AO21x1_ASAP7_75t_L g863 ( 
.A1(n_729),
.A2(n_574),
.B(n_572),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_L g864 ( 
.A(n_717),
.B(n_738),
.Y(n_864)
);

OAI21xp5_ASAP7_75t_L g865 ( 
.A1(n_721),
.A2(n_576),
.B(n_575),
.Y(n_865)
);

INVx2_ASAP7_75t_L g866 ( 
.A(n_702),
.Y(n_866)
);

AOI221xp5_ASAP7_75t_SL g867 ( 
.A1(n_738),
.A2(n_350),
.B1(n_278),
.B2(n_282),
.C(n_288),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_L g868 ( 
.A(n_717),
.B(n_627),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_SL g869 ( 
.A(n_691),
.B(n_541),
.Y(n_869)
);

NAND2xp5_ASAP7_75t_SL g870 ( 
.A(n_691),
.B(n_541),
.Y(n_870)
);

AOI21xp5_ASAP7_75t_L g871 ( 
.A1(n_827),
.A2(n_630),
.B(n_629),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_L g872 ( 
.A(n_679),
.B(n_628),
.Y(n_872)
);

AOI21xp5_ASAP7_75t_L g873 ( 
.A1(n_744),
.A2(n_642),
.B(n_644),
.Y(n_873)
);

AOI21x1_ASAP7_75t_L g874 ( 
.A1(n_769),
.A2(n_635),
.B(n_640),
.Y(n_874)
);

AOI21xp5_ASAP7_75t_L g875 ( 
.A1(n_695),
.A2(n_667),
.B(n_644),
.Y(n_875)
);

INVx3_ASAP7_75t_L g876 ( 
.A(n_775),
.Y(n_876)
);

AOI21xp5_ASAP7_75t_L g877 ( 
.A1(n_769),
.A2(n_642),
.B(n_631),
.Y(n_877)
);

A2O1A1Ixp33_ASAP7_75t_L g878 ( 
.A1(n_746),
.A2(n_639),
.B(n_628),
.C(n_635),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_L g879 ( 
.A(n_683),
.B(n_636),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_L g880 ( 
.A(n_675),
.B(n_636),
.Y(n_880)
);

AOI21xp5_ASAP7_75t_L g881 ( 
.A1(n_725),
.A2(n_657),
.B(n_631),
.Y(n_881)
);

A2O1A1Ixp33_ASAP7_75t_L g882 ( 
.A1(n_746),
.A2(n_639),
.B(n_646),
.C(n_576),
.Y(n_882)
);

AOI21xp5_ASAP7_75t_L g883 ( 
.A1(n_725),
.A2(n_732),
.B(n_703),
.Y(n_883)
);

BUFx12f_ASAP7_75t_L g884 ( 
.A(n_758),
.Y(n_884)
);

O2A1O1Ixp33_ASAP7_75t_L g885 ( 
.A1(n_739),
.A2(n_341),
.B(n_294),
.C(n_313),
.Y(n_885)
);

AOI22xp33_ASAP7_75t_L g886 ( 
.A1(n_712),
.A2(n_647),
.B1(n_650),
.B2(n_641),
.Y(n_886)
);

HB1xp67_ASAP7_75t_L g887 ( 
.A(n_712),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_SL g888 ( 
.A(n_776),
.B(n_541),
.Y(n_888)
);

NOR2x1_ASAP7_75t_L g889 ( 
.A(n_743),
.B(n_641),
.Y(n_889)
);

AOI21xp5_ASAP7_75t_L g890 ( 
.A1(n_732),
.A2(n_667),
.B(n_663),
.Y(n_890)
);

AOI21xp5_ASAP7_75t_L g891 ( 
.A1(n_700),
.A2(n_663),
.B(n_658),
.Y(n_891)
);

AOI21xp5_ASAP7_75t_L g892 ( 
.A1(n_714),
.A2(n_658),
.B(n_657),
.Y(n_892)
);

AOI21xp5_ASAP7_75t_L g893 ( 
.A1(n_714),
.A2(n_575),
.B(n_579),
.Y(n_893)
);

BUFx6f_ASAP7_75t_L g894 ( 
.A(n_775),
.Y(n_894)
);

AOI21xp5_ASAP7_75t_L g895 ( 
.A1(n_718),
.A2(n_579),
.B(n_583),
.Y(n_895)
);

AND2x4_ASAP7_75t_L g896 ( 
.A(n_765),
.B(n_646),
.Y(n_896)
);

INVx2_ASAP7_75t_SL g897 ( 
.A(n_673),
.Y(n_897)
);

AOI22xp33_ASAP7_75t_L g898 ( 
.A1(n_734),
.A2(n_650),
.B1(n_647),
.B2(n_333),
.Y(n_898)
);

AOI21xp5_ASAP7_75t_L g899 ( 
.A1(n_718),
.A2(n_583),
.B(n_656),
.Y(n_899)
);

INVx1_ASAP7_75t_L g900 ( 
.A(n_811),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_SL g901 ( 
.A(n_678),
.B(n_541),
.Y(n_901)
);

AOI22xp5_ASAP7_75t_L g902 ( 
.A1(n_688),
.A2(n_805),
.B1(n_742),
.B2(n_677),
.Y(n_902)
);

AOI21xp5_ASAP7_75t_L g903 ( 
.A1(n_719),
.A2(n_664),
.B(n_654),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_L g904 ( 
.A(n_740),
.B(n_742),
.Y(n_904)
);

AOI21xp5_ASAP7_75t_L g905 ( 
.A1(n_672),
.A2(n_664),
.B(n_654),
.Y(n_905)
);

AOI21xp5_ASAP7_75t_L g906 ( 
.A1(n_687),
.A2(n_664),
.B(n_652),
.Y(n_906)
);

AOI21xp5_ASAP7_75t_L g907 ( 
.A1(n_763),
.A2(n_664),
.B(n_652),
.Y(n_907)
);

AND2x4_ASAP7_75t_L g908 ( 
.A(n_771),
.B(n_664),
.Y(n_908)
);

NAND2x1p5_ASAP7_75t_L g909 ( 
.A(n_822),
.B(n_569),
.Y(n_909)
);

AOI21xp5_ASAP7_75t_L g910 ( 
.A1(n_723),
.A2(n_652),
.B(n_600),
.Y(n_910)
);

BUFx12f_ASAP7_75t_L g911 ( 
.A(n_758),
.Y(n_911)
);

AND2x2_ASAP7_75t_L g912 ( 
.A(n_705),
.B(n_294),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_L g913 ( 
.A(n_686),
.B(n_647),
.Y(n_913)
);

NOR2xp33_ASAP7_75t_L g914 ( 
.A(n_786),
.B(n_569),
.Y(n_914)
);

INVx5_ASAP7_75t_L g915 ( 
.A(n_773),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_L g916 ( 
.A(n_686),
.B(n_650),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_L g917 ( 
.A(n_728),
.B(n_650),
.Y(n_917)
);

NOR2xp33_ASAP7_75t_L g918 ( 
.A(n_728),
.B(n_569),
.Y(n_918)
);

INVx1_ASAP7_75t_L g919 ( 
.A(n_812),
.Y(n_919)
);

AOI21xp5_ASAP7_75t_L g920 ( 
.A1(n_731),
.A2(n_652),
.B(n_600),
.Y(n_920)
);

NAND2xp5_ASAP7_75t_L g921 ( 
.A(n_773),
.B(n_650),
.Y(n_921)
);

AOI21xp5_ASAP7_75t_L g922 ( 
.A1(n_724),
.A2(n_652),
.B(n_600),
.Y(n_922)
);

NOR2xp33_ASAP7_75t_L g923 ( 
.A(n_693),
.B(n_569),
.Y(n_923)
);

AOI21x1_ASAP7_75t_L g924 ( 
.A1(n_676),
.A2(n_217),
.B(n_292),
.Y(n_924)
);

AOI21xp5_ASAP7_75t_L g925 ( 
.A1(n_750),
.A2(n_569),
.B(n_600),
.Y(n_925)
);

AOI21xp5_ASAP7_75t_L g926 ( 
.A1(n_750),
.A2(n_591),
.B(n_600),
.Y(n_926)
);

NAND2xp5_ASAP7_75t_L g927 ( 
.A(n_773),
.B(n_650),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_L g928 ( 
.A(n_790),
.B(n_650),
.Y(n_928)
);

INVxp67_ASAP7_75t_L g929 ( 
.A(n_774),
.Y(n_929)
);

NOR2xp67_ASAP7_75t_L g930 ( 
.A(n_671),
.B(n_187),
.Y(n_930)
);

AOI21xp5_ASAP7_75t_L g931 ( 
.A1(n_754),
.A2(n_591),
.B(n_269),
.Y(n_931)
);

NAND2xp5_ASAP7_75t_L g932 ( 
.A(n_790),
.B(n_591),
.Y(n_932)
);

AOI21xp5_ASAP7_75t_L g933 ( 
.A1(n_676),
.A2(n_591),
.B(n_267),
.Y(n_933)
);

AND2x2_ASAP7_75t_L g934 ( 
.A(n_779),
.B(n_333),
.Y(n_934)
);

NAND2xp5_ASAP7_75t_L g935 ( 
.A(n_790),
.B(n_591),
.Y(n_935)
);

INVx3_ASAP7_75t_L g936 ( 
.A(n_792),
.Y(n_936)
);

AOI21xp5_ASAP7_75t_L g937 ( 
.A1(n_677),
.A2(n_264),
.B(n_342),
.Y(n_937)
);

NAND2xp5_ASAP7_75t_L g938 ( 
.A(n_768),
.B(n_341),
.Y(n_938)
);

INVx1_ASAP7_75t_L g939 ( 
.A(n_815),
.Y(n_939)
);

AO21x1_ASAP7_75t_L g940 ( 
.A1(n_704),
.A2(n_292),
.B(n_348),
.Y(n_940)
);

NOR2xp33_ASAP7_75t_L g941 ( 
.A(n_697),
.B(n_9),
.Y(n_941)
);

AOI21xp5_ASAP7_75t_L g942 ( 
.A1(n_755),
.A2(n_340),
.B(n_327),
.Y(n_942)
);

INVx2_ASAP7_75t_L g943 ( 
.A(n_713),
.Y(n_943)
);

NAND2x1_ASAP7_75t_L g944 ( 
.A(n_735),
.B(n_801),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_SL g945 ( 
.A(n_726),
.B(n_274),
.Y(n_945)
);

NAND2xp5_ASAP7_75t_L g946 ( 
.A(n_768),
.B(n_190),
.Y(n_946)
);

NAND2xp5_ASAP7_75t_L g947 ( 
.A(n_698),
.B(n_194),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_L g948 ( 
.A(n_706),
.B(n_196),
.Y(n_948)
);

NAND2xp5_ASAP7_75t_SL g949 ( 
.A(n_772),
.B(n_197),
.Y(n_949)
);

O2A1O1Ixp33_ASAP7_75t_L g950 ( 
.A1(n_739),
.A2(n_9),
.B(n_10),
.C(n_11),
.Y(n_950)
);

INVx1_ASAP7_75t_L g951 ( 
.A(n_824),
.Y(n_951)
);

AOI21x1_ASAP7_75t_L g952 ( 
.A1(n_823),
.A2(n_274),
.B(n_310),
.Y(n_952)
);

CKINVDCx10_ASAP7_75t_R g953 ( 
.A(n_758),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_SL g954 ( 
.A(n_709),
.B(n_212),
.Y(n_954)
);

A2O1A1Ixp33_ASAP7_75t_L g955 ( 
.A1(n_757),
.A2(n_320),
.B(n_319),
.C(n_315),
.Y(n_955)
);

AOI22xp5_ASAP7_75t_L g956 ( 
.A1(n_748),
.A2(n_781),
.B1(n_780),
.B2(n_727),
.Y(n_956)
);

INVx2_ASAP7_75t_L g957 ( 
.A(n_715),
.Y(n_957)
);

NOR2xp33_ASAP7_75t_L g958 ( 
.A(n_711),
.B(n_10),
.Y(n_958)
);

NAND2xp5_ASAP7_75t_SL g959 ( 
.A(n_780),
.B(n_221),
.Y(n_959)
);

NOR2xp33_ASAP7_75t_SL g960 ( 
.A(n_692),
.B(n_222),
.Y(n_960)
);

NOR2xp33_ASAP7_75t_L g961 ( 
.A(n_767),
.B(n_12),
.Y(n_961)
);

OAI21xp5_ASAP7_75t_L g962 ( 
.A1(n_721),
.A2(n_255),
.B(n_305),
.Y(n_962)
);

AOI22xp5_ASAP7_75t_L g963 ( 
.A1(n_752),
.A2(n_254),
.B1(n_302),
.B2(n_299),
.Y(n_963)
);

OAI21xp33_ASAP7_75t_L g964 ( 
.A1(n_809),
.A2(n_249),
.B(n_298),
.Y(n_964)
);

NOR2xp67_ASAP7_75t_L g965 ( 
.A(n_783),
.B(n_223),
.Y(n_965)
);

AOI22xp5_ASAP7_75t_L g966 ( 
.A1(n_785),
.A2(n_244),
.B1(n_286),
.B2(n_283),
.Y(n_966)
);

INVx2_ASAP7_75t_L g967 ( 
.A(n_715),
.Y(n_967)
);

AOI21xp5_ASAP7_75t_L g968 ( 
.A1(n_791),
.A2(n_242),
.B(n_279),
.Y(n_968)
);

O2A1O1Ixp33_ASAP7_75t_L g969 ( 
.A1(n_680),
.A2(n_13),
.B(n_14),
.C(n_17),
.Y(n_969)
);

NOR2xp33_ASAP7_75t_L g970 ( 
.A(n_735),
.B(n_21),
.Y(n_970)
);

OAI22xp5_ASAP7_75t_L g971 ( 
.A1(n_745),
.A2(n_231),
.B1(n_277),
.B2(n_225),
.Y(n_971)
);

AOI22xp5_ASAP7_75t_L g972 ( 
.A1(n_806),
.A2(n_230),
.B1(n_227),
.B2(n_270),
.Y(n_972)
);

AOI21xp5_ASAP7_75t_L g973 ( 
.A1(n_794),
.A2(n_257),
.B(n_229),
.Y(n_973)
);

AOI21xp5_ASAP7_75t_L g974 ( 
.A1(n_818),
.A2(n_224),
.B(n_310),
.Y(n_974)
);

INVx2_ASAP7_75t_L g975 ( 
.A(n_736),
.Y(n_975)
);

AOI21xp5_ASAP7_75t_L g976 ( 
.A1(n_756),
.A2(n_310),
.B(n_274),
.Y(n_976)
);

BUFx12f_ASAP7_75t_L g977 ( 
.A(n_681),
.Y(n_977)
);

NAND2xp5_ASAP7_75t_SL g978 ( 
.A(n_820),
.B(n_310),
.Y(n_978)
);

NAND2xp5_ASAP7_75t_L g979 ( 
.A(n_747),
.B(n_21),
.Y(n_979)
);

BUFx2_ASAP7_75t_L g980 ( 
.A(n_673),
.Y(n_980)
);

AOI21xp5_ASAP7_75t_L g981 ( 
.A1(n_764),
.A2(n_310),
.B(n_274),
.Y(n_981)
);

AOI21xp5_ASAP7_75t_L g982 ( 
.A1(n_784),
.A2(n_274),
.B(n_171),
.Y(n_982)
);

A2O1A1Ixp33_ASAP7_75t_L g983 ( 
.A1(n_802),
.A2(n_22),
.B(n_23),
.C(n_24),
.Y(n_983)
);

OAI22xp5_ASAP7_75t_L g984 ( 
.A1(n_821),
.A2(n_22),
.B1(n_25),
.B2(n_26),
.Y(n_984)
);

AOI21xp5_ASAP7_75t_L g985 ( 
.A1(n_822),
.A2(n_65),
.B(n_167),
.Y(n_985)
);

AOI21x1_ASAP7_75t_L g986 ( 
.A1(n_823),
.A2(n_168),
.B(n_160),
.Y(n_986)
);

AND2x2_ASAP7_75t_L g987 ( 
.A(n_751),
.B(n_28),
.Y(n_987)
);

AOI21xp5_ASAP7_75t_L g988 ( 
.A1(n_801),
.A2(n_154),
.B(n_152),
.Y(n_988)
);

NAND2xp5_ASAP7_75t_L g989 ( 
.A(n_788),
.B(n_29),
.Y(n_989)
);

AOI21xp5_ASAP7_75t_L g990 ( 
.A1(n_814),
.A2(n_136),
.B(n_133),
.Y(n_990)
);

AOI21xp5_ASAP7_75t_L g991 ( 
.A1(n_814),
.A2(n_123),
.B(n_119),
.Y(n_991)
);

AND2x2_ASAP7_75t_L g992 ( 
.A(n_828),
.B(n_31),
.Y(n_992)
);

A2O1A1Ixp33_ASAP7_75t_L g993 ( 
.A1(n_741),
.A2(n_33),
.B(n_34),
.C(n_35),
.Y(n_993)
);

AOI21xp5_ASAP7_75t_L g994 ( 
.A1(n_830),
.A2(n_116),
.B(n_110),
.Y(n_994)
);

NAND2xp5_ASAP7_75t_SL g995 ( 
.A(n_788),
.B(n_35),
.Y(n_995)
);

OAI21xp5_ASAP7_75t_L g996 ( 
.A1(n_682),
.A2(n_104),
.B(n_102),
.Y(n_996)
);

AOI21xp5_ASAP7_75t_L g997 ( 
.A1(n_830),
.A2(n_89),
.B(n_88),
.Y(n_997)
);

NAND2xp5_ASAP7_75t_L g998 ( 
.A(n_753),
.B(n_39),
.Y(n_998)
);

AOI21xp5_ASAP7_75t_L g999 ( 
.A1(n_804),
.A2(n_80),
.B(n_69),
.Y(n_999)
);

NOR2xp33_ASAP7_75t_L g1000 ( 
.A(n_778),
.B(n_792),
.Y(n_1000)
);

INVx3_ASAP7_75t_L g1001 ( 
.A(n_782),
.Y(n_1001)
);

AOI21xp5_ASAP7_75t_L g1002 ( 
.A1(n_804),
.A2(n_68),
.B(n_45),
.Y(n_1002)
);

AOI21xp5_ASAP7_75t_L g1003 ( 
.A1(n_782),
.A2(n_62),
.B(n_45),
.Y(n_1003)
);

AOI21xp5_ASAP7_75t_L g1004 ( 
.A1(n_787),
.A2(n_60),
.B(n_46),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_L g1005 ( 
.A(n_753),
.B(n_43),
.Y(n_1005)
);

INVx2_ASAP7_75t_SL g1006 ( 
.A(n_825),
.Y(n_1006)
);

NOR2x1_ASAP7_75t_L g1007 ( 
.A(n_793),
.B(n_46),
.Y(n_1007)
);

NAND2xp5_ASAP7_75t_SL g1008 ( 
.A(n_796),
.B(n_48),
.Y(n_1008)
);

OR2x6_ASAP7_75t_L g1009 ( 
.A(n_777),
.B(n_48),
.Y(n_1009)
);

AOI21xp5_ASAP7_75t_L g1010 ( 
.A1(n_787),
.A2(n_800),
.B(n_826),
.Y(n_1010)
);

NOR2xp33_ASAP7_75t_L g1011 ( 
.A(n_777),
.B(n_49),
.Y(n_1011)
);

BUFx2_ASAP7_75t_L g1012 ( 
.A(n_803),
.Y(n_1012)
);

INVx1_ASAP7_75t_L g1013 ( 
.A(n_829),
.Y(n_1013)
);

AOI21xp5_ASAP7_75t_L g1014 ( 
.A1(n_795),
.A2(n_800),
.B(n_826),
.Y(n_1014)
);

INVx3_ASAP7_75t_L g1015 ( 
.A(n_795),
.Y(n_1015)
);

BUFx3_ASAP7_75t_L g1016 ( 
.A(n_797),
.Y(n_1016)
);

INVx2_ASAP7_75t_L g1017 ( 
.A(n_766),
.Y(n_1017)
);

NAND2xp5_ASAP7_75t_L g1018 ( 
.A(n_864),
.B(n_770),
.Y(n_1018)
);

AOI22xp5_ASAP7_75t_L g1019 ( 
.A1(n_1012),
.A2(n_813),
.B1(n_833),
.B2(n_799),
.Y(n_1019)
);

INVx1_ASAP7_75t_SL g1020 ( 
.A(n_980),
.Y(n_1020)
);

INVx1_ASAP7_75t_L g1021 ( 
.A(n_858),
.Y(n_1021)
);

NAND2xp5_ASAP7_75t_L g1022 ( 
.A(n_904),
.B(n_761),
.Y(n_1022)
);

NOR2xp33_ASAP7_75t_L g1023 ( 
.A(n_838),
.B(n_807),
.Y(n_1023)
);

INVx4_ASAP7_75t_L g1024 ( 
.A(n_915),
.Y(n_1024)
);

CKINVDCx5p33_ASAP7_75t_R g1025 ( 
.A(n_953),
.Y(n_1025)
);

NOR2xp33_ASAP7_75t_L g1026 ( 
.A(n_838),
.B(n_929),
.Y(n_1026)
);

OAI21x1_ASAP7_75t_L g1027 ( 
.A1(n_844),
.A2(n_857),
.B(n_865),
.Y(n_1027)
);

AOI21xp5_ASAP7_75t_L g1028 ( 
.A1(n_849),
.A2(n_832),
.B(n_808),
.Y(n_1028)
);

BUFx2_ASAP7_75t_L g1029 ( 
.A(n_897),
.Y(n_1029)
);

AOI21xp5_ASAP7_75t_L g1030 ( 
.A1(n_843),
.A2(n_789),
.B(n_834),
.Y(n_1030)
);

NOR2xp33_ASAP7_75t_L g1031 ( 
.A(n_929),
.B(n_858),
.Y(n_1031)
);

INVx1_ASAP7_75t_L g1032 ( 
.A(n_840),
.Y(n_1032)
);

NAND2xp5_ASAP7_75t_L g1033 ( 
.A(n_887),
.B(n_759),
.Y(n_1033)
);

CKINVDCx5p33_ASAP7_75t_R g1034 ( 
.A(n_884),
.Y(n_1034)
);

BUFx3_ASAP7_75t_L g1035 ( 
.A(n_850),
.Y(n_1035)
);

OAI22xp5_ASAP7_75t_SL g1036 ( 
.A1(n_977),
.A2(n_762),
.B1(n_749),
.B2(n_810),
.Y(n_1036)
);

OAI22xp5_ASAP7_75t_SL g1037 ( 
.A1(n_961),
.A2(n_762),
.B1(n_797),
.B2(n_807),
.Y(n_1037)
);

INVx1_ASAP7_75t_L g1038 ( 
.A(n_866),
.Y(n_1038)
);

BUFx8_ASAP7_75t_SL g1039 ( 
.A(n_911),
.Y(n_1039)
);

AOI21x1_ASAP7_75t_L g1040 ( 
.A1(n_924),
.A2(n_831),
.B(n_798),
.Y(n_1040)
);

BUFx3_ASAP7_75t_L g1041 ( 
.A(n_850),
.Y(n_1041)
);

INVx1_ASAP7_75t_L g1042 ( 
.A(n_943),
.Y(n_1042)
);

NOR2xp33_ASAP7_75t_L g1043 ( 
.A(n_861),
.B(n_817),
.Y(n_1043)
);

OAI21xp33_ASAP7_75t_L g1044 ( 
.A1(n_1011),
.A2(n_674),
.B(n_819),
.Y(n_1044)
);

NAND2xp5_ASAP7_75t_L g1045 ( 
.A(n_934),
.B(n_816),
.Y(n_1045)
);

NAND2xp5_ASAP7_75t_L g1046 ( 
.A(n_912),
.B(n_836),
.Y(n_1046)
);

NOR2xp33_ASAP7_75t_L g1047 ( 
.A(n_861),
.B(n_872),
.Y(n_1047)
);

AOI21xp5_ASAP7_75t_L g1048 ( 
.A1(n_862),
.A2(n_853),
.B(n_871),
.Y(n_1048)
);

OR2x2_ASAP7_75t_L g1049 ( 
.A(n_856),
.B(n_819),
.Y(n_1049)
);

AOI21xp5_ASAP7_75t_L g1050 ( 
.A1(n_910),
.A2(n_798),
.B(n_831),
.Y(n_1050)
);

BUFx2_ASAP7_75t_L g1051 ( 
.A(n_915),
.Y(n_1051)
);

BUFx3_ASAP7_75t_L g1052 ( 
.A(n_850),
.Y(n_1052)
);

CKINVDCx11_ASAP7_75t_R g1053 ( 
.A(n_850),
.Y(n_1053)
);

AOI21xp5_ASAP7_75t_L g1054 ( 
.A1(n_920),
.A2(n_56),
.B(n_57),
.Y(n_1054)
);

AND2x2_ASAP7_75t_L g1055 ( 
.A(n_856),
.B(n_961),
.Y(n_1055)
);

OR2x2_ASAP7_75t_L g1056 ( 
.A(n_938),
.B(n_896),
.Y(n_1056)
);

AOI21xp5_ASAP7_75t_L g1057 ( 
.A1(n_907),
.A2(n_883),
.B(n_925),
.Y(n_1057)
);

INVx4_ASAP7_75t_L g1058 ( 
.A(n_915),
.Y(n_1058)
);

AOI22xp5_ASAP7_75t_L g1059 ( 
.A1(n_960),
.A2(n_1011),
.B1(n_1009),
.B2(n_956),
.Y(n_1059)
);

O2A1O1Ixp5_ASAP7_75t_L g1060 ( 
.A1(n_863),
.A2(n_839),
.B(n_940),
.C(n_962),
.Y(n_1060)
);

NAND2xp5_ASAP7_75t_L g1061 ( 
.A(n_842),
.B(n_845),
.Y(n_1061)
);

AOI21xp5_ASAP7_75t_L g1062 ( 
.A1(n_926),
.A2(n_922),
.B(n_873),
.Y(n_1062)
);

A2O1A1Ixp33_ASAP7_75t_L g1063 ( 
.A1(n_902),
.A2(n_842),
.B(n_845),
.C(n_885),
.Y(n_1063)
);

NOR2xp33_ASAP7_75t_L g1064 ( 
.A(n_896),
.B(n_1006),
.Y(n_1064)
);

O2A1O1Ixp33_ASAP7_75t_L g1065 ( 
.A1(n_969),
.A2(n_993),
.B(n_995),
.C(n_1009),
.Y(n_1065)
);

O2A1O1Ixp33_ASAP7_75t_L g1066 ( 
.A1(n_969),
.A2(n_995),
.B(n_1009),
.C(n_950),
.Y(n_1066)
);

NOR3xp33_ASAP7_75t_SL g1067 ( 
.A(n_984),
.B(n_983),
.C(n_955),
.Y(n_1067)
);

OAI22xp5_ASAP7_75t_L g1068 ( 
.A1(n_879),
.A2(n_915),
.B1(n_880),
.B2(n_847),
.Y(n_1068)
);

NAND2xp5_ASAP7_75t_L g1069 ( 
.A(n_900),
.B(n_919),
.Y(n_1069)
);

AND2x2_ASAP7_75t_L g1070 ( 
.A(n_992),
.B(n_987),
.Y(n_1070)
);

INVx4_ASAP7_75t_L g1071 ( 
.A(n_859),
.Y(n_1071)
);

INVx1_ASAP7_75t_L g1072 ( 
.A(n_957),
.Y(n_1072)
);

AOI22xp5_ASAP7_75t_L g1073 ( 
.A1(n_914),
.A2(n_930),
.B1(n_1000),
.B2(n_958),
.Y(n_1073)
);

OAI22xp33_ASAP7_75t_L g1074 ( 
.A1(n_989),
.A2(n_966),
.B1(n_916),
.B2(n_913),
.Y(n_1074)
);

AOI21xp5_ASAP7_75t_L g1075 ( 
.A1(n_881),
.A2(n_890),
.B(n_854),
.Y(n_1075)
);

NAND2xp5_ASAP7_75t_SL g1076 ( 
.A(n_894),
.B(n_908),
.Y(n_1076)
);

BUFx2_ASAP7_75t_L g1077 ( 
.A(n_835),
.Y(n_1077)
);

INVx8_ASAP7_75t_L g1078 ( 
.A(n_835),
.Y(n_1078)
);

OAI22xp5_ASAP7_75t_L g1079 ( 
.A1(n_932),
.A2(n_935),
.B1(n_837),
.B2(n_889),
.Y(n_1079)
);

NAND2xp5_ASAP7_75t_L g1080 ( 
.A(n_939),
.B(n_951),
.Y(n_1080)
);

AND2x4_ASAP7_75t_L g1081 ( 
.A(n_908),
.B(n_835),
.Y(n_1081)
);

O2A1O1Ixp5_ASAP7_75t_L g1082 ( 
.A1(n_882),
.A2(n_878),
.B(n_1008),
.C(n_979),
.Y(n_1082)
);

NOR2xp33_ASAP7_75t_L g1083 ( 
.A(n_959),
.B(n_1013),
.Y(n_1083)
);

A2O1A1Ixp33_ASAP7_75t_L g1084 ( 
.A1(n_885),
.A2(n_941),
.B(n_958),
.C(n_1000),
.Y(n_1084)
);

O2A1O1Ixp33_ASAP7_75t_L g1085 ( 
.A1(n_950),
.A2(n_941),
.B(n_1008),
.C(n_855),
.Y(n_1085)
);

INVx2_ASAP7_75t_L g1086 ( 
.A(n_967),
.Y(n_1086)
);

AOI21xp5_ASAP7_75t_L g1087 ( 
.A1(n_851),
.A2(n_860),
.B(n_906),
.Y(n_1087)
);

BUFx6f_ASAP7_75t_L g1088 ( 
.A(n_894),
.Y(n_1088)
);

BUFx2_ASAP7_75t_L g1089 ( 
.A(n_859),
.Y(n_1089)
);

NAND2xp5_ASAP7_75t_L g1090 ( 
.A(n_914),
.B(n_946),
.Y(n_1090)
);

BUFx2_ASAP7_75t_L g1091 ( 
.A(n_859),
.Y(n_1091)
);

NOR2xp33_ASAP7_75t_L g1092 ( 
.A(n_848),
.B(n_869),
.Y(n_1092)
);

NAND2xp5_ASAP7_75t_L g1093 ( 
.A(n_868),
.B(n_970),
.Y(n_1093)
);

INVx1_ASAP7_75t_L g1094 ( 
.A(n_975),
.Y(n_1094)
);

OAI22xp5_ASAP7_75t_L g1095 ( 
.A1(n_876),
.A2(n_936),
.B1(n_894),
.B2(n_970),
.Y(n_1095)
);

OAI21xp33_ASAP7_75t_L g1096 ( 
.A1(n_964),
.A2(n_963),
.B(n_972),
.Y(n_1096)
);

AOI21xp5_ASAP7_75t_L g1097 ( 
.A1(n_877),
.A2(n_905),
.B(n_846),
.Y(n_1097)
);

AOI21xp5_ASAP7_75t_L g1098 ( 
.A1(n_899),
.A2(n_895),
.B(n_893),
.Y(n_1098)
);

CKINVDCx16_ASAP7_75t_R g1099 ( 
.A(n_1007),
.Y(n_1099)
);

AND2x2_ASAP7_75t_L g1100 ( 
.A(n_965),
.B(n_867),
.Y(n_1100)
);

NAND3xp33_ASAP7_75t_L g1101 ( 
.A(n_1003),
.B(n_1004),
.C(n_971),
.Y(n_1101)
);

AOI21xp5_ASAP7_75t_L g1102 ( 
.A1(n_891),
.A2(n_892),
.B(n_875),
.Y(n_1102)
);

OAI22xp5_ASAP7_75t_L g1103 ( 
.A1(n_876),
.A2(n_936),
.B1(n_894),
.B2(n_928),
.Y(n_1103)
);

AOI22xp33_ASAP7_75t_L g1104 ( 
.A1(n_1017),
.A2(n_945),
.B1(n_1016),
.B2(n_949),
.Y(n_1104)
);

NAND2xp5_ASAP7_75t_L g1105 ( 
.A(n_870),
.B(n_918),
.Y(n_1105)
);

NAND2xp5_ASAP7_75t_L g1106 ( 
.A(n_918),
.B(n_1015),
.Y(n_1106)
);

NAND2xp5_ASAP7_75t_SL g1107 ( 
.A(n_921),
.B(n_927),
.Y(n_1107)
);

OAI21xp5_ASAP7_75t_L g1108 ( 
.A1(n_923),
.A2(n_1005),
.B(n_998),
.Y(n_1108)
);

NOR3xp33_ASAP7_75t_SL g1109 ( 
.A(n_954),
.B(n_968),
.C(n_973),
.Y(n_1109)
);

NAND2x1p5_ASAP7_75t_L g1110 ( 
.A(n_944),
.B(n_1015),
.Y(n_1110)
);

INVx1_ASAP7_75t_L g1111 ( 
.A(n_1001),
.Y(n_1111)
);

BUFx2_ASAP7_75t_L g1112 ( 
.A(n_909),
.Y(n_1112)
);

OAI21xp5_ASAP7_75t_L g1113 ( 
.A1(n_923),
.A2(n_933),
.B(n_931),
.Y(n_1113)
);

BUFx2_ASAP7_75t_L g1114 ( 
.A(n_909),
.Y(n_1114)
);

AOI21xp5_ASAP7_75t_L g1115 ( 
.A1(n_903),
.A2(n_888),
.B(n_1014),
.Y(n_1115)
);

AOI21xp5_ASAP7_75t_L g1116 ( 
.A1(n_1010),
.A2(n_942),
.B(n_996),
.Y(n_1116)
);

AOI21xp5_ASAP7_75t_L g1117 ( 
.A1(n_945),
.A2(n_901),
.B(n_974),
.Y(n_1117)
);

HB1xp67_ASAP7_75t_L g1118 ( 
.A(n_1001),
.Y(n_1118)
);

AOI21xp5_ASAP7_75t_L g1119 ( 
.A1(n_917),
.A2(n_947),
.B(n_948),
.Y(n_1119)
);

INVx2_ASAP7_75t_L g1120 ( 
.A(n_841),
.Y(n_1120)
);

INVx1_ASAP7_75t_L g1121 ( 
.A(n_852),
.Y(n_1121)
);

NOR2xp33_ASAP7_75t_L g1122 ( 
.A(n_978),
.B(n_937),
.Y(n_1122)
);

CKINVDCx5p33_ASAP7_75t_R g1123 ( 
.A(n_1002),
.Y(n_1123)
);

AND2x2_ASAP7_75t_L g1124 ( 
.A(n_898),
.B(n_886),
.Y(n_1124)
);

O2A1O1Ixp33_ASAP7_75t_L g1125 ( 
.A1(n_982),
.A2(n_985),
.B(n_990),
.C(n_997),
.Y(n_1125)
);

AOI21xp5_ASAP7_75t_L g1126 ( 
.A1(n_988),
.A2(n_994),
.B(n_991),
.Y(n_1126)
);

NAND2xp5_ASAP7_75t_L g1127 ( 
.A(n_898),
.B(n_886),
.Y(n_1127)
);

NAND2xp5_ASAP7_75t_L g1128 ( 
.A(n_874),
.B(n_976),
.Y(n_1128)
);

AND2x2_ASAP7_75t_L g1129 ( 
.A(n_986),
.B(n_999),
.Y(n_1129)
);

INVx1_ASAP7_75t_SL g1130 ( 
.A(n_981),
.Y(n_1130)
);

A2O1A1Ixp33_ASAP7_75t_L g1131 ( 
.A1(n_952),
.A2(n_699),
.B(n_539),
.C(n_729),
.Y(n_1131)
);

NOR2xp33_ASAP7_75t_L g1132 ( 
.A(n_1012),
.B(n_737),
.Y(n_1132)
);

AO21x1_ASAP7_75t_L g1133 ( 
.A1(n_888),
.A2(n_853),
.B(n_979),
.Y(n_1133)
);

BUFx6f_ASAP7_75t_L g1134 ( 
.A(n_850),
.Y(n_1134)
);

AOI21xp5_ASAP7_75t_L g1135 ( 
.A1(n_849),
.A2(n_904),
.B(n_843),
.Y(n_1135)
);

OAI22xp5_ASAP7_75t_L g1136 ( 
.A1(n_864),
.A2(n_690),
.B1(n_707),
.B2(n_689),
.Y(n_1136)
);

AND2x2_ASAP7_75t_L g1137 ( 
.A(n_838),
.B(n_730),
.Y(n_1137)
);

NOR2xp33_ASAP7_75t_L g1138 ( 
.A(n_1012),
.B(n_737),
.Y(n_1138)
);

INVx3_ASAP7_75t_L g1139 ( 
.A(n_861),
.Y(n_1139)
);

NOR2xp67_ASAP7_75t_L g1140 ( 
.A(n_897),
.B(n_593),
.Y(n_1140)
);

O2A1O1Ixp33_ASAP7_75t_L g1141 ( 
.A1(n_904),
.A2(n_684),
.B(n_737),
.C(n_710),
.Y(n_1141)
);

NAND2xp5_ASAP7_75t_SL g1142 ( 
.A(n_915),
.B(n_730),
.Y(n_1142)
);

INVx1_ASAP7_75t_L g1143 ( 
.A(n_858),
.Y(n_1143)
);

INVx3_ASAP7_75t_L g1144 ( 
.A(n_861),
.Y(n_1144)
);

NAND3xp33_ASAP7_75t_SL g1145 ( 
.A(n_961),
.B(n_737),
.C(n_684),
.Y(n_1145)
);

INVx3_ASAP7_75t_L g1146 ( 
.A(n_861),
.Y(n_1146)
);

O2A1O1Ixp33_ASAP7_75t_L g1147 ( 
.A1(n_904),
.A2(n_684),
.B(n_737),
.C(n_710),
.Y(n_1147)
);

A2O1A1Ixp33_ASAP7_75t_SL g1148 ( 
.A1(n_970),
.A2(n_567),
.B(n_608),
.C(n_573),
.Y(n_1148)
);

AOI21xp5_ASAP7_75t_L g1149 ( 
.A1(n_849),
.A2(n_904),
.B(n_843),
.Y(n_1149)
);

AND2x2_ASAP7_75t_L g1150 ( 
.A(n_838),
.B(n_730),
.Y(n_1150)
);

AND2x4_ASAP7_75t_L g1151 ( 
.A(n_861),
.B(n_850),
.Y(n_1151)
);

A2O1A1Ixp33_ASAP7_75t_L g1152 ( 
.A1(n_1011),
.A2(n_699),
.B(n_539),
.C(n_729),
.Y(n_1152)
);

A2O1A1Ixp33_ASAP7_75t_L g1153 ( 
.A1(n_1011),
.A2(n_699),
.B(n_539),
.C(n_729),
.Y(n_1153)
);

AND2x2_ASAP7_75t_L g1154 ( 
.A(n_838),
.B(n_730),
.Y(n_1154)
);

OAI22xp5_ASAP7_75t_L g1155 ( 
.A1(n_864),
.A2(n_690),
.B1(n_707),
.B2(n_689),
.Y(n_1155)
);

AOI21xp5_ASAP7_75t_L g1156 ( 
.A1(n_849),
.A2(n_904),
.B(n_843),
.Y(n_1156)
);

CKINVDCx5p33_ASAP7_75t_R g1157 ( 
.A(n_980),
.Y(n_1157)
);

A2O1A1Ixp33_ASAP7_75t_L g1158 ( 
.A1(n_1011),
.A2(n_699),
.B(n_539),
.C(n_729),
.Y(n_1158)
);

AOI21xp5_ASAP7_75t_L g1159 ( 
.A1(n_849),
.A2(n_904),
.B(n_843),
.Y(n_1159)
);

HB1xp67_ASAP7_75t_L g1160 ( 
.A(n_887),
.Y(n_1160)
);

OR2x2_ASAP7_75t_L g1161 ( 
.A(n_838),
.B(n_538),
.Y(n_1161)
);

OAI22xp5_ASAP7_75t_L g1162 ( 
.A1(n_864),
.A2(n_690),
.B1(n_707),
.B2(n_689),
.Y(n_1162)
);

O2A1O1Ixp33_ASAP7_75t_L g1163 ( 
.A1(n_904),
.A2(n_684),
.B(n_737),
.C(n_710),
.Y(n_1163)
);

OAI21x1_ASAP7_75t_L g1164 ( 
.A1(n_844),
.A2(n_857),
.B(n_865),
.Y(n_1164)
);

O2A1O1Ixp5_ASAP7_75t_L g1165 ( 
.A1(n_863),
.A2(n_839),
.B(n_940),
.C(n_962),
.Y(n_1165)
);

AND2x6_ASAP7_75t_L g1166 ( 
.A(n_850),
.B(n_691),
.Y(n_1166)
);

BUFx2_ASAP7_75t_L g1167 ( 
.A(n_980),
.Y(n_1167)
);

NAND2xp33_ASAP7_75t_SL g1168 ( 
.A(n_861),
.B(n_588),
.Y(n_1168)
);

AND2x2_ASAP7_75t_L g1169 ( 
.A(n_838),
.B(n_730),
.Y(n_1169)
);

AOI21xp5_ASAP7_75t_L g1170 ( 
.A1(n_849),
.A2(n_904),
.B(n_843),
.Y(n_1170)
);

INVx1_ASAP7_75t_L g1171 ( 
.A(n_858),
.Y(n_1171)
);

O2A1O1Ixp33_ASAP7_75t_L g1172 ( 
.A1(n_1152),
.A2(n_1158),
.B(n_1153),
.C(n_1148),
.Y(n_1172)
);

O2A1O1Ixp33_ASAP7_75t_L g1173 ( 
.A1(n_1084),
.A2(n_1145),
.B(n_1055),
.C(n_1163),
.Y(n_1173)
);

AOI21xp5_ASAP7_75t_L g1174 ( 
.A1(n_1135),
.A2(n_1156),
.B(n_1149),
.Y(n_1174)
);

AND2x2_ASAP7_75t_L g1175 ( 
.A(n_1132),
.B(n_1138),
.Y(n_1175)
);

INVx1_ASAP7_75t_SL g1176 ( 
.A(n_1020),
.Y(n_1176)
);

CKINVDCx5p33_ASAP7_75t_R g1177 ( 
.A(n_1025),
.Y(n_1177)
);

INVx2_ASAP7_75t_SL g1178 ( 
.A(n_1157),
.Y(n_1178)
);

OAI21xp5_ASAP7_75t_L g1179 ( 
.A1(n_1060),
.A2(n_1165),
.B(n_1082),
.Y(n_1179)
);

NAND2x1p5_ASAP7_75t_L g1180 ( 
.A(n_1024),
.B(n_1058),
.Y(n_1180)
);

NAND2xp5_ASAP7_75t_L g1181 ( 
.A(n_1132),
.B(n_1138),
.Y(n_1181)
);

AND2x2_ASAP7_75t_L g1182 ( 
.A(n_1137),
.B(n_1150),
.Y(n_1182)
);

INVxp67_ASAP7_75t_L g1183 ( 
.A(n_1154),
.Y(n_1183)
);

INVx1_ASAP7_75t_L g1184 ( 
.A(n_1032),
.Y(n_1184)
);

OAI21xp5_ASAP7_75t_L g1185 ( 
.A1(n_1060),
.A2(n_1165),
.B(n_1082),
.Y(n_1185)
);

OAI21x1_ASAP7_75t_L g1186 ( 
.A1(n_1097),
.A2(n_1115),
.B(n_1102),
.Y(n_1186)
);

OAI21x1_ASAP7_75t_L g1187 ( 
.A1(n_1057),
.A2(n_1062),
.B(n_1087),
.Y(n_1187)
);

BUFx4_ASAP7_75t_R g1188 ( 
.A(n_1039),
.Y(n_1188)
);

BUFx10_ASAP7_75t_L g1189 ( 
.A(n_1026),
.Y(n_1189)
);

NOR2xp67_ASAP7_75t_L g1190 ( 
.A(n_1069),
.B(n_1080),
.Y(n_1190)
);

BUFx6f_ASAP7_75t_L g1191 ( 
.A(n_1053),
.Y(n_1191)
);

AOI21xp5_ASAP7_75t_L g1192 ( 
.A1(n_1159),
.A2(n_1170),
.B(n_1126),
.Y(n_1192)
);

INVxp67_ASAP7_75t_L g1193 ( 
.A(n_1169),
.Y(n_1193)
);

AO32x2_ASAP7_75t_L g1194 ( 
.A1(n_1079),
.A2(n_1068),
.A3(n_1037),
.B1(n_1036),
.B2(n_1155),
.Y(n_1194)
);

NAND2xp5_ASAP7_75t_L g1195 ( 
.A(n_1031),
.B(n_1026),
.Y(n_1195)
);

A2O1A1Ixp33_ASAP7_75t_L g1196 ( 
.A1(n_1059),
.A2(n_1066),
.B(n_1065),
.C(n_1085),
.Y(n_1196)
);

INVxp67_ASAP7_75t_SL g1197 ( 
.A(n_1031),
.Y(n_1197)
);

OAI21xp5_ASAP7_75t_L g1198 ( 
.A1(n_1063),
.A2(n_1027),
.B(n_1164),
.Y(n_1198)
);

AOI21xp5_ASAP7_75t_L g1199 ( 
.A1(n_1048),
.A2(n_1028),
.B(n_1061),
.Y(n_1199)
);

NAND2xp5_ASAP7_75t_SL g1200 ( 
.A(n_1019),
.B(n_1073),
.Y(n_1200)
);

INVx1_ASAP7_75t_L g1201 ( 
.A(n_1038),
.Y(n_1201)
);

AOI21xp5_ASAP7_75t_L g1202 ( 
.A1(n_1125),
.A2(n_1090),
.B(n_1116),
.Y(n_1202)
);

AND2x2_ASAP7_75t_L g1203 ( 
.A(n_1070),
.B(n_1161),
.Y(n_1203)
);

OAI22xp33_ASAP7_75t_L g1204 ( 
.A1(n_1145),
.A2(n_1049),
.B1(n_1127),
.B2(n_1046),
.Y(n_1204)
);

CKINVDCx20_ASAP7_75t_R g1205 ( 
.A(n_1034),
.Y(n_1205)
);

BUFx3_ASAP7_75t_L g1206 ( 
.A(n_1167),
.Y(n_1206)
);

AOI22xp5_ASAP7_75t_L g1207 ( 
.A1(n_1124),
.A2(n_1136),
.B1(n_1162),
.B2(n_1096),
.Y(n_1207)
);

AOI21xp5_ASAP7_75t_L g1208 ( 
.A1(n_1093),
.A2(n_1075),
.B(n_1108),
.Y(n_1208)
);

AOI21xp5_ASAP7_75t_L g1209 ( 
.A1(n_1098),
.A2(n_1119),
.B(n_1131),
.Y(n_1209)
);

O2A1O1Ixp33_ASAP7_75t_SL g1210 ( 
.A1(n_1095),
.A2(n_1074),
.B(n_1022),
.C(n_1141),
.Y(n_1210)
);

OAI21xp5_ASAP7_75t_L g1211 ( 
.A1(n_1030),
.A2(n_1074),
.B(n_1101),
.Y(n_1211)
);

BUFx3_ASAP7_75t_L g1212 ( 
.A(n_1029),
.Y(n_1212)
);

INVxp67_ASAP7_75t_L g1213 ( 
.A(n_1064),
.Y(n_1213)
);

OAI21xp5_ASAP7_75t_SL g1214 ( 
.A1(n_1147),
.A2(n_1044),
.B(n_1083),
.Y(n_1214)
);

BUFx12f_ASAP7_75t_L g1215 ( 
.A(n_1134),
.Y(n_1215)
);

INVx6_ASAP7_75t_L g1216 ( 
.A(n_1071),
.Y(n_1216)
);

AOI21xp5_ASAP7_75t_L g1217 ( 
.A1(n_1113),
.A2(n_1128),
.B(n_1129),
.Y(n_1217)
);

OR2x6_ASAP7_75t_L g1218 ( 
.A(n_1078),
.B(n_1024),
.Y(n_1218)
);

NAND2x1_ASAP7_75t_L g1219 ( 
.A(n_1088),
.B(n_1058),
.Y(n_1219)
);

AOI21xp5_ASAP7_75t_L g1220 ( 
.A1(n_1123),
.A2(n_1133),
.B(n_1050),
.Y(n_1220)
);

AND2x6_ASAP7_75t_L g1221 ( 
.A(n_1081),
.B(n_1151),
.Y(n_1221)
);

AOI21xp5_ASAP7_75t_L g1222 ( 
.A1(n_1117),
.A2(n_1122),
.B(n_1047),
.Y(n_1222)
);

A2O1A1Ixp33_ASAP7_75t_L g1223 ( 
.A1(n_1083),
.A2(n_1067),
.B(n_1092),
.C(n_1047),
.Y(n_1223)
);

AO31x2_ASAP7_75t_L g1224 ( 
.A1(n_1120),
.A2(n_1121),
.A3(n_1122),
.B(n_1094),
.Y(n_1224)
);

INVx2_ASAP7_75t_SL g1225 ( 
.A(n_1035),
.Y(n_1225)
);

AND2x4_ASAP7_75t_L g1226 ( 
.A(n_1071),
.B(n_1166),
.Y(n_1226)
);

BUFx3_ASAP7_75t_L g1227 ( 
.A(n_1089),
.Y(n_1227)
);

AND2x4_ASAP7_75t_L g1228 ( 
.A(n_1166),
.B(n_1052),
.Y(n_1228)
);

OAI22xp5_ASAP7_75t_L g1229 ( 
.A1(n_1056),
.A2(n_1067),
.B1(n_1140),
.B2(n_1146),
.Y(n_1229)
);

OAI22xp5_ASAP7_75t_L g1230 ( 
.A1(n_1139),
.A2(n_1146),
.B1(n_1144),
.B2(n_1092),
.Y(n_1230)
);

AOI21xp5_ASAP7_75t_L g1231 ( 
.A1(n_1130),
.A2(n_1018),
.B(n_1103),
.Y(n_1231)
);

O2A1O1Ixp33_ASAP7_75t_L g1232 ( 
.A1(n_1100),
.A2(n_1160),
.B(n_1054),
.C(n_1107),
.Y(n_1232)
);

OAI22x1_ASAP7_75t_L g1233 ( 
.A1(n_1077),
.A2(n_1142),
.B1(n_1160),
.B2(n_1064),
.Y(n_1233)
);

AND2x2_ASAP7_75t_L g1234 ( 
.A(n_1021),
.B(n_1171),
.Y(n_1234)
);

NAND2xp5_ASAP7_75t_L g1235 ( 
.A(n_1023),
.B(n_1143),
.Y(n_1235)
);

NAND2xp5_ASAP7_75t_L g1236 ( 
.A(n_1023),
.B(n_1045),
.Y(n_1236)
);

AO31x2_ASAP7_75t_L g1237 ( 
.A1(n_1042),
.A2(n_1072),
.A3(n_1106),
.B(n_1111),
.Y(n_1237)
);

BUFx3_ASAP7_75t_L g1238 ( 
.A(n_1091),
.Y(n_1238)
);

AOI21xp5_ASAP7_75t_L g1239 ( 
.A1(n_1043),
.A2(n_1076),
.B(n_1105),
.Y(n_1239)
);

AOI22xp5_ASAP7_75t_L g1240 ( 
.A1(n_1168),
.A2(n_1099),
.B1(n_1043),
.B2(n_1166),
.Y(n_1240)
);

NOR2xp33_ASAP7_75t_L g1241 ( 
.A(n_1139),
.B(n_1144),
.Y(n_1241)
);

AND2x2_ASAP7_75t_L g1242 ( 
.A(n_1112),
.B(n_1114),
.Y(n_1242)
);

OAI21x1_ASAP7_75t_L g1243 ( 
.A1(n_1040),
.A2(n_1110),
.B(n_1104),
.Y(n_1243)
);

OAI21x1_ASAP7_75t_L g1244 ( 
.A1(n_1110),
.A2(n_1104),
.B(n_1033),
.Y(n_1244)
);

A2O1A1Ixp33_ASAP7_75t_L g1245 ( 
.A1(n_1109),
.A2(n_1118),
.B(n_1078),
.C(n_1051),
.Y(n_1245)
);

AOI21x1_ASAP7_75t_L g1246 ( 
.A1(n_1118),
.A2(n_1109),
.B(n_1078),
.Y(n_1246)
);

A2O1A1Ixp33_ASAP7_75t_L g1247 ( 
.A1(n_1041),
.A2(n_1088),
.B(n_1134),
.C(n_1166),
.Y(n_1247)
);

OAI21xp5_ASAP7_75t_L g1248 ( 
.A1(n_1166),
.A2(n_1088),
.B(n_1134),
.Y(n_1248)
);

INVx2_ASAP7_75t_L g1249 ( 
.A(n_1088),
.Y(n_1249)
);

AOI21xp5_ASAP7_75t_L g1250 ( 
.A1(n_1135),
.A2(n_1156),
.B(n_1149),
.Y(n_1250)
);

A2O1A1Ixp33_ASAP7_75t_L g1251 ( 
.A1(n_1152),
.A2(n_1158),
.B(n_1153),
.C(n_1059),
.Y(n_1251)
);

OAI21xp5_ASAP7_75t_L g1252 ( 
.A1(n_1152),
.A2(n_1158),
.B(n_1153),
.Y(n_1252)
);

AOI221xp5_ASAP7_75t_L g1253 ( 
.A1(n_1152),
.A2(n_489),
.B1(n_737),
.B2(n_684),
.C(n_1153),
.Y(n_1253)
);

A2O1A1Ixp33_ASAP7_75t_L g1254 ( 
.A1(n_1152),
.A2(n_1158),
.B(n_1153),
.C(n_1059),
.Y(n_1254)
);

NOR2xp33_ASAP7_75t_SL g1255 ( 
.A(n_1152),
.B(n_1153),
.Y(n_1255)
);

AOI21xp5_ASAP7_75t_L g1256 ( 
.A1(n_1135),
.A2(n_1156),
.B(n_1149),
.Y(n_1256)
);

INVx2_ASAP7_75t_L g1257 ( 
.A(n_1086),
.Y(n_1257)
);

O2A1O1Ixp33_ASAP7_75t_L g1258 ( 
.A1(n_1152),
.A2(n_1158),
.B(n_1153),
.C(n_737),
.Y(n_1258)
);

AOI221xp5_ASAP7_75t_L g1259 ( 
.A1(n_1152),
.A2(n_489),
.B1(n_737),
.B2(n_684),
.C(n_1153),
.Y(n_1259)
);

INVx1_ASAP7_75t_L g1260 ( 
.A(n_1032),
.Y(n_1260)
);

NAND2xp5_ASAP7_75t_L g1261 ( 
.A(n_1132),
.B(n_1138),
.Y(n_1261)
);

AOI22xp33_ASAP7_75t_L g1262 ( 
.A1(n_1055),
.A2(n_649),
.B1(n_651),
.B2(n_539),
.Y(n_1262)
);

NAND2xp5_ASAP7_75t_SL g1263 ( 
.A(n_1132),
.B(n_1138),
.Y(n_1263)
);

INVx1_ASAP7_75t_L g1264 ( 
.A(n_1032),
.Y(n_1264)
);

OAI22xp33_ASAP7_75t_L g1265 ( 
.A1(n_1059),
.A2(n_960),
.B1(n_1055),
.B2(n_737),
.Y(n_1265)
);

INVx3_ASAP7_75t_L g1266 ( 
.A(n_1024),
.Y(n_1266)
);

OAI21x1_ASAP7_75t_L g1267 ( 
.A1(n_1097),
.A2(n_1115),
.B(n_1102),
.Y(n_1267)
);

CKINVDCx5p33_ASAP7_75t_R g1268 ( 
.A(n_1025),
.Y(n_1268)
);

INVx2_ASAP7_75t_L g1269 ( 
.A(n_1086),
.Y(n_1269)
);

OAI22xp5_ASAP7_75t_L g1270 ( 
.A1(n_1152),
.A2(n_1153),
.B1(n_1158),
.B2(n_684),
.Y(n_1270)
);

OR2x6_ASAP7_75t_L g1271 ( 
.A(n_1078),
.B(n_701),
.Y(n_1271)
);

NAND2xp5_ASAP7_75t_SL g1272 ( 
.A(n_1132),
.B(n_1138),
.Y(n_1272)
);

OAI21x1_ASAP7_75t_L g1273 ( 
.A1(n_1097),
.A2(n_1115),
.B(n_1102),
.Y(n_1273)
);

AOI221x1_ASAP7_75t_L g1274 ( 
.A1(n_1152),
.A2(n_1153),
.B1(n_1158),
.B2(n_1084),
.C(n_1044),
.Y(n_1274)
);

NAND2xp5_ASAP7_75t_L g1275 ( 
.A(n_1132),
.B(n_1138),
.Y(n_1275)
);

INVx1_ASAP7_75t_L g1276 ( 
.A(n_1032),
.Y(n_1276)
);

O2A1O1Ixp33_ASAP7_75t_L g1277 ( 
.A1(n_1152),
.A2(n_1158),
.B(n_1153),
.C(n_737),
.Y(n_1277)
);

NAND2xp5_ASAP7_75t_L g1278 ( 
.A(n_1132),
.B(n_1138),
.Y(n_1278)
);

OAI21xp5_ASAP7_75t_L g1279 ( 
.A1(n_1152),
.A2(n_1158),
.B(n_1153),
.Y(n_1279)
);

HB1xp67_ASAP7_75t_L g1280 ( 
.A(n_1160),
.Y(n_1280)
);

AND2x4_ASAP7_75t_L g1281 ( 
.A(n_1081),
.B(n_861),
.Y(n_1281)
);

INVx2_ASAP7_75t_L g1282 ( 
.A(n_1086),
.Y(n_1282)
);

INVx1_ASAP7_75t_L g1283 ( 
.A(n_1032),
.Y(n_1283)
);

O2A1O1Ixp33_ASAP7_75t_SL g1284 ( 
.A1(n_1152),
.A2(n_1153),
.B(n_1158),
.C(n_1148),
.Y(n_1284)
);

AO21x1_ASAP7_75t_L g1285 ( 
.A1(n_1066),
.A2(n_1065),
.B(n_1085),
.Y(n_1285)
);

AO31x2_ASAP7_75t_L g1286 ( 
.A1(n_1133),
.A2(n_839),
.A3(n_863),
.B(n_1120),
.Y(n_1286)
);

OR2x2_ASAP7_75t_L g1287 ( 
.A(n_1132),
.B(n_1138),
.Y(n_1287)
);

OAI21xp5_ASAP7_75t_L g1288 ( 
.A1(n_1152),
.A2(n_1158),
.B(n_1153),
.Y(n_1288)
);

BUFx6f_ASAP7_75t_L g1289 ( 
.A(n_1053),
.Y(n_1289)
);

OAI22xp33_ASAP7_75t_L g1290 ( 
.A1(n_1059),
.A2(n_960),
.B1(n_1055),
.B2(n_737),
.Y(n_1290)
);

OAI21x1_ASAP7_75t_L g1291 ( 
.A1(n_1097),
.A2(n_1115),
.B(n_1102),
.Y(n_1291)
);

O2A1O1Ixp33_ASAP7_75t_SL g1292 ( 
.A1(n_1152),
.A2(n_1153),
.B(n_1158),
.C(n_1148),
.Y(n_1292)
);

O2A1O1Ixp33_ASAP7_75t_L g1293 ( 
.A1(n_1152),
.A2(n_1158),
.B(n_1153),
.C(n_737),
.Y(n_1293)
);

INVx1_ASAP7_75t_L g1294 ( 
.A(n_1032),
.Y(n_1294)
);

AO31x2_ASAP7_75t_L g1295 ( 
.A1(n_1133),
.A2(n_839),
.A3(n_863),
.B(n_1120),
.Y(n_1295)
);

INVx2_ASAP7_75t_L g1296 ( 
.A(n_1086),
.Y(n_1296)
);

NAND2xp5_ASAP7_75t_L g1297 ( 
.A(n_1132),
.B(n_1138),
.Y(n_1297)
);

OAI21x1_ASAP7_75t_L g1298 ( 
.A1(n_1097),
.A2(n_1115),
.B(n_1102),
.Y(n_1298)
);

CKINVDCx12_ASAP7_75t_R g1299 ( 
.A(n_1161),
.Y(n_1299)
);

OAI21x1_ASAP7_75t_L g1300 ( 
.A1(n_1097),
.A2(n_1115),
.B(n_1102),
.Y(n_1300)
);

O2A1O1Ixp33_ASAP7_75t_SL g1301 ( 
.A1(n_1152),
.A2(n_1153),
.B(n_1158),
.C(n_1148),
.Y(n_1301)
);

NAND2xp5_ASAP7_75t_L g1302 ( 
.A(n_1132),
.B(n_1138),
.Y(n_1302)
);

INVx2_ASAP7_75t_L g1303 ( 
.A(n_1086),
.Y(n_1303)
);

BUFx2_ASAP7_75t_L g1304 ( 
.A(n_1157),
.Y(n_1304)
);

AOI21xp5_ASAP7_75t_L g1305 ( 
.A1(n_1135),
.A2(n_1156),
.B(n_1149),
.Y(n_1305)
);

AOI22xp5_ASAP7_75t_L g1306 ( 
.A1(n_1055),
.A2(n_1138),
.B1(n_1132),
.B2(n_1152),
.Y(n_1306)
);

OAI21xp5_ASAP7_75t_L g1307 ( 
.A1(n_1152),
.A2(n_1158),
.B(n_1153),
.Y(n_1307)
);

OAI221xp5_ASAP7_75t_L g1308 ( 
.A1(n_1152),
.A2(n_737),
.B1(n_684),
.B2(n_1158),
.C(n_1153),
.Y(n_1308)
);

CKINVDCx6p67_ASAP7_75t_R g1309 ( 
.A(n_1053),
.Y(n_1309)
);

NOR2xp33_ASAP7_75t_L g1310 ( 
.A(n_1132),
.B(n_1138),
.Y(n_1310)
);

AO31x2_ASAP7_75t_L g1311 ( 
.A1(n_1133),
.A2(n_839),
.A3(n_863),
.B(n_1120),
.Y(n_1311)
);

INVx2_ASAP7_75t_L g1312 ( 
.A(n_1086),
.Y(n_1312)
);

INVx2_ASAP7_75t_L g1313 ( 
.A(n_1086),
.Y(n_1313)
);

NOR2xp33_ASAP7_75t_L g1314 ( 
.A(n_1132),
.B(n_1138),
.Y(n_1314)
);

NAND2xp5_ASAP7_75t_L g1315 ( 
.A(n_1132),
.B(n_1138),
.Y(n_1315)
);

INVx1_ASAP7_75t_L g1316 ( 
.A(n_1032),
.Y(n_1316)
);

OAI222xp33_ASAP7_75t_L g1317 ( 
.A1(n_1059),
.A2(n_392),
.B1(n_1124),
.B2(n_1055),
.C1(n_508),
.C2(n_489),
.Y(n_1317)
);

OAI21xp5_ASAP7_75t_SL g1318 ( 
.A1(n_1055),
.A2(n_1059),
.B(n_684),
.Y(n_1318)
);

BUFx2_ASAP7_75t_L g1319 ( 
.A(n_1157),
.Y(n_1319)
);

INVx2_ASAP7_75t_SL g1320 ( 
.A(n_1157),
.Y(n_1320)
);

AO22x2_ASAP7_75t_L g1321 ( 
.A1(n_1055),
.A2(n_1049),
.B1(n_1124),
.B2(n_1068),
.Y(n_1321)
);

INVx1_ASAP7_75t_SL g1322 ( 
.A(n_1020),
.Y(n_1322)
);

INVx2_ASAP7_75t_L g1323 ( 
.A(n_1086),
.Y(n_1323)
);

NAND3xp33_ASAP7_75t_L g1324 ( 
.A(n_1152),
.B(n_1158),
.C(n_1153),
.Y(n_1324)
);

O2A1O1Ixp33_ASAP7_75t_SL g1325 ( 
.A1(n_1152),
.A2(n_1153),
.B(n_1158),
.C(n_1148),
.Y(n_1325)
);

AOI21xp5_ASAP7_75t_L g1326 ( 
.A1(n_1135),
.A2(n_1156),
.B(n_1149),
.Y(n_1326)
);

BUFx2_ASAP7_75t_L g1327 ( 
.A(n_1157),
.Y(n_1327)
);

OAI22xp5_ASAP7_75t_SL g1328 ( 
.A1(n_1262),
.A2(n_1306),
.B1(n_1314),
.B2(n_1310),
.Y(n_1328)
);

OAI21xp5_ASAP7_75t_SL g1329 ( 
.A1(n_1306),
.A2(n_1173),
.B(n_1318),
.Y(n_1329)
);

CKINVDCx11_ASAP7_75t_R g1330 ( 
.A(n_1205),
.Y(n_1330)
);

AOI22xp33_ASAP7_75t_L g1331 ( 
.A1(n_1253),
.A2(n_1259),
.B1(n_1207),
.B2(n_1200),
.Y(n_1331)
);

CKINVDCx5p33_ASAP7_75t_R g1332 ( 
.A(n_1177),
.Y(n_1332)
);

OAI22xp33_ASAP7_75t_L g1333 ( 
.A1(n_1207),
.A2(n_1255),
.B1(n_1318),
.B2(n_1274),
.Y(n_1333)
);

BUFx12f_ASAP7_75t_L g1334 ( 
.A(n_1268),
.Y(n_1334)
);

INVx6_ASAP7_75t_L g1335 ( 
.A(n_1215),
.Y(n_1335)
);

AOI22xp33_ASAP7_75t_L g1336 ( 
.A1(n_1321),
.A2(n_1265),
.B1(n_1290),
.B2(n_1204),
.Y(n_1336)
);

AOI22xp33_ASAP7_75t_SL g1337 ( 
.A1(n_1255),
.A2(n_1321),
.B1(n_1317),
.B2(n_1324),
.Y(n_1337)
);

AOI22xp5_ASAP7_75t_L g1338 ( 
.A1(n_1214),
.A2(n_1229),
.B1(n_1299),
.B2(n_1175),
.Y(n_1338)
);

AOI22xp33_ASAP7_75t_L g1339 ( 
.A1(n_1324),
.A2(n_1252),
.B1(n_1307),
.B2(n_1279),
.Y(n_1339)
);

INVx1_ASAP7_75t_L g1340 ( 
.A(n_1201),
.Y(n_1340)
);

AOI22xp33_ASAP7_75t_L g1341 ( 
.A1(n_1252),
.A2(n_1279),
.B1(n_1288),
.B2(n_1307),
.Y(n_1341)
);

OAI21xp5_ASAP7_75t_SL g1342 ( 
.A1(n_1288),
.A2(n_1254),
.B(n_1251),
.Y(n_1342)
);

OAI22xp5_ASAP7_75t_L g1343 ( 
.A1(n_1308),
.A2(n_1223),
.B1(n_1196),
.B2(n_1302),
.Y(n_1343)
);

BUFx2_ASAP7_75t_L g1344 ( 
.A(n_1206),
.Y(n_1344)
);

BUFx10_ASAP7_75t_L g1345 ( 
.A(n_1289),
.Y(n_1345)
);

INVx1_ASAP7_75t_L g1346 ( 
.A(n_1260),
.Y(n_1346)
);

INVx1_ASAP7_75t_L g1347 ( 
.A(n_1264),
.Y(n_1347)
);

INVx3_ASAP7_75t_L g1348 ( 
.A(n_1226),
.Y(n_1348)
);

AOI22xp33_ASAP7_75t_L g1349 ( 
.A1(n_1190),
.A2(n_1285),
.B1(n_1270),
.B2(n_1313),
.Y(n_1349)
);

AOI22xp33_ASAP7_75t_L g1350 ( 
.A1(n_1190),
.A2(n_1296),
.B1(n_1312),
.B2(n_1323),
.Y(n_1350)
);

OAI22xp5_ASAP7_75t_L g1351 ( 
.A1(n_1181),
.A2(n_1261),
.B1(n_1315),
.B2(n_1297),
.Y(n_1351)
);

AOI22xp5_ASAP7_75t_L g1352 ( 
.A1(n_1214),
.A2(n_1197),
.B1(n_1272),
.B2(n_1263),
.Y(n_1352)
);

INVx6_ASAP7_75t_L g1353 ( 
.A(n_1281),
.Y(n_1353)
);

BUFx2_ASAP7_75t_R g1354 ( 
.A(n_1275),
.Y(n_1354)
);

AOI22xp33_ASAP7_75t_L g1355 ( 
.A1(n_1182),
.A2(n_1203),
.B1(n_1278),
.B2(n_1236),
.Y(n_1355)
);

AOI22xp33_ASAP7_75t_L g1356 ( 
.A1(n_1287),
.A2(n_1185),
.B1(n_1179),
.B2(n_1193),
.Y(n_1356)
);

BUFx3_ASAP7_75t_L g1357 ( 
.A(n_1289),
.Y(n_1357)
);

AOI22xp33_ASAP7_75t_SL g1358 ( 
.A1(n_1179),
.A2(n_1185),
.B1(n_1195),
.B2(n_1211),
.Y(n_1358)
);

OAI21xp5_ASAP7_75t_SL g1359 ( 
.A1(n_1258),
.A2(n_1293),
.B(n_1277),
.Y(n_1359)
);

AOI22xp33_ASAP7_75t_L g1360 ( 
.A1(n_1183),
.A2(n_1234),
.B1(n_1235),
.B2(n_1276),
.Y(n_1360)
);

AOI22xp33_ASAP7_75t_L g1361 ( 
.A1(n_1257),
.A2(n_1269),
.B1(n_1303),
.B2(n_1282),
.Y(n_1361)
);

AOI22xp33_ASAP7_75t_SL g1362 ( 
.A1(n_1211),
.A2(n_1194),
.B1(n_1221),
.B2(n_1189),
.Y(n_1362)
);

INVx4_ASAP7_75t_L g1363 ( 
.A(n_1216),
.Y(n_1363)
);

CKINVDCx11_ASAP7_75t_R g1364 ( 
.A(n_1309),
.Y(n_1364)
);

OAI22xp5_ASAP7_75t_L g1365 ( 
.A1(n_1240),
.A2(n_1172),
.B1(n_1280),
.B2(n_1212),
.Y(n_1365)
);

CKINVDCx5p33_ASAP7_75t_R g1366 ( 
.A(n_1304),
.Y(n_1366)
);

AOI22xp33_ASAP7_75t_SL g1367 ( 
.A1(n_1194),
.A2(n_1221),
.B1(n_1189),
.B2(n_1176),
.Y(n_1367)
);

BUFx2_ASAP7_75t_L g1368 ( 
.A(n_1227),
.Y(n_1368)
);

INVx1_ASAP7_75t_SL g1369 ( 
.A(n_1319),
.Y(n_1369)
);

BUFx3_ASAP7_75t_L g1370 ( 
.A(n_1327),
.Y(n_1370)
);

AOI22xp33_ASAP7_75t_L g1371 ( 
.A1(n_1283),
.A2(n_1294),
.B1(n_1316),
.B2(n_1322),
.Y(n_1371)
);

AND2x2_ASAP7_75t_L g1372 ( 
.A(n_1213),
.B(n_1322),
.Y(n_1372)
);

NAND2xp5_ASAP7_75t_L g1373 ( 
.A(n_1176),
.B(n_1242),
.Y(n_1373)
);

INVx4_ASAP7_75t_L g1374 ( 
.A(n_1238),
.Y(n_1374)
);

AOI22xp33_ASAP7_75t_SL g1375 ( 
.A1(n_1194),
.A2(n_1221),
.B1(n_1220),
.B2(n_1198),
.Y(n_1375)
);

CKINVDCx6p67_ASAP7_75t_R g1376 ( 
.A(n_1271),
.Y(n_1376)
);

BUFx8_ASAP7_75t_L g1377 ( 
.A(n_1178),
.Y(n_1377)
);

OAI22xp33_ASAP7_75t_SL g1378 ( 
.A1(n_1240),
.A2(n_1271),
.B1(n_1218),
.B2(n_1225),
.Y(n_1378)
);

BUFx3_ASAP7_75t_L g1379 ( 
.A(n_1320),
.Y(n_1379)
);

NAND2xp5_ASAP7_75t_L g1380 ( 
.A(n_1239),
.B(n_1241),
.Y(n_1380)
);

AOI22xp33_ASAP7_75t_SL g1381 ( 
.A1(n_1198),
.A2(n_1244),
.B1(n_1228),
.B2(n_1231),
.Y(n_1381)
);

BUFx2_ASAP7_75t_L g1382 ( 
.A(n_1228),
.Y(n_1382)
);

AOI21xp5_ASAP7_75t_SL g1383 ( 
.A1(n_1232),
.A2(n_1245),
.B(n_1247),
.Y(n_1383)
);

BUFx12f_ASAP7_75t_L g1384 ( 
.A(n_1180),
.Y(n_1384)
);

AOI22xp33_ASAP7_75t_L g1385 ( 
.A1(n_1233),
.A2(n_1174),
.B1(n_1305),
.B2(n_1256),
.Y(n_1385)
);

AOI22xp33_ASAP7_75t_SL g1386 ( 
.A1(n_1284),
.A2(n_1292),
.B1(n_1325),
.B2(n_1301),
.Y(n_1386)
);

AOI22xp33_ASAP7_75t_L g1387 ( 
.A1(n_1250),
.A2(n_1326),
.B1(n_1208),
.B2(n_1217),
.Y(n_1387)
);

AOI22xp33_ASAP7_75t_L g1388 ( 
.A1(n_1230),
.A2(n_1222),
.B1(n_1249),
.B2(n_1243),
.Y(n_1388)
);

NAND2xp5_ASAP7_75t_L g1389 ( 
.A(n_1210),
.B(n_1237),
.Y(n_1389)
);

AOI22xp33_ASAP7_75t_L g1390 ( 
.A1(n_1248),
.A2(n_1209),
.B1(n_1199),
.B2(n_1266),
.Y(n_1390)
);

BUFx2_ASAP7_75t_L g1391 ( 
.A(n_1180),
.Y(n_1391)
);

CKINVDCx20_ASAP7_75t_R g1392 ( 
.A(n_1266),
.Y(n_1392)
);

OAI22xp5_ASAP7_75t_L g1393 ( 
.A1(n_1202),
.A2(n_1192),
.B1(n_1246),
.B2(n_1219),
.Y(n_1393)
);

OAI22xp33_ASAP7_75t_L g1394 ( 
.A1(n_1286),
.A2(n_1311),
.B1(n_1295),
.B2(n_1224),
.Y(n_1394)
);

INVxp67_ASAP7_75t_L g1395 ( 
.A(n_1186),
.Y(n_1395)
);

AOI21xp5_ASAP7_75t_L g1396 ( 
.A1(n_1187),
.A2(n_1267),
.B(n_1273),
.Y(n_1396)
);

INVx3_ASAP7_75t_L g1397 ( 
.A(n_1295),
.Y(n_1397)
);

AOI22xp33_ASAP7_75t_L g1398 ( 
.A1(n_1291),
.A2(n_1298),
.B1(n_1300),
.B2(n_1311),
.Y(n_1398)
);

AOI22xp33_ASAP7_75t_SL g1399 ( 
.A1(n_1255),
.A2(n_1055),
.B1(n_1321),
.B2(n_1124),
.Y(n_1399)
);

NAND2xp5_ASAP7_75t_L g1400 ( 
.A(n_1310),
.B(n_1314),
.Y(n_1400)
);

BUFx10_ASAP7_75t_L g1401 ( 
.A(n_1177),
.Y(n_1401)
);

INVx1_ASAP7_75t_SL g1402 ( 
.A(n_1304),
.Y(n_1402)
);

INVx8_ASAP7_75t_L g1403 ( 
.A(n_1221),
.Y(n_1403)
);

BUFx4f_ASAP7_75t_L g1404 ( 
.A(n_1191),
.Y(n_1404)
);

BUFx2_ASAP7_75t_L g1405 ( 
.A(n_1206),
.Y(n_1405)
);

CKINVDCx8_ASAP7_75t_R g1406 ( 
.A(n_1177),
.Y(n_1406)
);

AND2x2_ASAP7_75t_L g1407 ( 
.A(n_1175),
.B(n_1310),
.Y(n_1407)
);

INVx4_ASAP7_75t_L g1408 ( 
.A(n_1188),
.Y(n_1408)
);

OAI22xp33_ASAP7_75t_L g1409 ( 
.A1(n_1306),
.A2(n_1207),
.B1(n_1059),
.B2(n_1255),
.Y(n_1409)
);

AOI22xp33_ASAP7_75t_L g1410 ( 
.A1(n_1262),
.A2(n_1055),
.B1(n_1200),
.B2(n_649),
.Y(n_1410)
);

BUFx6f_ASAP7_75t_SL g1411 ( 
.A(n_1191),
.Y(n_1411)
);

CKINVDCx20_ASAP7_75t_R g1412 ( 
.A(n_1177),
.Y(n_1412)
);

AOI22xp5_ASAP7_75t_L g1413 ( 
.A1(n_1262),
.A2(n_1055),
.B1(n_539),
.B2(n_1059),
.Y(n_1413)
);

INVx5_ASAP7_75t_L g1414 ( 
.A(n_1271),
.Y(n_1414)
);

OAI22xp5_ASAP7_75t_L g1415 ( 
.A1(n_1262),
.A2(n_1306),
.B1(n_1152),
.B2(n_1158),
.Y(n_1415)
);

NAND2xp5_ASAP7_75t_L g1416 ( 
.A(n_1310),
.B(n_1314),
.Y(n_1416)
);

BUFx4f_ASAP7_75t_L g1417 ( 
.A(n_1191),
.Y(n_1417)
);

INVx1_ASAP7_75t_L g1418 ( 
.A(n_1184),
.Y(n_1418)
);

AOI22xp5_ASAP7_75t_L g1419 ( 
.A1(n_1262),
.A2(n_1055),
.B1(n_539),
.B2(n_1059),
.Y(n_1419)
);

AOI22xp33_ASAP7_75t_L g1420 ( 
.A1(n_1262),
.A2(n_1055),
.B1(n_1200),
.B2(n_649),
.Y(n_1420)
);

AND2x2_ASAP7_75t_L g1421 ( 
.A(n_1175),
.B(n_1310),
.Y(n_1421)
);

BUFx3_ASAP7_75t_L g1422 ( 
.A(n_1191),
.Y(n_1422)
);

OAI22xp33_ASAP7_75t_L g1423 ( 
.A1(n_1306),
.A2(n_1207),
.B1(n_1059),
.B2(n_1255),
.Y(n_1423)
);

INVx1_ASAP7_75t_L g1424 ( 
.A(n_1184),
.Y(n_1424)
);

AOI22xp5_ASAP7_75t_L g1425 ( 
.A1(n_1262),
.A2(n_1055),
.B1(n_539),
.B2(n_1059),
.Y(n_1425)
);

AOI22xp33_ASAP7_75t_SL g1426 ( 
.A1(n_1255),
.A2(n_1055),
.B1(n_1321),
.B2(n_1124),
.Y(n_1426)
);

AOI22xp33_ASAP7_75t_SL g1427 ( 
.A1(n_1255),
.A2(n_1055),
.B1(n_1321),
.B2(n_1124),
.Y(n_1427)
);

BUFx3_ASAP7_75t_L g1428 ( 
.A(n_1191),
.Y(n_1428)
);

AOI22xp33_ASAP7_75t_L g1429 ( 
.A1(n_1262),
.A2(n_1055),
.B1(n_1259),
.B2(n_1253),
.Y(n_1429)
);

BUFx10_ASAP7_75t_L g1430 ( 
.A(n_1177),
.Y(n_1430)
);

NAND2xp5_ASAP7_75t_L g1431 ( 
.A(n_1310),
.B(n_1314),
.Y(n_1431)
);

INVx4_ASAP7_75t_L g1432 ( 
.A(n_1188),
.Y(n_1432)
);

CKINVDCx11_ASAP7_75t_R g1433 ( 
.A(n_1205),
.Y(n_1433)
);

CKINVDCx20_ASAP7_75t_R g1434 ( 
.A(n_1177),
.Y(n_1434)
);

AOI22xp33_ASAP7_75t_SL g1435 ( 
.A1(n_1255),
.A2(n_1055),
.B1(n_1321),
.B2(n_1124),
.Y(n_1435)
);

OAI22xp33_ASAP7_75t_L g1436 ( 
.A1(n_1306),
.A2(n_1207),
.B1(n_1059),
.B2(n_1255),
.Y(n_1436)
);

INVx1_ASAP7_75t_L g1437 ( 
.A(n_1184),
.Y(n_1437)
);

INVx1_ASAP7_75t_L g1438 ( 
.A(n_1184),
.Y(n_1438)
);

OAI21xp33_ASAP7_75t_L g1439 ( 
.A1(n_1255),
.A2(n_1262),
.B(n_1055),
.Y(n_1439)
);

NOR2xp33_ASAP7_75t_SL g1440 ( 
.A(n_1439),
.B(n_1409),
.Y(n_1440)
);

OAI21xp5_ASAP7_75t_L g1441 ( 
.A1(n_1331),
.A2(n_1342),
.B(n_1341),
.Y(n_1441)
);

AND2x2_ASAP7_75t_L g1442 ( 
.A(n_1341),
.B(n_1339),
.Y(n_1442)
);

AND2x2_ASAP7_75t_L g1443 ( 
.A(n_1358),
.B(n_1339),
.Y(n_1443)
);

BUFx2_ASAP7_75t_L g1444 ( 
.A(n_1395),
.Y(n_1444)
);

INVx3_ASAP7_75t_L g1445 ( 
.A(n_1397),
.Y(n_1445)
);

INVx1_ASAP7_75t_L g1446 ( 
.A(n_1389),
.Y(n_1446)
);

HB1xp67_ASAP7_75t_L g1447 ( 
.A(n_1395),
.Y(n_1447)
);

NAND2xp5_ASAP7_75t_L g1448 ( 
.A(n_1358),
.B(n_1351),
.Y(n_1448)
);

OAI21x1_ASAP7_75t_L g1449 ( 
.A1(n_1396),
.A2(n_1387),
.B(n_1385),
.Y(n_1449)
);

INVx1_ASAP7_75t_L g1450 ( 
.A(n_1340),
.Y(n_1450)
);

NAND2xp5_ASAP7_75t_L g1451 ( 
.A(n_1356),
.B(n_1333),
.Y(n_1451)
);

BUFx8_ASAP7_75t_L g1452 ( 
.A(n_1411),
.Y(n_1452)
);

HB1xp67_ASAP7_75t_L g1453 ( 
.A(n_1393),
.Y(n_1453)
);

OAI21x1_ASAP7_75t_L g1454 ( 
.A1(n_1396),
.A2(n_1387),
.B(n_1385),
.Y(n_1454)
);

AND2x4_ASAP7_75t_L g1455 ( 
.A(n_1348),
.B(n_1414),
.Y(n_1455)
);

INVx1_ASAP7_75t_L g1456 ( 
.A(n_1346),
.Y(n_1456)
);

INVx1_ASAP7_75t_L g1457 ( 
.A(n_1347),
.Y(n_1457)
);

AND2x2_ASAP7_75t_L g1458 ( 
.A(n_1407),
.B(n_1421),
.Y(n_1458)
);

INVx4_ASAP7_75t_L g1459 ( 
.A(n_1414),
.Y(n_1459)
);

AND2x2_ASAP7_75t_L g1460 ( 
.A(n_1355),
.B(n_1399),
.Y(n_1460)
);

OA21x2_ASAP7_75t_L g1461 ( 
.A1(n_1398),
.A2(n_1329),
.B(n_1388),
.Y(n_1461)
);

INVx1_ASAP7_75t_L g1462 ( 
.A(n_1418),
.Y(n_1462)
);

CKINVDCx5p33_ASAP7_75t_R g1463 ( 
.A(n_1330),
.Y(n_1463)
);

INVxp67_ASAP7_75t_L g1464 ( 
.A(n_1380),
.Y(n_1464)
);

INVx1_ASAP7_75t_L g1465 ( 
.A(n_1424),
.Y(n_1465)
);

CKINVDCx11_ASAP7_75t_R g1466 ( 
.A(n_1406),
.Y(n_1466)
);

OAI21x1_ASAP7_75t_L g1467 ( 
.A1(n_1390),
.A2(n_1415),
.B(n_1383),
.Y(n_1467)
);

BUFx2_ASAP7_75t_L g1468 ( 
.A(n_1348),
.Y(n_1468)
);

INVx2_ASAP7_75t_L g1469 ( 
.A(n_1437),
.Y(n_1469)
);

BUFx12f_ASAP7_75t_SL g1470 ( 
.A(n_1374),
.Y(n_1470)
);

OAI21x1_ASAP7_75t_L g1471 ( 
.A1(n_1349),
.A2(n_1336),
.B(n_1365),
.Y(n_1471)
);

INVx1_ASAP7_75t_L g1472 ( 
.A(n_1438),
.Y(n_1472)
);

AOI21xp5_ASAP7_75t_L g1473 ( 
.A1(n_1409),
.A2(n_1436),
.B(n_1423),
.Y(n_1473)
);

BUFx2_ASAP7_75t_L g1474 ( 
.A(n_1392),
.Y(n_1474)
);

INVx1_ASAP7_75t_L g1475 ( 
.A(n_1394),
.Y(n_1475)
);

INVx1_ASAP7_75t_L g1476 ( 
.A(n_1394),
.Y(n_1476)
);

BUFx4f_ASAP7_75t_SL g1477 ( 
.A(n_1412),
.Y(n_1477)
);

AND4x1_ASAP7_75t_SL g1478 ( 
.A(n_1400),
.B(n_1416),
.C(n_1431),
.D(n_1425),
.Y(n_1478)
);

HB1xp67_ASAP7_75t_L g1479 ( 
.A(n_1352),
.Y(n_1479)
);

AND2x2_ASAP7_75t_L g1480 ( 
.A(n_1355),
.B(n_1399),
.Y(n_1480)
);

INVx1_ASAP7_75t_L g1481 ( 
.A(n_1381),
.Y(n_1481)
);

INVx1_ASAP7_75t_L g1482 ( 
.A(n_1381),
.Y(n_1482)
);

NAND2xp5_ASAP7_75t_L g1483 ( 
.A(n_1333),
.B(n_1362),
.Y(n_1483)
);

AND2x2_ASAP7_75t_L g1484 ( 
.A(n_1426),
.B(n_1427),
.Y(n_1484)
);

INVx2_ASAP7_75t_SL g1485 ( 
.A(n_1414),
.Y(n_1485)
);

AOI22xp33_ASAP7_75t_L g1486 ( 
.A1(n_1337),
.A2(n_1426),
.B1(n_1435),
.B2(n_1427),
.Y(n_1486)
);

INVx3_ASAP7_75t_L g1487 ( 
.A(n_1384),
.Y(n_1487)
);

CKINVDCx11_ASAP7_75t_R g1488 ( 
.A(n_1433),
.Y(n_1488)
);

BUFx2_ASAP7_75t_L g1489 ( 
.A(n_1344),
.Y(n_1489)
);

AND2x2_ASAP7_75t_L g1490 ( 
.A(n_1375),
.B(n_1435),
.Y(n_1490)
);

INVx2_ASAP7_75t_SL g1491 ( 
.A(n_1335),
.Y(n_1491)
);

INVx1_ASAP7_75t_L g1492 ( 
.A(n_1375),
.Y(n_1492)
);

INVx1_ASAP7_75t_L g1493 ( 
.A(n_1423),
.Y(n_1493)
);

AND2x2_ASAP7_75t_L g1494 ( 
.A(n_1362),
.B(n_1367),
.Y(n_1494)
);

OAI21x1_ASAP7_75t_L g1495 ( 
.A1(n_1359),
.A2(n_1343),
.B(n_1331),
.Y(n_1495)
);

OAI21x1_ASAP7_75t_L g1496 ( 
.A1(n_1360),
.A2(n_1338),
.B(n_1350),
.Y(n_1496)
);

INVx1_ASAP7_75t_L g1497 ( 
.A(n_1436),
.Y(n_1497)
);

AND2x2_ASAP7_75t_L g1498 ( 
.A(n_1367),
.B(n_1360),
.Y(n_1498)
);

INVx1_ASAP7_75t_L g1499 ( 
.A(n_1378),
.Y(n_1499)
);

INVx2_ASAP7_75t_L g1500 ( 
.A(n_1382),
.Y(n_1500)
);

INVx1_ASAP7_75t_L g1501 ( 
.A(n_1371),
.Y(n_1501)
);

AND2x2_ASAP7_75t_L g1502 ( 
.A(n_1372),
.B(n_1337),
.Y(n_1502)
);

A2O1A1Ixp33_ASAP7_75t_L g1503 ( 
.A1(n_1413),
.A2(n_1419),
.B(n_1410),
.C(n_1420),
.Y(n_1503)
);

BUFx2_ASAP7_75t_L g1504 ( 
.A(n_1405),
.Y(n_1504)
);

INVx1_ASAP7_75t_L g1505 ( 
.A(n_1386),
.Y(n_1505)
);

INVx1_ASAP7_75t_L g1506 ( 
.A(n_1386),
.Y(n_1506)
);

OR2x2_ASAP7_75t_L g1507 ( 
.A(n_1373),
.B(n_1328),
.Y(n_1507)
);

OAI211xp5_ASAP7_75t_L g1508 ( 
.A1(n_1429),
.A2(n_1432),
.B(n_1408),
.C(n_1369),
.Y(n_1508)
);

BUFx3_ASAP7_75t_L g1509 ( 
.A(n_1376),
.Y(n_1509)
);

NAND3xp33_ASAP7_75t_L g1510 ( 
.A(n_1429),
.B(n_1377),
.C(n_1366),
.Y(n_1510)
);

INVx1_ASAP7_75t_L g1511 ( 
.A(n_1361),
.Y(n_1511)
);

AND2x2_ASAP7_75t_L g1512 ( 
.A(n_1368),
.B(n_1370),
.Y(n_1512)
);

BUFx2_ASAP7_75t_L g1513 ( 
.A(n_1391),
.Y(n_1513)
);

NAND2xp5_ASAP7_75t_L g1514 ( 
.A(n_1374),
.B(n_1363),
.Y(n_1514)
);

BUFx3_ASAP7_75t_L g1515 ( 
.A(n_1335),
.Y(n_1515)
);

HB1xp67_ASAP7_75t_L g1516 ( 
.A(n_1402),
.Y(n_1516)
);

NOR2xp33_ASAP7_75t_L g1517 ( 
.A(n_1354),
.B(n_1379),
.Y(n_1517)
);

INVx3_ASAP7_75t_L g1518 ( 
.A(n_1403),
.Y(n_1518)
);

AOI221xp5_ASAP7_75t_L g1519 ( 
.A1(n_1448),
.A2(n_1357),
.B1(n_1428),
.B2(n_1422),
.C(n_1411),
.Y(n_1519)
);

NOR2xp33_ASAP7_75t_SL g1520 ( 
.A(n_1463),
.B(n_1417),
.Y(n_1520)
);

AO32x1_ASAP7_75t_L g1521 ( 
.A1(n_1443),
.A2(n_1377),
.A3(n_1345),
.B1(n_1403),
.B2(n_1353),
.Y(n_1521)
);

AO21x2_ASAP7_75t_L g1522 ( 
.A1(n_1451),
.A2(n_1404),
.B(n_1364),
.Y(n_1522)
);

NAND4xp25_ASAP7_75t_L g1523 ( 
.A(n_1443),
.B(n_1401),
.C(n_1430),
.D(n_1334),
.Y(n_1523)
);

OA21x2_ASAP7_75t_L g1524 ( 
.A1(n_1449),
.A2(n_1332),
.B(n_1401),
.Y(n_1524)
);

AND2x2_ASAP7_75t_L g1525 ( 
.A(n_1512),
.B(n_1430),
.Y(n_1525)
);

AO32x2_ASAP7_75t_L g1526 ( 
.A1(n_1485),
.A2(n_1434),
.A3(n_1491),
.B1(n_1464),
.B2(n_1459),
.Y(n_1526)
);

AOI221xp5_ASAP7_75t_L g1527 ( 
.A1(n_1441),
.A2(n_1451),
.B1(n_1503),
.B2(n_1483),
.C(n_1492),
.Y(n_1527)
);

AOI22xp33_ASAP7_75t_L g1528 ( 
.A1(n_1440),
.A2(n_1473),
.B1(n_1441),
.B2(n_1483),
.Y(n_1528)
);

AOI22xp5_ASAP7_75t_L g1529 ( 
.A1(n_1490),
.A2(n_1473),
.B1(n_1442),
.B2(n_1484),
.Y(n_1529)
);

AND2x4_ASAP7_75t_L g1530 ( 
.A(n_1500),
.B(n_1468),
.Y(n_1530)
);

AND2x2_ASAP7_75t_L g1531 ( 
.A(n_1458),
.B(n_1489),
.Y(n_1531)
);

NOR2x1p5_ASAP7_75t_L g1532 ( 
.A(n_1510),
.B(n_1509),
.Y(n_1532)
);

AND2x2_ASAP7_75t_L g1533 ( 
.A(n_1458),
.B(n_1489),
.Y(n_1533)
);

CKINVDCx5p33_ASAP7_75t_R g1534 ( 
.A(n_1466),
.Y(n_1534)
);

NOR2xp33_ASAP7_75t_L g1535 ( 
.A(n_1495),
.B(n_1507),
.Y(n_1535)
);

AND2x2_ASAP7_75t_L g1536 ( 
.A(n_1504),
.B(n_1513),
.Y(n_1536)
);

HB1xp67_ASAP7_75t_L g1537 ( 
.A(n_1447),
.Y(n_1537)
);

AND2x2_ASAP7_75t_L g1538 ( 
.A(n_1516),
.B(n_1474),
.Y(n_1538)
);

NOR2x1_ASAP7_75t_SL g1539 ( 
.A(n_1508),
.B(n_1507),
.Y(n_1539)
);

A2O1A1Ixp33_ASAP7_75t_L g1540 ( 
.A1(n_1495),
.A2(n_1490),
.B(n_1471),
.C(n_1494),
.Y(n_1540)
);

OAI21x1_ASAP7_75t_L g1541 ( 
.A1(n_1449),
.A2(n_1454),
.B(n_1467),
.Y(n_1541)
);

NOR2xp33_ASAP7_75t_L g1542 ( 
.A(n_1495),
.B(n_1479),
.Y(n_1542)
);

AOI221xp5_ASAP7_75t_L g1543 ( 
.A1(n_1490),
.A2(n_1460),
.B1(n_1480),
.B2(n_1481),
.C(n_1482),
.Y(n_1543)
);

NAND4xp25_ASAP7_75t_L g1544 ( 
.A(n_1510),
.B(n_1442),
.C(n_1506),
.D(n_1505),
.Y(n_1544)
);

OA21x2_ASAP7_75t_L g1545 ( 
.A1(n_1449),
.A2(n_1454),
.B(n_1467),
.Y(n_1545)
);

OAI21xp5_ASAP7_75t_L g1546 ( 
.A1(n_1467),
.A2(n_1479),
.B(n_1506),
.Y(n_1546)
);

OAI21xp5_ASAP7_75t_L g1547 ( 
.A1(n_1505),
.A2(n_1471),
.B(n_1453),
.Y(n_1547)
);

OAI21xp5_ASAP7_75t_L g1548 ( 
.A1(n_1471),
.A2(n_1453),
.B(n_1494),
.Y(n_1548)
);

OAI22xp5_ASAP7_75t_L g1549 ( 
.A1(n_1486),
.A2(n_1493),
.B1(n_1497),
.B2(n_1484),
.Y(n_1549)
);

HB1xp67_ASAP7_75t_L g1550 ( 
.A(n_1447),
.Y(n_1550)
);

AND2x6_ASAP7_75t_L g1551 ( 
.A(n_1455),
.B(n_1518),
.Y(n_1551)
);

NAND2xp5_ASAP7_75t_L g1552 ( 
.A(n_1469),
.B(n_1450),
.Y(n_1552)
);

AND2x2_ASAP7_75t_L g1553 ( 
.A(n_1456),
.B(n_1457),
.Y(n_1553)
);

AND2x2_ASAP7_75t_L g1554 ( 
.A(n_1456),
.B(n_1457),
.Y(n_1554)
);

AND2x2_ASAP7_75t_L g1555 ( 
.A(n_1462),
.B(n_1465),
.Y(n_1555)
);

O2A1O1Ixp33_ASAP7_75t_SL g1556 ( 
.A1(n_1514),
.A2(n_1491),
.B(n_1493),
.C(n_1497),
.Y(n_1556)
);

AO32x2_ASAP7_75t_L g1557 ( 
.A1(n_1491),
.A2(n_1459),
.A3(n_1478),
.B1(n_1476),
.B2(n_1475),
.Y(n_1557)
);

OAI22xp5_ASAP7_75t_L g1558 ( 
.A1(n_1494),
.A2(n_1461),
.B1(n_1480),
.B2(n_1460),
.Y(n_1558)
);

AND2x2_ASAP7_75t_L g1559 ( 
.A(n_1545),
.B(n_1481),
.Y(n_1559)
);

AND2x2_ASAP7_75t_L g1560 ( 
.A(n_1545),
.B(n_1482),
.Y(n_1560)
);

BUFx3_ASAP7_75t_L g1561 ( 
.A(n_1551),
.Y(n_1561)
);

HB1xp67_ASAP7_75t_L g1562 ( 
.A(n_1537),
.Y(n_1562)
);

INVx1_ASAP7_75t_SL g1563 ( 
.A(n_1537),
.Y(n_1563)
);

NAND2xp5_ASAP7_75t_L g1564 ( 
.A(n_1535),
.B(n_1446),
.Y(n_1564)
);

AND2x2_ASAP7_75t_L g1565 ( 
.A(n_1541),
.B(n_1444),
.Y(n_1565)
);

AND2x2_ASAP7_75t_L g1566 ( 
.A(n_1541),
.B(n_1461),
.Y(n_1566)
);

AOI22xp33_ASAP7_75t_L g1567 ( 
.A1(n_1527),
.A2(n_1498),
.B1(n_1502),
.B2(n_1501),
.Y(n_1567)
);

AND2x2_ASAP7_75t_L g1568 ( 
.A(n_1531),
.B(n_1461),
.Y(n_1568)
);

HB1xp67_ASAP7_75t_L g1569 ( 
.A(n_1550),
.Y(n_1569)
);

NAND2xp5_ASAP7_75t_L g1570 ( 
.A(n_1535),
.B(n_1446),
.Y(n_1570)
);

AND2x2_ASAP7_75t_L g1571 ( 
.A(n_1533),
.B(n_1461),
.Y(n_1571)
);

AND2x2_ASAP7_75t_L g1572 ( 
.A(n_1524),
.B(n_1461),
.Y(n_1572)
);

AOI22xp33_ASAP7_75t_L g1573 ( 
.A1(n_1528),
.A2(n_1498),
.B1(n_1502),
.B2(n_1501),
.Y(n_1573)
);

AND2x2_ASAP7_75t_L g1574 ( 
.A(n_1524),
.B(n_1465),
.Y(n_1574)
);

AOI22xp33_ASAP7_75t_L g1575 ( 
.A1(n_1528),
.A2(n_1496),
.B1(n_1476),
.B2(n_1475),
.Y(n_1575)
);

INVx5_ASAP7_75t_L g1576 ( 
.A(n_1551),
.Y(n_1576)
);

OR2x2_ASAP7_75t_L g1577 ( 
.A(n_1542),
.B(n_1472),
.Y(n_1577)
);

BUFx2_ASAP7_75t_L g1578 ( 
.A(n_1526),
.Y(n_1578)
);

BUFx12f_ASAP7_75t_L g1579 ( 
.A(n_1534),
.Y(n_1579)
);

AOI22xp33_ASAP7_75t_L g1580 ( 
.A1(n_1558),
.A2(n_1496),
.B1(n_1499),
.B2(n_1511),
.Y(n_1580)
);

AND2x2_ASAP7_75t_L g1581 ( 
.A(n_1524),
.B(n_1472),
.Y(n_1581)
);

INVxp67_ASAP7_75t_SL g1582 ( 
.A(n_1552),
.Y(n_1582)
);

AOI211xp5_ASAP7_75t_L g1583 ( 
.A1(n_1544),
.A2(n_1517),
.B(n_1478),
.C(n_1499),
.Y(n_1583)
);

AND2x4_ASAP7_75t_L g1584 ( 
.A(n_1551),
.B(n_1445),
.Y(n_1584)
);

INVxp67_ASAP7_75t_L g1585 ( 
.A(n_1536),
.Y(n_1585)
);

HB1xp67_ASAP7_75t_L g1586 ( 
.A(n_1530),
.Y(n_1586)
);

NAND2xp5_ASAP7_75t_L g1587 ( 
.A(n_1582),
.B(n_1553),
.Y(n_1587)
);

AOI22xp33_ASAP7_75t_SL g1588 ( 
.A1(n_1578),
.A2(n_1539),
.B1(n_1548),
.B2(n_1549),
.Y(n_1588)
);

AND2x2_ASAP7_75t_L g1589 ( 
.A(n_1568),
.B(n_1557),
.Y(n_1589)
);

AND2x4_ASAP7_75t_L g1590 ( 
.A(n_1576),
.B(n_1551),
.Y(n_1590)
);

INVx5_ASAP7_75t_SL g1591 ( 
.A(n_1584),
.Y(n_1591)
);

NAND2xp5_ASAP7_75t_L g1592 ( 
.A(n_1582),
.B(n_1554),
.Y(n_1592)
);

HB1xp67_ASAP7_75t_L g1593 ( 
.A(n_1562),
.Y(n_1593)
);

AND2x2_ASAP7_75t_L g1594 ( 
.A(n_1568),
.B(n_1557),
.Y(n_1594)
);

OAI22xp5_ASAP7_75t_L g1595 ( 
.A1(n_1583),
.A2(n_1529),
.B1(n_1540),
.B2(n_1543),
.Y(n_1595)
);

INVx2_ASAP7_75t_L g1596 ( 
.A(n_1574),
.Y(n_1596)
);

BUFx2_ASAP7_75t_L g1597 ( 
.A(n_1561),
.Y(n_1597)
);

INVx2_ASAP7_75t_L g1598 ( 
.A(n_1574),
.Y(n_1598)
);

INVx2_ASAP7_75t_L g1599 ( 
.A(n_1574),
.Y(n_1599)
);

INVx2_ASAP7_75t_L g1600 ( 
.A(n_1581),
.Y(n_1600)
);

INVx2_ASAP7_75t_L g1601 ( 
.A(n_1581),
.Y(n_1601)
);

AND2x2_ASAP7_75t_L g1602 ( 
.A(n_1568),
.B(n_1557),
.Y(n_1602)
);

NAND2xp5_ASAP7_75t_L g1603 ( 
.A(n_1582),
.B(n_1555),
.Y(n_1603)
);

HB1xp67_ASAP7_75t_L g1604 ( 
.A(n_1562),
.Y(n_1604)
);

OAI221xp5_ASAP7_75t_L g1605 ( 
.A1(n_1583),
.A2(n_1540),
.B1(n_1547),
.B2(n_1546),
.C(n_1519),
.Y(n_1605)
);

AOI21xp5_ASAP7_75t_L g1606 ( 
.A1(n_1572),
.A2(n_1556),
.B(n_1521),
.Y(n_1606)
);

AND2x2_ASAP7_75t_L g1607 ( 
.A(n_1571),
.B(n_1557),
.Y(n_1607)
);

HB1xp67_ASAP7_75t_L g1608 ( 
.A(n_1569),
.Y(n_1608)
);

INVx2_ASAP7_75t_SL g1609 ( 
.A(n_1576),
.Y(n_1609)
);

OAI211xp5_ASAP7_75t_L g1610 ( 
.A1(n_1583),
.A2(n_1523),
.B(n_1488),
.C(n_1538),
.Y(n_1610)
);

AND2x2_ASAP7_75t_L g1611 ( 
.A(n_1571),
.B(n_1526),
.Y(n_1611)
);

AND2x2_ASAP7_75t_L g1612 ( 
.A(n_1571),
.B(n_1578),
.Y(n_1612)
);

INVx2_ASAP7_75t_L g1613 ( 
.A(n_1581),
.Y(n_1613)
);

INVx1_ASAP7_75t_SL g1614 ( 
.A(n_1563),
.Y(n_1614)
);

BUFx2_ASAP7_75t_SL g1615 ( 
.A(n_1590),
.Y(n_1615)
);

AND2x2_ASAP7_75t_L g1616 ( 
.A(n_1589),
.B(n_1578),
.Y(n_1616)
);

INVx1_ASAP7_75t_L g1617 ( 
.A(n_1593),
.Y(n_1617)
);

NAND2xp5_ASAP7_75t_L g1618 ( 
.A(n_1587),
.B(n_1564),
.Y(n_1618)
);

INVx2_ASAP7_75t_L g1619 ( 
.A(n_1596),
.Y(n_1619)
);

OR2x2_ASAP7_75t_L g1620 ( 
.A(n_1589),
.B(n_1564),
.Y(n_1620)
);

NAND2xp5_ASAP7_75t_L g1621 ( 
.A(n_1587),
.B(n_1564),
.Y(n_1621)
);

INVx1_ASAP7_75t_L g1622 ( 
.A(n_1593),
.Y(n_1622)
);

INVx1_ASAP7_75t_L g1623 ( 
.A(n_1604),
.Y(n_1623)
);

INVx2_ASAP7_75t_L g1624 ( 
.A(n_1596),
.Y(n_1624)
);

AND2x2_ASAP7_75t_L g1625 ( 
.A(n_1589),
.B(n_1571),
.Y(n_1625)
);

HB1xp67_ASAP7_75t_L g1626 ( 
.A(n_1604),
.Y(n_1626)
);

AND2x4_ASAP7_75t_L g1627 ( 
.A(n_1590),
.B(n_1576),
.Y(n_1627)
);

HB1xp67_ASAP7_75t_L g1628 ( 
.A(n_1608),
.Y(n_1628)
);

INVx1_ASAP7_75t_L g1629 ( 
.A(n_1608),
.Y(n_1629)
);

CKINVDCx16_ASAP7_75t_R g1630 ( 
.A(n_1595),
.Y(n_1630)
);

BUFx2_ASAP7_75t_L g1631 ( 
.A(n_1597),
.Y(n_1631)
);

NAND2xp5_ASAP7_75t_L g1632 ( 
.A(n_1592),
.B(n_1570),
.Y(n_1632)
);

NAND2xp5_ASAP7_75t_L g1633 ( 
.A(n_1592),
.B(n_1603),
.Y(n_1633)
);

AOI22xp5_ASAP7_75t_L g1634 ( 
.A1(n_1595),
.A2(n_1567),
.B1(n_1573),
.B2(n_1575),
.Y(n_1634)
);

AND2x2_ASAP7_75t_L g1635 ( 
.A(n_1594),
.B(n_1586),
.Y(n_1635)
);

INVx1_ASAP7_75t_L g1636 ( 
.A(n_1603),
.Y(n_1636)
);

INVxp67_ASAP7_75t_L g1637 ( 
.A(n_1605),
.Y(n_1637)
);

AND2x2_ASAP7_75t_L g1638 ( 
.A(n_1594),
.B(n_1586),
.Y(n_1638)
);

AOI22xp33_ASAP7_75t_L g1639 ( 
.A1(n_1605),
.A2(n_1567),
.B1(n_1580),
.B2(n_1575),
.Y(n_1639)
);

NOR2xp33_ASAP7_75t_L g1640 ( 
.A(n_1610),
.B(n_1579),
.Y(n_1640)
);

AND2x2_ASAP7_75t_L g1641 ( 
.A(n_1594),
.B(n_1565),
.Y(n_1641)
);

AND2x2_ASAP7_75t_L g1642 ( 
.A(n_1602),
.B(n_1565),
.Y(n_1642)
);

OR2x2_ASAP7_75t_L g1643 ( 
.A(n_1602),
.B(n_1570),
.Y(n_1643)
);

NAND2xp5_ASAP7_75t_L g1644 ( 
.A(n_1602),
.B(n_1570),
.Y(n_1644)
);

OR2x2_ASAP7_75t_L g1645 ( 
.A(n_1607),
.B(n_1563),
.Y(n_1645)
);

AND2x2_ASAP7_75t_L g1646 ( 
.A(n_1607),
.B(n_1565),
.Y(n_1646)
);

AND2x2_ASAP7_75t_L g1647 ( 
.A(n_1607),
.B(n_1565),
.Y(n_1647)
);

BUFx3_ASAP7_75t_L g1648 ( 
.A(n_1631),
.Y(n_1648)
);

NAND2xp5_ASAP7_75t_L g1649 ( 
.A(n_1637),
.B(n_1630),
.Y(n_1649)
);

NAND2xp5_ASAP7_75t_L g1650 ( 
.A(n_1637),
.B(n_1611),
.Y(n_1650)
);

AND2x2_ASAP7_75t_L g1651 ( 
.A(n_1625),
.B(n_1611),
.Y(n_1651)
);

INVx1_ASAP7_75t_L g1652 ( 
.A(n_1626),
.Y(n_1652)
);

INVx1_ASAP7_75t_L g1653 ( 
.A(n_1626),
.Y(n_1653)
);

OR2x2_ASAP7_75t_L g1654 ( 
.A(n_1633),
.B(n_1618),
.Y(n_1654)
);

INVxp67_ASAP7_75t_SL g1655 ( 
.A(n_1631),
.Y(n_1655)
);

INVx2_ASAP7_75t_L g1656 ( 
.A(n_1630),
.Y(n_1656)
);

INVx1_ASAP7_75t_L g1657 ( 
.A(n_1628),
.Y(n_1657)
);

INVx1_ASAP7_75t_L g1658 ( 
.A(n_1628),
.Y(n_1658)
);

NAND2xp5_ASAP7_75t_L g1659 ( 
.A(n_1636),
.B(n_1611),
.Y(n_1659)
);

INVx1_ASAP7_75t_L g1660 ( 
.A(n_1617),
.Y(n_1660)
);

NAND2xp5_ASAP7_75t_L g1661 ( 
.A(n_1636),
.B(n_1614),
.Y(n_1661)
);

NOR2xp33_ASAP7_75t_L g1662 ( 
.A(n_1640),
.B(n_1579),
.Y(n_1662)
);

OR2x2_ASAP7_75t_L g1663 ( 
.A(n_1633),
.B(n_1577),
.Y(n_1663)
);

NAND2xp5_ASAP7_75t_L g1664 ( 
.A(n_1634),
.B(n_1614),
.Y(n_1664)
);

OR2x2_ASAP7_75t_L g1665 ( 
.A(n_1618),
.B(n_1577),
.Y(n_1665)
);

INVx2_ASAP7_75t_L g1666 ( 
.A(n_1619),
.Y(n_1666)
);

CKINVDCx20_ASAP7_75t_R g1667 ( 
.A(n_1634),
.Y(n_1667)
);

INVx2_ASAP7_75t_L g1668 ( 
.A(n_1619),
.Y(n_1668)
);

INVx1_ASAP7_75t_L g1669 ( 
.A(n_1617),
.Y(n_1669)
);

OR2x2_ASAP7_75t_L g1670 ( 
.A(n_1621),
.B(n_1577),
.Y(n_1670)
);

AND2x2_ASAP7_75t_L g1671 ( 
.A(n_1625),
.B(n_1597),
.Y(n_1671)
);

INVx2_ASAP7_75t_L g1672 ( 
.A(n_1619),
.Y(n_1672)
);

OAI21xp5_ASAP7_75t_L g1673 ( 
.A1(n_1639),
.A2(n_1588),
.B(n_1606),
.Y(n_1673)
);

AND2x2_ASAP7_75t_L g1674 ( 
.A(n_1625),
.B(n_1597),
.Y(n_1674)
);

INVx2_ASAP7_75t_SL g1675 ( 
.A(n_1627),
.Y(n_1675)
);

OAI22xp33_ASAP7_75t_L g1676 ( 
.A1(n_1620),
.A2(n_1606),
.B1(n_1588),
.B2(n_1572),
.Y(n_1676)
);

INVx2_ASAP7_75t_L g1677 ( 
.A(n_1624),
.Y(n_1677)
);

AND2x4_ASAP7_75t_L g1678 ( 
.A(n_1627),
.B(n_1590),
.Y(n_1678)
);

OR2x2_ASAP7_75t_L g1679 ( 
.A(n_1621),
.B(n_1577),
.Y(n_1679)
);

INVx1_ASAP7_75t_L g1680 ( 
.A(n_1622),
.Y(n_1680)
);

OAI21xp5_ASAP7_75t_L g1681 ( 
.A1(n_1639),
.A2(n_1610),
.B(n_1572),
.Y(n_1681)
);

INVx1_ASAP7_75t_L g1682 ( 
.A(n_1622),
.Y(n_1682)
);

INVx1_ASAP7_75t_SL g1683 ( 
.A(n_1615),
.Y(n_1683)
);

AND2x4_ASAP7_75t_L g1684 ( 
.A(n_1627),
.B(n_1590),
.Y(n_1684)
);

OR2x2_ASAP7_75t_L g1685 ( 
.A(n_1632),
.B(n_1612),
.Y(n_1685)
);

AND2x2_ASAP7_75t_L g1686 ( 
.A(n_1616),
.B(n_1612),
.Y(n_1686)
);

AOI32xp33_ASAP7_75t_L g1687 ( 
.A1(n_1616),
.A2(n_1612),
.A3(n_1572),
.B1(n_1566),
.B2(n_1598),
.Y(n_1687)
);

INVxp33_ASAP7_75t_SL g1688 ( 
.A(n_1615),
.Y(n_1688)
);

AND2x2_ASAP7_75t_L g1689 ( 
.A(n_1616),
.B(n_1591),
.Y(n_1689)
);

INVx1_ASAP7_75t_L g1690 ( 
.A(n_1623),
.Y(n_1690)
);

INVx1_ASAP7_75t_L g1691 ( 
.A(n_1652),
.Y(n_1691)
);

INVx1_ASAP7_75t_SL g1692 ( 
.A(n_1656),
.Y(n_1692)
);

INVx1_ASAP7_75t_L g1693 ( 
.A(n_1652),
.Y(n_1693)
);

INVx1_ASAP7_75t_L g1694 ( 
.A(n_1660),
.Y(n_1694)
);

INVx1_ASAP7_75t_L g1695 ( 
.A(n_1660),
.Y(n_1695)
);

INVx1_ASAP7_75t_L g1696 ( 
.A(n_1680),
.Y(n_1696)
);

INVx2_ASAP7_75t_L g1697 ( 
.A(n_1671),
.Y(n_1697)
);

NOR2xp33_ASAP7_75t_L g1698 ( 
.A(n_1649),
.B(n_1673),
.Y(n_1698)
);

INVx2_ASAP7_75t_L g1699 ( 
.A(n_1671),
.Y(n_1699)
);

OR2x2_ASAP7_75t_L g1700 ( 
.A(n_1650),
.B(n_1664),
.Y(n_1700)
);

INVx1_ASAP7_75t_L g1701 ( 
.A(n_1680),
.Y(n_1701)
);

INVx1_ASAP7_75t_L g1702 ( 
.A(n_1690),
.Y(n_1702)
);

OR2x2_ASAP7_75t_L g1703 ( 
.A(n_1654),
.B(n_1632),
.Y(n_1703)
);

OR2x2_ASAP7_75t_L g1704 ( 
.A(n_1654),
.B(n_1620),
.Y(n_1704)
);

INVx1_ASAP7_75t_SL g1705 ( 
.A(n_1656),
.Y(n_1705)
);

OR2x2_ASAP7_75t_L g1706 ( 
.A(n_1685),
.B(n_1663),
.Y(n_1706)
);

AND2x2_ASAP7_75t_L g1707 ( 
.A(n_1689),
.B(n_1641),
.Y(n_1707)
);

NAND2xp5_ASAP7_75t_SL g1708 ( 
.A(n_1676),
.B(n_1579),
.Y(n_1708)
);

NAND2xp5_ASAP7_75t_L g1709 ( 
.A(n_1655),
.B(n_1644),
.Y(n_1709)
);

OAI21xp5_ASAP7_75t_L g1710 ( 
.A1(n_1681),
.A2(n_1667),
.B(n_1688),
.Y(n_1710)
);

NAND2xp5_ASAP7_75t_L g1711 ( 
.A(n_1653),
.B(n_1657),
.Y(n_1711)
);

AND2x4_ASAP7_75t_L g1712 ( 
.A(n_1689),
.B(n_1627),
.Y(n_1712)
);

XNOR2xp5_ASAP7_75t_L g1713 ( 
.A(n_1667),
.B(n_1532),
.Y(n_1713)
);

NAND2xp33_ASAP7_75t_L g1714 ( 
.A(n_1683),
.B(n_1534),
.Y(n_1714)
);

INVx2_ASAP7_75t_L g1715 ( 
.A(n_1674),
.Y(n_1715)
);

OR2x2_ASAP7_75t_L g1716 ( 
.A(n_1685),
.B(n_1620),
.Y(n_1716)
);

NAND2xp5_ASAP7_75t_SL g1717 ( 
.A(n_1688),
.B(n_1579),
.Y(n_1717)
);

NAND2xp5_ASAP7_75t_L g1718 ( 
.A(n_1658),
.B(n_1644),
.Y(n_1718)
);

INVx1_ASAP7_75t_L g1719 ( 
.A(n_1690),
.Y(n_1719)
);

OR2x2_ASAP7_75t_L g1720 ( 
.A(n_1663),
.B(n_1665),
.Y(n_1720)
);

INVx2_ASAP7_75t_L g1721 ( 
.A(n_1674),
.Y(n_1721)
);

NOR2xp33_ASAP7_75t_L g1722 ( 
.A(n_1662),
.B(n_1579),
.Y(n_1722)
);

NAND2xp5_ASAP7_75t_L g1723 ( 
.A(n_1648),
.B(n_1643),
.Y(n_1723)
);

INVx1_ASAP7_75t_L g1724 ( 
.A(n_1669),
.Y(n_1724)
);

NAND2xp5_ASAP7_75t_L g1725 ( 
.A(n_1648),
.B(n_1643),
.Y(n_1725)
);

INVx1_ASAP7_75t_L g1726 ( 
.A(n_1682),
.Y(n_1726)
);

INVx2_ASAP7_75t_L g1727 ( 
.A(n_1666),
.Y(n_1727)
);

NOR4xp25_ASAP7_75t_SL g1728 ( 
.A(n_1708),
.B(n_1629),
.C(n_1623),
.D(n_1687),
.Y(n_1728)
);

INVx1_ASAP7_75t_L g1729 ( 
.A(n_1694),
.Y(n_1729)
);

OAI211xp5_ASAP7_75t_SL g1730 ( 
.A1(n_1710),
.A2(n_1708),
.B(n_1698),
.C(n_1714),
.Y(n_1730)
);

INVx3_ASAP7_75t_L g1731 ( 
.A(n_1712),
.Y(n_1731)
);

NOR2xp33_ASAP7_75t_L g1732 ( 
.A(n_1698),
.B(n_1477),
.Y(n_1732)
);

AND2x2_ASAP7_75t_L g1733 ( 
.A(n_1712),
.B(n_1686),
.Y(n_1733)
);

OR2x2_ASAP7_75t_L g1734 ( 
.A(n_1700),
.B(n_1686),
.Y(n_1734)
);

INVx1_ASAP7_75t_L g1735 ( 
.A(n_1695),
.Y(n_1735)
);

INVx1_ASAP7_75t_L g1736 ( 
.A(n_1696),
.Y(n_1736)
);

NAND2xp5_ASAP7_75t_L g1737 ( 
.A(n_1692),
.B(n_1635),
.Y(n_1737)
);

NAND2x1_ASAP7_75t_L g1738 ( 
.A(n_1712),
.B(n_1675),
.Y(n_1738)
);

INVx1_ASAP7_75t_L g1739 ( 
.A(n_1701),
.Y(n_1739)
);

NOR2xp33_ASAP7_75t_L g1740 ( 
.A(n_1705),
.B(n_1477),
.Y(n_1740)
);

OAI222xp33_ASAP7_75t_L g1741 ( 
.A1(n_1713),
.A2(n_1580),
.B1(n_1651),
.B2(n_1643),
.C1(n_1645),
.C2(n_1659),
.Y(n_1741)
);

OAI22xp33_ASAP7_75t_SL g1742 ( 
.A1(n_1704),
.A2(n_1645),
.B1(n_1675),
.B2(n_1600),
.Y(n_1742)
);

INVx1_ASAP7_75t_L g1743 ( 
.A(n_1702),
.Y(n_1743)
);

NAND2xp5_ASAP7_75t_L g1744 ( 
.A(n_1697),
.B(n_1635),
.Y(n_1744)
);

INVxp67_ASAP7_75t_SL g1745 ( 
.A(n_1714),
.Y(n_1745)
);

INVx2_ASAP7_75t_L g1746 ( 
.A(n_1707),
.Y(n_1746)
);

AND2x4_ASAP7_75t_L g1747 ( 
.A(n_1697),
.B(n_1678),
.Y(n_1747)
);

INVx1_ASAP7_75t_L g1748 ( 
.A(n_1719),
.Y(n_1748)
);

O2A1O1Ixp33_ASAP7_75t_SL g1749 ( 
.A1(n_1717),
.A2(n_1661),
.B(n_1645),
.C(n_1585),
.Y(n_1749)
);

AOI221xp5_ASAP7_75t_L g1750 ( 
.A1(n_1709),
.A2(n_1672),
.B1(n_1666),
.B2(n_1668),
.C(n_1677),
.Y(n_1750)
);

HB1xp67_ASAP7_75t_L g1751 ( 
.A(n_1691),
.Y(n_1751)
);

INVxp67_ASAP7_75t_L g1752 ( 
.A(n_1693),
.Y(n_1752)
);

OAI21xp33_ASAP7_75t_L g1753 ( 
.A1(n_1723),
.A2(n_1670),
.B(n_1665),
.Y(n_1753)
);

AOI221xp5_ASAP7_75t_L g1754 ( 
.A1(n_1741),
.A2(n_1718),
.B1(n_1725),
.B2(n_1726),
.C(n_1724),
.Y(n_1754)
);

O2A1O1Ixp33_ASAP7_75t_L g1755 ( 
.A1(n_1730),
.A2(n_1711),
.B(n_1717),
.C(n_1704),
.Y(n_1755)
);

INVx1_ASAP7_75t_L g1756 ( 
.A(n_1751),
.Y(n_1756)
);

AOI211xp5_ASAP7_75t_L g1757 ( 
.A1(n_1745),
.A2(n_1722),
.B(n_1707),
.C(n_1716),
.Y(n_1757)
);

NAND2xp5_ASAP7_75t_L g1758 ( 
.A(n_1746),
.B(n_1699),
.Y(n_1758)
);

AOI21xp5_ASAP7_75t_L g1759 ( 
.A1(n_1728),
.A2(n_1722),
.B(n_1715),
.Y(n_1759)
);

NAND2xp33_ASAP7_75t_SL g1760 ( 
.A(n_1738),
.B(n_1699),
.Y(n_1760)
);

AOI211xp5_ASAP7_75t_L g1761 ( 
.A1(n_1745),
.A2(n_1706),
.B(n_1703),
.C(n_1715),
.Y(n_1761)
);

INVx1_ASAP7_75t_L g1762 ( 
.A(n_1751),
.Y(n_1762)
);

O2A1O1Ixp33_ASAP7_75t_L g1763 ( 
.A1(n_1752),
.A2(n_1703),
.B(n_1727),
.C(n_1721),
.Y(n_1763)
);

INVx1_ASAP7_75t_L g1764 ( 
.A(n_1729),
.Y(n_1764)
);

NAND2xp5_ASAP7_75t_L g1765 ( 
.A(n_1734),
.B(n_1721),
.Y(n_1765)
);

INVx1_ASAP7_75t_L g1766 ( 
.A(n_1735),
.Y(n_1766)
);

INVx1_ASAP7_75t_L g1767 ( 
.A(n_1736),
.Y(n_1767)
);

NAND2xp5_ASAP7_75t_L g1768 ( 
.A(n_1731),
.B(n_1706),
.Y(n_1768)
);

NAND3xp33_ASAP7_75t_SL g1769 ( 
.A(n_1732),
.B(n_1520),
.C(n_1720),
.Y(n_1769)
);

INVx1_ASAP7_75t_L g1770 ( 
.A(n_1739),
.Y(n_1770)
);

INVx1_ASAP7_75t_L g1771 ( 
.A(n_1743),
.Y(n_1771)
);

NOR2xp33_ASAP7_75t_L g1772 ( 
.A(n_1732),
.B(n_1678),
.Y(n_1772)
);

OAI21xp5_ASAP7_75t_L g1773 ( 
.A1(n_1752),
.A2(n_1727),
.B(n_1642),
.Y(n_1773)
);

INVx1_ASAP7_75t_L g1774 ( 
.A(n_1768),
.Y(n_1774)
);

O2A1O1Ixp33_ASAP7_75t_L g1775 ( 
.A1(n_1755),
.A2(n_1742),
.B(n_1749),
.C(n_1748),
.Y(n_1775)
);

AND2x2_ASAP7_75t_L g1776 ( 
.A(n_1772),
.B(n_1731),
.Y(n_1776)
);

INVx1_ASAP7_75t_L g1777 ( 
.A(n_1756),
.Y(n_1777)
);

NAND2xp5_ASAP7_75t_SL g1778 ( 
.A(n_1761),
.B(n_1740),
.Y(n_1778)
);

INVxp67_ASAP7_75t_SL g1779 ( 
.A(n_1762),
.Y(n_1779)
);

NAND2xp5_ASAP7_75t_L g1780 ( 
.A(n_1757),
.B(n_1765),
.Y(n_1780)
);

INVx1_ASAP7_75t_L g1781 ( 
.A(n_1758),
.Y(n_1781)
);

INVxp67_ASAP7_75t_L g1782 ( 
.A(n_1772),
.Y(n_1782)
);

INVx1_ASAP7_75t_L g1783 ( 
.A(n_1764),
.Y(n_1783)
);

INVx1_ASAP7_75t_L g1784 ( 
.A(n_1766),
.Y(n_1784)
);

NAND3xp33_ASAP7_75t_L g1785 ( 
.A(n_1754),
.B(n_1750),
.C(n_1740),
.Y(n_1785)
);

INVx1_ASAP7_75t_L g1786 ( 
.A(n_1767),
.Y(n_1786)
);

NAND2xp5_ASAP7_75t_L g1787 ( 
.A(n_1782),
.B(n_1763),
.Y(n_1787)
);

NAND3xp33_ASAP7_75t_L g1788 ( 
.A(n_1778),
.B(n_1760),
.C(n_1759),
.Y(n_1788)
);

NAND2xp5_ASAP7_75t_L g1789 ( 
.A(n_1781),
.B(n_1747),
.Y(n_1789)
);

BUFx2_ASAP7_75t_L g1790 ( 
.A(n_1776),
.Y(n_1790)
);

NAND4xp25_ASAP7_75t_L g1791 ( 
.A(n_1775),
.B(n_1760),
.C(n_1769),
.D(n_1770),
.Y(n_1791)
);

NAND2xp5_ASAP7_75t_L g1792 ( 
.A(n_1774),
.B(n_1747),
.Y(n_1792)
);

NOR4xp25_ASAP7_75t_SL g1793 ( 
.A(n_1778),
.B(n_1771),
.C(n_1753),
.D(n_1773),
.Y(n_1793)
);

NAND2xp5_ASAP7_75t_L g1794 ( 
.A(n_1779),
.B(n_1733),
.Y(n_1794)
);

OAI211xp5_ASAP7_75t_L g1795 ( 
.A1(n_1780),
.A2(n_1737),
.B(n_1744),
.C(n_1651),
.Y(n_1795)
);

NAND3xp33_ASAP7_75t_L g1796 ( 
.A(n_1785),
.B(n_1779),
.C(n_1777),
.Y(n_1796)
);

AND4x1_ASAP7_75t_L g1797 ( 
.A(n_1796),
.B(n_1786),
.C(n_1784),
.D(n_1783),
.Y(n_1797)
);

AOI221xp5_ASAP7_75t_L g1798 ( 
.A1(n_1788),
.A2(n_1677),
.B1(n_1672),
.B2(n_1668),
.C(n_1642),
.Y(n_1798)
);

AOI221xp5_ASAP7_75t_L g1799 ( 
.A1(n_1791),
.A2(n_1641),
.B1(n_1647),
.B2(n_1642),
.C(n_1646),
.Y(n_1799)
);

AOI222xp33_ASAP7_75t_L g1800 ( 
.A1(n_1787),
.A2(n_1641),
.B1(n_1647),
.B2(n_1646),
.C1(n_1560),
.C2(n_1559),
.Y(n_1800)
);

NOR2xp33_ASAP7_75t_L g1801 ( 
.A(n_1790),
.B(n_1629),
.Y(n_1801)
);

HB1xp67_ASAP7_75t_L g1802 ( 
.A(n_1797),
.Y(n_1802)
);

OAI21xp5_ASAP7_75t_L g1803 ( 
.A1(n_1801),
.A2(n_1794),
.B(n_1792),
.Y(n_1803)
);

AOI211x1_ASAP7_75t_SL g1804 ( 
.A1(n_1798),
.A2(n_1789),
.B(n_1793),
.C(n_1795),
.Y(n_1804)
);

AOI221xp5_ASAP7_75t_L g1805 ( 
.A1(n_1799),
.A2(n_1646),
.B1(n_1647),
.B2(n_1600),
.C(n_1613),
.Y(n_1805)
);

OAI211xp5_ASAP7_75t_L g1806 ( 
.A1(n_1800),
.A2(n_1635),
.B(n_1638),
.C(n_1670),
.Y(n_1806)
);

AOI221xp5_ASAP7_75t_L g1807 ( 
.A1(n_1798),
.A2(n_1600),
.B1(n_1601),
.B2(n_1599),
.C(n_1598),
.Y(n_1807)
);

NAND4xp75_ASAP7_75t_L g1808 ( 
.A(n_1803),
.B(n_1452),
.C(n_1638),
.D(n_1514),
.Y(n_1808)
);

INVx2_ASAP7_75t_L g1809 ( 
.A(n_1802),
.Y(n_1809)
);

AOI22xp5_ASAP7_75t_L g1810 ( 
.A1(n_1806),
.A2(n_1522),
.B1(n_1684),
.B2(n_1678),
.Y(n_1810)
);

NAND4xp75_ASAP7_75t_L g1811 ( 
.A(n_1804),
.B(n_1452),
.C(n_1638),
.D(n_1609),
.Y(n_1811)
);

NAND3xp33_ASAP7_75t_L g1812 ( 
.A(n_1805),
.B(n_1452),
.C(n_1679),
.Y(n_1812)
);

NAND3xp33_ASAP7_75t_L g1813 ( 
.A(n_1809),
.B(n_1810),
.C(n_1812),
.Y(n_1813)
);

NAND2xp5_ASAP7_75t_L g1814 ( 
.A(n_1811),
.B(n_1807),
.Y(n_1814)
);

NAND3xp33_ASAP7_75t_L g1815 ( 
.A(n_1808),
.B(n_1452),
.C(n_1684),
.Y(n_1815)
);

INVx4_ASAP7_75t_L g1816 ( 
.A(n_1813),
.Y(n_1816)
);

INVx1_ASAP7_75t_L g1817 ( 
.A(n_1816),
.Y(n_1817)
);

HB1xp67_ASAP7_75t_L g1818 ( 
.A(n_1817),
.Y(n_1818)
);

AOI21xp5_ASAP7_75t_L g1819 ( 
.A1(n_1817),
.A2(n_1814),
.B(n_1815),
.Y(n_1819)
);

CKINVDCx20_ASAP7_75t_R g1820 ( 
.A(n_1818),
.Y(n_1820)
);

INVx1_ASAP7_75t_L g1821 ( 
.A(n_1819),
.Y(n_1821)
);

INVx1_ASAP7_75t_L g1822 ( 
.A(n_1820),
.Y(n_1822)
);

NAND2xp5_ASAP7_75t_L g1823 ( 
.A(n_1821),
.B(n_1624),
.Y(n_1823)
);

NAND2xp5_ASAP7_75t_L g1824 ( 
.A(n_1822),
.B(n_1522),
.Y(n_1824)
);

OAI21xp5_ASAP7_75t_L g1825 ( 
.A1(n_1824),
.A2(n_1823),
.B(n_1684),
.Y(n_1825)
);

XNOR2xp5_ASAP7_75t_L g1826 ( 
.A(n_1825),
.B(n_1487),
.Y(n_1826)
);

OAI221xp5_ASAP7_75t_R g1827 ( 
.A1(n_1826),
.A2(n_1470),
.B1(n_1679),
.B2(n_1525),
.C(n_1591),
.Y(n_1827)
);

AOI211xp5_ASAP7_75t_L g1828 ( 
.A1(n_1827),
.A2(n_1487),
.B(n_1509),
.C(n_1515),
.Y(n_1828)
);


endmodule