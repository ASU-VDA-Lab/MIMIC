module fake_jpeg_24178_n_47 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_47);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;

output n_47;

wire n_13;
wire n_21;
wire n_33;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_22;
wire n_14;
wire n_40;
wire n_19;
wire n_20;
wire n_18;
wire n_35;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_43;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

BUFx12f_ASAP7_75t_L g7 ( 
.A(n_0),
.Y(n_7)
);

INVx2_ASAP7_75t_L g8 ( 
.A(n_0),
.Y(n_8)
);

INVx3_ASAP7_75t_L g9 ( 
.A(n_1),
.Y(n_9)
);

INVx2_ASAP7_75t_L g10 ( 
.A(n_3),
.Y(n_10)
);

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_1),
.Y(n_11)
);

BUFx6f_ASAP7_75t_L g12 ( 
.A(n_3),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_6),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_L g14 ( 
.A(n_5),
.B(n_2),
.Y(n_14)
);

INVx6_ASAP7_75t_L g15 ( 
.A(n_2),
.Y(n_15)
);

AOI21xp5_ASAP7_75t_L g16 ( 
.A1(n_8),
.A2(n_4),
.B(n_5),
.Y(n_16)
);

AOI21xp5_ASAP7_75t_L g24 ( 
.A1(n_16),
.A2(n_15),
.B(n_21),
.Y(n_24)
);

INVx6_ASAP7_75t_L g17 ( 
.A(n_12),
.Y(n_17)
);

AOI22xp33_ASAP7_75t_L g23 ( 
.A1(n_17),
.A2(n_15),
.B1(n_10),
.B2(n_13),
.Y(n_23)
);

INVx8_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

AOI21xp33_ASAP7_75t_SL g19 ( 
.A1(n_7),
.A2(n_4),
.B(n_6),
.Y(n_19)
);

A2O1A1O1Ixp25_ASAP7_75t_L g26 ( 
.A1(n_19),
.A2(n_7),
.B(n_21),
.C(n_16),
.D(n_14),
.Y(n_26)
);

OR2x2_ASAP7_75t_L g20 ( 
.A(n_11),
.B(n_7),
.Y(n_20)
);

XNOR2xp5_ASAP7_75t_SL g28 ( 
.A(n_20),
.B(n_21),
.Y(n_28)
);

OR2x2_ASAP7_75t_L g21 ( 
.A(n_14),
.B(n_9),
.Y(n_21)
);

INVx13_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_22),
.Y(n_30)
);

XNOR2xp5_ASAP7_75t_L g35 ( 
.A(n_24),
.B(n_25),
.Y(n_35)
);

AOI21xp5_ASAP7_75t_L g25 ( 
.A1(n_16),
.A2(n_20),
.B(n_22),
.Y(n_25)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_26),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_SL g27 ( 
.A(n_17),
.B(n_18),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_27),
.B(n_29),
.Y(n_33)
);

XNOR2xp5_ASAP7_75t_L g29 ( 
.A(n_21),
.B(n_16),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_30),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_31),
.Y(n_36)
);

CKINVDCx5p33_ASAP7_75t_R g32 ( 
.A(n_30),
.Y(n_32)
);

CKINVDCx16_ASAP7_75t_R g37 ( 
.A(n_32),
.Y(n_37)
);

MAJx2_ASAP7_75t_L g38 ( 
.A(n_35),
.B(n_28),
.C(n_23),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_38),
.B(n_35),
.Y(n_40)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_36),
.Y(n_39)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_39),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_L g42 ( 
.A1(n_40),
.A2(n_41),
.B1(n_34),
.B2(n_33),
.Y(n_42)
);

CKINVDCx5p33_ASAP7_75t_R g41 ( 
.A(n_37),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_SL g44 ( 
.A(n_42),
.B(n_38),
.Y(n_44)
);

MAJIxp5_ASAP7_75t_L g45 ( 
.A(n_44),
.B(n_43),
.C(n_41),
.Y(n_45)
);

XNOR2xp5_ASAP7_75t_L g46 ( 
.A(n_45),
.B(n_43),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_46),
.B(n_32),
.Y(n_47)
);


endmodule