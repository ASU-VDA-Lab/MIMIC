module fake_jpeg_15976_n_93 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_93);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_93;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_22;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;

INVx2_ASAP7_75t_L g12 ( 
.A(n_1),
.Y(n_12)
);

NOR2xp33_ASAP7_75t_L g13 ( 
.A(n_11),
.B(n_10),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_4),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_5),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_7),
.B(n_6),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_3),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_1),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_18),
.Y(n_23)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_23),
.Y(n_47)
);

OR2x2_ASAP7_75t_L g24 ( 
.A(n_12),
.B(n_0),
.Y(n_24)
);

INVx1_ASAP7_75t_SL g46 ( 
.A(n_24),
.Y(n_46)
);

INVx8_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_25),
.Y(n_44)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_21),
.Y(n_26)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_26),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_21),
.B(n_0),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_SL g36 ( 
.A(n_27),
.B(n_22),
.Y(n_36)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_20),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_28),
.B(n_32),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_L g29 ( 
.A1(n_14),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_29)
);

AOI22xp5_ASAP7_75t_L g34 ( 
.A1(n_29),
.A2(n_19),
.B1(n_22),
.B2(n_14),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_SL g30 ( 
.A(n_18),
.B(n_2),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_SL g50 ( 
.A(n_30),
.B(n_31),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_15),
.Y(n_31)
);

BUFx2_ASAP7_75t_L g32 ( 
.A(n_20),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_17),
.Y(n_33)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_33),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_L g52 ( 
.A1(n_34),
.A2(n_37),
.B1(n_41),
.B2(n_51),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_36),
.B(n_32),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_L g37 ( 
.A1(n_33),
.A2(n_19),
.B1(n_15),
.B2(n_17),
.Y(n_37)
);

INVxp67_ASAP7_75t_L g38 ( 
.A(n_26),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_38),
.B(n_48),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g40 ( 
.A1(n_28),
.A2(n_2),
.B1(n_3),
.B2(n_6),
.Y(n_40)
);

INVxp67_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g41 ( 
.A1(n_25),
.A2(n_3),
.B1(n_8),
.B2(n_9),
.Y(n_41)
);

XNOR2xp5_ASAP7_75t_L g42 ( 
.A(n_27),
.B(n_13),
.Y(n_42)
);

XOR2xp5_ASAP7_75t_L g64 ( 
.A(n_42),
.B(n_43),
.Y(n_64)
);

XOR2xp5_ASAP7_75t_L g43 ( 
.A(n_24),
.B(n_16),
.Y(n_43)
);

OAI21xp5_ASAP7_75t_SL g45 ( 
.A1(n_24),
.A2(n_8),
.B(n_9),
.Y(n_45)
);

MAJIxp5_ASAP7_75t_L g56 ( 
.A(n_45),
.B(n_30),
.C(n_31),
.Y(n_56)
);

FAx1_ASAP7_75t_SL g48 ( 
.A(n_24),
.B(n_10),
.CI(n_11),
.CON(n_48),
.SN(n_48)
);

AOI22xp5_ASAP7_75t_L g51 ( 
.A1(n_25),
.A2(n_29),
.B1(n_28),
.B2(n_23),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_47),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_54),
.B(n_55),
.Y(n_65)
);

CKINVDCx16_ASAP7_75t_R g55 ( 
.A(n_47),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_56),
.B(n_61),
.Y(n_67)
);

INVx2_ASAP7_75t_SL g57 ( 
.A(n_44),
.Y(n_57)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_57),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g58 ( 
.A1(n_46),
.A2(n_32),
.B1(n_51),
.B2(n_49),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_58),
.A2(n_44),
.B1(n_41),
.B2(n_38),
.Y(n_69)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_35),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_59),
.Y(n_74)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_39),
.Y(n_61)
);

MAJIxp5_ASAP7_75t_L g62 ( 
.A(n_43),
.B(n_32),
.C(n_42),
.Y(n_62)
);

MAJIxp5_ASAP7_75t_L g72 ( 
.A(n_62),
.B(n_64),
.C(n_56),
.Y(n_72)
);

XOR2xp5_ASAP7_75t_L g70 ( 
.A(n_63),
.B(n_48),
.Y(n_70)
);

AOI21xp5_ASAP7_75t_L g68 ( 
.A1(n_53),
.A2(n_45),
.B(n_46),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_68),
.A2(n_53),
.B1(n_52),
.B2(n_34),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_69),
.A2(n_57),
.B1(n_73),
.B2(n_67),
.Y(n_81)
);

XNOR2xp5_ASAP7_75t_L g75 ( 
.A(n_70),
.B(n_60),
.Y(n_75)
);

XOR2xp5_ASAP7_75t_L g71 ( 
.A(n_64),
.B(n_48),
.Y(n_71)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_71),
.B(n_72),
.C(n_73),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g73 ( 
.A(n_62),
.B(n_63),
.C(n_58),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_75),
.B(n_80),
.Y(n_86)
);

CKINVDCx16_ASAP7_75t_R g76 ( 
.A(n_65),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_76),
.B(n_80),
.Y(n_83)
);

AOI21xp5_ASAP7_75t_L g84 ( 
.A1(n_78),
.A2(n_71),
.B(n_70),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_74),
.B(n_50),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_79),
.B(n_66),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_72),
.B(n_52),
.C(n_57),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_81),
.B(n_69),
.Y(n_82)
);

AO21x1_ASAP7_75t_L g90 ( 
.A1(n_82),
.A2(n_86),
.B(n_77),
.Y(n_90)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_84),
.Y(n_88)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_85),
.Y(n_89)
);

AOI21xp5_ASAP7_75t_L g87 ( 
.A1(n_83),
.A2(n_75),
.B(n_77),
.Y(n_87)
);

AO21x1_ASAP7_75t_L g91 ( 
.A1(n_87),
.A2(n_90),
.B(n_88),
.Y(n_91)
);

AOI21xp5_ASAP7_75t_L g93 ( 
.A1(n_91),
.A2(n_92),
.B(n_90),
.Y(n_93)
);

HB1xp67_ASAP7_75t_L g92 ( 
.A(n_89),
.Y(n_92)
);


endmodule