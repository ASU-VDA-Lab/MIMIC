module fake_jpeg_17134_n_74 (n_13, n_21, n_1, n_10, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_74);

input n_13;
input n_21;
input n_1;
input n_10;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_74;

wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_23;
wire n_69;
wire n_27;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_40;
wire n_73;
wire n_59;
wire n_35;
wire n_48;
wire n_68;
wire n_52;
wire n_71;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_65;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_72;
wire n_24;
wire n_28;
wire n_44;
wire n_26;
wire n_38;
wire n_36;
wire n_62;
wire n_31;
wire n_25;
wire n_67;
wire n_56;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_32;
wire n_70;
wire n_66;

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_8),
.B(n_9),
.Y(n_23)
);

INVx11_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_11),
.Y(n_25)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_17),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_13),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_1),
.Y(n_30)
);

INVx5_ASAP7_75t_L g31 ( 
.A(n_24),
.Y(n_31)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_31),
.Y(n_45)
);

NAND3xp33_ASAP7_75t_L g32 ( 
.A(n_30),
.B(n_0),
.C(n_2),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_32),
.B(n_4),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_29),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_33),
.B(n_34),
.Y(n_38)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_29),
.Y(n_34)
);

NOR3xp33_ASAP7_75t_L g35 ( 
.A(n_30),
.B(n_15),
.C(n_22),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_35),
.B(n_37),
.Y(n_41)
);

MAJIxp5_ASAP7_75t_L g36 ( 
.A(n_25),
.B(n_0),
.C(n_3),
.Y(n_36)
);

MAJIxp5_ASAP7_75t_L g40 ( 
.A(n_36),
.B(n_27),
.C(n_5),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_25),
.B(n_3),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_L g39 ( 
.A1(n_32),
.A2(n_26),
.B1(n_27),
.B2(n_6),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_L g48 ( 
.A1(n_39),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_40),
.B(n_46),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_35),
.B(n_28),
.Y(n_42)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_42),
.Y(n_50)
);

MAJx2_ASAP7_75t_L g43 ( 
.A(n_32),
.B(n_26),
.C(n_19),
.Y(n_43)
);

MAJIxp5_ASAP7_75t_L g47 ( 
.A(n_43),
.B(n_23),
.C(n_24),
.Y(n_47)
);

INVx11_ASAP7_75t_L g44 ( 
.A(n_31),
.Y(n_44)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_44),
.Y(n_51)
);

AND2x2_ASAP7_75t_L g58 ( 
.A(n_47),
.B(n_48),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_38),
.B(n_10),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_49),
.B(n_52),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_41),
.B(n_12),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_45),
.Y(n_53)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_53),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_44),
.Y(n_55)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_55),
.Y(n_59)
);

INVx1_ASAP7_75t_SL g57 ( 
.A(n_51),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_57),
.B(n_60),
.Y(n_67)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_50),
.Y(n_60)
);

XNOR2xp5_ASAP7_75t_L g61 ( 
.A(n_54),
.B(n_40),
.Y(n_61)
);

MAJIxp5_ASAP7_75t_L g65 ( 
.A(n_61),
.B(n_62),
.C(n_63),
.Y(n_65)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_49),
.Y(n_62)
);

CKINVDCx16_ASAP7_75t_R g63 ( 
.A(n_47),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g66 ( 
.A1(n_58),
.A2(n_43),
.B1(n_16),
.B2(n_18),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_66),
.B(n_68),
.Y(n_69)
);

AOI21xp5_ASAP7_75t_SL g68 ( 
.A1(n_58),
.A2(n_14),
.B(n_20),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_69),
.Y(n_70)
);

MAJIxp5_ASAP7_75t_L g71 ( 
.A(n_70),
.B(n_67),
.C(n_59),
.Y(n_71)
);

MAJIxp5_ASAP7_75t_L g72 ( 
.A(n_71),
.B(n_64),
.C(n_56),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_L g73 ( 
.A1(n_72),
.A2(n_65),
.B1(n_60),
.B2(n_57),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_73),
.B(n_21),
.Y(n_74)
);


endmodule