module real_aes_1394_n_101 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_101);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_101;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_421;
wire n_364;
wire n_555;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_571;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_537;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_678;
wire n_548;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_815;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_816;
wire n_292;
wire n_539;
wire n_400;
wire n_626;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_781;
wire n_748;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_649;
wire n_651;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_455;
wire n_119;
wire n_504;
wire n_310;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_812;
wire n_817;
wire n_443;
wire n_565;
wire n_782;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_808;
wire n_770;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_527;
wire n_434;
wire n_502;
wire n_505;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_552;
wire n_402;
wire n_617;
wire n_733;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_807;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_785;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_810;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_749;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_765;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_809;
wire n_482;
wire n_633;
wire n_520;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_420;
wire n_336;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_753;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_521;
wire n_140;
wire n_418;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_103;
wire n_541;
wire n_224;
wire n_546;
wire n_151;
wire n_639;
wire n_587;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_710;
wire n_650;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_804;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_802;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_554;
wire n_475;
wire n_264;
wire n_798;
wire n_797;
wire n_237;
wire n_668;
NAND2xp5_ASAP7_75t_SL g198 ( .A(n_0), .B(n_141), .Y(n_198) );
AOI21xp5_ASAP7_75t_L g173 ( .A1(n_1), .A2(n_123), .B(n_174), .Y(n_173) );
NAND2xp5_ASAP7_75t_L g815 ( .A(n_2), .B(n_816), .Y(n_815) );
AOI22xp5_ASAP7_75t_L g804 ( .A1(n_3), .A2(n_11), .B1(n_805), .B2(n_806), .Y(n_804) );
CKINVDCx20_ASAP7_75t_R g806 ( .A(n_3), .Y(n_806) );
NAND2xp5_ASAP7_75t_SL g187 ( .A(n_4), .B(n_131), .Y(n_187) );
INVx1_ASAP7_75t_L g128 ( .A(n_5), .Y(n_128) );
NAND2xp5_ASAP7_75t_L g151 ( .A(n_6), .B(n_131), .Y(n_151) );
NAND2xp5_ASAP7_75t_SL g465 ( .A(n_7), .B(n_118), .Y(n_465) );
INVx1_ASAP7_75t_L g493 ( .A(n_8), .Y(n_493) );
CKINVDCx16_ASAP7_75t_R g816 ( .A(n_9), .Y(n_816) );
CKINVDCx5p33_ASAP7_75t_R g508 ( .A(n_10), .Y(n_508) );
CKINVDCx20_ASAP7_75t_R g805 ( .A(n_11), .Y(n_805) );
NAND2xp33_ASAP7_75t_L g168 ( .A(n_12), .B(n_135), .Y(n_168) );
INVx2_ASAP7_75t_L g120 ( .A(n_13), .Y(n_120) );
AOI221x1_ASAP7_75t_L g210 ( .A1(n_14), .A2(n_26), .B1(n_123), .B2(n_141), .C(n_211), .Y(n_210) );
CKINVDCx16_ASAP7_75t_R g431 ( .A(n_15), .Y(n_431) );
NAND2xp5_ASAP7_75t_SL g164 ( .A(n_16), .B(n_141), .Y(n_164) );
AO21x2_ASAP7_75t_L g161 ( .A1(n_17), .A2(n_162), .B(n_163), .Y(n_161) );
INVx1_ASAP7_75t_L g474 ( .A(n_18), .Y(n_474) );
NAND2xp5_ASAP7_75t_L g214 ( .A(n_19), .B(n_154), .Y(n_214) );
NAND2xp5_ASAP7_75t_L g130 ( .A(n_20), .B(n_131), .Y(n_130) );
AO21x1_ASAP7_75t_L g182 ( .A1(n_21), .A2(n_141), .B(n_183), .Y(n_182) );
INVx1_ASAP7_75t_L g434 ( .A(n_22), .Y(n_434) );
NOR2xp33_ASAP7_75t_SL g813 ( .A(n_22), .B(n_435), .Y(n_813) );
INVx1_ASAP7_75t_L g472 ( .A(n_23), .Y(n_472) );
INVx1_ASAP7_75t_SL g458 ( .A(n_24), .Y(n_458) );
NAND2xp5_ASAP7_75t_SL g552 ( .A(n_25), .B(n_142), .Y(n_552) );
NAND2x1_ASAP7_75t_L g196 ( .A(n_27), .B(n_131), .Y(n_196) );
AOI33xp33_ASAP7_75t_L g520 ( .A1(n_28), .A2(n_53), .A3(n_448), .B1(n_455), .B2(n_521), .B3(n_522), .Y(n_520) );
NAND2x1_ASAP7_75t_L g150 ( .A(n_29), .B(n_135), .Y(n_150) );
INVx1_ASAP7_75t_L g502 ( .A(n_30), .Y(n_502) );
OR2x2_ASAP7_75t_L g119 ( .A(n_31), .B(n_86), .Y(n_119) );
OA21x2_ASAP7_75t_L g159 ( .A1(n_31), .A2(n_86), .B(n_120), .Y(n_159) );
NAND2xp5_ASAP7_75t_L g445 ( .A(n_32), .B(n_446), .Y(n_445) );
NAND2xp5_ASAP7_75t_L g176 ( .A(n_33), .B(n_135), .Y(n_176) );
NAND2xp5_ASAP7_75t_L g167 ( .A(n_34), .B(n_131), .Y(n_167) );
NAND2xp5_ASAP7_75t_L g186 ( .A(n_35), .B(n_135), .Y(n_186) );
AOI21xp5_ASAP7_75t_L g228 ( .A1(n_36), .A2(n_123), .B(n_229), .Y(n_228) );
AND2x2_ASAP7_75t_L g124 ( .A(n_37), .B(n_125), .Y(n_124) );
AND2x2_ASAP7_75t_L g139 ( .A(n_37), .B(n_128), .Y(n_139) );
INVx1_ASAP7_75t_L g454 ( .A(n_37), .Y(n_454) );
OR2x6_ASAP7_75t_L g432 ( .A(n_38), .B(n_433), .Y(n_432) );
NOR3xp33_ASAP7_75t_L g814 ( .A(n_38), .B(n_431), .C(n_815), .Y(n_814) );
CKINVDCx20_ASAP7_75t_R g504 ( .A(n_39), .Y(n_504) );
NAND2xp5_ASAP7_75t_SL g232 ( .A(n_40), .B(n_141), .Y(n_232) );
NAND2xp5_ASAP7_75t_L g528 ( .A(n_41), .B(n_446), .Y(n_528) );
AOI22xp5_ASAP7_75t_L g545 ( .A1(n_42), .A2(n_118), .B1(n_158), .B2(n_546), .Y(n_545) );
NAND2xp5_ASAP7_75t_L g553 ( .A(n_43), .B(n_554), .Y(n_553) );
NAND2xp5_ASAP7_75t_L g460 ( .A(n_44), .B(n_142), .Y(n_460) );
INVxp33_ASAP7_75t_L g818 ( .A(n_45), .Y(n_818) );
CKINVDCx20_ASAP7_75t_R g144 ( .A(n_46), .Y(n_144) );
NAND2xp5_ASAP7_75t_L g230 ( .A(n_47), .B(n_135), .Y(n_230) );
NAND2xp5_ASAP7_75t_SL g495 ( .A(n_48), .B(n_162), .Y(n_495) );
NAND2xp5_ASAP7_75t_L g494 ( .A(n_49), .B(n_142), .Y(n_494) );
AOI21xp5_ASAP7_75t_L g148 ( .A1(n_50), .A2(n_123), .B(n_149), .Y(n_148) );
CKINVDCx5p33_ASAP7_75t_R g549 ( .A(n_51), .Y(n_549) );
NAND2xp5_ASAP7_75t_L g197 ( .A(n_52), .B(n_135), .Y(n_197) );
NAND2xp5_ASAP7_75t_L g532 ( .A(n_54), .B(n_142), .Y(n_532) );
INVx1_ASAP7_75t_L g127 ( .A(n_55), .Y(n_127) );
INVx1_ASAP7_75t_L g137 ( .A(n_55), .Y(n_137) );
AND2x2_ASAP7_75t_L g533 ( .A(n_56), .B(n_154), .Y(n_533) );
AOI221xp5_ASAP7_75t_L g491 ( .A1(n_57), .A2(n_75), .B1(n_446), .B2(n_452), .C(n_492), .Y(n_491) );
NAND2xp5_ASAP7_75t_L g486 ( .A(n_58), .B(n_446), .Y(n_486) );
NAND2xp5_ASAP7_75t_L g213 ( .A(n_59), .B(n_131), .Y(n_213) );
NAND2xp5_ASAP7_75t_L g510 ( .A(n_60), .B(n_158), .Y(n_510) );
CKINVDCx20_ASAP7_75t_R g796 ( .A(n_61), .Y(n_796) );
AOI21xp5_ASAP7_75t_SL g482 ( .A1(n_62), .A2(n_452), .B(n_483), .Y(n_482) );
AOI21xp5_ASAP7_75t_L g194 ( .A1(n_63), .A2(n_123), .B(n_195), .Y(n_194) );
INVx1_ASAP7_75t_L g468 ( .A(n_64), .Y(n_468) );
AO21x1_ASAP7_75t_L g184 ( .A1(n_65), .A2(n_123), .B(n_185), .Y(n_184) );
NAND2xp5_ASAP7_75t_SL g172 ( .A(n_66), .B(n_141), .Y(n_172) );
INVx1_ASAP7_75t_L g531 ( .A(n_67), .Y(n_531) );
NAND2xp5_ASAP7_75t_SL g152 ( .A(n_68), .B(n_141), .Y(n_152) );
AOI21xp5_ASAP7_75t_L g529 ( .A1(n_69), .A2(n_452), .B(n_530), .Y(n_529) );
AND2x2_ASAP7_75t_L g233 ( .A(n_70), .B(n_155), .Y(n_233) );
INVx1_ASAP7_75t_L g125 ( .A(n_71), .Y(n_125) );
INVx1_ASAP7_75t_L g133 ( .A(n_71), .Y(n_133) );
AOI22xp5_ASAP7_75t_L g104 ( .A1(n_72), .A2(n_97), .B1(n_105), .B2(n_106), .Y(n_104) );
CKINVDCx20_ASAP7_75t_R g105 ( .A(n_72), .Y(n_105) );
AND2x2_ASAP7_75t_L g156 ( .A(n_73), .B(n_157), .Y(n_156) );
NAND2xp5_ASAP7_75t_L g523 ( .A(n_74), .B(n_446), .Y(n_523) );
AND2x2_ASAP7_75t_L g461 ( .A(n_76), .B(n_157), .Y(n_461) );
INVx1_ASAP7_75t_L g469 ( .A(n_77), .Y(n_469) );
AOI21xp5_ASAP7_75t_L g451 ( .A1(n_78), .A2(n_452), .B(n_457), .Y(n_451) );
A2O1A1Ixp33_ASAP7_75t_L g550 ( .A1(n_79), .A2(n_452), .B(n_515), .C(n_551), .Y(n_550) );
INVx1_ASAP7_75t_L g435 ( .A(n_80), .Y(n_435) );
NAND2xp5_ASAP7_75t_SL g140 ( .A(n_81), .B(n_141), .Y(n_140) );
AND2x2_ASAP7_75t_L g170 ( .A(n_82), .B(n_157), .Y(n_170) );
AND2x2_ASAP7_75t_SL g480 ( .A(n_83), .B(n_157), .Y(n_480) );
AOI22xp5_ASAP7_75t_L g517 ( .A1(n_84), .A2(n_452), .B1(n_518), .B2(n_519), .Y(n_517) );
AND2x2_ASAP7_75t_L g183 ( .A(n_85), .B(n_118), .Y(n_183) );
NAND2xp5_ASAP7_75t_L g134 ( .A(n_87), .B(n_135), .Y(n_134) );
AND2x2_ASAP7_75t_L g200 ( .A(n_88), .B(n_157), .Y(n_200) );
INVx1_ASAP7_75t_L g484 ( .A(n_89), .Y(n_484) );
AOI22xp5_ASAP7_75t_L g776 ( .A1(n_90), .A2(n_104), .B1(n_777), .B2(n_781), .Y(n_776) );
NAND2xp5_ASAP7_75t_L g231 ( .A(n_91), .B(n_131), .Y(n_231) );
AOI21xp5_ASAP7_75t_L g122 ( .A1(n_92), .A2(n_123), .B(n_129), .Y(n_122) );
NAND2xp5_ASAP7_75t_L g212 ( .A(n_93), .B(n_135), .Y(n_212) );
AND2x2_ASAP7_75t_L g524 ( .A(n_94), .B(n_157), .Y(n_524) );
NAND2xp5_ASAP7_75t_L g175 ( .A(n_95), .B(n_131), .Y(n_175) );
A2O1A1Ixp33_ASAP7_75t_L g499 ( .A1(n_96), .A2(n_500), .B(n_501), .C(n_503), .Y(n_499) );
CKINVDCx20_ASAP7_75t_R g106 ( .A(n_97), .Y(n_106) );
BUFx2_ASAP7_75t_L g788 ( .A(n_98), .Y(n_788) );
BUFx2_ASAP7_75t_SL g801 ( .A(n_98), .Y(n_801) );
AOI21xp5_ASAP7_75t_L g165 ( .A1(n_99), .A2(n_123), .B(n_166), .Y(n_165) );
NAND2xp5_ASAP7_75t_L g485 ( .A(n_100), .B(n_142), .Y(n_485) );
AOI21xp33_ASAP7_75t_SL g101 ( .A1(n_102), .A2(n_810), .B(n_817), .Y(n_101) );
OA21x2_ASAP7_75t_L g102 ( .A1(n_103), .A2(n_785), .B(n_797), .Y(n_102) );
OAI21xp5_ASAP7_75t_L g103 ( .A1(n_104), .A2(n_107), .B(n_776), .Y(n_103) );
INVxp67_ASAP7_75t_L g107 ( .A(n_108), .Y(n_107) );
OAI22x1_ASAP7_75t_L g108 ( .A1(n_109), .A2(n_427), .B1(n_436), .B2(n_774), .Y(n_108) );
OAI22xp5_ASAP7_75t_SL g803 ( .A1(n_109), .A2(n_110), .B1(n_804), .B2(n_807), .Y(n_803) );
INVx2_ASAP7_75t_L g109 ( .A(n_110), .Y(n_109) );
OAI22xp5_ASAP7_75t_L g777 ( .A1(n_110), .A2(n_437), .B1(n_778), .B2(n_779), .Y(n_777) );
OR2x6_ASAP7_75t_L g110 ( .A(n_111), .B(n_325), .Y(n_110) );
NAND3xp33_ASAP7_75t_SL g111 ( .A(n_112), .B(n_237), .C(n_292), .Y(n_111) );
AOI221xp5_ASAP7_75t_L g112 ( .A1(n_113), .A2(n_177), .B1(n_201), .B2(n_205), .C(n_215), .Y(n_112) );
AND2x2_ASAP7_75t_L g113 ( .A(n_114), .B(n_160), .Y(n_113) );
AND2x2_ASAP7_75t_SL g203 ( .A(n_114), .B(n_204), .Y(n_203) );
INVx2_ASAP7_75t_L g236 ( .A(n_114), .Y(n_236) );
AND2x2_ASAP7_75t_L g281 ( .A(n_114), .B(n_218), .Y(n_281) );
AND2x4_ASAP7_75t_L g114 ( .A(n_115), .B(n_145), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_116), .Y(n_115) );
INVx2_ASAP7_75t_L g269 ( .A(n_116), .Y(n_269) );
INVx1_ASAP7_75t_L g279 ( .A(n_116), .Y(n_279) );
AO21x2_ASAP7_75t_L g116 ( .A1(n_117), .A2(n_121), .B(n_143), .Y(n_116) );
NOR2xp33_ASAP7_75t_L g143 ( .A(n_117), .B(n_144), .Y(n_143) );
AO21x2_ASAP7_75t_L g243 ( .A1(n_117), .A2(n_121), .B(n_143), .Y(n_243) );
INVx1_ASAP7_75t_SL g117 ( .A(n_118), .Y(n_117) );
AOI21xp5_ASAP7_75t_L g163 ( .A1(n_118), .A2(n_164), .B(n_165), .Y(n_163) );
NAND2xp5_ASAP7_75t_L g188 ( .A(n_118), .B(n_189), .Y(n_188) );
NOR2xp33_ASAP7_75t_L g476 ( .A(n_118), .B(n_138), .Y(n_476) );
AOI21xp5_ASAP7_75t_L g481 ( .A1(n_118), .A2(n_482), .B(n_486), .Y(n_481) );
AND2x4_ASAP7_75t_L g118 ( .A(n_119), .B(n_120), .Y(n_118) );
AND2x2_ASAP7_75t_SL g155 ( .A(n_119), .B(n_120), .Y(n_155) );
NAND2xp5_ASAP7_75t_L g121 ( .A(n_122), .B(n_140), .Y(n_121) );
AND2x6_ASAP7_75t_L g123 ( .A(n_124), .B(n_126), .Y(n_123) );
BUFx3_ASAP7_75t_L g450 ( .A(n_124), .Y(n_450) );
AND2x6_ASAP7_75t_L g135 ( .A(n_125), .B(n_136), .Y(n_135) );
INVx2_ASAP7_75t_L g456 ( .A(n_125), .Y(n_456) );
AND2x4_ASAP7_75t_L g452 ( .A(n_126), .B(n_453), .Y(n_452) );
AND2x2_ASAP7_75t_L g126 ( .A(n_127), .B(n_128), .Y(n_126) );
AND2x4_ASAP7_75t_L g131 ( .A(n_127), .B(n_132), .Y(n_131) );
INVx2_ASAP7_75t_L g448 ( .A(n_127), .Y(n_448) );
HB1xp67_ASAP7_75t_L g449 ( .A(n_128), .Y(n_449) );
AOI21xp5_ASAP7_75t_L g129 ( .A1(n_130), .A2(n_134), .B(n_138), .Y(n_129) );
INVxp67_ASAP7_75t_L g475 ( .A(n_131), .Y(n_475) );
AND2x4_ASAP7_75t_L g142 ( .A(n_132), .B(n_136), .Y(n_142) );
INVx2_ASAP7_75t_L g132 ( .A(n_133), .Y(n_132) );
INVxp67_ASAP7_75t_L g473 ( .A(n_135), .Y(n_473) );
INVx2_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
AOI21xp5_ASAP7_75t_L g149 ( .A1(n_138), .A2(n_150), .B(n_151), .Y(n_149) );
AOI21xp5_ASAP7_75t_L g166 ( .A1(n_138), .A2(n_167), .B(n_168), .Y(n_166) );
AOI21xp5_ASAP7_75t_L g174 ( .A1(n_138), .A2(n_175), .B(n_176), .Y(n_174) );
AOI21xp5_ASAP7_75t_L g185 ( .A1(n_138), .A2(n_186), .B(n_187), .Y(n_185) );
AOI21xp5_ASAP7_75t_L g195 ( .A1(n_138), .A2(n_196), .B(n_197), .Y(n_195) );
AOI21xp5_ASAP7_75t_L g211 ( .A1(n_138), .A2(n_212), .B(n_213), .Y(n_211) );
AOI21xp5_ASAP7_75t_L g229 ( .A1(n_138), .A2(n_230), .B(n_231), .Y(n_229) );
O2A1O1Ixp33_ASAP7_75t_SL g457 ( .A1(n_138), .A2(n_458), .B(n_459), .C(n_460), .Y(n_457) );
O2A1O1Ixp33_ASAP7_75t_L g483 ( .A1(n_138), .A2(n_459), .B(n_484), .C(n_485), .Y(n_483) );
O2A1O1Ixp33_ASAP7_75t_SL g492 ( .A1(n_138), .A2(n_459), .B(n_493), .C(n_494), .Y(n_492) );
INVx1_ASAP7_75t_L g518 ( .A(n_138), .Y(n_518) );
O2A1O1Ixp33_ASAP7_75t_L g530 ( .A1(n_138), .A2(n_459), .B(n_531), .C(n_532), .Y(n_530) );
AOI21xp5_ASAP7_75t_L g551 ( .A1(n_138), .A2(n_552), .B(n_553), .Y(n_551) );
INVx5_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
AND2x4_ASAP7_75t_L g141 ( .A(n_139), .B(n_142), .Y(n_141) );
HB1xp67_ASAP7_75t_L g503 ( .A(n_139), .Y(n_503) );
INVx1_ASAP7_75t_L g470 ( .A(n_142), .Y(n_470) );
OR2x2_ASAP7_75t_L g258 ( .A(n_145), .B(n_161), .Y(n_258) );
NAND2x1p5_ASAP7_75t_L g289 ( .A(n_145), .B(n_204), .Y(n_289) );
NAND2xp5_ASAP7_75t_L g302 ( .A(n_145), .B(n_169), .Y(n_302) );
INVx2_ASAP7_75t_L g311 ( .A(n_145), .Y(n_311) );
AND2x2_ASAP7_75t_L g332 ( .A(n_145), .B(n_333), .Y(n_332) );
AND2x2_ASAP7_75t_L g416 ( .A(n_145), .B(n_235), .Y(n_416) );
INVx4_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
AND2x2_ASAP7_75t_L g244 ( .A(n_146), .B(n_169), .Y(n_244) );
AND2x2_ASAP7_75t_L g377 ( .A(n_146), .B(n_204), .Y(n_377) );
HB1xp67_ASAP7_75t_L g403 ( .A(n_146), .Y(n_403) );
AO21x2_ASAP7_75t_L g146 ( .A1(n_147), .A2(n_153), .B(n_156), .Y(n_146) );
NAND2xp5_ASAP7_75t_L g147 ( .A(n_148), .B(n_152), .Y(n_147) );
AO21x2_ASAP7_75t_L g443 ( .A1(n_153), .A2(n_444), .B(n_461), .Y(n_443) );
CKINVDCx5p33_ASAP7_75t_R g153 ( .A(n_154), .Y(n_153) );
AOI21xp5_ASAP7_75t_L g171 ( .A1(n_154), .A2(n_172), .B(n_173), .Y(n_171) );
OA21x2_ASAP7_75t_L g209 ( .A1(n_154), .A2(n_210), .B(n_214), .Y(n_209) );
OA21x2_ASAP7_75t_L g221 ( .A1(n_154), .A2(n_210), .B(n_214), .Y(n_221) );
BUFx6f_ASAP7_75t_L g154 ( .A(n_155), .Y(n_154) );
INVx3_ASAP7_75t_L g199 ( .A(n_157), .Y(n_199) );
OAI22xp5_ASAP7_75t_L g498 ( .A1(n_157), .A2(n_199), .B1(n_499), .B2(n_504), .Y(n_498) );
INVx4_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
NAND2xp5_ASAP7_75t_L g506 ( .A(n_158), .B(n_507), .Y(n_506) );
INVx3_ASAP7_75t_L g158 ( .A(n_159), .Y(n_158) );
BUFx4f_ASAP7_75t_L g162 ( .A(n_159), .Y(n_162) );
AND2x4_ASAP7_75t_L g331 ( .A(n_160), .B(n_332), .Y(n_331) );
AOI321xp33_ASAP7_75t_L g345 ( .A1(n_160), .A2(n_274), .A3(n_275), .B1(n_307), .B2(n_346), .C(n_349), .Y(n_345) );
AND2x2_ASAP7_75t_L g160 ( .A(n_161), .B(n_169), .Y(n_160) );
BUFx3_ASAP7_75t_L g202 ( .A(n_161), .Y(n_202) );
INVx2_ASAP7_75t_L g235 ( .A(n_161), .Y(n_235) );
NAND2xp5_ASAP7_75t_L g242 ( .A(n_161), .B(n_243), .Y(n_242) );
AND2x2_ASAP7_75t_L g268 ( .A(n_161), .B(n_269), .Y(n_268) );
INVx1_ASAP7_75t_L g301 ( .A(n_161), .Y(n_301) );
OA21x2_ASAP7_75t_L g490 ( .A1(n_162), .A2(n_491), .B(n_495), .Y(n_490) );
INVx2_ASAP7_75t_SL g515 ( .A(n_162), .Y(n_515) );
INVx5_ASAP7_75t_L g204 ( .A(n_169), .Y(n_204) );
NOR2x1_ASAP7_75t_SL g253 ( .A(n_169), .B(n_243), .Y(n_253) );
BUFx2_ASAP7_75t_L g348 ( .A(n_169), .Y(n_348) );
OR2x6_ASAP7_75t_L g169 ( .A(n_170), .B(n_171), .Y(n_169) );
INVxp67_ASAP7_75t_L g177 ( .A(n_178), .Y(n_177) );
NAND2xp5_ASAP7_75t_L g178 ( .A(n_179), .B(n_190), .Y(n_178) );
NOR2xp33_ASAP7_75t_SL g246 ( .A(n_179), .B(n_247), .Y(n_246) );
NOR4xp25_ASAP7_75t_L g349 ( .A(n_179), .B(n_343), .C(n_347), .D(n_350), .Y(n_349) );
INVx1_ASAP7_75t_L g387 ( .A(n_179), .Y(n_387) );
AND2x2_ASAP7_75t_L g421 ( .A(n_179), .B(n_361), .Y(n_421) );
BUFx2_ASAP7_75t_L g179 ( .A(n_180), .Y(n_179) );
INVx2_ASAP7_75t_L g222 ( .A(n_180), .Y(n_222) );
INVx2_ASAP7_75t_L g180 ( .A(n_181), .Y(n_180) );
INVx2_ASAP7_75t_L g276 ( .A(n_181), .Y(n_276) );
OAI21x1_ASAP7_75t_SL g181 ( .A1(n_182), .A2(n_184), .B(n_188), .Y(n_181) );
INVx1_ASAP7_75t_L g189 ( .A(n_183), .Y(n_189) );
AOI33xp33_ASAP7_75t_L g417 ( .A1(n_190), .A2(n_219), .A3(n_250), .B1(n_266), .B2(n_372), .B3(n_418), .Y(n_417) );
INVx1_ASAP7_75t_SL g190 ( .A(n_191), .Y(n_190) );
AND2x2_ASAP7_75t_L g207 ( .A(n_191), .B(n_208), .Y(n_207) );
AND2x4_ASAP7_75t_L g217 ( .A(n_191), .B(n_218), .Y(n_217) );
BUFx3_ASAP7_75t_L g191 ( .A(n_192), .Y(n_191) );
INVx2_ASAP7_75t_L g224 ( .A(n_192), .Y(n_224) );
INVxp67_ASAP7_75t_L g305 ( .A(n_192), .Y(n_305) );
AND2x2_ASAP7_75t_L g361 ( .A(n_192), .B(n_226), .Y(n_361) );
AO21x2_ASAP7_75t_L g192 ( .A1(n_193), .A2(n_199), .B(n_200), .Y(n_192) );
AO21x2_ASAP7_75t_L g265 ( .A1(n_193), .A2(n_199), .B(n_200), .Y(n_265) );
NAND2xp5_ASAP7_75t_L g193 ( .A(n_194), .B(n_198), .Y(n_193) );
AO21x2_ASAP7_75t_L g226 ( .A1(n_199), .A2(n_227), .B(n_233), .Y(n_226) );
AO21x2_ASAP7_75t_L g262 ( .A1(n_199), .A2(n_227), .B(n_233), .Y(n_262) );
AO21x2_ASAP7_75t_L g526 ( .A1(n_199), .A2(n_527), .B(n_533), .Y(n_526) );
AO21x2_ASAP7_75t_L g564 ( .A1(n_199), .A2(n_527), .B(n_533), .Y(n_564) );
AOI21xp5_ASAP7_75t_L g382 ( .A1(n_201), .A2(n_383), .B(n_384), .Y(n_382) );
AND2x2_ASAP7_75t_L g201 ( .A(n_202), .B(n_203), .Y(n_201) );
AND2x2_ASAP7_75t_L g370 ( .A(n_202), .B(n_244), .Y(n_370) );
AND3x2_ASAP7_75t_L g372 ( .A(n_202), .B(n_256), .C(n_311), .Y(n_372) );
INVx3_ASAP7_75t_SL g324 ( .A(n_203), .Y(n_324) );
INVx4_ASAP7_75t_L g218 ( .A(n_204), .Y(n_218) );
AND2x2_ASAP7_75t_L g256 ( .A(n_204), .B(n_243), .Y(n_256) );
INVxp67_ASAP7_75t_L g205 ( .A(n_206), .Y(n_205) );
INVx1_ASAP7_75t_L g206 ( .A(n_207), .Y(n_206) );
BUFx2_ASAP7_75t_L g250 ( .A(n_208), .Y(n_250) );
AND2x4_ASAP7_75t_L g275 ( .A(n_208), .B(n_276), .Y(n_275) );
AND2x2_ASAP7_75t_L g338 ( .A(n_208), .B(n_226), .Y(n_338) );
INVx2_ASAP7_75t_L g208 ( .A(n_209), .Y(n_208) );
INVx2_ASAP7_75t_L g308 ( .A(n_209), .Y(n_308) );
HB1xp67_ASAP7_75t_L g330 ( .A(n_209), .Y(n_330) );
O2A1O1Ixp33_ASAP7_75t_R g215 ( .A1(n_216), .A2(n_219), .B(n_223), .C(n_234), .Y(n_215) );
CKINVDCx16_ASAP7_75t_R g216 ( .A(n_217), .Y(n_216) );
AND2x2_ASAP7_75t_L g267 ( .A(n_218), .B(n_268), .Y(n_267) );
NAND2xp5_ASAP7_75t_L g278 ( .A(n_218), .B(n_279), .Y(n_278) );
NAND2xp5_ASAP7_75t_L g396 ( .A(n_218), .B(n_235), .Y(n_396) );
INVx1_ASAP7_75t_SL g219 ( .A(n_220), .Y(n_219) );
AND2x2_ASAP7_75t_L g378 ( .A(n_220), .B(n_368), .Y(n_378) );
AND2x2_ASAP7_75t_SL g220 ( .A(n_221), .B(n_222), .Y(n_220) );
AND2x2_ASAP7_75t_L g225 ( .A(n_221), .B(n_226), .Y(n_225) );
AND2x2_ASAP7_75t_L g247 ( .A(n_221), .B(n_248), .Y(n_247) );
AND2x2_ASAP7_75t_L g263 ( .A(n_221), .B(n_264), .Y(n_263) );
AND2x4_ASAP7_75t_L g296 ( .A(n_221), .B(n_276), .Y(n_296) );
AND2x4_ASAP7_75t_L g261 ( .A(n_222), .B(n_262), .Y(n_261) );
OR2x2_ASAP7_75t_L g285 ( .A(n_222), .B(n_286), .Y(n_285) );
AND2x2_ASAP7_75t_L g323 ( .A(n_222), .B(n_248), .Y(n_323) );
NAND2xp5_ASAP7_75t_L g223 ( .A(n_224), .B(n_225), .Y(n_223) );
AND2x2_ASAP7_75t_L g251 ( .A(n_224), .B(n_248), .Y(n_251) );
AND2x2_ASAP7_75t_L g266 ( .A(n_224), .B(n_226), .Y(n_266) );
BUFx2_ASAP7_75t_L g322 ( .A(n_224), .Y(n_322) );
AND2x2_ASAP7_75t_L g336 ( .A(n_224), .B(n_247), .Y(n_336) );
INVx2_ASAP7_75t_L g248 ( .A(n_226), .Y(n_248) );
NAND2xp5_ASAP7_75t_SL g227 ( .A(n_228), .B(n_232), .Y(n_227) );
OAI22xp33_ASAP7_75t_L g284 ( .A1(n_234), .A2(n_285), .B1(n_287), .B2(n_291), .Y(n_284) );
INVx2_ASAP7_75t_SL g315 ( .A(n_234), .Y(n_315) );
OR2x2_ASAP7_75t_L g234 ( .A(n_235), .B(n_236), .Y(n_234) );
AND2x2_ASAP7_75t_L g290 ( .A(n_235), .B(n_243), .Y(n_290) );
INVx1_ASAP7_75t_L g397 ( .A(n_236), .Y(n_397) );
NOR3xp33_ASAP7_75t_L g237 ( .A(n_238), .B(n_270), .C(n_284), .Y(n_237) );
OAI221xp5_ASAP7_75t_SL g238 ( .A1(n_239), .A2(n_245), .B1(n_249), .B2(n_252), .C(n_254), .Y(n_238) );
INVx1_ASAP7_75t_SL g239 ( .A(n_240), .Y(n_239) );
AND2x2_ASAP7_75t_L g240 ( .A(n_241), .B(n_244), .Y(n_240) );
INVxp67_ASAP7_75t_SL g241 ( .A(n_242), .Y(n_241) );
INVx1_ASAP7_75t_L g298 ( .A(n_242), .Y(n_298) );
INVxp67_ASAP7_75t_SL g426 ( .A(n_242), .Y(n_426) );
INVx1_ASAP7_75t_L g389 ( .A(n_244), .Y(n_389) );
AND2x2_ASAP7_75t_SL g399 ( .A(n_244), .B(n_268), .Y(n_399) );
INVxp67_ASAP7_75t_L g245 ( .A(n_246), .Y(n_245) );
NAND2xp5_ASAP7_75t_L g304 ( .A(n_248), .B(n_276), .Y(n_304) );
NAND2xp5_ASAP7_75t_L g249 ( .A(n_250), .B(n_251), .Y(n_249) );
OR2x2_ASAP7_75t_L g282 ( .A(n_250), .B(n_283), .Y(n_282) );
INVx1_ASAP7_75t_L g360 ( .A(n_250), .Y(n_360) );
AND2x2_ASAP7_75t_L g295 ( .A(n_251), .B(n_296), .Y(n_295) );
INVx1_ASAP7_75t_L g252 ( .A(n_253), .Y(n_252) );
AND2x2_ASAP7_75t_L g341 ( .A(n_253), .B(n_301), .Y(n_341) );
AND2x2_ASAP7_75t_L g418 ( .A(n_253), .B(n_416), .Y(n_418) );
AOI22xp5_ASAP7_75t_L g254 ( .A1(n_255), .A2(n_259), .B1(n_266), .B2(n_267), .Y(n_254) );
AND2x4_ASAP7_75t_L g255 ( .A(n_256), .B(n_257), .Y(n_255) );
INVx2_ASAP7_75t_L g257 ( .A(n_258), .Y(n_257) );
OR2x2_ASAP7_75t_L g277 ( .A(n_258), .B(n_278), .Y(n_277) );
INVx1_ASAP7_75t_SL g259 ( .A(n_260), .Y(n_259) );
NAND2xp5_ASAP7_75t_L g260 ( .A(n_261), .B(n_263), .Y(n_260) );
INVx2_ASAP7_75t_L g283 ( .A(n_261), .Y(n_283) );
AND2x4_ASAP7_75t_L g307 ( .A(n_261), .B(n_308), .Y(n_307) );
OAI21xp33_ASAP7_75t_SL g337 ( .A1(n_261), .A2(n_338), .B(n_339), .Y(n_337) );
AND2x2_ASAP7_75t_L g364 ( .A(n_261), .B(n_322), .Y(n_364) );
INVx2_ASAP7_75t_L g286 ( .A(n_262), .Y(n_286) );
HB1xp67_ASAP7_75t_L g319 ( .A(n_262), .Y(n_319) );
INVx1_ASAP7_75t_SL g343 ( .A(n_263), .Y(n_343) );
INVx1_ASAP7_75t_L g264 ( .A(n_265), .Y(n_264) );
BUFx2_ASAP7_75t_L g274 ( .A(n_265), .Y(n_274) );
AND2x4_ASAP7_75t_SL g368 ( .A(n_265), .B(n_286), .Y(n_368) );
AND2x2_ASAP7_75t_L g365 ( .A(n_268), .B(n_311), .Y(n_365) );
AND2x2_ASAP7_75t_L g391 ( .A(n_268), .B(n_377), .Y(n_391) );
HB1xp67_ASAP7_75t_L g313 ( .A(n_269), .Y(n_313) );
INVx1_ASAP7_75t_L g333 ( .A(n_269), .Y(n_333) );
OAI22xp33_ASAP7_75t_L g270 ( .A1(n_271), .A2(n_277), .B1(n_280), .B2(n_282), .Y(n_270) );
INVx1_ASAP7_75t_L g271 ( .A(n_272), .Y(n_271) );
AND2x2_ASAP7_75t_L g272 ( .A(n_273), .B(n_275), .Y(n_272) );
INVx2_ASAP7_75t_L g273 ( .A(n_274), .Y(n_273) );
NAND2xp5_ASAP7_75t_SL g291 ( .A(n_275), .B(n_286), .Y(n_291) );
NAND2xp5_ASAP7_75t_L g367 ( .A(n_275), .B(n_368), .Y(n_367) );
INVx1_ASAP7_75t_L g414 ( .A(n_275), .Y(n_414) );
INVx2_ASAP7_75t_SL g339 ( .A(n_277), .Y(n_339) );
AND2x2_ASAP7_75t_L g351 ( .A(n_279), .B(n_311), .Y(n_351) );
INVx2_ASAP7_75t_L g357 ( .A(n_279), .Y(n_357) );
INVxp33_ASAP7_75t_L g280 ( .A(n_281), .Y(n_280) );
INVx2_ASAP7_75t_L g316 ( .A(n_282), .Y(n_316) );
NOR2xp33_ASAP7_75t_L g342 ( .A(n_285), .B(n_343), .Y(n_342) );
INVx1_ASAP7_75t_L g407 ( .A(n_285), .Y(n_407) );
INVx1_ASAP7_75t_L g335 ( .A(n_287), .Y(n_335) );
NAND2xp5_ASAP7_75t_L g287 ( .A(n_288), .B(n_290), .Y(n_287) );
NAND2xp5_ASAP7_75t_L g354 ( .A(n_288), .B(n_355), .Y(n_354) );
INVx2_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
AND2x2_ASAP7_75t_L g346 ( .A(n_290), .B(n_347), .Y(n_346) );
AOI22xp5_ASAP7_75t_L g419 ( .A1(n_290), .A2(n_420), .B1(n_421), .B2(n_422), .Y(n_419) );
NOR3xp33_ASAP7_75t_L g292 ( .A(n_293), .B(n_314), .C(n_317), .Y(n_292) );
OAI221xp5_ASAP7_75t_L g293 ( .A1(n_294), .A2(n_297), .B1(n_299), .B2(n_303), .C(n_306), .Y(n_293) );
INVx1_ASAP7_75t_SL g294 ( .A(n_295), .Y(n_294) );
INVx1_ASAP7_75t_SL g412 ( .A(n_297), .Y(n_412) );
INVx1_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
AND2x2_ASAP7_75t_L g381 ( .A(n_298), .B(n_347), .Y(n_381) );
OR2x2_ASAP7_75t_L g299 ( .A(n_300), .B(n_302), .Y(n_299) );
INVx1_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
AND2x2_ASAP7_75t_L g312 ( .A(n_301), .B(n_313), .Y(n_312) );
INVx1_ASAP7_75t_L g383 ( .A(n_303), .Y(n_383) );
OR2x2_ASAP7_75t_L g303 ( .A(n_304), .B(n_305), .Y(n_303) );
INVx1_ASAP7_75t_L g380 ( .A(n_304), .Y(n_380) );
INVx1_ASAP7_75t_L g386 ( .A(n_305), .Y(n_386) );
OR2x2_ASAP7_75t_L g409 ( .A(n_305), .B(n_410), .Y(n_409) );
NAND2xp5_ASAP7_75t_L g306 ( .A(n_307), .B(n_309), .Y(n_306) );
INVx1_ASAP7_75t_SL g318 ( .A(n_308), .Y(n_318) );
AND2x2_ASAP7_75t_L g388 ( .A(n_308), .B(n_368), .Y(n_388) );
AND2x2_ASAP7_75t_SL g420 ( .A(n_308), .B(n_321), .Y(n_420) );
INVx1_ASAP7_75t_SL g309 ( .A(n_310), .Y(n_309) );
NAND2xp5_ASAP7_75t_L g310 ( .A(n_311), .B(n_312), .Y(n_310) );
INVx1_ASAP7_75t_L g425 ( .A(n_311), .Y(n_425) );
INVx1_ASAP7_75t_L g375 ( .A(n_313), .Y(n_375) );
AND2x2_ASAP7_75t_L g314 ( .A(n_315), .B(n_316), .Y(n_314) );
O2A1O1Ixp33_ASAP7_75t_L g317 ( .A1(n_318), .A2(n_319), .B(n_320), .C(n_324), .Y(n_317) );
NAND2xp5_ASAP7_75t_L g392 ( .A(n_318), .B(n_368), .Y(n_392) );
INVx1_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
NAND2xp5_ASAP7_75t_L g371 ( .A(n_321), .B(n_372), .Y(n_371) );
AND2x2_ASAP7_75t_L g321 ( .A(n_322), .B(n_323), .Y(n_321) );
AND2x2_ASAP7_75t_L g329 ( .A(n_323), .B(n_330), .Y(n_329) );
INVx1_ASAP7_75t_L g410 ( .A(n_323), .Y(n_410) );
NAND4xp75_ASAP7_75t_L g325 ( .A(n_326), .B(n_382), .C(n_398), .D(n_419), .Y(n_325) );
NOR3x1_ASAP7_75t_L g326 ( .A(n_327), .B(n_344), .C(n_366), .Y(n_326) );
NAND4xp75_ASAP7_75t_L g327 ( .A(n_328), .B(n_334), .C(n_337), .D(n_340), .Y(n_327) );
NAND2xp5_ASAP7_75t_SL g328 ( .A(n_329), .B(n_331), .Y(n_328) );
AND2x2_ASAP7_75t_L g379 ( .A(n_330), .B(n_380), .Y(n_379) );
INVx1_ASAP7_75t_SL g404 ( .A(n_331), .Y(n_404) );
NAND2xp5_ASAP7_75t_SL g334 ( .A(n_335), .B(n_336), .Y(n_334) );
INVx1_ASAP7_75t_SL g393 ( .A(n_336), .Y(n_393) );
NAND2xp5_ASAP7_75t_L g340 ( .A(n_341), .B(n_342), .Y(n_340) );
NAND2xp5_ASAP7_75t_L g344 ( .A(n_345), .B(n_352), .Y(n_344) );
INVx2_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
NAND2xp5_ASAP7_75t_L g411 ( .A(n_348), .B(n_412), .Y(n_411) );
INVx1_ASAP7_75t_SL g350 ( .A(n_351), .Y(n_350) );
AOI21xp5_ASAP7_75t_L g352 ( .A1(n_353), .A2(n_358), .B(n_362), .Y(n_352) );
INVx1_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
INVx1_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
OAI322xp33_ASAP7_75t_L g384 ( .A1(n_356), .A2(n_385), .A3(n_389), .B1(n_390), .B2(n_392), .C1(n_393), .C2(n_394), .Y(n_384) );
INVx2_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
NAND2xp5_ASAP7_75t_L g402 ( .A(n_357), .B(n_403), .Y(n_402) );
INVx1_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
NAND2xp5_ASAP7_75t_L g359 ( .A(n_360), .B(n_361), .Y(n_359) );
NAND2xp5_ASAP7_75t_L g406 ( .A(n_360), .B(n_407), .Y(n_406) );
NAND2xp5_ASAP7_75t_L g413 ( .A(n_361), .B(n_414), .Y(n_413) );
INVx1_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
NAND2xp5_ASAP7_75t_L g363 ( .A(n_364), .B(n_365), .Y(n_363) );
OAI211xp5_ASAP7_75t_L g366 ( .A1(n_367), .A2(n_369), .B(n_371), .C(n_373), .Y(n_366) );
INVx1_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
AOI22xp5_ASAP7_75t_L g373 ( .A1(n_374), .A2(n_378), .B1(n_379), .B2(n_381), .Y(n_373) );
NOR2xp33_ASAP7_75t_SL g374 ( .A(n_375), .B(n_376), .Y(n_374) );
INVx2_ASAP7_75t_SL g376 ( .A(n_377), .Y(n_376) );
AOI21xp5_ASAP7_75t_L g385 ( .A1(n_386), .A2(n_387), .B(n_388), .Y(n_385) );
INVxp67_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
NOR2xp33_ASAP7_75t_L g423 ( .A(n_391), .B(n_424), .Y(n_423) );
NAND2xp5_ASAP7_75t_SL g394 ( .A(n_395), .B(n_397), .Y(n_394) );
INVx1_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
OR2x2_ASAP7_75t_L g401 ( .A(n_396), .B(n_402), .Y(n_401) );
O2A1O1Ixp5_ASAP7_75t_L g398 ( .A1(n_399), .A2(n_400), .B(n_405), .C(n_408), .Y(n_398) );
NAND2xp5_ASAP7_75t_SL g400 ( .A(n_401), .B(n_404), .Y(n_400) );
INVx1_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
OAI221xp5_ASAP7_75t_SL g408 ( .A1(n_409), .A2(n_411), .B1(n_413), .B2(n_415), .C(n_417), .Y(n_408) );
INVxp67_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
INVx1_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
AND2x2_ASAP7_75t_L g424 ( .A(n_425), .B(n_426), .Y(n_424) );
INVx4_ASAP7_75t_SL g427 ( .A(n_428), .Y(n_427) );
CKINVDCx6p67_ASAP7_75t_R g778 ( .A(n_428), .Y(n_778) );
INVx3_ASAP7_75t_SL g428 ( .A(n_429), .Y(n_428) );
CKINVDCx5p33_ASAP7_75t_R g429 ( .A(n_430), .Y(n_429) );
AND2x6_ASAP7_75t_SL g430 ( .A(n_431), .B(n_432), .Y(n_430) );
OR2x6_ASAP7_75t_SL g774 ( .A(n_431), .B(n_775), .Y(n_774) );
OR2x2_ASAP7_75t_L g784 ( .A(n_431), .B(n_432), .Y(n_784) );
NAND2xp5_ASAP7_75t_L g795 ( .A(n_431), .B(n_775), .Y(n_795) );
CKINVDCx5p33_ASAP7_75t_R g775 ( .A(n_432), .Y(n_775) );
NAND2xp5_ASAP7_75t_L g433 ( .A(n_434), .B(n_435), .Y(n_433) );
INVx1_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
OR3x2_ASAP7_75t_L g437 ( .A(n_438), .B(n_639), .C(n_710), .Y(n_437) );
NAND3x1_ASAP7_75t_SL g438 ( .A(n_439), .B(n_566), .C(n_588), .Y(n_438) );
AND2x2_ASAP7_75t_L g439 ( .A(n_440), .B(n_556), .Y(n_439) );
AOI22xp33_ASAP7_75t_SL g440 ( .A1(n_441), .A2(n_487), .B1(n_534), .B2(n_538), .Y(n_440) );
AOI22xp33_ASAP7_75t_L g741 ( .A1(n_441), .A2(n_742), .B1(n_743), .B2(n_745), .Y(n_741) );
AND2x2_ASAP7_75t_L g441 ( .A(n_442), .B(n_462), .Y(n_441) );
AND2x2_ASAP7_75t_L g557 ( .A(n_442), .B(n_558), .Y(n_557) );
NAND2xp5_ASAP7_75t_SL g623 ( .A(n_442), .B(n_604), .Y(n_623) );
INVx1_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
INVx2_ASAP7_75t_L g541 ( .A(n_443), .Y(n_541) );
AND2x2_ASAP7_75t_L g591 ( .A(n_443), .B(n_464), .Y(n_591) );
INVx1_ASAP7_75t_L g630 ( .A(n_443), .Y(n_630) );
OR2x2_ASAP7_75t_L g667 ( .A(n_443), .B(n_479), .Y(n_667) );
HB1xp67_ASAP7_75t_L g679 ( .A(n_443), .Y(n_679) );
HB1xp67_ASAP7_75t_L g703 ( .A(n_443), .Y(n_703) );
AND2x2_ASAP7_75t_L g760 ( .A(n_443), .B(n_587), .Y(n_760) );
NAND2xp5_ASAP7_75t_L g444 ( .A(n_445), .B(n_451), .Y(n_444) );
INVx1_ASAP7_75t_L g511 ( .A(n_446), .Y(n_511) );
AND2x4_ASAP7_75t_L g446 ( .A(n_447), .B(n_450), .Y(n_446) );
INVx1_ASAP7_75t_L g547 ( .A(n_447), .Y(n_547) );
AND2x2_ASAP7_75t_L g447 ( .A(n_448), .B(n_449), .Y(n_447) );
OR2x6_ASAP7_75t_L g459 ( .A(n_448), .B(n_456), .Y(n_459) );
INVxp33_ASAP7_75t_L g521 ( .A(n_448), .Y(n_521) );
INVx1_ASAP7_75t_L g548 ( .A(n_450), .Y(n_548) );
INVxp67_ASAP7_75t_L g509 ( .A(n_452), .Y(n_509) );
NOR2x1p5_ASAP7_75t_L g453 ( .A(n_454), .B(n_455), .Y(n_453) );
INVx1_ASAP7_75t_L g522 ( .A(n_455), .Y(n_522) );
INVx3_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
OAI22xp5_ASAP7_75t_L g467 ( .A1(n_459), .A2(n_468), .B1(n_469), .B2(n_470), .Y(n_467) );
INVxp67_ASAP7_75t_L g500 ( .A(n_459), .Y(n_500) );
INVx2_ASAP7_75t_L g554 ( .A(n_459), .Y(n_554) );
NOR2x1_ASAP7_75t_L g462 ( .A(n_463), .B(n_477), .Y(n_462) );
INVx1_ASAP7_75t_L g635 ( .A(n_463), .Y(n_635) );
AND2x2_ASAP7_75t_L g661 ( .A(n_463), .B(n_479), .Y(n_661) );
NAND2x1_ASAP7_75t_L g677 ( .A(n_463), .B(n_678), .Y(n_677) );
INVx2_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
AND2x2_ASAP7_75t_L g558 ( .A(n_464), .B(n_544), .Y(n_558) );
INVx3_ASAP7_75t_L g587 ( .A(n_464), .Y(n_587) );
NOR2x1_ASAP7_75t_SL g706 ( .A(n_464), .B(n_479), .Y(n_706) );
AND2x4_ASAP7_75t_L g464 ( .A(n_465), .B(n_466), .Y(n_464) );
OAI21xp5_ASAP7_75t_L g466 ( .A1(n_467), .A2(n_471), .B(n_476), .Y(n_466) );
NOR2xp33_ASAP7_75t_L g501 ( .A(n_470), .B(n_502), .Y(n_501) );
OAI22xp5_ASAP7_75t_L g471 ( .A1(n_472), .A2(n_473), .B1(n_474), .B2(n_475), .Y(n_471) );
NOR2x1_ASAP7_75t_L g614 ( .A(n_477), .B(n_615), .Y(n_614) );
INVx1_ASAP7_75t_L g477 ( .A(n_478), .Y(n_477) );
AND2x2_ASAP7_75t_L g585 ( .A(n_478), .B(n_586), .Y(n_585) );
INVx2_ASAP7_75t_L g478 ( .A(n_479), .Y(n_478) );
INVx4_ASAP7_75t_L g555 ( .A(n_479), .Y(n_555) );
BUFx6f_ASAP7_75t_L g600 ( .A(n_479), .Y(n_600) );
AND2x2_ASAP7_75t_L g672 ( .A(n_479), .B(n_544), .Y(n_672) );
AND2x4_ASAP7_75t_L g689 ( .A(n_479), .B(n_633), .Y(n_689) );
NAND2xp5_ASAP7_75t_SL g736 ( .A(n_479), .B(n_631), .Y(n_736) );
NAND2xp5_ASAP7_75t_L g765 ( .A(n_479), .B(n_540), .Y(n_765) );
OR2x6_ASAP7_75t_L g479 ( .A(n_480), .B(n_481), .Y(n_479) );
AOI22xp5_ASAP7_75t_L g694 ( .A1(n_487), .A2(n_582), .B1(n_653), .B2(n_695), .Y(n_694) );
AND2x2_ASAP7_75t_L g487 ( .A(n_488), .B(n_512), .Y(n_487) );
INVx2_ASAP7_75t_L g655 ( .A(n_488), .Y(n_655) );
AND2x2_ASAP7_75t_L g488 ( .A(n_489), .B(n_496), .Y(n_488) );
BUFx3_ASAP7_75t_L g645 ( .A(n_489), .Y(n_645) );
INVx1_ASAP7_75t_L g489 ( .A(n_490), .Y(n_489) );
NAND2xp5_ASAP7_75t_L g537 ( .A(n_490), .B(n_514), .Y(n_537) );
INVx2_ASAP7_75t_L g561 ( .A(n_490), .Y(n_561) );
INVx1_ASAP7_75t_L g573 ( .A(n_490), .Y(n_573) );
AND2x4_ASAP7_75t_L g580 ( .A(n_490), .B(n_581), .Y(n_580) );
AND2x2_ASAP7_75t_L g597 ( .A(n_490), .B(n_497), .Y(n_597) );
HB1xp67_ASAP7_75t_L g611 ( .A(n_490), .Y(n_611) );
INVxp67_ASAP7_75t_L g619 ( .A(n_490), .Y(n_619) );
AND2x2_ASAP7_75t_L g648 ( .A(n_496), .B(n_564), .Y(n_648) );
AND2x2_ASAP7_75t_L g664 ( .A(n_496), .B(n_565), .Y(n_664) );
NOR2xp67_ASAP7_75t_L g751 ( .A(n_496), .B(n_564), .Y(n_751) );
INVx2_ASAP7_75t_L g496 ( .A(n_497), .Y(n_496) );
AND2x4_ASAP7_75t_L g560 ( .A(n_497), .B(n_561), .Y(n_560) );
INVx1_ASAP7_75t_L g571 ( .A(n_497), .Y(n_571) );
INVx1_ASAP7_75t_L g584 ( .A(n_497), .Y(n_584) );
NAND2xp5_ASAP7_75t_L g621 ( .A(n_497), .B(n_526), .Y(n_621) );
OR2x2_ASAP7_75t_L g497 ( .A(n_498), .B(n_505), .Y(n_497) );
OAI22xp5_ASAP7_75t_L g505 ( .A1(n_506), .A2(n_509), .B1(n_510), .B2(n_511), .Y(n_505) );
INVx1_ASAP7_75t_L g507 ( .A(n_508), .Y(n_507) );
INVx1_ASAP7_75t_L g744 ( .A(n_512), .Y(n_744) );
AND2x4_ASAP7_75t_L g512 ( .A(n_513), .B(n_525), .Y(n_512) );
AND2x2_ASAP7_75t_L g618 ( .A(n_513), .B(n_619), .Y(n_618) );
INVx1_ASAP7_75t_L g647 ( .A(n_513), .Y(n_647) );
AND2x2_ASAP7_75t_L g749 ( .A(n_513), .B(n_564), .Y(n_749) );
INVx2_ASAP7_75t_L g513 ( .A(n_514), .Y(n_513) );
NAND2xp5_ASAP7_75t_L g609 ( .A(n_514), .B(n_526), .Y(n_609) );
AO21x2_ASAP7_75t_L g514 ( .A1(n_515), .A2(n_516), .B(n_524), .Y(n_514) );
AO21x2_ASAP7_75t_L g565 ( .A1(n_515), .A2(n_516), .B(n_524), .Y(n_565) );
NAND2xp5_ASAP7_75t_SL g516 ( .A(n_517), .B(n_523), .Y(n_516) );
INVx1_ASAP7_75t_L g519 ( .A(n_520), .Y(n_519) );
INVx3_ASAP7_75t_L g535 ( .A(n_525), .Y(n_535) );
NAND2x1p5_ASAP7_75t_L g724 ( .A(n_525), .B(n_645), .Y(n_724) );
INVx3_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
HB1xp67_ASAP7_75t_L g638 ( .A(n_526), .Y(n_638) );
AND2x2_ASAP7_75t_L g665 ( .A(n_526), .B(n_611), .Y(n_665) );
NAND2xp5_ASAP7_75t_L g527 ( .A(n_528), .B(n_529), .Y(n_527) );
AND2x2_ASAP7_75t_L g534 ( .A(n_535), .B(n_536), .Y(n_534) );
AND2x2_ASAP7_75t_L g579 ( .A(n_535), .B(n_580), .Y(n_579) );
INVx1_ASAP7_75t_L g595 ( .A(n_535), .Y(n_595) );
AND2x2_ASAP7_75t_L g683 ( .A(n_535), .B(n_560), .Y(n_683) );
NAND2xp5_ASAP7_75t_L g708 ( .A(n_535), .B(n_703), .Y(n_708) );
AND2x2_ASAP7_75t_L g718 ( .A(n_535), .B(n_597), .Y(n_718) );
OR2x2_ASAP7_75t_L g755 ( .A(n_535), .B(n_655), .Y(n_755) );
NAND2xp5_ASAP7_75t_L g594 ( .A(n_536), .B(n_595), .Y(n_594) );
AND2x2_ASAP7_75t_L g715 ( .A(n_536), .B(n_571), .Y(n_715) );
AND2x2_ASAP7_75t_L g731 ( .A(n_536), .B(n_732), .Y(n_731) );
INVx2_ASAP7_75t_L g536 ( .A(n_537), .Y(n_536) );
OR2x2_ASAP7_75t_L g725 ( .A(n_537), .B(n_621), .Y(n_725) );
AND2x2_ASAP7_75t_L g538 ( .A(n_539), .B(n_542), .Y(n_538) );
INVx1_ASAP7_75t_L g607 ( .A(n_539), .Y(n_607) );
NAND2xp5_ASAP7_75t_L g688 ( .A(n_539), .B(n_689), .Y(n_688) );
AND2x2_ASAP7_75t_L g705 ( .A(n_539), .B(n_706), .Y(n_705) );
NAND2xp5_ASAP7_75t_L g730 ( .A(n_539), .B(n_586), .Y(n_730) );
INVx3_ASAP7_75t_L g539 ( .A(n_540), .Y(n_539) );
HB1xp67_ASAP7_75t_L g577 ( .A(n_540), .Y(n_577) );
INVx2_ASAP7_75t_L g540 ( .A(n_541), .Y(n_540) );
HB1xp67_ASAP7_75t_L g686 ( .A(n_541), .Y(n_686) );
AOI22xp5_ASAP7_75t_L g592 ( .A1(n_542), .A2(n_575), .B1(n_593), .B2(n_596), .Y(n_592) );
NOR2xp33_ASAP7_75t_L g676 ( .A(n_542), .B(n_677), .Y(n_676) );
INVx2_ASAP7_75t_SL g709 ( .A(n_542), .Y(n_709) );
AND2x4_ASAP7_75t_SL g542 ( .A(n_543), .B(n_555), .Y(n_542) );
HB1xp67_ASAP7_75t_L g543 ( .A(n_544), .Y(n_543) );
AND2x4_ASAP7_75t_L g586 ( .A(n_544), .B(n_587), .Y(n_586) );
INVx2_ASAP7_75t_L g606 ( .A(n_544), .Y(n_606) );
INVx1_ASAP7_75t_L g633 ( .A(n_544), .Y(n_633) );
AND2x2_ASAP7_75t_L g544 ( .A(n_545), .B(n_550), .Y(n_544) );
NOR3xp33_ASAP7_75t_L g546 ( .A(n_547), .B(n_548), .C(n_549), .Y(n_546) );
HB1xp67_ASAP7_75t_L g575 ( .A(n_555), .Y(n_575) );
AND2x4_ASAP7_75t_L g632 ( .A(n_555), .B(n_633), .Y(n_632) );
NOR2x1_ASAP7_75t_L g693 ( .A(n_555), .B(n_662), .Y(n_693) );
NAND2xp5_ASAP7_75t_L g556 ( .A(n_557), .B(n_559), .Y(n_556) );
AND2x2_ASAP7_75t_L g657 ( .A(n_557), .B(n_600), .Y(n_657) );
OAI21xp5_ASAP7_75t_L g737 ( .A1(n_557), .A2(n_738), .B(n_739), .Y(n_737) );
INVx2_ASAP7_75t_L g615 ( .A(n_558), .Y(n_615) );
AOI22xp5_ASAP7_75t_L g668 ( .A1(n_559), .A2(n_669), .B1(n_673), .B2(n_676), .Y(n_668) );
AND2x2_ASAP7_75t_L g559 ( .A(n_560), .B(n_562), .Y(n_559) );
HB1xp67_ASAP7_75t_L g626 ( .A(n_560), .Y(n_626) );
AND2x2_ASAP7_75t_L g636 ( .A(n_560), .B(n_637), .Y(n_636) );
INVx3_ASAP7_75t_L g675 ( .A(n_560), .Y(n_675) );
NAND2x1_ASAP7_75t_SL g700 ( .A(n_560), .B(n_569), .Y(n_700) );
AND2x2_ASAP7_75t_L g596 ( .A(n_562), .B(n_597), .Y(n_596) );
AND2x4_ASAP7_75t_L g562 ( .A(n_563), .B(n_565), .Y(n_562) );
INVx2_ASAP7_75t_L g563 ( .A(n_564), .Y(n_563) );
NOR2x1_ASAP7_75t_L g572 ( .A(n_564), .B(n_573), .Y(n_572) );
INVx1_ASAP7_75t_L g569 ( .A(n_565), .Y(n_569) );
INVx2_ASAP7_75t_L g581 ( .A(n_565), .Y(n_581) );
AOI21xp5_ASAP7_75t_SL g566 ( .A1(n_567), .A2(n_574), .B(n_578), .Y(n_566) );
INVx1_ASAP7_75t_L g567 ( .A(n_568), .Y(n_567) );
NAND2xp5_ASAP7_75t_L g568 ( .A(n_569), .B(n_570), .Y(n_568) );
NAND2xp5_ASAP7_75t_L g762 ( .A(n_569), .B(n_763), .Y(n_762) );
AOI22xp5_ASAP7_75t_L g658 ( .A1(n_570), .A2(n_659), .B1(n_663), .B2(n_666), .Y(n_658) );
AND2x2_ASAP7_75t_L g570 ( .A(n_571), .B(n_572), .Y(n_570) );
BUFx2_ASAP7_75t_L g763 ( .A(n_571), .Y(n_763) );
INVx1_ASAP7_75t_SL g770 ( .A(n_571), .Y(n_770) );
HB1xp67_ASAP7_75t_L g733 ( .A(n_572), .Y(n_733) );
NOR2xp33_ASAP7_75t_L g574 ( .A(n_575), .B(n_576), .Y(n_574) );
HB1xp67_ASAP7_75t_L g576 ( .A(n_577), .Y(n_576) );
OA21x2_ASAP7_75t_L g578 ( .A1(n_579), .A2(n_582), .B(n_585), .Y(n_578) );
AND2x2_ASAP7_75t_L g582 ( .A(n_580), .B(n_583), .Y(n_582) );
AND2x2_ASAP7_75t_L g624 ( .A(n_580), .B(n_620), .Y(n_624) );
AND2x2_ASAP7_75t_L g739 ( .A(n_580), .B(n_637), .Y(n_739) );
AND2x2_ASAP7_75t_L g742 ( .A(n_580), .B(n_648), .Y(n_742) );
AND2x4_ASAP7_75t_L g750 ( .A(n_580), .B(n_751), .Y(n_750) );
OAI21xp33_ASAP7_75t_L g704 ( .A1(n_582), .A2(n_705), .B(n_707), .Y(n_704) );
INVx2_ASAP7_75t_L g583 ( .A(n_584), .Y(n_583) );
INVx1_ASAP7_75t_L g732 ( .A(n_584), .Y(n_732) );
AND2x2_ASAP7_75t_L g748 ( .A(n_584), .B(n_749), .Y(n_748) );
INVx4_ASAP7_75t_L g662 ( .A(n_586), .Y(n_662) );
INVx1_ASAP7_75t_L g631 ( .A(n_587), .Y(n_631) );
AND2x2_ASAP7_75t_L g653 ( .A(n_587), .B(n_606), .Y(n_653) );
NOR2x1_ASAP7_75t_L g588 ( .A(n_589), .B(n_612), .Y(n_588) );
OAI21xp5_ASAP7_75t_L g589 ( .A1(n_590), .A2(n_592), .B(n_598), .Y(n_589) );
INVx1_ASAP7_75t_L g590 ( .A(n_591), .Y(n_590) );
AND2x2_ASAP7_75t_L g599 ( .A(n_591), .B(n_600), .Y(n_599) );
AND2x2_ASAP7_75t_SL g752 ( .A(n_591), .B(n_604), .Y(n_752) );
AND2x2_ASAP7_75t_L g773 ( .A(n_591), .B(n_689), .Y(n_773) );
INVx1_ASAP7_75t_L g593 ( .A(n_594), .Y(n_593) );
INVx2_ASAP7_75t_L g699 ( .A(n_596), .Y(n_699) );
OAI21xp5_ASAP7_75t_SL g598 ( .A1(n_599), .A2(n_601), .B(n_608), .Y(n_598) );
OR2x6_ASAP7_75t_L g651 ( .A(n_600), .B(n_652), .Y(n_651) );
INVx1_ASAP7_75t_L g601 ( .A(n_602), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g602 ( .A(n_603), .B(n_607), .Y(n_602) );
INVx2_ASAP7_75t_SL g603 ( .A(n_604), .Y(n_603) );
INVx2_ASAP7_75t_L g604 ( .A(n_605), .Y(n_604) );
INVx1_ASAP7_75t_L g605 ( .A(n_606), .Y(n_605) );
NOR2xp33_ASAP7_75t_L g608 ( .A(n_609), .B(n_610), .Y(n_608) );
OR2x2_ASAP7_75t_L g674 ( .A(n_609), .B(n_675), .Y(n_674) );
INVx1_ASAP7_75t_L g771 ( .A(n_609), .Y(n_771) );
NOR2xp33_ASAP7_75t_L g743 ( .A(n_610), .B(n_744), .Y(n_743) );
HB1xp67_ASAP7_75t_L g610 ( .A(n_611), .Y(n_610) );
NAND2xp5_ASAP7_75t_L g612 ( .A(n_613), .B(n_625), .Y(n_612) );
AOI22xp5_ASAP7_75t_L g613 ( .A1(n_614), .A2(n_616), .B1(n_622), .B2(n_624), .Y(n_613) );
OR2x2_ASAP7_75t_L g685 ( .A(n_615), .B(n_686), .Y(n_685) );
INVx3_ASAP7_75t_L g616 ( .A(n_617), .Y(n_616) );
HB1xp67_ASAP7_75t_L g642 ( .A(n_617), .Y(n_642) );
NAND2x1p5_ASAP7_75t_L g617 ( .A(n_618), .B(n_620), .Y(n_617) );
INVx1_ASAP7_75t_L g691 ( .A(n_620), .Y(n_691) );
INVx2_ASAP7_75t_SL g620 ( .A(n_621), .Y(n_620) );
INVxp67_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
AOI22xp5_ASAP7_75t_L g625 ( .A1(n_626), .A2(n_627), .B1(n_634), .B2(n_636), .Y(n_625) );
INVx1_ASAP7_75t_L g627 ( .A(n_628), .Y(n_627) );
NAND2xp5_ASAP7_75t_L g628 ( .A(n_629), .B(n_632), .Y(n_628) );
AND2x4_ASAP7_75t_SL g629 ( .A(n_630), .B(n_631), .Y(n_629) );
AND2x2_ASAP7_75t_L g634 ( .A(n_632), .B(n_635), .Y(n_634) );
AND2x2_ASAP7_75t_L g695 ( .A(n_635), .B(n_689), .Y(n_695) );
INVx1_ASAP7_75t_L g637 ( .A(n_638), .Y(n_637) );
NAND2xp5_ASAP7_75t_SL g639 ( .A(n_640), .B(n_680), .Y(n_639) );
NOR2xp67_ASAP7_75t_L g640 ( .A(n_641), .B(n_654), .Y(n_640) );
AOI21xp33_ASAP7_75t_SL g641 ( .A1(n_642), .A2(n_643), .B(n_649), .Y(n_641) );
OR2x2_ASAP7_75t_L g643 ( .A(n_644), .B(n_646), .Y(n_643) );
INVx3_ASAP7_75t_L g644 ( .A(n_645), .Y(n_644) );
NAND2x1p5_ASAP7_75t_L g646 ( .A(n_647), .B(n_648), .Y(n_646) );
INVx1_ASAP7_75t_L g649 ( .A(n_650), .Y(n_649) );
INVx2_ASAP7_75t_L g650 ( .A(n_651), .Y(n_650) );
OAI22xp33_ASAP7_75t_SL g719 ( .A1(n_651), .A2(n_720), .B1(n_722), .B2(n_725), .Y(n_719) );
NOR2x1_ASAP7_75t_L g666 ( .A(n_652), .B(n_667), .Y(n_666) );
INVx2_ASAP7_75t_L g652 ( .A(n_653), .Y(n_652) );
AND2x2_ASAP7_75t_L g702 ( .A(n_653), .B(n_703), .Y(n_702) );
OAI211xp5_ASAP7_75t_L g654 ( .A1(n_655), .A2(n_656), .B(n_658), .C(n_668), .Y(n_654) );
INVx2_ASAP7_75t_L g656 ( .A(n_657), .Y(n_656) );
NAND2xp33_ASAP7_75t_SL g659 ( .A(n_660), .B(n_662), .Y(n_659) );
INVxp33_ASAP7_75t_L g660 ( .A(n_661), .Y(n_660) );
INVx2_ASAP7_75t_L g671 ( .A(n_662), .Y(n_671) );
AOI221xp5_ASAP7_75t_L g682 ( .A1(n_663), .A2(n_683), .B1(n_684), .B2(n_687), .C(n_690), .Y(n_682) );
AND2x4_ASAP7_75t_L g663 ( .A(n_664), .B(n_665), .Y(n_663) );
INVx1_ASAP7_75t_L g723 ( .A(n_664), .Y(n_723) );
INVx2_ASAP7_75t_SL g721 ( .A(n_667), .Y(n_721) );
INVx1_ASAP7_75t_L g669 ( .A(n_670), .Y(n_669) );
NOR2xp33_ASAP7_75t_L g670 ( .A(n_671), .B(n_672), .Y(n_670) );
NAND2x1_ASAP7_75t_L g720 ( .A(n_671), .B(n_721), .Y(n_720) );
INVx1_ASAP7_75t_L g673 ( .A(n_674), .Y(n_673) );
INVx1_ASAP7_75t_L g717 ( .A(n_677), .Y(n_717) );
INVx1_ASAP7_75t_L g746 ( .A(n_678), .Y(n_746) );
INVx1_ASAP7_75t_L g678 ( .A(n_679), .Y(n_678) );
NOR2x1_ASAP7_75t_L g680 ( .A(n_681), .B(n_696), .Y(n_680) );
NAND2xp5_ASAP7_75t_L g681 ( .A(n_682), .B(n_694), .Y(n_681) );
INVx1_ASAP7_75t_L g684 ( .A(n_685), .Y(n_684) );
INVx1_ASAP7_75t_L g735 ( .A(n_686), .Y(n_735) );
INVx1_ASAP7_75t_L g687 ( .A(n_688), .Y(n_687) );
AND2x2_ASAP7_75t_L g756 ( .A(n_689), .B(n_757), .Y(n_756) );
INVx2_ASAP7_75t_L g761 ( .A(n_689), .Y(n_761) );
NOR2xp33_ASAP7_75t_L g690 ( .A(n_691), .B(n_692), .Y(n_690) );
INVxp33_ASAP7_75t_L g692 ( .A(n_693), .Y(n_692) );
BUFx2_ASAP7_75t_L g714 ( .A(n_693), .Y(n_714) );
OAI21xp5_ASAP7_75t_SL g696 ( .A1(n_697), .A2(n_701), .B(n_704), .Y(n_696) );
INVxp67_ASAP7_75t_L g697 ( .A(n_698), .Y(n_697) );
NAND2xp5_ASAP7_75t_L g698 ( .A(n_699), .B(n_700), .Y(n_698) );
INVx2_ASAP7_75t_L g701 ( .A(n_702), .Y(n_701) );
BUFx2_ASAP7_75t_L g757 ( .A(n_703), .Y(n_757) );
AND2x2_ASAP7_75t_L g745 ( .A(n_706), .B(n_746), .Y(n_745) );
NOR2xp33_ASAP7_75t_R g707 ( .A(n_708), .B(n_709), .Y(n_707) );
NAND3xp33_ASAP7_75t_L g710 ( .A(n_711), .B(n_726), .C(n_753), .Y(n_710) );
NOR2xp33_ASAP7_75t_L g711 ( .A(n_712), .B(n_719), .Y(n_711) );
NAND2xp5_ASAP7_75t_SL g712 ( .A(n_713), .B(n_716), .Y(n_712) );
NAND2xp5_ASAP7_75t_L g713 ( .A(n_714), .B(n_715), .Y(n_713) );
NAND2xp5_ASAP7_75t_L g716 ( .A(n_717), .B(n_718), .Y(n_716) );
OR2x2_ASAP7_75t_L g722 ( .A(n_723), .B(n_724), .Y(n_722) );
NOR2xp33_ASAP7_75t_L g726 ( .A(n_727), .B(n_740), .Y(n_726) );
NAND2xp5_ASAP7_75t_SL g727 ( .A(n_728), .B(n_737), .Y(n_727) );
AOI22xp33_ASAP7_75t_SL g728 ( .A1(n_729), .A2(n_731), .B1(n_733), .B2(n_734), .Y(n_728) );
INVx1_ASAP7_75t_L g729 ( .A(n_730), .Y(n_729) );
NOR2x1_ASAP7_75t_L g734 ( .A(n_735), .B(n_736), .Y(n_734) );
INVxp67_ASAP7_75t_SL g738 ( .A(n_736), .Y(n_738) );
NAND2xp5_ASAP7_75t_SL g740 ( .A(n_741), .B(n_747), .Y(n_740) );
OAI21xp5_ASAP7_75t_L g747 ( .A1(n_748), .A2(n_750), .B(n_752), .Y(n_747) );
INVx1_ASAP7_75t_L g766 ( .A(n_750), .Y(n_766) );
AOI211xp5_ASAP7_75t_L g753 ( .A1(n_754), .A2(n_756), .B(n_758), .C(n_767), .Y(n_753) );
INVx1_ASAP7_75t_L g754 ( .A(n_755), .Y(n_754) );
OAI22xp5_ASAP7_75t_L g758 ( .A1(n_759), .A2(n_762), .B1(n_764), .B2(n_766), .Y(n_758) );
NAND2xp5_ASAP7_75t_L g759 ( .A(n_760), .B(n_761), .Y(n_759) );
HB1xp67_ASAP7_75t_L g764 ( .A(n_765), .Y(n_764) );
NOR2xp33_ASAP7_75t_L g767 ( .A(n_768), .B(n_772), .Y(n_767) );
INVx1_ASAP7_75t_L g768 ( .A(n_769), .Y(n_768) );
AND2x2_ASAP7_75t_L g769 ( .A(n_770), .B(n_771), .Y(n_769) );
INVxp67_ASAP7_75t_L g772 ( .A(n_773), .Y(n_772) );
CKINVDCx11_ASAP7_75t_R g780 ( .A(n_774), .Y(n_780) );
INVx2_ASAP7_75t_L g779 ( .A(n_780), .Y(n_779) );
INVx1_ASAP7_75t_L g781 ( .A(n_782), .Y(n_781) );
INVx1_ASAP7_75t_SL g782 ( .A(n_783), .Y(n_782) );
INVx2_ASAP7_75t_L g783 ( .A(n_784), .Y(n_783) );
NAND2xp5_ASAP7_75t_L g785 ( .A(n_786), .B(n_789), .Y(n_785) );
CKINVDCx5p33_ASAP7_75t_R g786 ( .A(n_787), .Y(n_786) );
CKINVDCx20_ASAP7_75t_R g787 ( .A(n_788), .Y(n_787) );
INVxp67_ASAP7_75t_L g789 ( .A(n_790), .Y(n_789) );
AOI21xp5_ASAP7_75t_L g802 ( .A1(n_790), .A2(n_803), .B(n_808), .Y(n_802) );
NOR2xp33_ASAP7_75t_SL g790 ( .A(n_791), .B(n_796), .Y(n_790) );
INVx1_ASAP7_75t_SL g791 ( .A(n_792), .Y(n_791) );
BUFx2_ASAP7_75t_L g792 ( .A(n_793), .Y(n_792) );
CKINVDCx20_ASAP7_75t_R g793 ( .A(n_794), .Y(n_793) );
BUFx3_ASAP7_75t_L g794 ( .A(n_795), .Y(n_794) );
BUFx2_ASAP7_75t_L g809 ( .A(n_795), .Y(n_809) );
NAND2xp5_ASAP7_75t_L g797 ( .A(n_798), .B(n_802), .Y(n_797) );
CKINVDCx5p33_ASAP7_75t_R g798 ( .A(n_799), .Y(n_798) );
CKINVDCx11_ASAP7_75t_R g799 ( .A(n_800), .Y(n_799) );
CKINVDCx8_ASAP7_75t_R g800 ( .A(n_801), .Y(n_800) );
CKINVDCx20_ASAP7_75t_R g807 ( .A(n_804), .Y(n_807) );
HB1xp67_ASAP7_75t_L g808 ( .A(n_809), .Y(n_808) );
INVx2_ASAP7_75t_L g810 ( .A(n_811), .Y(n_810) );
INVx2_ASAP7_75t_SL g819 ( .A(n_811), .Y(n_819) );
INVx2_ASAP7_75t_L g811 ( .A(n_812), .Y(n_811) );
AND2x2_ASAP7_75t_SL g812 ( .A(n_813), .B(n_814), .Y(n_812) );
NOR2xp33_ASAP7_75t_L g817 ( .A(n_818), .B(n_819), .Y(n_817) );
endmodule