module real_jpeg_5032_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_367;
wire n_127;
wire n_365;
wire n_356;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_215;
wire n_166;
wire n_176;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_330;
wire n_298;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_360;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;
wire n_364;

AND2x2_ASAP7_75t_L g54 ( 
.A(n_0),
.B(n_55),
.Y(n_54)
);

AND2x2_ASAP7_75t_L g73 ( 
.A(n_0),
.B(n_74),
.Y(n_73)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_0),
.Y(n_105)
);

AND2x2_ASAP7_75t_L g157 ( 
.A(n_0),
.B(n_158),
.Y(n_157)
);

AND2x2_ASAP7_75t_L g271 ( 
.A(n_0),
.B(n_272),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_0),
.B(n_294),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_SL g361 ( 
.A(n_0),
.B(n_362),
.Y(n_361)
);

INVx8_ASAP7_75t_L g67 ( 
.A(n_1),
.Y(n_67)
);

AND2x2_ASAP7_75t_L g78 ( 
.A(n_2),
.B(n_79),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_2),
.B(n_113),
.Y(n_112)
);

AND2x2_ASAP7_75t_L g156 ( 
.A(n_2),
.B(n_94),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_2),
.B(n_218),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_2),
.B(n_259),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_2),
.B(n_322),
.Y(n_321)
);

CKINVDCx16_ASAP7_75t_R g344 ( 
.A(n_2),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_3),
.B(n_206),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_3),
.B(n_186),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_3),
.B(n_320),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_3),
.B(n_84),
.Y(n_354)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_4),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g77 ( 
.A(n_4),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g167 ( 
.A(n_4),
.Y(n_167)
);

AND2x2_ASAP7_75t_L g168 ( 
.A(n_5),
.B(n_37),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_5),
.B(n_186),
.Y(n_185)
);

AND2x2_ASAP7_75t_L g265 ( 
.A(n_5),
.B(n_266),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_5),
.B(n_285),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_5),
.B(n_290),
.Y(n_353)
);

AND2x2_ASAP7_75t_L g309 ( 
.A(n_6),
.B(n_310),
.Y(n_309)
);

AND2x2_ASAP7_75t_L g341 ( 
.A(n_6),
.B(n_342),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_7),
.B(n_37),
.Y(n_36)
);

AND2x2_ASAP7_75t_L g51 ( 
.A(n_7),
.B(n_52),
.Y(n_51)
);

AND2x2_ASAP7_75t_L g93 ( 
.A(n_7),
.B(n_94),
.Y(n_93)
);

AND2x2_ASAP7_75t_L g121 ( 
.A(n_7),
.B(n_122),
.Y(n_121)
);

AND2x2_ASAP7_75t_L g154 ( 
.A(n_7),
.B(n_155),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_7),
.B(n_209),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_SL g262 ( 
.A(n_7),
.B(n_147),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_SL g301 ( 
.A(n_7),
.B(n_302),
.Y(n_301)
);

INVx6_ASAP7_75t_L g92 ( 
.A(n_8),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_9),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_9),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_9),
.Y(n_110)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_9),
.Y(n_207)
);

BUFx6f_ASAP7_75t_L g310 ( 
.A(n_9),
.Y(n_310)
);

BUFx5_ASAP7_75t_L g149 ( 
.A(n_10),
.Y(n_149)
);

INVx3_ASAP7_75t_L g193 ( 
.A(n_10),
.Y(n_193)
);

INVx3_ASAP7_75t_L g295 ( 
.A(n_10),
.Y(n_295)
);

INVx8_ASAP7_75t_L g130 ( 
.A(n_11),
.Y(n_130)
);

AND2x2_ASAP7_75t_SL g239 ( 
.A(n_12),
.B(n_240),
.Y(n_239)
);

AND2x2_ASAP7_75t_L g306 ( 
.A(n_12),
.B(n_307),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_12),
.B(n_350),
.Y(n_349)
);

BUFx6f_ASAP7_75t_L g215 ( 
.A(n_13),
.Y(n_215)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_13),
.Y(n_237)
);

BUFx5_ASAP7_75t_L g304 ( 
.A(n_13),
.Y(n_304)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_14),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_14),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_14),
.Y(n_94)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_14),
.Y(n_270)
);

BUFx5_ASAP7_75t_L g320 ( 
.A(n_14),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_15),
.B(n_41),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_15),
.B(n_39),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_15),
.B(n_65),
.Y(n_64)
);

AND2x2_ASAP7_75t_L g87 ( 
.A(n_15),
.B(n_88),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_15),
.B(n_126),
.Y(n_125)
);

AND2x2_ASAP7_75t_L g146 ( 
.A(n_15),
.B(n_147),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_15),
.B(n_215),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_16),
.B(n_110),
.Y(n_109)
);

AND2x2_ASAP7_75t_L g163 ( 
.A(n_16),
.B(n_164),
.Y(n_163)
);

AND2x2_ASAP7_75t_SL g219 ( 
.A(n_16),
.B(n_220),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_16),
.B(n_253),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_16),
.B(n_290),
.Y(n_289)
);

AND2x2_ASAP7_75t_L g364 ( 
.A(n_16),
.B(n_365),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_17),
.B(n_31),
.Y(n_30)
);

AND2x2_ASAP7_75t_L g59 ( 
.A(n_17),
.B(n_60),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_17),
.B(n_84),
.Y(n_83)
);

AND2x2_ASAP7_75t_L g131 ( 
.A(n_17),
.B(n_132),
.Y(n_131)
);

AND2x2_ASAP7_75t_L g142 ( 
.A(n_17),
.B(n_143),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_17),
.B(n_190),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_17),
.B(n_236),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_331),
.Y(n_18)
);

HB1xp67_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

OAI21x1_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_278),
.B(n_330),
.Y(n_20)
);

AOI21x1_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_229),
.B(n_277),
.Y(n_21)
);

OAI21x1_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_173),
.B(n_228),
.Y(n_22)
);

AOI21x1_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_137),
.B(n_172),
.Y(n_23)
);

OAI21xp5_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_97),
.B(n_136),
.Y(n_24)
);

AOI21xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_69),
.B(n_96),
.Y(n_25)
);

OAI21xp5_ASAP7_75t_L g26 ( 
.A1(n_27),
.A2(n_46),
.B(n_68),
.Y(n_26)
);

AOI21xp5_ASAP7_75t_L g27 ( 
.A1(n_28),
.A2(n_43),
.B(n_45),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_SL g28 ( 
.A(n_29),
.B(n_40),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_29),
.B(n_40),
.Y(n_45)
);

XNOR2xp5_ASAP7_75t_L g29 ( 
.A(n_30),
.B(n_36),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_30),
.B(n_44),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_30),
.B(n_36),
.Y(n_47)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx1_ASAP7_75t_SL g32 ( 
.A(n_33),
.Y(n_32)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_34),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_35),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g188 ( 
.A(n_35),
.Y(n_188)
);

INVx3_ASAP7_75t_SL g37 ( 
.A(n_38),
.Y(n_37)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g240 ( 
.A(n_39),
.Y(n_240)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g221 ( 
.A(n_42),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_47),
.B(n_48),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_47),
.B(n_48),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_49),
.A2(n_50),
.B1(n_56),
.B2(n_57),
.Y(n_48)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_49),
.B(n_59),
.C(n_63),
.Y(n_95)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

XNOR2xp5_ASAP7_75t_SL g50 ( 
.A(n_51),
.B(n_54),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_51),
.B(n_54),
.Y(n_81)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_55),
.Y(n_80)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_58),
.A2(n_59),
.B1(n_63),
.B2(n_64),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_62),
.Y(n_107)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_67),
.Y(n_85)
);

INVx11_ASAP7_75t_L g123 ( 
.A(n_67),
.Y(n_123)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_67),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_70),
.B(n_95),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_70),
.B(n_95),
.Y(n_96)
);

XNOR2xp5_ASAP7_75t_L g70 ( 
.A(n_71),
.B(n_82),
.Y(n_70)
);

XOR2xp5_ASAP7_75t_L g71 ( 
.A(n_72),
.B(n_81),
.Y(n_71)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_72),
.B(n_81),
.C(n_99),
.Y(n_98)
);

XNOR2xp5_ASAP7_75t_L g72 ( 
.A(n_73),
.B(n_78),
.Y(n_72)
);

AND2x2_ASAP7_75t_L g102 ( 
.A(n_73),
.B(n_78),
.Y(n_102)
);

HB1xp67_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

BUFx5_ASAP7_75t_L g342 ( 
.A(n_77),
.Y(n_342)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVxp67_ASAP7_75t_L g99 ( 
.A(n_82),
.Y(n_99)
);

XOR2xp5_ASAP7_75t_L g82 ( 
.A(n_83),
.B(n_86),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_83),
.B(n_118),
.C(n_119),
.Y(n_117)
);

INVx5_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

XNOR2xp5_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_93),
.Y(n_86)
);

INVxp67_ASAP7_75t_L g118 ( 
.A(n_87),
.Y(n_118)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g182 ( 
.A(n_91),
.Y(n_182)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

BUFx3_ASAP7_75t_L g133 ( 
.A(n_92),
.Y(n_133)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_92),
.Y(n_155)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_92),
.Y(n_261)
);

INVx3_ASAP7_75t_L g292 ( 
.A(n_92),
.Y(n_292)
);

CKINVDCx14_ASAP7_75t_R g119 ( 
.A(n_93),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_98),
.B(n_100),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_98),
.B(n_100),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_L g100 ( 
.A(n_101),
.B(n_116),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_101),
.B(n_117),
.C(n_120),
.Y(n_171)
);

XOR2xp5_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_103),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_102),
.B(n_104),
.C(n_108),
.Y(n_151)
);

XOR2xp5_ASAP7_75t_L g103 ( 
.A(n_104),
.B(n_108),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_105),
.B(n_106),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_105),
.B(n_181),
.Y(n_180)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_109),
.A2(n_111),
.B1(n_112),
.B2(n_115),
.Y(n_108)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_109),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_111),
.B(n_115),
.Y(n_150)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVx8_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVx4_ASAP7_75t_L g307 ( 
.A(n_114),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_L g116 ( 
.A(n_117),
.B(n_120),
.Y(n_116)
);

XNOR2xp5_ASAP7_75t_L g120 ( 
.A(n_121),
.B(n_124),
.Y(n_120)
);

MAJx2_ASAP7_75t_L g170 ( 
.A(n_121),
.B(n_131),
.C(n_134),
.Y(n_170)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g218 ( 
.A(n_123),
.Y(n_218)
);

INVx6_ASAP7_75t_L g256 ( 
.A(n_123),
.Y(n_256)
);

INVx6_ASAP7_75t_L g287 ( 
.A(n_123),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_125),
.A2(n_131),
.B1(n_134),
.B2(n_135),
.Y(n_124)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_125),
.Y(n_134)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

INVx4_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVx3_ASAP7_75t_L g323 ( 
.A(n_128),
.Y(n_323)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVx6_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

BUFx5_ASAP7_75t_L g145 ( 
.A(n_130),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g211 ( 
.A(n_130),
.Y(n_211)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_130),
.Y(n_274)
);

INVx1_ASAP7_75t_SL g135 ( 
.A(n_131),
.Y(n_135)
);

INVx6_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_138),
.B(n_171),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_138),
.B(n_171),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_SL g138 ( 
.A(n_139),
.B(n_152),
.Y(n_138)
);

XOR2xp5_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_151),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_140),
.B(n_151),
.C(n_227),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g140 ( 
.A(n_141),
.B(n_150),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_146),
.Y(n_141)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_142),
.Y(n_201)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

HB1xp67_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

INVx6_ASAP7_75t_L g365 ( 
.A(n_145),
.Y(n_365)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_146),
.Y(n_202)
);

INVx4_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

INVx6_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

INVx3_ASAP7_75t_SL g345 ( 
.A(n_149),
.Y(n_345)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_150),
.B(n_201),
.C(n_202),
.Y(n_200)
);

INVxp67_ASAP7_75t_L g227 ( 
.A(n_152),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_160),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_153),
.B(n_162),
.C(n_169),
.Y(n_176)
);

BUFx24_ASAP7_75t_SL g373 ( 
.A(n_153),
.Y(n_373)
);

FAx1_ASAP7_75t_SL g153 ( 
.A(n_154),
.B(n_156),
.CI(n_157),
.CON(n_153),
.SN(n_153)
);

MAJx2_ASAP7_75t_L g198 ( 
.A(n_154),
.B(n_156),
.C(n_157),
.Y(n_198)
);

BUFx3_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_161),
.A2(n_162),
.B1(n_169),
.B2(n_170),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_168),
.Y(n_162)
);

AND2x2_ASAP7_75t_L g197 ( 
.A(n_163),
.B(n_168),
.Y(n_197)
);

INVx3_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

INVx5_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

INVx1_ASAP7_75t_SL g169 ( 
.A(n_170),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_SL g173 ( 
.A(n_174),
.B(n_226),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_174),
.B(n_226),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g174 ( 
.A(n_175),
.B(n_199),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_L g175 ( 
.A(n_176),
.B(n_177),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_176),
.B(n_177),
.C(n_199),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_178),
.A2(n_179),
.B1(n_195),
.B2(n_196),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_178),
.B(n_248),
.C(n_249),
.Y(n_247)
);

INVx1_ASAP7_75t_SL g178 ( 
.A(n_179),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_183),
.Y(n_179)
);

MAJx2_ASAP7_75t_L g243 ( 
.A(n_180),
.B(n_184),
.C(n_194),
.Y(n_243)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_184),
.A2(n_185),
.B1(n_189),
.B2(n_194),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

BUFx6f_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

INVx5_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_189),
.Y(n_194)
);

INVx3_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

INVx6_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

INVx5_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_198),
.Y(n_196)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_197),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_198),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_SL g199 ( 
.A(n_200),
.B(n_203),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_200),
.B(n_204),
.C(n_225),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_204),
.A2(n_213),
.B1(n_224),
.B2(n_225),
.Y(n_203)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_204),
.Y(n_224)
);

OAI21xp5_ASAP7_75t_L g204 ( 
.A1(n_205),
.A2(n_208),
.B(n_212),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_205),
.B(n_208),
.Y(n_212)
);

INVx3_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

INVx5_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

BUFx6f_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_212),
.B(n_243),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_212),
.B(n_233),
.C(n_243),
.Y(n_313)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_213),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_214),
.B(n_216),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_214),
.B(n_219),
.C(n_222),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_217),
.A2(n_219),
.B1(n_222),
.B2(n_223),
.Y(n_216)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_217),
.Y(n_222)
);

INVx1_ASAP7_75t_SL g223 ( 
.A(n_219),
.Y(n_223)
);

INVx4_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_230),
.B(n_276),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_230),
.B(n_276),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_SL g230 ( 
.A(n_231),
.B(n_246),
.Y(n_230)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_232),
.B(n_245),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_232),
.B(n_245),
.C(n_329),
.Y(n_328)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_233),
.A2(n_234),
.B1(n_242),
.B2(n_244),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_SL g234 ( 
.A(n_235),
.B(n_238),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_235),
.B(n_239),
.C(n_325),
.Y(n_324)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

INVx2_ASAP7_75t_L g363 ( 
.A(n_237),
.Y(n_363)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_239),
.B(n_241),
.Y(n_238)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_241),
.Y(n_325)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_242),
.Y(n_244)
);

INVxp67_ASAP7_75t_L g329 ( 
.A(n_246),
.Y(n_329)
);

XNOR2xp5_ASAP7_75t_SL g246 ( 
.A(n_247),
.B(n_250),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_247),
.B(n_251),
.C(n_263),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_251),
.B(n_263),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_252),
.B(n_257),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_252),
.B(n_258),
.C(n_262),
.Y(n_298)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

INVx3_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

INVx6_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_258),
.B(n_262),
.Y(n_257)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g263 ( 
.A(n_264),
.B(n_275),
.Y(n_263)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_265),
.B(n_271),
.Y(n_264)
);

MAJx2_ASAP7_75t_L g315 ( 
.A(n_265),
.B(n_271),
.C(n_316),
.Y(n_315)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

INVx4_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

BUFx3_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

BUFx5_ASAP7_75t_L g351 ( 
.A(n_270),
.Y(n_351)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

INVx6_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

INVx1_ASAP7_75t_SL g316 ( 
.A(n_275),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_SL g278 ( 
.A(n_279),
.B(n_328),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_279),
.B(n_328),
.Y(n_330)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_280),
.B(n_281),
.Y(n_279)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_280),
.Y(n_370)
);

XOR2xp5_ASAP7_75t_L g281 ( 
.A(n_282),
.B(n_312),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g369 ( 
.A(n_282),
.B(n_312),
.C(n_370),
.Y(n_369)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_283),
.B(n_296),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g356 ( 
.A(n_283),
.B(n_297),
.C(n_300),
.Y(n_356)
);

XNOR2xp5_ASAP7_75t_SL g283 ( 
.A(n_284),
.B(n_288),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g368 ( 
.A(n_284),
.B(n_289),
.C(n_293),
.Y(n_368)
);

BUFx2_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

INVx8_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g288 ( 
.A(n_289),
.B(n_293),
.Y(n_288)
);

INVx6_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

INVx4_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

INVx6_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_L g296 ( 
.A1(n_297),
.A2(n_298),
.B1(n_299),
.B2(n_300),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_300),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_L g300 ( 
.A(n_301),
.B(n_305),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g347 ( 
.A(n_301),
.B(n_306),
.C(n_309),
.Y(n_347)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_303),
.Y(n_302)
);

INVx8_ASAP7_75t_L g303 ( 
.A(n_304),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_L g305 ( 
.A1(n_306),
.A2(n_308),
.B1(n_309),
.B2(n_311),
.Y(n_305)
);

CKINVDCx14_ASAP7_75t_R g311 ( 
.A(n_306),
.Y(n_311)
);

OAI22xp5_ASAP7_75t_SL g339 ( 
.A1(n_308),
.A2(n_309),
.B1(n_340),
.B2(n_341),
.Y(n_339)
);

CKINVDCx14_ASAP7_75t_R g308 ( 
.A(n_309),
.Y(n_308)
);

XOR2xp5_ASAP7_75t_L g312 ( 
.A(n_313),
.B(n_314),
.Y(n_312)
);

INVxp67_ASAP7_75t_L g335 ( 
.A(n_313),
.Y(n_335)
);

AOI22xp33_ASAP7_75t_L g314 ( 
.A1(n_315),
.A2(n_317),
.B1(n_326),
.B2(n_327),
.Y(n_314)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_315),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_315),
.B(n_327),
.C(n_335),
.Y(n_334)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_317),
.Y(n_327)
);

XNOR2xp5_ASAP7_75t_L g317 ( 
.A(n_318),
.B(n_324),
.Y(n_317)
);

XNOR2xp5_ASAP7_75t_L g318 ( 
.A(n_319),
.B(n_321),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g358 ( 
.A(n_319),
.B(n_321),
.C(n_324),
.Y(n_358)
);

INVx5_ASAP7_75t_L g322 ( 
.A(n_323),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_332),
.B(n_371),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_SL g332 ( 
.A(n_333),
.B(n_369),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g372 ( 
.A(n_333),
.B(n_369),
.Y(n_372)
);

XNOR2xp5_ASAP7_75t_L g333 ( 
.A(n_334),
.B(n_336),
.Y(n_333)
);

XNOR2xp5_ASAP7_75t_L g336 ( 
.A(n_337),
.B(n_355),
.Y(n_336)
);

XOR2xp5_ASAP7_75t_L g337 ( 
.A(n_338),
.B(n_346),
.Y(n_337)
);

XNOR2xp5_ASAP7_75t_SL g338 ( 
.A(n_339),
.B(n_343),
.Y(n_338)
);

CKINVDCx20_ASAP7_75t_R g340 ( 
.A(n_341),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_L g343 ( 
.A(n_344),
.B(n_345),
.Y(n_343)
);

XNOR2xp5_ASAP7_75t_L g346 ( 
.A(n_347),
.B(n_348),
.Y(n_346)
);

XNOR2xp5_ASAP7_75t_L g348 ( 
.A(n_349),
.B(n_352),
.Y(n_348)
);

INVx3_ASAP7_75t_L g350 ( 
.A(n_351),
.Y(n_350)
);

XNOR2xp5_ASAP7_75t_L g352 ( 
.A(n_353),
.B(n_354),
.Y(n_352)
);

XNOR2xp5_ASAP7_75t_SL g355 ( 
.A(n_356),
.B(n_357),
.Y(n_355)
);

XNOR2xp5_ASAP7_75t_L g357 ( 
.A(n_358),
.B(n_359),
.Y(n_357)
);

XNOR2xp5_ASAP7_75t_L g359 ( 
.A(n_360),
.B(n_368),
.Y(n_359)
);

AOI22xp5_ASAP7_75t_L g360 ( 
.A1(n_361),
.A2(n_364),
.B1(n_366),
.B2(n_367),
.Y(n_360)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_361),
.Y(n_366)
);

BUFx6f_ASAP7_75t_L g362 ( 
.A(n_363),
.Y(n_362)
);

CKINVDCx14_ASAP7_75t_R g367 ( 
.A(n_364),
.Y(n_367)
);

INVxp67_ASAP7_75t_L g371 ( 
.A(n_372),
.Y(n_371)
);


endmodule