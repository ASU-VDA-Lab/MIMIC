module real_jpeg_10940_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_68;
wire n_146;
wire n_247;
wire n_78;
wire n_83;
wire n_249;
wire n_166;
wire n_176;
wire n_221;
wire n_215;
wire n_194;
wire n_104;
wire n_153;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_173;
wire n_40;
wire n_105;
wire n_243;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_120;
wire n_113;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_242;
wire n_141;
wire n_65;
wire n_188;
wire n_33;
wire n_139;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_195;
wire n_205;
wire n_110;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_204;
wire n_158;
wire n_149;
wire n_144;
wire n_130;
wire n_241;
wire n_103;
wire n_225;
wire n_232;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_185;
wire n_125;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_187;
wire n_75;
wire n_97;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_167;
wire n_244;
wire n_213;
wire n_179;
wire n_202;
wire n_133;
wire n_216;
wire n_138;
wire n_25;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;

BUFx24_ASAP7_75t_L g54 ( 
.A(n_0),
.Y(n_54)
);

OAI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_1),
.A2(n_54),
.B1(n_55),
.B2(n_56),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_1),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_L g89 ( 
.A1(n_1),
.A2(n_38),
.B1(n_39),
.B2(n_55),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_L g163 ( 
.A1(n_1),
.A2(n_28),
.B1(n_32),
.B2(n_55),
.Y(n_163)
);

INVx2_ASAP7_75t_SL g67 ( 
.A(n_2),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_2),
.A2(n_54),
.B1(n_56),
.B2(n_67),
.Y(n_69)
);

AOI21xp33_ASAP7_75t_L g115 ( 
.A1(n_2),
.A2(n_3),
.B(n_54),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_3),
.Y(n_114)
);

OAI22xp33_ASAP7_75t_SL g139 ( 
.A1(n_3),
.A2(n_66),
.B1(n_71),
.B2(n_114),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_3),
.B(n_74),
.Y(n_160)
);

A2O1A1O1Ixp25_ASAP7_75t_L g172 ( 
.A1(n_3),
.A2(n_38),
.B(n_42),
.C(n_173),
.D(n_174),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_3),
.B(n_38),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_3),
.B(n_61),
.Y(n_182)
);

OAI21xp33_ASAP7_75t_L g207 ( 
.A1(n_3),
.A2(n_26),
.B(n_188),
.Y(n_207)
);

A2O1A1O1Ixp25_ASAP7_75t_L g220 ( 
.A1(n_3),
.A2(n_56),
.B(n_57),
.C(n_123),
.D(n_221),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_3),
.B(n_56),
.Y(n_221)
);

INVx2_ASAP7_75t_SL g27 ( 
.A(n_4),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_4),
.B(n_189),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_4),
.A2(n_194),
.B1(n_196),
.B2(n_197),
.Y(n_193)
);

AOI21xp5_ASAP7_75t_L g228 ( 
.A1(n_4),
.A2(n_205),
.B(n_229),
.Y(n_228)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

BUFx10_ASAP7_75t_L g44 ( 
.A(n_6),
.Y(n_44)
);

BUFx6f_ASAP7_75t_SL g59 ( 
.A(n_7),
.Y(n_59)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_8),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_L g31 ( 
.A1(n_9),
.A2(n_28),
.B1(n_32),
.B2(n_33),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_9),
.Y(n_33)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_9),
.A2(n_33),
.B1(n_38),
.B2(n_39),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_L g47 ( 
.A1(n_10),
.A2(n_38),
.B1(n_39),
.B2(n_48),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_10),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_10),
.A2(n_28),
.B1(n_32),
.B2(n_48),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_11),
.A2(n_66),
.B1(n_71),
.B2(n_93),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_11),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g143 ( 
.A1(n_11),
.A2(n_54),
.B1(n_56),
.B2(n_93),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_SL g185 ( 
.A1(n_11),
.A2(n_38),
.B1(n_39),
.B2(n_93),
.Y(n_185)
);

AOI22xp33_ASAP7_75t_SL g195 ( 
.A1(n_11),
.A2(n_28),
.B1(n_32),
.B2(n_93),
.Y(n_195)
);

OAI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_12),
.A2(n_66),
.B1(n_71),
.B2(n_76),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_12),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_L g100 ( 
.A1(n_12),
.A2(n_54),
.B1(n_56),
.B2(n_76),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_L g137 ( 
.A1(n_12),
.A2(n_38),
.B1(n_39),
.B2(n_76),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_12),
.A2(n_28),
.B1(n_32),
.B2(n_76),
.Y(n_190)
);

BUFx10_ASAP7_75t_L g66 ( 
.A(n_13),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g37 ( 
.A1(n_14),
.A2(n_38),
.B1(n_39),
.B2(n_40),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_14),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_14),
.A2(n_40),
.B1(n_54),
.B2(n_56),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_14),
.A2(n_28),
.B1(n_32),
.B2(n_40),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_15),
.A2(n_66),
.B1(n_71),
.B2(n_72),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_15),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_15),
.A2(n_54),
.B1(n_56),
.B2(n_72),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_SL g187 ( 
.A1(n_15),
.A2(n_28),
.B1(n_32),
.B2(n_72),
.Y(n_187)
);

AOI22xp33_ASAP7_75t_L g219 ( 
.A1(n_15),
.A2(n_38),
.B1(n_39),
.B2(n_72),
.Y(n_219)
);

AOI22xp33_ASAP7_75t_SL g34 ( 
.A1(n_16),
.A2(n_28),
.B1(n_32),
.B2(n_35),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_16),
.Y(n_35)
);

XNOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_126),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_124),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_SL g19 ( 
.A(n_20),
.B(n_101),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_20),
.B(n_101),
.Y(n_125)
);

XOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_84),
.Y(n_20)
);

OAI22xp5_ASAP7_75t_SL g21 ( 
.A1(n_22),
.A2(n_23),
.B1(n_77),
.B2(n_78),
.Y(n_21)
);

CKINVDCx16_ASAP7_75t_R g22 ( 
.A(n_23),
.Y(n_22)
);

XOR2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_50),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_36),
.Y(n_24)
);

XNOR2xp5_ASAP7_75t_L g104 ( 
.A(n_25),
.B(n_36),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_27),
.B1(n_31),
.B2(n_34),
.Y(n_25)
);

AOI21xp5_ASAP7_75t_L g80 ( 
.A1(n_26),
.A2(n_27),
.B(n_34),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_26),
.A2(n_27),
.B1(n_31),
.B2(n_87),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_26),
.A2(n_27),
.B1(n_87),
.B2(n_117),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_26),
.A2(n_27),
.B1(n_117),
.B2(n_163),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_SL g186 ( 
.A1(n_26),
.A2(n_187),
.B(n_188),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_26),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_26),
.B(n_190),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_28),
.Y(n_26)
);

OAI21xp5_ASAP7_75t_L g203 ( 
.A1(n_27),
.A2(n_195),
.B(n_204),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_27),
.B(n_114),
.Y(n_209)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_28),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_L g46 ( 
.A1(n_28),
.A2(n_32),
.B1(n_43),
.B2(n_44),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_28),
.A2(n_45),
.B1(n_177),
.B2(n_178),
.Y(n_176)
);

BUFx2_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

BUFx24_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_SL g177 ( 
.A(n_32),
.B(n_43),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_SL g208 ( 
.A(n_32),
.B(n_209),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_L g36 ( 
.A1(n_37),
.A2(n_41),
.B1(n_47),
.B2(n_49),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_37),
.A2(n_41),
.B1(n_49),
.B2(n_89),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_38),
.A2(n_39),
.B1(n_58),
.B2(n_59),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_38),
.A2(n_221),
.B1(n_226),
.B2(n_227),
.Y(n_225)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

O2A1O1Ixp33_ASAP7_75t_L g42 ( 
.A1(n_39),
.A2(n_43),
.B(n_45),
.C(n_46),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_39),
.B(n_43),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_39),
.B(n_59),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_41),
.A2(n_47),
.B1(n_49),
.B2(n_82),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g218 ( 
.A1(n_41),
.A2(n_49),
.B1(n_185),
.B2(n_219),
.Y(n_218)
);

OAI21xp5_ASAP7_75t_SL g241 ( 
.A1(n_41),
.A2(n_219),
.B(n_242),
.Y(n_241)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_42),
.B(n_136),
.Y(n_135)
);

CKINVDCx16_ASAP7_75t_R g43 ( 
.A(n_44),
.Y(n_43)
);

CKINVDCx16_ASAP7_75t_R g49 ( 
.A(n_46),
.Y(n_49)
);

OAI21xp5_ASAP7_75t_L g134 ( 
.A1(n_49),
.A2(n_89),
.B(n_135),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_49),
.B(n_137),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_L g184 ( 
.A1(n_49),
.A2(n_135),
.B(n_185),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_SL g202 ( 
.A(n_49),
.B(n_114),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_L g50 ( 
.A1(n_51),
.A2(n_52),
.B1(n_63),
.B2(n_64),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_52),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_L g52 ( 
.A1(n_53),
.A2(n_57),
.B1(n_61),
.B2(n_62),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_53),
.Y(n_96)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_54),
.Y(n_56)
);

O2A1O1Ixp33_ASAP7_75t_SL g57 ( 
.A1(n_54),
.A2(n_58),
.B(n_60),
.C(n_61),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_54),
.B(n_58),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_57),
.B(n_99),
.Y(n_98)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_57),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_59),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_60),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_61),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_64),
.Y(n_63)
);

OAI21xp5_ASAP7_75t_SL g64 ( 
.A1(n_65),
.A2(n_70),
.B(n_73),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_65),
.A2(n_69),
.B1(n_70),
.B2(n_92),
.Y(n_91)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_65),
.Y(n_110)
);

A2O1A1Ixp33_ASAP7_75t_L g65 ( 
.A1(n_66),
.A2(n_67),
.B(n_68),
.C(n_69),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_66),
.B(n_67),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_66),
.Y(n_71)
);

A2O1A1Ixp33_ASAP7_75t_L g113 ( 
.A1(n_66),
.A2(n_67),
.B(n_114),
.C(n_115),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_69),
.Y(n_74)
);

OAI21xp33_ASAP7_75t_L g108 ( 
.A1(n_69),
.A2(n_92),
.B(n_109),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_73),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_74),
.B(n_75),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_75),
.B(n_110),
.Y(n_109)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_79),
.A2(n_80),
.B1(n_81),
.B2(n_83),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_80),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_81),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_85),
.B(n_90),
.C(n_94),
.Y(n_84)
);

XOR2xp5_ASAP7_75t_L g102 ( 
.A(n_85),
.B(n_103),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_86),
.B(n_88),
.Y(n_85)
);

XOR2xp5_ASAP7_75t_L g131 ( 
.A(n_86),
.B(n_88),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_90),
.A2(n_91),
.B1(n_94),
.B2(n_95),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_91),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_95),
.Y(n_94)
);

OAI21xp5_ASAP7_75t_L g95 ( 
.A1(n_96),
.A2(n_97),
.B(n_98),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_97),
.B(n_100),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_97),
.A2(n_120),
.B1(n_121),
.B2(n_143),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_L g159 ( 
.A1(n_97),
.A2(n_98),
.B(n_143),
.Y(n_159)
);

CKINVDCx16_ASAP7_75t_R g99 ( 
.A(n_100),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_104),
.C(n_105),
.Y(n_101)
);

XOR2xp5_ASAP7_75t_L g148 ( 
.A(n_102),
.B(n_104),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_105),
.A2(n_106),
.B1(n_147),
.B2(n_148),
.Y(n_146)
);

CKINVDCx16_ASAP7_75t_R g105 ( 
.A(n_106),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_107),
.B(n_111),
.C(n_118),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_107),
.A2(n_108),
.B1(n_118),
.B2(n_119),
.Y(n_145)
);

CKINVDCx16_ASAP7_75t_R g107 ( 
.A(n_108),
.Y(n_107)
);

AOI21xp5_ASAP7_75t_L g138 ( 
.A1(n_110),
.A2(n_139),
.B(n_140),
.Y(n_138)
);

XOR2xp5_ASAP7_75t_L g144 ( 
.A(n_111),
.B(n_145),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_112),
.B(n_116),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_112),
.A2(n_113),
.B1(n_116),
.B2(n_155),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_113),
.Y(n_112)
);

CKINVDCx16_ASAP7_75t_R g155 ( 
.A(n_116),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_119),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_L g119 ( 
.A1(n_120),
.A2(n_121),
.B(n_122),
.Y(n_119)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_165),
.Y(n_126)
);

INVxp33_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

AOI21xp33_ASAP7_75t_L g128 ( 
.A1(n_129),
.A2(n_149),
.B(n_164),
.Y(n_128)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_129),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_146),
.Y(n_129)
);

CKINVDCx5p33_ASAP7_75t_R g150 ( 
.A(n_130),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_130),
.B(n_146),
.Y(n_164)
);

FAx1_ASAP7_75t_SL g130 ( 
.A(n_131),
.B(n_132),
.CI(n_144),
.CON(n_130),
.SN(n_130)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_133),
.B(n_138),
.C(n_141),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_133),
.A2(n_134),
.B1(n_141),
.B2(n_142),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_134),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_137),
.Y(n_136)
);

XOR2xp5_ASAP7_75t_L g152 ( 
.A(n_138),
.B(n_153),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_142),
.Y(n_141)
);

CKINVDCx16_ASAP7_75t_R g147 ( 
.A(n_148),
.Y(n_147)
);

AND2x2_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_151),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_150),
.B(n_151),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_154),
.C(n_156),
.Y(n_151)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_152),
.B(n_247),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_L g247 ( 
.A1(n_154),
.A2(n_156),
.B1(n_157),
.B2(n_248),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_154),
.Y(n_248)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_160),
.C(n_161),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_158),
.A2(n_159),
.B1(n_236),
.B2(n_238),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_159),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_160),
.A2(n_161),
.B1(n_162),
.B2(n_237),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_160),
.Y(n_237)
);

CKINVDCx16_ASAP7_75t_R g161 ( 
.A(n_162),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_163),
.Y(n_229)
);

NOR3xp33_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_250),
.C(n_251),
.Y(n_165)
);

AOI21xp5_ASAP7_75t_L g166 ( 
.A1(n_167),
.A2(n_244),
.B(n_249),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_SL g167 ( 
.A1(n_168),
.A2(n_232),
.B(n_243),
.Y(n_167)
);

AOI21xp5_ASAP7_75t_L g168 ( 
.A1(n_169),
.A2(n_213),
.B(n_231),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_SL g169 ( 
.A1(n_170),
.A2(n_191),
.B(n_212),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_179),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_171),
.B(n_179),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_SL g171 ( 
.A(n_172),
.B(n_175),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_172),
.A2(n_175),
.B1(n_176),
.B2(n_199),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_172),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_173),
.Y(n_178)
);

INVxp67_ASAP7_75t_L g242 ( 
.A(n_174),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_176),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_186),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_181),
.A2(n_182),
.B1(n_183),
.B2(n_184),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_181),
.B(n_184),
.C(n_186),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_182),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_184),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_187),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_190),
.Y(n_189)
);

AOI21xp5_ASAP7_75t_L g191 ( 
.A1(n_192),
.A2(n_200),
.B(n_211),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_193),
.B(n_198),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_SL g211 ( 
.A(n_193),
.B(n_198),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_195),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_SL g200 ( 
.A1(n_201),
.A2(n_206),
.B(n_210),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_202),
.B(n_203),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_202),
.B(n_203),
.Y(n_210)
);

INVxp67_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_207),
.B(n_208),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_214),
.B(n_215),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_SL g231 ( 
.A(n_214),
.B(n_215),
.Y(n_231)
);

AOI22xp33_ASAP7_75t_SL g215 ( 
.A1(n_216),
.A2(n_217),
.B1(n_224),
.B2(n_230),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_L g217 ( 
.A1(n_218),
.A2(n_220),
.B1(n_222),
.B2(n_223),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_218),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_220),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_220),
.B(n_223),
.C(n_230),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_224),
.Y(n_230)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_225),
.B(n_228),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_225),
.B(n_228),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_233),
.B(n_234),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_SL g243 ( 
.A(n_233),
.B(n_234),
.Y(n_243)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_235),
.B(n_239),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_235),
.B(n_240),
.C(n_241),
.Y(n_245)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_236),
.Y(n_238)
);

XOR2xp5_ASAP7_75t_L g239 ( 
.A(n_240),
.B(n_241),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_245),
.B(n_246),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_SL g249 ( 
.A(n_245),
.B(n_246),
.Y(n_249)
);


endmodule