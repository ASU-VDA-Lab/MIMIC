module real_jpeg_5117_n_14 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_2, n_13, n_6, n_7, n_3, n_10, n_9, n_14);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_2;
input n_13;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_14;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_18;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_16;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_15;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

INVx8_ASAP7_75t_L g49 ( 
.A(n_0),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_1),
.Y(n_70)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_1),
.Y(n_73)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_1),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_1),
.Y(n_83)
);

BUFx5_ASAP7_75t_L g91 ( 
.A(n_1),
.Y(n_91)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_1),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g172 ( 
.A(n_1),
.Y(n_172)
);

OAI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_2),
.A2(n_56),
.B1(n_59),
.B2(n_60),
.Y(n_55)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_2),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_L g144 ( 
.A1(n_2),
.A2(n_59),
.B1(n_145),
.B2(n_148),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_2),
.A2(n_59),
.B1(n_153),
.B2(n_157),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_2),
.A2(n_59),
.B1(n_91),
.B2(n_180),
.Y(n_179)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_3),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_3),
.Y(n_115)
);

BUFx3_ASAP7_75t_L g137 ( 
.A(n_3),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_4),
.A2(n_126),
.B1(n_127),
.B2(n_130),
.Y(n_125)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_4),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_4),
.A2(n_126),
.B1(n_208),
.B2(n_210),
.Y(n_207)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

INVx8_ASAP7_75t_L g140 ( 
.A(n_6),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g143 ( 
.A(n_6),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g163 ( 
.A(n_6),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g200 ( 
.A(n_6),
.Y(n_200)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_7),
.Y(n_79)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_7),
.Y(n_88)
);

BUFx5_ASAP7_75t_L g169 ( 
.A(n_7),
.Y(n_169)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_8),
.Y(n_35)
);

INVx3_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

AOI22xp5_ASAP7_75t_L g14 ( 
.A1(n_10),
.A2(n_15),
.B1(n_18),
.B2(n_19),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_11),
.Y(n_103)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_11),
.Y(n_106)
);

BUFx3_ASAP7_75t_L g117 ( 
.A(n_11),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_12),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_12),
.A2(n_47),
.B1(n_69),
.B2(n_121),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_12),
.A2(n_69),
.B1(n_187),
.B2(n_188),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_12),
.A2(n_69),
.B1(n_113),
.B2(n_203),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_12),
.B(n_84),
.Y(n_238)
);

O2A1O1Ixp33_ASAP7_75t_L g252 ( 
.A1(n_12),
.A2(n_253),
.B(n_255),
.C(n_263),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_12),
.B(n_281),
.C(n_283),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_12),
.B(n_65),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_12),
.B(n_163),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_12),
.B(n_110),
.Y(n_318)
);

OAI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_13),
.A2(n_56),
.B1(n_60),
.B2(n_64),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_13),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_13),
.A2(n_64),
.B1(n_91),
.B2(n_92),
.Y(n_90)
);

OAI22xp33_ASAP7_75t_SL g271 ( 
.A1(n_13),
.A2(n_64),
.B1(n_122),
.B2(n_259),
.Y(n_271)
);

AOI22xp33_ASAP7_75t_L g290 ( 
.A1(n_13),
.A2(n_64),
.B1(n_291),
.B2(n_295),
.Y(n_290)
);

INVx3_ASAP7_75t_L g15 ( 
.A(n_16),
.Y(n_15)
);

INVx5_ASAP7_75t_L g16 ( 
.A(n_17),
.Y(n_16)
);

INVx6_ASAP7_75t_L g18 ( 
.A(n_17),
.Y(n_18)
);

XNOR2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_225),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_223),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_192),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_SL g224 ( 
.A(n_22),
.B(n_192),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_22),
.B(n_227),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_22),
.B(n_227),
.Y(n_341)
);

FAx1_ASAP7_75t_SL g22 ( 
.A(n_23),
.B(n_123),
.CI(n_158),
.CON(n_22),
.SN(n_22)
);

MAJIxp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_66),
.C(n_96),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_L g229 ( 
.A1(n_24),
.A2(n_96),
.B1(n_230),
.B2(n_231),
.Y(n_229)
);

INVxp67_ASAP7_75t_L g231 ( 
.A(n_24),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_SL g24 ( 
.A(n_25),
.B(n_62),
.Y(n_24)
);

INVxp67_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_SL g26 ( 
.A(n_27),
.B(n_54),
.Y(n_26)
);

INVx1_ASAP7_75t_SL g191 ( 
.A(n_27),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_41),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_L g28 ( 
.A1(n_29),
.A2(n_32),
.B1(n_36),
.B2(n_38),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g254 ( 
.A(n_30),
.Y(n_254)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_31),
.Y(n_37)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_31),
.Y(n_44)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_31),
.Y(n_53)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_34),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_34),
.Y(n_87)
);

BUFx5_ASAP7_75t_L g167 ( 
.A(n_34),
.Y(n_167)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_35),
.Y(n_58)
);

BUFx5_ASAP7_75t_L g61 ( 
.A(n_35),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_35),
.Y(n_86)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx4_ASAP7_75t_SL g38 ( 
.A(n_39),
.Y(n_38)
);

INVx5_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_41),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_41),
.B(n_185),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g41 ( 
.A1(n_42),
.A2(n_45),
.B1(n_50),
.B2(n_52),
.Y(n_41)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx4_ASAP7_75t_L g258 ( 
.A(n_44),
.Y(n_258)
);

INVx3_ASAP7_75t_SL g45 ( 
.A(n_46),
.Y(n_45)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_48),
.Y(n_122)
);

INVx6_ASAP7_75t_L g156 ( 
.A(n_48),
.Y(n_156)
);

INVx5_ASAP7_75t_L g213 ( 
.A(n_48),
.Y(n_213)
);

INVx11_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_49),
.Y(n_51)
);

BUFx5_ASAP7_75t_L g101 ( 
.A(n_49),
.Y(n_101)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_49),
.Y(n_109)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_49),
.Y(n_262)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx3_ASAP7_75t_L g209 ( 
.A(n_51),
.Y(n_209)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_55),
.B(n_65),
.Y(n_236)
);

INVx5_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx3_ASAP7_75t_L g189 ( 
.A(n_58),
.Y(n_189)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_58),
.Y(n_264)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx5_ASAP7_75t_L g187 ( 
.A(n_61),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_62),
.B(n_329),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_63),
.B(n_65),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_63),
.B(n_191),
.Y(n_190)
);

OAI21xp5_ASAP7_75t_L g218 ( 
.A1(n_65),
.A2(n_186),
.B(n_191),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_SL g228 ( 
.A(n_66),
.B(n_229),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_67),
.B(n_89),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_68),
.B(n_74),
.Y(n_67)
);

OAI21xp5_ASAP7_75t_L g68 ( 
.A1(n_69),
.A2(n_70),
.B(n_71),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_69),
.B(n_72),
.Y(n_71)
);

OAI21xp33_ASAP7_75t_L g255 ( 
.A1(n_69),
.A2(n_256),
.B(n_259),
.Y(n_255)
);

INVxp33_ASAP7_75t_L g173 ( 
.A(n_71),
.Y(n_173)
);

INVx5_ASAP7_75t_L g180 ( 
.A(n_72),
.Y(n_180)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_74),
.B(n_90),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_74),
.B(n_179),
.Y(n_220)
);

NOR2x1_ASAP7_75t_L g74 ( 
.A(n_75),
.B(n_84),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_76),
.A2(n_78),
.B1(n_80),
.B2(n_82),
.Y(n_75)
);

INVx6_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_79),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_79),
.Y(n_85)
);

NAND2xp33_ASAP7_75t_SL g174 ( 
.A(n_80),
.B(n_175),
.Y(n_174)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_84),
.B(n_90),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_84),
.B(n_179),
.Y(n_178)
);

AO22x1_ASAP7_75t_SL g84 ( 
.A1(n_85),
.A2(n_86),
.B1(n_87),
.B2(n_88),
.Y(n_84)
);

INVx4_ASAP7_75t_L g175 ( 
.A(n_86),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_89),
.B(n_220),
.Y(n_219)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_96),
.Y(n_230)
);

AOI21xp5_ASAP7_75t_L g96 ( 
.A1(n_97),
.A2(n_118),
.B(n_119),
.Y(n_96)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_98),
.B(n_120),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_98),
.B(n_152),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_98),
.B(n_271),
.Y(n_270)
);

NOR2x1_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_110),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_100),
.A2(n_102),
.B1(n_104),
.B2(n_107),
.Y(n_99)
);

INVx5_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

AO22x1_ASAP7_75t_SL g110 ( 
.A1(n_103),
.A2(n_111),
.B1(n_113),
.B2(n_116),
.Y(n_110)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

BUFx3_ASAP7_75t_L g282 ( 
.A(n_106),
.Y(n_282)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVx4_ASAP7_75t_L g157 ( 
.A(n_109),
.Y(n_157)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_110),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_110),
.B(n_152),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g285 ( 
.A(n_110),
.B(n_271),
.Y(n_285)
);

INVx4_ASAP7_75t_L g295 ( 
.A(n_111),
.Y(n_295)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_112),
.Y(n_129)
);

BUFx3_ASAP7_75t_L g133 ( 
.A(n_112),
.Y(n_133)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_115),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g148 ( 
.A(n_115),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g204 ( 
.A(n_115),
.Y(n_204)
);

BUFx5_ASAP7_75t_L g283 ( 
.A(n_115),
.Y(n_283)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_L g206 ( 
.A1(n_118),
.A2(n_207),
.B(n_214),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_SL g269 ( 
.A(n_118),
.B(n_119),
.Y(n_269)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

BUFx3_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

XNOR2xp5_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_149),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_124),
.B(n_149),
.Y(n_216)
);

AOI21xp5_ASAP7_75t_L g124 ( 
.A1(n_125),
.A2(n_134),
.B(n_141),
.Y(n_124)
);

AOI21xp5_ASAP7_75t_L g160 ( 
.A1(n_125),
.A2(n_161),
.B(n_164),
.Y(n_160)
);

INVx6_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

BUFx3_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_135),
.B(n_144),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_135),
.B(n_202),
.Y(n_240)
);

AOI21xp5_ASAP7_75t_L g265 ( 
.A1(n_135),
.A2(n_199),
.B(n_202),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_135),
.B(n_290),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_136),
.B(n_138),
.Y(n_135)
);

INVx3_ASAP7_75t_L g313 ( 
.A(n_136),
.Y(n_313)
);

BUFx5_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_137),
.Y(n_294)
);

INVx3_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

OR2x2_ASAP7_75t_L g239 ( 
.A(n_141),
.B(n_240),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_SL g317 ( 
.A(n_141),
.B(n_289),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_144),
.Y(n_141)
);

INVx3_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

AND2x2_ASAP7_75t_SL g149 ( 
.A(n_150),
.B(n_151),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_150),
.B(n_285),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_151),
.B(n_270),
.Y(n_297)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

INVx3_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

INVx5_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

INVx6_ASAP7_75t_L g279 ( 
.A(n_156),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_SL g158 ( 
.A(n_159),
.B(n_176),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_159),
.B(n_177),
.C(n_182),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_SL g159 ( 
.A(n_160),
.B(n_165),
.Y(n_159)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_160),
.B(n_165),
.Y(n_233)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

INVx3_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_163),
.Y(n_308)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_164),
.Y(n_205)
);

AOI32xp33_ASAP7_75t_L g165 ( 
.A1(n_166),
.A2(n_168),
.A3(n_170),
.B1(n_173),
.B2(n_174),
.Y(n_165)
);

INVx3_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

INVx8_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

INVx8_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

XOR2xp5_ASAP7_75t_L g176 ( 
.A(n_177),
.B(n_182),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_181),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_190),
.Y(n_182)
);

INVxp67_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

INVxp67_ASAP7_75t_SL g185 ( 
.A(n_186),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g329 ( 
.A(n_186),
.B(n_191),
.Y(n_329)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_190),
.B(n_236),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g192 ( 
.A(n_193),
.B(n_194),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g194 ( 
.A(n_195),
.B(n_215),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_206),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_205),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_197),
.B(n_288),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_201),
.Y(n_197)
);

INVx4_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

INVx4_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

INVxp67_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

INVx3_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_205),
.B(n_306),
.Y(n_305)
);

INVx1_ASAP7_75t_SL g208 ( 
.A(n_209),
.Y(n_208)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

INVx5_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_214),
.B(n_285),
.Y(n_327)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_216),
.B(n_217),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_L g217 ( 
.A1(n_218),
.A2(n_219),
.B1(n_221),
.B2(n_222),
.Y(n_217)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_218),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_219),
.Y(n_222)
);

INVxp67_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_L g225 ( 
.A1(n_226),
.A2(n_241),
.B(n_341),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_228),
.B(n_232),
.C(n_234),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_228),
.B(n_245),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_232),
.A2(n_233),
.B1(n_234),
.B2(n_246),
.Y(n_245)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_234),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_235),
.B(n_237),
.C(n_239),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g248 ( 
.A(n_235),
.B(n_249),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_237),
.A2(n_238),
.B1(n_239),
.B2(n_250),
.Y(n_249)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

CKINVDCx16_ASAP7_75t_R g250 ( 
.A(n_239),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_240),
.B(n_307),
.Y(n_315)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

OAI21xp5_ASAP7_75t_L g242 ( 
.A1(n_243),
.A2(n_272),
.B(n_340),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_SL g243 ( 
.A(n_244),
.B(n_247),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_244),
.B(n_247),
.Y(n_340)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_248),
.B(n_251),
.C(n_266),
.Y(n_247)
);

XOR2xp5_ASAP7_75t_L g335 ( 
.A(n_248),
.B(n_336),
.Y(n_335)
);

OAI22xp5_ASAP7_75t_SL g336 ( 
.A1(n_251),
.A2(n_266),
.B1(n_267),
.B2(n_337),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_251),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_252),
.B(n_265),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_L g330 ( 
.A1(n_252),
.A2(n_265),
.B1(n_331),
.B2(n_332),
.Y(n_330)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_252),
.Y(n_332)
);

BUFx3_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

INVx4_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

INVx8_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

INVx4_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_265),
.Y(n_331)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_268),
.B(n_270),
.Y(n_267)
);

INVxp67_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

AOI21xp5_ASAP7_75t_L g272 ( 
.A1(n_273),
.A2(n_334),
.B(n_339),
.Y(n_272)
);

OAI21xp5_ASAP7_75t_SL g273 ( 
.A1(n_274),
.A2(n_322),
.B(n_333),
.Y(n_273)
);

AOI21xp5_ASAP7_75t_L g274 ( 
.A1(n_275),
.A2(n_301),
.B(n_321),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_276),
.B(n_286),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_276),
.B(n_286),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_277),
.B(n_284),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_L g303 ( 
.A1(n_277),
.A2(n_278),
.B1(n_284),
.B2(n_304),
.Y(n_303)
);

CKINVDCx16_ASAP7_75t_R g277 ( 
.A(n_278),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_279),
.B(n_280),
.Y(n_278)
);

INVx4_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_284),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_L g286 ( 
.A(n_287),
.B(n_296),
.Y(n_286)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_287),
.Y(n_324)
);

INVxp67_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_290),
.B(n_308),
.Y(n_307)
);

BUFx2_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

INVx2_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_297),
.A2(n_298),
.B1(n_299),
.B2(n_300),
.Y(n_296)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_297),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_298),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_298),
.B(n_299),
.C(n_324),
.Y(n_323)
);

OAI21xp5_ASAP7_75t_SL g301 ( 
.A1(n_302),
.A2(n_309),
.B(n_320),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_SL g302 ( 
.A(n_303),
.B(n_305),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_303),
.B(n_305),
.Y(n_320)
);

INVxp67_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

AOI21xp5_ASAP7_75t_L g309 ( 
.A1(n_310),
.A2(n_316),
.B(n_319),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_311),
.B(n_315),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_312),
.B(n_314),
.Y(n_311)
);

INVx1_ASAP7_75t_SL g312 ( 
.A(n_313),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_SL g316 ( 
.A(n_317),
.B(n_318),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_317),
.B(n_318),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_323),
.B(n_325),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_323),
.B(n_325),
.Y(n_333)
);

XOR2xp5_ASAP7_75t_L g325 ( 
.A(n_326),
.B(n_330),
.Y(n_325)
);

XOR2xp5_ASAP7_75t_L g326 ( 
.A(n_327),
.B(n_328),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_327),
.B(n_328),
.C(n_330),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_SL g334 ( 
.A(n_335),
.B(n_338),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_335),
.B(n_338),
.Y(n_339)
);


endmodule