module fake_jpeg_31389_n_321 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_321);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_321;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx10_ASAP7_75t_L g18 ( 
.A(n_15),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_10),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_9),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_3),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_16),
.Y(n_28)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_17),
.Y(n_30)
);

BUFx12_ASAP7_75t_L g31 ( 
.A(n_17),
.Y(n_31)
);

INVxp67_ASAP7_75t_L g32 ( 
.A(n_5),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_8),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_1),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_8),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_15),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_0),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_1),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_10),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_7),
.Y(n_40)
);

INVx11_ASAP7_75t_L g41 ( 
.A(n_20),
.Y(n_41)
);

INVx5_ASAP7_75t_L g68 ( 
.A(n_41),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_20),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_42),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_36),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_43),
.Y(n_78)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_36),
.Y(n_44)
);

INVx6_ASAP7_75t_L g86 ( 
.A(n_44),
.Y(n_86)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_29),
.Y(n_45)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_45),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_40),
.Y(n_46)
);

INVx11_ASAP7_75t_L g76 ( 
.A(n_46),
.Y(n_76)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_22),
.Y(n_47)
);

INVx5_ASAP7_75t_L g73 ( 
.A(n_47),
.Y(n_73)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_22),
.Y(n_48)
);

INVx8_ASAP7_75t_L g55 ( 
.A(n_48),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_40),
.Y(n_49)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_49),
.Y(n_74)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_29),
.Y(n_50)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_50),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_28),
.Y(n_51)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_51),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_28),
.Y(n_52)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_52),
.Y(n_85)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_25),
.Y(n_53)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_53),
.Y(n_91)
);

CKINVDCx5p33_ASAP7_75t_R g54 ( 
.A(n_47),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_54),
.B(n_62),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_45),
.B(n_24),
.Y(n_56)
);

NAND3xp33_ASAP7_75t_L g117 ( 
.A(n_56),
.B(n_58),
.C(n_61),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_47),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_SL g119 ( 
.A(n_57),
.B(n_64),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_50),
.B(n_24),
.Y(n_58)
);

MAJIxp5_ASAP7_75t_L g60 ( 
.A(n_53),
.B(n_32),
.C(n_39),
.Y(n_60)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_60),
.B(n_72),
.Y(n_100)
);

A2O1A1Ixp33_ASAP7_75t_L g61 ( 
.A1(n_53),
.A2(n_32),
.B(n_33),
.C(n_21),
.Y(n_61)
);

BUFx12_ASAP7_75t_L g62 ( 
.A(n_48),
.Y(n_62)
);

OAI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_44),
.A2(n_39),
.B1(n_35),
.B2(n_33),
.Y(n_63)
);

OAI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_63),
.A2(n_18),
.B1(n_23),
.B2(n_19),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_48),
.B(n_30),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_51),
.B(n_30),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_66),
.B(n_67),
.Y(n_126)
);

CKINVDCx14_ASAP7_75t_R g67 ( 
.A(n_41),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_51),
.B(n_38),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_70),
.B(n_75),
.Y(n_124)
);

INVx13_ASAP7_75t_L g71 ( 
.A(n_41),
.Y(n_71)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_71),
.Y(n_129)
);

INVx1_ASAP7_75t_SL g72 ( 
.A(n_42),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_52),
.B(n_38),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_52),
.B(n_37),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_77),
.Y(n_101)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_44),
.Y(n_79)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_79),
.Y(n_110)
);

OAI22xp33_ASAP7_75t_L g80 ( 
.A1(n_42),
.A2(n_35),
.B1(n_21),
.B2(n_18),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_L g122 ( 
.A1(n_80),
.A2(n_84),
.B1(n_34),
.B2(n_19),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_42),
.A2(n_34),
.B1(n_19),
.B2(n_23),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_82),
.A2(n_92),
.B1(n_0),
.B2(n_2),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_43),
.B(n_37),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_83),
.B(n_88),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_49),
.A2(n_26),
.B1(n_27),
.B2(n_25),
.Y(n_84)
);

INVx6_ASAP7_75t_SL g87 ( 
.A(n_43),
.Y(n_87)
);

AND2x2_ASAP7_75t_L g103 ( 
.A(n_87),
.B(n_90),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_43),
.B(n_27),
.Y(n_88)
);

BUFx4f_ASAP7_75t_SL g89 ( 
.A(n_46),
.Y(n_89)
);

BUFx2_ASAP7_75t_L g115 ( 
.A(n_89),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_46),
.B(n_26),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_46),
.A2(n_34),
.B1(n_23),
.B2(n_19),
.Y(n_92)
);

OR2x2_ASAP7_75t_L g93 ( 
.A(n_49),
.B(n_31),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_93),
.Y(n_102)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_49),
.Y(n_94)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_94),
.Y(n_104)
);

AND2x2_ASAP7_75t_L g95 ( 
.A(n_53),
.B(n_18),
.Y(n_95)
);

AND2x2_ASAP7_75t_L g113 ( 
.A(n_95),
.B(n_18),
.Y(n_113)
);

BUFx4f_ASAP7_75t_SL g96 ( 
.A(n_47),
.Y(n_96)
);

INVx4_ASAP7_75t_L g114 ( 
.A(n_96),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_53),
.B(n_31),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_97),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_53),
.B(n_31),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_98),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_53),
.B(n_31),
.Y(n_99)
);

AOI21xp33_ASAP7_75t_SL g121 ( 
.A1(n_99),
.A2(n_34),
.B(n_23),
.Y(n_121)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_91),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g162 ( 
.A(n_105),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_106),
.A2(n_55),
.B1(n_68),
.B2(n_89),
.Y(n_156)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_74),
.Y(n_107)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_107),
.Y(n_141)
);

AND2x2_ASAP7_75t_SL g108 ( 
.A(n_59),
.B(n_0),
.Y(n_108)
);

FAx1_ASAP7_75t_SL g139 ( 
.A(n_108),
.B(n_92),
.CI(n_96),
.CON(n_139),
.SN(n_139)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_74),
.Y(n_109)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_109),
.Y(n_151)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_69),
.Y(n_111)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_111),
.Y(n_160)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_72),
.Y(n_112)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_112),
.Y(n_161)
);

AND2x2_ASAP7_75t_L g150 ( 
.A(n_113),
.B(n_132),
.Y(n_150)
);

NAND3xp33_ASAP7_75t_L g146 ( 
.A(n_121),
.B(n_16),
.C(n_3),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_L g136 ( 
.A1(n_122),
.A2(n_73),
.B1(n_86),
.B2(n_82),
.Y(n_136)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_81),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_125),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_65),
.Y(n_127)
);

INVx2_ASAP7_75t_SL g144 ( 
.A(n_127),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_87),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_128)
);

INVxp67_ASAP7_75t_L g148 ( 
.A(n_128),
.Y(n_148)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_81),
.Y(n_131)
);

CKINVDCx16_ASAP7_75t_R g158 ( 
.A(n_131),
.Y(n_158)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_76),
.Y(n_132)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_76),
.Y(n_133)
);

AND2x2_ASAP7_75t_L g154 ( 
.A(n_133),
.B(n_73),
.Y(n_154)
);

AND2x2_ASAP7_75t_SL g134 ( 
.A(n_124),
.B(n_61),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_134),
.B(n_137),
.C(n_113),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_119),
.B(n_54),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_135),
.B(n_142),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_136),
.A2(n_166),
.B1(n_115),
.B2(n_114),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_100),
.B(n_60),
.C(n_95),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_124),
.B(n_93),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_138),
.B(n_157),
.Y(n_168)
);

AND2x2_ASAP7_75t_L g172 ( 
.A(n_139),
.B(n_154),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_130),
.A2(n_86),
.B1(n_85),
.B2(n_78),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_140),
.A2(n_149),
.B1(n_111),
.B2(n_110),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_101),
.B(n_62),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_101),
.B(n_62),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_143),
.B(n_145),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_130),
.B(n_63),
.Y(n_145)
);

OAI21xp33_ASAP7_75t_L g185 ( 
.A1(n_146),
.A2(n_114),
.B(n_129),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_126),
.B(n_96),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_147),
.B(n_152),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_102),
.A2(n_78),
.B1(n_65),
.B2(n_80),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_118),
.B(n_55),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_SL g153 ( 
.A(n_120),
.B(n_2),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_SL g188 ( 
.A(n_153),
.B(n_11),
.Y(n_188)
);

INVxp33_ASAP7_75t_L g155 ( 
.A(n_116),
.Y(n_155)
);

INVx11_ASAP7_75t_L g186 ( 
.A(n_155),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_L g184 ( 
.A1(n_156),
.A2(n_159),
.B1(n_164),
.B2(n_115),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_117),
.B(n_89),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_103),
.B(n_5),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_163),
.B(n_11),
.Y(n_189)
);

OAI22x1_ASAP7_75t_SL g164 ( 
.A1(n_103),
.A2(n_71),
.B1(n_68),
.B2(n_8),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_108),
.B(n_6),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_165),
.B(n_167),
.Y(n_171)
);

AOI22xp33_ASAP7_75t_L g166 ( 
.A1(n_112),
.A2(n_7),
.B1(n_9),
.B2(n_11),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_108),
.B(n_9),
.Y(n_167)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_162),
.Y(n_170)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_170),
.Y(n_209)
);

AOI21xp5_ASAP7_75t_L g173 ( 
.A1(n_164),
.A2(n_100),
.B(n_103),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_SL g216 ( 
.A1(n_173),
.A2(n_175),
.B(n_180),
.Y(n_216)
);

CKINVDCx16_ASAP7_75t_R g174 ( 
.A(n_154),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_174),
.B(n_176),
.Y(n_202)
);

AOI21xp5_ASAP7_75t_SL g175 ( 
.A1(n_157),
.A2(n_100),
.B(n_110),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_177),
.A2(n_195),
.B1(n_196),
.B2(n_200),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g213 ( 
.A(n_179),
.B(n_201),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_SL g180 ( 
.A1(n_137),
.A2(n_113),
.B(n_105),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_138),
.B(n_104),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_181),
.B(n_191),
.Y(n_215)
);

INVxp67_ASAP7_75t_L g182 ( 
.A(n_154),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_182),
.B(n_186),
.Y(n_222)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_160),
.Y(n_183)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_183),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_SL g218 ( 
.A1(n_184),
.A2(n_159),
.B(n_144),
.Y(n_218)
);

NAND3xp33_ASAP7_75t_L g225 ( 
.A(n_185),
.B(n_188),
.C(n_189),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_L g190 ( 
.A1(n_134),
.A2(n_127),
.B1(n_133),
.B2(n_132),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_190),
.B(n_193),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_134),
.B(n_104),
.Y(n_191)
);

O2A1O1Ixp33_ASAP7_75t_L g192 ( 
.A1(n_148),
.A2(n_131),
.B(n_123),
.C(n_107),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_L g224 ( 
.A1(n_192),
.A2(n_151),
.B(n_144),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_165),
.B(n_129),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_SL g194 ( 
.A(n_167),
.B(n_12),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_SL g204 ( 
.A(n_194),
.B(n_153),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_156),
.A2(n_109),
.B1(n_13),
.B2(n_14),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_148),
.A2(n_12),
.B1(n_13),
.B2(n_14),
.Y(n_196)
);

BUFx6f_ASAP7_75t_L g197 ( 
.A(n_162),
.Y(n_197)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_197),
.Y(n_214)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_160),
.Y(n_198)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_198),
.Y(n_210)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_161),
.Y(n_199)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_199),
.Y(n_211)
);

OAI22xp33_ASAP7_75t_SL g200 ( 
.A1(n_139),
.A2(n_13),
.B1(n_15),
.B2(n_149),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_150),
.B(n_139),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_179),
.B(n_150),
.C(n_158),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_203),
.B(n_206),
.C(n_220),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_204),
.B(n_205),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_187),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_180),
.B(n_150),
.C(n_140),
.Y(n_206)
);

CKINVDCx16_ASAP7_75t_R g207 ( 
.A(n_199),
.Y(n_207)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_207),
.Y(n_243)
);

OR2x4_ASAP7_75t_L g212 ( 
.A(n_172),
.B(n_161),
.Y(n_212)
);

AO21x1_ASAP7_75t_L g234 ( 
.A1(n_212),
.A2(n_218),
.B(n_224),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_SL g219 ( 
.A(n_169),
.B(n_141),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_SL g242 ( 
.A(n_219),
.B(n_226),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_201),
.B(n_141),
.Y(n_220)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_168),
.B(n_181),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_221),
.B(n_171),
.C(n_193),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_222),
.B(n_223),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_177),
.A2(n_144),
.B1(n_162),
.B2(n_151),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_186),
.B(n_178),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_213),
.B(n_168),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_SL g251 ( 
.A(n_228),
.B(n_229),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_213),
.B(n_172),
.Y(n_229)
);

OAI21xp5_ASAP7_75t_L g231 ( 
.A1(n_202),
.A2(n_172),
.B(n_173),
.Y(n_231)
);

OAI21xp5_ASAP7_75t_L g260 ( 
.A1(n_231),
.A2(n_225),
.B(n_236),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_215),
.B(n_191),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_232),
.B(n_236),
.Y(n_263)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_210),
.Y(n_233)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_233),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_215),
.B(n_198),
.Y(n_236)
);

XOR2xp5_ASAP7_75t_L g257 ( 
.A(n_238),
.B(n_239),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_221),
.B(n_175),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_206),
.A2(n_182),
.B1(n_176),
.B2(n_195),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_240),
.A2(n_246),
.B1(n_216),
.B2(n_196),
.Y(n_266)
);

CKINVDCx16_ASAP7_75t_R g241 ( 
.A(n_210),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_SL g256 ( 
.A(n_241),
.B(n_245),
.Y(n_256)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_211),
.Y(n_244)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_244),
.Y(n_259)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_211),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_227),
.A2(n_183),
.B1(n_171),
.B2(n_192),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_208),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_247),
.B(n_209),
.Y(n_264)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_223),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_248),
.B(n_227),
.Y(n_249)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_249),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_235),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_250),
.B(n_252),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_SL g252 ( 
.A(n_242),
.B(n_188),
.Y(n_252)
);

BUFx3_ASAP7_75t_L g253 ( 
.A(n_243),
.Y(n_253)
);

INVx1_ASAP7_75t_SL g277 ( 
.A(n_253),
.Y(n_277)
);

AND2x2_ASAP7_75t_L g254 ( 
.A(n_230),
.B(n_224),
.Y(n_254)
);

INVxp67_ASAP7_75t_L g271 ( 
.A(n_254),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_L g258 ( 
.A1(n_230),
.A2(n_217),
.B1(n_218),
.B2(n_212),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_L g272 ( 
.A1(n_258),
.A2(n_266),
.B1(n_265),
.B2(n_231),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_260),
.B(n_265),
.Y(n_269)
);

AOI21xp5_ASAP7_75t_SL g261 ( 
.A1(n_234),
.A2(n_216),
.B(n_220),
.Y(n_261)
);

INVxp67_ASAP7_75t_L g274 ( 
.A(n_261),
.Y(n_274)
);

INVxp67_ASAP7_75t_L g262 ( 
.A(n_247),
.Y(n_262)
);

CKINVDCx16_ASAP7_75t_R g268 ( 
.A(n_262),
.Y(n_268)
);

HB1xp67_ASAP7_75t_L g281 ( 
.A(n_264),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_232),
.B(n_217),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_257),
.B(n_237),
.C(n_251),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_270),
.B(n_278),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_SL g287 ( 
.A(n_272),
.B(n_275),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_257),
.B(n_237),
.C(n_228),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_273),
.B(n_240),
.C(n_263),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_SL g275 ( 
.A(n_251),
.B(n_229),
.Y(n_275)
);

XOR2xp5_ASAP7_75t_L g276 ( 
.A(n_266),
.B(n_239),
.Y(n_276)
);

XOR2xp5_ASAP7_75t_L g282 ( 
.A(n_276),
.B(n_254),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_260),
.B(n_203),
.C(n_238),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_261),
.B(n_234),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g286 ( 
.A(n_280),
.B(n_246),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g298 ( 
.A(n_282),
.B(n_285),
.Y(n_298)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_267),
.Y(n_283)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_283),
.Y(n_300)
);

XOR2xp5_ASAP7_75t_L g285 ( 
.A(n_273),
.B(n_254),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g299 ( 
.A(n_286),
.B(n_289),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_SL g288 ( 
.A(n_279),
.B(n_256),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_288),
.B(n_290),
.Y(n_301)
);

XOR2xp5_ASAP7_75t_L g289 ( 
.A(n_276),
.B(n_263),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_L g291 ( 
.A1(n_274),
.A2(n_255),
.B1(n_262),
.B2(n_259),
.Y(n_291)
);

OR2x2_ASAP7_75t_L g294 ( 
.A(n_291),
.B(n_292),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_269),
.B(n_253),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_282),
.B(n_268),
.Y(n_293)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_293),
.Y(n_304)
);

AOI322xp5_ASAP7_75t_SL g295 ( 
.A1(n_287),
.A2(n_274),
.A3(n_271),
.B1(n_275),
.B2(n_285),
.C1(n_284),
.C2(n_289),
.Y(n_295)
);

OAI21xp5_ASAP7_75t_SL g303 ( 
.A1(n_295),
.A2(n_277),
.B(n_264),
.Y(n_303)
);

OAI21xp5_ASAP7_75t_L g296 ( 
.A1(n_287),
.A2(n_271),
.B(n_281),
.Y(n_296)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_296),
.Y(n_305)
);

CKINVDCx16_ASAP7_75t_R g297 ( 
.A(n_283),
.Y(n_297)
);

INVx6_ASAP7_75t_L g308 ( 
.A(n_297),
.Y(n_308)
);

OR2x2_ASAP7_75t_L g302 ( 
.A(n_294),
.B(n_300),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_302),
.B(n_303),
.Y(n_309)
);

NAND2xp33_ASAP7_75t_SL g306 ( 
.A(n_295),
.B(n_277),
.Y(n_306)
);

HB1xp67_ASAP7_75t_L g312 ( 
.A(n_306),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_L g307 ( 
.A(n_299),
.B(n_233),
.Y(n_307)
);

XOR2xp5_ASAP7_75t_L g311 ( 
.A(n_307),
.B(n_194),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_L g310 ( 
.A1(n_305),
.A2(n_293),
.B1(n_298),
.B2(n_301),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_L g314 ( 
.A1(n_310),
.A2(n_302),
.B1(n_304),
.B2(n_306),
.Y(n_314)
);

XOR2xp5_ASAP7_75t_L g315 ( 
.A(n_311),
.B(n_308),
.Y(n_315)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_309),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_313),
.B(n_314),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_315),
.B(n_312),
.Y(n_316)
);

XOR2xp5_ASAP7_75t_L g318 ( 
.A(n_316),
.B(n_315),
.Y(n_318)
);

AOI21xp5_ASAP7_75t_SL g319 ( 
.A1(n_318),
.A2(n_317),
.B(n_311),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_319),
.B(n_308),
.C(n_214),
.Y(n_320)
);

XOR2xp5_ASAP7_75t_L g321 ( 
.A(n_320),
.B(n_214),
.Y(n_321)
);


endmodule