module fake_jpeg_22967_n_255 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_255);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_255;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_182;
wire n_19;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_122;
wire n_75;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_93;
wire n_54;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_213;
wire n_153;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx8_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_16),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

INVx11_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_13),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

BUFx4f_ASAP7_75t_SL g27 ( 
.A(n_9),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_8),
.Y(n_30)
);

INVx13_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_13),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

HB1xp67_ASAP7_75t_L g34 ( 
.A(n_8),
.Y(n_34)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_21),
.Y(n_35)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_35),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_27),
.Y(n_36)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_36),
.Y(n_53)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_24),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_37),
.B(n_41),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_31),
.B(n_0),
.Y(n_38)
);

AND2x2_ASAP7_75t_SL g62 ( 
.A(n_38),
.B(n_42),
.Y(n_62)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_21),
.Y(n_39)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_27),
.Y(n_40)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_40),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_25),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_25),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_31),
.B(n_0),
.Y(n_43)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_43),
.Y(n_50)
);

INVx6_ASAP7_75t_SL g44 ( 
.A(n_27),
.Y(n_44)
);

INVxp67_ASAP7_75t_L g56 ( 
.A(n_44),
.Y(n_56)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_39),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_45),
.B(n_52),
.Y(n_95)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_40),
.Y(n_46)
);

INVx5_ASAP7_75t_L g77 ( 
.A(n_46),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_L g47 ( 
.A1(n_35),
.A2(n_17),
.B1(n_34),
.B2(n_24),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_47),
.A2(n_58),
.B1(n_29),
.B2(n_23),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_39),
.A2(n_17),
.B1(n_24),
.B2(n_31),
.Y(n_48)
);

AOI21xp5_ASAP7_75t_L g69 ( 
.A1(n_48),
.A2(n_61),
.B(n_38),
.Y(n_69)
);

OA22x2_ASAP7_75t_L g51 ( 
.A1(n_40),
.A2(n_31),
.B1(n_27),
.B2(n_34),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_51),
.A2(n_55),
.B1(n_37),
.B2(n_35),
.Y(n_67)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_43),
.Y(n_52)
);

OA22x2_ASAP7_75t_L g55 ( 
.A1(n_40),
.A2(n_27),
.B1(n_19),
.B2(n_20),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_L g58 ( 
.A1(n_35),
.A2(n_17),
.B1(n_26),
.B2(n_33),
.Y(n_58)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_39),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_60),
.B(n_63),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_39),
.A2(n_17),
.B1(n_26),
.B2(n_29),
.Y(n_61)
);

INVxp67_ASAP7_75t_L g63 ( 
.A(n_40),
.Y(n_63)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_37),
.Y(n_64)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_64),
.Y(n_75)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_37),
.Y(n_65)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_65),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_62),
.B(n_38),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_66),
.B(n_73),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_67),
.A2(n_69),
.B1(n_90),
.B2(n_94),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g68 ( 
.A(n_46),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_68),
.B(n_70),
.Y(n_100)
);

OR2x2_ASAP7_75t_L g70 ( 
.A(n_49),
.B(n_42),
.Y(n_70)
);

AO22x1_ASAP7_75t_L g71 ( 
.A1(n_51),
.A2(n_44),
.B1(n_35),
.B2(n_36),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_71),
.A2(n_80),
.B1(n_88),
.B2(n_93),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_50),
.A2(n_26),
.B1(n_18),
.B2(n_23),
.Y(n_72)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_72),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_62),
.B(n_43),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_74),
.B(n_86),
.Y(n_101)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_64),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_78),
.B(n_79),
.Y(n_111)
);

CKINVDCx16_ASAP7_75t_R g79 ( 
.A(n_51),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_59),
.A2(n_19),
.B1(n_20),
.B2(n_41),
.Y(n_80)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_62),
.B(n_44),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_81),
.B(n_44),
.C(n_36),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_59),
.Y(n_82)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_82),
.Y(n_107)
);

OR2x2_ASAP7_75t_L g83 ( 
.A(n_56),
.B(n_42),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_83),
.B(n_84),
.Y(n_122)
);

OR2x2_ASAP7_75t_L g84 ( 
.A(n_56),
.B(n_41),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_51),
.B(n_36),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_85),
.B(n_89),
.Y(n_105)
);

CKINVDCx16_ASAP7_75t_R g86 ( 
.A(n_65),
.Y(n_86)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_53),
.Y(n_87)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_87),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_45),
.A2(n_19),
.B1(n_20),
.B2(n_18),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_63),
.B(n_36),
.Y(n_89)
);

CKINVDCx14_ASAP7_75t_R g90 ( 
.A(n_57),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_54),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_91),
.Y(n_119)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_53),
.Y(n_92)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_92),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_55),
.A2(n_29),
.B1(n_23),
.B2(n_18),
.Y(n_93)
);

OAI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_55),
.A2(n_33),
.B1(n_22),
.B2(n_30),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_L g96 ( 
.A1(n_55),
.A2(n_32),
.B1(n_30),
.B2(n_33),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_96),
.A2(n_32),
.B1(n_22),
.B2(n_28),
.Y(n_114)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_46),
.Y(n_97)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_97),
.Y(n_109)
);

XNOR2xp5_ASAP7_75t_L g142 ( 
.A(n_99),
.B(n_113),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_66),
.B(n_28),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_106),
.B(n_108),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_73),
.B(n_81),
.Y(n_108)
);

XOR2xp5_ASAP7_75t_L g113 ( 
.A(n_69),
.B(n_28),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_114),
.A2(n_116),
.B1(n_118),
.B2(n_88),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_81),
.B(n_28),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_115),
.B(n_82),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_85),
.A2(n_21),
.B1(n_16),
.B2(n_2),
.Y(n_116)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_95),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_117),
.B(n_120),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_71),
.A2(n_67),
.B1(n_74),
.B2(n_93),
.Y(n_118)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_98),
.Y(n_120)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_89),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_123),
.B(n_124),
.Y(n_132)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_80),
.Y(n_124)
);

AND2x6_ASAP7_75t_L g125 ( 
.A(n_113),
.B(n_71),
.Y(n_125)
);

XOR2xp5_ASAP7_75t_L g169 ( 
.A(n_125),
.B(n_141),
.Y(n_169)
);

INVx13_ASAP7_75t_L g126 ( 
.A(n_110),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_126),
.B(n_131),
.Y(n_153)
);

NAND3xp33_ASAP7_75t_SL g128 ( 
.A(n_108),
.B(n_84),
.C(n_83),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g157 ( 
.A(n_128),
.B(n_134),
.Y(n_157)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_107),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_129),
.B(n_130),
.Y(n_176)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_107),
.Y(n_130)
);

CKINVDCx14_ASAP7_75t_R g131 ( 
.A(n_100),
.Y(n_131)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_105),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_133),
.B(n_139),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_SL g134 ( 
.A(n_122),
.B(n_70),
.Y(n_134)
);

CKINVDCx16_ASAP7_75t_R g136 ( 
.A(n_105),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_136),
.B(n_137),
.Y(n_162)
);

INVxp67_ASAP7_75t_L g138 ( 
.A(n_99),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_138),
.B(n_147),
.Y(n_175)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_116),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_SL g171 ( 
.A1(n_140),
.A2(n_145),
.B(n_148),
.Y(n_171)
);

AND2x6_ASAP7_75t_L g141 ( 
.A(n_115),
.B(n_0),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_102),
.A2(n_78),
.B1(n_75),
.B2(n_76),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_143),
.A2(n_149),
.B1(n_150),
.B2(n_103),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_119),
.B(n_75),
.Y(n_144)
);

CKINVDCx16_ASAP7_75t_R g155 ( 
.A(n_144),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_L g145 ( 
.A1(n_103),
.A2(n_76),
.B(n_91),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_110),
.B(n_97),
.Y(n_146)
);

CKINVDCx16_ASAP7_75t_R g165 ( 
.A(n_146),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_109),
.B(n_87),
.Y(n_147)
);

OAI21xp33_ASAP7_75t_L g148 ( 
.A1(n_104),
.A2(n_1),
.B(n_2),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_102),
.A2(n_92),
.B1(n_77),
.B2(n_68),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_124),
.A2(n_77),
.B1(n_21),
.B2(n_3),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_109),
.B(n_1),
.Y(n_151)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_151),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_132),
.B(n_123),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_154),
.B(n_164),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_156),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_136),
.B(n_104),
.Y(n_158)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_158),
.Y(n_193)
);

O2A1O1Ixp33_ASAP7_75t_SL g159 ( 
.A1(n_143),
.A2(n_101),
.B(n_118),
.C(n_112),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_SL g179 ( 
.A1(n_159),
.A2(n_170),
.B(n_174),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_133),
.B(n_106),
.Y(n_160)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_160),
.Y(n_196)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_127),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_163),
.B(n_168),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_134),
.B(n_112),
.Y(n_164)
);

HB1xp67_ASAP7_75t_L g166 ( 
.A(n_126),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_166),
.B(n_172),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_135),
.B(n_120),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_167),
.B(n_173),
.Y(n_194)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_127),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_139),
.A2(n_111),
.B1(n_117),
.B2(n_114),
.Y(n_170)
);

HB1xp67_ASAP7_75t_L g172 ( 
.A(n_129),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_135),
.B(n_121),
.Y(n_173)
);

NAND2xp33_ASAP7_75t_L g174 ( 
.A(n_125),
.B(n_121),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_175),
.B(n_142),
.C(n_138),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_177),
.B(n_184),
.C(n_187),
.Y(n_200)
);

AND2x4_ASAP7_75t_L g180 ( 
.A(n_174),
.B(n_145),
.Y(n_180)
);

AND2x2_ASAP7_75t_L g199 ( 
.A(n_180),
.B(n_173),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_SL g182 ( 
.A(n_157),
.B(n_137),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_182),
.B(n_183),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_176),
.Y(n_183)
);

XOR2xp5_ASAP7_75t_L g184 ( 
.A(n_169),
.B(n_142),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_SL g185 ( 
.A(n_157),
.B(n_140),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_185),
.B(n_189),
.Y(n_211)
);

AOI21xp5_ASAP7_75t_L g186 ( 
.A1(n_162),
.A2(n_149),
.B(n_130),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_L g203 ( 
.A1(n_186),
.A2(n_191),
.B1(n_171),
.B2(n_170),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_158),
.B(n_141),
.C(n_150),
.Y(n_187)
);

OR2x2_ASAP7_75t_L g189 ( 
.A(n_154),
.B(n_2),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_155),
.B(n_12),
.Y(n_190)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_190),
.Y(n_202)
);

OR2x2_ASAP7_75t_L g192 ( 
.A(n_164),
.B(n_12),
.Y(n_192)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_192),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_169),
.B(n_3),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_195),
.B(n_171),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_180),
.A2(n_159),
.B1(n_156),
.B2(n_152),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g214 ( 
.A1(n_197),
.A2(n_198),
.B1(n_204),
.B2(n_209),
.Y(n_214)
);

AOI22xp33_ASAP7_75t_L g198 ( 
.A1(n_186),
.A2(n_165),
.B1(n_168),
.B2(n_163),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_199),
.A2(n_207),
.B1(n_188),
.B2(n_194),
.Y(n_217)
);

BUFx2_ASAP7_75t_L g201 ( 
.A(n_180),
.Y(n_201)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_201),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_203),
.B(n_210),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_180),
.A2(n_152),
.B1(n_159),
.B2(n_167),
.Y(n_204)
);

XOR2xp5_ASAP7_75t_L g219 ( 
.A(n_206),
.B(n_184),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_188),
.A2(n_193),
.B1(n_179),
.B2(n_196),
.Y(n_207)
);

OA22x2_ASAP7_75t_L g209 ( 
.A1(n_192),
.A2(n_165),
.B1(n_155),
.B2(n_176),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_181),
.Y(n_210)
);

BUFx2_ASAP7_75t_L g212 ( 
.A(n_178),
.Y(n_212)
);

HB1xp67_ASAP7_75t_L g222 ( 
.A(n_212),
.Y(n_222)
);

INVx1_ASAP7_75t_SL g213 ( 
.A(n_212),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_213),
.B(n_220),
.Y(n_226)
);

AOI21xp5_ASAP7_75t_SL g216 ( 
.A1(n_199),
.A2(n_179),
.B(n_205),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_L g231 ( 
.A1(n_216),
.A2(n_218),
.B(n_207),
.Y(n_231)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_217),
.B(n_219),
.Y(n_230)
);

AOI21xp5_ASAP7_75t_L g218 ( 
.A1(n_201),
.A2(n_187),
.B(n_194),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_200),
.B(n_177),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_200),
.B(n_195),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_221),
.B(n_206),
.Y(n_227)
);

NAND3xp33_ASAP7_75t_L g224 ( 
.A(n_208),
.B(n_193),
.C(n_196),
.Y(n_224)
);

AND2x2_ASAP7_75t_L g233 ( 
.A(n_224),
.B(n_209),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_SL g225 ( 
.A(n_215),
.B(n_202),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_225),
.B(n_227),
.Y(n_241)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_222),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_228),
.B(n_232),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_223),
.A2(n_204),
.B1(n_199),
.B2(n_197),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_229),
.A2(n_216),
.B1(n_191),
.B2(n_224),
.Y(n_235)
);

OAI21xp5_ASAP7_75t_L g238 ( 
.A1(n_231),
.A2(n_161),
.B(n_220),
.Y(n_238)
);

CKINVDCx16_ASAP7_75t_R g232 ( 
.A(n_214),
.Y(n_232)
);

AOI322xp5_ASAP7_75t_L g236 ( 
.A1(n_233),
.A2(n_234),
.A3(n_211),
.B1(n_209),
.B2(n_160),
.C1(n_189),
.C2(n_153),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_213),
.B(n_209),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_SL g244 ( 
.A(n_235),
.B(n_238),
.Y(n_244)
);

A2O1A1O1Ixp25_ASAP7_75t_L g242 ( 
.A1(n_236),
.A2(n_240),
.B(n_238),
.C(n_235),
.D(n_237),
.Y(n_242)
);

AOI322xp5_ASAP7_75t_L g239 ( 
.A1(n_231),
.A2(n_161),
.A3(n_5),
.B1(n_6),
.B2(n_7),
.C1(n_4),
.C2(n_9),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_SL g245 ( 
.A(n_239),
.B(n_240),
.Y(n_245)
);

NOR2x1_ASAP7_75t_L g240 ( 
.A(n_233),
.B(n_4),
.Y(n_240)
);

AOI21xp5_ASAP7_75t_L g250 ( 
.A1(n_242),
.A2(n_246),
.B(n_5),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_SL g243 ( 
.A(n_241),
.B(n_226),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_243),
.B(n_245),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_241),
.B(n_229),
.Y(n_246)
);

OAI21xp5_ASAP7_75t_L g248 ( 
.A1(n_244),
.A2(n_230),
.B(n_228),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_248),
.B(n_249),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_243),
.B(n_230),
.Y(n_249)
);

NAND3xp33_ASAP7_75t_L g251 ( 
.A(n_250),
.B(n_6),
.C(n_7),
.Y(n_251)
);

OAI221xp5_ASAP7_75t_L g254 ( 
.A1(n_251),
.A2(n_247),
.B1(n_9),
.B2(n_10),
.C(n_12),
.Y(n_254)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_252),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_253),
.B(n_254),
.Y(n_255)
);


endmodule