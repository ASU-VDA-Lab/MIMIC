module fake_jpeg_9717_n_315 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_315);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_315;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx3_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_4),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_1),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_11),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

INVx8_ASAP7_75t_SL g25 ( 
.A(n_14),
.Y(n_25)
);

BUFx12_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_13),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_14),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_12),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_26),
.B(n_15),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_34),
.B(n_39),
.Y(n_49)
);

INVx11_ASAP7_75t_L g35 ( 
.A(n_24),
.Y(n_35)
);

BUFx2_ASAP7_75t_L g53 ( 
.A(n_35),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g36 ( 
.A(n_24),
.B(n_0),
.Y(n_36)
);

AND2x2_ASAP7_75t_L g54 ( 
.A(n_36),
.B(n_27),
.Y(n_54)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_27),
.Y(n_37)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_18),
.Y(n_38)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_38),
.Y(n_51)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_27),
.Y(n_39)
);

INVx5_ASAP7_75t_L g40 ( 
.A(n_25),
.Y(n_40)
);

INVx5_ASAP7_75t_L g62 ( 
.A(n_40),
.Y(n_62)
);

OR2x2_ASAP7_75t_L g41 ( 
.A(n_26),
.B(n_0),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_SL g47 ( 
.A(n_41),
.B(n_19),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_18),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_42),
.Y(n_57)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_22),
.Y(n_43)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_43),
.Y(n_64)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_40),
.Y(n_44)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_44),
.Y(n_74)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_40),
.Y(n_45)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_45),
.Y(n_83)
);

OAI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_43),
.A2(n_16),
.B1(n_25),
.B2(n_32),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_46),
.A2(n_62),
.B1(n_35),
.B2(n_37),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_47),
.B(n_55),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g48 ( 
.A(n_41),
.B(n_21),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_SL g79 ( 
.A(n_48),
.B(n_58),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_41),
.B(n_21),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_52),
.B(n_59),
.Y(n_78)
);

AND2x2_ASAP7_75t_L g73 ( 
.A(n_54),
.B(n_36),
.Y(n_73)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_34),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_34),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_56),
.B(n_65),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_41),
.B(n_19),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_41),
.B(n_21),
.Y(n_59)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_40),
.Y(n_60)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_60),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_36),
.A2(n_16),
.B1(n_20),
.B2(n_33),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_61),
.A2(n_36),
.B1(n_20),
.B2(n_17),
.Y(n_75)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_40),
.Y(n_63)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_63),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_41),
.B(n_19),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_34),
.B(n_33),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_66),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_43),
.A2(n_16),
.B1(n_32),
.B2(n_33),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_67),
.A2(n_43),
.B1(n_39),
.B2(n_37),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_37),
.B(n_29),
.Y(n_68)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_68),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_L g120 ( 
.A1(n_69),
.A2(n_51),
.B1(n_30),
.B2(n_22),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_55),
.A2(n_32),
.B1(n_43),
.B2(n_37),
.Y(n_70)
);

CKINVDCx16_ASAP7_75t_R g111 ( 
.A(n_70),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_73),
.B(n_54),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_75),
.B(n_61),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g76 ( 
.A1(n_56),
.A2(n_35),
.B1(n_39),
.B2(n_37),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_76),
.A2(n_77),
.B1(n_80),
.B2(n_84),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_62),
.A2(n_39),
.B1(n_23),
.B2(n_29),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_L g81 ( 
.A(n_49),
.B(n_38),
.C(n_42),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_81),
.B(n_91),
.C(n_18),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_53),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_82),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_49),
.A2(n_35),
.B1(n_39),
.B2(n_23),
.Y(n_84)
);

BUFx3_ASAP7_75t_L g85 ( 
.A(n_57),
.Y(n_85)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_85),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_L g86 ( 
.A1(n_52),
.A2(n_35),
.B1(n_39),
.B2(n_30),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_86),
.A2(n_93),
.B1(n_50),
.B2(n_51),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_53),
.Y(n_87)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_87),
.Y(n_98)
);

AND2x2_ASAP7_75t_L g91 ( 
.A(n_48),
.B(n_0),
.Y(n_91)
);

A2O1A1Ixp33_ASAP7_75t_L g92 ( 
.A1(n_58),
.A2(n_20),
.B(n_17),
.C(n_28),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g102 ( 
.A(n_92),
.B(n_47),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_L g93 ( 
.A1(n_59),
.A2(n_22),
.B1(n_30),
.B2(n_31),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_73),
.A2(n_60),
.B1(n_45),
.B2(n_63),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_95),
.A2(n_97),
.B1(n_92),
.B2(n_83),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_73),
.A2(n_44),
.B1(n_54),
.B2(n_64),
.Y(n_97)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_76),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_100),
.B(n_110),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_101),
.B(n_121),
.C(n_90),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_102),
.B(n_104),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_84),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_103),
.B(n_105),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_86),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_88),
.B(n_65),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_SL g130 ( 
.A(n_106),
.B(n_107),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_SL g107 ( 
.A(n_88),
.B(n_66),
.Y(n_107)
);

OAI22xp33_ASAP7_75t_L g108 ( 
.A1(n_77),
.A2(n_50),
.B1(n_64),
.B2(n_51),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_108),
.A2(n_120),
.B1(n_71),
.B2(n_72),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_78),
.B(n_38),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_109),
.B(n_118),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_92),
.Y(n_110)
);

AND2x2_ASAP7_75t_L g127 ( 
.A(n_112),
.B(n_81),
.Y(n_127)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_94),
.Y(n_113)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_113),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_114),
.A2(n_72),
.B1(n_71),
.B2(n_83),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_89),
.B(n_94),
.Y(n_115)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_115),
.Y(n_134)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_93),
.Y(n_117)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_117),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_90),
.B(n_15),
.Y(n_118)
);

OA21x2_ASAP7_75t_L g119 ( 
.A1(n_74),
.A2(n_50),
.B(n_42),
.Y(n_119)
);

AOI21xp5_ASAP7_75t_L g137 ( 
.A1(n_119),
.A2(n_74),
.B(n_57),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_78),
.B(n_73),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_122),
.A2(n_143),
.B1(n_120),
.B2(n_95),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_123),
.B(n_127),
.C(n_42),
.Y(n_173)
);

OAI22xp33_ASAP7_75t_SL g161 ( 
.A1(n_124),
.A2(n_145),
.B1(n_146),
.B2(n_98),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_119),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_125),
.B(n_126),
.Y(n_148)
);

INVxp33_ASAP7_75t_L g126 ( 
.A(n_98),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_119),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_128),
.B(n_144),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_133),
.A2(n_99),
.B1(n_114),
.B2(n_117),
.Y(n_155)
);

INVx4_ASAP7_75t_L g135 ( 
.A(n_96),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_135),
.B(n_136),
.Y(n_150)
);

INVx3_ASAP7_75t_L g136 ( 
.A(n_116),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_SL g168 ( 
.A1(n_137),
.A2(n_138),
.B(n_139),
.Y(n_168)
);

AOI21xp5_ASAP7_75t_L g138 ( 
.A1(n_111),
.A2(n_91),
.B(n_79),
.Y(n_138)
);

AOI21xp5_ASAP7_75t_L g139 ( 
.A1(n_111),
.A2(n_91),
.B(n_79),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_100),
.A2(n_75),
.B1(n_89),
.B2(n_91),
.Y(n_143)
);

INVx8_ASAP7_75t_L g144 ( 
.A(n_116),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_SL g145 ( 
.A1(n_105),
.A2(n_103),
.B1(n_110),
.B2(n_96),
.Y(n_145)
);

INVx4_ASAP7_75t_SL g146 ( 
.A(n_116),
.Y(n_146)
);

AO221x1_ASAP7_75t_L g147 ( 
.A1(n_119),
.A2(n_42),
.B1(n_38),
.B2(n_87),
.C(n_82),
.Y(n_147)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_147),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_130),
.B(n_102),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_149),
.B(n_151),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_130),
.B(n_106),
.Y(n_151)
);

CKINVDCx16_ASAP7_75t_R g152 ( 
.A(n_132),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_152),
.B(n_153),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_140),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_SL g154 ( 
.A(n_134),
.B(n_131),
.Y(n_154)
);

CKINVDCx14_ASAP7_75t_R g188 ( 
.A(n_154),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_155),
.A2(n_158),
.B1(n_169),
.B2(n_171),
.Y(n_176)
);

NAND2x1p5_ASAP7_75t_L g156 ( 
.A(n_125),
.B(n_101),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_SL g194 ( 
.A1(n_156),
.A2(n_172),
.B(n_38),
.Y(n_194)
);

AND2x6_ASAP7_75t_L g157 ( 
.A(n_127),
.B(n_112),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_157),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_128),
.A2(n_99),
.B1(n_104),
.B2(n_113),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_140),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_160),
.B(n_170),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g199 ( 
.A1(n_161),
.A2(n_146),
.B1(n_144),
.B2(n_136),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_129),
.B(n_109),
.Y(n_162)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_162),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_134),
.B(n_115),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_164),
.B(n_167),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_129),
.B(n_121),
.Y(n_165)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_165),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_166),
.A2(n_144),
.B1(n_57),
.B2(n_53),
.Y(n_200)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_122),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_133),
.A2(n_107),
.B1(n_97),
.B2(n_118),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_SL g170 ( 
.A(n_131),
.B(n_12),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_137),
.A2(n_87),
.B1(n_82),
.B2(n_85),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_147),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_173),
.B(n_123),
.C(n_127),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_141),
.B(n_42),
.Y(n_174)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_174),
.Y(n_180)
);

CKINVDCx16_ASAP7_75t_R g178 ( 
.A(n_150),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_178),
.B(n_192),
.Y(n_203)
);

AOI21xp5_ASAP7_75t_L g181 ( 
.A1(n_168),
.A2(n_160),
.B(n_153),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_L g207 ( 
.A1(n_181),
.A2(n_199),
.B1(n_200),
.B2(n_172),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_158),
.A2(n_143),
.B1(n_142),
.B2(n_124),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_182),
.A2(n_167),
.B1(n_152),
.B2(n_159),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_183),
.B(n_184),
.C(n_186),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_173),
.B(n_139),
.C(n_138),
.Y(n_184)
);

INVxp67_ASAP7_75t_L g185 ( 
.A(n_163),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_185),
.B(n_187),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_168),
.B(n_141),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_148),
.Y(n_187)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_148),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_191),
.B(n_151),
.Y(n_209)
);

CKINVDCx16_ASAP7_75t_R g192 ( 
.A(n_163),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_156),
.B(n_142),
.Y(n_193)
);

XOR2xp5_ASAP7_75t_L g210 ( 
.A(n_193),
.B(n_196),
.Y(n_210)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_194),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_157),
.B(n_162),
.C(n_165),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_156),
.B(n_38),
.C(n_135),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_198),
.B(n_171),
.Y(n_211)
);

NAND3xp33_ASAP7_75t_L g204 ( 
.A(n_195),
.B(n_169),
.C(n_174),
.Y(n_204)
);

AOI21xp33_ASAP7_75t_L g229 ( 
.A1(n_204),
.A2(n_191),
.B(n_194),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_189),
.B(n_154),
.Y(n_205)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_205),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_196),
.B(n_164),
.Y(n_206)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_206),
.Y(n_236)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_207),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_208),
.A2(n_220),
.B1(n_200),
.B2(n_180),
.Y(n_233)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_209),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_211),
.B(n_212),
.C(n_183),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_L g212 ( 
.A(n_184),
.B(n_155),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_197),
.B(n_170),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_213),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_197),
.B(n_159),
.Y(n_214)
);

INVxp33_ASAP7_75t_L g245 ( 
.A(n_214),
.Y(n_245)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_195),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_215),
.B(n_217),
.Y(n_230)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_181),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_185),
.B(n_149),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_218),
.B(n_219),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_179),
.B(n_166),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_176),
.A2(n_146),
.B1(n_85),
.B2(n_31),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_SL g221 ( 
.A(n_186),
.B(n_28),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g232 ( 
.A(n_221),
.B(n_198),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_187),
.B(n_26),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_222),
.B(n_223),
.Y(n_239)
);

NOR3xp33_ASAP7_75t_L g223 ( 
.A(n_175),
.B(n_190),
.C(n_188),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_179),
.B(n_31),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_224),
.B(n_31),
.Y(n_238)
);

XOR2xp5_ASAP7_75t_L g261 ( 
.A(n_225),
.B(n_227),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_216),
.B(n_210),
.C(n_212),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_226),
.B(n_232),
.C(n_216),
.Y(n_247)
);

MAJx2_ASAP7_75t_L g227 ( 
.A(n_210),
.B(n_193),
.C(n_177),
.Y(n_227)
);

OAI21xp5_ASAP7_75t_SL g256 ( 
.A1(n_229),
.A2(n_237),
.B(n_240),
.Y(n_256)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_233),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_202),
.A2(n_176),
.B1(n_177),
.B2(n_182),
.Y(n_234)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_234),
.Y(n_262)
);

AOI21xp5_ASAP7_75t_L g237 ( 
.A1(n_201),
.A2(n_180),
.B(n_26),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_238),
.Y(n_260)
);

OAI21xp5_ASAP7_75t_SL g240 ( 
.A1(n_201),
.A2(n_1),
.B(n_2),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_211),
.A2(n_24),
.B1(n_30),
.B2(n_22),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_241),
.A2(n_243),
.B1(n_218),
.B2(n_209),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_219),
.A2(n_24),
.B1(n_2),
.B2(n_3),
.Y(n_243)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_246),
.Y(n_263)
);

XOR2xp5_ASAP7_75t_L g267 ( 
.A(n_247),
.B(n_261),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_242),
.A2(n_208),
.B1(n_220),
.B2(n_224),
.Y(n_248)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_248),
.Y(n_270)
);

FAx1_ASAP7_75t_SL g249 ( 
.A(n_228),
.B(n_221),
.CI(n_203),
.CON(n_249),
.SN(n_249)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_249),
.B(n_257),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_235),
.B(n_18),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_SL g271 ( 
.A(n_250),
.B(n_253),
.Y(n_271)
);

NOR2xp67_ASAP7_75t_SL g252 ( 
.A(n_230),
.B(n_9),
.Y(n_252)
);

OAI21xp5_ASAP7_75t_L g272 ( 
.A1(n_252),
.A2(n_238),
.B(n_13),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_245),
.B(n_18),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_225),
.B(n_18),
.C(n_28),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_254),
.B(n_255),
.C(n_244),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_226),
.B(n_236),
.C(n_232),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_240),
.B(n_26),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_SL g258 ( 
.A(n_231),
.B(n_15),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_258),
.B(n_259),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_243),
.B(n_13),
.Y(n_259)
);

AOI322xp5_ASAP7_75t_SL g264 ( 
.A1(n_252),
.A2(n_239),
.A3(n_231),
.B1(n_236),
.B2(n_227),
.C1(n_244),
.C2(n_234),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_SL g279 ( 
.A(n_264),
.B(n_274),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_265),
.B(n_260),
.C(n_262),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_255),
.B(n_237),
.C(n_228),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_266),
.B(n_267),
.C(n_269),
.Y(n_280)
);

NOR2x1_ASAP7_75t_L g268 ( 
.A(n_256),
.B(n_233),
.Y(n_268)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_268),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_247),
.B(n_242),
.C(n_241),
.Y(n_269)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_272),
.Y(n_281)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_251),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_251),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_275),
.A2(n_1),
.B1(n_4),
.B2(n_5),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_L g277 ( 
.A1(n_268),
.A2(n_262),
.B1(n_260),
.B2(n_248),
.Y(n_277)
);

AOI322xp5_ASAP7_75t_L g295 ( 
.A1(n_277),
.A2(n_8),
.A3(n_10),
.B1(n_9),
.B2(n_11),
.C1(n_7),
.C2(n_6),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_265),
.B(n_261),
.C(n_254),
.Y(n_282)
);

AOI21xp5_ASAP7_75t_L g296 ( 
.A1(n_282),
.A2(n_285),
.B(n_286),
.Y(n_296)
);

XOR2xp5_ASAP7_75t_L g283 ( 
.A(n_267),
.B(n_256),
.Y(n_283)
);

AND2x2_ASAP7_75t_L g291 ( 
.A(n_283),
.B(n_285),
.Y(n_291)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_284),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_266),
.B(n_246),
.C(n_249),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_269),
.B(n_249),
.C(n_3),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_270),
.A2(n_11),
.B1(n_10),
.B2(n_9),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_SL g289 ( 
.A(n_287),
.B(n_272),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g297 ( 
.A(n_288),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_289),
.B(n_292),
.Y(n_299)
);

AOI322xp5_ASAP7_75t_L g290 ( 
.A1(n_278),
.A2(n_270),
.A3(n_263),
.B1(n_273),
.B2(n_274),
.C1(n_271),
.C2(n_275),
.Y(n_290)
);

NOR2xp67_ASAP7_75t_SL g304 ( 
.A(n_290),
.B(n_295),
.Y(n_304)
);

AOI21xp5_ASAP7_75t_SL g300 ( 
.A1(n_291),
.A2(n_280),
.B(n_283),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_281),
.B(n_276),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_286),
.B(n_279),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_293),
.B(n_298),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_280),
.B(n_8),
.Y(n_298)
);

OAI21xp5_ASAP7_75t_SL g310 ( 
.A1(n_300),
.A2(n_301),
.B(n_302),
.Y(n_310)
);

NOR3xp33_ASAP7_75t_L g301 ( 
.A(n_296),
.B(n_282),
.C(n_5),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_297),
.B(n_4),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_294),
.B(n_5),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_305),
.B(n_306),
.C(n_290),
.Y(n_307)
);

INVx6_ASAP7_75t_L g306 ( 
.A(n_291),
.Y(n_306)
);

AOI21xp5_ASAP7_75t_L g311 ( 
.A1(n_307),
.A2(n_308),
.B(n_309),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_299),
.B(n_5),
.C(n_6),
.Y(n_308)
);

INVxp67_ASAP7_75t_L g309 ( 
.A(n_304),
.Y(n_309)
);

INVxp67_ASAP7_75t_L g312 ( 
.A(n_310),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_L g313 ( 
.A(n_312),
.B(n_303),
.Y(n_313)
);

MAJx2_ASAP7_75t_L g314 ( 
.A(n_313),
.B(n_311),
.C(n_6),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_L g315 ( 
.A(n_314),
.B(n_7),
.Y(n_315)
);


endmodule