module fake_ariane_2171_n_2612 (n_295, n_356, n_556, n_170, n_190, n_698, n_695, n_160, n_64, n_180, n_730, n_119, n_124, n_386, n_307, n_516, n_589, n_332, n_581, n_294, n_646, n_197, n_640, n_463, n_176, n_691, n_34, n_404, n_172, n_678, n_651, n_347, n_423, n_183, n_469, n_479, n_726, n_603, n_373, n_299, n_541, n_499, n_12, n_564, n_133, n_610, n_66, n_205, n_341, n_71, n_109, n_245, n_421, n_96, n_549, n_522, n_319, n_49, n_591, n_20, n_690, n_416, n_283, n_50, n_187, n_525, n_367, n_713, n_649, n_598, n_345, n_374, n_318, n_103, n_244, n_643, n_679, n_226, n_220, n_261, n_682, n_36, n_663, n_370, n_706, n_189, n_717, n_72, n_286, n_443, n_586, n_57, n_686, n_605, n_424, n_528, n_584, n_387, n_406, n_117, n_139, n_524, n_85, n_130, n_349, n_391, n_634, n_466, n_346, n_214, n_348, n_552, n_2, n_462, n_607, n_670, n_32, n_410, n_379, n_445, n_515, n_138, n_162, n_264, n_737, n_137, n_122, n_198, n_232, n_52, n_441, n_568, n_385, n_637, n_73, n_327, n_77, n_372, n_377, n_15, n_396, n_631, n_23, n_399, n_554, n_520, n_87, n_714, n_279, n_702, n_207, n_363, n_720, n_354, n_41, n_140, n_725, n_419, n_151, n_28, n_146, n_230, n_270, n_194, n_633, n_154, n_338, n_142, n_285, n_473, n_186, n_202, n_145, n_193, n_733, n_500, n_665, n_59, n_336, n_731, n_315, n_594, n_311, n_239, n_402, n_35, n_272, n_54, n_8, n_668, n_339, n_738, n_672, n_487, n_740, n_167, n_90, n_38, n_422, n_47, n_153, n_18, n_648, n_269, n_597, n_75, n_158, n_69, n_259, n_95, n_446, n_553, n_143, n_566, n_578, n_701, n_625, n_152, n_405, n_557, n_120, n_169, n_106, n_173, n_242, n_645, n_309, n_320, n_115, n_331, n_559, n_401, n_485, n_267, n_495, n_504, n_647, n_483, n_335, n_435, n_350, n_291, n_344, n_381, n_426, n_433, n_481, n_600, n_721, n_398, n_62, n_210, n_200, n_529, n_502, n_166, n_253, n_561, n_218, n_79, n_3, n_271, n_465, n_486, n_507, n_247, n_569, n_567, n_732, n_91, n_240, n_369, n_128, n_224, n_44, n_82, n_31, n_547, n_420, n_562, n_518, n_439, n_604, n_614, n_677, n_222, n_478, n_703, n_748, n_510, n_256, n_326, n_681, n_227, n_48, n_188, n_323, n_550, n_635, n_707, n_330, n_400, n_689, n_694, n_11, n_129, n_126, n_282, n_328, n_368, n_590, n_699, n_727, n_277, n_248, n_301, n_467, n_432, n_545, n_536, n_644, n_293, n_620, n_228, n_325, n_276, n_93, n_688, n_636, n_427, n_108, n_587, n_497, n_693, n_303, n_671, n_442, n_168, n_81, n_1, n_206, n_352, n_538, n_576, n_511, n_611, n_238, n_365, n_429, n_455, n_654, n_588, n_638, n_136, n_334, n_192, n_729, n_661, n_488, n_667, n_300, n_533, n_505, n_14, n_163, n_88, n_141, n_390, n_498, n_104, n_501, n_438, n_314, n_684, n_16, n_440, n_627, n_273, n_305, n_539, n_312, n_233, n_56, n_60, n_728, n_388, n_333, n_449, n_612, n_413, n_392, n_376, n_512, n_715, n_579, n_459, n_685, n_221, n_321, n_86, n_361, n_458, n_89, n_149, n_383, n_623, n_237, n_175, n_711, n_453, n_734, n_74, n_491, n_19, n_40, n_181, n_723, n_616, n_617, n_658, n_630, n_705, n_570, n_53, n_260, n_362, n_543, n_310, n_709, n_236, n_601, n_683, n_565, n_281, n_24, n_7, n_628, n_461, n_209, n_262, n_490, n_743, n_17, n_225, n_235, n_660, n_464, n_735, n_575, n_546, n_297, n_662, n_641, n_503, n_700, n_290, n_527, n_46, n_741, n_747, n_84, n_371, n_199, n_107, n_639, n_217, n_452, n_673, n_676, n_178, n_42, n_551, n_308, n_708, n_417, n_201, n_70, n_572, n_343, n_10, n_414, n_571, n_680, n_287, n_302, n_380, n_6, n_582, n_94, n_284, n_4, n_448, n_593, n_710, n_249, n_534, n_37, n_58, n_65, n_123, n_212, n_355, n_444, n_609, n_278, n_255, n_560, n_450, n_257, n_148, n_652, n_451, n_613, n_745, n_475, n_135, n_409, n_171, n_519, n_384, n_468, n_61, n_526, n_716, n_102, n_742, n_182, n_696, n_674, n_482, n_316, n_196, n_125, n_43, n_577, n_407, n_13, n_27, n_254, n_596, n_476, n_460, n_219, n_55, n_535, n_231, n_366, n_744, n_656, n_555, n_234, n_492, n_574, n_280, n_215, n_252, n_629, n_664, n_161, n_454, n_298, n_532, n_68, n_415, n_78, n_63, n_655, n_99, n_540, n_216, n_544, n_692, n_5, n_599, n_514, n_418, n_537, n_223, n_403, n_25, n_83, n_389, n_657, n_513, n_288, n_179, n_395, n_621, n_195, n_606, n_213, n_110, n_304, n_659, n_67, n_509, n_583, n_724, n_306, n_666, n_313, n_92, n_430, n_626, n_493, n_722, n_203, n_378, n_436, n_150, n_98, n_375, n_113, n_114, n_33, n_324, n_585, n_669, n_619, n_337, n_437, n_111, n_21, n_274, n_622, n_697, n_472, n_296, n_265, n_746, n_208, n_456, n_156, n_292, n_174, n_275, n_100, n_704, n_132, n_147, n_204, n_615, n_521, n_51, n_496, n_739, n_76, n_342, n_26, n_246, n_517, n_530, n_0, n_428, n_159, n_358, n_105, n_580, n_608, n_30, n_494, n_719, n_131, n_263, n_434, n_360, n_563, n_229, n_394, n_250, n_165, n_144, n_317, n_101, n_243, n_134, n_329, n_718, n_185, n_340, n_289, n_9, n_112, n_45, n_542, n_548, n_523, n_268, n_266, n_470, n_457, n_164, n_157, n_632, n_184, n_177, n_477, n_364, n_258, n_650, n_425, n_431, n_508, n_624, n_118, n_121, n_618, n_411, n_484, n_712, n_353, n_22, n_736, n_241, n_29, n_357, n_412, n_687, n_447, n_191, n_382, n_489, n_80, n_480, n_211, n_642, n_97, n_408, n_595, n_322, n_251, n_506, n_602, n_558, n_592, n_116, n_397, n_471, n_351, n_39, n_393, n_474, n_653, n_359, n_155, n_573, n_127, n_531, n_675, n_2612);

input n_295;
input n_356;
input n_556;
input n_170;
input n_190;
input n_698;
input n_695;
input n_160;
input n_64;
input n_180;
input n_730;
input n_119;
input n_124;
input n_386;
input n_307;
input n_516;
input n_589;
input n_332;
input n_581;
input n_294;
input n_646;
input n_197;
input n_640;
input n_463;
input n_176;
input n_691;
input n_34;
input n_404;
input n_172;
input n_678;
input n_651;
input n_347;
input n_423;
input n_183;
input n_469;
input n_479;
input n_726;
input n_603;
input n_373;
input n_299;
input n_541;
input n_499;
input n_12;
input n_564;
input n_133;
input n_610;
input n_66;
input n_205;
input n_341;
input n_71;
input n_109;
input n_245;
input n_421;
input n_96;
input n_549;
input n_522;
input n_319;
input n_49;
input n_591;
input n_20;
input n_690;
input n_416;
input n_283;
input n_50;
input n_187;
input n_525;
input n_367;
input n_713;
input n_649;
input n_598;
input n_345;
input n_374;
input n_318;
input n_103;
input n_244;
input n_643;
input n_679;
input n_226;
input n_220;
input n_261;
input n_682;
input n_36;
input n_663;
input n_370;
input n_706;
input n_189;
input n_717;
input n_72;
input n_286;
input n_443;
input n_586;
input n_57;
input n_686;
input n_605;
input n_424;
input n_528;
input n_584;
input n_387;
input n_406;
input n_117;
input n_139;
input n_524;
input n_85;
input n_130;
input n_349;
input n_391;
input n_634;
input n_466;
input n_346;
input n_214;
input n_348;
input n_552;
input n_2;
input n_462;
input n_607;
input n_670;
input n_32;
input n_410;
input n_379;
input n_445;
input n_515;
input n_138;
input n_162;
input n_264;
input n_737;
input n_137;
input n_122;
input n_198;
input n_232;
input n_52;
input n_441;
input n_568;
input n_385;
input n_637;
input n_73;
input n_327;
input n_77;
input n_372;
input n_377;
input n_15;
input n_396;
input n_631;
input n_23;
input n_399;
input n_554;
input n_520;
input n_87;
input n_714;
input n_279;
input n_702;
input n_207;
input n_363;
input n_720;
input n_354;
input n_41;
input n_140;
input n_725;
input n_419;
input n_151;
input n_28;
input n_146;
input n_230;
input n_270;
input n_194;
input n_633;
input n_154;
input n_338;
input n_142;
input n_285;
input n_473;
input n_186;
input n_202;
input n_145;
input n_193;
input n_733;
input n_500;
input n_665;
input n_59;
input n_336;
input n_731;
input n_315;
input n_594;
input n_311;
input n_239;
input n_402;
input n_35;
input n_272;
input n_54;
input n_8;
input n_668;
input n_339;
input n_738;
input n_672;
input n_487;
input n_740;
input n_167;
input n_90;
input n_38;
input n_422;
input n_47;
input n_153;
input n_18;
input n_648;
input n_269;
input n_597;
input n_75;
input n_158;
input n_69;
input n_259;
input n_95;
input n_446;
input n_553;
input n_143;
input n_566;
input n_578;
input n_701;
input n_625;
input n_152;
input n_405;
input n_557;
input n_120;
input n_169;
input n_106;
input n_173;
input n_242;
input n_645;
input n_309;
input n_320;
input n_115;
input n_331;
input n_559;
input n_401;
input n_485;
input n_267;
input n_495;
input n_504;
input n_647;
input n_483;
input n_335;
input n_435;
input n_350;
input n_291;
input n_344;
input n_381;
input n_426;
input n_433;
input n_481;
input n_600;
input n_721;
input n_398;
input n_62;
input n_210;
input n_200;
input n_529;
input n_502;
input n_166;
input n_253;
input n_561;
input n_218;
input n_79;
input n_3;
input n_271;
input n_465;
input n_486;
input n_507;
input n_247;
input n_569;
input n_567;
input n_732;
input n_91;
input n_240;
input n_369;
input n_128;
input n_224;
input n_44;
input n_82;
input n_31;
input n_547;
input n_420;
input n_562;
input n_518;
input n_439;
input n_604;
input n_614;
input n_677;
input n_222;
input n_478;
input n_703;
input n_748;
input n_510;
input n_256;
input n_326;
input n_681;
input n_227;
input n_48;
input n_188;
input n_323;
input n_550;
input n_635;
input n_707;
input n_330;
input n_400;
input n_689;
input n_694;
input n_11;
input n_129;
input n_126;
input n_282;
input n_328;
input n_368;
input n_590;
input n_699;
input n_727;
input n_277;
input n_248;
input n_301;
input n_467;
input n_432;
input n_545;
input n_536;
input n_644;
input n_293;
input n_620;
input n_228;
input n_325;
input n_276;
input n_93;
input n_688;
input n_636;
input n_427;
input n_108;
input n_587;
input n_497;
input n_693;
input n_303;
input n_671;
input n_442;
input n_168;
input n_81;
input n_1;
input n_206;
input n_352;
input n_538;
input n_576;
input n_511;
input n_611;
input n_238;
input n_365;
input n_429;
input n_455;
input n_654;
input n_588;
input n_638;
input n_136;
input n_334;
input n_192;
input n_729;
input n_661;
input n_488;
input n_667;
input n_300;
input n_533;
input n_505;
input n_14;
input n_163;
input n_88;
input n_141;
input n_390;
input n_498;
input n_104;
input n_501;
input n_438;
input n_314;
input n_684;
input n_16;
input n_440;
input n_627;
input n_273;
input n_305;
input n_539;
input n_312;
input n_233;
input n_56;
input n_60;
input n_728;
input n_388;
input n_333;
input n_449;
input n_612;
input n_413;
input n_392;
input n_376;
input n_512;
input n_715;
input n_579;
input n_459;
input n_685;
input n_221;
input n_321;
input n_86;
input n_361;
input n_458;
input n_89;
input n_149;
input n_383;
input n_623;
input n_237;
input n_175;
input n_711;
input n_453;
input n_734;
input n_74;
input n_491;
input n_19;
input n_40;
input n_181;
input n_723;
input n_616;
input n_617;
input n_658;
input n_630;
input n_705;
input n_570;
input n_53;
input n_260;
input n_362;
input n_543;
input n_310;
input n_709;
input n_236;
input n_601;
input n_683;
input n_565;
input n_281;
input n_24;
input n_7;
input n_628;
input n_461;
input n_209;
input n_262;
input n_490;
input n_743;
input n_17;
input n_225;
input n_235;
input n_660;
input n_464;
input n_735;
input n_575;
input n_546;
input n_297;
input n_662;
input n_641;
input n_503;
input n_700;
input n_290;
input n_527;
input n_46;
input n_741;
input n_747;
input n_84;
input n_371;
input n_199;
input n_107;
input n_639;
input n_217;
input n_452;
input n_673;
input n_676;
input n_178;
input n_42;
input n_551;
input n_308;
input n_708;
input n_417;
input n_201;
input n_70;
input n_572;
input n_343;
input n_10;
input n_414;
input n_571;
input n_680;
input n_287;
input n_302;
input n_380;
input n_6;
input n_582;
input n_94;
input n_284;
input n_4;
input n_448;
input n_593;
input n_710;
input n_249;
input n_534;
input n_37;
input n_58;
input n_65;
input n_123;
input n_212;
input n_355;
input n_444;
input n_609;
input n_278;
input n_255;
input n_560;
input n_450;
input n_257;
input n_148;
input n_652;
input n_451;
input n_613;
input n_745;
input n_475;
input n_135;
input n_409;
input n_171;
input n_519;
input n_384;
input n_468;
input n_61;
input n_526;
input n_716;
input n_102;
input n_742;
input n_182;
input n_696;
input n_674;
input n_482;
input n_316;
input n_196;
input n_125;
input n_43;
input n_577;
input n_407;
input n_13;
input n_27;
input n_254;
input n_596;
input n_476;
input n_460;
input n_219;
input n_55;
input n_535;
input n_231;
input n_366;
input n_744;
input n_656;
input n_555;
input n_234;
input n_492;
input n_574;
input n_280;
input n_215;
input n_252;
input n_629;
input n_664;
input n_161;
input n_454;
input n_298;
input n_532;
input n_68;
input n_415;
input n_78;
input n_63;
input n_655;
input n_99;
input n_540;
input n_216;
input n_544;
input n_692;
input n_5;
input n_599;
input n_514;
input n_418;
input n_537;
input n_223;
input n_403;
input n_25;
input n_83;
input n_389;
input n_657;
input n_513;
input n_288;
input n_179;
input n_395;
input n_621;
input n_195;
input n_606;
input n_213;
input n_110;
input n_304;
input n_659;
input n_67;
input n_509;
input n_583;
input n_724;
input n_306;
input n_666;
input n_313;
input n_92;
input n_430;
input n_626;
input n_493;
input n_722;
input n_203;
input n_378;
input n_436;
input n_150;
input n_98;
input n_375;
input n_113;
input n_114;
input n_33;
input n_324;
input n_585;
input n_669;
input n_619;
input n_337;
input n_437;
input n_111;
input n_21;
input n_274;
input n_622;
input n_697;
input n_472;
input n_296;
input n_265;
input n_746;
input n_208;
input n_456;
input n_156;
input n_292;
input n_174;
input n_275;
input n_100;
input n_704;
input n_132;
input n_147;
input n_204;
input n_615;
input n_521;
input n_51;
input n_496;
input n_739;
input n_76;
input n_342;
input n_26;
input n_246;
input n_517;
input n_530;
input n_0;
input n_428;
input n_159;
input n_358;
input n_105;
input n_580;
input n_608;
input n_30;
input n_494;
input n_719;
input n_131;
input n_263;
input n_434;
input n_360;
input n_563;
input n_229;
input n_394;
input n_250;
input n_165;
input n_144;
input n_317;
input n_101;
input n_243;
input n_134;
input n_329;
input n_718;
input n_185;
input n_340;
input n_289;
input n_9;
input n_112;
input n_45;
input n_542;
input n_548;
input n_523;
input n_268;
input n_266;
input n_470;
input n_457;
input n_164;
input n_157;
input n_632;
input n_184;
input n_177;
input n_477;
input n_364;
input n_258;
input n_650;
input n_425;
input n_431;
input n_508;
input n_624;
input n_118;
input n_121;
input n_618;
input n_411;
input n_484;
input n_712;
input n_353;
input n_22;
input n_736;
input n_241;
input n_29;
input n_357;
input n_412;
input n_687;
input n_447;
input n_191;
input n_382;
input n_489;
input n_80;
input n_480;
input n_211;
input n_642;
input n_97;
input n_408;
input n_595;
input n_322;
input n_251;
input n_506;
input n_602;
input n_558;
input n_592;
input n_116;
input n_397;
input n_471;
input n_351;
input n_39;
input n_393;
input n_474;
input n_653;
input n_359;
input n_155;
input n_573;
input n_127;
input n_531;
input n_675;

output n_2612;

wire n_913;
wire n_1681;
wire n_2163;
wire n_1486;
wire n_1507;
wire n_1938;
wire n_2484;
wire n_1174;
wire n_2346;
wire n_1469;
wire n_1353;
wire n_1355;
wire n_2131;
wire n_2559;
wire n_2500;
wire n_2509;
wire n_1383;
wire n_2182;
wire n_2135;
wire n_2334;
wire n_1250;
wire n_2030;
wire n_1169;
wire n_789;
wire n_850;
wire n_1916;
wire n_1713;
wire n_1436;
wire n_2407;
wire n_1109;
wire n_1430;
wire n_2537;
wire n_2002;
wire n_1463;
wire n_2243;
wire n_1238;
wire n_2011;
wire n_1515;
wire n_817;
wire n_1837;
wire n_924;
wire n_781;
wire n_2013;
wire n_1566;
wire n_2006;
wire n_952;
wire n_864;
wire n_2446;
wire n_1096;
wire n_1379;
wire n_2436;
wire n_2376;
wire n_2367;
wire n_1706;
wire n_2207;
wire n_2461;
wire n_1214;
wire n_1839;
wire n_1246;
wire n_1138;
wire n_2042;
wire n_2123;
wire n_1853;
wire n_764;
wire n_1503;
wire n_2238;
wire n_2529;
wire n_2374;
wire n_1196;
wire n_1181;
wire n_1999;
wire n_2380;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_1298;
wire n_1745;
wire n_1366;
wire n_2084;
wire n_2278;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1835;
wire n_1457;
wire n_2482;
wire n_1682;
wire n_1836;
wire n_870;
wire n_2547;
wire n_1453;
wire n_945;
wire n_958;
wire n_2554;
wire n_2248;
wire n_813;
wire n_1985;
wire n_2288;
wire n_995;
wire n_2579;
wire n_1909;
wire n_2156;
wire n_1184;
wire n_1961;
wire n_1535;
wire n_754;
wire n_903;
wire n_871;
wire n_2323;
wire n_1073;
wire n_1979;
wire n_1277;
wire n_2107;
wire n_1746;
wire n_829;
wire n_1761;
wire n_1062;
wire n_1690;
wire n_2221;
wire n_1283;
wire n_2317;
wire n_1974;
wire n_1736;
wire n_1018;
wire n_2342;
wire n_2200;
wire n_2442;
wire n_953;
wire n_1364;
wire n_2390;
wire n_1888;
wire n_1224;
wire n_2109;
wire n_1425;
wire n_2322;
wire n_1107;
wire n_1688;
wire n_989;
wire n_1944;
wire n_2233;
wire n_2370;
wire n_1988;
wire n_795;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_1936;
wire n_2149;
wire n_2277;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_770;
wire n_1514;
wire n_2539;
wire n_1528;
wire n_901;
wire n_2078;
wire n_1145;
wire n_971;
wire n_2359;
wire n_2201;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_2049;
wire n_1522;
wire n_1207;
wire n_786;
wire n_1404;
wire n_868;
wire n_2232;
wire n_1847;
wire n_2458;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_2227;
wire n_2301;
wire n_1539;
wire n_884;
wire n_1851;
wire n_2162;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_2192;
wire n_1676;
wire n_1085;
wire n_1636;
wire n_823;
wire n_1900;
wire n_1074;
wire n_859;
wire n_1765;
wire n_1889;
wire n_1977;
wire n_863;
wire n_1254;
wire n_929;
wire n_2433;
wire n_1703;
wire n_899;
wire n_2332;
wire n_2391;
wire n_1295;
wire n_2060;
wire n_1850;
wire n_2004;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_2571;
wire n_2427;
wire n_2098;
wire n_1751;
wire n_1917;
wire n_2456;
wire n_1924;
wire n_1560;
wire n_1654;
wire n_2341;
wire n_1548;
wire n_1811;
wire n_2045;
wire n_2575;
wire n_1396;
wire n_1230;
wire n_1840;
wire n_1597;
wire n_1771;
wire n_1544;
wire n_844;
wire n_1012;
wire n_1267;
wire n_2061;
wire n_2094;
wire n_2512;
wire n_1354;
wire n_1790;
wire n_1213;
wire n_2382;
wire n_2043;
wire n_780;
wire n_2349;
wire n_1918;
wire n_1443;
wire n_1021;
wire n_2595;
wire n_1465;
wire n_1949;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_942;
wire n_1437;
wire n_2077;
wire n_1378;
wire n_1121;
wire n_1416;
wire n_1461;
wire n_1391;
wire n_1947;
wire n_1599;
wire n_1876;
wire n_1006;
wire n_1830;
wire n_2527;
wire n_1112;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_2466;
wire n_2038;
wire n_2263;
wire n_2568;
wire n_2116;
wire n_2271;
wire n_2145;
wire n_2326;
wire n_1838;
wire n_1594;
wire n_1935;
wire n_1716;
wire n_1872;
wire n_1585;
wire n_2281;
wire n_1432;
wire n_2245;
wire n_1108;
wire n_851;
wire n_1590;
wire n_1351;
wire n_2216;
wire n_1274;
wire n_2426;
wire n_1819;
wire n_947;
wire n_2134;
wire n_1260;
wire n_930;
wire n_1179;
wire n_1442;
wire n_798;
wire n_1833;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_1884;
wire n_1555;
wire n_1842;
wire n_2499;
wire n_2549;
wire n_1253;
wire n_1468;
wire n_762;
wire n_1661;
wire n_804;
wire n_1656;
wire n_1382;
wire n_966;
wire n_992;
wire n_955;
wire n_1182;
wire n_794;
wire n_2166;
wire n_1692;
wire n_2611;
wire n_1562;
wire n_2185;
wire n_2398;
wire n_1376;
wire n_1292;
wire n_1178;
wire n_1972;
wire n_2015;
wire n_1435;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_2202;
wire n_2072;
wire n_2415;
wire n_2087;
wire n_1491;
wire n_931;
wire n_967;
wire n_1083;
wire n_2161;
wire n_1418;
wire n_1357;
wire n_1079;
wire n_1787;
wire n_2462;
wire n_1389;
wire n_2155;
wire n_1139;
wire n_2439;
wire n_1312;
wire n_1717;
wire n_1812;
wire n_824;
wire n_2172;
wire n_2601;
wire n_892;
wire n_1880;
wire n_959;
wire n_2365;
wire n_2257;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_2219;
wire n_1855;
wire n_2100;
wire n_2333;
wire n_990;
wire n_1623;
wire n_1903;
wire n_867;
wire n_2147;
wire n_2435;
wire n_1226;
wire n_2224;
wire n_944;
wire n_749;
wire n_1932;
wire n_1780;
wire n_1970;
wire n_1920;
wire n_2083;
wire n_815;
wire n_2167;
wire n_2293;
wire n_1340;
wire n_1240;
wire n_1087;
wire n_2400;
wire n_2388;
wire n_2273;
wire n_1433;
wire n_1911;
wire n_2567;
wire n_2557;
wire n_1825;
wire n_1908;
wire n_1155;
wire n_2598;
wire n_1071;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1832;
wire n_1841;
wire n_1680;
wire n_2066;
wire n_2302;
wire n_964;
wire n_1627;
wire n_2220;
wire n_2294;
wire n_2274;
wire n_974;
wire n_1731;
wire n_799;
wire n_1147;
wire n_2378;
wire n_2467;
wire n_965;
wire n_1914;
wire n_2253;
wire n_934;
wire n_2213;
wire n_1447;
wire n_2363;
wire n_1220;
wire n_2019;
wire n_2130;
wire n_1674;
wire n_2021;
wire n_2025;
wire n_2160;
wire n_1992;
wire n_1209;
wire n_1563;
wire n_1020;
wire n_2507;
wire n_2142;
wire n_1633;
wire n_1913;
wire n_2069;
wire n_2495;
wire n_1058;
wire n_2328;
wire n_2434;
wire n_1042;
wire n_1234;
wire n_2311;
wire n_1578;
wire n_2261;
wire n_1455;
wire n_2287;
wire n_836;
wire n_2223;
wire n_1279;
wire n_2473;
wire n_2144;
wire n_2511;
wire n_1029;
wire n_1247;
wire n_760;
wire n_2438;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_1111;
wire n_970;
wire n_1689;
wire n_2535;
wire n_1255;
wire n_1646;
wire n_2262;
wire n_2565;
wire n_1237;
wire n_927;
wire n_1095;
wire n_1728;
wire n_2335;
wire n_2120;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_2041;
wire n_2113;
wire n_1933;
wire n_1651;
wire n_1387;
wire n_1263;
wire n_1817;
wire n_2404;
wire n_2168;
wire n_2312;
wire n_1826;
wire n_2483;
wire n_1951;
wire n_2490;
wire n_1032;
wire n_1217;
wire n_2558;
wire n_1496;
wire n_1592;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_2132;
wire n_980;
wire n_1618;
wire n_1869;
wire n_1743;
wire n_905;
wire n_926;
wire n_1943;
wire n_2296;
wire n_1802;
wire n_2178;
wire n_2112;
wire n_1163;
wire n_1795;
wire n_1384;
wire n_2237;
wire n_2146;
wire n_1868;
wire n_1501;
wire n_2241;
wire n_2373;
wire n_1173;
wire n_2350;
wire n_1068;
wire n_1198;
wire n_2531;
wire n_1570;
wire n_2099;
wire n_1518;
wire n_1456;
wire n_1879;
wire n_1886;
wire n_1648;
wire n_2187;
wire n_1413;
wire n_2481;
wire n_2129;
wire n_855;
wire n_2327;
wire n_808;
wire n_1365;
wire n_2476;
wire n_2059;
wire n_2437;
wire n_1439;
wire n_814;
wire n_2074;
wire n_1665;
wire n_1287;
wire n_1611;
wire n_2122;
wire n_2399;
wire n_1414;
wire n_1134;
wire n_2067;
wire n_1484;
wire n_1901;
wire n_2055;
wire n_2027;
wire n_1423;
wire n_2117;
wire n_1609;
wire n_1053;
wire n_1939;
wire n_2308;
wire n_2242;
wire n_1906;
wire n_1899;
wire n_2195;
wire n_2194;
wire n_1467;
wire n_1828;
wire n_2159;
wire n_1798;
wire n_1304;
wire n_1608;
wire n_1744;
wire n_2267;
wire n_1105;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_2102;
wire n_874;
wire n_2286;
wire n_2023;
wire n_1278;
wire n_983;
wire n_2599;
wire n_2075;
wire n_1726;
wire n_2523;
wire n_1945;
wire n_1015;
wire n_2418;
wire n_1377;
wire n_1162;
wire n_1614;
wire n_2031;
wire n_2496;
wire n_2118;
wire n_1740;
wire n_1602;
wire n_1098;
wire n_1490;
wire n_2338;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_2225;
wire n_986;
wire n_1104;
wire n_1963;
wire n_887;
wire n_2057;
wire n_2218;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_2593;
wire n_1693;
wire n_2125;
wire n_1132;
wire n_1156;
wire n_2184;
wire n_1823;
wire n_1120;
wire n_1202;
wire n_2254;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_2033;
wire n_957;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_2217;
wire n_2226;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1863;
wire n_1763;
wire n_1666;
wire n_1500;
wire n_2214;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_2256;
wire n_1189;
wire n_1089;
wire n_1859;
wire n_1502;
wire n_1523;
wire n_2190;
wire n_1478;
wire n_1883;
wire n_2516;
wire n_2555;
wire n_1969;
wire n_1005;
wire n_2379;
wire n_1294;
wire n_1667;
wire n_845;
wire n_888;
wire n_2300;
wire n_1649;
wire n_2452;
wire n_1677;
wire n_2470;
wire n_1927;
wire n_1297;
wire n_1708;
wire n_1222;
wire n_2284;
wire n_1844;
wire n_2283;
wire n_2526;
wire n_1957;
wire n_1953;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_1919;
wire n_1791;
wire n_2508;
wire n_2124;
wire n_1894;
wire n_1460;
wire n_1239;
wire n_2594;
wire n_2266;
wire n_2449;
wire n_890;
wire n_842;
wire n_1898;
wire n_1741;
wire n_1572;
wire n_1907;
wire n_1793;
wire n_1373;
wire n_1081;
wire n_1975;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_2119;
wire n_769;
wire n_1797;
wire n_2366;
wire n_2493;
wire n_1753;
wire n_1990;
wire n_1372;
wire n_832;
wire n_1895;
wire n_2474;
wire n_982;
wire n_1800;
wire n_915;
wire n_1075;
wire n_2008;
wire n_1331;
wire n_1890;
wire n_1529;
wire n_1227;
wire n_2127;
wire n_1734;
wire n_1860;
wire n_2460;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_837;
wire n_812;
wire n_2448;
wire n_2211;
wire n_2292;
wire n_2480;
wire n_951;
wire n_862;
wire n_1700;
wire n_1332;
wire n_2306;
wire n_1854;
wire n_1747;
wire n_2071;
wire n_2424;
wire n_1206;
wire n_1729;
wire n_1508;
wire n_2414;
wire n_2082;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_2389;
wire n_1309;
wire n_999;
wire n_2280;
wire n_1766;
wire n_1338;
wire n_1342;
wire n_1867;
wire n_852;
wire n_1394;
wire n_2576;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_2140;
wire n_873;
wire n_1301;
wire n_1748;
wire n_2157;
wire n_1966;
wire n_1243;
wire n_2171;
wire n_2468;
wire n_1400;
wire n_2035;
wire n_1466;
wire n_1513;
wire n_1527;
wire n_2581;
wire n_1783;
wire n_2494;
wire n_1538;
wire n_2457;
wire n_2128;
wire n_1037;
wire n_1329;
wire n_1993;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1954;
wire n_1668;
wire n_1878;
wire n_2540;
wire n_1605;
wire n_1078;
wire n_2486;
wire n_1897;
wire n_2520;
wire n_2137;
wire n_1161;
wire n_2489;
wire n_811;
wire n_791;
wire n_876;
wire n_1191;
wire n_2492;
wire n_1025;
wire n_1215;
wire n_1449;
wire n_2337;
wire n_2265;
wire n_797;
wire n_2026;
wire n_1786;
wire n_1327;
wire n_1475;
wire n_1804;
wire n_2106;
wire n_1406;
wire n_1405;
wire n_2272;
wire n_1757;
wire n_1499;
wire n_1318;
wire n_854;
wire n_2091;
wire n_1632;
wire n_1769;
wire n_1929;
wire n_1950;
wire n_2264;
wire n_805;
wire n_2032;
wire n_2090;
wire n_1658;
wire n_2249;
wire n_1072;
wire n_1526;
wire n_1305;
wire n_1596;
wire n_2348;
wire n_1281;
wire n_2364;
wire n_1997;
wire n_2574;
wire n_1137;
wire n_1873;
wire n_1258;
wire n_1476;
wire n_1524;
wire n_1733;
wire n_1856;
wire n_2016;
wire n_1118;
wire n_943;
wire n_1874;
wire n_1293;
wire n_961;
wire n_1046;
wire n_1807;
wire n_1123;
wire n_1657;
wire n_878;
wire n_1784;
wire n_771;
wire n_1321;
wire n_752;
wire n_2307;
wire n_1488;
wire n_985;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_2295;
wire n_806;
wire n_1984;
wire n_1350;
wire n_1556;
wire n_1561;
wire n_2412;
wire n_1352;
wire n_2405;
wire n_1824;
wire n_2606;
wire n_1492;
wire n_2383;
wire n_1441;
wire n_1822;
wire n_1616;
wire n_2416;
wire n_819;
wire n_2386;
wire n_1971;
wire n_1429;
wire n_1324;
wire n_2064;
wire n_2353;
wire n_2528;
wire n_1778;
wire n_1776;
wire n_1154;
wire n_1557;
wire n_1759;
wire n_1829;
wire n_2325;
wire n_1130;
wire n_1450;
wire n_756;
wire n_2022;
wire n_1016;
wire n_2298;
wire n_1149;
wire n_1505;
wire n_2408;
wire n_2320;
wire n_979;
wire n_2329;
wire n_2570;
wire n_1642;
wire n_2417;
wire n_2525;
wire n_1815;
wire n_897;
wire n_2546;
wire n_949;
wire n_2454;
wire n_1493;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_2354;
wire n_1864;
wire n_1887;
wire n_1208;
wire n_1987;
wire n_2368;
wire n_802;
wire n_1151;
wire n_960;
wire n_2352;
wire n_2502;
wire n_1256;
wire n_2170;
wire n_790;
wire n_2244;
wire n_2143;
wire n_2393;
wire n_2377;
wire n_1577;
wire n_1448;
wire n_2198;
wire n_1009;
wire n_1133;
wire n_883;
wire n_1852;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_2410;
wire n_2314;
wire n_2477;
wire n_2279;
wire n_2222;
wire n_1995;
wire n_1877;
wire n_1397;
wire n_1052;
wire n_1333;
wire n_1306;
wire n_1849;
wire n_2076;
wire n_2133;
wire n_2203;
wire n_833;
wire n_1426;
wire n_2250;
wire n_2497;
wire n_2247;
wire n_2230;
wire n_879;
wire n_1117;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_2001;
wire n_1047;
wire n_2506;
wire n_1472;
wire n_2413;
wire n_1593;
wire n_2610;
wire n_1050;
wire n_2158;
wire n_2578;
wire n_2607;
wire n_2285;
wire n_1288;
wire n_1201;
wire n_2605;
wire n_858;
wire n_1185;
wire n_2475;
wire n_2173;
wire n_1035;
wire n_1143;
wire n_2070;
wire n_2136;
wire n_1090;
wire n_2403;
wire n_1367;
wire n_2044;
wire n_928;
wire n_1153;
wire n_1103;
wire n_825;
wire n_1565;
wire n_1192;
wire n_894;
wire n_1380;
wire n_1624;
wire n_1801;
wire n_1291;
wire n_2020;
wire n_2310;
wire n_1045;
wire n_1160;
wire n_1882;
wire n_1976;
wire n_1023;
wire n_1881;
wire n_988;
wire n_914;
wire n_1116;
wire n_1958;
wire n_1511;
wire n_2177;
wire n_1422;
wire n_1965;
wire n_1197;
wire n_1165;
wire n_1641;
wire n_1517;
wire n_2036;
wire n_843;
wire n_2003;
wire n_2533;
wire n_2210;
wire n_1307;
wire n_1128;
wire n_2053;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_2343;
wire n_775;
wire n_2419;
wire n_1049;
wire n_2330;
wire n_869;
wire n_846;
wire n_1398;
wire n_1921;
wire n_2450;
wire n_2411;
wire n_1356;
wire n_1341;
wire n_2234;
wire n_2309;
wire n_1504;
wire n_1955;
wire n_2110;
wire n_2431;
wire n_1773;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_2401;
wire n_889;
wire n_1549;
wire n_1066;
wire n_2588;
wire n_2331;
wire n_935;
wire n_2478;
wire n_911;
wire n_2608;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_1534;
wire n_1948;
wire n_810;
wire n_1290;
wire n_1959;
wire n_2396;
wire n_1362;
wire n_1559;
wire n_2121;
wire n_1300;
wire n_1960;
wire n_2068;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_2553;
wire n_907;
wire n_1454;
wire n_2592;
wire n_2459;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_1622;
wire n_1135;
wire n_2566;
wire n_918;
wire n_1968;
wire n_1885;
wire n_2196;
wire n_1038;
wire n_2371;
wire n_1978;
wire n_1521;
wire n_1694;
wire n_1940;
wire n_1695;
wire n_2560;
wire n_1164;
wire n_2313;
wire n_1193;
wire n_1345;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_1774;
wire n_2609;
wire n_2561;
wire n_1166;
wire n_1056;
wire n_2007;
wire n_1994;
wire n_1767;
wire n_1040;
wire n_1158;
wire n_1973;
wire n_1444;
wire n_1803;
wire n_820;
wire n_1749;
wire n_872;
wire n_1653;
wire n_2303;
wire n_1157;
wire n_1584;
wire n_848;
wire n_1664;
wire n_1739;
wire n_1814;
wire n_2154;
wire n_2441;
wire n_2236;
wire n_1789;
wire n_763;
wire n_1986;
wire n_2174;
wire n_2054;
wire n_1857;
wire n_2315;
wire n_984;
wire n_1687;
wire n_2073;
wire n_2150;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_2498;
wire n_800;
wire n_2046;
wire n_1816;
wire n_1910;
wire n_1756;
wire n_1606;
wire n_2189;
wire n_1587;
wire n_2093;
wire n_2340;
wire n_2018;
wire n_1772;
wire n_2444;
wire n_2602;
wire n_1014;
wire n_2204;
wire n_1427;
wire n_1481;
wire n_2040;
wire n_1311;
wire n_2199;
wire n_1956;
wire n_1589;
wire n_2151;
wire n_1100;
wire n_875;
wire n_1617;
wire n_2455;
wire n_827;
wire n_2600;
wire n_2231;
wire n_1626;
wire n_1962;
wire n_1335;
wire n_1715;
wire n_2305;
wire n_880;
wire n_793;
wire n_2114;
wire n_1175;
wire n_2289;
wire n_2530;
wire n_2299;
wire n_751;
wire n_1027;
wire n_1070;
wire n_2406;
wire n_1621;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_1785;
wire n_792;
wire n_1262;
wire n_1942;
wire n_2180;
wire n_1579;
wire n_2181;
wire n_2014;
wire n_975;
wire n_1645;
wire n_923;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1893;
wire n_1183;
wire n_1326;
wire n_2276;
wire n_1805;
wire n_2282;
wire n_981;
wire n_2141;
wire n_1110;
wire n_1758;
wire n_2503;
wire n_2270;
wire n_2443;
wire n_1407;
wire n_2465;
wire n_1204;
wire n_1554;
wire n_994;
wire n_2428;
wire n_2586;
wire n_1360;
wire n_973;
wire n_972;
wire n_2251;
wire n_856;
wire n_2572;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_2010;
wire n_1054;
wire n_1679;
wire n_2126;
wire n_1952;
wire n_2425;
wire n_2394;
wire n_1858;
wire n_1678;
wire n_2589;
wire n_1482;
wire n_1361;
wire n_2356;
wire n_1601;
wire n_1057;
wire n_2487;
wire n_1834;
wire n_1011;
wire n_978;
wire n_1520;
wire n_2534;
wire n_2488;
wire n_1509;
wire n_828;
wire n_1411;
wire n_1359;
wire n_1721;
wire n_2564;
wire n_2591;
wire n_1445;
wire n_1317;
wire n_2050;
wire n_2197;
wire n_783;
wire n_2550;
wire n_1127;
wire n_1536;
wire n_1471;
wire n_2385;
wire n_2387;
wire n_1008;
wire n_1024;
wire n_830;
wire n_2291;
wire n_1980;
wire n_2518;
wire n_987;
wire n_936;
wire n_2510;
wire n_1620;
wire n_2501;
wire n_2542;
wire n_1385;
wire n_1525;
wire n_1998;
wire n_2165;
wire n_2604;
wire n_1775;
wire n_788;
wire n_908;
wire n_1036;
wire n_2169;
wire n_2603;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_969;
wire n_2028;
wire n_919;
wire n_1663;
wire n_2092;
wire n_2175;
wire n_1625;
wire n_2086;
wire n_1926;
wire n_2402;
wire n_1458;
wire n_1630;
wire n_1720;
wire n_2409;
wire n_2176;
wire n_1412;
wire n_1738;
wire n_1550;
wire n_1358;
wire n_1200;
wire n_826;
wire n_2453;
wire n_2344;
wire n_1922;
wire n_1735;
wire n_1788;
wire n_940;
wire n_2392;
wire n_1537;
wire n_2138;
wire n_2065;
wire n_2543;
wire n_2321;
wire n_1077;
wire n_2597;
wire n_956;
wire n_1930;
wire n_765;
wire n_1809;
wire n_1843;
wire n_1904;
wire n_2000;
wire n_1268;
wire n_2395;
wire n_917;
wire n_1271;
wire n_2096;
wire n_2440;
wire n_2556;
wire n_2186;
wire n_1530;
wire n_2215;
wire n_1170;
wire n_2258;
wire n_1261;
wire n_2471;
wire n_898;
wire n_857;
wire n_968;
wire n_1067;
wire n_1235;
wire n_1323;
wire n_2584;
wire n_2375;
wire n_1462;
wire n_1937;
wire n_2012;
wire n_1064;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_2039;
wire n_1755;
wire n_1285;
wire n_761;
wire n_2212;
wire n_1813;
wire n_2268;
wire n_1452;
wire n_1573;
wire n_2569;
wire n_758;
wire n_2252;
wire n_2111;
wire n_2420;
wire n_1996;
wire n_1106;
wire n_2009;
wire n_784;
wire n_816;
wire n_1322;
wire n_2583;
wire n_1473;
wire n_835;
wire n_1076;
wire n_2024;
wire n_1348;
wire n_753;
wire n_2445;
wire n_1770;
wire n_1003;
wire n_2469;
wire n_1125;
wire n_2103;
wire n_2358;
wire n_1710;
wire n_1865;
wire n_2522;
wire n_2463;
wire n_1344;
wire n_2355;
wire n_1390;
wire n_2580;
wire n_1792;
wire n_2062;
wire n_1141;
wire n_1629;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_2153;
wire n_2324;
wire n_1510;
wire n_2505;
wire n_2139;
wire n_1099;
wire n_839;
wire n_1754;
wire n_759;
wire n_2397;
wire n_2521;
wire n_1727;
wire n_2235;
wire n_1991;
wire n_1575;
wire n_1848;
wire n_1892;
wire n_1172;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_2351;
wire n_2260;
wire n_1660;
wire n_1315;
wire n_1902;
wire n_997;
wire n_2206;
wire n_2541;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_2347;
wire n_1152;
wire n_2447;
wire n_2034;
wire n_1845;
wire n_2538;
wire n_1934;
wire n_2101;
wire n_2577;
wire n_921;
wire n_2362;
wire n_1615;
wire n_1236;
wire n_2104;
wire n_1265;
wire n_1576;
wire n_2105;
wire n_1470;
wire n_1533;
wire n_1806;
wire n_2372;
wire n_2552;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1684;
wire n_1673;
wire n_2422;
wire n_1334;
wire n_2290;
wire n_2088;
wire n_1275;
wire n_904;
wire n_2005;
wire n_2048;
wire n_1696;
wire n_1875;
wire n_1059;
wire n_2429;
wire n_2108;
wire n_1039;
wire n_2246;
wire n_1150;
wire n_977;
wire n_2339;
wire n_1628;
wire n_1289;
wire n_1831;
wire n_2532;
wire n_2191;
wire n_1497;
wire n_1866;
wire n_2472;
wire n_2056;
wire n_1136;
wire n_2515;
wire n_1782;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_838;
wire n_1558;
wire n_1941;
wire n_1316;
wire n_2519;
wire n_950;
wire n_1017;
wire n_1915;
wire n_2360;
wire n_1393;
wire n_2240;
wire n_1369;
wire n_1781;
wire n_2544;
wire n_809;
wire n_2085;
wire n_2432;
wire n_1686;
wire n_1964;
wire n_881;
wire n_1477;
wire n_1019;
wire n_1777;
wire n_2188;
wire n_1982;
wire n_2097;
wire n_2430;
wire n_2504;
wire n_910;
wire n_939;
wire n_1410;
wire n_2297;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_1223;
wire n_2545;
wire n_1768;
wire n_2513;
wire n_2193;
wire n_2369;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1983;
wire n_1041;
wire n_2451;
wire n_2115;
wire n_993;
wire n_1862;
wire n_948;
wire n_2017;
wire n_922;
wire n_1004;
wire n_1810;
wire n_2587;
wire n_1347;
wire n_860;
wire n_1043;
wire n_1923;
wire n_1764;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_1571;
wire n_1698;
wire n_1337;
wire n_774;
wire n_1946;
wire n_2148;
wire n_933;
wire n_1779;
wire n_2562;
wire n_954;
wire n_2051;
wire n_1168;
wire n_1821;
wire n_1310;
wire n_1591;
wire n_2585;
wire n_1229;
wire n_1683;
wire n_2582;
wire n_2548;
wire n_1896;
wire n_2164;
wire n_1732;
wire n_2381;
wire n_1967;
wire n_2384;
wire n_2179;
wire n_1280;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_768;
wire n_1091;
wire n_2052;
wire n_2485;
wire n_1063;
wire n_991;
wire n_2205;
wire n_2183;
wire n_2275;
wire n_2563;
wire n_1724;
wire n_1670;
wire n_1707;
wire n_1799;
wire n_2080;
wire n_2058;
wire n_1126;
wire n_2357;
wire n_2029;
wire n_1846;
wire n_1912;
wire n_938;
wire n_1891;
wire n_1328;
wire n_895;
wire n_1639;
wire n_2209;
wire n_2421;
wire n_1302;
wire n_1000;
wire n_1581;
wire n_1928;
wire n_946;
wire n_757;
wire n_2047;
wire n_1655;
wire n_1818;
wire n_1146;
wire n_1634;
wire n_2596;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_2269;
wire n_2081;
wire n_1474;
wire n_937;
wire n_2536;
wire n_2524;
wire n_1583;
wire n_1604;
wire n_1631;
wire n_1702;
wire n_1794;
wire n_1375;
wire n_1232;
wire n_1211;
wire n_996;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_2318;
wire n_1827;
wire n_866;
wire n_925;
wire n_1752;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_2361;
wire n_1115;
wire n_2229;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_2551;
wire n_1102;
wire n_2255;
wire n_1129;
wire n_1252;
wire n_2239;
wire n_1464;
wire n_1296;
wire n_773;
wire n_2316;
wire n_2464;
wire n_1010;
wire n_882;
wire n_2304;
wire n_1249;
wire n_803;
wire n_1871;
wire n_2514;
wire n_1434;
wire n_1905;
wire n_1569;
wire n_2573;
wire n_2336;
wire n_1662;
wire n_1299;
wire n_1870;
wire n_2063;
wire n_1925;
wire n_782;
wire n_2491;
wire n_1861;
wire n_2079;
wire n_1228;
wire n_2319;
wire n_2152;
wire n_2517;
wire n_1931;
wire n_1244;
wire n_1796;
wire n_2259;
wire n_849;
wire n_2095;
wire n_1820;
wire n_2590;
wire n_1251;
wire n_1989;
wire n_1421;
wire n_2208;
wire n_2423;
wire n_1762;
wire n_1233;
wire n_1808;
wire n_1574;
wire n_1672;
wire n_2228;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_2479;
wire n_886;
wire n_1069;
wire n_1981;
wire n_2037;
wire n_1308;
wire n_796;
wire n_2345;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_2089;
wire n_1487;

CKINVDCx5p33_ASAP7_75t_R g749 ( 
.A(n_201),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_238),
.Y(n_750)
);

BUFx8_ASAP7_75t_SL g751 ( 
.A(n_142),
.Y(n_751)
);

INVx2_ASAP7_75t_SL g752 ( 
.A(n_149),
.Y(n_752)
);

INVx1_ASAP7_75t_SL g753 ( 
.A(n_664),
.Y(n_753)
);

BUFx2_ASAP7_75t_L g754 ( 
.A(n_731),
.Y(n_754)
);

CKINVDCx5p33_ASAP7_75t_R g755 ( 
.A(n_631),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_259),
.Y(n_756)
);

BUFx3_ASAP7_75t_L g757 ( 
.A(n_391),
.Y(n_757)
);

CKINVDCx5p33_ASAP7_75t_R g758 ( 
.A(n_410),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_376),
.Y(n_759)
);

CKINVDCx5p33_ASAP7_75t_R g760 ( 
.A(n_224),
.Y(n_760)
);

CKINVDCx5p33_ASAP7_75t_R g761 ( 
.A(n_663),
.Y(n_761)
);

INVx2_ASAP7_75t_L g762 ( 
.A(n_702),
.Y(n_762)
);

BUFx10_ASAP7_75t_L g763 ( 
.A(n_734),
.Y(n_763)
);

CKINVDCx5p33_ASAP7_75t_R g764 ( 
.A(n_107),
.Y(n_764)
);

CKINVDCx5p33_ASAP7_75t_R g765 ( 
.A(n_732),
.Y(n_765)
);

CKINVDCx5p33_ASAP7_75t_R g766 ( 
.A(n_496),
.Y(n_766)
);

CKINVDCx20_ASAP7_75t_R g767 ( 
.A(n_670),
.Y(n_767)
);

CKINVDCx5p33_ASAP7_75t_R g768 ( 
.A(n_695),
.Y(n_768)
);

CKINVDCx5p33_ASAP7_75t_R g769 ( 
.A(n_687),
.Y(n_769)
);

CKINVDCx5p33_ASAP7_75t_R g770 ( 
.A(n_696),
.Y(n_770)
);

CKINVDCx20_ASAP7_75t_R g771 ( 
.A(n_216),
.Y(n_771)
);

CKINVDCx14_ASAP7_75t_R g772 ( 
.A(n_333),
.Y(n_772)
);

CKINVDCx5p33_ASAP7_75t_R g773 ( 
.A(n_673),
.Y(n_773)
);

CKINVDCx5p33_ASAP7_75t_R g774 ( 
.A(n_398),
.Y(n_774)
);

CKINVDCx5p33_ASAP7_75t_R g775 ( 
.A(n_627),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_274),
.Y(n_776)
);

CKINVDCx20_ASAP7_75t_R g777 ( 
.A(n_155),
.Y(n_777)
);

CKINVDCx5p33_ASAP7_75t_R g778 ( 
.A(n_660),
.Y(n_778)
);

CKINVDCx5p33_ASAP7_75t_R g779 ( 
.A(n_80),
.Y(n_779)
);

CKINVDCx5p33_ASAP7_75t_R g780 ( 
.A(n_706),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_355),
.Y(n_781)
);

CKINVDCx5p33_ASAP7_75t_R g782 ( 
.A(n_658),
.Y(n_782)
);

INVx2_ASAP7_75t_L g783 ( 
.A(n_203),
.Y(n_783)
);

INVx2_ASAP7_75t_L g784 ( 
.A(n_686),
.Y(n_784)
);

INVx2_ASAP7_75t_L g785 ( 
.A(n_640),
.Y(n_785)
);

INVx1_ASAP7_75t_SL g786 ( 
.A(n_10),
.Y(n_786)
);

BUFx10_ASAP7_75t_L g787 ( 
.A(n_520),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_86),
.Y(n_788)
);

INVx2_ASAP7_75t_L g789 ( 
.A(n_430),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_276),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_432),
.Y(n_791)
);

CKINVDCx5p33_ASAP7_75t_R g792 ( 
.A(n_182),
.Y(n_792)
);

CKINVDCx5p33_ASAP7_75t_R g793 ( 
.A(n_674),
.Y(n_793)
);

CKINVDCx5p33_ASAP7_75t_R g794 ( 
.A(n_165),
.Y(n_794)
);

CKINVDCx5p33_ASAP7_75t_R g795 ( 
.A(n_722),
.Y(n_795)
);

CKINVDCx5p33_ASAP7_75t_R g796 ( 
.A(n_676),
.Y(n_796)
);

CKINVDCx5p33_ASAP7_75t_R g797 ( 
.A(n_544),
.Y(n_797)
);

BUFx3_ASAP7_75t_L g798 ( 
.A(n_547),
.Y(n_798)
);

BUFx10_ASAP7_75t_L g799 ( 
.A(n_744),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_727),
.Y(n_800)
);

CKINVDCx5p33_ASAP7_75t_R g801 ( 
.A(n_291),
.Y(n_801)
);

BUFx10_ASAP7_75t_L g802 ( 
.A(n_724),
.Y(n_802)
);

BUFx2_ASAP7_75t_L g803 ( 
.A(n_654),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_649),
.Y(n_804)
);

CKINVDCx5p33_ASAP7_75t_R g805 ( 
.A(n_667),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_681),
.Y(n_806)
);

CKINVDCx5p33_ASAP7_75t_R g807 ( 
.A(n_321),
.Y(n_807)
);

CKINVDCx5p33_ASAP7_75t_R g808 ( 
.A(n_540),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_566),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_697),
.Y(n_810)
);

CKINVDCx5p33_ASAP7_75t_R g811 ( 
.A(n_128),
.Y(n_811)
);

BUFx6f_ASAP7_75t_L g812 ( 
.A(n_637),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_739),
.Y(n_813)
);

CKINVDCx5p33_ASAP7_75t_R g814 ( 
.A(n_353),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_52),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_684),
.Y(n_816)
);

CKINVDCx5p33_ASAP7_75t_R g817 ( 
.A(n_690),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_67),
.Y(n_818)
);

CKINVDCx5p33_ASAP7_75t_R g819 ( 
.A(n_469),
.Y(n_819)
);

CKINVDCx5p33_ASAP7_75t_R g820 ( 
.A(n_522),
.Y(n_820)
);

CKINVDCx5p33_ASAP7_75t_R g821 ( 
.A(n_244),
.Y(n_821)
);

CKINVDCx5p33_ASAP7_75t_R g822 ( 
.A(n_652),
.Y(n_822)
);

CKINVDCx5p33_ASAP7_75t_R g823 ( 
.A(n_64),
.Y(n_823)
);

INVx2_ASAP7_75t_SL g824 ( 
.A(n_719),
.Y(n_824)
);

CKINVDCx5p33_ASAP7_75t_R g825 ( 
.A(n_71),
.Y(n_825)
);

CKINVDCx5p33_ASAP7_75t_R g826 ( 
.A(n_682),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_645),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_591),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_200),
.Y(n_829)
);

INVxp33_ASAP7_75t_SL g830 ( 
.A(n_502),
.Y(n_830)
);

CKINVDCx5p33_ASAP7_75t_R g831 ( 
.A(n_471),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_211),
.Y(n_832)
);

BUFx2_ASAP7_75t_L g833 ( 
.A(n_151),
.Y(n_833)
);

CKINVDCx5p33_ASAP7_75t_R g834 ( 
.A(n_643),
.Y(n_834)
);

CKINVDCx5p33_ASAP7_75t_R g835 ( 
.A(n_705),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_526),
.Y(n_836)
);

CKINVDCx5p33_ASAP7_75t_R g837 ( 
.A(n_161),
.Y(n_837)
);

INVx1_ASAP7_75t_SL g838 ( 
.A(n_635),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_210),
.Y(n_839)
);

CKINVDCx5p33_ASAP7_75t_R g840 ( 
.A(n_205),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_11),
.Y(n_841)
);

CKINVDCx5p33_ASAP7_75t_R g842 ( 
.A(n_99),
.Y(n_842)
);

CKINVDCx5p33_ASAP7_75t_R g843 ( 
.A(n_608),
.Y(n_843)
);

CKINVDCx5p33_ASAP7_75t_R g844 ( 
.A(n_32),
.Y(n_844)
);

CKINVDCx20_ASAP7_75t_R g845 ( 
.A(n_668),
.Y(n_845)
);

CKINVDCx16_ASAP7_75t_R g846 ( 
.A(n_225),
.Y(n_846)
);

BUFx3_ASAP7_75t_L g847 ( 
.A(n_716),
.Y(n_847)
);

INVx1_ASAP7_75t_L g848 ( 
.A(n_219),
.Y(n_848)
);

CKINVDCx5p33_ASAP7_75t_R g849 ( 
.A(n_504),
.Y(n_849)
);

BUFx10_ASAP7_75t_L g850 ( 
.A(n_616),
.Y(n_850)
);

CKINVDCx5p33_ASAP7_75t_R g851 ( 
.A(n_735),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_694),
.Y(n_852)
);

CKINVDCx5p33_ASAP7_75t_R g853 ( 
.A(n_666),
.Y(n_853)
);

CKINVDCx5p33_ASAP7_75t_R g854 ( 
.A(n_636),
.Y(n_854)
);

INVx2_ASAP7_75t_SL g855 ( 
.A(n_490),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_177),
.Y(n_856)
);

CKINVDCx5p33_ASAP7_75t_R g857 ( 
.A(n_586),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_634),
.Y(n_858)
);

INVx2_ASAP7_75t_L g859 ( 
.A(n_273),
.Y(n_859)
);

CKINVDCx5p33_ASAP7_75t_R g860 ( 
.A(n_641),
.Y(n_860)
);

CKINVDCx20_ASAP7_75t_R g861 ( 
.A(n_462),
.Y(n_861)
);

CKINVDCx5p33_ASAP7_75t_R g862 ( 
.A(n_308),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_100),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_662),
.Y(n_864)
);

CKINVDCx14_ASAP7_75t_R g865 ( 
.A(n_90),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_357),
.Y(n_866)
);

CKINVDCx5p33_ASAP7_75t_R g867 ( 
.A(n_633),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_261),
.Y(n_868)
);

BUFx3_ASAP7_75t_L g869 ( 
.A(n_262),
.Y(n_869)
);

CKINVDCx20_ASAP7_75t_R g870 ( 
.A(n_601),
.Y(n_870)
);

CKINVDCx5p33_ASAP7_75t_R g871 ( 
.A(n_203),
.Y(n_871)
);

CKINVDCx5p33_ASAP7_75t_R g872 ( 
.A(n_335),
.Y(n_872)
);

CKINVDCx5p33_ASAP7_75t_R g873 ( 
.A(n_226),
.Y(n_873)
);

INVx2_ASAP7_75t_L g874 ( 
.A(n_251),
.Y(n_874)
);

CKINVDCx5p33_ASAP7_75t_R g875 ( 
.A(n_659),
.Y(n_875)
);

BUFx5_ASAP7_75t_L g876 ( 
.A(n_495),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_647),
.Y(n_877)
);

CKINVDCx5p33_ASAP7_75t_R g878 ( 
.A(n_653),
.Y(n_878)
);

CKINVDCx5p33_ASAP7_75t_R g879 ( 
.A(n_93),
.Y(n_879)
);

CKINVDCx5p33_ASAP7_75t_R g880 ( 
.A(n_34),
.Y(n_880)
);

INVx1_ASAP7_75t_L g881 ( 
.A(n_478),
.Y(n_881)
);

INVx1_ASAP7_75t_SL g882 ( 
.A(n_709),
.Y(n_882)
);

BUFx2_ASAP7_75t_L g883 ( 
.A(n_717),
.Y(n_883)
);

CKINVDCx5p33_ASAP7_75t_R g884 ( 
.A(n_743),
.Y(n_884)
);

INVx2_ASAP7_75t_L g885 ( 
.A(n_426),
.Y(n_885)
);

CKINVDCx14_ASAP7_75t_R g886 ( 
.A(n_310),
.Y(n_886)
);

CKINVDCx5p33_ASAP7_75t_R g887 ( 
.A(n_703),
.Y(n_887)
);

CKINVDCx5p33_ASAP7_75t_R g888 ( 
.A(n_707),
.Y(n_888)
);

CKINVDCx5p33_ASAP7_75t_R g889 ( 
.A(n_518),
.Y(n_889)
);

CKINVDCx5p33_ASAP7_75t_R g890 ( 
.A(n_114),
.Y(n_890)
);

CKINVDCx5p33_ASAP7_75t_R g891 ( 
.A(n_741),
.Y(n_891)
);

INVx1_ASAP7_75t_L g892 ( 
.A(n_491),
.Y(n_892)
);

CKINVDCx20_ASAP7_75t_R g893 ( 
.A(n_700),
.Y(n_893)
);

INVx1_ASAP7_75t_L g894 ( 
.A(n_699),
.Y(n_894)
);

INVx1_ASAP7_75t_L g895 ( 
.A(n_443),
.Y(n_895)
);

CKINVDCx5p33_ASAP7_75t_R g896 ( 
.A(n_737),
.Y(n_896)
);

INVx1_ASAP7_75t_L g897 ( 
.A(n_740),
.Y(n_897)
);

BUFx5_ASAP7_75t_L g898 ( 
.A(n_312),
.Y(n_898)
);

INVx1_ASAP7_75t_L g899 ( 
.A(n_711),
.Y(n_899)
);

CKINVDCx5p33_ASAP7_75t_R g900 ( 
.A(n_277),
.Y(n_900)
);

CKINVDCx5p33_ASAP7_75t_R g901 ( 
.A(n_255),
.Y(n_901)
);

CKINVDCx5p33_ASAP7_75t_R g902 ( 
.A(n_179),
.Y(n_902)
);

CKINVDCx5p33_ASAP7_75t_R g903 ( 
.A(n_536),
.Y(n_903)
);

INVx1_ASAP7_75t_L g904 ( 
.A(n_117),
.Y(n_904)
);

BUFx3_ASAP7_75t_L g905 ( 
.A(n_338),
.Y(n_905)
);

CKINVDCx5p33_ASAP7_75t_R g906 ( 
.A(n_714),
.Y(n_906)
);

INVx1_ASAP7_75t_SL g907 ( 
.A(n_215),
.Y(n_907)
);

INVx1_ASAP7_75t_SL g908 ( 
.A(n_594),
.Y(n_908)
);

INVx2_ASAP7_75t_L g909 ( 
.A(n_685),
.Y(n_909)
);

INVx2_ASAP7_75t_L g910 ( 
.A(n_427),
.Y(n_910)
);

CKINVDCx5p33_ASAP7_75t_R g911 ( 
.A(n_725),
.Y(n_911)
);

CKINVDCx5p33_ASAP7_75t_R g912 ( 
.A(n_59),
.Y(n_912)
);

INVx1_ASAP7_75t_L g913 ( 
.A(n_609),
.Y(n_913)
);

CKINVDCx5p33_ASAP7_75t_R g914 ( 
.A(n_140),
.Y(n_914)
);

CKINVDCx5p33_ASAP7_75t_R g915 ( 
.A(n_669),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_97),
.Y(n_916)
);

BUFx10_ASAP7_75t_L g917 ( 
.A(n_628),
.Y(n_917)
);

CKINVDCx5p33_ASAP7_75t_R g918 ( 
.A(n_6),
.Y(n_918)
);

HB1xp67_ASAP7_75t_L g919 ( 
.A(n_291),
.Y(n_919)
);

CKINVDCx5p33_ASAP7_75t_R g920 ( 
.A(n_644),
.Y(n_920)
);

CKINVDCx5p33_ASAP7_75t_R g921 ( 
.A(n_738),
.Y(n_921)
);

CKINVDCx5p33_ASAP7_75t_R g922 ( 
.A(n_569),
.Y(n_922)
);

CKINVDCx5p33_ASAP7_75t_R g923 ( 
.A(n_678),
.Y(n_923)
);

CKINVDCx5p33_ASAP7_75t_R g924 ( 
.A(n_688),
.Y(n_924)
);

INVx1_ASAP7_75t_L g925 ( 
.A(n_58),
.Y(n_925)
);

CKINVDCx5p33_ASAP7_75t_R g926 ( 
.A(n_265),
.Y(n_926)
);

INVx1_ASAP7_75t_L g927 ( 
.A(n_529),
.Y(n_927)
);

CKINVDCx5p33_ASAP7_75t_R g928 ( 
.A(n_392),
.Y(n_928)
);

HB1xp67_ASAP7_75t_L g929 ( 
.A(n_638),
.Y(n_929)
);

CKINVDCx5p33_ASAP7_75t_R g930 ( 
.A(n_715),
.Y(n_930)
);

CKINVDCx5p33_ASAP7_75t_R g931 ( 
.A(n_692),
.Y(n_931)
);

INVx1_ASAP7_75t_L g932 ( 
.A(n_425),
.Y(n_932)
);

CKINVDCx5p33_ASAP7_75t_R g933 ( 
.A(n_366),
.Y(n_933)
);

BUFx6f_ASAP7_75t_L g934 ( 
.A(n_708),
.Y(n_934)
);

CKINVDCx5p33_ASAP7_75t_R g935 ( 
.A(n_22),
.Y(n_935)
);

CKINVDCx5p33_ASAP7_75t_R g936 ( 
.A(n_312),
.Y(n_936)
);

CKINVDCx5p33_ASAP7_75t_R g937 ( 
.A(n_726),
.Y(n_937)
);

INVx1_ASAP7_75t_L g938 ( 
.A(n_401),
.Y(n_938)
);

CKINVDCx5p33_ASAP7_75t_R g939 ( 
.A(n_17),
.Y(n_939)
);

CKINVDCx5p33_ASAP7_75t_R g940 ( 
.A(n_657),
.Y(n_940)
);

INVx1_ASAP7_75t_L g941 ( 
.A(n_322),
.Y(n_941)
);

CKINVDCx20_ASAP7_75t_R g942 ( 
.A(n_172),
.Y(n_942)
);

CKINVDCx5p33_ASAP7_75t_R g943 ( 
.A(n_99),
.Y(n_943)
);

CKINVDCx5p33_ASAP7_75t_R g944 ( 
.A(n_97),
.Y(n_944)
);

INVx2_ASAP7_75t_L g945 ( 
.A(n_189),
.Y(n_945)
);

CKINVDCx5p33_ASAP7_75t_R g946 ( 
.A(n_571),
.Y(n_946)
);

CKINVDCx5p33_ASAP7_75t_R g947 ( 
.A(n_679),
.Y(n_947)
);

CKINVDCx5p33_ASAP7_75t_R g948 ( 
.A(n_27),
.Y(n_948)
);

INVx1_ASAP7_75t_SL g949 ( 
.A(n_325),
.Y(n_949)
);

INVx1_ASAP7_75t_L g950 ( 
.A(n_632),
.Y(n_950)
);

CKINVDCx5p33_ASAP7_75t_R g951 ( 
.A(n_481),
.Y(n_951)
);

INVx1_ASAP7_75t_L g952 ( 
.A(n_565),
.Y(n_952)
);

CKINVDCx5p33_ASAP7_75t_R g953 ( 
.A(n_256),
.Y(n_953)
);

INVx1_ASAP7_75t_L g954 ( 
.A(n_671),
.Y(n_954)
);

CKINVDCx5p33_ASAP7_75t_R g955 ( 
.A(n_144),
.Y(n_955)
);

INVx1_ASAP7_75t_L g956 ( 
.A(n_655),
.Y(n_956)
);

INVx1_ASAP7_75t_L g957 ( 
.A(n_639),
.Y(n_957)
);

INVx1_ASAP7_75t_L g958 ( 
.A(n_675),
.Y(n_958)
);

CKINVDCx16_ASAP7_75t_R g959 ( 
.A(n_172),
.Y(n_959)
);

CKINVDCx20_ASAP7_75t_R g960 ( 
.A(n_617),
.Y(n_960)
);

CKINVDCx5p33_ASAP7_75t_R g961 ( 
.A(n_733),
.Y(n_961)
);

CKINVDCx16_ASAP7_75t_R g962 ( 
.A(n_605),
.Y(n_962)
);

INVx1_ASAP7_75t_L g963 ( 
.A(n_720),
.Y(n_963)
);

CKINVDCx5p33_ASAP7_75t_R g964 ( 
.A(n_453),
.Y(n_964)
);

BUFx10_ASAP7_75t_L g965 ( 
.A(n_81),
.Y(n_965)
);

BUFx6f_ASAP7_75t_L g966 ( 
.A(n_650),
.Y(n_966)
);

INVx1_ASAP7_75t_L g967 ( 
.A(n_691),
.Y(n_967)
);

CKINVDCx20_ASAP7_75t_R g968 ( 
.A(n_386),
.Y(n_968)
);

INVx1_ASAP7_75t_L g969 ( 
.A(n_476),
.Y(n_969)
);

CKINVDCx5p33_ASAP7_75t_R g970 ( 
.A(n_197),
.Y(n_970)
);

INVx1_ASAP7_75t_L g971 ( 
.A(n_581),
.Y(n_971)
);

CKINVDCx5p33_ASAP7_75t_R g972 ( 
.A(n_729),
.Y(n_972)
);

CKINVDCx5p33_ASAP7_75t_R g973 ( 
.A(n_29),
.Y(n_973)
);

CKINVDCx5p33_ASAP7_75t_R g974 ( 
.A(n_710),
.Y(n_974)
);

INVx1_ASAP7_75t_L g975 ( 
.A(n_689),
.Y(n_975)
);

CKINVDCx20_ASAP7_75t_R g976 ( 
.A(n_288),
.Y(n_976)
);

INVx1_ASAP7_75t_L g977 ( 
.A(n_175),
.Y(n_977)
);

CKINVDCx5p33_ASAP7_75t_R g978 ( 
.A(n_177),
.Y(n_978)
);

CKINVDCx5p33_ASAP7_75t_R g979 ( 
.A(n_656),
.Y(n_979)
);

CKINVDCx5p33_ASAP7_75t_R g980 ( 
.A(n_100),
.Y(n_980)
);

INVx1_ASAP7_75t_L g981 ( 
.A(n_718),
.Y(n_981)
);

INVx1_ASAP7_75t_L g982 ( 
.A(n_567),
.Y(n_982)
);

CKINVDCx5p33_ASAP7_75t_R g983 ( 
.A(n_175),
.Y(n_983)
);

CKINVDCx5p33_ASAP7_75t_R g984 ( 
.A(n_169),
.Y(n_984)
);

CKINVDCx5p33_ASAP7_75t_R g985 ( 
.A(n_163),
.Y(n_985)
);

CKINVDCx16_ASAP7_75t_R g986 ( 
.A(n_272),
.Y(n_986)
);

BUFx6f_ASAP7_75t_L g987 ( 
.A(n_204),
.Y(n_987)
);

INVx1_ASAP7_75t_L g988 ( 
.A(n_742),
.Y(n_988)
);

INVx1_ASAP7_75t_L g989 ( 
.A(n_429),
.Y(n_989)
);

INVx1_ASAP7_75t_L g990 ( 
.A(n_219),
.Y(n_990)
);

CKINVDCx20_ASAP7_75t_R g991 ( 
.A(n_712),
.Y(n_991)
);

CKINVDCx5p33_ASAP7_75t_R g992 ( 
.A(n_389),
.Y(n_992)
);

CKINVDCx5p33_ASAP7_75t_R g993 ( 
.A(n_736),
.Y(n_993)
);

CKINVDCx5p33_ASAP7_75t_R g994 ( 
.A(n_721),
.Y(n_994)
);

INVx1_ASAP7_75t_L g995 ( 
.A(n_302),
.Y(n_995)
);

CKINVDCx5p33_ASAP7_75t_R g996 ( 
.A(n_135),
.Y(n_996)
);

CKINVDCx5p33_ASAP7_75t_R g997 ( 
.A(n_646),
.Y(n_997)
);

CKINVDCx5p33_ASAP7_75t_R g998 ( 
.A(n_465),
.Y(n_998)
);

CKINVDCx5p33_ASAP7_75t_R g999 ( 
.A(n_210),
.Y(n_999)
);

BUFx2_ASAP7_75t_L g1000 ( 
.A(n_538),
.Y(n_1000)
);

HB1xp67_ASAP7_75t_L g1001 ( 
.A(n_231),
.Y(n_1001)
);

BUFx3_ASAP7_75t_L g1002 ( 
.A(n_661),
.Y(n_1002)
);

INVx1_ASAP7_75t_L g1003 ( 
.A(n_713),
.Y(n_1003)
);

CKINVDCx5p33_ASAP7_75t_R g1004 ( 
.A(n_112),
.Y(n_1004)
);

CKINVDCx5p33_ASAP7_75t_R g1005 ( 
.A(n_365),
.Y(n_1005)
);

BUFx3_ASAP7_75t_L g1006 ( 
.A(n_36),
.Y(n_1006)
);

INVx1_ASAP7_75t_L g1007 ( 
.A(n_440),
.Y(n_1007)
);

INVx1_ASAP7_75t_L g1008 ( 
.A(n_16),
.Y(n_1008)
);

CKINVDCx5p33_ASAP7_75t_R g1009 ( 
.A(n_648),
.Y(n_1009)
);

INVx2_ASAP7_75t_L g1010 ( 
.A(n_474),
.Y(n_1010)
);

CKINVDCx5p33_ASAP7_75t_R g1011 ( 
.A(n_344),
.Y(n_1011)
);

INVx2_ASAP7_75t_L g1012 ( 
.A(n_642),
.Y(n_1012)
);

CKINVDCx16_ASAP7_75t_R g1013 ( 
.A(n_209),
.Y(n_1013)
);

CKINVDCx5p33_ASAP7_75t_R g1014 ( 
.A(n_231),
.Y(n_1014)
);

BUFx6f_ASAP7_75t_L g1015 ( 
.A(n_514),
.Y(n_1015)
);

BUFx2_ASAP7_75t_L g1016 ( 
.A(n_45),
.Y(n_1016)
);

CKINVDCx5p33_ASAP7_75t_R g1017 ( 
.A(n_300),
.Y(n_1017)
);

INVxp67_ASAP7_75t_L g1018 ( 
.A(n_378),
.Y(n_1018)
);

CKINVDCx5p33_ASAP7_75t_R g1019 ( 
.A(n_698),
.Y(n_1019)
);

CKINVDCx5p33_ASAP7_75t_R g1020 ( 
.A(n_747),
.Y(n_1020)
);

CKINVDCx5p33_ASAP7_75t_R g1021 ( 
.A(n_672),
.Y(n_1021)
);

INVx1_ASAP7_75t_L g1022 ( 
.A(n_533),
.Y(n_1022)
);

INVx1_ASAP7_75t_L g1023 ( 
.A(n_651),
.Y(n_1023)
);

CKINVDCx5p33_ASAP7_75t_R g1024 ( 
.A(n_693),
.Y(n_1024)
);

CKINVDCx5p33_ASAP7_75t_R g1025 ( 
.A(n_294),
.Y(n_1025)
);

CKINVDCx5p33_ASAP7_75t_R g1026 ( 
.A(n_62),
.Y(n_1026)
);

CKINVDCx20_ASAP7_75t_R g1027 ( 
.A(n_0),
.Y(n_1027)
);

CKINVDCx5p33_ASAP7_75t_R g1028 ( 
.A(n_267),
.Y(n_1028)
);

INVx3_ASAP7_75t_L g1029 ( 
.A(n_677),
.Y(n_1029)
);

CKINVDCx5p33_ASAP7_75t_R g1030 ( 
.A(n_227),
.Y(n_1030)
);

CKINVDCx5p33_ASAP7_75t_R g1031 ( 
.A(n_723),
.Y(n_1031)
);

INVx1_ASAP7_75t_L g1032 ( 
.A(n_483),
.Y(n_1032)
);

CKINVDCx5p33_ASAP7_75t_R g1033 ( 
.A(n_489),
.Y(n_1033)
);

INVx1_ASAP7_75t_L g1034 ( 
.A(n_294),
.Y(n_1034)
);

CKINVDCx5p33_ASAP7_75t_R g1035 ( 
.A(n_55),
.Y(n_1035)
);

CKINVDCx5p33_ASAP7_75t_R g1036 ( 
.A(n_151),
.Y(n_1036)
);

INVx1_ASAP7_75t_L g1037 ( 
.A(n_683),
.Y(n_1037)
);

CKINVDCx5p33_ASAP7_75t_R g1038 ( 
.A(n_704),
.Y(n_1038)
);

INVx2_ASAP7_75t_L g1039 ( 
.A(n_324),
.Y(n_1039)
);

INVx1_ASAP7_75t_L g1040 ( 
.A(n_54),
.Y(n_1040)
);

CKINVDCx5p33_ASAP7_75t_R g1041 ( 
.A(n_593),
.Y(n_1041)
);

INVx1_ASAP7_75t_L g1042 ( 
.A(n_446),
.Y(n_1042)
);

INVx1_ASAP7_75t_L g1043 ( 
.A(n_259),
.Y(n_1043)
);

CKINVDCx5p33_ASAP7_75t_R g1044 ( 
.A(n_367),
.Y(n_1044)
);

BUFx10_ASAP7_75t_L g1045 ( 
.A(n_56),
.Y(n_1045)
);

INVx1_ASAP7_75t_L g1046 ( 
.A(n_319),
.Y(n_1046)
);

CKINVDCx5p33_ASAP7_75t_R g1047 ( 
.A(n_198),
.Y(n_1047)
);

CKINVDCx5p33_ASAP7_75t_R g1048 ( 
.A(n_324),
.Y(n_1048)
);

CKINVDCx5p33_ASAP7_75t_R g1049 ( 
.A(n_20),
.Y(n_1049)
);

CKINVDCx5p33_ASAP7_75t_R g1050 ( 
.A(n_701),
.Y(n_1050)
);

INVx1_ASAP7_75t_SL g1051 ( 
.A(n_373),
.Y(n_1051)
);

INVx1_ASAP7_75t_SL g1052 ( 
.A(n_463),
.Y(n_1052)
);

CKINVDCx20_ASAP7_75t_R g1053 ( 
.A(n_508),
.Y(n_1053)
);

INVx1_ASAP7_75t_L g1054 ( 
.A(n_730),
.Y(n_1054)
);

CKINVDCx5p33_ASAP7_75t_R g1055 ( 
.A(n_503),
.Y(n_1055)
);

INVx1_ASAP7_75t_L g1056 ( 
.A(n_345),
.Y(n_1056)
);

INVx1_ASAP7_75t_L g1057 ( 
.A(n_680),
.Y(n_1057)
);

BUFx10_ASAP7_75t_L g1058 ( 
.A(n_55),
.Y(n_1058)
);

CKINVDCx5p33_ASAP7_75t_R g1059 ( 
.A(n_448),
.Y(n_1059)
);

INVx1_ASAP7_75t_L g1060 ( 
.A(n_137),
.Y(n_1060)
);

CKINVDCx20_ASAP7_75t_R g1061 ( 
.A(n_93),
.Y(n_1061)
);

CKINVDCx5p33_ASAP7_75t_R g1062 ( 
.A(n_220),
.Y(n_1062)
);

CKINVDCx5p33_ASAP7_75t_R g1063 ( 
.A(n_728),
.Y(n_1063)
);

CKINVDCx5p33_ASAP7_75t_R g1064 ( 
.A(n_265),
.Y(n_1064)
);

INVx1_ASAP7_75t_L g1065 ( 
.A(n_117),
.Y(n_1065)
);

CKINVDCx5p33_ASAP7_75t_R g1066 ( 
.A(n_745),
.Y(n_1066)
);

CKINVDCx5p33_ASAP7_75t_R g1067 ( 
.A(n_665),
.Y(n_1067)
);

INVx4_ASAP7_75t_L g1068 ( 
.A(n_1029),
.Y(n_1068)
);

BUFx12f_ASAP7_75t_L g1069 ( 
.A(n_763),
.Y(n_1069)
);

NOR2xp33_ASAP7_75t_L g1070 ( 
.A(n_754),
.B(n_1),
.Y(n_1070)
);

AND2x6_ASAP7_75t_L g1071 ( 
.A(n_757),
.B(n_358),
.Y(n_1071)
);

INVx2_ASAP7_75t_L g1072 ( 
.A(n_898),
.Y(n_1072)
);

INVx5_ASAP7_75t_L g1073 ( 
.A(n_763),
.Y(n_1073)
);

INVx1_ASAP7_75t_L g1074 ( 
.A(n_898),
.Y(n_1074)
);

NAND2xp5_ASAP7_75t_L g1075 ( 
.A(n_803),
.B(n_0),
.Y(n_1075)
);

INVx1_ASAP7_75t_L g1076 ( 
.A(n_898),
.Y(n_1076)
);

NAND2xp5_ASAP7_75t_SL g1077 ( 
.A(n_846),
.B(n_1),
.Y(n_1077)
);

BUFx6f_ASAP7_75t_L g1078 ( 
.A(n_987),
.Y(n_1078)
);

INVx5_ASAP7_75t_L g1079 ( 
.A(n_787),
.Y(n_1079)
);

INVx2_ASAP7_75t_L g1080 ( 
.A(n_898),
.Y(n_1080)
);

BUFx6f_ASAP7_75t_L g1081 ( 
.A(n_987),
.Y(n_1081)
);

NAND2xp5_ASAP7_75t_L g1082 ( 
.A(n_883),
.B(n_2),
.Y(n_1082)
);

BUFx12f_ASAP7_75t_L g1083 ( 
.A(n_787),
.Y(n_1083)
);

BUFx12f_ASAP7_75t_L g1084 ( 
.A(n_799),
.Y(n_1084)
);

BUFx6f_ASAP7_75t_L g1085 ( 
.A(n_987),
.Y(n_1085)
);

INVx5_ASAP7_75t_L g1086 ( 
.A(n_799),
.Y(n_1086)
);

NAND2xp5_ASAP7_75t_L g1087 ( 
.A(n_1000),
.B(n_2),
.Y(n_1087)
);

INVx2_ASAP7_75t_SL g1088 ( 
.A(n_965),
.Y(n_1088)
);

BUFx6f_ASAP7_75t_L g1089 ( 
.A(n_812),
.Y(n_1089)
);

NOR2x1_ASAP7_75t_L g1090 ( 
.A(n_798),
.B(n_359),
.Y(n_1090)
);

BUFx6f_ASAP7_75t_L g1091 ( 
.A(n_812),
.Y(n_1091)
);

BUFx3_ASAP7_75t_L g1092 ( 
.A(n_802),
.Y(n_1092)
);

NAND2xp5_ASAP7_75t_SL g1093 ( 
.A(n_959),
.B(n_3),
.Y(n_1093)
);

BUFx6f_ASAP7_75t_L g1094 ( 
.A(n_812),
.Y(n_1094)
);

NAND2xp5_ASAP7_75t_L g1095 ( 
.A(n_929),
.B(n_3),
.Y(n_1095)
);

AND2x2_ASAP7_75t_L g1096 ( 
.A(n_772),
.B(n_4),
.Y(n_1096)
);

AND2x4_ASAP7_75t_L g1097 ( 
.A(n_833),
.B(n_4),
.Y(n_1097)
);

BUFx6f_ASAP7_75t_L g1098 ( 
.A(n_934),
.Y(n_1098)
);

INVx2_ASAP7_75t_L g1099 ( 
.A(n_898),
.Y(n_1099)
);

AND2x2_ASAP7_75t_L g1100 ( 
.A(n_865),
.B(n_5),
.Y(n_1100)
);

NAND2xp5_ASAP7_75t_L g1101 ( 
.A(n_759),
.B(n_5),
.Y(n_1101)
);

NAND2xp5_ASAP7_75t_L g1102 ( 
.A(n_791),
.B(n_6),
.Y(n_1102)
);

NOR2xp33_ASAP7_75t_SL g1103 ( 
.A(n_962),
.B(n_360),
.Y(n_1103)
);

BUFx6f_ASAP7_75t_L g1104 ( 
.A(n_934),
.Y(n_1104)
);

HB1xp67_ASAP7_75t_L g1105 ( 
.A(n_919),
.Y(n_1105)
);

INVx1_ASAP7_75t_L g1106 ( 
.A(n_750),
.Y(n_1106)
);

AND2x4_ASAP7_75t_L g1107 ( 
.A(n_1016),
.B(n_7),
.Y(n_1107)
);

AND2x2_ASAP7_75t_L g1108 ( 
.A(n_886),
.B(n_7),
.Y(n_1108)
);

NOR2xp33_ASAP7_75t_L g1109 ( 
.A(n_986),
.B(n_1013),
.Y(n_1109)
);

HB1xp67_ASAP7_75t_L g1110 ( 
.A(n_1001),
.Y(n_1110)
);

NAND2xp5_ASAP7_75t_L g1111 ( 
.A(n_800),
.B(n_8),
.Y(n_1111)
);

NAND2xp5_ASAP7_75t_L g1112 ( 
.A(n_804),
.B(n_806),
.Y(n_1112)
);

AND2x2_ASAP7_75t_L g1113 ( 
.A(n_965),
.B(n_8),
.Y(n_1113)
);

INVx1_ASAP7_75t_L g1114 ( 
.A(n_756),
.Y(n_1114)
);

AND2x4_ASAP7_75t_L g1115 ( 
.A(n_869),
.B(n_9),
.Y(n_1115)
);

AND2x2_ASAP7_75t_L g1116 ( 
.A(n_1073),
.B(n_802),
.Y(n_1116)
);

AOI22xp5_ASAP7_75t_L g1117 ( 
.A1(n_1109),
.A2(n_976),
.B1(n_771),
.B2(n_942),
.Y(n_1117)
);

AND2x4_ASAP7_75t_L g1118 ( 
.A(n_1092),
.B(n_905),
.Y(n_1118)
);

AO22x2_ASAP7_75t_L g1119 ( 
.A1(n_1077),
.A2(n_786),
.B1(n_949),
.B2(n_907),
.Y(n_1119)
);

INVx3_ASAP7_75t_L g1120 ( 
.A(n_1078),
.Y(n_1120)
);

AOI22xp5_ASAP7_75t_L g1121 ( 
.A1(n_1096),
.A2(n_1061),
.B1(n_777),
.B2(n_1027),
.Y(n_1121)
);

AOI22xp5_ASAP7_75t_L g1122 ( 
.A1(n_1100),
.A2(n_845),
.B1(n_861),
.B2(n_767),
.Y(n_1122)
);

NOR2xp33_ASAP7_75t_L g1123 ( 
.A(n_1068),
.B(n_830),
.Y(n_1123)
);

OAI22xp33_ASAP7_75t_L g1124 ( 
.A1(n_1103),
.A2(n_752),
.B1(n_893),
.B2(n_870),
.Y(n_1124)
);

AOI22xp5_ASAP7_75t_L g1125 ( 
.A1(n_1108),
.A2(n_968),
.B1(n_991),
.B2(n_960),
.Y(n_1125)
);

NAND2xp5_ASAP7_75t_L g1126 ( 
.A(n_1073),
.B(n_809),
.Y(n_1126)
);

INVx2_ASAP7_75t_L g1127 ( 
.A(n_1078),
.Y(n_1127)
);

NAND2xp5_ASAP7_75t_SL g1128 ( 
.A(n_1079),
.B(n_850),
.Y(n_1128)
);

OR2x2_ASAP7_75t_L g1129 ( 
.A(n_1105),
.B(n_776),
.Y(n_1129)
);

INVx1_ASAP7_75t_L g1130 ( 
.A(n_1074),
.Y(n_1130)
);

INVx3_ASAP7_75t_L g1131 ( 
.A(n_1081),
.Y(n_1131)
);

AND2x2_ASAP7_75t_L g1132 ( 
.A(n_1079),
.B(n_850),
.Y(n_1132)
);

OAI22xp33_ASAP7_75t_L g1133 ( 
.A1(n_1110),
.A2(n_1053),
.B1(n_1006),
.B2(n_1062),
.Y(n_1133)
);

AO22x2_ASAP7_75t_L g1134 ( 
.A1(n_1093),
.A2(n_788),
.B1(n_790),
.B2(n_781),
.Y(n_1134)
);

OAI22xp33_ASAP7_75t_L g1135 ( 
.A1(n_1095),
.A2(n_760),
.B1(n_764),
.B2(n_749),
.Y(n_1135)
);

AO22x2_ASAP7_75t_L g1136 ( 
.A1(n_1113),
.A2(n_818),
.B1(n_829),
.B2(n_815),
.Y(n_1136)
);

CKINVDCx16_ASAP7_75t_R g1137 ( 
.A(n_1069),
.Y(n_1137)
);

INVx1_ASAP7_75t_L g1138 ( 
.A(n_1076),
.Y(n_1138)
);

AOI22xp5_ASAP7_75t_L g1139 ( 
.A1(n_1070),
.A2(n_792),
.B1(n_1011),
.B2(n_807),
.Y(n_1139)
);

XNOR2xp5_ASAP7_75t_SL g1140 ( 
.A(n_1083),
.B(n_751),
.Y(n_1140)
);

INVx1_ASAP7_75t_L g1141 ( 
.A(n_1072),
.Y(n_1141)
);

AOI22xp5_ASAP7_75t_L g1142 ( 
.A1(n_1075),
.A2(n_779),
.B1(n_811),
.B2(n_794),
.Y(n_1142)
);

AND2x2_ASAP7_75t_L g1143 ( 
.A(n_1086),
.B(n_917),
.Y(n_1143)
);

AOI22xp5_ASAP7_75t_L g1144 ( 
.A1(n_1082),
.A2(n_1087),
.B1(n_1088),
.B2(n_1097),
.Y(n_1144)
);

OAI22xp33_ASAP7_75t_L g1145 ( 
.A1(n_1086),
.A2(n_1064),
.B1(n_814),
.B2(n_821),
.Y(n_1145)
);

AO22x2_ASAP7_75t_L g1146 ( 
.A1(n_1107),
.A2(n_839),
.B1(n_841),
.B2(n_832),
.Y(n_1146)
);

INVx1_ASAP7_75t_SL g1147 ( 
.A(n_1084),
.Y(n_1147)
);

BUFx6f_ASAP7_75t_L g1148 ( 
.A(n_1089),
.Y(n_1148)
);

AND2x2_ASAP7_75t_L g1149 ( 
.A(n_1106),
.B(n_917),
.Y(n_1149)
);

OAI22xp33_ASAP7_75t_SL g1150 ( 
.A1(n_1112),
.A2(n_823),
.B1(n_825),
.B2(n_801),
.Y(n_1150)
);

AO22x2_ASAP7_75t_L g1151 ( 
.A1(n_1115),
.A2(n_1102),
.B1(n_1111),
.B2(n_1101),
.Y(n_1151)
);

OAI22xp33_ASAP7_75t_L g1152 ( 
.A1(n_1114),
.A2(n_840),
.B1(n_842),
.B2(n_837),
.Y(n_1152)
);

XNOR2xp5_ASAP7_75t_L g1153 ( 
.A(n_1124),
.B(n_1090),
.Y(n_1153)
);

INVx2_ASAP7_75t_SL g1154 ( 
.A(n_1116),
.Y(n_1154)
);

NOR2xp33_ASAP7_75t_L g1155 ( 
.A(n_1123),
.B(n_1080),
.Y(n_1155)
);

INVx2_ASAP7_75t_L g1156 ( 
.A(n_1141),
.Y(n_1156)
);

NOR2xp33_ASAP7_75t_L g1157 ( 
.A(n_1130),
.B(n_1099),
.Y(n_1157)
);

INVx1_ASAP7_75t_L g1158 ( 
.A(n_1138),
.Y(n_1158)
);

INVx1_ASAP7_75t_L g1159 ( 
.A(n_1149),
.Y(n_1159)
);

INVxp67_ASAP7_75t_L g1160 ( 
.A(n_1132),
.Y(n_1160)
);

INVx2_ASAP7_75t_L g1161 ( 
.A(n_1127),
.Y(n_1161)
);

NAND2x1p5_ASAP7_75t_L g1162 ( 
.A(n_1147),
.B(n_1081),
.Y(n_1162)
);

NAND2xp5_ASAP7_75t_L g1163 ( 
.A(n_1143),
.B(n_1071),
.Y(n_1163)
);

BUFx6f_ASAP7_75t_SL g1164 ( 
.A(n_1118),
.Y(n_1164)
);

AND2x2_ASAP7_75t_L g1165 ( 
.A(n_1137),
.B(n_1129),
.Y(n_1165)
);

INVx1_ASAP7_75t_L g1166 ( 
.A(n_1120),
.Y(n_1166)
);

CKINVDCx20_ASAP7_75t_R g1167 ( 
.A(n_1122),
.Y(n_1167)
);

AND2x2_ASAP7_75t_L g1168 ( 
.A(n_1125),
.B(n_1045),
.Y(n_1168)
);

INVx1_ASAP7_75t_L g1169 ( 
.A(n_1131),
.Y(n_1169)
);

NOR2xp33_ASAP7_75t_L g1170 ( 
.A(n_1139),
.B(n_1085),
.Y(n_1170)
);

NOR2xp67_ASAP7_75t_L g1171 ( 
.A(n_1126),
.B(n_1029),
.Y(n_1171)
);

INVx1_ASAP7_75t_L g1172 ( 
.A(n_1148),
.Y(n_1172)
);

INVx1_ASAP7_75t_L g1173 ( 
.A(n_1148),
.Y(n_1173)
);

INVx1_ASAP7_75t_L g1174 ( 
.A(n_1134),
.Y(n_1174)
);

INVx1_ASAP7_75t_L g1175 ( 
.A(n_1136),
.Y(n_1175)
);

INVx1_ASAP7_75t_L g1176 ( 
.A(n_1146),
.Y(n_1176)
);

AND2x4_ASAP7_75t_L g1177 ( 
.A(n_1128),
.B(n_1071),
.Y(n_1177)
);

INVx1_ASAP7_75t_L g1178 ( 
.A(n_1151),
.Y(n_1178)
);

INVx1_ASAP7_75t_L g1179 ( 
.A(n_1144),
.Y(n_1179)
);

INVx1_ASAP7_75t_L g1180 ( 
.A(n_1119),
.Y(n_1180)
);

AND2x6_ASAP7_75t_L g1181 ( 
.A(n_1142),
.B(n_810),
.Y(n_1181)
);

NOR2xp33_ASAP7_75t_L g1182 ( 
.A(n_1145),
.B(n_1085),
.Y(n_1182)
);

INVx1_ASAP7_75t_L g1183 ( 
.A(n_1152),
.Y(n_1183)
);

INVx1_ASAP7_75t_L g1184 ( 
.A(n_1150),
.Y(n_1184)
);

CKINVDCx20_ASAP7_75t_R g1185 ( 
.A(n_1117),
.Y(n_1185)
);

AND2x4_ASAP7_75t_L g1186 ( 
.A(n_1121),
.B(n_848),
.Y(n_1186)
);

INVxp67_ASAP7_75t_SL g1187 ( 
.A(n_1133),
.Y(n_1187)
);

INVx1_ASAP7_75t_L g1188 ( 
.A(n_1135),
.Y(n_1188)
);

OR2x2_ASAP7_75t_L g1189 ( 
.A(n_1140),
.B(n_977),
.Y(n_1189)
);

INVx1_ASAP7_75t_L g1190 ( 
.A(n_1130),
.Y(n_1190)
);

INVxp67_ASAP7_75t_SL g1191 ( 
.A(n_1130),
.Y(n_1191)
);

NAND2xp33_ASAP7_75t_R g1192 ( 
.A(n_1149),
.B(n_844),
.Y(n_1192)
);

INVx1_ASAP7_75t_L g1193 ( 
.A(n_1130),
.Y(n_1193)
);

INVx1_ASAP7_75t_L g1194 ( 
.A(n_1130),
.Y(n_1194)
);

INVx2_ASAP7_75t_SL g1195 ( 
.A(n_1116),
.Y(n_1195)
);

CKINVDCx20_ASAP7_75t_R g1196 ( 
.A(n_1137),
.Y(n_1196)
);

INVx1_ASAP7_75t_L g1197 ( 
.A(n_1130),
.Y(n_1197)
);

INVx1_ASAP7_75t_L g1198 ( 
.A(n_1130),
.Y(n_1198)
);

INVx2_ASAP7_75t_L g1199 ( 
.A(n_1141),
.Y(n_1199)
);

INVx1_ASAP7_75t_L g1200 ( 
.A(n_1130),
.Y(n_1200)
);

CKINVDCx20_ASAP7_75t_R g1201 ( 
.A(n_1137),
.Y(n_1201)
);

INVxp67_ASAP7_75t_L g1202 ( 
.A(n_1149),
.Y(n_1202)
);

INVx1_ASAP7_75t_L g1203 ( 
.A(n_1130),
.Y(n_1203)
);

AND2x2_ASAP7_75t_L g1204 ( 
.A(n_1149),
.B(n_1045),
.Y(n_1204)
);

XOR2xp5_ASAP7_75t_L g1205 ( 
.A(n_1140),
.B(n_862),
.Y(n_1205)
);

INVx2_ASAP7_75t_L g1206 ( 
.A(n_1141),
.Y(n_1206)
);

NAND2xp5_ASAP7_75t_L g1207 ( 
.A(n_1155),
.B(n_753),
.Y(n_1207)
);

INVx2_ASAP7_75t_L g1208 ( 
.A(n_1156),
.Y(n_1208)
);

HB1xp67_ASAP7_75t_L g1209 ( 
.A(n_1165),
.Y(n_1209)
);

BUFx6f_ASAP7_75t_L g1210 ( 
.A(n_1162),
.Y(n_1210)
);

AND2x4_ASAP7_75t_L g1211 ( 
.A(n_1196),
.B(n_856),
.Y(n_1211)
);

INVx1_ASAP7_75t_L g1212 ( 
.A(n_1158),
.Y(n_1212)
);

INVx2_ASAP7_75t_L g1213 ( 
.A(n_1199),
.Y(n_1213)
);

HB1xp67_ASAP7_75t_L g1214 ( 
.A(n_1204),
.Y(n_1214)
);

AND2x2_ASAP7_75t_L g1215 ( 
.A(n_1202),
.B(n_1168),
.Y(n_1215)
);

INVxp67_ASAP7_75t_L g1216 ( 
.A(n_1192),
.Y(n_1216)
);

INVx1_ASAP7_75t_L g1217 ( 
.A(n_1190),
.Y(n_1217)
);

INVx1_ASAP7_75t_L g1218 ( 
.A(n_1193),
.Y(n_1218)
);

AND2x4_ASAP7_75t_SL g1219 ( 
.A(n_1201),
.B(n_1058),
.Y(n_1219)
);

NAND2xp5_ASAP7_75t_L g1220 ( 
.A(n_1191),
.B(n_838),
.Y(n_1220)
);

AND2x2_ASAP7_75t_L g1221 ( 
.A(n_1187),
.B(n_1058),
.Y(n_1221)
);

INVx2_ASAP7_75t_SL g1222 ( 
.A(n_1154),
.Y(n_1222)
);

INVx1_ASAP7_75t_L g1223 ( 
.A(n_1194),
.Y(n_1223)
);

AND2x2_ASAP7_75t_L g1224 ( 
.A(n_1159),
.B(n_863),
.Y(n_1224)
);

AND2x6_ASAP7_75t_L g1225 ( 
.A(n_1179),
.B(n_1177),
.Y(n_1225)
);

INVx1_ASAP7_75t_L g1226 ( 
.A(n_1197),
.Y(n_1226)
);

HB1xp67_ASAP7_75t_L g1227 ( 
.A(n_1164),
.Y(n_1227)
);

INVx2_ASAP7_75t_L g1228 ( 
.A(n_1206),
.Y(n_1228)
);

OR2x2_ASAP7_75t_SL g1229 ( 
.A(n_1183),
.B(n_783),
.Y(n_1229)
);

AND2x2_ASAP7_75t_L g1230 ( 
.A(n_1186),
.B(n_866),
.Y(n_1230)
);

INVx3_ASAP7_75t_L g1231 ( 
.A(n_1161),
.Y(n_1231)
);

AND2x2_ASAP7_75t_L g1232 ( 
.A(n_1160),
.B(n_868),
.Y(n_1232)
);

NAND2xp5_ASAP7_75t_L g1233 ( 
.A(n_1188),
.B(n_882),
.Y(n_1233)
);

INVx2_ASAP7_75t_L g1234 ( 
.A(n_1198),
.Y(n_1234)
);

BUFx3_ASAP7_75t_L g1235 ( 
.A(n_1172),
.Y(n_1235)
);

NAND2xp5_ASAP7_75t_L g1236 ( 
.A(n_1200),
.B(n_1203),
.Y(n_1236)
);

INVx2_ASAP7_75t_SL g1237 ( 
.A(n_1195),
.Y(n_1237)
);

AND2x2_ASAP7_75t_L g1238 ( 
.A(n_1170),
.B(n_904),
.Y(n_1238)
);

INVxp67_ASAP7_75t_SL g1239 ( 
.A(n_1182),
.Y(n_1239)
);

INVx1_ASAP7_75t_L g1240 ( 
.A(n_1157),
.Y(n_1240)
);

NAND2xp5_ASAP7_75t_L g1241 ( 
.A(n_1153),
.B(n_908),
.Y(n_1241)
);

INVx1_ASAP7_75t_L g1242 ( 
.A(n_1166),
.Y(n_1242)
);

INVx1_ASAP7_75t_L g1243 ( 
.A(n_1169),
.Y(n_1243)
);

OAI21xp5_ASAP7_75t_L g1244 ( 
.A1(n_1163),
.A2(n_1018),
.B(n_816),
.Y(n_1244)
);

NAND2xp5_ASAP7_75t_L g1245 ( 
.A(n_1181),
.B(n_1051),
.Y(n_1245)
);

AND2x4_ASAP7_75t_L g1246 ( 
.A(n_1176),
.B(n_916),
.Y(n_1246)
);

AND2x2_ASAP7_75t_L g1247 ( 
.A(n_1175),
.B(n_1174),
.Y(n_1247)
);

INVx1_ASAP7_75t_L g1248 ( 
.A(n_1173),
.Y(n_1248)
);

NAND2xp5_ASAP7_75t_L g1249 ( 
.A(n_1181),
.B(n_1052),
.Y(n_1249)
);

INVxp67_ASAP7_75t_SL g1250 ( 
.A(n_1178),
.Y(n_1250)
);

INVx1_ASAP7_75t_L g1251 ( 
.A(n_1184),
.Y(n_1251)
);

INVx1_ASAP7_75t_L g1252 ( 
.A(n_1180),
.Y(n_1252)
);

INVx2_ASAP7_75t_L g1253 ( 
.A(n_1181),
.Y(n_1253)
);

INVx2_ASAP7_75t_SL g1254 ( 
.A(n_1189),
.Y(n_1254)
);

NAND2xp5_ASAP7_75t_SL g1255 ( 
.A(n_1171),
.B(n_871),
.Y(n_1255)
);

INVx1_ASAP7_75t_L g1256 ( 
.A(n_1167),
.Y(n_1256)
);

INVx2_ASAP7_75t_SL g1257 ( 
.A(n_1185),
.Y(n_1257)
);

INVx1_ASAP7_75t_L g1258 ( 
.A(n_1205),
.Y(n_1258)
);

NAND2xp5_ASAP7_75t_L g1259 ( 
.A(n_1155),
.B(n_872),
.Y(n_1259)
);

INVx2_ASAP7_75t_L g1260 ( 
.A(n_1156),
.Y(n_1260)
);

INVx3_ASAP7_75t_SL g1261 ( 
.A(n_1196),
.Y(n_1261)
);

NAND2xp5_ASAP7_75t_L g1262 ( 
.A(n_1155),
.B(n_873),
.Y(n_1262)
);

BUFx6f_ASAP7_75t_L g1263 ( 
.A(n_1162),
.Y(n_1263)
);

AND2x2_ASAP7_75t_L g1264 ( 
.A(n_1204),
.B(n_925),
.Y(n_1264)
);

INVx1_ASAP7_75t_L g1265 ( 
.A(n_1158),
.Y(n_1265)
);

INVx1_ASAP7_75t_L g1266 ( 
.A(n_1158),
.Y(n_1266)
);

INVx1_ASAP7_75t_L g1267 ( 
.A(n_1158),
.Y(n_1267)
);

INVx1_ASAP7_75t_L g1268 ( 
.A(n_1158),
.Y(n_1268)
);

BUFx3_ASAP7_75t_L g1269 ( 
.A(n_1196),
.Y(n_1269)
);

INVx2_ASAP7_75t_L g1270 ( 
.A(n_1156),
.Y(n_1270)
);

AND2x2_ASAP7_75t_L g1271 ( 
.A(n_1204),
.B(n_941),
.Y(n_1271)
);

BUFx6f_ASAP7_75t_L g1272 ( 
.A(n_1162),
.Y(n_1272)
);

INVx1_ASAP7_75t_L g1273 ( 
.A(n_1158),
.Y(n_1273)
);

INVx2_ASAP7_75t_L g1274 ( 
.A(n_1156),
.Y(n_1274)
);

BUFx6f_ASAP7_75t_L g1275 ( 
.A(n_1162),
.Y(n_1275)
);

AND2x6_ASAP7_75t_L g1276 ( 
.A(n_1204),
.B(n_813),
.Y(n_1276)
);

AND2x2_ASAP7_75t_L g1277 ( 
.A(n_1204),
.B(n_990),
.Y(n_1277)
);

AND2x2_ASAP7_75t_L g1278 ( 
.A(n_1204),
.B(n_995),
.Y(n_1278)
);

AND2x2_ASAP7_75t_L g1279 ( 
.A(n_1204),
.B(n_1008),
.Y(n_1279)
);

INVx1_ASAP7_75t_L g1280 ( 
.A(n_1158),
.Y(n_1280)
);

AND2x2_ASAP7_75t_L g1281 ( 
.A(n_1204),
.B(n_1034),
.Y(n_1281)
);

INVx2_ASAP7_75t_L g1282 ( 
.A(n_1156),
.Y(n_1282)
);

INVx3_ASAP7_75t_L g1283 ( 
.A(n_1164),
.Y(n_1283)
);

HB1xp67_ASAP7_75t_L g1284 ( 
.A(n_1165),
.Y(n_1284)
);

INVx4_ASAP7_75t_L g1285 ( 
.A(n_1164),
.Y(n_1285)
);

NAND2xp5_ASAP7_75t_L g1286 ( 
.A(n_1155),
.B(n_879),
.Y(n_1286)
);

BUFx6f_ASAP7_75t_L g1287 ( 
.A(n_1162),
.Y(n_1287)
);

AND2x4_ASAP7_75t_L g1288 ( 
.A(n_1196),
.B(n_1040),
.Y(n_1288)
);

AND2x2_ASAP7_75t_L g1289 ( 
.A(n_1204),
.B(n_1043),
.Y(n_1289)
);

INVx1_ASAP7_75t_L g1290 ( 
.A(n_1158),
.Y(n_1290)
);

INVx1_ASAP7_75t_L g1291 ( 
.A(n_1158),
.Y(n_1291)
);

INVx1_ASAP7_75t_L g1292 ( 
.A(n_1158),
.Y(n_1292)
);

INVx1_ASAP7_75t_L g1293 ( 
.A(n_1158),
.Y(n_1293)
);

INVx2_ASAP7_75t_L g1294 ( 
.A(n_1156),
.Y(n_1294)
);

AND2x2_ASAP7_75t_L g1295 ( 
.A(n_1204),
.B(n_1046),
.Y(n_1295)
);

INVxp67_ASAP7_75t_L g1296 ( 
.A(n_1204),
.Y(n_1296)
);

NAND2xp5_ASAP7_75t_L g1297 ( 
.A(n_1155),
.B(n_880),
.Y(n_1297)
);

INVx1_ASAP7_75t_L g1298 ( 
.A(n_1158),
.Y(n_1298)
);

NAND2xp5_ASAP7_75t_L g1299 ( 
.A(n_1155),
.B(n_890),
.Y(n_1299)
);

INVx1_ASAP7_75t_L g1300 ( 
.A(n_1158),
.Y(n_1300)
);

INVx2_ASAP7_75t_SL g1301 ( 
.A(n_1204),
.Y(n_1301)
);

BUFx3_ASAP7_75t_L g1302 ( 
.A(n_1196),
.Y(n_1302)
);

INVx2_ASAP7_75t_L g1303 ( 
.A(n_1156),
.Y(n_1303)
);

NOR2xp67_ASAP7_75t_R g1304 ( 
.A(n_1188),
.B(n_1056),
.Y(n_1304)
);

AND2x2_ASAP7_75t_L g1305 ( 
.A(n_1204),
.B(n_1060),
.Y(n_1305)
);

NAND2xp5_ASAP7_75t_L g1306 ( 
.A(n_1155),
.B(n_900),
.Y(n_1306)
);

INVx4_ASAP7_75t_L g1307 ( 
.A(n_1164),
.Y(n_1307)
);

INVx2_ASAP7_75t_SL g1308 ( 
.A(n_1204),
.Y(n_1308)
);

INVx1_ASAP7_75t_L g1309 ( 
.A(n_1158),
.Y(n_1309)
);

AND2x2_ASAP7_75t_L g1310 ( 
.A(n_1204),
.B(n_1065),
.Y(n_1310)
);

BUFx6f_ASAP7_75t_L g1311 ( 
.A(n_1162),
.Y(n_1311)
);

OAI21xp5_ASAP7_75t_L g1312 ( 
.A1(n_1155),
.A2(n_828),
.B(n_827),
.Y(n_1312)
);

AND2x2_ASAP7_75t_L g1313 ( 
.A(n_1204),
.B(n_901),
.Y(n_1313)
);

NOR2xp33_ASAP7_75t_L g1314 ( 
.A(n_1202),
.B(n_1049),
.Y(n_1314)
);

OAI21xp33_ASAP7_75t_L g1315 ( 
.A1(n_1155),
.A2(n_912),
.B(n_902),
.Y(n_1315)
);

INVx1_ASAP7_75t_L g1316 ( 
.A(n_1158),
.Y(n_1316)
);

AND2x4_ASAP7_75t_L g1317 ( 
.A(n_1196),
.B(n_859),
.Y(n_1317)
);

INVx2_ASAP7_75t_L g1318 ( 
.A(n_1208),
.Y(n_1318)
);

AND2x4_ASAP7_75t_L g1319 ( 
.A(n_1285),
.B(n_874),
.Y(n_1319)
);

NAND2xp5_ASAP7_75t_L g1320 ( 
.A(n_1239),
.B(n_914),
.Y(n_1320)
);

AND2x4_ASAP7_75t_L g1321 ( 
.A(n_1307),
.B(n_945),
.Y(n_1321)
);

OR2x2_ASAP7_75t_L g1322 ( 
.A(n_1209),
.B(n_918),
.Y(n_1322)
);

INVx2_ASAP7_75t_L g1323 ( 
.A(n_1213),
.Y(n_1323)
);

INVx1_ASAP7_75t_L g1324 ( 
.A(n_1250),
.Y(n_1324)
);

INVx2_ASAP7_75t_L g1325 ( 
.A(n_1228),
.Y(n_1325)
);

NAND2x1p5_ASAP7_75t_L g1326 ( 
.A(n_1283),
.B(n_847),
.Y(n_1326)
);

NAND2xp5_ASAP7_75t_L g1327 ( 
.A(n_1207),
.B(n_926),
.Y(n_1327)
);

NAND2xp5_ASAP7_75t_L g1328 ( 
.A(n_1240),
.B(n_935),
.Y(n_1328)
);

NAND2xp5_ASAP7_75t_L g1329 ( 
.A(n_1238),
.B(n_936),
.Y(n_1329)
);

OR2x6_ASAP7_75t_L g1330 ( 
.A(n_1227),
.B(n_1039),
.Y(n_1330)
);

INVx1_ASAP7_75t_L g1331 ( 
.A(n_1212),
.Y(n_1331)
);

NAND2x1_ASAP7_75t_SL g1332 ( 
.A(n_1261),
.B(n_836),
.Y(n_1332)
);

AND2x2_ASAP7_75t_L g1333 ( 
.A(n_1215),
.B(n_939),
.Y(n_1333)
);

INVx1_ASAP7_75t_L g1334 ( 
.A(n_1217),
.Y(n_1334)
);

BUFx6f_ASAP7_75t_L g1335 ( 
.A(n_1269),
.Y(n_1335)
);

AND2x2_ASAP7_75t_L g1336 ( 
.A(n_1313),
.B(n_943),
.Y(n_1336)
);

INVx1_ASAP7_75t_L g1337 ( 
.A(n_1218),
.Y(n_1337)
);

OR2x6_ASAP7_75t_L g1338 ( 
.A(n_1302),
.B(n_824),
.Y(n_1338)
);

AND2x4_ASAP7_75t_L g1339 ( 
.A(n_1257),
.B(n_852),
.Y(n_1339)
);

OR2x6_ASAP7_75t_L g1340 ( 
.A(n_1210),
.B(n_855),
.Y(n_1340)
);

NAND2xp5_ASAP7_75t_L g1341 ( 
.A(n_1259),
.B(n_944),
.Y(n_1341)
);

BUFx6f_ASAP7_75t_L g1342 ( 
.A(n_1210),
.Y(n_1342)
);

AND2x6_ASAP7_75t_L g1343 ( 
.A(n_1221),
.B(n_1002),
.Y(n_1343)
);

BUFx2_ASAP7_75t_L g1344 ( 
.A(n_1284),
.Y(n_1344)
);

NAND2xp5_ASAP7_75t_L g1345 ( 
.A(n_1262),
.B(n_948),
.Y(n_1345)
);

AND2x4_ASAP7_75t_L g1346 ( 
.A(n_1301),
.B(n_864),
.Y(n_1346)
);

INVx1_ASAP7_75t_L g1347 ( 
.A(n_1223),
.Y(n_1347)
);

AND2x2_ASAP7_75t_L g1348 ( 
.A(n_1264),
.B(n_953),
.Y(n_1348)
);

OR2x6_ASAP7_75t_L g1349 ( 
.A(n_1263),
.B(n_877),
.Y(n_1349)
);

INVx1_ASAP7_75t_L g1350 ( 
.A(n_1226),
.Y(n_1350)
);

AND2x4_ASAP7_75t_L g1351 ( 
.A(n_1308),
.B(n_881),
.Y(n_1351)
);

AND2x2_ASAP7_75t_L g1352 ( 
.A(n_1271),
.B(n_955),
.Y(n_1352)
);

INVx1_ASAP7_75t_L g1353 ( 
.A(n_1265),
.Y(n_1353)
);

NAND2x1p5_ASAP7_75t_L g1354 ( 
.A(n_1263),
.B(n_1089),
.Y(n_1354)
);

NAND2x1p5_ASAP7_75t_L g1355 ( 
.A(n_1272),
.B(n_1091),
.Y(n_1355)
);

BUFx2_ASAP7_75t_L g1356 ( 
.A(n_1317),
.Y(n_1356)
);

NAND2xp5_ASAP7_75t_L g1357 ( 
.A(n_1286),
.B(n_970),
.Y(n_1357)
);

INVx1_ASAP7_75t_L g1358 ( 
.A(n_1266),
.Y(n_1358)
);

INVx1_ASAP7_75t_L g1359 ( 
.A(n_1267),
.Y(n_1359)
);

INVx2_ASAP7_75t_L g1360 ( 
.A(n_1260),
.Y(n_1360)
);

NAND2xp5_ASAP7_75t_L g1361 ( 
.A(n_1297),
.B(n_973),
.Y(n_1361)
);

AND2x2_ASAP7_75t_L g1362 ( 
.A(n_1277),
.B(n_978),
.Y(n_1362)
);

NAND2xp5_ASAP7_75t_SL g1363 ( 
.A(n_1220),
.B(n_980),
.Y(n_1363)
);

BUFx6f_ASAP7_75t_L g1364 ( 
.A(n_1272),
.Y(n_1364)
);

NAND2xp5_ASAP7_75t_L g1365 ( 
.A(n_1299),
.B(n_1306),
.Y(n_1365)
);

AND2x2_ASAP7_75t_L g1366 ( 
.A(n_1278),
.B(n_983),
.Y(n_1366)
);

OR2x6_ASAP7_75t_L g1367 ( 
.A(n_1275),
.B(n_892),
.Y(n_1367)
);

CKINVDCx8_ASAP7_75t_R g1368 ( 
.A(n_1276),
.Y(n_1368)
);

NOR2xp33_ASAP7_75t_L g1369 ( 
.A(n_1216),
.B(n_984),
.Y(n_1369)
);

INVx6_ASAP7_75t_L g1370 ( 
.A(n_1211),
.Y(n_1370)
);

NAND2xp5_ASAP7_75t_L g1371 ( 
.A(n_1312),
.B(n_985),
.Y(n_1371)
);

INVx2_ASAP7_75t_SL g1372 ( 
.A(n_1219),
.Y(n_1372)
);

AND2x2_ASAP7_75t_L g1373 ( 
.A(n_1279),
.B(n_996),
.Y(n_1373)
);

NAND2xp5_ASAP7_75t_L g1374 ( 
.A(n_1233),
.B(n_999),
.Y(n_1374)
);

INVx1_ASAP7_75t_L g1375 ( 
.A(n_1268),
.Y(n_1375)
);

INVx5_ASAP7_75t_L g1376 ( 
.A(n_1275),
.Y(n_1376)
);

BUFx2_ASAP7_75t_L g1377 ( 
.A(n_1288),
.Y(n_1377)
);

INVxp67_ASAP7_75t_SL g1378 ( 
.A(n_1296),
.Y(n_1378)
);

INVx2_ASAP7_75t_L g1379 ( 
.A(n_1270),
.Y(n_1379)
);

NAND2xp5_ASAP7_75t_L g1380 ( 
.A(n_1281),
.B(n_1004),
.Y(n_1380)
);

OR2x2_ASAP7_75t_L g1381 ( 
.A(n_1241),
.B(n_1014),
.Y(n_1381)
);

OR2x2_ASAP7_75t_L g1382 ( 
.A(n_1214),
.B(n_1017),
.Y(n_1382)
);

AND2x4_ASAP7_75t_L g1383 ( 
.A(n_1254),
.B(n_894),
.Y(n_1383)
);

OR2x2_ASAP7_75t_L g1384 ( 
.A(n_1256),
.B(n_1025),
.Y(n_1384)
);

NAND2x1_ASAP7_75t_L g1385 ( 
.A(n_1234),
.B(n_858),
.Y(n_1385)
);

OR2x2_ASAP7_75t_L g1386 ( 
.A(n_1289),
.B(n_1026),
.Y(n_1386)
);

INVx4_ASAP7_75t_L g1387 ( 
.A(n_1287),
.Y(n_1387)
);

INVx2_ASAP7_75t_L g1388 ( 
.A(n_1274),
.Y(n_1388)
);

OR2x2_ASAP7_75t_L g1389 ( 
.A(n_1295),
.B(n_1028),
.Y(n_1389)
);

INVx1_ASAP7_75t_L g1390 ( 
.A(n_1273),
.Y(n_1390)
);

BUFx2_ASAP7_75t_L g1391 ( 
.A(n_1276),
.Y(n_1391)
);

INVx5_ASAP7_75t_L g1392 ( 
.A(n_1287),
.Y(n_1392)
);

NOR2xp33_ASAP7_75t_L g1393 ( 
.A(n_1245),
.B(n_1030),
.Y(n_1393)
);

INVx2_ASAP7_75t_L g1394 ( 
.A(n_1282),
.Y(n_1394)
);

INVx2_ASAP7_75t_L g1395 ( 
.A(n_1294),
.Y(n_1395)
);

NAND2xp5_ASAP7_75t_L g1396 ( 
.A(n_1305),
.B(n_1035),
.Y(n_1396)
);

NAND2xp5_ASAP7_75t_L g1397 ( 
.A(n_1310),
.B(n_1036),
.Y(n_1397)
);

AND2x2_ASAP7_75t_L g1398 ( 
.A(n_1230),
.B(n_1047),
.Y(n_1398)
);

BUFx6f_ASAP7_75t_L g1399 ( 
.A(n_1311),
.Y(n_1399)
);

NOR2xp33_ASAP7_75t_SL g1400 ( 
.A(n_1258),
.B(n_1048),
.Y(n_1400)
);

NAND2xp5_ASAP7_75t_L g1401 ( 
.A(n_1280),
.B(n_1054),
.Y(n_1401)
);

INVx1_ASAP7_75t_SL g1402 ( 
.A(n_1222),
.Y(n_1402)
);

AND2x4_ASAP7_75t_L g1403 ( 
.A(n_1311),
.B(n_1237),
.Y(n_1403)
);

OR2x2_ASAP7_75t_L g1404 ( 
.A(n_1229),
.B(n_9),
.Y(n_1404)
);

INVx1_ASAP7_75t_L g1405 ( 
.A(n_1290),
.Y(n_1405)
);

AND2x4_ASAP7_75t_L g1406 ( 
.A(n_1246),
.B(n_895),
.Y(n_1406)
);

NAND2xp5_ASAP7_75t_L g1407 ( 
.A(n_1291),
.B(n_897),
.Y(n_1407)
);

INVx2_ASAP7_75t_L g1408 ( 
.A(n_1303),
.Y(n_1408)
);

INVx3_ASAP7_75t_L g1409 ( 
.A(n_1235),
.Y(n_1409)
);

NOR2xp33_ASAP7_75t_L g1410 ( 
.A(n_1249),
.B(n_899),
.Y(n_1410)
);

INVx2_ASAP7_75t_L g1411 ( 
.A(n_1242),
.Y(n_1411)
);

AND2x4_ASAP7_75t_L g1412 ( 
.A(n_1247),
.B(n_927),
.Y(n_1412)
);

BUFx6f_ASAP7_75t_L g1413 ( 
.A(n_1252),
.Y(n_1413)
);

OR2x6_ASAP7_75t_L g1414 ( 
.A(n_1253),
.B(n_932),
.Y(n_1414)
);

BUFx8_ASAP7_75t_SL g1415 ( 
.A(n_1232),
.Y(n_1415)
);

AND2x4_ASAP7_75t_L g1416 ( 
.A(n_1225),
.B(n_938),
.Y(n_1416)
);

BUFx3_ASAP7_75t_L g1417 ( 
.A(n_1243),
.Y(n_1417)
);

INVx1_ASAP7_75t_L g1418 ( 
.A(n_1292),
.Y(n_1418)
);

INVx1_ASAP7_75t_SL g1419 ( 
.A(n_1276),
.Y(n_1419)
);

INVx1_ASAP7_75t_L g1420 ( 
.A(n_1293),
.Y(n_1420)
);

NAND2x1p5_ASAP7_75t_L g1421 ( 
.A(n_1298),
.B(n_1091),
.Y(n_1421)
);

INVx4_ASAP7_75t_L g1422 ( 
.A(n_1225),
.Y(n_1422)
);

NOR2xp33_ASAP7_75t_L g1423 ( 
.A(n_1315),
.B(n_913),
.Y(n_1423)
);

BUFx6f_ASAP7_75t_L g1424 ( 
.A(n_1231),
.Y(n_1424)
);

AND2x4_ASAP7_75t_L g1425 ( 
.A(n_1225),
.B(n_950),
.Y(n_1425)
);

NOR2xp33_ASAP7_75t_L g1426 ( 
.A(n_1314),
.B(n_952),
.Y(n_1426)
);

INVx1_ASAP7_75t_L g1427 ( 
.A(n_1300),
.Y(n_1427)
);

NAND2xp5_ASAP7_75t_L g1428 ( 
.A(n_1309),
.B(n_1037),
.Y(n_1428)
);

INVx2_ASAP7_75t_L g1429 ( 
.A(n_1248),
.Y(n_1429)
);

INVx1_ASAP7_75t_L g1430 ( 
.A(n_1316),
.Y(n_1430)
);

INVx2_ASAP7_75t_L g1431 ( 
.A(n_1236),
.Y(n_1431)
);

AND2x4_ASAP7_75t_L g1432 ( 
.A(n_1251),
.B(n_956),
.Y(n_1432)
);

NOR2xp33_ASAP7_75t_L g1433 ( 
.A(n_1244),
.B(n_954),
.Y(n_1433)
);

NAND2xp5_ASAP7_75t_L g1434 ( 
.A(n_1224),
.B(n_1042),
.Y(n_1434)
);

NOR2xp33_ASAP7_75t_L g1435 ( 
.A(n_1255),
.B(n_957),
.Y(n_1435)
);

AND2x2_ASAP7_75t_L g1436 ( 
.A(n_1304),
.B(n_1094),
.Y(n_1436)
);

NAND2xp5_ASAP7_75t_SL g1437 ( 
.A(n_1301),
.B(n_755),
.Y(n_1437)
);

NOR2xp33_ASAP7_75t_L g1438 ( 
.A(n_1239),
.B(n_958),
.Y(n_1438)
);

AND2x4_ASAP7_75t_L g1439 ( 
.A(n_1285),
.B(n_967),
.Y(n_1439)
);

BUFx8_ASAP7_75t_L g1440 ( 
.A(n_1269),
.Y(n_1440)
);

AND2x2_ASAP7_75t_L g1441 ( 
.A(n_1215),
.B(n_1094),
.Y(n_1441)
);

OR2x2_ASAP7_75t_L g1442 ( 
.A(n_1209),
.B(n_10),
.Y(n_1442)
);

BUFx6f_ASAP7_75t_L g1443 ( 
.A(n_1261),
.Y(n_1443)
);

NAND2xp5_ASAP7_75t_L g1444 ( 
.A(n_1239),
.B(n_963),
.Y(n_1444)
);

INVxp67_ASAP7_75t_L g1445 ( 
.A(n_1214),
.Y(n_1445)
);

BUFx6f_ASAP7_75t_L g1446 ( 
.A(n_1261),
.Y(n_1446)
);

AND2x2_ASAP7_75t_L g1447 ( 
.A(n_1215),
.B(n_1098),
.Y(n_1447)
);

INVx2_ASAP7_75t_L g1448 ( 
.A(n_1208),
.Y(n_1448)
);

INVx2_ASAP7_75t_L g1449 ( 
.A(n_1208),
.Y(n_1449)
);

BUFx3_ASAP7_75t_L g1450 ( 
.A(n_1269),
.Y(n_1450)
);

AND2x4_ASAP7_75t_L g1451 ( 
.A(n_1285),
.B(n_969),
.Y(n_1451)
);

BUFx3_ASAP7_75t_L g1452 ( 
.A(n_1269),
.Y(n_1452)
);

INVx6_ASAP7_75t_L g1453 ( 
.A(n_1285),
.Y(n_1453)
);

INVx1_ASAP7_75t_SL g1454 ( 
.A(n_1261),
.Y(n_1454)
);

INVx4_ASAP7_75t_L g1455 ( 
.A(n_1285),
.Y(n_1455)
);

AND2x6_ASAP7_75t_L g1456 ( 
.A(n_1221),
.B(n_971),
.Y(n_1456)
);

INVx2_ASAP7_75t_L g1457 ( 
.A(n_1208),
.Y(n_1457)
);

INVx5_ASAP7_75t_L g1458 ( 
.A(n_1285),
.Y(n_1458)
);

INVx1_ASAP7_75t_L g1459 ( 
.A(n_1250),
.Y(n_1459)
);

BUFx8_ASAP7_75t_SL g1460 ( 
.A(n_1269),
.Y(n_1460)
);

INVx2_ASAP7_75t_L g1461 ( 
.A(n_1208),
.Y(n_1461)
);

INVx1_ASAP7_75t_L g1462 ( 
.A(n_1250),
.Y(n_1462)
);

NOR2x1_ASAP7_75t_R g1463 ( 
.A(n_1269),
.B(n_758),
.Y(n_1463)
);

INVx1_ASAP7_75t_L g1464 ( 
.A(n_1250),
.Y(n_1464)
);

AND2x4_ASAP7_75t_L g1465 ( 
.A(n_1285),
.B(n_975),
.Y(n_1465)
);

NAND2xp5_ASAP7_75t_L g1466 ( 
.A(n_1239),
.B(n_981),
.Y(n_1466)
);

BUFx6f_ASAP7_75t_L g1467 ( 
.A(n_1269),
.Y(n_1467)
);

OR2x2_ASAP7_75t_L g1468 ( 
.A(n_1209),
.B(n_11),
.Y(n_1468)
);

NAND2xp5_ASAP7_75t_L g1469 ( 
.A(n_1239),
.B(n_1032),
.Y(n_1469)
);

AND2x4_ASAP7_75t_L g1470 ( 
.A(n_1285),
.B(n_982),
.Y(n_1470)
);

INVx2_ASAP7_75t_L g1471 ( 
.A(n_1208),
.Y(n_1471)
);

HB1xp67_ASAP7_75t_L g1472 ( 
.A(n_1209),
.Y(n_1472)
);

INVx3_ASAP7_75t_L g1473 ( 
.A(n_1285),
.Y(n_1473)
);

NAND2xp5_ASAP7_75t_L g1474 ( 
.A(n_1239),
.B(n_1057),
.Y(n_1474)
);

INVx6_ASAP7_75t_L g1475 ( 
.A(n_1285),
.Y(n_1475)
);

INVx1_ASAP7_75t_L g1476 ( 
.A(n_1331),
.Y(n_1476)
);

INVx4_ASAP7_75t_L g1477 ( 
.A(n_1458),
.Y(n_1477)
);

BUFx12f_ASAP7_75t_L g1478 ( 
.A(n_1440),
.Y(n_1478)
);

INVx8_ASAP7_75t_L g1479 ( 
.A(n_1460),
.Y(n_1479)
);

AOI22xp33_ASAP7_75t_L g1480 ( 
.A1(n_1433),
.A2(n_1456),
.B1(n_1426),
.B2(n_1398),
.Y(n_1480)
);

BUFx6f_ASAP7_75t_L g1481 ( 
.A(n_1467),
.Y(n_1481)
);

INVx2_ASAP7_75t_SL g1482 ( 
.A(n_1453),
.Y(n_1482)
);

OR2x6_ASAP7_75t_L g1483 ( 
.A(n_1475),
.B(n_988),
.Y(n_1483)
);

BUFx3_ASAP7_75t_L g1484 ( 
.A(n_1450),
.Y(n_1484)
);

AND2x2_ASAP7_75t_L g1485 ( 
.A(n_1348),
.B(n_12),
.Y(n_1485)
);

AND2x2_ASAP7_75t_L g1486 ( 
.A(n_1352),
.B(n_12),
.Y(n_1486)
);

BUFx6f_ASAP7_75t_L g1487 ( 
.A(n_1467),
.Y(n_1487)
);

INVx2_ASAP7_75t_SL g1488 ( 
.A(n_1376),
.Y(n_1488)
);

INVx5_ASAP7_75t_L g1489 ( 
.A(n_1443),
.Y(n_1489)
);

BUFx12f_ASAP7_75t_L g1490 ( 
.A(n_1446),
.Y(n_1490)
);

BUFx6f_ASAP7_75t_L g1491 ( 
.A(n_1335),
.Y(n_1491)
);

CKINVDCx16_ASAP7_75t_R g1492 ( 
.A(n_1452),
.Y(n_1492)
);

INVx1_ASAP7_75t_L g1493 ( 
.A(n_1334),
.Y(n_1493)
);

INVx4_ASAP7_75t_L g1494 ( 
.A(n_1458),
.Y(n_1494)
);

OR2x6_ASAP7_75t_L g1495 ( 
.A(n_1370),
.B(n_989),
.Y(n_1495)
);

BUFx2_ASAP7_75t_L g1496 ( 
.A(n_1344),
.Y(n_1496)
);

OR2x2_ASAP7_75t_L g1497 ( 
.A(n_1472),
.B(n_1098),
.Y(n_1497)
);

INVx1_ASAP7_75t_L g1498 ( 
.A(n_1337),
.Y(n_1498)
);

NAND2xp5_ASAP7_75t_L g1499 ( 
.A(n_1431),
.B(n_13),
.Y(n_1499)
);

BUFx3_ASAP7_75t_L g1500 ( 
.A(n_1376),
.Y(n_1500)
);

CKINVDCx20_ASAP7_75t_R g1501 ( 
.A(n_1415),
.Y(n_1501)
);

INVx3_ASAP7_75t_L g1502 ( 
.A(n_1455),
.Y(n_1502)
);

BUFx2_ASAP7_75t_SL g1503 ( 
.A(n_1392),
.Y(n_1503)
);

INVx3_ASAP7_75t_L g1504 ( 
.A(n_1392),
.Y(n_1504)
);

INVx5_ASAP7_75t_L g1505 ( 
.A(n_1349),
.Y(n_1505)
);

INVx1_ASAP7_75t_L g1506 ( 
.A(n_1347),
.Y(n_1506)
);

BUFx6f_ASAP7_75t_L g1507 ( 
.A(n_1342),
.Y(n_1507)
);

BUFx3_ASAP7_75t_L g1508 ( 
.A(n_1364),
.Y(n_1508)
);

BUFx6f_ASAP7_75t_L g1509 ( 
.A(n_1399),
.Y(n_1509)
);

AO21x2_ASAP7_75t_L g1510 ( 
.A1(n_1365),
.A2(n_1007),
.B(n_1003),
.Y(n_1510)
);

BUFx4_ASAP7_75t_R g1511 ( 
.A(n_1417),
.Y(n_1511)
);

INVx1_ASAP7_75t_SL g1512 ( 
.A(n_1377),
.Y(n_1512)
);

CKINVDCx5p33_ASAP7_75t_R g1513 ( 
.A(n_1454),
.Y(n_1513)
);

CKINVDCx5p33_ASAP7_75t_R g1514 ( 
.A(n_1424),
.Y(n_1514)
);

BUFx2_ASAP7_75t_L g1515 ( 
.A(n_1356),
.Y(n_1515)
);

BUFx3_ASAP7_75t_L g1516 ( 
.A(n_1403),
.Y(n_1516)
);

BUFx3_ASAP7_75t_L g1517 ( 
.A(n_1473),
.Y(n_1517)
);

INVx3_ASAP7_75t_L g1518 ( 
.A(n_1387),
.Y(n_1518)
);

BUFx12f_ASAP7_75t_L g1519 ( 
.A(n_1372),
.Y(n_1519)
);

BUFx4_ASAP7_75t_SL g1520 ( 
.A(n_1338),
.Y(n_1520)
);

INVx3_ASAP7_75t_L g1521 ( 
.A(n_1368),
.Y(n_1521)
);

INVx1_ASAP7_75t_L g1522 ( 
.A(n_1350),
.Y(n_1522)
);

INVx6_ASAP7_75t_L g1523 ( 
.A(n_1319),
.Y(n_1523)
);

INVx8_ASAP7_75t_L g1524 ( 
.A(n_1367),
.Y(n_1524)
);

INVx4_ASAP7_75t_L g1525 ( 
.A(n_1409),
.Y(n_1525)
);

INVx3_ASAP7_75t_L g1526 ( 
.A(n_1413),
.Y(n_1526)
);

INVx1_ASAP7_75t_L g1527 ( 
.A(n_1353),
.Y(n_1527)
);

INVx1_ASAP7_75t_SL g1528 ( 
.A(n_1402),
.Y(n_1528)
);

BUFx2_ASAP7_75t_L g1529 ( 
.A(n_1445),
.Y(n_1529)
);

INVx1_ASAP7_75t_SL g1530 ( 
.A(n_1441),
.Y(n_1530)
);

INVx1_ASAP7_75t_L g1531 ( 
.A(n_1358),
.Y(n_1531)
);

BUFx4_ASAP7_75t_SL g1532 ( 
.A(n_1330),
.Y(n_1532)
);

NAND2xp5_ASAP7_75t_L g1533 ( 
.A(n_1438),
.B(n_1456),
.Y(n_1533)
);

CKINVDCx16_ASAP7_75t_R g1534 ( 
.A(n_1400),
.Y(n_1534)
);

BUFx12f_ASAP7_75t_L g1535 ( 
.A(n_1340),
.Y(n_1535)
);

INVx2_ASAP7_75t_L g1536 ( 
.A(n_1429),
.Y(n_1536)
);

NAND2xp5_ASAP7_75t_L g1537 ( 
.A(n_1362),
.B(n_13),
.Y(n_1537)
);

INVx8_ASAP7_75t_L g1538 ( 
.A(n_1343),
.Y(n_1538)
);

BUFx6f_ASAP7_75t_L g1539 ( 
.A(n_1354),
.Y(n_1539)
);

AND2x4_ASAP7_75t_L g1540 ( 
.A(n_1422),
.B(n_1022),
.Y(n_1540)
);

BUFx3_ASAP7_75t_L g1541 ( 
.A(n_1355),
.Y(n_1541)
);

INVx2_ASAP7_75t_L g1542 ( 
.A(n_1411),
.Y(n_1542)
);

INVx5_ASAP7_75t_L g1543 ( 
.A(n_1343),
.Y(n_1543)
);

BUFx3_ASAP7_75t_L g1544 ( 
.A(n_1321),
.Y(n_1544)
);

INVx4_ASAP7_75t_L g1545 ( 
.A(n_1326),
.Y(n_1545)
);

AND2x2_ASAP7_75t_L g1546 ( 
.A(n_1366),
.B(n_14),
.Y(n_1546)
);

INVx5_ASAP7_75t_L g1547 ( 
.A(n_1414),
.Y(n_1547)
);

INVx2_ASAP7_75t_L g1548 ( 
.A(n_1318),
.Y(n_1548)
);

INVx3_ASAP7_75t_L g1549 ( 
.A(n_1439),
.Y(n_1549)
);

BUFx3_ASAP7_75t_L g1550 ( 
.A(n_1451),
.Y(n_1550)
);

NAND2x1p5_ASAP7_75t_L g1551 ( 
.A(n_1391),
.B(n_1104),
.Y(n_1551)
);

NAND2x1p5_ASAP7_75t_L g1552 ( 
.A(n_1419),
.B(n_1104),
.Y(n_1552)
);

BUFx8_ASAP7_75t_L g1553 ( 
.A(n_1465),
.Y(n_1553)
);

INVx1_ASAP7_75t_L g1554 ( 
.A(n_1359),
.Y(n_1554)
);

INVx2_ASAP7_75t_SL g1555 ( 
.A(n_1447),
.Y(n_1555)
);

NOR2xp33_ASAP7_75t_L g1556 ( 
.A(n_1378),
.B(n_761),
.Y(n_1556)
);

NAND2xp5_ASAP7_75t_L g1557 ( 
.A(n_1373),
.B(n_14),
.Y(n_1557)
);

BUFx5_ASAP7_75t_L g1558 ( 
.A(n_1324),
.Y(n_1558)
);

CKINVDCx5p33_ASAP7_75t_R g1559 ( 
.A(n_1369),
.Y(n_1559)
);

INVx2_ASAP7_75t_SL g1560 ( 
.A(n_1470),
.Y(n_1560)
);

INVx5_ASAP7_75t_L g1561 ( 
.A(n_1416),
.Y(n_1561)
);

INVx1_ASAP7_75t_SL g1562 ( 
.A(n_1442),
.Y(n_1562)
);

INVx6_ASAP7_75t_L g1563 ( 
.A(n_1339),
.Y(n_1563)
);

CKINVDCx16_ASAP7_75t_R g1564 ( 
.A(n_1336),
.Y(n_1564)
);

INVx1_ASAP7_75t_SL g1565 ( 
.A(n_1468),
.Y(n_1565)
);

BUFx3_ASAP7_75t_L g1566 ( 
.A(n_1406),
.Y(n_1566)
);

BUFx5_ASAP7_75t_L g1567 ( 
.A(n_1459),
.Y(n_1567)
);

INVx2_ASAP7_75t_L g1568 ( 
.A(n_1323),
.Y(n_1568)
);

INVx6_ASAP7_75t_L g1569 ( 
.A(n_1383),
.Y(n_1569)
);

AOI22xp5_ASAP7_75t_L g1570 ( 
.A1(n_1423),
.A2(n_1023),
.B1(n_765),
.B2(n_768),
.Y(n_1570)
);

BUFx12f_ASAP7_75t_L g1571 ( 
.A(n_1346),
.Y(n_1571)
);

INVx1_ASAP7_75t_L g1572 ( 
.A(n_1375),
.Y(n_1572)
);

BUFx12f_ASAP7_75t_L g1573 ( 
.A(n_1351),
.Y(n_1573)
);

NAND2xp5_ASAP7_75t_L g1574 ( 
.A(n_1462),
.B(n_15),
.Y(n_1574)
);

INVx1_ASAP7_75t_SL g1575 ( 
.A(n_1333),
.Y(n_1575)
);

INVxp33_ASAP7_75t_L g1576 ( 
.A(n_1463),
.Y(n_1576)
);

INVx4_ASAP7_75t_L g1577 ( 
.A(n_1425),
.Y(n_1577)
);

INVx4_ASAP7_75t_L g1578 ( 
.A(n_1436),
.Y(n_1578)
);

BUFx6f_ASAP7_75t_L g1579 ( 
.A(n_1412),
.Y(n_1579)
);

INVx2_ASAP7_75t_L g1580 ( 
.A(n_1325),
.Y(n_1580)
);

BUFx4_ASAP7_75t_SL g1581 ( 
.A(n_1404),
.Y(n_1581)
);

INVx1_ASAP7_75t_SL g1582 ( 
.A(n_1322),
.Y(n_1582)
);

INVx1_ASAP7_75t_SL g1583 ( 
.A(n_1384),
.Y(n_1583)
);

INVx2_ASAP7_75t_L g1584 ( 
.A(n_1360),
.Y(n_1584)
);

BUFx2_ASAP7_75t_SL g1585 ( 
.A(n_1464),
.Y(n_1585)
);

AOI22xp33_ASAP7_75t_SL g1586 ( 
.A1(n_1371),
.A2(n_784),
.B1(n_785),
.B2(n_762),
.Y(n_1586)
);

INVx3_ASAP7_75t_L g1587 ( 
.A(n_1421),
.Y(n_1587)
);

BUFx2_ASAP7_75t_L g1588 ( 
.A(n_1432),
.Y(n_1588)
);

BUFx12f_ASAP7_75t_L g1589 ( 
.A(n_1382),
.Y(n_1589)
);

NAND2x1p5_ASAP7_75t_L g1590 ( 
.A(n_1390),
.B(n_1405),
.Y(n_1590)
);

BUFx12f_ASAP7_75t_L g1591 ( 
.A(n_1386),
.Y(n_1591)
);

INVx8_ASAP7_75t_L g1592 ( 
.A(n_1332),
.Y(n_1592)
);

CKINVDCx6p67_ASAP7_75t_R g1593 ( 
.A(n_1478),
.Y(n_1593)
);

AOI22xp33_ASAP7_75t_SL g1594 ( 
.A1(n_1534),
.A2(n_1410),
.B1(n_1393),
.B2(n_1435),
.Y(n_1594)
);

INVx6_ASAP7_75t_L g1595 ( 
.A(n_1489),
.Y(n_1595)
);

BUFx6f_ASAP7_75t_L g1596 ( 
.A(n_1484),
.Y(n_1596)
);

INVx2_ASAP7_75t_L g1597 ( 
.A(n_1536),
.Y(n_1597)
);

AOI22xp33_ASAP7_75t_L g1598 ( 
.A1(n_1480),
.A2(n_1381),
.B1(n_1388),
.B2(n_1379),
.Y(n_1598)
);

AOI22xp33_ASAP7_75t_L g1599 ( 
.A1(n_1571),
.A2(n_1395),
.B1(n_1408),
.B2(n_1394),
.Y(n_1599)
);

NAND2xp5_ASAP7_75t_L g1600 ( 
.A(n_1575),
.B(n_1389),
.Y(n_1600)
);

INVx6_ASAP7_75t_L g1601 ( 
.A(n_1489),
.Y(n_1601)
);

INVx2_ASAP7_75t_L g1602 ( 
.A(n_1542),
.Y(n_1602)
);

AOI22xp33_ASAP7_75t_SL g1603 ( 
.A1(n_1533),
.A2(n_1434),
.B1(n_1329),
.B2(n_1444),
.Y(n_1603)
);

BUFx8_ASAP7_75t_L g1604 ( 
.A(n_1490),
.Y(n_1604)
);

INVx1_ASAP7_75t_L g1605 ( 
.A(n_1476),
.Y(n_1605)
);

BUFx2_ASAP7_75t_R g1606 ( 
.A(n_1503),
.Y(n_1606)
);

INVx1_ASAP7_75t_L g1607 ( 
.A(n_1493),
.Y(n_1607)
);

AOI22xp33_ASAP7_75t_SL g1608 ( 
.A1(n_1505),
.A2(n_1469),
.B1(n_1474),
.B2(n_1466),
.Y(n_1608)
);

AOI22xp5_ASAP7_75t_L g1609 ( 
.A1(n_1559),
.A2(n_1320),
.B1(n_1396),
.B2(n_1380),
.Y(n_1609)
);

INVxp67_ASAP7_75t_SL g1610 ( 
.A(n_1496),
.Y(n_1610)
);

OAI22xp33_ASAP7_75t_L g1611 ( 
.A1(n_1564),
.A2(n_1327),
.B1(n_1345),
.B2(n_1341),
.Y(n_1611)
);

INVx6_ASAP7_75t_L g1612 ( 
.A(n_1492),
.Y(n_1612)
);

NAND2xp5_ASAP7_75t_L g1613 ( 
.A(n_1583),
.B(n_1418),
.Y(n_1613)
);

CKINVDCx20_ASAP7_75t_R g1614 ( 
.A(n_1501),
.Y(n_1614)
);

INVx1_ASAP7_75t_L g1615 ( 
.A(n_1498),
.Y(n_1615)
);

AOI22xp33_ASAP7_75t_L g1616 ( 
.A1(n_1573),
.A2(n_1449),
.B1(n_1457),
.B2(n_1448),
.Y(n_1616)
);

BUFx2_ASAP7_75t_L g1617 ( 
.A(n_1589),
.Y(n_1617)
);

CKINVDCx11_ASAP7_75t_R g1618 ( 
.A(n_1479),
.Y(n_1618)
);

BUFx6f_ASAP7_75t_L g1619 ( 
.A(n_1500),
.Y(n_1619)
);

INVx1_ASAP7_75t_L g1620 ( 
.A(n_1506),
.Y(n_1620)
);

INVx1_ASAP7_75t_SL g1621 ( 
.A(n_1511),
.Y(n_1621)
);

CKINVDCx5p33_ASAP7_75t_R g1622 ( 
.A(n_1520),
.Y(n_1622)
);

AOI22xp33_ASAP7_75t_SL g1623 ( 
.A1(n_1505),
.A2(n_1397),
.B1(n_1357),
.B2(n_1361),
.Y(n_1623)
);

INVx2_ASAP7_75t_L g1624 ( 
.A(n_1548),
.Y(n_1624)
);

INVx1_ASAP7_75t_L g1625 ( 
.A(n_1522),
.Y(n_1625)
);

AOI22xp33_ASAP7_75t_SL g1626 ( 
.A1(n_1485),
.A2(n_1374),
.B1(n_1428),
.B2(n_1407),
.Y(n_1626)
);

OAI22xp5_ASAP7_75t_L g1627 ( 
.A1(n_1570),
.A2(n_1328),
.B1(n_1427),
.B2(n_1420),
.Y(n_1627)
);

NAND2xp5_ASAP7_75t_L g1628 ( 
.A(n_1582),
.B(n_1430),
.Y(n_1628)
);

INVx2_ASAP7_75t_L g1629 ( 
.A(n_1568),
.Y(n_1629)
);

INVx4_ASAP7_75t_SL g1630 ( 
.A(n_1563),
.Y(n_1630)
);

CKINVDCx5p33_ASAP7_75t_R g1631 ( 
.A(n_1513),
.Y(n_1631)
);

INVx1_ASAP7_75t_L g1632 ( 
.A(n_1527),
.Y(n_1632)
);

AOI22xp33_ASAP7_75t_L g1633 ( 
.A1(n_1569),
.A2(n_1471),
.B1(n_1461),
.B2(n_1437),
.Y(n_1633)
);

AOI22xp33_ASAP7_75t_L g1634 ( 
.A1(n_1591),
.A2(n_1363),
.B1(n_1401),
.B2(n_1385),
.Y(n_1634)
);

OAI22xp5_ASAP7_75t_L g1635 ( 
.A1(n_1529),
.A2(n_885),
.B1(n_909),
.B2(n_789),
.Y(n_1635)
);

BUFx3_ASAP7_75t_L g1636 ( 
.A(n_1481),
.Y(n_1636)
);

OAI21xp5_ASAP7_75t_SL g1637 ( 
.A1(n_1486),
.A2(n_1010),
.B(n_910),
.Y(n_1637)
);

BUFx2_ASAP7_75t_L g1638 ( 
.A(n_1516),
.Y(n_1638)
);

OAI21xp5_ASAP7_75t_SL g1639 ( 
.A1(n_1546),
.A2(n_1012),
.B(n_966),
.Y(n_1639)
);

INVx1_ASAP7_75t_L g1640 ( 
.A(n_1531),
.Y(n_1640)
);

NAND2xp5_ASAP7_75t_L g1641 ( 
.A(n_1530),
.B(n_15),
.Y(n_1641)
);

BUFx2_ASAP7_75t_L g1642 ( 
.A(n_1550),
.Y(n_1642)
);

NAND2xp5_ASAP7_75t_L g1643 ( 
.A(n_1528),
.B(n_16),
.Y(n_1643)
);

AOI22xp33_ASAP7_75t_SL g1644 ( 
.A1(n_1524),
.A2(n_1547),
.B1(n_1588),
.B2(n_1561),
.Y(n_1644)
);

OAI22xp33_ASAP7_75t_L g1645 ( 
.A1(n_1562),
.A2(n_769),
.B1(n_770),
.B2(n_766),
.Y(n_1645)
);

INVx1_ASAP7_75t_L g1646 ( 
.A(n_1554),
.Y(n_1646)
);

INVx1_ASAP7_75t_L g1647 ( 
.A(n_1572),
.Y(n_1647)
);

AOI22xp33_ASAP7_75t_SL g1648 ( 
.A1(n_1547),
.A2(n_934),
.B1(n_1015),
.B2(n_966),
.Y(n_1648)
);

NAND2x1p5_ASAP7_75t_L g1649 ( 
.A(n_1482),
.B(n_1543),
.Y(n_1649)
);

BUFx2_ASAP7_75t_L g1650 ( 
.A(n_1579),
.Y(n_1650)
);

BUFx12f_ASAP7_75t_L g1651 ( 
.A(n_1553),
.Y(n_1651)
);

AOI22xp33_ASAP7_75t_L g1652 ( 
.A1(n_1566),
.A2(n_966),
.B1(n_1015),
.B2(n_876),
.Y(n_1652)
);

CKINVDCx20_ASAP7_75t_R g1653 ( 
.A(n_1514),
.Y(n_1653)
);

BUFx3_ASAP7_75t_L g1654 ( 
.A(n_1487),
.Y(n_1654)
);

CKINVDCx5p33_ASAP7_75t_R g1655 ( 
.A(n_1532),
.Y(n_1655)
);

AOI22xp33_ASAP7_75t_L g1656 ( 
.A1(n_1560),
.A2(n_1015),
.B1(n_876),
.B2(n_774),
.Y(n_1656)
);

OAI22xp5_ASAP7_75t_L g1657 ( 
.A1(n_1537),
.A2(n_1557),
.B1(n_1590),
.B2(n_1556),
.Y(n_1657)
);

AOI22xp33_ASAP7_75t_L g1658 ( 
.A1(n_1549),
.A2(n_876),
.B1(n_775),
.B2(n_778),
.Y(n_1658)
);

INVx1_ASAP7_75t_SL g1659 ( 
.A(n_1512),
.Y(n_1659)
);

AOI22xp33_ASAP7_75t_SL g1660 ( 
.A1(n_1561),
.A2(n_876),
.B1(n_831),
.B2(n_857),
.Y(n_1660)
);

INVx1_ASAP7_75t_L g1661 ( 
.A(n_1580),
.Y(n_1661)
);

OAI22xp33_ASAP7_75t_L g1662 ( 
.A1(n_1565),
.A2(n_780),
.B1(n_782),
.B2(n_773),
.Y(n_1662)
);

AOI22xp33_ASAP7_75t_SL g1663 ( 
.A1(n_1543),
.A2(n_876),
.B1(n_849),
.B2(n_817),
.Y(n_1663)
);

CKINVDCx20_ASAP7_75t_R g1664 ( 
.A(n_1538),
.Y(n_1664)
);

AOI22xp33_ASAP7_75t_L g1665 ( 
.A1(n_1495),
.A2(n_795),
.B1(n_796),
.B2(n_793),
.Y(n_1665)
);

INVx1_ASAP7_75t_L g1666 ( 
.A(n_1584),
.Y(n_1666)
);

OAI22xp5_ASAP7_75t_L g1667 ( 
.A1(n_1585),
.A2(n_805),
.B1(n_808),
.B2(n_797),
.Y(n_1667)
);

INVx1_ASAP7_75t_L g1668 ( 
.A(n_1499),
.Y(n_1668)
);

INVx2_ASAP7_75t_L g1669 ( 
.A(n_1558),
.Y(n_1669)
);

BUFx6f_ASAP7_75t_L g1670 ( 
.A(n_1507),
.Y(n_1670)
);

AOI22xp5_ASAP7_75t_L g1671 ( 
.A1(n_1577),
.A2(n_820),
.B1(n_822),
.B2(n_819),
.Y(n_1671)
);

INVx1_ASAP7_75t_L g1672 ( 
.A(n_1574),
.Y(n_1672)
);

INVx1_ASAP7_75t_L g1673 ( 
.A(n_1555),
.Y(n_1673)
);

INVx1_ASAP7_75t_L g1674 ( 
.A(n_1497),
.Y(n_1674)
);

INVx1_ASAP7_75t_L g1675 ( 
.A(n_1558),
.Y(n_1675)
);

AND2x2_ASAP7_75t_L g1676 ( 
.A(n_1515),
.B(n_17),
.Y(n_1676)
);

INVx6_ASAP7_75t_L g1677 ( 
.A(n_1491),
.Y(n_1677)
);

INVx1_ASAP7_75t_L g1678 ( 
.A(n_1558),
.Y(n_1678)
);

INVx1_ASAP7_75t_L g1679 ( 
.A(n_1567),
.Y(n_1679)
);

BUFx12f_ASAP7_75t_L g1680 ( 
.A(n_1535),
.Y(n_1680)
);

INVx4_ASAP7_75t_L g1681 ( 
.A(n_1509),
.Y(n_1681)
);

INVx1_ASAP7_75t_L g1682 ( 
.A(n_1567),
.Y(n_1682)
);

CKINVDCx11_ASAP7_75t_R g1683 ( 
.A(n_1519),
.Y(n_1683)
);

CKINVDCx20_ASAP7_75t_R g1684 ( 
.A(n_1508),
.Y(n_1684)
);

INVx1_ASAP7_75t_L g1685 ( 
.A(n_1567),
.Y(n_1685)
);

INVx3_ASAP7_75t_L g1686 ( 
.A(n_1477),
.Y(n_1686)
);

INVx2_ASAP7_75t_L g1687 ( 
.A(n_1510),
.Y(n_1687)
);

INVx1_ASAP7_75t_L g1688 ( 
.A(n_1587),
.Y(n_1688)
);

BUFx6f_ASAP7_75t_L g1689 ( 
.A(n_1488),
.Y(n_1689)
);

BUFx2_ASAP7_75t_SL g1690 ( 
.A(n_1521),
.Y(n_1690)
);

AOI22xp33_ASAP7_75t_L g1691 ( 
.A1(n_1544),
.A2(n_834),
.B1(n_835),
.B2(n_826),
.Y(n_1691)
);

OAI22xp5_ASAP7_75t_L g1692 ( 
.A1(n_1525),
.A2(n_851),
.B1(n_853),
.B2(n_843),
.Y(n_1692)
);

INVx6_ASAP7_75t_L g1693 ( 
.A(n_1494),
.Y(n_1693)
);

OAI22xp5_ASAP7_75t_L g1694 ( 
.A1(n_1586),
.A2(n_860),
.B1(n_867),
.B2(n_854),
.Y(n_1694)
);

BUFx2_ASAP7_75t_L g1695 ( 
.A(n_1526),
.Y(n_1695)
);

BUFx2_ASAP7_75t_SL g1696 ( 
.A(n_1504),
.Y(n_1696)
);

INVx1_ASAP7_75t_L g1697 ( 
.A(n_1552),
.Y(n_1697)
);

CKINVDCx5p33_ASAP7_75t_R g1698 ( 
.A(n_1581),
.Y(n_1698)
);

INVx2_ASAP7_75t_L g1699 ( 
.A(n_1541),
.Y(n_1699)
);

AOI22xp33_ASAP7_75t_SL g1700 ( 
.A1(n_1592),
.A2(n_923),
.B1(n_946),
.B2(n_896),
.Y(n_1700)
);

INVx1_ASAP7_75t_SL g1701 ( 
.A(n_1523),
.Y(n_1701)
);

BUFx8_ASAP7_75t_L g1702 ( 
.A(n_1517),
.Y(n_1702)
);

AOI22xp5_ASAP7_75t_SL g1703 ( 
.A1(n_1576),
.A2(n_878),
.B1(n_884),
.B2(n_875),
.Y(n_1703)
);

INVx6_ASAP7_75t_L g1704 ( 
.A(n_1545),
.Y(n_1704)
);

AOI22xp33_ASAP7_75t_L g1705 ( 
.A1(n_1483),
.A2(n_888),
.B1(n_889),
.B2(n_887),
.Y(n_1705)
);

INVx2_ASAP7_75t_L g1706 ( 
.A(n_1539),
.Y(n_1706)
);

AOI22xp33_ASAP7_75t_L g1707 ( 
.A1(n_1540),
.A2(n_903),
.B1(n_906),
.B2(n_891),
.Y(n_1707)
);

BUFx3_ASAP7_75t_L g1708 ( 
.A(n_1502),
.Y(n_1708)
);

CKINVDCx11_ASAP7_75t_R g1709 ( 
.A(n_1578),
.Y(n_1709)
);

OAI21xp5_ASAP7_75t_SL g1710 ( 
.A1(n_1551),
.A2(n_18),
.B(n_19),
.Y(n_1710)
);

AOI22xp33_ASAP7_75t_SL g1711 ( 
.A1(n_1518),
.A2(n_964),
.B1(n_998),
.B2(n_930),
.Y(n_1711)
);

INVx1_ASAP7_75t_L g1712 ( 
.A(n_1476),
.Y(n_1712)
);

NAND2xp5_ASAP7_75t_L g1713 ( 
.A(n_1480),
.B(n_18),
.Y(n_1713)
);

BUFx2_ASAP7_75t_SL g1714 ( 
.A(n_1489),
.Y(n_1714)
);

OAI21xp33_ASAP7_75t_L g1715 ( 
.A1(n_1480),
.A2(n_1021),
.B(n_1020),
.Y(n_1715)
);

CKINVDCx5p33_ASAP7_75t_R g1716 ( 
.A(n_1478),
.Y(n_1716)
);

NAND2xp5_ASAP7_75t_L g1717 ( 
.A(n_1480),
.B(n_19),
.Y(n_1717)
);

INVx2_ASAP7_75t_SL g1718 ( 
.A(n_1492),
.Y(n_1718)
);

OAI22xp5_ASAP7_75t_L g1719 ( 
.A1(n_1480),
.A2(n_915),
.B1(n_920),
.B2(n_911),
.Y(n_1719)
);

INVx1_ASAP7_75t_L g1720 ( 
.A(n_1476),
.Y(n_1720)
);

AOI22xp33_ASAP7_75t_SL g1721 ( 
.A1(n_1657),
.A2(n_1717),
.B1(n_1713),
.B2(n_1635),
.Y(n_1721)
);

AOI22xp33_ASAP7_75t_L g1722 ( 
.A1(n_1594),
.A2(n_922),
.B1(n_924),
.B2(n_921),
.Y(n_1722)
);

BUFx6f_ASAP7_75t_L g1723 ( 
.A(n_1709),
.Y(n_1723)
);

OAI21xp5_ASAP7_75t_L g1724 ( 
.A1(n_1609),
.A2(n_933),
.B(n_928),
.Y(n_1724)
);

BUFx3_ASAP7_75t_L g1725 ( 
.A(n_1702),
.Y(n_1725)
);

CKINVDCx5p33_ASAP7_75t_R g1726 ( 
.A(n_1618),
.Y(n_1726)
);

OAI22xp5_ASAP7_75t_L g1727 ( 
.A1(n_1626),
.A2(n_940),
.B1(n_947),
.B2(n_931),
.Y(n_1727)
);

AOI22xp33_ASAP7_75t_L g1728 ( 
.A1(n_1715),
.A2(n_951),
.B1(n_961),
.B2(n_937),
.Y(n_1728)
);

CKINVDCx20_ASAP7_75t_R g1729 ( 
.A(n_1614),
.Y(n_1729)
);

OAI22xp5_ASAP7_75t_L g1730 ( 
.A1(n_1603),
.A2(n_979),
.B1(n_992),
.B2(n_972),
.Y(n_1730)
);

OAI22xp5_ASAP7_75t_L g1731 ( 
.A1(n_1611),
.A2(n_994),
.B1(n_997),
.B2(n_974),
.Y(n_1731)
);

BUFx12f_ASAP7_75t_L g1732 ( 
.A(n_1622),
.Y(n_1732)
);

BUFx8_ASAP7_75t_SL g1733 ( 
.A(n_1651),
.Y(n_1733)
);

BUFx2_ASAP7_75t_L g1734 ( 
.A(n_1610),
.Y(n_1734)
);

NAND2xp5_ASAP7_75t_L g1735 ( 
.A(n_1659),
.B(n_20),
.Y(n_1735)
);

INVx2_ASAP7_75t_SL g1736 ( 
.A(n_1595),
.Y(n_1736)
);

AOI211xp5_ASAP7_75t_L g1737 ( 
.A1(n_1637),
.A2(n_1005),
.B(n_1009),
.C(n_993),
.Y(n_1737)
);

INVx1_ASAP7_75t_SL g1738 ( 
.A(n_1701),
.Y(n_1738)
);

OAI22x1_ASAP7_75t_L g1739 ( 
.A1(n_1672),
.A2(n_1024),
.B1(n_1031),
.B2(n_1019),
.Y(n_1739)
);

INVx5_ASAP7_75t_L g1740 ( 
.A(n_1601),
.Y(n_1740)
);

OAI22xp33_ASAP7_75t_L g1741 ( 
.A1(n_1600),
.A2(n_1038),
.B1(n_1041),
.B2(n_1033),
.Y(n_1741)
);

INVx1_ASAP7_75t_L g1742 ( 
.A(n_1605),
.Y(n_1742)
);

INVx2_ASAP7_75t_L g1743 ( 
.A(n_1597),
.Y(n_1743)
);

NAND2xp5_ASAP7_75t_L g1744 ( 
.A(n_1613),
.B(n_21),
.Y(n_1744)
);

AOI22xp33_ASAP7_75t_L g1745 ( 
.A1(n_1608),
.A2(n_1668),
.B1(n_1623),
.B2(n_1598),
.Y(n_1745)
);

INVx1_ASAP7_75t_L g1746 ( 
.A(n_1607),
.Y(n_1746)
);

INVx1_ASAP7_75t_L g1747 ( 
.A(n_1615),
.Y(n_1747)
);

AOI22xp33_ASAP7_75t_L g1748 ( 
.A1(n_1624),
.A2(n_1050),
.B1(n_1055),
.B2(n_1044),
.Y(n_1748)
);

INVx2_ASAP7_75t_L g1749 ( 
.A(n_1602),
.Y(n_1749)
);

INVx1_ASAP7_75t_L g1750 ( 
.A(n_1620),
.Y(n_1750)
);

BUFx6f_ASAP7_75t_L g1751 ( 
.A(n_1596),
.Y(n_1751)
);

AOI22xp33_ASAP7_75t_SL g1752 ( 
.A1(n_1627),
.A2(n_1063),
.B1(n_1066),
.B2(n_1059),
.Y(n_1752)
);

AOI22xp33_ASAP7_75t_SL g1753 ( 
.A1(n_1703),
.A2(n_1067),
.B1(n_23),
.B2(n_24),
.Y(n_1753)
);

INVx2_ASAP7_75t_SL g1754 ( 
.A(n_1612),
.Y(n_1754)
);

AOI22xp33_ASAP7_75t_L g1755 ( 
.A1(n_1629),
.A2(n_23),
.B1(n_21),
.B2(n_22),
.Y(n_1755)
);

AND2x2_ASAP7_75t_L g1756 ( 
.A(n_1676),
.B(n_24),
.Y(n_1756)
);

BUFx4f_ASAP7_75t_SL g1757 ( 
.A(n_1653),
.Y(n_1757)
);

OAI21xp33_ASAP7_75t_L g1758 ( 
.A1(n_1710),
.A2(n_25),
.B(n_26),
.Y(n_1758)
);

INVx1_ASAP7_75t_L g1759 ( 
.A(n_1625),
.Y(n_1759)
);

INVx1_ASAP7_75t_L g1760 ( 
.A(n_1632),
.Y(n_1760)
);

OAI22xp33_ASAP7_75t_L g1761 ( 
.A1(n_1639),
.A2(n_1621),
.B1(n_1641),
.B2(n_1643),
.Y(n_1761)
);

OAI21xp33_ASAP7_75t_L g1762 ( 
.A1(n_1705),
.A2(n_25),
.B(n_26),
.Y(n_1762)
);

AOI22xp33_ASAP7_75t_L g1763 ( 
.A1(n_1674),
.A2(n_29),
.B1(n_27),
.B2(n_28),
.Y(n_1763)
);

INVx1_ASAP7_75t_L g1764 ( 
.A(n_1640),
.Y(n_1764)
);

INVx1_ASAP7_75t_L g1765 ( 
.A(n_1646),
.Y(n_1765)
);

BUFx12f_ASAP7_75t_L g1766 ( 
.A(n_1655),
.Y(n_1766)
);

HB1xp67_ASAP7_75t_L g1767 ( 
.A(n_1647),
.Y(n_1767)
);

INVx1_ASAP7_75t_L g1768 ( 
.A(n_1712),
.Y(n_1768)
);

AOI22xp33_ASAP7_75t_L g1769 ( 
.A1(n_1661),
.A2(n_1666),
.B1(n_1616),
.B2(n_1599),
.Y(n_1769)
);

AOI22xp5_ASAP7_75t_L g1770 ( 
.A1(n_1719),
.A2(n_31),
.B1(n_28),
.B2(n_30),
.Y(n_1770)
);

OAI21xp33_ASAP7_75t_L g1771 ( 
.A1(n_1665),
.A2(n_30),
.B(n_31),
.Y(n_1771)
);

INVx2_ASAP7_75t_L g1772 ( 
.A(n_1720),
.Y(n_1772)
);

AND2x2_ASAP7_75t_L g1773 ( 
.A(n_1628),
.B(n_32),
.Y(n_1773)
);

OAI21xp33_ASAP7_75t_L g1774 ( 
.A1(n_1707),
.A2(n_33),
.B(n_34),
.Y(n_1774)
);

AOI22xp33_ASAP7_75t_L g1775 ( 
.A1(n_1650),
.A2(n_36),
.B1(n_33),
.B2(n_35),
.Y(n_1775)
);

OAI222xp33_ASAP7_75t_L g1776 ( 
.A1(n_1644),
.A2(n_38),
.B1(n_40),
.B2(n_35),
.C1(n_37),
.C2(n_39),
.Y(n_1776)
);

BUFx2_ASAP7_75t_L g1777 ( 
.A(n_1612),
.Y(n_1777)
);

INVx1_ASAP7_75t_L g1778 ( 
.A(n_1673),
.Y(n_1778)
);

INVx2_ASAP7_75t_L g1779 ( 
.A(n_1688),
.Y(n_1779)
);

HB1xp67_ASAP7_75t_L g1780 ( 
.A(n_1695),
.Y(n_1780)
);

AOI21xp33_ASAP7_75t_L g1781 ( 
.A1(n_1687),
.A2(n_37),
.B(n_38),
.Y(n_1781)
);

NAND2xp5_ASAP7_75t_L g1782 ( 
.A(n_1638),
.B(n_39),
.Y(n_1782)
);

BUFx2_ASAP7_75t_L g1783 ( 
.A(n_1718),
.Y(n_1783)
);

AOI22xp5_ASAP7_75t_L g1784 ( 
.A1(n_1642),
.A2(n_42),
.B1(n_40),
.B2(n_41),
.Y(n_1784)
);

OAI22xp5_ASAP7_75t_L g1785 ( 
.A1(n_1634),
.A2(n_43),
.B1(n_41),
.B2(n_42),
.Y(n_1785)
);

NAND2xp5_ASAP7_75t_L g1786 ( 
.A(n_1690),
.B(n_43),
.Y(n_1786)
);

AOI22xp33_ASAP7_75t_L g1787 ( 
.A1(n_1633),
.A2(n_46),
.B1(n_44),
.B2(n_45),
.Y(n_1787)
);

INVx1_ASAP7_75t_L g1788 ( 
.A(n_1669),
.Y(n_1788)
);

AOI22xp33_ASAP7_75t_L g1789 ( 
.A1(n_1699),
.A2(n_47),
.B1(n_44),
.B2(n_46),
.Y(n_1789)
);

OAI22xp5_ASAP7_75t_L g1790 ( 
.A1(n_1671),
.A2(n_1658),
.B1(n_1711),
.B2(n_1660),
.Y(n_1790)
);

AOI22xp33_ASAP7_75t_L g1791 ( 
.A1(n_1706),
.A2(n_1617),
.B1(n_1667),
.B2(n_1694),
.Y(n_1791)
);

AOI22xp33_ASAP7_75t_L g1792 ( 
.A1(n_1656),
.A2(n_49),
.B1(n_47),
.B2(n_48),
.Y(n_1792)
);

OAI21xp33_ASAP7_75t_L g1793 ( 
.A1(n_1700),
.A2(n_48),
.B(n_49),
.Y(n_1793)
);

BUFx6f_ASAP7_75t_SL g1794 ( 
.A(n_1596),
.Y(n_1794)
);

NAND2xp5_ASAP7_75t_SL g1795 ( 
.A(n_1675),
.B(n_50),
.Y(n_1795)
);

AOI22xp33_ASAP7_75t_L g1796 ( 
.A1(n_1645),
.A2(n_52),
.B1(n_50),
.B2(n_51),
.Y(n_1796)
);

AND2x2_ASAP7_75t_L g1797 ( 
.A(n_1696),
.B(n_51),
.Y(n_1797)
);

INVx2_ASAP7_75t_L g1798 ( 
.A(n_1697),
.Y(n_1798)
);

OAI222xp33_ASAP7_75t_L g1799 ( 
.A1(n_1648),
.A2(n_56),
.B1(n_58),
.B2(n_53),
.C1(n_54),
.C2(n_57),
.Y(n_1799)
);

AOI22xp33_ASAP7_75t_L g1800 ( 
.A1(n_1662),
.A2(n_59),
.B1(n_53),
.B2(n_57),
.Y(n_1800)
);

INVx1_ASAP7_75t_L g1801 ( 
.A(n_1678),
.Y(n_1801)
);

INVx2_ASAP7_75t_L g1802 ( 
.A(n_1772),
.Y(n_1802)
);

NAND2xp5_ASAP7_75t_L g1803 ( 
.A(n_1734),
.B(n_1631),
.Y(n_1803)
);

AOI22xp33_ASAP7_75t_L g1804 ( 
.A1(n_1758),
.A2(n_1652),
.B1(n_1683),
.B2(n_1680),
.Y(n_1804)
);

AOI22xp33_ASAP7_75t_L g1805 ( 
.A1(n_1774),
.A2(n_1762),
.B1(n_1771),
.B2(n_1721),
.Y(n_1805)
);

AOI22xp33_ASAP7_75t_SL g1806 ( 
.A1(n_1731),
.A2(n_1790),
.B1(n_1724),
.B2(n_1785),
.Y(n_1806)
);

AOI22xp33_ASAP7_75t_L g1807 ( 
.A1(n_1793),
.A2(n_1682),
.B1(n_1685),
.B2(n_1679),
.Y(n_1807)
);

OAI222xp33_ASAP7_75t_L g1808 ( 
.A1(n_1745),
.A2(n_1663),
.B1(n_1684),
.B2(n_1649),
.C1(n_1698),
.C2(n_1716),
.Y(n_1808)
);

OAI22xp5_ASAP7_75t_L g1809 ( 
.A1(n_1752),
.A2(n_1606),
.B1(n_1708),
.B2(n_1691),
.Y(n_1809)
);

NAND2xp5_ASAP7_75t_L g1810 ( 
.A(n_1767),
.B(n_1714),
.Y(n_1810)
);

NAND2xp5_ASAP7_75t_L g1811 ( 
.A(n_1780),
.B(n_1689),
.Y(n_1811)
);

AOI221xp5_ASAP7_75t_L g1812 ( 
.A1(n_1776),
.A2(n_1692),
.B1(n_1689),
.B2(n_1670),
.C(n_1654),
.Y(n_1812)
);

AOI22xp5_ASAP7_75t_L g1813 ( 
.A1(n_1761),
.A2(n_1593),
.B1(n_1664),
.B2(n_1630),
.Y(n_1813)
);

AOI222xp33_ASAP7_75t_L g1814 ( 
.A1(n_1722),
.A2(n_1630),
.B1(n_1636),
.B2(n_1604),
.C1(n_1670),
.C2(n_1681),
.Y(n_1814)
);

AOI22xp33_ASAP7_75t_L g1815 ( 
.A1(n_1769),
.A2(n_1677),
.B1(n_1619),
.B2(n_1704),
.Y(n_1815)
);

OAI21xp5_ASAP7_75t_SL g1816 ( 
.A1(n_1753),
.A2(n_1686),
.B(n_1619),
.Y(n_1816)
);

AOI22xp5_ASAP7_75t_L g1817 ( 
.A1(n_1784),
.A2(n_1693),
.B1(n_62),
.B2(n_60),
.Y(n_1817)
);

OAI22xp5_ASAP7_75t_L g1818 ( 
.A1(n_1770),
.A2(n_63),
.B1(n_60),
.B2(n_61),
.Y(n_1818)
);

NAND2xp5_ASAP7_75t_L g1819 ( 
.A(n_1742),
.B(n_61),
.Y(n_1819)
);

NAND2xp5_ASAP7_75t_L g1820 ( 
.A(n_1746),
.B(n_63),
.Y(n_1820)
);

AOI22xp33_ASAP7_75t_SL g1821 ( 
.A1(n_1727),
.A2(n_72),
.B1(n_80),
.B2(n_64),
.Y(n_1821)
);

AOI22xp33_ASAP7_75t_L g1822 ( 
.A1(n_1743),
.A2(n_67),
.B1(n_65),
.B2(n_66),
.Y(n_1822)
);

OAI22xp5_ASAP7_75t_L g1823 ( 
.A1(n_1796),
.A2(n_68),
.B1(n_65),
.B2(n_66),
.Y(n_1823)
);

OAI22xp33_ASAP7_75t_L g1824 ( 
.A1(n_1786),
.A2(n_1744),
.B1(n_1782),
.B2(n_1730),
.Y(n_1824)
);

NAND2xp5_ASAP7_75t_L g1825 ( 
.A(n_1747),
.B(n_68),
.Y(n_1825)
);

OAI222xp33_ASAP7_75t_L g1826 ( 
.A1(n_1800),
.A2(n_1787),
.B1(n_1763),
.B2(n_1755),
.C1(n_1775),
.C2(n_1789),
.Y(n_1826)
);

AOI22xp33_ASAP7_75t_SL g1827 ( 
.A1(n_1756),
.A2(n_77),
.B1(n_86),
.B2(n_69),
.Y(n_1827)
);

OAI211xp5_ASAP7_75t_L g1828 ( 
.A1(n_1792),
.A2(n_71),
.B(n_69),
.C(n_70),
.Y(n_1828)
);

NAND2xp5_ASAP7_75t_L g1829 ( 
.A(n_1750),
.B(n_70),
.Y(n_1829)
);

OAI22xp5_ASAP7_75t_L g1830 ( 
.A1(n_1737),
.A2(n_74),
.B1(n_72),
.B2(n_73),
.Y(n_1830)
);

AOI22xp33_ASAP7_75t_L g1831 ( 
.A1(n_1749),
.A2(n_75),
.B1(n_73),
.B2(n_74),
.Y(n_1831)
);

NAND2xp5_ASAP7_75t_L g1832 ( 
.A(n_1759),
.B(n_75),
.Y(n_1832)
);

NAND2xp5_ASAP7_75t_L g1833 ( 
.A(n_1760),
.B(n_76),
.Y(n_1833)
);

OAI22xp5_ASAP7_75t_L g1834 ( 
.A1(n_1791),
.A2(n_1728),
.B1(n_1795),
.B2(n_1783),
.Y(n_1834)
);

AND2x2_ASAP7_75t_L g1835 ( 
.A(n_1773),
.B(n_76),
.Y(n_1835)
);

AOI22xp33_ASAP7_75t_L g1836 ( 
.A1(n_1798),
.A2(n_79),
.B1(n_77),
.B2(n_78),
.Y(n_1836)
);

AOI22xp33_ASAP7_75t_L g1837 ( 
.A1(n_1779),
.A2(n_81),
.B1(n_78),
.B2(n_79),
.Y(n_1837)
);

AOI22xp33_ASAP7_75t_SL g1838 ( 
.A1(n_1797),
.A2(n_91),
.B1(n_103),
.B2(n_82),
.Y(n_1838)
);

NAND3xp33_ASAP7_75t_SL g1839 ( 
.A(n_1729),
.B(n_82),
.C(n_83),
.Y(n_1839)
);

OAI222xp33_ASAP7_75t_L g1840 ( 
.A1(n_1778),
.A2(n_1735),
.B1(n_1764),
.B2(n_1768),
.C1(n_1765),
.C2(n_1738),
.Y(n_1840)
);

AOI22xp33_ASAP7_75t_SL g1841 ( 
.A1(n_1740),
.A2(n_1794),
.B1(n_1723),
.B2(n_1777),
.Y(n_1841)
);

AOI22xp33_ASAP7_75t_L g1842 ( 
.A1(n_1739),
.A2(n_85),
.B1(n_83),
.B2(n_84),
.Y(n_1842)
);

OAI22xp5_ASAP7_75t_L g1843 ( 
.A1(n_1754),
.A2(n_87),
.B1(n_84),
.B2(n_85),
.Y(n_1843)
);

OAI22xp5_ASAP7_75t_L g1844 ( 
.A1(n_1741),
.A2(n_89),
.B1(n_87),
.B2(n_88),
.Y(n_1844)
);

INVx2_ASAP7_75t_L g1845 ( 
.A(n_1788),
.Y(n_1845)
);

OAI22xp5_ASAP7_75t_L g1846 ( 
.A1(n_1723),
.A2(n_90),
.B1(n_88),
.B2(n_89),
.Y(n_1846)
);

CKINVDCx5p33_ASAP7_75t_R g1847 ( 
.A(n_1733),
.Y(n_1847)
);

INVx1_ASAP7_75t_L g1848 ( 
.A(n_1801),
.Y(n_1848)
);

OAI21xp5_ASAP7_75t_SL g1849 ( 
.A1(n_1799),
.A2(n_1723),
.B(n_1781),
.Y(n_1849)
);

AND2x2_ASAP7_75t_L g1850 ( 
.A(n_1751),
.B(n_91),
.Y(n_1850)
);

OAI221xp5_ASAP7_75t_SL g1851 ( 
.A1(n_1849),
.A2(n_1748),
.B1(n_1725),
.B2(n_1736),
.C(n_95),
.Y(n_1851)
);

NAND2xp5_ASAP7_75t_SL g1852 ( 
.A(n_1824),
.B(n_1740),
.Y(n_1852)
);

NAND3xp33_ASAP7_75t_L g1853 ( 
.A(n_1806),
.B(n_1740),
.C(n_1751),
.Y(n_1853)
);

OAI21xp5_ASAP7_75t_SL g1854 ( 
.A1(n_1817),
.A2(n_1757),
.B(n_1726),
.Y(n_1854)
);

NAND2xp5_ASAP7_75t_L g1855 ( 
.A(n_1848),
.B(n_92),
.Y(n_1855)
);

HB1xp67_ASAP7_75t_L g1856 ( 
.A(n_1810),
.Y(n_1856)
);

AND2x2_ASAP7_75t_SL g1857 ( 
.A(n_1805),
.B(n_1732),
.Y(n_1857)
);

NAND2xp5_ASAP7_75t_L g1858 ( 
.A(n_1825),
.B(n_92),
.Y(n_1858)
);

OAI221xp5_ASAP7_75t_SL g1859 ( 
.A1(n_1842),
.A2(n_1827),
.B1(n_1838),
.B2(n_1804),
.C(n_1828),
.Y(n_1859)
);

AOI221xp5_ASAP7_75t_L g1860 ( 
.A1(n_1839),
.A2(n_96),
.B1(n_94),
.B2(n_95),
.C(n_98),
.Y(n_1860)
);

OAI21xp5_ASAP7_75t_SL g1861 ( 
.A1(n_1808),
.A2(n_1809),
.B(n_1846),
.Y(n_1861)
);

AND2x2_ASAP7_75t_L g1862 ( 
.A(n_1803),
.B(n_1766),
.Y(n_1862)
);

INVx1_ASAP7_75t_L g1863 ( 
.A(n_1845),
.Y(n_1863)
);

NAND2xp5_ASAP7_75t_L g1864 ( 
.A(n_1825),
.B(n_94),
.Y(n_1864)
);

NAND2xp5_ASAP7_75t_L g1865 ( 
.A(n_1819),
.B(n_96),
.Y(n_1865)
);

AND2x2_ASAP7_75t_SL g1866 ( 
.A(n_1813),
.B(n_98),
.Y(n_1866)
);

NAND2xp5_ASAP7_75t_L g1867 ( 
.A(n_1820),
.B(n_101),
.Y(n_1867)
);

AOI22xp33_ASAP7_75t_L g1868 ( 
.A1(n_1830),
.A2(n_103),
.B1(n_101),
.B2(n_102),
.Y(n_1868)
);

NAND2xp5_ASAP7_75t_L g1869 ( 
.A(n_1829),
.B(n_102),
.Y(n_1869)
);

AOI221xp5_ASAP7_75t_L g1870 ( 
.A1(n_1818),
.A2(n_106),
.B1(n_104),
.B2(n_105),
.C(n_107),
.Y(n_1870)
);

AND2x2_ASAP7_75t_L g1871 ( 
.A(n_1811),
.B(n_104),
.Y(n_1871)
);

AND2x2_ASAP7_75t_L g1872 ( 
.A(n_1835),
.B(n_105),
.Y(n_1872)
);

AOI22xp33_ASAP7_75t_L g1873 ( 
.A1(n_1807),
.A2(n_109),
.B1(n_106),
.B2(n_108),
.Y(n_1873)
);

NAND3xp33_ASAP7_75t_L g1874 ( 
.A(n_1821),
.B(n_108),
.C(n_109),
.Y(n_1874)
);

NAND2xp5_ASAP7_75t_L g1875 ( 
.A(n_1832),
.B(n_110),
.Y(n_1875)
);

AND2x2_ASAP7_75t_L g1876 ( 
.A(n_1850),
.B(n_1841),
.Y(n_1876)
);

OAI211xp5_ASAP7_75t_SL g1877 ( 
.A1(n_1833),
.A2(n_112),
.B(n_110),
.C(n_111),
.Y(n_1877)
);

NAND3xp33_ASAP7_75t_L g1878 ( 
.A(n_1844),
.B(n_111),
.C(n_113),
.Y(n_1878)
);

OAI21xp5_ASAP7_75t_SL g1879 ( 
.A1(n_1816),
.A2(n_113),
.B(n_114),
.Y(n_1879)
);

NAND3xp33_ASAP7_75t_L g1880 ( 
.A(n_1836),
.B(n_115),
.C(n_116),
.Y(n_1880)
);

NAND2xp5_ASAP7_75t_L g1881 ( 
.A(n_1802),
.B(n_115),
.Y(n_1881)
);

OAI21xp33_ASAP7_75t_L g1882 ( 
.A1(n_1837),
.A2(n_1831),
.B(n_1822),
.Y(n_1882)
);

AND2x2_ASAP7_75t_L g1883 ( 
.A(n_1814),
.B(n_116),
.Y(n_1883)
);

AND2x2_ASAP7_75t_L g1884 ( 
.A(n_1834),
.B(n_118),
.Y(n_1884)
);

NAND4xp25_ASAP7_75t_L g1885 ( 
.A(n_1843),
.B(n_1823),
.C(n_1812),
.D(n_1815),
.Y(n_1885)
);

NAND2xp5_ASAP7_75t_SL g1886 ( 
.A(n_1847),
.B(n_118),
.Y(n_1886)
);

OAI21xp5_ASAP7_75t_SL g1887 ( 
.A1(n_1826),
.A2(n_119),
.B(n_120),
.Y(n_1887)
);

OAI211xp5_ASAP7_75t_L g1888 ( 
.A1(n_1840),
.A2(n_121),
.B(n_119),
.C(n_120),
.Y(n_1888)
);

NAND3xp33_ASAP7_75t_L g1889 ( 
.A(n_1806),
.B(n_121),
.C(n_122),
.Y(n_1889)
);

OAI221xp5_ASAP7_75t_L g1890 ( 
.A1(n_1806),
.A2(n_124),
.B1(n_122),
.B2(n_123),
.C(n_125),
.Y(n_1890)
);

AND2x2_ASAP7_75t_L g1891 ( 
.A(n_1803),
.B(n_123),
.Y(n_1891)
);

OAI21xp33_ASAP7_75t_SL g1892 ( 
.A1(n_1810),
.A2(n_132),
.B(n_124),
.Y(n_1892)
);

OAI21xp5_ASAP7_75t_SL g1893 ( 
.A1(n_1806),
.A2(n_125),
.B(n_126),
.Y(n_1893)
);

NAND2xp5_ASAP7_75t_L g1894 ( 
.A(n_1848),
.B(n_126),
.Y(n_1894)
);

OAI221xp5_ASAP7_75t_L g1895 ( 
.A1(n_1806),
.A2(n_129),
.B1(n_127),
.B2(n_128),
.C(n_130),
.Y(n_1895)
);

OAI21xp33_ASAP7_75t_SL g1896 ( 
.A1(n_1825),
.A2(n_127),
.B(n_129),
.Y(n_1896)
);

AND2x2_ASAP7_75t_L g1897 ( 
.A(n_1803),
.B(n_130),
.Y(n_1897)
);

AND2x2_ASAP7_75t_L g1898 ( 
.A(n_1803),
.B(n_131),
.Y(n_1898)
);

INVx1_ASAP7_75t_L g1899 ( 
.A(n_1848),
.Y(n_1899)
);

AND2x2_ASAP7_75t_L g1900 ( 
.A(n_1803),
.B(n_131),
.Y(n_1900)
);

NAND2xp5_ASAP7_75t_L g1901 ( 
.A(n_1848),
.B(n_132),
.Y(n_1901)
);

AO21x2_ASAP7_75t_L g1902 ( 
.A1(n_1881),
.A2(n_133),
.B(n_134),
.Y(n_1902)
);

NAND2x1_ASAP7_75t_L g1903 ( 
.A(n_1899),
.B(n_133),
.Y(n_1903)
);

INVx3_ASAP7_75t_L g1904 ( 
.A(n_1863),
.Y(n_1904)
);

NAND3xp33_ASAP7_75t_L g1905 ( 
.A(n_1889),
.B(n_134),
.C(n_135),
.Y(n_1905)
);

AOI22xp33_ASAP7_75t_L g1906 ( 
.A1(n_1882),
.A2(n_138),
.B1(n_136),
.B2(n_137),
.Y(n_1906)
);

NOR3xp33_ASAP7_75t_L g1907 ( 
.A(n_1879),
.B(n_136),
.C(n_138),
.Y(n_1907)
);

OR2x2_ASAP7_75t_L g1908 ( 
.A(n_1856),
.B(n_139),
.Y(n_1908)
);

BUFx3_ASAP7_75t_L g1909 ( 
.A(n_1862),
.Y(n_1909)
);

OR2x2_ASAP7_75t_L g1910 ( 
.A(n_1855),
.B(n_139),
.Y(n_1910)
);

NOR3xp33_ASAP7_75t_L g1911 ( 
.A(n_1893),
.B(n_1887),
.C(n_1861),
.Y(n_1911)
);

AND2x2_ASAP7_75t_L g1912 ( 
.A(n_1876),
.B(n_140),
.Y(n_1912)
);

OR2x2_ASAP7_75t_L g1913 ( 
.A(n_1894),
.B(n_1901),
.Y(n_1913)
);

NAND3xp33_ASAP7_75t_L g1914 ( 
.A(n_1896),
.B(n_141),
.C(n_142),
.Y(n_1914)
);

OR2x2_ASAP7_75t_L g1915 ( 
.A(n_1858),
.B(n_141),
.Y(n_1915)
);

OR2x2_ASAP7_75t_L g1916 ( 
.A(n_1864),
.B(n_143),
.Y(n_1916)
);

INVx1_ASAP7_75t_L g1917 ( 
.A(n_1865),
.Y(n_1917)
);

INVx1_ASAP7_75t_L g1918 ( 
.A(n_1867),
.Y(n_1918)
);

AOI221xp5_ASAP7_75t_L g1919 ( 
.A1(n_1896),
.A2(n_145),
.B1(n_143),
.B2(n_144),
.C(n_146),
.Y(n_1919)
);

INVx1_ASAP7_75t_L g1920 ( 
.A(n_1869),
.Y(n_1920)
);

AOI21x1_ASAP7_75t_L g1921 ( 
.A1(n_1852),
.A2(n_145),
.B(n_146),
.Y(n_1921)
);

NAND3xp33_ASAP7_75t_L g1922 ( 
.A(n_1860),
.B(n_147),
.C(n_148),
.Y(n_1922)
);

NAND2xp5_ASAP7_75t_L g1923 ( 
.A(n_1884),
.B(n_147),
.Y(n_1923)
);

NOR3xp33_ASAP7_75t_L g1924 ( 
.A(n_1890),
.B(n_148),
.C(n_149),
.Y(n_1924)
);

INVx2_ASAP7_75t_L g1925 ( 
.A(n_1871),
.Y(n_1925)
);

AOI22xp5_ASAP7_75t_L g1926 ( 
.A1(n_1853),
.A2(n_153),
.B1(n_150),
.B2(n_152),
.Y(n_1926)
);

AOI22xp33_ASAP7_75t_L g1927 ( 
.A1(n_1885),
.A2(n_153),
.B1(n_150),
.B2(n_152),
.Y(n_1927)
);

AOI22xp5_ASAP7_75t_L g1928 ( 
.A1(n_1888),
.A2(n_156),
.B1(n_154),
.B2(n_155),
.Y(n_1928)
);

NOR2xp33_ASAP7_75t_L g1929 ( 
.A(n_1886),
.B(n_154),
.Y(n_1929)
);

AND2x2_ASAP7_75t_L g1930 ( 
.A(n_1891),
.B(n_156),
.Y(n_1930)
);

AND2x2_ASAP7_75t_L g1931 ( 
.A(n_1897),
.B(n_157),
.Y(n_1931)
);

NOR3xp33_ASAP7_75t_L g1932 ( 
.A(n_1895),
.B(n_157),
.C(n_158),
.Y(n_1932)
);

NAND2xp5_ASAP7_75t_L g1933 ( 
.A(n_1875),
.B(n_158),
.Y(n_1933)
);

INVx1_ASAP7_75t_L g1934 ( 
.A(n_1900),
.Y(n_1934)
);

NAND2xp5_ASAP7_75t_L g1935 ( 
.A(n_1898),
.B(n_159),
.Y(n_1935)
);

NAND2xp5_ASAP7_75t_L g1936 ( 
.A(n_1872),
.B(n_159),
.Y(n_1936)
);

INVx1_ASAP7_75t_L g1937 ( 
.A(n_1877),
.Y(n_1937)
);

NOR2xp33_ASAP7_75t_L g1938 ( 
.A(n_1854),
.B(n_160),
.Y(n_1938)
);

NOR4xp75_ASAP7_75t_L g1939 ( 
.A(n_1883),
.B(n_162),
.C(n_160),
.D(n_161),
.Y(n_1939)
);

AND2x2_ASAP7_75t_L g1940 ( 
.A(n_1857),
.B(n_162),
.Y(n_1940)
);

NOR2x1p5_ASAP7_75t_L g1941 ( 
.A(n_1878),
.B(n_1874),
.Y(n_1941)
);

NOR2xp33_ASAP7_75t_L g1942 ( 
.A(n_1866),
.B(n_163),
.Y(n_1942)
);

NAND3xp33_ASAP7_75t_L g1943 ( 
.A(n_1870),
.B(n_164),
.C(n_165),
.Y(n_1943)
);

NOR3xp33_ASAP7_75t_L g1944 ( 
.A(n_1851),
.B(n_164),
.C(n_166),
.Y(n_1944)
);

BUFx3_ASAP7_75t_L g1945 ( 
.A(n_1880),
.Y(n_1945)
);

AOI211xp5_ASAP7_75t_L g1946 ( 
.A1(n_1892),
.A2(n_168),
.B(n_166),
.C(n_167),
.Y(n_1946)
);

NOR3xp33_ASAP7_75t_L g1947 ( 
.A(n_1859),
.B(n_167),
.C(n_168),
.Y(n_1947)
);

NAND3xp33_ASAP7_75t_L g1948 ( 
.A(n_1868),
.B(n_169),
.C(n_170),
.Y(n_1948)
);

NAND2xp5_ASAP7_75t_L g1949 ( 
.A(n_1873),
.B(n_170),
.Y(n_1949)
);

OR2x2_ASAP7_75t_L g1950 ( 
.A(n_1856),
.B(n_171),
.Y(n_1950)
);

NAND2x1_ASAP7_75t_L g1951 ( 
.A(n_1899),
.B(n_171),
.Y(n_1951)
);

OAI211xp5_ASAP7_75t_SL g1952 ( 
.A1(n_1886),
.A2(n_176),
.B(n_173),
.C(n_174),
.Y(n_1952)
);

NAND3xp33_ASAP7_75t_L g1953 ( 
.A(n_1889),
.B(n_173),
.C(n_174),
.Y(n_1953)
);

INVx1_ASAP7_75t_L g1954 ( 
.A(n_1899),
.Y(n_1954)
);

NOR3xp33_ASAP7_75t_SL g1955 ( 
.A(n_1854),
.B(n_176),
.C(n_178),
.Y(n_1955)
);

INVx1_ASAP7_75t_L g1956 ( 
.A(n_1899),
.Y(n_1956)
);

NAND2xp33_ASAP7_75t_R g1957 ( 
.A(n_1876),
.B(n_178),
.Y(n_1957)
);

AND2x2_ASAP7_75t_L g1958 ( 
.A(n_1856),
.B(n_179),
.Y(n_1958)
);

OR2x2_ASAP7_75t_L g1959 ( 
.A(n_1856),
.B(n_180),
.Y(n_1959)
);

NAND2xp5_ASAP7_75t_L g1960 ( 
.A(n_1856),
.B(n_180),
.Y(n_1960)
);

OR2x2_ASAP7_75t_L g1961 ( 
.A(n_1856),
.B(n_181),
.Y(n_1961)
);

OAI211xp5_ASAP7_75t_SL g1962 ( 
.A1(n_1886),
.A2(n_183),
.B(n_181),
.C(n_182),
.Y(n_1962)
);

INVx1_ASAP7_75t_L g1963 ( 
.A(n_1899),
.Y(n_1963)
);

OAI211xp5_ASAP7_75t_SL g1964 ( 
.A1(n_1886),
.A2(n_185),
.B(n_183),
.C(n_184),
.Y(n_1964)
);

AND2x2_ASAP7_75t_L g1965 ( 
.A(n_1856),
.B(n_184),
.Y(n_1965)
);

NAND4xp75_ASAP7_75t_L g1966 ( 
.A(n_1857),
.B(n_187),
.C(n_185),
.D(n_186),
.Y(n_1966)
);

INVx2_ASAP7_75t_L g1967 ( 
.A(n_1863),
.Y(n_1967)
);

INVx2_ASAP7_75t_L g1968 ( 
.A(n_1863),
.Y(n_1968)
);

NAND4xp75_ASAP7_75t_L g1969 ( 
.A(n_1857),
.B(n_188),
.C(n_186),
.D(n_187),
.Y(n_1969)
);

NOR3xp33_ASAP7_75t_L g1970 ( 
.A(n_1889),
.B(n_188),
.C(n_189),
.Y(n_1970)
);

NAND2xp5_ASAP7_75t_L g1971 ( 
.A(n_1856),
.B(n_190),
.Y(n_1971)
);

INVx1_ASAP7_75t_L g1972 ( 
.A(n_1899),
.Y(n_1972)
);

NOR2xp33_ASAP7_75t_L g1973 ( 
.A(n_1856),
.B(n_190),
.Y(n_1973)
);

OAI21xp5_ASAP7_75t_L g1974 ( 
.A1(n_1887),
.A2(n_191),
.B(n_192),
.Y(n_1974)
);

XNOR2x2_ASAP7_75t_L g1975 ( 
.A(n_1974),
.B(n_191),
.Y(n_1975)
);

XNOR2x2_ASAP7_75t_L g1976 ( 
.A(n_1957),
.B(n_192),
.Y(n_1976)
);

XOR2x2_ASAP7_75t_L g1977 ( 
.A(n_1911),
.B(n_193),
.Y(n_1977)
);

AND2x2_ASAP7_75t_L g1978 ( 
.A(n_1909),
.B(n_193),
.Y(n_1978)
);

NAND3xp33_ASAP7_75t_L g1979 ( 
.A(n_1947),
.B(n_194),
.C(n_195),
.Y(n_1979)
);

NAND4xp75_ASAP7_75t_L g1980 ( 
.A(n_1942),
.B(n_196),
.C(n_194),
.D(n_195),
.Y(n_1980)
);

NAND2xp5_ASAP7_75t_L g1981 ( 
.A(n_1917),
.B(n_1918),
.Y(n_1981)
);

NAND2xp5_ASAP7_75t_L g1982 ( 
.A(n_1920),
.B(n_196),
.Y(n_1982)
);

NAND2xp5_ASAP7_75t_L g1983 ( 
.A(n_1904),
.B(n_1913),
.Y(n_1983)
);

INVx1_ASAP7_75t_SL g1984 ( 
.A(n_1908),
.Y(n_1984)
);

INVx1_ASAP7_75t_L g1985 ( 
.A(n_1954),
.Y(n_1985)
);

INVx1_ASAP7_75t_L g1986 ( 
.A(n_1956),
.Y(n_1986)
);

INVx2_ASAP7_75t_L g1987 ( 
.A(n_1904),
.Y(n_1987)
);

NOR2xp33_ASAP7_75t_L g1988 ( 
.A(n_1933),
.B(n_197),
.Y(n_1988)
);

NAND2xp5_ASAP7_75t_L g1989 ( 
.A(n_1963),
.B(n_198),
.Y(n_1989)
);

INVx1_ASAP7_75t_L g1990 ( 
.A(n_1972),
.Y(n_1990)
);

INVx1_ASAP7_75t_L g1991 ( 
.A(n_1967),
.Y(n_1991)
);

AOI22xp5_ASAP7_75t_L g1992 ( 
.A1(n_1907),
.A2(n_201),
.B1(n_199),
.B2(n_200),
.Y(n_1992)
);

CKINVDCx8_ASAP7_75t_R g1993 ( 
.A(n_1973),
.Y(n_1993)
);

AND2x2_ASAP7_75t_L g1994 ( 
.A(n_1934),
.B(n_199),
.Y(n_1994)
);

INVx2_ASAP7_75t_L g1995 ( 
.A(n_1968),
.Y(n_1995)
);

INVx2_ASAP7_75t_L g1996 ( 
.A(n_1950),
.Y(n_1996)
);

INVx2_ASAP7_75t_L g1997 ( 
.A(n_1959),
.Y(n_1997)
);

INVx4_ASAP7_75t_L g1998 ( 
.A(n_1958),
.Y(n_1998)
);

XNOR2xp5_ASAP7_75t_L g1999 ( 
.A(n_1939),
.B(n_202),
.Y(n_1999)
);

NOR2x1_ASAP7_75t_L g2000 ( 
.A(n_1961),
.B(n_1960),
.Y(n_2000)
);

AND2x2_ASAP7_75t_L g2001 ( 
.A(n_1925),
.B(n_1965),
.Y(n_2001)
);

BUFx6f_ASAP7_75t_L g2002 ( 
.A(n_1903),
.Y(n_2002)
);

INVx2_ASAP7_75t_SL g2003 ( 
.A(n_1971),
.Y(n_2003)
);

NAND3xp33_ASAP7_75t_L g2004 ( 
.A(n_1924),
.B(n_202),
.C(n_204),
.Y(n_2004)
);

NOR3xp33_ASAP7_75t_L g2005 ( 
.A(n_1905),
.B(n_205),
.C(n_206),
.Y(n_2005)
);

INVx1_ASAP7_75t_L g2006 ( 
.A(n_1902),
.Y(n_2006)
);

NOR3xp33_ASAP7_75t_L g2007 ( 
.A(n_1953),
.B(n_206),
.C(n_207),
.Y(n_2007)
);

INVx1_ASAP7_75t_L g2008 ( 
.A(n_1910),
.Y(n_2008)
);

NAND2xp5_ASAP7_75t_L g2009 ( 
.A(n_1945),
.B(n_1937),
.Y(n_2009)
);

INVx2_ASAP7_75t_L g2010 ( 
.A(n_1951),
.Y(n_2010)
);

INVx2_ASAP7_75t_L g2011 ( 
.A(n_1912),
.Y(n_2011)
);

INVx1_ASAP7_75t_L g2012 ( 
.A(n_1915),
.Y(n_2012)
);

INVx2_ASAP7_75t_SL g2013 ( 
.A(n_1916),
.Y(n_2013)
);

NAND2xp5_ASAP7_75t_L g2014 ( 
.A(n_1923),
.B(n_207),
.Y(n_2014)
);

AND2x4_ASAP7_75t_L g2015 ( 
.A(n_1940),
.B(n_208),
.Y(n_2015)
);

INVx1_ASAP7_75t_L g2016 ( 
.A(n_1914),
.Y(n_2016)
);

INVx2_ASAP7_75t_L g2017 ( 
.A(n_1921),
.Y(n_2017)
);

INVx2_ASAP7_75t_SL g2018 ( 
.A(n_1930),
.Y(n_2018)
);

NOR3xp33_ASAP7_75t_L g2019 ( 
.A(n_1938),
.B(n_208),
.C(n_209),
.Y(n_2019)
);

AND2x2_ASAP7_75t_L g2020 ( 
.A(n_1931),
.B(n_211),
.Y(n_2020)
);

AND2x4_ASAP7_75t_L g2021 ( 
.A(n_1941),
.B(n_1955),
.Y(n_2021)
);

AND2x2_ASAP7_75t_L g2022 ( 
.A(n_1936),
.B(n_212),
.Y(n_2022)
);

NAND2xp5_ASAP7_75t_L g2023 ( 
.A(n_1935),
.B(n_212),
.Y(n_2023)
);

INVx2_ASAP7_75t_SL g2024 ( 
.A(n_1949),
.Y(n_2024)
);

XOR2x2_ASAP7_75t_L g2025 ( 
.A(n_1966),
.B(n_213),
.Y(n_2025)
);

INVx1_ASAP7_75t_L g2026 ( 
.A(n_1926),
.Y(n_2026)
);

INVx1_ASAP7_75t_L g2027 ( 
.A(n_1929),
.Y(n_2027)
);

XNOR2xp5_ASAP7_75t_L g2028 ( 
.A(n_1969),
.B(n_213),
.Y(n_2028)
);

NAND4xp75_ASAP7_75t_SL g2029 ( 
.A(n_1952),
.B(n_216),
.C(n_214),
.D(n_215),
.Y(n_2029)
);

NAND3xp33_ASAP7_75t_SL g2030 ( 
.A(n_1946),
.B(n_214),
.C(n_217),
.Y(n_2030)
);

INVx3_ASAP7_75t_L g2031 ( 
.A(n_1962),
.Y(n_2031)
);

NOR2xp33_ASAP7_75t_L g2032 ( 
.A(n_1964),
.B(n_217),
.Y(n_2032)
);

NAND4xp75_ASAP7_75t_L g2033 ( 
.A(n_1928),
.B(n_221),
.C(n_218),
.D(n_220),
.Y(n_2033)
);

NAND4xp75_ASAP7_75t_L g2034 ( 
.A(n_1919),
.B(n_222),
.C(n_218),
.D(n_221),
.Y(n_2034)
);

OR2x2_ASAP7_75t_L g2035 ( 
.A(n_1922),
.B(n_222),
.Y(n_2035)
);

HB1xp67_ASAP7_75t_L g2036 ( 
.A(n_1970),
.Y(n_2036)
);

INVx1_ASAP7_75t_L g2037 ( 
.A(n_1943),
.Y(n_2037)
);

OR2x2_ASAP7_75t_L g2038 ( 
.A(n_1906),
.B(n_223),
.Y(n_2038)
);

NAND2xp5_ASAP7_75t_L g2039 ( 
.A(n_1932),
.B(n_223),
.Y(n_2039)
);

BUFx2_ASAP7_75t_L g2040 ( 
.A(n_1948),
.Y(n_2040)
);

OAI22xp33_ASAP7_75t_SL g2041 ( 
.A1(n_1944),
.A2(n_1927),
.B1(n_226),
.B2(n_224),
.Y(n_2041)
);

AND2x4_ASAP7_75t_L g2042 ( 
.A(n_1909),
.B(n_225),
.Y(n_2042)
);

NAND4xp75_ASAP7_75t_SL g2043 ( 
.A(n_1938),
.B(n_229),
.C(n_227),
.D(n_228),
.Y(n_2043)
);

NAND2xp5_ASAP7_75t_L g2044 ( 
.A(n_1917),
.B(n_228),
.Y(n_2044)
);

NAND4xp75_ASAP7_75t_L g2045 ( 
.A(n_1974),
.B(n_232),
.C(n_229),
.D(n_230),
.Y(n_2045)
);

INVx1_ASAP7_75t_L g2046 ( 
.A(n_1954),
.Y(n_2046)
);

AND2x2_ASAP7_75t_L g2047 ( 
.A(n_1909),
.B(n_230),
.Y(n_2047)
);

XNOR2xp5_ASAP7_75t_L g2048 ( 
.A(n_1930),
.B(n_232),
.Y(n_2048)
);

NAND4xp75_ASAP7_75t_L g2049 ( 
.A(n_1974),
.B(n_235),
.C(n_233),
.D(n_234),
.Y(n_2049)
);

INVx2_ASAP7_75t_L g2050 ( 
.A(n_1904),
.Y(n_2050)
);

NAND4xp75_ASAP7_75t_L g2051 ( 
.A(n_1974),
.B(n_235),
.C(n_233),
.D(n_234),
.Y(n_2051)
);

AND2x2_ASAP7_75t_L g2052 ( 
.A(n_1909),
.B(n_236),
.Y(n_2052)
);

XOR2x2_ASAP7_75t_L g2053 ( 
.A(n_1911),
.B(n_236),
.Y(n_2053)
);

AND2x2_ASAP7_75t_L g2054 ( 
.A(n_1909),
.B(n_237),
.Y(n_2054)
);

XOR2x2_ASAP7_75t_L g2055 ( 
.A(n_1911),
.B(n_237),
.Y(n_2055)
);

OR2x2_ASAP7_75t_L g2056 ( 
.A(n_1904),
.B(n_238),
.Y(n_2056)
);

INVx1_ASAP7_75t_L g2057 ( 
.A(n_1954),
.Y(n_2057)
);

INVx2_ASAP7_75t_L g2058 ( 
.A(n_1904),
.Y(n_2058)
);

INVx2_ASAP7_75t_SL g2059 ( 
.A(n_1909),
.Y(n_2059)
);

INVxp67_ASAP7_75t_SL g2060 ( 
.A(n_1904),
.Y(n_2060)
);

INVxp67_ASAP7_75t_SL g2061 ( 
.A(n_1904),
.Y(n_2061)
);

INVx2_ASAP7_75t_L g2062 ( 
.A(n_1904),
.Y(n_2062)
);

XNOR2xp5_ASAP7_75t_L g2063 ( 
.A(n_1930),
.B(n_239),
.Y(n_2063)
);

NAND4xp75_ASAP7_75t_L g2064 ( 
.A(n_1974),
.B(n_241),
.C(n_239),
.D(n_240),
.Y(n_2064)
);

NOR3xp33_ASAP7_75t_L g2065 ( 
.A(n_1911),
.B(n_240),
.C(n_241),
.Y(n_2065)
);

AND2x2_ASAP7_75t_L g2066 ( 
.A(n_1909),
.B(n_242),
.Y(n_2066)
);

AND2x2_ASAP7_75t_L g2067 ( 
.A(n_1909),
.B(n_242),
.Y(n_2067)
);

OAI22xp5_ASAP7_75t_L g2068 ( 
.A1(n_1911),
.A2(n_245),
.B1(n_243),
.B2(n_244),
.Y(n_2068)
);

INVx2_ASAP7_75t_L g2069 ( 
.A(n_1904),
.Y(n_2069)
);

INVx1_ASAP7_75t_L g2070 ( 
.A(n_1985),
.Y(n_2070)
);

AOI22x1_ASAP7_75t_SL g2071 ( 
.A1(n_2037),
.A2(n_246),
.B1(n_243),
.B2(n_245),
.Y(n_2071)
);

XNOR2x2_ASAP7_75t_L g2072 ( 
.A(n_1976),
.B(n_246),
.Y(n_2072)
);

NOR2x1_ASAP7_75t_L g2073 ( 
.A(n_2009),
.B(n_247),
.Y(n_2073)
);

INVx1_ASAP7_75t_L g2074 ( 
.A(n_1986),
.Y(n_2074)
);

INVx1_ASAP7_75t_SL g2075 ( 
.A(n_1984),
.Y(n_2075)
);

INVx1_ASAP7_75t_L g2076 ( 
.A(n_1990),
.Y(n_2076)
);

AOI22xp5_ASAP7_75t_L g2077 ( 
.A1(n_2019),
.A2(n_249),
.B1(n_247),
.B2(n_248),
.Y(n_2077)
);

INVx1_ASAP7_75t_L g2078 ( 
.A(n_2046),
.Y(n_2078)
);

CKINVDCx8_ASAP7_75t_R g2079 ( 
.A(n_2042),
.Y(n_2079)
);

AOI22xp33_ASAP7_75t_SL g2080 ( 
.A1(n_1975),
.A2(n_256),
.B1(n_266),
.B2(n_248),
.Y(n_2080)
);

AND2x2_ASAP7_75t_L g2081 ( 
.A(n_2059),
.B(n_249),
.Y(n_2081)
);

OA22x2_ASAP7_75t_L g2082 ( 
.A1(n_2015),
.A2(n_252),
.B1(n_250),
.B2(n_251),
.Y(n_2082)
);

INVxp67_ASAP7_75t_L g2083 ( 
.A(n_2036),
.Y(n_2083)
);

INVx1_ASAP7_75t_L g2084 ( 
.A(n_2057),
.Y(n_2084)
);

AND2x2_ASAP7_75t_L g2085 ( 
.A(n_1998),
.B(n_250),
.Y(n_2085)
);

AOI22xp5_ASAP7_75t_L g2086 ( 
.A1(n_2030),
.A2(n_254),
.B1(n_252),
.B2(n_253),
.Y(n_2086)
);

XNOR2xp5_ASAP7_75t_L g2087 ( 
.A(n_2048),
.B(n_2063),
.Y(n_2087)
);

XNOR2xp5_ASAP7_75t_L g2088 ( 
.A(n_1977),
.B(n_253),
.Y(n_2088)
);

INVx1_ASAP7_75t_L g2089 ( 
.A(n_1981),
.Y(n_2089)
);

XNOR2xp5_ASAP7_75t_L g2090 ( 
.A(n_2053),
.B(n_254),
.Y(n_2090)
);

INVx1_ASAP7_75t_L g2091 ( 
.A(n_2006),
.Y(n_2091)
);

AND2x2_ASAP7_75t_L g2092 ( 
.A(n_2018),
.B(n_2060),
.Y(n_2092)
);

INVx2_ASAP7_75t_L g2093 ( 
.A(n_2010),
.Y(n_2093)
);

XOR2x2_ASAP7_75t_L g2094 ( 
.A(n_2055),
.B(n_2025),
.Y(n_2094)
);

OA22x2_ASAP7_75t_L g2095 ( 
.A1(n_2040),
.A2(n_2016),
.B1(n_2024),
.B2(n_2003),
.Y(n_2095)
);

INVx1_ASAP7_75t_L g2096 ( 
.A(n_1991),
.Y(n_2096)
);

XNOR2xp5_ASAP7_75t_L g2097 ( 
.A(n_1999),
.B(n_255),
.Y(n_2097)
);

INVxp67_ASAP7_75t_L g2098 ( 
.A(n_2021),
.Y(n_2098)
);

OA22x2_ASAP7_75t_L g2099 ( 
.A1(n_2027),
.A2(n_260),
.B1(n_257),
.B2(n_258),
.Y(n_2099)
);

XNOR2xp5_ASAP7_75t_L g2100 ( 
.A(n_1999),
.B(n_2028),
.Y(n_2100)
);

AND2x2_ASAP7_75t_L g2101 ( 
.A(n_2061),
.B(n_257),
.Y(n_2101)
);

XNOR2x2_ASAP7_75t_L g2102 ( 
.A(n_2000),
.B(n_258),
.Y(n_2102)
);

INVx1_ASAP7_75t_SL g2103 ( 
.A(n_2001),
.Y(n_2103)
);

XOR2x2_ASAP7_75t_L g2104 ( 
.A(n_1980),
.B(n_260),
.Y(n_2104)
);

XNOR2xp5_ASAP7_75t_L g2105 ( 
.A(n_2020),
.B(n_261),
.Y(n_2105)
);

INVx2_ASAP7_75t_L g2106 ( 
.A(n_1995),
.Y(n_2106)
);

AO22x2_ASAP7_75t_L g2107 ( 
.A1(n_1996),
.A2(n_264),
.B1(n_262),
.B2(n_263),
.Y(n_2107)
);

OA22x2_ASAP7_75t_L g2108 ( 
.A1(n_2011),
.A2(n_266),
.B1(n_263),
.B2(n_264),
.Y(n_2108)
);

INVx1_ASAP7_75t_L g2109 ( 
.A(n_1983),
.Y(n_2109)
);

INVx1_ASAP7_75t_L g2110 ( 
.A(n_2012),
.Y(n_2110)
);

NOR2xp33_ASAP7_75t_R g2111 ( 
.A(n_1993),
.B(n_267),
.Y(n_2111)
);

INVxp67_ASAP7_75t_L g2112 ( 
.A(n_1988),
.Y(n_2112)
);

CKINVDCx16_ASAP7_75t_R g2113 ( 
.A(n_1978),
.Y(n_2113)
);

XOR2x2_ASAP7_75t_L g2114 ( 
.A(n_2045),
.B(n_268),
.Y(n_2114)
);

INVx1_ASAP7_75t_L g2115 ( 
.A(n_1989),
.Y(n_2115)
);

XNOR2xp5_ASAP7_75t_L g2116 ( 
.A(n_2047),
.B(n_268),
.Y(n_2116)
);

OAI22xp5_ASAP7_75t_L g2117 ( 
.A1(n_1992),
.A2(n_271),
.B1(n_269),
.B2(n_270),
.Y(n_2117)
);

INVx1_ASAP7_75t_L g2118 ( 
.A(n_2008),
.Y(n_2118)
);

INVx1_ASAP7_75t_L g2119 ( 
.A(n_1997),
.Y(n_2119)
);

INVx1_ASAP7_75t_L g2120 ( 
.A(n_2056),
.Y(n_2120)
);

XOR2xp5_ASAP7_75t_L g2121 ( 
.A(n_2043),
.B(n_269),
.Y(n_2121)
);

XOR2x2_ASAP7_75t_L g2122 ( 
.A(n_2049),
.B(n_270),
.Y(n_2122)
);

OR2x2_ASAP7_75t_L g2123 ( 
.A(n_2013),
.B(n_271),
.Y(n_2123)
);

INVx2_ASAP7_75t_SL g2124 ( 
.A(n_2052),
.Y(n_2124)
);

XOR2x2_ASAP7_75t_L g2125 ( 
.A(n_2051),
.B(n_272),
.Y(n_2125)
);

INVx1_ASAP7_75t_L g2126 ( 
.A(n_1982),
.Y(n_2126)
);

NAND2xp5_ASAP7_75t_L g2127 ( 
.A(n_1987),
.B(n_273),
.Y(n_2127)
);

INVx1_ASAP7_75t_L g2128 ( 
.A(n_2044),
.Y(n_2128)
);

OAI22xp5_ASAP7_75t_L g2129 ( 
.A1(n_2004),
.A2(n_276),
.B1(n_274),
.B2(n_275),
.Y(n_2129)
);

INVx1_ASAP7_75t_L g2130 ( 
.A(n_2050),
.Y(n_2130)
);

INVx1_ASAP7_75t_L g2131 ( 
.A(n_2058),
.Y(n_2131)
);

OA22x2_ASAP7_75t_L g2132 ( 
.A1(n_2026),
.A2(n_278),
.B1(n_275),
.B2(n_277),
.Y(n_2132)
);

XOR2x2_ASAP7_75t_L g2133 ( 
.A(n_2064),
.B(n_278),
.Y(n_2133)
);

XOR2xp5_ASAP7_75t_L g2134 ( 
.A(n_2029),
.B(n_279),
.Y(n_2134)
);

INVx1_ASAP7_75t_L g2135 ( 
.A(n_2062),
.Y(n_2135)
);

AND2x4_ASAP7_75t_L g2136 ( 
.A(n_2002),
.B(n_279),
.Y(n_2136)
);

XNOR2xp5_ASAP7_75t_L g2137 ( 
.A(n_2054),
.B(n_280),
.Y(n_2137)
);

AOI22xp5_ASAP7_75t_L g2138 ( 
.A1(n_2065),
.A2(n_282),
.B1(n_280),
.B2(n_281),
.Y(n_2138)
);

INVx1_ASAP7_75t_SL g2139 ( 
.A(n_2066),
.Y(n_2139)
);

INVx1_ASAP7_75t_SL g2140 ( 
.A(n_2067),
.Y(n_2140)
);

INVxp67_ASAP7_75t_L g2141 ( 
.A(n_2002),
.Y(n_2141)
);

INVx1_ASAP7_75t_L g2142 ( 
.A(n_2069),
.Y(n_2142)
);

XOR2xp5_ASAP7_75t_L g2143 ( 
.A(n_2068),
.B(n_281),
.Y(n_2143)
);

NOR2xp33_ASAP7_75t_L g2144 ( 
.A(n_2014),
.B(n_282),
.Y(n_2144)
);

INVx1_ASAP7_75t_SL g2145 ( 
.A(n_2022),
.Y(n_2145)
);

INVxp67_ASAP7_75t_L g2146 ( 
.A(n_2039),
.Y(n_2146)
);

INVx2_ASAP7_75t_L g2147 ( 
.A(n_2017),
.Y(n_2147)
);

AND2x2_ASAP7_75t_L g2148 ( 
.A(n_1994),
.B(n_283),
.Y(n_2148)
);

XOR2x2_ASAP7_75t_L g2149 ( 
.A(n_1979),
.B(n_283),
.Y(n_2149)
);

INVx2_ASAP7_75t_L g2150 ( 
.A(n_2035),
.Y(n_2150)
);

XNOR2xp5_ASAP7_75t_L g2151 ( 
.A(n_2023),
.B(n_284),
.Y(n_2151)
);

INVx1_ASAP7_75t_SL g2152 ( 
.A(n_2031),
.Y(n_2152)
);

XOR2x2_ASAP7_75t_L g2153 ( 
.A(n_2033),
.B(n_284),
.Y(n_2153)
);

INVx1_ASAP7_75t_SL g2154 ( 
.A(n_2038),
.Y(n_2154)
);

INVxp67_ASAP7_75t_L g2155 ( 
.A(n_2032),
.Y(n_2155)
);

XOR2x2_ASAP7_75t_L g2156 ( 
.A(n_2034),
.B(n_285),
.Y(n_2156)
);

XOR2x2_ASAP7_75t_L g2157 ( 
.A(n_2041),
.B(n_2005),
.Y(n_2157)
);

INVx1_ASAP7_75t_L g2158 ( 
.A(n_2007),
.Y(n_2158)
);

INVx1_ASAP7_75t_SL g2159 ( 
.A(n_1984),
.Y(n_2159)
);

OR2x2_ASAP7_75t_L g2160 ( 
.A(n_1983),
.B(n_285),
.Y(n_2160)
);

AND2x2_ASAP7_75t_L g2161 ( 
.A(n_2059),
.B(n_286),
.Y(n_2161)
);

AND2x2_ASAP7_75t_L g2162 ( 
.A(n_2059),
.B(n_286),
.Y(n_2162)
);

INVx1_ASAP7_75t_L g2163 ( 
.A(n_1985),
.Y(n_2163)
);

INVx1_ASAP7_75t_L g2164 ( 
.A(n_1985),
.Y(n_2164)
);

XOR2x2_ASAP7_75t_L g2165 ( 
.A(n_1976),
.B(n_287),
.Y(n_2165)
);

NOR2xp33_ASAP7_75t_L g2166 ( 
.A(n_1993),
.B(n_287),
.Y(n_2166)
);

INVx1_ASAP7_75t_L g2167 ( 
.A(n_1985),
.Y(n_2167)
);

INVx2_ASAP7_75t_L g2168 ( 
.A(n_2010),
.Y(n_2168)
);

INVxp67_ASAP7_75t_L g2169 ( 
.A(n_2009),
.Y(n_2169)
);

INVx1_ASAP7_75t_L g2170 ( 
.A(n_1985),
.Y(n_2170)
);

INVx2_ASAP7_75t_L g2171 ( 
.A(n_2010),
.Y(n_2171)
);

XNOR2xp5_ASAP7_75t_L g2172 ( 
.A(n_2048),
.B(n_288),
.Y(n_2172)
);

INVx1_ASAP7_75t_L g2173 ( 
.A(n_1985),
.Y(n_2173)
);

INVxp67_ASAP7_75t_L g2174 ( 
.A(n_2009),
.Y(n_2174)
);

AND2x2_ASAP7_75t_L g2175 ( 
.A(n_2059),
.B(n_289),
.Y(n_2175)
);

INVx2_ASAP7_75t_L g2176 ( 
.A(n_2010),
.Y(n_2176)
);

INVx2_ASAP7_75t_SL g2177 ( 
.A(n_2059),
.Y(n_2177)
);

BUFx2_ASAP7_75t_L g2178 ( 
.A(n_2010),
.Y(n_2178)
);

INVx1_ASAP7_75t_L g2179 ( 
.A(n_1985),
.Y(n_2179)
);

INVx1_ASAP7_75t_SL g2180 ( 
.A(n_1984),
.Y(n_2180)
);

XNOR2xp5_ASAP7_75t_L g2181 ( 
.A(n_2048),
.B(n_289),
.Y(n_2181)
);

INVx1_ASAP7_75t_SL g2182 ( 
.A(n_1984),
.Y(n_2182)
);

HB1xp67_ASAP7_75t_L g2183 ( 
.A(n_2083),
.Y(n_2183)
);

INVx2_ASAP7_75t_L g2184 ( 
.A(n_2093),
.Y(n_2184)
);

XOR2x2_ASAP7_75t_L g2185 ( 
.A(n_2094),
.B(n_290),
.Y(n_2185)
);

XOR2x2_ASAP7_75t_L g2186 ( 
.A(n_2088),
.B(n_290),
.Y(n_2186)
);

OA22x2_ASAP7_75t_L g2187 ( 
.A1(n_2152),
.A2(n_295),
.B1(n_292),
.B2(n_293),
.Y(n_2187)
);

INVx2_ASAP7_75t_SL g2188 ( 
.A(n_2113),
.Y(n_2188)
);

OAI22xp5_ASAP7_75t_L g2189 ( 
.A1(n_2095),
.A2(n_295),
.B1(n_292),
.B2(n_293),
.Y(n_2189)
);

OAI22x1_ASAP7_75t_L g2190 ( 
.A1(n_2169),
.A2(n_2174),
.B1(n_2124),
.B2(n_2140),
.Y(n_2190)
);

BUFx3_ASAP7_75t_L g2191 ( 
.A(n_2079),
.Y(n_2191)
);

INVx2_ASAP7_75t_L g2192 ( 
.A(n_2168),
.Y(n_2192)
);

INVx2_ASAP7_75t_SL g2193 ( 
.A(n_2177),
.Y(n_2193)
);

AOI22x1_ASAP7_75t_L g2194 ( 
.A1(n_2134),
.A2(n_298),
.B1(n_296),
.B2(n_297),
.Y(n_2194)
);

INVx1_ASAP7_75t_L g2195 ( 
.A(n_2070),
.Y(n_2195)
);

OA22x2_ASAP7_75t_L g2196 ( 
.A1(n_2155),
.A2(n_298),
.B1(n_296),
.B2(n_297),
.Y(n_2196)
);

OAI22xp5_ASAP7_75t_L g2197 ( 
.A1(n_2146),
.A2(n_301),
.B1(n_299),
.B2(n_300),
.Y(n_2197)
);

OA22x2_ASAP7_75t_L g2198 ( 
.A1(n_2098),
.A2(n_302),
.B1(n_299),
.B2(n_301),
.Y(n_2198)
);

XNOR2x1_ASAP7_75t_L g2199 ( 
.A(n_2165),
.B(n_303),
.Y(n_2199)
);

INVx2_ASAP7_75t_SL g2200 ( 
.A(n_2136),
.Y(n_2200)
);

OA22x2_ASAP7_75t_L g2201 ( 
.A1(n_2139),
.A2(n_305),
.B1(n_303),
.B2(n_304),
.Y(n_2201)
);

INVx2_ASAP7_75t_L g2202 ( 
.A(n_2171),
.Y(n_2202)
);

INVx1_ASAP7_75t_L g2203 ( 
.A(n_2074),
.Y(n_2203)
);

BUFx2_ASAP7_75t_L g2204 ( 
.A(n_2141),
.Y(n_2204)
);

INVx1_ASAP7_75t_L g2205 ( 
.A(n_2076),
.Y(n_2205)
);

INVx2_ASAP7_75t_SL g2206 ( 
.A(n_2085),
.Y(n_2206)
);

AOI22x1_ASAP7_75t_L g2207 ( 
.A1(n_2158),
.A2(n_306),
.B1(n_304),
.B2(n_305),
.Y(n_2207)
);

XOR2x2_ASAP7_75t_L g2208 ( 
.A(n_2090),
.B(n_306),
.Y(n_2208)
);

AOI22x1_ASAP7_75t_L g2209 ( 
.A1(n_2121),
.A2(n_309),
.B1(n_307),
.B2(n_308),
.Y(n_2209)
);

INVx2_ASAP7_75t_L g2210 ( 
.A(n_2176),
.Y(n_2210)
);

AOI22xp5_ASAP7_75t_L g2211 ( 
.A1(n_2157),
.A2(n_2132),
.B1(n_2099),
.B2(n_2108),
.Y(n_2211)
);

INVx2_ASAP7_75t_L g2212 ( 
.A(n_2147),
.Y(n_2212)
);

OR2x2_ASAP7_75t_L g2213 ( 
.A(n_2109),
.B(n_307),
.Y(n_2213)
);

OA22x2_ASAP7_75t_L g2214 ( 
.A1(n_2145),
.A2(n_311),
.B1(n_309),
.B2(n_310),
.Y(n_2214)
);

XOR2x2_ASAP7_75t_L g2215 ( 
.A(n_2072),
.B(n_311),
.Y(n_2215)
);

INVx1_ASAP7_75t_L g2216 ( 
.A(n_2078),
.Y(n_2216)
);

INVx2_ASAP7_75t_L g2217 ( 
.A(n_2178),
.Y(n_2217)
);

INVx2_ASAP7_75t_L g2218 ( 
.A(n_2106),
.Y(n_2218)
);

XNOR2xp5_ASAP7_75t_L g2219 ( 
.A(n_2087),
.B(n_313),
.Y(n_2219)
);

OA22x2_ASAP7_75t_L g2220 ( 
.A1(n_2116),
.A2(n_2137),
.B1(n_2150),
.B2(n_2075),
.Y(n_2220)
);

XOR2xp5_ASAP7_75t_L g2221 ( 
.A(n_2100),
.B(n_313),
.Y(n_2221)
);

INVx1_ASAP7_75t_SL g2222 ( 
.A(n_2111),
.Y(n_2222)
);

INVx3_ASAP7_75t_L g2223 ( 
.A(n_2159),
.Y(n_2223)
);

XNOR2x1_ASAP7_75t_L g2224 ( 
.A(n_2097),
.B(n_314),
.Y(n_2224)
);

BUFx2_ASAP7_75t_L g2225 ( 
.A(n_2092),
.Y(n_2225)
);

INVx2_ASAP7_75t_L g2226 ( 
.A(n_2103),
.Y(n_2226)
);

INVx2_ASAP7_75t_L g2227 ( 
.A(n_2110),
.Y(n_2227)
);

BUFx3_ASAP7_75t_L g2228 ( 
.A(n_2148),
.Y(n_2228)
);

INVx2_ASAP7_75t_L g2229 ( 
.A(n_2118),
.Y(n_2229)
);

OA22x2_ASAP7_75t_L g2230 ( 
.A1(n_2180),
.A2(n_316),
.B1(n_314),
.B2(n_315),
.Y(n_2230)
);

OAI22xp5_ASAP7_75t_SL g2231 ( 
.A1(n_2112),
.A2(n_323),
.B1(n_332),
.B2(n_315),
.Y(n_2231)
);

OA22x2_ASAP7_75t_L g2232 ( 
.A1(n_2182),
.A2(n_318),
.B1(n_316),
.B2(n_317),
.Y(n_2232)
);

INVx2_ASAP7_75t_L g2233 ( 
.A(n_2084),
.Y(n_2233)
);

AOI22x1_ASAP7_75t_L g2234 ( 
.A1(n_2101),
.A2(n_319),
.B1(n_317),
.B2(n_318),
.Y(n_2234)
);

AO22x2_ASAP7_75t_L g2235 ( 
.A1(n_2115),
.A2(n_322),
.B1(n_320),
.B2(n_321),
.Y(n_2235)
);

OA22x2_ASAP7_75t_L g2236 ( 
.A1(n_2154),
.A2(n_325),
.B1(n_320),
.B2(n_323),
.Y(n_2236)
);

AO22x2_ASAP7_75t_L g2237 ( 
.A1(n_2126),
.A2(n_328),
.B1(n_326),
.B2(n_327),
.Y(n_2237)
);

INVx1_ASAP7_75t_L g2238 ( 
.A(n_2163),
.Y(n_2238)
);

OA22x2_ASAP7_75t_L g2239 ( 
.A1(n_2105),
.A2(n_328),
.B1(n_326),
.B2(n_327),
.Y(n_2239)
);

OAI22x1_ASAP7_75t_SL g2240 ( 
.A1(n_2128),
.A2(n_331),
.B1(n_329),
.B2(n_330),
.Y(n_2240)
);

OA22x2_ASAP7_75t_L g2241 ( 
.A1(n_2077),
.A2(n_331),
.B1(n_329),
.B2(n_330),
.Y(n_2241)
);

INVx1_ASAP7_75t_L g2242 ( 
.A(n_2164),
.Y(n_2242)
);

INVx2_ASAP7_75t_SL g2243 ( 
.A(n_2123),
.Y(n_2243)
);

OAI22xp5_ASAP7_75t_L g2244 ( 
.A1(n_2138),
.A2(n_334),
.B1(n_332),
.B2(n_333),
.Y(n_2244)
);

AOI22xp5_ASAP7_75t_L g2245 ( 
.A1(n_2071),
.A2(n_336),
.B1(n_334),
.B2(n_335),
.Y(n_2245)
);

INVx3_ASAP7_75t_SL g2246 ( 
.A(n_2149),
.Y(n_2246)
);

XNOR2x1_ASAP7_75t_L g2247 ( 
.A(n_2172),
.B(n_336),
.Y(n_2247)
);

AO22x2_ASAP7_75t_L g2248 ( 
.A1(n_2119),
.A2(n_339),
.B1(n_337),
.B2(n_338),
.Y(n_2248)
);

AOI22x1_ASAP7_75t_L g2249 ( 
.A1(n_2143),
.A2(n_340),
.B1(n_337),
.B2(n_339),
.Y(n_2249)
);

INVx1_ASAP7_75t_L g2250 ( 
.A(n_2167),
.Y(n_2250)
);

OA22x2_ASAP7_75t_L g2251 ( 
.A1(n_2086),
.A2(n_342),
.B1(n_340),
.B2(n_341),
.Y(n_2251)
);

INVx1_ASAP7_75t_L g2252 ( 
.A(n_2170),
.Y(n_2252)
);

INVx2_ASAP7_75t_L g2253 ( 
.A(n_2173),
.Y(n_2253)
);

AO22x1_ASAP7_75t_L g2254 ( 
.A1(n_2073),
.A2(n_343),
.B1(n_341),
.B2(n_342),
.Y(n_2254)
);

AOI22xp5_ASAP7_75t_L g2255 ( 
.A1(n_2082),
.A2(n_345),
.B1(n_343),
.B2(n_344),
.Y(n_2255)
);

OA22x2_ASAP7_75t_L g2256 ( 
.A1(n_2181),
.A2(n_348),
.B1(n_346),
.B2(n_347),
.Y(n_2256)
);

INVx1_ASAP7_75t_SL g2257 ( 
.A(n_2081),
.Y(n_2257)
);

HB1xp67_ASAP7_75t_L g2258 ( 
.A(n_2089),
.Y(n_2258)
);

INVx1_ASAP7_75t_L g2259 ( 
.A(n_2179),
.Y(n_2259)
);

AND2x4_ASAP7_75t_L g2260 ( 
.A(n_2120),
.B(n_346),
.Y(n_2260)
);

INVx2_ASAP7_75t_L g2261 ( 
.A(n_2091),
.Y(n_2261)
);

XOR2x2_ASAP7_75t_L g2262 ( 
.A(n_2102),
.B(n_347),
.Y(n_2262)
);

INVx2_ASAP7_75t_L g2263 ( 
.A(n_2130),
.Y(n_2263)
);

AOI22x1_ASAP7_75t_L g2264 ( 
.A1(n_2161),
.A2(n_350),
.B1(n_348),
.B2(n_349),
.Y(n_2264)
);

INVx2_ASAP7_75t_L g2265 ( 
.A(n_2131),
.Y(n_2265)
);

XNOR2xp5_ASAP7_75t_L g2266 ( 
.A(n_2151),
.B(n_349),
.Y(n_2266)
);

INVx1_ASAP7_75t_L g2267 ( 
.A(n_2096),
.Y(n_2267)
);

OA22x2_ASAP7_75t_L g2268 ( 
.A1(n_2162),
.A2(n_352),
.B1(n_350),
.B2(n_351),
.Y(n_2268)
);

AOI22x1_ASAP7_75t_L g2269 ( 
.A1(n_2175),
.A2(n_353),
.B1(n_351),
.B2(n_352),
.Y(n_2269)
);

OA22x2_ASAP7_75t_L g2270 ( 
.A1(n_2127),
.A2(n_356),
.B1(n_354),
.B2(n_355),
.Y(n_2270)
);

INVx1_ASAP7_75t_L g2271 ( 
.A(n_2107),
.Y(n_2271)
);

OA22x2_ASAP7_75t_L g2272 ( 
.A1(n_2135),
.A2(n_357),
.B1(n_354),
.B2(n_356),
.Y(n_2272)
);

INVx1_ASAP7_75t_L g2273 ( 
.A(n_2107),
.Y(n_2273)
);

OA22x2_ASAP7_75t_L g2274 ( 
.A1(n_2142),
.A2(n_363),
.B1(n_361),
.B2(n_362),
.Y(n_2274)
);

OAI22xp5_ASAP7_75t_L g2275 ( 
.A1(n_2080),
.A2(n_369),
.B1(n_364),
.B2(n_368),
.Y(n_2275)
);

INVx2_ASAP7_75t_L g2276 ( 
.A(n_2160),
.Y(n_2276)
);

AOI22x1_ASAP7_75t_L g2277 ( 
.A1(n_2114),
.A2(n_372),
.B1(n_370),
.B2(n_371),
.Y(n_2277)
);

INVx2_ASAP7_75t_L g2278 ( 
.A(n_2104),
.Y(n_2278)
);

INVx1_ASAP7_75t_L g2279 ( 
.A(n_2144),
.Y(n_2279)
);

INVx5_ASAP7_75t_L g2280 ( 
.A(n_2153),
.Y(n_2280)
);

INVx2_ASAP7_75t_L g2281 ( 
.A(n_2122),
.Y(n_2281)
);

INVx2_ASAP7_75t_L g2282 ( 
.A(n_2125),
.Y(n_2282)
);

HB1xp67_ASAP7_75t_L g2283 ( 
.A(n_2166),
.Y(n_2283)
);

XNOR2xp5_ASAP7_75t_L g2284 ( 
.A(n_2133),
.B(n_374),
.Y(n_2284)
);

XNOR2x1_ASAP7_75t_L g2285 ( 
.A(n_2156),
.B(n_375),
.Y(n_2285)
);

INVx1_ASAP7_75t_SL g2286 ( 
.A(n_2117),
.Y(n_2286)
);

INVxp67_ASAP7_75t_L g2287 ( 
.A(n_2129),
.Y(n_2287)
);

INVx5_ASAP7_75t_L g2288 ( 
.A(n_2165),
.Y(n_2288)
);

OA22x2_ASAP7_75t_L g2289 ( 
.A1(n_2152),
.A2(n_380),
.B1(n_377),
.B2(n_379),
.Y(n_2289)
);

XNOR2xp5_ASAP7_75t_L g2290 ( 
.A(n_2087),
.B(n_381),
.Y(n_2290)
);

INVx2_ASAP7_75t_SL g2291 ( 
.A(n_2113),
.Y(n_2291)
);

INVx2_ASAP7_75t_L g2292 ( 
.A(n_2093),
.Y(n_2292)
);

OA22x2_ASAP7_75t_L g2293 ( 
.A1(n_2152),
.A2(n_384),
.B1(n_382),
.B2(n_383),
.Y(n_2293)
);

OA22x2_ASAP7_75t_L g2294 ( 
.A1(n_2152),
.A2(n_388),
.B1(n_385),
.B2(n_387),
.Y(n_2294)
);

INVx2_ASAP7_75t_L g2295 ( 
.A(n_2093),
.Y(n_2295)
);

CKINVDCx20_ASAP7_75t_R g2296 ( 
.A(n_2113),
.Y(n_2296)
);

INVx1_ASAP7_75t_L g2297 ( 
.A(n_2070),
.Y(n_2297)
);

AOI22xp5_ASAP7_75t_L g2298 ( 
.A1(n_2157),
.A2(n_394),
.B1(n_390),
.B2(n_393),
.Y(n_2298)
);

INVx1_ASAP7_75t_L g2299 ( 
.A(n_2070),
.Y(n_2299)
);

NAND2xp5_ASAP7_75t_L g2300 ( 
.A(n_2169),
.B(n_395),
.Y(n_2300)
);

INVx3_ASAP7_75t_L g2301 ( 
.A(n_2079),
.Y(n_2301)
);

AOI22xp5_ASAP7_75t_L g2302 ( 
.A1(n_2157),
.A2(n_399),
.B1(n_396),
.B2(n_397),
.Y(n_2302)
);

OAI22xp5_ASAP7_75t_L g2303 ( 
.A1(n_2095),
.A2(n_403),
.B1(n_400),
.B2(n_402),
.Y(n_2303)
);

INVx2_ASAP7_75t_SL g2304 ( 
.A(n_2113),
.Y(n_2304)
);

INVx2_ASAP7_75t_SL g2305 ( 
.A(n_2113),
.Y(n_2305)
);

INVx3_ASAP7_75t_SL g2306 ( 
.A(n_2165),
.Y(n_2306)
);

XOR2x2_ASAP7_75t_L g2307 ( 
.A(n_2094),
.B(n_404),
.Y(n_2307)
);

INVx1_ASAP7_75t_L g2308 ( 
.A(n_2070),
.Y(n_2308)
);

AOI22x1_ASAP7_75t_L g2309 ( 
.A1(n_2152),
.A2(n_407),
.B1(n_405),
.B2(n_406),
.Y(n_2309)
);

XNOR2x1_ASAP7_75t_L g2310 ( 
.A(n_2094),
.B(n_408),
.Y(n_2310)
);

BUFx3_ASAP7_75t_L g2311 ( 
.A(n_2079),
.Y(n_2311)
);

OA22x2_ASAP7_75t_L g2312 ( 
.A1(n_2152),
.A2(n_412),
.B1(n_409),
.B2(n_411),
.Y(n_2312)
);

INVx2_ASAP7_75t_L g2313 ( 
.A(n_2093),
.Y(n_2313)
);

INVxp67_ASAP7_75t_SL g2314 ( 
.A(n_2102),
.Y(n_2314)
);

HB1xp67_ASAP7_75t_L g2315 ( 
.A(n_2083),
.Y(n_2315)
);

INVx2_ASAP7_75t_L g2316 ( 
.A(n_2093),
.Y(n_2316)
);

INVx1_ASAP7_75t_L g2317 ( 
.A(n_2070),
.Y(n_2317)
);

INVx1_ASAP7_75t_L g2318 ( 
.A(n_2070),
.Y(n_2318)
);

INVx1_ASAP7_75t_SL g2319 ( 
.A(n_2111),
.Y(n_2319)
);

INVx2_ASAP7_75t_L g2320 ( 
.A(n_2093),
.Y(n_2320)
);

INVx2_ASAP7_75t_L g2321 ( 
.A(n_2093),
.Y(n_2321)
);

AND2x4_ASAP7_75t_L g2322 ( 
.A(n_2141),
.B(n_413),
.Y(n_2322)
);

INVx1_ASAP7_75t_L g2323 ( 
.A(n_2070),
.Y(n_2323)
);

AOI22x1_ASAP7_75t_L g2324 ( 
.A1(n_2152),
.A2(n_416),
.B1(n_414),
.B2(n_415),
.Y(n_2324)
);

INVx1_ASAP7_75t_L g2325 ( 
.A(n_2070),
.Y(n_2325)
);

INVx1_ASAP7_75t_L g2326 ( 
.A(n_2070),
.Y(n_2326)
);

INVx1_ASAP7_75t_L g2327 ( 
.A(n_2070),
.Y(n_2327)
);

XNOR2xp5_ASAP7_75t_L g2328 ( 
.A(n_2087),
.B(n_417),
.Y(n_2328)
);

XNOR2xp5_ASAP7_75t_L g2329 ( 
.A(n_2087),
.B(n_418),
.Y(n_2329)
);

XOR2x2_ASAP7_75t_L g2330 ( 
.A(n_2094),
.B(n_419),
.Y(n_2330)
);

INVx1_ASAP7_75t_L g2331 ( 
.A(n_2070),
.Y(n_2331)
);

OA22x2_ASAP7_75t_L g2332 ( 
.A1(n_2152),
.A2(n_422),
.B1(n_420),
.B2(n_421),
.Y(n_2332)
);

OA22x2_ASAP7_75t_L g2333 ( 
.A1(n_2152),
.A2(n_428),
.B1(n_423),
.B2(n_424),
.Y(n_2333)
);

AOI22x1_ASAP7_75t_L g2334 ( 
.A1(n_2152),
.A2(n_434),
.B1(n_431),
.B2(n_433),
.Y(n_2334)
);

AOI22x1_ASAP7_75t_L g2335 ( 
.A1(n_2152),
.A2(n_437),
.B1(n_435),
.B2(n_436),
.Y(n_2335)
);

OA22x2_ASAP7_75t_L g2336 ( 
.A1(n_2152),
.A2(n_441),
.B1(n_438),
.B2(n_439),
.Y(n_2336)
);

XOR2x2_ASAP7_75t_L g2337 ( 
.A(n_2094),
.B(n_442),
.Y(n_2337)
);

OA22x2_ASAP7_75t_L g2338 ( 
.A1(n_2152),
.A2(n_447),
.B1(n_444),
.B2(n_445),
.Y(n_2338)
);

OAI22xp5_ASAP7_75t_L g2339 ( 
.A1(n_2095),
.A2(n_451),
.B1(n_449),
.B2(n_450),
.Y(n_2339)
);

AND2x4_ASAP7_75t_L g2340 ( 
.A(n_2141),
.B(n_452),
.Y(n_2340)
);

XNOR2xp5_ASAP7_75t_L g2341 ( 
.A(n_2087),
.B(n_454),
.Y(n_2341)
);

OA22x2_ASAP7_75t_L g2342 ( 
.A1(n_2152),
.A2(n_457),
.B1(n_455),
.B2(n_456),
.Y(n_2342)
);

INVx1_ASAP7_75t_L g2343 ( 
.A(n_2070),
.Y(n_2343)
);

BUFx3_ASAP7_75t_L g2344 ( 
.A(n_2079),
.Y(n_2344)
);

XOR2x2_ASAP7_75t_L g2345 ( 
.A(n_2094),
.B(n_458),
.Y(n_2345)
);

INVx1_ASAP7_75t_L g2346 ( 
.A(n_2070),
.Y(n_2346)
);

INVx1_ASAP7_75t_L g2347 ( 
.A(n_2070),
.Y(n_2347)
);

INVx1_ASAP7_75t_L g2348 ( 
.A(n_2070),
.Y(n_2348)
);

INVxp67_ASAP7_75t_L g2349 ( 
.A(n_2191),
.Y(n_2349)
);

INVx1_ASAP7_75t_L g2350 ( 
.A(n_2258),
.Y(n_2350)
);

INVx1_ASAP7_75t_L g2351 ( 
.A(n_2195),
.Y(n_2351)
);

INVx2_ASAP7_75t_L g2352 ( 
.A(n_2296),
.Y(n_2352)
);

INVx2_ASAP7_75t_L g2353 ( 
.A(n_2188),
.Y(n_2353)
);

INVx1_ASAP7_75t_L g2354 ( 
.A(n_2203),
.Y(n_2354)
);

OAI322xp33_ASAP7_75t_L g2355 ( 
.A1(n_2314),
.A2(n_467),
.A3(n_466),
.B1(n_461),
.B2(n_459),
.C1(n_460),
.C2(n_464),
.Y(n_2355)
);

BUFx2_ASAP7_75t_L g2356 ( 
.A(n_2311),
.Y(n_2356)
);

INVx1_ASAP7_75t_L g2357 ( 
.A(n_2205),
.Y(n_2357)
);

INVx1_ASAP7_75t_L g2358 ( 
.A(n_2216),
.Y(n_2358)
);

INVxp67_ASAP7_75t_L g2359 ( 
.A(n_2344),
.Y(n_2359)
);

INVx1_ASAP7_75t_L g2360 ( 
.A(n_2238),
.Y(n_2360)
);

INVx1_ASAP7_75t_L g2361 ( 
.A(n_2242),
.Y(n_2361)
);

INVx1_ASAP7_75t_L g2362 ( 
.A(n_2250),
.Y(n_2362)
);

INVx1_ASAP7_75t_L g2363 ( 
.A(n_2252),
.Y(n_2363)
);

NAND2xp5_ASAP7_75t_SL g2364 ( 
.A(n_2303),
.B(n_468),
.Y(n_2364)
);

INVx2_ASAP7_75t_L g2365 ( 
.A(n_2291),
.Y(n_2365)
);

INVx1_ASAP7_75t_SL g2366 ( 
.A(n_2222),
.Y(n_2366)
);

OA22x2_ASAP7_75t_L g2367 ( 
.A1(n_2211),
.A2(n_473),
.B1(n_470),
.B2(n_472),
.Y(n_2367)
);

INVx1_ASAP7_75t_L g2368 ( 
.A(n_2259),
.Y(n_2368)
);

INVx1_ASAP7_75t_L g2369 ( 
.A(n_2297),
.Y(n_2369)
);

CKINVDCx5p33_ASAP7_75t_R g2370 ( 
.A(n_2306),
.Y(n_2370)
);

INVxp67_ASAP7_75t_L g2371 ( 
.A(n_2301),
.Y(n_2371)
);

INVx1_ASAP7_75t_L g2372 ( 
.A(n_2299),
.Y(n_2372)
);

XNOR2x2_ASAP7_75t_L g2373 ( 
.A(n_2220),
.B(n_748),
.Y(n_2373)
);

INVx2_ASAP7_75t_L g2374 ( 
.A(n_2304),
.Y(n_2374)
);

AO22x2_ASAP7_75t_L g2375 ( 
.A1(n_2189),
.A2(n_479),
.B1(n_475),
.B2(n_477),
.Y(n_2375)
);

INVx1_ASAP7_75t_L g2376 ( 
.A(n_2308),
.Y(n_2376)
);

INVxp33_ASAP7_75t_L g2377 ( 
.A(n_2283),
.Y(n_2377)
);

INVx1_ASAP7_75t_L g2378 ( 
.A(n_2317),
.Y(n_2378)
);

INVx1_ASAP7_75t_L g2379 ( 
.A(n_2318),
.Y(n_2379)
);

BUFx2_ASAP7_75t_L g2380 ( 
.A(n_2305),
.Y(n_2380)
);

INVx1_ASAP7_75t_L g2381 ( 
.A(n_2323),
.Y(n_2381)
);

AOI22xp5_ASAP7_75t_SL g2382 ( 
.A1(n_2187),
.A2(n_484),
.B1(n_480),
.B2(n_482),
.Y(n_2382)
);

INVx2_ASAP7_75t_L g2383 ( 
.A(n_2228),
.Y(n_2383)
);

HB1xp67_ASAP7_75t_L g2384 ( 
.A(n_2183),
.Y(n_2384)
);

INVx2_ASAP7_75t_L g2385 ( 
.A(n_2223),
.Y(n_2385)
);

INVx1_ASAP7_75t_L g2386 ( 
.A(n_2325),
.Y(n_2386)
);

INVx1_ASAP7_75t_L g2387 ( 
.A(n_2326),
.Y(n_2387)
);

INVx1_ASAP7_75t_L g2388 ( 
.A(n_2327),
.Y(n_2388)
);

INVx2_ASAP7_75t_L g2389 ( 
.A(n_2204),
.Y(n_2389)
);

INVxp67_ASAP7_75t_L g2390 ( 
.A(n_2278),
.Y(n_2390)
);

INVx1_ASAP7_75t_L g2391 ( 
.A(n_2331),
.Y(n_2391)
);

BUFx2_ASAP7_75t_L g2392 ( 
.A(n_2225),
.Y(n_2392)
);

INVxp67_ASAP7_75t_L g2393 ( 
.A(n_2281),
.Y(n_2393)
);

INVx1_ASAP7_75t_L g2394 ( 
.A(n_2343),
.Y(n_2394)
);

INVx2_ASAP7_75t_L g2395 ( 
.A(n_2206),
.Y(n_2395)
);

AOI22xp5_ASAP7_75t_L g2396 ( 
.A1(n_2339),
.A2(n_2185),
.B1(n_2245),
.B2(n_2255),
.Y(n_2396)
);

INVx1_ASAP7_75t_L g2397 ( 
.A(n_2346),
.Y(n_2397)
);

INVx1_ASAP7_75t_L g2398 ( 
.A(n_2347),
.Y(n_2398)
);

INVx1_ASAP7_75t_L g2399 ( 
.A(n_2348),
.Y(n_2399)
);

INVx1_ASAP7_75t_L g2400 ( 
.A(n_2267),
.Y(n_2400)
);

INVx1_ASAP7_75t_L g2401 ( 
.A(n_2233),
.Y(n_2401)
);

INVx1_ASAP7_75t_SL g2402 ( 
.A(n_2319),
.Y(n_2402)
);

INVx1_ASAP7_75t_L g2403 ( 
.A(n_2253),
.Y(n_2403)
);

INVx2_ASAP7_75t_L g2404 ( 
.A(n_2257),
.Y(n_2404)
);

INVx1_ASAP7_75t_L g2405 ( 
.A(n_2315),
.Y(n_2405)
);

AOI322xp5_ASAP7_75t_L g2406 ( 
.A1(n_2288),
.A2(n_493),
.A3(n_492),
.B1(n_487),
.B2(n_485),
.C1(n_486),
.C2(n_488),
.Y(n_2406)
);

NOR2xp33_ASAP7_75t_L g2407 ( 
.A(n_2288),
.B(n_494),
.Y(n_2407)
);

INVx1_ASAP7_75t_L g2408 ( 
.A(n_2227),
.Y(n_2408)
);

INVx1_ASAP7_75t_L g2409 ( 
.A(n_2229),
.Y(n_2409)
);

INVx1_ASAP7_75t_L g2410 ( 
.A(n_2261),
.Y(n_2410)
);

INVx1_ASAP7_75t_L g2411 ( 
.A(n_2276),
.Y(n_2411)
);

OAI322xp33_ASAP7_75t_L g2412 ( 
.A1(n_2287),
.A2(n_2199),
.A3(n_2246),
.B1(n_2230),
.B2(n_2232),
.C1(n_2214),
.C2(n_2231),
.Y(n_2412)
);

INVx1_ASAP7_75t_L g2413 ( 
.A(n_2271),
.Y(n_2413)
);

INVx1_ASAP7_75t_L g2414 ( 
.A(n_2273),
.Y(n_2414)
);

INVx2_ASAP7_75t_L g2415 ( 
.A(n_2243),
.Y(n_2415)
);

INVx1_ASAP7_75t_L g2416 ( 
.A(n_2213),
.Y(n_2416)
);

INVx1_ASAP7_75t_L g2417 ( 
.A(n_2226),
.Y(n_2417)
);

INVx1_ASAP7_75t_L g2418 ( 
.A(n_2263),
.Y(n_2418)
);

INVx1_ASAP7_75t_L g2419 ( 
.A(n_2265),
.Y(n_2419)
);

OAI322xp33_ASAP7_75t_L g2420 ( 
.A1(n_2201),
.A2(n_505),
.A3(n_501),
.B1(n_499),
.B2(n_497),
.C1(n_498),
.C2(n_500),
.Y(n_2420)
);

INVx1_ASAP7_75t_L g2421 ( 
.A(n_2248),
.Y(n_2421)
);

OA22x2_ASAP7_75t_L g2422 ( 
.A1(n_2190),
.A2(n_509),
.B1(n_506),
.B2(n_507),
.Y(n_2422)
);

OAI22xp5_ASAP7_75t_L g2423 ( 
.A1(n_2286),
.A2(n_512),
.B1(n_510),
.B2(n_511),
.Y(n_2423)
);

HB1xp67_ASAP7_75t_L g2424 ( 
.A(n_2217),
.Y(n_2424)
);

BUFx2_ASAP7_75t_L g2425 ( 
.A(n_2193),
.Y(n_2425)
);

INVx1_ASAP7_75t_L g2426 ( 
.A(n_2212),
.Y(n_2426)
);

INVx1_ASAP7_75t_L g2427 ( 
.A(n_2236),
.Y(n_2427)
);

BUFx2_ASAP7_75t_L g2428 ( 
.A(n_2279),
.Y(n_2428)
);

INVx1_ASAP7_75t_L g2429 ( 
.A(n_2235),
.Y(n_2429)
);

INVx1_ASAP7_75t_L g2430 ( 
.A(n_2237),
.Y(n_2430)
);

INVx1_ASAP7_75t_L g2431 ( 
.A(n_2300),
.Y(n_2431)
);

INVx2_ASAP7_75t_L g2432 ( 
.A(n_2184),
.Y(n_2432)
);

INVx1_ASAP7_75t_L g2433 ( 
.A(n_2272),
.Y(n_2433)
);

INVxp67_ASAP7_75t_L g2434 ( 
.A(n_2282),
.Y(n_2434)
);

INVx1_ASAP7_75t_L g2435 ( 
.A(n_2192),
.Y(n_2435)
);

INVx1_ASAP7_75t_L g2436 ( 
.A(n_2202),
.Y(n_2436)
);

INVx1_ASAP7_75t_L g2437 ( 
.A(n_2210),
.Y(n_2437)
);

INVx2_ASAP7_75t_SL g2438 ( 
.A(n_2260),
.Y(n_2438)
);

INVx1_ASAP7_75t_L g2439 ( 
.A(n_2292),
.Y(n_2439)
);

INVx2_ASAP7_75t_SL g2440 ( 
.A(n_2200),
.Y(n_2440)
);

INVx1_ASAP7_75t_L g2441 ( 
.A(n_2295),
.Y(n_2441)
);

INVx2_ASAP7_75t_L g2442 ( 
.A(n_2313),
.Y(n_2442)
);

INVx2_ASAP7_75t_L g2443 ( 
.A(n_2316),
.Y(n_2443)
);

INVxp67_ASAP7_75t_SL g2444 ( 
.A(n_2240),
.Y(n_2444)
);

INVx1_ASAP7_75t_L g2445 ( 
.A(n_2320),
.Y(n_2445)
);

INVx1_ASAP7_75t_SL g2446 ( 
.A(n_2221),
.Y(n_2446)
);

INVx1_ASAP7_75t_L g2447 ( 
.A(n_2321),
.Y(n_2447)
);

INVx1_ASAP7_75t_L g2448 ( 
.A(n_2218),
.Y(n_2448)
);

INVx1_ASAP7_75t_L g2449 ( 
.A(n_2270),
.Y(n_2449)
);

INVx1_ASAP7_75t_L g2450 ( 
.A(n_2268),
.Y(n_2450)
);

INVx1_ASAP7_75t_L g2451 ( 
.A(n_2196),
.Y(n_2451)
);

INVx1_ASAP7_75t_L g2452 ( 
.A(n_2197),
.Y(n_2452)
);

INVx1_ASAP7_75t_L g2453 ( 
.A(n_2254),
.Y(n_2453)
);

INVx1_ASAP7_75t_L g2454 ( 
.A(n_2251),
.Y(n_2454)
);

INVx1_ASAP7_75t_L g2455 ( 
.A(n_2198),
.Y(n_2455)
);

OA22x2_ASAP7_75t_L g2456 ( 
.A1(n_2298),
.A2(n_516),
.B1(n_513),
.B2(n_515),
.Y(n_2456)
);

INVx1_ASAP7_75t_L g2457 ( 
.A(n_2241),
.Y(n_2457)
);

INVx1_ASAP7_75t_L g2458 ( 
.A(n_2234),
.Y(n_2458)
);

XNOR2xp5_ASAP7_75t_L g2459 ( 
.A(n_2186),
.B(n_517),
.Y(n_2459)
);

NAND2xp33_ASAP7_75t_SL g2460 ( 
.A(n_2310),
.B(n_519),
.Y(n_2460)
);

INVx2_ASAP7_75t_SL g2461 ( 
.A(n_2262),
.Y(n_2461)
);

INVx1_ASAP7_75t_L g2462 ( 
.A(n_2264),
.Y(n_2462)
);

INVx2_ASAP7_75t_L g2463 ( 
.A(n_2289),
.Y(n_2463)
);

INVx3_ASAP7_75t_L g2464 ( 
.A(n_2215),
.Y(n_2464)
);

INVx1_ASAP7_75t_SL g2465 ( 
.A(n_2208),
.Y(n_2465)
);

INVx1_ASAP7_75t_L g2466 ( 
.A(n_2269),
.Y(n_2466)
);

INVx1_ASAP7_75t_L g2467 ( 
.A(n_2293),
.Y(n_2467)
);

INVx1_ASAP7_75t_L g2468 ( 
.A(n_2294),
.Y(n_2468)
);

XNOR2xp5_ASAP7_75t_L g2469 ( 
.A(n_2307),
.B(n_521),
.Y(n_2469)
);

INVx2_ASAP7_75t_L g2470 ( 
.A(n_2312),
.Y(n_2470)
);

NOR2xp33_ASAP7_75t_L g2471 ( 
.A(n_2280),
.B(n_523),
.Y(n_2471)
);

INVx1_ASAP7_75t_L g2472 ( 
.A(n_2384),
.Y(n_2472)
);

INVx1_ASAP7_75t_L g2473 ( 
.A(n_2413),
.Y(n_2473)
);

INVx1_ASAP7_75t_L g2474 ( 
.A(n_2414),
.Y(n_2474)
);

AOI22xp5_ASAP7_75t_L g2475 ( 
.A1(n_2444),
.A2(n_2239),
.B1(n_2256),
.B2(n_2280),
.Y(n_2475)
);

OAI22xp33_ASAP7_75t_L g2476 ( 
.A1(n_2422),
.A2(n_2302),
.B1(n_2333),
.B2(n_2332),
.Y(n_2476)
);

AO22x2_ASAP7_75t_L g2477 ( 
.A1(n_2429),
.A2(n_2224),
.B1(n_2285),
.B2(n_2247),
.Y(n_2477)
);

INVxp67_ASAP7_75t_L g2478 ( 
.A(n_2356),
.Y(n_2478)
);

AOI221xp5_ASAP7_75t_L g2479 ( 
.A1(n_2412),
.A2(n_2244),
.B1(n_2275),
.B2(n_2219),
.C(n_2266),
.Y(n_2479)
);

HB1xp67_ASAP7_75t_L g2480 ( 
.A(n_2349),
.Y(n_2480)
);

INVx1_ASAP7_75t_L g2481 ( 
.A(n_2411),
.Y(n_2481)
);

AND4x1_ASAP7_75t_L g2482 ( 
.A(n_2453),
.B(n_2209),
.C(n_2194),
.D(n_2249),
.Y(n_2482)
);

INVxp67_ASAP7_75t_SL g2483 ( 
.A(n_2464),
.Y(n_2483)
);

OAI22xp5_ASAP7_75t_SL g2484 ( 
.A1(n_2370),
.A2(n_2284),
.B1(n_2328),
.B2(n_2290),
.Y(n_2484)
);

INVxp67_ASAP7_75t_L g2485 ( 
.A(n_2352),
.Y(n_2485)
);

INVx1_ASAP7_75t_L g2486 ( 
.A(n_2351),
.Y(n_2486)
);

A2O1A1Ixp33_ASAP7_75t_L g2487 ( 
.A1(n_2396),
.A2(n_2337),
.B(n_2345),
.C(n_2330),
.Y(n_2487)
);

INVx1_ASAP7_75t_L g2488 ( 
.A(n_2354),
.Y(n_2488)
);

AOI22xp5_ASAP7_75t_L g2489 ( 
.A1(n_2367),
.A2(n_2433),
.B1(n_2451),
.B2(n_2457),
.Y(n_2489)
);

AOI22xp5_ASAP7_75t_L g2490 ( 
.A1(n_2455),
.A2(n_2338),
.B1(n_2342),
.B2(n_2336),
.Y(n_2490)
);

INVx2_ASAP7_75t_L g2491 ( 
.A(n_2380),
.Y(n_2491)
);

INVx2_ASAP7_75t_L g2492 ( 
.A(n_2353),
.Y(n_2492)
);

INVx2_ASAP7_75t_L g2493 ( 
.A(n_2365),
.Y(n_2493)
);

INVx1_ASAP7_75t_L g2494 ( 
.A(n_2357),
.Y(n_2494)
);

INVx1_ASAP7_75t_L g2495 ( 
.A(n_2358),
.Y(n_2495)
);

AOI22x1_ASAP7_75t_L g2496 ( 
.A1(n_2392),
.A2(n_2341),
.B1(n_2329),
.B2(n_2340),
.Y(n_2496)
);

AOI221xp5_ASAP7_75t_L g2497 ( 
.A1(n_2377),
.A2(n_2207),
.B1(n_2322),
.B2(n_2274),
.C(n_2277),
.Y(n_2497)
);

AOI22xp5_ASAP7_75t_L g2498 ( 
.A1(n_2454),
.A2(n_2324),
.B1(n_2334),
.B2(n_2309),
.Y(n_2498)
);

INVx1_ASAP7_75t_L g2499 ( 
.A(n_2360),
.Y(n_2499)
);

AOI22xp5_ASAP7_75t_L g2500 ( 
.A1(n_2449),
.A2(n_2450),
.B1(n_2427),
.B2(n_2467),
.Y(n_2500)
);

OA22x2_ASAP7_75t_L g2501 ( 
.A1(n_2390),
.A2(n_2335),
.B1(n_527),
.B2(n_524),
.Y(n_2501)
);

INVx1_ASAP7_75t_L g2502 ( 
.A(n_2361),
.Y(n_2502)
);

AOI22xp5_ASAP7_75t_L g2503 ( 
.A1(n_2468),
.A2(n_530),
.B1(n_525),
.B2(n_528),
.Y(n_2503)
);

AOI221xp5_ASAP7_75t_L g2504 ( 
.A1(n_2393),
.A2(n_746),
.B1(n_534),
.B2(n_531),
.C(n_532),
.Y(n_2504)
);

AOI22x1_ASAP7_75t_L g2505 ( 
.A1(n_2425),
.A2(n_539),
.B1(n_535),
.B2(n_537),
.Y(n_2505)
);

AOI22x1_ASAP7_75t_L g2506 ( 
.A1(n_2389),
.A2(n_543),
.B1(n_541),
.B2(n_542),
.Y(n_2506)
);

INVx1_ASAP7_75t_SL g2507 ( 
.A(n_2446),
.Y(n_2507)
);

AOI22xp5_ASAP7_75t_L g2508 ( 
.A1(n_2463),
.A2(n_548),
.B1(n_545),
.B2(n_546),
.Y(n_2508)
);

AOI22xp5_ASAP7_75t_L g2509 ( 
.A1(n_2470),
.A2(n_551),
.B1(n_549),
.B2(n_550),
.Y(n_2509)
);

OAI22xp5_ASAP7_75t_L g2510 ( 
.A1(n_2452),
.A2(n_554),
.B1(n_552),
.B2(n_553),
.Y(n_2510)
);

OAI222xp33_ASAP7_75t_L g2511 ( 
.A1(n_2421),
.A2(n_557),
.B1(n_559),
.B2(n_555),
.C1(n_556),
.C2(n_558),
.Y(n_2511)
);

OAI322xp33_ASAP7_75t_L g2512 ( 
.A1(n_2405),
.A2(n_560),
.A3(n_561),
.B1(n_562),
.B2(n_563),
.C1(n_564),
.C2(n_568),
.Y(n_2512)
);

AOI31xp33_ASAP7_75t_L g2513 ( 
.A1(n_2371),
.A2(n_573),
.A3(n_570),
.B(n_572),
.Y(n_2513)
);

INVx1_ASAP7_75t_L g2514 ( 
.A(n_2362),
.Y(n_2514)
);

AOI22xp5_ASAP7_75t_L g2515 ( 
.A1(n_2375),
.A2(n_576),
.B1(n_574),
.B2(n_575),
.Y(n_2515)
);

CKINVDCx20_ASAP7_75t_R g2516 ( 
.A(n_2459),
.Y(n_2516)
);

NAND4xp25_ASAP7_75t_SL g2517 ( 
.A(n_2458),
.B(n_579),
.C(n_577),
.D(n_578),
.Y(n_2517)
);

INVx1_ASAP7_75t_SL g2518 ( 
.A(n_2366),
.Y(n_2518)
);

CKINVDCx20_ASAP7_75t_R g2519 ( 
.A(n_2469),
.Y(n_2519)
);

AOI221xp5_ASAP7_75t_L g2520 ( 
.A1(n_2434),
.A2(n_583),
.B1(n_580),
.B2(n_582),
.C(n_584),
.Y(n_2520)
);

OAI22x1_ASAP7_75t_L g2521 ( 
.A1(n_2385),
.A2(n_588),
.B1(n_585),
.B2(n_587),
.Y(n_2521)
);

OAI322xp33_ASAP7_75t_L g2522 ( 
.A1(n_2461),
.A2(n_589),
.A3(n_590),
.B1(n_592),
.B2(n_595),
.C1(n_596),
.C2(n_597),
.Y(n_2522)
);

AOI22xp5_ASAP7_75t_L g2523 ( 
.A1(n_2375),
.A2(n_600),
.B1(n_598),
.B2(n_599),
.Y(n_2523)
);

INVx3_ASAP7_75t_L g2524 ( 
.A(n_2374),
.Y(n_2524)
);

AOI22xp5_ASAP7_75t_L g2525 ( 
.A1(n_2430),
.A2(n_604),
.B1(n_602),
.B2(n_603),
.Y(n_2525)
);

INVx1_ASAP7_75t_L g2526 ( 
.A(n_2363),
.Y(n_2526)
);

INVx1_ASAP7_75t_L g2527 ( 
.A(n_2368),
.Y(n_2527)
);

INVx1_ASAP7_75t_L g2528 ( 
.A(n_2369),
.Y(n_2528)
);

OAI322xp33_ASAP7_75t_L g2529 ( 
.A1(n_2350),
.A2(n_606),
.A3(n_607),
.B1(n_610),
.B2(n_611),
.C1(n_612),
.C2(n_613),
.Y(n_2529)
);

INVx1_ASAP7_75t_L g2530 ( 
.A(n_2372),
.Y(n_2530)
);

NOR2xp33_ASAP7_75t_L g2531 ( 
.A(n_2359),
.B(n_614),
.Y(n_2531)
);

INVx1_ASAP7_75t_L g2532 ( 
.A(n_2480),
.Y(n_2532)
);

OAI22xp5_ASAP7_75t_L g2533 ( 
.A1(n_2518),
.A2(n_2466),
.B1(n_2462),
.B2(n_2428),
.Y(n_2533)
);

AOI22xp5_ASAP7_75t_L g2534 ( 
.A1(n_2477),
.A2(n_2460),
.B1(n_2364),
.B2(n_2416),
.Y(n_2534)
);

AOI221xp5_ASAP7_75t_SL g2535 ( 
.A1(n_2483),
.A2(n_2402),
.B1(n_2417),
.B2(n_2404),
.C(n_2395),
.Y(n_2535)
);

OAI211xp5_ASAP7_75t_L g2536 ( 
.A1(n_2478),
.A2(n_2424),
.B(n_2383),
.C(n_2440),
.Y(n_2536)
);

INVx1_ASAP7_75t_L g2537 ( 
.A(n_2472),
.Y(n_2537)
);

INVx1_ASAP7_75t_L g2538 ( 
.A(n_2473),
.Y(n_2538)
);

BUFx2_ASAP7_75t_L g2539 ( 
.A(n_2485),
.Y(n_2539)
);

A2O1A1Ixp33_ASAP7_75t_L g2540 ( 
.A1(n_2475),
.A2(n_2407),
.B(n_2382),
.C(n_2471),
.Y(n_2540)
);

INVx2_ASAP7_75t_L g2541 ( 
.A(n_2524),
.Y(n_2541)
);

AOI221xp5_ASAP7_75t_L g2542 ( 
.A1(n_2477),
.A2(n_2465),
.B1(n_2431),
.B2(n_2408),
.C(n_2409),
.Y(n_2542)
);

AOI221xp5_ASAP7_75t_L g2543 ( 
.A1(n_2500),
.A2(n_2410),
.B1(n_2403),
.B2(n_2401),
.C(n_2418),
.Y(n_2543)
);

O2A1O1Ixp33_ASAP7_75t_L g2544 ( 
.A1(n_2479),
.A2(n_2415),
.B(n_2378),
.C(n_2379),
.Y(n_2544)
);

OAI22xp5_ASAP7_75t_L g2545 ( 
.A1(n_2490),
.A2(n_2438),
.B1(n_2381),
.B2(n_2386),
.Y(n_2545)
);

INVx1_ASAP7_75t_L g2546 ( 
.A(n_2474),
.Y(n_2546)
);

AOI22xp5_ASAP7_75t_L g2547 ( 
.A1(n_2476),
.A2(n_2456),
.B1(n_2426),
.B2(n_2436),
.Y(n_2547)
);

INVx1_ASAP7_75t_L g2548 ( 
.A(n_2507),
.Y(n_2548)
);

INVx2_ASAP7_75t_L g2549 ( 
.A(n_2524),
.Y(n_2549)
);

OAI221xp5_ASAP7_75t_L g2550 ( 
.A1(n_2489),
.A2(n_2373),
.B1(n_2419),
.B2(n_2437),
.C(n_2435),
.Y(n_2550)
);

INVx1_ASAP7_75t_L g2551 ( 
.A(n_2486),
.Y(n_2551)
);

INVx1_ASAP7_75t_L g2552 ( 
.A(n_2488),
.Y(n_2552)
);

HB1xp67_ASAP7_75t_L g2553 ( 
.A(n_2491),
.Y(n_2553)
);

HB1xp67_ASAP7_75t_L g2554 ( 
.A(n_2492),
.Y(n_2554)
);

INVx2_ASAP7_75t_L g2555 ( 
.A(n_2493),
.Y(n_2555)
);

AOI22xp5_ASAP7_75t_L g2556 ( 
.A1(n_2501),
.A2(n_2448),
.B1(n_2441),
.B2(n_2445),
.Y(n_2556)
);

AOI22xp33_ASAP7_75t_SL g2557 ( 
.A1(n_2496),
.A2(n_2423),
.B1(n_2447),
.B2(n_2439),
.Y(n_2557)
);

INVx1_ASAP7_75t_L g2558 ( 
.A(n_2494),
.Y(n_2558)
);

INVx1_ASAP7_75t_L g2559 ( 
.A(n_2495),
.Y(n_2559)
);

OAI22xp5_ASAP7_75t_L g2560 ( 
.A1(n_2497),
.A2(n_2376),
.B1(n_2388),
.B2(n_2387),
.Y(n_2560)
);

HB1xp67_ASAP7_75t_L g2561 ( 
.A(n_2482),
.Y(n_2561)
);

AOI22xp5_ASAP7_75t_L g2562 ( 
.A1(n_2498),
.A2(n_2442),
.B1(n_2443),
.B2(n_2432),
.Y(n_2562)
);

AOI22xp33_ASAP7_75t_L g2563 ( 
.A1(n_2515),
.A2(n_2420),
.B1(n_2355),
.B2(n_2394),
.Y(n_2563)
);

INVx1_ASAP7_75t_L g2564 ( 
.A(n_2539),
.Y(n_2564)
);

AOI31xp33_ASAP7_75t_L g2565 ( 
.A1(n_2561),
.A2(n_2499),
.A3(n_2514),
.B(n_2502),
.Y(n_2565)
);

INVx1_ASAP7_75t_L g2566 ( 
.A(n_2548),
.Y(n_2566)
);

AOI22xp5_ASAP7_75t_L g2567 ( 
.A1(n_2550),
.A2(n_2516),
.B1(n_2519),
.B2(n_2523),
.Y(n_2567)
);

INVx1_ASAP7_75t_L g2568 ( 
.A(n_2553),
.Y(n_2568)
);

AOI22xp5_ASAP7_75t_L g2569 ( 
.A1(n_2542),
.A2(n_2503),
.B1(n_2509),
.B2(n_2508),
.Y(n_2569)
);

AOI22xp5_ASAP7_75t_L g2570 ( 
.A1(n_2547),
.A2(n_2556),
.B1(n_2534),
.B2(n_2563),
.Y(n_2570)
);

NOR4xp25_ASAP7_75t_L g2571 ( 
.A(n_2544),
.B(n_2526),
.C(n_2528),
.D(n_2527),
.Y(n_2571)
);

AOI22xp5_ASAP7_75t_L g2572 ( 
.A1(n_2545),
.A2(n_2510),
.B1(n_2525),
.B2(n_2484),
.Y(n_2572)
);

INVx1_ASAP7_75t_L g2573 ( 
.A(n_2532),
.Y(n_2573)
);

NOR2xp33_ASAP7_75t_L g2574 ( 
.A(n_2536),
.B(n_2531),
.Y(n_2574)
);

AOI22xp5_ASAP7_75t_L g2575 ( 
.A1(n_2560),
.A2(n_2487),
.B1(n_2517),
.B2(n_2481),
.Y(n_2575)
);

INVx1_ASAP7_75t_L g2576 ( 
.A(n_2554),
.Y(n_2576)
);

NOR2xp33_ASAP7_75t_L g2577 ( 
.A(n_2541),
.B(n_2530),
.Y(n_2577)
);

AOI22xp5_ASAP7_75t_L g2578 ( 
.A1(n_2543),
.A2(n_2562),
.B1(n_2540),
.B2(n_2557),
.Y(n_2578)
);

AO22x2_ASAP7_75t_L g2579 ( 
.A1(n_2533),
.A2(n_2549),
.B1(n_2537),
.B2(n_2555),
.Y(n_2579)
);

NOR2xp33_ASAP7_75t_L g2580 ( 
.A(n_2538),
.B(n_2546),
.Y(n_2580)
);

INVx1_ASAP7_75t_L g2581 ( 
.A(n_2551),
.Y(n_2581)
);

AOI22xp5_ASAP7_75t_L g2582 ( 
.A1(n_2570),
.A2(n_2535),
.B1(n_2558),
.B2(n_2552),
.Y(n_2582)
);

AOI22xp5_ASAP7_75t_L g2583 ( 
.A1(n_2578),
.A2(n_2535),
.B1(n_2559),
.B2(n_2521),
.Y(n_2583)
);

NOR2x1_ASAP7_75t_L g2584 ( 
.A(n_2564),
.B(n_2391),
.Y(n_2584)
);

AOI22xp33_ASAP7_75t_L g2585 ( 
.A1(n_2569),
.A2(n_2505),
.B1(n_2506),
.B2(n_2504),
.Y(n_2585)
);

INVx2_ASAP7_75t_L g2586 ( 
.A(n_2568),
.Y(n_2586)
);

AOI22xp5_ASAP7_75t_L g2587 ( 
.A1(n_2567),
.A2(n_2398),
.B1(n_2399),
.B2(n_2397),
.Y(n_2587)
);

NOR2x1_ASAP7_75t_L g2588 ( 
.A(n_2565),
.B(n_2400),
.Y(n_2588)
);

NAND2xp5_ASAP7_75t_L g2589 ( 
.A(n_2576),
.B(n_2513),
.Y(n_2589)
);

NOR2x1_ASAP7_75t_L g2590 ( 
.A(n_2566),
.B(n_2522),
.Y(n_2590)
);

INVx2_ASAP7_75t_L g2591 ( 
.A(n_2588),
.Y(n_2591)
);

AO22x2_ASAP7_75t_L g2592 ( 
.A1(n_2586),
.A2(n_2573),
.B1(n_2581),
.B2(n_2589),
.Y(n_2592)
);

OA22x2_ASAP7_75t_L g2593 ( 
.A1(n_2582),
.A2(n_2575),
.B1(n_2572),
.B2(n_2571),
.Y(n_2593)
);

NOR2x1_ASAP7_75t_L g2594 ( 
.A(n_2584),
.B(n_2574),
.Y(n_2594)
);

NOR2x1_ASAP7_75t_L g2595 ( 
.A(n_2590),
.B(n_2580),
.Y(n_2595)
);

AND4x1_ASAP7_75t_L g2596 ( 
.A(n_2583),
.B(n_2577),
.C(n_2520),
.D(n_2579),
.Y(n_2596)
);

AOI22xp5_ASAP7_75t_L g2597 ( 
.A1(n_2585),
.A2(n_2511),
.B1(n_2406),
.B2(n_2529),
.Y(n_2597)
);

OAI22xp5_ASAP7_75t_L g2598 ( 
.A1(n_2587),
.A2(n_2512),
.B1(n_619),
.B2(n_615),
.Y(n_2598)
);

INVx1_ASAP7_75t_L g2599 ( 
.A(n_2595),
.Y(n_2599)
);

OR2x2_ASAP7_75t_L g2600 ( 
.A(n_2591),
.B(n_618),
.Y(n_2600)
);

INVx1_ASAP7_75t_L g2601 ( 
.A(n_2592),
.Y(n_2601)
);

HB1xp67_ASAP7_75t_L g2602 ( 
.A(n_2594),
.Y(n_2602)
);

INVx1_ASAP7_75t_L g2603 ( 
.A(n_2593),
.Y(n_2603)
);

OAI22xp5_ASAP7_75t_L g2604 ( 
.A1(n_2599),
.A2(n_2602),
.B1(n_2601),
.B2(n_2597),
.Y(n_2604)
);

HB1xp67_ASAP7_75t_L g2605 ( 
.A(n_2603),
.Y(n_2605)
);

HB1xp67_ASAP7_75t_L g2606 ( 
.A(n_2605),
.Y(n_2606)
);

AOI22xp5_ASAP7_75t_L g2607 ( 
.A1(n_2606),
.A2(n_2604),
.B1(n_2598),
.B2(n_2600),
.Y(n_2607)
);

INVx2_ASAP7_75t_L g2608 ( 
.A(n_2607),
.Y(n_2608)
);

AOI22xp33_ASAP7_75t_L g2609 ( 
.A1(n_2608),
.A2(n_2596),
.B1(n_622),
.B2(n_620),
.Y(n_2609)
);

INVx1_ASAP7_75t_L g2610 ( 
.A(n_2609),
.Y(n_2610)
);

OAI221xp5_ASAP7_75t_L g2611 ( 
.A1(n_2610),
.A2(n_624),
.B1(n_621),
.B2(n_623),
.C(n_625),
.Y(n_2611)
);

AOI211xp5_ASAP7_75t_L g2612 ( 
.A1(n_2611),
.A2(n_630),
.B(n_626),
.C(n_629),
.Y(n_2612)
);


endmodule