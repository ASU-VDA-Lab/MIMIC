module real_aes_4478_n_16 (n_13, n_4, n_0, n_3, n_5, n_2, n_15, n_7, n_8, n_6, n_9, n_12, n_1, n_14, n_10, n_11, n_16);
input n_13;
input n_4;
input n_0;
input n_3;
input n_5;
input n_2;
input n_15;
input n_7;
input n_8;
input n_6;
input n_9;
input n_12;
input n_1;
input n_14;
input n_10;
input n_11;
output n_16;
wire n_17;
wire n_28;
wire n_22;
wire n_24;
wire n_41;
wire n_34;
wire n_19;
wire n_40;
wire n_49;
wire n_46;
wire n_25;
wire n_47;
wire n_48;
wire n_43;
wire n_32;
wire n_30;
wire n_37;
wire n_35;
wire n_42;
wire n_39;
wire n_45;
wire n_27;
wire n_23;
wire n_38;
wire n_50;
wire n_29;
wire n_20;
wire n_44;
wire n_26;
wire n_18;
wire n_21;
wire n_31;
wire n_33;
wire n_36;
CKINVDCx5p33_ASAP7_75t_R g27 ( .A(n_0), .Y(n_27) );
AOI221xp5_ASAP7_75t_R g34 ( .A1(n_1), .A2(n_10), .B1(n_35), .B2(n_41), .C(n_43), .Y(n_34) );
CKINVDCx5p33_ASAP7_75t_R g26 ( .A(n_2), .Y(n_26) );
NOR2xp33_ASAP7_75t_R g45 ( .A(n_2), .B(n_6), .Y(n_45) );
NOR2xp33_ASAP7_75t_R g21 ( .A(n_3), .B(n_22), .Y(n_21) );
HB1xp67_ASAP7_75t_L g47 ( .A(n_4), .Y(n_47) );
NOR4xp25_ASAP7_75t_SL g19 ( .A(n_5), .B(n_20), .C(n_26), .D(n_27), .Y(n_19) );
CKINVDCx5p33_ASAP7_75t_R g33 ( .A(n_5), .Y(n_33) );
NAND2xp33_ASAP7_75t_R g39 ( .A(n_5), .B(n_21), .Y(n_39) );
NAND2xp33_ASAP7_75t_R g18 ( .A(n_6), .B(n_19), .Y(n_18) );
NAND3xp33_ASAP7_75t_SL g29 ( .A(n_6), .B(n_26), .C(n_30), .Y(n_29) );
NAND2xp33_ASAP7_75t_R g37 ( .A(n_6), .B(n_38), .Y(n_37) );
NOR2xp33_ASAP7_75t_R g41 ( .A(n_6), .B(n_42), .Y(n_41) );
CKINVDCx5p33_ASAP7_75t_R g49 ( .A(n_6), .Y(n_49) );
CKINVDCx5p33_ASAP7_75t_R g17 ( .A(n_7), .Y(n_17) );
CKINVDCx5p33_ASAP7_75t_R g28 ( .A(n_8), .Y(n_28) );
NAND3xp33_ASAP7_75t_SL g22 ( .A(n_9), .B(n_23), .C(n_24), .Y(n_22) );
CKINVDCx5p33_ASAP7_75t_R g50 ( .A(n_11), .Y(n_50) );
NOR2xp33_ASAP7_75t_R g25 ( .A(n_12), .B(n_13), .Y(n_25) );
NOR3xp33_ASAP7_75t_SL g30 ( .A(n_12), .B(n_31), .C(n_32), .Y(n_30) );
CKINVDCx5p33_ASAP7_75t_R g31 ( .A(n_13), .Y(n_31) );
CKINVDCx5p33_ASAP7_75t_R g23 ( .A(n_14), .Y(n_23) );
CKINVDCx5p33_ASAP7_75t_R g24 ( .A(n_15), .Y(n_24) );
OAI221xp5_ASAP7_75t_R g16 ( .A1(n_17), .A2(n_18), .B1(n_28), .B2(n_29), .C(n_34), .Y(n_16) );
NAND2xp33_ASAP7_75t_R g48 ( .A(n_19), .B(n_49), .Y(n_48) );
NAND2xp33_ASAP7_75t_R g20 ( .A(n_21), .B(n_25), .Y(n_20) );
NAND3xp33_ASAP7_75t_SL g32 ( .A(n_21), .B(n_27), .C(n_33), .Y(n_32) );
CKINVDCx5p33_ASAP7_75t_R g40 ( .A(n_25), .Y(n_40) );
NOR4xp25_ASAP7_75t_SL g38 ( .A(n_26), .B(n_27), .C(n_39), .D(n_40), .Y(n_38) );
NAND2xp33_ASAP7_75t_R g44 ( .A(n_30), .B(n_45), .Y(n_44) );
HB1xp67_ASAP7_75t_L g35 ( .A(n_36), .Y(n_35) );
CKINVDCx5p33_ASAP7_75t_R g36 ( .A(n_37), .Y(n_36) );
CKINVDCx5p33_ASAP7_75t_R g42 ( .A(n_38), .Y(n_42) );
OAI22xp33_ASAP7_75t_L g43 ( .A1(n_44), .A2(n_46), .B1(n_48), .B2(n_50), .Y(n_43) );
CKINVDCx5p33_ASAP7_75t_R g46 ( .A(n_47), .Y(n_46) );
endmodule