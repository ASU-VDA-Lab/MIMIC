module fake_jpeg_16107_n_167 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_167);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_167;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g48 ( 
.A(n_0),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_4),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_29),
.Y(n_50)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_40),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_37),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_47),
.Y(n_53)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_44),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_46),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_36),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_13),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_39),
.Y(n_58)
);

BUFx2_ASAP7_75t_L g59 ( 
.A(n_41),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_3),
.Y(n_60)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_38),
.Y(n_61)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_34),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_18),
.Y(n_63)
);

INVx6_ASAP7_75t_SL g64 ( 
.A(n_0),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_31),
.Y(n_65)
);

BUFx8_ASAP7_75t_L g66 ( 
.A(n_8),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_10),
.Y(n_67)
);

BUFx8_ASAP7_75t_L g68 ( 
.A(n_59),
.Y(n_68)
);

INVx1_ASAP7_75t_SL g82 ( 
.A(n_68),
.Y(n_82)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_51),
.Y(n_69)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_69),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_63),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_70),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_62),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_71),
.A2(n_62),
.B1(n_61),
.B2(n_48),
.Y(n_85)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_51),
.Y(n_72)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_72),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_63),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_73),
.Y(n_90)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_51),
.Y(n_74)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_74),
.Y(n_84)
);

BUFx5_ASAP7_75t_L g75 ( 
.A(n_54),
.Y(n_75)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_75),
.Y(n_77)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_54),
.Y(n_76)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_76),
.Y(n_86)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_70),
.Y(n_79)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_79),
.Y(n_97)
);

BUFx2_ASAP7_75t_L g83 ( 
.A(n_68),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_83),
.B(n_67),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_L g99 ( 
.A1(n_85),
.A2(n_66),
.B1(n_67),
.B2(n_57),
.Y(n_99)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_73),
.Y(n_87)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_87),
.Y(n_103)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_71),
.Y(n_88)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_88),
.Y(n_107)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_70),
.Y(n_89)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_89),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_70),
.Y(n_91)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_91),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_68),
.B(n_49),
.Y(n_92)
);

AND2x2_ASAP7_75t_L g102 ( 
.A(n_92),
.B(n_1),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_70),
.Y(n_93)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_93),
.Y(n_104)
);

O2A1O1Ixp33_ASAP7_75t_SL g94 ( 
.A1(n_92),
.A2(n_54),
.B(n_66),
.C(n_59),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_94),
.A2(n_108),
.B1(n_60),
.B2(n_5),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_80),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_96),
.B(n_105),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_78),
.A2(n_64),
.B1(n_65),
.B2(n_50),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_98),
.A2(n_101),
.B1(n_90),
.B2(n_6),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_99),
.A2(n_111),
.B1(n_112),
.B2(n_91),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_77),
.A2(n_65),
.B1(n_50),
.B2(n_66),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_102),
.B(n_113),
.Y(n_117)
);

CKINVDCx16_ASAP7_75t_R g105 ( 
.A(n_83),
.Y(n_105)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_84),
.Y(n_106)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_106),
.Y(n_114)
);

AND2x2_ASAP7_75t_L g108 ( 
.A(n_82),
.B(n_2),
.Y(n_108)
);

CKINVDCx16_ASAP7_75t_R g119 ( 
.A(n_109),
.Y(n_119)
);

BUFx5_ASAP7_75t_L g110 ( 
.A(n_86),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_110),
.Y(n_116)
);

OAI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_81),
.A2(n_60),
.B1(n_57),
.B2(n_55),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_81),
.A2(n_58),
.B1(n_56),
.B2(n_53),
.Y(n_112)
);

OR2x2_ASAP7_75t_L g113 ( 
.A(n_93),
.B(n_52),
.Y(n_113)
);

XNOR2xp5_ASAP7_75t_L g133 ( 
.A(n_115),
.B(n_111),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_102),
.B(n_4),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_120),
.B(n_123),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_107),
.A2(n_21),
.B1(n_45),
.B2(n_43),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_121),
.A2(n_124),
.B1(n_108),
.B2(n_104),
.Y(n_127)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_100),
.Y(n_122)
);

INVxp67_ASAP7_75t_L g132 ( 
.A(n_122),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_113),
.Y(n_123)
);

INVx3_ASAP7_75t_L g125 ( 
.A(n_95),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_125),
.B(n_104),
.Y(n_131)
);

AOI21xp5_ASAP7_75t_L g130 ( 
.A1(n_126),
.A2(n_101),
.B(n_98),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_127),
.A2(n_99),
.B1(n_121),
.B2(n_119),
.Y(n_135)
);

AND2x2_ASAP7_75t_SL g128 ( 
.A(n_117),
.B(n_94),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_128),
.B(n_130),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_131),
.Y(n_138)
);

XOR2xp5_ASAP7_75t_L g134 ( 
.A(n_133),
.B(n_115),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_134),
.B(n_128),
.C(n_118),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_135),
.A2(n_128),
.B1(n_124),
.B2(n_129),
.Y(n_139)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_132),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_136),
.B(n_132),
.Y(n_140)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_139),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_140),
.B(n_141),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_138),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_SL g149 ( 
.A1(n_142),
.A2(n_143),
.B(n_19),
.Y(n_149)
);

AOI32xp33_ASAP7_75t_L g143 ( 
.A1(n_137),
.A2(n_116),
.A3(n_27),
.B1(n_23),
.B2(n_42),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_135),
.A2(n_125),
.B1(n_122),
.B2(n_116),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_144),
.A2(n_136),
.B1(n_114),
.B2(n_103),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_144),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_SL g150 ( 
.A(n_146),
.B(n_134),
.Y(n_150)
);

AOI322xp5_ASAP7_75t_L g151 ( 
.A1(n_147),
.A2(n_149),
.A3(n_97),
.B1(n_17),
.B2(n_35),
.C1(n_33),
.C2(n_32),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_150),
.A2(n_148),
.B1(n_141),
.B2(n_145),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_151),
.B(n_152),
.C(n_90),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_147),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_153),
.A2(n_154),
.B1(n_30),
.B2(n_28),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_155),
.B(n_26),
.Y(n_156)
);

XOR2xp5_ASAP7_75t_L g157 ( 
.A(n_156),
.B(n_25),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_157),
.B(n_24),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_158),
.A2(n_22),
.B1(n_20),
.B2(n_16),
.Y(n_159)
);

AOI21xp5_ASAP7_75t_L g160 ( 
.A1(n_159),
.A2(n_15),
.B(n_6),
.Y(n_160)
);

AOI21xp5_ASAP7_75t_L g161 ( 
.A1(n_160),
.A2(n_5),
.B(n_7),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_161),
.B(n_7),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_162),
.B(n_8),
.Y(n_163)
);

AOI21x1_ASAP7_75t_L g164 ( 
.A1(n_163),
.A2(n_9),
.B(n_10),
.Y(n_164)
);

AO21x1_ASAP7_75t_L g165 ( 
.A1(n_164),
.A2(n_9),
.B(n_11),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_165),
.B(n_11),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_L g167 ( 
.A1(n_166),
.A2(n_12),
.B1(n_13),
.B2(n_14),
.Y(n_167)
);


endmodule