module fake_jpeg_12932_n_383 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_383);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_383;

wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx11_ASAP7_75t_L g15 ( 
.A(n_6),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

INVx6_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

INVx3_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

INVx8_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

INVx11_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

INVx6_ASAP7_75t_SL g33 ( 
.A(n_2),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_9),
.Y(n_34)
);

INVxp67_ASAP7_75t_L g35 ( 
.A(n_7),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_33),
.Y(n_36)
);

INVx5_ASAP7_75t_L g61 ( 
.A(n_36),
.Y(n_61)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_18),
.Y(n_37)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_37),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_18),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_38),
.Y(n_86)
);

BUFx12_ASAP7_75t_L g39 ( 
.A(n_33),
.Y(n_39)
);

INVx5_ASAP7_75t_L g66 ( 
.A(n_39),
.Y(n_66)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_18),
.Y(n_40)
);

INVx5_ASAP7_75t_L g81 ( 
.A(n_40),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_35),
.B(n_7),
.Y(n_41)
);

AND2x2_ASAP7_75t_L g70 ( 
.A(n_41),
.B(n_48),
.Y(n_70)
);

BUFx16f_ASAP7_75t_L g42 ( 
.A(n_33),
.Y(n_42)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_42),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_18),
.Y(n_43)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_43),
.Y(n_74)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_19),
.Y(n_44)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_44),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_26),
.Y(n_45)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_45),
.Y(n_91)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_20),
.Y(n_46)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_46),
.Y(n_85)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_22),
.Y(n_47)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_47),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_34),
.B(n_7),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_SL g49 ( 
.A(n_22),
.B(n_6),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_49),
.B(n_0),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_15),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_50),
.B(n_58),
.Y(n_88)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_20),
.Y(n_51)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_51),
.Y(n_62)
);

HB1xp67_ASAP7_75t_L g52 ( 
.A(n_22),
.Y(n_52)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_52),
.Y(n_64)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_23),
.Y(n_53)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_53),
.Y(n_65)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_20),
.Y(n_54)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_54),
.Y(n_71)
);

INVx4_ASAP7_75t_SL g55 ( 
.A(n_15),
.Y(n_55)
);

INVx11_ASAP7_75t_L g87 ( 
.A(n_55),
.Y(n_87)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_19),
.Y(n_56)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_56),
.Y(n_73)
);

INVx11_ASAP7_75t_L g57 ( 
.A(n_15),
.Y(n_57)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_57),
.Y(n_82)
);

BUFx16f_ASAP7_75t_L g58 ( 
.A(n_15),
.Y(n_58)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_23),
.Y(n_59)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_59),
.Y(n_77)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_63),
.B(n_0),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g67 ( 
.A1(n_49),
.A2(n_23),
.B1(n_19),
.B2(n_34),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_67),
.A2(n_31),
.B1(n_28),
.B2(n_25),
.Y(n_101)
);

OR2x2_ASAP7_75t_SL g69 ( 
.A(n_41),
.B(n_32),
.Y(n_69)
);

OR2x2_ASAP7_75t_L g114 ( 
.A(n_69),
.B(n_89),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_48),
.B(n_34),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g107 ( 
.A(n_75),
.B(n_76),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_47),
.B(n_16),
.Y(n_76)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_53),
.Y(n_78)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_78),
.Y(n_99)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_59),
.Y(n_80)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_80),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_36),
.A2(n_26),
.B1(n_32),
.B2(n_19),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_83),
.A2(n_84),
.B1(n_32),
.B2(n_31),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_L g84 ( 
.A1(n_37),
.A2(n_26),
.B1(n_31),
.B2(n_30),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_46),
.B(n_16),
.Y(n_89)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_37),
.Y(n_90)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_90),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_70),
.B(n_36),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g140 ( 
.A(n_92),
.B(n_94),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_83),
.A2(n_40),
.B1(n_43),
.B2(n_38),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_93),
.A2(n_98),
.B1(n_112),
.B2(n_57),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_70),
.B(n_36),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_69),
.B(n_50),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_95),
.B(n_97),
.Y(n_130)
);

BUFx12f_ASAP7_75t_L g96 ( 
.A(n_87),
.Y(n_96)
);

INVx3_ASAP7_75t_L g146 ( 
.A(n_96),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_88),
.B(n_27),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_64),
.A2(n_40),
.B1(n_43),
.B2(n_38),
.Y(n_98)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_85),
.Y(n_100)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_100),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_101),
.A2(n_126),
.B1(n_28),
.B2(n_24),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_60),
.B(n_17),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_102),
.B(n_115),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_87),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_103),
.B(n_104),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_68),
.Y(n_104)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_73),
.Y(n_105)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_105),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_L g158 ( 
.A(n_106),
.B(n_21),
.Y(n_158)
);

AND2x2_ASAP7_75t_L g108 ( 
.A(n_65),
.B(n_54),
.Y(n_108)
);

CKINVDCx16_ASAP7_75t_R g147 ( 
.A(n_108),
.Y(n_147)
);

INVx1_ASAP7_75t_SL g109 ( 
.A(n_62),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_109),
.B(n_117),
.Y(n_134)
);

OA22x2_ASAP7_75t_L g111 ( 
.A1(n_91),
.A2(n_56),
.B1(n_44),
.B2(n_45),
.Y(n_111)
);

INVx3_ASAP7_75t_SL g150 ( 
.A(n_111),
.Y(n_150)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_79),
.Y(n_113)
);

BUFx2_ASAP7_75t_L g160 ( 
.A(n_113),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_77),
.B(n_25),
.Y(n_115)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_61),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_71),
.B(n_62),
.C(n_73),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_118),
.B(n_122),
.C(n_125),
.Y(n_135)
);

BUFx3_ASAP7_75t_L g119 ( 
.A(n_68),
.Y(n_119)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_119),
.Y(n_138)
);

AOI21xp5_ASAP7_75t_SL g120 ( 
.A1(n_61),
.A2(n_25),
.B(n_17),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_L g148 ( 
.A1(n_120),
.A2(n_29),
.B(n_24),
.Y(n_148)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_74),
.Y(n_121)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_121),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_71),
.B(n_45),
.C(n_51),
.Y(n_122)
);

BUFx8_ASAP7_75t_L g123 ( 
.A(n_66),
.Y(n_123)
);

INVxp67_ASAP7_75t_L g141 ( 
.A(n_123),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_66),
.B(n_42),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_124),
.B(n_96),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_90),
.B(n_21),
.C(n_17),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_L g126 ( 
.A1(n_74),
.A2(n_44),
.B1(n_56),
.B2(n_26),
.Y(n_126)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_81),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_127),
.B(n_79),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_114),
.A2(n_72),
.B1(n_91),
.B2(n_86),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_128),
.A2(n_154),
.B1(n_156),
.B2(n_100),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_SL g129 ( 
.A(n_95),
.B(n_32),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_129),
.B(n_120),
.C(n_111),
.Y(n_176)
);

CKINVDCx14_ASAP7_75t_R g182 ( 
.A(n_131),
.Y(n_182)
);

OAI22xp33_ASAP7_75t_SL g187 ( 
.A1(n_133),
.A2(n_55),
.B1(n_117),
.B2(n_21),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_93),
.A2(n_72),
.B1(n_81),
.B2(n_86),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_136),
.A2(n_133),
.B1(n_150),
.B2(n_144),
.Y(n_164)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_139),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_102),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_142),
.B(n_159),
.Y(n_161)
);

NAND2xp33_ASAP7_75t_SL g143 ( 
.A(n_115),
.B(n_16),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_SL g185 ( 
.A1(n_143),
.A2(n_153),
.B(n_157),
.Y(n_185)
);

AOI22xp33_ASAP7_75t_L g144 ( 
.A1(n_98),
.A2(n_82),
.B1(n_30),
.B2(n_29),
.Y(n_144)
);

AO21x2_ASAP7_75t_L g191 ( 
.A1(n_144),
.A2(n_96),
.B(n_58),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_107),
.B(n_82),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_145),
.B(n_155),
.Y(n_170)
);

CKINVDCx16_ASAP7_75t_R g190 ( 
.A(n_148),
.Y(n_190)
);

AOI21xp5_ASAP7_75t_L g153 ( 
.A1(n_114),
.A2(n_103),
.B(n_125),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_101),
.A2(n_29),
.B1(n_24),
.B2(n_27),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_106),
.B(n_30),
.Y(n_155)
);

AOI21xp5_ASAP7_75t_L g157 ( 
.A1(n_97),
.A2(n_28),
.B(n_27),
.Y(n_157)
);

MAJx2_ASAP7_75t_L g181 ( 
.A(n_158),
.B(n_109),
.C(n_110),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_108),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g219 ( 
.A1(n_162),
.A2(n_166),
.B1(n_168),
.B2(n_172),
.Y(n_219)
);

INVxp67_ASAP7_75t_L g163 ( 
.A(n_134),
.Y(n_163)
);

HB1xp67_ASAP7_75t_L g204 ( 
.A(n_163),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_164),
.A2(n_187),
.B1(n_156),
.B2(n_147),
.Y(n_202)
);

INVxp67_ASAP7_75t_L g165 ( 
.A(n_134),
.Y(n_165)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_165),
.Y(n_205)
);

AOI22xp33_ASAP7_75t_L g166 ( 
.A1(n_150),
.A2(n_111),
.B1(n_108),
.B2(n_121),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_150),
.A2(n_107),
.B1(n_106),
.B2(n_122),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_140),
.B(n_104),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_SL g210 ( 
.A(n_169),
.B(n_174),
.Y(n_210)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_149),
.Y(n_171)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_171),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_142),
.A2(n_111),
.B1(n_118),
.B2(n_99),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_132),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_173),
.B(n_175),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_140),
.B(n_119),
.Y(n_174)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_152),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_176),
.B(n_181),
.Y(n_200)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_152),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_177),
.B(n_194),
.Y(n_208)
);

INVxp67_ASAP7_75t_L g178 ( 
.A(n_131),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_178),
.B(n_193),
.Y(n_209)
);

AO22x1_ASAP7_75t_L g179 ( 
.A1(n_148),
.A2(n_105),
.B1(n_99),
.B2(n_110),
.Y(n_179)
);

AOI21xp5_ASAP7_75t_SL g223 ( 
.A1(n_179),
.A2(n_191),
.B(n_176),
.Y(n_223)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_149),
.Y(n_180)
);

AND2x2_ASAP7_75t_L g230 ( 
.A(n_180),
.B(n_186),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_128),
.A2(n_113),
.B1(n_116),
.B2(n_127),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_183),
.A2(n_191),
.B1(n_195),
.B2(n_147),
.Y(n_199)
);

FAx1_ASAP7_75t_SL g184 ( 
.A(n_130),
.B(n_116),
.CI(n_55),
.CON(n_184),
.SN(n_184)
);

AOI31xp33_ASAP7_75t_SL g225 ( 
.A1(n_184),
.A2(n_146),
.A3(n_8),
.B(n_2),
.Y(n_225)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_151),
.Y(n_186)
);

OAI22x1_ASAP7_75t_L g188 ( 
.A1(n_136),
.A2(n_39),
.B1(n_42),
.B2(n_123),
.Y(n_188)
);

AOI22xp33_ASAP7_75t_SL g220 ( 
.A1(n_188),
.A2(n_192),
.B1(n_146),
.B2(n_138),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_135),
.B(n_123),
.C(n_96),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_189),
.B(n_146),
.C(n_1),
.Y(n_221)
);

AOI22xp33_ASAP7_75t_L g192 ( 
.A1(n_159),
.A2(n_39),
.B1(n_58),
.B2(n_123),
.Y(n_192)
);

INVxp67_ASAP7_75t_L g193 ( 
.A(n_160),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_137),
.B(n_0),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_137),
.A2(n_39),
.B1(n_8),
.B2(n_2),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_151),
.Y(n_196)
);

INVxp67_ASAP7_75t_L g222 ( 
.A(n_196),
.Y(n_222)
);

AOI22x1_ASAP7_75t_SL g197 ( 
.A1(n_190),
.A2(n_153),
.B1(n_129),
.B2(n_130),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_SL g255 ( 
.A1(n_197),
.A2(n_223),
.B(n_225),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_L g198 ( 
.A(n_189),
.B(n_135),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_198),
.B(n_207),
.C(n_214),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_199),
.A2(n_163),
.B1(n_184),
.B2(n_179),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_202),
.B(n_212),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_161),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g262 ( 
.A(n_203),
.B(n_211),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_164),
.A2(n_154),
.B1(n_129),
.B2(n_145),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_206),
.A2(n_172),
.B1(n_184),
.B2(n_183),
.Y(n_244)
);

XOR2xp5_ASAP7_75t_L g207 ( 
.A(n_170),
.B(n_132),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_171),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_173),
.B(n_143),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_167),
.B(n_155),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_213),
.B(n_216),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g214 ( 
.A(n_170),
.B(n_158),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g215 ( 
.A(n_185),
.B(n_157),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_215),
.B(n_221),
.C(n_231),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_167),
.B(n_139),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_194),
.B(n_160),
.Y(n_217)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_217),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_168),
.A2(n_160),
.B1(n_141),
.B2(n_138),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_218),
.A2(n_229),
.B1(n_199),
.B2(n_227),
.Y(n_232)
);

CKINVDCx16_ASAP7_75t_R g236 ( 
.A(n_220),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_180),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_224),
.B(n_226),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_186),
.Y(n_226)
);

OAI21xp5_ASAP7_75t_L g227 ( 
.A1(n_178),
.A2(n_8),
.B(n_12),
.Y(n_227)
);

CKINVDCx16_ASAP7_75t_R g257 ( 
.A(n_227),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_162),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_185),
.B(n_10),
.Y(n_231)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_232),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_SL g234 ( 
.A(n_210),
.B(n_165),
.Y(n_234)
);

NAND3xp33_ASAP7_75t_L g269 ( 
.A(n_234),
.B(n_213),
.C(n_208),
.Y(n_269)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_228),
.Y(n_237)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_237),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_SL g238 ( 
.A(n_200),
.B(n_182),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_238),
.B(n_240),
.C(n_247),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_230),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_SL g270 ( 
.A(n_239),
.B(n_241),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_SL g240 ( 
.A(n_200),
.B(n_181),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_230),
.Y(n_241)
);

CKINVDCx14_ASAP7_75t_R g242 ( 
.A(n_209),
.Y(n_242)
);

CKINVDCx14_ASAP7_75t_R g286 ( 
.A(n_242),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_243),
.A2(n_250),
.B1(n_202),
.B2(n_201),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_244),
.A2(n_256),
.B1(n_229),
.B2(n_231),
.Y(n_275)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_198),
.B(n_196),
.Y(n_247)
);

INVx6_ASAP7_75t_L g248 ( 
.A(n_204),
.Y(n_248)
);

INVx3_ASAP7_75t_L g272 ( 
.A(n_248),
.Y(n_272)
);

INVx3_ASAP7_75t_L g249 ( 
.A(n_205),
.Y(n_249)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_249),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_219),
.A2(n_179),
.B1(n_191),
.B2(n_177),
.Y(n_250)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_228),
.Y(n_251)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_251),
.Y(n_266)
);

OAI32xp33_ASAP7_75t_L g252 ( 
.A1(n_216),
.A2(n_175),
.A3(n_191),
.B1(n_195),
.B2(n_188),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_252),
.B(n_218),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_206),
.A2(n_191),
.B1(n_193),
.B2(n_1),
.Y(n_256)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_207),
.B(n_10),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_258),
.B(n_260),
.C(n_221),
.Y(n_287)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_230),
.Y(n_259)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_259),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_197),
.B(n_10),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_201),
.Y(n_261)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_261),
.Y(n_281)
);

AO21x1_ASAP7_75t_L g264 ( 
.A1(n_233),
.A2(n_212),
.B(n_223),
.Y(n_264)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_264),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_235),
.B(n_215),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_L g302 ( 
.A(n_268),
.B(n_285),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_269),
.B(n_260),
.Y(n_290)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_271),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_245),
.B(n_254),
.Y(n_273)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_273),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_262),
.B(n_253),
.Y(n_274)
);

NAND3xp33_ASAP7_75t_L g292 ( 
.A(n_274),
.B(n_283),
.C(n_289),
.Y(n_292)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_275),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_245),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_SL g298 ( 
.A(n_276),
.B(n_287),
.Y(n_298)
);

INVxp67_ASAP7_75t_SL g277 ( 
.A(n_237),
.Y(n_277)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_277),
.Y(n_296)
);

INVxp67_ASAP7_75t_L g278 ( 
.A(n_233),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_278),
.B(n_232),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_279),
.A2(n_263),
.B1(n_278),
.B2(n_271),
.Y(n_304)
);

OAI21xp5_ASAP7_75t_L g282 ( 
.A1(n_243),
.A2(n_225),
.B(n_222),
.Y(n_282)
);

OAI21xp5_ASAP7_75t_SL g310 ( 
.A1(n_282),
.A2(n_257),
.B(n_250),
.Y(n_310)
);

AOI31xp33_ASAP7_75t_L g283 ( 
.A1(n_238),
.A2(n_208),
.A3(n_217),
.B(n_222),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_235),
.B(n_214),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g288 ( 
.A(n_247),
.B(n_10),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_288),
.B(n_246),
.C(n_258),
.Y(n_291)
);

NAND3xp33_ASAP7_75t_L g289 ( 
.A(n_255),
.B(n_14),
.C(n_4),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_SL g317 ( 
.A(n_290),
.B(n_291),
.Y(n_317)
);

XNOR2xp5_ASAP7_75t_L g294 ( 
.A(n_285),
.B(n_240),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_L g315 ( 
.A(n_294),
.B(n_303),
.Y(n_315)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_300),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_268),
.B(n_246),
.C(n_244),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_301),
.B(n_312),
.C(n_287),
.Y(n_318)
);

XNOR2xp5_ASAP7_75t_SL g303 ( 
.A(n_284),
.B(n_255),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_SL g321 ( 
.A1(n_304),
.A2(n_264),
.B1(n_281),
.B2(n_282),
.Y(n_321)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_270),
.Y(n_305)
);

BUFx2_ASAP7_75t_L g319 ( 
.A(n_305),
.Y(n_319)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_266),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_306),
.B(n_311),
.Y(n_324)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_280),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_307),
.B(n_308),
.Y(n_316)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_273),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_286),
.B(n_248),
.Y(n_309)
);

INVxp67_ASAP7_75t_L g322 ( 
.A(n_309),
.Y(n_322)
);

OR2x2_ASAP7_75t_L g320 ( 
.A(n_310),
.B(n_275),
.Y(n_320)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_267),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_284),
.B(n_249),
.C(n_251),
.Y(n_312)
);

OAI21xp5_ASAP7_75t_L g313 ( 
.A1(n_300),
.A2(n_279),
.B(n_263),
.Y(n_313)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_313),
.Y(n_336)
);

INVx13_ASAP7_75t_L g314 ( 
.A(n_296),
.Y(n_314)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_314),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_SL g332 ( 
.A(n_318),
.B(n_323),
.Y(n_332)
);

OAI21xp5_ASAP7_75t_SL g335 ( 
.A1(n_320),
.A2(n_293),
.B(n_297),
.Y(n_335)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_321),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_302),
.B(n_288),
.C(n_267),
.Y(n_323)
);

OAI322xp33_ASAP7_75t_L g325 ( 
.A1(n_292),
.A2(n_265),
.A3(n_236),
.B1(n_252),
.B2(n_256),
.C1(n_272),
.C2(n_12),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_SL g344 ( 
.A(n_325),
.B(n_326),
.Y(n_344)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_302),
.B(n_272),
.C(n_1),
.Y(n_326)
);

OAI22xp5_ASAP7_75t_L g327 ( 
.A1(n_304),
.A2(n_4),
.B1(n_5),
.B2(n_9),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_327),
.B(n_311),
.Y(n_338)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_312),
.B(n_1),
.C(n_4),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_328),
.B(n_291),
.C(n_298),
.Y(n_331)
);

FAx1_ASAP7_75t_SL g329 ( 
.A(n_301),
.B(n_4),
.CI(n_5),
.CON(n_329),
.SN(n_329)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_329),
.B(n_319),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_331),
.B(n_333),
.Y(n_353)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_318),
.B(n_294),
.C(n_299),
.Y(n_333)
);

OAI22xp5_ASAP7_75t_L g334 ( 
.A1(n_319),
.A2(n_297),
.B1(n_299),
.B2(n_295),
.Y(n_334)
);

AOI22xp5_ASAP7_75t_L g354 ( 
.A1(n_334),
.A2(n_340),
.B1(n_330),
.B2(n_327),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_SL g346 ( 
.A(n_335),
.B(n_339),
.Y(n_346)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_338),
.Y(n_349)
);

OAI22xp5_ASAP7_75t_SL g340 ( 
.A1(n_320),
.A2(n_293),
.B1(n_310),
.B2(n_306),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_L g341 ( 
.A(n_319),
.B(n_303),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_SL g352 ( 
.A(n_341),
.B(n_342),
.Y(n_352)
);

NOR2xp33_ASAP7_75t_L g342 ( 
.A(n_316),
.B(n_5),
.Y(n_342)
);

XNOR2x1_ASAP7_75t_L g345 ( 
.A(n_315),
.B(n_14),
.Y(n_345)
);

MAJIxp5_ASAP7_75t_L g350 ( 
.A(n_345),
.B(n_328),
.C(n_322),
.Y(n_350)
);

AOI22xp5_ASAP7_75t_SL g347 ( 
.A1(n_336),
.A2(n_321),
.B1(n_330),
.B2(n_322),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_347),
.B(n_350),
.Y(n_359)
);

AND2x2_ASAP7_75t_L g348 ( 
.A(n_344),
.B(n_326),
.Y(n_348)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_348),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_SL g351 ( 
.A(n_336),
.B(n_340),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_351),
.B(n_354),
.Y(n_366)
);

OAI21x1_ASAP7_75t_L g355 ( 
.A1(n_331),
.A2(n_324),
.B(n_329),
.Y(n_355)
);

OAI21xp5_ASAP7_75t_SL g360 ( 
.A1(n_355),
.A2(n_356),
.B(n_343),
.Y(n_360)
);

AOI21xp5_ASAP7_75t_SL g356 ( 
.A1(n_335),
.A2(n_317),
.B(n_313),
.Y(n_356)
);

MAJIxp5_ASAP7_75t_L g357 ( 
.A(n_332),
.B(n_323),
.C(n_315),
.Y(n_357)
);

NOR2xp33_ASAP7_75t_L g361 ( 
.A(n_357),
.B(n_329),
.Y(n_361)
);

OAI21xp5_ASAP7_75t_SL g358 ( 
.A1(n_346),
.A2(n_343),
.B(n_333),
.Y(n_358)
);

NAND2x1p5_ASAP7_75t_L g370 ( 
.A(n_358),
.B(n_360),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_361),
.B(n_362),
.Y(n_367)
);

NOR2xp33_ASAP7_75t_L g362 ( 
.A(n_352),
.B(n_337),
.Y(n_362)
);

OAI21xp5_ASAP7_75t_SL g363 ( 
.A1(n_353),
.A2(n_337),
.B(n_324),
.Y(n_363)
);

AOI21xp5_ASAP7_75t_SL g372 ( 
.A1(n_363),
.A2(n_5),
.B(n_11),
.Y(n_372)
);

OAI22xp5_ASAP7_75t_SL g365 ( 
.A1(n_349),
.A2(n_338),
.B1(n_345),
.B2(n_314),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_365),
.B(n_11),
.Y(n_373)
);

OAI21xp5_ASAP7_75t_L g368 ( 
.A1(n_359),
.A2(n_346),
.B(n_348),
.Y(n_368)
);

HB1xp67_ASAP7_75t_L g375 ( 
.A(n_368),
.Y(n_375)
);

OAI21xp5_ASAP7_75t_SL g369 ( 
.A1(n_364),
.A2(n_351),
.B(n_9),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_L g374 ( 
.A(n_369),
.B(n_371),
.Y(n_374)
);

CKINVDCx20_ASAP7_75t_R g371 ( 
.A(n_366),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_L g376 ( 
.A(n_372),
.B(n_373),
.Y(n_376)
);

OAI31xp67_ASAP7_75t_L g377 ( 
.A1(n_370),
.A2(n_358),
.A3(n_365),
.B(n_12),
.Y(n_377)
);

INVxp33_ASAP7_75t_L g379 ( 
.A(n_377),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_375),
.B(n_367),
.Y(n_378)
);

MAJIxp5_ASAP7_75t_L g380 ( 
.A(n_378),
.B(n_369),
.C(n_376),
.Y(n_380)
);

NAND3xp33_ASAP7_75t_L g381 ( 
.A(n_380),
.B(n_374),
.C(n_379),
.Y(n_381)
);

XOR2xp5_ASAP7_75t_L g382 ( 
.A(n_381),
.B(n_14),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_382),
.B(n_14),
.Y(n_383)
);


endmodule