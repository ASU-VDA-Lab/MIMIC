module fake_jpeg_9186_n_259 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_259);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_259;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_223;
wire n_187;
wire n_21;
wire n_57;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_212;
wire n_131;
wire n_56;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_192;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_96;

INVx6_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_5),
.Y(n_19)
);

INVx1_ASAP7_75t_SL g20 ( 
.A(n_2),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_15),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_9),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_16),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

INVx2_ASAP7_75t_SL g26 ( 
.A(n_1),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_10),
.Y(n_27)
);

CKINVDCx14_ASAP7_75t_R g28 ( 
.A(n_4),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_3),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_16),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_20),
.B(n_0),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_SL g50 ( 
.A(n_34),
.B(n_35),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_20),
.B(n_1),
.Y(n_35)
);

BUFx12_ASAP7_75t_L g36 ( 
.A(n_25),
.Y(n_36)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_36),
.Y(n_42)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_25),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_37),
.B(n_38),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_20),
.B(n_1),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_25),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_39),
.Y(n_52)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_33),
.Y(n_40)
);

INVx8_ASAP7_75t_L g49 ( 
.A(n_40),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_33),
.Y(n_41)
);

INVx5_ASAP7_75t_L g43 ( 
.A(n_41),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_L g44 ( 
.A1(n_37),
.A2(n_17),
.B1(n_18),
.B2(n_26),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_44),
.A2(n_45),
.B1(n_55),
.B2(n_31),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g45 ( 
.A1(n_37),
.A2(n_18),
.B1(n_17),
.B2(n_26),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_34),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_46),
.B(n_28),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_34),
.B(n_32),
.Y(n_48)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_48),
.Y(n_59)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_41),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_51),
.B(n_36),
.Y(n_82)
);

BUFx2_ASAP7_75t_L g53 ( 
.A(n_41),
.Y(n_53)
);

INVx5_ASAP7_75t_SL g72 ( 
.A(n_53),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_35),
.B(n_21),
.Y(n_54)
);

AND2x2_ASAP7_75t_L g71 ( 
.A(n_54),
.B(n_2),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g55 ( 
.A1(n_40),
.A2(n_17),
.B1(n_26),
.B2(n_31),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_38),
.B(n_32),
.Y(n_56)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_56),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_39),
.B(n_30),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_57),
.B(n_39),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g58 ( 
.A(n_56),
.B(n_24),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_58),
.B(n_63),
.Y(n_94)
);

INVxp67_ASAP7_75t_L g60 ( 
.A(n_57),
.Y(n_60)
);

CKINVDCx16_ASAP7_75t_R g113 ( 
.A(n_60),
.Y(n_113)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_53),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_61),
.Y(n_106)
);

INVx5_ASAP7_75t_L g62 ( 
.A(n_43),
.Y(n_62)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_62),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_SL g63 ( 
.A(n_48),
.B(n_24),
.Y(n_63)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_64),
.Y(n_95)
);

BUFx12f_ASAP7_75t_L g65 ( 
.A(n_53),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_65),
.B(n_66),
.Y(n_108)
);

HB1xp67_ASAP7_75t_L g66 ( 
.A(n_51),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_46),
.B(n_21),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_67),
.B(n_69),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_51),
.Y(n_68)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_68),
.Y(n_115)
);

INVx5_ASAP7_75t_L g69 ( 
.A(n_43),
.Y(n_69)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_43),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_70),
.Y(n_109)
);

AND2x2_ASAP7_75t_L g114 ( 
.A(n_71),
.B(n_78),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_46),
.A2(n_26),
.B1(n_40),
.B2(n_23),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_73),
.A2(n_79),
.B1(n_84),
.B2(n_88),
.Y(n_101)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_45),
.Y(n_74)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_74),
.Y(n_96)
);

INVx8_ASAP7_75t_L g75 ( 
.A(n_42),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_75),
.A2(n_86),
.B1(n_89),
.B2(n_90),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_50),
.B(n_19),
.Y(n_76)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_76),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_54),
.B(n_19),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_77),
.B(n_87),
.Y(n_100)
);

AND2x2_ASAP7_75t_L g78 ( 
.A(n_47),
.B(n_50),
.Y(n_78)
);

OAI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_57),
.A2(n_40),
.B1(n_28),
.B2(n_23),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_80),
.A2(n_22),
.B1(n_49),
.B2(n_30),
.Y(n_92)
);

INVx1_ASAP7_75t_SL g81 ( 
.A(n_42),
.Y(n_81)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_81),
.Y(n_105)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_82),
.Y(n_107)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_55),
.Y(n_83)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_83),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_L g84 ( 
.A1(n_47),
.A2(n_27),
.B1(n_22),
.B2(n_30),
.Y(n_84)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_44),
.Y(n_86)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_53),
.Y(n_87)
);

OAI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_49),
.A2(n_27),
.B1(n_22),
.B2(n_29),
.Y(n_88)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_49),
.Y(n_89)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_49),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_91),
.B(n_52),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_92),
.A2(n_110),
.B1(n_72),
.B2(n_81),
.Y(n_124)
);

NAND2x1_ASAP7_75t_L g97 ( 
.A(n_60),
.B(n_41),
.Y(n_97)
);

A2O1A1Ixp33_ASAP7_75t_SL g120 ( 
.A1(n_97),
.A2(n_72),
.B(n_69),
.C(n_62),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_SL g98 ( 
.A1(n_91),
.A2(n_39),
.B(n_36),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_98),
.B(n_99),
.C(n_36),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_78),
.B(n_39),
.C(n_52),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_83),
.A2(n_42),
.B1(n_30),
.B2(n_22),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_103),
.A2(n_70),
.B1(n_87),
.B2(n_75),
.Y(n_123)
);

O2A1O1Ixp33_ASAP7_75t_L g104 ( 
.A1(n_80),
.A2(n_39),
.B(n_52),
.C(n_29),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_104),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_74),
.A2(n_29),
.B1(n_33),
.B2(n_36),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_112),
.B(n_118),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_78),
.B(n_52),
.Y(n_118)
);

NOR2xp67_ASAP7_75t_L g119 ( 
.A(n_114),
.B(n_71),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_SL g157 ( 
.A(n_119),
.B(n_133),
.Y(n_157)
);

XOR2xp5_ASAP7_75t_SL g169 ( 
.A(n_120),
.B(n_141),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_106),
.Y(n_121)
);

HB1xp67_ASAP7_75t_L g163 ( 
.A(n_121),
.Y(n_163)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_100),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_122),
.B(n_125),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_123),
.A2(n_124),
.B1(n_126),
.B2(n_131),
.Y(n_158)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_100),
.Y(n_125)
);

OAI22xp33_ASAP7_75t_L g126 ( 
.A1(n_117),
.A2(n_68),
.B1(n_61),
.B2(n_59),
.Y(n_126)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_108),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_127),
.B(n_128),
.Y(n_162)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_116),
.Y(n_128)
);

INVx1_ASAP7_75t_SL g130 ( 
.A(n_97),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_130),
.B(n_132),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_117),
.A2(n_85),
.B1(n_71),
.B2(n_33),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_118),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_95),
.B(n_33),
.Y(n_133)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_112),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_134),
.B(n_137),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_96),
.A2(n_36),
.B1(n_65),
.B2(n_4),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_135),
.A2(n_140),
.B1(n_145),
.B2(n_104),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_136),
.B(n_92),
.C(n_107),
.Y(n_159)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_93),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_111),
.B(n_65),
.Y(n_138)
);

INVxp67_ASAP7_75t_L g151 ( 
.A(n_138),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_98),
.B(n_114),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_139),
.B(n_144),
.Y(n_146)
);

NOR4xp25_ASAP7_75t_L g141 ( 
.A(n_97),
.B(n_14),
.C(n_5),
.D(n_6),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_111),
.B(n_14),
.Y(n_142)
);

INVxp67_ASAP7_75t_L g156 ( 
.A(n_142),
.Y(n_156)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_109),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_143),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_114),
.B(n_3),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_L g145 ( 
.A1(n_96),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_126),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_148),
.B(n_149),
.Y(n_191)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_129),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_143),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_150),
.B(n_161),
.Y(n_173)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_129),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_152),
.B(n_164),
.Y(n_172)
);

AOI21xp5_ASAP7_75t_L g153 ( 
.A1(n_139),
.A2(n_99),
.B(n_113),
.Y(n_153)
);

AND2x2_ASAP7_75t_L g189 ( 
.A(n_153),
.B(n_154),
.Y(n_189)
);

AOI21xp5_ASAP7_75t_L g154 ( 
.A1(n_136),
.A2(n_107),
.B(n_105),
.Y(n_154)
);

XOR2xp5_ASAP7_75t_L g177 ( 
.A(n_159),
.B(n_171),
.Y(n_177)
);

INVxp67_ASAP7_75t_L g164 ( 
.A(n_135),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_123),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_165),
.B(n_166),
.Y(n_174)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_124),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_131),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_167),
.B(n_168),
.Y(n_186)
);

AOI21xp5_ASAP7_75t_L g168 ( 
.A1(n_130),
.A2(n_105),
.B(n_109),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_L g171 ( 
.A1(n_144),
.A2(n_95),
.B(n_93),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_SL g175 ( 
.A(n_162),
.B(n_102),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g204 ( 
.A(n_175),
.B(n_176),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_160),
.Y(n_176)
);

XOR2x1_ASAP7_75t_L g178 ( 
.A(n_169),
.B(n_120),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_L g202 ( 
.A1(n_178),
.A2(n_146),
.B(n_154),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_166),
.A2(n_103),
.B1(n_120),
.B2(n_101),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_179),
.A2(n_167),
.B1(n_165),
.B2(n_164),
.Y(n_193)
);

XOR2xp5_ASAP7_75t_L g180 ( 
.A(n_153),
.B(n_120),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_180),
.B(n_158),
.C(n_161),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_147),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_181),
.B(n_187),
.Y(n_196)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_170),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_182),
.B(n_184),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_149),
.B(n_140),
.Y(n_183)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_183),
.Y(n_197)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_147),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_155),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_185),
.B(n_190),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_168),
.Y(n_187)
);

AOI221xp5_ASAP7_75t_L g188 ( 
.A1(n_169),
.A2(n_102),
.B1(n_94),
.B2(n_110),
.C(n_115),
.Y(n_188)
);

AOI322xp5_ASAP7_75t_L g201 ( 
.A1(n_188),
.A2(n_178),
.A3(n_189),
.B1(n_171),
.B2(n_185),
.C1(n_176),
.C2(n_182),
.Y(n_201)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_158),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_152),
.B(n_115),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_192),
.B(n_151),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_193),
.A2(n_209),
.B1(n_174),
.B2(n_172),
.Y(n_218)
);

AOI21xp5_ASAP7_75t_L g194 ( 
.A1(n_187),
.A2(n_151),
.B(n_148),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_L g213 ( 
.A1(n_194),
.A2(n_203),
.B(n_172),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_177),
.B(n_159),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_195),
.B(n_177),
.C(n_189),
.Y(n_214)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_200),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_SL g223 ( 
.A(n_201),
.B(n_202),
.Y(n_223)
);

AOI21xp5_ASAP7_75t_SL g203 ( 
.A1(n_186),
.A2(n_146),
.B(n_157),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_192),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_205),
.B(n_208),
.Y(n_210)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_206),
.B(n_174),
.Y(n_217)
);

NAND3xp33_ASAP7_75t_L g207 ( 
.A(n_183),
.B(n_156),
.C(n_7),
.Y(n_207)
);

NOR3xp33_ASAP7_75t_L g220 ( 
.A(n_207),
.B(n_6),
.C(n_8),
.Y(n_220)
);

OR2x2_ASAP7_75t_L g208 ( 
.A(n_173),
.B(n_156),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_190),
.A2(n_163),
.B1(n_121),
.B2(n_106),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_204),
.B(n_198),
.Y(n_211)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_211),
.Y(n_231)
);

AND2x2_ASAP7_75t_L g212 ( 
.A(n_197),
.B(n_180),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_212),
.B(n_215),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_213),
.A2(n_218),
.B1(n_193),
.B2(n_209),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_214),
.B(n_219),
.C(n_199),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_198),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_217),
.B(n_221),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_195),
.B(n_189),
.C(n_184),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_220),
.B(n_8),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_202),
.B(n_191),
.Y(n_221)
);

AOI21xp5_ASAP7_75t_L g222 ( 
.A1(n_196),
.A2(n_179),
.B(n_9),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_222),
.B(n_8),
.Y(n_232)
);

NOR4xp25_ASAP7_75t_L g224 ( 
.A(n_210),
.B(n_200),
.C(n_199),
.D(n_203),
.Y(n_224)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_224),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g239 ( 
.A(n_225),
.B(n_230),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_219),
.B(n_206),
.C(n_194),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_227),
.B(n_233),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_SL g228 ( 
.A(n_213),
.B(n_208),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_228),
.B(n_229),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_232),
.B(n_11),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_214),
.B(n_10),
.C(n_11),
.Y(n_233)
);

AOI31xp67_ASAP7_75t_SL g235 ( 
.A1(n_231),
.A2(n_226),
.A3(n_216),
.B(n_221),
.Y(n_235)
);

OAI321xp33_ASAP7_75t_L g247 ( 
.A1(n_235),
.A2(n_212),
.A3(n_223),
.B1(n_13),
.B2(n_11),
.C(n_12),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_225),
.B(n_218),
.Y(n_237)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_237),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_238),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_234),
.B(n_217),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_240),
.B(n_227),
.C(n_234),
.Y(n_243)
);

XOR2xp5_ASAP7_75t_L g252 ( 
.A(n_243),
.B(n_240),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_SL g246 ( 
.A(n_242),
.B(n_233),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_246),
.B(n_241),
.Y(n_249)
);

AOI21xp5_ASAP7_75t_L g251 ( 
.A1(n_247),
.A2(n_248),
.B(n_13),
.Y(n_251)
);

OAI21xp5_ASAP7_75t_L g248 ( 
.A1(n_236),
.A2(n_223),
.B(n_12),
.Y(n_248)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_249),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_SL g250 ( 
.A(n_245),
.B(n_239),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_250),
.B(n_251),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_252),
.B(n_243),
.C(n_244),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_254),
.B(n_239),
.Y(n_256)
);

NAND3xp33_ASAP7_75t_L g258 ( 
.A(n_256),
.B(n_257),
.C(n_253),
.Y(n_258)
);

INVxp67_ASAP7_75t_L g257 ( 
.A(n_255),
.Y(n_257)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_258),
.B(n_13),
.Y(n_259)
);


endmodule