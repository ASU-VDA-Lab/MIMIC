module real_jpeg_6303_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_498;
wire n_369;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_366;
wire n_456;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_483;
wire n_367;
wire n_127;
wire n_365;
wire n_356;
wire n_423;
wire n_464;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_422;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_469;
wire n_378;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_338;
wire n_175;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_470;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_21;
wire n_476;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_195;
wire n_110;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_25;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_323;
wire n_166;
wire n_176;
wire n_215;
wire n_286;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_487;
wire n_242;
wire n_493;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_501;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_204;
wire n_158;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_299;
wire n_243;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

INVx8_ASAP7_75t_L g63 ( 
.A(n_0),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_1),
.B(n_128),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_1),
.B(n_183),
.Y(n_182)
);

AND2x2_ASAP7_75t_L g220 ( 
.A(n_1),
.B(n_221),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_SL g249 ( 
.A(n_1),
.B(n_250),
.Y(n_249)
);

AND2x2_ASAP7_75t_SL g298 ( 
.A(n_1),
.B(n_299),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_1),
.B(n_362),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_1),
.B(n_365),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_1),
.B(n_391),
.Y(n_390)
);

AND2x2_ASAP7_75t_SL g24 ( 
.A(n_2),
.B(n_25),
.Y(n_24)
);

INVx1_ASAP7_75t_SL g36 ( 
.A(n_2),
.Y(n_36)
);

AND2x2_ASAP7_75t_L g41 ( 
.A(n_2),
.B(n_42),
.Y(n_41)
);

AND2x2_ASAP7_75t_L g195 ( 
.A(n_2),
.B(n_196),
.Y(n_195)
);

AND2x2_ASAP7_75t_SL g240 ( 
.A(n_2),
.B(n_241),
.Y(n_240)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_3),
.Y(n_504)
);

BUFx3_ASAP7_75t_L g125 ( 
.A(n_4),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g141 ( 
.A(n_4),
.Y(n_141)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_4),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_5),
.B(n_56),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_5),
.B(n_78),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_5),
.B(n_87),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_5),
.B(n_159),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_5),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_5),
.B(n_232),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_5),
.B(n_295),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_5),
.B(n_334),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_6),
.B(n_144),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_6),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g267 ( 
.A(n_6),
.B(n_268),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_6),
.B(n_183),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_6),
.B(n_401),
.Y(n_400)
);

AND2x2_ASAP7_75t_L g153 ( 
.A(n_7),
.B(n_154),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_7),
.B(n_144),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_7),
.B(n_204),
.Y(n_203)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_7),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_7),
.B(n_403),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_7),
.B(n_408),
.Y(n_407)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_8),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g151 ( 
.A(n_9),
.Y(n_151)
);

INVx8_ASAP7_75t_L g162 ( 
.A(n_9),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g241 ( 
.A(n_9),
.Y(n_241)
);

BUFx6f_ASAP7_75t_L g393 ( 
.A(n_9),
.Y(n_393)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

BUFx5_ASAP7_75t_L g42 ( 
.A(n_10),
.Y(n_42)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_10),
.Y(n_80)
);

BUFx5_ASAP7_75t_L g95 ( 
.A(n_10),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g173 ( 
.A(n_10),
.Y(n_173)
);

INVx8_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

INVx3_ASAP7_75t_L g500 ( 
.A(n_12),
.Y(n_500)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_13),
.Y(n_47)
);

BUFx5_ASAP7_75t_L g56 ( 
.A(n_13),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_13),
.Y(n_82)
);

BUFx5_ASAP7_75t_L g154 ( 
.A(n_13),
.Y(n_154)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_13),
.Y(n_180)
);

BUFx6f_ASAP7_75t_L g235 ( 
.A(n_13),
.Y(n_235)
);

BUFx6f_ASAP7_75t_L g327 ( 
.A(n_13),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_14),
.B(n_30),
.Y(n_29)
);

AND2x2_ASAP7_75t_SL g45 ( 
.A(n_14),
.B(n_46),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_14),
.B(n_66),
.Y(n_65)
);

AND2x2_ASAP7_75t_L g89 ( 
.A(n_14),
.B(n_90),
.Y(n_89)
);

AND2x2_ASAP7_75t_L g138 ( 
.A(n_14),
.B(n_139),
.Y(n_138)
);

AND2x2_ASAP7_75t_L g150 ( 
.A(n_14),
.B(n_151),
.Y(n_150)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_14),
.Y(n_188)
);

AND2x2_ASAP7_75t_SL g216 ( 
.A(n_14),
.B(n_217),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_15),
.B(n_118),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_15),
.B(n_132),
.Y(n_131)
);

INVx1_ASAP7_75t_SL g170 ( 
.A(n_15),
.Y(n_170)
);

AND2x2_ASAP7_75t_L g233 ( 
.A(n_15),
.B(n_234),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_15),
.B(n_365),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_15),
.B(n_387),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_SL g413 ( 
.A(n_15),
.B(n_414),
.Y(n_413)
);

BUFx3_ASAP7_75t_L g75 ( 
.A(n_16),
.Y(n_75)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_16),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g428 ( 
.A(n_16),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_17),
.B(n_82),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_17),
.B(n_93),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_17),
.B(n_121),
.Y(n_120)
);

CKINVDCx14_ASAP7_75t_R g165 ( 
.A(n_17),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_17),
.B(n_201),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_17),
.B(n_252),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_17),
.B(n_311),
.Y(n_310)
);

AND2x2_ASAP7_75t_L g350 ( 
.A(n_17),
.B(n_87),
.Y(n_350)
);

AOI21xp5_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_499),
.B(n_501),
.Y(n_18)
);

XNOR2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_106),
.Y(n_19)
);

OAI21xp33_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_68),
.B(n_105),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_21),
.B(n_68),
.Y(n_105)
);

XNOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_48),
.Y(n_21)
);

XNOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_37),
.Y(n_22)
);

MAJIxp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_28),
.C(n_32),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_SL g39 ( 
.A1(n_24),
.A2(n_40),
.B1(n_41),
.B2(n_43),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_24),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_L g52 ( 
.A1(n_24),
.A2(n_32),
.B1(n_43),
.B2(n_53),
.Y(n_52)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_24),
.B(n_230),
.Y(n_229)
);

INVx5_ASAP7_75t_L g67 ( 
.A(n_25),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_26),
.Y(n_87)
);

INVx6_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g205 ( 
.A(n_27),
.Y(n_205)
);

INVx3_ASAP7_75t_L g268 ( 
.A(n_27),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_28),
.A2(n_29),
.B1(n_51),
.B2(n_52),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g331 ( 
.A1(n_28),
.A2(n_29),
.B1(n_332),
.B2(n_338),
.Y(n_331)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

MAJIxp5_ASAP7_75t_L g480 ( 
.A(n_29),
.B(n_333),
.C(n_337),
.Y(n_480)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx3_ASAP7_75t_L g250 ( 
.A(n_31),
.Y(n_250)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_32),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_32),
.A2(n_53),
.B1(n_58),
.B2(n_99),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_32),
.A2(n_53),
.B1(n_147),
.B2(n_148),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_32),
.B(n_149),
.C(n_153),
.Y(n_254)
);

OR2x2_ASAP7_75t_SL g32 ( 
.A(n_33),
.B(n_36),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_35),
.Y(n_91)
);

INVx3_ASAP7_75t_L g135 ( 
.A(n_35),
.Y(n_135)
);

INVx3_ASAP7_75t_L g185 ( 
.A(n_35),
.Y(n_185)
);

BUFx3_ASAP7_75t_L g335 ( 
.A(n_35),
.Y(n_335)
);

OR2x2_ASAP7_75t_L g58 ( 
.A(n_36),
.B(n_59),
.Y(n_58)
);

OR2x2_ASAP7_75t_SL g73 ( 
.A(n_36),
.B(n_74),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_36),
.B(n_326),
.Y(n_325)
);

AOI22xp5_ASAP7_75t_SL g37 ( 
.A1(n_38),
.A2(n_39),
.B1(n_44),
.B2(n_45),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_39),
.Y(n_38)
);

AOI22xp33_ASAP7_75t_L g308 ( 
.A1(n_40),
.A2(n_41),
.B1(n_309),
.B2(n_310),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_SL g349 ( 
.A1(n_40),
.A2(n_41),
.B1(n_350),
.B2(n_351),
.Y(n_349)
);

MAJIxp5_ASAP7_75t_L g467 ( 
.A(n_40),
.B(n_346),
.C(n_351),
.Y(n_467)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_41),
.Y(n_40)
);

MAJIxp5_ASAP7_75t_L g344 ( 
.A(n_41),
.B(n_310),
.C(n_313),
.Y(n_344)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_43),
.B(n_231),
.C(n_233),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_SL g476 ( 
.A1(n_44),
.A2(n_45),
.B1(n_72),
.B2(n_73),
.Y(n_476)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_45),
.Y(n_44)
);

MAJIxp5_ASAP7_75t_L g71 ( 
.A(n_45),
.B(n_58),
.C(n_72),
.Y(n_71)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

MAJIxp5_ASAP7_75t_L g48 ( 
.A(n_49),
.B(n_54),
.C(n_57),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_49),
.A2(n_50),
.B1(n_102),
.B2(n_103),
.Y(n_101)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

CKINVDCx16_ASAP7_75t_R g51 ( 
.A(n_52),
.Y(n_51)
);

MAJIxp5_ASAP7_75t_L g57 ( 
.A(n_53),
.B(n_58),
.C(n_64),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_54),
.A2(n_55),
.B1(n_57),
.B2(n_104),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_55),
.Y(n_54)
);

CKINVDCx16_ASAP7_75t_R g104 ( 
.A(n_57),
.Y(n_104)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_58),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_58),
.A2(n_99),
.B1(n_117),
.B2(n_119),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_58),
.B(n_117),
.C(n_120),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g474 ( 
.A1(n_58),
.A2(n_99),
.B1(n_475),
.B2(n_476),
.Y(n_474)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx4_ASAP7_75t_L g130 ( 
.A(n_61),
.Y(n_130)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx11_ASAP7_75t_L g219 ( 
.A(n_63),
.Y(n_219)
);

BUFx3_ASAP7_75t_L g253 ( 
.A(n_63),
.Y(n_253)
);

BUFx5_ASAP7_75t_L g372 ( 
.A(n_63),
.Y(n_372)
);

INVx3_ASAP7_75t_L g401 ( 
.A(n_63),
.Y(n_401)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_64),
.A2(n_65),
.B1(n_97),
.B2(n_98),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_64),
.A2(n_65),
.B1(n_293),
.B2(n_294),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_64),
.B(n_195),
.C(n_293),
.Y(n_330)
);

INVx1_ASAP7_75t_SL g64 ( 
.A(n_65),
.Y(n_64)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

MAJIxp5_ASAP7_75t_L g68 ( 
.A(n_69),
.B(n_100),
.C(n_101),
.Y(n_68)
);

XOR2xp5_ASAP7_75t_L g495 ( 
.A(n_69),
.B(n_496),
.Y(n_495)
);

MAJIxp5_ASAP7_75t_L g69 ( 
.A(n_70),
.B(n_85),
.C(n_96),
.Y(n_69)
);

XOR2xp5_ASAP7_75t_L g486 ( 
.A(n_70),
.B(n_487),
.Y(n_486)
);

XOR2xp5_ASAP7_75t_L g70 ( 
.A(n_71),
.B(n_76),
.Y(n_70)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_71),
.B(n_81),
.C(n_83),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_72),
.A2(n_73),
.B1(n_131),
.B2(n_264),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g322 ( 
.A1(n_72),
.A2(n_73),
.B1(n_323),
.B2(n_324),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_73),
.Y(n_72)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_73),
.B(n_127),
.C(n_131),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g479 ( 
.A(n_73),
.B(n_195),
.C(n_325),
.Y(n_479)
);

OR2x2_ASAP7_75t_L g187 ( 
.A(n_74),
.B(n_188),
.Y(n_187)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_74),
.Y(n_232)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g403 ( 
.A(n_75),
.Y(n_403)
);

OAI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_77),
.A2(n_81),
.B1(n_83),
.B2(n_84),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_77),
.Y(n_83)
);

INVx6_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVx3_ASAP7_75t_L g144 ( 
.A(n_80),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_81),
.Y(n_84)
);

XNOR2xp5_ASAP7_75t_L g487 ( 
.A(n_85),
.B(n_96),
.Y(n_487)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_86),
.B(n_88),
.C(n_92),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g469 ( 
.A1(n_86),
.A2(n_88),
.B1(n_89),
.B2(n_470),
.Y(n_469)
);

CKINVDCx16_ASAP7_75t_R g470 ( 
.A(n_86),
.Y(n_470)
);

BUFx12f_ASAP7_75t_L g118 ( 
.A(n_87),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_88),
.A2(n_89),
.B1(n_237),
.B2(n_238),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_89),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_89),
.B(n_138),
.C(n_240),
.Y(n_313)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

XOR2xp5_ASAP7_75t_L g468 ( 
.A(n_92),
.B(n_469),
.Y(n_468)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

XNOR2xp5_ASAP7_75t_L g496 ( 
.A(n_100),
.B(n_101),
.Y(n_496)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

OAI21xp5_ASAP7_75t_SL g106 ( 
.A1(n_107),
.A2(n_494),
.B(n_498),
.Y(n_106)
);

AOI21xp5_ASAP7_75t_L g107 ( 
.A1(n_108),
.A2(n_462),
.B(n_491),
.Y(n_107)
);

OR2x2_ASAP7_75t_L g108 ( 
.A(n_109),
.B(n_352),
.Y(n_108)
);

O2A1O1Ixp33_ASAP7_75t_L g109 ( 
.A1(n_110),
.A2(n_282),
.B(n_315),
.C(n_316),
.Y(n_109)
);

AOI21xp5_ASAP7_75t_L g110 ( 
.A1(n_111),
.A2(n_255),
.B(n_281),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_111),
.B(n_460),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_112),
.B(n_223),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_112),
.B(n_223),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_113),
.B(n_174),
.C(n_206),
.Y(n_112)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_113),
.B(n_280),
.Y(n_279)
);

XOR2xp5_ASAP7_75t_L g113 ( 
.A(n_114),
.B(n_145),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_114),
.B(n_146),
.C(n_155),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_115),
.B(n_126),
.C(n_136),
.Y(n_114)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_115),
.B(n_277),
.Y(n_276)
);

XOR2xp5_ASAP7_75t_L g115 ( 
.A(n_116),
.B(n_120),
.Y(n_115)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_117),
.Y(n_119)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

BUFx8_ASAP7_75t_L g362 ( 
.A(n_125),
.Y(n_362)
);

BUFx5_ASAP7_75t_L g420 ( 
.A(n_125),
.Y(n_420)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_126),
.A2(n_136),
.B1(n_137),
.B2(n_278),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_126),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_SL g262 ( 
.A(n_127),
.B(n_263),
.Y(n_262)
);

INVx3_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_129),
.B(n_170),
.Y(n_269)
);

INVx5_ASAP7_75t_SL g129 ( 
.A(n_130),
.Y(n_129)
);

INVxp67_ASAP7_75t_L g264 ( 
.A(n_131),
.Y(n_264)
);

INVx5_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

INVx5_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx4_ASAP7_75t_L g274 ( 
.A(n_135),
.Y(n_274)
);

INVx3_ASAP7_75t_L g312 ( 
.A(n_135),
.Y(n_312)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_142),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_138),
.A2(n_239),
.B1(n_240),
.B2(n_242),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_138),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_138),
.A2(n_142),
.B1(n_143),
.B2(n_242),
.Y(n_275)
);

INVx3_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

INVx3_ASAP7_75t_L g388 ( 
.A(n_141),
.Y(n_388)
);

INVx2_ASAP7_75t_L g411 ( 
.A(n_141),
.Y(n_411)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

XNOR2xp5_ASAP7_75t_L g145 ( 
.A(n_146),
.B(n_155),
.Y(n_145)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_149),
.A2(n_150),
.B1(n_152),
.B2(n_153),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_150),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_150),
.B(n_195),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g366 ( 
.A(n_150),
.B(n_195),
.Y(n_366)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_153),
.Y(n_152)
);

XOR2xp5_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_163),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_L g191 ( 
.A1(n_156),
.A2(n_157),
.B(n_158),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_156),
.B(n_164),
.C(n_169),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_157),
.B(n_158),
.Y(n_156)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_160),
.Y(n_201)
);

INVx4_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g415 ( 
.A(n_162),
.Y(n_415)
);

XNOR2xp5_ASAP7_75t_L g163 ( 
.A(n_164),
.B(n_169),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_165),
.B(n_166),
.Y(n_164)
);

HB1xp67_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

INVx3_ASAP7_75t_L g365 ( 
.A(n_167),
.Y(n_365)
);

BUFx6f_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_171),
.Y(n_169)
);

INVx8_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

BUFx6f_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_174),
.B(n_206),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_175),
.B(n_190),
.C(n_192),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_175),
.A2(n_190),
.B1(n_191),
.B2(n_260),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_175),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g175 ( 
.A(n_176),
.B(n_181),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_176),
.B(n_182),
.C(n_187),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_177),
.B(n_178),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g418 ( 
.A(n_177),
.B(n_419),
.Y(n_418)
);

NOR2xp33_ASAP7_75t_L g426 ( 
.A(n_177),
.B(n_427),
.Y(n_426)
);

INVx5_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

INVx3_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

INVx3_ASAP7_75t_L g299 ( 
.A(n_180),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_182),
.A2(n_186),
.B1(n_187),
.B2(n_189),
.Y(n_181)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_182),
.Y(n_189)
);

INVx4_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

INVx6_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_L g296 ( 
.A1(n_186),
.A2(n_187),
.B1(n_297),
.B2(n_301),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_187),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g347 ( 
.A(n_187),
.B(n_240),
.C(n_298),
.Y(n_347)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_SL g258 ( 
.A(n_192),
.B(n_259),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_193),
.B(n_199),
.C(n_202),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g448 ( 
.A1(n_193),
.A2(n_194),
.B1(n_449),
.B2(n_450),
.Y(n_448)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g289 ( 
.A1(n_195),
.A2(n_290),
.B1(n_291),
.B2(n_292),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_195),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_SL g324 ( 
.A1(n_195),
.A2(n_290),
.B1(n_325),
.B2(n_328),
.Y(n_324)
);

INVx3_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

BUFx3_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

BUFx6f_ASAP7_75t_L g214 ( 
.A(n_198),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g450 ( 
.A1(n_199),
.A2(n_200),
.B1(n_202),
.B2(n_203),
.Y(n_450)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

INVx3_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_205),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g206 ( 
.A(n_207),
.B(n_222),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_209),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_208),
.B(n_209),
.C(n_222),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_SL g209 ( 
.A(n_210),
.B(n_215),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_210),
.B(n_216),
.C(n_220),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_211),
.B(n_212),
.Y(n_210)
);

INVx3_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

INVx4_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_216),
.B(n_220),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g332 ( 
.A1(n_216),
.A2(n_333),
.B1(n_336),
.B2(n_337),
.Y(n_332)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_216),
.Y(n_337)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

INVx6_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

BUFx6f_ASAP7_75t_L g295 ( 
.A(n_219),
.Y(n_295)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_224),
.B(n_225),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_224),
.B(n_226),
.C(n_243),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_243),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_227),
.B(n_236),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_228),
.B(n_229),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_228),
.B(n_229),
.C(n_236),
.Y(n_303)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_231),
.B(n_233),
.Y(n_230)
);

BUFx3_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_L g297 ( 
.A1(n_239),
.A2(n_240),
.B1(n_298),
.B2(n_300),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_SL g394 ( 
.A1(n_239),
.A2(n_240),
.B1(n_360),
.B2(n_361),
.Y(n_394)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_240),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_SL g359 ( 
.A(n_240),
.B(n_360),
.Y(n_359)
);

INVx4_ASAP7_75t_L g424 ( 
.A(n_241),
.Y(n_424)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_244),
.B(n_245),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_244),
.B(n_246),
.C(n_247),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_246),
.B(n_247),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_248),
.B(n_254),
.Y(n_247)
);

XOR2xp5_ASAP7_75t_L g248 ( 
.A(n_249),
.B(n_251),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_249),
.B(n_251),
.C(n_306),
.Y(n_305)
);

INVx3_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

INVxp67_ASAP7_75t_L g306 ( 
.A(n_254),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_256),
.B(n_279),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_SL g460 ( 
.A(n_256),
.B(n_279),
.Y(n_460)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_257),
.B(n_261),
.C(n_276),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g453 ( 
.A1(n_257),
.A2(n_258),
.B1(n_454),
.B2(n_455),
.Y(n_453)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_SL g454 ( 
.A(n_261),
.B(n_276),
.Y(n_454)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_262),
.B(n_265),
.C(n_275),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_SL g443 ( 
.A(n_262),
.B(n_444),
.Y(n_443)
);

XNOR2xp5_ASAP7_75t_L g444 ( 
.A(n_265),
.B(n_275),
.Y(n_444)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_266),
.B(n_269),
.C(n_270),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g378 ( 
.A1(n_266),
.A2(n_267),
.B1(n_270),
.B2(n_379),
.Y(n_378)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

XOR2xp5_ASAP7_75t_L g377 ( 
.A(n_269),
.B(n_378),
.Y(n_377)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_270),
.Y(n_379)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_271),
.B(n_272),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g369 ( 
.A(n_271),
.B(n_370),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_L g421 ( 
.A(n_271),
.B(n_422),
.Y(n_421)
);

INVx3_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

INVx6_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_283),
.B(n_317),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_284),
.B(n_285),
.Y(n_283)
);

OR2x2_ASAP7_75t_L g315 ( 
.A(n_284),
.B(n_285),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_285),
.B(n_318),
.Y(n_317)
);

OR2x2_ASAP7_75t_L g461 ( 
.A(n_285),
.B(n_318),
.Y(n_461)
);

FAx1_ASAP7_75t_L g285 ( 
.A(n_286),
.B(n_302),
.CI(n_314),
.CON(n_285),
.SN(n_285)
);

XNOR2xp5_ASAP7_75t_L g286 ( 
.A(n_287),
.B(n_296),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_288),
.B(n_289),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_288),
.B(n_289),
.C(n_296),
.Y(n_341)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_297),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g300 ( 
.A(n_298),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_SL g302 ( 
.A(n_303),
.B(n_304),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_303),
.B(n_305),
.C(n_307),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_L g304 ( 
.A(n_305),
.B(n_307),
.Y(n_304)
);

XOR2xp5_ASAP7_75t_L g307 ( 
.A(n_308),
.B(n_313),
.Y(n_307)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_310),
.Y(n_309)
);

INVx6_ASAP7_75t_L g311 ( 
.A(n_312),
.Y(n_311)
);

INVxp67_ASAP7_75t_L g316 ( 
.A(n_317),
.Y(n_316)
);

XNOR2xp5_ASAP7_75t_L g318 ( 
.A(n_319),
.B(n_320),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g489 ( 
.A(n_319),
.B(n_321),
.C(n_339),
.Y(n_489)
);

XNOR2xp5_ASAP7_75t_L g320 ( 
.A(n_321),
.B(n_339),
.Y(n_320)
);

XNOR2xp5_ASAP7_75t_L g321 ( 
.A(n_322),
.B(n_329),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g471 ( 
.A(n_322),
.B(n_330),
.C(n_331),
.Y(n_471)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_324),
.Y(n_323)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_325),
.Y(n_328)
);

INVx8_ASAP7_75t_L g326 ( 
.A(n_327),
.Y(n_326)
);

XNOR2xp5_ASAP7_75t_L g329 ( 
.A(n_330),
.B(n_331),
.Y(n_329)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_332),
.Y(n_338)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_333),
.Y(n_336)
);

INVx6_ASAP7_75t_L g334 ( 
.A(n_335),
.Y(n_334)
);

AOI22xp5_ASAP7_75t_L g339 ( 
.A1(n_340),
.A2(n_341),
.B1(n_342),
.B2(n_343),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_L g481 ( 
.A(n_340),
.B(n_344),
.C(n_345),
.Y(n_481)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_341),
.Y(n_340)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_343),
.Y(n_342)
);

XOR2xp5_ASAP7_75t_L g343 ( 
.A(n_344),
.B(n_345),
.Y(n_343)
);

AO22x1_ASAP7_75t_SL g345 ( 
.A1(n_346),
.A2(n_347),
.B1(n_348),
.B2(n_349),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_347),
.Y(n_346)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_349),
.Y(n_348)
);

CKINVDCx20_ASAP7_75t_R g351 ( 
.A(n_350),
.Y(n_351)
);

OAI31xp33_ASAP7_75t_L g352 ( 
.A1(n_353),
.A2(n_458),
.A3(n_459),
.B(n_461),
.Y(n_352)
);

AOI21xp5_ASAP7_75t_L g353 ( 
.A1(n_354),
.A2(n_452),
.B(n_457),
.Y(n_353)
);

OAI21xp5_ASAP7_75t_SL g354 ( 
.A1(n_355),
.A2(n_439),
.B(n_451),
.Y(n_354)
);

AOI21xp5_ASAP7_75t_L g355 ( 
.A1(n_356),
.A2(n_395),
.B(n_438),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_SL g356 ( 
.A(n_357),
.B(n_380),
.Y(n_356)
);

NOR2xp33_ASAP7_75t_L g438 ( 
.A(n_357),
.B(n_380),
.Y(n_438)
);

XNOR2xp5_ASAP7_75t_L g357 ( 
.A(n_358),
.B(n_367),
.Y(n_357)
);

MAJIxp5_ASAP7_75t_L g440 ( 
.A(n_358),
.B(n_368),
.C(n_377),
.Y(n_440)
);

XNOR2xp5_ASAP7_75t_SL g358 ( 
.A(n_359),
.B(n_363),
.Y(n_358)
);

MAJIxp5_ASAP7_75t_L g447 ( 
.A(n_359),
.B(n_364),
.C(n_366),
.Y(n_447)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_361),
.Y(n_360)
);

XNOR2xp5_ASAP7_75t_L g363 ( 
.A(n_364),
.B(n_366),
.Y(n_363)
);

XNOR2xp5_ASAP7_75t_L g367 ( 
.A(n_368),
.B(n_377),
.Y(n_367)
);

MAJIxp5_ASAP7_75t_L g368 ( 
.A(n_369),
.B(n_373),
.C(n_375),
.Y(n_368)
);

XNOR2xp5_ASAP7_75t_SL g381 ( 
.A(n_369),
.B(n_382),
.Y(n_381)
);

INVx2_ASAP7_75t_L g370 ( 
.A(n_371),
.Y(n_370)
);

INVx5_ASAP7_75t_L g371 ( 
.A(n_372),
.Y(n_371)
);

AOI22xp5_ASAP7_75t_L g382 ( 
.A1(n_373),
.A2(n_374),
.B1(n_375),
.B2(n_376),
.Y(n_382)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_374),
.Y(n_373)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_376),
.Y(n_375)
);

MAJIxp5_ASAP7_75t_L g380 ( 
.A(n_381),
.B(n_383),
.C(n_394),
.Y(n_380)
);

XNOR2xp5_ASAP7_75t_L g434 ( 
.A(n_381),
.B(n_435),
.Y(n_434)
);

AOI22xp5_ASAP7_75t_L g435 ( 
.A1(n_383),
.A2(n_384),
.B1(n_394),
.B2(n_436),
.Y(n_435)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_384),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_385),
.B(n_389),
.Y(n_384)
);

AOI22xp5_ASAP7_75t_L g404 ( 
.A1(n_385),
.A2(n_386),
.B1(n_389),
.B2(n_390),
.Y(n_404)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_386),
.Y(n_385)
);

INVx2_ASAP7_75t_L g387 ( 
.A(n_388),
.Y(n_387)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_390),
.Y(n_389)
);

INVx2_ASAP7_75t_L g391 ( 
.A(n_392),
.Y(n_391)
);

INVx2_ASAP7_75t_L g392 ( 
.A(n_393),
.Y(n_392)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_394),
.Y(n_436)
);

OAI21xp5_ASAP7_75t_L g395 ( 
.A1(n_396),
.A2(n_432),
.B(n_437),
.Y(n_395)
);

AOI21xp5_ASAP7_75t_L g396 ( 
.A1(n_397),
.A2(n_416),
.B(n_431),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_SL g397 ( 
.A(n_398),
.B(n_405),
.Y(n_397)
);

NOR2xp33_ASAP7_75t_L g431 ( 
.A(n_398),
.B(n_405),
.Y(n_431)
);

XNOR2xp5_ASAP7_75t_L g398 ( 
.A(n_399),
.B(n_404),
.Y(n_398)
);

XNOR2xp5_ASAP7_75t_L g399 ( 
.A(n_400),
.B(n_402),
.Y(n_399)
);

MAJIxp5_ASAP7_75t_L g433 ( 
.A(n_400),
.B(n_402),
.C(n_404),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_406),
.B(n_412),
.Y(n_405)
);

OAI22xp5_ASAP7_75t_L g429 ( 
.A1(n_406),
.A2(n_407),
.B1(n_412),
.B2(n_413),
.Y(n_429)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_407),
.Y(n_406)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_409),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_410),
.Y(n_409)
);

INVx6_ASAP7_75t_L g410 ( 
.A(n_411),
.Y(n_410)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_413),
.Y(n_412)
);

INVx8_ASAP7_75t_L g414 ( 
.A(n_415),
.Y(n_414)
);

OAI21xp5_ASAP7_75t_L g416 ( 
.A1(n_417),
.A2(n_425),
.B(n_430),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g417 ( 
.A(n_418),
.B(n_421),
.Y(n_417)
);

INVx3_ASAP7_75t_L g419 ( 
.A(n_420),
.Y(n_419)
);

INVx1_ASAP7_75t_SL g422 ( 
.A(n_423),
.Y(n_422)
);

INVx4_ASAP7_75t_L g423 ( 
.A(n_424),
.Y(n_423)
);

NOR2xp33_ASAP7_75t_L g425 ( 
.A(n_426),
.B(n_429),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_426),
.B(n_429),
.Y(n_430)
);

INVx4_ASAP7_75t_L g427 ( 
.A(n_428),
.Y(n_427)
);

NOR2xp33_ASAP7_75t_L g432 ( 
.A(n_433),
.B(n_434),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_433),
.B(n_434),
.Y(n_437)
);

NOR2xp33_ASAP7_75t_L g439 ( 
.A(n_440),
.B(n_441),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_440),
.B(n_441),
.Y(n_451)
);

OAI22xp5_ASAP7_75t_SL g441 ( 
.A1(n_442),
.A2(n_443),
.B1(n_445),
.B2(n_446),
.Y(n_441)
);

MAJIxp5_ASAP7_75t_L g456 ( 
.A(n_442),
.B(n_447),
.C(n_448),
.Y(n_456)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_443),
.Y(n_442)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_446),
.Y(n_445)
);

XOR2xp5_ASAP7_75t_L g446 ( 
.A(n_447),
.B(n_448),
.Y(n_446)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_450),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_SL g452 ( 
.A(n_453),
.B(n_456),
.Y(n_452)
);

NOR2xp33_ASAP7_75t_L g457 ( 
.A(n_453),
.B(n_456),
.Y(n_457)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_454),
.Y(n_455)
);

NOR2xp33_ASAP7_75t_L g462 ( 
.A(n_463),
.B(n_488),
.Y(n_462)
);

OAI21xp33_ASAP7_75t_L g491 ( 
.A1(n_463),
.A2(n_492),
.B(n_493),
.Y(n_491)
);

NOR2xp33_ASAP7_75t_L g463 ( 
.A(n_464),
.B(n_482),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_L g493 ( 
.A(n_464),
.B(n_482),
.Y(n_493)
);

MAJIxp5_ASAP7_75t_L g464 ( 
.A(n_465),
.B(n_472),
.C(n_481),
.Y(n_464)
);

FAx1_ASAP7_75t_SL g490 ( 
.A(n_465),
.B(n_472),
.CI(n_481),
.CON(n_490),
.SN(n_490)
);

XNOR2xp5_ASAP7_75t_SL g465 ( 
.A(n_466),
.B(n_471),
.Y(n_465)
);

XOR2xp5_ASAP7_75t_L g466 ( 
.A(n_467),
.B(n_468),
.Y(n_466)
);

MAJIxp5_ASAP7_75t_L g483 ( 
.A(n_467),
.B(n_468),
.C(n_471),
.Y(n_483)
);

AOI22xp5_ASAP7_75t_L g472 ( 
.A1(n_473),
.A2(n_474),
.B1(n_477),
.B2(n_478),
.Y(n_472)
);

MAJIxp5_ASAP7_75t_L g485 ( 
.A(n_473),
.B(n_479),
.C(n_480),
.Y(n_485)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_474),
.Y(n_473)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_476),
.Y(n_475)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_478),
.Y(n_477)
);

XOR2xp5_ASAP7_75t_L g478 ( 
.A(n_479),
.B(n_480),
.Y(n_478)
);

XOR2xp5_ASAP7_75t_L g482 ( 
.A(n_483),
.B(n_484),
.Y(n_482)
);

MAJIxp5_ASAP7_75t_L g497 ( 
.A(n_483),
.B(n_485),
.C(n_486),
.Y(n_497)
);

XNOR2xp5_ASAP7_75t_L g484 ( 
.A(n_485),
.B(n_486),
.Y(n_484)
);

NOR2xp33_ASAP7_75t_L g488 ( 
.A(n_489),
.B(n_490),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_L g492 ( 
.A(n_489),
.B(n_490),
.Y(n_492)
);

BUFx24_ASAP7_75t_SL g506 ( 
.A(n_490),
.Y(n_506)
);

NOR2xp33_ASAP7_75t_L g494 ( 
.A(n_495),
.B(n_497),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_L g498 ( 
.A(n_495),
.B(n_497),
.Y(n_498)
);

INVx8_ASAP7_75t_L g499 ( 
.A(n_500),
.Y(n_499)
);

INVx13_ASAP7_75t_L g503 ( 
.A(n_500),
.Y(n_503)
);

NOR2xp33_ASAP7_75t_L g501 ( 
.A(n_502),
.B(n_504),
.Y(n_501)
);

BUFx12f_ASAP7_75t_L g502 ( 
.A(n_503),
.Y(n_502)
);


endmodule