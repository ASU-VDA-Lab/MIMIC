module fake_aes_8980_n_1840 (n_117, n_44, n_361, n_185, n_22, n_57, n_26, n_407, n_284, n_278, n_60, n_114, n_41, n_94, n_125, n_9, n_161, n_177, n_130, n_189, n_311, n_19, n_292, n_309, n_160, n_154, n_7, n_29, n_328, n_229, n_336, n_348, n_252, n_152, n_113, n_353, n_206, n_17, n_288, n_383, n_6, n_400, n_296, n_157, n_79, n_202, n_386, n_38, n_142, n_232, n_316, n_31, n_211, n_334, n_389, n_275, n_0, n_131, n_112, n_205, n_330, n_162, n_387, n_163, n_105, n_227, n_384, n_231, n_298, n_411, n_144, n_27, n_53, n_183, n_199, n_351, n_83, n_401, n_28, n_48, n_100, n_305, n_228, n_345, n_360, n_236, n_340, n_150, n_373, n_3, n_18, n_301, n_66, n_222, n_234, n_366, n_286, n_15, n_190, n_246, n_321, n_324, n_392, n_39, n_279, n_303, n_326, n_289, n_333, n_249, n_244, n_50, n_73, n_49, n_119, n_141, n_97, n_167, n_171, n_65, n_196, n_192, n_312, n_137, n_277, n_367, n_45, n_85, n_250, n_314, n_237, n_181, n_101, n_62, n_255, n_36, n_37, n_91, n_108, n_116, n_230, n_209, n_274, n_16, n_282, n_319, n_417, n_241, n_95, n_238, n_318, n_293, n_135, n_42, n_393, n_24, n_247, n_381, n_304, n_399, n_294, n_313, n_210, n_184, n_322, n_310, n_191, n_307, n_46, n_354, n_402, n_32, n_413, n_391, n_235, n_243, n_415, n_394, n_331, n_352, n_268, n_174, n_248, n_72, n_299, n_43, n_89, n_338, n_256, n_67, n_77, n_20, n_404, n_54, n_369, n_172, n_329, n_251, n_59, n_218, n_1, n_271, n_302, n_270, n_362, n_153, n_61, n_259, n_308, n_93, n_412, n_140, n_207, n_224, n_96, n_219, n_133, n_149, n_81, n_69, n_214, n_204, n_88, n_33, n_107, n_403, n_254, n_262, n_10, n_239, n_87, n_379, n_98, n_276, n_320, n_285, n_195, n_165, n_420, n_423, n_342, n_370, n_34, n_5, n_23, n_8, n_217, n_139, n_388, n_193, n_273, n_390, n_120, n_70, n_245, n_90, n_357, n_260, n_78, n_197, n_201, n_317, n_416, n_4, n_374, n_40, n_111, n_64, n_265, n_264, n_200, n_208, n_126, n_178, n_118, n_365, n_179, n_315, n_363, n_409, n_86, n_143, n_295, n_263, n_166, n_186, n_364, n_75, n_376, n_344, n_136, n_283, n_76, n_216, n_147, n_148, n_212, n_92, n_11, n_419, n_396, n_168, n_398, n_134, n_233, n_82, n_106, n_173, n_422, n_327, n_325, n_349, n_51, n_225, n_220, n_358, n_267, n_221, n_203, n_52, n_102, n_115, n_80, n_300, n_158, n_121, n_35, n_339, n_240, n_378, n_359, n_346, n_103, n_180, n_104, n_74, n_335, n_272, n_146, n_397, n_306, n_47, n_215, n_242, n_155, n_13, n_198, n_169, n_424, n_156, n_124, n_297, n_128, n_129, n_410, n_63, n_14, n_71, n_56, n_188, n_377, n_343, n_127, n_291, n_170, n_418, n_380, n_356, n_281, n_341, n_58, n_122, n_187, n_375, n_138, n_371, n_323, n_347, n_258, n_253, n_84, n_266, n_55, n_12, n_213, n_182, n_368, n_355, n_226, n_382, n_159, n_337, n_176, n_68, n_2, n_123, n_223, n_25, n_30, n_372, n_194, n_287, n_110, n_261, n_425, n_332, n_414, n_350, n_164, n_421, n_175, n_145, n_408, n_290, n_405, n_280, n_21, n_99, n_109, n_132, n_395, n_406, n_151, n_385, n_257, n_269, n_1840);
input n_117;
input n_44;
input n_361;
input n_185;
input n_22;
input n_57;
input n_26;
input n_407;
input n_284;
input n_278;
input n_60;
input n_114;
input n_41;
input n_94;
input n_125;
input n_9;
input n_161;
input n_177;
input n_130;
input n_189;
input n_311;
input n_19;
input n_292;
input n_309;
input n_160;
input n_154;
input n_7;
input n_29;
input n_328;
input n_229;
input n_336;
input n_348;
input n_252;
input n_152;
input n_113;
input n_353;
input n_206;
input n_17;
input n_288;
input n_383;
input n_6;
input n_400;
input n_296;
input n_157;
input n_79;
input n_202;
input n_386;
input n_38;
input n_142;
input n_232;
input n_316;
input n_31;
input n_211;
input n_334;
input n_389;
input n_275;
input n_0;
input n_131;
input n_112;
input n_205;
input n_330;
input n_162;
input n_387;
input n_163;
input n_105;
input n_227;
input n_384;
input n_231;
input n_298;
input n_411;
input n_144;
input n_27;
input n_53;
input n_183;
input n_199;
input n_351;
input n_83;
input n_401;
input n_28;
input n_48;
input n_100;
input n_305;
input n_228;
input n_345;
input n_360;
input n_236;
input n_340;
input n_150;
input n_373;
input n_3;
input n_18;
input n_301;
input n_66;
input n_222;
input n_234;
input n_366;
input n_286;
input n_15;
input n_190;
input n_246;
input n_321;
input n_324;
input n_392;
input n_39;
input n_279;
input n_303;
input n_326;
input n_289;
input n_333;
input n_249;
input n_244;
input n_50;
input n_73;
input n_49;
input n_119;
input n_141;
input n_97;
input n_167;
input n_171;
input n_65;
input n_196;
input n_192;
input n_312;
input n_137;
input n_277;
input n_367;
input n_45;
input n_85;
input n_250;
input n_314;
input n_237;
input n_181;
input n_101;
input n_62;
input n_255;
input n_36;
input n_37;
input n_91;
input n_108;
input n_116;
input n_230;
input n_209;
input n_274;
input n_16;
input n_282;
input n_319;
input n_417;
input n_241;
input n_95;
input n_238;
input n_318;
input n_293;
input n_135;
input n_42;
input n_393;
input n_24;
input n_247;
input n_381;
input n_304;
input n_399;
input n_294;
input n_313;
input n_210;
input n_184;
input n_322;
input n_310;
input n_191;
input n_307;
input n_46;
input n_354;
input n_402;
input n_32;
input n_413;
input n_391;
input n_235;
input n_243;
input n_415;
input n_394;
input n_331;
input n_352;
input n_268;
input n_174;
input n_248;
input n_72;
input n_299;
input n_43;
input n_89;
input n_338;
input n_256;
input n_67;
input n_77;
input n_20;
input n_404;
input n_54;
input n_369;
input n_172;
input n_329;
input n_251;
input n_59;
input n_218;
input n_1;
input n_271;
input n_302;
input n_270;
input n_362;
input n_153;
input n_61;
input n_259;
input n_308;
input n_93;
input n_412;
input n_140;
input n_207;
input n_224;
input n_96;
input n_219;
input n_133;
input n_149;
input n_81;
input n_69;
input n_214;
input n_204;
input n_88;
input n_33;
input n_107;
input n_403;
input n_254;
input n_262;
input n_10;
input n_239;
input n_87;
input n_379;
input n_98;
input n_276;
input n_320;
input n_285;
input n_195;
input n_165;
input n_420;
input n_423;
input n_342;
input n_370;
input n_34;
input n_5;
input n_23;
input n_8;
input n_217;
input n_139;
input n_388;
input n_193;
input n_273;
input n_390;
input n_120;
input n_70;
input n_245;
input n_90;
input n_357;
input n_260;
input n_78;
input n_197;
input n_201;
input n_317;
input n_416;
input n_4;
input n_374;
input n_40;
input n_111;
input n_64;
input n_265;
input n_264;
input n_200;
input n_208;
input n_126;
input n_178;
input n_118;
input n_365;
input n_179;
input n_315;
input n_363;
input n_409;
input n_86;
input n_143;
input n_295;
input n_263;
input n_166;
input n_186;
input n_364;
input n_75;
input n_376;
input n_344;
input n_136;
input n_283;
input n_76;
input n_216;
input n_147;
input n_148;
input n_212;
input n_92;
input n_11;
input n_419;
input n_396;
input n_168;
input n_398;
input n_134;
input n_233;
input n_82;
input n_106;
input n_173;
input n_422;
input n_327;
input n_325;
input n_349;
input n_51;
input n_225;
input n_220;
input n_358;
input n_267;
input n_221;
input n_203;
input n_52;
input n_102;
input n_115;
input n_80;
input n_300;
input n_158;
input n_121;
input n_35;
input n_339;
input n_240;
input n_378;
input n_359;
input n_346;
input n_103;
input n_180;
input n_104;
input n_74;
input n_335;
input n_272;
input n_146;
input n_397;
input n_306;
input n_47;
input n_215;
input n_242;
input n_155;
input n_13;
input n_198;
input n_169;
input n_424;
input n_156;
input n_124;
input n_297;
input n_128;
input n_129;
input n_410;
input n_63;
input n_14;
input n_71;
input n_56;
input n_188;
input n_377;
input n_343;
input n_127;
input n_291;
input n_170;
input n_418;
input n_380;
input n_356;
input n_281;
input n_341;
input n_58;
input n_122;
input n_187;
input n_375;
input n_138;
input n_371;
input n_323;
input n_347;
input n_258;
input n_253;
input n_84;
input n_266;
input n_55;
input n_12;
input n_213;
input n_182;
input n_368;
input n_355;
input n_226;
input n_382;
input n_159;
input n_337;
input n_176;
input n_68;
input n_2;
input n_123;
input n_223;
input n_25;
input n_30;
input n_372;
input n_194;
input n_287;
input n_110;
input n_261;
input n_425;
input n_332;
input n_414;
input n_350;
input n_164;
input n_421;
input n_175;
input n_145;
input n_408;
input n_290;
input n_405;
input n_280;
input n_21;
input n_99;
input n_109;
input n_132;
input n_395;
input n_406;
input n_151;
input n_385;
input n_257;
input n_269;
output n_1840;
wire n_1309;
wire n_1497;
wire n_963;
wire n_1034;
wire n_949;
wire n_1277;
wire n_1312;
wire n_858;
wire n_1671;
wire n_646;
wire n_1334;
wire n_1698;
wire n_1627;
wire n_829;
wire n_1603;
wire n_1198;
wire n_1571;
wire n_1382;
wire n_667;
wire n_988;
wire n_1618;
wire n_1477;
wire n_1363;
wire n_1594;
wire n_1812;
wire n_655;
wire n_1298;
wire n_1391;
wire n_903;
wire n_1785;
wire n_965;
wire n_1646;
wire n_918;
wire n_770;
wire n_1211;
wire n_878;
wire n_1667;
wire n_637;
wire n_564;
wire n_779;
wire n_528;
wire n_1128;
wire n_850;
wire n_672;
wire n_627;
wire n_1118;
wire n_1527;
wire n_1161;
wire n_1030;
wire n_807;
wire n_1782;
wire n_877;
wire n_1663;
wire n_1445;
wire n_545;
wire n_896;
wire n_588;
wire n_1743;
wire n_1019;
wire n_1714;
wire n_940;
wire n_1528;
wire n_789;
wire n_1197;
wire n_1163;
wire n_1404;
wire n_452;
wire n_518;
wire n_1336;
wire n_1341;
wire n_1381;
wire n_1760;
wire n_860;
wire n_1208;
wire n_1201;
wire n_1672;
wire n_1342;
wire n_1619;
wire n_1194;
wire n_922;
wire n_465;
wire n_636;
wire n_914;
wire n_1598;
wire n_1352;
wire n_1503;
wire n_1005;
wire n_1097;
wire n_1125;
wire n_1017;
wire n_773;
wire n_847;
wire n_668;
wire n_437;
wire n_680;
wire n_642;
wire n_1267;
wire n_1631;
wire n_830;
wire n_1112;
wire n_517;
wire n_1295;
wire n_1297;
wire n_502;
wire n_543;
wire n_1159;
wire n_1250;
wire n_1002;
wire n_1355;
wire n_915;
wire n_1536;
wire n_1661;
wire n_999;
wire n_769;
wire n_624;
wire n_1597;
wire n_725;
wire n_1407;
wire n_1475;
wire n_1505;
wire n_1018;
wire n_979;
wire n_499;
wire n_1683;
wire n_1349;
wire n_1573;
wire n_1580;
wire n_1605;
wire n_1033;
wire n_1063;
wire n_533;
wire n_1010;
wire n_490;
wire n_648;
wire n_613;
wire n_892;
wire n_1656;
wire n_571;
wire n_1595;
wire n_1604;
wire n_610;
wire n_771;
wire n_1561;
wire n_1337;
wire n_474;
wire n_676;
wire n_950;
wire n_995;
wire n_938;
wire n_746;
wire n_1307;
wire n_619;
wire n_1744;
wire n_501;
wire n_699;
wire n_1654;
wire n_551;
wire n_1061;
wire n_509;
wire n_849;
wire n_1732;
wire n_864;
wire n_1772;
wire n_961;
wire n_1525;
wire n_1718;
wire n_1448;
wire n_1140;
wire n_611;
wire n_990;
wire n_800;
wire n_626;
wire n_1414;
wire n_1500;
wire n_1209;
wire n_1739;
wire n_1399;
wire n_1441;
wire n_926;
wire n_1274;
wire n_1569;
wire n_1775;
wire n_1620;
wire n_537;
wire n_1764;
wire n_660;
wire n_839;
wire n_1210;
wire n_1001;
wire n_1129;
wire n_450;
wire n_1758;
wire n_1406;
wire n_1789;
wire n_1099;
wire n_1328;
wire n_1369;
wire n_1623;
wire n_1831;
wire n_556;
wire n_1214;
wire n_641;
wire n_966;
wire n_527;
wire n_797;
wire n_666;
wire n_1443;
wire n_1313;
wire n_954;
wire n_574;
wire n_1707;
wire n_823;
wire n_706;
wire n_822;
wire n_1181;
wire n_1438;
wire n_1731;
wire n_514;
wire n_1693;
wire n_1690;
wire n_486;
wire n_568;
wire n_716;
wire n_899;
wire n_1547;
wire n_1066;
wire n_1251;
wire n_1199;
wire n_883;
wire n_573;
wire n_1308;
wire n_1790;
wire n_1613;
wire n_673;
wire n_1071;
wire n_1323;
wire n_1703;
wire n_1377;
wire n_1079;
wire n_1582;
wire n_1321;
wire n_1801;
wire n_1838;
wire n_677;
wire n_1354;
wire n_1242;
wire n_756;
wire n_1728;
wire n_1385;
wire n_1711;
wire n_1240;
wire n_1139;
wire n_577;
wire n_1394;
wire n_870;
wire n_1324;
wire n_1716;
wire n_1662;
wire n_790;
wire n_761;
wire n_1660;
wire n_1287;
wire n_472;
wire n_1100;
wire n_1648;
wire n_1193;
wire n_1119;
wire n_825;
wire n_477;
wire n_815;
wire n_1695;
wire n_908;
wire n_429;
wire n_1551;
wire n_488;
wire n_821;
wire n_745;
wire n_684;
wire n_1281;
wire n_1388;
wire n_1102;
wire n_1819;
wire n_723;
wire n_972;
wire n_1522;
wire n_1499;
wire n_1437;
wire n_997;
wire n_1788;
wire n_1387;
wire n_1244;
wire n_1464;
wire n_1184;
wire n_947;
wire n_620;
wire n_1141;
wire n_1740;
wire n_1682;
wire n_1213;
wire n_1452;
wire n_1402;
wire n_1826;
wire n_1189;
wire n_1316;
wire n_923;
wire n_1205;
wire n_1172;
wire n_741;
wire n_1142;
wire n_1447;
wire n_1228;
wire n_1639;
wire n_1730;
wire n_831;
wire n_859;
wire n_1165;
wire n_1300;
wire n_1510;
wire n_1467;
wire n_930;
wire n_994;
wire n_1413;
wire n_774;
wire n_1207;
wire n_1463;
wire n_510;
wire n_1075;
wire n_1615;
wire n_1282;
wire n_493;
wire n_1768;
wire n_855;
wire n_722;
wire n_1590;
wire n_1083;
wire n_690;
wire n_1365;
wire n_1802;
wire n_1164;
wire n_1628;
wire n_1533;
wire n_1611;
wire n_451;
wire n_487;
wire n_748;
wire n_1373;
wire n_1694;
wire n_1563;
wire n_1642;
wire n_824;
wire n_793;
wire n_1792;
wire n_753;
wire n_1753;
wire n_658;
wire n_691;
wire n_444;
wire n_1461;
wire n_1600;
wire n_1226;
wire n_1233;
wire n_1067;
wire n_866;
wire n_1108;
wire n_433;
wire n_1542;
wire n_1311;
wire n_1558;
wire n_483;
wire n_992;
wire n_1748;
wire n_1754;
wire n_1077;
wire n_838;
wire n_705;
wire n_1741;
wire n_964;
wire n_590;
wire n_1229;
wire n_792;
wire n_1412;
wire n_1502;
wire n_925;
wire n_1681;
wire n_1289;
wire n_957;
wire n_808;
wire n_431;
wire n_484;
wire n_852;
wire n_862;
wire n_1602;
wire n_1769;
wire n_1306;
wire n_958;
wire n_468;
wire n_1453;
wire n_917;
wire n_523;
wire n_920;
wire n_1202;
wire n_1361;
wire n_1333;
wire n_1557;
wire n_1733;
wire n_911;
wire n_980;
wire n_1675;
wire n_817;
wire n_1056;
wire n_856;
wire n_1345;
wire n_661;
wire n_1709;
wire n_1606;
wire n_890;
wire n_787;
wire n_1488;
wire n_1015;
wire n_548;
wire n_1048;
wire n_1564;
wire n_1625;
wire n_1521;
wire n_1825;
wire n_973;
wire n_587;
wire n_1818;
wire n_1468;
wire n_476;
wire n_434;
wire n_1725;
wire n_489;
wire n_752;
wire n_1098;
wire n_1012;
wire n_1787;
wire n_461;
wire n_857;
wire n_1090;
wire n_786;
wire n_1121;
wire n_576;
wire n_1179;
wire n_1435;
wire n_1539;
wire n_1629;
wire n_796;
wire n_1216;
wire n_927;
wire n_1405;
wire n_1433;
wire n_1829;
wire n_840;
wire n_846;
wire n_968;
wire n_1543;
wire n_512;
wire n_1834;
wire n_1670;
wire n_1330;
wire n_586;
wire n_1246;
wire n_1276;
wire n_560;
wire n_697;
wire n_780;
wire n_1581;
wire n_447;
wire n_1515;
wire n_897;
wire n_1810;
wire n_1188;
wire n_1496;
wire n_580;
wire n_1009;
wire n_921;
wire n_854;
wire n_1011;
wire n_1807;
wire n_1791;
wire n_1155;
wire n_511;
wire n_467;
wire n_692;
wire n_1415;
wire n_1643;
wire n_1687;
wire n_644;
wire n_1116;
wire n_818;
wire n_738;
wire n_1225;
wire n_575;
wire n_711;
wire n_977;
wire n_884;
wire n_1811;
wire n_767;
wire n_550;
wire n_826;
wire n_1235;
wire n_1171;
wire n_459;
wire n_907;
wire n_1062;
wire n_708;
wire n_1271;
wire n_634;
wire n_1537;
wire n_1520;
wire n_696;
wire n_1608;
wire n_1203;
wire n_1546;
wire n_1524;
wire n_1013;
wire n_1000;
wire n_1370;
wire n_939;
wire n_953;
wire n_478;
wire n_482;
wire n_442;
wire n_485;
wire n_1248;
wire n_1828;
wire n_519;
wire n_1465;
wire n_1777;
wire n_1020;
wire n_1106;
wire n_635;
wire n_731;
wire n_986;
wire n_507;
wire n_605;
wire n_704;
wire n_633;
wire n_873;
wire n_1322;
wire n_751;
wire n_1147;
wire n_466;
wire n_900;
wire n_1540;
wire n_952;
wire n_685;
wire n_565;
wire n_1778;
wire n_1035;
wire n_475;
wire n_578;
wire n_542;
wire n_430;
wire n_1472;
wire n_943;
wire n_1326;
wire n_557;
wire n_1710;
wire n_1781;
wire n_842;
wire n_1269;
wire n_439;
wire n_614;
wire n_1346;
wire n_1107;
wire n_446;
wire n_799;
wire n_1427;
wire n_1765;
wire n_1050;
wire n_1593;
wire n_1763;
wire n_643;
wire n_874;
wire n_1049;
wire n_454;
wire n_687;
wire n_970;
wire n_984;
wire n_1647;
wire n_1621;
wire n_720;
wire n_1157;
wire n_806;
wire n_539;
wire n_1668;
wire n_1692;
wire n_1153;
wire n_1797;
wire n_1657;
wire n_1655;
wire n_1771;
wire n_816;
wire n_522;
wire n_898;
wire n_1562;
wire n_1135;
wire n_669;
wire n_541;
wire n_733;
wire n_894;
wire n_744;
wire n_1514;
wire n_520;
wire n_681;
wire n_1762;
wire n_942;
wire n_1029;
wire n_1665;
wire n_508;
wire n_721;
wire n_1060;
wire n_438;
wire n_640;
wire n_1766;
wire n_1037;
wire n_686;
wire n_944;
wire n_1110;
wire n_498;
wire n_1069;
wire n_1123;
wire n_1817;
wire n_811;
wire n_530;
wire n_737;
wire n_1696;
wire n_1832;
wire n_1266;
wire n_795;
wire n_1232;
wire n_449;
wire n_1796;
wire n_734;
wire n_919;
wire n_763;
wire n_1724;
wire n_1174;
wire n_657;
wire n_583;
wire n_841;
wire n_582;
wire n_1440;
wire n_1541;
wire n_1397;
wire n_1356;
wire n_836;
wire n_1638;
wire n_561;
wire n_1096;
wire n_1553;
wire n_594;
wire n_531;
wire n_1136;
wire n_1752;
wire n_1645;
wire n_1007;
wire n_1117;
wire n_1408;
wire n_1633;
wire n_1784;
wire n_714;
wire n_932;
wire n_837;
wire n_1339;
wire n_1432;
wire n_1315;
wire n_1490;
wire n_867;
wire n_1070;
wire n_1529;
wire n_1270;
wire n_1474;
wire n_1512;
wire n_675;
wire n_504;
wire n_581;
wire n_698;
wire n_555;
wire n_901;
wire n_834;
wire n_727;
wire n_1626;
wire n_1837;
wire n_1038;
wire n_1507;
wire n_1162;
wire n_1103;
wire n_785;
wire n_688;
wire n_1800;
wire n_515;
wire n_1577;
wire n_1719;
wire n_1290;
wire n_1813;
wire n_1234;
wire n_592;
wire n_1045;
wire n_1449;
wire n_1641;
wire n_1798;
wire n_1115;
wire n_521;
wire n_625;
wire n_585;
wire n_1190;
wire n_1237;
wire n_713;
wire n_1705;
wire n_457;
wire n_1799;
wire n_1757;
wire n_736;
wire n_1495;
wire n_1822;
wire n_1583;
wire n_606;
wire n_1729;
wire n_1585;
wire n_1292;
wire n_1425;
wire n_1148;
wire n_1586;
wire n_739;
wire n_1166;
wire n_987;
wire n_1086;
wire n_1697;
wire n_1416;
wire n_1566;
wire n_1236;
wire n_791;
wire n_707;
wire n_1599;
wire n_603;
wire n_1261;
wire n_885;
wire n_500;
wire n_1720;
wire n_607;
wire n_1559;
wire n_1483;
wire n_496;
wire n_1362;
wire n_801;
wire n_1059;
wire n_701;
wire n_1530;
wire n_612;
wire n_1513;
wire n_1679;
wire n_1418;
wire n_1032;
wire n_1284;
wire n_1358;
wire n_1688;
wire n_1767;
wire n_464;
wire n_1243;
wire n_1196;
wire n_1338;
wire n_1634;
wire n_814;
wire n_985;
wire n_1191;
wire n_971;
wire n_904;
wire n_1301;
wire n_532;
wire n_1554;
wire n_1455;
wire n_659;
wire n_432;
wire n_1329;
wire n_1750;
wire n_1572;
wire n_1509;
wire n_1185;
wire n_1511;
wire n_436;
wire n_1653;
wire n_1217;
wire n_715;
wire n_1087;
wire n_662;
wire n_1460;
wire n_1372;
wire n_1640;
wire n_1451;
wire n_617;
wire n_598;
wire n_732;
wire n_724;
wire n_599;
wire n_1459;
wire n_1579;
wire n_609;
wire n_909;
wire n_1273;
wire n_1319;
wire n_596;
wire n_1215;
wire n_951;
wire n_1024;
wire n_1016;
wire n_652;
wire n_1658;
wire n_1417;
wire n_1357;
wire n_638;
wire n_563;
wire n_479;
wire n_623;
wire n_1222;
wire n_593;
wire n_872;
wire n_809;
wire n_1830;
wire n_1101;
wire n_1072;
wire n_1761;
wire n_865;
wire n_1064;
wire n_1380;
wire n_1254;
wire n_1575;
wire n_764;
wire n_426;
wire n_1508;
wire n_1375;
wire n_969;
wire n_1835;
wire n_1253;
wire n_632;
wire n_1182;
wire n_828;
wire n_1138;
wire n_506;
wire n_1458;
wire n_1795;
wire n_1659;
wire n_1816;
wire n_1255;
wire n_1299;
wire n_1450;
wire n_1734;
wire n_1701;
wire n_1480;
wire n_1332;
wire n_427;
wire n_703;
wire n_1272;
wire n_928;
wire n_882;
wire n_1635;
wire n_871;
wire n_803;
wire n_1704;
wire n_1429;
wire n_729;
wire n_805;
wire n_693;
wire n_1036;
wire n_1145;
wire n_651;
wire n_1303;
wire n_1320;
wire n_747;
wire n_1470;
wire n_905;
wire n_525;
wire n_876;
wire n_886;
wire n_959;
wire n_719;
wire n_1206;
wire n_1257;
wire n_710;
wire n_1178;
wire n_1823;
wire n_546;
wire n_664;
wire n_1249;
wire n_1526;
wire n_788;
wire n_1759;
wire n_1774;
wire n_1454;
wire n_1471;
wire n_1383;
wire n_516;
wire n_549;
wire n_1609;
wire n_1576;
wire n_832;
wire n_996;
wire n_1578;
wire n_1794;
wire n_1684;
wire n_1089;
wire n_1717;
wire n_1434;
wire n_1058;
wire n_1396;
wire n_1400;
wire n_1517;
wire n_1610;
wire n_1082;
wire n_1052;
wire n_1055;
wire n_974;
wire n_591;
wire n_933;
wire n_1252;
wire n_1706;
wire n_1473;
wire n_1678;
wire n_536;
wire n_1256;
wire n_1259;
wire n_1674;
wire n_1351;
wire n_1318;
wire n_956;
wire n_1622;
wire n_1755;
wire n_1804;
wire n_1773;
wire n_1614;
wire n_989;
wire n_754;
wire n_775;
wire n_616;
wire n_1227;
wire n_495;
wire n_566;
wire n_1144;
wire n_503;
wire n_1279;
wire n_1152;
wire n_1478;
wire n_1068;
wire n_1565;
wire n_1712;
wire n_1149;
wire n_1430;
wire n_615;
wire n_1386;
wire n_1552;
wire n_1779;
wire n_1170;
wire n_1523;
wire n_1700;
wire n_804;
wire n_570;
wire n_1133;
wire n_1317;
wire n_1492;
wire n_440;
wire n_1550;
wire n_1827;
wire n_679;
wire n_1131;
wire n_597;
wire n_1612;
wire n_1636;
wire n_1039;
wire n_1395;
wire n_835;
wire n_778;
wire n_1156;
wire n_1722;
wire n_1288;
wire n_1340;
wire n_1042;
wire n_1130;
wire n_584;
wire n_912;
wire n_1325;
wire n_1043;
wire n_1283;
wire n_1587;
wire n_1489;
wire n_1726;
wire n_1008;
wire n_1109;
wire n_1026;
wire n_1516;
wire n_1027;
wire n_1040;
wire n_1735;
wire n_1367;
wire n_569;
wire n_946;
wire n_960;
wire n_1689;
wire n_1756;
wire n_1805;
wire n_1592;
wire n_1168;
wire n_1574;
wire n_458;
wire n_1084;
wire n_1824;
wire n_1624;
wire n_618;
wire n_1596;
wire n_470;
wire n_1085;
wire n_1538;
wire n_1073;
wire n_868;
wire n_1466;
wire n_473;
wire n_1699;
wire n_991;
wire n_843;
wire n_1263;
wire n_1393;
wire n_538;
wire n_492;
wire n_1426;
wire n_1555;
wire n_1150;
wire n_1462;
wire n_1327;
wire n_1444;
wire n_650;
wire n_469;
wire n_1187;
wire n_742;
wire n_1713;
wire n_913;
wire n_845;
wire n_1776;
wire n_891;
wire n_1134;
wire n_494;
wire n_631;
wire n_1780;
wire n_934;
wire n_1737;
wire n_562;
wire n_1436;
wire n_1192;
wire n_983;
wire n_781;
wire n_709;
wire n_1105;
wire n_1616;
wire n_1378;
wire n_1570;
wire n_1127;
wire n_1348;
wire n_1173;
wire n_663;
wire n_513;
wire n_1092;
wire n_1124;
wire n_1278;
wire n_998;
wire n_604;
wire n_1260;
wire n_755;
wire n_1409;
wire n_848;
wire n_1031;
wire n_1293;
wire n_1749;
wire n_1280;
wire n_1158;
wire n_1493;
wire n_1544;
wire n_743;
wire n_1786;
wire n_757;
wire n_1568;
wire n_750;
wire n_448;
wire n_645;
wire n_1022;
wire n_802;
wire n_993;
wire n_1122;
wire n_1498;
wire n_1224;
wire n_1806;
wire n_762;
wire n_1422;
wire n_981;
wire n_1095;
wire n_1821;
wire n_758;
wire n_544;
wire n_1175;
wire n_853;
wire n_1376;
wire n_765;
wire n_1177;
wire n_1545;
wire n_1310;
wire n_462;
wire n_1347;
wire n_1384;
wire n_783;
wire n_1074;
wire n_1374;
wire n_463;
wire n_1833;
wire n_1379;
wire n_1003;
wire n_1676;
wire n_678;
wire n_1200;
wire n_1534;
wire n_978;
wire n_547;
wire n_1247;
wire n_628;
wire n_812;
wire n_1501;
wire n_777;
wire n_1504;
wire n_1708;
wire n_481;
wire n_443;
wire n_694;
wire n_1601;
wire n_1262;
wire n_1479;
wire n_1360;
wire n_1486;
wire n_1078;
wire n_702;
wire n_572;
wire n_1094;
wire n_1204;
wire n_1666;
wire n_1169;
wire n_975;
wire n_1721;
wire n_1081;
wire n_1680;
wire n_1644;
wire n_1457;
wire n_671;
wire n_540;
wire n_937;
wire n_1093;
wire n_955;
wire n_1275;
wire n_1669;
wire n_945;
wire n_1518;
wire n_554;
wire n_726;
wire n_1519;
wire n_712;
wire n_608;
wire n_567;
wire n_888;
wire n_1815;
wire n_455;
wire n_529;
wire n_1025;
wire n_1132;
wire n_1389;
wire n_630;
wire n_1673;
wire n_1180;
wire n_647;
wire n_1839;
wire n_1364;
wire n_1350;
wire n_844;
wire n_1742;
wire n_1403;
wire n_1160;
wire n_1420;
wire n_1736;
wire n_1245;
wire n_1195;
wire n_1241;
wire n_1302;
wire n_1589;
wire n_895;
wire n_1481;
wire n_798;
wire n_887;
wire n_471;
wire n_1476;
wire n_1014;
wire n_1410;
wire n_1442;
wire n_665;
wire n_1154;
wire n_1560;
wire n_863;
wire n_1265;
wire n_730;
wire n_1212;
wire n_735;
wire n_1091;
wire n_1630;
wire n_784;
wire n_1491;
wire n_1220;
wire n_893;
wire n_1028;
wire n_910;
wire n_935;
wire n_1046;
wire n_1183;
wire n_460;
wire n_813;
wire n_1485;
wire n_1076;
wire n_1808;
wire n_1186;
wire n_1167;
wire n_674;
wire n_810;
wire n_982;
wire n_1532;
wire n_889;
wire n_689;
wire n_902;
wire n_1423;
wire n_1113;
wire n_1264;
wire n_760;
wire n_941;
wire n_1368;
wire n_931;
wire n_827;
wire n_1218;
wire n_1482;
wire n_1343;
wire n_1793;
wire n_1041;
wire n_1745;
wire n_1080;
wire n_1727;
wire n_1637;
wire n_1126;
wire n_1151;
wire n_936;
wire n_579;
wire n_776;
wire n_879;
wire n_1617;
wire n_1632;
wire n_1738;
wire n_1065;
wire n_1494;
wire n_622;
wire n_601;
wire n_1331;
wire n_1176;
wire n_649;
wire n_526;
wire n_1047;
wire n_768;
wire n_869;
wire n_880;
wire n_621;
wire n_589;
wire n_1809;
wire n_1506;
wire n_1469;
wire n_505;
wire n_1664;
wire n_682;
wire n_1607;
wire n_906;
wire n_1650;
wire n_653;
wire n_881;
wire n_1820;
wire n_1535;
wire n_1439;
wire n_718;
wire n_1484;
wire n_1567;
wire n_1238;
wire n_1411;
wire n_1814;
wire n_1114;
wire n_1304;
wire n_948;
wire n_1286;
wire n_1314;
wire n_717;
wire n_861;
wire n_654;
wire n_1221;
wire n_428;
wire n_794;
wire n_1268;
wire n_639;
wire n_1305;
wire n_552;
wire n_1591;
wire n_1023;
wire n_1057;
wire n_435;
wire n_1702;
wire n_1359;
wire n_1294;
wire n_1051;
wire n_1088;
wire n_851;
wire n_445;
wire n_656;
wire n_1230;
wire n_553;
wire n_1431;
wire n_1685;
wire n_1021;
wire n_1456;
wire n_749;
wire n_535;
wire n_1006;
wire n_1054;
wire n_1353;
wire n_1231;
wire n_456;
wire n_962;
wire n_1424;
wire n_782;
wire n_524;
wire n_1044;
wire n_875;
wire n_497;
wire n_728;
wire n_1239;
wire n_1335;
wire n_924;
wire n_1836;
wire n_441;
wire n_1285;
wire n_1344;
wire n_700;
wire n_534;
wire n_1401;
wire n_1677;
wire n_1296;
wire n_1751;
wire n_1428;
wire n_766;
wire n_602;
wire n_1649;
wire n_1143;
wire n_629;
wire n_1723;
wire n_1549;
wire n_1053;
wire n_1223;
wire n_1421;
wire n_1783;
wire n_1390;
wire n_1691;
wire n_1715;
wire n_967;
wire n_1419;
wire n_1258;
wire n_1487;
wire n_1747;
wire n_1686;
wire n_600;
wire n_1531;
wire n_1548;
wire n_1651;
wire n_1584;
wire n_820;
wire n_558;
wire n_670;
wire n_1004;
wire n_683;
wire n_1371;
wire n_929;
wire n_1111;
wire n_976;
wire n_1446;
wire n_695;
wire n_1104;
wire n_1392;
wire n_1219;
wire n_1120;
wire n_595;
wire n_759;
wire n_1770;
wire n_559;
wire n_1366;
wire n_1588;
wire n_480;
wire n_453;
wire n_833;
wire n_1556;
wire n_1146;
wire n_1652;
wire n_1137;
wire n_916;
wire n_740;
wire n_772;
wire n_819;
wire n_1803;
wire n_1398;
wire n_491;
wire n_1746;
wire n_1291;
INVx1_ASAP7_75t_L g426 ( .A(n_164), .Y(n_426) );
INVx2_ASAP7_75t_L g427 ( .A(n_376), .Y(n_427) );
BUFx2_ASAP7_75t_L g428 ( .A(n_313), .Y(n_428) );
INVx1_ASAP7_75t_L g429 ( .A(n_57), .Y(n_429) );
INVx1_ASAP7_75t_L g430 ( .A(n_265), .Y(n_430) );
INVxp33_ASAP7_75t_SL g431 ( .A(n_7), .Y(n_431) );
INVx1_ASAP7_75t_L g432 ( .A(n_104), .Y(n_432) );
INVx2_ASAP7_75t_L g433 ( .A(n_199), .Y(n_433) );
INVx2_ASAP7_75t_L g434 ( .A(n_73), .Y(n_434) );
CKINVDCx20_ASAP7_75t_R g435 ( .A(n_107), .Y(n_435) );
INVx1_ASAP7_75t_L g436 ( .A(n_251), .Y(n_436) );
CKINVDCx20_ASAP7_75t_R g437 ( .A(n_397), .Y(n_437) );
INVx2_ASAP7_75t_L g438 ( .A(n_270), .Y(n_438) );
INVx1_ASAP7_75t_L g439 ( .A(n_119), .Y(n_439) );
INVx1_ASAP7_75t_L g440 ( .A(n_340), .Y(n_440) );
INVx1_ASAP7_75t_L g441 ( .A(n_210), .Y(n_441) );
INVx1_ASAP7_75t_L g442 ( .A(n_250), .Y(n_442) );
INVxp33_ASAP7_75t_L g443 ( .A(n_399), .Y(n_443) );
INVx1_ASAP7_75t_L g444 ( .A(n_119), .Y(n_444) );
CKINVDCx20_ASAP7_75t_R g445 ( .A(n_335), .Y(n_445) );
CKINVDCx5p33_ASAP7_75t_R g446 ( .A(n_18), .Y(n_446) );
CKINVDCx5p33_ASAP7_75t_R g447 ( .A(n_105), .Y(n_447) );
CKINVDCx5p33_ASAP7_75t_R g448 ( .A(n_204), .Y(n_448) );
INVx1_ASAP7_75t_L g449 ( .A(n_416), .Y(n_449) );
INVx2_ASAP7_75t_L g450 ( .A(n_239), .Y(n_450) );
INVxp33_ASAP7_75t_L g451 ( .A(n_31), .Y(n_451) );
INVx1_ASAP7_75t_L g452 ( .A(n_135), .Y(n_452) );
BUFx10_ASAP7_75t_L g453 ( .A(n_127), .Y(n_453) );
NOR2xp67_ASAP7_75t_L g454 ( .A(n_146), .B(n_184), .Y(n_454) );
CKINVDCx5p33_ASAP7_75t_R g455 ( .A(n_400), .Y(n_455) );
HB1xp67_ASAP7_75t_L g456 ( .A(n_154), .Y(n_456) );
INVx1_ASAP7_75t_L g457 ( .A(n_102), .Y(n_457) );
INVx1_ASAP7_75t_L g458 ( .A(n_417), .Y(n_458) );
INVxp33_ASAP7_75t_L g459 ( .A(n_41), .Y(n_459) );
INVx1_ASAP7_75t_L g460 ( .A(n_218), .Y(n_460) );
INVx1_ASAP7_75t_L g461 ( .A(n_23), .Y(n_461) );
INVx1_ASAP7_75t_L g462 ( .A(n_419), .Y(n_462) );
INVx1_ASAP7_75t_L g463 ( .A(n_55), .Y(n_463) );
INVx1_ASAP7_75t_L g464 ( .A(n_246), .Y(n_464) );
INVxp67_ASAP7_75t_SL g465 ( .A(n_352), .Y(n_465) );
CKINVDCx5p33_ASAP7_75t_R g466 ( .A(n_124), .Y(n_466) );
INVx1_ASAP7_75t_L g467 ( .A(n_120), .Y(n_467) );
INVx1_ASAP7_75t_L g468 ( .A(n_342), .Y(n_468) );
INVx1_ASAP7_75t_L g469 ( .A(n_49), .Y(n_469) );
CKINVDCx5p33_ASAP7_75t_R g470 ( .A(n_235), .Y(n_470) );
INVx1_ASAP7_75t_L g471 ( .A(n_366), .Y(n_471) );
INVx1_ASAP7_75t_L g472 ( .A(n_88), .Y(n_472) );
CKINVDCx5p33_ASAP7_75t_R g473 ( .A(n_163), .Y(n_473) );
INVx1_ASAP7_75t_L g474 ( .A(n_58), .Y(n_474) );
CKINVDCx5p33_ASAP7_75t_R g475 ( .A(n_345), .Y(n_475) );
CKINVDCx5p33_ASAP7_75t_R g476 ( .A(n_54), .Y(n_476) );
INVx1_ASAP7_75t_L g477 ( .A(n_123), .Y(n_477) );
CKINVDCx5p33_ASAP7_75t_R g478 ( .A(n_98), .Y(n_478) );
CKINVDCx20_ASAP7_75t_R g479 ( .A(n_247), .Y(n_479) );
INVx1_ASAP7_75t_L g480 ( .A(n_326), .Y(n_480) );
CKINVDCx5p33_ASAP7_75t_R g481 ( .A(n_414), .Y(n_481) );
INVx1_ASAP7_75t_L g482 ( .A(n_206), .Y(n_482) );
INVx1_ASAP7_75t_SL g483 ( .A(n_401), .Y(n_483) );
CKINVDCx20_ASAP7_75t_R g484 ( .A(n_145), .Y(n_484) );
INVx1_ASAP7_75t_L g485 ( .A(n_163), .Y(n_485) );
INVxp67_ASAP7_75t_SL g486 ( .A(n_290), .Y(n_486) );
INVx1_ASAP7_75t_L g487 ( .A(n_34), .Y(n_487) );
INVx1_ASAP7_75t_SL g488 ( .A(n_226), .Y(n_488) );
INVx1_ASAP7_75t_L g489 ( .A(n_244), .Y(n_489) );
INVx1_ASAP7_75t_L g490 ( .A(n_13), .Y(n_490) );
BUFx3_ASAP7_75t_L g491 ( .A(n_148), .Y(n_491) );
INVx1_ASAP7_75t_L g492 ( .A(n_317), .Y(n_492) );
INVx1_ASAP7_75t_L g493 ( .A(n_208), .Y(n_493) );
INVx1_ASAP7_75t_L g494 ( .A(n_387), .Y(n_494) );
INVx1_ASAP7_75t_L g495 ( .A(n_287), .Y(n_495) );
INVx1_ASAP7_75t_SL g496 ( .A(n_341), .Y(n_496) );
INVx1_ASAP7_75t_L g497 ( .A(n_112), .Y(n_497) );
CKINVDCx5p33_ASAP7_75t_R g498 ( .A(n_172), .Y(n_498) );
INVx1_ASAP7_75t_L g499 ( .A(n_415), .Y(n_499) );
INVx1_ASAP7_75t_L g500 ( .A(n_30), .Y(n_500) );
INVx2_ASAP7_75t_L g501 ( .A(n_47), .Y(n_501) );
INVx2_ASAP7_75t_L g502 ( .A(n_219), .Y(n_502) );
INVx1_ASAP7_75t_L g503 ( .A(n_319), .Y(n_503) );
INVxp67_ASAP7_75t_L g504 ( .A(n_112), .Y(n_504) );
INVx1_ASAP7_75t_L g505 ( .A(n_289), .Y(n_505) );
CKINVDCx20_ASAP7_75t_R g506 ( .A(n_308), .Y(n_506) );
CKINVDCx20_ASAP7_75t_R g507 ( .A(n_252), .Y(n_507) );
INVxp33_ASAP7_75t_L g508 ( .A(n_310), .Y(n_508) );
INVxp67_ASAP7_75t_SL g509 ( .A(n_368), .Y(n_509) );
INVx1_ASAP7_75t_L g510 ( .A(n_198), .Y(n_510) );
CKINVDCx20_ASAP7_75t_R g511 ( .A(n_105), .Y(n_511) );
INVx1_ASAP7_75t_L g512 ( .A(n_46), .Y(n_512) );
INVx1_ASAP7_75t_L g513 ( .A(n_90), .Y(n_513) );
HB1xp67_ASAP7_75t_L g514 ( .A(n_254), .Y(n_514) );
INVx1_ASAP7_75t_L g515 ( .A(n_273), .Y(n_515) );
INVx1_ASAP7_75t_L g516 ( .A(n_279), .Y(n_516) );
CKINVDCx5p33_ASAP7_75t_R g517 ( .A(n_79), .Y(n_517) );
INVx1_ASAP7_75t_L g518 ( .A(n_62), .Y(n_518) );
INVx1_ASAP7_75t_L g519 ( .A(n_348), .Y(n_519) );
INVx1_ASAP7_75t_L g520 ( .A(n_33), .Y(n_520) );
CKINVDCx5p33_ASAP7_75t_R g521 ( .A(n_237), .Y(n_521) );
INVxp67_ASAP7_75t_SL g522 ( .A(n_11), .Y(n_522) );
CKINVDCx5p33_ASAP7_75t_R g523 ( .A(n_190), .Y(n_523) );
INVx1_ASAP7_75t_L g524 ( .A(n_172), .Y(n_524) );
CKINVDCx5p33_ASAP7_75t_R g525 ( .A(n_223), .Y(n_525) );
INVx2_ASAP7_75t_L g526 ( .A(n_302), .Y(n_526) );
INVx1_ASAP7_75t_L g527 ( .A(n_222), .Y(n_527) );
INVxp67_ASAP7_75t_SL g528 ( .A(n_201), .Y(n_528) );
INVx1_ASAP7_75t_L g529 ( .A(n_375), .Y(n_529) );
INVx1_ASAP7_75t_L g530 ( .A(n_363), .Y(n_530) );
BUFx3_ASAP7_75t_L g531 ( .A(n_395), .Y(n_531) );
INVx1_ASAP7_75t_L g532 ( .A(n_10), .Y(n_532) );
INVx1_ASAP7_75t_SL g533 ( .A(n_281), .Y(n_533) );
CKINVDCx5p33_ASAP7_75t_R g534 ( .A(n_39), .Y(n_534) );
INVx1_ASAP7_75t_L g535 ( .A(n_257), .Y(n_535) );
INVx1_ASAP7_75t_SL g536 ( .A(n_132), .Y(n_536) );
INVx2_ASAP7_75t_L g537 ( .A(n_120), .Y(n_537) );
CKINVDCx16_ASAP7_75t_R g538 ( .A(n_286), .Y(n_538) );
INVx1_ASAP7_75t_L g539 ( .A(n_421), .Y(n_539) );
CKINVDCx5p33_ASAP7_75t_R g540 ( .A(n_346), .Y(n_540) );
CKINVDCx5p33_ASAP7_75t_R g541 ( .A(n_374), .Y(n_541) );
CKINVDCx16_ASAP7_75t_R g542 ( .A(n_282), .Y(n_542) );
INVx2_ASAP7_75t_L g543 ( .A(n_8), .Y(n_543) );
INVxp33_ASAP7_75t_L g544 ( .A(n_8), .Y(n_544) );
INVx1_ASAP7_75t_L g545 ( .A(n_338), .Y(n_545) );
BUFx6f_ASAP7_75t_L g546 ( .A(n_267), .Y(n_546) );
INVx1_ASAP7_75t_L g547 ( .A(n_48), .Y(n_547) );
INVx1_ASAP7_75t_L g548 ( .A(n_283), .Y(n_548) );
INVx2_ASAP7_75t_L g549 ( .A(n_135), .Y(n_549) );
INVx2_ASAP7_75t_L g550 ( .A(n_409), .Y(n_550) );
INVx1_ASAP7_75t_L g551 ( .A(n_255), .Y(n_551) );
BUFx6f_ASAP7_75t_L g552 ( .A(n_406), .Y(n_552) );
CKINVDCx5p33_ASAP7_75t_R g553 ( .A(n_336), .Y(n_553) );
INVxp67_ASAP7_75t_SL g554 ( .A(n_284), .Y(n_554) );
INVx1_ASAP7_75t_L g555 ( .A(n_159), .Y(n_555) );
INVx1_ASAP7_75t_L g556 ( .A(n_180), .Y(n_556) );
INVx1_ASAP7_75t_L g557 ( .A(n_134), .Y(n_557) );
INVxp67_ASAP7_75t_L g558 ( .A(n_407), .Y(n_558) );
INVx1_ASAP7_75t_L g559 ( .A(n_422), .Y(n_559) );
NOR2xp67_ASAP7_75t_L g560 ( .A(n_307), .B(n_292), .Y(n_560) );
CKINVDCx20_ASAP7_75t_R g561 ( .A(n_268), .Y(n_561) );
INVx2_ASAP7_75t_L g562 ( .A(n_309), .Y(n_562) );
INVx1_ASAP7_75t_L g563 ( .A(n_382), .Y(n_563) );
CKINVDCx5p33_ASAP7_75t_R g564 ( .A(n_328), .Y(n_564) );
BUFx6f_ASAP7_75t_L g565 ( .A(n_122), .Y(n_565) );
NOR2xp67_ASAP7_75t_L g566 ( .A(n_424), .B(n_107), .Y(n_566) );
INVx1_ASAP7_75t_L g567 ( .A(n_10), .Y(n_567) );
CKINVDCx5p33_ASAP7_75t_R g568 ( .A(n_304), .Y(n_568) );
INVx1_ASAP7_75t_L g569 ( .A(n_79), .Y(n_569) );
INVx1_ASAP7_75t_L g570 ( .A(n_116), .Y(n_570) );
CKINVDCx5p33_ASAP7_75t_R g571 ( .A(n_94), .Y(n_571) );
INVxp67_ASAP7_75t_SL g572 ( .A(n_102), .Y(n_572) );
CKINVDCx5p33_ASAP7_75t_R g573 ( .A(n_325), .Y(n_573) );
INVx1_ASAP7_75t_L g574 ( .A(n_353), .Y(n_574) );
INVx1_ASAP7_75t_L g575 ( .A(n_22), .Y(n_575) );
BUFx10_ASAP7_75t_L g576 ( .A(n_329), .Y(n_576) );
INVxp67_ASAP7_75t_SL g577 ( .A(n_271), .Y(n_577) );
INVx1_ASAP7_75t_L g578 ( .A(n_360), .Y(n_578) );
INVx2_ASAP7_75t_L g579 ( .A(n_331), .Y(n_579) );
CKINVDCx5p33_ASAP7_75t_R g580 ( .A(n_57), .Y(n_580) );
CKINVDCx20_ASAP7_75t_R g581 ( .A(n_211), .Y(n_581) );
INVx1_ASAP7_75t_L g582 ( .A(n_40), .Y(n_582) );
INVxp67_ASAP7_75t_SL g583 ( .A(n_362), .Y(n_583) );
INVx1_ASAP7_75t_L g584 ( .A(n_258), .Y(n_584) );
BUFx3_ASAP7_75t_L g585 ( .A(n_18), .Y(n_585) );
INVx1_ASAP7_75t_L g586 ( .A(n_48), .Y(n_586) );
CKINVDCx5p33_ASAP7_75t_R g587 ( .A(n_4), .Y(n_587) );
CKINVDCx5p33_ASAP7_75t_R g588 ( .A(n_306), .Y(n_588) );
INVx1_ASAP7_75t_L g589 ( .A(n_408), .Y(n_589) );
CKINVDCx20_ASAP7_75t_R g590 ( .A(n_285), .Y(n_590) );
INVx1_ASAP7_75t_L g591 ( .A(n_214), .Y(n_591) );
CKINVDCx20_ASAP7_75t_R g592 ( .A(n_77), .Y(n_592) );
BUFx2_ASAP7_75t_SL g593 ( .A(n_101), .Y(n_593) );
INVx1_ASAP7_75t_L g594 ( .A(n_56), .Y(n_594) );
INVx1_ASAP7_75t_L g595 ( .A(n_148), .Y(n_595) );
INVx1_ASAP7_75t_L g596 ( .A(n_327), .Y(n_596) );
NOR2xp67_ASAP7_75t_L g597 ( .A(n_133), .B(n_248), .Y(n_597) );
INVx1_ASAP7_75t_L g598 ( .A(n_36), .Y(n_598) );
CKINVDCx14_ASAP7_75t_R g599 ( .A(n_243), .Y(n_599) );
INVx1_ASAP7_75t_L g600 ( .A(n_26), .Y(n_600) );
BUFx8_ASAP7_75t_SL g601 ( .A(n_127), .Y(n_601) );
INVx1_ASAP7_75t_L g602 ( .A(n_183), .Y(n_602) );
CKINVDCx20_ASAP7_75t_R g603 ( .A(n_404), .Y(n_603) );
INVx1_ASAP7_75t_L g604 ( .A(n_41), .Y(n_604) );
INVx1_ASAP7_75t_L g605 ( .A(n_98), .Y(n_605) );
CKINVDCx20_ASAP7_75t_R g606 ( .A(n_185), .Y(n_606) );
CKINVDCx5p33_ASAP7_75t_R g607 ( .A(n_358), .Y(n_607) );
INVx1_ASAP7_75t_L g608 ( .A(n_165), .Y(n_608) );
CKINVDCx16_ASAP7_75t_R g609 ( .A(n_405), .Y(n_609) );
INVxp67_ASAP7_75t_L g610 ( .A(n_191), .Y(n_610) );
INVxp33_ASAP7_75t_SL g611 ( .A(n_274), .Y(n_611) );
INVx1_ASAP7_75t_L g612 ( .A(n_212), .Y(n_612) );
INVx1_ASAP7_75t_L g613 ( .A(n_249), .Y(n_613) );
CKINVDCx5p33_ASAP7_75t_R g614 ( .A(n_12), .Y(n_614) );
INVx1_ASAP7_75t_L g615 ( .A(n_398), .Y(n_615) );
INVx1_ASAP7_75t_L g616 ( .A(n_396), .Y(n_616) );
INVx2_ASAP7_75t_L g617 ( .A(n_333), .Y(n_617) );
BUFx3_ASAP7_75t_L g618 ( .A(n_69), .Y(n_618) );
INVx1_ASAP7_75t_L g619 ( .A(n_115), .Y(n_619) );
INVxp33_ASAP7_75t_L g620 ( .A(n_192), .Y(n_620) );
CKINVDCx20_ASAP7_75t_R g621 ( .A(n_425), .Y(n_621) );
INVx1_ASAP7_75t_L g622 ( .A(n_224), .Y(n_622) );
CKINVDCx5p33_ASAP7_75t_R g623 ( .A(n_322), .Y(n_623) );
INVx1_ASAP7_75t_L g624 ( .A(n_121), .Y(n_624) );
CKINVDCx5p33_ASAP7_75t_R g625 ( .A(n_95), .Y(n_625) );
INVx1_ASAP7_75t_L g626 ( .A(n_316), .Y(n_626) );
INVx1_ASAP7_75t_L g627 ( .A(n_225), .Y(n_627) );
NOR2xp67_ASAP7_75t_L g628 ( .A(n_89), .B(n_47), .Y(n_628) );
INVx1_ASAP7_75t_L g629 ( .A(n_85), .Y(n_629) );
INVx1_ASAP7_75t_L g630 ( .A(n_1), .Y(n_630) );
BUFx2_ASAP7_75t_L g631 ( .A(n_221), .Y(n_631) );
INVxp67_ASAP7_75t_SL g632 ( .A(n_402), .Y(n_632) );
INVx1_ASAP7_75t_L g633 ( .A(n_74), .Y(n_633) );
INVx1_ASAP7_75t_L g634 ( .A(n_203), .Y(n_634) );
INVx1_ASAP7_75t_L g635 ( .A(n_385), .Y(n_635) );
INVx1_ASAP7_75t_L g636 ( .A(n_312), .Y(n_636) );
BUFx6f_ASAP7_75t_L g637 ( .A(n_403), .Y(n_637) );
CKINVDCx5p33_ASAP7_75t_R g638 ( .A(n_303), .Y(n_638) );
INVx1_ASAP7_75t_L g639 ( .A(n_217), .Y(n_639) );
INVx1_ASAP7_75t_L g640 ( .A(n_108), .Y(n_640) );
INVx1_ASAP7_75t_L g641 ( .A(n_52), .Y(n_641) );
CKINVDCx5p33_ASAP7_75t_R g642 ( .A(n_118), .Y(n_642) );
INVx1_ASAP7_75t_L g643 ( .A(n_83), .Y(n_643) );
INVx1_ASAP7_75t_L g644 ( .A(n_394), .Y(n_644) );
INVx2_ASAP7_75t_L g645 ( .A(n_171), .Y(n_645) );
INVx1_ASAP7_75t_L g646 ( .A(n_220), .Y(n_646) );
CKINVDCx16_ASAP7_75t_R g647 ( .A(n_314), .Y(n_647) );
INVx2_ASAP7_75t_L g648 ( .A(n_213), .Y(n_648) );
INVx1_ASAP7_75t_L g649 ( .A(n_370), .Y(n_649) );
BUFx6f_ASAP7_75t_L g650 ( .A(n_546), .Y(n_650) );
INVx1_ASAP7_75t_L g651 ( .A(n_434), .Y(n_651) );
OAI22xp5_ASAP7_75t_SL g652 ( .A1(n_435), .A2(n_2), .B1(n_0), .B2(n_1), .Y(n_652) );
INVx3_ASAP7_75t_L g653 ( .A(n_576), .Y(n_653) );
INVx2_ASAP7_75t_L g654 ( .A(n_546), .Y(n_654) );
INVxp33_ASAP7_75t_L g655 ( .A(n_456), .Y(n_655) );
AND2x2_ASAP7_75t_L g656 ( .A(n_451), .B(n_0), .Y(n_656) );
AND2x4_ASAP7_75t_L g657 ( .A(n_491), .B(n_2), .Y(n_657) );
AND2x4_ASAP7_75t_L g658 ( .A(n_491), .B(n_3), .Y(n_658) );
INVx1_ASAP7_75t_L g659 ( .A(n_434), .Y(n_659) );
NAND2xp33_ASAP7_75t_L g660 ( .A(n_443), .B(n_186), .Y(n_660) );
CKINVDCx20_ASAP7_75t_R g661 ( .A(n_435), .Y(n_661) );
INVx1_ASAP7_75t_L g662 ( .A(n_501), .Y(n_662) );
BUFx6f_ASAP7_75t_L g663 ( .A(n_546), .Y(n_663) );
BUFx12f_ASAP7_75t_L g664 ( .A(n_576), .Y(n_664) );
INVx1_ASAP7_75t_L g665 ( .A(n_501), .Y(n_665) );
OAI22xp5_ASAP7_75t_SL g666 ( .A1(n_484), .A2(n_5), .B1(n_3), .B2(n_4), .Y(n_666) );
INVx2_ASAP7_75t_L g667 ( .A(n_546), .Y(n_667) );
INVx2_ASAP7_75t_L g668 ( .A(n_552), .Y(n_668) );
BUFx6f_ASAP7_75t_L g669 ( .A(n_552), .Y(n_669) );
CKINVDCx5p33_ASAP7_75t_R g670 ( .A(n_538), .Y(n_670) );
NOR2xp67_ASAP7_75t_L g671 ( .A(n_514), .B(n_504), .Y(n_671) );
INVx2_ASAP7_75t_L g672 ( .A(n_552), .Y(n_672) );
INVx2_ASAP7_75t_L g673 ( .A(n_552), .Y(n_673) );
INVx1_ASAP7_75t_L g674 ( .A(n_537), .Y(n_674) );
INVx1_ASAP7_75t_L g675 ( .A(n_537), .Y(n_675) );
INVx1_ASAP7_75t_L g676 ( .A(n_543), .Y(n_676) );
INVx1_ASAP7_75t_L g677 ( .A(n_543), .Y(n_677) );
INVx2_ASAP7_75t_L g678 ( .A(n_637), .Y(n_678) );
BUFx6f_ASAP7_75t_L g679 ( .A(n_637), .Y(n_679) );
INVx1_ASAP7_75t_L g680 ( .A(n_549), .Y(n_680) );
INVx6_ASAP7_75t_L g681 ( .A(n_576), .Y(n_681) );
OAI22xp5_ASAP7_75t_L g682 ( .A1(n_451), .A2(n_7), .B1(n_5), .B2(n_6), .Y(n_682) );
AOI22xp5_ASAP7_75t_L g683 ( .A1(n_431), .A2(n_11), .B1(n_6), .B2(n_9), .Y(n_683) );
OA21x2_ASAP7_75t_L g684 ( .A1(n_427), .A2(n_188), .B(n_187), .Y(n_684) );
NAND2xp5_ASAP7_75t_L g685 ( .A(n_428), .B(n_9), .Y(n_685) );
INVx1_ASAP7_75t_L g686 ( .A(n_549), .Y(n_686) );
INVx1_ASAP7_75t_L g687 ( .A(n_645), .Y(n_687) );
NAND2xp5_ASAP7_75t_L g688 ( .A(n_631), .B(n_12), .Y(n_688) );
INVx2_ASAP7_75t_L g689 ( .A(n_637), .Y(n_689) );
BUFx6f_ASAP7_75t_L g690 ( .A(n_637), .Y(n_690) );
INVx1_ASAP7_75t_L g691 ( .A(n_645), .Y(n_691) );
INVx1_ASAP7_75t_L g692 ( .A(n_657), .Y(n_692) );
INVx1_ASAP7_75t_L g693 ( .A(n_657), .Y(n_693) );
INVx1_ASAP7_75t_L g694 ( .A(n_657), .Y(n_694) );
NAND2x1p5_ASAP7_75t_L g695 ( .A(n_657), .B(n_585), .Y(n_695) );
AO22x1_ASAP7_75t_L g696 ( .A1(n_658), .A2(n_508), .B1(n_620), .B2(n_443), .Y(n_696) );
INVx2_ASAP7_75t_L g697 ( .A(n_650), .Y(n_697) );
AND2x6_ASAP7_75t_L g698 ( .A(n_658), .B(n_531), .Y(n_698) );
INVxp33_ASAP7_75t_L g699 ( .A(n_655), .Y(n_699) );
AND2x6_ASAP7_75t_L g700 ( .A(n_658), .B(n_531), .Y(n_700) );
AOI22xp33_ASAP7_75t_L g701 ( .A1(n_658), .A2(n_429), .B1(n_432), .B2(n_426), .Y(n_701) );
INVx1_ASAP7_75t_L g702 ( .A(n_654), .Y(n_702) );
NAND2xp5_ASAP7_75t_SL g703 ( .A(n_653), .B(n_542), .Y(n_703) );
AND2x4_ASAP7_75t_L g704 ( .A(n_653), .B(n_585), .Y(n_704) );
BUFx6f_ASAP7_75t_L g705 ( .A(n_650), .Y(n_705) );
INVx2_ASAP7_75t_L g706 ( .A(n_650), .Y(n_706) );
INVx2_ASAP7_75t_L g707 ( .A(n_650), .Y(n_707) );
NOR2xp33_ASAP7_75t_L g708 ( .A(n_681), .B(n_508), .Y(n_708) );
NAND2xp5_ASAP7_75t_L g709 ( .A(n_653), .B(n_620), .Y(n_709) );
INVx1_ASAP7_75t_L g710 ( .A(n_654), .Y(n_710) );
NAND2xp33_ASAP7_75t_L g711 ( .A(n_653), .B(n_475), .Y(n_711) );
INVx1_ASAP7_75t_L g712 ( .A(n_654), .Y(n_712) );
INVx2_ASAP7_75t_L g713 ( .A(n_650), .Y(n_713) );
AND2x2_ASAP7_75t_L g714 ( .A(n_656), .B(n_459), .Y(n_714) );
AND2x2_ASAP7_75t_SL g715 ( .A(n_660), .B(n_609), .Y(n_715) );
AND2x2_ASAP7_75t_L g716 ( .A(n_656), .B(n_459), .Y(n_716) );
INVx4_ASAP7_75t_L g717 ( .A(n_684), .Y(n_717) );
BUFx10_ASAP7_75t_L g718 ( .A(n_681), .Y(n_718) );
CKINVDCx8_ASAP7_75t_R g719 ( .A(n_670), .Y(n_719) );
INVx5_ASAP7_75t_L g720 ( .A(n_650), .Y(n_720) );
CKINVDCx5p33_ASAP7_75t_R g721 ( .A(n_664), .Y(n_721) );
INVx1_ASAP7_75t_SL g722 ( .A(n_681), .Y(n_722) );
AND2x6_ASAP7_75t_L g723 ( .A(n_685), .B(n_430), .Y(n_723) );
INVx2_ASAP7_75t_L g724 ( .A(n_663), .Y(n_724) );
INVx3_ASAP7_75t_L g725 ( .A(n_663), .Y(n_725) );
AND2x2_ASAP7_75t_L g726 ( .A(n_681), .B(n_544), .Y(n_726) );
INVx1_ASAP7_75t_L g727 ( .A(n_667), .Y(n_727) );
AND2x4_ASAP7_75t_L g728 ( .A(n_671), .B(n_618), .Y(n_728) );
NAND2x1p5_ASAP7_75t_L g729 ( .A(n_684), .B(n_618), .Y(n_729) );
INVx1_ASAP7_75t_L g730 ( .A(n_667), .Y(n_730) );
NOR2x1p5_ASAP7_75t_L g731 ( .A(n_664), .B(n_446), .Y(n_731) );
NAND2xp5_ASAP7_75t_SL g732 ( .A(n_692), .B(n_647), .Y(n_732) );
NAND2xp5_ASAP7_75t_L g733 ( .A(n_709), .B(n_681), .Y(n_733) );
NAND2xp5_ASAP7_75t_L g734 ( .A(n_709), .B(n_664), .Y(n_734) );
INVx2_ASAP7_75t_L g735 ( .A(n_702), .Y(n_735) );
INVx1_ASAP7_75t_L g736 ( .A(n_704), .Y(n_736) );
AND2x4_ASAP7_75t_L g737 ( .A(n_731), .B(n_671), .Y(n_737) );
INVx5_ASAP7_75t_L g738 ( .A(n_698), .Y(n_738) );
AOI22xp5_ASAP7_75t_L g739 ( .A1(n_696), .A2(n_685), .B1(n_688), .B2(n_682), .Y(n_739) );
NAND2xp5_ASAP7_75t_SL g740 ( .A(n_692), .B(n_688), .Y(n_740) );
AND2x2_ASAP7_75t_L g741 ( .A(n_699), .B(n_544), .Y(n_741) );
BUFx3_ASAP7_75t_L g742 ( .A(n_698), .Y(n_742) );
NAND2xp5_ASAP7_75t_L g743 ( .A(n_726), .B(n_448), .Y(n_743) );
NAND2xp5_ASAP7_75t_L g744 ( .A(n_726), .B(n_448), .Y(n_744) );
INVx2_ASAP7_75t_L g745 ( .A(n_710), .Y(n_745) );
CKINVDCx5p33_ASAP7_75t_R g746 ( .A(n_721), .Y(n_746) );
AND3x2_ASAP7_75t_SL g747 ( .A(n_696), .B(n_661), .C(n_652), .Y(n_747) );
AND3x1_ASAP7_75t_L g748 ( .A(n_714), .B(n_683), .C(n_666), .Y(n_748) );
NOR2x1_ASAP7_75t_L g749 ( .A(n_731), .B(n_703), .Y(n_749) );
INVx1_ASAP7_75t_L g750 ( .A(n_704), .Y(n_750) );
INVx2_ASAP7_75t_L g751 ( .A(n_695), .Y(n_751) );
AOI22xp33_ASAP7_75t_L g752 ( .A1(n_698), .A2(n_682), .B1(n_431), .B2(n_659), .Y(n_752) );
INVx1_ASAP7_75t_L g753 ( .A(n_695), .Y(n_753) );
INVx1_ASAP7_75t_L g754 ( .A(n_695), .Y(n_754) );
NAND2xp5_ASAP7_75t_L g755 ( .A(n_708), .B(n_455), .Y(n_755) );
INVx4_ASAP7_75t_L g756 ( .A(n_718), .Y(n_756) );
NOR2x2_ASAP7_75t_L g757 ( .A(n_719), .B(n_601), .Y(n_757) );
NAND2xp5_ASAP7_75t_L g758 ( .A(n_714), .B(n_455), .Y(n_758) );
INVx2_ASAP7_75t_L g759 ( .A(n_693), .Y(n_759) );
CKINVDCx5p33_ASAP7_75t_R g760 ( .A(n_719), .Y(n_760) );
NAND2xp5_ASAP7_75t_L g761 ( .A(n_716), .B(n_470), .Y(n_761) );
CKINVDCx5p33_ASAP7_75t_R g762 ( .A(n_719), .Y(n_762) );
BUFx6f_ASAP7_75t_L g763 ( .A(n_698), .Y(n_763) );
OAI22xp33_ASAP7_75t_L g764 ( .A1(n_693), .A2(n_683), .B1(n_437), .B2(n_479), .Y(n_764) );
INVx1_ASAP7_75t_L g765 ( .A(n_728), .Y(n_765) );
INVx4_ASAP7_75t_L g766 ( .A(n_718), .Y(n_766) );
NAND2xp5_ASAP7_75t_L g767 ( .A(n_716), .B(n_470), .Y(n_767) );
NAND2xp5_ASAP7_75t_SL g768 ( .A(n_694), .B(n_436), .Y(n_768) );
NAND2xp5_ASAP7_75t_L g769 ( .A(n_722), .B(n_553), .Y(n_769) );
NOR2x1_ASAP7_75t_L g770 ( .A(n_728), .B(n_437), .Y(n_770) );
NAND2x1p5_ASAP7_75t_L g771 ( .A(n_722), .B(n_439), .Y(n_771) );
AOI22xp33_ASAP7_75t_L g772 ( .A1(n_698), .A2(n_659), .B1(n_662), .B2(n_651), .Y(n_772) );
INVx2_ASAP7_75t_L g773 ( .A(n_710), .Y(n_773) );
OR2x6_ASAP7_75t_L g774 ( .A(n_728), .B(n_652), .Y(n_774) );
AOI22xp5_ASAP7_75t_L g775 ( .A1(n_715), .A2(n_445), .B1(n_506), .B2(n_479), .Y(n_775) );
BUFx3_ASAP7_75t_L g776 ( .A(n_698), .Y(n_776) );
NAND2xp5_ASAP7_75t_L g777 ( .A(n_723), .B(n_553), .Y(n_777) );
NAND2xp5_ASAP7_75t_L g778 ( .A(n_723), .B(n_564), .Y(n_778) );
AND2x4_ASAP7_75t_L g779 ( .A(n_728), .B(n_445), .Y(n_779) );
HB1xp67_ASAP7_75t_L g780 ( .A(n_698), .Y(n_780) );
INVx2_ASAP7_75t_L g781 ( .A(n_712), .Y(n_781) );
NAND2xp5_ASAP7_75t_L g782 ( .A(n_723), .B(n_564), .Y(n_782) );
INVxp67_ASAP7_75t_L g783 ( .A(n_723), .Y(n_783) );
CKINVDCx5p33_ASAP7_75t_R g784 ( .A(n_715), .Y(n_784) );
NAND2xp5_ASAP7_75t_L g785 ( .A(n_723), .B(n_568), .Y(n_785) );
INVx3_ASAP7_75t_L g786 ( .A(n_718), .Y(n_786) );
HB1xp67_ASAP7_75t_L g787 ( .A(n_698), .Y(n_787) );
AOI22xp5_ASAP7_75t_L g788 ( .A1(n_715), .A2(n_507), .B1(n_561), .B2(n_506), .Y(n_788) );
NAND2xp5_ASAP7_75t_L g789 ( .A(n_723), .B(n_568), .Y(n_789) );
INVx1_ASAP7_75t_SL g790 ( .A(n_723), .Y(n_790) );
AOI22xp5_ASAP7_75t_L g791 ( .A1(n_723), .A2(n_561), .B1(n_581), .B2(n_507), .Y(n_791) );
NAND2xp5_ASAP7_75t_SL g792 ( .A(n_694), .B(n_440), .Y(n_792) );
NAND2xp5_ASAP7_75t_SL g793 ( .A(n_701), .B(n_441), .Y(n_793) );
HB1xp67_ASAP7_75t_L g794 ( .A(n_700), .Y(n_794) );
OR2x6_ASAP7_75t_L g795 ( .A(n_729), .B(n_666), .Y(n_795) );
NAND2xp5_ASAP7_75t_SL g796 ( .A(n_701), .B(n_442), .Y(n_796) );
NOR2x1_ASAP7_75t_L g797 ( .A(n_711), .B(n_581), .Y(n_797) );
NAND2xp5_ASAP7_75t_L g798 ( .A(n_700), .B(n_573), .Y(n_798) );
CKINVDCx20_ASAP7_75t_R g799 ( .A(n_718), .Y(n_799) );
AOI22xp33_ASAP7_75t_L g800 ( .A1(n_700), .A2(n_662), .B1(n_665), .B2(n_651), .Y(n_800) );
INVx3_ASAP7_75t_L g801 ( .A(n_700), .Y(n_801) );
AOI21xp5_ASAP7_75t_L g802 ( .A1(n_717), .A2(n_684), .B(n_433), .Y(n_802) );
AND2x4_ASAP7_75t_L g803 ( .A(n_700), .B(n_590), .Y(n_803) );
AOI22xp5_ASAP7_75t_L g804 ( .A1(n_700), .A2(n_603), .B1(n_606), .B2(n_590), .Y(n_804) );
BUFx6f_ASAP7_75t_L g805 ( .A(n_700), .Y(n_805) );
INVx1_ASAP7_75t_L g806 ( .A(n_700), .Y(n_806) );
NOR2x1p5_ASAP7_75t_L g807 ( .A(n_717), .B(n_446), .Y(n_807) );
HB1xp67_ASAP7_75t_L g808 ( .A(n_729), .Y(n_808) );
NAND2xp5_ASAP7_75t_L g809 ( .A(n_717), .B(n_588), .Y(n_809) );
INVx1_ASAP7_75t_L g810 ( .A(n_712), .Y(n_810) );
OR2x6_ASAP7_75t_L g811 ( .A(n_803), .B(n_593), .Y(n_811) );
A2O1A1Ixp33_ASAP7_75t_L g812 ( .A1(n_759), .A2(n_452), .B(n_457), .C(n_444), .Y(n_812) );
INVx4_ASAP7_75t_SL g813 ( .A(n_763), .Y(n_813) );
AND2x4_ASAP7_75t_L g814 ( .A(n_749), .B(n_522), .Y(n_814) );
AND2x2_ASAP7_75t_L g815 ( .A(n_741), .B(n_484), .Y(n_815) );
NAND2xp5_ASAP7_75t_L g816 ( .A(n_739), .B(n_729), .Y(n_816) );
CKINVDCx20_ASAP7_75t_R g817 ( .A(n_746), .Y(n_817) );
INVx2_ASAP7_75t_L g818 ( .A(n_736), .Y(n_818) );
NOR2xp33_ASAP7_75t_L g819 ( .A(n_734), .B(n_601), .Y(n_819) );
NAND2xp5_ASAP7_75t_L g820 ( .A(n_740), .B(n_447), .Y(n_820) );
BUFx6f_ASAP7_75t_L g821 ( .A(n_763), .Y(n_821) );
O2A1O1Ixp33_ASAP7_75t_L g822 ( .A1(n_793), .A2(n_674), .B(n_675), .C(n_665), .Y(n_822) );
BUFx2_ASAP7_75t_L g823 ( .A(n_799), .Y(n_823) );
BUFx12f_ASAP7_75t_L g824 ( .A(n_760), .Y(n_824) );
BUFx6f_ASAP7_75t_L g825 ( .A(n_763), .Y(n_825) );
BUFx6f_ASAP7_75t_L g826 ( .A(n_763), .Y(n_826) );
AND2x2_ASAP7_75t_L g827 ( .A(n_779), .B(n_511), .Y(n_827) );
HB1xp67_ASAP7_75t_L g828 ( .A(n_771), .Y(n_828) );
INVx3_ASAP7_75t_L g829 ( .A(n_756), .Y(n_829) );
AND2x4_ASAP7_75t_L g830 ( .A(n_765), .B(n_572), .Y(n_830) );
INVx3_ASAP7_75t_L g831 ( .A(n_756), .Y(n_831) );
CKINVDCx8_ASAP7_75t_R g832 ( .A(n_762), .Y(n_832) );
BUFx3_ASAP7_75t_L g833 ( .A(n_753), .Y(n_833) );
OR2x2_ASAP7_75t_L g834 ( .A(n_764), .B(n_447), .Y(n_834) );
AOI21xp5_ASAP7_75t_L g835 ( .A1(n_802), .A2(n_684), .B(n_727), .Y(n_835) );
BUFx6f_ASAP7_75t_L g836 ( .A(n_805), .Y(n_836) );
INVx1_ASAP7_75t_L g837 ( .A(n_750), .Y(n_837) );
INVxp67_ASAP7_75t_L g838 ( .A(n_758), .Y(n_838) );
INVx2_ASAP7_75t_L g839 ( .A(n_735), .Y(n_839) );
HB1xp67_ASAP7_75t_L g840 ( .A(n_771), .Y(n_840) );
CKINVDCx20_ASAP7_75t_R g841 ( .A(n_804), .Y(n_841) );
NAND2xp5_ASAP7_75t_SL g842 ( .A(n_766), .B(n_588), .Y(n_842) );
INVxp67_ASAP7_75t_L g843 ( .A(n_761), .Y(n_843) );
BUFx6f_ASAP7_75t_L g844 ( .A(n_805), .Y(n_844) );
O2A1O1Ixp5_ASAP7_75t_L g845 ( .A1(n_793), .A2(n_486), .B(n_509), .C(n_465), .Y(n_845) );
BUFx3_ASAP7_75t_L g846 ( .A(n_754), .Y(n_846) );
NAND2xp5_ASAP7_75t_SL g847 ( .A(n_766), .B(n_607), .Y(n_847) );
INVx2_ASAP7_75t_SL g848 ( .A(n_803), .Y(n_848) );
A2O1A1Ixp33_ASAP7_75t_L g849 ( .A1(n_752), .A2(n_463), .B(n_467), .C(n_461), .Y(n_849) );
OR2x2_ASAP7_75t_L g850 ( .A(n_764), .B(n_466), .Y(n_850) );
BUFx3_ASAP7_75t_L g851 ( .A(n_779), .Y(n_851) );
AOI21xp5_ASAP7_75t_L g852 ( .A1(n_809), .A2(n_730), .B(n_554), .Y(n_852) );
INVx1_ASAP7_75t_L g853 ( .A(n_751), .Y(n_853) );
INVx2_ASAP7_75t_L g854 ( .A(n_735), .Y(n_854) );
NAND2xp5_ASAP7_75t_L g855 ( .A(n_740), .B(n_466), .Y(n_855) );
INVx1_ASAP7_75t_L g856 ( .A(n_810), .Y(n_856) );
OR2x2_ASAP7_75t_L g857 ( .A(n_775), .B(n_498), .Y(n_857) );
AOI21xp5_ASAP7_75t_L g858 ( .A1(n_768), .A2(n_730), .B(n_577), .Y(n_858) );
AND2x2_ASAP7_75t_L g859 ( .A(n_791), .B(n_511), .Y(n_859) );
BUFx2_ASAP7_75t_L g860 ( .A(n_757), .Y(n_860) );
INVx1_ASAP7_75t_L g861 ( .A(n_767), .Y(n_861) );
AOI222xp33_ASAP7_75t_L g862 ( .A1(n_784), .A2(n_592), .B1(n_580), .B2(n_517), .C1(n_587), .C2(n_571), .Y(n_862) );
CKINVDCx5p33_ASAP7_75t_R g863 ( .A(n_788), .Y(n_863) );
O2A1O1Ixp33_ASAP7_75t_L g864 ( .A1(n_796), .A2(n_675), .B(n_676), .C(n_674), .Y(n_864) );
INVxp67_ASAP7_75t_L g865 ( .A(n_743), .Y(n_865) );
INVx2_ASAP7_75t_SL g866 ( .A(n_807), .Y(n_866) );
HB1xp67_ASAP7_75t_L g867 ( .A(n_805), .Y(n_867) );
BUFx6f_ASAP7_75t_L g868 ( .A(n_805), .Y(n_868) );
AND2x4_ASAP7_75t_L g869 ( .A(n_738), .B(n_454), .Y(n_869) );
INVx2_ASAP7_75t_L g870 ( .A(n_745), .Y(n_870) );
INVx1_ASAP7_75t_L g871 ( .A(n_733), .Y(n_871) );
INVx2_ASAP7_75t_L g872 ( .A(n_745), .Y(n_872) );
NAND2xp5_ASAP7_75t_L g873 ( .A(n_752), .B(n_498), .Y(n_873) );
BUFx6f_ASAP7_75t_L g874 ( .A(n_742), .Y(n_874) );
CKINVDCx20_ASAP7_75t_R g875 ( .A(n_795), .Y(n_875) );
BUFx12f_ASAP7_75t_L g876 ( .A(n_774), .Y(n_876) );
AOI22xp5_ASAP7_75t_L g877 ( .A1(n_770), .A2(n_606), .B1(n_621), .B2(n_603), .Y(n_877) );
INVx2_ASAP7_75t_L g878 ( .A(n_773), .Y(n_878) );
AOI21xp5_ASAP7_75t_L g879 ( .A1(n_768), .A2(n_583), .B(n_528), .Y(n_879) );
INVx1_ASAP7_75t_L g880 ( .A(n_773), .Y(n_880) );
INVx2_ASAP7_75t_L g881 ( .A(n_781), .Y(n_881) );
NAND2xp5_ASAP7_75t_L g882 ( .A(n_772), .B(n_517), .Y(n_882) );
INVx1_ASAP7_75t_L g883 ( .A(n_781), .Y(n_883) );
NOR2xp33_ASAP7_75t_L g884 ( .A(n_732), .B(n_611), .Y(n_884) );
AOI22xp33_ASAP7_75t_L g885 ( .A1(n_795), .A2(n_611), .B1(n_599), .B2(n_592), .Y(n_885) );
A2O1A1Ixp33_ASAP7_75t_L g886 ( .A1(n_792), .A2(n_472), .B(n_474), .C(n_469), .Y(n_886) );
BUFx3_ASAP7_75t_L g887 ( .A(n_737), .Y(n_887) );
NOR2x1_ASAP7_75t_L g888 ( .A(n_797), .B(n_621), .Y(n_888) );
NOR2xp33_ASAP7_75t_L g889 ( .A(n_732), .B(n_571), .Y(n_889) );
INVx1_ASAP7_75t_SL g890 ( .A(n_738), .Y(n_890) );
INVx1_ASAP7_75t_L g891 ( .A(n_744), .Y(n_891) );
BUFx6f_ASAP7_75t_L g892 ( .A(n_742), .Y(n_892) );
A2O1A1Ixp33_ASAP7_75t_L g893 ( .A1(n_792), .A2(n_485), .B(n_487), .C(n_477), .Y(n_893) );
INVx1_ASAP7_75t_L g894 ( .A(n_796), .Y(n_894) );
INVxp67_ASAP7_75t_SL g895 ( .A(n_808), .Y(n_895) );
INVx2_ASAP7_75t_L g896 ( .A(n_808), .Y(n_896) );
AOI21xp5_ASAP7_75t_L g897 ( .A1(n_755), .A2(n_632), .B(n_458), .Y(n_897) );
NAND2xp5_ASAP7_75t_L g898 ( .A(n_772), .B(n_580), .Y(n_898) );
INVx2_ASAP7_75t_L g899 ( .A(n_801), .Y(n_899) );
NAND2xp5_ASAP7_75t_L g900 ( .A(n_800), .B(n_587), .Y(n_900) );
OAI22xp33_ASAP7_75t_L g901 ( .A1(n_795), .A2(n_774), .B1(n_776), .B2(n_747), .Y(n_901) );
AND2x2_ASAP7_75t_L g902 ( .A(n_748), .B(n_774), .Y(n_902) );
INVx1_ASAP7_75t_SL g903 ( .A(n_738), .Y(n_903) );
NAND2xp5_ASAP7_75t_L g904 ( .A(n_800), .B(n_614), .Y(n_904) );
INVx2_ASAP7_75t_L g905 ( .A(n_801), .Y(n_905) );
INVx1_ASAP7_75t_SL g906 ( .A(n_738), .Y(n_906) );
CKINVDCx20_ASAP7_75t_R g907 ( .A(n_776), .Y(n_907) );
AND2x2_ASAP7_75t_L g908 ( .A(n_737), .B(n_614), .Y(n_908) );
A2O1A1Ixp33_ASAP7_75t_L g909 ( .A1(n_783), .A2(n_497), .B(n_500), .C(n_490), .Y(n_909) );
BUFx2_ASAP7_75t_L g910 ( .A(n_780), .Y(n_910) );
INVx1_ASAP7_75t_L g911 ( .A(n_777), .Y(n_911) );
INVx2_ASAP7_75t_L g912 ( .A(n_806), .Y(n_912) );
CKINVDCx11_ASAP7_75t_R g913 ( .A(n_747), .Y(n_913) );
INVx2_ASAP7_75t_L g914 ( .A(n_786), .Y(n_914) );
NAND2xp5_ASAP7_75t_L g915 ( .A(n_780), .B(n_642), .Y(n_915) );
INVx2_ASAP7_75t_L g916 ( .A(n_786), .Y(n_916) );
HB1xp67_ASAP7_75t_L g917 ( .A(n_787), .Y(n_917) );
INVx5_ASAP7_75t_L g918 ( .A(n_787), .Y(n_918) );
O2A1O1Ixp33_ASAP7_75t_L g919 ( .A1(n_778), .A2(n_677), .B(n_680), .C(n_676), .Y(n_919) );
AOI21xp5_ASAP7_75t_L g920 ( .A1(n_782), .A2(n_789), .B(n_785), .Y(n_920) );
NOR2xp33_ASAP7_75t_L g921 ( .A(n_794), .B(n_642), .Y(n_921) );
BUFx2_ASAP7_75t_L g922 ( .A(n_794), .Y(n_922) );
CKINVDCx5p33_ASAP7_75t_R g923 ( .A(n_769), .Y(n_923) );
AND2x2_ASAP7_75t_L g924 ( .A(n_798), .B(n_453), .Y(n_924) );
OAI22xp5_ASAP7_75t_L g925 ( .A1(n_790), .A2(n_513), .B1(n_518), .B2(n_512), .Y(n_925) );
INVx1_ASAP7_75t_L g926 ( .A(n_736), .Y(n_926) );
BUFx3_ASAP7_75t_L g927 ( .A(n_799), .Y(n_927) );
O2A1O1Ixp33_ASAP7_75t_L g928 ( .A1(n_793), .A2(n_680), .B(n_686), .C(n_677), .Y(n_928) );
AND2x4_ASAP7_75t_L g929 ( .A(n_749), .B(n_628), .Y(n_929) );
INVx3_ASAP7_75t_L g930 ( .A(n_756), .Y(n_930) );
NOR2xp67_ASAP7_75t_L g931 ( .A(n_746), .B(n_607), .Y(n_931) );
BUFx6f_ASAP7_75t_L g932 ( .A(n_763), .Y(n_932) );
INVx1_ASAP7_75t_L g933 ( .A(n_736), .Y(n_933) );
INVx2_ASAP7_75t_L g934 ( .A(n_736), .Y(n_934) );
INVx4_ASAP7_75t_L g935 ( .A(n_738), .Y(n_935) );
AOI21xp5_ASAP7_75t_L g936 ( .A1(n_802), .A2(n_460), .B(n_449), .Y(n_936) );
INVx2_ASAP7_75t_SL g937 ( .A(n_741), .Y(n_937) );
OAI22xp5_ASAP7_75t_SL g938 ( .A1(n_748), .A2(n_476), .B1(n_478), .B2(n_473), .Y(n_938) );
AOI22xp33_ASAP7_75t_SL g939 ( .A1(n_803), .A2(n_453), .B1(n_625), .B2(n_534), .Y(n_939) );
INVx1_ASAP7_75t_L g940 ( .A(n_736), .Y(n_940) );
O2A1O1Ixp33_ASAP7_75t_L g941 ( .A1(n_793), .A2(n_687), .B(n_691), .C(n_686), .Y(n_941) );
AO21x2_ASAP7_75t_L g942 ( .A1(n_835), .A2(n_560), .B(n_566), .Y(n_942) );
NAND2xp5_ASAP7_75t_L g943 ( .A(n_861), .B(n_520), .Y(n_943) );
BUFx12f_ASAP7_75t_L g944 ( .A(n_860), .Y(n_944) );
AOI22x1_ASAP7_75t_L g945 ( .A1(n_936), .A2(n_667), .B1(n_672), .B2(n_668), .Y(n_945) );
INVx2_ASAP7_75t_L g946 ( .A(n_839), .Y(n_946) );
INVx2_ASAP7_75t_SL g947 ( .A(n_927), .Y(n_947) );
OAI21x1_ASAP7_75t_L g948 ( .A1(n_835), .A2(n_450), .B(n_438), .Y(n_948) );
NAND2xp5_ASAP7_75t_L g949 ( .A(n_891), .B(n_524), .Y(n_949) );
O2A1O1Ixp33_ASAP7_75t_SL g950 ( .A1(n_816), .A2(n_464), .B(n_468), .C(n_462), .Y(n_950) );
A2O1A1Ixp33_ASAP7_75t_L g951 ( .A1(n_852), .A2(n_597), .B(n_471), .C(n_482), .Y(n_951) );
AND2x4_ASAP7_75t_L g952 ( .A(n_896), .B(n_687), .Y(n_952) );
INVx1_ASAP7_75t_L g953 ( .A(n_856), .Y(n_953) );
OAI21x1_ASAP7_75t_L g954 ( .A1(n_936), .A2(n_920), .B(n_852), .Y(n_954) );
OA21x2_ASAP7_75t_L g955 ( .A1(n_816), .A2(n_526), .B(n_502), .Y(n_955) );
INVx1_ASAP7_75t_SL g956 ( .A(n_828), .Y(n_956) );
NAND3xp33_ASAP7_75t_L g957 ( .A(n_819), .B(n_691), .C(n_599), .Y(n_957) );
INVx1_ASAP7_75t_L g958 ( .A(n_853), .Y(n_958) );
OAI21x1_ASAP7_75t_L g959 ( .A1(n_920), .A2(n_562), .B(n_550), .Y(n_959) );
INVxp67_ASAP7_75t_SL g960 ( .A(n_895), .Y(n_960) );
INVxp67_ASAP7_75t_L g961 ( .A(n_840), .Y(n_961) );
AO21x2_ASAP7_75t_L g962 ( .A1(n_894), .A2(n_489), .B(n_480), .Y(n_962) );
BUFx4_ASAP7_75t_SL g963 ( .A(n_817), .Y(n_963) );
OAI21x1_ASAP7_75t_L g964 ( .A1(n_912), .A2(n_562), .B(n_550), .Y(n_964) );
BUFx6f_ASAP7_75t_L g965 ( .A(n_821), .Y(n_965) );
INVx2_ASAP7_75t_SL g966 ( .A(n_833), .Y(n_966) );
OA21x2_ASAP7_75t_L g967 ( .A1(n_845), .A2(n_617), .B(n_579), .Y(n_967) );
AO21x2_ASAP7_75t_L g968 ( .A1(n_919), .A2(n_493), .B(n_492), .Y(n_968) );
INVx1_ASAP7_75t_L g969 ( .A(n_818), .Y(n_969) );
OAI21x1_ASAP7_75t_L g970 ( .A1(n_854), .A2(n_617), .B(n_579), .Y(n_970) );
AO21x2_ASAP7_75t_L g971 ( .A1(n_919), .A2(n_495), .B(n_494), .Y(n_971) );
AOI22xp33_ASAP7_75t_L g972 ( .A1(n_902), .A2(n_565), .B1(n_532), .B2(n_555), .Y(n_972) );
OAI21xp5_ASAP7_75t_L g973 ( .A1(n_911), .A2(n_503), .B(n_499), .Y(n_973) );
INVx1_ASAP7_75t_SL g974 ( .A(n_846), .Y(n_974) );
INVx1_ASAP7_75t_L g975 ( .A(n_934), .Y(n_975) );
NAND2xp5_ASAP7_75t_SL g976 ( .A(n_923), .B(n_623), .Y(n_976) );
BUFx6f_ASAP7_75t_L g977 ( .A(n_821), .Y(n_977) );
O2A1O1Ixp33_ASAP7_75t_L g978 ( .A1(n_849), .A2(n_547), .B(n_557), .C(n_556), .Y(n_978) );
AOI21x1_ASAP7_75t_L g979 ( .A1(n_897), .A2(n_648), .B(n_510), .Y(n_979) );
NOR2xp33_ASAP7_75t_L g980 ( .A(n_838), .B(n_536), .Y(n_980) );
BUFx3_ASAP7_75t_L g981 ( .A(n_823), .Y(n_981) );
AO21x2_ASAP7_75t_L g982 ( .A1(n_897), .A2(n_515), .B(n_505), .Y(n_982) );
OAI21x1_ASAP7_75t_L g983 ( .A1(n_870), .A2(n_648), .B(n_519), .Y(n_983) );
AOI21xp5_ASAP7_75t_L g984 ( .A1(n_858), .A2(n_706), .B(n_697), .Y(n_984) );
AOI22xp33_ASAP7_75t_L g985 ( .A1(n_901), .A2(n_565), .B1(n_569), .B2(n_567), .Y(n_985) );
INVx2_ASAP7_75t_L g986 ( .A(n_872), .Y(n_986) );
AOI22xp33_ASAP7_75t_L g987 ( .A1(n_873), .A2(n_565), .B1(n_575), .B2(n_570), .Y(n_987) );
NAND2xp5_ASAP7_75t_L g988 ( .A(n_871), .B(n_582), .Y(n_988) );
INVx1_ASAP7_75t_L g989 ( .A(n_837), .Y(n_989) );
OAI21x1_ASAP7_75t_L g990 ( .A1(n_878), .A2(n_527), .B(n_516), .Y(n_990) );
OAI21x1_ASAP7_75t_L g991 ( .A1(n_881), .A2(n_530), .B(n_529), .Y(n_991) );
NOR2xp33_ASAP7_75t_L g992 ( .A(n_843), .B(n_453), .Y(n_992) );
AOI22xp33_ASAP7_75t_L g993 ( .A1(n_873), .A2(n_565), .B1(n_594), .B2(n_586), .Y(n_993) );
O2A1O1Ixp33_ASAP7_75t_SL g994 ( .A1(n_880), .A2(n_539), .B(n_545), .C(n_535), .Y(n_994) );
AOI22xp33_ASAP7_75t_L g995 ( .A1(n_830), .A2(n_598), .B1(n_600), .B2(n_595), .Y(n_995) );
AND2x4_ASAP7_75t_L g996 ( .A(n_866), .B(n_602), .Y(n_996) );
INVx1_ASAP7_75t_L g997 ( .A(n_926), .Y(n_997) );
AND2x4_ASAP7_75t_L g998 ( .A(n_865), .B(n_604), .Y(n_998) );
OAI21x1_ASAP7_75t_L g999 ( .A1(n_883), .A2(n_551), .B(n_548), .Y(n_999) );
INVx2_ASAP7_75t_SL g1000 ( .A(n_824), .Y(n_1000) );
BUFx2_ASAP7_75t_SL g1001 ( .A(n_832), .Y(n_1001) );
A2O1A1Ixp33_ASAP7_75t_L g1002 ( .A1(n_822), .A2(n_559), .B(n_574), .C(n_563), .Y(n_1002) );
INVx1_ASAP7_75t_SL g1003 ( .A(n_910), .Y(n_1003) );
INVx1_ASAP7_75t_L g1004 ( .A(n_933), .Y(n_1004) );
OAI22xp33_ASAP7_75t_L g1005 ( .A1(n_811), .A2(n_608), .B1(n_619), .B2(n_605), .Y(n_1005) );
OAI21x1_ASAP7_75t_SL g1006 ( .A1(n_822), .A2(n_584), .B(n_578), .Y(n_1006) );
INVx2_ASAP7_75t_L g1007 ( .A(n_940), .Y(n_1007) );
INVx1_ASAP7_75t_L g1008 ( .A(n_830), .Y(n_1008) );
AO31x2_ASAP7_75t_L g1009 ( .A1(n_925), .A2(n_672), .A3(n_673), .B(n_668), .Y(n_1009) );
AND2x4_ASAP7_75t_SL g1010 ( .A(n_811), .B(n_624), .Y(n_1010) );
AOI21xp5_ASAP7_75t_L g1011 ( .A1(n_858), .A2(n_706), .B(n_697), .Y(n_1011) );
OAI21xp5_ASAP7_75t_L g1012 ( .A1(n_864), .A2(n_591), .B(n_589), .Y(n_1012) );
OAI21x1_ASAP7_75t_L g1013 ( .A1(n_864), .A2(n_612), .B(n_596), .Y(n_1013) );
INVx1_ASAP7_75t_L g1014 ( .A(n_937), .Y(n_1014) );
OA21x2_ASAP7_75t_L g1015 ( .A1(n_909), .A2(n_615), .B(n_613), .Y(n_1015) );
NOR2xp67_ASAP7_75t_L g1016 ( .A(n_876), .B(n_13), .Y(n_1016) );
OR2x6_ASAP7_75t_L g1017 ( .A(n_811), .B(n_629), .Y(n_1017) );
BUFx3_ASAP7_75t_L g1018 ( .A(n_887), .Y(n_1018) );
OR2x2_ASAP7_75t_L g1019 ( .A(n_834), .B(n_630), .Y(n_1019) );
NAND2x1p5_ASAP7_75t_L g1020 ( .A(n_829), .B(n_831), .Y(n_1020) );
OA21x2_ASAP7_75t_L g1021 ( .A1(n_812), .A2(n_622), .B(n_616), .Y(n_1021) );
AOI22xp5_ASAP7_75t_L g1022 ( .A1(n_815), .A2(n_638), .B1(n_623), .B2(n_633), .Y(n_1022) );
OAI21x1_ASAP7_75t_SL g1023 ( .A1(n_928), .A2(n_627), .B(n_626), .Y(n_1023) );
AO21x2_ASAP7_75t_L g1024 ( .A1(n_925), .A2(n_635), .B(n_634), .Y(n_1024) );
OA21x2_ASAP7_75t_L g1025 ( .A1(n_879), .A2(n_639), .B(n_636), .Y(n_1025) );
INVx2_ASAP7_75t_L g1026 ( .A(n_914), .Y(n_1026) );
OR2x6_ASAP7_75t_L g1027 ( .A(n_848), .B(n_640), .Y(n_1027) );
OA21x2_ASAP7_75t_L g1028 ( .A1(n_879), .A2(n_646), .B(n_644), .Y(n_1028) );
OAI21x1_ASAP7_75t_L g1029 ( .A1(n_928), .A2(n_649), .B(n_707), .Y(n_1029) );
O2A1O1Ixp5_ASAP7_75t_L g1030 ( .A1(n_869), .A2(n_672), .B(n_673), .C(n_668), .Y(n_1030) );
OAI21x1_ASAP7_75t_L g1031 ( .A1(n_941), .A2(n_713), .B(n_707), .Y(n_1031) );
AND2x4_ASAP7_75t_L g1032 ( .A(n_829), .B(n_641), .Y(n_1032) );
INVx1_ASAP7_75t_L g1033 ( .A(n_820), .Y(n_1033) );
NAND2xp5_ASAP7_75t_L g1034 ( .A(n_884), .B(n_643), .Y(n_1034) );
AOI22xp33_ASAP7_75t_L g1035 ( .A1(n_938), .A2(n_638), .B1(n_610), .B2(n_558), .Y(n_1035) );
INVx1_ASAP7_75t_L g1036 ( .A(n_820), .Y(n_1036) );
INVx3_ASAP7_75t_L g1037 ( .A(n_831), .Y(n_1037) );
INVx2_ASAP7_75t_L g1038 ( .A(n_916), .Y(n_1038) );
INVx2_ASAP7_75t_L g1039 ( .A(n_930), .Y(n_1039) );
O2A1O1Ixp33_ASAP7_75t_L g1040 ( .A1(n_886), .A2(n_678), .B(n_689), .C(n_673), .Y(n_1040) );
INVx1_ASAP7_75t_SL g1041 ( .A(n_922), .Y(n_1041) );
AOI21x1_ASAP7_75t_L g1042 ( .A1(n_869), .A2(n_689), .B(n_678), .Y(n_1042) );
OAI21x1_ASAP7_75t_SL g1043 ( .A1(n_941), .A2(n_689), .B(n_678), .Y(n_1043) );
INVx1_ASAP7_75t_L g1044 ( .A(n_855), .Y(n_1044) );
CKINVDCx5p33_ASAP7_75t_R g1045 ( .A(n_913), .Y(n_1045) );
A2O1A1Ixp33_ASAP7_75t_L g1046 ( .A1(n_889), .A2(n_483), .B(n_496), .C(n_488), .Y(n_1046) );
AND2x4_ASAP7_75t_L g1047 ( .A(n_930), .B(n_851), .Y(n_1047) );
NOR2xp33_ASAP7_75t_L g1048 ( .A(n_857), .B(n_533), .Y(n_1048) );
BUFx2_ASAP7_75t_R g1049 ( .A(n_863), .Y(n_1049) );
OAI22xp5_ASAP7_75t_L g1050 ( .A1(n_875), .A2(n_521), .B1(n_523), .B2(n_481), .Y(n_1050) );
AND2x4_ASAP7_75t_L g1051 ( .A(n_918), .B(n_14), .Y(n_1051) );
OR2x2_ASAP7_75t_L g1052 ( .A(n_850), .B(n_14), .Y(n_1052) );
NAND2xp5_ASAP7_75t_L g1053 ( .A(n_855), .B(n_525), .Y(n_1053) );
NOR2xp33_ASAP7_75t_L g1054 ( .A(n_877), .B(n_15), .Y(n_1054) );
NAND2x1p5_ASAP7_75t_L g1055 ( .A(n_918), .B(n_663), .Y(n_1055) );
INVx1_ASAP7_75t_L g1056 ( .A(n_893), .Y(n_1056) );
OAI22xp5_ASAP7_75t_L g1057 ( .A1(n_841), .A2(n_541), .B1(n_540), .B2(n_663), .Y(n_1057) );
O2A1O1Ixp33_ASAP7_75t_L g1058 ( .A1(n_882), .A2(n_725), .B(n_713), .C(n_724), .Y(n_1058) );
OAI21x1_ASAP7_75t_L g1059 ( .A1(n_899), .A2(n_713), .B(n_707), .Y(n_1059) );
OAI21x1_ASAP7_75t_SL g1060 ( .A1(n_915), .A2(n_15), .B(n_16), .Y(n_1060) );
INVx2_ASAP7_75t_L g1061 ( .A(n_905), .Y(n_1061) );
INVx1_ASAP7_75t_L g1062 ( .A(n_924), .Y(n_1062) );
OAI21x1_ASAP7_75t_L g1063 ( .A1(n_842), .A2(n_847), .B(n_915), .Y(n_1063) );
AOI22xp5_ASAP7_75t_L g1064 ( .A1(n_827), .A2(n_669), .B1(n_679), .B2(n_663), .Y(n_1064) );
INVx3_ASAP7_75t_L g1065 ( .A(n_935), .Y(n_1065) );
NAND2xp5_ASAP7_75t_L g1066 ( .A(n_882), .B(n_16), .Y(n_1066) );
OA21x2_ASAP7_75t_L g1067 ( .A1(n_929), .A2(n_724), .B(n_669), .Y(n_1067) );
INVx2_ASAP7_75t_SL g1068 ( .A(n_908), .Y(n_1068) );
CKINVDCx5p33_ASAP7_75t_R g1069 ( .A(n_939), .Y(n_1069) );
AO21x2_ASAP7_75t_L g1070 ( .A1(n_929), .A2(n_724), .B(n_669), .Y(n_1070) );
OAI21xp5_ASAP7_75t_L g1071 ( .A1(n_898), .A2(n_725), .B(n_720), .Y(n_1071) );
INVx1_ASAP7_75t_L g1072 ( .A(n_898), .Y(n_1072) );
INVx4_ASAP7_75t_L g1073 ( .A(n_813), .Y(n_1073) );
NAND2xp5_ASAP7_75t_L g1074 ( .A(n_900), .B(n_17), .Y(n_1074) );
OAI22xp5_ASAP7_75t_L g1075 ( .A1(n_885), .A2(n_669), .B1(n_679), .B2(n_663), .Y(n_1075) );
AOI22xp33_ASAP7_75t_L g1076 ( .A1(n_900), .A2(n_679), .B1(n_690), .B2(n_669), .Y(n_1076) );
INVxp67_ASAP7_75t_L g1077 ( .A(n_917), .Y(n_1077) );
OA21x2_ASAP7_75t_L g1078 ( .A1(n_904), .A2(n_679), .B(n_669), .Y(n_1078) );
OAI222xp33_ASAP7_75t_L g1079 ( .A1(n_859), .A2(n_17), .B1(n_19), .B2(n_20), .C1(n_21), .C2(n_22), .Y(n_1079) );
AO21x2_ASAP7_75t_L g1080 ( .A1(n_904), .A2(n_690), .B(n_679), .Y(n_1080) );
INVx1_ASAP7_75t_L g1081 ( .A(n_814), .Y(n_1081) );
INVx2_ASAP7_75t_L g1082 ( .A(n_874), .Y(n_1082) );
A2O1A1Ixp33_ASAP7_75t_L g1083 ( .A1(n_921), .A2(n_690), .B(n_679), .C(n_725), .Y(n_1083) );
OAI21xp5_ASAP7_75t_L g1084 ( .A1(n_814), .A2(n_720), .B(n_690), .Y(n_1084) );
AO31x2_ASAP7_75t_L g1085 ( .A1(n_935), .A2(n_690), .A3(n_705), .B(n_21), .Y(n_1085) );
INVx1_ASAP7_75t_L g1086 ( .A(n_888), .Y(n_1086) );
AOI21x1_ASAP7_75t_L g1087 ( .A1(n_867), .A2(n_690), .B(n_705), .Y(n_1087) );
BUFx6f_ASAP7_75t_L g1088 ( .A(n_821), .Y(n_1088) );
INVx6_ASAP7_75t_L g1089 ( .A(n_813), .Y(n_1089) );
OAI21x1_ASAP7_75t_L g1090 ( .A1(n_931), .A2(n_193), .B(n_189), .Y(n_1090) );
NOR2x1_ASAP7_75t_SL g1091 ( .A(n_918), .B(n_19), .Y(n_1091) );
AO31x2_ASAP7_75t_L g1092 ( .A1(n_813), .A2(n_705), .A3(n_24), .B(n_20), .Y(n_1092) );
A2O1A1Ixp33_ASAP7_75t_L g1093 ( .A1(n_890), .A2(n_720), .B(n_705), .C(n_25), .Y(n_1093) );
BUFx6f_ASAP7_75t_L g1094 ( .A(n_825), .Y(n_1094) );
INVx2_ASAP7_75t_L g1095 ( .A(n_874), .Y(n_1095) );
AOI22xp33_ASAP7_75t_L g1096 ( .A1(n_918), .A2(n_705), .B1(n_720), .B2(n_25), .Y(n_1096) );
OAI21x1_ASAP7_75t_SL g1097 ( .A1(n_825), .A2(n_23), .B(n_24), .Y(n_1097) );
OR2x6_ASAP7_75t_L g1098 ( .A(n_892), .B(n_26), .Y(n_1098) );
NOR2xp33_ASAP7_75t_L g1099 ( .A(n_907), .B(n_27), .Y(n_1099) );
AO21x2_ASAP7_75t_L g1100 ( .A1(n_825), .A2(n_705), .B(n_195), .Y(n_1100) );
AO21x2_ASAP7_75t_L g1101 ( .A1(n_826), .A2(n_196), .B(n_194), .Y(n_1101) );
OAI21x1_ASAP7_75t_L g1102 ( .A1(n_826), .A2(n_200), .B(n_197), .Y(n_1102) );
AOI221xp5_ASAP7_75t_L g1103 ( .A1(n_903), .A2(n_720), .B1(n_29), .B2(n_27), .C(n_28), .Y(n_1103) );
INVx2_ASAP7_75t_L g1104 ( .A(n_892), .Y(n_1104) );
OAI21x1_ASAP7_75t_L g1105 ( .A1(n_826), .A2(n_205), .B(n_202), .Y(n_1105) );
AOI22xp33_ASAP7_75t_L g1106 ( .A1(n_1017), .A2(n_862), .B1(n_892), .B2(n_903), .Y(n_1106) );
AND2x2_ASAP7_75t_L g1107 ( .A(n_1019), .B(n_862), .Y(n_1107) );
AOI22xp5_ASAP7_75t_L g1108 ( .A1(n_960), .A2(n_906), .B1(n_836), .B2(n_868), .Y(n_1108) );
OR2x2_ASAP7_75t_L g1109 ( .A(n_956), .B(n_906), .Y(n_1109) );
AOI22xp5_ASAP7_75t_L g1110 ( .A1(n_960), .A2(n_836), .B1(n_868), .B2(n_844), .Y(n_1110) );
OAI221xp5_ASAP7_75t_L g1111 ( .A1(n_1048), .A2(n_844), .B1(n_932), .B2(n_868), .C(n_836), .Y(n_1111) );
AOI222xp33_ASAP7_75t_L g1112 ( .A1(n_1054), .A2(n_932), .B1(n_29), .B2(n_30), .C1(n_31), .C2(n_32), .Y(n_1112) );
INVx1_ASAP7_75t_L g1113 ( .A(n_953), .Y(n_1113) );
OR2x2_ASAP7_75t_L g1114 ( .A(n_956), .B(n_28), .Y(n_1114) );
AND2x2_ASAP7_75t_L g1115 ( .A(n_998), .B(n_32), .Y(n_1115) );
AOI22xp33_ASAP7_75t_L g1116 ( .A1(n_1017), .A2(n_720), .B1(n_35), .B2(n_33), .Y(n_1116) );
OAI22xp5_ASAP7_75t_L g1117 ( .A1(n_985), .A2(n_36), .B1(n_34), .B2(n_35), .Y(n_1117) );
NAND2xp5_ASAP7_75t_L g1118 ( .A(n_1033), .B(n_37), .Y(n_1118) );
AOI22xp5_ASAP7_75t_L g1119 ( .A1(n_980), .A2(n_720), .B1(n_39), .B2(n_37), .Y(n_1119) );
AND2x2_ASAP7_75t_L g1120 ( .A(n_998), .B(n_38), .Y(n_1120) );
NAND3xp33_ASAP7_75t_L g1121 ( .A(n_957), .B(n_38), .C(n_40), .Y(n_1121) );
AOI22xp33_ASAP7_75t_SL g1122 ( .A1(n_1010), .A2(n_44), .B1(n_42), .B2(n_43), .Y(n_1122) );
NAND2xp5_ASAP7_75t_L g1123 ( .A(n_1036), .B(n_42), .Y(n_1123) );
CKINVDCx14_ASAP7_75t_R g1124 ( .A(n_963), .Y(n_1124) );
OR2x2_ASAP7_75t_L g1125 ( .A(n_1052), .B(n_43), .Y(n_1125) );
OAI211xp5_ASAP7_75t_L g1126 ( .A1(n_1035), .A2(n_46), .B(n_44), .C(n_45), .Y(n_1126) );
INVx2_ASAP7_75t_L g1127 ( .A(n_1007), .Y(n_1127) );
INVx1_ASAP7_75t_L g1128 ( .A(n_958), .Y(n_1128) );
AO21x2_ASAP7_75t_L g1129 ( .A1(n_942), .A2(n_209), .B(n_207), .Y(n_1129) );
AND2x2_ASAP7_75t_L g1130 ( .A(n_980), .B(n_45), .Y(n_1130) );
INVx3_ASAP7_75t_L g1131 ( .A(n_1089), .Y(n_1131) );
INVx1_ASAP7_75t_L g1132 ( .A(n_1008), .Y(n_1132) );
OAI211xp5_ASAP7_75t_L g1133 ( .A1(n_1035), .A2(n_51), .B(n_49), .C(n_50), .Y(n_1133) );
AND2x4_ASAP7_75t_L g1134 ( .A(n_974), .B(n_50), .Y(n_1134) );
OAI22xp5_ASAP7_75t_L g1135 ( .A1(n_985), .A2(n_53), .B1(n_51), .B2(n_52), .Y(n_1135) );
OAI211xp5_ASAP7_75t_SL g1136 ( .A1(n_995), .A2(n_55), .B(n_53), .C(n_54), .Y(n_1136) );
AOI221xp5_ASAP7_75t_L g1137 ( .A1(n_1005), .A2(n_56), .B1(n_58), .B2(n_59), .C(n_60), .Y(n_1137) );
INVx1_ASAP7_75t_L g1138 ( .A(n_989), .Y(n_1138) );
AND2x4_ASAP7_75t_L g1139 ( .A(n_974), .B(n_59), .Y(n_1139) );
AOI22xp5_ASAP7_75t_L g1140 ( .A1(n_1069), .A2(n_62), .B1(n_60), .B2(n_61), .Y(n_1140) );
AOI22xp33_ASAP7_75t_L g1141 ( .A1(n_1017), .A2(n_64), .B1(n_61), .B2(n_63), .Y(n_1141) );
AOI22xp33_ASAP7_75t_SL g1142 ( .A1(n_1054), .A2(n_65), .B1(n_63), .B2(n_64), .Y(n_1142) );
AOI22xp33_ASAP7_75t_L g1143 ( .A1(n_1005), .A2(n_67), .B1(n_65), .B2(n_66), .Y(n_1143) );
AOI31xp33_ASAP7_75t_L g1144 ( .A1(n_1103), .A2(n_68), .A3(n_66), .B(n_67), .Y(n_1144) );
AND2x2_ASAP7_75t_L g1145 ( .A(n_1027), .B(n_68), .Y(n_1145) );
BUFx2_ASAP7_75t_L g1146 ( .A(n_961), .Y(n_1146) );
AOI22xp33_ASAP7_75t_SL g1147 ( .A1(n_1099), .A2(n_71), .B1(n_69), .B2(n_70), .Y(n_1147) );
OAI21xp5_ASAP7_75t_L g1148 ( .A1(n_954), .A2(n_70), .B(n_71), .Y(n_1148) );
INVxp67_ASAP7_75t_L g1149 ( .A(n_1099), .Y(n_1149) );
AND2x2_ASAP7_75t_L g1150 ( .A(n_1027), .B(n_72), .Y(n_1150) );
AOI222xp33_ASAP7_75t_L g1151 ( .A1(n_1044), .A2(n_72), .B1(n_73), .B2(n_74), .C1(n_75), .C2(n_76), .Y(n_1151) );
AOI22xp33_ASAP7_75t_L g1152 ( .A1(n_1068), .A2(n_77), .B1(n_75), .B2(n_76), .Y(n_1152) );
AOI221xp5_ASAP7_75t_L g1153 ( .A1(n_1034), .A2(n_78), .B1(n_80), .B2(n_81), .C(n_82), .Y(n_1153) );
AOI21xp5_ASAP7_75t_L g1154 ( .A1(n_1058), .A2(n_216), .B(n_215), .Y(n_1154) );
OAI22xp5_ASAP7_75t_L g1155 ( .A1(n_1098), .A2(n_81), .B1(n_78), .B2(n_80), .Y(n_1155) );
INVx2_ASAP7_75t_L g1156 ( .A(n_946), .Y(n_1156) );
OR2x2_ASAP7_75t_L g1157 ( .A(n_961), .B(n_82), .Y(n_1157) );
AOI221xp5_ASAP7_75t_L g1158 ( .A1(n_1034), .A2(n_83), .B1(n_84), .B2(n_85), .C(n_86), .Y(n_1158) );
AOI22xp33_ASAP7_75t_L g1159 ( .A1(n_1048), .A2(n_87), .B1(n_84), .B2(n_86), .Y(n_1159) );
AOI22xp33_ASAP7_75t_SL g1160 ( .A1(n_1091), .A2(n_89), .B1(n_87), .B2(n_88), .Y(n_1160) );
AOI21xp5_ASAP7_75t_L g1161 ( .A1(n_948), .A2(n_228), .B(n_227), .Y(n_1161) );
OAI22xp5_ASAP7_75t_L g1162 ( .A1(n_1098), .A2(n_92), .B1(n_90), .B2(n_91), .Y(n_1162) );
AOI21xp5_ASAP7_75t_L g1163 ( .A1(n_959), .A2(n_230), .B(n_229), .Y(n_1163) );
A2O1A1Ixp33_ASAP7_75t_L g1164 ( .A1(n_978), .A2(n_93), .B(n_91), .C(n_92), .Y(n_1164) );
NAND2xp5_ASAP7_75t_L g1165 ( .A(n_1081), .B(n_93), .Y(n_1165) );
AOI221xp5_ASAP7_75t_L g1166 ( .A1(n_995), .A2(n_94), .B1(n_95), .B2(n_96), .C(n_97), .Y(n_1166) );
AOI21xp5_ASAP7_75t_L g1167 ( .A1(n_984), .A2(n_232), .B(n_231), .Y(n_1167) );
AND2x2_ASAP7_75t_L g1168 ( .A(n_1027), .B(n_96), .Y(n_1168) );
AOI221xp5_ASAP7_75t_L g1169 ( .A1(n_978), .A2(n_97), .B1(n_99), .B2(n_100), .C(n_101), .Y(n_1169) );
AOI221xp5_ASAP7_75t_L g1170 ( .A1(n_1062), .A2(n_99), .B1(n_100), .B2(n_103), .C(n_104), .Y(n_1170) );
AOI22xp33_ASAP7_75t_L g1171 ( .A1(n_996), .A2(n_103), .B1(n_106), .B2(n_108), .Y(n_1171) );
A2O1A1Ixp33_ASAP7_75t_L g1172 ( .A1(n_1072), .A2(n_106), .B(n_109), .C(n_110), .Y(n_1172) );
OAI22xp5_ASAP7_75t_L g1173 ( .A1(n_1098), .A2(n_109), .B1(n_110), .B2(n_111), .Y(n_1173) );
O2A1O1Ixp33_ASAP7_75t_L g1174 ( .A1(n_1046), .A2(n_111), .B(n_113), .C(n_114), .Y(n_1174) );
AOI22xp33_ASAP7_75t_L g1175 ( .A1(n_996), .A2(n_113), .B1(n_114), .B2(n_115), .Y(n_1175) );
A2O1A1Ixp33_ASAP7_75t_L g1176 ( .A1(n_1056), .A2(n_116), .B(n_117), .C(n_118), .Y(n_1176) );
BUFx3_ASAP7_75t_L g1177 ( .A(n_981), .Y(n_1177) );
OAI22xp33_ASAP7_75t_L g1178 ( .A1(n_1003), .A2(n_117), .B1(n_121), .B2(n_122), .Y(n_1178) );
AOI221xp5_ASAP7_75t_L g1179 ( .A1(n_992), .A2(n_123), .B1(n_124), .B2(n_125), .C(n_126), .Y(n_1179) );
CKINVDCx5p33_ASAP7_75t_R g1180 ( .A(n_963), .Y(n_1180) );
NAND2xp5_ASAP7_75t_L g1181 ( .A(n_1003), .B(n_125), .Y(n_1181) );
AO21x2_ASAP7_75t_L g1182 ( .A1(n_942), .A2(n_234), .B(n_233), .Y(n_1182) );
OR2x2_ASAP7_75t_L g1183 ( .A(n_1050), .B(n_126), .Y(n_1183) );
AND2x2_ASAP7_75t_L g1184 ( .A(n_1041), .B(n_128), .Y(n_1184) );
AOI22xp33_ASAP7_75t_L g1185 ( .A1(n_992), .A2(n_128), .B1(n_129), .B2(n_130), .Y(n_1185) );
AND2x2_ASAP7_75t_L g1186 ( .A(n_1041), .B(n_129), .Y(n_1186) );
NOR3xp33_ASAP7_75t_SL g1187 ( .A(n_1045), .B(n_130), .C(n_131), .Y(n_1187) );
OAI221xp5_ASAP7_75t_L g1188 ( .A1(n_1022), .A2(n_131), .B1(n_132), .B2(n_133), .C(n_134), .Y(n_1188) );
INVx1_ASAP7_75t_L g1189 ( .A(n_997), .Y(n_1189) );
NAND3xp33_ASAP7_75t_L g1190 ( .A(n_951), .B(n_136), .C(n_137), .Y(n_1190) );
AND2x2_ASAP7_75t_L g1191 ( .A(n_952), .B(n_136), .Y(n_1191) );
INVx1_ASAP7_75t_L g1192 ( .A(n_1004), .Y(n_1192) );
OAI211xp5_ASAP7_75t_L g1193 ( .A1(n_972), .A2(n_137), .B(n_138), .C(n_139), .Y(n_1193) );
OAI22xp5_ASAP7_75t_L g1194 ( .A1(n_987), .A2(n_138), .B1(n_139), .B2(n_140), .Y(n_1194) );
AOI221xp5_ASAP7_75t_L g1195 ( .A1(n_943), .A2(n_140), .B1(n_141), .B2(n_142), .C(n_143), .Y(n_1195) );
OR2x2_ASAP7_75t_L g1196 ( .A(n_1050), .B(n_141), .Y(n_1196) );
OAI22xp33_ASAP7_75t_L g1197 ( .A1(n_1077), .A2(n_142), .B1(n_143), .B2(n_144), .Y(n_1197) );
OAI22xp33_ASAP7_75t_L g1198 ( .A1(n_1077), .A2(n_146), .B1(n_147), .B2(n_149), .Y(n_1198) );
HB1xp67_ASAP7_75t_L g1199 ( .A(n_1051), .Y(n_1199) );
AOI22xp33_ASAP7_75t_L g1200 ( .A1(n_1086), .A2(n_147), .B1(n_149), .B2(n_150), .Y(n_1200) );
INVx1_ASAP7_75t_L g1201 ( .A(n_969), .Y(n_1201) );
OAI211xp5_ASAP7_75t_L g1202 ( .A1(n_972), .A2(n_150), .B(n_151), .C(n_152), .Y(n_1202) );
INVx2_ASAP7_75t_L g1203 ( .A(n_986), .Y(n_1203) );
CKINVDCx8_ASAP7_75t_R g1204 ( .A(n_1001), .Y(n_1204) );
INVx4_ASAP7_75t_SL g1205 ( .A(n_1089), .Y(n_1205) );
AOI22xp33_ASAP7_75t_SL g1206 ( .A1(n_1051), .A2(n_151), .B1(n_152), .B2(n_153), .Y(n_1206) );
AOI22xp33_ASAP7_75t_L g1207 ( .A1(n_1075), .A2(n_1032), .B1(n_1057), .B2(n_1014), .Y(n_1207) );
OAI22xp5_ASAP7_75t_L g1208 ( .A1(n_987), .A2(n_153), .B1(n_154), .B2(n_155), .Y(n_1208) );
AOI22xp33_ASAP7_75t_L g1209 ( .A1(n_1075), .A2(n_1032), .B1(n_1084), .B2(n_1024), .Y(n_1209) );
INVx2_ASAP7_75t_L g1210 ( .A(n_975), .Y(n_1210) );
AND2x2_ASAP7_75t_L g1211 ( .A(n_952), .B(n_155), .Y(n_1211) );
AOI21xp5_ASAP7_75t_L g1212 ( .A1(n_984), .A2(n_238), .B(n_236), .Y(n_1212) );
OAI221xp5_ASAP7_75t_L g1213 ( .A1(n_943), .A2(n_156), .B1(n_157), .B2(n_158), .C(n_159), .Y(n_1213) );
INVx2_ASAP7_75t_L g1214 ( .A(n_1067), .Y(n_1214) );
INVx1_ASAP7_75t_SL g1215 ( .A(n_966), .Y(n_1215) );
BUFx12f_ASAP7_75t_L g1216 ( .A(n_1000), .Y(n_1216) );
OR2x2_ASAP7_75t_L g1217 ( .A(n_988), .B(n_156), .Y(n_1217) );
INVx2_ASAP7_75t_L g1218 ( .A(n_1067), .Y(n_1218) );
INVx1_ASAP7_75t_L g1219 ( .A(n_988), .Y(n_1219) );
CKINVDCx5p33_ASAP7_75t_R g1220 ( .A(n_944), .Y(n_1220) );
OR2x2_ASAP7_75t_SL g1221 ( .A(n_1049), .B(n_157), .Y(n_1221) );
BUFx3_ASAP7_75t_L g1222 ( .A(n_947), .Y(n_1222) );
OA21x2_ASAP7_75t_L g1223 ( .A1(n_970), .A2(n_241), .B(n_240), .Y(n_1223) );
INVx2_ASAP7_75t_L g1224 ( .A(n_1070), .Y(n_1224) );
NOR2xp33_ASAP7_75t_L g1225 ( .A(n_976), .B(n_158), .Y(n_1225) );
HB1xp67_ASAP7_75t_L g1226 ( .A(n_1047), .Y(n_1226) );
CKINVDCx20_ASAP7_75t_R g1227 ( .A(n_1018), .Y(n_1227) );
OR2x2_ASAP7_75t_L g1228 ( .A(n_949), .B(n_160), .Y(n_1228) );
OAI22xp5_ASAP7_75t_L g1229 ( .A1(n_1066), .A2(n_160), .B1(n_161), .B2(n_162), .Y(n_1229) );
AOI211xp5_ASAP7_75t_SL g1230 ( .A1(n_1079), .A2(n_161), .B(n_162), .C(n_164), .Y(n_1230) );
NOR2xp33_ASAP7_75t_L g1231 ( .A(n_1049), .B(n_1053), .Y(n_1231) );
CKINVDCx12_ASAP7_75t_R g1232 ( .A(n_1026), .Y(n_1232) );
HB1xp67_ASAP7_75t_L g1233 ( .A(n_1047), .Y(n_1233) );
OAI21xp5_ASAP7_75t_L g1234 ( .A1(n_1066), .A2(n_165), .B(n_166), .Y(n_1234) );
HB1xp67_ASAP7_75t_L g1235 ( .A(n_1084), .Y(n_1235) );
AOI21xp5_ASAP7_75t_L g1236 ( .A1(n_1011), .A2(n_330), .B(n_420), .Y(n_1236) );
AOI221xp5_ASAP7_75t_L g1237 ( .A1(n_949), .A2(n_166), .B1(n_167), .B2(n_168), .C(n_169), .Y(n_1237) );
INVx2_ASAP7_75t_L g1238 ( .A(n_1070), .Y(n_1238) );
BUFx2_ASAP7_75t_L g1239 ( .A(n_1020), .Y(n_1239) );
AND2x2_ASAP7_75t_L g1240 ( .A(n_973), .B(n_167), .Y(n_1240) );
AND2x4_ASAP7_75t_L g1241 ( .A(n_1073), .B(n_168), .Y(n_1241) );
AO21x2_ASAP7_75t_L g1242 ( .A1(n_1080), .A2(n_332), .B(n_418), .Y(n_1242) );
OR2x6_ASAP7_75t_L g1243 ( .A(n_1089), .B(n_169), .Y(n_1243) );
INVx1_ASAP7_75t_L g1244 ( .A(n_1074), .Y(n_1244) );
AND2x2_ASAP7_75t_L g1245 ( .A(n_973), .B(n_170), .Y(n_1245) );
INVx4_ASAP7_75t_L g1246 ( .A(n_1073), .Y(n_1246) );
AOI22xp33_ASAP7_75t_L g1247 ( .A1(n_1024), .A2(n_170), .B1(n_171), .B2(n_173), .Y(n_1247) );
INVxp67_ASAP7_75t_L g1248 ( .A(n_1016), .Y(n_1248) );
AOI21xp5_ASAP7_75t_L g1249 ( .A1(n_1011), .A2(n_334), .B(n_413), .Y(n_1249) );
OAI21xp5_ASAP7_75t_L g1250 ( .A1(n_1074), .A2(n_173), .B(n_174), .Y(n_1250) );
AND2x4_ASAP7_75t_L g1251 ( .A(n_1065), .B(n_174), .Y(n_1251) );
OR2x2_ASAP7_75t_L g1252 ( .A(n_1053), .B(n_175), .Y(n_1252) );
INVx1_ASAP7_75t_L g1253 ( .A(n_1060), .Y(n_1253) );
AOI22xp33_ASAP7_75t_L g1254 ( .A1(n_1006), .A2(n_175), .B1(n_176), .B2(n_177), .Y(n_1254) );
AND2x2_ASAP7_75t_L g1255 ( .A(n_993), .B(n_176), .Y(n_1255) );
INVx5_ASAP7_75t_L g1256 ( .A(n_965), .Y(n_1256) );
AOI222xp33_ASAP7_75t_L g1257 ( .A1(n_1079), .A2(n_177), .B1(n_178), .B2(n_179), .C1(n_180), .C2(n_181), .Y(n_1257) );
AOI21xp5_ASAP7_75t_L g1258 ( .A1(n_1080), .A2(n_343), .B(n_412), .Y(n_1258) );
AOI221xp5_ASAP7_75t_L g1259 ( .A1(n_993), .A2(n_178), .B1(n_179), .B2(n_181), .C(n_182), .Y(n_1259) );
AOI222xp33_ASAP7_75t_L g1260 ( .A1(n_1103), .A2(n_182), .B1(n_183), .B2(n_184), .C1(n_242), .C2(n_245), .Y(n_1260) );
OAI22xp5_ASAP7_75t_L g1261 ( .A1(n_1096), .A2(n_253), .B1(n_256), .B2(n_259), .Y(n_1261) );
OR2x2_ASAP7_75t_L g1262 ( .A(n_1038), .B(n_260), .Y(n_1262) );
OAI22xp33_ASAP7_75t_L g1263 ( .A1(n_1012), .A2(n_261), .B1(n_262), .B2(n_263), .Y(n_1263) );
AOI21xp5_ASAP7_75t_L g1264 ( .A1(n_1078), .A2(n_264), .B(n_266), .Y(n_1264) );
NAND2xp5_ASAP7_75t_L g1265 ( .A(n_982), .B(n_423), .Y(n_1265) );
AOI22xp33_ASAP7_75t_SL g1266 ( .A1(n_1023), .A2(n_269), .B1(n_272), .B2(n_275), .Y(n_1266) );
A2O1A1Ixp33_ASAP7_75t_L g1267 ( .A1(n_1040), .A2(n_276), .B(n_277), .C(n_278), .Y(n_1267) );
CKINVDCx5p33_ASAP7_75t_R g1268 ( .A(n_1065), .Y(n_1268) );
AND2x2_ASAP7_75t_L g1269 ( .A(n_1021), .B(n_280), .Y(n_1269) );
AOI221xp5_ASAP7_75t_L g1270 ( .A1(n_994), .A2(n_950), .B1(n_1012), .B2(n_1002), .C(n_1040), .Y(n_1270) );
HB1xp67_ASAP7_75t_L g1271 ( .A(n_1020), .Y(n_1271) );
OAI22xp5_ASAP7_75t_L g1272 ( .A1(n_1096), .A2(n_288), .B1(n_291), .B2(n_293), .Y(n_1272) );
INVx1_ASAP7_75t_L g1273 ( .A(n_1021), .Y(n_1273) );
AOI22xp33_ASAP7_75t_SL g1274 ( .A1(n_1097), .A2(n_294), .B1(n_295), .B2(n_296), .Y(n_1274) );
BUFx3_ASAP7_75t_L g1275 ( .A(n_1227), .Y(n_1275) );
INVx1_ASAP7_75t_L g1276 ( .A(n_1113), .Y(n_1276) );
NAND2xp5_ASAP7_75t_L g1277 ( .A(n_1107), .B(n_982), .Y(n_1277) );
AND2x2_ASAP7_75t_L g1278 ( .A(n_1127), .B(n_962), .Y(n_1278) );
AOI22xp33_ASAP7_75t_L g1279 ( .A1(n_1106), .A2(n_1015), .B1(n_962), .B2(n_968), .Y(n_1279) );
OR2x2_ASAP7_75t_L g1280 ( .A(n_1219), .B(n_968), .Y(n_1280) );
AND2x2_ASAP7_75t_L g1281 ( .A(n_1240), .B(n_1025), .Y(n_1281) );
HB1xp67_ASAP7_75t_L g1282 ( .A(n_1146), .Y(n_1282) );
AND2x2_ASAP7_75t_L g1283 ( .A(n_1245), .B(n_1025), .Y(n_1283) );
INVx2_ASAP7_75t_L g1284 ( .A(n_1214), .Y(n_1284) );
INVx2_ASAP7_75t_L g1285 ( .A(n_1218), .Y(n_1285) );
HB1xp67_ASAP7_75t_L g1286 ( .A(n_1232), .Y(n_1286) );
AND2x2_ASAP7_75t_L g1287 ( .A(n_1156), .B(n_1028), .Y(n_1287) );
NAND2xp5_ASAP7_75t_L g1288 ( .A(n_1138), .B(n_1015), .Y(n_1288) );
BUFx4f_ASAP7_75t_L g1289 ( .A(n_1243), .Y(n_1289) );
BUFx3_ASAP7_75t_L g1290 ( .A(n_1177), .Y(n_1290) );
INVx1_ASAP7_75t_SL g1291 ( .A(n_1215), .Y(n_1291) );
AND2x2_ASAP7_75t_L g1292 ( .A(n_1203), .B(n_1028), .Y(n_1292) );
INVx2_ASAP7_75t_L g1293 ( .A(n_1224), .Y(n_1293) );
OAI222xp33_ASAP7_75t_L g1294 ( .A1(n_1155), .A2(n_1064), .B1(n_979), .B2(n_1037), .C1(n_1055), .C2(n_1076), .Y(n_1294) );
AND2x2_ASAP7_75t_L g1295 ( .A(n_1210), .B(n_1244), .Y(n_1295) );
INVx1_ASAP7_75t_L g1296 ( .A(n_1189), .Y(n_1296) );
AND2x2_ASAP7_75t_L g1297 ( .A(n_1192), .B(n_971), .Y(n_1297) );
AND2x2_ASAP7_75t_L g1298 ( .A(n_1201), .B(n_971), .Y(n_1298) );
INVx1_ASAP7_75t_L g1299 ( .A(n_1128), .Y(n_1299) );
INVx1_ASAP7_75t_L g1300 ( .A(n_1132), .Y(n_1300) );
HB1xp67_ASAP7_75t_L g1301 ( .A(n_1109), .Y(n_1301) );
INVx1_ASAP7_75t_L g1302 ( .A(n_1157), .Y(n_1302) );
OR2x2_ASAP7_75t_L g1303 ( .A(n_1217), .B(n_955), .Y(n_1303) );
INVxp67_ASAP7_75t_SL g1304 ( .A(n_1199), .Y(n_1304) );
AND2x2_ASAP7_75t_L g1305 ( .A(n_1257), .B(n_1009), .Y(n_1305) );
HB1xp67_ASAP7_75t_L g1306 ( .A(n_1191), .Y(n_1306) );
AND2x2_ASAP7_75t_L g1307 ( .A(n_1257), .B(n_1230), .Y(n_1307) );
INVx1_ASAP7_75t_L g1308 ( .A(n_1251), .Y(n_1308) );
INVx2_ASAP7_75t_SL g1309 ( .A(n_1256), .Y(n_1309) );
INVx2_ASAP7_75t_L g1310 ( .A(n_1238), .Y(n_1310) );
INVx1_ASAP7_75t_L g1311 ( .A(n_1251), .Y(n_1311) );
INVx1_ASAP7_75t_L g1312 ( .A(n_1211), .Y(n_1312) );
INVx1_ASAP7_75t_L g1313 ( .A(n_1114), .Y(n_1313) );
NAND2xp5_ASAP7_75t_L g1314 ( .A(n_1149), .B(n_1061), .Y(n_1314) );
AND2x2_ASAP7_75t_L g1315 ( .A(n_1230), .B(n_1009), .Y(n_1315) );
INVx1_ASAP7_75t_L g1316 ( .A(n_1273), .Y(n_1316) );
INVx1_ASAP7_75t_L g1317 ( .A(n_1148), .Y(n_1317) );
AND2x2_ASAP7_75t_L g1318 ( .A(n_1234), .B(n_1009), .Y(n_1318) );
INVx1_ASAP7_75t_L g1319 ( .A(n_1148), .Y(n_1319) );
BUFx2_ASAP7_75t_L g1320 ( .A(n_1243), .Y(n_1320) );
INVx3_ASAP7_75t_L g1321 ( .A(n_1256), .Y(n_1321) );
INVx1_ASAP7_75t_L g1322 ( .A(n_1253), .Y(n_1322) );
AND2x2_ASAP7_75t_L g1323 ( .A(n_1234), .B(n_1092), .Y(n_1323) );
INVx3_ASAP7_75t_L g1324 ( .A(n_1256), .Y(n_1324) );
AND2x2_ASAP7_75t_L g1325 ( .A(n_1250), .B(n_1092), .Y(n_1325) );
OR2x2_ASAP7_75t_L g1326 ( .A(n_1228), .B(n_1037), .Y(n_1326) );
AND2x2_ASAP7_75t_L g1327 ( .A(n_1250), .B(n_1092), .Y(n_1327) );
INVx1_ASAP7_75t_L g1328 ( .A(n_1235), .Y(n_1328) );
INVx1_ASAP7_75t_L g1329 ( .A(n_1129), .Y(n_1329) );
AND2x2_ASAP7_75t_L g1330 ( .A(n_1243), .B(n_1085), .Y(n_1330) );
NOR2xp67_ASAP7_75t_L g1331 ( .A(n_1180), .B(n_1039), .Y(n_1331) );
INVx1_ASAP7_75t_L g1332 ( .A(n_1129), .Y(n_1332) );
OR2x2_ASAP7_75t_L g1333 ( .A(n_1125), .B(n_999), .Y(n_1333) );
INVx1_ASAP7_75t_L g1334 ( .A(n_1182), .Y(n_1334) );
INVx1_ASAP7_75t_L g1335 ( .A(n_1182), .Y(n_1335) );
INVx1_ASAP7_75t_L g1336 ( .A(n_1181), .Y(n_1336) );
AND2x2_ASAP7_75t_L g1337 ( .A(n_1255), .B(n_1085), .Y(n_1337) );
INVx1_ASAP7_75t_L g1338 ( .A(n_1184), .Y(n_1338) );
AND2x2_ASAP7_75t_L g1339 ( .A(n_1134), .B(n_1085), .Y(n_1339) );
NAND3xp33_ASAP7_75t_SL g1340 ( .A(n_1151), .B(n_1093), .C(n_1076), .Y(n_1340) );
HB1xp67_ASAP7_75t_L g1341 ( .A(n_1268), .Y(n_1341) );
INVx1_ASAP7_75t_L g1342 ( .A(n_1186), .Y(n_1342) );
NOR2x1_ASAP7_75t_L g1343 ( .A(n_1155), .B(n_1101), .Y(n_1343) );
INVx1_ASAP7_75t_L g1344 ( .A(n_1165), .Y(n_1344) );
AOI222xp33_ASAP7_75t_L g1345 ( .A1(n_1231), .A2(n_1071), .B1(n_1063), .B2(n_1043), .C1(n_1013), .C2(n_990), .Y(n_1345) );
NOR2xp67_ASAP7_75t_L g1346 ( .A(n_1246), .B(n_1082), .Y(n_1346) );
AND2x2_ASAP7_75t_L g1347 ( .A(n_1134), .B(n_1095), .Y(n_1347) );
OR2x2_ASAP7_75t_L g1348 ( .A(n_1183), .B(n_1078), .Y(n_1348) );
NAND2xp5_ASAP7_75t_L g1349 ( .A(n_1130), .B(n_1104), .Y(n_1349) );
INVx1_ASAP7_75t_L g1350 ( .A(n_1118), .Y(n_1350) );
NAND2xp5_ASAP7_75t_L g1351 ( .A(n_1252), .B(n_991), .Y(n_1351) );
INVx2_ASAP7_75t_R g1352 ( .A(n_1256), .Y(n_1352) );
AND2x2_ASAP7_75t_L g1353 ( .A(n_1139), .B(n_1071), .Y(n_1353) );
INVxp67_ASAP7_75t_L g1354 ( .A(n_1145), .Y(n_1354) );
INVx1_ASAP7_75t_L g1355 ( .A(n_1123), .Y(n_1355) );
HB1xp67_ASAP7_75t_L g1356 ( .A(n_1150), .Y(n_1356) );
AND2x2_ASAP7_75t_L g1357 ( .A(n_1139), .B(n_964), .Y(n_1357) );
AND2x2_ASAP7_75t_L g1358 ( .A(n_1112), .B(n_967), .Y(n_1358) );
INVx1_ASAP7_75t_L g1359 ( .A(n_1196), .Y(n_1359) );
INVx2_ASAP7_75t_L g1360 ( .A(n_1223), .Y(n_1360) );
OR2x2_ASAP7_75t_L g1361 ( .A(n_1215), .B(n_1055), .Y(n_1361) );
INVx1_ASAP7_75t_L g1362 ( .A(n_1241), .Y(n_1362) );
BUFx2_ASAP7_75t_L g1363 ( .A(n_1108), .Y(n_1363) );
INVx1_ASAP7_75t_L g1364 ( .A(n_1241), .Y(n_1364) );
INVx1_ASAP7_75t_L g1365 ( .A(n_1162), .Y(n_1365) );
INVx4_ASAP7_75t_L g1366 ( .A(n_1205), .Y(n_1366) );
BUFx12f_ASAP7_75t_L g1367 ( .A(n_1220), .Y(n_1367) );
AND2x2_ASAP7_75t_L g1368 ( .A(n_1112), .B(n_967), .Y(n_1368) );
HB1xp67_ASAP7_75t_L g1369 ( .A(n_1168), .Y(n_1369) );
INVx1_ASAP7_75t_L g1370 ( .A(n_1162), .Y(n_1370) );
INVx2_ASAP7_75t_L g1371 ( .A(n_1223), .Y(n_1371) );
NAND2xp5_ASAP7_75t_L g1372 ( .A(n_1115), .B(n_983), .Y(n_1372) );
AND2x2_ASAP7_75t_L g1373 ( .A(n_1151), .B(n_1029), .Y(n_1373) );
NAND2xp5_ASAP7_75t_L g1374 ( .A(n_1120), .B(n_1083), .Y(n_1374) );
AND2x2_ASAP7_75t_L g1375 ( .A(n_1173), .B(n_965), .Y(n_1375) );
AND2x2_ASAP7_75t_L g1376 ( .A(n_1173), .B(n_965), .Y(n_1376) );
AND2x4_ASAP7_75t_L g1377 ( .A(n_1205), .B(n_1101), .Y(n_1377) );
INVx1_ASAP7_75t_L g1378 ( .A(n_1229), .Y(n_1378) );
INVx1_ASAP7_75t_L g1379 ( .A(n_1117), .Y(n_1379) );
AND2x2_ASAP7_75t_L g1380 ( .A(n_1271), .B(n_977), .Y(n_1380) );
AND2x2_ASAP7_75t_L g1381 ( .A(n_1260), .B(n_977), .Y(n_1381) );
INVx1_ASAP7_75t_L g1382 ( .A(n_1117), .Y(n_1382) );
OR2x2_ASAP7_75t_L g1383 ( .A(n_1207), .B(n_977), .Y(n_1383) );
BUFx2_ASAP7_75t_L g1384 ( .A(n_1110), .Y(n_1384) );
INVx1_ASAP7_75t_L g1385 ( .A(n_1135), .Y(n_1385) );
AND2x2_ASAP7_75t_L g1386 ( .A(n_1260), .B(n_1088), .Y(n_1386) );
INVx1_ASAP7_75t_L g1387 ( .A(n_1135), .Y(n_1387) );
INVx1_ASAP7_75t_L g1388 ( .A(n_1225), .Y(n_1388) );
NAND2xp5_ASAP7_75t_L g1389 ( .A(n_1226), .B(n_1042), .Y(n_1389) );
INVx1_ASAP7_75t_L g1390 ( .A(n_1194), .Y(n_1390) );
HB1xp67_ASAP7_75t_L g1391 ( .A(n_1233), .Y(n_1391) );
INVx1_ASAP7_75t_L g1392 ( .A(n_1208), .Y(n_1392) );
INVx1_ASAP7_75t_L g1393 ( .A(n_1197), .Y(n_1393) );
INVx1_ASAP7_75t_L g1394 ( .A(n_1242), .Y(n_1394) );
INVx1_ASAP7_75t_L g1395 ( .A(n_1242), .Y(n_1395) );
INVx1_ASAP7_75t_L g1396 ( .A(n_1269), .Y(n_1396) );
INVxp67_ASAP7_75t_L g1397 ( .A(n_1222), .Y(n_1397) );
INVx1_ASAP7_75t_L g1398 ( .A(n_1198), .Y(n_1398) );
AND2x2_ASAP7_75t_L g1399 ( .A(n_1239), .B(n_1088), .Y(n_1399) );
AND2x2_ASAP7_75t_L g1400 ( .A(n_1206), .B(n_1088), .Y(n_1400) );
INVx3_ASAP7_75t_L g1401 ( .A(n_1246), .Y(n_1401) );
NAND2xp5_ASAP7_75t_L g1402 ( .A(n_1179), .B(n_945), .Y(n_1402) );
OR2x2_ASAP7_75t_L g1403 ( .A(n_1209), .B(n_1094), .Y(n_1403) );
HB1xp67_ASAP7_75t_L g1404 ( .A(n_1124), .Y(n_1404) );
NAND2xp5_ASAP7_75t_L g1405 ( .A(n_1185), .B(n_1090), .Y(n_1405) );
AND2x2_ASAP7_75t_L g1406 ( .A(n_1247), .B(n_1094), .Y(n_1406) );
INVxp67_ASAP7_75t_L g1407 ( .A(n_1144), .Y(n_1407) );
INVx2_ASAP7_75t_L g1408 ( .A(n_1265), .Y(n_1408) );
AND2x2_ASAP7_75t_L g1409 ( .A(n_1143), .B(n_1094), .Y(n_1409) );
AND2x2_ASAP7_75t_L g1410 ( .A(n_1172), .B(n_1102), .Y(n_1410) );
HB1xp67_ASAP7_75t_L g1411 ( .A(n_1204), .Y(n_1411) );
AND2x4_ASAP7_75t_L g1412 ( .A(n_1131), .B(n_1100), .Y(n_1412) );
INVx1_ASAP7_75t_L g1413 ( .A(n_1213), .Y(n_1413) );
INVx2_ASAP7_75t_L g1414 ( .A(n_1262), .Y(n_1414) );
NAND2xp5_ASAP7_75t_L g1415 ( .A(n_1142), .B(n_1031), .Y(n_1415) );
AND2x2_ASAP7_75t_L g1416 ( .A(n_1176), .B(n_1105), .Y(n_1416) );
CKINVDCx6p67_ASAP7_75t_R g1417 ( .A(n_1216), .Y(n_1417) );
OR2x2_ASAP7_75t_L g1418 ( .A(n_1144), .B(n_1059), .Y(n_1418) );
INVx2_ASAP7_75t_L g1419 ( .A(n_1111), .Y(n_1419) );
AO21x2_ASAP7_75t_L g1420 ( .A1(n_1264), .A2(n_1087), .B(n_1030), .Y(n_1420) );
AND2x4_ASAP7_75t_L g1421 ( .A(n_1131), .B(n_297), .Y(n_1421) );
NAND4xp25_ASAP7_75t_L g1422 ( .A(n_1147), .B(n_1030), .C(n_299), .D(n_300), .Y(n_1422) );
INVx1_ASAP7_75t_L g1423 ( .A(n_1193), .Y(n_1423) );
INVx2_ASAP7_75t_L g1424 ( .A(n_1261), .Y(n_1424) );
NAND2xp5_ASAP7_75t_L g1425 ( .A(n_1359), .B(n_1140), .Y(n_1425) );
OR2x2_ASAP7_75t_L g1426 ( .A(n_1328), .B(n_1164), .Y(n_1426) );
OR2x6_ASAP7_75t_L g1427 ( .A(n_1320), .B(n_1261), .Y(n_1427) );
INVx4_ASAP7_75t_L g1428 ( .A(n_1289), .Y(n_1428) );
NOR2xp33_ASAP7_75t_L g1429 ( .A(n_1397), .B(n_1221), .Y(n_1429) );
INVx3_ASAP7_75t_L g1430 ( .A(n_1377), .Y(n_1430) );
AOI221xp5_ASAP7_75t_L g1431 ( .A1(n_1388), .A2(n_1178), .B1(n_1188), .B2(n_1137), .C(n_1166), .Y(n_1431) );
INVxp67_ASAP7_75t_L g1432 ( .A(n_1282), .Y(n_1432) );
INVx1_ASAP7_75t_L g1433 ( .A(n_1276), .Y(n_1433) );
NAND2xp5_ASAP7_75t_L g1434 ( .A(n_1295), .B(n_1301), .Y(n_1434) );
AND2x4_ASAP7_75t_L g1435 ( .A(n_1322), .B(n_1258), .Y(n_1435) );
AND2x2_ASAP7_75t_L g1436 ( .A(n_1337), .B(n_1187), .Y(n_1436) );
INVx2_ASAP7_75t_L g1437 ( .A(n_1284), .Y(n_1437) );
INVx1_ASAP7_75t_SL g1438 ( .A(n_1290), .Y(n_1438) );
INVxp67_ASAP7_75t_SL g1439 ( .A(n_1289), .Y(n_1439) );
NAND2xp5_ASAP7_75t_L g1440 ( .A(n_1295), .B(n_1159), .Y(n_1440) );
INVx2_ASAP7_75t_L g1441 ( .A(n_1284), .Y(n_1441) );
HB1xp67_ASAP7_75t_L g1442 ( .A(n_1361), .Y(n_1442) );
NAND2xp5_ASAP7_75t_L g1443 ( .A(n_1407), .B(n_1169), .Y(n_1443) );
AND2x4_ASAP7_75t_L g1444 ( .A(n_1322), .B(n_1190), .Y(n_1444) );
NAND2xp5_ASAP7_75t_L g1445 ( .A(n_1296), .B(n_1153), .Y(n_1445) );
OR2x2_ASAP7_75t_L g1446 ( .A(n_1328), .B(n_1119), .Y(n_1446) );
HB1xp67_ASAP7_75t_L g1447 ( .A(n_1361), .Y(n_1447) );
AND2x2_ASAP7_75t_L g1448 ( .A(n_1337), .B(n_1141), .Y(n_1448) );
AND3x2_ASAP7_75t_L g1449 ( .A(n_1404), .B(n_1248), .C(n_1158), .Y(n_1449) );
AOI22xp5_ASAP7_75t_L g1450 ( .A1(n_1307), .A2(n_1122), .B1(n_1136), .B2(n_1126), .Y(n_1450) );
OR2x2_ASAP7_75t_L g1451 ( .A(n_1285), .B(n_1133), .Y(n_1451) );
INVx1_ASAP7_75t_L g1452 ( .A(n_1299), .Y(n_1452) );
AOI22xp33_ASAP7_75t_L g1453 ( .A1(n_1307), .A2(n_1160), .B1(n_1195), .B2(n_1237), .Y(n_1453) );
INVx4_ASAP7_75t_L g1454 ( .A(n_1289), .Y(n_1454) );
NAND2xp5_ASAP7_75t_L g1455 ( .A(n_1302), .B(n_1171), .Y(n_1455) );
BUFx3_ASAP7_75t_L g1456 ( .A(n_1290), .Y(n_1456) );
AND2x2_ASAP7_75t_L g1457 ( .A(n_1297), .B(n_1254), .Y(n_1457) );
NAND2x1_ASAP7_75t_L g1458 ( .A(n_1401), .B(n_1121), .Y(n_1458) );
AND2x2_ASAP7_75t_L g1459 ( .A(n_1297), .B(n_1175), .Y(n_1459) );
INVx1_ASAP7_75t_L g1460 ( .A(n_1300), .Y(n_1460) );
INVx2_ASAP7_75t_L g1461 ( .A(n_1285), .Y(n_1461) );
OR2x2_ASAP7_75t_L g1462 ( .A(n_1365), .B(n_1202), .Y(n_1462) );
NAND2xp5_ASAP7_75t_L g1463 ( .A(n_1313), .B(n_1170), .Y(n_1463) );
AND2x2_ASAP7_75t_L g1464 ( .A(n_1318), .B(n_1200), .Y(n_1464) );
NOR2x1_ASAP7_75t_L g1465 ( .A(n_1401), .B(n_1263), .Y(n_1465) );
NAND2xp5_ASAP7_75t_L g1466 ( .A(n_1338), .B(n_1152), .Y(n_1466) );
INVx2_ASAP7_75t_L g1467 ( .A(n_1316), .Y(n_1467) );
INVx1_ASAP7_75t_L g1468 ( .A(n_1314), .Y(n_1468) );
HB1xp67_ASAP7_75t_L g1469 ( .A(n_1291), .Y(n_1469) );
AND2x2_ASAP7_75t_L g1470 ( .A(n_1318), .B(n_1259), .Y(n_1470) );
OR2x2_ASAP7_75t_L g1471 ( .A(n_1370), .B(n_1116), .Y(n_1471) );
AND2x2_ASAP7_75t_L g1472 ( .A(n_1298), .B(n_1270), .Y(n_1472) );
AND2x2_ASAP7_75t_L g1473 ( .A(n_1298), .B(n_1274), .Y(n_1473) );
AND2x2_ASAP7_75t_L g1474 ( .A(n_1316), .B(n_1266), .Y(n_1474) );
INVx1_ASAP7_75t_L g1475 ( .A(n_1342), .Y(n_1475) );
INVx2_ASAP7_75t_SL g1476 ( .A(n_1401), .Y(n_1476) );
NAND2xp5_ASAP7_75t_L g1477 ( .A(n_1393), .B(n_1174), .Y(n_1477) );
INVx3_ASAP7_75t_L g1478 ( .A(n_1377), .Y(n_1478) );
AOI22xp33_ASAP7_75t_L g1479 ( .A1(n_1373), .A2(n_1272), .B1(n_1154), .B2(n_1249), .Y(n_1479) );
INVx1_ASAP7_75t_L g1480 ( .A(n_1288), .Y(n_1480) );
AND2x4_ASAP7_75t_L g1481 ( .A(n_1330), .B(n_1163), .Y(n_1481) );
AND2x2_ASAP7_75t_L g1482 ( .A(n_1323), .B(n_1267), .Y(n_1482) );
INVxp67_ASAP7_75t_SL g1483 ( .A(n_1320), .Y(n_1483) );
INVx4_ASAP7_75t_L g1484 ( .A(n_1366), .Y(n_1484) );
INVx2_ASAP7_75t_L g1485 ( .A(n_1293), .Y(n_1485) );
INVx2_ASAP7_75t_L g1486 ( .A(n_1293), .Y(n_1486) );
INVx2_ASAP7_75t_L g1487 ( .A(n_1310), .Y(n_1487) );
CKINVDCx5p33_ASAP7_75t_R g1488 ( .A(n_1417), .Y(n_1488) );
INVx1_ASAP7_75t_L g1489 ( .A(n_1312), .Y(n_1489) );
AND2x2_ASAP7_75t_L g1490 ( .A(n_1323), .B(n_1167), .Y(n_1490) );
HB1xp67_ASAP7_75t_L g1491 ( .A(n_1391), .Y(n_1491) );
AND2x2_ASAP7_75t_L g1492 ( .A(n_1325), .B(n_1212), .Y(n_1492) );
AND2x2_ASAP7_75t_L g1493 ( .A(n_1325), .B(n_1236), .Y(n_1493) );
INVx1_ASAP7_75t_L g1494 ( .A(n_1362), .Y(n_1494) );
INVx1_ASAP7_75t_L g1495 ( .A(n_1364), .Y(n_1495) );
OAI21x1_ASAP7_75t_L g1496 ( .A1(n_1360), .A2(n_1161), .B(n_301), .Y(n_1496) );
BUFx3_ASAP7_75t_L g1497 ( .A(n_1321), .Y(n_1497) );
BUFx2_ASAP7_75t_L g1498 ( .A(n_1321), .Y(n_1498) );
AND2x2_ASAP7_75t_L g1499 ( .A(n_1327), .B(n_298), .Y(n_1499) );
OAI31xp33_ASAP7_75t_L g1500 ( .A1(n_1398), .A2(n_305), .A3(n_311), .B(n_315), .Y(n_1500) );
HB1xp67_ASAP7_75t_L g1501 ( .A(n_1356), .Y(n_1501) );
NAND2xp5_ASAP7_75t_L g1502 ( .A(n_1306), .B(n_411), .Y(n_1502) );
INVx2_ASAP7_75t_L g1503 ( .A(n_1310), .Y(n_1503) );
OAI22xp5_ASAP7_75t_L g1504 ( .A1(n_1373), .A2(n_318), .B1(n_320), .B2(n_321), .Y(n_1504) );
INVx1_ASAP7_75t_L g1505 ( .A(n_1336), .Y(n_1505) );
AND2x2_ASAP7_75t_L g1506 ( .A(n_1327), .B(n_323), .Y(n_1506) );
BUFx2_ASAP7_75t_L g1507 ( .A(n_1330), .Y(n_1507) );
BUFx3_ASAP7_75t_L g1508 ( .A(n_1321), .Y(n_1508) );
CKINVDCx20_ASAP7_75t_R g1509 ( .A(n_1417), .Y(n_1509) );
INVx1_ASAP7_75t_L g1510 ( .A(n_1308), .Y(n_1510) );
NAND2xp5_ASAP7_75t_L g1511 ( .A(n_1369), .B(n_324), .Y(n_1511) );
AND2x2_ASAP7_75t_L g1512 ( .A(n_1339), .B(n_337), .Y(n_1512) );
AOI22xp33_ASAP7_75t_L g1513 ( .A1(n_1413), .A2(n_339), .B1(n_344), .B2(n_347), .Y(n_1513) );
INVx1_ASAP7_75t_L g1514 ( .A(n_1311), .Y(n_1514) );
INVx2_ASAP7_75t_L g1515 ( .A(n_1287), .Y(n_1515) );
OAI31xp33_ASAP7_75t_L g1516 ( .A1(n_1378), .A2(n_349), .A3(n_350), .B(n_351), .Y(n_1516) );
AND2x2_ASAP7_75t_L g1517 ( .A(n_1339), .B(n_354), .Y(n_1517) );
NAND2xp5_ASAP7_75t_L g1518 ( .A(n_1277), .B(n_410), .Y(n_1518) );
HB1xp67_ASAP7_75t_L g1519 ( .A(n_1304), .Y(n_1519) );
OAI221xp5_ASAP7_75t_L g1520 ( .A1(n_1354), .A2(n_355), .B1(n_356), .B2(n_357), .C(n_359), .Y(n_1520) );
OAI22xp5_ASAP7_75t_L g1521 ( .A1(n_1333), .A2(n_361), .B1(n_364), .B2(n_365), .Y(n_1521) );
INVx2_ASAP7_75t_L g1522 ( .A(n_1287), .Y(n_1522) );
INVx1_ASAP7_75t_L g1523 ( .A(n_1278), .Y(n_1523) );
AND2x2_ASAP7_75t_L g1524 ( .A(n_1281), .B(n_367), .Y(n_1524) );
AND2x2_ASAP7_75t_L g1525 ( .A(n_1281), .B(n_369), .Y(n_1525) );
NOR2x1_ASAP7_75t_SL g1526 ( .A(n_1366), .B(n_371), .Y(n_1526) );
AND2x2_ASAP7_75t_L g1527 ( .A(n_1283), .B(n_372), .Y(n_1527) );
BUFx2_ASAP7_75t_L g1528 ( .A(n_1377), .Y(n_1528) );
INVx2_ASAP7_75t_L g1529 ( .A(n_1292), .Y(n_1529) );
INVx1_ASAP7_75t_SL g1530 ( .A(n_1275), .Y(n_1530) );
INVxp67_ASAP7_75t_SL g1531 ( .A(n_1348), .Y(n_1531) );
INVx1_ASAP7_75t_L g1532 ( .A(n_1278), .Y(n_1532) );
INVxp67_ASAP7_75t_L g1533 ( .A(n_1341), .Y(n_1533) );
NAND2x1p5_ASAP7_75t_L g1534 ( .A(n_1366), .B(n_373), .Y(n_1534) );
OAI33xp33_ASAP7_75t_L g1535 ( .A1(n_1423), .A2(n_377), .A3(n_378), .B1(n_379), .B2(n_380), .B3(n_381), .Y(n_1535) );
NAND2xp5_ASAP7_75t_L g1536 ( .A(n_1350), .B(n_383), .Y(n_1536) );
AND2x2_ASAP7_75t_L g1537 ( .A(n_1283), .B(n_384), .Y(n_1537) );
AND2x2_ASAP7_75t_SL g1538 ( .A(n_1375), .B(n_386), .Y(n_1538) );
AND2x2_ASAP7_75t_L g1539 ( .A(n_1396), .B(n_388), .Y(n_1539) );
INVx1_ASAP7_75t_SL g1540 ( .A(n_1275), .Y(n_1540) );
AND2x2_ASAP7_75t_SL g1541 ( .A(n_1375), .B(n_389), .Y(n_1541) );
AND2x2_ASAP7_75t_L g1542 ( .A(n_1396), .B(n_390), .Y(n_1542) );
NAND2x1p5_ASAP7_75t_L g1543 ( .A(n_1324), .B(n_391), .Y(n_1543) );
INVx2_ASAP7_75t_L g1544 ( .A(n_1292), .Y(n_1544) );
INVx2_ASAP7_75t_SL g1545 ( .A(n_1324), .Y(n_1545) );
INVx1_ASAP7_75t_L g1546 ( .A(n_1280), .Y(n_1546) );
AO21x2_ASAP7_75t_L g1547 ( .A1(n_1394), .A2(n_392), .B(n_393), .Y(n_1547) );
INVx2_ASAP7_75t_L g1548 ( .A(n_1371), .Y(n_1548) );
BUFx2_ASAP7_75t_L g1549 ( .A(n_1324), .Y(n_1549) );
INVx3_ASAP7_75t_L g1550 ( .A(n_1412), .Y(n_1550) );
AND2x2_ASAP7_75t_L g1551 ( .A(n_1434), .B(n_1353), .Y(n_1551) );
AND2x2_ASAP7_75t_L g1552 ( .A(n_1436), .B(n_1353), .Y(n_1552) );
OR2x2_ASAP7_75t_L g1553 ( .A(n_1519), .B(n_1348), .Y(n_1553) );
NOR2x1_ASAP7_75t_L g1554 ( .A(n_1509), .B(n_1346), .Y(n_1554) );
INVx1_ASAP7_75t_L g1555 ( .A(n_1433), .Y(n_1555) );
AND2x2_ASAP7_75t_L g1556 ( .A(n_1436), .B(n_1347), .Y(n_1556) );
OR2x2_ASAP7_75t_L g1557 ( .A(n_1491), .B(n_1280), .Y(n_1557) );
NAND2xp5_ASAP7_75t_L g1558 ( .A(n_1546), .B(n_1379), .Y(n_1558) );
OR2x2_ASAP7_75t_L g1559 ( .A(n_1501), .B(n_1303), .Y(n_1559) );
CKINVDCx5p33_ASAP7_75t_R g1560 ( .A(n_1509), .Y(n_1560) );
NAND2xp5_ASAP7_75t_L g1561 ( .A(n_1472), .B(n_1382), .Y(n_1561) );
NOR2xp33_ASAP7_75t_L g1562 ( .A(n_1438), .B(n_1286), .Y(n_1562) );
INVx1_ASAP7_75t_L g1563 ( .A(n_1452), .Y(n_1563) );
AND2x2_ASAP7_75t_L g1564 ( .A(n_1456), .B(n_1347), .Y(n_1564) );
INVx1_ASAP7_75t_L g1565 ( .A(n_1460), .Y(n_1565) );
INVx1_ASAP7_75t_L g1566 ( .A(n_1505), .Y(n_1566) );
NAND2xp5_ASAP7_75t_L g1567 ( .A(n_1468), .B(n_1385), .Y(n_1567) );
NOR2xp67_ASAP7_75t_L g1568 ( .A(n_1484), .B(n_1309), .Y(n_1568) );
INVx1_ASAP7_75t_L g1569 ( .A(n_1475), .Y(n_1569) );
CKINVDCx5p33_ASAP7_75t_R g1570 ( .A(n_1488), .Y(n_1570) );
NAND2xp5_ASAP7_75t_L g1571 ( .A(n_1472), .B(n_1387), .Y(n_1571) );
OR2x2_ASAP7_75t_L g1572 ( .A(n_1442), .B(n_1303), .Y(n_1572) );
AND2x4_ASAP7_75t_L g1573 ( .A(n_1483), .B(n_1403), .Y(n_1573) );
AND2x2_ASAP7_75t_L g1574 ( .A(n_1456), .B(n_1380), .Y(n_1574) );
INVx3_ASAP7_75t_L g1575 ( .A(n_1484), .Y(n_1575) );
NAND2xp5_ASAP7_75t_L g1576 ( .A(n_1523), .B(n_1317), .Y(n_1576) );
INVxp67_ASAP7_75t_L g1577 ( .A(n_1469), .Y(n_1577) );
HB1xp67_ASAP7_75t_L g1578 ( .A(n_1447), .Y(n_1578) );
AND2x2_ASAP7_75t_L g1579 ( .A(n_1507), .B(n_1380), .Y(n_1579) );
NOR2xp33_ASAP7_75t_R g1580 ( .A(n_1488), .B(n_1367), .Y(n_1580) );
INVx2_ASAP7_75t_L g1581 ( .A(n_1437), .Y(n_1581) );
INVx1_ASAP7_75t_L g1582 ( .A(n_1489), .Y(n_1582) );
NAND2xp5_ASAP7_75t_L g1583 ( .A(n_1532), .B(n_1317), .Y(n_1583) );
AND2x2_ASAP7_75t_L g1584 ( .A(n_1507), .B(n_1399), .Y(n_1584) );
OR2x6_ASAP7_75t_L g1585 ( .A(n_1427), .B(n_1376), .Y(n_1585) );
OR2x2_ASAP7_75t_L g1586 ( .A(n_1432), .B(n_1333), .Y(n_1586) );
NAND2xp5_ASAP7_75t_L g1587 ( .A(n_1510), .B(n_1305), .Y(n_1587) );
INVxp67_ASAP7_75t_L g1588 ( .A(n_1498), .Y(n_1588) );
NAND2xp5_ASAP7_75t_L g1589 ( .A(n_1467), .B(n_1319), .Y(n_1589) );
INVx2_ASAP7_75t_L g1590 ( .A(n_1437), .Y(n_1590) );
INVx1_ASAP7_75t_L g1591 ( .A(n_1467), .Y(n_1591) );
INVx3_ASAP7_75t_L g1592 ( .A(n_1484), .Y(n_1592) );
AOI22xp33_ASAP7_75t_L g1593 ( .A1(n_1427), .A2(n_1305), .B1(n_1381), .B2(n_1386), .Y(n_1593) );
INVxp67_ASAP7_75t_SL g1594 ( .A(n_1531), .Y(n_1594) );
NAND2xp5_ASAP7_75t_L g1595 ( .A(n_1480), .B(n_1319), .Y(n_1595) );
INVx2_ASAP7_75t_L g1596 ( .A(n_1441), .Y(n_1596) );
AOI22xp5_ASAP7_75t_L g1597 ( .A1(n_1450), .A2(n_1381), .B1(n_1386), .B2(n_1358), .Y(n_1597) );
AND2x2_ASAP7_75t_L g1598 ( .A(n_1549), .B(n_1399), .Y(n_1598) );
INVx2_ASAP7_75t_SL g1599 ( .A(n_1497), .Y(n_1599) );
HB1xp67_ASAP7_75t_L g1600 ( .A(n_1476), .Y(n_1600) );
INVx1_ASAP7_75t_L g1601 ( .A(n_1494), .Y(n_1601) );
AND2x2_ASAP7_75t_L g1602 ( .A(n_1512), .B(n_1376), .Y(n_1602) );
OR2x2_ASAP7_75t_L g1603 ( .A(n_1515), .B(n_1403), .Y(n_1603) );
NOR2xp33_ASAP7_75t_L g1604 ( .A(n_1530), .B(n_1367), .Y(n_1604) );
AOI221xp5_ASAP7_75t_L g1605 ( .A1(n_1425), .A2(n_1355), .B1(n_1344), .B2(n_1340), .C(n_1374), .Y(n_1605) );
OR2x2_ASAP7_75t_L g1606 ( .A(n_1515), .B(n_1383), .Y(n_1606) );
NAND2xp5_ASAP7_75t_L g1607 ( .A(n_1457), .B(n_1315), .Y(n_1607) );
INVx1_ASAP7_75t_L g1608 ( .A(n_1495), .Y(n_1608) );
OR2x2_ASAP7_75t_L g1609 ( .A(n_1522), .B(n_1383), .Y(n_1609) );
INVxp67_ASAP7_75t_L g1610 ( .A(n_1429), .Y(n_1610) );
OR2x2_ASAP7_75t_L g1611 ( .A(n_1522), .B(n_1414), .Y(n_1611) );
OR2x2_ASAP7_75t_L g1612 ( .A(n_1529), .B(n_1414), .Y(n_1612) );
OR2x2_ASAP7_75t_L g1613 ( .A(n_1529), .B(n_1372), .Y(n_1613) );
NAND2xp5_ASAP7_75t_L g1614 ( .A(n_1457), .B(n_1315), .Y(n_1614) );
AND2x4_ASAP7_75t_L g1615 ( .A(n_1430), .B(n_1363), .Y(n_1615) );
INVxp67_ASAP7_75t_SL g1616 ( .A(n_1476), .Y(n_1616) );
OR2x2_ASAP7_75t_L g1617 ( .A(n_1544), .B(n_1418), .Y(n_1617) );
INVx1_ASAP7_75t_L g1618 ( .A(n_1514), .Y(n_1618) );
AND2x4_ASAP7_75t_L g1619 ( .A(n_1430), .B(n_1363), .Y(n_1619) );
NAND2xp5_ASAP7_75t_L g1620 ( .A(n_1544), .B(n_1424), .Y(n_1620) );
INVx2_ASAP7_75t_L g1621 ( .A(n_1461), .Y(n_1621) );
INVx1_ASAP7_75t_L g1622 ( .A(n_1461), .Y(n_1622) );
INVx1_ASAP7_75t_SL g1623 ( .A(n_1497), .Y(n_1623) );
INVx1_ASAP7_75t_L g1624 ( .A(n_1485), .Y(n_1624) );
AND2x2_ASAP7_75t_L g1625 ( .A(n_1512), .B(n_1357), .Y(n_1625) );
AND2x2_ASAP7_75t_L g1626 ( .A(n_1517), .B(n_1357), .Y(n_1626) );
OAI33xp33_ASAP7_75t_L g1627 ( .A1(n_1533), .A2(n_1349), .A3(n_1392), .B1(n_1390), .B2(n_1326), .B3(n_1418), .Y(n_1627) );
INVx1_ASAP7_75t_L g1628 ( .A(n_1486), .Y(n_1628) );
AOI22xp33_ASAP7_75t_SL g1629 ( .A1(n_1538), .A2(n_1358), .B1(n_1368), .B2(n_1400), .Y(n_1629) );
AND2x2_ASAP7_75t_L g1630 ( .A(n_1517), .B(n_1524), .Y(n_1630) );
INVx1_ASAP7_75t_L g1631 ( .A(n_1486), .Y(n_1631) );
NAND2xp5_ASAP7_75t_L g1632 ( .A(n_1459), .B(n_1424), .Y(n_1632) );
OAI22xp5_ASAP7_75t_L g1633 ( .A1(n_1538), .A2(n_1368), .B1(n_1279), .B2(n_1351), .Y(n_1633) );
AOI21xp5_ASAP7_75t_L g1634 ( .A1(n_1541), .A2(n_1343), .B(n_1405), .Y(n_1634) );
AND2x2_ASAP7_75t_L g1635 ( .A(n_1524), .B(n_1309), .Y(n_1635) );
INVx5_ASAP7_75t_L g1636 ( .A(n_1428), .Y(n_1636) );
INVx2_ASAP7_75t_SL g1637 ( .A(n_1508), .Y(n_1637) );
AND2x2_ASAP7_75t_L g1638 ( .A(n_1525), .B(n_1400), .Y(n_1638) );
INVx1_ASAP7_75t_L g1639 ( .A(n_1487), .Y(n_1639) );
HB1xp67_ASAP7_75t_L g1640 ( .A(n_1508), .Y(n_1640) );
AOI22xp5_ASAP7_75t_L g1641 ( .A1(n_1453), .A2(n_1422), .B1(n_1406), .B2(n_1409), .Y(n_1641) );
NAND2xp33_ASAP7_75t_L g1642 ( .A(n_1534), .B(n_1411), .Y(n_1642) );
INVx1_ASAP7_75t_L g1643 ( .A(n_1487), .Y(n_1643) );
NAND2xp5_ASAP7_75t_L g1644 ( .A(n_1459), .B(n_1448), .Y(n_1644) );
NAND3xp33_ASAP7_75t_L g1645 ( .A(n_1449), .B(n_1345), .C(n_1329), .Y(n_1645) );
INVx1_ASAP7_75t_L g1646 ( .A(n_1503), .Y(n_1646) );
INVx1_ASAP7_75t_L g1647 ( .A(n_1503), .Y(n_1647) );
AND2x2_ASAP7_75t_L g1648 ( .A(n_1552), .B(n_1550), .Y(n_1648) );
NAND2xp5_ASAP7_75t_SL g1649 ( .A(n_1575), .B(n_1541), .Y(n_1649) );
AND2x2_ASAP7_75t_L g1650 ( .A(n_1585), .B(n_1550), .Y(n_1650) );
INVx1_ASAP7_75t_L g1651 ( .A(n_1555), .Y(n_1651) );
OR2x2_ASAP7_75t_L g1652 ( .A(n_1553), .B(n_1448), .Y(n_1652) );
OR2x2_ASAP7_75t_L g1653 ( .A(n_1557), .B(n_1550), .Y(n_1653) );
AND2x2_ASAP7_75t_L g1654 ( .A(n_1585), .B(n_1528), .Y(n_1654) );
INVx1_ASAP7_75t_L g1655 ( .A(n_1563), .Y(n_1655) );
OR2x2_ASAP7_75t_L g1656 ( .A(n_1559), .B(n_1528), .Y(n_1656) );
NAND2xp5_ASAP7_75t_L g1657 ( .A(n_1644), .B(n_1464), .Y(n_1657) );
AND2x2_ASAP7_75t_L g1658 ( .A(n_1585), .B(n_1490), .Y(n_1658) );
INVx1_ASAP7_75t_L g1659 ( .A(n_1565), .Y(n_1659) );
AND2x2_ASAP7_75t_L g1660 ( .A(n_1625), .B(n_1490), .Y(n_1660) );
NOR2xp33_ASAP7_75t_L g1661 ( .A(n_1610), .B(n_1540), .Y(n_1661) );
AND2x2_ASAP7_75t_L g1662 ( .A(n_1626), .B(n_1492), .Y(n_1662) );
AND2x2_ASAP7_75t_L g1663 ( .A(n_1632), .B(n_1492), .Y(n_1663) );
INVx1_ASAP7_75t_L g1664 ( .A(n_1566), .Y(n_1664) );
OR2x2_ASAP7_75t_L g1665 ( .A(n_1606), .B(n_1430), .Y(n_1665) );
NAND2xp5_ASAP7_75t_L g1666 ( .A(n_1644), .B(n_1464), .Y(n_1666) );
INVx1_ASAP7_75t_L g1667 ( .A(n_1569), .Y(n_1667) );
AND2x2_ASAP7_75t_L g1668 ( .A(n_1632), .B(n_1493), .Y(n_1668) );
NAND2xp5_ASAP7_75t_L g1669 ( .A(n_1561), .B(n_1470), .Y(n_1669) );
INVx2_ASAP7_75t_L g1670 ( .A(n_1591), .Y(n_1670) );
HB1xp67_ASAP7_75t_L g1671 ( .A(n_1594), .Y(n_1671) );
NOR2xp33_ASAP7_75t_L g1672 ( .A(n_1560), .B(n_1428), .Y(n_1672) );
INVx1_ASAP7_75t_L g1673 ( .A(n_1582), .Y(n_1673) );
INVx2_ASAP7_75t_L g1674 ( .A(n_1581), .Y(n_1674) );
NAND2xp33_ASAP7_75t_L g1675 ( .A(n_1554), .B(n_1636), .Y(n_1675) );
AND2x2_ASAP7_75t_L g1676 ( .A(n_1551), .B(n_1493), .Y(n_1676) );
OR2x2_ASAP7_75t_L g1677 ( .A(n_1586), .B(n_1446), .Y(n_1677) );
NAND2xp5_ASAP7_75t_L g1678 ( .A(n_1561), .B(n_1470), .Y(n_1678) );
INVx2_ASAP7_75t_L g1679 ( .A(n_1590), .Y(n_1679) );
INVx1_ASAP7_75t_L g1680 ( .A(n_1601), .Y(n_1680) );
INVx1_ASAP7_75t_L g1681 ( .A(n_1608), .Y(n_1681) );
INVx1_ASAP7_75t_L g1682 ( .A(n_1618), .Y(n_1682) );
NAND2xp5_ASAP7_75t_L g1683 ( .A(n_1571), .B(n_1474), .Y(n_1683) );
OR2x2_ASAP7_75t_L g1684 ( .A(n_1609), .B(n_1478), .Y(n_1684) );
AND2x2_ASAP7_75t_L g1685 ( .A(n_1607), .B(n_1478), .Y(n_1685) );
AND2x2_ASAP7_75t_L g1686 ( .A(n_1607), .B(n_1478), .Y(n_1686) );
INVx2_ASAP7_75t_SL g1687 ( .A(n_1575), .Y(n_1687) );
NAND2xp5_ASAP7_75t_L g1688 ( .A(n_1571), .B(n_1474), .Y(n_1688) );
NAND2x1_ASAP7_75t_L g1689 ( .A(n_1592), .B(n_1428), .Y(n_1689) );
INVx1_ASAP7_75t_SL g1690 ( .A(n_1580), .Y(n_1690) );
NAND2xp5_ASAP7_75t_L g1691 ( .A(n_1578), .B(n_1556), .Y(n_1691) );
NAND2xp33_ASAP7_75t_L g1692 ( .A(n_1636), .B(n_1534), .Y(n_1692) );
AND2x2_ASAP7_75t_L g1693 ( .A(n_1614), .B(n_1481), .Y(n_1693) );
NAND2xp5_ASAP7_75t_L g1694 ( .A(n_1577), .B(n_1614), .Y(n_1694) );
OR2x2_ASAP7_75t_L g1695 ( .A(n_1617), .B(n_1481), .Y(n_1695) );
INVx1_ASAP7_75t_L g1696 ( .A(n_1611), .Y(n_1696) );
AND2x4_ASAP7_75t_L g1697 ( .A(n_1615), .B(n_1481), .Y(n_1697) );
NAND2xp5_ASAP7_75t_L g1698 ( .A(n_1567), .B(n_1462), .Y(n_1698) );
OR2x2_ASAP7_75t_L g1699 ( .A(n_1572), .B(n_1548), .Y(n_1699) );
NAND2x1p5_ASAP7_75t_L g1700 ( .A(n_1568), .B(n_1454), .Y(n_1700) );
AND3x2_ASAP7_75t_L g1701 ( .A(n_1604), .B(n_1439), .C(n_1499), .Y(n_1701) );
AND2x2_ASAP7_75t_L g1702 ( .A(n_1602), .B(n_1603), .Y(n_1702) );
NAND2xp5_ASAP7_75t_L g1703 ( .A(n_1558), .B(n_1462), .Y(n_1703) );
AND2x2_ASAP7_75t_L g1704 ( .A(n_1613), .B(n_1473), .Y(n_1704) );
AND2x2_ASAP7_75t_L g1705 ( .A(n_1579), .B(n_1473), .Y(n_1705) );
AND2x2_ASAP7_75t_L g1706 ( .A(n_1584), .B(n_1482), .Y(n_1706) );
NAND2xp5_ASAP7_75t_SL g1707 ( .A(n_1592), .B(n_1545), .Y(n_1707) );
AND2x2_ASAP7_75t_L g1708 ( .A(n_1620), .B(n_1482), .Y(n_1708) );
NAND2xp5_ASAP7_75t_L g1709 ( .A(n_1558), .B(n_1446), .Y(n_1709) );
OR2x2_ASAP7_75t_L g1710 ( .A(n_1612), .B(n_1545), .Y(n_1710) );
INVx1_ASAP7_75t_L g1711 ( .A(n_1595), .Y(n_1711) );
AOI21xp33_ASAP7_75t_SL g1712 ( .A1(n_1570), .A2(n_1427), .B(n_1504), .Y(n_1712) );
AND2x2_ASAP7_75t_L g1713 ( .A(n_1620), .B(n_1548), .Y(n_1713) );
NOR2x1_ASAP7_75t_L g1714 ( .A(n_1675), .B(n_1642), .Y(n_1714) );
INVxp67_ASAP7_75t_L g1715 ( .A(n_1671), .Y(n_1715) );
AND2x2_ASAP7_75t_L g1716 ( .A(n_1702), .B(n_1615), .Y(n_1716) );
NAND2xp5_ASAP7_75t_L g1717 ( .A(n_1708), .B(n_1576), .Y(n_1717) );
OR2x2_ASAP7_75t_L g1718 ( .A(n_1652), .B(n_1576), .Y(n_1718) );
OAI221xp5_ASAP7_75t_SL g1719 ( .A1(n_1669), .A2(n_1597), .B1(n_1593), .B2(n_1605), .C(n_1641), .Y(n_1719) );
A2O1A1Ixp33_ASAP7_75t_L g1720 ( .A1(n_1649), .A2(n_1645), .B(n_1331), .C(n_1629), .Y(n_1720) );
OAI31xp33_ASAP7_75t_L g1721 ( .A1(n_1649), .A2(n_1645), .A3(n_1633), .B(n_1623), .Y(n_1721) );
INVx2_ASAP7_75t_SL g1722 ( .A(n_1690), .Y(n_1722) );
OR2x2_ASAP7_75t_L g1723 ( .A(n_1677), .B(n_1583), .Y(n_1723) );
NAND2xp5_ASAP7_75t_L g1724 ( .A(n_1708), .B(n_1587), .Y(n_1724) );
AOI321xp33_ASAP7_75t_L g1725 ( .A1(n_1712), .A2(n_1633), .A3(n_1638), .B1(n_1443), .B2(n_1562), .C(n_1634), .Y(n_1725) );
INVx1_ASAP7_75t_L g1726 ( .A(n_1651), .Y(n_1726) );
AOI22xp5_ASAP7_75t_L g1727 ( .A1(n_1698), .A2(n_1627), .B1(n_1427), .B2(n_1619), .Y(n_1727) );
NAND2xp5_ASAP7_75t_L g1728 ( .A(n_1663), .B(n_1583), .Y(n_1728) );
A2O1A1Ixp33_ASAP7_75t_L g1729 ( .A1(n_1675), .A2(n_1588), .B(n_1599), .C(n_1637), .Y(n_1729) );
OR2x2_ASAP7_75t_L g1730 ( .A(n_1694), .B(n_1595), .Y(n_1730) );
OAI22xp33_ASAP7_75t_SL g1731 ( .A1(n_1689), .A2(n_1454), .B1(n_1623), .B2(n_1636), .Y(n_1731) );
NOR2x1_ASAP7_75t_L g1732 ( .A(n_1692), .B(n_1454), .Y(n_1732) );
NOR2xp33_ASAP7_75t_L g1733 ( .A(n_1691), .B(n_1574), .Y(n_1733) );
OAI322xp33_ASAP7_75t_L g1734 ( .A1(n_1683), .A2(n_1471), .A3(n_1426), .B1(n_1463), .B2(n_1455), .C1(n_1477), .C2(n_1466), .Y(n_1734) );
INVxp67_ASAP7_75t_L g1735 ( .A(n_1661), .Y(n_1735) );
NAND2xp5_ASAP7_75t_L g1736 ( .A(n_1663), .B(n_1564), .Y(n_1736) );
AOI22xp5_ASAP7_75t_L g1737 ( .A1(n_1703), .A2(n_1619), .B1(n_1630), .B2(n_1598), .Y(n_1737) );
OR2x2_ASAP7_75t_L g1738 ( .A(n_1696), .B(n_1573), .Y(n_1738) );
O2A1O1Ixp33_ASAP7_75t_L g1739 ( .A1(n_1692), .A2(n_1445), .B(n_1502), .C(n_1511), .Y(n_1739) );
OAI21xp5_ASAP7_75t_L g1740 ( .A1(n_1707), .A2(n_1465), .B(n_1616), .Y(n_1740) );
NAND2xp5_ASAP7_75t_L g1741 ( .A(n_1711), .B(n_1589), .Y(n_1741) );
AOI32xp33_ASAP7_75t_L g1742 ( .A1(n_1654), .A2(n_1635), .A3(n_1499), .B1(n_1506), .B2(n_1537), .Y(n_1742) );
OAI21xp33_ASAP7_75t_L g1743 ( .A1(n_1658), .A2(n_1573), .B(n_1600), .Y(n_1743) );
AOI22xp33_ASAP7_75t_SL g1744 ( .A1(n_1654), .A2(n_1640), .B1(n_1636), .B2(n_1506), .Y(n_1744) );
AOI22xp5_ASAP7_75t_L g1745 ( .A1(n_1709), .A2(n_1444), .B1(n_1431), .B2(n_1471), .Y(n_1745) );
INVx1_ASAP7_75t_L g1746 ( .A(n_1655), .Y(n_1746) );
INVx2_ASAP7_75t_L g1747 ( .A(n_1699), .Y(n_1747) );
NAND2xp5_ASAP7_75t_L g1748 ( .A(n_1668), .B(n_1589), .Y(n_1748) );
AOI22xp33_ASAP7_75t_L g1749 ( .A1(n_1658), .A2(n_1444), .B1(n_1426), .B2(n_1435), .Y(n_1749) );
OAI32xp33_ASAP7_75t_L g1750 ( .A1(n_1700), .A2(n_1543), .A3(n_1451), .B1(n_1537), .B2(n_1525), .Y(n_1750) );
AOI21xp33_ASAP7_75t_L g1751 ( .A1(n_1707), .A2(n_1458), .B(n_1536), .Y(n_1751) );
OAI332xp33_ASAP7_75t_L g1752 ( .A1(n_1678), .A2(n_1440), .A3(n_1451), .B1(n_1326), .B2(n_1639), .B3(n_1631), .C1(n_1628), .C2(n_1624), .Y(n_1752) );
INVx1_ASAP7_75t_L g1753 ( .A(n_1659), .Y(n_1753) );
OAI22xp33_ASAP7_75t_L g1754 ( .A1(n_1700), .A2(n_1543), .B1(n_1384), .B2(n_1520), .Y(n_1754) );
XNOR2xp5_ASAP7_75t_L g1755 ( .A(n_1722), .B(n_1701), .Y(n_1755) );
INVx1_ASAP7_75t_L g1756 ( .A(n_1726), .Y(n_1756) );
NAND2xp5_ASAP7_75t_L g1757 ( .A(n_1752), .B(n_1676), .Y(n_1757) );
INVxp67_ASAP7_75t_L g1758 ( .A(n_1714), .Y(n_1758) );
AO22x2_ASAP7_75t_L g1759 ( .A1(n_1715), .A2(n_1673), .B1(n_1667), .B2(n_1680), .Y(n_1759) );
AOI22xp5_ASAP7_75t_L g1760 ( .A1(n_1745), .A2(n_1693), .B1(n_1688), .B2(n_1686), .Y(n_1760) );
INVx1_ASAP7_75t_L g1761 ( .A(n_1746), .Y(n_1761) );
NOR2xp33_ASAP7_75t_L g1762 ( .A(n_1735), .B(n_1664), .Y(n_1762) );
AOI21xp33_ASAP7_75t_SL g1763 ( .A1(n_1721), .A2(n_1687), .B(n_1672), .Y(n_1763) );
NOR2xp33_ASAP7_75t_L g1764 ( .A(n_1734), .B(n_1681), .Y(n_1764) );
AOI322xp5_ASAP7_75t_L g1765 ( .A1(n_1720), .A2(n_1705), .A3(n_1676), .B1(n_1704), .B2(n_1657), .C1(n_1666), .C2(n_1706), .Y(n_1765) );
OAI21xp5_ASAP7_75t_L g1766 ( .A1(n_1740), .A2(n_1687), .B(n_1682), .Y(n_1766) );
AND2x2_ASAP7_75t_L g1767 ( .A(n_1716), .B(n_1702), .Y(n_1767) );
XNOR2xp5_ASAP7_75t_L g1768 ( .A(n_1737), .B(n_1706), .Y(n_1768) );
AOI21xp33_ASAP7_75t_L g1769 ( .A1(n_1739), .A2(n_1650), .B(n_1653), .Y(n_1769) );
NAND2xp5_ASAP7_75t_L g1770 ( .A(n_1717), .B(n_1668), .Y(n_1770) );
O2A1O1Ixp33_ASAP7_75t_L g1771 ( .A1(n_1719), .A2(n_1294), .B(n_1521), .C(n_1653), .Y(n_1771) );
NOR2x1_ASAP7_75t_L g1772 ( .A(n_1732), .B(n_1547), .Y(n_1772) );
NAND3xp33_ASAP7_75t_L g1773 ( .A(n_1725), .B(n_1516), .C(n_1500), .Y(n_1773) );
OAI22xp5_ASAP7_75t_L g1774 ( .A1(n_1729), .A2(n_1656), .B1(n_1710), .B2(n_1695), .Y(n_1774) );
NAND2xp5_ASAP7_75t_SL g1775 ( .A(n_1731), .B(n_1674), .Y(n_1775) );
INVx2_ASAP7_75t_L g1776 ( .A(n_1753), .Y(n_1776) );
INVx1_ASAP7_75t_SL g1777 ( .A(n_1738), .Y(n_1777) );
INVx1_ASAP7_75t_L g1778 ( .A(n_1741), .Y(n_1778) );
AOI22xp5_ASAP7_75t_SL g1779 ( .A1(n_1733), .A2(n_1650), .B1(n_1697), .B2(n_1648), .Y(n_1779) );
OAI21xp33_ASAP7_75t_L g1780 ( .A1(n_1727), .A2(n_1693), .B(n_1704), .Y(n_1780) );
AND2x2_ASAP7_75t_L g1781 ( .A(n_1747), .B(n_1648), .Y(n_1781) );
AOI21xp33_ASAP7_75t_L g1782 ( .A1(n_1758), .A2(n_1740), .B(n_1754), .Y(n_1782) );
AOI221xp5_ASAP7_75t_L g1783 ( .A1(n_1764), .A2(n_1717), .B1(n_1728), .B2(n_1743), .C(n_1748), .Y(n_1783) );
OAI32xp33_ASAP7_75t_L g1784 ( .A1(n_1758), .A2(n_1730), .A3(n_1718), .B1(n_1723), .B2(n_1736), .Y(n_1784) );
A2O1A1Ixp33_ASAP7_75t_L g1785 ( .A1(n_1779), .A2(n_1742), .B(n_1750), .C(n_1744), .Y(n_1785) );
NOR2xp33_ASAP7_75t_L g1786 ( .A(n_1757), .B(n_1724), .Y(n_1786) );
XNOR2xp5_ASAP7_75t_L g1787 ( .A(n_1755), .B(n_1705), .Y(n_1787) );
NOR2x1_ASAP7_75t_L g1788 ( .A(n_1775), .B(n_1547), .Y(n_1788) );
AOI332xp33_ASAP7_75t_L g1789 ( .A1(n_1760), .A2(n_1749), .A3(n_1741), .B1(n_1662), .B2(n_1660), .B3(n_1685), .C1(n_1686), .C2(n_1713), .Y(n_1789) );
NOR2xp67_ASAP7_75t_L g1790 ( .A(n_1763), .B(n_1775), .Y(n_1790) );
AOI221xp5_ASAP7_75t_L g1791 ( .A1(n_1764), .A2(n_1660), .B1(n_1662), .B2(n_1685), .C(n_1751), .Y(n_1791) );
INVx1_ASAP7_75t_L g1792 ( .A(n_1759), .Y(n_1792) );
AOI22xp33_ASAP7_75t_L g1793 ( .A1(n_1780), .A2(n_1773), .B1(n_1769), .B2(n_1774), .Y(n_1793) );
OAI22xp5_ASAP7_75t_L g1794 ( .A1(n_1768), .A2(n_1656), .B1(n_1697), .B2(n_1695), .Y(n_1794) );
OAI21xp33_ASAP7_75t_L g1795 ( .A1(n_1765), .A2(n_1697), .B(n_1713), .Y(n_1795) );
AOI21xp33_ASAP7_75t_L g1796 ( .A1(n_1771), .A2(n_1751), .B(n_1518), .Y(n_1796) );
OAI21xp33_ASAP7_75t_L g1797 ( .A1(n_1759), .A2(n_1684), .B(n_1665), .Y(n_1797) );
OAI22xp5_ASAP7_75t_L g1798 ( .A1(n_1777), .A2(n_1665), .B1(n_1684), .B2(n_1670), .Y(n_1798) );
NAND2xp5_ASAP7_75t_L g1799 ( .A(n_1778), .B(n_1670), .Y(n_1799) );
AOI221xp5_ASAP7_75t_L g1800 ( .A1(n_1762), .A2(n_1535), .B1(n_1674), .B2(n_1679), .C(n_1444), .Y(n_1800) );
OAI21xp33_ASAP7_75t_SL g1801 ( .A1(n_1766), .A2(n_1527), .B(n_1679), .Y(n_1801) );
OAI22xp5_ASAP7_75t_L g1802 ( .A1(n_1785), .A2(n_1770), .B1(n_1767), .B2(n_1772), .Y(n_1802) );
INVx2_ASAP7_75t_SL g1803 ( .A(n_1798), .Y(n_1803) );
AOI211x1_ASAP7_75t_SL g1804 ( .A1(n_1790), .A2(n_1782), .B(n_1794), .C(n_1796), .Y(n_1804) );
AOI211xp5_ASAP7_75t_L g1805 ( .A1(n_1784), .A2(n_1762), .B(n_1756), .C(n_1761), .Y(n_1805) );
BUFx6f_ASAP7_75t_L g1806 ( .A(n_1799), .Y(n_1806) );
AOI221xp5_ASAP7_75t_L g1807 ( .A1(n_1791), .A2(n_1776), .B1(n_1781), .B2(n_1527), .C(n_1479), .Y(n_1807) );
AOI221xp5_ASAP7_75t_L g1808 ( .A1(n_1783), .A2(n_1435), .B1(n_1539), .B2(n_1542), .C(n_1647), .Y(n_1808) );
NAND2xp5_ASAP7_75t_SL g1809 ( .A(n_1797), .B(n_1596), .Y(n_1809) );
NAND2xp5_ASAP7_75t_L g1810 ( .A(n_1786), .B(n_1539), .Y(n_1810) );
NOR3xp33_ASAP7_75t_L g1811 ( .A(n_1792), .B(n_1402), .C(n_1389), .Y(n_1811) );
AOI31xp33_ASAP7_75t_L g1812 ( .A1(n_1793), .A2(n_1542), .A3(n_1421), .B(n_1415), .Y(n_1812) );
INVx1_ASAP7_75t_L g1813 ( .A(n_1795), .Y(n_1813) );
AND2x2_ASAP7_75t_L g1814 ( .A(n_1787), .B(n_1435), .Y(n_1814) );
OAI22xp5_ASAP7_75t_L g1815 ( .A1(n_1813), .A2(n_1788), .B1(n_1789), .B2(n_1800), .Y(n_1815) );
NAND2xp5_ASAP7_75t_SL g1816 ( .A(n_1805), .B(n_1801), .Y(n_1816) );
NOR2x1_ASAP7_75t_L g1817 ( .A(n_1802), .B(n_1547), .Y(n_1817) );
NOR2xp67_ASAP7_75t_L g1818 ( .A(n_1803), .B(n_1646), .Y(n_1818) );
NOR2xp67_ASAP7_75t_L g1819 ( .A(n_1809), .B(n_1643), .Y(n_1819) );
AOI22xp5_ASAP7_75t_L g1820 ( .A1(n_1807), .A2(n_1421), .B1(n_1384), .B2(n_1419), .Y(n_1820) );
AOI221xp5_ASAP7_75t_L g1821 ( .A1(n_1812), .A2(n_1622), .B1(n_1329), .B2(n_1332), .C(n_1335), .Y(n_1821) );
AOI31xp33_ASAP7_75t_L g1822 ( .A1(n_1804), .A2(n_1513), .A3(n_1410), .B(n_1406), .Y(n_1822) );
NOR3xp33_ASAP7_75t_SL g1823 ( .A(n_1808), .B(n_1335), .C(n_1334), .Y(n_1823) );
NAND4xp75_ASAP7_75t_L g1824 ( .A(n_1817), .B(n_1814), .C(n_1810), .D(n_1811), .Y(n_1824) );
NAND4xp25_ASAP7_75t_L g1825 ( .A(n_1815), .B(n_1816), .C(n_1820), .D(n_1818), .Y(n_1825) );
AOI22xp33_ASAP7_75t_L g1826 ( .A1(n_1821), .A2(n_1806), .B1(n_1352), .B2(n_1621), .Y(n_1826) );
XNOR2xp5_ASAP7_75t_L g1827 ( .A(n_1823), .B(n_1819), .Y(n_1827) );
INVx2_ASAP7_75t_L g1828 ( .A(n_1822), .Y(n_1828) );
NAND3xp33_ASAP7_75t_SL g1829 ( .A(n_1815), .B(n_1416), .C(n_1526), .Y(n_1829) );
OR3x1_ASAP7_75t_L g1830 ( .A(n_1829), .B(n_1334), .C(n_1332), .Y(n_1830) );
INVx1_ASAP7_75t_L g1831 ( .A(n_1827), .Y(n_1831) );
AOI222xp33_ASAP7_75t_L g1832 ( .A1(n_1828), .A2(n_1394), .B1(n_1395), .B2(n_1409), .C1(n_1408), .C2(n_1412), .Y(n_1832) );
OAI22x1_ASAP7_75t_SL g1833 ( .A1(n_1825), .A2(n_1395), .B1(n_1352), .B2(n_1408), .Y(n_1833) );
AOI22xp33_ASAP7_75t_L g1834 ( .A1(n_1831), .A2(n_1825), .B1(n_1826), .B2(n_1824), .Y(n_1834) );
INVx1_ASAP7_75t_L g1835 ( .A(n_1830), .Y(n_1835) );
INVx1_ASAP7_75t_L g1836 ( .A(n_1833), .Y(n_1836) );
INVx1_ASAP7_75t_L g1837 ( .A(n_1835), .Y(n_1837) );
AO22x2_ASAP7_75t_L g1838 ( .A1(n_1837), .A2(n_1836), .B1(n_1834), .B2(n_1832), .Y(n_1838) );
INVxp67_ASAP7_75t_L g1839 ( .A(n_1838), .Y(n_1839) );
AOI21xp5_ASAP7_75t_L g1840 ( .A1(n_1839), .A2(n_1496), .B(n_1420), .Y(n_1840) );
endmodule