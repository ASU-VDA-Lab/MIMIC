module fake_jpeg_28110_n_102 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_102);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_102;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_0),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_0),
.Y(n_12)
);

INVx6_ASAP7_75t_L g13 ( 
.A(n_2),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_4),
.Y(n_14)
);

BUFx12f_ASAP7_75t_L g15 ( 
.A(n_6),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g16 ( 
.A(n_6),
.B(n_10),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_8),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

INVx11_ASAP7_75t_L g22 ( 
.A(n_15),
.Y(n_22)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_22),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_16),
.B(n_0),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_23),
.B(n_26),
.Y(n_32)
);

INVx5_ASAP7_75t_L g24 ( 
.A(n_15),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_24),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_15),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_25),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_SL g26 ( 
.A(n_16),
.B(n_1),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_21),
.Y(n_27)
);

INVx11_ASAP7_75t_L g30 ( 
.A(n_27),
.Y(n_30)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_21),
.Y(n_28)
);

BUFx2_ASAP7_75t_L g36 ( 
.A(n_28),
.Y(n_36)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_18),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_29),
.Y(n_34)
);

OAI22xp33_ASAP7_75t_SL g33 ( 
.A1(n_29),
.A2(n_13),
.B1(n_12),
.B2(n_14),
.Y(n_33)
);

AOI22xp33_ASAP7_75t_L g44 ( 
.A1(n_33),
.A2(n_29),
.B1(n_11),
.B2(n_28),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_26),
.B(n_19),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_38),
.B(n_14),
.Y(n_41)
);

AO22x2_ASAP7_75t_SL g39 ( 
.A1(n_29),
.A2(n_13),
.B1(n_18),
.B2(n_17),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_39),
.A2(n_24),
.B1(n_22),
.B2(n_28),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_32),
.B(n_26),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_SL g52 ( 
.A(n_40),
.B(n_41),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_35),
.B(n_23),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_SL g50 ( 
.A(n_42),
.B(n_46),
.Y(n_50)
);

AND2x2_ASAP7_75t_L g43 ( 
.A(n_39),
.B(n_23),
.Y(n_43)
);

OAI21xp5_ASAP7_75t_L g55 ( 
.A1(n_43),
.A2(n_39),
.B(n_34),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_44),
.B(n_39),
.Y(n_53)
);

BUFx2_ASAP7_75t_L g45 ( 
.A(n_31),
.Y(n_45)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_45),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_35),
.B(n_11),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_36),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_SL g56 ( 
.A(n_47),
.B(n_31),
.Y(n_56)
);

HAxp5_ASAP7_75t_SL g58 ( 
.A(n_48),
.B(n_27),
.CON(n_58),
.SN(n_58)
);

NAND2xp5_ASAP7_75t_SL g49 ( 
.A(n_34),
.B(n_27),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_49),
.B(n_42),
.Y(n_54)
);

CKINVDCx16_ASAP7_75t_R g51 ( 
.A(n_49),
.Y(n_51)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_51),
.Y(n_62)
);

AND2x2_ASAP7_75t_L g66 ( 
.A(n_53),
.B(n_54),
.Y(n_66)
);

XNOR2xp5_ASAP7_75t_L g67 ( 
.A(n_55),
.B(n_48),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_56),
.Y(n_64)
);

NAND2x1p5_ASAP7_75t_R g70 ( 
.A(n_58),
.B(n_27),
.Y(n_70)
);

INVxp67_ASAP7_75t_L g59 ( 
.A(n_46),
.Y(n_59)
);

NOR3xp33_ASAP7_75t_L g68 ( 
.A(n_59),
.B(n_27),
.C(n_37),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_41),
.B(n_21),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_60),
.A2(n_24),
.B1(n_22),
.B2(n_30),
.Y(n_65)
);

XOR2xp5_ASAP7_75t_L g61 ( 
.A(n_54),
.B(n_43),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_61),
.B(n_65),
.Y(n_73)
);

AOI21xp5_ASAP7_75t_L g63 ( 
.A1(n_55),
.A2(n_59),
.B(n_50),
.Y(n_63)
);

OAI21xp5_ASAP7_75t_SL g76 ( 
.A1(n_63),
.A2(n_68),
.B(n_70),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_67),
.B(n_69),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g69 ( 
.A(n_50),
.B(n_43),
.C(n_58),
.Y(n_69)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_66),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_71),
.B(n_74),
.Y(n_84)
);

HB1xp67_ASAP7_75t_L g72 ( 
.A(n_70),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_72),
.Y(n_80)
);

INVxp67_ASAP7_75t_L g74 ( 
.A(n_66),
.Y(n_74)
);

AOI21xp33_ASAP7_75t_L g75 ( 
.A1(n_69),
.A2(n_52),
.B(n_5),
.Y(n_75)
);

AOI21xp5_ASAP7_75t_L g85 ( 
.A1(n_75),
.A2(n_1),
.B(n_2),
.Y(n_85)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_64),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_78),
.B(n_79),
.Y(n_83)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_67),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g81 ( 
.A(n_77),
.B(n_61),
.C(n_62),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_SL g89 ( 
.A(n_81),
.B(n_83),
.Y(n_89)
);

OAI321xp33_ASAP7_75t_L g82 ( 
.A1(n_73),
.A2(n_17),
.A3(n_5),
.B1(n_7),
.B2(n_9),
.C(n_10),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_82),
.A2(n_57),
.B1(n_30),
.B2(n_4),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_85),
.B(n_1),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_74),
.A2(n_20),
.B1(n_47),
.B2(n_57),
.Y(n_86)
);

AND2x2_ASAP7_75t_L g88 ( 
.A(n_86),
.B(n_84),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_87),
.B(n_90),
.Y(n_95)
);

AOI322xp5_ASAP7_75t_L g92 ( 
.A1(n_88),
.A2(n_76),
.A3(n_83),
.B1(n_36),
.B2(n_45),
.C1(n_20),
.C2(n_25),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_89),
.B(n_91),
.C(n_25),
.Y(n_93)
);

FAx1_ASAP7_75t_L g90 ( 
.A(n_80),
.B(n_76),
.CI(n_27),
.CON(n_90),
.SN(n_90)
);

XNOR2xp5_ASAP7_75t_L g97 ( 
.A(n_92),
.B(n_93),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_90),
.B(n_25),
.C(n_37),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_94),
.Y(n_98)
);

AOI211xp5_ASAP7_75t_SL g96 ( 
.A1(n_95),
.A2(n_87),
.B(n_45),
.C(n_3),
.Y(n_96)
);

OAI321xp33_ASAP7_75t_L g100 ( 
.A1(n_96),
.A2(n_3),
.A3(n_36),
.B1(n_37),
.B2(n_98),
.C(n_97),
.Y(n_100)
);

OAI21x1_ASAP7_75t_L g99 ( 
.A1(n_96),
.A2(n_2),
.B(n_3),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_99),
.B(n_100),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_101),
.B(n_37),
.Y(n_102)
);


endmodule