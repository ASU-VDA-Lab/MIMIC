module real_jpeg_17678_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_215;
wire n_166;
wire n_176;
wire n_221;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_164;
wire n_48;
wire n_200;
wire n_140;
wire n_227;
wire n_126;
wire n_214;
wire n_13;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_93;
wire n_141;
wire n_95;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_208;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_203;
wire n_192;
wire n_100;
wire n_198;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_110;
wire n_61;
wire n_195;
wire n_205;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_30;
wire n_204;
wire n_158;
wire n_149;
wire n_144;
wire n_15;
wire n_130;
wire n_103;
wire n_225;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_185;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_97;
wire n_75;
wire n_187;
wire n_34;
wire n_190;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_167;
wire n_128;
wire n_202;
wire n_179;
wire n_213;
wire n_216;
wire n_133;
wire n_138;
wire n_25;
wire n_217;
wire n_53;
wire n_206;
wire n_127;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;
wire n_16;

AND2x4_ASAP7_75t_L g28 ( 
.A(n_0),
.B(n_29),
.Y(n_28)
);

AND2x2_ASAP7_75t_L g38 ( 
.A(n_0),
.B(n_39),
.Y(n_38)
);

AND2x2_ASAP7_75t_L g54 ( 
.A(n_0),
.B(n_55),
.Y(n_54)
);

AND2x4_ASAP7_75t_SL g66 ( 
.A(n_0),
.B(n_67),
.Y(n_66)
);

AND2x4_ASAP7_75t_L g92 ( 
.A(n_0),
.B(n_93),
.Y(n_92)
);

AND2x2_ASAP7_75t_L g110 ( 
.A(n_0),
.B(n_49),
.Y(n_110)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_0),
.Y(n_133)
);

NAND2x1p5_ASAP7_75t_L g174 ( 
.A(n_0),
.B(n_175),
.Y(n_174)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_1),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_1),
.Y(n_40)
);

BUFx5_ASAP7_75t_L g49 ( 
.A(n_2),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_2),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_3),
.B(n_179),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_3),
.B(n_219),
.Y(n_218)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_4),
.Y(n_61)
);

BUFx5_ASAP7_75t_L g67 ( 
.A(n_4),
.Y(n_67)
);

BUFx5_ASAP7_75t_L g84 ( 
.A(n_4),
.Y(n_84)
);

BUFx3_ASAP7_75t_L g183 ( 
.A(n_4),
.Y(n_183)
);

AND2x2_ASAP7_75t_L g22 ( 
.A(n_5),
.B(n_23),
.Y(n_22)
);

INVx2_ASAP7_75t_SL g47 ( 
.A(n_5),
.Y(n_47)
);

AND2x2_ASAP7_75t_L g96 ( 
.A(n_5),
.B(n_97),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g142 ( 
.A(n_5),
.B(n_33),
.Y(n_142)
);

AND2x2_ASAP7_75t_L g205 ( 
.A(n_5),
.B(n_206),
.Y(n_205)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_6),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_7),
.B(n_32),
.Y(n_31)
);

AND2x2_ASAP7_75t_SL g42 ( 
.A(n_7),
.B(n_43),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_7),
.B(n_59),
.Y(n_58)
);

AND2x2_ASAP7_75t_L g63 ( 
.A(n_7),
.B(n_64),
.Y(n_63)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_7),
.B(n_78),
.Y(n_77)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_7),
.Y(n_126)
);

AND2x2_ASAP7_75t_SL g163 ( 
.A(n_7),
.B(n_164),
.Y(n_163)
);

AND2x2_ASAP7_75t_SL g214 ( 
.A(n_7),
.B(n_215),
.Y(n_214)
);

INVx6_ASAP7_75t_L g136 ( 
.A(n_8),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g166 ( 
.A(n_8),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_9),
.Y(n_130)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_10),
.Y(n_57)
);

BUFx12f_ASAP7_75t_L g80 ( 
.A(n_10),
.Y(n_80)
);

BUFx4f_ASAP7_75t_L g221 ( 
.A(n_10),
.Y(n_221)
);

BUFx5_ASAP7_75t_L g175 ( 
.A(n_11),
.Y(n_175)
);

BUFx8_ASAP7_75t_L g215 ( 
.A(n_11),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_190),
.Y(n_12)
);

HB1xp67_ASAP7_75t_L g13 ( 
.A(n_14),
.Y(n_13)
);

OAI21xp5_ASAP7_75t_SL g14 ( 
.A1(n_15),
.A2(n_152),
.B(n_189),
.Y(n_14)
);

AOI21xp5_ASAP7_75t_L g15 ( 
.A1(n_16),
.A2(n_119),
.B(n_151),
.Y(n_15)
);

OAI21x1_ASAP7_75t_L g16 ( 
.A1(n_17),
.A2(n_89),
.B(n_118),
.Y(n_16)
);

NOR2xp67_ASAP7_75t_SL g17 ( 
.A(n_18),
.B(n_71),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_18),
.B(n_71),
.Y(n_118)
);

XOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_50),
.Y(n_18)
);

OAI22xp5_ASAP7_75t_SL g19 ( 
.A1(n_20),
.A2(n_21),
.B1(n_35),
.B2(n_36),
.Y(n_19)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_20),
.B(n_36),
.C(n_50),
.Y(n_120)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_26),
.B1(n_27),
.B2(n_34),
.Y(n_21)
);

INVx1_ASAP7_75t_SL g34 ( 
.A(n_22),
.Y(n_34)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_22),
.B(n_28),
.C(n_148),
.Y(n_147)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g94 ( 
.A(n_25),
.Y(n_94)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

XNOR2xp5_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_31),
.Y(n_27)
);

BUFx2_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_31),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_31),
.A2(n_148),
.B1(n_162),
.B2(n_168),
.Y(n_161)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

MAJIxp5_ASAP7_75t_L g36 ( 
.A(n_37),
.B(n_41),
.C(n_46),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_37),
.A2(n_38),
.B1(n_46),
.B2(n_74),
.Y(n_73)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

XNOR2xp5_ASAP7_75t_L g203 ( 
.A(n_38),
.B(n_204),
.Y(n_203)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_41),
.A2(n_42),
.B1(n_73),
.B2(n_75),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_41),
.A2(n_42),
.B1(n_141),
.B2(n_144),
.Y(n_140)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

O2A1O1Ixp33_ASAP7_75t_L g158 ( 
.A1(n_42),
.A2(n_101),
.B(n_110),
.C(n_142),
.Y(n_158)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx1_ASAP7_75t_SL g74 ( 
.A(n_46),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_46),
.A2(n_74),
.B1(n_125),
.B2(n_137),
.Y(n_200)
);

OR2x2_ASAP7_75t_L g46 ( 
.A(n_47),
.B(n_48),
.Y(n_46)
);

OR2x2_ASAP7_75t_L g82 ( 
.A(n_47),
.B(n_83),
.Y(n_82)
);

OR2x2_ASAP7_75t_L g184 ( 
.A(n_47),
.B(n_185),
.Y(n_184)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

XNOR2xp5_ASAP7_75t_L g50 ( 
.A(n_51),
.B(n_62),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

AOI21xp5_ASAP7_75t_L g106 ( 
.A1(n_52),
.A2(n_107),
.B(n_111),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_SL g138 ( 
.A1(n_52),
.A2(n_63),
.B(n_70),
.Y(n_138)
);

NOR2x1_ASAP7_75t_R g52 ( 
.A(n_53),
.B(n_58),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_53),
.A2(n_54),
.B1(n_81),
.B2(n_82),
.Y(n_150)
);

INVx2_ASAP7_75t_SL g53 ( 
.A(n_54),
.Y(n_53)
);

OAI21xp5_ASAP7_75t_L g65 ( 
.A1(n_54),
.A2(n_66),
.B(n_68),
.Y(n_65)
);

NAND2x1p5_ASAP7_75t_L g68 ( 
.A(n_54),
.B(n_66),
.Y(n_68)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_57),
.Y(n_98)
);

OAI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_58),
.A2(n_96),
.B1(n_99),
.B2(n_100),
.Y(n_95)
);

INVxp33_ASAP7_75t_L g100 ( 
.A(n_58),
.Y(n_100)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_63),
.A2(n_65),
.B1(n_69),
.B2(n_70),
.Y(n_62)
);

CKINVDCx16_ASAP7_75t_R g69 ( 
.A(n_63),
.Y(n_69)
);

O2A1O1Ixp33_ASAP7_75t_SL g91 ( 
.A1(n_63),
.A2(n_92),
.B(n_95),
.C(n_101),
.Y(n_91)
);

AND2x2_ASAP7_75t_L g101 ( 
.A(n_63),
.B(n_92),
.Y(n_101)
);

OAI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_63),
.A2(n_69),
.B1(n_92),
.B2(n_115),
.Y(n_114)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_65),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_66),
.A2(n_77),
.B1(n_87),
.B2(n_88),
.Y(n_86)
);

INVx1_ASAP7_75t_SL g87 ( 
.A(n_66),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_66),
.B(n_96),
.Y(n_160)
);

XOR2xp5_ASAP7_75t_L g123 ( 
.A(n_68),
.B(n_124),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_68),
.B(n_125),
.C(n_132),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g71 ( 
.A(n_72),
.B(n_76),
.C(n_85),
.Y(n_71)
);

XOR2xp5_ASAP7_75t_L g102 ( 
.A(n_72),
.B(n_103),
.Y(n_102)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_73),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_76),
.A2(n_85),
.B1(n_86),
.B2(n_104),
.Y(n_103)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_76),
.Y(n_104)
);

OAI21xp5_ASAP7_75t_SL g108 ( 
.A1(n_76),
.A2(n_77),
.B(n_81),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_77),
.B(n_81),
.Y(n_76)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_77),
.Y(n_88)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_81),
.A2(n_82),
.B1(n_217),
.B2(n_218),
.Y(n_216)
);

INVx1_ASAP7_75t_SL g81 ( 
.A(n_82),
.Y(n_81)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

AOI21xp5_ASAP7_75t_L g89 ( 
.A1(n_90),
.A2(n_105),
.B(n_117),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_102),
.Y(n_90)
);

NOR2xp67_ASAP7_75t_L g117 ( 
.A(n_91),
.B(n_102),
.Y(n_117)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_92),
.Y(n_115)
);

XNOR2xp5_ASAP7_75t_L g172 ( 
.A(n_92),
.B(n_109),
.Y(n_172)
);

MAJx2_ASAP7_75t_L g199 ( 
.A(n_92),
.B(n_110),
.C(n_174),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_92),
.A2(n_115),
.B1(n_203),
.B2(n_207),
.Y(n_202)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

XOR2xp5_ASAP7_75t_L g113 ( 
.A(n_95),
.B(n_114),
.Y(n_113)
);

INVx1_ASAP7_75t_SL g99 ( 
.A(n_96),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_96),
.A2(n_99),
.B1(n_163),
.B2(n_167),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_96),
.B(n_148),
.C(n_163),
.Y(n_224)
);

INVx4_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_104),
.B(n_113),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_104),
.B(n_113),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_L g105 ( 
.A1(n_106),
.A2(n_112),
.B(n_116),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_108),
.B(n_109),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_108),
.B(n_109),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_109),
.A2(n_110),
.B1(n_142),
.B2(n_143),
.Y(n_141)
);

INVx2_ASAP7_75t_SL g109 ( 
.A(n_110),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_120),
.B(n_121),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_120),
.B(n_121),
.Y(n_151)
);

XOR2x2_ASAP7_75t_L g121 ( 
.A(n_122),
.B(n_139),
.Y(n_121)
);

XOR2xp5_ASAP7_75t_L g122 ( 
.A(n_123),
.B(n_138),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_123),
.B(n_138),
.C(n_139),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_125),
.A2(n_131),
.B1(n_132),
.B2(n_137),
.Y(n_124)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_125),
.Y(n_137)
);

OR2x2_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_127),
.Y(n_125)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVx3_ASAP7_75t_L g185 ( 
.A(n_129),
.Y(n_185)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

INVx1_ASAP7_75t_SL g131 ( 
.A(n_132),
.Y(n_131)
);

OR2x2_ASAP7_75t_L g132 ( 
.A(n_133),
.B(n_134),
.Y(n_132)
);

INVx6_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx4_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_136),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_SL g139 ( 
.A(n_140),
.B(n_145),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_140),
.B(n_146),
.C(n_150),
.Y(n_155)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_141),
.Y(n_144)
);

INVxp67_ASAP7_75t_L g143 ( 
.A(n_142),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_146),
.A2(n_147),
.B1(n_149),
.B2(n_150),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_188),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_153),
.B(n_188),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_169),
.Y(n_153)
);

XOR2xp5_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_156),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_155),
.B(n_156),
.C(n_169),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_161),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_159),
.Y(n_157)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_158),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_159),
.B(n_161),
.C(n_209),
.Y(n_208)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_162),
.Y(n_168)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_163),
.Y(n_167)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_SL g169 ( 
.A(n_170),
.B(n_187),
.Y(n_169)
);

XOR2xp5_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_177),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_171),
.B(n_177),
.C(n_187),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_172),
.A2(n_173),
.B1(n_174),
.B2(n_176),
.Y(n_171)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_172),
.Y(n_176)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_L g177 ( 
.A1(n_178),
.A2(n_184),
.B(n_186),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_178),
.B(n_184),
.Y(n_186)
);

INVx5_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

INVx6_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

INVx5_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

INVx3_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_186),
.A2(n_223),
.B1(n_224),
.B2(n_225),
.Y(n_222)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_186),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_191),
.B(n_227),
.Y(n_190)
);

HB1xp67_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_193),
.B(n_194),
.Y(n_192)
);

OR2x2_ASAP7_75t_L g227 ( 
.A(n_193),
.B(n_194),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g194 ( 
.A(n_195),
.B(n_210),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_208),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_197),
.A2(n_198),
.B1(n_201),
.B2(n_202),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

XNOR2x2_ASAP7_75t_L g198 ( 
.A(n_199),
.B(n_200),
.Y(n_198)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_203),
.Y(n_207)
);

INVx1_ASAP7_75t_SL g204 ( 
.A(n_205),
.Y(n_204)
);

XOR2xp5_ASAP7_75t_L g210 ( 
.A(n_211),
.B(n_226),
.Y(n_210)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_212),
.B(n_222),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g212 ( 
.A(n_213),
.B(n_216),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);


endmodule