module fake_jpeg_7400_n_63 (n_13, n_21, n_1, n_10, n_23, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_63);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_63;

wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_27;
wire n_55;
wire n_51;
wire n_47;
wire n_40;
wire n_59;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_62;
wire n_31;
wire n_25;
wire n_56;
wire n_37;
wire n_29;
wire n_43;
wire n_50;
wire n_32;

NAND2xp5_ASAP7_75t_SL g24 ( 
.A(n_3),
.B(n_11),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_21),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_15),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_16),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_20),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_2),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_24),
.Y(n_33)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_33),
.Y(n_42)
);

INVx2_ASAP7_75t_SL g34 ( 
.A(n_27),
.Y(n_34)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_34),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_31),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_SL g51 ( 
.A(n_35),
.B(n_13),
.Y(n_51)
);

OAI21xp33_ASAP7_75t_L g36 ( 
.A1(n_30),
.A2(n_0),
.B(n_23),
.Y(n_36)
);

OAI21xp5_ASAP7_75t_SL g46 ( 
.A1(n_36),
.A2(n_38),
.B(n_8),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_26),
.Y(n_37)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_37),
.Y(n_48)
);

CKINVDCx14_ASAP7_75t_R g38 ( 
.A(n_25),
.Y(n_38)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_29),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_SL g43 ( 
.A(n_39),
.B(n_4),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_SL g40 ( 
.A(n_28),
.B(n_1),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_40),
.B(n_12),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g41 ( 
.A1(n_38),
.A2(n_32),
.B1(n_5),
.B2(n_7),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_41),
.A2(n_51),
.B1(n_52),
.B2(n_53),
.Y(n_57)
);

AND2x2_ASAP7_75t_L g55 ( 
.A(n_43),
.B(n_50),
.Y(n_55)
);

INVxp67_ASAP7_75t_L g45 ( 
.A(n_34),
.Y(n_45)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_45),
.Y(n_56)
);

FAx1_ASAP7_75t_SL g54 ( 
.A(n_46),
.B(n_47),
.CI(n_49),
.CON(n_54),
.SN(n_54)
);

MAJx2_ASAP7_75t_L g47 ( 
.A(n_33),
.B(n_9),
.C(n_10),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_SL g50 ( 
.A(n_33),
.B(n_22),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_33),
.B(n_17),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_SL g53 ( 
.A(n_33),
.B(n_18),
.Y(n_53)
);

XOR2xp5_ASAP7_75t_L g58 ( 
.A(n_57),
.B(n_42),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_SL g59 ( 
.A(n_58),
.B(n_54),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_59),
.B(n_55),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_60),
.Y(n_61)
);

MAJIxp5_ASAP7_75t_L g62 ( 
.A(n_61),
.B(n_56),
.C(n_44),
.Y(n_62)
);

OAI21xp5_ASAP7_75t_L g63 ( 
.A1(n_62),
.A2(n_48),
.B(n_19),
.Y(n_63)
);


endmodule