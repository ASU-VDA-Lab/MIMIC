module fake_jpeg_3395_n_228 (n_13, n_21, n_53, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_51, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_52, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_228);

input n_13;
input n_21;
input n_53;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_51;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_52;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_228;

wire n_159;
wire n_117;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_155;
wire n_207;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_223;
wire n_171;
wire n_119;
wire n_69;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_143;
wire n_202;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_91;
wire n_54;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_149;
wire n_157;
wire n_87;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_29),
.Y(n_54)
);

CKINVDCx16_ASAP7_75t_R g55 ( 
.A(n_42),
.Y(n_55)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_27),
.Y(n_56)
);

BUFx24_ASAP7_75t_L g57 ( 
.A(n_0),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_25),
.Y(n_58)
);

INVx1_ASAP7_75t_SL g59 ( 
.A(n_45),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_39),
.Y(n_60)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_36),
.Y(n_61)
);

BUFx16f_ASAP7_75t_L g62 ( 
.A(n_2),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_9),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_47),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_51),
.Y(n_65)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_38),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_10),
.Y(n_67)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_24),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_6),
.Y(n_69)
);

BUFx5_ASAP7_75t_L g70 ( 
.A(n_35),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_40),
.B(n_44),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_13),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_41),
.Y(n_73)
);

BUFx12_ASAP7_75t_L g74 ( 
.A(n_23),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_53),
.Y(n_75)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_31),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_13),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_6),
.Y(n_78)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_19),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_62),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_80),
.B(n_82),
.Y(n_91)
);

BUFx12f_ASAP7_75t_L g81 ( 
.A(n_74),
.Y(n_81)
);

BUFx12f_ASAP7_75t_L g93 ( 
.A(n_81),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_79),
.B(n_52),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_SL g83 ( 
.A(n_63),
.B(n_0),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_83),
.B(n_84),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_59),
.B(n_1),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_60),
.Y(n_85)
);

BUFx3_ASAP7_75t_L g88 ( 
.A(n_85),
.Y(n_88)
);

BUFx3_ASAP7_75t_L g86 ( 
.A(n_62),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_86),
.Y(n_89)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_62),
.Y(n_87)
);

BUFx12f_ASAP7_75t_L g99 ( 
.A(n_87),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_87),
.A2(n_79),
.B1(n_57),
.B2(n_67),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_90),
.A2(n_100),
.B1(n_55),
.B2(n_70),
.Y(n_116)
);

CKINVDCx12_ASAP7_75t_R g94 ( 
.A(n_80),
.Y(n_94)
);

CKINVDCx16_ASAP7_75t_R g102 ( 
.A(n_94),
.Y(n_102)
);

CKINVDCx9p33_ASAP7_75t_R g95 ( 
.A(n_81),
.Y(n_95)
);

CKINVDCx16_ASAP7_75t_R g120 ( 
.A(n_95),
.Y(n_120)
);

AO22x2_ASAP7_75t_L g96 ( 
.A1(n_86),
.A2(n_68),
.B1(n_66),
.B2(n_76),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g110 ( 
.A(n_96),
.B(n_81),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_82),
.A2(n_66),
.B1(n_76),
.B2(n_77),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_97),
.B(n_58),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_85),
.Y(n_98)
);

BUFx3_ASAP7_75t_L g115 ( 
.A(n_98),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_81),
.A2(n_57),
.B1(n_68),
.B2(n_61),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_L g101 ( 
.A1(n_84),
.A2(n_69),
.B1(n_72),
.B2(n_78),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_L g117 ( 
.A1(n_101),
.A2(n_58),
.B1(n_96),
.B2(n_54),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_91),
.B(n_83),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_SL g134 ( 
.A(n_103),
.B(n_105),
.Y(n_134)
);

OR2x2_ASAP7_75t_SL g104 ( 
.A(n_101),
.B(n_61),
.Y(n_104)
);

CKINVDCx16_ASAP7_75t_R g121 ( 
.A(n_104),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_92),
.B(n_65),
.Y(n_105)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_98),
.Y(n_106)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_106),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_89),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_107),
.B(n_108),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_88),
.B(n_65),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_SL g109 ( 
.A1(n_100),
.A2(n_59),
.B(n_57),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_109),
.B(n_110),
.C(n_116),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_110),
.A2(n_111),
.B1(n_116),
.B2(n_117),
.Y(n_131)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_99),
.Y(n_112)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_112),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_96),
.B(n_73),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_113),
.B(n_56),
.Y(n_130)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_89),
.Y(n_114)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_114),
.Y(n_125)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_99),
.Y(n_118)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_118),
.Y(n_129)
);

HB1xp67_ASAP7_75t_L g119 ( 
.A(n_99),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_119),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_102),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_126),
.B(n_127),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_111),
.B(n_64),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_130),
.B(n_132),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_120),
.B(n_75),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_114),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_133),
.B(n_135),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_118),
.B(n_71),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_112),
.B(n_56),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_136),
.B(n_139),
.Y(n_160)
);

INVx6_ASAP7_75t_L g137 ( 
.A(n_115),
.Y(n_137)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_137),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_L g138 ( 
.A1(n_110),
.A2(n_93),
.B(n_70),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_SL g164 ( 
.A1(n_138),
.A2(n_4),
.B(n_5),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_106),
.B(n_1),
.Y(n_139)
);

INVxp67_ASAP7_75t_L g149 ( 
.A(n_140),
.Y(n_149)
);

BUFx5_ASAP7_75t_L g141 ( 
.A(n_109),
.Y(n_141)
);

INVx13_ASAP7_75t_L g148 ( 
.A(n_141),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_104),
.B(n_34),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_142),
.B(n_5),
.Y(n_165)
);

BUFx3_ASAP7_75t_L g143 ( 
.A(n_137),
.Y(n_143)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_143),
.Y(n_175)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_125),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_145),
.B(n_151),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_126),
.B(n_115),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_SL g170 ( 
.A(n_146),
.B(n_163),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_124),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_125),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_152),
.B(n_161),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_L g153 ( 
.A(n_127),
.B(n_93),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_153),
.B(n_155),
.C(n_158),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_121),
.A2(n_93),
.B1(n_74),
.B2(n_4),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_154),
.A2(n_8),
.B1(n_11),
.B2(n_12),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_140),
.B(n_74),
.C(n_50),
.Y(n_155)
);

INVxp67_ASAP7_75t_L g156 ( 
.A(n_138),
.Y(n_156)
);

INVxp67_ASAP7_75t_L g186 ( 
.A(n_156),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_131),
.B(n_49),
.C(n_48),
.Y(n_158)
);

AOI21xp5_ASAP7_75t_L g159 ( 
.A1(n_141),
.A2(n_2),
.B(n_3),
.Y(n_159)
);

AOI21xp5_ASAP7_75t_L g185 ( 
.A1(n_159),
.A2(n_164),
.B(n_15),
.Y(n_185)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_123),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_122),
.B(n_129),
.C(n_142),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_162),
.B(n_128),
.C(n_46),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_134),
.B(n_3),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_165),
.B(n_166),
.Y(n_184)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_123),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_156),
.A2(n_122),
.B1(n_129),
.B2(n_128),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_167),
.A2(n_16),
.B1(n_17),
.B2(n_18),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_162),
.B(n_150),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_168),
.B(n_171),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_SL g171 ( 
.A(n_147),
.B(n_7),
.Y(n_171)
);

A2O1A1O1Ixp25_ASAP7_75t_L g172 ( 
.A1(n_149),
.A2(n_144),
.B(n_148),
.C(n_155),
.D(n_153),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_SL g193 ( 
.A1(n_172),
.A2(n_176),
.B(n_185),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_173),
.B(n_22),
.C(n_32),
.Y(n_189)
);

AOI221xp5_ASAP7_75t_L g176 ( 
.A1(n_149),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.C(n_10),
.Y(n_176)
);

CKINVDCx16_ASAP7_75t_R g178 ( 
.A(n_160),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_178),
.B(n_179),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_158),
.B(n_164),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_180),
.B(n_183),
.Y(n_199)
);

OAI22x1_ASAP7_75t_L g181 ( 
.A1(n_148),
.A2(n_21),
.B1(n_37),
.B2(n_33),
.Y(n_181)
);

OA21x2_ASAP7_75t_L g192 ( 
.A1(n_181),
.A2(n_43),
.B(n_30),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_154),
.A2(n_11),
.B1(n_12),
.B2(n_14),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_182),
.A2(n_16),
.B1(n_17),
.B2(n_18),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_159),
.B(n_14),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_157),
.B(n_15),
.Y(n_187)
);

CKINVDCx16_ASAP7_75t_R g190 ( 
.A(n_187),
.Y(n_190)
);

AO21x1_ASAP7_75t_L g188 ( 
.A1(n_186),
.A2(n_157),
.B(n_143),
.Y(n_188)
);

INVxp67_ASAP7_75t_L g205 ( 
.A(n_188),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_189),
.B(n_196),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_191),
.A2(n_200),
.B1(n_181),
.B2(n_184),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_192),
.A2(n_195),
.B1(n_182),
.B2(n_180),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_177),
.Y(n_196)
);

CKINVDCx16_ASAP7_75t_R g197 ( 
.A(n_174),
.Y(n_197)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_197),
.Y(n_209)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_175),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_L g214 ( 
.A1(n_201),
.A2(n_206),
.B1(n_210),
.B2(n_192),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_188),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_202),
.B(n_207),
.Y(n_212)
);

XOR2xp5_ASAP7_75t_L g204 ( 
.A(n_194),
.B(n_173),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_204),
.B(n_169),
.C(n_189),
.Y(n_211)
);

NOR3xp33_ASAP7_75t_SL g207 ( 
.A(n_199),
.B(n_186),
.C(n_172),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_198),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_208),
.B(n_190),
.Y(n_213)
);

AOI21xp5_ASAP7_75t_L g210 ( 
.A1(n_193),
.A2(n_170),
.B(n_169),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_211),
.B(n_213),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_214),
.B(n_215),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_204),
.B(n_195),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_209),
.Y(n_216)
);

OAI22xp33_ASAP7_75t_SL g219 ( 
.A1(n_216),
.A2(n_205),
.B1(n_203),
.B2(n_207),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_205),
.A2(n_191),
.B1(n_192),
.B2(n_19),
.Y(n_217)
);

INVx6_ASAP7_75t_L g221 ( 
.A(n_217),
.Y(n_221)
);

INVxp67_ASAP7_75t_L g222 ( 
.A(n_219),
.Y(n_222)
);

OAI21xp5_ASAP7_75t_SL g223 ( 
.A1(n_220),
.A2(n_212),
.B(n_211),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_223),
.B(n_218),
.C(n_215),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_224),
.B(n_219),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_225),
.A2(n_222),
.B1(n_221),
.B2(n_28),
.Y(n_226)
);

OAI21xp5_ASAP7_75t_L g227 ( 
.A1(n_226),
.A2(n_26),
.B(n_20),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_227),
.B(n_20),
.Y(n_228)
);


endmodule