module real_jpeg_30490_n_19 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_16, n_15, n_689, n_13, n_19);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_689;
input n_13;

output n_19;

wire n_661;
wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_598;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_630;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_663;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_648;
wire n_95;
wire n_541;
wire n_441;
wire n_657;
wire n_643;
wire n_656;
wire n_557;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_669;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_679;
wire n_239;
wire n_290;
wire n_553;
wire n_121;
wire n_234;
wire n_640;
wire n_666;
wire n_160;
wire n_211;
wire n_574;
wire n_627;
wire n_595;
wire n_490;
wire n_39;
wire n_685;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_680;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_203;
wire n_198;
wire n_500;
wire n_562;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_678;
wire n_30;
wire n_332;
wire n_149;
wire n_366;
wire n_328;
wire n_578;
wire n_456;
wire n_620;
wire n_259;
wire n_556;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_560;
wire n_538;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_565;
wire n_466;
wire n_623;
wire n_353;
wire n_668;
wire n_453;
wire n_551;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_605;
wire n_483;
wire n_367;
wire n_639;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_464;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_422;
wire n_682;
wire n_317;
wire n_658;
wire n_506;
wire n_108;
wire n_550;
wire n_233;
wire n_73;
wire n_621;
wire n_532;
wire n_348;
wire n_516;
wire n_473;
wire n_674;
wire n_252;
wire n_601;
wire n_655;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_525;
wire n_221;
wire n_393;
wire n_489;
wire n_611;
wire n_104;
wire n_153;
wire n_634;
wire n_599;
wire n_443;
wire n_337;
wire n_544;
wire n_131;
wire n_439;
wire n_607;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_561;
wire n_684;
wire n_378;
wire n_98;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_569;
wire n_335;
wire n_646;
wire n_214;
wire n_671;
wire n_113;
wire n_566;
wire n_543;
wire n_251;
wire n_459;
wire n_576;
wire n_139;
wire n_33;
wire n_631;
wire n_673;
wire n_175;
wire n_338;
wire n_653;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_577;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_650;
wire n_564;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_470;
wire n_372;
wire n_219;
wire n_122;
wire n_262;
wire n_652;
wire n_334;
wire n_647;
wire n_383;
wire n_593;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_590;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_612;
wire n_110;
wire n_195;
wire n_592;
wire n_533;
wire n_289;
wire n_117;
wire n_614;
wire n_193;
wire n_651;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_559;
wire n_232;
wire n_582;
wire n_448;
wire n_615;
wire n_212;
wire n_284;
wire n_579;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_583;
wire n_60;
wire n_263;
wire n_46;
wire n_672;
wire n_59;
wire n_452;
wire n_213;
wire n_670;
wire n_511;
wire n_524;
wire n_589;
wire n_25;
wire n_480;
wire n_542;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_644;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_632;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_638;
wire n_497;
wire n_633;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_596;
wire n_617;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_594;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_604;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_412;
wire n_120;
wire n_155;
wire n_405;
wire n_572;
wire n_586;
wire n_548;
wire n_319;
wire n_664;
wire n_93;
wire n_487;
wire n_242;
wire n_493;
wire n_637;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_613;
wire n_231;
wire n_44;
wire n_635;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_642;
wire n_172;
wire n_285;
wire n_531;
wire n_546;
wire n_112;
wire n_554;
wire n_508;
wire n_145;
wire n_266;
wire n_654;
wire n_616;
wire n_377;
wire n_686;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_536;
wire n_148;
wire n_373;
wire n_563;
wire n_558;
wire n_510;
wire n_396;
wire n_501;
wire n_600;
wire n_392;
wire n_575;
wire n_196;
wire n_375;
wire n_667;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_584;
wire n_270;
wire n_683;
wire n_159;
wire n_429;
wire n_347;
wire n_622;
wire n_183;
wire n_248;
wire n_192;
wire n_624;
wire n_537;
wire n_318;
wire n_603;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_677;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_628;
wire n_413;
wire n_585;
wire n_494;
wire n_539;
wire n_512;
wire n_75;
wire n_581;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_675;
wire n_138;
wire n_662;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_534;
wire n_256;
wire n_520;
wire n_253;
wire n_273;
wire n_649;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_545;
wire n_484;
wire n_587;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_502;
wire n_418;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_608;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_681;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_602;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_571;
wire n_610;
wire n_573;
wire n_379;
wire n_141;
wire n_555;
wire n_65;
wire n_188;
wire n_636;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_570;
wire n_28;
wire n_606;
wire n_245;
wire n_451;
wire n_626;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_597;
wire n_618;
wire n_609;
wire n_94;
wire n_645;
wire n_687;
wire n_547;
wire n_309;
wire n_294;
wire n_619;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_588;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_540;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_567;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_530;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_549;
wire n_70;
wire n_568;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_580;
wire n_144;
wire n_130;
wire n_641;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_676;
wire n_187;
wire n_436;
wire n_629;
wire n_88;
wire n_169;
wire n_167;
wire n_659;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_660;
wire n_210;
wire n_206;
wire n_552;
wire n_408;
wire n_85;
wire n_591;
wire n_625;
wire n_96;
wire n_665;
wire n_308;
wire n_433;
wire n_364;

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_0),
.Y(n_134)
);

BUFx12f_ASAP7_75t_L g144 ( 
.A(n_0),
.Y(n_144)
);

HB1xp67_ASAP7_75t_L g254 ( 
.A(n_0),
.Y(n_254)
);

INVx2_ASAP7_75t_L g347 ( 
.A(n_0),
.Y(n_347)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_1),
.A2(n_96),
.B1(n_101),
.B2(n_102),
.Y(n_95)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_1),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g209 ( 
.A1(n_1),
.A2(n_101),
.B1(n_210),
.B2(n_214),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_1),
.A2(n_101),
.B1(n_276),
.B2(n_282),
.Y(n_275)
);

AOI22xp33_ASAP7_75t_L g636 ( 
.A1(n_1),
.A2(n_101),
.B1(n_637),
.B2(n_638),
.Y(n_636)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_2),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_L g23 ( 
.A1(n_3),
.A2(n_24),
.B1(n_25),
.B2(n_32),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_3),
.A2(n_24),
.B1(n_126),
.B2(n_128),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_L g256 ( 
.A1(n_3),
.A2(n_24),
.B1(n_257),
.B2(n_260),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g616 ( 
.A1(n_3),
.A2(n_24),
.B1(n_617),
.B2(n_621),
.Y(n_616)
);

OAI22xp5_ASAP7_75t_L g59 ( 
.A1(n_4),
.A2(n_60),
.B1(n_61),
.B2(n_65),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_4),
.Y(n_60)
);

AO22x1_ASAP7_75t_L g139 ( 
.A1(n_4),
.A2(n_60),
.B1(n_140),
.B2(n_141),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g291 ( 
.A1(n_4),
.A2(n_60),
.B1(n_260),
.B2(n_292),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_L g645 ( 
.A1(n_4),
.A2(n_60),
.B1(n_646),
.B2(n_648),
.Y(n_645)
);

OAI22xp5_ASAP7_75t_L g242 ( 
.A1(n_5),
.A2(n_243),
.B1(n_244),
.B2(n_247),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_5),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g395 ( 
.A1(n_5),
.A2(n_243),
.B1(n_396),
.B2(n_399),
.Y(n_395)
);

AOI22xp33_ASAP7_75t_SL g495 ( 
.A1(n_5),
.A2(n_243),
.B1(n_260),
.B2(n_496),
.Y(n_495)
);

AOI22xp33_ASAP7_75t_L g536 ( 
.A1(n_5),
.A2(n_243),
.B1(n_537),
.B2(n_540),
.Y(n_536)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_6),
.A2(n_171),
.B1(n_175),
.B2(n_176),
.Y(n_170)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_6),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_6),
.A2(n_175),
.B1(n_221),
.B2(n_225),
.Y(n_220)
);

OAI22xp33_ASAP7_75t_L g305 ( 
.A1(n_6),
.A2(n_175),
.B1(n_194),
.B2(n_306),
.Y(n_305)
);

AOI22x1_ASAP7_75t_L g409 ( 
.A1(n_6),
.A2(n_175),
.B1(n_410),
.B2(n_412),
.Y(n_409)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_7),
.A2(n_194),
.B1(n_197),
.B2(n_202),
.Y(n_193)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_7),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g320 ( 
.A1(n_7),
.A2(n_202),
.B1(n_321),
.B2(n_326),
.Y(n_320)
);

AOI22xp33_ASAP7_75t_SL g478 ( 
.A1(n_7),
.A2(n_202),
.B1(n_260),
.B2(n_479),
.Y(n_478)
);

AOI22xp33_ASAP7_75t_SL g517 ( 
.A1(n_7),
.A2(n_202),
.B1(n_518),
.B2(n_522),
.Y(n_517)
);

AOI22xp5_ASAP7_75t_L g19 ( 
.A1(n_8),
.A2(n_15),
.B1(n_20),
.B2(n_687),
.Y(n_19)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_9),
.A2(n_115),
.B1(n_116),
.B2(n_119),
.Y(n_114)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_9),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_9),
.A2(n_54),
.B1(n_115),
.B2(n_180),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g337 ( 
.A1(n_9),
.A2(n_115),
.B1(n_338),
.B2(n_339),
.Y(n_337)
);

OAI22xp5_ASAP7_75t_SL g609 ( 
.A1(n_9),
.A2(n_115),
.B1(n_244),
.B2(n_610),
.Y(n_609)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_10),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_10),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g151 ( 
.A(n_11),
.Y(n_151)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_11),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_12),
.Y(n_85)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_12),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_12),
.Y(n_137)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_12),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_L g366 ( 
.A(n_13),
.B(n_367),
.Y(n_366)
);

CKINVDCx20_ASAP7_75t_R g380 ( 
.A(n_13),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_13),
.B(n_67),
.Y(n_406)
);

OAI32xp33_ASAP7_75t_L g447 ( 
.A1(n_13),
.A2(n_448),
.A3(n_451),
.B1(n_453),
.B2(n_461),
.Y(n_447)
);

AOI22xp33_ASAP7_75t_SL g500 ( 
.A1(n_13),
.A2(n_380),
.B1(n_501),
.B2(n_502),
.Y(n_500)
);

OAI21xp33_ASAP7_75t_L g575 ( 
.A1(n_13),
.A2(n_131),
.B(n_527),
.Y(n_575)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_14),
.Y(n_88)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_14),
.Y(n_111)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_14),
.Y(n_556)
);

INVx1_ASAP7_75t_SL g687 ( 
.A(n_15),
.Y(n_687)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_16),
.A2(n_27),
.B1(n_187),
.B2(n_188),
.Y(n_186)
);

INVx1_ASAP7_75t_SL g187 ( 
.A(n_16),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_16),
.A2(n_54),
.B1(n_187),
.B2(n_232),
.Y(n_231)
);

OAI22x1_ASAP7_75t_SL g384 ( 
.A1(n_16),
.A2(n_187),
.B1(n_385),
.B2(n_389),
.Y(n_384)
);

OAI22xp5_ASAP7_75t_SL g469 ( 
.A1(n_16),
.A2(n_187),
.B1(n_470),
.B2(n_474),
.Y(n_469)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_17),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_17),
.Y(n_105)
);

BUFx3_ASAP7_75t_L g123 ( 
.A(n_17),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g159 ( 
.A(n_17),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_18),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_18),
.Y(n_55)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_18),
.Y(n_174)
);

BUFx6f_ASAP7_75t_L g281 ( 
.A(n_18),
.Y(n_281)
);

AOI21xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_70),
.B(n_684),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_68),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g676 ( 
.A(n_22),
.B(n_677),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_L g683 ( 
.A(n_22),
.B(n_677),
.Y(n_683)
);

INVxp67_ASAP7_75t_L g686 ( 
.A(n_22),
.Y(n_686)
);

AOI22xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_36),
.B1(n_59),
.B2(n_66),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_L g669 ( 
.A1(n_23),
.A2(n_36),
.B1(n_66),
.B2(n_670),
.Y(n_669)
);

INVxp67_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVx3_ASAP7_75t_SL g27 ( 
.A(n_28),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_29),
.Y(n_246)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g308 ( 
.A(n_31),
.Y(n_308)
);

INVx2_ASAP7_75t_SL g32 ( 
.A(n_33),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx4_ASAP7_75t_SL g39 ( 
.A(n_34),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_35),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g191 ( 
.A(n_35),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_L g69 ( 
.A1(n_36),
.A2(n_59),
.B(n_66),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_SL g608 ( 
.A1(n_36),
.A2(n_66),
.B1(n_305),
.B2(n_609),
.Y(n_608)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_36),
.Y(n_640)
);

HB1xp67_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_37),
.B(n_193),
.Y(n_192)
);

AO22x1_ASAP7_75t_L g241 ( 
.A1(n_37),
.A2(n_67),
.B1(n_193),
.B2(n_242),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_SL g303 ( 
.A(n_37),
.B(n_186),
.Y(n_303)
);

OAI21xp33_ASAP7_75t_L g377 ( 
.A1(n_37),
.A2(n_366),
.B(n_378),
.Y(n_377)
);

AND2x2_ASAP7_75t_L g37 ( 
.A(n_38),
.B(n_48),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_L g38 ( 
.A1(n_39),
.A2(n_40),
.B1(n_44),
.B2(n_46),
.Y(n_38)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx2_ASAP7_75t_L g355 ( 
.A(n_42),
.Y(n_355)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_43),
.Y(n_47)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_43),
.Y(n_50)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_43),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g365 ( 
.A(n_43),
.Y(n_365)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_48),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g48 ( 
.A1(n_49),
.A2(n_51),
.B1(n_54),
.B2(n_56),
.Y(n_48)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_51),
.Y(n_502)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_52),
.Y(n_169)
);

INVx2_ASAP7_75t_L g650 ( 
.A(n_52),
.Y(n_650)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g162 ( 
.A(n_53),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g183 ( 
.A(n_53),
.Y(n_183)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_53),
.Y(n_236)
);

BUFx6f_ASAP7_75t_L g325 ( 
.A(n_53),
.Y(n_325)
);

BUFx12f_ASAP7_75t_L g452 ( 
.A(n_53),
.Y(n_452)
);

INVx2_ASAP7_75t_L g362 ( 
.A(n_54),
.Y(n_362)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g398 ( 
.A(n_55),
.Y(n_398)
);

INVx8_ASAP7_75t_L g620 ( 
.A(n_55),
.Y(n_620)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_61),
.Y(n_65)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g196 ( 
.A(n_64),
.Y(n_196)
);

INVx3_ASAP7_75t_L g201 ( 
.A(n_64),
.Y(n_201)
);

BUFx3_ASAP7_75t_L g248 ( 
.A(n_64),
.Y(n_248)
);

BUFx6f_ASAP7_75t_L g612 ( 
.A(n_64),
.Y(n_612)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_66),
.Y(n_639)
);

HB1xp67_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_67),
.B(n_186),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_67),
.B(n_305),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_67),
.B(n_242),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_69),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g685 ( 
.A(n_69),
.B(n_686),
.Y(n_685)
);

AO21x2_ASAP7_75t_L g70 ( 
.A1(n_71),
.A2(n_602),
.B(n_678),
.Y(n_70)
);

NAND2x1_ASAP7_75t_L g71 ( 
.A(n_72),
.B(n_437),
.Y(n_71)
);

AOI21xp5_ASAP7_75t_L g72 ( 
.A1(n_73),
.A2(n_372),
.B(n_433),
.Y(n_72)
);

INVxp67_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g599 ( 
.A(n_74),
.B(n_600),
.Y(n_599)
);

OAI21xp5_ASAP7_75t_SL g74 ( 
.A1(n_75),
.A2(n_262),
.B(n_309),
.Y(n_74)
);

NOR2xp67_ASAP7_75t_L g434 ( 
.A(n_75),
.B(n_262),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g436 ( 
.A(n_75),
.B(n_262),
.Y(n_436)
);

MAJx2_ASAP7_75t_L g75 ( 
.A(n_76),
.B(n_203),
.C(n_249),
.Y(n_75)
);

HB1xp67_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g370 ( 
.A1(n_77),
.A2(n_78),
.B1(n_249),
.B2(n_371),
.Y(n_370)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

XNOR2xp5_ASAP7_75t_L g78 ( 
.A(n_79),
.B(n_145),
.Y(n_78)
);

INVxp33_ASAP7_75t_L g265 ( 
.A(n_79),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_80),
.B(n_124),
.Y(n_79)
);

XOR2xp5_ASAP7_75t_L g313 ( 
.A(n_80),
.B(n_124),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_81),
.A2(n_95),
.B1(n_106),
.B2(n_114),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g219 ( 
.A1(n_81),
.A2(n_106),
.B1(n_114),
.B2(n_220),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_L g255 ( 
.A1(n_81),
.A2(n_95),
.B1(n_106),
.B2(n_256),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_SL g494 ( 
.A1(n_81),
.A2(n_106),
.B1(n_478),
.B2(n_495),
.Y(n_494)
);

INVxp67_ASAP7_75t_R g81 ( 
.A(n_82),
.Y(n_81)
);

OR2x2_ASAP7_75t_L g106 ( 
.A(n_82),
.B(n_107),
.Y(n_106)
);

INVxp33_ASAP7_75t_L g297 ( 
.A(n_82),
.Y(n_297)
);

OAI22x1_ASAP7_75t_L g82 ( 
.A1(n_83),
.A2(n_86),
.B1(n_89),
.B2(n_92),
.Y(n_82)
);

INVx3_ASAP7_75t_L g558 ( 
.A(n_83),
.Y(n_558)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_84),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

BUFx2_ASAP7_75t_L g127 ( 
.A(n_85),
.Y(n_127)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_85),
.Y(n_411)
);

INVx2_ASAP7_75t_L g415 ( 
.A(n_85),
.Y(n_415)
);

INVx2_ASAP7_75t_L g550 ( 
.A(n_85),
.Y(n_550)
);

AOI22xp33_ASAP7_75t_L g107 ( 
.A1(n_86),
.A2(n_108),
.B1(n_109),
.B2(n_112),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_88),
.Y(n_91)
);

INVx4_ASAP7_75t_L g560 ( 
.A(n_88),
.Y(n_560)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVx2_ASAP7_75t_L g474 ( 
.A(n_92),
.Y(n_474)
);

BUFx12f_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_93),
.Y(n_130)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g142 ( 
.A(n_94),
.Y(n_142)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_99),
.Y(n_118)
);

BUFx5_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g295 ( 
.A(n_100),
.Y(n_295)
);

BUFx3_ASAP7_75t_L g392 ( 
.A(n_100),
.Y(n_392)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_102),
.Y(n_260)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_105),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_105),
.Y(n_113)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_105),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g224 ( 
.A(n_105),
.Y(n_224)
);

BUFx6f_ASAP7_75t_L g259 ( 
.A(n_105),
.Y(n_259)
);

INVx2_ASAP7_75t_SL g290 ( 
.A(n_106),
.Y(n_290)
);

HB1xp67_ASAP7_75t_L g477 ( 
.A(n_106),
.Y(n_477)
);

HB1xp67_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g551 ( 
.A(n_119),
.B(n_552),
.Y(n_551)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

BUFx4f_ASAP7_75t_SL g120 ( 
.A(n_121),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g227 ( 
.A(n_123),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_125),
.A2(n_131),
.B1(n_138),
.B2(n_143),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g207 ( 
.A1(n_125),
.A2(n_131),
.B1(n_208),
.B2(n_217),
.Y(n_207)
);

INVx2_ASAP7_75t_SL g126 ( 
.A(n_127),
.Y(n_126)
);

BUFx3_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g408 ( 
.A1(n_131),
.A2(n_337),
.B1(n_409),
.B2(n_416),
.Y(n_408)
);

OAI21x1_ASAP7_75t_SL g516 ( 
.A1(n_131),
.A2(n_517),
.B(n_527),
.Y(n_516)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

OA21x2_ASAP7_75t_L g252 ( 
.A1(n_132),
.A2(n_139),
.B(n_253),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_SL g335 ( 
.A(n_132),
.B(n_336),
.Y(n_335)
);

AOI22xp33_ASAP7_75t_SL g419 ( 
.A1(n_132),
.A2(n_209),
.B1(n_336),
.B2(n_344),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g468 ( 
.A(n_132),
.B(n_469),
.Y(n_468)
);

AOI22xp5_ASAP7_75t_L g534 ( 
.A1(n_132),
.A2(n_417),
.B1(n_535),
.B2(n_544),
.Y(n_534)
);

AND2x4_ASAP7_75t_L g132 ( 
.A(n_133),
.B(n_135),
.Y(n_132)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g218 ( 
.A(n_134),
.Y(n_218)
);

BUFx3_ASAP7_75t_L g467 ( 
.A(n_134),
.Y(n_467)
);

BUFx6f_ASAP7_75t_L g529 ( 
.A(n_134),
.Y(n_529)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g213 ( 
.A(n_136),
.Y(n_213)
);

INVx6_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

INVx2_ASAP7_75t_L g473 ( 
.A(n_137),
.Y(n_473)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_137),
.Y(n_539)
);

BUFx6f_ASAP7_75t_L g543 ( 
.A(n_137),
.Y(n_543)
);

BUFx6f_ASAP7_75t_L g585 ( 
.A(n_137),
.Y(n_585)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

HB1xp67_ASAP7_75t_L g216 ( 
.A(n_142),
.Y(n_216)
);

INVx2_ASAP7_75t_L g338 ( 
.A(n_142),
.Y(n_338)
);

INVx5_ASAP7_75t_L g417 ( 
.A(n_143),
.Y(n_417)
);

INVx8_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

XOR2xp5_ASAP7_75t_L g145 ( 
.A(n_146),
.B(n_184),
.Y(n_145)
);

INVxp67_ASAP7_75t_SL g267 ( 
.A(n_146),
.Y(n_267)
);

AOI22x1_ASAP7_75t_L g146 ( 
.A1(n_147),
.A2(n_170),
.B1(n_178),
.B2(n_179),
.Y(n_146)
);

INVx3_ASAP7_75t_SL g237 ( 
.A(n_147),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_147),
.A2(n_179),
.B1(n_275),
.B2(n_287),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_SL g393 ( 
.A1(n_147),
.A2(n_287),
.B1(n_394),
.B2(n_395),
.Y(n_393)
);

NAND2xp33_ASAP7_75t_SL g404 ( 
.A(n_147),
.B(n_231),
.Y(n_404)
);

AOI22xp5_ASAP7_75t_L g615 ( 
.A1(n_147),
.A2(n_275),
.B1(n_287),
.B2(n_616),
.Y(n_615)
);

AOI22xp5_ASAP7_75t_L g644 ( 
.A1(n_147),
.A2(n_287),
.B1(n_616),
.B2(n_645),
.Y(n_644)
);

AND2x2_ASAP7_75t_L g147 ( 
.A(n_148),
.B(n_160),
.Y(n_147)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_148),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_R g514 ( 
.A(n_148),
.B(n_380),
.Y(n_514)
);

AOI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_149),
.A2(n_152),
.B1(n_154),
.B2(n_157),
.Y(n_148)
);

INVx5_ASAP7_75t_SL g149 ( 
.A(n_150),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g167 ( 
.A(n_151),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g460 ( 
.A(n_151),
.Y(n_460)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

INVx3_ASAP7_75t_L g498 ( 
.A(n_153),
.Y(n_498)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

INVx4_ASAP7_75t_L g165 ( 
.A(n_155),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

INVx5_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g450 ( 
.A(n_159),
.Y(n_450)
);

INVx2_ASAP7_75t_L g482 ( 
.A(n_159),
.Y(n_482)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_161),
.A2(n_163),
.B1(n_166),
.B2(n_168),
.Y(n_160)
);

BUFx4f_ASAP7_75t_L g501 ( 
.A(n_161),
.Y(n_501)
);

INVx2_ASAP7_75t_SL g161 ( 
.A(n_162),
.Y(n_161)
);

INVx2_ASAP7_75t_SL g163 ( 
.A(n_164),
.Y(n_163)
);

INVx3_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

INVx3_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_170),
.Y(n_238)
);

BUFx3_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_173),
.Y(n_177)
);

BUFx5_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

BUFx6f_ASAP7_75t_L g286 ( 
.A(n_174),
.Y(n_286)
);

BUFx3_ASAP7_75t_L g331 ( 
.A(n_174),
.Y(n_331)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_178),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_178),
.B(n_231),
.Y(n_332)
);

INVx2_ASAP7_75t_L g647 ( 
.A(n_180),
.Y(n_647)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

INVxp67_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_182),
.Y(n_400)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

HB1xp67_ASAP7_75t_L g269 ( 
.A(n_184),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_192),
.Y(n_184)
);

AND2x2_ASAP7_75t_L g376 ( 
.A(n_185),
.B(n_377),
.Y(n_376)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

INVx4_ASAP7_75t_SL g190 ( 
.A(n_191),
.Y(n_190)
);

BUFx3_ASAP7_75t_L g638 ( 
.A(n_191),
.Y(n_638)
);

INVx11_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

BUFx12f_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

INVx2_ASAP7_75t_SL g637 ( 
.A(n_197),
.Y(n_637)
);

BUFx3_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

INVxp67_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_199),
.Y(n_368)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_L g369 ( 
.A(n_204),
.B(n_370),
.Y(n_369)
);

MAJx2_ASAP7_75t_L g204 ( 
.A(n_205),
.B(n_228),
.C(n_240),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

XNOR2x1_ASAP7_75t_L g311 ( 
.A(n_206),
.B(n_312),
.Y(n_311)
);

AND2x2_ASAP7_75t_L g206 ( 
.A(n_207),
.B(n_219),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_SL g423 ( 
.A(n_207),
.B(n_219),
.Y(n_423)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

NAND2xp33_ASAP7_75t_R g343 ( 
.A(n_209),
.B(n_344),
.Y(n_343)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

INVx8_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_220),
.Y(n_383)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

INVx2_ASAP7_75t_SL g222 ( 
.A(n_223),
.Y(n_222)
);

INVx4_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

INVx4_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

INVxp33_ASAP7_75t_SL g228 ( 
.A(n_229),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g312 ( 
.A(n_229),
.B(n_241),
.Y(n_312)
);

OAI22x1_ASAP7_75t_L g229 ( 
.A1(n_230),
.A2(n_237),
.B1(n_238),
.B2(n_239),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

OAI21xp5_ASAP7_75t_L g319 ( 
.A1(n_237),
.A2(n_320),
.B(n_332),
.Y(n_319)
);

OAI21xp5_ASAP7_75t_SL g499 ( 
.A1(n_237),
.A2(n_332),
.B(n_500),
.Y(n_499)
);

AO21x1_ASAP7_75t_L g667 ( 
.A1(n_237),
.A2(n_239),
.B(n_668),
.Y(n_667)
);

INVx2_ASAP7_75t_L g287 ( 
.A(n_239),
.Y(n_287)
);

OAI21xp5_ASAP7_75t_SL g402 ( 
.A1(n_239),
.A2(n_403),
.B(n_404),
.Y(n_402)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

INVx4_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

INVx3_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

INVxp67_ASAP7_75t_SL g247 ( 
.A(n_248),
.Y(n_247)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_249),
.Y(n_371)
);

OAI22xp5_ASAP7_75t_L g249 ( 
.A1(n_250),
.A2(n_251),
.B1(n_255),
.B2(n_261),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g301 ( 
.A(n_250),
.B(n_302),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_L g630 ( 
.A1(n_250),
.A2(n_300),
.B1(n_631),
.B2(n_689),
.Y(n_630)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

AND2x2_ASAP7_75t_L g300 ( 
.A(n_251),
.B(n_255),
.Y(n_300)
);

BUFx4f_ASAP7_75t_SL g251 ( 
.A(n_252),
.Y(n_251)
);

INVx2_ASAP7_75t_L g572 ( 
.A(n_253),
.Y(n_572)
);

BUFx4f_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

INVxp67_ASAP7_75t_SL g261 ( 
.A(n_255),
.Y(n_261)
);

INVxp67_ASAP7_75t_L g289 ( 
.A(n_256),
.Y(n_289)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

BUFx2_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

XOR2x2_ASAP7_75t_L g262 ( 
.A(n_263),
.B(n_270),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g653 ( 
.A(n_263),
.B(n_654),
.C(n_655),
.Y(n_653)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_264),
.B(n_266),
.C(n_268),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_267),
.Y(n_266)
);

INVx1_ASAP7_75t_SL g268 ( 
.A(n_269),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_L g270 ( 
.A(n_271),
.B(n_299),
.Y(n_270)
);

HB1xp67_ASAP7_75t_L g655 ( 
.A(n_271),
.Y(n_655)
);

NAND2x1p5_ASAP7_75t_L g271 ( 
.A(n_272),
.B(n_298),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g605 ( 
.A(n_272),
.B(n_606),
.C(n_629),
.Y(n_605)
);

AOI22xp5_ASAP7_75t_L g658 ( 
.A1(n_272),
.A2(n_273),
.B1(n_608),
.B2(n_659),
.Y(n_658)
);

INVx3_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

AND2x2_ASAP7_75t_L g273 ( 
.A(n_274),
.B(n_288),
.Y(n_273)
);

OR2x2_ASAP7_75t_L g298 ( 
.A(n_274),
.B(n_288),
.Y(n_298)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

INVx4_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

BUFx6f_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

INVx2_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

INVx2_ASAP7_75t_L g359 ( 
.A(n_280),
.Y(n_359)
);

INVx8_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

INVx2_ASAP7_75t_SL g283 ( 
.A(n_284),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

INVx2_ASAP7_75t_SL g285 ( 
.A(n_286),
.Y(n_285)
);

INVx4_ASAP7_75t_L g456 ( 
.A(n_286),
.Y(n_456)
);

INVx2_ASAP7_75t_L g623 ( 
.A(n_286),
.Y(n_623)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_289),
.A2(n_290),
.B1(n_291),
.B2(n_296),
.Y(n_288)
);

AOI22x1_ASAP7_75t_L g382 ( 
.A1(n_290),
.A2(n_296),
.B1(n_383),
.B2(n_384),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g512 ( 
.A(n_290),
.B(n_384),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_L g564 ( 
.A(n_290),
.B(n_565),
.Y(n_564)
);

OA21x2_ASAP7_75t_L g625 ( 
.A1(n_290),
.A2(n_291),
.B(n_296),
.Y(n_625)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

HB1xp67_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

INVx2_ASAP7_75t_L g388 ( 
.A(n_295),
.Y(n_388)
);

INVx3_ASAP7_75t_L g464 ( 
.A(n_295),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_L g483 ( 
.A(n_296),
.B(n_384),
.Y(n_483)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_296),
.Y(n_510)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_297),
.Y(n_296)
);

HB1xp67_ASAP7_75t_L g654 ( 
.A(n_299),
.Y(n_654)
);

XNOR2xp5_ASAP7_75t_L g299 ( 
.A(n_300),
.B(n_301),
.Y(n_299)
);

HB1xp67_ASAP7_75t_L g631 ( 
.A(n_302),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_SL g302 ( 
.A(n_303),
.B(n_304),
.Y(n_302)
);

NAND2xp33_ASAP7_75t_SL g316 ( 
.A(n_303),
.B(n_317),
.Y(n_316)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

INVx1_ASAP7_75t_SL g307 ( 
.A(n_308),
.Y(n_307)
);

INVx2_ASAP7_75t_L g352 ( 
.A(n_308),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_310),
.B(n_369),
.Y(n_309)
);

OR2x2_ASAP7_75t_L g435 ( 
.A(n_310),
.B(n_369),
.Y(n_435)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_311),
.B(n_313),
.C(n_314),
.Y(n_310)
);

XNOR2x1_ASAP7_75t_L g432 ( 
.A(n_311),
.B(n_313),
.Y(n_432)
);

XNOR2x1_ASAP7_75t_L g431 ( 
.A(n_314),
.B(n_432),
.Y(n_431)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_315),
.B(n_318),
.C(n_333),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_L g425 ( 
.A1(n_315),
.A2(n_316),
.B1(n_318),
.B2(n_319),
.Y(n_425)
);

INVxp67_ASAP7_75t_SL g315 ( 
.A(n_316),
.Y(n_315)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_319),
.Y(n_318)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_320),
.Y(n_394)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_322),
.Y(n_321)
);

HB1xp67_ASAP7_75t_L g322 ( 
.A(n_323),
.Y(n_322)
);

INVx3_ASAP7_75t_L g323 ( 
.A(n_324),
.Y(n_323)
);

INVx2_ASAP7_75t_L g324 ( 
.A(n_325),
.Y(n_324)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_327),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_328),
.Y(n_327)
);

INVxp67_ASAP7_75t_L g328 ( 
.A(n_329),
.Y(n_328)
);

INVx3_ASAP7_75t_L g329 ( 
.A(n_330),
.Y(n_329)
);

INVx2_ASAP7_75t_L g330 ( 
.A(n_331),
.Y(n_330)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_334),
.Y(n_333)
);

XNOR2xp5_ASAP7_75t_L g424 ( 
.A(n_334),
.B(n_425),
.Y(n_424)
);

AOI21xp5_ASAP7_75t_L g334 ( 
.A1(n_335),
.A2(n_343),
.B(n_348),
.Y(n_334)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_337),
.Y(n_336)
);

BUFx2_ASAP7_75t_L g339 ( 
.A(n_340),
.Y(n_339)
);

INVx2_ASAP7_75t_L g340 ( 
.A(n_341),
.Y(n_340)
);

INVx2_ASAP7_75t_L g341 ( 
.A(n_342),
.Y(n_341)
);

INVx2_ASAP7_75t_L g526 ( 
.A(n_342),
.Y(n_526)
);

INVx4_ASAP7_75t_L g344 ( 
.A(n_345),
.Y(n_344)
);

INVx2_ASAP7_75t_SL g345 ( 
.A(n_346),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_347),
.Y(n_346)
);

XOR2xp5_ASAP7_75t_L g418 ( 
.A(n_348),
.B(n_419),
.Y(n_418)
);

AOI32xp33_ASAP7_75t_L g348 ( 
.A1(n_349),
.A2(n_353),
.A3(n_356),
.B1(n_360),
.B2(n_366),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_350),
.Y(n_349)
);

INVx2_ASAP7_75t_L g350 ( 
.A(n_351),
.Y(n_350)
);

INVx2_ASAP7_75t_L g351 ( 
.A(n_352),
.Y(n_351)
);

INVx1_ASAP7_75t_SL g353 ( 
.A(n_354),
.Y(n_353)
);

INVx2_ASAP7_75t_L g354 ( 
.A(n_355),
.Y(n_354)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_357),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_358),
.Y(n_357)
);

INVx2_ASAP7_75t_L g358 ( 
.A(n_359),
.Y(n_358)
);

NAND2xp33_ASAP7_75t_SL g360 ( 
.A(n_361),
.B(n_363),
.Y(n_360)
);

INVx1_ASAP7_75t_SL g361 ( 
.A(n_362),
.Y(n_361)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_364),
.Y(n_363)
);

INVx2_ASAP7_75t_L g364 ( 
.A(n_365),
.Y(n_364)
);

INVx2_ASAP7_75t_L g379 ( 
.A(n_367),
.Y(n_379)
);

INVx2_ASAP7_75t_L g367 ( 
.A(n_368),
.Y(n_367)
);

MAJIxp5_ASAP7_75t_L g372 ( 
.A(n_373),
.B(n_426),
.C(n_430),
.Y(n_372)
);

OR2x2_ASAP7_75t_L g373 ( 
.A(n_374),
.B(n_420),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g601 ( 
.A(n_374),
.B(n_420),
.Y(n_601)
);

MAJIxp5_ASAP7_75t_L g374 ( 
.A(n_375),
.B(n_401),
.C(n_418),
.Y(n_374)
);

XNOR2xp5_ASAP7_75t_L g484 ( 
.A(n_375),
.B(n_485),
.Y(n_484)
);

XOR2xp5_ASAP7_75t_L g375 ( 
.A(n_376),
.B(n_381),
.Y(n_375)
);

MAJx2_ASAP7_75t_L g422 ( 
.A(n_376),
.B(n_382),
.C(n_393),
.Y(n_422)
);

NOR2xp33_ASAP7_75t_L g378 ( 
.A(n_379),
.B(n_380),
.Y(n_378)
);

NOR2xp33_ASAP7_75t_L g461 ( 
.A(n_380),
.B(n_462),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_L g561 ( 
.A(n_380),
.B(n_562),
.Y(n_561)
);

OAI21xp33_ASAP7_75t_L g565 ( 
.A1(n_380),
.A2(n_561),
.B(n_566),
.Y(n_565)
);

NOR2xp33_ASAP7_75t_SL g573 ( 
.A(n_380),
.B(n_510),
.Y(n_573)
);

NOR2xp33_ASAP7_75t_L g577 ( 
.A(n_380),
.B(n_578),
.Y(n_577)
);

XNOR2xp5_ASAP7_75t_L g381 ( 
.A(n_382),
.B(n_393),
.Y(n_381)
);

BUFx3_ASAP7_75t_L g385 ( 
.A(n_386),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_387),
.Y(n_386)
);

INVx2_ASAP7_75t_L g387 ( 
.A(n_388),
.Y(n_387)
);

INVx3_ASAP7_75t_L g566 ( 
.A(n_389),
.Y(n_566)
);

INVx3_ASAP7_75t_L g389 ( 
.A(n_390),
.Y(n_389)
);

INVx4_ASAP7_75t_L g390 ( 
.A(n_391),
.Y(n_390)
);

BUFx3_ASAP7_75t_L g391 ( 
.A(n_392),
.Y(n_391)
);

INVx5_ASAP7_75t_L g562 ( 
.A(n_392),
.Y(n_562)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_395),
.Y(n_403)
);

INVx5_ASAP7_75t_L g396 ( 
.A(n_397),
.Y(n_396)
);

INVx8_ASAP7_75t_L g397 ( 
.A(n_398),
.Y(n_397)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_400),
.Y(n_399)
);

XOR2xp5_ASAP7_75t_L g485 ( 
.A(n_401),
.B(n_418),
.Y(n_485)
);

MAJx2_ASAP7_75t_L g401 ( 
.A(n_402),
.B(n_405),
.C(n_407),
.Y(n_401)
);

XNOR2xp5_ASAP7_75t_SL g443 ( 
.A(n_402),
.B(n_444),
.Y(n_443)
);

AOI22xp5_ASAP7_75t_L g444 ( 
.A1(n_405),
.A2(n_406),
.B1(n_408),
.B2(n_445),
.Y(n_444)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_406),
.Y(n_405)
);

HB1xp67_ASAP7_75t_L g407 ( 
.A(n_408),
.Y(n_407)
);

INVxp67_ASAP7_75t_L g445 ( 
.A(n_408),
.Y(n_445)
);

OAI21xp5_ASAP7_75t_L g465 ( 
.A1(n_409),
.A2(n_466),
.B(n_468),
.Y(n_465)
);

INVx2_ASAP7_75t_L g410 ( 
.A(n_411),
.Y(n_410)
);

INVx3_ASAP7_75t_L g412 ( 
.A(n_413),
.Y(n_412)
);

BUFx2_ASAP7_75t_SL g413 ( 
.A(n_414),
.Y(n_413)
);

INVx2_ASAP7_75t_L g414 ( 
.A(n_415),
.Y(n_414)
);

INVx4_ASAP7_75t_L g521 ( 
.A(n_415),
.Y(n_521)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_417),
.Y(n_416)
);

XNOR2xp5_ASAP7_75t_L g420 ( 
.A(n_421),
.B(n_424),
.Y(n_420)
);

XNOR2xp5_ASAP7_75t_L g421 ( 
.A(n_422),
.B(n_423),
.Y(n_421)
);

HB1xp67_ASAP7_75t_L g428 ( 
.A(n_422),
.Y(n_428)
);

HB1xp67_ASAP7_75t_L g429 ( 
.A(n_423),
.Y(n_429)
);

MAJIxp5_ASAP7_75t_L g427 ( 
.A(n_424),
.B(n_428),
.C(n_429),
.Y(n_427)
);

INVx1_ASAP7_75t_SL g426 ( 
.A(n_427),
.Y(n_426)
);

OAI21xp5_ASAP7_75t_L g600 ( 
.A1(n_427),
.A2(n_431),
.B(n_601),
.Y(n_600)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_431),
.Y(n_430)
);

OAI21xp5_ASAP7_75t_L g433 ( 
.A1(n_434),
.A2(n_435),
.B(n_436),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_438),
.B(n_599),
.Y(n_437)
);

OAI21x1_ASAP7_75t_L g438 ( 
.A1(n_439),
.A2(n_486),
.B(n_597),
.Y(n_438)
);

AND2x2_ASAP7_75t_L g439 ( 
.A(n_440),
.B(n_484),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_441),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_L g597 ( 
.A(n_441),
.B(n_598),
.Y(n_597)
);

MAJIxp5_ASAP7_75t_L g441 ( 
.A(n_442),
.B(n_446),
.C(n_475),
.Y(n_441)
);

INVxp67_ASAP7_75t_L g442 ( 
.A(n_443),
.Y(n_442)
);

XNOR2xp5_ASAP7_75t_L g489 ( 
.A(n_443),
.B(n_490),
.Y(n_489)
);

OAI22xp5_ASAP7_75t_L g490 ( 
.A1(n_446),
.A2(n_475),
.B1(n_476),
.B2(n_491),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_446),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_L g446 ( 
.A(n_447),
.B(n_465),
.Y(n_446)
);

XOR2xp5_ASAP7_75t_L g493 ( 
.A(n_447),
.B(n_465),
.Y(n_493)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_449),
.Y(n_448)
);

INVxp67_ASAP7_75t_L g449 ( 
.A(n_450),
.Y(n_449)
);

INVx4_ASAP7_75t_L g451 ( 
.A(n_452),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_454),
.B(n_457),
.Y(n_453)
);

INVx3_ASAP7_75t_L g454 ( 
.A(n_455),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_456),
.Y(n_455)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_458),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_459),
.Y(n_458)
);

INVx3_ASAP7_75t_L g459 ( 
.A(n_460),
.Y(n_459)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_463),
.Y(n_462)
);

HB1xp67_ASAP7_75t_L g463 ( 
.A(n_464),
.Y(n_463)
);

INVx3_ASAP7_75t_L g466 ( 
.A(n_467),
.Y(n_466)
);

OAI21xp5_ASAP7_75t_SL g571 ( 
.A1(n_468),
.A2(n_536),
.B(n_572),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_L g527 ( 
.A(n_469),
.B(n_528),
.Y(n_527)
);

INVx2_ASAP7_75t_L g470 ( 
.A(n_471),
.Y(n_470)
);

INVx2_ASAP7_75t_L g471 ( 
.A(n_472),
.Y(n_471)
);

INVx2_ASAP7_75t_L g472 ( 
.A(n_473),
.Y(n_472)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_476),
.Y(n_475)
);

OAI21xp33_ASAP7_75t_SL g476 ( 
.A1(n_477),
.A2(n_478),
.B(n_483),
.Y(n_476)
);

INVx2_ASAP7_75t_L g479 ( 
.A(n_480),
.Y(n_479)
);

BUFx3_ASAP7_75t_L g480 ( 
.A(n_481),
.Y(n_480)
);

INVx2_ASAP7_75t_L g481 ( 
.A(n_482),
.Y(n_481)
);

AND2x2_ASAP7_75t_L g563 ( 
.A(n_483),
.B(n_564),
.Y(n_563)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_484),
.Y(n_598)
);

AOI21x1_ASAP7_75t_L g486 ( 
.A1(n_487),
.A2(n_530),
.B(n_596),
.Y(n_486)
);

AND2x2_ASAP7_75t_L g487 ( 
.A(n_488),
.B(n_503),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_SL g488 ( 
.A(n_489),
.B(n_492),
.Y(n_488)
);

NOR2xp33_ASAP7_75t_L g596 ( 
.A(n_489),
.B(n_492),
.Y(n_596)
);

MAJIxp5_ASAP7_75t_L g492 ( 
.A(n_493),
.B(n_494),
.C(n_499),
.Y(n_492)
);

XNOR2xp5_ASAP7_75t_L g504 ( 
.A(n_493),
.B(n_505),
.Y(n_504)
);

XNOR2xp5_ASAP7_75t_L g505 ( 
.A(n_494),
.B(n_499),
.Y(n_505)
);

HB1xp67_ASAP7_75t_L g511 ( 
.A(n_495),
.Y(n_511)
);

INVx1_ASAP7_75t_SL g496 ( 
.A(n_497),
.Y(n_496)
);

BUFx2_ASAP7_75t_L g497 ( 
.A(n_498),
.Y(n_497)
);

OR2x2_ASAP7_75t_L g503 ( 
.A(n_504),
.B(n_506),
.Y(n_503)
);

AND2x2_ASAP7_75t_L g594 ( 
.A(n_504),
.B(n_506),
.Y(n_594)
);

MAJIxp5_ASAP7_75t_L g506 ( 
.A(n_507),
.B(n_513),
.C(n_515),
.Y(n_506)
);

HB1xp67_ASAP7_75t_L g507 ( 
.A(n_508),
.Y(n_507)
);

OAI22xp5_ASAP7_75t_L g590 ( 
.A1(n_508),
.A2(n_509),
.B1(n_513),
.B2(n_514),
.Y(n_590)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_509),
.Y(n_508)
);

OAI21xp5_ASAP7_75t_L g509 ( 
.A1(n_510),
.A2(n_511),
.B(n_512),
.Y(n_509)
);

INVxp33_ASAP7_75t_L g513 ( 
.A(n_514),
.Y(n_513)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_516),
.Y(n_515)
);

XNOR2xp5_ASAP7_75t_L g589 ( 
.A(n_516),
.B(n_590),
.Y(n_589)
);

INVxp67_ASAP7_75t_L g544 ( 
.A(n_517),
.Y(n_544)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_519),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_520),
.Y(n_519)
);

INVx4_ASAP7_75t_L g520 ( 
.A(n_521),
.Y(n_520)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_523),
.Y(n_522)
);

HB1xp67_ASAP7_75t_L g523 ( 
.A(n_524),
.Y(n_523)
);

BUFx3_ASAP7_75t_L g524 ( 
.A(n_525),
.Y(n_524)
);

INVx2_ASAP7_75t_L g525 ( 
.A(n_526),
.Y(n_525)
);

BUFx2_ASAP7_75t_L g528 ( 
.A(n_529),
.Y(n_528)
);

BUFx2_ASAP7_75t_L g580 ( 
.A(n_529),
.Y(n_580)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_531),
.B(n_593),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_L g531 ( 
.A(n_532),
.B(n_587),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_L g532 ( 
.A(n_533),
.B(n_567),
.Y(n_532)
);

OR2x2_ASAP7_75t_L g533 ( 
.A(n_534),
.B(n_545),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_L g568 ( 
.A(n_534),
.B(n_545),
.Y(n_568)
);

INVxp67_ASAP7_75t_L g535 ( 
.A(n_536),
.Y(n_535)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_538),
.Y(n_537)
);

INVx2_ASAP7_75t_L g538 ( 
.A(n_539),
.Y(n_538)
);

BUFx2_ASAP7_75t_SL g540 ( 
.A(n_541),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_542),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_543),
.Y(n_542)
);

XNOR2xp5_ASAP7_75t_L g545 ( 
.A(n_546),
.B(n_563),
.Y(n_545)
);

NOR2xp33_ASAP7_75t_L g592 ( 
.A(n_546),
.B(n_563),
.Y(n_592)
);

AOI21xp33_ASAP7_75t_L g546 ( 
.A1(n_547),
.A2(n_551),
.B(n_557),
.Y(n_546)
);

BUFx2_ASAP7_75t_L g547 ( 
.A(n_548),
.Y(n_547)
);

INVx2_ASAP7_75t_L g548 ( 
.A(n_549),
.Y(n_548)
);

INVx4_ASAP7_75t_L g549 ( 
.A(n_550),
.Y(n_549)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_553),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_554),
.Y(n_553)
);

INVx3_ASAP7_75t_L g554 ( 
.A(n_555),
.Y(n_554)
);

BUFx3_ASAP7_75t_L g555 ( 
.A(n_556),
.Y(n_555)
);

AOI21xp5_ASAP7_75t_L g557 ( 
.A1(n_558),
.A2(n_559),
.B(n_561),
.Y(n_557)
);

BUFx3_ASAP7_75t_L g559 ( 
.A(n_560),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_L g567 ( 
.A(n_568),
.B(n_569),
.Y(n_567)
);

OAI21x1_ASAP7_75t_L g569 ( 
.A1(n_570),
.A2(n_574),
.B(n_586),
.Y(n_569)
);

NOR2xp33_ASAP7_75t_L g570 ( 
.A(n_571),
.B(n_573),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_SL g586 ( 
.A(n_571),
.B(n_573),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_SL g574 ( 
.A(n_575),
.B(n_576),
.Y(n_574)
);

NOR2xp33_ASAP7_75t_SL g576 ( 
.A(n_577),
.B(n_581),
.Y(n_576)
);

BUFx6f_ASAP7_75t_L g578 ( 
.A(n_579),
.Y(n_578)
);

INVx2_ASAP7_75t_L g579 ( 
.A(n_580),
.Y(n_579)
);

INVx1_ASAP7_75t_SL g581 ( 
.A(n_582),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_583),
.Y(n_582)
);

HB1xp67_ASAP7_75t_L g583 ( 
.A(n_584),
.Y(n_583)
);

INVx3_ASAP7_75t_L g584 ( 
.A(n_585),
.Y(n_584)
);

NAND2xp5_ASAP7_75t_L g587 ( 
.A(n_588),
.B(n_591),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_589),
.Y(n_588)
);

AND2x2_ASAP7_75t_L g595 ( 
.A(n_589),
.B(n_592),
.Y(n_595)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_592),
.Y(n_591)
);

NOR2x1_ASAP7_75t_SL g593 ( 
.A(n_594),
.B(n_595),
.Y(n_593)
);

NOR3xp33_ASAP7_75t_L g602 ( 
.A(n_603),
.B(n_660),
.C(n_676),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_SL g603 ( 
.A(n_604),
.B(n_652),
.Y(n_603)
);

A2O1A1Ixp33_ASAP7_75t_L g680 ( 
.A1(n_604),
.A2(n_661),
.B(n_681),
.C(n_682),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_L g604 ( 
.A(n_605),
.B(n_632),
.Y(n_604)
);

NOR2xp67_ASAP7_75t_SL g682 ( 
.A(n_605),
.B(n_632),
.Y(n_682)
);

OAI22xp5_ASAP7_75t_L g606 ( 
.A1(n_607),
.A2(n_613),
.B1(n_627),
.B2(n_628),
.Y(n_606)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_607),
.Y(n_627)
);

XOR2xp5_ASAP7_75t_L g633 ( 
.A(n_607),
.B(n_634),
.Y(n_633)
);

MAJIxp5_ASAP7_75t_L g651 ( 
.A(n_607),
.B(n_614),
.C(n_626),
.Y(n_651)
);

BUFx2_ASAP7_75t_L g607 ( 
.A(n_608),
.Y(n_607)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_608),
.Y(n_659)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_609),
.Y(n_641)
);

BUFx2_ASAP7_75t_L g610 ( 
.A(n_611),
.Y(n_610)
);

INVx3_ASAP7_75t_L g611 ( 
.A(n_612),
.Y(n_611)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_613),
.Y(n_628)
);

XNOR2xp5_ASAP7_75t_L g657 ( 
.A(n_613),
.B(n_658),
.Y(n_657)
);

AOI22xp5_ASAP7_75t_L g613 ( 
.A1(n_614),
.A2(n_615),
.B1(n_624),
.B2(n_626),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_615),
.Y(n_614)
);

INVx2_ASAP7_75t_L g617 ( 
.A(n_618),
.Y(n_617)
);

INVx2_ASAP7_75t_L g618 ( 
.A(n_619),
.Y(n_618)
);

INVx5_ASAP7_75t_L g619 ( 
.A(n_620),
.Y(n_619)
);

INVx3_ASAP7_75t_L g621 ( 
.A(n_622),
.Y(n_621)
);

BUFx3_ASAP7_75t_L g622 ( 
.A(n_623),
.Y(n_622)
);

OAI22xp5_ASAP7_75t_L g642 ( 
.A1(n_624),
.A2(n_625),
.B1(n_643),
.B2(n_644),
.Y(n_642)
);

MAJIxp5_ASAP7_75t_SL g663 ( 
.A(n_624),
.B(n_664),
.C(n_665),
.Y(n_663)
);

INVx2_ASAP7_75t_SL g624 ( 
.A(n_625),
.Y(n_624)
);

BUFx3_ASAP7_75t_L g626 ( 
.A(n_625),
.Y(n_626)
);

MAJIxp5_ASAP7_75t_L g673 ( 
.A(n_627),
.B(n_674),
.C(n_675),
.Y(n_673)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_630),
.Y(n_629)
);

XNOR2xp5_ASAP7_75t_L g656 ( 
.A(n_630),
.B(n_657),
.Y(n_656)
);

XNOR2xp5_ASAP7_75t_L g632 ( 
.A(n_633),
.B(n_651),
.Y(n_632)
);

HB1xp67_ASAP7_75t_L g674 ( 
.A(n_634),
.Y(n_674)
);

XNOR2xp5_ASAP7_75t_L g634 ( 
.A(n_635),
.B(n_642),
.Y(n_634)
);

OAI22x1_ASAP7_75t_SL g635 ( 
.A1(n_636),
.A2(n_639),
.B1(n_640),
.B2(n_641),
.Y(n_635)
);

OAI22xp5_ASAP7_75t_L g664 ( 
.A1(n_636),
.A2(n_639),
.B1(n_640),
.B2(n_641),
.Y(n_664)
);

INVxp67_ASAP7_75t_L g670 ( 
.A(n_636),
.Y(n_670)
);

HB1xp67_ASAP7_75t_L g665 ( 
.A(n_643),
.Y(n_665)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_644),
.Y(n_643)
);

INVxp67_ASAP7_75t_SL g668 ( 
.A(n_645),
.Y(n_668)
);

INVx2_ASAP7_75t_L g646 ( 
.A(n_647),
.Y(n_646)
);

INVx1_ASAP7_75t_SL g648 ( 
.A(n_649),
.Y(n_648)
);

BUFx3_ASAP7_75t_L g649 ( 
.A(n_650),
.Y(n_649)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_651),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_L g652 ( 
.A(n_653),
.B(n_656),
.Y(n_652)
);

NOR2xp33_ASAP7_75t_L g681 ( 
.A(n_653),
.B(n_656),
.Y(n_681)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_661),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_L g661 ( 
.A(n_662),
.B(n_673),
.Y(n_661)
);

OR2x2_ASAP7_75t_L g679 ( 
.A(n_662),
.B(n_673),
.Y(n_679)
);

XNOR2xp5_ASAP7_75t_L g662 ( 
.A(n_663),
.B(n_666),
.Y(n_662)
);

MAJIxp5_ASAP7_75t_L g677 ( 
.A(n_663),
.B(n_669),
.C(n_671),
.Y(n_677)
);

AOI22xp5_ASAP7_75t_SL g666 ( 
.A1(n_667),
.A2(n_669),
.B1(n_671),
.B2(n_672),
.Y(n_666)
);

CKINVDCx12_ASAP7_75t_R g671 ( 
.A(n_667),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_669),
.Y(n_672)
);

A2O1A1Ixp33_ASAP7_75t_L g678 ( 
.A1(n_676),
.A2(n_679),
.B(n_680),
.C(n_683),
.Y(n_678)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_685),
.Y(n_684)
);


endmodule