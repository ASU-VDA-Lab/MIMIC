module fake_jpeg_1154_n_176 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_176);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_176;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g43 ( 
.A(n_16),
.Y(n_43)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_18),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_41),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_25),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_20),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_28),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_27),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_34),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_4),
.Y(n_51)
);

BUFx5_ASAP7_75t_L g52 ( 
.A(n_31),
.Y(n_52)
);

INVx13_ASAP7_75t_L g53 ( 
.A(n_10),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_3),
.B(n_39),
.Y(n_54)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_24),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_20),
.Y(n_56)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_13),
.Y(n_57)
);

BUFx12_ASAP7_75t_L g58 ( 
.A(n_26),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_0),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_44),
.Y(n_60)
);

INVx5_ASAP7_75t_L g70 ( 
.A(n_60),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_45),
.B(n_50),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_61),
.B(n_63),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_46),
.Y(n_62)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_62),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_45),
.B(n_0),
.Y(n_63)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_57),
.Y(n_64)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_64),
.Y(n_78)
);

BUFx2_ASAP7_75t_L g65 ( 
.A(n_44),
.Y(n_65)
);

OR2x2_ASAP7_75t_L g77 ( 
.A(n_65),
.B(n_53),
.Y(n_77)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_57),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_66),
.B(n_55),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_65),
.A2(n_53),
.B1(n_46),
.B2(n_56),
.Y(n_67)
);

OA22x2_ASAP7_75t_L g90 ( 
.A1(n_67),
.A2(n_69),
.B1(n_58),
.B2(n_42),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_65),
.A2(n_53),
.B1(n_46),
.B2(n_56),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g71 ( 
.A1(n_64),
.A2(n_48),
.B1(n_51),
.B2(n_43),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_71),
.A2(n_73),
.B1(n_76),
.B2(n_47),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_72),
.B(n_40),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_66),
.A2(n_55),
.B1(n_51),
.B2(n_59),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_60),
.B(n_59),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g89 ( 
.A(n_74),
.B(n_58),
.Y(n_89)
);

OAI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_62),
.A2(n_50),
.B1(n_49),
.B2(n_48),
.Y(n_76)
);

NAND2xp33_ASAP7_75t_SL g86 ( 
.A(n_77),
.B(n_52),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_79),
.A2(n_81),
.B1(n_85),
.B2(n_75),
.Y(n_103)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_70),
.Y(n_80)
);

BUFx3_ASAP7_75t_L g98 ( 
.A(n_80),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_L g81 ( 
.A1(n_76),
.A2(n_62),
.B1(n_47),
.B2(n_43),
.Y(n_81)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_74),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_82),
.B(n_83),
.Y(n_95)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_71),
.Y(n_83)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_78),
.Y(n_84)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_84),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_73),
.A2(n_49),
.B1(n_54),
.B2(n_52),
.Y(n_85)
);

CKINVDCx16_ASAP7_75t_R g106 ( 
.A(n_86),
.Y(n_106)
);

INVxp67_ASAP7_75t_L g87 ( 
.A(n_77),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_87),
.B(n_89),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_77),
.A2(n_58),
.B1(n_2),
.B2(n_3),
.Y(n_88)
);

OAI21xp5_ASAP7_75t_L g96 ( 
.A1(n_88),
.A2(n_69),
.B(n_67),
.Y(n_96)
);

INVx11_ASAP7_75t_L g110 ( 
.A(n_90),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_91),
.B(n_38),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_68),
.B(n_1),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_92),
.B(n_68),
.Y(n_101)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_78),
.Y(n_93)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_93),
.Y(n_105)
);

BUFx12f_ASAP7_75t_L g94 ( 
.A(n_70),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_94),
.Y(n_100)
);

AND2x2_ASAP7_75t_L g123 ( 
.A(n_96),
.B(n_111),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_101),
.B(n_104),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_87),
.B(n_72),
.Y(n_102)
);

XNOR2xp5_ASAP7_75t_L g127 ( 
.A(n_102),
.B(n_108),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_103),
.A2(n_95),
.B1(n_107),
.B2(n_112),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_85),
.B(n_78),
.C(n_75),
.Y(n_107)
);

XNOR2xp5_ASAP7_75t_L g114 ( 
.A(n_107),
.B(n_90),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_86),
.B(n_70),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_80),
.B(n_1),
.Y(n_109)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_109),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_94),
.B(n_2),
.Y(n_111)
);

AOI21xp5_ASAP7_75t_L g112 ( 
.A1(n_79),
.A2(n_90),
.B(n_94),
.Y(n_112)
);

INVxp33_ASAP7_75t_L g126 ( 
.A(n_112),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_95),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_113),
.B(n_115),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_L g145 ( 
.A(n_114),
.B(n_30),
.Y(n_145)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_99),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_116),
.A2(n_125),
.B1(n_96),
.B2(n_98),
.Y(n_135)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_99),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_117),
.B(n_120),
.Y(n_139)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_100),
.Y(n_118)
);

INVx3_ASAP7_75t_L g131 ( 
.A(n_118),
.Y(n_131)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_105),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_105),
.Y(n_121)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_121),
.Y(n_134)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_102),
.Y(n_122)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_122),
.Y(n_136)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_98),
.Y(n_124)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_124),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_103),
.A2(n_58),
.B1(n_5),
.B2(n_6),
.Y(n_125)
);

AO22x1_ASAP7_75t_L g128 ( 
.A1(n_110),
.A2(n_37),
.B1(n_36),
.B2(n_35),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_L g143 ( 
.A1(n_128),
.A2(n_7),
.B(n_8),
.Y(n_143)
);

OAI32xp33_ASAP7_75t_L g130 ( 
.A1(n_97),
.A2(n_4),
.A3(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_L g133 ( 
.A1(n_130),
.A2(n_101),
.B(n_100),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_SL g132 ( 
.A(n_127),
.B(n_108),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_L g149 ( 
.A(n_132),
.B(n_145),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_133),
.B(n_141),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_135),
.B(n_137),
.Y(n_156)
);

OAI32xp33_ASAP7_75t_SL g137 ( 
.A1(n_114),
.A2(n_106),
.A3(n_110),
.B1(n_33),
.B2(n_32),
.Y(n_137)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_118),
.Y(n_141)
);

FAx1_ASAP7_75t_L g142 ( 
.A(n_126),
.B(n_106),
.CI(n_100),
.CON(n_142),
.SN(n_142)
);

AOI21xp5_ASAP7_75t_L g157 ( 
.A1(n_142),
.A2(n_22),
.B(n_15),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_143),
.B(n_144),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_119),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_SL g146 ( 
.A(n_129),
.B(n_8),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_SL g151 ( 
.A(n_146),
.B(n_147),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_123),
.B(n_29),
.C(n_23),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_142),
.A2(n_126),
.B1(n_123),
.B2(n_128),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_148),
.A2(n_150),
.B1(n_152),
.B2(n_155),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_142),
.A2(n_119),
.B1(n_10),
.B2(n_11),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_136),
.A2(n_9),
.B1(n_11),
.B2(n_12),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_138),
.A2(n_9),
.B1(n_12),
.B2(n_13),
.Y(n_155)
);

OAI21xp33_ASAP7_75t_L g160 ( 
.A1(n_157),
.A2(n_147),
.B(n_137),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_139),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_158),
.B(n_154),
.Y(n_165)
);

AOI21xp5_ASAP7_75t_L g159 ( 
.A1(n_153),
.A2(n_143),
.B(n_140),
.Y(n_159)
);

AOI31xp67_ASAP7_75t_L g168 ( 
.A1(n_159),
.A2(n_163),
.A3(n_155),
.B(n_152),
.Y(n_168)
);

AOI21xp5_ASAP7_75t_SL g167 ( 
.A1(n_160),
.A2(n_165),
.B(n_151),
.Y(n_167)
);

AOI322xp5_ASAP7_75t_L g162 ( 
.A1(n_156),
.A2(n_132),
.A3(n_145),
.B1(n_134),
.B2(n_131),
.C1(n_18),
.C2(n_14),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_162),
.B(n_164),
.Y(n_166)
);

AOI321xp33_ASAP7_75t_L g163 ( 
.A1(n_149),
.A2(n_14),
.A3(n_15),
.B1(n_16),
.B2(n_17),
.C(n_19),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_149),
.B(n_131),
.C(n_19),
.Y(n_164)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_167),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_168),
.B(n_169),
.Y(n_171)
);

XOR2xp5_ASAP7_75t_L g169 ( 
.A(n_160),
.B(n_148),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_170),
.B(n_166),
.C(n_150),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_172),
.B(n_171),
.Y(n_173)
);

AOI31xp33_ASAP7_75t_L g174 ( 
.A1(n_173),
.A2(n_161),
.A3(n_17),
.B(n_21),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_174),
.B(n_21),
.Y(n_175)
);

BUFx24_ASAP7_75t_SL g176 ( 
.A(n_175),
.Y(n_176)
);


endmodule