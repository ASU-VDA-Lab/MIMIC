module fake_jpeg_13851_n_361 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_361);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_361;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_256;
wire n_221;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

INVx3_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

INVx1_ASAP7_75t_SL g18 ( 
.A(n_11),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_6),
.Y(n_19)
);

BUFx12_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

INVx13_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_6),
.Y(n_24)
);

INVx6_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_0),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

CKINVDCx16_ASAP7_75t_R g32 ( 
.A(n_14),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_10),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_6),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_16),
.Y(n_35)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_35),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_20),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_36),
.B(n_27),
.Y(n_58)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_22),
.Y(n_37)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_37),
.Y(n_57)
);

INVx11_ASAP7_75t_L g38 ( 
.A(n_23),
.Y(n_38)
);

INVx11_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

INVx2_ASAP7_75t_SL g39 ( 
.A(n_16),
.Y(n_39)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_39),
.Y(n_62)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_21),
.Y(n_40)
);

INVx5_ASAP7_75t_L g77 ( 
.A(n_40),
.Y(n_77)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_21),
.Y(n_41)
);

INVx1_ASAP7_75t_SL g79 ( 
.A(n_41),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_21),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_42),
.Y(n_60)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_16),
.Y(n_43)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_43),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_21),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_44),
.Y(n_80)
);

INVx11_ASAP7_75t_L g45 ( 
.A(n_23),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g72 ( 
.A(n_45),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_30),
.Y(n_46)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_46),
.Y(n_70)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_22),
.Y(n_47)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_47),
.Y(n_61)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_30),
.Y(n_48)
);

INVx6_ASAP7_75t_L g76 ( 
.A(n_48),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_28),
.B(n_0),
.Y(n_49)
);

MAJIxp5_ASAP7_75t_L g78 ( 
.A(n_49),
.B(n_52),
.C(n_32),
.Y(n_78)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_16),
.Y(n_50)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_50),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_30),
.Y(n_51)
);

INVx8_ASAP7_75t_L g66 ( 
.A(n_51),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_28),
.B(n_0),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_39),
.A2(n_18),
.B1(n_28),
.B2(n_17),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_53),
.A2(n_75),
.B1(n_81),
.B2(n_38),
.Y(n_82)
);

OAI21xp33_ASAP7_75t_SL g55 ( 
.A1(n_49),
.A2(n_18),
.B(n_52),
.Y(n_55)
);

OR2x4_ASAP7_75t_L g113 ( 
.A(n_55),
.B(n_45),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_L g56 ( 
.A1(n_48),
.A2(n_18),
.B1(n_25),
.B2(n_24),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_56),
.A2(n_65),
.B1(n_68),
.B2(n_31),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_58),
.B(n_67),
.Y(n_87)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_37),
.Y(n_64)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_64),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_L g65 ( 
.A1(n_48),
.A2(n_25),
.B1(n_19),
.B2(n_24),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_36),
.B(n_33),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g68 ( 
.A1(n_52),
.A2(n_25),
.B1(n_34),
.B2(n_33),
.Y(n_68)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_47),
.Y(n_69)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_69),
.Y(n_97)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_35),
.Y(n_71)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_71),
.Y(n_104)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_38),
.Y(n_74)
);

BUFx2_ASAP7_75t_L g101 ( 
.A(n_74),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_39),
.A2(n_17),
.B1(n_22),
.B2(n_29),
.Y(n_75)
);

AND2x2_ASAP7_75t_L g103 ( 
.A(n_78),
.B(n_27),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_39),
.A2(n_17),
.B1(n_29),
.B2(n_16),
.Y(n_81)
);

INVxp67_ASAP7_75t_L g142 ( 
.A(n_82),
.Y(n_142)
);

INVx6_ASAP7_75t_L g83 ( 
.A(n_60),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g146 ( 
.A(n_83),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_L g84 ( 
.A1(n_57),
.A2(n_40),
.B1(n_29),
.B2(n_26),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_84),
.A2(n_31),
.B1(n_79),
.B2(n_70),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_78),
.B(n_49),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_85),
.B(n_86),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_57),
.B(n_35),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_54),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_88),
.B(n_89),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_54),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_61),
.B(n_24),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_SL g125 ( 
.A(n_90),
.B(n_98),
.Y(n_125)
);

INVxp67_ASAP7_75t_L g91 ( 
.A(n_62),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_91),
.B(n_102),
.Y(n_139)
);

INVx1_ASAP7_75t_SL g92 ( 
.A(n_62),
.Y(n_92)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_92),
.Y(n_121)
);

CKINVDCx14_ASAP7_75t_R g93 ( 
.A(n_72),
.Y(n_93)
);

INVx11_ASAP7_75t_L g128 ( 
.A(n_93),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_61),
.B(n_26),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_94),
.B(n_99),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_64),
.A2(n_31),
.B1(n_19),
.B2(n_16),
.Y(n_95)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_95),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_SL g98 ( 
.A(n_69),
.B(n_19),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_59),
.B(n_43),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_59),
.B(n_71),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_100),
.B(n_105),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_63),
.Y(n_102)
);

XNOR2xp5_ASAP7_75t_L g123 ( 
.A(n_103),
.B(n_108),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_72),
.B(n_32),
.Y(n_105)
);

INVxp67_ASAP7_75t_L g106 ( 
.A(n_66),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_106),
.B(n_110),
.Y(n_140)
);

OR2x2_ASAP7_75t_SL g107 ( 
.A(n_63),
.B(n_45),
.Y(n_107)
);

AOI21xp33_ASAP7_75t_L g117 ( 
.A1(n_107),
.A2(n_113),
.B(n_23),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_76),
.B(n_43),
.Y(n_108)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_74),
.Y(n_109)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_109),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_77),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_76),
.B(n_27),
.Y(n_111)
);

XNOR2xp5_ASAP7_75t_L g144 ( 
.A(n_111),
.B(n_116),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_112),
.A2(n_44),
.B1(n_42),
.B2(n_51),
.Y(n_136)
);

INVx11_ASAP7_75t_L g114 ( 
.A(n_72),
.Y(n_114)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_114),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_77),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_115),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_66),
.B(n_27),
.Y(n_116)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_117),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_119),
.A2(n_135),
.B1(n_137),
.B2(n_92),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_L g122 ( 
.A1(n_90),
.A2(n_40),
.B1(n_70),
.B2(n_80),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_122),
.A2(n_136),
.B1(n_141),
.B2(n_60),
.Y(n_166)
);

INVx4_ASAP7_75t_L g129 ( 
.A(n_114),
.Y(n_129)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_129),
.Y(n_148)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_104),
.Y(n_130)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_130),
.Y(n_158)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_86),
.Y(n_131)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_131),
.Y(n_167)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_97),
.Y(n_132)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_132),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_85),
.A2(n_25),
.B1(n_34),
.B2(n_80),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_113),
.A2(n_44),
.B1(n_42),
.B2(n_46),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_94),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_138),
.B(n_27),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_112),
.A2(n_44),
.B1(n_51),
.B2(n_42),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_103),
.B(n_73),
.C(n_79),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_143),
.B(n_50),
.C(n_72),
.Y(n_171)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_104),
.Y(n_147)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_147),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_127),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_149),
.B(n_168),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_L g150 ( 
.A1(n_145),
.A2(n_98),
.B(n_87),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_L g185 ( 
.A1(n_150),
.A2(n_118),
.B(n_121),
.Y(n_185)
);

OAI22xp33_ASAP7_75t_SL g194 ( 
.A1(n_151),
.A2(n_162),
.B1(n_156),
.B2(n_141),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_131),
.A2(n_103),
.B1(n_116),
.B2(n_111),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_152),
.A2(n_153),
.B1(n_156),
.B2(n_161),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_138),
.A2(n_108),
.B1(n_100),
.B2(n_92),
.Y(n_153)
);

INVxp67_ASAP7_75t_L g154 ( 
.A(n_128),
.Y(n_154)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_154),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_125),
.B(n_120),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_SL g183 ( 
.A(n_155),
.B(n_163),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_137),
.A2(n_97),
.B1(n_99),
.B2(n_115),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_120),
.A2(n_87),
.B1(n_105),
.B2(n_46),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_157),
.A2(n_160),
.B1(n_166),
.B2(n_129),
.Y(n_200)
);

AOI22xp33_ASAP7_75t_SL g159 ( 
.A1(n_142),
.A2(n_101),
.B1(n_110),
.B2(n_114),
.Y(n_159)
);

AOI22xp33_ASAP7_75t_SL g214 ( 
.A1(n_159),
.A2(n_165),
.B1(n_41),
.B2(n_2),
.Y(n_214)
);

OAI22xp33_ASAP7_75t_SL g160 ( 
.A1(n_142),
.A2(n_107),
.B1(n_96),
.B2(n_101),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_133),
.A2(n_96),
.B1(n_88),
.B2(n_89),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_133),
.A2(n_83),
.B1(n_102),
.B2(n_46),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_162),
.A2(n_169),
.B1(n_170),
.B2(n_41),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_125),
.B(n_109),
.Y(n_163)
);

INVxp67_ASAP7_75t_L g164 ( 
.A(n_128),
.Y(n_164)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_164),
.Y(n_193)
);

INVx3_ASAP7_75t_SL g165 ( 
.A(n_146),
.Y(n_165)
);

CKINVDCx14_ASAP7_75t_R g168 ( 
.A(n_140),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_145),
.A2(n_83),
.B1(n_51),
.B2(n_101),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_143),
.A2(n_93),
.B1(n_34),
.B2(n_73),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_171),
.B(n_178),
.C(n_124),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_134),
.B(n_12),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_SL g206 ( 
.A(n_172),
.B(n_176),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_175),
.B(n_182),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_139),
.B(n_27),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_123),
.B(n_50),
.C(n_34),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_132),
.Y(n_179)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_179),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_SL g180 ( 
.A(n_123),
.B(n_10),
.Y(n_180)
);

OR2x2_ASAP7_75t_L g201 ( 
.A(n_180),
.B(n_124),
.Y(n_201)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_147),
.Y(n_181)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_181),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_144),
.B(n_9),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_185),
.B(n_195),
.Y(n_227)
);

CKINVDCx14_ASAP7_75t_R g186 ( 
.A(n_149),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_186),
.B(n_201),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_L g188 ( 
.A(n_167),
.B(n_144),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_188),
.B(n_190),
.C(n_196),
.Y(n_224)
);

OAI21xp5_ASAP7_75t_SL g189 ( 
.A1(n_173),
.A2(n_118),
.B(n_121),
.Y(n_189)
);

OR2x2_ASAP7_75t_L g219 ( 
.A(n_189),
.B(n_169),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g190 ( 
.A(n_152),
.B(n_126),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_167),
.B(n_130),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_192),
.B(n_194),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_161),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g198 ( 
.A(n_173),
.B(n_126),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_198),
.B(n_202),
.C(n_215),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_L g218 ( 
.A1(n_200),
.A2(n_207),
.B1(n_209),
.B2(n_214),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_178),
.B(n_136),
.C(n_146),
.Y(n_202)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_203),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_151),
.A2(n_41),
.B1(n_30),
.B2(n_23),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_204),
.B(n_205),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_157),
.B(n_0),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_150),
.A2(n_41),
.B1(n_20),
.B2(n_9),
.Y(n_207)
);

NOR2xp67_ASAP7_75t_L g208 ( 
.A(n_180),
.B(n_9),
.Y(n_208)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_208),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_153),
.A2(n_41),
.B1(n_20),
.B2(n_8),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_174),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_210),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_174),
.B(n_8),
.Y(n_211)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_211),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_179),
.B(n_8),
.Y(n_212)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_212),
.Y(n_238)
);

XOR2xp5_ASAP7_75t_L g215 ( 
.A(n_171),
.B(n_20),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_177),
.Y(n_216)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_216),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_170),
.B(n_181),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_217),
.B(n_20),
.C(n_2),
.Y(n_235)
);

INVx1_ASAP7_75t_SL g254 ( 
.A(n_219),
.Y(n_254)
);

OA21x2_ASAP7_75t_L g220 ( 
.A1(n_200),
.A2(n_164),
.B(n_154),
.Y(n_220)
);

INVxp67_ASAP7_75t_L g264 ( 
.A(n_220),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_L g222 ( 
.A1(n_199),
.A2(n_165),
.B1(n_177),
.B2(n_158),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_L g251 ( 
.A1(n_222),
.A2(n_207),
.B1(n_216),
.B2(n_193),
.Y(n_251)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_192),
.Y(n_223)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_223),
.Y(n_252)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_197),
.Y(n_225)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_225),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_202),
.A2(n_165),
.B1(n_158),
.B2(n_148),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_229),
.A2(n_236),
.B1(n_239),
.B2(n_241),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_191),
.B(n_148),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_230),
.B(n_245),
.Y(n_249)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_197),
.Y(n_231)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_231),
.Y(n_265)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_213),
.Y(n_232)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_232),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_235),
.B(n_240),
.C(n_15),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_205),
.A2(n_7),
.B1(n_14),
.B2(n_13),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_185),
.A2(n_191),
.B1(n_196),
.B2(n_209),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_198),
.B(n_15),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_183),
.A2(n_190),
.B1(n_217),
.B2(n_201),
.Y(n_241)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_213),
.Y(n_244)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_244),
.Y(n_269)
);

BUFx2_ASAP7_75t_L g245 ( 
.A(n_187),
.Y(n_245)
);

AND2x2_ASAP7_75t_SL g246 ( 
.A(n_189),
.B(n_1),
.Y(n_246)
);

CKINVDCx14_ASAP7_75t_R g267 ( 
.A(n_246),
.Y(n_267)
);

XOR2xp5_ASAP7_75t_L g248 ( 
.A(n_224),
.B(n_215),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_248),
.B(n_250),
.C(n_257),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_233),
.B(n_188),
.Y(n_250)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_251),
.Y(n_276)
);

AOI21xp5_ASAP7_75t_L g253 ( 
.A1(n_227),
.A2(n_219),
.B(n_242),
.Y(n_253)
);

AOI21xp5_ASAP7_75t_L g281 ( 
.A1(n_253),
.A2(n_259),
.B(n_234),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_239),
.A2(n_203),
.B1(n_204),
.B2(n_206),
.Y(n_256)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_256),
.Y(n_284)
);

XOR2xp5_ASAP7_75t_L g257 ( 
.A(n_224),
.B(n_184),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_258),
.B(n_271),
.Y(n_279)
);

AOI21xp5_ASAP7_75t_L g259 ( 
.A1(n_233),
.A2(n_15),
.B(n_13),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_241),
.B(n_7),
.C(n_11),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_260),
.B(n_266),
.C(n_270),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_221),
.A2(n_7),
.B1(n_2),
.B2(n_3),
.Y(n_262)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_262),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_229),
.B(n_1),
.C(n_3),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_247),
.B(n_1),
.Y(n_268)
);

CKINVDCx14_ASAP7_75t_R g280 ( 
.A(n_268),
.Y(n_280)
);

XOR2xp5_ASAP7_75t_L g270 ( 
.A(n_240),
.B(n_230),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_246),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_225),
.Y(n_272)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_272),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_223),
.B(n_3),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_273),
.B(n_235),
.C(n_246),
.Y(n_289)
);

INVxp67_ASAP7_75t_L g275 ( 
.A(n_253),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_275),
.B(n_277),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_249),
.Y(n_277)
);

AOI22xp33_ASAP7_75t_L g278 ( 
.A1(n_254),
.A2(n_221),
.B1(n_237),
.B2(n_238),
.Y(n_278)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_278),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_SL g296 ( 
.A(n_281),
.B(n_289),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_252),
.B(n_232),
.Y(n_282)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_282),
.Y(n_308)
);

INVx1_ASAP7_75t_SL g283 ( 
.A(n_254),
.Y(n_283)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_283),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_273),
.B(n_245),
.Y(n_286)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_286),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_263),
.B(n_226),
.Y(n_287)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_287),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_269),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_SL g305 ( 
.A(n_290),
.B(n_295),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_250),
.B(n_248),
.C(n_257),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_291),
.B(n_255),
.C(n_260),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_265),
.B(n_226),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g303 ( 
.A(n_293),
.Y(n_303)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_261),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_294),
.B(n_231),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_270),
.B(n_236),
.Y(n_295)
);

XOR2xp5_ASAP7_75t_L g297 ( 
.A(n_274),
.B(n_255),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_L g320 ( 
.A(n_297),
.B(n_300),
.Y(n_320)
);

XOR2xp5_ASAP7_75t_L g301 ( 
.A(n_274),
.B(n_256),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_301),
.B(n_302),
.C(n_276),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_291),
.B(n_264),
.C(n_220),
.Y(n_302)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_304),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_L g306 ( 
.A1(n_284),
.A2(n_264),
.B1(n_220),
.B2(n_218),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_L g324 ( 
.A1(n_306),
.A2(n_267),
.B1(n_228),
.B2(n_266),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_SL g309 ( 
.A(n_275),
.B(n_258),
.Y(n_309)
);

CKINVDCx14_ASAP7_75t_R g325 ( 
.A(n_309),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_282),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_310),
.B(n_285),
.Y(n_323)
);

OAI22xp5_ASAP7_75t_SL g314 ( 
.A1(n_298),
.A2(n_306),
.B1(n_284),
.B2(n_283),
.Y(n_314)
);

AOI22xp33_ASAP7_75t_L g335 ( 
.A1(n_314),
.A2(n_322),
.B1(n_323),
.B2(n_312),
.Y(n_335)
);

AOI22xp5_ASAP7_75t_L g315 ( 
.A1(n_298),
.A2(n_276),
.B1(n_277),
.B2(n_293),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_SL g334 ( 
.A1(n_315),
.A2(n_308),
.B1(n_312),
.B2(n_307),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_316),
.B(n_318),
.C(n_319),
.Y(n_327)
);

OAI21xp5_ASAP7_75t_SL g317 ( 
.A1(n_296),
.A2(n_281),
.B(n_279),
.Y(n_317)
);

XNOR2xp5_ASAP7_75t_L g328 ( 
.A(n_317),
.B(n_326),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_301),
.B(n_288),
.C(n_286),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_297),
.B(n_288),
.C(n_287),
.Y(n_319)
);

HB1xp67_ASAP7_75t_L g321 ( 
.A(n_305),
.Y(n_321)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_321),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_SL g322 ( 
.A1(n_303),
.A2(n_285),
.B1(n_262),
.B2(n_228),
.Y(n_322)
);

AOI22xp5_ASAP7_75t_SL g338 ( 
.A1(n_324),
.A2(n_292),
.B1(n_294),
.B2(n_243),
.Y(n_338)
);

OAI21xp5_ASAP7_75t_SL g326 ( 
.A1(n_299),
.A2(n_280),
.B(n_292),
.Y(n_326)
);

XOR2xp5_ASAP7_75t_L g329 ( 
.A(n_316),
.B(n_302),
.Y(n_329)
);

AND2x2_ASAP7_75t_L g343 ( 
.A(n_329),
.B(n_337),
.Y(n_343)
);

AND2x2_ASAP7_75t_L g331 ( 
.A(n_319),
.B(n_299),
.Y(n_331)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_331),
.Y(n_339)
);

AND2x2_ASAP7_75t_L g332 ( 
.A(n_318),
.B(n_300),
.Y(n_332)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_332),
.Y(n_346)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_320),
.B(n_307),
.C(n_311),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_333),
.B(n_334),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_335),
.B(n_314),
.Y(n_341)
);

NOR2xp67_ASAP7_75t_L g336 ( 
.A(n_313),
.B(n_289),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_336),
.B(n_4),
.Y(n_345)
);

XOR2xp5_ASAP7_75t_L g337 ( 
.A(n_320),
.B(n_311),
.Y(n_337)
);

OAI22xp5_ASAP7_75t_L g344 ( 
.A1(n_338),
.A2(n_326),
.B1(n_322),
.B2(n_5),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_341),
.B(n_342),
.Y(n_350)
);

MAJIxp5_ASAP7_75t_L g342 ( 
.A(n_327),
.B(n_325),
.C(n_315),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_344),
.B(n_347),
.Y(n_353)
);

OAI21xp5_ASAP7_75t_SL g348 ( 
.A1(n_345),
.A2(n_4),
.B(n_5),
.Y(n_348)
);

OAI22xp33_ASAP7_75t_SL g347 ( 
.A1(n_330),
.A2(n_335),
.B1(n_328),
.B2(n_331),
.Y(n_347)
);

OR2x2_ASAP7_75t_L g356 ( 
.A(n_348),
.B(n_352),
.Y(n_356)
);

NOR2xp33_ASAP7_75t_L g349 ( 
.A(n_346),
.B(n_337),
.Y(n_349)
);

AOI21xp5_ASAP7_75t_L g354 ( 
.A1(n_349),
.A2(n_351),
.B(n_343),
.Y(n_354)
);

AND2x2_ASAP7_75t_L g351 ( 
.A(n_343),
.B(n_332),
.Y(n_351)
);

MAJIxp5_ASAP7_75t_L g352 ( 
.A(n_339),
.B(n_329),
.C(n_5),
.Y(n_352)
);

OAI21xp5_ASAP7_75t_SL g357 ( 
.A1(n_354),
.A2(n_355),
.B(n_340),
.Y(n_357)
);

BUFx24_ASAP7_75t_SL g355 ( 
.A(n_350),
.Y(n_355)
);

INVxp67_ASAP7_75t_L g358 ( 
.A(n_357),
.Y(n_358)
);

AOI21xp5_ASAP7_75t_L g359 ( 
.A1(n_358),
.A2(n_353),
.B(n_345),
.Y(n_359)
);

XNOR2xp5_ASAP7_75t_L g360 ( 
.A(n_359),
.B(n_349),
.Y(n_360)
);

XOR2xp5_ASAP7_75t_L g361 ( 
.A(n_360),
.B(n_356),
.Y(n_361)
);


endmodule