module fake_jpeg_6763_n_56 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_7, n_56);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;
input n_7;

output n_56;

wire n_13;
wire n_21;
wire n_53;
wire n_33;
wire n_54;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_55;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_31;
wire n_25;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_8;
wire n_15;

INVx2_ASAP7_75t_L g8 ( 
.A(n_0),
.Y(n_8)
);

INVx8_ASAP7_75t_L g9 ( 
.A(n_1),
.Y(n_9)
);

BUFx12f_ASAP7_75t_L g10 ( 
.A(n_3),
.Y(n_10)
);

INVx3_ASAP7_75t_L g11 ( 
.A(n_7),
.Y(n_11)
);

BUFx6f_ASAP7_75t_L g12 ( 
.A(n_7),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_6),
.Y(n_13)
);

NOR2xp67_ASAP7_75t_L g14 ( 
.A(n_2),
.B(n_1),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_2),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_3),
.B(n_0),
.Y(n_16)
);

OR2x2_ASAP7_75t_L g17 ( 
.A(n_14),
.B(n_0),
.Y(n_17)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_17),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_13),
.B(n_15),
.Y(n_18)
);

MAJIxp5_ASAP7_75t_L g23 ( 
.A(n_18),
.B(n_20),
.C(n_16),
.Y(n_23)
);

INVx3_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_19),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_13),
.B(n_1),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_SL g21 ( 
.A(n_15),
.B(n_6),
.Y(n_21)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_21),
.Y(n_29)
);

INVx6_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_22),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_23),
.B(n_27),
.Y(n_30)
);

AOI22xp33_ASAP7_75t_SL g26 ( 
.A1(n_19),
.A2(n_11),
.B1(n_8),
.B2(n_9),
.Y(n_26)
);

AOI22xp33_ASAP7_75t_SL g37 ( 
.A1(n_26),
.A2(n_11),
.B1(n_9),
.B2(n_19),
.Y(n_37)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_22),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_24),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_31),
.B(n_34),
.Y(n_39)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_24),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_32),
.B(n_35),
.Y(n_42)
);

OAI21xp5_ASAP7_75t_L g33 ( 
.A1(n_28),
.A2(n_20),
.B(n_18),
.Y(n_33)
);

MAJIxp5_ASAP7_75t_L g41 ( 
.A(n_33),
.B(n_23),
.C(n_29),
.Y(n_41)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_27),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_27),
.B(n_21),
.Y(n_35)
);

CKINVDCx16_ASAP7_75t_R g36 ( 
.A(n_25),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_SL g40 ( 
.A(n_36),
.B(n_4),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_SL g38 ( 
.A1(n_37),
.A2(n_8),
.B1(n_28),
.B2(n_22),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_L g45 ( 
.A1(n_38),
.A2(n_41),
.B1(n_29),
.B2(n_17),
.Y(n_45)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_40),
.Y(n_44)
);

NAND3xp33_ASAP7_75t_SL g43 ( 
.A(n_41),
.B(n_30),
.C(n_33),
.Y(n_43)
);

MAJIxp5_ASAP7_75t_L g47 ( 
.A(n_43),
.B(n_45),
.C(n_46),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_42),
.B(n_34),
.Y(n_46)
);

MAJIxp5_ASAP7_75t_L g48 ( 
.A(n_46),
.B(n_39),
.C(n_32),
.Y(n_48)
);

MAJIxp5_ASAP7_75t_L g51 ( 
.A(n_48),
.B(n_49),
.C(n_10),
.Y(n_51)
);

MAJIxp5_ASAP7_75t_L g49 ( 
.A(n_44),
.B(n_25),
.C(n_31),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_L g50 ( 
.A1(n_47),
.A2(n_44),
.B1(n_25),
.B2(n_12),
.Y(n_50)
);

INVxp67_ASAP7_75t_L g52 ( 
.A(n_50),
.Y(n_52)
);

MAJIxp5_ASAP7_75t_L g53 ( 
.A(n_51),
.B(n_10),
.C(n_17),
.Y(n_53)
);

MAJIxp5_ASAP7_75t_L g54 ( 
.A(n_53),
.B(n_4),
.C(n_5),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_54),
.B(n_5),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_55),
.B(n_52),
.Y(n_56)
);


endmodule