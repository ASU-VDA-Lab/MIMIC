module fake_jpeg_21779_n_72 (n_3, n_2, n_1, n_0, n_4, n_8, n_6, n_5, n_7, n_72);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_6;
input n_5;
input n_7;

output n_72;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_23;
wire n_10;
wire n_69;
wire n_27;
wire n_55;
wire n_64;
wire n_47;
wire n_22;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_20;
wire n_18;
wire n_59;
wire n_35;
wire n_48;
wire n_68;
wire n_52;
wire n_71;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_65;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_16;
wire n_24;
wire n_44;
wire n_38;
wire n_26;
wire n_28;
wire n_9;
wire n_36;
wire n_11;
wire n_62;
wire n_25;
wire n_17;
wire n_31;
wire n_56;
wire n_67;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_70;
wire n_15;
wire n_66;

CKINVDCx20_ASAP7_75t_R g9 ( 
.A(n_8),
.Y(n_9)
);

CKINVDCx20_ASAP7_75t_R g10 ( 
.A(n_1),
.Y(n_10)
);

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_5),
.Y(n_11)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_3),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_0),
.B(n_3),
.Y(n_13)
);

INVx6_ASAP7_75t_L g14 ( 
.A(n_8),
.Y(n_14)
);

INVx4_ASAP7_75t_L g15 ( 
.A(n_7),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_2),
.B(n_1),
.Y(n_16)
);

CKINVDCx16_ASAP7_75t_R g17 ( 
.A(n_4),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_7),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_13),
.B(n_0),
.Y(n_20)
);

NAND2xp33_ASAP7_75t_SL g34 ( 
.A(n_20),
.B(n_25),
.Y(n_34)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_19),
.Y(n_21)
);

INVx5_ASAP7_75t_L g39 ( 
.A(n_21),
.Y(n_39)
);

INVx4_ASAP7_75t_L g22 ( 
.A(n_19),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_22),
.B(n_23),
.Y(n_28)
);

BUFx16f_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_19),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_24),
.B(n_14),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_13),
.B(n_0),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_9),
.B(n_1),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_SL g35 ( 
.A(n_26),
.B(n_27),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_9),
.B(n_2),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_L g29 ( 
.A1(n_20),
.A2(n_14),
.B1(n_15),
.B2(n_10),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_SL g49 ( 
.A1(n_29),
.A2(n_12),
.B1(n_11),
.B2(n_17),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_21),
.Y(n_30)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_30),
.Y(n_43)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_31),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_25),
.B(n_18),
.Y(n_32)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_32),
.Y(n_41)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_23),
.Y(n_33)
);

INVxp67_ASAP7_75t_L g47 ( 
.A(n_33),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_23),
.B(n_14),
.Y(n_36)
);

AND2x2_ASAP7_75t_L g42 ( 
.A(n_36),
.B(n_10),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_24),
.Y(n_37)
);

INVxp67_ASAP7_75t_L g48 ( 
.A(n_37),
.Y(n_48)
);

INVxp67_ASAP7_75t_L g38 ( 
.A(n_22),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_38),
.B(n_17),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_42),
.B(n_44),
.Y(n_50)
);

OR2x2_ASAP7_75t_L g44 ( 
.A(n_34),
.B(n_11),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_45),
.B(n_33),
.Y(n_55)
);

AND2x2_ASAP7_75t_L g46 ( 
.A(n_36),
.B(n_18),
.Y(n_46)
);

HAxp5_ASAP7_75t_SL g51 ( 
.A(n_46),
.B(n_12),
.CON(n_51),
.SN(n_51)
);

XNOR2xp5_ASAP7_75t_L g52 ( 
.A(n_49),
.B(n_35),
.Y(n_52)
);

AND2x2_ASAP7_75t_L g60 ( 
.A(n_51),
.B(n_52),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_42),
.B(n_30),
.Y(n_53)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_53),
.Y(n_59)
);

MAJIxp5_ASAP7_75t_L g54 ( 
.A(n_40),
.B(n_28),
.C(n_37),
.Y(n_54)
);

MAJIxp5_ASAP7_75t_L g57 ( 
.A(n_54),
.B(n_56),
.C(n_37),
.Y(n_57)
);

INVx13_ASAP7_75t_L g61 ( 
.A(n_55),
.Y(n_61)
);

MAJIxp5_ASAP7_75t_L g56 ( 
.A(n_44),
.B(n_37),
.C(n_39),
.Y(n_56)
);

MAJIxp5_ASAP7_75t_L g64 ( 
.A(n_57),
.B(n_58),
.C(n_41),
.Y(n_64)
);

OAI21xp5_ASAP7_75t_L g58 ( 
.A1(n_56),
.A2(n_46),
.B(n_48),
.Y(n_58)
);

AO221x1_ASAP7_75t_L g62 ( 
.A1(n_61),
.A2(n_43),
.B1(n_39),
.B2(n_48),
.C(n_47),
.Y(n_62)
);

INVxp67_ASAP7_75t_L g66 ( 
.A(n_62),
.Y(n_66)
);

AOI21xp33_ASAP7_75t_L g63 ( 
.A1(n_59),
.A2(n_50),
.B(n_51),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_63),
.B(n_64),
.Y(n_67)
);

MAJIxp5_ASAP7_75t_L g65 ( 
.A(n_57),
.B(n_47),
.C(n_16),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_66),
.B(n_61),
.Y(n_68)
);

OAI21xp5_ASAP7_75t_L g70 ( 
.A1(n_68),
.A2(n_69),
.B(n_60),
.Y(n_70)
);

OAI21xp5_ASAP7_75t_SL g69 ( 
.A1(n_67),
.A2(n_65),
.B(n_58),
.Y(n_69)
);

OAI32xp33_ASAP7_75t_SL g71 ( 
.A1(n_70),
.A2(n_60),
.A3(n_6),
.B1(n_5),
.B2(n_38),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g72 ( 
.A1(n_71),
.A2(n_60),
.B1(n_6),
.B2(n_43),
.Y(n_72)
);


endmodule