module fake_jpeg_155_n_443 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_443);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_443;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_433;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_11),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_7),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_4),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_14),
.B(n_4),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_0),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_8),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_11),
.Y(n_35)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_1),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_14),
.Y(n_37)
);

BUFx5_ASAP7_75t_L g38 ( 
.A(n_0),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_1),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_9),
.Y(n_40)
);

INVx5_ASAP7_75t_L g41 ( 
.A(n_1),
.Y(n_41)
);

BUFx12_ASAP7_75t_L g42 ( 
.A(n_8),
.Y(n_42)
);

CKINVDCx16_ASAP7_75t_R g43 ( 
.A(n_13),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_6),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_2),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_13),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_17),
.Y(n_47)
);

INVx11_ASAP7_75t_L g48 ( 
.A(n_2),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_3),
.Y(n_49)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_2),
.Y(n_50)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_2),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_5),
.Y(n_52)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_15),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_24),
.Y(n_54)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_54),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_27),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_55),
.B(n_57),
.Y(n_116)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_41),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g172 ( 
.A(n_56),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_53),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_53),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_58),
.B(n_59),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_23),
.Y(n_59)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_39),
.Y(n_60)
);

INVx4_ASAP7_75t_SL g122 ( 
.A(n_60),
.Y(n_122)
);

INVx4_ASAP7_75t_SL g61 ( 
.A(n_39),
.Y(n_61)
);

INVx1_ASAP7_75t_SL g129 ( 
.A(n_61),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_23),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_62),
.B(n_71),
.Y(n_139)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_23),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g178 ( 
.A(n_63),
.Y(n_178)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_32),
.Y(n_64)
);

INVx6_ASAP7_75t_L g151 ( 
.A(n_64),
.Y(n_151)
);

INVx8_ASAP7_75t_L g65 ( 
.A(n_39),
.Y(n_65)
);

INVx5_ASAP7_75t_L g120 ( 
.A(n_65),
.Y(n_120)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_39),
.Y(n_66)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_66),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_20),
.B(n_9),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_67),
.B(n_73),
.Y(n_125)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_41),
.Y(n_68)
);

BUFx2_ASAP7_75t_L g130 ( 
.A(n_68),
.Y(n_130)
);

INVx8_ASAP7_75t_L g69 ( 
.A(n_19),
.Y(n_69)
);

INVx5_ASAP7_75t_L g135 ( 
.A(n_69),
.Y(n_135)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_19),
.Y(n_70)
);

INVx5_ASAP7_75t_L g160 ( 
.A(n_70),
.Y(n_160)
);

CKINVDCx14_ASAP7_75t_R g71 ( 
.A(n_43),
.Y(n_71)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_34),
.Y(n_72)
);

BUFx2_ASAP7_75t_L g186 ( 
.A(n_72),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_18),
.B(n_10),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_32),
.Y(n_74)
);

INVx6_ASAP7_75t_L g175 ( 
.A(n_74),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_24),
.A2(n_10),
.B1(n_3),
.B2(n_5),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_75),
.A2(n_52),
.B1(n_25),
.B2(n_22),
.Y(n_123)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_33),
.Y(n_76)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_76),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_32),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_77),
.B(n_78),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_35),
.Y(n_78)
);

BUFx12_ASAP7_75t_L g79 ( 
.A(n_42),
.Y(n_79)
);

BUFx12f_ASAP7_75t_L g156 ( 
.A(n_79),
.Y(n_156)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_33),
.Y(n_80)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_80),
.Y(n_136)
);

CKINVDCx16_ASAP7_75t_R g81 ( 
.A(n_35),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_81),
.B(n_99),
.Y(n_148)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_44),
.Y(n_82)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_82),
.Y(n_137)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_34),
.Y(n_83)
);

INVx4_ASAP7_75t_L g121 ( 
.A(n_83),
.Y(n_121)
);

BUFx12f_ASAP7_75t_L g84 ( 
.A(n_42),
.Y(n_84)
);

INVx5_ASAP7_75t_L g187 ( 
.A(n_84),
.Y(n_187)
);

INVx5_ASAP7_75t_L g85 ( 
.A(n_19),
.Y(n_85)
);

INVx4_ASAP7_75t_L g124 ( 
.A(n_85),
.Y(n_124)
);

BUFx12f_ASAP7_75t_L g86 ( 
.A(n_42),
.Y(n_86)
);

INVx5_ASAP7_75t_L g177 ( 
.A(n_86),
.Y(n_177)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_35),
.Y(n_87)
);

INVx3_ASAP7_75t_SL g145 ( 
.A(n_87),
.Y(n_145)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_26),
.Y(n_88)
);

INVx4_ASAP7_75t_L g140 ( 
.A(n_88),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_20),
.B(n_10),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_89),
.B(n_107),
.Y(n_131)
);

INVx11_ASAP7_75t_L g90 ( 
.A(n_19),
.Y(n_90)
);

INVx11_ASAP7_75t_L g185 ( 
.A(n_90),
.Y(n_185)
);

BUFx5_ASAP7_75t_L g91 ( 
.A(n_26),
.Y(n_91)
);

INVx4_ASAP7_75t_L g154 ( 
.A(n_91),
.Y(n_154)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_44),
.Y(n_92)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_92),
.Y(n_138)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_18),
.Y(n_93)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_93),
.Y(n_181)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_50),
.Y(n_94)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_94),
.Y(n_155)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_50),
.Y(n_95)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_95),
.Y(n_158)
);

BUFx12f_ASAP7_75t_L g96 ( 
.A(n_42),
.Y(n_96)
);

INVx4_ASAP7_75t_L g180 ( 
.A(n_96),
.Y(n_180)
);

INVx5_ASAP7_75t_L g97 ( 
.A(n_36),
.Y(n_97)
);

HB1xp67_ASAP7_75t_L g117 ( 
.A(n_97),
.Y(n_117)
);

NAND2x1_ASAP7_75t_SL g98 ( 
.A(n_21),
.B(n_1),
.Y(n_98)
);

AND2x2_ASAP7_75t_L g162 ( 
.A(n_98),
.B(n_101),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_36),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_51),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_100),
.B(n_106),
.Y(n_153)
);

INVx1_ASAP7_75t_SL g101 ( 
.A(n_28),
.Y(n_101)
);

CKINVDCx6p67_ASAP7_75t_R g102 ( 
.A(n_38),
.Y(n_102)
);

BUFx12f_ASAP7_75t_L g165 ( 
.A(n_102),
.Y(n_165)
);

AOI21xp33_ASAP7_75t_L g103 ( 
.A1(n_21),
.A2(n_5),
.B(n_6),
.Y(n_103)
);

AOI21xp33_ASAP7_75t_L g141 ( 
.A1(n_103),
.A2(n_105),
.B(n_49),
.Y(n_141)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_30),
.Y(n_104)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_104),
.Y(n_184)
);

BUFx8_ASAP7_75t_L g105 ( 
.A(n_38),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_51),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_30),
.B(n_17),
.Y(n_107)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_31),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_108),
.B(n_110),
.Y(n_167)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_28),
.Y(n_109)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_109),
.Y(n_166)
);

BUFx4f_ASAP7_75t_SL g110 ( 
.A(n_31),
.Y(n_110)
);

BUFx5_ASAP7_75t_L g111 ( 
.A(n_48),
.Y(n_111)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_111),
.Y(n_173)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_37),
.Y(n_112)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_112),
.Y(n_174)
);

INVx6_ASAP7_75t_SL g113 ( 
.A(n_22),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_113),
.B(n_16),
.Y(n_168)
);

INVx5_ASAP7_75t_L g114 ( 
.A(n_48),
.Y(n_114)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_114),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_112),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_SL g210 ( 
.A(n_119),
.B(n_128),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_123),
.A2(n_132),
.B1(n_144),
.B2(n_189),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_SL g128 ( 
.A(n_101),
.B(n_52),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_63),
.A2(n_25),
.B1(n_47),
.B2(n_46),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_64),
.A2(n_37),
.B1(n_47),
.B2(n_46),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g228 ( 
.A1(n_133),
.A2(n_134),
.B1(n_147),
.B2(n_149),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_74),
.A2(n_49),
.B1(n_40),
.B2(n_45),
.Y(n_134)
);

AOI21xp33_ASAP7_75t_SL g226 ( 
.A1(n_141),
.A2(n_172),
.B(n_179),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_98),
.B(n_40),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_143),
.B(n_152),
.Y(n_238)
);

OAI22xp33_ASAP7_75t_SL g144 ( 
.A1(n_87),
.A2(n_45),
.B1(n_29),
.B2(n_15),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_110),
.B(n_29),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_SL g235 ( 
.A(n_146),
.B(n_150),
.Y(n_235)
);

AOI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_102),
.A2(n_105),
.B1(n_61),
.B2(n_88),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_97),
.A2(n_7),
.B1(n_12),
.B2(n_15),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_110),
.B(n_72),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_83),
.B(n_7),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_85),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_SL g239 ( 
.A(n_157),
.B(n_163),
.Y(n_239)
);

OR2x2_ASAP7_75t_L g159 ( 
.A(n_102),
.B(n_12),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_159),
.B(n_168),
.Y(n_193)
);

AOI22xp33_ASAP7_75t_SL g161 ( 
.A1(n_105),
.A2(n_16),
.B1(n_17),
.B2(n_56),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g243 ( 
.A1(n_161),
.A2(n_164),
.B1(n_169),
.B2(n_171),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_114),
.Y(n_163)
);

AOI22xp33_ASAP7_75t_SL g164 ( 
.A1(n_68),
.A2(n_16),
.B1(n_90),
.B2(n_60),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_66),
.A2(n_69),
.B1(n_70),
.B2(n_65),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_84),
.B(n_86),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_170),
.B(n_129),
.Y(n_194)
);

AOI22xp33_ASAP7_75t_SL g171 ( 
.A1(n_84),
.A2(n_86),
.B1(n_96),
.B2(n_111),
.Y(n_171)
);

AOI22xp33_ASAP7_75t_SL g176 ( 
.A1(n_96),
.A2(n_102),
.B1(n_105),
.B2(n_61),
.Y(n_176)
);

AOI22xp33_ASAP7_75t_SL g213 ( 
.A1(n_176),
.A2(n_182),
.B1(n_165),
.B2(n_154),
.Y(n_213)
);

AOI22xp33_ASAP7_75t_SL g182 ( 
.A1(n_79),
.A2(n_102),
.B1(n_105),
.B2(n_61),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_79),
.B(n_55),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_183),
.B(n_165),
.Y(n_218)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_109),
.Y(n_188)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_188),
.Y(n_223)
);

OAI22xp33_ASAP7_75t_L g189 ( 
.A1(n_99),
.A2(n_106),
.B1(n_100),
.B2(n_57),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_L g190 ( 
.A1(n_75),
.A2(n_57),
.B1(n_58),
.B2(n_100),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_190),
.A2(n_117),
.B1(n_130),
.B2(n_120),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_167),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g264 ( 
.A(n_191),
.B(n_196),
.Y(n_264)
);

INVx4_ASAP7_75t_L g192 ( 
.A(n_135),
.Y(n_192)
);

INVx4_ASAP7_75t_L g258 ( 
.A(n_192),
.Y(n_258)
);

INVxp67_ASAP7_75t_L g265 ( 
.A(n_194),
.Y(n_265)
);

BUFx6f_ASAP7_75t_L g195 ( 
.A(n_151),
.Y(n_195)
);

INVx4_ASAP7_75t_L g289 ( 
.A(n_195),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_142),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_116),
.B(n_184),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_197),
.B(n_199),
.Y(n_257)
);

INVx8_ASAP7_75t_L g198 ( 
.A(n_165),
.Y(n_198)
);

INVx3_ASAP7_75t_L g290 ( 
.A(n_198),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_181),
.B(n_125),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_131),
.B(n_139),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_200),
.B(n_208),
.Y(n_261)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_115),
.B(n_137),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_201),
.B(n_216),
.C(n_249),
.Y(n_259)
);

BUFx3_ASAP7_75t_L g202 ( 
.A(n_129),
.Y(n_202)
);

HB1xp67_ASAP7_75t_L g293 ( 
.A(n_202),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_127),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g276 ( 
.A(n_203),
.B(n_218),
.Y(n_276)
);

INVxp67_ASAP7_75t_L g204 ( 
.A(n_182),
.Y(n_204)
);

INVxp33_ASAP7_75t_L g283 ( 
.A(n_204),
.Y(n_283)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_174),
.Y(n_205)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_205),
.Y(n_254)
);

INVx3_ASAP7_75t_L g206 ( 
.A(n_135),
.Y(n_206)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_206),
.Y(n_280)
);

INVxp67_ASAP7_75t_L g208 ( 
.A(n_176),
.Y(n_208)
);

BUFx6f_ASAP7_75t_L g209 ( 
.A(n_151),
.Y(n_209)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_209),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_R g211 ( 
.A(n_162),
.B(n_153),
.Y(n_211)
);

CKINVDCx14_ASAP7_75t_R g271 ( 
.A(n_211),
.Y(n_271)
);

OAI22xp33_ASAP7_75t_SL g212 ( 
.A1(n_159),
.A2(n_189),
.B1(n_148),
.B2(n_161),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_212),
.A2(n_220),
.B1(n_253),
.B2(n_218),
.Y(n_273)
);

OAI21xp33_ASAP7_75t_SL g267 ( 
.A1(n_213),
.A2(n_226),
.B(n_241),
.Y(n_267)
);

INVx13_ASAP7_75t_L g214 ( 
.A(n_156),
.Y(n_214)
);

INVx13_ASAP7_75t_L g266 ( 
.A(n_214),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_136),
.B(n_138),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_215),
.B(n_219),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_126),
.B(n_166),
.C(n_155),
.Y(n_216)
);

AND2x2_ASAP7_75t_L g217 ( 
.A(n_162),
.B(n_121),
.Y(n_217)
);

AND2x2_ASAP7_75t_L g274 ( 
.A(n_217),
.B(n_229),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_122),
.B(n_118),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_158),
.A2(n_178),
.B1(n_175),
.B2(n_144),
.Y(n_220)
);

BUFx5_ASAP7_75t_L g221 ( 
.A(n_173),
.Y(n_221)
);

INVx13_ASAP7_75t_L g279 ( 
.A(n_221),
.Y(n_279)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_145),
.Y(n_222)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_222),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_186),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_224),
.B(n_225),
.Y(n_281)
);

INVxp67_ASAP7_75t_L g225 ( 
.A(n_147),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_178),
.B(n_140),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_227),
.B(n_245),
.Y(n_262)
);

AND2x2_ASAP7_75t_L g229 ( 
.A(n_121),
.B(n_186),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_122),
.B(n_140),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_230),
.B(n_237),
.Y(n_284)
);

INVx6_ASAP7_75t_L g231 ( 
.A(n_172),
.Y(n_231)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_231),
.Y(n_256)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_145),
.Y(n_232)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_232),
.Y(n_269)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_175),
.Y(n_233)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_233),
.Y(n_278)
);

BUFx6f_ASAP7_75t_L g234 ( 
.A(n_160),
.Y(n_234)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_234),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_L g263 ( 
.A1(n_236),
.A2(n_225),
.B1(n_207),
.B2(n_208),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_130),
.B(n_124),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_124),
.B(n_160),
.Y(n_240)
);

BUFx24_ASAP7_75t_SL g270 ( 
.A(n_240),
.Y(n_270)
);

AOI22xp33_ASAP7_75t_SL g241 ( 
.A1(n_154),
.A2(n_120),
.B1(n_180),
.B2(n_177),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_177),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_242),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_187),
.Y(n_244)
);

INVx13_ASAP7_75t_L g291 ( 
.A(n_244),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_180),
.B(n_156),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_164),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_246),
.B(n_248),
.Y(n_272)
);

AND2x6_ASAP7_75t_L g247 ( 
.A(n_171),
.B(n_156),
.Y(n_247)
);

AND2x6_ASAP7_75t_L g299 ( 
.A(n_247),
.B(n_204),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_185),
.B(n_162),
.Y(n_248)
);

AND2x2_ASAP7_75t_L g249 ( 
.A(n_185),
.B(n_150),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_174),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_250),
.B(n_251),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_162),
.B(n_152),
.Y(n_251)
);

BUFx12f_ASAP7_75t_L g252 ( 
.A(n_118),
.Y(n_252)
);

INVx13_ASAP7_75t_L g292 ( 
.A(n_252),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_152),
.A2(n_106),
.B1(n_100),
.B2(n_99),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g260 ( 
.A(n_201),
.B(n_251),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g329 ( 
.A(n_260),
.B(n_282),
.Y(n_329)
);

AOI22xp33_ASAP7_75t_L g321 ( 
.A1(n_263),
.A2(n_283),
.B1(n_261),
.B2(n_262),
.Y(n_321)
);

AOI22xp5_ASAP7_75t_L g306 ( 
.A1(n_273),
.A2(n_297),
.B1(n_233),
.B2(n_206),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_217),
.B(n_216),
.C(n_248),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_238),
.B(n_253),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_285),
.B(n_286),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_227),
.B(n_249),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_249),
.B(n_211),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_288),
.B(n_252),
.Y(n_313)
);

OA21x2_ASAP7_75t_L g295 ( 
.A1(n_207),
.A2(n_246),
.B(n_220),
.Y(n_295)
);

OR2x2_ASAP7_75t_L g301 ( 
.A(n_295),
.B(n_239),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_217),
.B(n_196),
.C(n_223),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_296),
.B(n_298),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_L g297 ( 
.A1(n_228),
.A2(n_235),
.B1(n_236),
.B2(n_243),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_223),
.B(n_250),
.C(n_205),
.Y(n_298)
);

BUFx5_ASAP7_75t_L g324 ( 
.A(n_299),
.Y(n_324)
);

INVxp67_ASAP7_75t_L g300 ( 
.A(n_293),
.Y(n_300)
);

AOI21xp5_ASAP7_75t_L g336 ( 
.A1(n_301),
.A2(n_314),
.B(n_322),
.Y(n_336)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_254),
.Y(n_302)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_302),
.Y(n_356)
);

OAI22xp5_ASAP7_75t_L g304 ( 
.A1(n_295),
.A2(n_247),
.B1(n_210),
.B2(n_193),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_L g340 ( 
.A1(n_304),
.A2(n_312),
.B1(n_319),
.B2(n_333),
.Y(n_340)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_254),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g338 ( 
.A(n_305),
.B(n_317),
.Y(n_338)
);

OAI22xp5_ASAP7_75t_SL g348 ( 
.A1(n_306),
.A2(n_309),
.B1(n_310),
.B2(n_311),
.Y(n_348)
);

INVx2_ASAP7_75t_L g308 ( 
.A(n_278),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_L g309 ( 
.A1(n_295),
.A2(n_222),
.B1(n_195),
.B2(n_209),
.Y(n_309)
);

AOI22xp5_ASAP7_75t_L g310 ( 
.A1(n_273),
.A2(n_224),
.B1(n_232),
.B2(n_229),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_L g311 ( 
.A1(n_272),
.A2(n_229),
.B1(n_192),
.B2(n_234),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_L g312 ( 
.A1(n_272),
.A2(n_202),
.B1(n_198),
.B2(n_231),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_SL g355 ( 
.A(n_313),
.B(n_315),
.Y(n_355)
);

AOI21xp5_ASAP7_75t_L g314 ( 
.A1(n_281),
.A2(n_214),
.B(n_252),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_265),
.B(n_221),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_262),
.B(n_286),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_316),
.B(n_258),
.Y(n_346)
);

CKINVDCx20_ASAP7_75t_R g317 ( 
.A(n_264),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_265),
.B(n_257),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_SL g358 ( 
.A(n_318),
.B(n_332),
.Y(n_358)
);

OAI22xp5_ASAP7_75t_L g319 ( 
.A1(n_259),
.A2(n_282),
.B1(n_271),
.B2(n_288),
.Y(n_319)
);

INVxp33_ASAP7_75t_L g320 ( 
.A(n_284),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g350 ( 
.A(n_320),
.B(n_325),
.Y(n_350)
);

OAI21xp5_ASAP7_75t_SL g337 ( 
.A1(n_321),
.A2(n_323),
.B(n_316),
.Y(n_337)
);

AOI21xp5_ASAP7_75t_L g322 ( 
.A1(n_283),
.A2(n_267),
.B(n_274),
.Y(n_322)
);

OAI21xp5_ASAP7_75t_L g323 ( 
.A1(n_276),
.A2(n_274),
.B(n_285),
.Y(n_323)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_255),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_269),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_SL g342 ( 
.A(n_326),
.B(n_327),
.Y(n_342)
);

CKINVDCx16_ASAP7_75t_R g327 ( 
.A(n_275),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_298),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_SL g345 ( 
.A(n_328),
.B(n_330),
.Y(n_345)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_280),
.Y(n_330)
);

INVxp67_ASAP7_75t_L g331 ( 
.A(n_290),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g335 ( 
.A(n_331),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_270),
.B(n_268),
.Y(n_332)
);

AOI22xp5_ASAP7_75t_L g333 ( 
.A1(n_259),
.A2(n_277),
.B1(n_260),
.B2(n_274),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_280),
.Y(n_334)
);

OAI21xp33_ASAP7_75t_SL g368 ( 
.A1(n_337),
.A2(n_339),
.B(n_343),
.Y(n_368)
);

OAI21xp5_ASAP7_75t_SL g339 ( 
.A1(n_322),
.A2(n_299),
.B(n_277),
.Y(n_339)
);

XOR2xp5_ASAP7_75t_L g341 ( 
.A(n_329),
.B(n_296),
.Y(n_341)
);

MAJIxp5_ASAP7_75t_L g370 ( 
.A(n_341),
.B(n_344),
.C(n_311),
.Y(n_370)
);

OAI21xp5_ASAP7_75t_SL g343 ( 
.A1(n_301),
.A2(n_291),
.B(n_256),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g344 ( 
.A(n_329),
.B(n_258),
.C(n_290),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_346),
.B(n_353),
.Y(n_363)
);

AOI22xp5_ASAP7_75t_L g347 ( 
.A1(n_306),
.A2(n_294),
.B1(n_287),
.B2(n_289),
.Y(n_347)
);

OAI22xp5_ASAP7_75t_SL g371 ( 
.A1(n_347),
.A2(n_352),
.B1(n_354),
.B2(n_302),
.Y(n_371)
);

AOI21xp5_ASAP7_75t_L g349 ( 
.A1(n_301),
.A2(n_266),
.B(n_291),
.Y(n_349)
);

AOI21xp5_ASAP7_75t_L g360 ( 
.A1(n_349),
.A2(n_314),
.B(n_312),
.Y(n_360)
);

OAI21xp5_ASAP7_75t_SL g351 ( 
.A1(n_313),
.A2(n_266),
.B(n_294),
.Y(n_351)
);

CKINVDCx14_ASAP7_75t_R g359 ( 
.A(n_351),
.Y(n_359)
);

AOI22xp5_ASAP7_75t_L g352 ( 
.A1(n_307),
.A2(n_279),
.B1(n_292),
.B2(n_304),
.Y(n_352)
);

CKINVDCx20_ASAP7_75t_R g353 ( 
.A(n_331),
.Y(n_353)
);

AOI22xp5_ASAP7_75t_L g354 ( 
.A1(n_307),
.A2(n_279),
.B1(n_292),
.B2(n_310),
.Y(n_354)
);

CKINVDCx20_ASAP7_75t_R g357 ( 
.A(n_300),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_357),
.B(n_325),
.Y(n_365)
);

OAI21xp5_ASAP7_75t_SL g395 ( 
.A1(n_360),
.A2(n_336),
.B(n_351),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_SL g361 ( 
.A(n_343),
.B(n_323),
.Y(n_361)
);

CKINVDCx14_ASAP7_75t_R g391 ( 
.A(n_361),
.Y(n_391)
);

CKINVDCx20_ASAP7_75t_R g362 ( 
.A(n_338),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_362),
.B(n_371),
.Y(n_380)
);

AOI22xp5_ASAP7_75t_L g364 ( 
.A1(n_348),
.A2(n_309),
.B1(n_319),
.B2(n_328),
.Y(n_364)
);

OAI22xp5_ASAP7_75t_SL g383 ( 
.A1(n_364),
.A2(n_369),
.B1(n_340),
.B2(n_345),
.Y(n_383)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_365),
.Y(n_381)
);

CKINVDCx16_ASAP7_75t_R g366 ( 
.A(n_342),
.Y(n_366)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_366),
.Y(n_392)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_356),
.Y(n_367)
);

INVx1_ASAP7_75t_SL g386 ( 
.A(n_367),
.Y(n_386)
);

AOI22xp5_ASAP7_75t_L g369 ( 
.A1(n_348),
.A2(n_303),
.B1(n_333),
.B2(n_317),
.Y(n_369)
);

MAJIxp5_ASAP7_75t_L g379 ( 
.A(n_370),
.B(n_372),
.C(n_374),
.Y(n_379)
);

MAJIxp5_ASAP7_75t_L g372 ( 
.A(n_341),
.B(n_324),
.C(n_305),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_338),
.B(n_326),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_373),
.B(n_375),
.Y(n_390)
);

MAJIxp5_ASAP7_75t_L g374 ( 
.A(n_341),
.B(n_324),
.C(n_330),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_356),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_SL g376 ( 
.A(n_355),
.B(n_334),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_SL g393 ( 
.A(n_376),
.B(n_378),
.Y(n_393)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_346),
.Y(n_377)
);

INVxp67_ASAP7_75t_L g387 ( 
.A(n_377),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_357),
.B(n_308),
.Y(n_378)
);

XNOR2xp5_ASAP7_75t_L g382 ( 
.A(n_369),
.B(n_337),
.Y(n_382)
);

MAJIxp5_ASAP7_75t_L g408 ( 
.A(n_382),
.B(n_388),
.C(n_370),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_SL g398 ( 
.A(n_383),
.B(n_362),
.Y(n_398)
);

OAI22xp5_ASAP7_75t_SL g384 ( 
.A1(n_364),
.A2(n_340),
.B1(n_359),
.B2(n_377),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_384),
.B(n_394),
.Y(n_402)
);

CKINVDCx16_ASAP7_75t_R g385 ( 
.A(n_365),
.Y(n_385)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_385),
.Y(n_396)
);

MAJIxp5_ASAP7_75t_L g388 ( 
.A(n_370),
.B(n_344),
.C(n_345),
.Y(n_388)
);

AOI21xp5_ASAP7_75t_L g389 ( 
.A1(n_359),
.A2(n_349),
.B(n_336),
.Y(n_389)
);

INVxp67_ASAP7_75t_L g404 ( 
.A(n_389),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_SL g394 ( 
.A(n_366),
.B(n_355),
.Y(n_394)
);

MAJIxp5_ASAP7_75t_SL g399 ( 
.A(n_395),
.B(n_368),
.C(n_371),
.Y(n_399)
);

INVx13_ASAP7_75t_L g397 ( 
.A(n_386),
.Y(n_397)
);

HB1xp67_ASAP7_75t_L g412 ( 
.A(n_397),
.Y(n_412)
);

OAI22xp5_ASAP7_75t_SL g415 ( 
.A1(n_398),
.A2(n_391),
.B1(n_381),
.B2(n_387),
.Y(n_415)
);

XNOR2x1_ASAP7_75t_L g413 ( 
.A(n_399),
.B(n_389),
.Y(n_413)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_390),
.Y(n_400)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_400),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_SL g401 ( 
.A(n_394),
.B(n_358),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_SL g410 ( 
.A(n_401),
.B(n_358),
.Y(n_410)
);

BUFx4f_ASAP7_75t_SL g403 ( 
.A(n_392),
.Y(n_403)
);

NOR2xp33_ASAP7_75t_L g414 ( 
.A(n_403),
.B(n_405),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_385),
.B(n_373),
.Y(n_405)
);

OAI22xp5_ASAP7_75t_L g406 ( 
.A1(n_380),
.A2(n_363),
.B1(n_372),
.B2(n_374),
.Y(n_406)
);

AOI22xp5_ASAP7_75t_SL g409 ( 
.A1(n_406),
.A2(n_407),
.B1(n_383),
.B2(n_384),
.Y(n_409)
);

OAI22xp5_ASAP7_75t_SL g407 ( 
.A1(n_380),
.A2(n_363),
.B1(n_361),
.B2(n_352),
.Y(n_407)
);

MAJIxp5_ASAP7_75t_L g411 ( 
.A(n_408),
.B(n_379),
.C(n_388),
.Y(n_411)
);

XNOR2xp5_ASAP7_75t_L g424 ( 
.A(n_409),
.B(n_413),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_410),
.B(n_411),
.Y(n_421)
);

NOR2xp33_ASAP7_75t_L g419 ( 
.A(n_415),
.B(n_416),
.Y(n_419)
);

NOR2xp33_ASAP7_75t_L g416 ( 
.A(n_402),
.B(n_350),
.Y(n_416)
);

XOR2xp5_ASAP7_75t_L g418 ( 
.A(n_406),
.B(n_379),
.Y(n_418)
);

MAJIxp5_ASAP7_75t_L g426 ( 
.A(n_418),
.B(n_408),
.C(n_374),
.Y(n_426)
);

AO21x1_ASAP7_75t_L g420 ( 
.A1(n_409),
.A2(n_402),
.B(n_404),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_420),
.B(n_422),
.Y(n_431)
);

NOR2xp33_ASAP7_75t_L g422 ( 
.A(n_411),
.B(n_342),
.Y(n_422)
);

NOR2xp33_ASAP7_75t_L g423 ( 
.A(n_415),
.B(n_350),
.Y(n_423)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_423),
.Y(n_427)
);

NOR2xp33_ASAP7_75t_L g425 ( 
.A(n_418),
.B(n_335),
.Y(n_425)
);

OAI21xp5_ASAP7_75t_SL g432 ( 
.A1(n_425),
.A2(n_376),
.B(n_414),
.Y(n_432)
);

INVxp67_ASAP7_75t_L g430 ( 
.A(n_426),
.Y(n_430)
);

OAI22xp5_ASAP7_75t_SL g428 ( 
.A1(n_419),
.A2(n_417),
.B1(n_400),
.B2(n_396),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_428),
.B(n_429),
.Y(n_433)
);

AOI22xp5_ASAP7_75t_SL g429 ( 
.A1(n_424),
.A2(n_404),
.B1(n_391),
.B2(n_413),
.Y(n_429)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_432),
.Y(n_434)
);

NAND3xp33_ASAP7_75t_L g435 ( 
.A(n_430),
.B(n_421),
.C(n_426),
.Y(n_435)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_435),
.Y(n_437)
);

AOI21xp5_ASAP7_75t_SL g436 ( 
.A1(n_431),
.A2(n_396),
.B(n_405),
.Y(n_436)
);

AOI322xp5_ASAP7_75t_L g438 ( 
.A1(n_436),
.A2(n_403),
.A3(n_397),
.B1(n_392),
.B2(n_393),
.C1(n_381),
.C2(n_390),
.Y(n_438)
);

INVxp67_ASAP7_75t_L g439 ( 
.A(n_438),
.Y(n_439)
);

NOR2xp33_ASAP7_75t_L g440 ( 
.A(n_437),
.B(n_427),
.Y(n_440)
);

MAJIxp5_ASAP7_75t_L g441 ( 
.A(n_440),
.B(n_430),
.C(n_434),
.Y(n_441)
);

O2A1O1Ixp33_ASAP7_75t_L g442 ( 
.A1(n_441),
.A2(n_439),
.B(n_433),
.C(n_412),
.Y(n_442)
);

XNOR2xp5_ASAP7_75t_L g443 ( 
.A(n_442),
.B(n_403),
.Y(n_443)
);


endmodule