module fake_jpeg_25965_n_182 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_182);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_182;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_175;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_145;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx12_ASAP7_75t_L g14 ( 
.A(n_8),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_2),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

BUFx10_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_25),
.Y(n_29)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_29),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_21),
.B(n_0),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_SL g56 ( 
.A(n_30),
.B(n_37),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_21),
.Y(n_31)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_31),
.Y(n_43)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_21),
.Y(n_32)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_32),
.Y(n_49)
);

INVx11_ASAP7_75t_L g33 ( 
.A(n_21),
.Y(n_33)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_33),
.Y(n_46)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_25),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_34),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_14),
.Y(n_35)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_35),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_25),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_36),
.B(n_27),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_SL g37 ( 
.A(n_18),
.B(n_0),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_25),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_38),
.Y(n_47)
);

BUFx2_ASAP7_75t_L g39 ( 
.A(n_25),
.Y(n_39)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_39),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_30),
.B(n_24),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_40),
.B(n_50),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_37),
.B(n_28),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_42),
.B(n_44),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_36),
.B(n_28),
.Y(n_44)
);

AND2x2_ASAP7_75t_L g50 ( 
.A(n_38),
.B(n_24),
.Y(n_50)
);

OR2x2_ASAP7_75t_L g65 ( 
.A(n_50),
.B(n_57),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_33),
.Y(n_51)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_51),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_36),
.B(n_19),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_52),
.B(n_18),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_33),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_53),
.Y(n_66)
);

BUFx2_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_54),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_58),
.B(n_60),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_56),
.B(n_19),
.Y(n_60)
);

INVxp67_ASAP7_75t_L g61 ( 
.A(n_50),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_61),
.B(n_62),
.Y(n_92)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_49),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_SL g80 ( 
.A(n_64),
.B(n_32),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g67 ( 
.A1(n_40),
.A2(n_34),
.B1(n_22),
.B2(n_29),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_67),
.A2(n_70),
.B1(n_71),
.B2(n_48),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_41),
.B(n_31),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_68),
.B(n_73),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_43),
.A2(n_34),
.B1(n_22),
.B2(n_29),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_43),
.A2(n_29),
.B1(n_32),
.B2(n_55),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_54),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_72),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_49),
.B(n_31),
.Y(n_73)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_45),
.Y(n_74)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_74),
.Y(n_82)
);

AND2x2_ASAP7_75t_SL g76 ( 
.A(n_67),
.B(n_31),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_76),
.B(n_81),
.Y(n_101)
);

INVxp33_ASAP7_75t_SL g77 ( 
.A(n_68),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_77),
.B(n_78),
.Y(n_98)
);

INVxp67_ASAP7_75t_L g78 ( 
.A(n_73),
.Y(n_78)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_79),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_80),
.B(n_89),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_65),
.A2(n_48),
.B1(n_55),
.B2(n_46),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_64),
.B(n_38),
.C(n_45),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_83),
.B(n_86),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_65),
.A2(n_46),
.B1(n_39),
.B2(n_16),
.Y(n_86)
);

AOI21xp5_ASAP7_75t_SL g87 ( 
.A1(n_65),
.A2(n_16),
.B(n_15),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_L g96 ( 
.A1(n_87),
.A2(n_27),
.B(n_23),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_70),
.A2(n_71),
.B1(n_74),
.B2(n_62),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_88),
.B(n_91),
.Y(n_105)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_72),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_SL g90 ( 
.A(n_69),
.B(n_15),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_SL g100 ( 
.A(n_90),
.B(n_23),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_69),
.B(n_35),
.Y(n_91)
);

O2A1O1Ixp33_ASAP7_75t_L g93 ( 
.A1(n_78),
.A2(n_66),
.B(n_59),
.C(n_63),
.Y(n_93)
);

OAI21xp5_ASAP7_75t_SL g115 ( 
.A1(n_93),
.A2(n_76),
.B(n_92),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_85),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_95),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_SL g125 ( 
.A(n_96),
.B(n_100),
.Y(n_125)
);

BUFx24_ASAP7_75t_SL g97 ( 
.A(n_90),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_97),
.B(n_104),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_85),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_99),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_75),
.B(n_59),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_103),
.B(n_106),
.Y(n_116)
);

NOR3xp33_ASAP7_75t_L g104 ( 
.A(n_91),
.B(n_17),
.C(n_47),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_81),
.B(n_89),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_84),
.B(n_66),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_107),
.B(n_80),
.Y(n_113)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_84),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_108),
.B(n_109),
.Y(n_118)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_88),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_113),
.B(n_115),
.Y(n_130)
);

XOR2xp5_ASAP7_75t_L g114 ( 
.A(n_102),
.B(n_83),
.Y(n_114)
);

XOR2xp5_ASAP7_75t_L g133 ( 
.A(n_114),
.B(n_98),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_95),
.B(n_86),
.Y(n_117)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_117),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_L g119 ( 
.A1(n_102),
.A2(n_87),
.B(n_76),
.Y(n_119)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_119),
.Y(n_134)
);

A2O1A1O1Ixp25_ASAP7_75t_L g121 ( 
.A1(n_101),
.A2(n_76),
.B(n_79),
.C(n_39),
.D(n_38),
.Y(n_121)
);

OAI221xp5_ASAP7_75t_L g141 ( 
.A1(n_121),
.A2(n_94),
.B1(n_38),
.B2(n_51),
.C(n_35),
.Y(n_141)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_93),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_122),
.B(n_124),
.Y(n_131)
);

INVxp67_ASAP7_75t_SL g123 ( 
.A(n_99),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_123),
.B(n_126),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_107),
.B(n_82),
.Y(n_124)
);

AOI21xp5_ASAP7_75t_L g126 ( 
.A1(n_101),
.A2(n_82),
.B(n_63),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_105),
.B(n_53),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_105),
.B(n_26),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_128),
.B(n_35),
.Y(n_143)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_124),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_129),
.B(n_132),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_111),
.Y(n_132)
);

XOR2xp5_ASAP7_75t_L g150 ( 
.A(n_133),
.B(n_141),
.Y(n_150)
);

NOR2xp67_ASAP7_75t_SL g135 ( 
.A(n_111),
.B(n_96),
.Y(n_135)
);

AOI21xp5_ASAP7_75t_L g149 ( 
.A1(n_135),
.A2(n_125),
.B(n_118),
.Y(n_149)
);

INVx2_ASAP7_75t_SL g136 ( 
.A(n_120),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_120),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_137),
.B(n_140),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_114),
.B(n_108),
.C(n_110),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_138),
.B(n_119),
.C(n_116),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_122),
.A2(n_94),
.B1(n_109),
.B2(n_17),
.Y(n_140)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_143),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_118),
.A2(n_38),
.B1(n_26),
.B2(n_14),
.Y(n_144)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_144),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_L g161 ( 
.A(n_145),
.B(n_148),
.Y(n_161)
);

NAND3xp33_ASAP7_75t_L g146 ( 
.A(n_130),
.B(n_131),
.C(n_113),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_SL g164 ( 
.A1(n_146),
.A2(n_149),
.B(n_14),
.Y(n_164)
);

MAJx2_ASAP7_75t_L g148 ( 
.A(n_138),
.B(n_115),
.C(n_116),
.Y(n_148)
);

INVxp67_ASAP7_75t_SL g152 ( 
.A(n_136),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_152),
.B(n_47),
.Y(n_165)
);

NOR3xp33_ASAP7_75t_SL g153 ( 
.A(n_139),
.B(n_125),
.C(n_112),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_153),
.B(n_147),
.Y(n_162)
);

XOR2xp5_ASAP7_75t_L g156 ( 
.A(n_133),
.B(n_130),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_156),
.B(n_157),
.C(n_158),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_129),
.B(n_126),
.C(n_127),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_144),
.B(n_121),
.C(n_47),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_155),
.A2(n_134),
.B1(n_131),
.B2(n_142),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_SL g160 ( 
.A(n_154),
.B(n_136),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_160),
.B(n_165),
.Y(n_170)
);

BUFx24_ASAP7_75t_SL g171 ( 
.A(n_162),
.Y(n_171)
);

AOI21xp5_ASAP7_75t_L g168 ( 
.A1(n_164),
.A2(n_1),
.B(n_3),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_151),
.B(n_9),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_L g167 ( 
.A(n_166),
.B(n_150),
.Y(n_167)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_167),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_168),
.B(n_169),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_159),
.A2(n_11),
.B1(n_20),
.B2(n_4),
.Y(n_169)
);

OR2x2_ASAP7_75t_L g173 ( 
.A(n_171),
.B(n_163),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_SL g176 ( 
.A(n_173),
.B(n_175),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_170),
.B(n_161),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_L g177 ( 
.A1(n_172),
.A2(n_7),
.B(n_5),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_177),
.B(n_178),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_174),
.B(n_6),
.C(n_7),
.Y(n_178)
);

INVxp67_ASAP7_75t_L g179 ( 
.A(n_176),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_179),
.B(n_7),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g182 ( 
.A(n_181),
.B(n_180),
.Y(n_182)
);


endmodule