module fake_netlist_6_3376_n_5237 (n_52, n_591, n_435, n_1, n_91, n_326, n_256, n_440, n_587, n_695, n_507, n_580, n_209, n_367, n_465, n_680, n_590, n_625, n_63, n_661, n_223, n_278, n_341, n_362, n_148, n_226, n_161, n_22, n_208, n_462, n_68, n_607, n_671, n_316, n_419, n_28, n_304, n_212, n_50, n_694, n_7, n_578, n_144, n_365, n_125, n_168, n_384, n_297, n_595, n_627, n_524, n_342, n_77, n_106, n_358, n_160, n_449, n_131, n_188, n_310, n_509, n_186, n_245, n_0, n_368, n_575, n_677, n_396, n_495, n_350, n_78, n_84, n_585, n_568, n_392, n_442, n_480, n_142, n_143, n_382, n_673, n_180, n_62, n_628, n_557, n_349, n_643, n_233, n_617, n_698, n_255, n_284, n_400, n_140, n_337, n_214, n_485, n_67, n_15, n_443, n_246, n_38, n_471, n_289, n_421, n_424, n_615, n_59, n_181, n_182, n_238, n_573, n_202, n_320, n_108, n_639, n_676, n_327, n_369, n_597, n_685, n_280, n_287, n_353, n_610, n_555, n_389, n_415, n_65, n_230, n_605, n_461, n_141, n_383, n_669, n_200, n_447, n_176, n_114, n_86, n_198, n_104, n_222, n_179, n_248, n_300, n_517, n_667, n_71, n_74, n_229, n_542, n_644, n_682, n_621, n_305, n_72, n_532, n_173, n_535, n_691, n_250, n_372, n_468, n_544, n_111, n_504, n_314, n_378, n_413, n_377, n_35, n_183, n_510, n_79, n_375, n_601, n_338, n_522, n_466, n_506, n_56, n_360, n_603, n_119, n_235, n_536, n_622, n_147, n_191, n_340, n_387, n_452, n_616, n_658, n_39, n_344, n_73, n_581, n_428, n_609, n_432, n_641, n_693, n_101, n_167, n_631, n_174, n_127, n_516, n_153, n_525, n_611, n_156, n_491, n_145, n_42, n_133, n_656, n_96, n_8, n_666, n_371, n_567, n_189, n_405, n_213, n_538, n_294, n_302, n_499, n_380, n_129, n_647, n_197, n_11, n_137, n_17, n_343, n_448, n_20, n_494, n_539, n_493, n_397, n_155, n_109, n_614, n_529, n_445, n_425, n_684, n_122, n_45, n_454, n_34, n_218, n_638, n_70, n_234, n_37, n_486, n_381, n_82, n_27, n_236, n_653, n_112, n_172, n_648, n_657, n_576, n_472, n_270, n_239, n_126, n_414, n_97, n_563, n_58, n_490, n_290, n_220, n_118, n_224, n_48, n_25, n_93, n_80, n_196, n_402, n_352, n_668, n_478, n_626, n_574, n_9, n_460, n_107, n_6, n_417, n_14, n_446, n_498, n_662, n_89, n_374, n_659, n_366, n_407, n_450, n_103, n_272, n_526, n_185, n_348, n_579, n_69, n_376, n_390, n_473, n_293, n_31, n_334, n_559, n_53, n_370, n_44, n_458, n_232, n_650, n_16, n_163, n_46, n_330, n_470, n_475, n_298, n_18, n_492, n_281, n_258, n_551, n_154, n_456, n_564, n_98, n_260, n_265, n_313, n_451, n_624, n_279, n_686, n_252, n_228, n_565, n_594, n_356, n_577, n_166, n_184, n_552, n_619, n_216, n_455, n_83, n_521, n_363, n_572, n_395, n_592, n_654, n_323, n_606, n_393, n_411, n_503, n_152, n_623, n_92, n_599, n_513, n_321, n_645, n_331, n_105, n_227, n_132, n_570, n_406, n_483, n_102, n_204, n_482, n_474, n_527, n_261, n_608, n_620, n_420, n_683, n_630, n_312, n_394, n_32, n_66, n_130, n_519, n_541, n_512, n_164, n_292, n_100, n_121, n_307, n_469, n_433, n_500, n_23, n_476, n_2, n_291, n_219, n_543, n_357, n_150, n_264, n_263, n_589, n_481, n_325, n_329, n_464, n_600, n_561, n_33, n_477, n_549, n_533, n_408, n_61, n_237, n_584, n_244, n_399, n_76, n_243, n_124, n_548, n_94, n_282, n_436, n_116, n_211, n_523, n_117, n_175, n_322, n_345, n_409, n_231, n_354, n_689, n_40, n_505, n_240, n_139, n_319, n_41, n_134, n_547, n_537, n_273, n_558, n_635, n_95, n_311, n_10, n_403, n_253, n_634, n_583, n_596, n_123, n_136, n_546, n_562, n_249, n_201, n_386, n_556, n_159, n_157, n_162, n_692, n_115, n_487, n_550, n_128, n_241, n_30, n_275, n_553, n_43, n_652, n_560, n_642, n_276, n_569, n_441, n_221, n_444, n_586, n_423, n_146, n_318, n_303, n_511, n_467, n_306, n_21, n_193, n_269, n_359, n_346, n_88, n_3, n_416, n_530, n_277, n_520, n_418, n_113, n_618, n_582, n_4, n_199, n_138, n_266, n_296, n_674, n_571, n_268, n_271, n_404, n_651, n_439, n_158, n_217, n_49, n_210, n_299, n_518, n_206, n_679, n_5, n_453, n_612, n_633, n_665, n_333, n_588, n_215, n_178, n_247, n_225, n_308, n_309, n_355, n_426, n_317, n_149, n_632, n_431, n_90, n_347, n_24, n_459, n_54, n_502, n_328, n_672, n_534, n_488, n_429, n_373, n_87, n_195, n_285, n_497, n_675, n_85, n_99, n_257, n_655, n_13, n_670, n_203, n_286, n_254, n_207, n_242, n_19, n_47, n_690, n_29, n_75, n_401, n_324, n_335, n_430, n_463, n_545, n_489, n_205, n_604, n_120, n_251, n_301, n_274, n_636, n_681, n_110, n_151, n_412, n_640, n_81, n_660, n_36, n_26, n_55, n_267, n_438, n_339, n_315, n_434, n_515, n_64, n_288, n_427, n_479, n_496, n_598, n_422, n_696, n_688, n_135, n_165, n_351, n_437, n_259, n_177, n_540, n_593, n_514, n_646, n_528, n_391, n_457, n_687, n_697, n_364, n_637, n_295, n_385, n_629, n_388, n_190, n_262, n_484, n_613, n_187, n_501, n_531, n_60, n_361, n_508, n_663, n_379, n_170, n_332, n_336, n_12, n_398, n_410, n_566, n_554, n_602, n_194, n_664, n_171, n_678, n_192, n_57, n_169, n_51, n_649, n_283, n_5237);

input n_52;
input n_591;
input n_435;
input n_1;
input n_91;
input n_326;
input n_256;
input n_440;
input n_587;
input n_695;
input n_507;
input n_580;
input n_209;
input n_367;
input n_465;
input n_680;
input n_590;
input n_625;
input n_63;
input n_661;
input n_223;
input n_278;
input n_341;
input n_362;
input n_148;
input n_226;
input n_161;
input n_22;
input n_208;
input n_462;
input n_68;
input n_607;
input n_671;
input n_316;
input n_419;
input n_28;
input n_304;
input n_212;
input n_50;
input n_694;
input n_7;
input n_578;
input n_144;
input n_365;
input n_125;
input n_168;
input n_384;
input n_297;
input n_595;
input n_627;
input n_524;
input n_342;
input n_77;
input n_106;
input n_358;
input n_160;
input n_449;
input n_131;
input n_188;
input n_310;
input n_509;
input n_186;
input n_245;
input n_0;
input n_368;
input n_575;
input n_677;
input n_396;
input n_495;
input n_350;
input n_78;
input n_84;
input n_585;
input n_568;
input n_392;
input n_442;
input n_480;
input n_142;
input n_143;
input n_382;
input n_673;
input n_180;
input n_62;
input n_628;
input n_557;
input n_349;
input n_643;
input n_233;
input n_617;
input n_698;
input n_255;
input n_284;
input n_400;
input n_140;
input n_337;
input n_214;
input n_485;
input n_67;
input n_15;
input n_443;
input n_246;
input n_38;
input n_471;
input n_289;
input n_421;
input n_424;
input n_615;
input n_59;
input n_181;
input n_182;
input n_238;
input n_573;
input n_202;
input n_320;
input n_108;
input n_639;
input n_676;
input n_327;
input n_369;
input n_597;
input n_685;
input n_280;
input n_287;
input n_353;
input n_610;
input n_555;
input n_389;
input n_415;
input n_65;
input n_230;
input n_605;
input n_461;
input n_141;
input n_383;
input n_669;
input n_200;
input n_447;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_222;
input n_179;
input n_248;
input n_300;
input n_517;
input n_667;
input n_71;
input n_74;
input n_229;
input n_542;
input n_644;
input n_682;
input n_621;
input n_305;
input n_72;
input n_532;
input n_173;
input n_535;
input n_691;
input n_250;
input n_372;
input n_468;
input n_544;
input n_111;
input n_504;
input n_314;
input n_378;
input n_413;
input n_377;
input n_35;
input n_183;
input n_510;
input n_79;
input n_375;
input n_601;
input n_338;
input n_522;
input n_466;
input n_506;
input n_56;
input n_360;
input n_603;
input n_119;
input n_235;
input n_536;
input n_622;
input n_147;
input n_191;
input n_340;
input n_387;
input n_452;
input n_616;
input n_658;
input n_39;
input n_344;
input n_73;
input n_581;
input n_428;
input n_609;
input n_432;
input n_641;
input n_693;
input n_101;
input n_167;
input n_631;
input n_174;
input n_127;
input n_516;
input n_153;
input n_525;
input n_611;
input n_156;
input n_491;
input n_145;
input n_42;
input n_133;
input n_656;
input n_96;
input n_8;
input n_666;
input n_371;
input n_567;
input n_189;
input n_405;
input n_213;
input n_538;
input n_294;
input n_302;
input n_499;
input n_380;
input n_129;
input n_647;
input n_197;
input n_11;
input n_137;
input n_17;
input n_343;
input n_448;
input n_20;
input n_494;
input n_539;
input n_493;
input n_397;
input n_155;
input n_109;
input n_614;
input n_529;
input n_445;
input n_425;
input n_684;
input n_122;
input n_45;
input n_454;
input n_34;
input n_218;
input n_638;
input n_70;
input n_234;
input n_37;
input n_486;
input n_381;
input n_82;
input n_27;
input n_236;
input n_653;
input n_112;
input n_172;
input n_648;
input n_657;
input n_576;
input n_472;
input n_270;
input n_239;
input n_126;
input n_414;
input n_97;
input n_563;
input n_58;
input n_490;
input n_290;
input n_220;
input n_118;
input n_224;
input n_48;
input n_25;
input n_93;
input n_80;
input n_196;
input n_402;
input n_352;
input n_668;
input n_478;
input n_626;
input n_574;
input n_9;
input n_460;
input n_107;
input n_6;
input n_417;
input n_14;
input n_446;
input n_498;
input n_662;
input n_89;
input n_374;
input n_659;
input n_366;
input n_407;
input n_450;
input n_103;
input n_272;
input n_526;
input n_185;
input n_348;
input n_579;
input n_69;
input n_376;
input n_390;
input n_473;
input n_293;
input n_31;
input n_334;
input n_559;
input n_53;
input n_370;
input n_44;
input n_458;
input n_232;
input n_650;
input n_16;
input n_163;
input n_46;
input n_330;
input n_470;
input n_475;
input n_298;
input n_18;
input n_492;
input n_281;
input n_258;
input n_551;
input n_154;
input n_456;
input n_564;
input n_98;
input n_260;
input n_265;
input n_313;
input n_451;
input n_624;
input n_279;
input n_686;
input n_252;
input n_228;
input n_565;
input n_594;
input n_356;
input n_577;
input n_166;
input n_184;
input n_552;
input n_619;
input n_216;
input n_455;
input n_83;
input n_521;
input n_363;
input n_572;
input n_395;
input n_592;
input n_654;
input n_323;
input n_606;
input n_393;
input n_411;
input n_503;
input n_152;
input n_623;
input n_92;
input n_599;
input n_513;
input n_321;
input n_645;
input n_331;
input n_105;
input n_227;
input n_132;
input n_570;
input n_406;
input n_483;
input n_102;
input n_204;
input n_482;
input n_474;
input n_527;
input n_261;
input n_608;
input n_620;
input n_420;
input n_683;
input n_630;
input n_312;
input n_394;
input n_32;
input n_66;
input n_130;
input n_519;
input n_541;
input n_512;
input n_164;
input n_292;
input n_100;
input n_121;
input n_307;
input n_469;
input n_433;
input n_500;
input n_23;
input n_476;
input n_2;
input n_291;
input n_219;
input n_543;
input n_357;
input n_150;
input n_264;
input n_263;
input n_589;
input n_481;
input n_325;
input n_329;
input n_464;
input n_600;
input n_561;
input n_33;
input n_477;
input n_549;
input n_533;
input n_408;
input n_61;
input n_237;
input n_584;
input n_244;
input n_399;
input n_76;
input n_243;
input n_124;
input n_548;
input n_94;
input n_282;
input n_436;
input n_116;
input n_211;
input n_523;
input n_117;
input n_175;
input n_322;
input n_345;
input n_409;
input n_231;
input n_354;
input n_689;
input n_40;
input n_505;
input n_240;
input n_139;
input n_319;
input n_41;
input n_134;
input n_547;
input n_537;
input n_273;
input n_558;
input n_635;
input n_95;
input n_311;
input n_10;
input n_403;
input n_253;
input n_634;
input n_583;
input n_596;
input n_123;
input n_136;
input n_546;
input n_562;
input n_249;
input n_201;
input n_386;
input n_556;
input n_159;
input n_157;
input n_162;
input n_692;
input n_115;
input n_487;
input n_550;
input n_128;
input n_241;
input n_30;
input n_275;
input n_553;
input n_43;
input n_652;
input n_560;
input n_642;
input n_276;
input n_569;
input n_441;
input n_221;
input n_444;
input n_586;
input n_423;
input n_146;
input n_318;
input n_303;
input n_511;
input n_467;
input n_306;
input n_21;
input n_193;
input n_269;
input n_359;
input n_346;
input n_88;
input n_3;
input n_416;
input n_530;
input n_277;
input n_520;
input n_418;
input n_113;
input n_618;
input n_582;
input n_4;
input n_199;
input n_138;
input n_266;
input n_296;
input n_674;
input n_571;
input n_268;
input n_271;
input n_404;
input n_651;
input n_439;
input n_158;
input n_217;
input n_49;
input n_210;
input n_299;
input n_518;
input n_206;
input n_679;
input n_5;
input n_453;
input n_612;
input n_633;
input n_665;
input n_333;
input n_588;
input n_215;
input n_178;
input n_247;
input n_225;
input n_308;
input n_309;
input n_355;
input n_426;
input n_317;
input n_149;
input n_632;
input n_431;
input n_90;
input n_347;
input n_24;
input n_459;
input n_54;
input n_502;
input n_328;
input n_672;
input n_534;
input n_488;
input n_429;
input n_373;
input n_87;
input n_195;
input n_285;
input n_497;
input n_675;
input n_85;
input n_99;
input n_257;
input n_655;
input n_13;
input n_670;
input n_203;
input n_286;
input n_254;
input n_207;
input n_242;
input n_19;
input n_47;
input n_690;
input n_29;
input n_75;
input n_401;
input n_324;
input n_335;
input n_430;
input n_463;
input n_545;
input n_489;
input n_205;
input n_604;
input n_120;
input n_251;
input n_301;
input n_274;
input n_636;
input n_681;
input n_110;
input n_151;
input n_412;
input n_640;
input n_81;
input n_660;
input n_36;
input n_26;
input n_55;
input n_267;
input n_438;
input n_339;
input n_315;
input n_434;
input n_515;
input n_64;
input n_288;
input n_427;
input n_479;
input n_496;
input n_598;
input n_422;
input n_696;
input n_688;
input n_135;
input n_165;
input n_351;
input n_437;
input n_259;
input n_177;
input n_540;
input n_593;
input n_514;
input n_646;
input n_528;
input n_391;
input n_457;
input n_687;
input n_697;
input n_364;
input n_637;
input n_295;
input n_385;
input n_629;
input n_388;
input n_190;
input n_262;
input n_484;
input n_613;
input n_187;
input n_501;
input n_531;
input n_60;
input n_361;
input n_508;
input n_663;
input n_379;
input n_170;
input n_332;
input n_336;
input n_12;
input n_398;
input n_410;
input n_566;
input n_554;
input n_602;
input n_194;
input n_664;
input n_171;
input n_678;
input n_192;
input n_57;
input n_169;
input n_51;
input n_649;
input n_283;

output n_5237;

wire n_2542;
wire n_1671;
wire n_2817;
wire n_801;
wire n_4452;
wire n_2576;
wire n_5172;
wire n_4649;
wire n_1674;
wire n_741;
wire n_1351;
wire n_1212;
wire n_4251;
wire n_2157;
wire n_5019;
wire n_2332;
wire n_3849;
wire n_5138;
wire n_4388;
wire n_4395;
wire n_1061;
wire n_3089;
wire n_783;
wire n_4978;
wire n_1854;
wire n_3088;
wire n_3257;
wire n_1342;
wire n_4829;
wire n_1387;
wire n_3222;
wire n_4699;
wire n_1151;
wire n_4686;
wire n_2317;
wire n_1975;
wire n_1930;
wire n_3706;
wire n_2179;
wire n_5055;
wire n_1547;
wire n_3376;
wire n_4868;
wire n_893;
wire n_3801;
wire n_4249;
wire n_1192;
wire n_3564;
wire n_1844;
wire n_1555;
wire n_5057;
wire n_3030;
wire n_830;
wire n_2838;
wire n_5229;
wire n_3427;
wire n_852;
wire n_5101;
wire n_2628;
wire n_3071;
wire n_2926;
wire n_1078;
wire n_4273;
wire n_2321;
wire n_2019;
wire n_5102;
wire n_3345;
wire n_2074;
wire n_2919;
wire n_4501;
wire n_2129;
wire n_4724;
wire n_945;
wire n_4997;
wire n_2399;
wire n_4843;
wire n_1232;
wire n_4696;
wire n_4347;
wire n_2480;
wire n_3877;
wire n_3929;
wire n_3048;
wire n_1455;
wire n_2786;
wire n_1781;
wire n_1971;
wire n_2004;
wire n_1106;
wire n_4814;
wire n_953;
wire n_3979;
wire n_3077;
wire n_2873;
wire n_3452;
wire n_3107;
wire n_4956;
wire n_1421;
wire n_3664;
wire n_1936;
wire n_5129;
wire n_1660;
wire n_5070;
wire n_3047;
wire n_4414;
wire n_713;
wire n_1400;
wire n_2625;
wire n_4646;
wire n_2843;
wire n_3760;
wire n_1560;
wire n_4262;
wire n_734;
wire n_1088;
wire n_1894;
wire n_3347;
wire n_5136;
wire n_907;
wire n_4110;
wire n_1658;
wire n_4950;
wire n_4729;
wire n_4268;
wire n_1967;
wire n_3999;
wire n_3928;
wire n_2613;
wire n_3535;
wire n_4751;
wire n_2708;
wire n_1648;
wire n_5151;
wire n_1911;
wire n_2011;
wire n_4102;
wire n_1641;
wire n_3871;
wire n_2735;
wire n_4662;
wire n_4671;
wire n_3959;
wire n_2268;
wire n_1367;
wire n_1336;
wire n_4314;
wire n_2080;
wire n_5099;
wire n_1381;
wire n_1699;
wire n_2093;
wire n_4296;
wire n_2770;
wire n_2101;
wire n_4507;
wire n_3484;
wire n_4677;
wire n_792;
wire n_5063;
wire n_1328;
wire n_2917;
wire n_2616;
wire n_3923;
wire n_3900;
wire n_3488;
wire n_939;
wire n_2811;
wire n_3732;
wire n_2832;
wire n_4226;
wire n_1762;
wire n_1910;
wire n_1075;
wire n_3980;
wire n_2998;
wire n_4366;
wire n_3446;
wire n_1895;
wire n_4294;
wire n_4698;
wire n_4445;
wire n_4810;
wire n_3859;
wire n_2692;
wire n_3914;
wire n_4456;
wire n_3397;
wire n_3575;
wire n_2469;
wire n_3927;
wire n_3888;
wire n_764;
wire n_2764;
wire n_2895;
wire n_733;
wire n_2922;
wire n_3882;
wire n_4856;
wire n_3492;
wire n_4369;
wire n_2068;
wire n_4331;
wire n_4972;
wire n_1290;
wire n_4993;
wire n_2072;
wire n_1354;
wire n_4375;
wire n_1701;
wire n_2678;
wire n_3935;
wire n_5130;
wire n_4291;
wire n_1726;
wire n_4613;
wire n_2434;
wire n_2878;
wire n_3012;
wire n_3875;
wire n_1167;
wire n_2428;
wire n_4717;
wire n_4877;
wire n_3247;
wire n_871;
wire n_2641;
wire n_4731;
wire n_3052;
wire n_5046;
wire n_2749;
wire n_3298;
wire n_2254;
wire n_5058;
wire n_1926;
wire n_3273;
wire n_4467;
wire n_1747;
wire n_780;
wire n_2624;
wire n_2350;
wire n_5042;
wire n_4681;
wire n_4072;
wire n_4752;
wire n_4220;
wire n_835;
wire n_928;
wire n_2092;
wire n_1654;
wire n_1750;
wire n_1462;
wire n_2514;
wire n_1588;
wire n_3942;
wire n_3997;
wire n_2468;
wire n_4381;
wire n_5144;
wire n_2096;
wire n_3968;
wire n_4466;
wire n_4418;
wire n_3434;
wire n_4510;
wire n_4473;
wire n_5226;
wire n_890;
wire n_2812;
wire n_4518;
wire n_1709;
wire n_2393;
wire n_2657;
wire n_2921;
wire n_2136;
wire n_2409;
wire n_2252;
wire n_3237;
wire n_949;
wire n_3500;
wire n_3834;
wire n_4589;
wire n_2075;
wire n_2972;
wire n_3542;
wire n_2763;
wire n_2762;
wire n_3192;
wire n_760;
wire n_1546;
wire n_4394;
wire n_2279;
wire n_1296;
wire n_3352;
wire n_3073;
wire n_2150;
wire n_1294;
wire n_3696;
wire n_1420;
wire n_4082;
wire n_1779;
wire n_4921;
wire n_1858;
wire n_4329;
wire n_5135;
wire n_3021;
wire n_2558;
wire n_1164;
wire n_4697;
wire n_4288;
wire n_4289;
wire n_3763;
wire n_2712;
wire n_3733;
wire n_1487;
wire n_3614;
wire n_874;
wire n_5183;
wire n_2145;
wire n_898;
wire n_4964;
wire n_4228;
wire n_3423;
wire n_925;
wire n_1932;
wire n_1101;
wire n_4636;
wire n_4322;
wire n_3644;
wire n_1249;
wire n_4946;
wire n_2706;
wire n_4767;
wire n_4287;
wire n_2693;
wire n_4137;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_963;
wire n_2767;
wire n_4576;
wire n_4615;
wire n_1139;
wire n_3179;
wire n_1018;
wire n_3400;
wire n_1521;
wire n_1366;
wire n_4000;
wire n_2897;
wire n_4389;
wire n_3970;
wire n_4345;
wire n_996;
wire n_1376;
wire n_4664;
wire n_2170;
wire n_4156;
wire n_948;
wire n_977;
wire n_3158;
wire n_1788;
wire n_4873;
wire n_2643;
wire n_3782;
wire n_1835;
wire n_3470;
wire n_5076;
wire n_4713;
wire n_4098;
wire n_5026;
wire n_4476;
wire n_3700;
wire n_4995;
wire n_3166;
wire n_3104;
wire n_3435;
wire n_842;
wire n_2239;
wire n_4310;
wire n_1432;
wire n_5212;
wire n_989;
wire n_2689;
wire n_1473;
wire n_2191;
wire n_1246;
wire n_4528;
wire n_899;
wire n_1035;
wire n_4914;
wire n_4939;
wire n_1426;
wire n_3418;
wire n_705;
wire n_1004;
wire n_1529;
wire n_2473;
wire n_4634;
wire n_2069;
wire n_2362;
wire n_4096;
wire n_2539;
wire n_2698;
wire n_4123;
wire n_3119;
wire n_3735;
wire n_2297;
wire n_4379;
wire n_4718;
wire n_1448;
wire n_3631;
wire n_2445;
wire n_2057;
wire n_2103;
wire n_3770;
wire n_2772;
wire n_4440;
wire n_4402;
wire n_927;
wire n_5052;
wire n_4541;
wire n_5009;
wire n_4872;
wire n_929;
wire n_4551;
wire n_2857;
wire n_1183;
wire n_4627;
wire n_4079;
wire n_2494;
wire n_3342;
wire n_998;
wire n_5035;
wire n_717;
wire n_1383;
wire n_3390;
wire n_3656;
wire n_1424;
wire n_1000;
wire n_3025;
wire n_2137;
wire n_1626;
wire n_1507;
wire n_2482;
wire n_3810;
wire n_4798;
wire n_2532;
wire n_1388;
wire n_3006;
wire n_912;
wire n_5010;
wire n_2296;
wire n_3633;
wire n_5089;
wire n_2849;
wire n_1201;
wire n_1398;
wire n_884;
wire n_4592;
wire n_1395;
wire n_2199;
wire n_2661;
wire n_731;
wire n_1955;
wire n_931;
wire n_1791;
wire n_958;
wire n_5137;
wire n_3331;
wire n_5104;
wire n_1897;
wire n_2064;
wire n_2773;
wire n_3606;
wire n_1310;
wire n_819;
wire n_1334;
wire n_3591;
wire n_2788;
wire n_964;
wire n_4756;
wire n_2797;
wire n_4746;
wire n_3892;
wire n_4970;
wire n_4069;
wire n_2748;
wire n_5194;
wire n_1834;
wire n_2331;
wire n_2292;
wire n_3441;
wire n_3534;
wire n_3964;
wire n_2416;
wire n_1877;
wire n_3944;
wire n_1939;
wire n_2030;
wire n_1769;
wire n_2209;
wire n_3605;
wire n_1602;
wire n_4633;
wire n_3306;
wire n_3026;
wire n_4584;
wire n_3090;
wire n_5232;
wire n_3724;
wire n_4276;
wire n_5116;
wire n_2990;
wire n_3847;
wire n_1773;
wire n_5001;
wire n_2552;
wire n_1053;
wire n_5176;
wire n_4428;
wire n_1533;
wire n_3323;
wire n_2274;
wire n_4618;
wire n_4679;
wire n_1745;
wire n_914;
wire n_3479;
wire n_4496;
wire n_4805;
wire n_1679;
wire n_3454;
wire n_2160;
wire n_2146;
wire n_2131;
wire n_3547;
wire n_2575;
wire n_5100;
wire n_4410;
wire n_1933;
wire n_1179;
wire n_3816;
wire n_4807;
wire n_4411;
wire n_3214;
wire n_1243;
wire n_2928;
wire n_5166;
wire n_1917;
wire n_1580;
wire n_2822;
wire n_4180;
wire n_1281;
wire n_3109;
wire n_3354;
wire n_2572;
wire n_1520;
wire n_3126;
wire n_3663;
wire n_2863;
wire n_1419;
wire n_3299;
wire n_1731;
wire n_2135;
wire n_4707;
wire n_1645;
wire n_1832;
wire n_4676;
wire n_5180;
wire n_858;
wire n_2049;
wire n_5182;
wire n_956;
wire n_4880;
wire n_3566;
wire n_2781;
wire n_4126;
wire n_2829;
wire n_1696;
wire n_3845;
wire n_1594;
wire n_1869;
wire n_3804;
wire n_4207;
wire n_5196;
wire n_2016;
wire n_5171;
wire n_4470;
wire n_4813;
wire n_1030;
wire n_3901;
wire n_1937;
wire n_1790;
wire n_4014;
wire n_4704;
wire n_1744;
wire n_828;
wire n_2142;
wire n_4252;
wire n_4028;
wire n_2448;
wire n_4048;
wire n_4596;
wire n_4444;
wire n_3756;
wire n_3406;
wire n_820;
wire n_951;
wire n_952;
wire n_3919;
wire n_2263;
wire n_5185;
wire n_974;
wire n_4952;
wire n_2656;
wire n_5023;
wire n_2375;
wire n_1934;
wire n_1434;
wire n_1573;
wire n_3981;
wire n_3973;
wire n_2756;
wire n_807;
wire n_4761;
wire n_1275;
wire n_2884;
wire n_1510;
wire n_3120;
wire n_3797;
wire n_2024;
wire n_1595;
wire n_4770;
wire n_1749;
wire n_3474;
wire n_2549;
wire n_4690;
wire n_1669;
wire n_1024;
wire n_3864;
wire n_4932;
wire n_2302;
wire n_1667;
wire n_1037;
wire n_5143;
wire n_3592;
wire n_4230;
wire n_2637;
wire n_1639;
wire n_3967;
wire n_3195;
wire n_2526;
wire n_4274;
wire n_5215;
wire n_3277;
wire n_2548;
wire n_991;
wire n_4189;
wire n_3817;
wire n_1108;
wire n_3659;
wire n_2559;
wire n_2177;
wire n_2595;
wire n_5003;
wire n_4827;
wire n_1601;
wire n_1960;
wire n_2694;
wire n_3648;
wire n_1686;
wire n_3042;
wire n_5094;
wire n_4610;
wire n_4472;
wire n_3228;
wire n_3657;
wire n_3081;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1586;
wire n_2264;
wire n_3464;
wire n_3723;
wire n_1190;
wire n_4380;
wire n_4990;
wire n_4996;
wire n_4398;
wire n_2498;
wire n_4515;
wire n_1891;
wire n_5031;
wire n_1213;
wire n_2235;
wire n_4193;
wire n_3570;
wire n_5082;
wire n_1673;
wire n_3828;
wire n_2392;
wire n_3424;
wire n_4131;
wire n_2298;
wire n_2326;
wire n_1539;
wire n_3594;
wire n_1043;
wire n_4090;
wire n_4165;
wire n_2305;
wire n_2120;
wire n_4626;
wire n_4144;
wire n_2964;
wire n_2169;
wire n_3485;
wire n_4077;
wire n_2371;
wire n_1361;
wire n_3262;
wire n_4008;
wire n_3356;
wire n_5221;
wire n_1642;
wire n_3210;
wire n_937;
wire n_4689;
wire n_1682;
wire n_4547;
wire n_3329;
wire n_3826;
wire n_4905;
wire n_1406;
wire n_4601;
wire n_962;
wire n_3647;
wire n_3681;
wire n_1883;
wire n_4300;
wire n_1288;
wire n_1186;
wire n_4623;
wire n_5007;
wire n_3320;
wire n_2518;
wire n_3988;
wire n_1720;
wire n_3476;
wire n_4842;
wire n_3439;
wire n_4135;
wire n_2688;
wire n_1845;
wire n_1489;
wire n_942;
wire n_2798;
wire n_2852;
wire n_1524;
wire n_1964;
wire n_1920;
wire n_2753;
wire n_1496;
wire n_3292;
wire n_2007;
wire n_2039;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_1846;
wire n_3437;
wire n_4111;
wire n_3712;
wire n_4608;
wire n_879;
wire n_2310;
wire n_2506;
wire n_4859;
wire n_2626;
wire n_1567;
wire n_4037;
wire n_3562;
wire n_2973;
wire n_5218;
wire n_3665;
wire n_3007;
wire n_3528;
wire n_4571;
wire n_3698;
wire n_3355;
wire n_2454;
wire n_2114;
wire n_3174;
wire n_1066;
wire n_1948;
wire n_4215;
wire n_2154;
wire n_1484;
wire n_4185;
wire n_3752;
wire n_2283;
wire n_5145;
wire n_4219;
wire n_1229;
wire n_1373;
wire n_3958;
wire n_3985;
wire n_2427;
wire n_4196;
wire n_1447;
wire n_4774;
wire n_2056;
wire n_5210;
wire n_4242;
wire n_5109;
wire n_3389;
wire n_4232;
wire n_4190;
wire n_4902;
wire n_3000;
wire n_5149;
wire n_2680;
wire n_1047;
wire n_3375;
wire n_3899;
wire n_1385;
wire n_3713;
wire n_1931;
wire n_2668;
wire n_1257;
wire n_3197;
wire n_4987;
wire n_2128;
wire n_4736;
wire n_2398;
wire n_1725;
wire n_3743;
wire n_834;
wire n_5033;
wire n_2695;
wire n_4035;
wire n_3818;
wire n_3124;
wire n_1741;
wire n_1002;
wire n_1949;
wire n_3759;
wire n_2671;
wire n_4516;
wire n_2715;
wire n_1804;
wire n_2508;
wire n_3511;
wire n_2054;
wire n_1337;
wire n_1477;
wire n_2614;
wire n_4492;
wire n_2833;
wire n_2758;
wire n_3694;
wire n_2937;
wire n_4789;
wire n_4376;
wire n_1001;
wire n_2241;
wire n_4708;
wire n_4657;
wire n_1690;
wire n_1191;
wire n_1076;
wire n_4512;
wire n_1378;
wire n_855;
wire n_1377;
wire n_4081;
wire n_1542;
wire n_4542;
wire n_4462;
wire n_1716;
wire n_4931;
wire n_4536;
wire n_3303;
wire n_978;
wire n_4324;
wire n_1976;
wire n_4382;
wire n_2905;
wire n_1291;
wire n_749;
wire n_1824;
wire n_3954;
wire n_2122;
wire n_2140;
wire n_3503;
wire n_3160;
wire n_1065;
wire n_1255;
wire n_5124;
wire n_3951;
wire n_823;
wire n_1074;
wire n_3569;
wire n_739;
wire n_3874;
wire n_2528;
wire n_5123;
wire n_4639;
wire n_1338;
wire n_1097;
wire n_3027;
wire n_781;
wire n_4083;
wire n_1810;
wire n_1583;
wire n_4480;
wire n_1730;
wire n_2295;
wire n_2746;
wire n_814;
wire n_1643;
wire n_2020;
wire n_4171;
wire n_3652;
wire n_4023;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_3617;
wire n_2076;
wire n_3567;
wire n_1598;
wire n_4344;
wire n_2935;
wire n_4705;
wire n_4046;
wire n_3807;
wire n_918;
wire n_1114;
wire n_763;
wire n_4027;
wire n_3154;
wire n_1227;
wire n_2485;
wire n_3898;
wire n_3520;
wire n_4391;
wire n_946;
wire n_1303;
wire n_4095;
wire n_2881;
wire n_1116;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_3551;
wire n_4947;
wire n_3064;
wire n_1780;
wire n_3897;
wire n_1689;
wire n_3372;
wire n_1944;
wire n_1347;
wire n_795;
wire n_1221;
wire n_1245;
wire n_3215;
wire n_3853;
wire n_4740;
wire n_4631;
wire n_1561;
wire n_1112;
wire n_2081;
wire n_2168;
wire n_5068;
wire n_1460;
wire n_911;
wire n_5159;
wire n_2862;
wire n_2615;
wire n_4068;
wire n_4625;
wire n_2474;
wire n_3703;
wire n_2437;
wire n_2444;
wire n_3962;
wire n_2743;
wire n_4766;
wire n_4863;
wire n_2267;
wire n_3035;
wire n_4166;
wire n_1821;
wire n_1058;
wire n_3378;
wire n_3745;
wire n_3362;
wire n_4744;
wire n_4188;
wire n_2934;
wire n_3667;
wire n_3523;
wire n_2222;
wire n_712;
wire n_3176;
wire n_2505;
wire n_4817;
wire n_4115;
wire n_2999;
wire n_2014;
wire n_1239;
wire n_3697;
wire n_1584;
wire n_3680;
wire n_2408;
wire n_3468;
wire n_5045;
wire n_1972;
wire n_4383;
wire n_4491;
wire n_4486;
wire n_1816;
wire n_3024;
wire n_4612;
wire n_2531;
wire n_5163;
wire n_4529;
wire n_3361;
wire n_714;
wire n_3478;
wire n_3936;
wire n_1349;
wire n_2723;
wire n_2800;
wire n_3496;
wire n_4390;
wire n_3096;
wire n_2651;
wire n_2095;
wire n_3239;
wire n_3161;
wire n_2799;
wire n_3902;
wire n_4062;
wire n_3295;
wire n_4396;
wire n_1998;
wire n_1574;
wire n_3101;
wire n_756;
wire n_1981;
wire n_4233;
wire n_1606;
wire n_3374;
wire n_2640;
wire n_1552;
wire n_2918;
wire n_3288;
wire n_4307;
wire n_3992;
wire n_3876;
wire n_3125;
wire n_4293;
wire n_941;
wire n_3552;
wire n_1031;
wire n_849;
wire n_4684;
wire n_3116;
wire n_4091;
wire n_1753;
wire n_5027;
wire n_3095;
wire n_2471;
wire n_4412;
wire n_2807;
wire n_1921;
wire n_3618;
wire n_4580;
wire n_1055;
wire n_2217;
wire n_2197;
wire n_4758;
wire n_4781;
wire n_4148;
wire n_2461;
wire n_4057;
wire n_1170;
wire n_3444;
wire n_1040;
wire n_3059;
wire n_2634;
wire n_1761;
wire n_1890;
wire n_3017;
wire n_1805;
wire n_2477;
wire n_2308;
wire n_2333;
wire n_3001;
wire n_1089;
wire n_3795;
wire n_3852;
wire n_1365;
wire n_4138;
wire n_5018;
wire n_3815;
wire n_3896;
wire n_3274;
wire n_4457;
wire n_4093;
wire n_1616;
wire n_1862;
wire n_4928;
wire n_4794;
wire n_722;
wire n_2223;
wire n_4197;
wire n_4482;
wire n_1621;
wire n_2547;
wire n_2415;
wire n_5073;
wire n_827;
wire n_4834;
wire n_4762;
wire n_3113;
wire n_992;
wire n_3813;
wire n_3660;
wire n_3766;
wire n_1613;
wire n_1458;
wire n_1027;
wire n_3266;
wire n_3574;
wire n_1189;
wire n_4154;
wire n_4907;
wire n_5077;
wire n_5034;
wire n_726;
wire n_4504;
wire n_3844;
wire n_1237;
wire n_2534;
wire n_4975;
wire n_3741;
wire n_2451;
wire n_2243;
wire n_4815;
wire n_4898;
wire n_3443;
wire n_4819;
wire n_1209;
wire n_1708;
wire n_805;
wire n_2051;
wire n_4370;
wire n_2359;
wire n_5112;
wire n_1402;
wire n_1691;
wire n_3332;
wire n_4134;
wire n_1238;
wire n_2570;
wire n_4092;
wire n_4645;
wire n_3668;
wire n_2491;
wire n_1264;
wire n_4755;
wire n_4359;
wire n_4960;
wire n_4087;
wire n_1700;
wire n_4933;
wire n_5091;
wire n_3487;
wire n_4591;
wire n_4302;
wire n_5111;
wire n_3340;
wire n_5227;
wire n_873;
wire n_3946;
wire n_2989;
wire n_3395;
wire n_4474;
wire n_2509;
wire n_2513;
wire n_3757;
wire n_4178;
wire n_5165;
wire n_1704;
wire n_2247;
wire n_1711;
wire n_4884;
wire n_1579;
wire n_3275;
wire n_836;
wire n_3678;
wire n_3440;
wire n_2094;
wire n_1511;
wire n_2356;
wire n_1422;
wire n_1772;
wire n_4692;
wire n_3165;
wire n_1119;
wire n_1433;
wire n_1902;
wire n_1842;
wire n_1620;
wire n_2739;
wire n_1735;
wire n_3890;
wire n_1541;
wire n_1300;
wire n_3750;
wire n_1313;
wire n_3607;
wire n_3316;
wire n_2418;
wire n_2864;
wire n_4311;
wire n_1180;
wire n_2703;
wire n_3371;
wire n_4722;
wire n_4606;
wire n_3261;
wire n_4187;
wire n_940;
wire n_2058;
wire n_2660;
wire n_1094;
wire n_4962;
wire n_4563;
wire n_5056;
wire n_4820;
wire n_2394;
wire n_3532;
wire n_3948;
wire n_2124;
wire n_4619;
wire n_4327;
wire n_1961;
wire n_5211;
wire n_3765;
wire n_4125;
wire n_5036;
wire n_4221;
wire n_3297;
wire n_976;
wire n_3067;
wire n_2155;
wire n_2686;
wire n_2364;
wire n_4392;
wire n_2996;
wire n_3803;
wire n_2085;
wire n_917;
wire n_5014;
wire n_3639;
wire n_5192;
wire n_4334;
wire n_3351;
wire n_808;
wire n_4047;
wire n_3413;
wire n_1193;
wire n_5233;
wire n_3412;
wire n_3791;
wire n_3164;
wire n_4575;
wire n_699;
wire n_4320;
wire n_3884;
wire n_5139;
wire n_757;
wire n_5231;
wire n_2190;
wire n_3438;
wire n_4141;
wire n_5193;
wire n_2850;
wire n_1481;
wire n_1441;
wire n_3373;
wire n_2104;
wire n_3883;
wire n_3728;
wire n_2925;
wire n_4499;
wire n_5195;
wire n_3949;
wire n_2792;
wire n_3315;
wire n_3798;
wire n_788;
wire n_1543;
wire n_1599;
wire n_4257;
wire n_4458;
wire n_2674;
wire n_5103;
wire n_4641;
wire n_4720;
wire n_4893;
wire n_3857;
wire n_1876;
wire n_4107;
wire n_1873;
wire n_3630;
wire n_3518;
wire n_1866;
wire n_2130;
wire n_1413;
wire n_1330;
wire n_3714;
wire n_2228;
wire n_5039;
wire n_2455;
wire n_2876;
wire n_4772;
wire n_3099;
wire n_5198;
wire n_4468;
wire n_4161;
wire n_1663;
wire n_4172;
wire n_3403;
wire n_2714;
wire n_2245;
wire n_4961;
wire n_4454;
wire n_1107;
wire n_2457;
wire n_3294;
wire n_4119;
wire n_3686;
wire n_4502;
wire n_2971;
wire n_1713;
wire n_715;
wire n_4277;
wire n_4526;
wire n_1265;
wire n_3490;
wire n_4849;
wire n_4319;
wire n_3369;
wire n_3581;
wire n_3069;
wire n_2028;
wire n_3715;
wire n_1069;
wire n_3725;
wire n_3933;
wire n_1175;
wire n_2311;
wire n_1012;
wire n_3691;
wire n_4485;
wire n_4066;
wire n_903;
wire n_4146;
wire n_1802;
wire n_1504;
wire n_4340;
wire n_3961;
wire n_4855;
wire n_1801;
wire n_2347;
wire n_3917;
wire n_816;
wire n_1188;
wire n_2206;
wire n_4004;
wire n_2967;
wire n_2916;
wire n_4292;
wire n_2467;
wire n_3145;
wire n_1124;
wire n_1624;
wire n_3983;
wire n_4940;
wire n_3538;
wire n_3280;
wire n_1515;
wire n_961;
wire n_4356;
wire n_3510;
wire n_2824;
wire n_2377;
wire n_701;
wire n_950;
wire n_3009;
wire n_3719;
wire n_2525;
wire n_4361;
wire n_3827;
wire n_891;
wire n_5154;
wire n_2067;
wire n_3889;
wire n_2687;
wire n_1630;
wire n_2887;
wire n_4245;
wire n_4136;
wire n_3526;
wire n_2194;
wire n_2619;
wire n_4367;
wire n_1987;
wire n_968;
wire n_2271;
wire n_1008;
wire n_2583;
wire n_4560;
wire n_2606;
wire n_4899;
wire n_1033;
wire n_1052;
wire n_2794;
wire n_5164;
wire n_2391;
wire n_2431;
wire n_2078;
wire n_2932;
wire n_1767;
wire n_3431;
wire n_3450;
wire n_4663;
wire n_2893;
wire n_1208;
wire n_2954;
wire n_2728;
wire n_1072;
wire n_815;
wire n_3421;
wire n_3183;
wire n_2493;
wire n_4802;
wire n_2705;
wire n_1067;
wire n_3405;
wire n_1952;
wire n_5074;
wire n_4044;
wire n_3436;
wire n_1026;
wire n_1880;
wire n_3442;
wire n_3366;
wire n_2631;
wire n_3937;
wire n_1293;
wire n_3159;
wire n_4701;
wire n_794;
wire n_727;
wire n_894;
wire n_3240;
wire n_3576;
wire n_1863;
wire n_3385;
wire n_4851;
wire n_3293;
wire n_872;
wire n_3922;
wire n_5204;
wire n_847;
wire n_851;
wire n_4991;
wire n_2554;
wire n_1513;
wire n_1913;
wire n_4934;
wire n_837;
wire n_5087;
wire n_2517;
wire n_2713;
wire n_5000;
wire n_2765;
wire n_2590;
wire n_3150;
wire n_2060;
wire n_4479;
wire n_2608;
wire n_4011;
wire n_5131;
wire n_1959;
wire n_3133;
wire n_765;
wire n_1492;
wire n_1340;
wire n_4688;
wire n_4753;
wire n_4058;
wire n_2262;
wire n_3611;
wire n_3082;
wire n_4848;
wire n_5059;
wire n_843;
wire n_2604;
wire n_2407;
wire n_1277;
wire n_2816;
wire n_3799;
wire n_2574;
wire n_4475;
wire n_5219;
wire n_2675;
wire n_3537;
wire n_4443;
wire n_3887;
wire n_1022;
wire n_2667;
wire n_4587;
wire n_1615;
wire n_4114;
wire n_1474;
wire n_1571;
wire n_2948;
wire n_1577;
wire n_2119;
wire n_947;
wire n_1117;
wire n_1992;
wire n_3223;
wire n_3140;
wire n_3185;
wire n_4749;
wire n_2605;
wire n_5155;
wire n_926;
wire n_3654;
wire n_1849;
wire n_2848;
wire n_919;
wire n_1698;
wire n_4100;
wire n_4264;
wire n_3788;
wire n_4891;
wire n_777;
wire n_1299;
wire n_3837;
wire n_2718;
wire n_1436;
wire n_1384;
wire n_3325;
wire n_2238;
wire n_4085;
wire n_4464;
wire n_4624;
wire n_4818;
wire n_4659;
wire n_3600;
wire n_5217;
wire n_5015;
wire n_4339;
wire n_1178;
wire n_2338;
wire n_3324;
wire n_796;
wire n_1195;
wire n_1811;
wire n_1857;
wire n_3987;
wire n_1519;
wire n_2144;
wire n_1284;
wire n_1604;
wire n_4487;
wire n_4889;
wire n_4866;
wire n_1142;
wire n_1048;
wire n_3638;
wire n_4816;
wire n_2110;
wire n_1502;
wire n_1659;
wire n_3393;
wire n_3451;
wire n_1418;
wire n_1250;
wire n_4937;
wire n_3615;
wire n_3072;
wire n_3087;
wire n_2053;
wire n_2259;
wire n_2121;
wire n_4222;
wire n_4874;
wire n_4401;
wire n_889;
wire n_2710;
wire n_3142;
wire n_4015;
wire n_1966;
wire n_1110;
wire n_4709;
wire n_2213;
wire n_4976;
wire n_2389;
wire n_2132;
wire n_2892;
wire n_4120;
wire n_1564;
wire n_4658;
wire n_2860;
wire n_2330;
wire n_1457;
wire n_3718;
wire n_1787;
wire n_1993;
wire n_2281;
wire n_2617;
wire n_2776;
wire n_1466;
wire n_1919;
wire n_5207;
wire n_3705;
wire n_3211;
wire n_3909;
wire n_1220;
wire n_1893;
wire n_2301;
wire n_4665;
wire n_3582;
wire n_4223;
wire n_2387;
wire n_3270;
wire n_2846;
wire n_970;
wire n_2488;
wire n_1980;
wire n_2237;
wire n_1060;
wire n_1951;
wire n_4362;
wire n_1252;
wire n_3311;
wire n_3913;
wire n_1223;
wire n_5121;
wire n_1286;
wire n_2115;
wire n_4430;
wire n_3302;
wire n_4348;
wire n_5013;
wire n_1597;
wire n_4489;
wire n_4839;
wire n_2596;
wire n_3163;
wire n_775;
wire n_4404;
wire n_1153;
wire n_1531;
wire n_2828;
wire n_2384;
wire n_4261;
wire n_4204;
wire n_759;
wire n_2724;
wire n_2585;
wire n_4825;
wire n_2352;
wire n_1625;
wire n_3986;
wire n_5006;
wire n_4513;
wire n_4006;
wire n_2226;
wire n_2801;
wire n_1901;
wire n_3869;
wire n_2556;
wire n_4747;
wire n_1647;
wire n_3753;
wire n_2306;
wire n_1614;
wire n_1892;
wire n_3742;
wire n_3683;
wire n_4801;
wire n_3260;
wire n_2550;
wire n_3175;
wire n_3736;
wire n_4448;
wire n_1096;
wire n_2227;
wire n_5216;
wire n_3284;
wire n_4869;
wire n_2159;
wire n_4386;
wire n_1077;
wire n_2315;
wire n_4132;
wire n_2995;
wire n_1437;
wire n_4438;
wire n_4844;
wire n_4836;
wire n_4955;
wire n_4149;
wire n_4355;
wire n_3234;
wire n_2276;
wire n_856;
wire n_2803;
wire n_1668;
wire n_2777;
wire n_3202;
wire n_2830;
wire n_3220;
wire n_1129;
wire n_2181;
wire n_2911;
wire n_4655;
wire n_1429;
wire n_2826;
wire n_3429;
wire n_2379;
wire n_3554;
wire n_1593;
wire n_1202;
wire n_1635;
wire n_4067;
wire n_4357;
wire n_3462;
wire n_2851;
wire n_4374;
wire n_5132;
wire n_2420;
wire n_3722;
wire n_4400;
wire n_4846;
wire n_2984;
wire n_5187;
wire n_4024;
wire n_1508;
wire n_732;
wire n_2983;
wire n_2240;
wire n_2538;
wire n_724;
wire n_3250;
wire n_1042;
wire n_4582;
wire n_1728;
wire n_1871;
wire n_4860;
wire n_845;
wire n_3414;
wire n_1549;
wire n_4870;
wire n_768;
wire n_3651;
wire n_2102;
wire n_2563;
wire n_4989;
wire n_3449;
wire n_1683;
wire n_1916;
wire n_2598;
wire n_1187;
wire n_4304;
wire n_4558;
wire n_1403;
wire n_4488;
wire n_3767;
wire n_2544;
wire n_3550;
wire n_4211;
wire n_1206;
wire n_4016;
wire n_750;
wire n_4656;
wire n_3839;
wire n_2823;
wire n_4915;
wire n_4328;
wire n_1057;
wire n_2785;
wire n_1997;
wire n_2636;
wire n_3131;
wire n_710;
wire n_1818;
wire n_3730;
wire n_1298;
wire n_4397;
wire n_3399;
wire n_2088;
wire n_1611;
wire n_5050;
wire n_2740;
wire n_746;
wire n_4808;
wire n_3416;
wire n_3498;
wire n_2401;
wire n_1589;
wire n_4712;
wire n_2309;
wire n_2900;
wire n_2957;
wire n_1740;
wire n_2737;
wire n_3994;
wire n_1497;
wire n_3672;
wire n_3533;
wire n_1622;
wire n_4725;
wire n_4406;
wire n_1694;
wire n_1535;
wire n_3382;
wire n_3132;
wire n_2571;
wire n_3138;
wire n_5053;
wire n_2171;
wire n_2988;
wire n_4908;
wire n_3136;
wire n_1350;
wire n_4192;
wire n_4109;
wire n_4824;
wire n_2037;
wire n_2808;
wire n_4567;
wire n_5150;
wire n_782;
wire n_809;
wire n_3819;
wire n_4778;
wire n_1797;
wire n_5175;
wire n_986;
wire n_2050;
wire n_4595;
wire n_2164;
wire n_4174;
wire n_1870;
wire n_1171;
wire n_5179;
wire n_1827;
wire n_4904;
wire n_2187;
wire n_1152;
wire n_3544;
wire n_4150;
wire n_2904;
wire n_711;
wire n_3105;
wire n_2872;
wire n_3692;
wire n_4616;
wire n_4982;
wire n_1695;
wire n_2046;
wire n_2272;
wire n_2760;
wire n_1979;
wire n_4643;
wire n_2738;
wire n_972;
wire n_1332;
wire n_4323;
wire n_2346;
wire n_4831;
wire n_936;
wire n_3045;
wire n_3821;
wire n_885;
wire n_2342;
wire n_2167;
wire n_2970;
wire n_3676;
wire n_4896;
wire n_2882;
wire n_3666;
wire n_3675;
wire n_4017;
wire n_4260;
wire n_4916;
wire n_2541;
wire n_2940;
wire n_4739;
wire n_1974;
wire n_4122;
wire n_934;
wire n_4209;
wire n_2768;
wire n_3858;
wire n_1341;
wire n_4298;
wire n_2314;
wire n_3502;
wire n_3003;
wire n_4128;
wire n_5147;
wire n_4271;
wire n_4644;
wire n_1355;
wire n_2258;
wire n_804;
wire n_2390;
wire n_959;
wire n_2562;
wire n_4716;
wire n_4312;
wire n_1343;
wire n_1522;
wire n_2734;
wire n_1782;
wire n_707;
wire n_1900;
wire n_5048;
wire n_3246;
wire n_1548;
wire n_3381;
wire n_1155;
wire n_2195;
wire n_3208;
wire n_4944;
wire n_4343;
wire n_4715;
wire n_4935;
wire n_4694;
wire n_4672;
wire n_5054;
wire n_2962;
wire n_2939;
wire n_1672;
wire n_1925;
wire n_4407;
wire n_737;
wire n_3517;
wire n_4045;
wire n_3893;
wire n_4598;
wire n_2945;
wire n_3061;
wire n_3932;
wire n_3469;
wire n_2960;
wire n_3258;
wire n_4524;
wire n_3143;
wire n_4084;
wire n_3149;
wire n_3365;
wire n_3379;
wire n_4850;
wire n_4424;
wire n_3008;
wire n_1751;
wire n_2840;
wire n_3939;
wire n_4776;
wire n_1375;
wire n_3972;
wire n_4153;
wire n_3506;
wire n_1650;
wire n_1962;
wire n_3855;
wire n_1928;
wire n_3091;
wire n_4317;
wire n_4723;
wire n_4269;
wire n_4088;
wire n_3398;
wire n_2761;
wire n_2793;
wire n_3776;
wire n_3711;
wire n_4235;
wire n_1019;
wire n_4143;
wire n_4170;
wire n_729;
wire n_876;
wire n_774;
wire n_3642;
wire n_2845;
wire n_4650;
wire n_4719;
wire n_5173;
wire n_1860;
wire n_5016;
wire n_1904;
wire n_2874;
wire n_1200;
wire n_2588;
wire n_1353;
wire n_1777;
wire n_4967;
wire n_3308;
wire n_1600;
wire n_1113;
wire n_2253;
wire n_2366;
wire n_4912;
wire n_4799;
wire n_2261;
wire n_4423;
wire n_5086;
wire n_2210;
wire n_4735;
wire n_3602;
wire n_3300;
wire n_2978;
wire n_2516;
wire n_1050;
wire n_1411;
wire n_5170;
wire n_2827;
wire n_1177;
wire n_3515;
wire n_1150;
wire n_1023;
wire n_2951;
wire n_1118;
wire n_2949;
wire n_1807;
wire n_5028;
wire n_1814;
wire n_1631;
wire n_1879;
wire n_3806;
wire n_2931;
wire n_2569;
wire n_3866;
wire n_4543;
wire n_740;
wire n_703;
wire n_4157;
wire n_4229;
wire n_3865;
wire n_4073;
wire n_1324;
wire n_3629;
wire n_1435;
wire n_3920;
wire n_969;
wire n_4892;
wire n_3255;
wire n_1401;
wire n_1516;
wire n_3846;
wire n_3512;
wire n_5201;
wire n_2029;
wire n_4439;
wire n_1394;
wire n_1326;
wire n_4783;
wire n_1379;
wire n_935;
wire n_4910;
wire n_1130;
wire n_3083;
wire n_832;
wire n_3049;
wire n_5142;
wire n_3830;
wire n_3679;
wire n_3541;
wire n_3117;
wire n_4930;
wire n_1283;
wire n_2385;
wire n_4112;
wire n_2149;
wire n_2396;
wire n_4557;
wire n_4917;
wire n_895;
wire n_2450;
wire n_3739;
wire n_4432;
wire n_2284;
wire n_4352;
wire n_4416;
wire n_4593;
wire n_2769;
wire n_4465;
wire n_3622;
wire n_5114;
wire n_4980;
wire n_1392;
wire n_4495;
wire n_5117;
wire n_1924;
wire n_2463;
wire n_3363;
wire n_1677;
wire n_3721;
wire n_3062;
wire n_2679;
wire n_5024;
wire n_4559;
wire n_838;
wire n_3969;
wire n_3336;
wire n_4160;
wire n_4231;
wire n_2952;
wire n_1017;
wire n_4256;
wire n_2779;
wire n_4938;
wire n_5203;
wire n_930;
wire n_2620;
wire n_5162;
wire n_1945;
wire n_1656;
wire n_2112;
wire n_1464;
wire n_2430;
wire n_1414;
wire n_2721;
wire n_944;
wire n_4335;
wire n_2034;
wire n_2683;
wire n_2744;
wire n_1011;
wire n_4521;
wire n_1566;
wire n_990;
wire n_3204;
wire n_1104;
wire n_4920;
wire n_870;
wire n_1253;
wire n_1693;
wire n_3256;
wire n_3802;
wire n_2118;
wire n_2111;
wire n_2915;
wire n_1148;
wire n_2188;
wire n_1989;
wire n_2802;
wire n_3643;
wire n_2425;
wire n_4265;
wire n_2950;
wire n_719;
wire n_3060;
wire n_3098;
wire n_4105;
wire n_1851;
wire n_1090;
wire n_4861;
wire n_4064;
wire n_4926;
wire n_1518;
wire n_1362;
wire n_3123;
wire n_3380;
wire n_1829;
wire n_1450;
wire n_4828;
wire n_1638;
wire n_3038;
wire n_1789;
wire n_2523;
wire n_2413;
wire n_3769;
wire n_1482;
wire n_3863;
wire n_3669;
wire n_3130;
wire n_4316;
wire n_4640;
wire n_5122;
wire n_1710;
wire n_2161;
wire n_1301;
wire n_2805;
wire n_4769;
wire n_2282;
wire n_4628;
wire n_2047;
wire n_1609;
wire n_3344;
wire n_2334;
wire n_5133;
wire n_1763;
wire n_3989;
wire n_2490;
wire n_4460;
wire n_4108;
wire n_3786;
wire n_3841;
wire n_4254;
wire n_1996;
wire n_2867;
wire n_1442;
wire n_2726;
wire n_4303;
wire n_1158;
wire n_2248;
wire n_5011;
wire n_2662;
wire n_3147;
wire n_4909;
wire n_753;
wire n_3925;
wire n_3180;
wire n_2795;
wire n_3472;
wire n_5106;
wire n_1479;
wire n_4768;
wire n_1675;
wire n_3717;
wire n_2215;
wire n_1884;
wire n_2055;
wire n_5156;
wire n_2553;
wire n_2038;
wire n_4447;
wire n_4826;
wire n_3445;
wire n_1833;
wire n_3903;
wire n_1494;
wire n_2325;
wire n_1850;
wire n_3854;
wire n_3235;
wire n_1417;
wire n_3673;
wire n_4281;
wire n_4648;
wire n_3094;
wire n_965;
wire n_1428;
wire n_1576;
wire n_1856;
wire n_2077;
wire n_1059;
wire n_4951;
wire n_4957;
wire n_3079;
wire n_4360;
wire n_4039;
wire n_3070;
wire n_3800;
wire n_4566;
wire n_3263;
wire n_4853;
wire n_1748;
wire n_3504;
wire n_4272;
wire n_2930;
wire n_1025;
wire n_3111;
wire n_1885;
wire n_3054;
wire n_1538;
wire n_1240;
wire n_4730;
wire n_1234;
wire n_3254;
wire n_3684;
wire n_4670;
wire n_4882;
wire n_4620;
wire n_3152;
wire n_4738;
wire n_3579;
wire n_3335;
wire n_4177;
wire n_3783;
wire n_700;
wire n_1307;
wire n_3178;
wire n_4127;
wire n_5206;
wire n_1003;
wire n_2353;
wire n_4099;
wire n_4517;
wire n_4168;
wire n_5188;
wire n_1738;
wire n_4490;
wire n_1575;
wire n_1923;
wire n_2260;
wire n_3952;
wire n_3911;
wire n_1688;
wire n_4285;
wire n_3465;
wire n_1743;
wire n_2997;
wire n_1991;
wire n_2386;
wire n_5161;
wire n_1724;
wire n_3708;
wire n_4078;
wire n_3046;
wire n_2956;
wire n_1553;
wire n_3619;
wire n_1415;
wire n_1370;
wire n_1786;
wire n_4198;
wire n_2382;
wire n_3754;
wire n_2291;
wire n_1371;
wire n_2886;
wire n_2974;
wire n_4213;
wire n_2184;
wire n_2982;
wire n_1803;
wire n_4065;
wire n_2645;
wire n_3904;
wire n_1393;
wire n_1517;
wire n_1867;
wire n_2630;
wire n_1444;
wire n_1603;
wire n_2470;
wire n_4446;
wire n_1263;
wire n_4417;
wire n_4733;
wire n_4764;
wire n_1261;
wire n_3879;
wire n_2286;
wire n_4743;
wire n_2018;
wire n_3080;
wire n_1903;
wire n_1143;
wire n_1874;
wire n_2865;
wire n_2825;
wire n_2013;
wire n_2044;
wire n_3023;
wire n_3232;
wire n_1056;
wire n_758;
wire n_2256;
wire n_943;
wire n_4060;
wire n_5110;
wire n_4879;
wire n_772;
wire n_2806;
wire n_770;
wire n_3028;
wire n_3662;
wire n_2981;
wire n_3076;
wire n_886;
wire n_3624;
wire n_1345;
wire n_1820;
wire n_4556;
wire n_4117;
wire n_4687;
wire n_2836;
wire n_1404;
wire n_2378;
wire n_887;
wire n_2655;
wire n_4600;
wire n_1467;
wire n_4250;
wire n_3906;
wire n_4954;
wire n_5191;
wire n_1231;
wire n_2599;
wire n_3963;
wire n_3368;
wire n_2370;
wire n_2612;
wire n_2591;
wire n_4881;
wire n_1815;
wire n_2214;
wire n_4253;
wire n_913;
wire n_2593;
wire n_4255;
wire n_867;
wire n_4071;
wire n_3568;
wire n_1230;
wire n_3850;
wire n_1333;
wire n_2496;
wire n_3313;
wire n_4605;
wire n_3189;
wire n_1644;
wire n_2725;
wire n_2277;
wire n_4691;
wire n_1558;
wire n_1732;
wire n_2300;
wire n_3943;
wire n_4305;
wire n_824;
wire n_4297;
wire n_2907;
wire n_1843;
wire n_4227;
wire n_2778;
wire n_1909;
wire n_5020;
wire n_1123;
wire n_1309;
wire n_2961;
wire n_916;
wire n_3934;
wire n_4033;
wire n_4415;
wire n_1970;
wire n_2059;
wire n_2669;
wire n_4094;
wire n_4765;
wire n_2546;
wire n_3193;
wire n_2522;
wire n_4364;
wire n_1957;
wire n_4354;
wire n_4732;
wire n_3912;
wire n_3118;
wire n_3720;
wire n_1907;
wire n_2529;
wire n_860;
wire n_1530;
wire n_4745;
wire n_938;
wire n_1302;
wire n_4581;
wire n_4377;
wire n_2143;
wire n_905;
wire n_4792;
wire n_1680;
wire n_3842;
wire n_993;
wire n_2031;
wire n_4878;
wire n_1605;
wire n_3514;
wire n_4979;
wire n_1988;
wire n_2654;
wire n_3036;
wire n_966;
wire n_4511;
wire n_2908;
wire n_3357;
wire n_1233;
wire n_3895;
wire n_4520;
wire n_3455;
wire n_4118;
wire n_4503;
wire n_2176;
wire n_2459;
wire n_1111;
wire n_3599;
wire n_1251;
wire n_2711;
wire n_4199;
wire n_1912;
wire n_4441;
wire n_1982;
wire n_3872;
wire n_3772;
wire n_1312;
wire n_5038;
wire n_1760;
wire n_4585;
wire n_2664;
wire n_1664;
wire n_1722;
wire n_3022;
wire n_1165;
wire n_4773;
wire n_2008;
wire n_2192;
wire n_3281;
wire n_2345;
wire n_1386;
wire n_4427;
wire n_5113;
wire n_3549;
wire n_2804;
wire n_2453;
wire n_2676;
wire n_3940;
wire n_4822;
wire n_1214;
wire n_850;
wire n_4800;
wire n_1157;
wire n_3453;
wire n_3410;
wire n_1752;
wire n_1813;
wire n_3768;
wire n_4958;
wire n_2810;
wire n_4043;
wire n_2319;
wire n_825;
wire n_3785;
wire n_2963;
wire n_2602;
wire n_3873;
wire n_2980;
wire n_4886;
wire n_1317;
wire n_1082;
wire n_3227;
wire n_2733;
wire n_3289;
wire n_4055;
wire n_2178;
wire n_2644;
wire n_2036;
wire n_3326;
wire n_4200;
wire n_3460;
wire n_2411;
wire n_1796;
wire n_2082;
wire n_3519;
wire n_5078;
wire n_3707;
wire n_3578;
wire n_909;
wire n_4737;
wire n_4925;
wire n_4116;
wire n_1990;
wire n_3805;
wire n_2943;
wire n_5205;
wire n_1634;
wire n_3252;
wire n_3253;
wire n_1465;
wire n_2622;
wire n_2658;
wire n_2665;
wire n_2133;
wire n_1712;
wire n_4603;
wire n_1523;
wire n_1627;
wire n_5080;
wire n_3128;
wire n_1527;
wire n_2691;
wire n_840;
wire n_2913;
wire n_4471;
wire n_2230;
wire n_1969;
wire n_2690;
wire n_5208;
wire n_1565;
wire n_1493;
wire n_2573;
wire n_2646;
wire n_2535;
wire n_1364;
wire n_3078;
wire n_2436;
wire n_3838;
wire n_4651;
wire n_3941;
wire n_3793;
wire n_4854;
wire n_5071;
wire n_3789;
wire n_1514;
wire n_3037;
wire n_1646;
wire n_3729;
wire n_4994;
wire n_2537;
wire n_4483;
wire n_5168;
wire n_4661;
wire n_1308;
wire n_4988;
wire n_3171;
wire n_3608;
wire n_4540;
wire n_2097;
wire n_3459;
wire n_2853;
wire n_1808;
wire n_3053;
wire n_3358;
wire n_3499;
wire n_4284;
wire n_1005;
wire n_1947;
wire n_3426;
wire n_4971;
wire n_1469;
wire n_5125;
wire n_2650;
wire n_987;
wire n_720;
wire n_3229;
wire n_3348;
wire n_1707;
wire n_5228;
wire n_797;
wire n_2933;
wire n_2717;
wire n_1723;
wire n_1878;
wire n_738;
wire n_2012;
wire n_3497;
wire n_5066;
wire n_2842;
wire n_3580;
wire n_2335;
wire n_2307;
wire n_3704;
wire n_1809;
wire n_4280;
wire n_1181;
wire n_5190;
wire n_3173;
wire n_3677;
wire n_3996;
wire n_1049;
wire n_4097;
wire n_1666;
wire n_803;
wire n_4218;
wire n_1717;
wire n_1817;
wire n_2449;
wire n_3880;
wire n_3685;
wire n_2868;
wire n_2231;
wire n_3609;
wire n_1228;
wire n_4459;
wire n_4545;
wire n_2896;
wire n_3019;
wire n_2639;
wire n_3471;
wire n_2898;
wire n_2368;
wire n_4175;
wire n_3200;
wire n_4771;
wire n_3259;
wire n_2524;
wire n_3167;
wire n_2460;
wire n_3867;
wire n_3593;
wire n_4455;
wire n_1073;
wire n_4514;
wire n_3191;
wire n_4140;
wire n_2481;
wire n_3561;
wire n_4806;
wire n_2682;
wire n_3032;
wire n_5160;
wire n_2877;
wire n_5098;
wire n_1021;
wire n_811;
wire n_1207;
wire n_5140;
wire n_4992;
wire n_5197;
wire n_880;
wire n_3505;
wire n_3577;
wire n_3540;
wire n_2432;
wire n_1478;
wire n_4796;
wire n_3598;
wire n_4442;
wire n_2581;
wire n_1363;
wire n_3641;
wire n_3777;
wire n_4203;
wire n_767;
wire n_1837;
wire n_2218;
wire n_4533;
wire n_831;
wire n_3590;
wire n_2435;
wire n_954;
wire n_4419;
wire n_1410;
wire n_5184;
wire n_1382;
wire n_1736;
wire n_4053;
wire n_1483;
wire n_3848;
wire n_1372;
wire n_3327;
wire n_1719;
wire n_2701;
wire n_2511;
wire n_4167;
wire n_1427;
wire n_2745;
wire n_1080;
wire n_2323;
wire n_2784;
wire n_5234;
wire n_4431;
wire n_2421;
wire n_1136;
wire n_4387;
wire n_2618;
wire n_3265;
wire n_2464;
wire n_1125;
wire n_3755;
wire n_4042;
wire n_5128;
wire n_2224;
wire n_2329;
wire n_1092;
wire n_4299;
wire n_4890;
wire n_1784;
wire n_3571;
wire n_1775;
wire n_2410;
wire n_1093;
wire n_1783;
wire n_2929;
wire n_4176;
wire n_5199;
wire n_3407;
wire n_1185;
wire n_3856;
wire n_4236;
wire n_3425;
wire n_3894;
wire n_3127;
wire n_1831;
wire n_2621;
wire n_3623;
wire n_5079;
wire n_1453;
wire n_2502;
wire n_3646;
wire n_4830;
wire n_4706;
wire n_1315;
wire n_5225;
wire n_4570;
wire n_2754;
wire n_1224;
wire n_2783;
wire n_3188;
wire n_1459;
wire n_2462;
wire n_3243;
wire n_1135;
wire n_2889;
wire n_4034;
wire n_4056;
wire n_4622;
wire n_3960;
wire n_1470;
wire n_4887;
wire n_2732;
wire n_4693;
wire n_4206;
wire n_2249;
wire n_1091;
wire n_2000;
wire n_3862;
wire n_4267;
wire n_2270;
wire n_1425;
wire n_5049;
wire n_983;
wire n_906;
wire n_1390;
wire n_2289;
wire n_1733;
wire n_2955;
wire n_2158;
wire n_4609;
wire n_1855;
wire n_3051;
wire n_3367;
wire n_1687;
wire n_1439;
wire n_2328;
wire n_2859;
wire n_2202;
wire n_1331;
wire n_736;
wire n_3314;
wire n_3525;
wire n_2100;
wire n_5157;
wire n_2993;
wire n_3016;
wire n_4754;
wire n_4647;
wire n_1134;
wire n_3688;
wire n_4003;
wire n_1995;
wire n_3751;
wire n_5223;
wire n_4894;
wire n_4113;
wire n_1889;
wire n_4760;
wire n_1905;
wire n_3466;
wire n_762;
wire n_4983;
wire n_1778;
wire n_1079;
wire n_2139;
wire n_5083;
wire n_4509;
wire n_2875;
wire n_1103;
wire n_3907;
wire n_3338;
wire n_4217;
wire n_4906;
wire n_2219;
wire n_1203;
wire n_3636;
wire n_2327;
wire n_999;
wire n_1254;
wire n_2841;
wire n_4897;
wire n_3539;
wire n_3291;
wire n_4399;
wire n_2304;
wire n_2487;
wire n_3276;
wire n_2597;
wire n_3194;
wire n_5084;
wire n_3572;
wire n_3886;
wire n_4710;
wire n_4420;
wire n_892;
wire n_3637;
wire n_4574;
wire n_1468;
wire n_2855;
wire n_1859;
wire n_2156;
wire n_1718;
wire n_5174;
wire n_4234;
wire n_4101;
wire n_3548;
wire n_5017;
wire n_1768;
wire n_3974;
wire n_1847;
wire n_3634;
wire n_1397;
wire n_3236;
wire n_901;
wire n_2755;
wire n_3141;
wire n_923;
wire n_5096;
wire n_1841;
wire n_4660;
wire n_1623;
wire n_1015;
wire n_3112;
wire n_4797;
wire n_3108;
wire n_4270;
wire n_4151;
wire n_4945;
wire n_3417;
wire n_4124;
wire n_785;
wire n_5153;
wire n_4611;
wire n_2337;
wire n_1356;
wire n_3213;
wire n_4333;
wire n_3820;
wire n_5200;
wire n_2607;
wire n_2890;
wire n_1168;
wire n_5115;
wire n_1943;
wire n_3249;
wire n_1320;
wire n_2722;
wire n_1452;
wire n_2854;
wire n_2499;
wire n_4152;
wire n_1596;
wire n_5092;
wire n_1734;
wire n_3172;
wire n_4832;
wire n_2902;
wire n_3217;
wire n_1983;
wire n_1938;
wire n_2472;
wire n_3394;
wire n_1715;
wire n_3536;
wire n_1443;
wire n_1272;
wire n_2894;
wire n_3957;
wire n_3710;
wire n_4195;
wire n_4554;
wire n_3040;
wire n_3279;
wire n_2402;
wire n_2225;
wire n_1081;
wire n_1692;
wire n_1084;
wire n_1864;
wire n_2006;
wire n_3402;
wire n_3475;
wire n_3501;
wire n_1705;
wire n_3905;
wire n_4680;
wire n_3013;
wire n_921;
wire n_2789;
wire n_5152;
wire n_2257;
wire n_4927;
wire n_4258;
wire n_1828;
wire n_2699;
wire n_2200;
wire n_1940;
wire n_4548;
wire n_4862;
wire n_1405;
wire n_2376;
wire n_3878;
wire n_2670;
wire n_2700;
wire n_1041;
wire n_3134;
wire n_1569;
wire n_3115;
wire n_1062;
wire n_896;
wire n_4553;
wire n_3278;
wire n_2084;
wire n_4875;
wire n_2458;
wire n_1222;
wire n_3050;
wire n_2673;
wire n_2456;
wire n_2527;
wire n_2635;
wire n_1637;
wire n_3307;
wire n_1407;
wire n_1795;
wire n_2871;
wire n_4321;
wire n_4183;
wire n_1271;
wire n_4901;
wire n_1545;
wire n_4821;
wire n_4145;
wire n_3121;
wire n_1640;
wire n_4040;
wire n_2406;
wire n_806;
wire n_2141;
wire n_833;
wire n_3930;
wire n_4943;
wire n_799;
wire n_3044;
wire n_4757;
wire n_2196;
wire n_2629;
wire n_2809;
wire n_787;
wire n_2172;
wire n_4682;
wire n_4530;
wire n_1528;
wire n_1146;
wire n_2021;
wire n_4942;
wire n_1086;
wire n_2125;
wire n_2561;
wire n_4604;
wire n_1906;
wire n_3305;
wire n_2992;
wire n_1241;
wire n_3157;
wire n_4841;
wire n_1758;
wire n_3221;
wire n_3267;
wire n_2422;
wire n_1914;
wire n_1318;
wire n_4338;
wire n_3457;
wire n_3762;
wire n_3005;
wire n_3151;
wire n_3411;
wire n_4840;
wire n_1029;
wire n_4519;
wire n_3779;
wire n_2388;
wire n_3984;
wire n_1706;
wire n_5186;
wire n_1498;
wire n_2417;
wire n_1210;
wire n_5093;
wire n_1556;
wire n_4052;
wire n_3558;
wire n_1984;
wire n_2236;
wire n_4326;
wire n_1269;
wire n_2083;
wire n_2834;
wire n_3207;
wire n_2441;
wire n_3401;
wire n_3242;
wire n_3613;
wire n_4726;
wire n_1045;
wire n_786;
wire n_1559;
wire n_1872;
wire n_5040;
wire n_1325;
wire n_3761;
wire n_4315;
wire n_2923;
wire n_2888;
wire n_1727;
wire n_4301;
wire n_3744;
wire n_4788;
wire n_2041;
wire n_1360;
wire n_3814;
wire n_3781;
wire n_1908;
wire n_2484;
wire n_2126;
wire n_3843;
wire n_1098;
wire n_2045;
wire n_817;
wire n_3687;
wire n_2216;
wire n_3543;
wire n_3621;
wire n_2903;
wire n_3216;
wire n_3808;
wire n_4365;
wire n_1882;
wire n_3726;
wire n_1007;
wire n_1929;
wire n_2369;
wire n_1592;
wire n_2719;
wire n_3758;
wire n_2587;
wire n_3199;
wire n_3339;
wire n_4923;
wire n_2400;
wire n_1953;
wire n_4741;
wire n_3343;
wire n_2752;
wire n_4885;
wire n_751;
wire n_1399;
wire n_4550;
wire n_4652;
wire n_2358;
wire n_3658;
wire n_4900;
wire n_2186;
wire n_2163;
wire n_2815;
wire n_3034;
wire n_4408;
wire n_4577;
wire n_4748;
wire n_2814;
wire n_5209;
wire n_789;
wire n_3231;
wire n_4212;
wire n_2979;
wire n_2953;
wire n_4295;
wire n_2946;
wire n_2500;
wire n_3430;
wire n_2269;
wire n_1729;
wire n_4225;
wire n_747;
wire n_2565;
wire n_1389;
wire n_3583;
wire n_3860;
wire n_3851;
wire n_5064;
wire n_3015;
wire n_2175;
wire n_2182;
wire n_4009;
wire n_1848;
wire n_5002;
wire n_1506;
wire n_3473;
wire n_1652;
wire n_957;
wire n_1994;
wire n_2566;
wire n_744;
wire n_971;
wire n_2702;
wire n_3241;
wire n_2906;
wire n_4342;
wire n_4568;
wire n_1205;
wire n_1258;
wire n_2438;
wire n_2914;
wire n_3100;
wire n_2180;
wire n_2858;
wire n_3573;
wire n_1016;
wire n_4106;
wire n_1501;
wire n_3604;
wire n_4373;
wire n_4711;
wire n_3068;
wire n_2685;
wire n_1083;
wire n_3553;
wire n_2275;
wire n_2465;
wire n_2568;
wire n_2022;
wire n_3811;
wire n_910;
wire n_3494;
wire n_1721;
wire n_1737;
wire n_3486;
wire n_4086;
wire n_908;
wire n_752;
wire n_1028;
wire n_2106;
wire n_2265;
wire n_2032;
wire n_4812;
wire n_4409;
wire n_4629;
wire n_4638;
wire n_708;
wire n_1973;
wire n_3181;
wire n_1500;
wire n_3699;
wire n_854;
wire n_4913;
wire n_2312;
wire n_904;
wire n_1266;
wire n_709;
wire n_2242;
wire n_3328;
wire n_3868;
wire n_1276;
wire n_4266;
wire n_2466;
wire n_2530;
wire n_1085;
wire n_2042;
wire n_771;
wire n_924;
wire n_1582;
wire n_2318;
wire n_3286;
wire n_4012;
wire n_1149;
wire n_3170;
wire n_3645;
wire n_5075;
wire n_3682;
wire n_3304;
wire n_2592;
wire n_4968;
wire n_3771;
wire n_2666;
wire n_1585;
wire n_1799;
wire n_2564;
wire n_5085;
wire n_4259;
wire n_2433;
wire n_829;
wire n_2035;
wire n_3422;
wire n_4572;
wire n_859;
wire n_3086;
wire n_2033;
wire n_4104;
wire n_4845;
wire n_1770;
wire n_878;
wire n_5120;
wire n_3285;
wire n_4208;
wire n_981;
wire n_4089;
wire n_1144;
wire n_2071;
wire n_3219;
wire n_3702;
wire n_2233;
wire n_4779;
wire n_3233;
wire n_4599;
wire n_997;
wire n_4437;
wire n_5222;
wire n_3310;
wire n_1306;
wire n_3264;
wire n_2010;
wire n_1198;
wire n_4061;
wire n_2174;
wire n_3881;
wire n_4508;
wire n_4727;
wire n_4594;
wire n_2426;
wire n_2478;
wire n_1133;
wire n_4429;
wire n_4642;
wire n_4051;
wire n_1051;
wire n_4865;
wire n_1039;
wire n_2043;
wire n_1480;
wire n_3206;
wire n_1305;
wire n_2363;
wire n_2578;
wire n_4562;
wire n_3383;
wire n_4903;
wire n_3709;
wire n_3738;
wire n_4186;
wire n_2540;
wire n_973;
wire n_3610;
wire n_4998;
wire n_3330;
wire n_2065;
wire n_2879;
wire n_967;
wire n_4522;
wire n_2001;
wire n_4341;
wire n_1629;
wire n_4263;
wire n_1260;
wire n_1819;
wire n_3555;
wire n_915;
wire n_812;
wire n_1131;
wire n_3155;
wire n_1006;
wire n_3110;
wire n_1632;
wire n_1888;
wire n_1311;
wire n_4780;
wire n_2697;
wire n_3908;
wire n_4973;
wire n_3467;
wire n_1887;
wire n_1587;
wire n_3916;
wire n_3527;
wire n_4803;
wire n_2512;
wire n_3950;
wire n_1242;
wire n_2086;
wire n_2927;
wire n_4750;
wire n_3039;
wire n_1226;
wire n_3740;
wire n_2166;
wire n_2899;
wire n_3186;
wire n_1322;
wire n_1958;
wire n_1197;
wire n_3065;
wire n_2632;
wire n_4984;
wire n_2579;
wire n_2105;
wire n_1423;
wire n_3387;
wire n_3420;
wire n_5041;
wire n_1915;
wire n_4275;
wire n_4283;
wire n_4959;
wire n_900;
wire n_4426;
wire n_2912;
wire n_2659;
wire n_4425;
wire n_3409;
wire n_4449;
wire n_2116;
wire n_2320;
wire n_1013;
wire n_1259;
wire n_2183;
wire n_3002;
wire n_1612;
wire n_4809;
wire n_1199;
wire n_3392;
wire n_3773;
wire n_2003;
wire n_1038;
wire n_1581;
wire n_3301;
wire n_1357;
wire n_4241;
wire n_1853;
wire n_798;
wire n_2324;
wire n_1348;
wire n_2977;
wire n_1739;
wire n_1380;
wire n_2847;
wire n_2557;
wire n_1009;
wire n_2405;
wire n_4050;
wire n_1160;
wire n_883;
wire n_2647;
wire n_1032;
wire n_2336;
wire n_1247;
wire n_2521;
wire n_1099;
wire n_4578;
wire n_2211;
wire n_4777;
wire n_2672;
wire n_4702;
wire n_2299;
wire n_4179;
wire n_4895;
wire n_1285;
wire n_1985;
wire n_1172;
wire n_4026;
wire n_4531;
wire n_3282;
wire n_1590;
wire n_3626;
wire n_1532;
wire n_2313;
wire n_5072;
wire n_3106;
wire n_1140;
wire n_1670;
wire n_2344;
wire n_2365;
wire n_4666;
wire n_3031;
wire n_4029;
wire n_2447;
wire n_4617;
wire n_2340;
wire n_4010;
wire n_1649;
wire n_4555;
wire n_4969;
wire n_5105;
wire n_1572;
wire n_4308;
wire n_5021;
wire n_3463;
wire n_2510;
wire n_1954;
wire n_822;
wire n_2791;
wire n_4325;
wire n_3251;
wire n_4602;
wire n_5044;
wire n_5134;
wire n_2212;
wire n_3063;
wire n_1163;
wire n_2729;
wire n_2582;
wire n_1798;
wire n_1550;
wire n_3998;
wire n_1591;
wire n_3632;
wire n_3122;
wire n_1344;
wire n_2730;
wire n_2495;
wire n_2090;
wire n_2603;
wire n_3829;
wire n_4164;
wire n_2173;
wire n_1471;
wire n_4919;
wire n_3737;
wire n_3655;
wire n_3825;
wire n_2880;
wire n_3225;
wire n_2108;
wire n_5158;
wire n_1211;
wire n_5022;
wire n_1280;
wire n_3296;
wire n_1445;
wire n_2551;
wire n_1526;
wire n_5047;
wire n_2985;
wire n_1978;
wire n_3792;
wire n_4202;
wire n_1446;
wire n_3938;
wire n_4791;
wire n_3507;
wire n_4403;
wire n_3269;
wire n_3531;
wire n_1054;
wire n_1956;
wire n_4139;
wire n_4549;
wire n_1986;
wire n_2397;
wire n_3931;
wire n_4349;
wire n_5141;
wire n_2113;
wire n_1918;
wire n_3603;
wire n_813;
wire n_3822;
wire n_4163;
wire n_818;
wire n_3812;
wire n_3910;
wire n_2633;
wire n_2207;
wire n_4948;
wire n_2696;
wire n_3482;
wire n_4080;
wire n_2198;
wire n_3319;
wire n_2073;
wire n_2273;
wire n_3748;
wire n_3272;
wire n_4941;
wire n_3396;
wire n_4393;
wire n_1162;
wire n_4372;
wire n_821;
wire n_1068;
wire n_982;
wire n_932;
wire n_2831;
wire n_4318;
wire n_4158;
wire n_3317;
wire n_3978;
wire n_2123;
wire n_1697;
wire n_979;
wire n_4074;
wire n_3716;
wire n_4795;
wire n_4918;
wire n_3824;
wire n_5067;
wire n_4013;
wire n_4544;
wire n_3248;
wire n_2941;
wire n_1278;
wire n_5108;
wire n_4032;
wire n_1064;
wire n_1396;
wire n_2355;
wire n_4147;
wire n_4477;
wire n_3168;
wire n_2751;
wire n_4337;
wire n_4130;
wire n_2009;
wire n_1793;
wire n_3601;
wire n_3092;
wire n_1289;
wire n_3055;
wire n_3966;
wire n_2866;
wire n_4742;
wire n_1014;
wire n_3734;
wire n_1703;
wire n_2580;
wire n_882;
wire n_3649;
wire n_2821;
wire n_1875;
wire n_1865;
wire n_3746;
wire n_3384;
wire n_1950;
wire n_1563;
wire n_3419;
wire n_1297;
wire n_1662;
wire n_4478;
wire n_1359;
wire n_2818;
wire n_3794;
wire n_3921;
wire n_922;
wire n_1335;
wire n_1927;
wire n_4838;
wire n_5202;
wire n_702;
wire n_4965;
wire n_3346;
wire n_1896;
wire n_2965;
wire n_3058;
wire n_3861;
wire n_1540;
wire n_1977;
wire n_3891;
wire n_2193;
wire n_4523;
wire n_1655;
wire n_1886;
wire n_4371;
wire n_2994;
wire n_3428;
wire n_3153;
wire n_4552;
wire n_3689;
wire n_877;
wire n_4673;
wire n_2519;
wire n_728;
wire n_3415;
wire n_1063;
wire n_4607;
wire n_4041;
wire n_2947;
wire n_3918;
wire n_1965;
wire n_4837;
wire n_2476;
wire n_4169;
wire n_3271;
wire n_5088;
wire n_4248;
wire n_2976;
wire n_2152;
wire n_2652;
wire n_1825;
wire n_1757;
wire n_1792;
wire n_1412;
wire n_2497;
wire n_3809;
wire n_3139;
wire n_4070;
wire n_3545;
wire n_3885;
wire n_1369;
wire n_881;
wire n_3993;
wire n_4685;
wire n_4031;
wire n_4675;
wire n_2663;
wire n_4018;
wire n_2987;
wire n_2938;
wire n_3780;
wire n_3337;
wire n_4002;
wire n_3209;
wire n_5178;
wire n_1044;
wire n_2165;
wire n_1391;
wire n_2750;
wire n_2775;
wire n_1295;
wire n_3477;
wire n_2349;
wire n_2684;
wire n_3146;
wire n_1495;
wire n_1438;
wire n_3953;
wire n_4588;
wire n_1100;
wire n_4653;
wire n_4435;
wire n_1756;
wire n_1128;
wire n_4019;
wire n_1071;
wire n_1968;
wire n_4728;
wire n_4999;
wire n_4385;
wire n_4922;
wire n_865;
wire n_3616;
wire n_4191;
wire n_2870;
wire n_2151;
wire n_1839;
wire n_2341;
wire n_1765;
wire n_3727;
wire n_5235;
wire n_2707;
wire n_826;
wire n_4350;
wire n_3747;
wire n_1714;
wire n_718;
wire n_4330;
wire n_2089;
wire n_3522;
wire n_2747;
wire n_3924;
wire n_791;
wire n_4621;
wire n_4216;
wire n_4240;
wire n_3491;
wire n_1488;
wire n_704;
wire n_2148;
wire n_4162;
wire n_2339;
wire n_2861;
wire n_1999;
wire n_2731;
wire n_3353;
wire n_3018;
wire n_3975;
wire n_1838;
wire n_2638;
wire n_4785;
wire n_4683;
wire n_1766;
wire n_1776;
wire n_2002;
wire n_2138;
wire n_4021;
wire n_2414;
wire n_3014;
wire n_1771;
wire n_2316;
wire n_4103;
wire n_5060;
wire n_3148;
wire n_4022;
wire n_4986;
wire n_2208;
wire n_4775;
wire n_4864;
wire n_4674;
wire n_4481;
wire n_1304;
wire n_3775;
wire n_4669;
wire n_2134;
wire n_1176;
wire n_1431;
wire n_3312;
wire n_3835;
wire n_4286;
wire n_2958;
wire n_3731;
wire n_1822;
wire n_2936;
wire n_3224;
wire n_2489;
wire n_1087;
wire n_2771;
wire n_3020;
wire n_4525;
wire n_1505;
wire n_3557;
wire n_2610;
wire n_3129;
wire n_3620;
wire n_3832;
wire n_2520;
wire n_4484;
wire n_3693;
wire n_4497;
wire n_1568;
wire n_2372;
wire n_1490;
wire n_2251;
wire n_3674;
wire n_2959;
wire n_2501;
wire n_3203;
wire n_4871;
wire n_1070;
wire n_2403;
wire n_2837;
wire n_4700;
wire n_4883;
wire n_1665;
wire n_4306;
wire n_4224;
wire n_2127;
wire n_3341;
wire n_4453;
wire n_3559;
wire n_4005;
wire n_3546;
wire n_1358;
wire n_3661;
wire n_4564;
wire n_5146;
wire n_3056;
wire n_745;
wire n_2424;
wire n_3201;
wire n_3447;
wire n_3971;
wire n_716;
wire n_1475;
wire n_1774;
wire n_2354;
wire n_3103;
wire n_4573;
wire n_2589;
wire n_4535;
wire n_755;
wire n_2442;
wire n_3627;
wire n_3480;
wire n_1368;
wire n_1137;
wire n_3612;
wire n_4695;
wire n_2545;
wire n_3509;
wire n_4368;
wire n_2966;
wire n_2294;
wire n_1942;
wire n_1314;
wire n_3196;
wire n_864;
wire n_2504;
wire n_2623;
wire n_1440;
wire n_2063;
wire n_1534;
wire n_5005;
wire n_1339;
wire n_2475;
wire n_5181;
wire n_723;
wire n_3144;
wire n_3244;
wire n_1141;
wire n_1268;
wire n_3287;
wire n_3322;
wire n_1755;
wire n_5043;
wire n_2025;
wire n_2357;
wire n_4654;
wire n_3640;
wire n_995;
wire n_1159;
wire n_3481;
wire n_2250;
wire n_3033;
wire n_2374;
wire n_1681;
wire n_4597;
wire n_3364;
wire n_3226;
wire n_2780;
wire n_4020;
wire n_5220;
wire n_1618;
wire n_4867;
wire n_5061;
wire n_1653;
wire n_4063;
wire n_4237;
wire n_2601;
wire n_5029;
wire n_5127;
wire n_2920;
wire n_773;
wire n_920;
wire n_1374;
wire n_2648;
wire n_3212;
wire n_1169;
wire n_1617;
wire n_3370;
wire n_3386;
wire n_4721;
wire n_3093;
wire n_848;
wire n_4247;
wire n_3169;
wire n_3205;
wire n_1881;
wire n_1267;
wire n_1806;
wire n_2023;
wire n_2204;
wire n_2720;
wire n_4614;
wire n_3360;
wire n_2087;
wire n_1636;
wire n_3956;
wire n_4001;
wire n_1323;
wire n_2627;
wire n_4422;
wire n_960;
wire n_778;
wire n_3004;
wire n_3870;
wire n_5177;
wire n_3625;
wire n_1764;
wire n_4632;
wire n_1610;
wire n_3084;
wire n_2343;
wire n_793;
wire n_4546;
wire n_4583;
wire n_4963;
wire n_3749;
wire n_2942;
wire n_4966;
wire n_4714;
wire n_5037;
wire n_2515;
wire n_1551;
wire n_4847;
wire n_4054;
wire n_2555;
wire n_3586;
wire n_3653;
wire n_2201;
wire n_725;
wire n_3349;
wire n_4668;
wire n_5213;
wire n_4635;
wire n_994;
wire n_2278;
wire n_1020;
wire n_1273;
wire n_4214;
wire n_3448;
wire n_2924;
wire n_1036;
wire n_3595;
wire n_1138;
wire n_1661;
wire n_3991;
wire n_3516;
wire n_3926;
wire n_1095;
wire n_1270;
wire n_4405;
wire n_4413;
wire n_1852;
wire n_4036;
wire n_4759;
wire n_2153;
wire n_3670;
wire n_2381;
wire n_2052;
wire n_4667;
wire n_5081;
wire n_4182;
wire n_3230;
wire n_1279;
wire n_1115;
wire n_1499;
wire n_1409;
wire n_5189;
wire n_1503;
wire n_2819;
wire n_3041;
wire n_4637;
wire n_2423;
wire n_1657;
wire n_1126;
wire n_2412;
wire n_2439;
wire n_2404;
wire n_1182;
wire n_3635;
wire n_5118;
wire n_4155;
wire n_4238;
wire n_3011;
wire n_2061;
wire n_2757;
wire n_4977;
wire n_1216;
wire n_2716;
wire n_2452;
wire n_3650;
wire n_3010;
wire n_3043;
wire n_5224;
wire n_4590;
wire n_2543;
wire n_5090;
wire n_3137;
wire n_2486;
wire n_3560;
wire n_3177;
wire n_4929;
wire n_2220;
wire n_2577;
wire n_1262;
wire n_3238;
wire n_3529;
wire n_4835;
wire n_2232;
wire n_4038;
wire n_2790;
wire n_4565;
wire n_4159;
wire n_3784;
wire n_4586;
wire n_1608;
wire n_2373;
wire n_1472;
wire n_3628;
wire n_800;
wire n_4734;
wire n_1491;
wire n_1840;
wire n_4434;
wire n_2244;
wire n_4290;
wire n_2586;
wire n_1684;
wire n_2446;
wire n_1346;
wire n_1352;
wire n_2017;
wire n_3029;
wire n_3597;
wire n_1046;
wire n_2560;
wire n_2704;
wire n_1145;
wire n_1121;
wire n_1102;
wire n_1963;
wire n_3790;
wire n_2766;
wire n_3318;
wire n_4833;
wire n_5062;
wire n_5230;
wire n_4888;
wire n_776;
wire n_1823;
wire n_2479;
wire n_3350;
wire n_2782;
wire n_3977;
wire n_3588;
wire n_4279;
wire n_5008;
wire n_1456;
wire n_5004;
wire n_2229;
wire n_4133;
wire n_4527;
wire n_2288;
wire n_2099;
wire n_3388;
wire n_4790;
wire n_1946;
wire n_4181;
wire n_3184;
wire n_4561;
wire n_4461;
wire n_3245;
wire n_3075;
wire n_4007;
wire n_4949;
wire n_2642;
wire n_4239;
wire n_2383;
wire n_4184;
wire n_1676;
wire n_1830;
wire n_2351;
wire n_1319;
wire n_5069;
wire n_2986;
wire n_2536;
wire n_3915;
wire n_1633;
wire n_3489;
wire n_2835;
wire n_1416;
wire n_2820;
wire n_2293;
wire n_3074;
wire n_3102;
wire n_2026;
wire n_1282;
wire n_3321;
wire n_2567;
wire n_2322;
wire n_2727;
wire n_3377;
wire n_4782;
wire n_1321;
wire n_2533;
wire n_3530;
wire n_2869;
wire n_4378;
wire n_1235;
wire n_2759;
wire n_2361;
wire n_1292;
wire n_2266;
wire n_4876;
wire n_790;
wire n_2611;
wire n_2901;
wire n_4358;
wire n_2653;
wire n_1248;
wire n_902;
wire n_2189;
wire n_2246;
wire n_4469;
wire n_5169;
wire n_3156;
wire n_1941;
wire n_3483;
wire n_706;
wire n_1794;
wire n_1236;
wire n_4493;
wire n_4924;
wire n_743;
wire n_766;
wire n_1746;
wire n_3524;
wire n_2885;
wire n_3097;
wire n_2062;
wire n_4539;
wire n_2975;
wire n_4421;
wire n_2839;
wire n_2856;
wire n_4793;
wire n_4498;
wire n_2070;
wire n_1607;
wire n_1454;
wire n_4953;
wire n_2348;
wire n_2944;
wire n_3831;
wire n_869;
wire n_1154;
wire n_1329;
wire n_5167;
wire n_3589;
wire n_897;
wire n_846;
wire n_2066;
wire n_841;
wire n_1476;
wire n_3391;
wire n_1800;
wire n_1463;
wire n_3458;
wire n_4505;
wire n_3190;
wire n_1562;
wire n_1826;
wire n_5126;
wire n_1759;
wire n_5051;
wire n_5236;
wire n_853;
wire n_875;
wire n_5012;
wire n_1678;
wire n_3787;
wire n_1256;
wire n_3585;
wire n_3565;
wire n_4450;
wire n_5025;
wire n_933;
wire n_4173;
wire n_3135;
wire n_4630;
wire n_1217;
wire n_3990;
wire n_1628;
wire n_2109;
wire n_988;
wire n_2796;
wire n_2507;
wire n_4534;
wire n_1536;
wire n_1204;
wire n_1132;
wire n_1327;
wire n_955;
wire n_2787;
wire n_2969;
wire n_2395;
wire n_1554;
wire n_4494;
wire n_769;
wire n_2380;
wire n_4786;
wire n_1120;
wire n_4579;
wire n_2290;
wire n_4811;
wire n_2048;
wire n_2005;
wire n_4857;
wire n_3432;
wire n_2736;
wire n_2883;
wire n_1408;
wire n_4282;
wire n_1196;
wire n_3493;
wire n_863;
wire n_3774;
wire n_2910;
wire n_748;
wire n_3268;
wire n_1785;
wire n_1147;
wire n_1754;
wire n_3057;
wire n_3701;
wire n_5148;
wire n_2584;
wire n_1812;
wire n_866;
wire n_2287;
wire n_761;
wire n_2492;
wire n_3778;
wire n_1173;
wire n_4974;
wire n_4911;
wire n_4436;
wire n_5119;
wire n_4569;
wire n_1174;
wire n_3334;
wire n_5097;
wire n_844;
wire n_4985;
wire n_2117;
wire n_2234;
wire n_3823;
wire n_4384;
wire n_2741;
wire n_3114;
wire n_888;
wire n_2203;
wire n_2255;
wire n_3584;
wire n_4858;
wire n_4678;
wire n_2649;
wire n_3556;
wire n_3836;
wire n_1922;
wire n_4823;
wire n_4309;
wire n_4363;
wire n_1215;
wire n_839;
wire n_5107;
wire n_3456;
wire n_5095;
wire n_779;
wire n_1537;
wire n_2205;
wire n_4243;
wire n_4025;
wire n_3404;
wire n_1122;
wire n_4059;
wire n_1509;
wire n_4121;
wire n_3290;
wire n_1109;
wire n_4313;
wire n_3309;
wire n_3671;
wire n_4142;
wire n_2015;
wire n_3982;
wire n_2609;
wire n_1161;
wire n_3796;
wire n_3840;
wire n_3461;
wire n_3408;
wire n_4246;
wire n_3513;
wire n_3690;
wire n_1184;
wire n_2483;
wire n_4532;
wire n_1525;
wire n_3995;
wire n_4076;
wire n_2594;
wire n_4244;
wire n_2147;
wire n_2503;
wire n_4049;
wire n_1156;
wire n_2600;
wire n_984;
wire n_3508;
wire n_868;
wire n_4353;
wire n_735;
wire n_4787;
wire n_1218;
wire n_3596;
wire n_4537;
wire n_4346;
wire n_4351;
wire n_2429;
wire n_985;
wire n_2440;
wire n_3521;
wire n_802;
wire n_980;
wire n_2681;
wire n_1651;
wire n_2360;
wire n_3764;
wire n_4784;
wire n_4075;
wire n_3947;
wire n_1244;
wire n_1685;
wire n_3066;
wire n_2844;
wire n_2303;
wire n_1619;
wire n_2285;
wire n_4451;
wire n_4332;
wire n_810;
wire n_1194;
wire n_4538;
wire n_4506;
wire n_2742;
wire n_3695;
wire n_3976;
wire n_3563;
wire n_2367;
wire n_3198;
wire n_3495;
wire n_1034;
wire n_2909;
wire n_754;
wire n_975;
wire n_3359;
wire n_3187;
wire n_3218;
wire n_861;
wire n_857;
wire n_2107;
wire n_2040;
wire n_2968;
wire n_4201;
wire n_4336;
wire n_2221;
wire n_4852;
wire n_1010;
wire n_4210;
wire n_4981;
wire n_1166;
wire n_2891;
wire n_2709;
wire n_1578;
wire n_1861;
wire n_3955;
wire n_1557;
wire n_2280;
wire n_3945;
wire n_730;
wire n_5214;
wire n_1898;
wire n_2443;
wire n_4936;
wire n_4205;
wire n_2162;
wire n_1868;
wire n_2079;
wire n_4763;
wire n_3587;
wire n_4278;
wire n_3433;
wire n_4463;
wire n_2185;
wire n_1836;
wire n_3833;
wire n_2774;
wire n_3162;
wire n_1274;
wire n_1486;
wire n_3333;
wire n_4129;
wire n_5032;
wire n_1899;
wire n_784;
wire n_4804;
wire n_3965;
wire n_4500;
wire n_5065;
wire n_862;
wire n_2098;
wire n_3085;
wire n_4433;
wire n_2813;
wire n_1935;
wire n_2027;
wire n_2091;
wire n_2991;
wire n_5030;
wire n_4194;
wire n_1449;
wire n_4703;
wire n_2419;
wire n_2677;
wire n_3182;
wire n_3283;
wire n_1742;
wire n_4030;

CKINVDCx5p33_ASAP7_75t_R g699 ( 
.A(n_624),
.Y(n_699)
);

CKINVDCx5p33_ASAP7_75t_R g700 ( 
.A(n_271),
.Y(n_700)
);

CKINVDCx5p33_ASAP7_75t_R g701 ( 
.A(n_554),
.Y(n_701)
);

CKINVDCx5p33_ASAP7_75t_R g702 ( 
.A(n_194),
.Y(n_702)
);

BUFx10_ASAP7_75t_L g703 ( 
.A(n_93),
.Y(n_703)
);

CKINVDCx5p33_ASAP7_75t_R g704 ( 
.A(n_642),
.Y(n_704)
);

CKINVDCx5p33_ASAP7_75t_R g705 ( 
.A(n_379),
.Y(n_705)
);

CKINVDCx5p33_ASAP7_75t_R g706 ( 
.A(n_395),
.Y(n_706)
);

CKINVDCx5p33_ASAP7_75t_R g707 ( 
.A(n_192),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_618),
.Y(n_708)
);

CKINVDCx5p33_ASAP7_75t_R g709 ( 
.A(n_618),
.Y(n_709)
);

BUFx6f_ASAP7_75t_L g710 ( 
.A(n_560),
.Y(n_710)
);

CKINVDCx5p33_ASAP7_75t_R g711 ( 
.A(n_24),
.Y(n_711)
);

CKINVDCx5p33_ASAP7_75t_R g712 ( 
.A(n_547),
.Y(n_712)
);

CKINVDCx5p33_ASAP7_75t_R g713 ( 
.A(n_8),
.Y(n_713)
);

BUFx5_ASAP7_75t_L g714 ( 
.A(n_173),
.Y(n_714)
);

INVx2_ASAP7_75t_L g715 ( 
.A(n_80),
.Y(n_715)
);

CKINVDCx5p33_ASAP7_75t_R g716 ( 
.A(n_50),
.Y(n_716)
);

HB1xp67_ASAP7_75t_L g717 ( 
.A(n_12),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_641),
.Y(n_718)
);

INVx2_ASAP7_75t_SL g719 ( 
.A(n_131),
.Y(n_719)
);

CKINVDCx5p33_ASAP7_75t_R g720 ( 
.A(n_140),
.Y(n_720)
);

CKINVDCx20_ASAP7_75t_R g721 ( 
.A(n_139),
.Y(n_721)
);

CKINVDCx5p33_ASAP7_75t_R g722 ( 
.A(n_379),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_625),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_649),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_371),
.Y(n_725)
);

BUFx2_ASAP7_75t_L g726 ( 
.A(n_539),
.Y(n_726)
);

INVx2_ASAP7_75t_L g727 ( 
.A(n_246),
.Y(n_727)
);

CKINVDCx5p33_ASAP7_75t_R g728 ( 
.A(n_118),
.Y(n_728)
);

CKINVDCx16_ASAP7_75t_R g729 ( 
.A(n_61),
.Y(n_729)
);

CKINVDCx5p33_ASAP7_75t_R g730 ( 
.A(n_86),
.Y(n_730)
);

CKINVDCx5p33_ASAP7_75t_R g731 ( 
.A(n_309),
.Y(n_731)
);

CKINVDCx5p33_ASAP7_75t_R g732 ( 
.A(n_487),
.Y(n_732)
);

CKINVDCx5p33_ASAP7_75t_R g733 ( 
.A(n_235),
.Y(n_733)
);

CKINVDCx5p33_ASAP7_75t_R g734 ( 
.A(n_277),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_435),
.Y(n_735)
);

CKINVDCx20_ASAP7_75t_R g736 ( 
.A(n_515),
.Y(n_736)
);

CKINVDCx5p33_ASAP7_75t_R g737 ( 
.A(n_569),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_363),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_374),
.Y(n_739)
);

CKINVDCx5p33_ASAP7_75t_R g740 ( 
.A(n_256),
.Y(n_740)
);

CKINVDCx5p33_ASAP7_75t_R g741 ( 
.A(n_120),
.Y(n_741)
);

CKINVDCx5p33_ASAP7_75t_R g742 ( 
.A(n_634),
.Y(n_742)
);

CKINVDCx5p33_ASAP7_75t_R g743 ( 
.A(n_87),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_600),
.Y(n_744)
);

CKINVDCx5p33_ASAP7_75t_R g745 ( 
.A(n_389),
.Y(n_745)
);

CKINVDCx5p33_ASAP7_75t_R g746 ( 
.A(n_280),
.Y(n_746)
);

CKINVDCx5p33_ASAP7_75t_R g747 ( 
.A(n_408),
.Y(n_747)
);

CKINVDCx5p33_ASAP7_75t_R g748 ( 
.A(n_20),
.Y(n_748)
);

CKINVDCx5p33_ASAP7_75t_R g749 ( 
.A(n_291),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_101),
.Y(n_750)
);

CKINVDCx5p33_ASAP7_75t_R g751 ( 
.A(n_480),
.Y(n_751)
);

CKINVDCx5p33_ASAP7_75t_R g752 ( 
.A(n_257),
.Y(n_752)
);

CKINVDCx5p33_ASAP7_75t_R g753 ( 
.A(n_664),
.Y(n_753)
);

CKINVDCx14_ASAP7_75t_R g754 ( 
.A(n_530),
.Y(n_754)
);

CKINVDCx5p33_ASAP7_75t_R g755 ( 
.A(n_538),
.Y(n_755)
);

CKINVDCx5p33_ASAP7_75t_R g756 ( 
.A(n_126),
.Y(n_756)
);

CKINVDCx20_ASAP7_75t_R g757 ( 
.A(n_385),
.Y(n_757)
);

CKINVDCx5p33_ASAP7_75t_R g758 ( 
.A(n_467),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_392),
.Y(n_759)
);

CKINVDCx5p33_ASAP7_75t_R g760 ( 
.A(n_483),
.Y(n_760)
);

HB1xp67_ASAP7_75t_L g761 ( 
.A(n_619),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_362),
.Y(n_762)
);

INVx2_ASAP7_75t_L g763 ( 
.A(n_675),
.Y(n_763)
);

CKINVDCx5p33_ASAP7_75t_R g764 ( 
.A(n_698),
.Y(n_764)
);

CKINVDCx5p33_ASAP7_75t_R g765 ( 
.A(n_319),
.Y(n_765)
);

CKINVDCx5p33_ASAP7_75t_R g766 ( 
.A(n_462),
.Y(n_766)
);

CKINVDCx5p33_ASAP7_75t_R g767 ( 
.A(n_78),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_271),
.Y(n_768)
);

CKINVDCx5p33_ASAP7_75t_R g769 ( 
.A(n_341),
.Y(n_769)
);

CKINVDCx20_ASAP7_75t_R g770 ( 
.A(n_198),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_21),
.Y(n_771)
);

BUFx10_ASAP7_75t_L g772 ( 
.A(n_295),
.Y(n_772)
);

CKINVDCx5p33_ASAP7_75t_R g773 ( 
.A(n_167),
.Y(n_773)
);

CKINVDCx5p33_ASAP7_75t_R g774 ( 
.A(n_163),
.Y(n_774)
);

CKINVDCx20_ASAP7_75t_R g775 ( 
.A(n_249),
.Y(n_775)
);

CKINVDCx5p33_ASAP7_75t_R g776 ( 
.A(n_169),
.Y(n_776)
);

CKINVDCx5p33_ASAP7_75t_R g777 ( 
.A(n_41),
.Y(n_777)
);

CKINVDCx12_ASAP7_75t_R g778 ( 
.A(n_273),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_566),
.Y(n_779)
);

CKINVDCx12_ASAP7_75t_R g780 ( 
.A(n_392),
.Y(n_780)
);

CKINVDCx20_ASAP7_75t_R g781 ( 
.A(n_53),
.Y(n_781)
);

CKINVDCx5p33_ASAP7_75t_R g782 ( 
.A(n_595),
.Y(n_782)
);

CKINVDCx5p33_ASAP7_75t_R g783 ( 
.A(n_423),
.Y(n_783)
);

CKINVDCx5p33_ASAP7_75t_R g784 ( 
.A(n_583),
.Y(n_784)
);

CKINVDCx5p33_ASAP7_75t_R g785 ( 
.A(n_648),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_206),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_571),
.Y(n_787)
);

CKINVDCx20_ASAP7_75t_R g788 ( 
.A(n_437),
.Y(n_788)
);

CKINVDCx5p33_ASAP7_75t_R g789 ( 
.A(n_601),
.Y(n_789)
);

CKINVDCx5p33_ASAP7_75t_R g790 ( 
.A(n_293),
.Y(n_790)
);

BUFx3_ASAP7_75t_L g791 ( 
.A(n_267),
.Y(n_791)
);

INVx2_ASAP7_75t_L g792 ( 
.A(n_527),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_337),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_595),
.Y(n_794)
);

CKINVDCx5p33_ASAP7_75t_R g795 ( 
.A(n_530),
.Y(n_795)
);

CKINVDCx5p33_ASAP7_75t_R g796 ( 
.A(n_593),
.Y(n_796)
);

CKINVDCx5p33_ASAP7_75t_R g797 ( 
.A(n_7),
.Y(n_797)
);

CKINVDCx5p33_ASAP7_75t_R g798 ( 
.A(n_274),
.Y(n_798)
);

CKINVDCx5p33_ASAP7_75t_R g799 ( 
.A(n_435),
.Y(n_799)
);

CKINVDCx5p33_ASAP7_75t_R g800 ( 
.A(n_310),
.Y(n_800)
);

CKINVDCx5p33_ASAP7_75t_R g801 ( 
.A(n_666),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_539),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_61),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_6),
.Y(n_804)
);

HB1xp67_ASAP7_75t_L g805 ( 
.A(n_401),
.Y(n_805)
);

CKINVDCx5p33_ASAP7_75t_R g806 ( 
.A(n_241),
.Y(n_806)
);

CKINVDCx5p33_ASAP7_75t_R g807 ( 
.A(n_186),
.Y(n_807)
);

INVx1_ASAP7_75t_SL g808 ( 
.A(n_204),
.Y(n_808)
);

CKINVDCx5p33_ASAP7_75t_R g809 ( 
.A(n_51),
.Y(n_809)
);

INVx2_ASAP7_75t_L g810 ( 
.A(n_470),
.Y(n_810)
);

CKINVDCx5p33_ASAP7_75t_R g811 ( 
.A(n_184),
.Y(n_811)
);

BUFx10_ASAP7_75t_L g812 ( 
.A(n_124),
.Y(n_812)
);

CKINVDCx5p33_ASAP7_75t_R g813 ( 
.A(n_668),
.Y(n_813)
);

BUFx3_ASAP7_75t_L g814 ( 
.A(n_159),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_165),
.Y(n_815)
);

CKINVDCx5p33_ASAP7_75t_R g816 ( 
.A(n_408),
.Y(n_816)
);

CKINVDCx5p33_ASAP7_75t_R g817 ( 
.A(n_682),
.Y(n_817)
);

BUFx3_ASAP7_75t_L g818 ( 
.A(n_111),
.Y(n_818)
);

CKINVDCx5p33_ASAP7_75t_R g819 ( 
.A(n_94),
.Y(n_819)
);

CKINVDCx5p33_ASAP7_75t_R g820 ( 
.A(n_454),
.Y(n_820)
);

INVx1_ASAP7_75t_SL g821 ( 
.A(n_592),
.Y(n_821)
);

CKINVDCx5p33_ASAP7_75t_R g822 ( 
.A(n_266),
.Y(n_822)
);

BUFx10_ASAP7_75t_L g823 ( 
.A(n_693),
.Y(n_823)
);

CKINVDCx5p33_ASAP7_75t_R g824 ( 
.A(n_22),
.Y(n_824)
);

CKINVDCx5p33_ASAP7_75t_R g825 ( 
.A(n_284),
.Y(n_825)
);

CKINVDCx5p33_ASAP7_75t_R g826 ( 
.A(n_686),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_77),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_447),
.Y(n_828)
);

CKINVDCx5p33_ASAP7_75t_R g829 ( 
.A(n_375),
.Y(n_829)
);

CKINVDCx5p33_ASAP7_75t_R g830 ( 
.A(n_545),
.Y(n_830)
);

CKINVDCx20_ASAP7_75t_R g831 ( 
.A(n_331),
.Y(n_831)
);

CKINVDCx5p33_ASAP7_75t_R g832 ( 
.A(n_29),
.Y(n_832)
);

CKINVDCx5p33_ASAP7_75t_R g833 ( 
.A(n_670),
.Y(n_833)
);

CKINVDCx5p33_ASAP7_75t_R g834 ( 
.A(n_332),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_607),
.Y(n_835)
);

INVx1_ASAP7_75t_SL g836 ( 
.A(n_437),
.Y(n_836)
);

CKINVDCx20_ASAP7_75t_R g837 ( 
.A(n_134),
.Y(n_837)
);

CKINVDCx5p33_ASAP7_75t_R g838 ( 
.A(n_70),
.Y(n_838)
);

CKINVDCx5p33_ASAP7_75t_R g839 ( 
.A(n_495),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_182),
.Y(n_840)
);

CKINVDCx14_ASAP7_75t_R g841 ( 
.A(n_404),
.Y(n_841)
);

CKINVDCx5p33_ASAP7_75t_R g842 ( 
.A(n_555),
.Y(n_842)
);

CKINVDCx5p33_ASAP7_75t_R g843 ( 
.A(n_91),
.Y(n_843)
);

INVx1_ASAP7_75t_SL g844 ( 
.A(n_645),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_594),
.Y(n_845)
);

CKINVDCx5p33_ASAP7_75t_R g846 ( 
.A(n_602),
.Y(n_846)
);

CKINVDCx5p33_ASAP7_75t_R g847 ( 
.A(n_192),
.Y(n_847)
);

INVx1_ASAP7_75t_L g848 ( 
.A(n_547),
.Y(n_848)
);

INVx1_ASAP7_75t_SL g849 ( 
.A(n_337),
.Y(n_849)
);

BUFx3_ASAP7_75t_L g850 ( 
.A(n_303),
.Y(n_850)
);

CKINVDCx5p33_ASAP7_75t_R g851 ( 
.A(n_296),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_146),
.Y(n_852)
);

CKINVDCx5p33_ASAP7_75t_R g853 ( 
.A(n_196),
.Y(n_853)
);

CKINVDCx5p33_ASAP7_75t_R g854 ( 
.A(n_151),
.Y(n_854)
);

CKINVDCx5p33_ASAP7_75t_R g855 ( 
.A(n_86),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_40),
.Y(n_856)
);

CKINVDCx5p33_ASAP7_75t_R g857 ( 
.A(n_36),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_226),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_242),
.Y(n_859)
);

CKINVDCx5p33_ASAP7_75t_R g860 ( 
.A(n_25),
.Y(n_860)
);

BUFx6f_ASAP7_75t_L g861 ( 
.A(n_587),
.Y(n_861)
);

CKINVDCx5p33_ASAP7_75t_R g862 ( 
.A(n_280),
.Y(n_862)
);

CKINVDCx5p33_ASAP7_75t_R g863 ( 
.A(n_248),
.Y(n_863)
);

CKINVDCx5p33_ASAP7_75t_R g864 ( 
.A(n_290),
.Y(n_864)
);

BUFx6f_ASAP7_75t_L g865 ( 
.A(n_199),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_19),
.Y(n_866)
);

CKINVDCx16_ASAP7_75t_R g867 ( 
.A(n_642),
.Y(n_867)
);

CKINVDCx5p33_ASAP7_75t_R g868 ( 
.A(n_0),
.Y(n_868)
);

CKINVDCx5p33_ASAP7_75t_R g869 ( 
.A(n_52),
.Y(n_869)
);

INVx2_ASAP7_75t_L g870 ( 
.A(n_662),
.Y(n_870)
);

CKINVDCx5p33_ASAP7_75t_R g871 ( 
.A(n_173),
.Y(n_871)
);

CKINVDCx5p33_ASAP7_75t_R g872 ( 
.A(n_492),
.Y(n_872)
);

BUFx6f_ASAP7_75t_L g873 ( 
.A(n_554),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_629),
.Y(n_874)
);

INVx1_ASAP7_75t_L g875 ( 
.A(n_473),
.Y(n_875)
);

CKINVDCx5p33_ASAP7_75t_R g876 ( 
.A(n_158),
.Y(n_876)
);

HB1xp67_ASAP7_75t_L g877 ( 
.A(n_174),
.Y(n_877)
);

CKINVDCx5p33_ASAP7_75t_R g878 ( 
.A(n_449),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_11),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_548),
.Y(n_880)
);

CKINVDCx5p33_ASAP7_75t_R g881 ( 
.A(n_398),
.Y(n_881)
);

CKINVDCx5p33_ASAP7_75t_R g882 ( 
.A(n_30),
.Y(n_882)
);

INVx1_ASAP7_75t_SL g883 ( 
.A(n_105),
.Y(n_883)
);

CKINVDCx5p33_ASAP7_75t_R g884 ( 
.A(n_497),
.Y(n_884)
);

INVx2_ASAP7_75t_L g885 ( 
.A(n_313),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_1),
.Y(n_886)
);

INVx2_ASAP7_75t_L g887 ( 
.A(n_44),
.Y(n_887)
);

CKINVDCx5p33_ASAP7_75t_R g888 ( 
.A(n_620),
.Y(n_888)
);

CKINVDCx5p33_ASAP7_75t_R g889 ( 
.A(n_265),
.Y(n_889)
);

CKINVDCx20_ASAP7_75t_R g890 ( 
.A(n_106),
.Y(n_890)
);

CKINVDCx5p33_ASAP7_75t_R g891 ( 
.A(n_89),
.Y(n_891)
);

INVx2_ASAP7_75t_L g892 ( 
.A(n_568),
.Y(n_892)
);

CKINVDCx5p33_ASAP7_75t_R g893 ( 
.A(n_338),
.Y(n_893)
);

CKINVDCx20_ASAP7_75t_R g894 ( 
.A(n_67),
.Y(n_894)
);

INVx1_ASAP7_75t_L g895 ( 
.A(n_587),
.Y(n_895)
);

INVx1_ASAP7_75t_L g896 ( 
.A(n_665),
.Y(n_896)
);

CKINVDCx5p33_ASAP7_75t_R g897 ( 
.A(n_370),
.Y(n_897)
);

CKINVDCx5p33_ASAP7_75t_R g898 ( 
.A(n_663),
.Y(n_898)
);

CKINVDCx5p33_ASAP7_75t_R g899 ( 
.A(n_278),
.Y(n_899)
);

CKINVDCx5p33_ASAP7_75t_R g900 ( 
.A(n_181),
.Y(n_900)
);

CKINVDCx5p33_ASAP7_75t_R g901 ( 
.A(n_691),
.Y(n_901)
);

CKINVDCx5p33_ASAP7_75t_R g902 ( 
.A(n_619),
.Y(n_902)
);

CKINVDCx5p33_ASAP7_75t_R g903 ( 
.A(n_589),
.Y(n_903)
);

INVx3_ASAP7_75t_L g904 ( 
.A(n_35),
.Y(n_904)
);

INVx1_ASAP7_75t_SL g905 ( 
.A(n_51),
.Y(n_905)
);

CKINVDCx5p33_ASAP7_75t_R g906 ( 
.A(n_343),
.Y(n_906)
);

INVx1_ASAP7_75t_L g907 ( 
.A(n_99),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_285),
.Y(n_908)
);

CKINVDCx5p33_ASAP7_75t_R g909 ( 
.A(n_119),
.Y(n_909)
);

CKINVDCx5p33_ASAP7_75t_R g910 ( 
.A(n_678),
.Y(n_910)
);

CKINVDCx5p33_ASAP7_75t_R g911 ( 
.A(n_22),
.Y(n_911)
);

CKINVDCx5p33_ASAP7_75t_R g912 ( 
.A(n_67),
.Y(n_912)
);

INVx1_ASAP7_75t_L g913 ( 
.A(n_611),
.Y(n_913)
);

INVx1_ASAP7_75t_L g914 ( 
.A(n_37),
.Y(n_914)
);

CKINVDCx20_ASAP7_75t_R g915 ( 
.A(n_376),
.Y(n_915)
);

CKINVDCx5p33_ASAP7_75t_R g916 ( 
.A(n_300),
.Y(n_916)
);

CKINVDCx5p33_ASAP7_75t_R g917 ( 
.A(n_290),
.Y(n_917)
);

CKINVDCx20_ASAP7_75t_R g918 ( 
.A(n_42),
.Y(n_918)
);

CKINVDCx5p33_ASAP7_75t_R g919 ( 
.A(n_9),
.Y(n_919)
);

BUFx10_ASAP7_75t_L g920 ( 
.A(n_174),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_242),
.Y(n_921)
);

CKINVDCx5p33_ASAP7_75t_R g922 ( 
.A(n_166),
.Y(n_922)
);

CKINVDCx5p33_ASAP7_75t_R g923 ( 
.A(n_188),
.Y(n_923)
);

BUFx5_ASAP7_75t_L g924 ( 
.A(n_508),
.Y(n_924)
);

CKINVDCx5p33_ASAP7_75t_R g925 ( 
.A(n_485),
.Y(n_925)
);

CKINVDCx20_ASAP7_75t_R g926 ( 
.A(n_351),
.Y(n_926)
);

CKINVDCx20_ASAP7_75t_R g927 ( 
.A(n_646),
.Y(n_927)
);

CKINVDCx5p33_ASAP7_75t_R g928 ( 
.A(n_3),
.Y(n_928)
);

CKINVDCx5p33_ASAP7_75t_R g929 ( 
.A(n_209),
.Y(n_929)
);

CKINVDCx5p33_ASAP7_75t_R g930 ( 
.A(n_579),
.Y(n_930)
);

CKINVDCx5p33_ASAP7_75t_R g931 ( 
.A(n_407),
.Y(n_931)
);

CKINVDCx5p33_ASAP7_75t_R g932 ( 
.A(n_442),
.Y(n_932)
);

INVx2_ASAP7_75t_SL g933 ( 
.A(n_360),
.Y(n_933)
);

BUFx3_ASAP7_75t_L g934 ( 
.A(n_485),
.Y(n_934)
);

CKINVDCx5p33_ASAP7_75t_R g935 ( 
.A(n_368),
.Y(n_935)
);

CKINVDCx5p33_ASAP7_75t_R g936 ( 
.A(n_567),
.Y(n_936)
);

CKINVDCx5p33_ASAP7_75t_R g937 ( 
.A(n_15),
.Y(n_937)
);

INVx2_ASAP7_75t_L g938 ( 
.A(n_251),
.Y(n_938)
);

INVx1_ASAP7_75t_L g939 ( 
.A(n_171),
.Y(n_939)
);

CKINVDCx20_ASAP7_75t_R g940 ( 
.A(n_125),
.Y(n_940)
);

CKINVDCx5p33_ASAP7_75t_R g941 ( 
.A(n_272),
.Y(n_941)
);

INVx2_ASAP7_75t_SL g942 ( 
.A(n_270),
.Y(n_942)
);

CKINVDCx5p33_ASAP7_75t_R g943 ( 
.A(n_573),
.Y(n_943)
);

BUFx3_ASAP7_75t_L g944 ( 
.A(n_80),
.Y(n_944)
);

INVx1_ASAP7_75t_L g945 ( 
.A(n_671),
.Y(n_945)
);

INVx1_ASAP7_75t_SL g946 ( 
.A(n_96),
.Y(n_946)
);

CKINVDCx5p33_ASAP7_75t_R g947 ( 
.A(n_404),
.Y(n_947)
);

CKINVDCx5p33_ASAP7_75t_R g948 ( 
.A(n_107),
.Y(n_948)
);

CKINVDCx5p33_ASAP7_75t_R g949 ( 
.A(n_111),
.Y(n_949)
);

CKINVDCx5p33_ASAP7_75t_R g950 ( 
.A(n_656),
.Y(n_950)
);

CKINVDCx5p33_ASAP7_75t_R g951 ( 
.A(n_115),
.Y(n_951)
);

CKINVDCx5p33_ASAP7_75t_R g952 ( 
.A(n_336),
.Y(n_952)
);

CKINVDCx5p33_ASAP7_75t_R g953 ( 
.A(n_613),
.Y(n_953)
);

INVx1_ASAP7_75t_L g954 ( 
.A(n_385),
.Y(n_954)
);

CKINVDCx20_ASAP7_75t_R g955 ( 
.A(n_527),
.Y(n_955)
);

CKINVDCx5p33_ASAP7_75t_R g956 ( 
.A(n_245),
.Y(n_956)
);

CKINVDCx5p33_ASAP7_75t_R g957 ( 
.A(n_646),
.Y(n_957)
);

CKINVDCx5p33_ASAP7_75t_R g958 ( 
.A(n_397),
.Y(n_958)
);

CKINVDCx16_ASAP7_75t_R g959 ( 
.A(n_416),
.Y(n_959)
);

CKINVDCx5p33_ASAP7_75t_R g960 ( 
.A(n_139),
.Y(n_960)
);

INVxp67_ASAP7_75t_L g961 ( 
.A(n_584),
.Y(n_961)
);

CKINVDCx5p33_ASAP7_75t_R g962 ( 
.A(n_586),
.Y(n_962)
);

CKINVDCx5p33_ASAP7_75t_R g963 ( 
.A(n_142),
.Y(n_963)
);

BUFx3_ASAP7_75t_L g964 ( 
.A(n_351),
.Y(n_964)
);

INVx1_ASAP7_75t_L g965 ( 
.A(n_333),
.Y(n_965)
);

INVx1_ASAP7_75t_L g966 ( 
.A(n_628),
.Y(n_966)
);

INVx1_ASAP7_75t_L g967 ( 
.A(n_364),
.Y(n_967)
);

INVx1_ASAP7_75t_L g968 ( 
.A(n_601),
.Y(n_968)
);

BUFx5_ASAP7_75t_L g969 ( 
.A(n_138),
.Y(n_969)
);

INVx1_ASAP7_75t_L g970 ( 
.A(n_662),
.Y(n_970)
);

INVx2_ASAP7_75t_L g971 ( 
.A(n_247),
.Y(n_971)
);

INVx1_ASAP7_75t_L g972 ( 
.A(n_245),
.Y(n_972)
);

CKINVDCx5p33_ASAP7_75t_R g973 ( 
.A(n_426),
.Y(n_973)
);

BUFx2_ASAP7_75t_L g974 ( 
.A(n_7),
.Y(n_974)
);

CKINVDCx5p33_ASAP7_75t_R g975 ( 
.A(n_119),
.Y(n_975)
);

CKINVDCx5p33_ASAP7_75t_R g976 ( 
.A(n_643),
.Y(n_976)
);

INVx2_ASAP7_75t_L g977 ( 
.A(n_396),
.Y(n_977)
);

CKINVDCx5p33_ASAP7_75t_R g978 ( 
.A(n_262),
.Y(n_978)
);

CKINVDCx5p33_ASAP7_75t_R g979 ( 
.A(n_443),
.Y(n_979)
);

INVx1_ASAP7_75t_L g980 ( 
.A(n_617),
.Y(n_980)
);

CKINVDCx5p33_ASAP7_75t_R g981 ( 
.A(n_57),
.Y(n_981)
);

BUFx10_ASAP7_75t_L g982 ( 
.A(n_163),
.Y(n_982)
);

INVx1_ASAP7_75t_SL g983 ( 
.A(n_467),
.Y(n_983)
);

INVx2_ASAP7_75t_L g984 ( 
.A(n_18),
.Y(n_984)
);

INVx1_ASAP7_75t_L g985 ( 
.A(n_158),
.Y(n_985)
);

CKINVDCx5p33_ASAP7_75t_R g986 ( 
.A(n_575),
.Y(n_986)
);

BUFx3_ASAP7_75t_L g987 ( 
.A(n_405),
.Y(n_987)
);

INVx1_ASAP7_75t_L g988 ( 
.A(n_516),
.Y(n_988)
);

INVx1_ASAP7_75t_L g989 ( 
.A(n_672),
.Y(n_989)
);

INVx2_ASAP7_75t_L g990 ( 
.A(n_194),
.Y(n_990)
);

CKINVDCx5p33_ASAP7_75t_R g991 ( 
.A(n_243),
.Y(n_991)
);

BUFx2_ASAP7_75t_SL g992 ( 
.A(n_679),
.Y(n_992)
);

CKINVDCx5p33_ASAP7_75t_R g993 ( 
.A(n_32),
.Y(n_993)
);

CKINVDCx20_ASAP7_75t_R g994 ( 
.A(n_557),
.Y(n_994)
);

CKINVDCx20_ASAP7_75t_R g995 ( 
.A(n_536),
.Y(n_995)
);

INVx1_ASAP7_75t_L g996 ( 
.A(n_57),
.Y(n_996)
);

CKINVDCx20_ASAP7_75t_R g997 ( 
.A(n_236),
.Y(n_997)
);

INVx1_ASAP7_75t_L g998 ( 
.A(n_694),
.Y(n_998)
);

CKINVDCx5p33_ASAP7_75t_R g999 ( 
.A(n_559),
.Y(n_999)
);

CKINVDCx5p33_ASAP7_75t_R g1000 ( 
.A(n_597),
.Y(n_1000)
);

CKINVDCx20_ASAP7_75t_R g1001 ( 
.A(n_332),
.Y(n_1001)
);

CKINVDCx5p33_ASAP7_75t_R g1002 ( 
.A(n_514),
.Y(n_1002)
);

CKINVDCx5p33_ASAP7_75t_R g1003 ( 
.A(n_667),
.Y(n_1003)
);

CKINVDCx16_ASAP7_75t_R g1004 ( 
.A(n_688),
.Y(n_1004)
);

CKINVDCx5p33_ASAP7_75t_R g1005 ( 
.A(n_204),
.Y(n_1005)
);

CKINVDCx5p33_ASAP7_75t_R g1006 ( 
.A(n_227),
.Y(n_1006)
);

CKINVDCx5p33_ASAP7_75t_R g1007 ( 
.A(n_669),
.Y(n_1007)
);

CKINVDCx5p33_ASAP7_75t_R g1008 ( 
.A(n_324),
.Y(n_1008)
);

INVx1_ASAP7_75t_L g1009 ( 
.A(n_150),
.Y(n_1009)
);

CKINVDCx5p33_ASAP7_75t_R g1010 ( 
.A(n_648),
.Y(n_1010)
);

CKINVDCx5p33_ASAP7_75t_R g1011 ( 
.A(n_336),
.Y(n_1011)
);

CKINVDCx5p33_ASAP7_75t_R g1012 ( 
.A(n_323),
.Y(n_1012)
);

CKINVDCx20_ASAP7_75t_R g1013 ( 
.A(n_562),
.Y(n_1013)
);

CKINVDCx5p33_ASAP7_75t_R g1014 ( 
.A(n_148),
.Y(n_1014)
);

CKINVDCx5p33_ASAP7_75t_R g1015 ( 
.A(n_631),
.Y(n_1015)
);

INVx1_ASAP7_75t_L g1016 ( 
.A(n_608),
.Y(n_1016)
);

CKINVDCx20_ASAP7_75t_R g1017 ( 
.A(n_406),
.Y(n_1017)
);

CKINVDCx5p33_ASAP7_75t_R g1018 ( 
.A(n_233),
.Y(n_1018)
);

CKINVDCx5p33_ASAP7_75t_R g1019 ( 
.A(n_315),
.Y(n_1019)
);

CKINVDCx20_ASAP7_75t_R g1020 ( 
.A(n_411),
.Y(n_1020)
);

BUFx3_ASAP7_75t_L g1021 ( 
.A(n_611),
.Y(n_1021)
);

INVx1_ASAP7_75t_L g1022 ( 
.A(n_101),
.Y(n_1022)
);

CKINVDCx5p33_ASAP7_75t_R g1023 ( 
.A(n_300),
.Y(n_1023)
);

INVxp67_ASAP7_75t_L g1024 ( 
.A(n_70),
.Y(n_1024)
);

INVx1_ASAP7_75t_L g1025 ( 
.A(n_74),
.Y(n_1025)
);

INVx1_ASAP7_75t_L g1026 ( 
.A(n_630),
.Y(n_1026)
);

CKINVDCx5p33_ASAP7_75t_R g1027 ( 
.A(n_371),
.Y(n_1027)
);

CKINVDCx5p33_ASAP7_75t_R g1028 ( 
.A(n_306),
.Y(n_1028)
);

INVx1_ASAP7_75t_L g1029 ( 
.A(n_411),
.Y(n_1029)
);

INVx1_ASAP7_75t_L g1030 ( 
.A(n_94),
.Y(n_1030)
);

CKINVDCx5p33_ASAP7_75t_R g1031 ( 
.A(n_609),
.Y(n_1031)
);

CKINVDCx5p33_ASAP7_75t_R g1032 ( 
.A(n_434),
.Y(n_1032)
);

INVx1_ASAP7_75t_L g1033 ( 
.A(n_621),
.Y(n_1033)
);

CKINVDCx5p33_ASAP7_75t_R g1034 ( 
.A(n_448),
.Y(n_1034)
);

INVx1_ASAP7_75t_L g1035 ( 
.A(n_714),
.Y(n_1035)
);

CKINVDCx5p33_ASAP7_75t_R g1036 ( 
.A(n_754),
.Y(n_1036)
);

INVx1_ASAP7_75t_L g1037 ( 
.A(n_714),
.Y(n_1037)
);

CKINVDCx5p33_ASAP7_75t_R g1038 ( 
.A(n_729),
.Y(n_1038)
);

INVx1_ASAP7_75t_L g1039 ( 
.A(n_714),
.Y(n_1039)
);

CKINVDCx5p33_ASAP7_75t_R g1040 ( 
.A(n_841),
.Y(n_1040)
);

CKINVDCx5p33_ASAP7_75t_R g1041 ( 
.A(n_867),
.Y(n_1041)
);

INVx1_ASAP7_75t_L g1042 ( 
.A(n_714),
.Y(n_1042)
);

INVx2_ASAP7_75t_L g1043 ( 
.A(n_714),
.Y(n_1043)
);

INVx1_ASAP7_75t_L g1044 ( 
.A(n_714),
.Y(n_1044)
);

INVxp33_ASAP7_75t_L g1045 ( 
.A(n_717),
.Y(n_1045)
);

BUFx2_ASAP7_75t_L g1046 ( 
.A(n_974),
.Y(n_1046)
);

INVx1_ASAP7_75t_L g1047 ( 
.A(n_714),
.Y(n_1047)
);

CKINVDCx5p33_ASAP7_75t_R g1048 ( 
.A(n_959),
.Y(n_1048)
);

CKINVDCx5p33_ASAP7_75t_R g1049 ( 
.A(n_1004),
.Y(n_1049)
);

INVxp67_ASAP7_75t_L g1050 ( 
.A(n_726),
.Y(n_1050)
);

INVxp67_ASAP7_75t_L g1051 ( 
.A(n_761),
.Y(n_1051)
);

CKINVDCx5p33_ASAP7_75t_R g1052 ( 
.A(n_769),
.Y(n_1052)
);

HB1xp67_ASAP7_75t_L g1053 ( 
.A(n_778),
.Y(n_1053)
);

INVx1_ASAP7_75t_L g1054 ( 
.A(n_714),
.Y(n_1054)
);

INVx1_ASAP7_75t_L g1055 ( 
.A(n_924),
.Y(n_1055)
);

CKINVDCx5p33_ASAP7_75t_R g1056 ( 
.A(n_773),
.Y(n_1056)
);

CKINVDCx5p33_ASAP7_75t_R g1057 ( 
.A(n_774),
.Y(n_1057)
);

INVx1_ASAP7_75t_L g1058 ( 
.A(n_924),
.Y(n_1058)
);

INVx1_ASAP7_75t_L g1059 ( 
.A(n_924),
.Y(n_1059)
);

CKINVDCx5p33_ASAP7_75t_R g1060 ( 
.A(n_776),
.Y(n_1060)
);

INVx1_ASAP7_75t_L g1061 ( 
.A(n_924),
.Y(n_1061)
);

INVx1_ASAP7_75t_L g1062 ( 
.A(n_924),
.Y(n_1062)
);

INVx1_ASAP7_75t_L g1063 ( 
.A(n_924),
.Y(n_1063)
);

INVx1_ASAP7_75t_L g1064 ( 
.A(n_924),
.Y(n_1064)
);

INVx1_ASAP7_75t_L g1065 ( 
.A(n_924),
.Y(n_1065)
);

INVx1_ASAP7_75t_L g1066 ( 
.A(n_969),
.Y(n_1066)
);

INVx1_ASAP7_75t_L g1067 ( 
.A(n_969),
.Y(n_1067)
);

INVx1_ASAP7_75t_L g1068 ( 
.A(n_969),
.Y(n_1068)
);

CKINVDCx20_ASAP7_75t_R g1069 ( 
.A(n_721),
.Y(n_1069)
);

INVx1_ASAP7_75t_L g1070 ( 
.A(n_969),
.Y(n_1070)
);

CKINVDCx5p33_ASAP7_75t_R g1071 ( 
.A(n_782),
.Y(n_1071)
);

INVx1_ASAP7_75t_SL g1072 ( 
.A(n_781),
.Y(n_1072)
);

CKINVDCx16_ASAP7_75t_R g1073 ( 
.A(n_703),
.Y(n_1073)
);

CKINVDCx5p33_ASAP7_75t_R g1074 ( 
.A(n_783),
.Y(n_1074)
);

INVx1_ASAP7_75t_L g1075 ( 
.A(n_969),
.Y(n_1075)
);

INVx1_ASAP7_75t_L g1076 ( 
.A(n_969),
.Y(n_1076)
);

INVx1_ASAP7_75t_L g1077 ( 
.A(n_969),
.Y(n_1077)
);

CKINVDCx5p33_ASAP7_75t_R g1078 ( 
.A(n_784),
.Y(n_1078)
);

CKINVDCx20_ASAP7_75t_R g1079 ( 
.A(n_736),
.Y(n_1079)
);

CKINVDCx5p33_ASAP7_75t_R g1080 ( 
.A(n_785),
.Y(n_1080)
);

CKINVDCx16_ASAP7_75t_R g1081 ( 
.A(n_703),
.Y(n_1081)
);

INVx1_ASAP7_75t_L g1082 ( 
.A(n_969),
.Y(n_1082)
);

CKINVDCx20_ASAP7_75t_R g1083 ( 
.A(n_757),
.Y(n_1083)
);

INVx1_ASAP7_75t_L g1084 ( 
.A(n_904),
.Y(n_1084)
);

INVx1_ASAP7_75t_SL g1085 ( 
.A(n_890),
.Y(n_1085)
);

CKINVDCx5p33_ASAP7_75t_R g1086 ( 
.A(n_789),
.Y(n_1086)
);

INVx1_ASAP7_75t_L g1087 ( 
.A(n_904),
.Y(n_1087)
);

CKINVDCx20_ASAP7_75t_R g1088 ( 
.A(n_770),
.Y(n_1088)
);

CKINVDCx16_ASAP7_75t_R g1089 ( 
.A(n_703),
.Y(n_1089)
);

CKINVDCx5p33_ASAP7_75t_R g1090 ( 
.A(n_790),
.Y(n_1090)
);

INVxp67_ASAP7_75t_L g1091 ( 
.A(n_805),
.Y(n_1091)
);

INVx1_ASAP7_75t_L g1092 ( 
.A(n_904),
.Y(n_1092)
);

BUFx3_ASAP7_75t_L g1093 ( 
.A(n_944),
.Y(n_1093)
);

INVxp33_ASAP7_75t_SL g1094 ( 
.A(n_877),
.Y(n_1094)
);

CKINVDCx5p33_ASAP7_75t_R g1095 ( 
.A(n_795),
.Y(n_1095)
);

CKINVDCx5p33_ASAP7_75t_R g1096 ( 
.A(n_796),
.Y(n_1096)
);

CKINVDCx5p33_ASAP7_75t_R g1097 ( 
.A(n_798),
.Y(n_1097)
);

CKINVDCx5p33_ASAP7_75t_R g1098 ( 
.A(n_799),
.Y(n_1098)
);

INVx1_ASAP7_75t_L g1099 ( 
.A(n_750),
.Y(n_1099)
);

CKINVDCx5p33_ASAP7_75t_R g1100 ( 
.A(n_800),
.Y(n_1100)
);

INVx1_ASAP7_75t_L g1101 ( 
.A(n_771),
.Y(n_1101)
);

CKINVDCx20_ASAP7_75t_R g1102 ( 
.A(n_775),
.Y(n_1102)
);

CKINVDCx5p33_ASAP7_75t_R g1103 ( 
.A(n_801),
.Y(n_1103)
);

CKINVDCx20_ASAP7_75t_R g1104 ( 
.A(n_788),
.Y(n_1104)
);

INVx1_ASAP7_75t_L g1105 ( 
.A(n_803),
.Y(n_1105)
);

INVx1_ASAP7_75t_L g1106 ( 
.A(n_804),
.Y(n_1106)
);

INVx1_ASAP7_75t_L g1107 ( 
.A(n_827),
.Y(n_1107)
);

INVx1_ASAP7_75t_L g1108 ( 
.A(n_856),
.Y(n_1108)
);

CKINVDCx5p33_ASAP7_75t_R g1109 ( 
.A(n_806),
.Y(n_1109)
);

CKINVDCx5p33_ASAP7_75t_R g1110 ( 
.A(n_807),
.Y(n_1110)
);

INVx1_ASAP7_75t_L g1111 ( 
.A(n_866),
.Y(n_1111)
);

CKINVDCx5p33_ASAP7_75t_R g1112 ( 
.A(n_811),
.Y(n_1112)
);

INVxp67_ASAP7_75t_L g1113 ( 
.A(n_879),
.Y(n_1113)
);

CKINVDCx5p33_ASAP7_75t_R g1114 ( 
.A(n_813),
.Y(n_1114)
);

INVx1_ASAP7_75t_L g1115 ( 
.A(n_886),
.Y(n_1115)
);

CKINVDCx5p33_ASAP7_75t_R g1116 ( 
.A(n_816),
.Y(n_1116)
);

CKINVDCx5p33_ASAP7_75t_R g1117 ( 
.A(n_817),
.Y(n_1117)
);

CKINVDCx20_ASAP7_75t_R g1118 ( 
.A(n_831),
.Y(n_1118)
);

CKINVDCx5p33_ASAP7_75t_R g1119 ( 
.A(n_820),
.Y(n_1119)
);

NOR2xp33_ASAP7_75t_L g1120 ( 
.A(n_944),
.B(n_0),
.Y(n_1120)
);

CKINVDCx5p33_ASAP7_75t_R g1121 ( 
.A(n_822),
.Y(n_1121)
);

CKINVDCx5p33_ASAP7_75t_R g1122 ( 
.A(n_825),
.Y(n_1122)
);

BUFx3_ASAP7_75t_L g1123 ( 
.A(n_791),
.Y(n_1123)
);

BUFx3_ASAP7_75t_L g1124 ( 
.A(n_791),
.Y(n_1124)
);

INVx1_ASAP7_75t_L g1125 ( 
.A(n_907),
.Y(n_1125)
);

CKINVDCx20_ASAP7_75t_R g1126 ( 
.A(n_837),
.Y(n_1126)
);

INVx1_ASAP7_75t_L g1127 ( 
.A(n_914),
.Y(n_1127)
);

CKINVDCx14_ASAP7_75t_R g1128 ( 
.A(n_772),
.Y(n_1128)
);

INVx2_ASAP7_75t_L g1129 ( 
.A(n_710),
.Y(n_1129)
);

CKINVDCx5p33_ASAP7_75t_R g1130 ( 
.A(n_777),
.Y(n_1130)
);

BUFx6f_ASAP7_75t_L g1131 ( 
.A(n_710),
.Y(n_1131)
);

INVx1_ASAP7_75t_L g1132 ( 
.A(n_996),
.Y(n_1132)
);

INVx1_ASAP7_75t_L g1133 ( 
.A(n_1022),
.Y(n_1133)
);

CKINVDCx20_ASAP7_75t_R g1134 ( 
.A(n_915),
.Y(n_1134)
);

INVx1_ASAP7_75t_L g1135 ( 
.A(n_1025),
.Y(n_1135)
);

HB1xp67_ASAP7_75t_L g1136 ( 
.A(n_780),
.Y(n_1136)
);

CKINVDCx5p33_ASAP7_75t_R g1137 ( 
.A(n_797),
.Y(n_1137)
);

CKINVDCx20_ASAP7_75t_R g1138 ( 
.A(n_926),
.Y(n_1138)
);

INVx1_ASAP7_75t_L g1139 ( 
.A(n_1030),
.Y(n_1139)
);

CKINVDCx20_ASAP7_75t_R g1140 ( 
.A(n_927),
.Y(n_1140)
);

INVx1_ASAP7_75t_L g1141 ( 
.A(n_814),
.Y(n_1141)
);

INVxp67_ASAP7_75t_L g1142 ( 
.A(n_772),
.Y(n_1142)
);

INVxp67_ASAP7_75t_L g1143 ( 
.A(n_772),
.Y(n_1143)
);

INVx1_ASAP7_75t_L g1144 ( 
.A(n_814),
.Y(n_1144)
);

CKINVDCx5p33_ASAP7_75t_R g1145 ( 
.A(n_809),
.Y(n_1145)
);

CKINVDCx5p33_ASAP7_75t_R g1146 ( 
.A(n_819),
.Y(n_1146)
);

INVx1_ASAP7_75t_L g1147 ( 
.A(n_818),
.Y(n_1147)
);

INVx1_ASAP7_75t_L g1148 ( 
.A(n_818),
.Y(n_1148)
);

CKINVDCx5p33_ASAP7_75t_R g1149 ( 
.A(n_824),
.Y(n_1149)
);

CKINVDCx5p33_ASAP7_75t_R g1150 ( 
.A(n_832),
.Y(n_1150)
);

INVx1_ASAP7_75t_L g1151 ( 
.A(n_850),
.Y(n_1151)
);

INVx1_ASAP7_75t_L g1152 ( 
.A(n_850),
.Y(n_1152)
);

INVx1_ASAP7_75t_L g1153 ( 
.A(n_934),
.Y(n_1153)
);

CKINVDCx5p33_ASAP7_75t_R g1154 ( 
.A(n_838),
.Y(n_1154)
);

INVx1_ASAP7_75t_L g1155 ( 
.A(n_934),
.Y(n_1155)
);

CKINVDCx5p33_ASAP7_75t_R g1156 ( 
.A(n_843),
.Y(n_1156)
);

BUFx2_ASAP7_75t_L g1157 ( 
.A(n_711),
.Y(n_1157)
);

INVx1_ASAP7_75t_L g1158 ( 
.A(n_964),
.Y(n_1158)
);

BUFx6f_ASAP7_75t_L g1159 ( 
.A(n_710),
.Y(n_1159)
);

INVx1_ASAP7_75t_L g1160 ( 
.A(n_964),
.Y(n_1160)
);

INVx1_ASAP7_75t_L g1161 ( 
.A(n_987),
.Y(n_1161)
);

CKINVDCx5p33_ASAP7_75t_R g1162 ( 
.A(n_855),
.Y(n_1162)
);

INVxp67_ASAP7_75t_SL g1163 ( 
.A(n_710),
.Y(n_1163)
);

CKINVDCx5p33_ASAP7_75t_R g1164 ( 
.A(n_826),
.Y(n_1164)
);

INVx2_ASAP7_75t_L g1165 ( 
.A(n_710),
.Y(n_1165)
);

INVx2_ASAP7_75t_L g1166 ( 
.A(n_861),
.Y(n_1166)
);

INVx1_ASAP7_75t_L g1167 ( 
.A(n_987),
.Y(n_1167)
);

CKINVDCx5p33_ASAP7_75t_R g1168 ( 
.A(n_829),
.Y(n_1168)
);

BUFx10_ASAP7_75t_L g1169 ( 
.A(n_861),
.Y(n_1169)
);

INVx1_ASAP7_75t_L g1170 ( 
.A(n_1021),
.Y(n_1170)
);

INVx1_ASAP7_75t_SL g1171 ( 
.A(n_894),
.Y(n_1171)
);

INVx1_ASAP7_75t_L g1172 ( 
.A(n_1021),
.Y(n_1172)
);

NOR2xp67_ASAP7_75t_L g1173 ( 
.A(n_961),
.B(n_0),
.Y(n_1173)
);

INVx1_ASAP7_75t_L g1174 ( 
.A(n_861),
.Y(n_1174)
);

CKINVDCx5p33_ASAP7_75t_R g1175 ( 
.A(n_830),
.Y(n_1175)
);

CKINVDCx5p33_ASAP7_75t_R g1176 ( 
.A(n_833),
.Y(n_1176)
);

BUFx3_ASAP7_75t_L g1177 ( 
.A(n_861),
.Y(n_1177)
);

CKINVDCx5p33_ASAP7_75t_R g1178 ( 
.A(n_834),
.Y(n_1178)
);

INVx1_ASAP7_75t_L g1179 ( 
.A(n_861),
.Y(n_1179)
);

INVx1_ASAP7_75t_L g1180 ( 
.A(n_865),
.Y(n_1180)
);

INVx2_ASAP7_75t_L g1181 ( 
.A(n_865),
.Y(n_1181)
);

BUFx2_ASAP7_75t_L g1182 ( 
.A(n_711),
.Y(n_1182)
);

INVx2_ASAP7_75t_L g1183 ( 
.A(n_865),
.Y(n_1183)
);

INVx1_ASAP7_75t_L g1184 ( 
.A(n_865),
.Y(n_1184)
);

INVx1_ASAP7_75t_L g1185 ( 
.A(n_865),
.Y(n_1185)
);

BUFx6f_ASAP7_75t_L g1186 ( 
.A(n_873),
.Y(n_1186)
);

INVx1_ASAP7_75t_L g1187 ( 
.A(n_873),
.Y(n_1187)
);

INVxp33_ASAP7_75t_SL g1188 ( 
.A(n_713),
.Y(n_1188)
);

HB1xp67_ASAP7_75t_L g1189 ( 
.A(n_713),
.Y(n_1189)
);

CKINVDCx5p33_ASAP7_75t_R g1190 ( 
.A(n_839),
.Y(n_1190)
);

INVx1_ASAP7_75t_L g1191 ( 
.A(n_873),
.Y(n_1191)
);

INVx1_ASAP7_75t_L g1192 ( 
.A(n_873),
.Y(n_1192)
);

INVx1_ASAP7_75t_L g1193 ( 
.A(n_873),
.Y(n_1193)
);

INVx2_ASAP7_75t_L g1194 ( 
.A(n_715),
.Y(n_1194)
);

CKINVDCx5p33_ASAP7_75t_R g1195 ( 
.A(n_842),
.Y(n_1195)
);

INVx1_ASAP7_75t_L g1196 ( 
.A(n_715),
.Y(n_1196)
);

INVx1_ASAP7_75t_L g1197 ( 
.A(n_887),
.Y(n_1197)
);

INVx2_ASAP7_75t_SL g1198 ( 
.A(n_812),
.Y(n_1198)
);

INVx1_ASAP7_75t_L g1199 ( 
.A(n_887),
.Y(n_1199)
);

CKINVDCx5p33_ASAP7_75t_R g1200 ( 
.A(n_857),
.Y(n_1200)
);

CKINVDCx5p33_ASAP7_75t_R g1201 ( 
.A(n_860),
.Y(n_1201)
);

INVx1_ASAP7_75t_L g1202 ( 
.A(n_984),
.Y(n_1202)
);

INVx2_ASAP7_75t_L g1203 ( 
.A(n_984),
.Y(n_1203)
);

CKINVDCx5p33_ASAP7_75t_R g1204 ( 
.A(n_868),
.Y(n_1204)
);

INVx1_ASAP7_75t_L g1205 ( 
.A(n_708),
.Y(n_1205)
);

BUFx3_ASAP7_75t_L g1206 ( 
.A(n_812),
.Y(n_1206)
);

BUFx3_ASAP7_75t_L g1207 ( 
.A(n_812),
.Y(n_1207)
);

BUFx6f_ASAP7_75t_L g1208 ( 
.A(n_727),
.Y(n_1208)
);

INVx1_ASAP7_75t_L g1209 ( 
.A(n_718),
.Y(n_1209)
);

BUFx2_ASAP7_75t_L g1210 ( 
.A(n_716),
.Y(n_1210)
);

CKINVDCx5p33_ASAP7_75t_R g1211 ( 
.A(n_869),
.Y(n_1211)
);

INVx1_ASAP7_75t_L g1212 ( 
.A(n_723),
.Y(n_1212)
);

INVx1_ASAP7_75t_L g1213 ( 
.A(n_724),
.Y(n_1213)
);

INVx1_ASAP7_75t_L g1214 ( 
.A(n_725),
.Y(n_1214)
);

INVx1_ASAP7_75t_L g1215 ( 
.A(n_735),
.Y(n_1215)
);

INVx1_ASAP7_75t_L g1216 ( 
.A(n_738),
.Y(n_1216)
);

INVx2_ASAP7_75t_L g1217 ( 
.A(n_727),
.Y(n_1217)
);

CKINVDCx5p33_ASAP7_75t_R g1218 ( 
.A(n_882),
.Y(n_1218)
);

INVxp67_ASAP7_75t_SL g1219 ( 
.A(n_1024),
.Y(n_1219)
);

INVx1_ASAP7_75t_L g1220 ( 
.A(n_739),
.Y(n_1220)
);

CKINVDCx5p33_ASAP7_75t_R g1221 ( 
.A(n_891),
.Y(n_1221)
);

BUFx6f_ASAP7_75t_L g1222 ( 
.A(n_763),
.Y(n_1222)
);

CKINVDCx5p33_ASAP7_75t_R g1223 ( 
.A(n_911),
.Y(n_1223)
);

CKINVDCx5p33_ASAP7_75t_R g1224 ( 
.A(n_912),
.Y(n_1224)
);

INVx1_ASAP7_75t_L g1225 ( 
.A(n_744),
.Y(n_1225)
);

NAND2xp5_ASAP7_75t_L g1226 ( 
.A(n_719),
.B(n_1),
.Y(n_1226)
);

BUFx2_ASAP7_75t_L g1227 ( 
.A(n_716),
.Y(n_1227)
);

INVx1_ASAP7_75t_L g1228 ( 
.A(n_759),
.Y(n_1228)
);

INVx1_ASAP7_75t_L g1229 ( 
.A(n_762),
.Y(n_1229)
);

CKINVDCx5p33_ASAP7_75t_R g1230 ( 
.A(n_919),
.Y(n_1230)
);

INVxp67_ASAP7_75t_L g1231 ( 
.A(n_823),
.Y(n_1231)
);

INVx1_ASAP7_75t_L g1232 ( 
.A(n_768),
.Y(n_1232)
);

INVx1_ASAP7_75t_L g1233 ( 
.A(n_779),
.Y(n_1233)
);

CKINVDCx5p33_ASAP7_75t_R g1234 ( 
.A(n_928),
.Y(n_1234)
);

INVx2_ASAP7_75t_L g1235 ( 
.A(n_763),
.Y(n_1235)
);

CKINVDCx5p33_ASAP7_75t_R g1236 ( 
.A(n_937),
.Y(n_1236)
);

NOR2xp67_ASAP7_75t_L g1237 ( 
.A(n_719),
.B(n_1),
.Y(n_1237)
);

OR2x2_ASAP7_75t_L g1238 ( 
.A(n_883),
.B(n_3),
.Y(n_1238)
);

INVx1_ASAP7_75t_L g1239 ( 
.A(n_786),
.Y(n_1239)
);

INVx2_ASAP7_75t_L g1240 ( 
.A(n_792),
.Y(n_1240)
);

CKINVDCx5p33_ASAP7_75t_R g1241 ( 
.A(n_846),
.Y(n_1241)
);

OR2x2_ASAP7_75t_L g1242 ( 
.A(n_905),
.B(n_3),
.Y(n_1242)
);

INVx1_ASAP7_75t_L g1243 ( 
.A(n_787),
.Y(n_1243)
);

INVx1_ASAP7_75t_L g1244 ( 
.A(n_793),
.Y(n_1244)
);

INVx1_ASAP7_75t_L g1245 ( 
.A(n_794),
.Y(n_1245)
);

INVx1_ASAP7_75t_L g1246 ( 
.A(n_802),
.Y(n_1246)
);

BUFx2_ASAP7_75t_L g1247 ( 
.A(n_730),
.Y(n_1247)
);

INVx1_ASAP7_75t_L g1248 ( 
.A(n_815),
.Y(n_1248)
);

INVx1_ASAP7_75t_L g1249 ( 
.A(n_828),
.Y(n_1249)
);

INVx1_ASAP7_75t_L g1250 ( 
.A(n_835),
.Y(n_1250)
);

CKINVDCx5p33_ASAP7_75t_R g1251 ( 
.A(n_847),
.Y(n_1251)
);

INVx1_ASAP7_75t_L g1252 ( 
.A(n_840),
.Y(n_1252)
);

CKINVDCx5p33_ASAP7_75t_R g1253 ( 
.A(n_851),
.Y(n_1253)
);

INVx1_ASAP7_75t_L g1254 ( 
.A(n_845),
.Y(n_1254)
);

INVx1_ASAP7_75t_L g1255 ( 
.A(n_848),
.Y(n_1255)
);

CKINVDCx5p33_ASAP7_75t_R g1256 ( 
.A(n_853),
.Y(n_1256)
);

INVxp67_ASAP7_75t_L g1257 ( 
.A(n_823),
.Y(n_1257)
);

INVx2_ASAP7_75t_L g1258 ( 
.A(n_792),
.Y(n_1258)
);

CKINVDCx5p33_ASAP7_75t_R g1259 ( 
.A(n_854),
.Y(n_1259)
);

CKINVDCx5p33_ASAP7_75t_R g1260 ( 
.A(n_862),
.Y(n_1260)
);

INVx1_ASAP7_75t_L g1261 ( 
.A(n_852),
.Y(n_1261)
);

INVx1_ASAP7_75t_L g1262 ( 
.A(n_858),
.Y(n_1262)
);

BUFx6f_ASAP7_75t_L g1263 ( 
.A(n_810),
.Y(n_1263)
);

INVx1_ASAP7_75t_L g1264 ( 
.A(n_859),
.Y(n_1264)
);

INVx1_ASAP7_75t_SL g1265 ( 
.A(n_918),
.Y(n_1265)
);

INVxp67_ASAP7_75t_L g1266 ( 
.A(n_823),
.Y(n_1266)
);

INVx1_ASAP7_75t_L g1267 ( 
.A(n_874),
.Y(n_1267)
);

INVx1_ASAP7_75t_L g1268 ( 
.A(n_875),
.Y(n_1268)
);

INVx1_ASAP7_75t_L g1269 ( 
.A(n_880),
.Y(n_1269)
);

CKINVDCx5p33_ASAP7_75t_R g1270 ( 
.A(n_863),
.Y(n_1270)
);

INVx1_ASAP7_75t_L g1271 ( 
.A(n_895),
.Y(n_1271)
);

CKINVDCx20_ASAP7_75t_R g1272 ( 
.A(n_940),
.Y(n_1272)
);

CKINVDCx5p33_ASAP7_75t_R g1273 ( 
.A(n_864),
.Y(n_1273)
);

CKINVDCx20_ASAP7_75t_R g1274 ( 
.A(n_955),
.Y(n_1274)
);

BUFx6f_ASAP7_75t_L g1275 ( 
.A(n_810),
.Y(n_1275)
);

CKINVDCx5p33_ASAP7_75t_R g1276 ( 
.A(n_871),
.Y(n_1276)
);

INVx1_ASAP7_75t_L g1277 ( 
.A(n_896),
.Y(n_1277)
);

INVxp33_ASAP7_75t_L g1278 ( 
.A(n_908),
.Y(n_1278)
);

INVx1_ASAP7_75t_L g1279 ( 
.A(n_913),
.Y(n_1279)
);

BUFx10_ASAP7_75t_L g1280 ( 
.A(n_730),
.Y(n_1280)
);

CKINVDCx5p33_ASAP7_75t_R g1281 ( 
.A(n_872),
.Y(n_1281)
);

NOR2xp67_ASAP7_75t_L g1282 ( 
.A(n_933),
.B(n_2),
.Y(n_1282)
);

INVx1_ASAP7_75t_L g1283 ( 
.A(n_921),
.Y(n_1283)
);

INVx1_ASAP7_75t_L g1284 ( 
.A(n_939),
.Y(n_1284)
);

INVx1_ASAP7_75t_L g1285 ( 
.A(n_945),
.Y(n_1285)
);

CKINVDCx5p33_ASAP7_75t_R g1286 ( 
.A(n_876),
.Y(n_1286)
);

INVx1_ASAP7_75t_L g1287 ( 
.A(n_954),
.Y(n_1287)
);

CKINVDCx5p33_ASAP7_75t_R g1288 ( 
.A(n_878),
.Y(n_1288)
);

CKINVDCx5p33_ASAP7_75t_R g1289 ( 
.A(n_881),
.Y(n_1289)
);

CKINVDCx5p33_ASAP7_75t_R g1290 ( 
.A(n_884),
.Y(n_1290)
);

INVx1_ASAP7_75t_L g1291 ( 
.A(n_965),
.Y(n_1291)
);

CKINVDCx5p33_ASAP7_75t_R g1292 ( 
.A(n_888),
.Y(n_1292)
);

CKINVDCx16_ASAP7_75t_R g1293 ( 
.A(n_920),
.Y(n_1293)
);

INVx1_ASAP7_75t_L g1294 ( 
.A(n_966),
.Y(n_1294)
);

INVx1_ASAP7_75t_L g1295 ( 
.A(n_967),
.Y(n_1295)
);

CKINVDCx20_ASAP7_75t_R g1296 ( 
.A(n_994),
.Y(n_1296)
);

INVx1_ASAP7_75t_L g1297 ( 
.A(n_968),
.Y(n_1297)
);

CKINVDCx20_ASAP7_75t_R g1298 ( 
.A(n_995),
.Y(n_1298)
);

BUFx8_ASAP7_75t_SL g1299 ( 
.A(n_997),
.Y(n_1299)
);

INVx1_ASAP7_75t_L g1300 ( 
.A(n_970),
.Y(n_1300)
);

CKINVDCx5p33_ASAP7_75t_R g1301 ( 
.A(n_889),
.Y(n_1301)
);

INVx1_ASAP7_75t_L g1302 ( 
.A(n_972),
.Y(n_1302)
);

INVx1_ASAP7_75t_L g1303 ( 
.A(n_980),
.Y(n_1303)
);

BUFx3_ASAP7_75t_L g1304 ( 
.A(n_920),
.Y(n_1304)
);

INVx2_ASAP7_75t_L g1305 ( 
.A(n_870),
.Y(n_1305)
);

INVx1_ASAP7_75t_L g1306 ( 
.A(n_985),
.Y(n_1306)
);

HB1xp67_ASAP7_75t_L g1307 ( 
.A(n_743),
.Y(n_1307)
);

INVxp67_ASAP7_75t_L g1308 ( 
.A(n_920),
.Y(n_1308)
);

INVx1_ASAP7_75t_L g1309 ( 
.A(n_988),
.Y(n_1309)
);

INVx1_ASAP7_75t_L g1310 ( 
.A(n_989),
.Y(n_1310)
);

CKINVDCx5p33_ASAP7_75t_R g1311 ( 
.A(n_893),
.Y(n_1311)
);

CKINVDCx16_ASAP7_75t_R g1312 ( 
.A(n_982),
.Y(n_1312)
);

INVx2_ASAP7_75t_L g1313 ( 
.A(n_870),
.Y(n_1313)
);

CKINVDCx5p33_ASAP7_75t_R g1314 ( 
.A(n_897),
.Y(n_1314)
);

INVx1_ASAP7_75t_L g1315 ( 
.A(n_998),
.Y(n_1315)
);

BUFx3_ASAP7_75t_L g1316 ( 
.A(n_982),
.Y(n_1316)
);

CKINVDCx16_ASAP7_75t_R g1317 ( 
.A(n_982),
.Y(n_1317)
);

CKINVDCx5p33_ASAP7_75t_R g1318 ( 
.A(n_898),
.Y(n_1318)
);

INVx2_ASAP7_75t_L g1319 ( 
.A(n_885),
.Y(n_1319)
);

INVx1_ASAP7_75t_L g1320 ( 
.A(n_1009),
.Y(n_1320)
);

INVx1_ASAP7_75t_L g1321 ( 
.A(n_1016),
.Y(n_1321)
);

INVx1_ASAP7_75t_L g1322 ( 
.A(n_1026),
.Y(n_1322)
);

CKINVDCx5p33_ASAP7_75t_R g1323 ( 
.A(n_899),
.Y(n_1323)
);

INVx1_ASAP7_75t_L g1324 ( 
.A(n_1029),
.Y(n_1324)
);

CKINVDCx5p33_ASAP7_75t_R g1325 ( 
.A(n_900),
.Y(n_1325)
);

OR2x2_ASAP7_75t_L g1326 ( 
.A(n_946),
.B(n_4),
.Y(n_1326)
);

INVx1_ASAP7_75t_L g1327 ( 
.A(n_1033),
.Y(n_1327)
);

CKINVDCx5p33_ASAP7_75t_R g1328 ( 
.A(n_901),
.Y(n_1328)
);

CKINVDCx5p33_ASAP7_75t_R g1329 ( 
.A(n_902),
.Y(n_1329)
);

CKINVDCx5p33_ASAP7_75t_R g1330 ( 
.A(n_903),
.Y(n_1330)
);

INVx1_ASAP7_75t_L g1331 ( 
.A(n_885),
.Y(n_1331)
);

CKINVDCx5p33_ASAP7_75t_R g1332 ( 
.A(n_906),
.Y(n_1332)
);

INVx1_ASAP7_75t_L g1333 ( 
.A(n_892),
.Y(n_1333)
);

INVx1_ASAP7_75t_L g1334 ( 
.A(n_892),
.Y(n_1334)
);

CKINVDCx16_ASAP7_75t_R g1335 ( 
.A(n_1001),
.Y(n_1335)
);

CKINVDCx16_ASAP7_75t_R g1336 ( 
.A(n_1013),
.Y(n_1336)
);

INVx1_ASAP7_75t_L g1337 ( 
.A(n_938),
.Y(n_1337)
);

NOR2xp67_ASAP7_75t_L g1338 ( 
.A(n_933),
.B(n_2),
.Y(n_1338)
);

INVx1_ASAP7_75t_L g1339 ( 
.A(n_938),
.Y(n_1339)
);

INVx2_ASAP7_75t_L g1340 ( 
.A(n_971),
.Y(n_1340)
);

INVx1_ASAP7_75t_L g1341 ( 
.A(n_971),
.Y(n_1341)
);

INVx1_ASAP7_75t_L g1342 ( 
.A(n_977),
.Y(n_1342)
);

INVx1_ASAP7_75t_L g1343 ( 
.A(n_977),
.Y(n_1343)
);

CKINVDCx5p33_ASAP7_75t_R g1344 ( 
.A(n_909),
.Y(n_1344)
);

INVx1_ASAP7_75t_L g1345 ( 
.A(n_990),
.Y(n_1345)
);

INVx1_ASAP7_75t_L g1346 ( 
.A(n_990),
.Y(n_1346)
);

CKINVDCx16_ASAP7_75t_R g1347 ( 
.A(n_1017),
.Y(n_1347)
);

INVx1_ASAP7_75t_L g1348 ( 
.A(n_992),
.Y(n_1348)
);

INVx1_ASAP7_75t_L g1349 ( 
.A(n_942),
.Y(n_1349)
);

BUFx6f_ASAP7_75t_L g1350 ( 
.A(n_942),
.Y(n_1350)
);

INVx1_ASAP7_75t_L g1351 ( 
.A(n_910),
.Y(n_1351)
);

CKINVDCx5p33_ASAP7_75t_R g1352 ( 
.A(n_916),
.Y(n_1352)
);

CKINVDCx5p33_ASAP7_75t_R g1353 ( 
.A(n_917),
.Y(n_1353)
);

INVx2_ASAP7_75t_L g1354 ( 
.A(n_922),
.Y(n_1354)
);

CKINVDCx20_ASAP7_75t_R g1355 ( 
.A(n_1020),
.Y(n_1355)
);

INVx1_ASAP7_75t_L g1356 ( 
.A(n_923),
.Y(n_1356)
);

CKINVDCx5p33_ASAP7_75t_R g1357 ( 
.A(n_925),
.Y(n_1357)
);

INVx1_ASAP7_75t_L g1358 ( 
.A(n_929),
.Y(n_1358)
);

INVxp67_ASAP7_75t_L g1359 ( 
.A(n_743),
.Y(n_1359)
);

INVx1_ASAP7_75t_L g1360 ( 
.A(n_930),
.Y(n_1360)
);

INVx2_ASAP7_75t_SL g1361 ( 
.A(n_748),
.Y(n_1361)
);

BUFx6f_ASAP7_75t_L g1362 ( 
.A(n_931),
.Y(n_1362)
);

INVxp67_ASAP7_75t_L g1363 ( 
.A(n_748),
.Y(n_1363)
);

INVx1_ASAP7_75t_L g1364 ( 
.A(n_932),
.Y(n_1364)
);

CKINVDCx5p33_ASAP7_75t_R g1365 ( 
.A(n_935),
.Y(n_1365)
);

INVx1_ASAP7_75t_L g1366 ( 
.A(n_936),
.Y(n_1366)
);

INVx1_ASAP7_75t_L g1367 ( 
.A(n_941),
.Y(n_1367)
);

CKINVDCx20_ASAP7_75t_R g1368 ( 
.A(n_767),
.Y(n_1368)
);

CKINVDCx20_ASAP7_75t_R g1369 ( 
.A(n_767),
.Y(n_1369)
);

BUFx6f_ASAP7_75t_L g1370 ( 
.A(n_943),
.Y(n_1370)
);

INVx1_ASAP7_75t_L g1371 ( 
.A(n_947),
.Y(n_1371)
);

INVx1_ASAP7_75t_L g1372 ( 
.A(n_948),
.Y(n_1372)
);

INVx1_ASAP7_75t_SL g1373 ( 
.A(n_981),
.Y(n_1373)
);

CKINVDCx5p33_ASAP7_75t_R g1374 ( 
.A(n_949),
.Y(n_1374)
);

CKINVDCx20_ASAP7_75t_R g1375 ( 
.A(n_981),
.Y(n_1375)
);

INVx1_ASAP7_75t_L g1376 ( 
.A(n_950),
.Y(n_1376)
);

INVx1_ASAP7_75t_L g1377 ( 
.A(n_951),
.Y(n_1377)
);

CKINVDCx5p33_ASAP7_75t_R g1378 ( 
.A(n_952),
.Y(n_1378)
);

INVx1_ASAP7_75t_L g1379 ( 
.A(n_953),
.Y(n_1379)
);

CKINVDCx20_ASAP7_75t_R g1380 ( 
.A(n_993),
.Y(n_1380)
);

INVx1_ASAP7_75t_L g1381 ( 
.A(n_956),
.Y(n_1381)
);

CKINVDCx5p33_ASAP7_75t_R g1382 ( 
.A(n_957),
.Y(n_1382)
);

INVx1_ASAP7_75t_L g1383 ( 
.A(n_958),
.Y(n_1383)
);

CKINVDCx5p33_ASAP7_75t_R g1384 ( 
.A(n_960),
.Y(n_1384)
);

INVx1_ASAP7_75t_L g1385 ( 
.A(n_962),
.Y(n_1385)
);

CKINVDCx5p33_ASAP7_75t_R g1386 ( 
.A(n_963),
.Y(n_1386)
);

CKINVDCx5p33_ASAP7_75t_R g1387 ( 
.A(n_973),
.Y(n_1387)
);

CKINVDCx16_ASAP7_75t_R g1388 ( 
.A(n_808),
.Y(n_1388)
);

INVx1_ASAP7_75t_L g1389 ( 
.A(n_1034),
.Y(n_1389)
);

HB1xp67_ASAP7_75t_L g1390 ( 
.A(n_993),
.Y(n_1390)
);

INVx1_ASAP7_75t_L g1391 ( 
.A(n_699),
.Y(n_1391)
);

INVx1_ASAP7_75t_SL g1392 ( 
.A(n_821),
.Y(n_1392)
);

INVx1_ASAP7_75t_L g1393 ( 
.A(n_1032),
.Y(n_1393)
);

INVx1_ASAP7_75t_L g1394 ( 
.A(n_1032),
.Y(n_1394)
);

INVx1_ASAP7_75t_L g1395 ( 
.A(n_699),
.Y(n_1395)
);

INVx1_ASAP7_75t_L g1396 ( 
.A(n_1031),
.Y(n_1396)
);

INVx1_ASAP7_75t_L g1397 ( 
.A(n_1031),
.Y(n_1397)
);

BUFx6f_ASAP7_75t_L g1398 ( 
.A(n_700),
.Y(n_1398)
);

INVx1_ASAP7_75t_L g1399 ( 
.A(n_1163),
.Y(n_1399)
);

INVx1_ASAP7_75t_L g1400 ( 
.A(n_1174),
.Y(n_1400)
);

INVx1_ASAP7_75t_SL g1401 ( 
.A(n_1072),
.Y(n_1401)
);

INVx2_ASAP7_75t_L g1402 ( 
.A(n_1131),
.Y(n_1402)
);

INVx1_ASAP7_75t_L g1403 ( 
.A(n_1179),
.Y(n_1403)
);

INVx1_ASAP7_75t_L g1404 ( 
.A(n_1180),
.Y(n_1404)
);

CKINVDCx5p33_ASAP7_75t_R g1405 ( 
.A(n_1040),
.Y(n_1405)
);

CKINVDCx20_ASAP7_75t_R g1406 ( 
.A(n_1069),
.Y(n_1406)
);

CKINVDCx5p33_ASAP7_75t_R g1407 ( 
.A(n_1036),
.Y(n_1407)
);

CKINVDCx5p33_ASAP7_75t_R g1408 ( 
.A(n_1036),
.Y(n_1408)
);

CKINVDCx20_ASAP7_75t_R g1409 ( 
.A(n_1069),
.Y(n_1409)
);

NOR2xp67_ASAP7_75t_L g1410 ( 
.A(n_1241),
.B(n_1251),
.Y(n_1410)
);

CKINVDCx5p33_ASAP7_75t_R g1411 ( 
.A(n_1299),
.Y(n_1411)
);

CKINVDCx5p33_ASAP7_75t_R g1412 ( 
.A(n_1299),
.Y(n_1412)
);

INVx1_ASAP7_75t_L g1413 ( 
.A(n_1184),
.Y(n_1413)
);

CKINVDCx5p33_ASAP7_75t_R g1414 ( 
.A(n_1253),
.Y(n_1414)
);

BUFx2_ASAP7_75t_L g1415 ( 
.A(n_1041),
.Y(n_1415)
);

INVx1_ASAP7_75t_L g1416 ( 
.A(n_1185),
.Y(n_1416)
);

NOR2xp67_ASAP7_75t_L g1417 ( 
.A(n_1256),
.B(n_2),
.Y(n_1417)
);

CKINVDCx5p33_ASAP7_75t_R g1418 ( 
.A(n_1259),
.Y(n_1418)
);

INVxp67_ASAP7_75t_SL g1419 ( 
.A(n_1362),
.Y(n_1419)
);

NOR2xp33_ASAP7_75t_L g1420 ( 
.A(n_1386),
.B(n_700),
.Y(n_1420)
);

CKINVDCx20_ASAP7_75t_R g1421 ( 
.A(n_1079),
.Y(n_1421)
);

CKINVDCx5p33_ASAP7_75t_R g1422 ( 
.A(n_1387),
.Y(n_1422)
);

INVx1_ASAP7_75t_L g1423 ( 
.A(n_1187),
.Y(n_1423)
);

INVx2_ASAP7_75t_L g1424 ( 
.A(n_1131),
.Y(n_1424)
);

INVx1_ASAP7_75t_L g1425 ( 
.A(n_1191),
.Y(n_1425)
);

HB1xp67_ASAP7_75t_L g1426 ( 
.A(n_1038),
.Y(n_1426)
);

CKINVDCx5p33_ASAP7_75t_R g1427 ( 
.A(n_1130),
.Y(n_1427)
);

CKINVDCx5p33_ASAP7_75t_R g1428 ( 
.A(n_1137),
.Y(n_1428)
);

INVxp67_ASAP7_75t_L g1429 ( 
.A(n_1392),
.Y(n_1429)
);

INVxp67_ASAP7_75t_L g1430 ( 
.A(n_1189),
.Y(n_1430)
);

NOR2xp33_ASAP7_75t_L g1431 ( 
.A(n_1362),
.B(n_701),
.Y(n_1431)
);

CKINVDCx20_ASAP7_75t_R g1432 ( 
.A(n_1079),
.Y(n_1432)
);

CKINVDCx20_ASAP7_75t_R g1433 ( 
.A(n_1083),
.Y(n_1433)
);

INVxp67_ASAP7_75t_L g1434 ( 
.A(n_1307),
.Y(n_1434)
);

CKINVDCx5p33_ASAP7_75t_R g1435 ( 
.A(n_1145),
.Y(n_1435)
);

CKINVDCx5p33_ASAP7_75t_R g1436 ( 
.A(n_1146),
.Y(n_1436)
);

BUFx2_ASAP7_75t_L g1437 ( 
.A(n_1048),
.Y(n_1437)
);

CKINVDCx20_ASAP7_75t_R g1438 ( 
.A(n_1083),
.Y(n_1438)
);

CKINVDCx5p33_ASAP7_75t_R g1439 ( 
.A(n_1149),
.Y(n_1439)
);

INVxp67_ASAP7_75t_L g1440 ( 
.A(n_1390),
.Y(n_1440)
);

INVx1_ASAP7_75t_L g1441 ( 
.A(n_1192),
.Y(n_1441)
);

BUFx3_ASAP7_75t_L g1442 ( 
.A(n_1169),
.Y(n_1442)
);

CKINVDCx20_ASAP7_75t_R g1443 ( 
.A(n_1088),
.Y(n_1443)
);

INVx1_ASAP7_75t_L g1444 ( 
.A(n_1193),
.Y(n_1444)
);

CKINVDCx20_ASAP7_75t_R g1445 ( 
.A(n_1088),
.Y(n_1445)
);

INVx1_ASAP7_75t_L g1446 ( 
.A(n_1177),
.Y(n_1446)
);

INVxp67_ASAP7_75t_SL g1447 ( 
.A(n_1362),
.Y(n_1447)
);

BUFx6f_ASAP7_75t_L g1448 ( 
.A(n_1131),
.Y(n_1448)
);

CKINVDCx5p33_ASAP7_75t_R g1449 ( 
.A(n_1150),
.Y(n_1449)
);

CKINVDCx16_ASAP7_75t_R g1450 ( 
.A(n_1335),
.Y(n_1450)
);

CKINVDCx5p33_ASAP7_75t_R g1451 ( 
.A(n_1154),
.Y(n_1451)
);

CKINVDCx5p33_ASAP7_75t_R g1452 ( 
.A(n_1156),
.Y(n_1452)
);

INVx1_ASAP7_75t_L g1453 ( 
.A(n_1177),
.Y(n_1453)
);

INVx1_ASAP7_75t_L g1454 ( 
.A(n_1084),
.Y(n_1454)
);

CKINVDCx5p33_ASAP7_75t_R g1455 ( 
.A(n_1162),
.Y(n_1455)
);

INVxp33_ASAP7_75t_L g1456 ( 
.A(n_1157),
.Y(n_1456)
);

CKINVDCx16_ASAP7_75t_R g1457 ( 
.A(n_1336),
.Y(n_1457)
);

INVx1_ASAP7_75t_L g1458 ( 
.A(n_1087),
.Y(n_1458)
);

CKINVDCx5p33_ASAP7_75t_R g1459 ( 
.A(n_1200),
.Y(n_1459)
);

NOR2xp33_ASAP7_75t_L g1460 ( 
.A(n_1362),
.B(n_701),
.Y(n_1460)
);

INVx1_ASAP7_75t_L g1461 ( 
.A(n_1092),
.Y(n_1461)
);

NOR2xp33_ASAP7_75t_L g1462 ( 
.A(n_1370),
.B(n_702),
.Y(n_1462)
);

INVxp33_ASAP7_75t_SL g1463 ( 
.A(n_1048),
.Y(n_1463)
);

INVx2_ASAP7_75t_L g1464 ( 
.A(n_1131),
.Y(n_1464)
);

INVx1_ASAP7_75t_L g1465 ( 
.A(n_1129),
.Y(n_1465)
);

CKINVDCx5p33_ASAP7_75t_R g1466 ( 
.A(n_1201),
.Y(n_1466)
);

CKINVDCx5p33_ASAP7_75t_R g1467 ( 
.A(n_1204),
.Y(n_1467)
);

NOR2xp33_ASAP7_75t_L g1468 ( 
.A(n_1370),
.B(n_702),
.Y(n_1468)
);

CKINVDCx16_ASAP7_75t_R g1469 ( 
.A(n_1347),
.Y(n_1469)
);

NOR2xp33_ASAP7_75t_L g1470 ( 
.A(n_1370),
.B(n_704),
.Y(n_1470)
);

INVx1_ASAP7_75t_L g1471 ( 
.A(n_1129),
.Y(n_1471)
);

INVx2_ASAP7_75t_L g1472 ( 
.A(n_1159),
.Y(n_1472)
);

CKINVDCx5p33_ASAP7_75t_R g1473 ( 
.A(n_1211),
.Y(n_1473)
);

CKINVDCx5p33_ASAP7_75t_R g1474 ( 
.A(n_1218),
.Y(n_1474)
);

INVx2_ASAP7_75t_L g1475 ( 
.A(n_1159),
.Y(n_1475)
);

CKINVDCx20_ASAP7_75t_R g1476 ( 
.A(n_1102),
.Y(n_1476)
);

NOR2xp33_ASAP7_75t_L g1477 ( 
.A(n_1370),
.B(n_704),
.Y(n_1477)
);

INVxp67_ASAP7_75t_SL g1478 ( 
.A(n_1398),
.Y(n_1478)
);

BUFx3_ASAP7_75t_L g1479 ( 
.A(n_1169),
.Y(n_1479)
);

INVx1_ASAP7_75t_L g1480 ( 
.A(n_1165),
.Y(n_1480)
);

CKINVDCx5p33_ASAP7_75t_R g1481 ( 
.A(n_1221),
.Y(n_1481)
);

CKINVDCx20_ASAP7_75t_R g1482 ( 
.A(n_1102),
.Y(n_1482)
);

INVx1_ASAP7_75t_L g1483 ( 
.A(n_1165),
.Y(n_1483)
);

INVxp33_ASAP7_75t_L g1484 ( 
.A(n_1182),
.Y(n_1484)
);

INVx1_ASAP7_75t_L g1485 ( 
.A(n_1166),
.Y(n_1485)
);

CKINVDCx5p33_ASAP7_75t_R g1486 ( 
.A(n_1223),
.Y(n_1486)
);

INVxp67_ASAP7_75t_L g1487 ( 
.A(n_1210),
.Y(n_1487)
);

HB1xp67_ASAP7_75t_L g1488 ( 
.A(n_1049),
.Y(n_1488)
);

NOR2xp33_ASAP7_75t_L g1489 ( 
.A(n_1224),
.B(n_705),
.Y(n_1489)
);

INVx1_ASAP7_75t_L g1490 ( 
.A(n_1166),
.Y(n_1490)
);

INVx1_ASAP7_75t_L g1491 ( 
.A(n_1181),
.Y(n_1491)
);

INVx1_ASAP7_75t_L g1492 ( 
.A(n_1181),
.Y(n_1492)
);

INVxp67_ASAP7_75t_SL g1493 ( 
.A(n_1398),
.Y(n_1493)
);

CKINVDCx5p33_ASAP7_75t_R g1494 ( 
.A(n_1230),
.Y(n_1494)
);

CKINVDCx5p33_ASAP7_75t_R g1495 ( 
.A(n_1234),
.Y(n_1495)
);

HB1xp67_ASAP7_75t_L g1496 ( 
.A(n_1049),
.Y(n_1496)
);

OR2x2_ASAP7_75t_L g1497 ( 
.A(n_1388),
.B(n_1373),
.Y(n_1497)
);

INVxp67_ASAP7_75t_SL g1498 ( 
.A(n_1398),
.Y(n_1498)
);

INVx1_ASAP7_75t_L g1499 ( 
.A(n_1183),
.Y(n_1499)
);

CKINVDCx20_ASAP7_75t_R g1500 ( 
.A(n_1104),
.Y(n_1500)
);

CKINVDCx20_ASAP7_75t_R g1501 ( 
.A(n_1104),
.Y(n_1501)
);

CKINVDCx5p33_ASAP7_75t_R g1502 ( 
.A(n_1236),
.Y(n_1502)
);

INVx1_ASAP7_75t_L g1503 ( 
.A(n_1183),
.Y(n_1503)
);

CKINVDCx5p33_ASAP7_75t_R g1504 ( 
.A(n_1052),
.Y(n_1504)
);

CKINVDCx5p33_ASAP7_75t_R g1505 ( 
.A(n_1052),
.Y(n_1505)
);

INVx1_ASAP7_75t_L g1506 ( 
.A(n_1169),
.Y(n_1506)
);

CKINVDCx20_ASAP7_75t_R g1507 ( 
.A(n_1118),
.Y(n_1507)
);

INVxp67_ASAP7_75t_SL g1508 ( 
.A(n_1398),
.Y(n_1508)
);

CKINVDCx5p33_ASAP7_75t_R g1509 ( 
.A(n_1056),
.Y(n_1509)
);

CKINVDCx5p33_ASAP7_75t_R g1510 ( 
.A(n_1056),
.Y(n_1510)
);

BUFx3_ASAP7_75t_L g1511 ( 
.A(n_1093),
.Y(n_1511)
);

INVx1_ASAP7_75t_L g1512 ( 
.A(n_1205),
.Y(n_1512)
);

INVx1_ASAP7_75t_L g1513 ( 
.A(n_1209),
.Y(n_1513)
);

INVx1_ASAP7_75t_L g1514 ( 
.A(n_1212),
.Y(n_1514)
);

CKINVDCx5p33_ASAP7_75t_R g1515 ( 
.A(n_1057),
.Y(n_1515)
);

INVxp67_ASAP7_75t_SL g1516 ( 
.A(n_1354),
.Y(n_1516)
);

CKINVDCx5p33_ASAP7_75t_R g1517 ( 
.A(n_1057),
.Y(n_1517)
);

INVx1_ASAP7_75t_L g1518 ( 
.A(n_1213),
.Y(n_1518)
);

CKINVDCx5p33_ASAP7_75t_R g1519 ( 
.A(n_1060),
.Y(n_1519)
);

NAND2xp33_ASAP7_75t_R g1520 ( 
.A(n_1060),
.B(n_705),
.Y(n_1520)
);

CKINVDCx5p33_ASAP7_75t_R g1521 ( 
.A(n_1071),
.Y(n_1521)
);

INVx2_ASAP7_75t_L g1522 ( 
.A(n_1159),
.Y(n_1522)
);

CKINVDCx16_ASAP7_75t_R g1523 ( 
.A(n_1128),
.Y(n_1523)
);

CKINVDCx5p33_ASAP7_75t_R g1524 ( 
.A(n_1071),
.Y(n_1524)
);

CKINVDCx5p33_ASAP7_75t_R g1525 ( 
.A(n_1074),
.Y(n_1525)
);

CKINVDCx5p33_ASAP7_75t_R g1526 ( 
.A(n_1074),
.Y(n_1526)
);

BUFx2_ASAP7_75t_L g1527 ( 
.A(n_1078),
.Y(n_1527)
);

INVx1_ASAP7_75t_L g1528 ( 
.A(n_1214),
.Y(n_1528)
);

CKINVDCx20_ASAP7_75t_R g1529 ( 
.A(n_1118),
.Y(n_1529)
);

CKINVDCx5p33_ASAP7_75t_R g1530 ( 
.A(n_1078),
.Y(n_1530)
);

CKINVDCx5p33_ASAP7_75t_R g1531 ( 
.A(n_1080),
.Y(n_1531)
);

CKINVDCx5p33_ASAP7_75t_R g1532 ( 
.A(n_1080),
.Y(n_1532)
);

CKINVDCx5p33_ASAP7_75t_R g1533 ( 
.A(n_1086),
.Y(n_1533)
);

CKINVDCx20_ASAP7_75t_R g1534 ( 
.A(n_1126),
.Y(n_1534)
);

CKINVDCx20_ASAP7_75t_R g1535 ( 
.A(n_1126),
.Y(n_1535)
);

INVxp33_ASAP7_75t_SL g1536 ( 
.A(n_1086),
.Y(n_1536)
);

NOR2xp67_ASAP7_75t_L g1537 ( 
.A(n_1359),
.B(n_4),
.Y(n_1537)
);

CKINVDCx20_ASAP7_75t_R g1538 ( 
.A(n_1134),
.Y(n_1538)
);

CKINVDCx5p33_ASAP7_75t_R g1539 ( 
.A(n_1090),
.Y(n_1539)
);

CKINVDCx20_ASAP7_75t_R g1540 ( 
.A(n_1134),
.Y(n_1540)
);

INVx1_ASAP7_75t_SL g1541 ( 
.A(n_1085),
.Y(n_1541)
);

CKINVDCx20_ASAP7_75t_R g1542 ( 
.A(n_1138),
.Y(n_1542)
);

INVx2_ASAP7_75t_L g1543 ( 
.A(n_1159),
.Y(n_1543)
);

INVx1_ASAP7_75t_L g1544 ( 
.A(n_1215),
.Y(n_1544)
);

BUFx2_ASAP7_75t_L g1545 ( 
.A(n_1090),
.Y(n_1545)
);

CKINVDCx5p33_ASAP7_75t_R g1546 ( 
.A(n_1095),
.Y(n_1546)
);

NAND2xp5_ASAP7_75t_L g1547 ( 
.A(n_1351),
.B(n_706),
.Y(n_1547)
);

CKINVDCx5p33_ASAP7_75t_R g1548 ( 
.A(n_1095),
.Y(n_1548)
);

INVxp67_ASAP7_75t_L g1549 ( 
.A(n_1227),
.Y(n_1549)
);

CKINVDCx5p33_ASAP7_75t_R g1550 ( 
.A(n_1096),
.Y(n_1550)
);

INVx1_ASAP7_75t_L g1551 ( 
.A(n_1216),
.Y(n_1551)
);

HB1xp67_ASAP7_75t_L g1552 ( 
.A(n_1096),
.Y(n_1552)
);

CKINVDCx20_ASAP7_75t_R g1553 ( 
.A(n_1138),
.Y(n_1553)
);

INVxp67_ASAP7_75t_SL g1554 ( 
.A(n_1354),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_1220),
.Y(n_1555)
);

CKINVDCx5p33_ASAP7_75t_R g1556 ( 
.A(n_1097),
.Y(n_1556)
);

CKINVDCx5p33_ASAP7_75t_R g1557 ( 
.A(n_1097),
.Y(n_1557)
);

NOR2xp33_ASAP7_75t_L g1558 ( 
.A(n_1098),
.B(n_706),
.Y(n_1558)
);

CKINVDCx5p33_ASAP7_75t_R g1559 ( 
.A(n_1098),
.Y(n_1559)
);

CKINVDCx20_ASAP7_75t_R g1560 ( 
.A(n_1140),
.Y(n_1560)
);

CKINVDCx5p33_ASAP7_75t_R g1561 ( 
.A(n_1100),
.Y(n_1561)
);

INVx1_ASAP7_75t_L g1562 ( 
.A(n_1225),
.Y(n_1562)
);

INVxp67_ASAP7_75t_L g1563 ( 
.A(n_1247),
.Y(n_1563)
);

INVx1_ASAP7_75t_L g1564 ( 
.A(n_1228),
.Y(n_1564)
);

HB1xp67_ASAP7_75t_L g1565 ( 
.A(n_1100),
.Y(n_1565)
);

INVx1_ASAP7_75t_L g1566 ( 
.A(n_1229),
.Y(n_1566)
);

INVx1_ASAP7_75t_L g1567 ( 
.A(n_1232),
.Y(n_1567)
);

INVx1_ASAP7_75t_L g1568 ( 
.A(n_1233),
.Y(n_1568)
);

INVx1_ASAP7_75t_L g1569 ( 
.A(n_1239),
.Y(n_1569)
);

CKINVDCx20_ASAP7_75t_R g1570 ( 
.A(n_1140),
.Y(n_1570)
);

NOR2xp33_ASAP7_75t_L g1571 ( 
.A(n_1103),
.B(n_707),
.Y(n_1571)
);

INVx1_ASAP7_75t_L g1572 ( 
.A(n_1243),
.Y(n_1572)
);

INVx1_ASAP7_75t_L g1573 ( 
.A(n_1244),
.Y(n_1573)
);

INVx1_ASAP7_75t_L g1574 ( 
.A(n_1245),
.Y(n_1574)
);

INVx1_ASAP7_75t_L g1575 ( 
.A(n_1246),
.Y(n_1575)
);

HB1xp67_ASAP7_75t_L g1576 ( 
.A(n_1103),
.Y(n_1576)
);

INVx1_ASAP7_75t_L g1577 ( 
.A(n_1248),
.Y(n_1577)
);

INVx1_ASAP7_75t_L g1578 ( 
.A(n_1249),
.Y(n_1578)
);

CKINVDCx20_ASAP7_75t_R g1579 ( 
.A(n_1272),
.Y(n_1579)
);

HB1xp67_ASAP7_75t_L g1580 ( 
.A(n_1109),
.Y(n_1580)
);

INVx1_ASAP7_75t_L g1581 ( 
.A(n_1250),
.Y(n_1581)
);

CKINVDCx5p33_ASAP7_75t_R g1582 ( 
.A(n_1109),
.Y(n_1582)
);

BUFx3_ASAP7_75t_L g1583 ( 
.A(n_1093),
.Y(n_1583)
);

CKINVDCx20_ASAP7_75t_R g1584 ( 
.A(n_1272),
.Y(n_1584)
);

CKINVDCx20_ASAP7_75t_R g1585 ( 
.A(n_1274),
.Y(n_1585)
);

CKINVDCx20_ASAP7_75t_R g1586 ( 
.A(n_1274),
.Y(n_1586)
);

INVx1_ASAP7_75t_L g1587 ( 
.A(n_1252),
.Y(n_1587)
);

CKINVDCx5p33_ASAP7_75t_R g1588 ( 
.A(n_1110),
.Y(n_1588)
);

NOR2xp67_ASAP7_75t_L g1589 ( 
.A(n_1363),
.B(n_1110),
.Y(n_1589)
);

CKINVDCx5p33_ASAP7_75t_R g1590 ( 
.A(n_1112),
.Y(n_1590)
);

CKINVDCx5p33_ASAP7_75t_R g1591 ( 
.A(n_1112),
.Y(n_1591)
);

BUFx2_ASAP7_75t_L g1592 ( 
.A(n_1114),
.Y(n_1592)
);

CKINVDCx5p33_ASAP7_75t_R g1593 ( 
.A(n_1114),
.Y(n_1593)
);

INVx1_ASAP7_75t_L g1594 ( 
.A(n_1254),
.Y(n_1594)
);

INVx1_ASAP7_75t_L g1595 ( 
.A(n_1255),
.Y(n_1595)
);

CKINVDCx5p33_ASAP7_75t_R g1596 ( 
.A(n_1116),
.Y(n_1596)
);

CKINVDCx5p33_ASAP7_75t_R g1597 ( 
.A(n_1116),
.Y(n_1597)
);

INVx1_ASAP7_75t_L g1598 ( 
.A(n_1261),
.Y(n_1598)
);

NOR2xp33_ASAP7_75t_L g1599 ( 
.A(n_1117),
.B(n_707),
.Y(n_1599)
);

INVxp67_ASAP7_75t_SL g1600 ( 
.A(n_1356),
.Y(n_1600)
);

CKINVDCx20_ASAP7_75t_R g1601 ( 
.A(n_1296),
.Y(n_1601)
);

INVx1_ASAP7_75t_L g1602 ( 
.A(n_1262),
.Y(n_1602)
);

INVx1_ASAP7_75t_L g1603 ( 
.A(n_1264),
.Y(n_1603)
);

CKINVDCx5p33_ASAP7_75t_R g1604 ( 
.A(n_1117),
.Y(n_1604)
);

NOR2xp33_ASAP7_75t_L g1605 ( 
.A(n_1119),
.B(n_709),
.Y(n_1605)
);

CKINVDCx5p33_ASAP7_75t_R g1606 ( 
.A(n_1119),
.Y(n_1606)
);

INVx2_ASAP7_75t_L g1607 ( 
.A(n_1186),
.Y(n_1607)
);

CKINVDCx5p33_ASAP7_75t_R g1608 ( 
.A(n_1121),
.Y(n_1608)
);

CKINVDCx5p33_ASAP7_75t_R g1609 ( 
.A(n_1121),
.Y(n_1609)
);

INVx1_ASAP7_75t_L g1610 ( 
.A(n_1267),
.Y(n_1610)
);

INVx1_ASAP7_75t_L g1611 ( 
.A(n_1268),
.Y(n_1611)
);

INVx2_ASAP7_75t_L g1612 ( 
.A(n_1186),
.Y(n_1612)
);

NOR2xp67_ASAP7_75t_L g1613 ( 
.A(n_1122),
.B(n_4),
.Y(n_1613)
);

INVx1_ASAP7_75t_L g1614 ( 
.A(n_1269),
.Y(n_1614)
);

CKINVDCx20_ASAP7_75t_R g1615 ( 
.A(n_1296),
.Y(n_1615)
);

CKINVDCx20_ASAP7_75t_R g1616 ( 
.A(n_1298),
.Y(n_1616)
);

AND2x2_ASAP7_75t_L g1617 ( 
.A(n_1350),
.B(n_1141),
.Y(n_1617)
);

CKINVDCx20_ASAP7_75t_R g1618 ( 
.A(n_1298),
.Y(n_1618)
);

INVx1_ASAP7_75t_L g1619 ( 
.A(n_1271),
.Y(n_1619)
);

CKINVDCx5p33_ASAP7_75t_R g1620 ( 
.A(n_1122),
.Y(n_1620)
);

CKINVDCx5p33_ASAP7_75t_R g1621 ( 
.A(n_1164),
.Y(n_1621)
);

INVx1_ASAP7_75t_L g1622 ( 
.A(n_1277),
.Y(n_1622)
);

CKINVDCx20_ASAP7_75t_R g1623 ( 
.A(n_1355),
.Y(n_1623)
);

INVx1_ASAP7_75t_L g1624 ( 
.A(n_1279),
.Y(n_1624)
);

INVx1_ASAP7_75t_L g1625 ( 
.A(n_1283),
.Y(n_1625)
);

INVx1_ASAP7_75t_L g1626 ( 
.A(n_1284),
.Y(n_1626)
);

INVxp33_ASAP7_75t_SL g1627 ( 
.A(n_1164),
.Y(n_1627)
);

INVx2_ASAP7_75t_L g1628 ( 
.A(n_1186),
.Y(n_1628)
);

INVx1_ASAP7_75t_L g1629 ( 
.A(n_1285),
.Y(n_1629)
);

CKINVDCx16_ASAP7_75t_R g1630 ( 
.A(n_1073),
.Y(n_1630)
);

INVx1_ASAP7_75t_L g1631 ( 
.A(n_1287),
.Y(n_1631)
);

INVx2_ASAP7_75t_L g1632 ( 
.A(n_1186),
.Y(n_1632)
);

BUFx3_ASAP7_75t_L g1633 ( 
.A(n_1123),
.Y(n_1633)
);

BUFx3_ASAP7_75t_L g1634 ( 
.A(n_1123),
.Y(n_1634)
);

CKINVDCx20_ASAP7_75t_R g1635 ( 
.A(n_1355),
.Y(n_1635)
);

INVx1_ASAP7_75t_L g1636 ( 
.A(n_1291),
.Y(n_1636)
);

CKINVDCx5p33_ASAP7_75t_R g1637 ( 
.A(n_1168),
.Y(n_1637)
);

NOR2xp67_ASAP7_75t_L g1638 ( 
.A(n_1168),
.B(n_5),
.Y(n_1638)
);

INVx1_ASAP7_75t_L g1639 ( 
.A(n_1294),
.Y(n_1639)
);

INVx1_ASAP7_75t_L g1640 ( 
.A(n_1295),
.Y(n_1640)
);

HB1xp67_ASAP7_75t_L g1641 ( 
.A(n_1175),
.Y(n_1641)
);

INVx2_ASAP7_75t_L g1642 ( 
.A(n_1208),
.Y(n_1642)
);

HB1xp67_ASAP7_75t_L g1643 ( 
.A(n_1175),
.Y(n_1643)
);

INVx1_ASAP7_75t_L g1644 ( 
.A(n_1297),
.Y(n_1644)
);

INVx1_ASAP7_75t_L g1645 ( 
.A(n_1300),
.Y(n_1645)
);

CKINVDCx5p33_ASAP7_75t_R g1646 ( 
.A(n_1176),
.Y(n_1646)
);

INVxp33_ASAP7_75t_SL g1647 ( 
.A(n_1176),
.Y(n_1647)
);

CKINVDCx5p33_ASAP7_75t_R g1648 ( 
.A(n_1178),
.Y(n_1648)
);

INVxp67_ASAP7_75t_L g1649 ( 
.A(n_1206),
.Y(n_1649)
);

INVx1_ASAP7_75t_L g1650 ( 
.A(n_1302),
.Y(n_1650)
);

INVx1_ASAP7_75t_L g1651 ( 
.A(n_1303),
.Y(n_1651)
);

INVx1_ASAP7_75t_L g1652 ( 
.A(n_1306),
.Y(n_1652)
);

CKINVDCx20_ASAP7_75t_R g1653 ( 
.A(n_1368),
.Y(n_1653)
);

NOR2xp33_ASAP7_75t_L g1654 ( 
.A(n_1178),
.B(n_709),
.Y(n_1654)
);

INVx1_ASAP7_75t_L g1655 ( 
.A(n_1309),
.Y(n_1655)
);

CKINVDCx5p33_ASAP7_75t_R g1656 ( 
.A(n_1190),
.Y(n_1656)
);

CKINVDCx5p33_ASAP7_75t_R g1657 ( 
.A(n_1190),
.Y(n_1657)
);

CKINVDCx5p33_ASAP7_75t_R g1658 ( 
.A(n_1195),
.Y(n_1658)
);

INVx1_ASAP7_75t_L g1659 ( 
.A(n_1310),
.Y(n_1659)
);

INVxp33_ASAP7_75t_L g1660 ( 
.A(n_1045),
.Y(n_1660)
);

CKINVDCx20_ASAP7_75t_R g1661 ( 
.A(n_1368),
.Y(n_1661)
);

CKINVDCx5p33_ASAP7_75t_R g1662 ( 
.A(n_1195),
.Y(n_1662)
);

INVx1_ASAP7_75t_L g1663 ( 
.A(n_1315),
.Y(n_1663)
);

INVx2_ASAP7_75t_L g1664 ( 
.A(n_1208),
.Y(n_1664)
);

INVxp33_ASAP7_75t_SL g1665 ( 
.A(n_1260),
.Y(n_1665)
);

CKINVDCx16_ASAP7_75t_R g1666 ( 
.A(n_1081),
.Y(n_1666)
);

BUFx2_ASAP7_75t_SL g1667 ( 
.A(n_1369),
.Y(n_1667)
);

INVx1_ASAP7_75t_L g1668 ( 
.A(n_1320),
.Y(n_1668)
);

INVx1_ASAP7_75t_L g1669 ( 
.A(n_1321),
.Y(n_1669)
);

INVx1_ASAP7_75t_L g1670 ( 
.A(n_1322),
.Y(n_1670)
);

CKINVDCx20_ASAP7_75t_R g1671 ( 
.A(n_1369),
.Y(n_1671)
);

INVx1_ASAP7_75t_L g1672 ( 
.A(n_1324),
.Y(n_1672)
);

INVx1_ASAP7_75t_L g1673 ( 
.A(n_1327),
.Y(n_1673)
);

INVx1_ASAP7_75t_L g1674 ( 
.A(n_1144),
.Y(n_1674)
);

CKINVDCx5p33_ASAP7_75t_R g1675 ( 
.A(n_1260),
.Y(n_1675)
);

NAND2xp5_ASAP7_75t_L g1676 ( 
.A(n_1358),
.B(n_712),
.Y(n_1676)
);

CKINVDCx5p33_ASAP7_75t_R g1677 ( 
.A(n_1270),
.Y(n_1677)
);

CKINVDCx5p33_ASAP7_75t_R g1678 ( 
.A(n_1270),
.Y(n_1678)
);

CKINVDCx5p33_ASAP7_75t_R g1679 ( 
.A(n_1273),
.Y(n_1679)
);

INVx1_ASAP7_75t_L g1680 ( 
.A(n_1147),
.Y(n_1680)
);

CKINVDCx5p33_ASAP7_75t_R g1681 ( 
.A(n_1273),
.Y(n_1681)
);

INVx1_ASAP7_75t_L g1682 ( 
.A(n_1148),
.Y(n_1682)
);

INVx1_ASAP7_75t_L g1683 ( 
.A(n_1151),
.Y(n_1683)
);

INVxp67_ASAP7_75t_SL g1684 ( 
.A(n_1360),
.Y(n_1684)
);

CKINVDCx20_ASAP7_75t_R g1685 ( 
.A(n_1375),
.Y(n_1685)
);

CKINVDCx5p33_ASAP7_75t_R g1686 ( 
.A(n_1276),
.Y(n_1686)
);

BUFx2_ASAP7_75t_SL g1687 ( 
.A(n_1375),
.Y(n_1687)
);

INVx1_ASAP7_75t_L g1688 ( 
.A(n_1152),
.Y(n_1688)
);

CKINVDCx20_ASAP7_75t_R g1689 ( 
.A(n_1380),
.Y(n_1689)
);

BUFx3_ASAP7_75t_L g1690 ( 
.A(n_1124),
.Y(n_1690)
);

INVx1_ASAP7_75t_L g1691 ( 
.A(n_1153),
.Y(n_1691)
);

INVxp67_ASAP7_75t_SL g1692 ( 
.A(n_1364),
.Y(n_1692)
);

CKINVDCx5p33_ASAP7_75t_R g1693 ( 
.A(n_1276),
.Y(n_1693)
);

CKINVDCx16_ASAP7_75t_R g1694 ( 
.A(n_1089),
.Y(n_1694)
);

CKINVDCx20_ASAP7_75t_R g1695 ( 
.A(n_1380),
.Y(n_1695)
);

INVx1_ASAP7_75t_L g1696 ( 
.A(n_1155),
.Y(n_1696)
);

CKINVDCx16_ASAP7_75t_R g1697 ( 
.A(n_1293),
.Y(n_1697)
);

CKINVDCx5p33_ASAP7_75t_R g1698 ( 
.A(n_1281),
.Y(n_1698)
);

CKINVDCx5p33_ASAP7_75t_R g1699 ( 
.A(n_1281),
.Y(n_1699)
);

CKINVDCx16_ASAP7_75t_R g1700 ( 
.A(n_1312),
.Y(n_1700)
);

CKINVDCx20_ASAP7_75t_R g1701 ( 
.A(n_1171),
.Y(n_1701)
);

INVx1_ASAP7_75t_L g1702 ( 
.A(n_1158),
.Y(n_1702)
);

INVx1_ASAP7_75t_L g1703 ( 
.A(n_1160),
.Y(n_1703)
);

INVxp67_ASAP7_75t_SL g1704 ( 
.A(n_1366),
.Y(n_1704)
);

INVx1_ASAP7_75t_L g1705 ( 
.A(n_1617),
.Y(n_1705)
);

OA21x2_ASAP7_75t_L g1706 ( 
.A1(n_1400),
.A2(n_1037),
.B(n_1035),
.Y(n_1706)
);

INVx2_ASAP7_75t_L g1707 ( 
.A(n_1465),
.Y(n_1707)
);

INVx2_ASAP7_75t_L g1708 ( 
.A(n_1471),
.Y(n_1708)
);

NAND2xp5_ASAP7_75t_L g1709 ( 
.A(n_1478),
.B(n_1367),
.Y(n_1709)
);

BUFx6f_ASAP7_75t_L g1710 ( 
.A(n_1448),
.Y(n_1710)
);

INVx2_ASAP7_75t_L g1711 ( 
.A(n_1480),
.Y(n_1711)
);

INVx1_ASAP7_75t_L g1712 ( 
.A(n_1617),
.Y(n_1712)
);

INVx2_ASAP7_75t_L g1713 ( 
.A(n_1483),
.Y(n_1713)
);

BUFx6f_ASAP7_75t_L g1714 ( 
.A(n_1448),
.Y(n_1714)
);

INVx3_ASAP7_75t_L g1715 ( 
.A(n_1448),
.Y(n_1715)
);

NAND2xp5_ASAP7_75t_L g1716 ( 
.A(n_1493),
.B(n_1371),
.Y(n_1716)
);

INVx2_ASAP7_75t_L g1717 ( 
.A(n_1485),
.Y(n_1717)
);

INVx1_ASAP7_75t_L g1718 ( 
.A(n_1674),
.Y(n_1718)
);

BUFx6f_ASAP7_75t_L g1719 ( 
.A(n_1448),
.Y(n_1719)
);

AOI22xp5_ASAP7_75t_L g1720 ( 
.A1(n_1589),
.A2(n_1094),
.B1(n_1288),
.B2(n_1286),
.Y(n_1720)
);

OAI21x1_ASAP7_75t_L g1721 ( 
.A1(n_1547),
.A2(n_1043),
.B(n_1042),
.Y(n_1721)
);

NAND2xp5_ASAP7_75t_L g1722 ( 
.A(n_1498),
.B(n_1508),
.Y(n_1722)
);

INVxp67_ASAP7_75t_L g1723 ( 
.A(n_1429),
.Y(n_1723)
);

INVx2_ASAP7_75t_L g1724 ( 
.A(n_1490),
.Y(n_1724)
);

INVx4_ASAP7_75t_L g1725 ( 
.A(n_1448),
.Y(n_1725)
);

BUFx8_ASAP7_75t_L g1726 ( 
.A(n_1437),
.Y(n_1726)
);

INVx2_ASAP7_75t_L g1727 ( 
.A(n_1491),
.Y(n_1727)
);

INVx3_ASAP7_75t_L g1728 ( 
.A(n_1402),
.Y(n_1728)
);

AND2x2_ASAP7_75t_L g1729 ( 
.A(n_1660),
.B(n_1198),
.Y(n_1729)
);

NAND2xp5_ASAP7_75t_L g1730 ( 
.A(n_1516),
.B(n_1372),
.Y(n_1730)
);

HB1xp67_ASAP7_75t_L g1731 ( 
.A(n_1401),
.Y(n_1731)
);

INVx1_ASAP7_75t_L g1732 ( 
.A(n_1680),
.Y(n_1732)
);

OAI22xp5_ASAP7_75t_L g1733 ( 
.A1(n_1600),
.A2(n_1094),
.B1(n_1188),
.B2(n_1050),
.Y(n_1733)
);

INVx2_ASAP7_75t_L g1734 ( 
.A(n_1492),
.Y(n_1734)
);

NAND2xp5_ASAP7_75t_L g1735 ( 
.A(n_1554),
.B(n_1376),
.Y(n_1735)
);

NAND2xp33_ASAP7_75t_L g1736 ( 
.A(n_1676),
.B(n_1226),
.Y(n_1736)
);

INVx3_ASAP7_75t_L g1737 ( 
.A(n_1402),
.Y(n_1737)
);

BUFx3_ASAP7_75t_L g1738 ( 
.A(n_1511),
.Y(n_1738)
);

OAI22xp5_ASAP7_75t_L g1739 ( 
.A1(n_1684),
.A2(n_1188),
.B1(n_1288),
.B2(n_1286),
.Y(n_1739)
);

BUFx6f_ASAP7_75t_L g1740 ( 
.A(n_1424),
.Y(n_1740)
);

OAI22xp5_ASAP7_75t_L g1741 ( 
.A1(n_1692),
.A2(n_1290),
.B1(n_1292),
.B2(n_1289),
.Y(n_1741)
);

OA21x2_ASAP7_75t_L g1742 ( 
.A1(n_1403),
.A2(n_1044),
.B(n_1039),
.Y(n_1742)
);

INVx1_ASAP7_75t_L g1743 ( 
.A(n_1682),
.Y(n_1743)
);

BUFx6f_ASAP7_75t_L g1744 ( 
.A(n_1424),
.Y(n_1744)
);

BUFx2_ASAP7_75t_L g1745 ( 
.A(n_1701),
.Y(n_1745)
);

INVx1_ASAP7_75t_L g1746 ( 
.A(n_1683),
.Y(n_1746)
);

AND2x4_ASAP7_75t_L g1747 ( 
.A(n_1446),
.B(n_1217),
.Y(n_1747)
);

AND2x2_ASAP7_75t_L g1748 ( 
.A(n_1541),
.B(n_1198),
.Y(n_1748)
);

INVx2_ASAP7_75t_SL g1749 ( 
.A(n_1497),
.Y(n_1749)
);

AOI22xp5_ASAP7_75t_L g1750 ( 
.A1(n_1520),
.A2(n_1289),
.B1(n_1292),
.B2(n_1290),
.Y(n_1750)
);

AND2x4_ASAP7_75t_L g1751 ( 
.A(n_1453),
.B(n_1217),
.Y(n_1751)
);

INVx1_ASAP7_75t_L g1752 ( 
.A(n_1688),
.Y(n_1752)
);

AND2x4_ASAP7_75t_L g1753 ( 
.A(n_1419),
.B(n_1235),
.Y(n_1753)
);

OA21x2_ASAP7_75t_L g1754 ( 
.A1(n_1404),
.A2(n_1054),
.B(n_1047),
.Y(n_1754)
);

AND2x4_ASAP7_75t_L g1755 ( 
.A(n_1447),
.B(n_1235),
.Y(n_1755)
);

AND2x4_ASAP7_75t_L g1756 ( 
.A(n_1633),
.B(n_1240),
.Y(n_1756)
);

BUFx6f_ASAP7_75t_L g1757 ( 
.A(n_1464),
.Y(n_1757)
);

AND2x4_ASAP7_75t_L g1758 ( 
.A(n_1633),
.B(n_1240),
.Y(n_1758)
);

INVx1_ASAP7_75t_L g1759 ( 
.A(n_1691),
.Y(n_1759)
);

BUFx8_ASAP7_75t_L g1760 ( 
.A(n_1415),
.Y(n_1760)
);

NAND2xp5_ASAP7_75t_L g1761 ( 
.A(n_1704),
.B(n_1377),
.Y(n_1761)
);

CKINVDCx5p33_ASAP7_75t_R g1762 ( 
.A(n_1523),
.Y(n_1762)
);

INVx1_ASAP7_75t_L g1763 ( 
.A(n_1696),
.Y(n_1763)
);

OAI22xp5_ASAP7_75t_SL g1764 ( 
.A1(n_1653),
.A2(n_1265),
.B1(n_1317),
.B2(n_720),
.Y(n_1764)
);

OA21x2_ASAP7_75t_L g1765 ( 
.A1(n_1413),
.A2(n_1058),
.B(n_1055),
.Y(n_1765)
);

INVx2_ASAP7_75t_L g1766 ( 
.A(n_1499),
.Y(n_1766)
);

BUFx6f_ASAP7_75t_L g1767 ( 
.A(n_1464),
.Y(n_1767)
);

OAI22x1_ASAP7_75t_L g1768 ( 
.A1(n_1430),
.A2(n_1046),
.B1(n_1143),
.B2(n_1142),
.Y(n_1768)
);

INVx2_ASAP7_75t_L g1769 ( 
.A(n_1503),
.Y(n_1769)
);

INVx1_ASAP7_75t_L g1770 ( 
.A(n_1702),
.Y(n_1770)
);

INVx1_ASAP7_75t_L g1771 ( 
.A(n_1703),
.Y(n_1771)
);

INVx1_ASAP7_75t_L g1772 ( 
.A(n_1512),
.Y(n_1772)
);

NOR2xp33_ASAP7_75t_L g1773 ( 
.A(n_1399),
.B(n_1558),
.Y(n_1773)
);

NOR2xp33_ASAP7_75t_L g1774 ( 
.A(n_1571),
.B(n_1599),
.Y(n_1774)
);

NOR2xp33_ASAP7_75t_SL g1775 ( 
.A(n_1414),
.B(n_1418),
.Y(n_1775)
);

BUFx12f_ASAP7_75t_L g1776 ( 
.A(n_1411),
.Y(n_1776)
);

BUFx6f_ASAP7_75t_L g1777 ( 
.A(n_1472),
.Y(n_1777)
);

INVx1_ASAP7_75t_L g1778 ( 
.A(n_1513),
.Y(n_1778)
);

BUFx3_ASAP7_75t_L g1779 ( 
.A(n_1511),
.Y(n_1779)
);

BUFx6f_ASAP7_75t_L g1780 ( 
.A(n_1472),
.Y(n_1780)
);

INVx1_ASAP7_75t_L g1781 ( 
.A(n_1514),
.Y(n_1781)
);

AND2x4_ASAP7_75t_L g1782 ( 
.A(n_1634),
.B(n_1258),
.Y(n_1782)
);

NOR2xp33_ASAP7_75t_L g1783 ( 
.A(n_1605),
.B(n_1301),
.Y(n_1783)
);

INVx2_ASAP7_75t_L g1784 ( 
.A(n_1642),
.Y(n_1784)
);

BUFx2_ASAP7_75t_L g1785 ( 
.A(n_1649),
.Y(n_1785)
);

BUFx6f_ASAP7_75t_L g1786 ( 
.A(n_1475),
.Y(n_1786)
);

AND2x2_ASAP7_75t_L g1787 ( 
.A(n_1489),
.B(n_1301),
.Y(n_1787)
);

INVx1_ASAP7_75t_L g1788 ( 
.A(n_1518),
.Y(n_1788)
);

INVx2_ASAP7_75t_L g1789 ( 
.A(n_1642),
.Y(n_1789)
);

INVx1_ASAP7_75t_L g1790 ( 
.A(n_1528),
.Y(n_1790)
);

BUFx6f_ASAP7_75t_L g1791 ( 
.A(n_1475),
.Y(n_1791)
);

INVx3_ASAP7_75t_L g1792 ( 
.A(n_1522),
.Y(n_1792)
);

AND2x4_ASAP7_75t_L g1793 ( 
.A(n_1634),
.B(n_1258),
.Y(n_1793)
);

INVx1_ASAP7_75t_L g1794 ( 
.A(n_1544),
.Y(n_1794)
);

AND2x6_ASAP7_75t_L g1795 ( 
.A(n_1431),
.B(n_1379),
.Y(n_1795)
);

INVx1_ASAP7_75t_L g1796 ( 
.A(n_1551),
.Y(n_1796)
);

INVx3_ASAP7_75t_L g1797 ( 
.A(n_1522),
.Y(n_1797)
);

OAI21x1_ASAP7_75t_L g1798 ( 
.A1(n_1506),
.A2(n_1043),
.B(n_1059),
.Y(n_1798)
);

HB1xp67_ASAP7_75t_L g1799 ( 
.A(n_1583),
.Y(n_1799)
);

OAI22xp5_ASAP7_75t_L g1800 ( 
.A1(n_1434),
.A2(n_1314),
.B1(n_1318),
.B2(n_1311),
.Y(n_1800)
);

AND2x2_ASAP7_75t_L g1801 ( 
.A(n_1420),
.B(n_1311),
.Y(n_1801)
);

INVx3_ASAP7_75t_L g1802 ( 
.A(n_1543),
.Y(n_1802)
);

AND2x6_ASAP7_75t_L g1803 ( 
.A(n_1460),
.B(n_1383),
.Y(n_1803)
);

HB1xp67_ASAP7_75t_L g1804 ( 
.A(n_1583),
.Y(n_1804)
);

OA21x2_ASAP7_75t_L g1805 ( 
.A1(n_1416),
.A2(n_1062),
.B(n_1061),
.Y(n_1805)
);

BUFx8_ASAP7_75t_L g1806 ( 
.A(n_1527),
.Y(n_1806)
);

OA21x2_ASAP7_75t_L g1807 ( 
.A1(n_1423),
.A2(n_1064),
.B(n_1063),
.Y(n_1807)
);

INVx6_ASAP7_75t_L g1808 ( 
.A(n_1690),
.Y(n_1808)
);

BUFx6f_ASAP7_75t_L g1809 ( 
.A(n_1543),
.Y(n_1809)
);

INVx1_ASAP7_75t_L g1810 ( 
.A(n_1555),
.Y(n_1810)
);

BUFx6f_ASAP7_75t_L g1811 ( 
.A(n_1607),
.Y(n_1811)
);

NOR2xp33_ASAP7_75t_SL g1812 ( 
.A(n_1414),
.B(n_1314),
.Y(n_1812)
);

INVx2_ASAP7_75t_L g1813 ( 
.A(n_1664),
.Y(n_1813)
);

AND2x6_ASAP7_75t_L g1814 ( 
.A(n_1462),
.B(n_1381),
.Y(n_1814)
);

INVx1_ASAP7_75t_L g1815 ( 
.A(n_1562),
.Y(n_1815)
);

NOR2xp33_ASAP7_75t_L g1816 ( 
.A(n_1654),
.B(n_1318),
.Y(n_1816)
);

INVx3_ASAP7_75t_L g1817 ( 
.A(n_1607),
.Y(n_1817)
);

AND2x2_ASAP7_75t_L g1818 ( 
.A(n_1440),
.B(n_1323),
.Y(n_1818)
);

INVx2_ASAP7_75t_L g1819 ( 
.A(n_1664),
.Y(n_1819)
);

INVx3_ASAP7_75t_L g1820 ( 
.A(n_1612),
.Y(n_1820)
);

BUFx6f_ASAP7_75t_L g1821 ( 
.A(n_1612),
.Y(n_1821)
);

HB1xp67_ASAP7_75t_L g1822 ( 
.A(n_1690),
.Y(n_1822)
);

BUFx6f_ASAP7_75t_L g1823 ( 
.A(n_1628),
.Y(n_1823)
);

CKINVDCx5p33_ASAP7_75t_R g1824 ( 
.A(n_1450),
.Y(n_1824)
);

INVx2_ASAP7_75t_L g1825 ( 
.A(n_1628),
.Y(n_1825)
);

INVx1_ASAP7_75t_L g1826 ( 
.A(n_1564),
.Y(n_1826)
);

INVx4_ASAP7_75t_L g1827 ( 
.A(n_1632),
.Y(n_1827)
);

INVx2_ASAP7_75t_L g1828 ( 
.A(n_1632),
.Y(n_1828)
);

INVxp67_ASAP7_75t_L g1829 ( 
.A(n_1468),
.Y(n_1829)
);

INVx1_ASAP7_75t_L g1830 ( 
.A(n_1566),
.Y(n_1830)
);

INVx1_ASAP7_75t_L g1831 ( 
.A(n_1567),
.Y(n_1831)
);

INVx1_ASAP7_75t_L g1832 ( 
.A(n_1568),
.Y(n_1832)
);

INVx1_ASAP7_75t_L g1833 ( 
.A(n_1569),
.Y(n_1833)
);

INVx1_ASAP7_75t_L g1834 ( 
.A(n_1572),
.Y(n_1834)
);

OA21x2_ASAP7_75t_L g1835 ( 
.A1(n_1425),
.A2(n_1066),
.B(n_1065),
.Y(n_1835)
);

AND2x6_ASAP7_75t_L g1836 ( 
.A(n_1470),
.B(n_1385),
.Y(n_1836)
);

BUFx2_ASAP7_75t_L g1837 ( 
.A(n_1661),
.Y(n_1837)
);

BUFx8_ASAP7_75t_SL g1838 ( 
.A(n_1411),
.Y(n_1838)
);

NAND2xp5_ASAP7_75t_L g1839 ( 
.A(n_1477),
.B(n_1389),
.Y(n_1839)
);

INVx1_ASAP7_75t_L g1840 ( 
.A(n_1573),
.Y(n_1840)
);

INVx1_ASAP7_75t_L g1841 ( 
.A(n_1574),
.Y(n_1841)
);

INVx1_ASAP7_75t_L g1842 ( 
.A(n_1575),
.Y(n_1842)
);

HB1xp67_ASAP7_75t_L g1843 ( 
.A(n_1417),
.Y(n_1843)
);

INVx3_ASAP7_75t_L g1844 ( 
.A(n_1441),
.Y(n_1844)
);

INVx1_ASAP7_75t_L g1845 ( 
.A(n_1577),
.Y(n_1845)
);

AND2x2_ASAP7_75t_L g1846 ( 
.A(n_1456),
.B(n_1323),
.Y(n_1846)
);

INVx2_ASAP7_75t_L g1847 ( 
.A(n_1444),
.Y(n_1847)
);

OAI21x1_ASAP7_75t_L g1848 ( 
.A1(n_1454),
.A2(n_1068),
.B(n_1067),
.Y(n_1848)
);

INVx2_ASAP7_75t_L g1849 ( 
.A(n_1458),
.Y(n_1849)
);

HB1xp67_ASAP7_75t_L g1850 ( 
.A(n_1487),
.Y(n_1850)
);

BUFx6f_ASAP7_75t_L g1851 ( 
.A(n_1461),
.Y(n_1851)
);

AND2x4_ASAP7_75t_L g1852 ( 
.A(n_1578),
.B(n_1305),
.Y(n_1852)
);

INVxp67_ASAP7_75t_L g1853 ( 
.A(n_1488),
.Y(n_1853)
);

AND2x4_ASAP7_75t_L g1854 ( 
.A(n_1581),
.B(n_1305),
.Y(n_1854)
);

INVx2_ASAP7_75t_L g1855 ( 
.A(n_1587),
.Y(n_1855)
);

AND2x4_ASAP7_75t_L g1856 ( 
.A(n_1594),
.B(n_1313),
.Y(n_1856)
);

OAI22xp5_ASAP7_75t_L g1857 ( 
.A1(n_1549),
.A2(n_1563),
.B1(n_1410),
.B2(n_1537),
.Y(n_1857)
);

INVx1_ASAP7_75t_L g1858 ( 
.A(n_1595),
.Y(n_1858)
);

BUFx6f_ASAP7_75t_L g1859 ( 
.A(n_1598),
.Y(n_1859)
);

INVx1_ASAP7_75t_L g1860 ( 
.A(n_1602),
.Y(n_1860)
);

NAND2xp5_ASAP7_75t_SL g1861 ( 
.A(n_1613),
.B(n_1325),
.Y(n_1861)
);

BUFx2_ASAP7_75t_L g1862 ( 
.A(n_1671),
.Y(n_1862)
);

NAND2xp5_ASAP7_75t_L g1863 ( 
.A(n_1442),
.B(n_1070),
.Y(n_1863)
);

OA21x2_ASAP7_75t_L g1864 ( 
.A1(n_1603),
.A2(n_1076),
.B(n_1075),
.Y(n_1864)
);

OAI22xp5_ASAP7_75t_L g1865 ( 
.A1(n_1638),
.A2(n_1328),
.B1(n_1329),
.B2(n_1325),
.Y(n_1865)
);

NAND2xp5_ASAP7_75t_L g1866 ( 
.A(n_1442),
.B(n_1077),
.Y(n_1866)
);

INVx1_ASAP7_75t_L g1867 ( 
.A(n_1610),
.Y(n_1867)
);

NAND2xp5_ASAP7_75t_L g1868 ( 
.A(n_1479),
.B(n_1082),
.Y(n_1868)
);

OA21x2_ASAP7_75t_L g1869 ( 
.A1(n_1611),
.A2(n_1319),
.B(n_1313),
.Y(n_1869)
);

INVx1_ASAP7_75t_L g1870 ( 
.A(n_1614),
.Y(n_1870)
);

BUFx6f_ASAP7_75t_L g1871 ( 
.A(n_1619),
.Y(n_1871)
);

AND2x4_ASAP7_75t_L g1872 ( 
.A(n_1622),
.B(n_1319),
.Y(n_1872)
);

INVx2_ASAP7_75t_L g1873 ( 
.A(n_1624),
.Y(n_1873)
);

INVx3_ASAP7_75t_L g1874 ( 
.A(n_1625),
.Y(n_1874)
);

AND2x4_ASAP7_75t_L g1875 ( 
.A(n_1626),
.B(n_1340),
.Y(n_1875)
);

INVx1_ASAP7_75t_L g1876 ( 
.A(n_1629),
.Y(n_1876)
);

INVx2_ASAP7_75t_L g1877 ( 
.A(n_1631),
.Y(n_1877)
);

HB1xp67_ASAP7_75t_L g1878 ( 
.A(n_1496),
.Y(n_1878)
);

OA21x2_ASAP7_75t_L g1879 ( 
.A1(n_1636),
.A2(n_1340),
.B(n_1203),
.Y(n_1879)
);

NAND2xp5_ASAP7_75t_L g1880 ( 
.A(n_1479),
.B(n_1328),
.Y(n_1880)
);

NAND2xp33_ASAP7_75t_L g1881 ( 
.A(n_1639),
.B(n_1329),
.Y(n_1881)
);

BUFx3_ASAP7_75t_L g1882 ( 
.A(n_1640),
.Y(n_1882)
);

HB1xp67_ASAP7_75t_L g1883 ( 
.A(n_1552),
.Y(n_1883)
);

NOR2x1_ASAP7_75t_L g1884 ( 
.A(n_1644),
.B(n_1645),
.Y(n_1884)
);

CKINVDCx5p33_ASAP7_75t_R g1885 ( 
.A(n_1457),
.Y(n_1885)
);

INVx3_ASAP7_75t_L g1886 ( 
.A(n_1650),
.Y(n_1886)
);

INVx3_ASAP7_75t_L g1887 ( 
.A(n_1651),
.Y(n_1887)
);

INVx1_ASAP7_75t_L g1888 ( 
.A(n_1652),
.Y(n_1888)
);

INVx2_ASAP7_75t_L g1889 ( 
.A(n_1655),
.Y(n_1889)
);

INVx2_ASAP7_75t_L g1890 ( 
.A(n_1659),
.Y(n_1890)
);

INVx6_ASAP7_75t_L g1891 ( 
.A(n_1469),
.Y(n_1891)
);

BUFx6f_ASAP7_75t_L g1892 ( 
.A(n_1663),
.Y(n_1892)
);

INVx1_ASAP7_75t_L g1893 ( 
.A(n_1668),
.Y(n_1893)
);

INVx6_ASAP7_75t_L g1894 ( 
.A(n_1697),
.Y(n_1894)
);

OAI21x1_ASAP7_75t_L g1895 ( 
.A1(n_1669),
.A2(n_1203),
.B(n_1194),
.Y(n_1895)
);

BUFx8_ASAP7_75t_L g1896 ( 
.A(n_1545),
.Y(n_1896)
);

NAND2xp5_ASAP7_75t_L g1897 ( 
.A(n_1670),
.B(n_1330),
.Y(n_1897)
);

BUFx2_ASAP7_75t_L g1898 ( 
.A(n_1685),
.Y(n_1898)
);

CKINVDCx20_ASAP7_75t_R g1899 ( 
.A(n_1406),
.Y(n_1899)
);

INVx2_ASAP7_75t_L g1900 ( 
.A(n_1672),
.Y(n_1900)
);

OAI21x1_ASAP7_75t_L g1901 ( 
.A1(n_1673),
.A2(n_1194),
.B(n_1391),
.Y(n_1901)
);

AOI22xp5_ASAP7_75t_L g1902 ( 
.A1(n_1536),
.A2(n_1330),
.B1(n_1344),
.B2(n_1332),
.Y(n_1902)
);

NAND2xp5_ASAP7_75t_L g1903 ( 
.A(n_1473),
.B(n_1332),
.Y(n_1903)
);

INVx2_ASAP7_75t_L g1904 ( 
.A(n_1565),
.Y(n_1904)
);

OAI22xp5_ASAP7_75t_L g1905 ( 
.A1(n_1407),
.A2(n_1352),
.B1(n_1353),
.B2(n_1344),
.Y(n_1905)
);

INVx2_ASAP7_75t_L g1906 ( 
.A(n_1576),
.Y(n_1906)
);

INVx2_ASAP7_75t_L g1907 ( 
.A(n_1580),
.Y(n_1907)
);

AND2x2_ASAP7_75t_L g1908 ( 
.A(n_1484),
.B(n_1352),
.Y(n_1908)
);

AND2x2_ASAP7_75t_L g1909 ( 
.A(n_1592),
.B(n_1353),
.Y(n_1909)
);

AOI22xp5_ASAP7_75t_L g1910 ( 
.A1(n_1536),
.A2(n_1357),
.B1(n_1374),
.B2(n_1365),
.Y(n_1910)
);

INVx2_ASAP7_75t_L g1911 ( 
.A(n_1641),
.Y(n_1911)
);

INVx2_ASAP7_75t_L g1912 ( 
.A(n_1643),
.Y(n_1912)
);

AOI22xp5_ASAP7_75t_L g1913 ( 
.A1(n_1627),
.A2(n_1357),
.B1(n_1374),
.B2(n_1365),
.Y(n_1913)
);

INVx1_ASAP7_75t_L g1914 ( 
.A(n_1426),
.Y(n_1914)
);

BUFx6f_ASAP7_75t_L g1915 ( 
.A(n_1474),
.Y(n_1915)
);

AOI22xp5_ASAP7_75t_L g1916 ( 
.A1(n_1627),
.A2(n_1378),
.B1(n_1384),
.B2(n_1382),
.Y(n_1916)
);

OA21x2_ASAP7_75t_L g1917 ( 
.A1(n_1504),
.A2(n_1167),
.B(n_1161),
.Y(n_1917)
);

NAND2xp33_ASAP7_75t_L g1918 ( 
.A(n_1504),
.B(n_1378),
.Y(n_1918)
);

AND2x4_ASAP7_75t_L g1919 ( 
.A(n_1481),
.B(n_1099),
.Y(n_1919)
);

INVx2_ASAP7_75t_L g1920 ( 
.A(n_1418),
.Y(n_1920)
);

CKINVDCx5p33_ASAP7_75t_R g1921 ( 
.A(n_1667),
.Y(n_1921)
);

AOI22xp5_ASAP7_75t_L g1922 ( 
.A1(n_1647),
.A2(n_1382),
.B1(n_1384),
.B2(n_1219),
.Y(n_1922)
);

INVx1_ASAP7_75t_L g1923 ( 
.A(n_1509),
.Y(n_1923)
);

INVx2_ASAP7_75t_L g1924 ( 
.A(n_1422),
.Y(n_1924)
);

HB1xp67_ASAP7_75t_L g1925 ( 
.A(n_1510),
.Y(n_1925)
);

NOR2xp33_ASAP7_75t_L g1926 ( 
.A(n_1647),
.B(n_1393),
.Y(n_1926)
);

BUFx6f_ASAP7_75t_L g1927 ( 
.A(n_1422),
.Y(n_1927)
);

BUFx6f_ASAP7_75t_L g1928 ( 
.A(n_1515),
.Y(n_1928)
);

INVx1_ASAP7_75t_L g1929 ( 
.A(n_1517),
.Y(n_1929)
);

INVx1_ASAP7_75t_L g1930 ( 
.A(n_1519),
.Y(n_1930)
);

INVx1_ASAP7_75t_L g1931 ( 
.A(n_1621),
.Y(n_1931)
);

INVx2_ASAP7_75t_L g1932 ( 
.A(n_1427),
.Y(n_1932)
);

BUFx8_ASAP7_75t_L g1933 ( 
.A(n_1630),
.Y(n_1933)
);

INVx1_ASAP7_75t_L g1934 ( 
.A(n_1662),
.Y(n_1934)
);

INVx3_ASAP7_75t_L g1935 ( 
.A(n_1427),
.Y(n_1935)
);

NAND2xp5_ASAP7_75t_SL g1936 ( 
.A(n_1428),
.B(n_1280),
.Y(n_1936)
);

OAI21x1_ASAP7_75t_L g1937 ( 
.A1(n_1665),
.A2(n_1395),
.B(n_1394),
.Y(n_1937)
);

NAND2xp5_ASAP7_75t_L g1938 ( 
.A(n_1428),
.B(n_1208),
.Y(n_1938)
);

INVx2_ASAP7_75t_L g1939 ( 
.A(n_1435),
.Y(n_1939)
);

AOI22xp5_ASAP7_75t_L g1940 ( 
.A1(n_1665),
.A2(n_1396),
.B1(n_1397),
.B2(n_1361),
.Y(n_1940)
);

OA21x2_ASAP7_75t_L g1941 ( 
.A1(n_1505),
.A2(n_1172),
.B(n_1170),
.Y(n_1941)
);

INVx3_ASAP7_75t_L g1942 ( 
.A(n_1435),
.Y(n_1942)
);

INVx4_ASAP7_75t_L g1943 ( 
.A(n_1436),
.Y(n_1943)
);

HB1xp67_ASAP7_75t_L g1944 ( 
.A(n_1675),
.Y(n_1944)
);

INVx1_ASAP7_75t_L g1945 ( 
.A(n_1677),
.Y(n_1945)
);

BUFx6f_ASAP7_75t_L g1946 ( 
.A(n_1678),
.Y(n_1946)
);

NAND2xp5_ASAP7_75t_SL g1947 ( 
.A(n_1436),
.B(n_1280),
.Y(n_1947)
);

INVx1_ASAP7_75t_L g1948 ( 
.A(n_1505),
.Y(n_1948)
);

AND2x4_ASAP7_75t_L g1949 ( 
.A(n_1439),
.B(n_1101),
.Y(n_1949)
);

INVx2_ASAP7_75t_L g1950 ( 
.A(n_1439),
.Y(n_1950)
);

INVx3_ASAP7_75t_L g1951 ( 
.A(n_1449),
.Y(n_1951)
);

OAI21x1_ASAP7_75t_L g1952 ( 
.A1(n_1463),
.A2(n_1348),
.B(n_1282),
.Y(n_1952)
);

INVx2_ASAP7_75t_L g1953 ( 
.A(n_1449),
.Y(n_1953)
);

AND2x2_ASAP7_75t_L g1954 ( 
.A(n_1451),
.B(n_1280),
.Y(n_1954)
);

BUFx6f_ASAP7_75t_L g1955 ( 
.A(n_1451),
.Y(n_1955)
);

INVx1_ASAP7_75t_L g1956 ( 
.A(n_1521),
.Y(n_1956)
);

NAND2x1_ASAP7_75t_L g1957 ( 
.A(n_1463),
.B(n_1208),
.Y(n_1957)
);

OA21x2_ASAP7_75t_L g1958 ( 
.A1(n_1521),
.A2(n_1333),
.B(n_1331),
.Y(n_1958)
);

INVx5_ASAP7_75t_L g1959 ( 
.A(n_1700),
.Y(n_1959)
);

AND2x4_ASAP7_75t_L g1960 ( 
.A(n_1452),
.B(n_1105),
.Y(n_1960)
);

AND2x2_ASAP7_75t_SL g1961 ( 
.A(n_1666),
.B(n_1238),
.Y(n_1961)
);

INVx6_ASAP7_75t_L g1962 ( 
.A(n_1694),
.Y(n_1962)
);

INVx3_ASAP7_75t_L g1963 ( 
.A(n_1452),
.Y(n_1963)
);

NAND2xp5_ASAP7_75t_L g1964 ( 
.A(n_1455),
.B(n_1222),
.Y(n_1964)
);

BUFx6f_ASAP7_75t_L g1965 ( 
.A(n_1455),
.Y(n_1965)
);

INVx3_ASAP7_75t_L g1966 ( 
.A(n_1459),
.Y(n_1966)
);

BUFx6f_ASAP7_75t_L g1967 ( 
.A(n_1459),
.Y(n_1967)
);

BUFx6f_ASAP7_75t_L g1968 ( 
.A(n_1466),
.Y(n_1968)
);

INVx1_ASAP7_75t_L g1969 ( 
.A(n_1524),
.Y(n_1969)
);

AND2x4_ASAP7_75t_L g1970 ( 
.A(n_1466),
.B(n_1106),
.Y(n_1970)
);

AND2x4_ASAP7_75t_L g1971 ( 
.A(n_1467),
.B(n_1107),
.Y(n_1971)
);

NOR2x1_ASAP7_75t_L g1972 ( 
.A(n_1687),
.B(n_1124),
.Y(n_1972)
);

OAI22xp5_ASAP7_75t_L g1973 ( 
.A1(n_1407),
.A2(n_1242),
.B1(n_1326),
.B2(n_1173),
.Y(n_1973)
);

INVx2_ASAP7_75t_L g1974 ( 
.A(n_1467),
.Y(n_1974)
);

INVx1_ASAP7_75t_L g1975 ( 
.A(n_1524),
.Y(n_1975)
);

NAND2xp5_ASAP7_75t_L g1976 ( 
.A(n_1486),
.B(n_1222),
.Y(n_1976)
);

NAND2xp5_ASAP7_75t_L g1977 ( 
.A(n_1486),
.B(n_1222),
.Y(n_1977)
);

NAND2xp5_ASAP7_75t_SL g1978 ( 
.A(n_1494),
.B(n_1237),
.Y(n_1978)
);

NOR2x1_ASAP7_75t_L g1979 ( 
.A(n_1409),
.B(n_1206),
.Y(n_1979)
);

NOR2xp33_ASAP7_75t_L g1980 ( 
.A(n_1494),
.B(n_1361),
.Y(n_1980)
);

AND2x4_ASAP7_75t_L g1981 ( 
.A(n_1495),
.B(n_1108),
.Y(n_1981)
);

HB1xp67_ASAP7_75t_L g1982 ( 
.A(n_1525),
.Y(n_1982)
);

BUFx6f_ASAP7_75t_L g1983 ( 
.A(n_1495),
.Y(n_1983)
);

INVx2_ASAP7_75t_L g1984 ( 
.A(n_1502),
.Y(n_1984)
);

BUFx3_ASAP7_75t_L g1985 ( 
.A(n_1502),
.Y(n_1985)
);

INVx2_ASAP7_75t_L g1986 ( 
.A(n_1525),
.Y(n_1986)
);

INVx1_ASAP7_75t_L g1987 ( 
.A(n_1526),
.Y(n_1987)
);

INVx2_ASAP7_75t_L g1988 ( 
.A(n_1526),
.Y(n_1988)
);

INVx1_ASAP7_75t_L g1989 ( 
.A(n_1530),
.Y(n_1989)
);

AOI22xp5_ASAP7_75t_L g1990 ( 
.A1(n_1530),
.A2(n_1091),
.B1(n_1051),
.B2(n_1231),
.Y(n_1990)
);

INVx1_ASAP7_75t_L g1991 ( 
.A(n_1531),
.Y(n_1991)
);

AND2x4_ASAP7_75t_L g1992 ( 
.A(n_1531),
.B(n_1111),
.Y(n_1992)
);

NAND2xp5_ASAP7_75t_L g1993 ( 
.A(n_1532),
.B(n_1222),
.Y(n_1993)
);

INVx2_ASAP7_75t_L g1994 ( 
.A(n_1879),
.Y(n_1994)
);

INVx1_ASAP7_75t_L g1995 ( 
.A(n_1879),
.Y(n_1995)
);

OAI22xp33_ASAP7_75t_SL g1996 ( 
.A1(n_1774),
.A2(n_1533),
.B1(n_1539),
.B2(n_1532),
.Y(n_1996)
);

AND2x2_ASAP7_75t_SL g1997 ( 
.A(n_1961),
.B(n_1120),
.Y(n_1997)
);

INVx1_ASAP7_75t_L g1998 ( 
.A(n_1879),
.Y(n_1998)
);

AND2x2_ASAP7_75t_SL g1999 ( 
.A(n_1961),
.B(n_1053),
.Y(n_1999)
);

AND2x2_ASAP7_75t_L g2000 ( 
.A(n_1748),
.B(n_1533),
.Y(n_2000)
);

BUFx3_ASAP7_75t_L g2001 ( 
.A(n_1738),
.Y(n_2001)
);

NAND2xp33_ASAP7_75t_SL g2002 ( 
.A(n_1843),
.B(n_1539),
.Y(n_2002)
);

INVx1_ASAP7_75t_L g2003 ( 
.A(n_1869),
.Y(n_2003)
);

AOI22xp5_ASAP7_75t_L g2004 ( 
.A1(n_1774),
.A2(n_1546),
.B1(n_1550),
.B2(n_1548),
.Y(n_2004)
);

OR2x2_ASAP7_75t_L g2005 ( 
.A(n_1731),
.B(n_1637),
.Y(n_2005)
);

AOI22xp5_ASAP7_75t_L g2006 ( 
.A1(n_1736),
.A2(n_1546),
.B1(n_1550),
.B2(n_1548),
.Y(n_2006)
);

OR2x2_ASAP7_75t_L g2007 ( 
.A(n_1723),
.B(n_1749),
.Y(n_2007)
);

OAI22xp33_ASAP7_75t_SL g2008 ( 
.A1(n_1839),
.A2(n_1557),
.B1(n_1559),
.B2(n_1556),
.Y(n_2008)
);

AOI22xp5_ASAP7_75t_L g2009 ( 
.A1(n_1736),
.A2(n_1556),
.B1(n_1559),
.B2(n_1557),
.Y(n_2009)
);

AND2x2_ASAP7_75t_L g2010 ( 
.A(n_1729),
.B(n_1561),
.Y(n_2010)
);

OAI22xp33_ASAP7_75t_L g2011 ( 
.A1(n_1829),
.A2(n_1561),
.B1(n_1588),
.B2(n_1582),
.Y(n_2011)
);

OAI22xp33_ASAP7_75t_SL g2012 ( 
.A1(n_1897),
.A2(n_1588),
.B1(n_1590),
.B2(n_1582),
.Y(n_2012)
);

INVx8_ASAP7_75t_L g2013 ( 
.A(n_1959),
.Y(n_2013)
);

OAI22xp33_ASAP7_75t_SL g2014 ( 
.A1(n_1861),
.A2(n_1591),
.B1(n_1593),
.B2(n_1590),
.Y(n_2014)
);

NOR2xp33_ASAP7_75t_L g2015 ( 
.A(n_1783),
.B(n_1591),
.Y(n_2015)
);

NOR2xp33_ASAP7_75t_L g2016 ( 
.A(n_1783),
.B(n_1593),
.Y(n_2016)
);

AO22x2_ASAP7_75t_L g2017 ( 
.A1(n_1973),
.A2(n_844),
.B1(n_849),
.B2(n_836),
.Y(n_2017)
);

INVx1_ASAP7_75t_L g2018 ( 
.A(n_1869),
.Y(n_2018)
);

NOR2xp33_ASAP7_75t_L g2019 ( 
.A(n_1816),
.B(n_1926),
.Y(n_2019)
);

AND2x2_ASAP7_75t_L g2020 ( 
.A(n_1749),
.B(n_1596),
.Y(n_2020)
);

NAND2xp5_ASAP7_75t_L g2021 ( 
.A(n_1795),
.B(n_1803),
.Y(n_2021)
);

OAI22xp33_ASAP7_75t_SL g2022 ( 
.A1(n_1861),
.A2(n_1597),
.B1(n_1604),
.B2(n_1596),
.Y(n_2022)
);

AO22x2_ASAP7_75t_L g2023 ( 
.A1(n_1733),
.A2(n_983),
.B1(n_1266),
.B2(n_1257),
.Y(n_2023)
);

NAND2xp33_ASAP7_75t_SL g2024 ( 
.A(n_1954),
.B(n_1597),
.Y(n_2024)
);

INVx1_ASAP7_75t_L g2025 ( 
.A(n_1756),
.Y(n_2025)
);

BUFx2_ASAP7_75t_L g2026 ( 
.A(n_1745),
.Y(n_2026)
);

OR2x2_ASAP7_75t_L g2027 ( 
.A(n_1993),
.B(n_1657),
.Y(n_2027)
);

INVx1_ASAP7_75t_L g2028 ( 
.A(n_1756),
.Y(n_2028)
);

OR2x2_ASAP7_75t_L g2029 ( 
.A(n_1904),
.B(n_1657),
.Y(n_2029)
);

OA22x2_ASAP7_75t_L g2030 ( 
.A1(n_1940),
.A2(n_1308),
.B1(n_1606),
.B2(n_1604),
.Y(n_2030)
);

OAI22xp33_ASAP7_75t_L g2031 ( 
.A1(n_1761),
.A2(n_1606),
.B1(n_1609),
.B2(n_1608),
.Y(n_2031)
);

NAND3x1_ASAP7_75t_L g2032 ( 
.A(n_1979),
.B(n_1349),
.C(n_1125),
.Y(n_2032)
);

OAI22xp5_ASAP7_75t_SL g2033 ( 
.A1(n_1764),
.A2(n_1695),
.B1(n_1689),
.B2(n_1432),
.Y(n_2033)
);

INVx1_ASAP7_75t_L g2034 ( 
.A(n_1869),
.Y(n_2034)
);

AOI22xp5_ASAP7_75t_L g2035 ( 
.A1(n_1795),
.A2(n_1803),
.B1(n_1836),
.B2(n_1814),
.Y(n_2035)
);

AND2x2_ASAP7_75t_L g2036 ( 
.A(n_1846),
.B(n_1908),
.Y(n_2036)
);

AND2x2_ASAP7_75t_L g2037 ( 
.A(n_1909),
.B(n_1608),
.Y(n_2037)
);

AND2x2_ASAP7_75t_L g2038 ( 
.A(n_1980),
.B(n_1609),
.Y(n_2038)
);

AND2x2_ASAP7_75t_L g2039 ( 
.A(n_1980),
.B(n_1620),
.Y(n_2039)
);

OAI22xp5_ASAP7_75t_SL g2040 ( 
.A1(n_1899),
.A2(n_1433),
.B1(n_1438),
.B2(n_1421),
.Y(n_2040)
);

AO22x2_ASAP7_75t_L g2041 ( 
.A1(n_1800),
.A2(n_1207),
.B1(n_1316),
.B2(n_1304),
.Y(n_2041)
);

OAI22xp33_ASAP7_75t_L g2042 ( 
.A1(n_1730),
.A2(n_1620),
.B1(n_1646),
.B2(n_1637),
.Y(n_2042)
);

INVx2_ASAP7_75t_L g2043 ( 
.A(n_1849),
.Y(n_2043)
);

OAI22xp33_ASAP7_75t_SL g2044 ( 
.A1(n_1978),
.A2(n_1648),
.B1(n_1656),
.B2(n_1646),
.Y(n_2044)
);

AOI22x1_ASAP7_75t_SL g2045 ( 
.A1(n_1899),
.A2(n_1443),
.B1(n_1476),
.B2(n_1445),
.Y(n_2045)
);

AND2x2_ASAP7_75t_L g2046 ( 
.A(n_1785),
.B(n_1648),
.Y(n_2046)
);

NAND2xp5_ASAP7_75t_SL g2047 ( 
.A(n_1949),
.B(n_1656),
.Y(n_2047)
);

OAI22xp5_ASAP7_75t_SL g2048 ( 
.A1(n_1837),
.A2(n_1500),
.B1(n_1501),
.B2(n_1482),
.Y(n_2048)
);

AND2x2_ASAP7_75t_L g2049 ( 
.A(n_1773),
.B(n_1658),
.Y(n_2049)
);

INVx1_ASAP7_75t_L g2050 ( 
.A(n_1895),
.Y(n_2050)
);

OAI22xp5_ASAP7_75t_SL g2051 ( 
.A1(n_1862),
.A2(n_1529),
.B1(n_1534),
.B2(n_1507),
.Y(n_2051)
);

INVx1_ASAP7_75t_L g2052 ( 
.A(n_1895),
.Y(n_2052)
);

INVx2_ASAP7_75t_L g2053 ( 
.A(n_1849),
.Y(n_2053)
);

OAI22xp33_ASAP7_75t_SL g2054 ( 
.A1(n_1978),
.A2(n_1816),
.B1(n_1964),
.B2(n_1938),
.Y(n_2054)
);

BUFx6f_ASAP7_75t_L g2055 ( 
.A(n_1738),
.Y(n_2055)
);

AND2x2_ASAP7_75t_SL g2056 ( 
.A(n_1918),
.B(n_1136),
.Y(n_2056)
);

AND2x2_ASAP7_75t_L g2057 ( 
.A(n_1773),
.B(n_1658),
.Y(n_2057)
);

NOR2xp33_ASAP7_75t_L g2058 ( 
.A(n_1926),
.B(n_1679),
.Y(n_2058)
);

AOI22xp5_ASAP7_75t_L g2059 ( 
.A1(n_1795),
.A2(n_1681),
.B1(n_1686),
.B2(n_1679),
.Y(n_2059)
);

OAI22xp33_ASAP7_75t_L g2060 ( 
.A1(n_1735),
.A2(n_1681),
.B1(n_1693),
.B2(n_1686),
.Y(n_2060)
);

OR2x2_ASAP7_75t_L g2061 ( 
.A(n_1904),
.B(n_1693),
.Y(n_2061)
);

CKINVDCx5p33_ASAP7_75t_R g2062 ( 
.A(n_1915),
.Y(n_2062)
);

INVx1_ASAP7_75t_L g2063 ( 
.A(n_1901),
.Y(n_2063)
);

AO22x1_ASAP7_75t_L g2064 ( 
.A1(n_1992),
.A2(n_1698),
.B1(n_1699),
.B2(n_1408),
.Y(n_2064)
);

AND2x2_ASAP7_75t_L g2065 ( 
.A(n_1818),
.B(n_1698),
.Y(n_2065)
);

BUFx6f_ASAP7_75t_L g2066 ( 
.A(n_1779),
.Y(n_2066)
);

NAND2xp5_ASAP7_75t_L g2067 ( 
.A(n_1795),
.B(n_1699),
.Y(n_2067)
);

INVx2_ASAP7_75t_L g2068 ( 
.A(n_1707),
.Y(n_2068)
);

AO22x1_ASAP7_75t_SL g2069 ( 
.A1(n_1948),
.A2(n_1127),
.B1(n_1132),
.B2(n_1115),
.Y(n_2069)
);

INVx2_ASAP7_75t_L g2070 ( 
.A(n_1707),
.Y(n_2070)
);

OAI22xp33_ASAP7_75t_L g2071 ( 
.A1(n_1705),
.A2(n_1408),
.B1(n_1405),
.B2(n_1338),
.Y(n_2071)
);

OAI22xp33_ASAP7_75t_L g2072 ( 
.A1(n_1712),
.A2(n_1405),
.B1(n_1278),
.B2(n_1304),
.Y(n_2072)
);

INVx2_ASAP7_75t_L g2073 ( 
.A(n_1708),
.Y(n_2073)
);

AND2x2_ASAP7_75t_L g2074 ( 
.A(n_1992),
.B(n_1207),
.Y(n_2074)
);

OAI22xp5_ASAP7_75t_SL g2075 ( 
.A1(n_1898),
.A2(n_1535),
.B1(n_1540),
.B2(n_1538),
.Y(n_2075)
);

INVx2_ASAP7_75t_L g2076 ( 
.A(n_1708),
.Y(n_2076)
);

OAI22xp5_ASAP7_75t_SL g2077 ( 
.A1(n_1824),
.A2(n_1542),
.B1(n_1560),
.B2(n_1553),
.Y(n_2077)
);

NAND2xp5_ASAP7_75t_L g2078 ( 
.A(n_1795),
.B(n_1263),
.Y(n_2078)
);

AND2x2_ASAP7_75t_L g2079 ( 
.A(n_1992),
.B(n_1316),
.Y(n_2079)
);

AOI22xp5_ASAP7_75t_L g2080 ( 
.A1(n_1803),
.A2(n_1113),
.B1(n_1135),
.B2(n_1133),
.Y(n_2080)
);

XOR2xp5_ASAP7_75t_L g2081 ( 
.A(n_1824),
.B(n_1570),
.Y(n_2081)
);

INVx3_ASAP7_75t_L g2082 ( 
.A(n_1747),
.Y(n_2082)
);

OAI22xp33_ASAP7_75t_SL g2083 ( 
.A1(n_1976),
.A2(n_720),
.B1(n_722),
.B2(n_712),
.Y(n_2083)
);

CKINVDCx5p33_ASAP7_75t_R g2084 ( 
.A(n_1915),
.Y(n_2084)
);

AOI22xp5_ASAP7_75t_L g2085 ( 
.A1(n_1803),
.A2(n_1139),
.B1(n_1275),
.B2(n_1263),
.Y(n_2085)
);

OAI22xp5_ASAP7_75t_SL g2086 ( 
.A1(n_1885),
.A2(n_1579),
.B1(n_1585),
.B2(n_1584),
.Y(n_2086)
);

OAI22xp33_ASAP7_75t_L g2087 ( 
.A1(n_1750),
.A2(n_728),
.B1(n_731),
.B2(n_722),
.Y(n_2087)
);

INVx1_ASAP7_75t_L g2088 ( 
.A(n_1901),
.Y(n_2088)
);

AOI22xp5_ASAP7_75t_L g2089 ( 
.A1(n_1803),
.A2(n_1275),
.B1(n_1263),
.B2(n_1334),
.Y(n_2089)
);

OAI22xp33_ASAP7_75t_L g2090 ( 
.A1(n_1709),
.A2(n_731),
.B1(n_732),
.B2(n_728),
.Y(n_2090)
);

AOI22xp5_ASAP7_75t_L g2091 ( 
.A1(n_1814),
.A2(n_1275),
.B1(n_1263),
.B2(n_1337),
.Y(n_2091)
);

OAI22xp33_ASAP7_75t_L g2092 ( 
.A1(n_1716),
.A2(n_733),
.B1(n_734),
.B2(n_732),
.Y(n_2092)
);

OA22x2_ASAP7_75t_L g2093 ( 
.A1(n_1990),
.A2(n_752),
.B1(n_766),
.B2(n_740),
.Y(n_2093)
);

BUFx6f_ASAP7_75t_SL g2094 ( 
.A(n_1915),
.Y(n_2094)
);

AOI22xp5_ASAP7_75t_L g2095 ( 
.A1(n_1814),
.A2(n_1275),
.B1(n_1341),
.B2(n_1339),
.Y(n_2095)
);

AOI22xp5_ASAP7_75t_L g2096 ( 
.A1(n_1814),
.A2(n_1343),
.B1(n_1345),
.B2(n_1342),
.Y(n_2096)
);

OAI22xp33_ASAP7_75t_L g2097 ( 
.A1(n_1958),
.A2(n_734),
.B1(n_737),
.B2(n_733),
.Y(n_2097)
);

BUFx2_ASAP7_75t_L g2098 ( 
.A(n_1949),
.Y(n_2098)
);

OAI22xp33_ASAP7_75t_SL g2099 ( 
.A1(n_1977),
.A2(n_740),
.B1(n_741),
.B2(n_737),
.Y(n_2099)
);

OAI22xp33_ASAP7_75t_SL g2100 ( 
.A1(n_1880),
.A2(n_742),
.B1(n_745),
.B2(n_741),
.Y(n_2100)
);

INVx2_ASAP7_75t_L g2101 ( 
.A(n_1711),
.Y(n_2101)
);

BUFx6f_ASAP7_75t_L g2102 ( 
.A(n_1779),
.Y(n_2102)
);

INVx1_ASAP7_75t_L g2103 ( 
.A(n_1798),
.Y(n_2103)
);

NOR2xp33_ASAP7_75t_L g2104 ( 
.A(n_1903),
.B(n_1586),
.Y(n_2104)
);

OAI22xp33_ASAP7_75t_SL g2105 ( 
.A1(n_1772),
.A2(n_745),
.B1(n_746),
.B2(n_742),
.Y(n_2105)
);

OAI22xp33_ASAP7_75t_L g2106 ( 
.A1(n_1958),
.A2(n_747),
.B1(n_749),
.B2(n_746),
.Y(n_2106)
);

AND2x2_ASAP7_75t_SL g2107 ( 
.A(n_1918),
.B(n_1350),
.Y(n_2107)
);

AOI22xp5_ASAP7_75t_L g2108 ( 
.A1(n_1814),
.A2(n_1346),
.B1(n_1197),
.B2(n_1199),
.Y(n_2108)
);

OR2x6_ASAP7_75t_L g2109 ( 
.A(n_1891),
.B(n_1350),
.Y(n_2109)
);

OAI22xp33_ASAP7_75t_SL g2110 ( 
.A1(n_1778),
.A2(n_749),
.B1(n_751),
.B2(n_747),
.Y(n_2110)
);

INVx2_ASAP7_75t_L g2111 ( 
.A(n_1711),
.Y(n_2111)
);

AND2x2_ASAP7_75t_L g2112 ( 
.A(n_1949),
.B(n_1350),
.Y(n_2112)
);

AND2x2_ASAP7_75t_L g2113 ( 
.A(n_1960),
.B(n_1196),
.Y(n_2113)
);

AOI22xp5_ASAP7_75t_L g2114 ( 
.A1(n_1836),
.A2(n_1202),
.B1(n_752),
.B2(n_753),
.Y(n_2114)
);

OAI22xp33_ASAP7_75t_L g2115 ( 
.A1(n_1958),
.A2(n_753),
.B1(n_755),
.B2(n_751),
.Y(n_2115)
);

OAI22xp33_ASAP7_75t_L g2116 ( 
.A1(n_1917),
.A2(n_1941),
.B1(n_1863),
.B2(n_1868),
.Y(n_2116)
);

AND2x2_ASAP7_75t_L g2117 ( 
.A(n_1960),
.B(n_1412),
.Y(n_2117)
);

AND2x2_ASAP7_75t_L g2118 ( 
.A(n_1960),
.B(n_1412),
.Y(n_2118)
);

NOR2xp33_ASAP7_75t_L g2119 ( 
.A(n_1787),
.B(n_1601),
.Y(n_2119)
);

AOI22xp5_ASAP7_75t_L g2120 ( 
.A1(n_1836),
.A2(n_756),
.B1(n_758),
.B2(n_755),
.Y(n_2120)
);

OAI22xp33_ASAP7_75t_SL g2121 ( 
.A1(n_1781),
.A2(n_1790),
.B1(n_1794),
.B2(n_1788),
.Y(n_2121)
);

OAI22xp5_ASAP7_75t_SL g2122 ( 
.A1(n_1885),
.A2(n_1616),
.B1(n_1618),
.B2(n_1615),
.Y(n_2122)
);

INVx8_ASAP7_75t_L g2123 ( 
.A(n_1959),
.Y(n_2123)
);

INVx8_ASAP7_75t_L g2124 ( 
.A(n_1959),
.Y(n_2124)
);

INVx1_ASAP7_75t_L g2125 ( 
.A(n_1798),
.Y(n_2125)
);

INVx1_ASAP7_75t_L g2126 ( 
.A(n_1756),
.Y(n_2126)
);

AND2x2_ASAP7_75t_SL g2127 ( 
.A(n_1927),
.B(n_1623),
.Y(n_2127)
);

AND2x2_ASAP7_75t_L g2128 ( 
.A(n_1970),
.B(n_1635),
.Y(n_2128)
);

OR2x2_ASAP7_75t_L g2129 ( 
.A(n_1906),
.B(n_1023),
.Y(n_2129)
);

AOI22xp5_ASAP7_75t_L g2130 ( 
.A1(n_1836),
.A2(n_758),
.B1(n_760),
.B2(n_756),
.Y(n_2130)
);

NAND2xp5_ASAP7_75t_L g2131 ( 
.A(n_1836),
.B(n_760),
.Y(n_2131)
);

NOR2xp33_ASAP7_75t_L g2132 ( 
.A(n_1801),
.B(n_1741),
.Y(n_2132)
);

AND2x2_ASAP7_75t_SL g2133 ( 
.A(n_1927),
.B(n_764),
.Y(n_2133)
);

BUFx4f_ASAP7_75t_L g2134 ( 
.A(n_1891),
.Y(n_2134)
);

OAI22xp33_ASAP7_75t_SL g2135 ( 
.A1(n_1796),
.A2(n_765),
.B1(n_766),
.B2(n_764),
.Y(n_2135)
);

AOI22xp5_ASAP7_75t_L g2136 ( 
.A1(n_1917),
.A2(n_975),
.B1(n_976),
.B2(n_765),
.Y(n_2136)
);

CKINVDCx5p33_ASAP7_75t_R g2137 ( 
.A(n_1915),
.Y(n_2137)
);

OAI22xp33_ASAP7_75t_L g2138 ( 
.A1(n_1917),
.A2(n_976),
.B1(n_978),
.B2(n_975),
.Y(n_2138)
);

INVx1_ASAP7_75t_L g2139 ( 
.A(n_1784),
.Y(n_2139)
);

INVx1_ASAP7_75t_SL g2140 ( 
.A(n_1891),
.Y(n_2140)
);

AO22x2_ASAP7_75t_L g2141 ( 
.A1(n_1857),
.A2(n_7),
.B1(n_5),
.B2(n_6),
.Y(n_2141)
);

AOI22xp5_ASAP7_75t_L g2142 ( 
.A1(n_1941),
.A2(n_979),
.B1(n_986),
.B2(n_978),
.Y(n_2142)
);

OAI22xp33_ASAP7_75t_L g2143 ( 
.A1(n_1941),
.A2(n_986),
.B1(n_991),
.B2(n_979),
.Y(n_2143)
);

AOI22xp5_ASAP7_75t_L g2144 ( 
.A1(n_1970),
.A2(n_999),
.B1(n_1000),
.B2(n_991),
.Y(n_2144)
);

AO22x2_ASAP7_75t_L g2145 ( 
.A1(n_1739),
.A2(n_1905),
.B1(n_1988),
.B2(n_1986),
.Y(n_2145)
);

XNOR2xp5_ASAP7_75t_L g2146 ( 
.A(n_1762),
.B(n_999),
.Y(n_2146)
);

OAI22xp33_ASAP7_75t_SL g2147 ( 
.A1(n_1810),
.A2(n_1002),
.B1(n_1003),
.B2(n_1000),
.Y(n_2147)
);

AND2x2_ASAP7_75t_L g2148 ( 
.A(n_1970),
.B(n_1002),
.Y(n_2148)
);

INVx2_ASAP7_75t_L g2149 ( 
.A(n_1713),
.Y(n_2149)
);

AND2x2_ASAP7_75t_L g2150 ( 
.A(n_1971),
.B(n_1003),
.Y(n_2150)
);

AND2x2_ASAP7_75t_L g2151 ( 
.A(n_1971),
.B(n_1005),
.Y(n_2151)
);

AND2x2_ASAP7_75t_L g2152 ( 
.A(n_1971),
.B(n_1005),
.Y(n_2152)
);

AND2x2_ASAP7_75t_L g2153 ( 
.A(n_1981),
.B(n_1006),
.Y(n_2153)
);

AOI22xp5_ASAP7_75t_L g2154 ( 
.A1(n_1981),
.A2(n_1007),
.B1(n_1008),
.B2(n_1006),
.Y(n_2154)
);

BUFx6f_ASAP7_75t_L g2155 ( 
.A(n_1758),
.Y(n_2155)
);

INVx1_ASAP7_75t_L g2156 ( 
.A(n_1784),
.Y(n_2156)
);

OR2x2_ASAP7_75t_L g2157 ( 
.A(n_1906),
.B(n_1007),
.Y(n_2157)
);

AND2x2_ASAP7_75t_L g2158 ( 
.A(n_1981),
.B(n_1008),
.Y(n_2158)
);

INVx2_ASAP7_75t_L g2159 ( 
.A(n_1713),
.Y(n_2159)
);

NAND2xp33_ASAP7_75t_SL g2160 ( 
.A(n_1986),
.B(n_1010),
.Y(n_2160)
);

OR2x6_ASAP7_75t_L g2161 ( 
.A(n_1894),
.B(n_1010),
.Y(n_2161)
);

AND2x2_ASAP7_75t_L g2162 ( 
.A(n_1919),
.B(n_1011),
.Y(n_2162)
);

AOI22xp5_ASAP7_75t_L g2163 ( 
.A1(n_1881),
.A2(n_1012),
.B1(n_1014),
.B2(n_1011),
.Y(n_2163)
);

INVx1_ASAP7_75t_L g2164 ( 
.A(n_1789),
.Y(n_2164)
);

AOI22xp5_ASAP7_75t_L g2165 ( 
.A1(n_1881),
.A2(n_1014),
.B1(n_1015),
.B2(n_1012),
.Y(n_2165)
);

INVx4_ASAP7_75t_L g2166 ( 
.A(n_1808),
.Y(n_2166)
);

INVx1_ASAP7_75t_L g2167 ( 
.A(n_1789),
.Y(n_2167)
);

OAI22xp33_ASAP7_75t_R g2168 ( 
.A1(n_1988),
.A2(n_1907),
.B1(n_1912),
.B2(n_1911),
.Y(n_2168)
);

OR2x6_ASAP7_75t_L g2169 ( 
.A(n_1894),
.B(n_1015),
.Y(n_2169)
);

OAI22xp5_ASAP7_75t_L g2170 ( 
.A1(n_1722),
.A2(n_1019),
.B1(n_1023),
.B2(n_1018),
.Y(n_2170)
);

OAI22xp33_ASAP7_75t_SL g2171 ( 
.A1(n_1815),
.A2(n_1019),
.B1(n_1027),
.B2(n_1018),
.Y(n_2171)
);

NAND2xp33_ASAP7_75t_SL g2172 ( 
.A(n_1768),
.B(n_1027),
.Y(n_2172)
);

OAI22xp33_ASAP7_75t_L g2173 ( 
.A1(n_1866),
.A2(n_1028),
.B1(n_8),
.B2(n_5),
.Y(n_2173)
);

AOI22xp5_ASAP7_75t_L g2174 ( 
.A1(n_1919),
.A2(n_1755),
.B1(n_1753),
.B2(n_1826),
.Y(n_2174)
);

OAI22xp33_ASAP7_75t_SL g2175 ( 
.A1(n_1830),
.A2(n_1028),
.B1(n_9),
.B2(n_6),
.Y(n_2175)
);

NAND2xp5_ASAP7_75t_SL g2176 ( 
.A(n_1919),
.B(n_1859),
.Y(n_2176)
);

INVx2_ASAP7_75t_L g2177 ( 
.A(n_1717),
.Y(n_2177)
);

AOI22xp5_ASAP7_75t_L g2178 ( 
.A1(n_1753),
.A2(n_108),
.B1(n_109),
.B2(n_107),
.Y(n_2178)
);

OAI22xp33_ASAP7_75t_L g2179 ( 
.A1(n_1874),
.A2(n_10),
.B1(n_8),
.B2(n_9),
.Y(n_2179)
);

INVx2_ASAP7_75t_L g2180 ( 
.A(n_1717),
.Y(n_2180)
);

INVx1_ASAP7_75t_L g2181 ( 
.A(n_1813),
.Y(n_2181)
);

AO22x2_ASAP7_75t_L g2182 ( 
.A1(n_1956),
.A2(n_12),
.B1(n_10),
.B2(n_11),
.Y(n_2182)
);

OAI22xp33_ASAP7_75t_SL g2183 ( 
.A1(n_1831),
.A2(n_12),
.B1(n_10),
.B2(n_11),
.Y(n_2183)
);

AND2x2_ASAP7_75t_L g2184 ( 
.A(n_1907),
.B(n_687),
.Y(n_2184)
);

AO22x2_ASAP7_75t_L g2185 ( 
.A1(n_1969),
.A2(n_15),
.B1(n_13),
.B2(n_14),
.Y(n_2185)
);

OAI22xp33_ASAP7_75t_SL g2186 ( 
.A1(n_1832),
.A2(n_15),
.B1(n_13),
.B2(n_14),
.Y(n_2186)
);

OAI22xp33_ASAP7_75t_SL g2187 ( 
.A1(n_1833),
.A2(n_1840),
.B1(n_1841),
.B2(n_1834),
.Y(n_2187)
);

CKINVDCx5p33_ASAP7_75t_R g2188 ( 
.A(n_1838),
.Y(n_2188)
);

INVx2_ASAP7_75t_L g2189 ( 
.A(n_1724),
.Y(n_2189)
);

AOI22xp5_ASAP7_75t_L g2190 ( 
.A1(n_1753),
.A2(n_109),
.B1(n_110),
.B2(n_108),
.Y(n_2190)
);

AO22x2_ASAP7_75t_L g2191 ( 
.A1(n_1975),
.A2(n_16),
.B1(n_13),
.B2(n_14),
.Y(n_2191)
);

OR2x6_ASAP7_75t_L g2192 ( 
.A(n_1894),
.B(n_1962),
.Y(n_2192)
);

AOI22xp5_ASAP7_75t_L g2193 ( 
.A1(n_1755),
.A2(n_112),
.B1(n_113),
.B2(n_110),
.Y(n_2193)
);

BUFx6f_ASAP7_75t_SL g2194 ( 
.A(n_1927),
.Y(n_2194)
);

OAI22xp5_ASAP7_75t_SL g2195 ( 
.A1(n_1987),
.A2(n_24),
.B1(n_32),
.B2(n_16),
.Y(n_2195)
);

AOI22xp5_ASAP7_75t_L g2196 ( 
.A1(n_1755),
.A2(n_113),
.B1(n_114),
.B2(n_112),
.Y(n_2196)
);

INVx1_ASAP7_75t_L g2197 ( 
.A(n_1813),
.Y(n_2197)
);

BUFx10_ASAP7_75t_L g2198 ( 
.A(n_1962),
.Y(n_2198)
);

AO22x2_ASAP7_75t_L g2199 ( 
.A1(n_1989),
.A2(n_18),
.B1(n_16),
.B2(n_17),
.Y(n_2199)
);

INVx2_ASAP7_75t_SL g2200 ( 
.A(n_1758),
.Y(n_2200)
);

AO22x2_ASAP7_75t_L g2201 ( 
.A1(n_1991),
.A2(n_19),
.B1(n_17),
.B2(n_18),
.Y(n_2201)
);

NAND2xp5_ASAP7_75t_SL g2202 ( 
.A(n_1859),
.B(n_17),
.Y(n_2202)
);

AND2x4_ASAP7_75t_L g2203 ( 
.A(n_1758),
.B(n_19),
.Y(n_2203)
);

INVx2_ASAP7_75t_L g2204 ( 
.A(n_1724),
.Y(n_2204)
);

AND2x2_ASAP7_75t_SL g2205 ( 
.A(n_1927),
.B(n_20),
.Y(n_2205)
);

NOR2xp33_ASAP7_75t_L g2206 ( 
.A(n_1850),
.B(n_20),
.Y(n_2206)
);

NOR2xp33_ASAP7_75t_L g2207 ( 
.A(n_1902),
.B(n_21),
.Y(n_2207)
);

INVx1_ASAP7_75t_L g2208 ( 
.A(n_1819),
.Y(n_2208)
);

AND2x2_ASAP7_75t_L g2209 ( 
.A(n_1911),
.B(n_684),
.Y(n_2209)
);

AOI22xp5_ASAP7_75t_L g2210 ( 
.A1(n_1842),
.A2(n_115),
.B1(n_116),
.B2(n_114),
.Y(n_2210)
);

AO22x2_ASAP7_75t_L g2211 ( 
.A1(n_1865),
.A2(n_23),
.B1(n_21),
.B2(n_22),
.Y(n_2211)
);

INVx1_ASAP7_75t_L g2212 ( 
.A(n_1782),
.Y(n_2212)
);

AOI22xp5_ASAP7_75t_L g2213 ( 
.A1(n_1845),
.A2(n_117),
.B1(n_118),
.B2(n_116),
.Y(n_2213)
);

NAND3x1_ASAP7_75t_L g2214 ( 
.A(n_1910),
.B(n_23),
.C(n_24),
.Y(n_2214)
);

OAI22xp33_ASAP7_75t_SL g2215 ( 
.A1(n_1858),
.A2(n_26),
.B1(n_23),
.B2(n_25),
.Y(n_2215)
);

INVx1_ASAP7_75t_SL g2216 ( 
.A(n_1962),
.Y(n_2216)
);

INVx3_ASAP7_75t_L g2217 ( 
.A(n_1747),
.Y(n_2217)
);

OAI22xp33_ASAP7_75t_SL g2218 ( 
.A1(n_1860),
.A2(n_27),
.B1(n_25),
.B2(n_26),
.Y(n_2218)
);

INVx2_ASAP7_75t_L g2219 ( 
.A(n_1727),
.Y(n_2219)
);

INVxp33_ASAP7_75t_L g2220 ( 
.A(n_1878),
.Y(n_2220)
);

INVx2_ASAP7_75t_SL g2221 ( 
.A(n_1782),
.Y(n_2221)
);

OAI22xp33_ASAP7_75t_SL g2222 ( 
.A1(n_1867),
.A2(n_1876),
.B1(n_1888),
.B2(n_1870),
.Y(n_2222)
);

INVx2_ASAP7_75t_L g2223 ( 
.A(n_1727),
.Y(n_2223)
);

OAI22xp33_ASAP7_75t_L g2224 ( 
.A1(n_1874),
.A2(n_28),
.B1(n_26),
.B2(n_27),
.Y(n_2224)
);

AO22x2_ASAP7_75t_L g2225 ( 
.A1(n_1936),
.A2(n_29),
.B1(n_27),
.B2(n_28),
.Y(n_2225)
);

INVx2_ASAP7_75t_L g2226 ( 
.A(n_1734),
.Y(n_2226)
);

OAI22xp5_ASAP7_75t_SL g2227 ( 
.A1(n_1920),
.A2(n_36),
.B1(n_44),
.B2(n_28),
.Y(n_2227)
);

BUFx10_ASAP7_75t_L g2228 ( 
.A(n_1762),
.Y(n_2228)
);

INVx3_ASAP7_75t_L g2229 ( 
.A(n_1747),
.Y(n_2229)
);

AOI22xp5_ASAP7_75t_L g2230 ( 
.A1(n_1893),
.A2(n_120),
.B1(n_121),
.B2(n_117),
.Y(n_2230)
);

INVx2_ASAP7_75t_L g2231 ( 
.A(n_1734),
.Y(n_2231)
);

AND2x2_ASAP7_75t_L g2232 ( 
.A(n_1912),
.B(n_698),
.Y(n_2232)
);

OAI22xp33_ASAP7_75t_SL g2233 ( 
.A1(n_1936),
.A2(n_31),
.B1(n_29),
.B2(n_30),
.Y(n_2233)
);

OAI22xp5_ASAP7_75t_SL g2234 ( 
.A1(n_1920),
.A2(n_38),
.B1(n_46),
.B2(n_30),
.Y(n_2234)
);

NAND2xp5_ASAP7_75t_L g2235 ( 
.A(n_1874),
.B(n_31),
.Y(n_2235)
);

AO22x2_ASAP7_75t_L g2236 ( 
.A1(n_1947),
.A2(n_33),
.B1(n_31),
.B2(n_32),
.Y(n_2236)
);

INVx1_ASAP7_75t_SL g2237 ( 
.A(n_1921),
.Y(n_2237)
);

OAI22xp5_ASAP7_75t_L g2238 ( 
.A1(n_1886),
.A2(n_35),
.B1(n_33),
.B2(n_34),
.Y(n_2238)
);

AOI22xp5_ASAP7_75t_L g2239 ( 
.A1(n_1886),
.A2(n_122),
.B1(n_123),
.B2(n_121),
.Y(n_2239)
);

BUFx6f_ASAP7_75t_SL g2240 ( 
.A(n_1955),
.Y(n_2240)
);

AO22x2_ASAP7_75t_L g2241 ( 
.A1(n_1947),
.A2(n_35),
.B1(n_33),
.B2(n_34),
.Y(n_2241)
);

AOI22xp5_ASAP7_75t_L g2242 ( 
.A1(n_1886),
.A2(n_123),
.B1(n_124),
.B2(n_122),
.Y(n_2242)
);

BUFx10_ASAP7_75t_L g2243 ( 
.A(n_1955),
.Y(n_2243)
);

OAI22xp33_ASAP7_75t_L g2244 ( 
.A1(n_1887),
.A2(n_37),
.B1(n_34),
.B2(n_36),
.Y(n_2244)
);

OAI22xp33_ASAP7_75t_SL g2245 ( 
.A1(n_1718),
.A2(n_39),
.B1(n_37),
.B2(n_38),
.Y(n_2245)
);

INVx2_ASAP7_75t_L g2246 ( 
.A(n_1766),
.Y(n_2246)
);

AOI22xp5_ASAP7_75t_L g2247 ( 
.A1(n_1887),
.A2(n_126),
.B1(n_127),
.B2(n_125),
.Y(n_2247)
);

AND2x2_ASAP7_75t_L g2248 ( 
.A(n_1935),
.B(n_697),
.Y(n_2248)
);

BUFx2_ASAP7_75t_L g2249 ( 
.A(n_1921),
.Y(n_2249)
);

AND2x2_ASAP7_75t_L g2250 ( 
.A(n_1935),
.B(n_697),
.Y(n_2250)
);

AO22x2_ASAP7_75t_L g2251 ( 
.A1(n_1924),
.A2(n_40),
.B1(n_38),
.B2(n_39),
.Y(n_2251)
);

XNOR2xp5_ASAP7_75t_L g2252 ( 
.A(n_1925),
.B(n_39),
.Y(n_2252)
);

OA22x2_ASAP7_75t_L g2253 ( 
.A1(n_1768),
.A2(n_1720),
.B1(n_1922),
.B2(n_1916),
.Y(n_2253)
);

OAI22xp33_ASAP7_75t_R g2254 ( 
.A1(n_1924),
.A2(n_48),
.B1(n_56),
.B2(n_40),
.Y(n_2254)
);

AOI22xp5_ASAP7_75t_L g2255 ( 
.A1(n_1887),
.A2(n_128),
.B1(n_129),
.B2(n_127),
.Y(n_2255)
);

AND2x2_ASAP7_75t_L g2256 ( 
.A(n_1935),
.B(n_685),
.Y(n_2256)
);

AO22x2_ASAP7_75t_L g2257 ( 
.A1(n_1932),
.A2(n_43),
.B1(n_41),
.B2(n_42),
.Y(n_2257)
);

NOR2xp33_ASAP7_75t_L g2258 ( 
.A(n_1913),
.B(n_41),
.Y(n_2258)
);

INVx2_ASAP7_75t_L g2259 ( 
.A(n_1766),
.Y(n_2259)
);

INVx2_ASAP7_75t_L g2260 ( 
.A(n_1769),
.Y(n_2260)
);

NAND2xp5_ASAP7_75t_L g2261 ( 
.A(n_1844),
.B(n_42),
.Y(n_2261)
);

AND2x4_ASAP7_75t_L g2262 ( 
.A(n_1782),
.B(n_43),
.Y(n_2262)
);

AND2x2_ASAP7_75t_L g2263 ( 
.A(n_1942),
.B(n_1951),
.Y(n_2263)
);

AOI22xp5_ASAP7_75t_L g2264 ( 
.A1(n_1884),
.A2(n_129),
.B1(n_130),
.B2(n_128),
.Y(n_2264)
);

AO22x2_ASAP7_75t_L g2265 ( 
.A1(n_1932),
.A2(n_45),
.B1(n_43),
.B2(n_44),
.Y(n_2265)
);

NAND2xp5_ASAP7_75t_L g2266 ( 
.A(n_1844),
.B(n_45),
.Y(n_2266)
);

INVx2_ASAP7_75t_L g2267 ( 
.A(n_1769),
.Y(n_2267)
);

OAI22xp33_ASAP7_75t_L g2268 ( 
.A1(n_1812),
.A2(n_47),
.B1(n_45),
.B2(n_46),
.Y(n_2268)
);

AND2x2_ASAP7_75t_L g2269 ( 
.A(n_1942),
.B(n_692),
.Y(n_2269)
);

NOR2xp33_ASAP7_75t_L g2270 ( 
.A(n_1853),
.B(n_1808),
.Y(n_2270)
);

NAND2xp5_ASAP7_75t_L g2271 ( 
.A(n_1844),
.B(n_46),
.Y(n_2271)
);

OA22x2_ASAP7_75t_L g2272 ( 
.A1(n_1914),
.A2(n_49),
.B1(n_47),
.B2(n_48),
.Y(n_2272)
);

INVx1_ASAP7_75t_L g2273 ( 
.A(n_1819),
.Y(n_2273)
);

INVx1_ASAP7_75t_L g2274 ( 
.A(n_1825),
.Y(n_2274)
);

AOI22xp5_ASAP7_75t_L g2275 ( 
.A1(n_1732),
.A2(n_131),
.B1(n_132),
.B2(n_130),
.Y(n_2275)
);

AOI22xp5_ASAP7_75t_L g2276 ( 
.A1(n_1743),
.A2(n_133),
.B1(n_134),
.B2(n_132),
.Y(n_2276)
);

AND2x2_ASAP7_75t_L g2277 ( 
.A(n_1942),
.B(n_133),
.Y(n_2277)
);

CKINVDCx5p33_ASAP7_75t_R g2278 ( 
.A(n_1838),
.Y(n_2278)
);

OR2x2_ASAP7_75t_L g2279 ( 
.A(n_1883),
.B(n_47),
.Y(n_2279)
);

AO22x2_ASAP7_75t_L g2280 ( 
.A1(n_1939),
.A2(n_50),
.B1(n_48),
.B2(n_49),
.Y(n_2280)
);

OAI22xp33_ASAP7_75t_R g2281 ( 
.A1(n_1939),
.A2(n_57),
.B1(n_65),
.B2(n_49),
.Y(n_2281)
);

AND2x2_ASAP7_75t_L g2282 ( 
.A(n_1951),
.B(n_686),
.Y(n_2282)
);

AND2x6_ASAP7_75t_L g2283 ( 
.A(n_1950),
.B(n_50),
.Y(n_2283)
);

AND2x2_ASAP7_75t_L g2284 ( 
.A(n_1951),
.B(n_688),
.Y(n_2284)
);

AOI22xp5_ASAP7_75t_L g2285 ( 
.A1(n_1746),
.A2(n_136),
.B1(n_137),
.B2(n_135),
.Y(n_2285)
);

AOI22xp5_ASAP7_75t_L g2286 ( 
.A1(n_1752),
.A2(n_136),
.B1(n_137),
.B2(n_135),
.Y(n_2286)
);

INVx2_ASAP7_75t_SL g2287 ( 
.A(n_1793),
.Y(n_2287)
);

INVx1_ASAP7_75t_L g2288 ( 
.A(n_1825),
.Y(n_2288)
);

AO22x2_ASAP7_75t_L g2289 ( 
.A1(n_1950),
.A2(n_53),
.B1(n_51),
.B2(n_52),
.Y(n_2289)
);

AND2x2_ASAP7_75t_L g2290 ( 
.A(n_1963),
.B(n_1966),
.Y(n_2290)
);

AOI22xp5_ASAP7_75t_L g2291 ( 
.A1(n_1759),
.A2(n_140),
.B1(n_141),
.B2(n_138),
.Y(n_2291)
);

AND2x2_ASAP7_75t_L g2292 ( 
.A(n_1963),
.B(n_695),
.Y(n_2292)
);

OAI22xp5_ASAP7_75t_L g2293 ( 
.A1(n_1953),
.A2(n_54),
.B1(n_52),
.B2(n_53),
.Y(n_2293)
);

INVx1_ASAP7_75t_L g2294 ( 
.A(n_1793),
.Y(n_2294)
);

OAI22xp33_ASAP7_75t_L g2295 ( 
.A1(n_1855),
.A2(n_56),
.B1(n_54),
.B2(n_55),
.Y(n_2295)
);

INVx2_ASAP7_75t_L g2296 ( 
.A(n_1847),
.Y(n_2296)
);

AOI22xp5_ASAP7_75t_L g2297 ( 
.A1(n_1763),
.A2(n_142),
.B1(n_143),
.B2(n_141),
.Y(n_2297)
);

OAI22xp33_ASAP7_75t_L g2298 ( 
.A1(n_1855),
.A2(n_1877),
.B1(n_1889),
.B2(n_1873),
.Y(n_2298)
);

INVx4_ASAP7_75t_L g2299 ( 
.A(n_1808),
.Y(n_2299)
);

INVx3_ASAP7_75t_L g2300 ( 
.A(n_1751),
.Y(n_2300)
);

INVx2_ASAP7_75t_SL g2301 ( 
.A(n_1793),
.Y(n_2301)
);

NAND3x1_ASAP7_75t_L g2302 ( 
.A(n_1972),
.B(n_54),
.C(n_55),
.Y(n_2302)
);

AND2x2_ASAP7_75t_L g2303 ( 
.A(n_1963),
.B(n_682),
.Y(n_2303)
);

AND2x2_ASAP7_75t_L g2304 ( 
.A(n_1966),
.B(n_683),
.Y(n_2304)
);

AND2x2_ASAP7_75t_L g2305 ( 
.A(n_1966),
.B(n_683),
.Y(n_2305)
);

NAND3x1_ASAP7_75t_L g2306 ( 
.A(n_1923),
.B(n_55),
.C(n_56),
.Y(n_2306)
);

INVx1_ASAP7_75t_L g2307 ( 
.A(n_1828),
.Y(n_2307)
);

INVx2_ASAP7_75t_L g2308 ( 
.A(n_1847),
.Y(n_2308)
);

AND2x2_ASAP7_75t_L g2309 ( 
.A(n_1953),
.B(n_687),
.Y(n_2309)
);

AND2x2_ASAP7_75t_L g2310 ( 
.A(n_1974),
.B(n_689),
.Y(n_2310)
);

AOI22xp5_ASAP7_75t_L g2311 ( 
.A1(n_1770),
.A2(n_144),
.B1(n_145),
.B2(n_143),
.Y(n_2311)
);

INVx1_ASAP7_75t_L g2312 ( 
.A(n_1828),
.Y(n_2312)
);

AND2x2_ASAP7_75t_L g2313 ( 
.A(n_1974),
.B(n_690),
.Y(n_2313)
);

INVx2_ASAP7_75t_SL g2314 ( 
.A(n_1799),
.Y(n_2314)
);

AND2x6_ASAP7_75t_L g2315 ( 
.A(n_2035),
.B(n_1955),
.Y(n_2315)
);

INVx2_ASAP7_75t_L g2316 ( 
.A(n_1994),
.Y(n_2316)
);

INVx2_ASAP7_75t_L g2317 ( 
.A(n_1995),
.Y(n_2317)
);

INVx3_ASAP7_75t_L g2318 ( 
.A(n_2155),
.Y(n_2318)
);

INVx2_ASAP7_75t_L g2319 ( 
.A(n_1995),
.Y(n_2319)
);

NAND2xp5_ASAP7_75t_SL g2320 ( 
.A(n_2054),
.B(n_1965),
.Y(n_2320)
);

INVx6_ASAP7_75t_L g2321 ( 
.A(n_2198),
.Y(n_2321)
);

INVx2_ASAP7_75t_L g2322 ( 
.A(n_1998),
.Y(n_2322)
);

BUFx6f_ASAP7_75t_L g2323 ( 
.A(n_2155),
.Y(n_2323)
);

INVx2_ASAP7_75t_L g2324 ( 
.A(n_1998),
.Y(n_2324)
);

INVx2_ASAP7_75t_L g2325 ( 
.A(n_2003),
.Y(n_2325)
);

OR2x6_ASAP7_75t_L g2326 ( 
.A(n_2192),
.B(n_1955),
.Y(n_2326)
);

INVx1_ASAP7_75t_L g2327 ( 
.A(n_2025),
.Y(n_2327)
);

OR2x6_ASAP7_75t_L g2328 ( 
.A(n_2192),
.B(n_1965),
.Y(n_2328)
);

INVx2_ASAP7_75t_L g2329 ( 
.A(n_2003),
.Y(n_2329)
);

NAND2xp5_ASAP7_75t_SL g2330 ( 
.A(n_2019),
.B(n_1965),
.Y(n_2330)
);

BUFx10_ASAP7_75t_L g2331 ( 
.A(n_2094),
.Y(n_2331)
);

INVx2_ASAP7_75t_L g2332 ( 
.A(n_2018),
.Y(n_2332)
);

AND2x2_ASAP7_75t_L g2333 ( 
.A(n_2263),
.B(n_1965),
.Y(n_2333)
);

INVx2_ASAP7_75t_L g2334 ( 
.A(n_2018),
.Y(n_2334)
);

BUFx3_ASAP7_75t_L g2335 ( 
.A(n_2198),
.Y(n_2335)
);

CKINVDCx5p33_ASAP7_75t_R g2336 ( 
.A(n_2062),
.Y(n_2336)
);

NAND2xp5_ASAP7_75t_SL g2337 ( 
.A(n_2067),
.B(n_2107),
.Y(n_2337)
);

NAND2xp5_ASAP7_75t_L g2338 ( 
.A(n_2015),
.B(n_1871),
.Y(n_2338)
);

BUFx6f_ASAP7_75t_L g2339 ( 
.A(n_2155),
.Y(n_2339)
);

INVx4_ASAP7_75t_L g2340 ( 
.A(n_2166),
.Y(n_2340)
);

INVx1_ASAP7_75t_L g2341 ( 
.A(n_2028),
.Y(n_2341)
);

INVxp33_ASAP7_75t_SL g2342 ( 
.A(n_2040),
.Y(n_2342)
);

AND2x2_ASAP7_75t_L g2343 ( 
.A(n_2290),
.B(n_1967),
.Y(n_2343)
);

HB1xp67_ASAP7_75t_L g2344 ( 
.A(n_2098),
.Y(n_2344)
);

NAND2xp5_ASAP7_75t_SL g2345 ( 
.A(n_2021),
.B(n_1967),
.Y(n_2345)
);

INVx3_ASAP7_75t_L g2346 ( 
.A(n_2082),
.Y(n_2346)
);

INVx2_ASAP7_75t_SL g2347 ( 
.A(n_2243),
.Y(n_2347)
);

INVx1_ASAP7_75t_L g2348 ( 
.A(n_2126),
.Y(n_2348)
);

NAND2xp5_ASAP7_75t_L g2349 ( 
.A(n_2016),
.B(n_2112),
.Y(n_2349)
);

BUFx3_ASAP7_75t_L g2350 ( 
.A(n_2243),
.Y(n_2350)
);

INVx2_ASAP7_75t_L g2351 ( 
.A(n_2034),
.Y(n_2351)
);

BUFx6f_ASAP7_75t_SL g2352 ( 
.A(n_2127),
.Y(n_2352)
);

CKINVDCx20_ASAP7_75t_R g2353 ( 
.A(n_2077),
.Y(n_2353)
);

NOR3xp33_ASAP7_75t_L g2354 ( 
.A(n_2058),
.B(n_1943),
.C(n_1984),
.Y(n_2354)
);

AND2x4_ASAP7_75t_L g2355 ( 
.A(n_2203),
.B(n_1873),
.Y(n_2355)
);

INVx1_ASAP7_75t_L g2356 ( 
.A(n_2212),
.Y(n_2356)
);

INVx4_ASAP7_75t_L g2357 ( 
.A(n_2166),
.Y(n_2357)
);

NAND2xp5_ASAP7_75t_L g2358 ( 
.A(n_2082),
.B(n_1871),
.Y(n_2358)
);

NAND2xp5_ASAP7_75t_L g2359 ( 
.A(n_2217),
.B(n_1871),
.Y(n_2359)
);

INVx2_ASAP7_75t_L g2360 ( 
.A(n_2034),
.Y(n_2360)
);

NOR2xp33_ASAP7_75t_L g2361 ( 
.A(n_2049),
.B(n_1984),
.Y(n_2361)
);

INVxp33_ASAP7_75t_L g2362 ( 
.A(n_2000),
.Y(n_2362)
);

INVx1_ASAP7_75t_L g2363 ( 
.A(n_2294),
.Y(n_2363)
);

INVx2_ASAP7_75t_SL g2364 ( 
.A(n_2007),
.Y(n_2364)
);

AND3x2_ASAP7_75t_L g2365 ( 
.A(n_2207),
.B(n_1775),
.C(n_1982),
.Y(n_2365)
);

INVx2_ASAP7_75t_L g2366 ( 
.A(n_2139),
.Y(n_2366)
);

INVx1_ASAP7_75t_L g2367 ( 
.A(n_2217),
.Y(n_2367)
);

INVx2_ASAP7_75t_L g2368 ( 
.A(n_2139),
.Y(n_2368)
);

INVx3_ASAP7_75t_L g2369 ( 
.A(n_2229),
.Y(n_2369)
);

BUFx3_ASAP7_75t_L g2370 ( 
.A(n_2134),
.Y(n_2370)
);

BUFx6f_ASAP7_75t_L g2371 ( 
.A(n_2055),
.Y(n_2371)
);

BUFx2_ASAP7_75t_L g2372 ( 
.A(n_2026),
.Y(n_2372)
);

INVx5_ASAP7_75t_L g2373 ( 
.A(n_2013),
.Y(n_2373)
);

INVx1_ASAP7_75t_L g2374 ( 
.A(n_2229),
.Y(n_2374)
);

INVx1_ASAP7_75t_L g2375 ( 
.A(n_2300),
.Y(n_2375)
);

BUFx3_ASAP7_75t_L g2376 ( 
.A(n_2134),
.Y(n_2376)
);

INVx1_ASAP7_75t_L g2377 ( 
.A(n_2300),
.Y(n_2377)
);

NOR2xp33_ASAP7_75t_L g2378 ( 
.A(n_2057),
.B(n_1943),
.Y(n_2378)
);

INVx1_ASAP7_75t_L g2379 ( 
.A(n_2156),
.Y(n_2379)
);

INVx4_ASAP7_75t_L g2380 ( 
.A(n_2299),
.Y(n_2380)
);

NAND2xp5_ASAP7_75t_SL g2381 ( 
.A(n_2116),
.B(n_1968),
.Y(n_2381)
);

HB1xp67_ASAP7_75t_L g2382 ( 
.A(n_2109),
.Y(n_2382)
);

INVx2_ASAP7_75t_L g2383 ( 
.A(n_2156),
.Y(n_2383)
);

INVx2_ASAP7_75t_SL g2384 ( 
.A(n_2036),
.Y(n_2384)
);

AND2x2_ASAP7_75t_SL g2385 ( 
.A(n_2205),
.B(n_1967),
.Y(n_2385)
);

INVx1_ASAP7_75t_L g2386 ( 
.A(n_2164),
.Y(n_2386)
);

INVx1_ASAP7_75t_L g2387 ( 
.A(n_2164),
.Y(n_2387)
);

INVx2_ASAP7_75t_L g2388 ( 
.A(n_2167),
.Y(n_2388)
);

OR2x2_ASAP7_75t_L g2389 ( 
.A(n_2005),
.B(n_1944),
.Y(n_2389)
);

NAND2xp5_ASAP7_75t_L g2390 ( 
.A(n_2113),
.B(n_1859),
.Y(n_2390)
);

INVx2_ASAP7_75t_L g2391 ( 
.A(n_2167),
.Y(n_2391)
);

NAND2xp5_ASAP7_75t_L g2392 ( 
.A(n_2200),
.B(n_1859),
.Y(n_2392)
);

INVx1_ASAP7_75t_L g2393 ( 
.A(n_2181),
.Y(n_2393)
);

NOR2xp33_ASAP7_75t_L g2394 ( 
.A(n_2038),
.B(n_1943),
.Y(n_2394)
);

INVx2_ASAP7_75t_L g2395 ( 
.A(n_2181),
.Y(n_2395)
);

AOI22xp33_ASAP7_75t_L g2396 ( 
.A1(n_2258),
.A2(n_2132),
.B1(n_1997),
.B2(n_2203),
.Y(n_2396)
);

NOR2x1p5_ASAP7_75t_L g2397 ( 
.A(n_2084),
.B(n_1985),
.Y(n_2397)
);

AOI22xp33_ASAP7_75t_L g2398 ( 
.A1(n_2262),
.A2(n_1937),
.B1(n_1877),
.B2(n_1890),
.Y(n_2398)
);

AND2x6_ASAP7_75t_L g2399 ( 
.A(n_2103),
.B(n_1967),
.Y(n_2399)
);

NAND2xp5_ASAP7_75t_SL g2400 ( 
.A(n_2174),
.B(n_1968),
.Y(n_2400)
);

AND2x2_ASAP7_75t_L g2401 ( 
.A(n_2309),
.B(n_1968),
.Y(n_2401)
);

CKINVDCx5p33_ASAP7_75t_R g2402 ( 
.A(n_2137),
.Y(n_2402)
);

NAND2xp33_ASAP7_75t_SL g2403 ( 
.A(n_2194),
.B(n_1968),
.Y(n_2403)
);

BUFx3_ASAP7_75t_L g2404 ( 
.A(n_2013),
.Y(n_2404)
);

BUFx3_ASAP7_75t_L g2405 ( 
.A(n_2123),
.Y(n_2405)
);

NAND2xp5_ASAP7_75t_L g2406 ( 
.A(n_2221),
.B(n_1871),
.Y(n_2406)
);

INVx2_ASAP7_75t_L g2407 ( 
.A(n_2197),
.Y(n_2407)
);

INVx2_ASAP7_75t_L g2408 ( 
.A(n_2197),
.Y(n_2408)
);

INVx1_ASAP7_75t_L g2409 ( 
.A(n_2208),
.Y(n_2409)
);

INVx1_ASAP7_75t_L g2410 ( 
.A(n_2208),
.Y(n_2410)
);

INVx1_ASAP7_75t_L g2411 ( 
.A(n_2273),
.Y(n_2411)
);

OR2x6_ASAP7_75t_L g2412 ( 
.A(n_2123),
.B(n_1983),
.Y(n_2412)
);

INVx2_ASAP7_75t_L g2413 ( 
.A(n_2273),
.Y(n_2413)
);

INVx4_ASAP7_75t_L g2414 ( 
.A(n_2299),
.Y(n_2414)
);

INVx1_ASAP7_75t_L g2415 ( 
.A(n_2274),
.Y(n_2415)
);

NAND2xp5_ASAP7_75t_SL g2416 ( 
.A(n_2027),
.B(n_1983),
.Y(n_2416)
);

INVx4_ASAP7_75t_L g2417 ( 
.A(n_2055),
.Y(n_2417)
);

INVx1_ASAP7_75t_L g2418 ( 
.A(n_2274),
.Y(n_2418)
);

INVx1_ASAP7_75t_L g2419 ( 
.A(n_2288),
.Y(n_2419)
);

INVx1_ASAP7_75t_L g2420 ( 
.A(n_2288),
.Y(n_2420)
);

INVx3_ASAP7_75t_L g2421 ( 
.A(n_2103),
.Y(n_2421)
);

BUFx10_ASAP7_75t_L g2422 ( 
.A(n_2094),
.Y(n_2422)
);

INVx2_ASAP7_75t_L g2423 ( 
.A(n_2307),
.Y(n_2423)
);

NOR2xp33_ASAP7_75t_L g2424 ( 
.A(n_2039),
.B(n_1983),
.Y(n_2424)
);

INVx2_ASAP7_75t_SL g2425 ( 
.A(n_2109),
.Y(n_2425)
);

INVx3_ASAP7_75t_L g2426 ( 
.A(n_2125),
.Y(n_2426)
);

INVx2_ASAP7_75t_L g2427 ( 
.A(n_2307),
.Y(n_2427)
);

OR2x6_ASAP7_75t_L g2428 ( 
.A(n_2124),
.B(n_1983),
.Y(n_2428)
);

AOI22xp5_ASAP7_75t_L g2429 ( 
.A1(n_2168),
.A2(n_1937),
.B1(n_1892),
.B2(n_1931),
.Y(n_2429)
);

INVx2_ASAP7_75t_L g2430 ( 
.A(n_2312),
.Y(n_2430)
);

INVx2_ASAP7_75t_L g2431 ( 
.A(n_2312),
.Y(n_2431)
);

INVx1_ASAP7_75t_L g2432 ( 
.A(n_2068),
.Y(n_2432)
);

NOR2xp33_ASAP7_75t_L g2433 ( 
.A(n_2004),
.B(n_1929),
.Y(n_2433)
);

BUFx3_ASAP7_75t_L g2434 ( 
.A(n_2124),
.Y(n_2434)
);

INVx2_ASAP7_75t_L g2435 ( 
.A(n_2125),
.Y(n_2435)
);

OR2x6_ASAP7_75t_L g2436 ( 
.A(n_2176),
.B(n_1928),
.Y(n_2436)
);

INVx2_ASAP7_75t_L g2437 ( 
.A(n_2050),
.Y(n_2437)
);

BUFx3_ASAP7_75t_L g2438 ( 
.A(n_2001),
.Y(n_2438)
);

INVx2_ASAP7_75t_L g2439 ( 
.A(n_2050),
.Y(n_2439)
);

AND2x6_ASAP7_75t_L g2440 ( 
.A(n_2063),
.B(n_1928),
.Y(n_2440)
);

AOI22xp33_ASAP7_75t_L g2441 ( 
.A1(n_2262),
.A2(n_2248),
.B1(n_2256),
.B2(n_2250),
.Y(n_2441)
);

INVx1_ASAP7_75t_L g2442 ( 
.A(n_2070),
.Y(n_2442)
);

INVx2_ASAP7_75t_L g2443 ( 
.A(n_2052),
.Y(n_2443)
);

BUFx10_ASAP7_75t_L g2444 ( 
.A(n_2194),
.Y(n_2444)
);

INVx1_ASAP7_75t_L g2445 ( 
.A(n_2073),
.Y(n_2445)
);

INVx1_ASAP7_75t_L g2446 ( 
.A(n_2076),
.Y(n_2446)
);

INVx1_ASAP7_75t_L g2447 ( 
.A(n_2101),
.Y(n_2447)
);

NOR2xp33_ASAP7_75t_L g2448 ( 
.A(n_2029),
.B(n_1930),
.Y(n_2448)
);

NAND2xp5_ASAP7_75t_L g2449 ( 
.A(n_2287),
.B(n_1892),
.Y(n_2449)
);

INVx2_ASAP7_75t_L g2450 ( 
.A(n_2052),
.Y(n_2450)
);

INVx1_ASAP7_75t_L g2451 ( 
.A(n_2111),
.Y(n_2451)
);

NAND2xp5_ASAP7_75t_L g2452 ( 
.A(n_2301),
.B(n_1892),
.Y(n_2452)
);

INVx2_ASAP7_75t_L g2453 ( 
.A(n_2063),
.Y(n_2453)
);

INVx2_ASAP7_75t_L g2454 ( 
.A(n_2088),
.Y(n_2454)
);

NAND2xp5_ASAP7_75t_L g2455 ( 
.A(n_2043),
.B(n_1892),
.Y(n_2455)
);

NAND2xp5_ASAP7_75t_L g2456 ( 
.A(n_2053),
.B(n_1889),
.Y(n_2456)
);

INVx4_ASAP7_75t_L g2457 ( 
.A(n_2055),
.Y(n_2457)
);

INVx1_ASAP7_75t_L g2458 ( 
.A(n_2149),
.Y(n_2458)
);

INVx2_ASAP7_75t_L g2459 ( 
.A(n_2088),
.Y(n_2459)
);

INVx2_ASAP7_75t_L g2460 ( 
.A(n_2159),
.Y(n_2460)
);

INVx2_ASAP7_75t_L g2461 ( 
.A(n_2177),
.Y(n_2461)
);

INVx2_ASAP7_75t_L g2462 ( 
.A(n_2180),
.Y(n_2462)
);

INVx1_ASAP7_75t_L g2463 ( 
.A(n_2189),
.Y(n_2463)
);

INVx2_ASAP7_75t_L g2464 ( 
.A(n_2204),
.Y(n_2464)
);

NAND3xp33_ASAP7_75t_L g2465 ( 
.A(n_2061),
.B(n_1945),
.C(n_1934),
.Y(n_2465)
);

INVx1_ASAP7_75t_L g2466 ( 
.A(n_2219),
.Y(n_2466)
);

INVx2_ASAP7_75t_L g2467 ( 
.A(n_2223),
.Y(n_2467)
);

INVx4_ASAP7_75t_L g2468 ( 
.A(n_2066),
.Y(n_2468)
);

INVx4_ASAP7_75t_L g2469 ( 
.A(n_2066),
.Y(n_2469)
);

INVx4_ASAP7_75t_L g2470 ( 
.A(n_2066),
.Y(n_2470)
);

INVx3_ASAP7_75t_L g2471 ( 
.A(n_2226),
.Y(n_2471)
);

NAND2xp5_ASAP7_75t_L g2472 ( 
.A(n_2296),
.B(n_1890),
.Y(n_2472)
);

INVx5_ASAP7_75t_L g2473 ( 
.A(n_2283),
.Y(n_2473)
);

INVx1_ASAP7_75t_L g2474 ( 
.A(n_2231),
.Y(n_2474)
);

INVx1_ASAP7_75t_L g2475 ( 
.A(n_2246),
.Y(n_2475)
);

AND2x6_ASAP7_75t_L g2476 ( 
.A(n_2269),
.B(n_1928),
.Y(n_2476)
);

BUFx6f_ASAP7_75t_L g2477 ( 
.A(n_2102),
.Y(n_2477)
);

NOR2xp33_ASAP7_75t_L g2478 ( 
.A(n_2220),
.B(n_1928),
.Y(n_2478)
);

INVx1_ASAP7_75t_L g2479 ( 
.A(n_2259),
.Y(n_2479)
);

INVx2_ASAP7_75t_L g2480 ( 
.A(n_2260),
.Y(n_2480)
);

BUFx3_ASAP7_75t_L g2481 ( 
.A(n_2102),
.Y(n_2481)
);

AND2x2_ASAP7_75t_L g2482 ( 
.A(n_2310),
.B(n_1946),
.Y(n_2482)
);

AOI22xp33_ASAP7_75t_L g2483 ( 
.A1(n_2277),
.A2(n_2282),
.B1(n_2292),
.B2(n_2284),
.Y(n_2483)
);

NOR2xp33_ASAP7_75t_L g2484 ( 
.A(n_2011),
.B(n_1946),
.Y(n_2484)
);

INVx2_ASAP7_75t_L g2485 ( 
.A(n_2267),
.Y(n_2485)
);

INVx3_ASAP7_75t_L g2486 ( 
.A(n_2308),
.Y(n_2486)
);

OR2x2_ASAP7_75t_L g2487 ( 
.A(n_2129),
.B(n_1985),
.Y(n_2487)
);

INVx5_ASAP7_75t_L g2488 ( 
.A(n_2283),
.Y(n_2488)
);

INVx2_ASAP7_75t_L g2489 ( 
.A(n_2235),
.Y(n_2489)
);

AND2x2_ASAP7_75t_L g2490 ( 
.A(n_2313),
.B(n_2184),
.Y(n_2490)
);

NOR2xp33_ASAP7_75t_L g2491 ( 
.A(n_2031),
.B(n_1946),
.Y(n_2491)
);

NAND2xp5_ASAP7_75t_SL g2492 ( 
.A(n_2059),
.B(n_1946),
.Y(n_2492)
);

INVx2_ASAP7_75t_SL g2493 ( 
.A(n_2074),
.Y(n_2493)
);

AND2x2_ASAP7_75t_L g2494 ( 
.A(n_2209),
.B(n_2232),
.Y(n_2494)
);

NAND2xp5_ASAP7_75t_SL g2495 ( 
.A(n_2133),
.B(n_1851),
.Y(n_2495)
);

AOI22xp33_ASAP7_75t_L g2496 ( 
.A1(n_2303),
.A2(n_1900),
.B1(n_1952),
.B2(n_1851),
.Y(n_2496)
);

INVx2_ASAP7_75t_L g2497 ( 
.A(n_2261),
.Y(n_2497)
);

BUFx6f_ASAP7_75t_L g2498 ( 
.A(n_2102),
.Y(n_2498)
);

INVx1_ASAP7_75t_L g2499 ( 
.A(n_2298),
.Y(n_2499)
);

NAND2xp5_ASAP7_75t_L g2500 ( 
.A(n_2304),
.B(n_1900),
.Y(n_2500)
);

INVx1_ASAP7_75t_L g2501 ( 
.A(n_2266),
.Y(n_2501)
);

AOI22xp33_ASAP7_75t_L g2502 ( 
.A1(n_2305),
.A2(n_1952),
.B1(n_1851),
.B2(n_1882),
.Y(n_2502)
);

NOR2xp33_ASAP7_75t_L g2503 ( 
.A(n_2042),
.B(n_1804),
.Y(n_2503)
);

AOI22xp33_ASAP7_75t_L g2504 ( 
.A1(n_2131),
.A2(n_1851),
.B1(n_1882),
.B2(n_1864),
.Y(n_2504)
);

NAND2xp5_ASAP7_75t_L g2505 ( 
.A(n_2080),
.B(n_1771),
.Y(n_2505)
);

INVx2_ASAP7_75t_L g2506 ( 
.A(n_2271),
.Y(n_2506)
);

OR2x2_ASAP7_75t_L g2507 ( 
.A(n_2157),
.B(n_1822),
.Y(n_2507)
);

INVxp67_ASAP7_75t_SL g2508 ( 
.A(n_2078),
.Y(n_2508)
);

INVx2_ASAP7_75t_L g2509 ( 
.A(n_2251),
.Y(n_2509)
);

INVx1_ASAP7_75t_L g2510 ( 
.A(n_2121),
.Y(n_2510)
);

INVx1_ASAP7_75t_L g2511 ( 
.A(n_2187),
.Y(n_2511)
);

INVx2_ASAP7_75t_L g2512 ( 
.A(n_2251),
.Y(n_2512)
);

INVx1_ASAP7_75t_L g2513 ( 
.A(n_2222),
.Y(n_2513)
);

NAND2xp5_ASAP7_75t_L g2514 ( 
.A(n_2270),
.B(n_2079),
.Y(n_2514)
);

AOI22xp33_ASAP7_75t_L g2515 ( 
.A1(n_2253),
.A2(n_1864),
.B1(n_1742),
.B2(n_1754),
.Y(n_2515)
);

BUFx10_ASAP7_75t_L g2516 ( 
.A(n_2240),
.Y(n_2516)
);

NAND2xp5_ASAP7_75t_SL g2517 ( 
.A(n_2014),
.B(n_1959),
.Y(n_2517)
);

INVx2_ASAP7_75t_SL g2518 ( 
.A(n_2314),
.Y(n_2518)
);

OR2x6_ASAP7_75t_L g2519 ( 
.A(n_2069),
.B(n_1957),
.Y(n_2519)
);

INVx5_ASAP7_75t_L g2520 ( 
.A(n_2283),
.Y(n_2520)
);

INVx1_ASAP7_75t_L g2521 ( 
.A(n_2202),
.Y(n_2521)
);

INVx1_ASAP7_75t_L g2522 ( 
.A(n_2168),
.Y(n_2522)
);

INVx1_ASAP7_75t_L g2523 ( 
.A(n_2095),
.Y(n_2523)
);

BUFx4f_ASAP7_75t_L g2524 ( 
.A(n_2283),
.Y(n_2524)
);

INVxp67_ASAP7_75t_SL g2525 ( 
.A(n_2085),
.Y(n_2525)
);

NOR2xp33_ASAP7_75t_L g2526 ( 
.A(n_2060),
.B(n_1896),
.Y(n_2526)
);

INVx1_ASAP7_75t_L g2527 ( 
.A(n_2257),
.Y(n_2527)
);

INVx3_ASAP7_75t_L g2528 ( 
.A(n_2032),
.Y(n_2528)
);

INVx2_ASAP7_75t_L g2529 ( 
.A(n_2257),
.Y(n_2529)
);

NOR2xp33_ASAP7_75t_L g2530 ( 
.A(n_2065),
.B(n_1896),
.Y(n_2530)
);

INVx4_ASAP7_75t_L g2531 ( 
.A(n_2240),
.Y(n_2531)
);

INVx2_ASAP7_75t_L g2532 ( 
.A(n_2265),
.Y(n_2532)
);

INVx1_ASAP7_75t_L g2533 ( 
.A(n_2265),
.Y(n_2533)
);

INVx2_ASAP7_75t_L g2534 ( 
.A(n_2280),
.Y(n_2534)
);

INVx2_ASAP7_75t_L g2535 ( 
.A(n_2280),
.Y(n_2535)
);

INVx1_ASAP7_75t_L g2536 ( 
.A(n_2289),
.Y(n_2536)
);

OA22x2_ASAP7_75t_L g2537 ( 
.A1(n_2227),
.A2(n_1854),
.B1(n_1856),
.B2(n_1852),
.Y(n_2537)
);

NOR2xp33_ASAP7_75t_L g2538 ( 
.A(n_2237),
.B(n_1896),
.Y(n_2538)
);

AND2x4_ASAP7_75t_L g2539 ( 
.A(n_2140),
.B(n_1751),
.Y(n_2539)
);

INVx2_ASAP7_75t_L g2540 ( 
.A(n_2289),
.Y(n_2540)
);

INVx1_ASAP7_75t_L g2541 ( 
.A(n_2272),
.Y(n_2541)
);

AOI22xp33_ASAP7_75t_L g2542 ( 
.A1(n_2225),
.A2(n_1864),
.B1(n_1742),
.B2(n_1754),
.Y(n_2542)
);

BUFx3_ASAP7_75t_L g2543 ( 
.A(n_2216),
.Y(n_2543)
);

INVx2_ASAP7_75t_L g2544 ( 
.A(n_2089),
.Y(n_2544)
);

INVx1_ASAP7_75t_L g2545 ( 
.A(n_2145),
.Y(n_2545)
);

INVxp33_ASAP7_75t_L g2546 ( 
.A(n_2020),
.Y(n_2546)
);

INVx1_ASAP7_75t_L g2547 ( 
.A(n_2145),
.Y(n_2547)
);

NAND2xp5_ASAP7_75t_SL g2548 ( 
.A(n_2022),
.B(n_1740),
.Y(n_2548)
);

BUFx3_ASAP7_75t_L g2549 ( 
.A(n_2249),
.Y(n_2549)
);

INVx2_ASAP7_75t_L g2550 ( 
.A(n_2091),
.Y(n_2550)
);

NAND2xp5_ASAP7_75t_L g2551 ( 
.A(n_2148),
.B(n_2150),
.Y(n_2551)
);

INVx4_ASAP7_75t_L g2552 ( 
.A(n_2225),
.Y(n_2552)
);

NAND2xp33_ASAP7_75t_L g2553 ( 
.A(n_2108),
.B(n_1740),
.Y(n_2553)
);

INVx2_ASAP7_75t_L g2554 ( 
.A(n_2141),
.Y(n_2554)
);

INVx1_ASAP7_75t_L g2555 ( 
.A(n_2279),
.Y(n_2555)
);

INVx2_ASAP7_75t_L g2556 ( 
.A(n_2141),
.Y(n_2556)
);

INVx2_ASAP7_75t_L g2557 ( 
.A(n_2236),
.Y(n_2557)
);

NAND2xp5_ASAP7_75t_L g2558 ( 
.A(n_2151),
.B(n_1827),
.Y(n_2558)
);

INVx1_ASAP7_75t_L g2559 ( 
.A(n_2152),
.Y(n_2559)
);

INVx1_ASAP7_75t_L g2560 ( 
.A(n_2153),
.Y(n_2560)
);

INVx1_ASAP7_75t_L g2561 ( 
.A(n_2158),
.Y(n_2561)
);

OAI21xp33_ASAP7_75t_SL g2562 ( 
.A1(n_2096),
.A2(n_1721),
.B(n_1848),
.Y(n_2562)
);

BUFx3_ASAP7_75t_L g2563 ( 
.A(n_2228),
.Y(n_2563)
);

INVx3_ASAP7_75t_L g2564 ( 
.A(n_2302),
.Y(n_2564)
);

INVx2_ASAP7_75t_L g2565 ( 
.A(n_2236),
.Y(n_2565)
);

AND2x6_ASAP7_75t_L g2566 ( 
.A(n_2178),
.B(n_1740),
.Y(n_2566)
);

INVx3_ASAP7_75t_L g2567 ( 
.A(n_2214),
.Y(n_2567)
);

OR2x2_ASAP7_75t_L g2568 ( 
.A(n_2037),
.B(n_1751),
.Y(n_2568)
);

INVx2_ASAP7_75t_L g2569 ( 
.A(n_2241),
.Y(n_2569)
);

AND2x6_ASAP7_75t_L g2570 ( 
.A(n_2190),
.B(n_1740),
.Y(n_2570)
);

INVx3_ASAP7_75t_L g2571 ( 
.A(n_2241),
.Y(n_2571)
);

AND2x2_ASAP7_75t_L g2572 ( 
.A(n_2010),
.B(n_1852),
.Y(n_2572)
);

AO21x2_ASAP7_75t_L g2573 ( 
.A1(n_2114),
.A2(n_1721),
.B(n_1848),
.Y(n_2573)
);

NOR2xp33_ASAP7_75t_L g2574 ( 
.A(n_2104),
.B(n_1806),
.Y(n_2574)
);

INVx2_ASAP7_75t_L g2575 ( 
.A(n_2182),
.Y(n_2575)
);

INVx2_ASAP7_75t_L g2576 ( 
.A(n_2182),
.Y(n_2576)
);

INVxp67_ASAP7_75t_SL g2577 ( 
.A(n_2046),
.Y(n_2577)
);

INVx3_ASAP7_75t_L g2578 ( 
.A(n_2306),
.Y(n_2578)
);

AO22x2_ASAP7_75t_L g2579 ( 
.A1(n_2293),
.A2(n_1827),
.B1(n_1854),
.B2(n_1852),
.Y(n_2579)
);

NAND2xp5_ASAP7_75t_L g2580 ( 
.A(n_2162),
.B(n_1827),
.Y(n_2580)
);

NAND2xp5_ASAP7_75t_SL g2581 ( 
.A(n_2056),
.B(n_1744),
.Y(n_2581)
);

AND2x2_ASAP7_75t_SL g2582 ( 
.A(n_1999),
.B(n_1706),
.Y(n_2582)
);

NOR2xp33_ASAP7_75t_L g2583 ( 
.A(n_2006),
.B(n_1806),
.Y(n_2583)
);

AOI22xp33_ASAP7_75t_L g2584 ( 
.A1(n_2090),
.A2(n_1742),
.B1(n_1754),
.B2(n_1706),
.Y(n_2584)
);

AND2x4_ASAP7_75t_L g2585 ( 
.A(n_2047),
.B(n_1854),
.Y(n_2585)
);

INVx2_ASAP7_75t_L g2586 ( 
.A(n_2185),
.Y(n_2586)
);

INVx1_ASAP7_75t_L g2587 ( 
.A(n_2238),
.Y(n_2587)
);

BUFx10_ASAP7_75t_L g2588 ( 
.A(n_2119),
.Y(n_2588)
);

INVx5_ASAP7_75t_L g2589 ( 
.A(n_2161),
.Y(n_2589)
);

INVx1_ASAP7_75t_L g2590 ( 
.A(n_2193),
.Y(n_2590)
);

INVx1_ASAP7_75t_L g2591 ( 
.A(n_2196),
.Y(n_2591)
);

INVx4_ASAP7_75t_L g2592 ( 
.A(n_2185),
.Y(n_2592)
);

OR2x2_ASAP7_75t_L g2593 ( 
.A(n_2128),
.B(n_1856),
.Y(n_2593)
);

INVx1_ASAP7_75t_L g2594 ( 
.A(n_2239),
.Y(n_2594)
);

NAND2xp5_ASAP7_75t_SL g2595 ( 
.A(n_2044),
.B(n_1744),
.Y(n_2595)
);

NOR2xp33_ASAP7_75t_L g2596 ( 
.A(n_2009),
.B(n_1806),
.Y(n_2596)
);

NAND2xp5_ASAP7_75t_SL g2597 ( 
.A(n_2008),
.B(n_1744),
.Y(n_2597)
);

INVx2_ASAP7_75t_L g2598 ( 
.A(n_2191),
.Y(n_2598)
);

INVx1_ASAP7_75t_L g2599 ( 
.A(n_2242),
.Y(n_2599)
);

INVx1_ASAP7_75t_L g2600 ( 
.A(n_2247),
.Y(n_2600)
);

INVx1_ASAP7_75t_L g2601 ( 
.A(n_2255),
.Y(n_2601)
);

INVx1_ASAP7_75t_L g2602 ( 
.A(n_2206),
.Y(n_2602)
);

NAND3xp33_ASAP7_75t_L g2603 ( 
.A(n_2120),
.B(n_1760),
.C(n_1726),
.Y(n_2603)
);

INVx2_ASAP7_75t_SL g2604 ( 
.A(n_2161),
.Y(n_2604)
);

NOR2xp33_ASAP7_75t_L g2605 ( 
.A(n_2072),
.B(n_1776),
.Y(n_2605)
);

AND2x2_ASAP7_75t_L g2606 ( 
.A(n_2136),
.B(n_1856),
.Y(n_2606)
);

OR2x6_ASAP7_75t_L g2607 ( 
.A(n_2064),
.B(n_1776),
.Y(n_2607)
);

INVx2_ASAP7_75t_L g2608 ( 
.A(n_2191),
.Y(n_2608)
);

HB1xp67_ASAP7_75t_L g2609 ( 
.A(n_2169),
.Y(n_2609)
);

INVx2_ASAP7_75t_L g2610 ( 
.A(n_2199),
.Y(n_2610)
);

INVx4_ASAP7_75t_L g2611 ( 
.A(n_2199),
.Y(n_2611)
);

AO22x2_ASAP7_75t_L g2612 ( 
.A1(n_2254),
.A2(n_1875),
.B1(n_1872),
.B2(n_60),
.Y(n_2612)
);

BUFx4f_ASAP7_75t_L g2613 ( 
.A(n_2117),
.Y(n_2613)
);

AND2x6_ASAP7_75t_L g2614 ( 
.A(n_2264),
.B(n_1744),
.Y(n_2614)
);

OAI22xp33_ASAP7_75t_L g2615 ( 
.A1(n_2142),
.A2(n_1765),
.B1(n_1805),
.B2(n_1706),
.Y(n_2615)
);

NAND2xp5_ASAP7_75t_L g2616 ( 
.A(n_2097),
.B(n_1765),
.Y(n_2616)
);

INVx2_ASAP7_75t_L g2617 ( 
.A(n_2201),
.Y(n_2617)
);

INVx3_ASAP7_75t_L g2618 ( 
.A(n_2201),
.Y(n_2618)
);

INVxp67_ASAP7_75t_SL g2619 ( 
.A(n_2048),
.Y(n_2619)
);

INVx1_ASAP7_75t_L g2620 ( 
.A(n_2211),
.Y(n_2620)
);

AND2x2_ASAP7_75t_L g2621 ( 
.A(n_2017),
.B(n_1872),
.Y(n_2621)
);

AND2x2_ASAP7_75t_L g2622 ( 
.A(n_2017),
.B(n_2041),
.Y(n_2622)
);

NAND2xp5_ASAP7_75t_L g2623 ( 
.A(n_2106),
.B(n_1765),
.Y(n_2623)
);

INVx4_ASAP7_75t_L g2624 ( 
.A(n_2211),
.Y(n_2624)
);

INVx1_ASAP7_75t_L g2625 ( 
.A(n_2233),
.Y(n_2625)
);

NAND2xp5_ASAP7_75t_L g2626 ( 
.A(n_2115),
.B(n_1805),
.Y(n_2626)
);

NOR2xp33_ASAP7_75t_L g2627 ( 
.A(n_2071),
.B(n_1760),
.Y(n_2627)
);

NOR2xp33_ASAP7_75t_L g2628 ( 
.A(n_2087),
.B(n_1760),
.Y(n_2628)
);

XOR2xp5_ASAP7_75t_L g2629 ( 
.A(n_2081),
.B(n_1933),
.Y(n_2629)
);

OR2x2_ASAP7_75t_L g2630 ( 
.A(n_2169),
.B(n_1872),
.Y(n_2630)
);

NAND2xp5_ASAP7_75t_L g2631 ( 
.A(n_2138),
.B(n_1805),
.Y(n_2631)
);

INVx1_ASAP7_75t_L g2632 ( 
.A(n_2093),
.Y(n_2632)
);

INVx1_ASAP7_75t_L g2633 ( 
.A(n_2179),
.Y(n_2633)
);

BUFx2_ASAP7_75t_L g2634 ( 
.A(n_2051),
.Y(n_2634)
);

BUFx4f_ASAP7_75t_L g2635 ( 
.A(n_2118),
.Y(n_2635)
);

INVx4_ASAP7_75t_L g2636 ( 
.A(n_2228),
.Y(n_2636)
);

INVx3_ASAP7_75t_L g2637 ( 
.A(n_2030),
.Y(n_2637)
);

INVx3_ASAP7_75t_L g2638 ( 
.A(n_2041),
.Y(n_2638)
);

BUFx10_ASAP7_75t_L g2639 ( 
.A(n_2188),
.Y(n_2639)
);

INVx2_ASAP7_75t_L g2640 ( 
.A(n_2210),
.Y(n_2640)
);

NOR2xp33_ASAP7_75t_L g2641 ( 
.A(n_2130),
.B(n_2146),
.Y(n_2641)
);

INVx3_ASAP7_75t_L g2642 ( 
.A(n_2023),
.Y(n_2642)
);

NAND2xp5_ASAP7_75t_SL g2643 ( 
.A(n_2012),
.B(n_1757),
.Y(n_2643)
);

INVx2_ASAP7_75t_SL g2644 ( 
.A(n_2252),
.Y(n_2644)
);

NOR2xp33_ASAP7_75t_L g2645 ( 
.A(n_1996),
.B(n_1726),
.Y(n_2645)
);

INVx3_ASAP7_75t_L g2646 ( 
.A(n_2023),
.Y(n_2646)
);

INVx1_ASAP7_75t_L g2647 ( 
.A(n_2224),
.Y(n_2647)
);

INVx1_ASAP7_75t_L g2648 ( 
.A(n_2244),
.Y(n_2648)
);

OAI22xp5_ASAP7_75t_L g2649 ( 
.A1(n_2144),
.A2(n_1835),
.B1(n_1807),
.B2(n_1728),
.Y(n_2649)
);

INVx2_ASAP7_75t_L g2650 ( 
.A(n_2213),
.Y(n_2650)
);

NAND2xp5_ASAP7_75t_SL g2651 ( 
.A(n_2083),
.B(n_1757),
.Y(n_2651)
);

BUFx4f_ASAP7_75t_L g2652 ( 
.A(n_2183),
.Y(n_2652)
);

NAND2xp5_ASAP7_75t_SL g2653 ( 
.A(n_2099),
.B(n_1757),
.Y(n_2653)
);

INVx5_ASAP7_75t_L g2654 ( 
.A(n_2186),
.Y(n_2654)
);

NAND2xp5_ASAP7_75t_SL g2655 ( 
.A(n_2143),
.B(n_2100),
.Y(n_2655)
);

INVx2_ASAP7_75t_SL g2656 ( 
.A(n_2170),
.Y(n_2656)
);

AND2x2_ASAP7_75t_L g2657 ( 
.A(n_2154),
.B(n_1875),
.Y(n_2657)
);

INVx2_ASAP7_75t_L g2658 ( 
.A(n_2230),
.Y(n_2658)
);

INVx2_ASAP7_75t_SL g2659 ( 
.A(n_2275),
.Y(n_2659)
);

AOI22xp33_ASAP7_75t_L g2660 ( 
.A1(n_2092),
.A2(n_1835),
.B1(n_1807),
.B2(n_1875),
.Y(n_2660)
);

INVx1_ASAP7_75t_L g2661 ( 
.A(n_2276),
.Y(n_2661)
);

NOR2xp33_ASAP7_75t_L g2662 ( 
.A(n_2002),
.B(n_1726),
.Y(n_2662)
);

INVx2_ASAP7_75t_L g2663 ( 
.A(n_2285),
.Y(n_2663)
);

INVx2_ASAP7_75t_L g2664 ( 
.A(n_2286),
.Y(n_2664)
);

INVx1_ASAP7_75t_L g2665 ( 
.A(n_2291),
.Y(n_2665)
);

INVx4_ASAP7_75t_L g2666 ( 
.A(n_2278),
.Y(n_2666)
);

NAND2xp5_ASAP7_75t_L g2667 ( 
.A(n_2163),
.B(n_1807),
.Y(n_2667)
);

NAND2xp5_ASAP7_75t_L g2668 ( 
.A(n_2165),
.B(n_1835),
.Y(n_2668)
);

NAND2xp5_ASAP7_75t_SL g2669 ( 
.A(n_2024),
.B(n_1757),
.Y(n_2669)
);

NAND2xp5_ASAP7_75t_SL g2670 ( 
.A(n_2424),
.B(n_2075),
.Y(n_2670)
);

AND2x6_ASAP7_75t_L g2671 ( 
.A(n_2571),
.B(n_2297),
.Y(n_2671)
);

HB1xp67_ASAP7_75t_L g2672 ( 
.A(n_2372),
.Y(n_2672)
);

INVx4_ASAP7_75t_L g2673 ( 
.A(n_2321),
.Y(n_2673)
);

INVx2_ASAP7_75t_L g2674 ( 
.A(n_2366),
.Y(n_2674)
);

INVx2_ASAP7_75t_L g2675 ( 
.A(n_2366),
.Y(n_2675)
);

NOR2xp33_ASAP7_75t_L g2676 ( 
.A(n_2546),
.B(n_2045),
.Y(n_2676)
);

BUFx10_ASAP7_75t_L g2677 ( 
.A(n_2538),
.Y(n_2677)
);

NOR2x1p5_ASAP7_75t_L g2678 ( 
.A(n_2619),
.B(n_2045),
.Y(n_2678)
);

INVx1_ASAP7_75t_L g2679 ( 
.A(n_2368),
.Y(n_2679)
);

INVx3_ASAP7_75t_L g2680 ( 
.A(n_2340),
.Y(n_2680)
);

INVx1_ASAP7_75t_L g2681 ( 
.A(n_2368),
.Y(n_2681)
);

INVx1_ASAP7_75t_L g2682 ( 
.A(n_2383),
.Y(n_2682)
);

BUFx6f_ASAP7_75t_L g2683 ( 
.A(n_2371),
.Y(n_2683)
);

NAND2xp5_ASAP7_75t_L g2684 ( 
.A(n_2501),
.B(n_2268),
.Y(n_2684)
);

NAND2x1p5_ASAP7_75t_L g2685 ( 
.A(n_2473),
.B(n_1725),
.Y(n_2685)
);

INVx1_ASAP7_75t_L g2686 ( 
.A(n_2383),
.Y(n_2686)
);

INVx2_ASAP7_75t_L g2687 ( 
.A(n_2388),
.Y(n_2687)
);

INVx1_ASAP7_75t_L g2688 ( 
.A(n_2388),
.Y(n_2688)
);

AOI22xp33_ASAP7_75t_L g2689 ( 
.A1(n_2612),
.A2(n_2254),
.B1(n_2281),
.B2(n_2234),
.Y(n_2689)
);

NAND2xp5_ASAP7_75t_L g2690 ( 
.A(n_2333),
.B(n_2173),
.Y(n_2690)
);

NOR2xp33_ASAP7_75t_L g2691 ( 
.A(n_2361),
.B(n_2086),
.Y(n_2691)
);

AND2x4_ASAP7_75t_L g2692 ( 
.A(n_2384),
.B(n_2311),
.Y(n_2692)
);

INVxp67_ASAP7_75t_L g2693 ( 
.A(n_2401),
.Y(n_2693)
);

BUFx10_ASAP7_75t_L g2694 ( 
.A(n_2530),
.Y(n_2694)
);

NAND2xp5_ASAP7_75t_SL g2695 ( 
.A(n_2385),
.B(n_2122),
.Y(n_2695)
);

BUFx6f_ASAP7_75t_L g2696 ( 
.A(n_2371),
.Y(n_2696)
);

AND2x4_ASAP7_75t_L g2697 ( 
.A(n_2384),
.B(n_2481),
.Y(n_2697)
);

INVx1_ASAP7_75t_L g2698 ( 
.A(n_2391),
.Y(n_2698)
);

NOR2xp33_ASAP7_75t_L g2699 ( 
.A(n_2378),
.B(n_2033),
.Y(n_2699)
);

NAND2xp5_ASAP7_75t_L g2700 ( 
.A(n_2333),
.B(n_2295),
.Y(n_2700)
);

AND2x2_ASAP7_75t_L g2701 ( 
.A(n_2577),
.B(n_2160),
.Y(n_2701)
);

INVx1_ASAP7_75t_L g2702 ( 
.A(n_2391),
.Y(n_2702)
);

NAND2xp33_ASAP7_75t_L g2703 ( 
.A(n_2315),
.B(n_1767),
.Y(n_2703)
);

AOI22xp5_ASAP7_75t_L g2704 ( 
.A1(n_2396),
.A2(n_2281),
.B1(n_2195),
.B2(n_2172),
.Y(n_2704)
);

BUFx2_ASAP7_75t_L g2705 ( 
.A(n_2549),
.Y(n_2705)
);

INVx2_ASAP7_75t_L g2706 ( 
.A(n_2395),
.Y(n_2706)
);

INVx1_ASAP7_75t_L g2707 ( 
.A(n_2395),
.Y(n_2707)
);

AO22x2_ASAP7_75t_L g2708 ( 
.A1(n_2552),
.A2(n_2175),
.B1(n_2218),
.B2(n_2215),
.Y(n_2708)
);

OR2x2_ASAP7_75t_L g2709 ( 
.A(n_2389),
.B(n_1817),
.Y(n_2709)
);

NAND2x1_ASAP7_75t_L g2710 ( 
.A(n_2340),
.B(n_1728),
.Y(n_2710)
);

INVx1_ASAP7_75t_L g2711 ( 
.A(n_2407),
.Y(n_2711)
);

INVx2_ASAP7_75t_L g2712 ( 
.A(n_2407),
.Y(n_2712)
);

INVx8_ASAP7_75t_L g2713 ( 
.A(n_2326),
.Y(n_2713)
);

BUFx6f_ASAP7_75t_L g2714 ( 
.A(n_2371),
.Y(n_2714)
);

NAND2xp5_ASAP7_75t_SL g2715 ( 
.A(n_2385),
.B(n_2105),
.Y(n_2715)
);

BUFx10_ASAP7_75t_L g2716 ( 
.A(n_2662),
.Y(n_2716)
);

INVx2_ASAP7_75t_L g2717 ( 
.A(n_2408),
.Y(n_2717)
);

BUFx3_ASAP7_75t_L g2718 ( 
.A(n_2543),
.Y(n_2718)
);

INVx1_ASAP7_75t_L g2719 ( 
.A(n_2408),
.Y(n_2719)
);

BUFx3_ASAP7_75t_L g2720 ( 
.A(n_2543),
.Y(n_2720)
);

AND2x4_ASAP7_75t_L g2721 ( 
.A(n_2481),
.B(n_1767),
.Y(n_2721)
);

AND2x6_ASAP7_75t_L g2722 ( 
.A(n_2571),
.B(n_1767),
.Y(n_2722)
);

OR2x2_ASAP7_75t_L g2723 ( 
.A(n_2389),
.B(n_1817),
.Y(n_2723)
);

NAND2x1p5_ASAP7_75t_L g2724 ( 
.A(n_2473),
.B(n_1725),
.Y(n_2724)
);

INVx1_ASAP7_75t_L g2725 ( 
.A(n_2413),
.Y(n_2725)
);

INVx1_ASAP7_75t_L g2726 ( 
.A(n_2413),
.Y(n_2726)
);

INVx1_ASAP7_75t_L g2727 ( 
.A(n_2423),
.Y(n_2727)
);

INVxp67_ASAP7_75t_L g2728 ( 
.A(n_2401),
.Y(n_2728)
);

AND2x4_ASAP7_75t_L g2729 ( 
.A(n_2493),
.B(n_1767),
.Y(n_2729)
);

CKINVDCx20_ASAP7_75t_R g2730 ( 
.A(n_2336),
.Y(n_2730)
);

INVx1_ASAP7_75t_L g2731 ( 
.A(n_2423),
.Y(n_2731)
);

INVx2_ASAP7_75t_L g2732 ( 
.A(n_2427),
.Y(n_2732)
);

INVx1_ASAP7_75t_L g2733 ( 
.A(n_2427),
.Y(n_2733)
);

INVxp67_ASAP7_75t_L g2734 ( 
.A(n_2551),
.Y(n_2734)
);

INVx1_ASAP7_75t_L g2735 ( 
.A(n_2430),
.Y(n_2735)
);

INVx1_ASAP7_75t_L g2736 ( 
.A(n_2430),
.Y(n_2736)
);

INVx1_ASAP7_75t_L g2737 ( 
.A(n_2431),
.Y(n_2737)
);

AND2x2_ASAP7_75t_L g2738 ( 
.A(n_2494),
.B(n_2110),
.Y(n_2738)
);

NAND2xp5_ASAP7_75t_SL g2739 ( 
.A(n_2394),
.B(n_2135),
.Y(n_2739)
);

INVx1_ASAP7_75t_L g2740 ( 
.A(n_2431),
.Y(n_2740)
);

INVx2_ASAP7_75t_L g2741 ( 
.A(n_2379),
.Y(n_2741)
);

AOI22xp5_ASAP7_75t_L g2742 ( 
.A1(n_2490),
.A2(n_2171),
.B1(n_2147),
.B2(n_2245),
.Y(n_2742)
);

BUFx6f_ASAP7_75t_L g2743 ( 
.A(n_2371),
.Y(n_2743)
);

INVx1_ASAP7_75t_L g2744 ( 
.A(n_2386),
.Y(n_2744)
);

OR2x2_ASAP7_75t_SL g2745 ( 
.A(n_2603),
.B(n_1933),
.Y(n_2745)
);

AND2x2_ASAP7_75t_L g2746 ( 
.A(n_2494),
.B(n_2362),
.Y(n_2746)
);

OAI22xp5_ASAP7_75t_L g2747 ( 
.A1(n_2552),
.A2(n_1728),
.B1(n_1792),
.B2(n_1737),
.Y(n_2747)
);

INVx1_ASAP7_75t_L g2748 ( 
.A(n_2387),
.Y(n_2748)
);

AND2x4_ASAP7_75t_L g2749 ( 
.A(n_2493),
.B(n_1777),
.Y(n_2749)
);

INVx3_ASAP7_75t_L g2750 ( 
.A(n_2340),
.Y(n_2750)
);

CKINVDCx20_ASAP7_75t_R g2751 ( 
.A(n_2336),
.Y(n_2751)
);

INVx1_ASAP7_75t_L g2752 ( 
.A(n_2393),
.Y(n_2752)
);

INVx1_ASAP7_75t_L g2753 ( 
.A(n_2409),
.Y(n_2753)
);

INVx1_ASAP7_75t_L g2754 ( 
.A(n_2410),
.Y(n_2754)
);

AND2x4_ASAP7_75t_L g2755 ( 
.A(n_2482),
.B(n_1777),
.Y(n_2755)
);

BUFx6f_ASAP7_75t_L g2756 ( 
.A(n_2477),
.Y(n_2756)
);

BUFx6f_ASAP7_75t_L g2757 ( 
.A(n_2477),
.Y(n_2757)
);

AO22x2_ASAP7_75t_L g2758 ( 
.A1(n_2552),
.A2(n_60),
.B1(n_58),
.B2(n_59),
.Y(n_2758)
);

AND2x4_ASAP7_75t_L g2759 ( 
.A(n_2482),
.B(n_1777),
.Y(n_2759)
);

NOR2xp33_ASAP7_75t_L g2760 ( 
.A(n_2546),
.B(n_1933),
.Y(n_2760)
);

INVx1_ASAP7_75t_L g2761 ( 
.A(n_2411),
.Y(n_2761)
);

INVx1_ASAP7_75t_L g2762 ( 
.A(n_2415),
.Y(n_2762)
);

HB1xp67_ASAP7_75t_L g2763 ( 
.A(n_2343),
.Y(n_2763)
);

NOR2xp33_ASAP7_75t_L g2764 ( 
.A(n_2362),
.B(n_1777),
.Y(n_2764)
);

INVx1_ASAP7_75t_L g2765 ( 
.A(n_2418),
.Y(n_2765)
);

AND2x4_ASAP7_75t_L g2766 ( 
.A(n_2438),
.B(n_1780),
.Y(n_2766)
);

OAI221xp5_ASAP7_75t_L g2767 ( 
.A1(n_2659),
.A2(n_1737),
.B1(n_1802),
.B2(n_1797),
.C(n_1792),
.Y(n_2767)
);

HB1xp67_ASAP7_75t_L g2768 ( 
.A(n_2343),
.Y(n_2768)
);

NAND2xp5_ASAP7_75t_L g2769 ( 
.A(n_2349),
.B(n_1737),
.Y(n_2769)
);

INVx2_ASAP7_75t_L g2770 ( 
.A(n_2419),
.Y(n_2770)
);

BUFx6f_ASAP7_75t_L g2771 ( 
.A(n_2477),
.Y(n_2771)
);

INVx1_ASAP7_75t_L g2772 ( 
.A(n_2420),
.Y(n_2772)
);

INVx1_ASAP7_75t_SL g2773 ( 
.A(n_2507),
.Y(n_2773)
);

AO22x2_ASAP7_75t_L g2774 ( 
.A1(n_2557),
.A2(n_60),
.B1(n_58),
.B2(n_59),
.Y(n_2774)
);

BUFx2_ASAP7_75t_L g2775 ( 
.A(n_2549),
.Y(n_2775)
);

AND2x4_ASAP7_75t_L g2776 ( 
.A(n_2438),
.B(n_1780),
.Y(n_2776)
);

INVx1_ASAP7_75t_L g2777 ( 
.A(n_2327),
.Y(n_2777)
);

OAI22xp5_ASAP7_75t_L g2778 ( 
.A1(n_2545),
.A2(n_1792),
.B1(n_1802),
.B2(n_1797),
.Y(n_2778)
);

AND2x4_ASAP7_75t_L g2779 ( 
.A(n_2539),
.B(n_1780),
.Y(n_2779)
);

INVx1_ASAP7_75t_L g2780 ( 
.A(n_2341),
.Y(n_2780)
);

NAND2xp5_ASAP7_75t_L g2781 ( 
.A(n_2489),
.B(n_2497),
.Y(n_2781)
);

INVxp33_ASAP7_75t_L g2782 ( 
.A(n_2478),
.Y(n_2782)
);

NAND3xp33_ASAP7_75t_SL g2783 ( 
.A(n_2354),
.B(n_1725),
.C(n_58),
.Y(n_2783)
);

INVx1_ASAP7_75t_L g2784 ( 
.A(n_2348),
.Y(n_2784)
);

NAND3xp33_ASAP7_75t_L g2785 ( 
.A(n_2448),
.B(n_1786),
.C(n_1780),
.Y(n_2785)
);

INVx1_ASAP7_75t_SL g2786 ( 
.A(n_2507),
.Y(n_2786)
);

BUFx3_ASAP7_75t_L g2787 ( 
.A(n_2335),
.Y(n_2787)
);

AND2x4_ASAP7_75t_L g2788 ( 
.A(n_2539),
.B(n_1786),
.Y(n_2788)
);

NAND2xp5_ASAP7_75t_L g2789 ( 
.A(n_2489),
.B(n_1797),
.Y(n_2789)
);

NAND2xp5_ASAP7_75t_SL g2790 ( 
.A(n_2514),
.B(n_1786),
.Y(n_2790)
);

BUFx6f_ASAP7_75t_L g2791 ( 
.A(n_2477),
.Y(n_2791)
);

OAI22xp33_ASAP7_75t_L g2792 ( 
.A1(n_2537),
.A2(n_2659),
.B1(n_2591),
.B2(n_2590),
.Y(n_2792)
);

AND2x2_ASAP7_75t_L g2793 ( 
.A(n_2490),
.B(n_1802),
.Y(n_2793)
);

BUFx6f_ASAP7_75t_L g2794 ( 
.A(n_2498),
.Y(n_2794)
);

INVx1_ASAP7_75t_L g2795 ( 
.A(n_2356),
.Y(n_2795)
);

AND2x4_ASAP7_75t_L g2796 ( 
.A(n_2539),
.B(n_1786),
.Y(n_2796)
);

INVx1_ASAP7_75t_L g2797 ( 
.A(n_2363),
.Y(n_2797)
);

INVx1_ASAP7_75t_L g2798 ( 
.A(n_2317),
.Y(n_2798)
);

BUFx6f_ASAP7_75t_L g2799 ( 
.A(n_2498),
.Y(n_2799)
);

AND2x6_ASAP7_75t_L g2800 ( 
.A(n_2571),
.B(n_1791),
.Y(n_2800)
);

NOR2xp33_ASAP7_75t_L g2801 ( 
.A(n_2330),
.B(n_2433),
.Y(n_2801)
);

INVx1_ASAP7_75t_L g2802 ( 
.A(n_2317),
.Y(n_2802)
);

AND2x2_ASAP7_75t_L g2803 ( 
.A(n_2572),
.B(n_1817),
.Y(n_2803)
);

INVx1_ASAP7_75t_L g2804 ( 
.A(n_2319),
.Y(n_2804)
);

INVx3_ASAP7_75t_L g2805 ( 
.A(n_2357),
.Y(n_2805)
);

INVx1_ASAP7_75t_L g2806 ( 
.A(n_2319),
.Y(n_2806)
);

BUFx6f_ASAP7_75t_L g2807 ( 
.A(n_2498),
.Y(n_2807)
);

INVx2_ASAP7_75t_L g2808 ( 
.A(n_2460),
.Y(n_2808)
);

NAND2xp5_ASAP7_75t_SL g2809 ( 
.A(n_2330),
.B(n_1791),
.Y(n_2809)
);

NAND2xp5_ASAP7_75t_L g2810 ( 
.A(n_2497),
.B(n_1820),
.Y(n_2810)
);

INVx2_ASAP7_75t_L g2811 ( 
.A(n_2460),
.Y(n_2811)
);

NAND2xp5_ASAP7_75t_SL g2812 ( 
.A(n_2613),
.B(n_1791),
.Y(n_2812)
);

BUFx3_ASAP7_75t_L g2813 ( 
.A(n_2335),
.Y(n_2813)
);

AO22x2_ASAP7_75t_L g2814 ( 
.A1(n_2557),
.A2(n_62),
.B1(n_59),
.B2(n_61),
.Y(n_2814)
);

NOR2xp33_ASAP7_75t_L g2815 ( 
.A(n_2364),
.B(n_1791),
.Y(n_2815)
);

NAND2xp5_ASAP7_75t_L g2816 ( 
.A(n_2506),
.B(n_1820),
.Y(n_2816)
);

BUFx2_ASAP7_75t_L g2817 ( 
.A(n_2402),
.Y(n_2817)
);

INVx2_ASAP7_75t_SL g2818 ( 
.A(n_2518),
.Y(n_2818)
);

INVx4_ASAP7_75t_L g2819 ( 
.A(n_2321),
.Y(n_2819)
);

BUFx6f_ASAP7_75t_L g2820 ( 
.A(n_2498),
.Y(n_2820)
);

AND2x4_ASAP7_75t_L g2821 ( 
.A(n_2572),
.B(n_1809),
.Y(n_2821)
);

BUFx3_ASAP7_75t_L g2822 ( 
.A(n_2321),
.Y(n_2822)
);

INVx2_ASAP7_75t_L g2823 ( 
.A(n_2461),
.Y(n_2823)
);

NAND3xp33_ASAP7_75t_L g2824 ( 
.A(n_2491),
.B(n_1811),
.C(n_1809),
.Y(n_2824)
);

BUFx6f_ASAP7_75t_L g2825 ( 
.A(n_2350),
.Y(n_2825)
);

AND2x4_ASAP7_75t_L g2826 ( 
.A(n_2585),
.B(n_1809),
.Y(n_2826)
);

BUFx6f_ASAP7_75t_L g2827 ( 
.A(n_2350),
.Y(n_2827)
);

AO22x2_ASAP7_75t_L g2828 ( 
.A1(n_2565),
.A2(n_64),
.B1(n_62),
.B2(n_63),
.Y(n_2828)
);

INVx1_ASAP7_75t_SL g2829 ( 
.A(n_2487),
.Y(n_2829)
);

OAI22xp33_ASAP7_75t_L g2830 ( 
.A1(n_2537),
.A2(n_1820),
.B1(n_1811),
.B2(n_1809),
.Y(n_2830)
);

INVxp67_ASAP7_75t_L g2831 ( 
.A(n_2364),
.Y(n_2831)
);

INVx2_ASAP7_75t_SL g2832 ( 
.A(n_2518),
.Y(n_2832)
);

INVxp33_ASAP7_75t_L g2833 ( 
.A(n_2487),
.Y(n_2833)
);

AND2x4_ASAP7_75t_L g2834 ( 
.A(n_2585),
.B(n_1811),
.Y(n_2834)
);

INVx2_ASAP7_75t_L g2835 ( 
.A(n_2461),
.Y(n_2835)
);

NAND2xp5_ASAP7_75t_SL g2836 ( 
.A(n_2613),
.B(n_1811),
.Y(n_2836)
);

AO22x2_ASAP7_75t_L g2837 ( 
.A1(n_2565),
.A2(n_2569),
.B1(n_2611),
.B2(n_2592),
.Y(n_2837)
);

INVx1_ASAP7_75t_L g2838 ( 
.A(n_2322),
.Y(n_2838)
);

NAND2xp5_ASAP7_75t_SL g2839 ( 
.A(n_2613),
.B(n_1821),
.Y(n_2839)
);

INVx2_ASAP7_75t_L g2840 ( 
.A(n_2462),
.Y(n_2840)
);

INVx1_ASAP7_75t_L g2841 ( 
.A(n_2322),
.Y(n_2841)
);

INVx1_ASAP7_75t_L g2842 ( 
.A(n_2324),
.Y(n_2842)
);

INVx8_ASAP7_75t_L g2843 ( 
.A(n_2326),
.Y(n_2843)
);

AND3x1_ASAP7_75t_L g2844 ( 
.A(n_2641),
.B(n_1715),
.C(n_62),
.Y(n_2844)
);

NAND2x1p5_ASAP7_75t_L g2845 ( 
.A(n_2473),
.B(n_1821),
.Y(n_2845)
);

INVx2_ASAP7_75t_L g2846 ( 
.A(n_2462),
.Y(n_2846)
);

INVx4_ASAP7_75t_L g2847 ( 
.A(n_2323),
.Y(n_2847)
);

AND2x2_ASAP7_75t_L g2848 ( 
.A(n_2555),
.B(n_1821),
.Y(n_2848)
);

CKINVDCx5p33_ASAP7_75t_R g2849 ( 
.A(n_2402),
.Y(n_2849)
);

AND2x2_ASAP7_75t_L g2850 ( 
.A(n_2602),
.B(n_1821),
.Y(n_2850)
);

INVx1_ASAP7_75t_L g2851 ( 
.A(n_2324),
.Y(n_2851)
);

INVx2_ASAP7_75t_L g2852 ( 
.A(n_2464),
.Y(n_2852)
);

INVx1_ASAP7_75t_L g2853 ( 
.A(n_2325),
.Y(n_2853)
);

INVx2_ASAP7_75t_L g2854 ( 
.A(n_2464),
.Y(n_2854)
);

AND2x2_ASAP7_75t_L g2855 ( 
.A(n_2559),
.B(n_1823),
.Y(n_2855)
);

INVxp67_ASAP7_75t_L g2856 ( 
.A(n_2568),
.Y(n_2856)
);

INVx1_ASAP7_75t_L g2857 ( 
.A(n_2325),
.Y(n_2857)
);

NAND2x1p5_ASAP7_75t_L g2858 ( 
.A(n_2473),
.B(n_1823),
.Y(n_2858)
);

AND2x2_ASAP7_75t_L g2859 ( 
.A(n_2560),
.B(n_1823),
.Y(n_2859)
);

NAND2xp5_ASAP7_75t_L g2860 ( 
.A(n_2506),
.B(n_1823),
.Y(n_2860)
);

INVx2_ASAP7_75t_L g2861 ( 
.A(n_2467),
.Y(n_2861)
);

INVx2_ASAP7_75t_L g2862 ( 
.A(n_2467),
.Y(n_2862)
);

BUFx3_ASAP7_75t_L g2863 ( 
.A(n_2563),
.Y(n_2863)
);

INVx2_ASAP7_75t_L g2864 ( 
.A(n_2480),
.Y(n_2864)
);

AND2x2_ASAP7_75t_L g2865 ( 
.A(n_2561),
.B(n_695),
.Y(n_2865)
);

INVx1_ASAP7_75t_L g2866 ( 
.A(n_2329),
.Y(n_2866)
);

INVxp67_ASAP7_75t_SL g2867 ( 
.A(n_2329),
.Y(n_2867)
);

OR2x2_ASAP7_75t_L g2868 ( 
.A(n_2568),
.B(n_1715),
.Y(n_2868)
);

INVx4_ASAP7_75t_L g2869 ( 
.A(n_2323),
.Y(n_2869)
);

HB1xp67_ASAP7_75t_L g2870 ( 
.A(n_2344),
.Y(n_2870)
);

INVx2_ASAP7_75t_L g2871 ( 
.A(n_2480),
.Y(n_2871)
);

NAND2xp5_ASAP7_75t_L g2872 ( 
.A(n_2547),
.B(n_1715),
.Y(n_2872)
);

INVxp67_ASAP7_75t_L g2873 ( 
.A(n_2593),
.Y(n_2873)
);

INVx1_ASAP7_75t_L g2874 ( 
.A(n_2332),
.Y(n_2874)
);

NAND2xp5_ASAP7_75t_L g2875 ( 
.A(n_2332),
.B(n_1710),
.Y(n_2875)
);

NAND2x1p5_ASAP7_75t_L g2876 ( 
.A(n_2473),
.B(n_1710),
.Y(n_2876)
);

OR2x2_ASAP7_75t_SL g2877 ( 
.A(n_2465),
.B(n_63),
.Y(n_2877)
);

AND2x2_ASAP7_75t_L g2878 ( 
.A(n_2657),
.B(n_696),
.Y(n_2878)
);

BUFx3_ASAP7_75t_L g2879 ( 
.A(n_2563),
.Y(n_2879)
);

OAI22xp5_ASAP7_75t_L g2880 ( 
.A1(n_2441),
.A2(n_1714),
.B1(n_1719),
.B2(n_1710),
.Y(n_2880)
);

INVx1_ASAP7_75t_L g2881 ( 
.A(n_2334),
.Y(n_2881)
);

INVx2_ASAP7_75t_L g2882 ( 
.A(n_2485),
.Y(n_2882)
);

NAND2xp5_ASAP7_75t_L g2883 ( 
.A(n_2334),
.B(n_1710),
.Y(n_2883)
);

INVx4_ASAP7_75t_L g2884 ( 
.A(n_2323),
.Y(n_2884)
);

INVx1_ASAP7_75t_L g2885 ( 
.A(n_2351),
.Y(n_2885)
);

INVx1_ASAP7_75t_L g2886 ( 
.A(n_2351),
.Y(n_2886)
);

INVx1_ASAP7_75t_L g2887 ( 
.A(n_2360),
.Y(n_2887)
);

INVx2_ASAP7_75t_L g2888 ( 
.A(n_2485),
.Y(n_2888)
);

INVx1_ASAP7_75t_SL g2889 ( 
.A(n_2593),
.Y(n_2889)
);

CKINVDCx5p33_ASAP7_75t_R g2890 ( 
.A(n_2352),
.Y(n_2890)
);

INVx1_ASAP7_75t_L g2891 ( 
.A(n_2360),
.Y(n_2891)
);

AND2x2_ASAP7_75t_L g2892 ( 
.A(n_2657),
.B(n_696),
.Y(n_2892)
);

INVx1_ASAP7_75t_L g2893 ( 
.A(n_2456),
.Y(n_2893)
);

AND2x4_ASAP7_75t_L g2894 ( 
.A(n_2585),
.B(n_1714),
.Y(n_2894)
);

BUFx6f_ASAP7_75t_L g2895 ( 
.A(n_2323),
.Y(n_2895)
);

INVx2_ASAP7_75t_L g2896 ( 
.A(n_2316),
.Y(n_2896)
);

INVx2_ASAP7_75t_L g2897 ( 
.A(n_2316),
.Y(n_2897)
);

INVx1_ASAP7_75t_L g2898 ( 
.A(n_2472),
.Y(n_2898)
);

AO22x2_ASAP7_75t_L g2899 ( 
.A1(n_2569),
.A2(n_65),
.B1(n_63),
.B2(n_64),
.Y(n_2899)
);

INVx1_ASAP7_75t_L g2900 ( 
.A(n_2432),
.Y(n_2900)
);

INVxp67_ASAP7_75t_L g2901 ( 
.A(n_2510),
.Y(n_2901)
);

INVx1_ASAP7_75t_L g2902 ( 
.A(n_2442),
.Y(n_2902)
);

AND2x4_ASAP7_75t_L g2903 ( 
.A(n_2417),
.B(n_1714),
.Y(n_2903)
);

BUFx6f_ASAP7_75t_L g2904 ( 
.A(n_2339),
.Y(n_2904)
);

INVx2_ASAP7_75t_L g2905 ( 
.A(n_2471),
.Y(n_2905)
);

BUFx6f_ASAP7_75t_L g2906 ( 
.A(n_2339),
.Y(n_2906)
);

INVx1_ASAP7_75t_L g2907 ( 
.A(n_2445),
.Y(n_2907)
);

INVx2_ASAP7_75t_L g2908 ( 
.A(n_2471),
.Y(n_2908)
);

BUFx3_ASAP7_75t_L g2909 ( 
.A(n_2331),
.Y(n_2909)
);

INVx1_ASAP7_75t_L g2910 ( 
.A(n_2446),
.Y(n_2910)
);

INVx1_ASAP7_75t_L g2911 ( 
.A(n_2447),
.Y(n_2911)
);

NAND2xp5_ASAP7_75t_L g2912 ( 
.A(n_2656),
.B(n_2594),
.Y(n_2912)
);

INVx2_ASAP7_75t_SL g2913 ( 
.A(n_2630),
.Y(n_2913)
);

NAND2xp5_ASAP7_75t_L g2914 ( 
.A(n_2656),
.B(n_1714),
.Y(n_2914)
);

NAND2xp33_ASAP7_75t_R g2915 ( 
.A(n_2365),
.B(n_64),
.Y(n_2915)
);

INVx1_ASAP7_75t_L g2916 ( 
.A(n_2451),
.Y(n_2916)
);

BUFx3_ASAP7_75t_L g2917 ( 
.A(n_2331),
.Y(n_2917)
);

BUFx2_ASAP7_75t_L g2918 ( 
.A(n_2326),
.Y(n_2918)
);

AND2x4_ASAP7_75t_L g2919 ( 
.A(n_2417),
.B(n_1719),
.Y(n_2919)
);

INVx4_ASAP7_75t_L g2920 ( 
.A(n_2339),
.Y(n_2920)
);

INVx3_ASAP7_75t_L g2921 ( 
.A(n_2357),
.Y(n_2921)
);

BUFx6f_ASAP7_75t_L g2922 ( 
.A(n_2339),
.Y(n_2922)
);

INVx4_ASAP7_75t_L g2923 ( 
.A(n_2373),
.Y(n_2923)
);

NOR2xp33_ASAP7_75t_L g2924 ( 
.A(n_2484),
.B(n_1719),
.Y(n_2924)
);

INVx2_ASAP7_75t_L g2925 ( 
.A(n_2471),
.Y(n_2925)
);

NAND2xp5_ASAP7_75t_L g2926 ( 
.A(n_2599),
.B(n_2600),
.Y(n_2926)
);

AND2x4_ASAP7_75t_L g2927 ( 
.A(n_2417),
.B(n_1719),
.Y(n_2927)
);

BUFx6f_ASAP7_75t_L g2928 ( 
.A(n_2404),
.Y(n_2928)
);

INVx3_ASAP7_75t_L g2929 ( 
.A(n_2357),
.Y(n_2929)
);

OR2x2_ASAP7_75t_L g2930 ( 
.A(n_2522),
.B(n_144),
.Y(n_2930)
);

INVx1_ASAP7_75t_L g2931 ( 
.A(n_2458),
.Y(n_2931)
);

BUFx6f_ASAP7_75t_L g2932 ( 
.A(n_2404),
.Y(n_2932)
);

INVxp67_ASAP7_75t_L g2933 ( 
.A(n_2511),
.Y(n_2933)
);

OAI22xp5_ASAP7_75t_L g2934 ( 
.A1(n_2612),
.A2(n_67),
.B1(n_65),
.B2(n_66),
.Y(n_2934)
);

INVx1_ASAP7_75t_L g2935 ( 
.A(n_2463),
.Y(n_2935)
);

BUFx6f_ASAP7_75t_L g2936 ( 
.A(n_2405),
.Y(n_2936)
);

INVx2_ASAP7_75t_L g2937 ( 
.A(n_2486),
.Y(n_2937)
);

INVx1_ASAP7_75t_L g2938 ( 
.A(n_2466),
.Y(n_2938)
);

BUFx2_ASAP7_75t_L g2939 ( 
.A(n_2326),
.Y(n_2939)
);

AND2x4_ASAP7_75t_L g2940 ( 
.A(n_2457),
.B(n_145),
.Y(n_2940)
);

AND2x2_ASAP7_75t_L g2941 ( 
.A(n_2588),
.B(n_680),
.Y(n_2941)
);

AND2x2_ASAP7_75t_L g2942 ( 
.A(n_2588),
.B(n_680),
.Y(n_2942)
);

INVx1_ASAP7_75t_L g2943 ( 
.A(n_2474),
.Y(n_2943)
);

INVx1_ASAP7_75t_L g2944 ( 
.A(n_2475),
.Y(n_2944)
);

INVx2_ASAP7_75t_L g2945 ( 
.A(n_2486),
.Y(n_2945)
);

INVx2_ASAP7_75t_L g2946 ( 
.A(n_2486),
.Y(n_2946)
);

HB1xp67_ASAP7_75t_L g2947 ( 
.A(n_2509),
.Y(n_2947)
);

BUFx6f_ASAP7_75t_L g2948 ( 
.A(n_2405),
.Y(n_2948)
);

NOR2xp33_ASAP7_75t_L g2949 ( 
.A(n_2416),
.B(n_681),
.Y(n_2949)
);

BUFx6f_ASAP7_75t_L g2950 ( 
.A(n_2434),
.Y(n_2950)
);

INVx1_ASAP7_75t_L g2951 ( 
.A(n_2479),
.Y(n_2951)
);

INVx2_ASAP7_75t_L g2952 ( 
.A(n_2437),
.Y(n_2952)
);

AND2x4_ASAP7_75t_L g2953 ( 
.A(n_2457),
.B(n_146),
.Y(n_2953)
);

INVx3_ASAP7_75t_L g2954 ( 
.A(n_2380),
.Y(n_2954)
);

AO22x1_ASAP7_75t_L g2955 ( 
.A1(n_2578),
.A2(n_2628),
.B1(n_2342),
.B2(n_2526),
.Y(n_2955)
);

AND2x4_ASAP7_75t_L g2956 ( 
.A(n_2457),
.B(n_147),
.Y(n_2956)
);

AND2x6_ASAP7_75t_L g2957 ( 
.A(n_2509),
.B(n_66),
.Y(n_2957)
);

INVx1_ASAP7_75t_L g2958 ( 
.A(n_2437),
.Y(n_2958)
);

AND2x4_ASAP7_75t_L g2959 ( 
.A(n_2468),
.B(n_147),
.Y(n_2959)
);

AND2x6_ASAP7_75t_L g2960 ( 
.A(n_2512),
.B(n_66),
.Y(n_2960)
);

OR2x2_ASAP7_75t_SL g2961 ( 
.A(n_2609),
.B(n_68),
.Y(n_2961)
);

BUFx3_ASAP7_75t_L g2962 ( 
.A(n_2331),
.Y(n_2962)
);

NAND2xp5_ASAP7_75t_L g2963 ( 
.A(n_2801),
.B(n_2661),
.Y(n_2963)
);

AOI22xp33_ASAP7_75t_L g2964 ( 
.A1(n_2699),
.A2(n_2564),
.B1(n_2567),
.B2(n_2652),
.Y(n_2964)
);

INVx2_ASAP7_75t_L g2965 ( 
.A(n_2674),
.Y(n_2965)
);

NAND2xp5_ASAP7_75t_SL g2966 ( 
.A(n_2829),
.B(n_2588),
.Y(n_2966)
);

INVx2_ASAP7_75t_L g2967 ( 
.A(n_2675),
.Y(n_2967)
);

NAND2xp5_ASAP7_75t_L g2968 ( 
.A(n_2781),
.B(n_2601),
.Y(n_2968)
);

INVx1_ASAP7_75t_L g2969 ( 
.A(n_2947),
.Y(n_2969)
);

NOR2xp67_ASAP7_75t_L g2970 ( 
.A(n_2673),
.B(n_2636),
.Y(n_2970)
);

NOR2xp33_ASAP7_75t_L g2971 ( 
.A(n_2782),
.B(n_2416),
.Y(n_2971)
);

AOI22xp33_ASAP7_75t_L g2972 ( 
.A1(n_2691),
.A2(n_2564),
.B1(n_2567),
.B2(n_2652),
.Y(n_2972)
);

NAND2xp5_ASAP7_75t_SL g2973 ( 
.A(n_2829),
.B(n_2635),
.Y(n_2973)
);

INVxp67_ASAP7_75t_L g2974 ( 
.A(n_2870),
.Y(n_2974)
);

INVx2_ASAP7_75t_L g2975 ( 
.A(n_2687),
.Y(n_2975)
);

INVx5_ASAP7_75t_L g2976 ( 
.A(n_2923),
.Y(n_2976)
);

INVx4_ASAP7_75t_L g2977 ( 
.A(n_2673),
.Y(n_2977)
);

AOI22xp33_ASAP7_75t_L g2978 ( 
.A1(n_2671),
.A2(n_2564),
.B1(n_2567),
.B2(n_2652),
.Y(n_2978)
);

INVx1_ASAP7_75t_L g2979 ( 
.A(n_2947),
.Y(n_2979)
);

NAND2xp5_ASAP7_75t_L g2980 ( 
.A(n_2781),
.B(n_2625),
.Y(n_2980)
);

BUFx3_ASAP7_75t_L g2981 ( 
.A(n_2822),
.Y(n_2981)
);

INVx3_ASAP7_75t_L g2982 ( 
.A(n_2680),
.Y(n_2982)
);

INVx1_ASAP7_75t_L g2983 ( 
.A(n_2958),
.Y(n_2983)
);

NAND2xp5_ASAP7_75t_L g2984 ( 
.A(n_2867),
.B(n_2587),
.Y(n_2984)
);

AND2x2_ASAP7_75t_L g2985 ( 
.A(n_2746),
.B(n_2621),
.Y(n_2985)
);

AOI22xp5_ASAP7_75t_L g2986 ( 
.A1(n_2670),
.A2(n_2574),
.B1(n_2352),
.B2(n_2635),
.Y(n_2986)
);

AND2x4_ASAP7_75t_L g2987 ( 
.A(n_2697),
.B(n_2397),
.Y(n_2987)
);

NAND2xp5_ASAP7_75t_L g2988 ( 
.A(n_2734),
.B(n_2665),
.Y(n_2988)
);

NAND2xp5_ASAP7_75t_L g2989 ( 
.A(n_2734),
.B(n_2640),
.Y(n_2989)
);

NOR2xp33_ASAP7_75t_L g2990 ( 
.A(n_2833),
.B(n_2342),
.Y(n_2990)
);

NOR2xp33_ASAP7_75t_R g2991 ( 
.A(n_2849),
.B(n_2403),
.Y(n_2991)
);

NAND2xp5_ASAP7_75t_L g2992 ( 
.A(n_2926),
.B(n_2640),
.Y(n_2992)
);

INVx1_ASAP7_75t_SL g2993 ( 
.A(n_2773),
.Y(n_2993)
);

NOR2xp33_ASAP7_75t_L g2994 ( 
.A(n_2889),
.B(n_2503),
.Y(n_2994)
);

INVx4_ASAP7_75t_L g2995 ( 
.A(n_2819),
.Y(n_2995)
);

AND2x6_ASAP7_75t_SL g2996 ( 
.A(n_2676),
.B(n_2645),
.Y(n_2996)
);

INVx2_ASAP7_75t_SL g2997 ( 
.A(n_2825),
.Y(n_2997)
);

NAND2xp5_ASAP7_75t_L g2998 ( 
.A(n_2926),
.B(n_2650),
.Y(n_2998)
);

NAND2x1_ASAP7_75t_L g2999 ( 
.A(n_2923),
.B(n_2380),
.Y(n_2999)
);

INVx2_ASAP7_75t_L g3000 ( 
.A(n_2706),
.Y(n_3000)
);

NOR2xp33_ASAP7_75t_L g3001 ( 
.A(n_2889),
.B(n_2773),
.Y(n_3001)
);

INVx1_ASAP7_75t_L g3002 ( 
.A(n_2744),
.Y(n_3002)
);

NAND2xp5_ASAP7_75t_L g3003 ( 
.A(n_2693),
.B(n_2650),
.Y(n_3003)
);

NOR2x2_ASAP7_75t_L g3004 ( 
.A(n_2741),
.B(n_2554),
.Y(n_3004)
);

AOI22xp33_ASAP7_75t_L g3005 ( 
.A1(n_2671),
.A2(n_2352),
.B1(n_2578),
.B2(n_2612),
.Y(n_3005)
);

INVx1_ASAP7_75t_L g3006 ( 
.A(n_2748),
.Y(n_3006)
);

NAND2xp5_ASAP7_75t_L g3007 ( 
.A(n_2693),
.B(n_2658),
.Y(n_3007)
);

NOR2xp33_ASAP7_75t_L g3008 ( 
.A(n_2786),
.B(n_2634),
.Y(n_3008)
);

AOI22xp5_ASAP7_75t_L g3009 ( 
.A1(n_2760),
.A2(n_2635),
.B1(n_2583),
.B2(n_2596),
.Y(n_3009)
);

AND2x2_ASAP7_75t_L g3010 ( 
.A(n_2786),
.B(n_2621),
.Y(n_3010)
);

BUFx3_ASAP7_75t_L g3011 ( 
.A(n_2718),
.Y(n_3011)
);

NAND2xp5_ASAP7_75t_SL g3012 ( 
.A(n_2720),
.B(n_2589),
.Y(n_3012)
);

NAND2xp5_ASAP7_75t_SL g3013 ( 
.A(n_2856),
.B(n_2589),
.Y(n_3013)
);

NOR2xp33_ASAP7_75t_SL g3014 ( 
.A(n_2819),
.B(n_2531),
.Y(n_3014)
);

INVx8_ASAP7_75t_L g3015 ( 
.A(n_2713),
.Y(n_3015)
);

AND2x2_ASAP7_75t_L g3016 ( 
.A(n_2738),
.B(n_2612),
.Y(n_3016)
);

NOR2xp33_ASAP7_75t_L g3017 ( 
.A(n_2856),
.B(n_2644),
.Y(n_3017)
);

AOI21xp5_ASAP7_75t_L g3018 ( 
.A1(n_2703),
.A2(n_2338),
.B(n_2508),
.Y(n_3018)
);

INVx1_ASAP7_75t_L g3019 ( 
.A(n_2752),
.Y(n_3019)
);

INVx1_ASAP7_75t_L g3020 ( 
.A(n_2753),
.Y(n_3020)
);

OAI22xp33_ASAP7_75t_L g3021 ( 
.A1(n_2704),
.A2(n_2578),
.B1(n_2589),
.B2(n_2328),
.Y(n_3021)
);

NAND2xp5_ASAP7_75t_L g3022 ( 
.A(n_2728),
.B(n_2658),
.Y(n_3022)
);

INVx2_ASAP7_75t_L g3023 ( 
.A(n_2712),
.Y(n_3023)
);

OR2x2_ASAP7_75t_L g3024 ( 
.A(n_2672),
.B(n_2644),
.Y(n_3024)
);

NAND2xp5_ASAP7_75t_L g3025 ( 
.A(n_2728),
.B(n_2663),
.Y(n_3025)
);

AND2x2_ASAP7_75t_L g3026 ( 
.A(n_2873),
.B(n_2632),
.Y(n_3026)
);

NAND2xp5_ASAP7_75t_L g3027 ( 
.A(n_2912),
.B(n_2663),
.Y(n_3027)
);

A2O1A1Ixp33_ASAP7_75t_L g3028 ( 
.A1(n_2901),
.A2(n_2320),
.B(n_2492),
.C(n_2513),
.Y(n_3028)
);

NOR2xp33_ASAP7_75t_L g3029 ( 
.A(n_2873),
.B(n_2624),
.Y(n_3029)
);

NAND2xp5_ASAP7_75t_L g3030 ( 
.A(n_2912),
.B(n_2664),
.Y(n_3030)
);

NAND2xp5_ASAP7_75t_L g3031 ( 
.A(n_2901),
.B(n_2664),
.Y(n_3031)
);

INVx1_ASAP7_75t_L g3032 ( 
.A(n_2754),
.Y(n_3032)
);

NOR2xp33_ASAP7_75t_L g3033 ( 
.A(n_2672),
.B(n_2624),
.Y(n_3033)
);

NAND2xp5_ASAP7_75t_L g3034 ( 
.A(n_2933),
.B(n_2541),
.Y(n_3034)
);

NAND2xp5_ASAP7_75t_L g3035 ( 
.A(n_2933),
.B(n_2633),
.Y(n_3035)
);

NAND2xp5_ASAP7_75t_L g3036 ( 
.A(n_2867),
.B(n_2390),
.Y(n_3036)
);

INVx2_ASAP7_75t_SL g3037 ( 
.A(n_2825),
.Y(n_3037)
);

NAND2xp5_ASAP7_75t_L g3038 ( 
.A(n_2684),
.B(n_2647),
.Y(n_3038)
);

INVxp67_ASAP7_75t_L g3039 ( 
.A(n_2870),
.Y(n_3039)
);

NAND2xp5_ASAP7_75t_L g3040 ( 
.A(n_2684),
.B(n_2648),
.Y(n_3040)
);

INVx2_ASAP7_75t_L g3041 ( 
.A(n_2717),
.Y(n_3041)
);

A2O1A1Ixp33_ASAP7_75t_L g3042 ( 
.A1(n_2924),
.A2(n_2320),
.B(n_2492),
.C(n_2429),
.Y(n_3042)
);

NAND2xp5_ASAP7_75t_L g3043 ( 
.A(n_2763),
.B(n_2521),
.Y(n_3043)
);

BUFx6f_ASAP7_75t_L g3044 ( 
.A(n_2825),
.Y(n_3044)
);

AOI22xp33_ASAP7_75t_L g3045 ( 
.A1(n_2671),
.A2(n_2655),
.B1(n_2582),
.B2(n_2637),
.Y(n_3045)
);

OR2x2_ASAP7_75t_L g3046 ( 
.A(n_2913),
.B(n_2709),
.Y(n_3046)
);

NAND2xp5_ASAP7_75t_L g3047 ( 
.A(n_2763),
.B(n_2654),
.Y(n_3047)
);

NAND2xp5_ASAP7_75t_SL g3048 ( 
.A(n_2705),
.B(n_2589),
.Y(n_3048)
);

NAND2xp5_ASAP7_75t_L g3049 ( 
.A(n_2768),
.B(n_2893),
.Y(n_3049)
);

OAI22xp33_ASAP7_75t_L g3050 ( 
.A1(n_2704),
.A2(n_2589),
.B1(n_2328),
.B2(n_2654),
.Y(n_3050)
);

NOR2xp33_ASAP7_75t_L g3051 ( 
.A(n_2695),
.B(n_2624),
.Y(n_3051)
);

INVx3_ASAP7_75t_L g3052 ( 
.A(n_2680),
.Y(n_3052)
);

NAND2xp5_ASAP7_75t_SL g3053 ( 
.A(n_2775),
.B(n_2403),
.Y(n_3053)
);

NAND2xp5_ASAP7_75t_L g3054 ( 
.A(n_2768),
.B(n_2654),
.Y(n_3054)
);

INVx1_ASAP7_75t_L g3055 ( 
.A(n_2761),
.Y(n_3055)
);

NAND2xp5_ASAP7_75t_SL g3056 ( 
.A(n_2818),
.B(n_2370),
.Y(n_3056)
);

O2A1O1Ixp33_ASAP7_75t_L g3057 ( 
.A1(n_2739),
.A2(n_2655),
.B(n_2517),
.C(n_2400),
.Y(n_3057)
);

INVx1_ASAP7_75t_L g3058 ( 
.A(n_2762),
.Y(n_3058)
);

NAND2xp5_ASAP7_75t_SL g3059 ( 
.A(n_2832),
.B(n_2370),
.Y(n_3059)
);

AOI22xp5_ASAP7_75t_L g3060 ( 
.A1(n_2676),
.A2(n_2605),
.B1(n_2627),
.B2(n_2581),
.Y(n_3060)
);

NOR3x1_ASAP7_75t_L g3061 ( 
.A(n_2955),
.B(n_2604),
.C(n_2620),
.Y(n_3061)
);

INVx2_ASAP7_75t_L g3062 ( 
.A(n_2732),
.Y(n_3062)
);

INVx2_ASAP7_75t_SL g3063 ( 
.A(n_2827),
.Y(n_3063)
);

AOI22xp5_ASAP7_75t_L g3064 ( 
.A1(n_2692),
.A2(n_2581),
.B1(n_2400),
.B2(n_2353),
.Y(n_3064)
);

NAND2xp5_ASAP7_75t_L g3065 ( 
.A(n_2898),
.B(n_2654),
.Y(n_3065)
);

INVx2_ASAP7_75t_L g3066 ( 
.A(n_2896),
.Y(n_3066)
);

O2A1O1Ixp33_ASAP7_75t_L g3067 ( 
.A1(n_2715),
.A2(n_2517),
.B(n_2495),
.C(n_2642),
.Y(n_3067)
);

NAND2xp5_ASAP7_75t_L g3068 ( 
.A(n_2690),
.B(n_2654),
.Y(n_3068)
);

NAND2xp5_ASAP7_75t_L g3069 ( 
.A(n_2690),
.B(n_2527),
.Y(n_3069)
);

NAND2xp5_ASAP7_75t_SL g3070 ( 
.A(n_2827),
.B(n_2376),
.Y(n_3070)
);

AOI22xp5_ASAP7_75t_L g3071 ( 
.A1(n_2692),
.A2(n_2353),
.B1(n_2528),
.B2(n_2495),
.Y(n_3071)
);

AOI22xp5_ASAP7_75t_L g3072 ( 
.A1(n_2701),
.A2(n_2528),
.B1(n_2604),
.B2(n_2519),
.Y(n_3072)
);

NAND2xp5_ASAP7_75t_L g3073 ( 
.A(n_2878),
.B(n_2533),
.Y(n_3073)
);

AOI22xp33_ASAP7_75t_L g3074 ( 
.A1(n_2671),
.A2(n_2582),
.B1(n_2637),
.B2(n_2528),
.Y(n_3074)
);

INVx1_ASAP7_75t_L g3075 ( 
.A(n_2765),
.Y(n_3075)
);

NAND2xp5_ASAP7_75t_L g3076 ( 
.A(n_2892),
.B(n_2536),
.Y(n_3076)
);

NAND2xp5_ASAP7_75t_SL g3077 ( 
.A(n_2827),
.B(n_2376),
.Y(n_3077)
);

INVx1_ASAP7_75t_L g3078 ( 
.A(n_2772),
.Y(n_3078)
);

XNOR2xp5_ASAP7_75t_L g3079 ( 
.A(n_2730),
.B(n_2629),
.Y(n_3079)
);

NOR2xp33_ASAP7_75t_L g3080 ( 
.A(n_2831),
.B(n_2592),
.Y(n_3080)
);

AND2x2_ASAP7_75t_L g3081 ( 
.A(n_2865),
.B(n_2355),
.Y(n_3081)
);

AOI22xp33_ASAP7_75t_L g3082 ( 
.A1(n_2689),
.A2(n_2637),
.B1(n_2611),
.B2(n_2592),
.Y(n_3082)
);

INVx1_ASAP7_75t_L g3083 ( 
.A(n_2952),
.Y(n_3083)
);

INVx1_ASAP7_75t_L g3084 ( 
.A(n_2777),
.Y(n_3084)
);

NAND2xp5_ASAP7_75t_SL g3085 ( 
.A(n_2817),
.B(n_2831),
.Y(n_3085)
);

NAND2xp5_ASAP7_75t_L g3086 ( 
.A(n_2700),
.B(n_2512),
.Y(n_3086)
);

CKINVDCx5p33_ASAP7_75t_R g3087 ( 
.A(n_2751),
.Y(n_3087)
);

NAND2xp5_ASAP7_75t_L g3088 ( 
.A(n_2700),
.B(n_2529),
.Y(n_3088)
);

NAND2xp5_ASAP7_75t_L g3089 ( 
.A(n_2793),
.B(n_2529),
.Y(n_3089)
);

NAND2xp5_ASAP7_75t_L g3090 ( 
.A(n_2792),
.B(n_2499),
.Y(n_3090)
);

NAND2xp5_ASAP7_75t_L g3091 ( 
.A(n_2792),
.B(n_2532),
.Y(n_3091)
);

AOI22xp5_ASAP7_75t_L g3092 ( 
.A1(n_2915),
.A2(n_2519),
.B1(n_2315),
.B2(n_2606),
.Y(n_3092)
);

NAND2xp5_ASAP7_75t_L g3093 ( 
.A(n_2798),
.B(n_2532),
.Y(n_3093)
);

NAND2xp5_ASAP7_75t_L g3094 ( 
.A(n_2802),
.B(n_2534),
.Y(n_3094)
);

INVx2_ASAP7_75t_L g3095 ( 
.A(n_2897),
.Y(n_3095)
);

BUFx3_ASAP7_75t_L g3096 ( 
.A(n_2787),
.Y(n_3096)
);

NAND2xp5_ASAP7_75t_L g3097 ( 
.A(n_2804),
.B(n_2534),
.Y(n_3097)
);

NAND2xp5_ASAP7_75t_L g3098 ( 
.A(n_2806),
.B(n_2535),
.Y(n_3098)
);

INVx1_ASAP7_75t_L g3099 ( 
.A(n_2780),
.Y(n_3099)
);

NAND2xp5_ASAP7_75t_L g3100 ( 
.A(n_2838),
.B(n_2535),
.Y(n_3100)
);

AND2x2_ASAP7_75t_L g3101 ( 
.A(n_2689),
.B(n_2355),
.Y(n_3101)
);

NAND2xp5_ASAP7_75t_L g3102 ( 
.A(n_2841),
.B(n_2540),
.Y(n_3102)
);

INVx3_ASAP7_75t_L g3103 ( 
.A(n_2750),
.Y(n_3103)
);

NAND2xp5_ASAP7_75t_SL g3104 ( 
.A(n_2697),
.B(n_2347),
.Y(n_3104)
);

NAND2xp5_ASAP7_75t_L g3105 ( 
.A(n_2784),
.B(n_2540),
.Y(n_3105)
);

AND2x2_ASAP7_75t_L g3106 ( 
.A(n_2941),
.B(n_2355),
.Y(n_3106)
);

NOR2xp67_ASAP7_75t_L g3107 ( 
.A(n_2723),
.B(n_2636),
.Y(n_3107)
);

INVx2_ASAP7_75t_SL g3108 ( 
.A(n_2813),
.Y(n_3108)
);

CKINVDCx5p33_ASAP7_75t_R g3109 ( 
.A(n_2890),
.Y(n_3109)
);

NAND2xp5_ASAP7_75t_L g3110 ( 
.A(n_2842),
.B(n_2554),
.Y(n_3110)
);

NAND2xp5_ASAP7_75t_SL g3111 ( 
.A(n_2677),
.B(n_2347),
.Y(n_3111)
);

NAND2xp5_ASAP7_75t_L g3112 ( 
.A(n_2795),
.B(n_2556),
.Y(n_3112)
);

INVx2_ASAP7_75t_SL g3113 ( 
.A(n_2863),
.Y(n_3113)
);

NAND2xp5_ASAP7_75t_L g3114 ( 
.A(n_2851),
.B(n_2556),
.Y(n_3114)
);

NOR2xp33_ASAP7_75t_L g3115 ( 
.A(n_2677),
.B(n_2611),
.Y(n_3115)
);

INVx1_ASAP7_75t_L g3116 ( 
.A(n_2797),
.Y(n_3116)
);

NAND2xp5_ASAP7_75t_SL g3117 ( 
.A(n_2694),
.B(n_2531),
.Y(n_3117)
);

NAND2xp5_ASAP7_75t_L g3118 ( 
.A(n_2764),
.B(n_2618),
.Y(n_3118)
);

AOI22xp33_ASAP7_75t_L g3119 ( 
.A1(n_2949),
.A2(n_2606),
.B1(n_2646),
.B2(n_2642),
.Y(n_3119)
);

NAND2xp5_ASAP7_75t_L g3120 ( 
.A(n_2742),
.B(n_2618),
.Y(n_3120)
);

OAI22xp33_ASAP7_75t_L g3121 ( 
.A1(n_2742),
.A2(n_2328),
.B1(n_2428),
.B2(n_2412),
.Y(n_3121)
);

NAND2xp5_ASAP7_75t_L g3122 ( 
.A(n_2708),
.B(n_2618),
.Y(n_3122)
);

NAND2xp33_ASAP7_75t_L g3123 ( 
.A(n_2713),
.B(n_2315),
.Y(n_3123)
);

AOI22xp5_ASAP7_75t_L g3124 ( 
.A1(n_2678),
.A2(n_2519),
.B1(n_2315),
.B2(n_2436),
.Y(n_3124)
);

INVxp67_ASAP7_75t_L g3125 ( 
.A(n_2930),
.Y(n_3125)
);

INVx1_ASAP7_75t_L g3126 ( 
.A(n_2853),
.Y(n_3126)
);

NAND2xp5_ASAP7_75t_L g3127 ( 
.A(n_2708),
.B(n_2575),
.Y(n_3127)
);

OR2x6_ASAP7_75t_L g3128 ( 
.A(n_2713),
.B(n_2328),
.Y(n_3128)
);

INVx1_ASAP7_75t_L g3129 ( 
.A(n_2857),
.Y(n_3129)
);

NOR2xp33_ASAP7_75t_R g3130 ( 
.A(n_2879),
.B(n_2422),
.Y(n_3130)
);

BUFx6f_ASAP7_75t_L g3131 ( 
.A(n_2928),
.Y(n_3131)
);

INVx1_ASAP7_75t_L g3132 ( 
.A(n_2866),
.Y(n_3132)
);

INVx8_ASAP7_75t_L g3133 ( 
.A(n_2843),
.Y(n_3133)
);

INVx5_ASAP7_75t_L g3134 ( 
.A(n_2895),
.Y(n_3134)
);

INVx2_ASAP7_75t_L g3135 ( 
.A(n_2679),
.Y(n_3135)
);

AOI22xp33_ASAP7_75t_L g3136 ( 
.A1(n_2783),
.A2(n_2646),
.B1(n_2642),
.B2(n_2622),
.Y(n_3136)
);

INVx1_ASAP7_75t_L g3137 ( 
.A(n_2874),
.Y(n_3137)
);

OAI22xp5_ASAP7_75t_L g3138 ( 
.A1(n_2758),
.A2(n_2483),
.B1(n_2576),
.B2(n_2575),
.Y(n_3138)
);

INVx1_ASAP7_75t_L g3139 ( 
.A(n_2881),
.Y(n_3139)
);

INVx1_ASAP7_75t_L g3140 ( 
.A(n_2885),
.Y(n_3140)
);

INVx1_ASAP7_75t_L g3141 ( 
.A(n_2886),
.Y(n_3141)
);

NAND2xp5_ASAP7_75t_L g3142 ( 
.A(n_2848),
.B(n_2576),
.Y(n_3142)
);

INVx2_ASAP7_75t_L g3143 ( 
.A(n_2681),
.Y(n_3143)
);

OAI22xp5_ASAP7_75t_L g3144 ( 
.A1(n_2758),
.A2(n_2586),
.B1(n_2608),
.B2(n_2598),
.Y(n_3144)
);

NAND2xp5_ASAP7_75t_L g3145 ( 
.A(n_2887),
.B(n_2315),
.Y(n_3145)
);

AOI22xp33_ASAP7_75t_L g3146 ( 
.A1(n_2783),
.A2(n_2646),
.B1(n_2622),
.B2(n_2638),
.Y(n_3146)
);

NAND2xp5_ASAP7_75t_SL g3147 ( 
.A(n_2694),
.B(n_2531),
.Y(n_3147)
);

INVx2_ASAP7_75t_L g3148 ( 
.A(n_2682),
.Y(n_3148)
);

NAND2xp5_ASAP7_75t_L g3149 ( 
.A(n_2755),
.B(n_2586),
.Y(n_3149)
);

INVx1_ASAP7_75t_L g3150 ( 
.A(n_2891),
.Y(n_3150)
);

NAND2xp5_ASAP7_75t_L g3151 ( 
.A(n_2755),
.B(n_2598),
.Y(n_3151)
);

INVx2_ASAP7_75t_L g3152 ( 
.A(n_2686),
.Y(n_3152)
);

OAI22xp5_ASAP7_75t_L g3153 ( 
.A1(n_2830),
.A2(n_2608),
.B1(n_2617),
.B2(n_2610),
.Y(n_3153)
);

NOR3xp33_ASAP7_75t_L g3154 ( 
.A(n_2934),
.B(n_2643),
.C(n_2597),
.Y(n_3154)
);

NOR2xp33_ASAP7_75t_L g3155 ( 
.A(n_2716),
.B(n_2638),
.Y(n_3155)
);

INVx1_ASAP7_75t_L g3156 ( 
.A(n_2688),
.Y(n_3156)
);

NAND2xp5_ASAP7_75t_L g3157 ( 
.A(n_2759),
.B(n_2610),
.Y(n_3157)
);

INVx1_ASAP7_75t_L g3158 ( 
.A(n_2698),
.Y(n_3158)
);

AOI22xp33_ASAP7_75t_L g3159 ( 
.A1(n_2934),
.A2(n_2638),
.B1(n_2653),
.B2(n_2651),
.Y(n_3159)
);

NAND2xp5_ASAP7_75t_L g3160 ( 
.A(n_2759),
.B(n_2617),
.Y(n_3160)
);

INVx2_ASAP7_75t_L g3161 ( 
.A(n_2702),
.Y(n_3161)
);

INVx1_ASAP7_75t_L g3162 ( 
.A(n_2707),
.Y(n_3162)
);

INVx2_ASAP7_75t_L g3163 ( 
.A(n_2711),
.Y(n_3163)
);

INVx2_ASAP7_75t_L g3164 ( 
.A(n_2719),
.Y(n_3164)
);

INVx1_ASAP7_75t_SL g3165 ( 
.A(n_2850),
.Y(n_3165)
);

NAND2xp5_ASAP7_75t_L g3166 ( 
.A(n_2725),
.B(n_2315),
.Y(n_3166)
);

INVx2_ASAP7_75t_SL g3167 ( 
.A(n_2928),
.Y(n_3167)
);

CKINVDCx5p33_ASAP7_75t_R g3168 ( 
.A(n_2716),
.Y(n_3168)
);

NAND2xp5_ASAP7_75t_L g3169 ( 
.A(n_2726),
.B(n_2580),
.Y(n_3169)
);

OAI22xp33_ASAP7_75t_L g3170 ( 
.A1(n_2770),
.A2(n_2412),
.B1(n_2428),
.B2(n_2630),
.Y(n_3170)
);

INVx1_ASAP7_75t_L g3171 ( 
.A(n_2727),
.Y(n_3171)
);

AOI22xp33_ASAP7_75t_L g3172 ( 
.A1(n_2821),
.A2(n_2960),
.B1(n_2957),
.B2(n_2653),
.Y(n_3172)
);

INVx1_ASAP7_75t_L g3173 ( 
.A(n_2731),
.Y(n_3173)
);

NAND2xp5_ASAP7_75t_L g3174 ( 
.A(n_2733),
.B(n_2558),
.Y(n_3174)
);

AO22x1_ASAP7_75t_L g3175 ( 
.A1(n_2957),
.A2(n_2488),
.B1(n_2520),
.B2(n_2636),
.Y(n_3175)
);

AO22x1_ASAP7_75t_L g3176 ( 
.A1(n_2957),
.A2(n_2960),
.B1(n_2953),
.B2(n_2956),
.Y(n_3176)
);

INVx3_ASAP7_75t_L g3177 ( 
.A(n_2750),
.Y(n_3177)
);

INVx1_ASAP7_75t_L g3178 ( 
.A(n_2735),
.Y(n_3178)
);

INVx1_ASAP7_75t_L g3179 ( 
.A(n_2736),
.Y(n_3179)
);

INVx1_ASAP7_75t_L g3180 ( 
.A(n_2737),
.Y(n_3180)
);

INVx1_ASAP7_75t_L g3181 ( 
.A(n_2740),
.Y(n_3181)
);

AND2x4_ASAP7_75t_L g3182 ( 
.A(n_2918),
.B(n_2468),
.Y(n_3182)
);

NOR3x1_ASAP7_75t_L g3183 ( 
.A(n_2939),
.B(n_2425),
.C(n_2597),
.Y(n_3183)
);

INVx1_ASAP7_75t_L g3184 ( 
.A(n_2808),
.Y(n_3184)
);

NOR2xp33_ASAP7_75t_L g3185 ( 
.A(n_2942),
.B(n_2666),
.Y(n_3185)
);

INVx2_ASAP7_75t_SL g3186 ( 
.A(n_2928),
.Y(n_3186)
);

AOI211xp5_ASAP7_75t_L g3187 ( 
.A1(n_3021),
.A2(n_2381),
.B(n_2830),
.C(n_2877),
.Y(n_3187)
);

INVx1_ASAP7_75t_L g3188 ( 
.A(n_3084),
.Y(n_3188)
);

HB1xp67_ASAP7_75t_L g3189 ( 
.A(n_2993),
.Y(n_3189)
);

BUFx12f_ASAP7_75t_SL g3190 ( 
.A(n_3044),
.Y(n_3190)
);

INVx2_ASAP7_75t_L g3191 ( 
.A(n_2965),
.Y(n_3191)
);

NOR2xp67_ASAP7_75t_L g3192 ( 
.A(n_2976),
.B(n_2488),
.Y(n_3192)
);

AOI22xp33_ASAP7_75t_L g3193 ( 
.A1(n_3154),
.A2(n_2651),
.B1(n_2519),
.B2(n_2821),
.Y(n_3193)
);

AOI22xp33_ASAP7_75t_L g3194 ( 
.A1(n_3050),
.A2(n_3051),
.B1(n_2964),
.B2(n_2972),
.Y(n_3194)
);

INVx1_ASAP7_75t_L g3195 ( 
.A(n_3099),
.Y(n_3195)
);

INVx1_ASAP7_75t_L g3196 ( 
.A(n_3116),
.Y(n_3196)
);

INVx1_ASAP7_75t_L g3197 ( 
.A(n_3002),
.Y(n_3197)
);

AOI22xp5_ASAP7_75t_L g3198 ( 
.A1(n_2994),
.A2(n_2844),
.B1(n_2960),
.B2(n_2957),
.Y(n_3198)
);

INVx2_ASAP7_75t_L g3199 ( 
.A(n_2967),
.Y(n_3199)
);

AND2x4_ASAP7_75t_L g3200 ( 
.A(n_3128),
.B(n_2766),
.Y(n_3200)
);

NAND2xp5_ASAP7_75t_L g3201 ( 
.A(n_2963),
.B(n_2837),
.Y(n_3201)
);

NAND2xp5_ASAP7_75t_SL g3202 ( 
.A(n_2986),
.B(n_3060),
.Y(n_3202)
);

INVx5_ASAP7_75t_L g3203 ( 
.A(n_3128),
.Y(n_3203)
);

HB1xp67_ASAP7_75t_L g3204 ( 
.A(n_2993),
.Y(n_3204)
);

CKINVDCx5p33_ASAP7_75t_R g3205 ( 
.A(n_3087),
.Y(n_3205)
);

AOI22xp33_ASAP7_75t_L g3206 ( 
.A1(n_2985),
.A2(n_2643),
.B1(n_2595),
.B2(n_2524),
.Y(n_3206)
);

AND2x6_ASAP7_75t_L g3207 ( 
.A(n_3183),
.B(n_2805),
.Y(n_3207)
);

AND2x2_ASAP7_75t_L g3208 ( 
.A(n_3010),
.B(n_3016),
.Y(n_3208)
);

CKINVDCx20_ASAP7_75t_R g3209 ( 
.A(n_3109),
.Y(n_3209)
);

NAND2xp5_ASAP7_75t_L g3210 ( 
.A(n_2988),
.B(n_2837),
.Y(n_3210)
);

NAND2xp5_ASAP7_75t_SL g3211 ( 
.A(n_3009),
.B(n_2524),
.Y(n_3211)
);

AOI22xp33_ASAP7_75t_SL g3212 ( 
.A1(n_3008),
.A2(n_2774),
.B1(n_2828),
.B2(n_2814),
.Y(n_3212)
);

AND2x2_ASAP7_75t_SL g3213 ( 
.A(n_3123),
.B(n_2844),
.Y(n_3213)
);

OR2x2_ASAP7_75t_L g3214 ( 
.A(n_3024),
.B(n_2900),
.Y(n_3214)
);

BUFx3_ASAP7_75t_L g3215 ( 
.A(n_3011),
.Y(n_3215)
);

INVx1_ASAP7_75t_L g3216 ( 
.A(n_3006),
.Y(n_3216)
);

OR2x2_ASAP7_75t_L g3217 ( 
.A(n_2989),
.B(n_2902),
.Y(n_3217)
);

INVx2_ASAP7_75t_L g3218 ( 
.A(n_2975),
.Y(n_3218)
);

AOI22xp5_ASAP7_75t_L g3219 ( 
.A1(n_3064),
.A2(n_2960),
.B1(n_2774),
.B2(n_2828),
.Y(n_3219)
);

INVx1_ASAP7_75t_L g3220 ( 
.A(n_3019),
.Y(n_3220)
);

NOR2xp33_ASAP7_75t_L g3221 ( 
.A(n_3017),
.B(n_2666),
.Y(n_3221)
);

NAND2xp5_ASAP7_75t_L g3222 ( 
.A(n_2992),
.B(n_2855),
.Y(n_3222)
);

INVx1_ASAP7_75t_L g3223 ( 
.A(n_3020),
.Y(n_3223)
);

AOI22xp33_ASAP7_75t_L g3224 ( 
.A1(n_3005),
.A2(n_2595),
.B1(n_2524),
.B2(n_2337),
.Y(n_3224)
);

NAND2xp5_ASAP7_75t_L g3225 ( 
.A(n_2998),
.B(n_2859),
.Y(n_3225)
);

INVx2_ASAP7_75t_L g3226 ( 
.A(n_3000),
.Y(n_3226)
);

HB1xp67_ASAP7_75t_L g3227 ( 
.A(n_3001),
.Y(n_3227)
);

BUFx12f_ASAP7_75t_L g3228 ( 
.A(n_3044),
.Y(n_3228)
);

CKINVDCx11_ASAP7_75t_R g3229 ( 
.A(n_2996),
.Y(n_3229)
);

CKINVDCx5p33_ASAP7_75t_R g3230 ( 
.A(n_3168),
.Y(n_3230)
);

NAND2xp5_ASAP7_75t_L g3231 ( 
.A(n_2968),
.B(n_2907),
.Y(n_3231)
);

NAND2xp5_ASAP7_75t_L g3232 ( 
.A(n_2968),
.B(n_2910),
.Y(n_3232)
);

BUFx6f_ASAP7_75t_L g3233 ( 
.A(n_3044),
.Y(n_3233)
);

INVx2_ASAP7_75t_L g3234 ( 
.A(n_3023),
.Y(n_3234)
);

INVx2_ASAP7_75t_SL g3235 ( 
.A(n_2981),
.Y(n_3235)
);

AND2x2_ASAP7_75t_L g3236 ( 
.A(n_3106),
.B(n_2940),
.Y(n_3236)
);

INVx1_ASAP7_75t_L g3237 ( 
.A(n_3032),
.Y(n_3237)
);

INVx1_ASAP7_75t_L g3238 ( 
.A(n_3055),
.Y(n_3238)
);

NAND2xp5_ASAP7_75t_L g3239 ( 
.A(n_3038),
.B(n_2911),
.Y(n_3239)
);

INVx1_ASAP7_75t_L g3240 ( 
.A(n_3058),
.Y(n_3240)
);

INVx1_ASAP7_75t_L g3241 ( 
.A(n_3075),
.Y(n_3241)
);

O2A1O1Ixp33_ASAP7_75t_L g3242 ( 
.A1(n_3035),
.A2(n_2337),
.B(n_2548),
.C(n_2381),
.Y(n_3242)
);

INVxp67_ASAP7_75t_L g3243 ( 
.A(n_3033),
.Y(n_3243)
);

NAND2xp5_ASAP7_75t_SL g3244 ( 
.A(n_2971),
.B(n_3071),
.Y(n_3244)
);

INVx2_ASAP7_75t_SL g3245 ( 
.A(n_3096),
.Y(n_3245)
);

INVx1_ASAP7_75t_L g3246 ( 
.A(n_3078),
.Y(n_3246)
);

NAND2xp5_ASAP7_75t_L g3247 ( 
.A(n_3040),
.B(n_2916),
.Y(n_3247)
);

BUFx3_ASAP7_75t_L g3248 ( 
.A(n_3131),
.Y(n_3248)
);

NOR2xp33_ASAP7_75t_L g3249 ( 
.A(n_2990),
.B(n_2666),
.Y(n_3249)
);

BUFx4f_ASAP7_75t_L g3250 ( 
.A(n_3015),
.Y(n_3250)
);

NOR2xp33_ASAP7_75t_L g3251 ( 
.A(n_3185),
.B(n_2961),
.Y(n_3251)
);

INVx2_ASAP7_75t_L g3252 ( 
.A(n_3041),
.Y(n_3252)
);

INVx1_ASAP7_75t_L g3253 ( 
.A(n_3112),
.Y(n_3253)
);

AOI22xp33_ASAP7_75t_L g3254 ( 
.A1(n_3045),
.A2(n_2548),
.B1(n_2436),
.B2(n_2940),
.Y(n_3254)
);

NAND2xp5_ASAP7_75t_L g3255 ( 
.A(n_3027),
.B(n_2931),
.Y(n_3255)
);

INVx2_ASAP7_75t_L g3256 ( 
.A(n_3062),
.Y(n_3256)
);

INVx2_ASAP7_75t_L g3257 ( 
.A(n_3135),
.Y(n_3257)
);

INVx4_ASAP7_75t_L g3258 ( 
.A(n_3134),
.Y(n_3258)
);

AND3x1_ASAP7_75t_L g3259 ( 
.A(n_3115),
.B(n_2425),
.C(n_2935),
.Y(n_3259)
);

AND2x2_ASAP7_75t_L g3260 ( 
.A(n_3101),
.B(n_2953),
.Y(n_3260)
);

INVx1_ASAP7_75t_L g3261 ( 
.A(n_2969),
.Y(n_3261)
);

NAND2xp5_ASAP7_75t_SL g3262 ( 
.A(n_3031),
.B(n_2488),
.Y(n_3262)
);

BUFx4f_ASAP7_75t_L g3263 ( 
.A(n_3015),
.Y(n_3263)
);

NAND2xp5_ASAP7_75t_L g3264 ( 
.A(n_2984),
.B(n_2769),
.Y(n_3264)
);

AND2x4_ASAP7_75t_L g3265 ( 
.A(n_3128),
.B(n_2766),
.Y(n_3265)
);

HB1xp67_ASAP7_75t_L g3266 ( 
.A(n_2974),
.Y(n_3266)
);

CKINVDCx5p33_ASAP7_75t_R g3267 ( 
.A(n_3130),
.Y(n_3267)
);

AOI22xp33_ASAP7_75t_L g3268 ( 
.A1(n_3068),
.A2(n_2436),
.B1(n_2959),
.B2(n_2956),
.Y(n_3268)
);

INVx2_ASAP7_75t_L g3269 ( 
.A(n_3143),
.Y(n_3269)
);

BUFx6f_ASAP7_75t_L g3270 ( 
.A(n_3131),
.Y(n_3270)
);

NAND2xp5_ASAP7_75t_L g3271 ( 
.A(n_3030),
.B(n_2938),
.Y(n_3271)
);

INVx5_ASAP7_75t_L g3272 ( 
.A(n_3134),
.Y(n_3272)
);

NAND2xp5_ASAP7_75t_SL g3273 ( 
.A(n_3125),
.B(n_2488),
.Y(n_3273)
);

INVx1_ASAP7_75t_L g3274 ( 
.A(n_2979),
.Y(n_3274)
);

AND2x4_ASAP7_75t_L g3275 ( 
.A(n_2987),
.B(n_2776),
.Y(n_3275)
);

INVx1_ASAP7_75t_L g3276 ( 
.A(n_3105),
.Y(n_3276)
);

BUFx6f_ASAP7_75t_L g3277 ( 
.A(n_3131),
.Y(n_3277)
);

INVxp67_ASAP7_75t_SL g3278 ( 
.A(n_3036),
.Y(n_3278)
);

INVx3_ASAP7_75t_L g3279 ( 
.A(n_3015),
.Y(n_3279)
);

INVx1_ASAP7_75t_L g3280 ( 
.A(n_3083),
.Y(n_3280)
);

NAND2xp5_ASAP7_75t_L g3281 ( 
.A(n_2980),
.B(n_3003),
.Y(n_3281)
);

INVx2_ASAP7_75t_L g3282 ( 
.A(n_3148),
.Y(n_3282)
);

INVx2_ASAP7_75t_SL g3283 ( 
.A(n_3108),
.Y(n_3283)
);

INVx1_ASAP7_75t_L g3284 ( 
.A(n_2983),
.Y(n_3284)
);

A2O1A1Ixp33_ASAP7_75t_L g3285 ( 
.A1(n_3057),
.A2(n_2505),
.B(n_2525),
.C(n_2824),
.Y(n_3285)
);

BUFx12f_ASAP7_75t_L g3286 ( 
.A(n_3113),
.Y(n_3286)
);

AND2x6_ASAP7_75t_L g3287 ( 
.A(n_3124),
.B(n_2805),
.Y(n_3287)
);

NAND2xp5_ASAP7_75t_SL g3288 ( 
.A(n_3092),
.B(n_2488),
.Y(n_3288)
);

INVxp67_ASAP7_75t_L g3289 ( 
.A(n_3046),
.Y(n_3289)
);

BUFx6f_ASAP7_75t_L g3290 ( 
.A(n_3134),
.Y(n_3290)
);

BUFx6f_ASAP7_75t_L g3291 ( 
.A(n_3134),
.Y(n_3291)
);

OR2x6_ASAP7_75t_L g3292 ( 
.A(n_3176),
.B(n_2843),
.Y(n_3292)
);

BUFx2_ASAP7_75t_L g3293 ( 
.A(n_3004),
.Y(n_3293)
);

AOI211xp5_ASAP7_75t_L g3294 ( 
.A1(n_3121),
.A2(n_2382),
.B(n_2944),
.C(n_2943),
.Y(n_3294)
);

NAND2xp5_ASAP7_75t_L g3295 ( 
.A(n_2980),
.B(n_2951),
.Y(n_3295)
);

INVx1_ASAP7_75t_L g3296 ( 
.A(n_3126),
.Y(n_3296)
);

INVx2_ASAP7_75t_L g3297 ( 
.A(n_3152),
.Y(n_3297)
);

INVx1_ASAP7_75t_L g3298 ( 
.A(n_3129),
.Y(n_3298)
);

INVx2_ASAP7_75t_L g3299 ( 
.A(n_3161),
.Y(n_3299)
);

INVx2_ASAP7_75t_L g3300 ( 
.A(n_3163),
.Y(n_3300)
);

AND2x4_ASAP7_75t_L g3301 ( 
.A(n_2987),
.B(n_2776),
.Y(n_3301)
);

INVx2_ASAP7_75t_SL g3302 ( 
.A(n_2997),
.Y(n_3302)
);

NOR2xp33_ASAP7_75t_L g3303 ( 
.A(n_3085),
.B(n_2639),
.Y(n_3303)
);

INVx1_ASAP7_75t_L g3304 ( 
.A(n_3132),
.Y(n_3304)
);

AND2x4_ASAP7_75t_L g3305 ( 
.A(n_3182),
.B(n_2468),
.Y(n_3305)
);

AND2x4_ASAP7_75t_L g3306 ( 
.A(n_3182),
.B(n_2469),
.Y(n_3306)
);

INVx2_ASAP7_75t_L g3307 ( 
.A(n_3164),
.Y(n_3307)
);

BUFx2_ASAP7_75t_L g3308 ( 
.A(n_3039),
.Y(n_3308)
);

INVx1_ASAP7_75t_L g3309 ( 
.A(n_3137),
.Y(n_3309)
);

INVx1_ASAP7_75t_L g3310 ( 
.A(n_3139),
.Y(n_3310)
);

INVx2_ASAP7_75t_L g3311 ( 
.A(n_3066),
.Y(n_3311)
);

BUFx4f_ASAP7_75t_L g3312 ( 
.A(n_3133),
.Y(n_3312)
);

NAND2xp5_ASAP7_75t_L g3313 ( 
.A(n_3007),
.B(n_2803),
.Y(n_3313)
);

INVx3_ASAP7_75t_L g3314 ( 
.A(n_3133),
.Y(n_3314)
);

INVx3_ASAP7_75t_L g3315 ( 
.A(n_3133),
.Y(n_3315)
);

BUFx8_ASAP7_75t_SL g3316 ( 
.A(n_3026),
.Y(n_3316)
);

BUFx6f_ASAP7_75t_L g3317 ( 
.A(n_3037),
.Y(n_3317)
);

INVx1_ASAP7_75t_L g3318 ( 
.A(n_3140),
.Y(n_3318)
);

INVx1_ASAP7_75t_L g3319 ( 
.A(n_3141),
.Y(n_3319)
);

AOI22xp5_ASAP7_75t_L g3320 ( 
.A1(n_3119),
.A2(n_2814),
.B1(n_2899),
.B2(n_2436),
.Y(n_3320)
);

INVx1_ASAP7_75t_L g3321 ( 
.A(n_3150),
.Y(n_3321)
);

INVx5_ASAP7_75t_L g3322 ( 
.A(n_2976),
.Y(n_3322)
);

INVx3_ASAP7_75t_L g3323 ( 
.A(n_2977),
.Y(n_3323)
);

AOI22xp5_ASAP7_75t_L g3324 ( 
.A1(n_3120),
.A2(n_3072),
.B1(n_2978),
.B2(n_3136),
.Y(n_3324)
);

INVx2_ASAP7_75t_L g3325 ( 
.A(n_3095),
.Y(n_3325)
);

INVx4_ASAP7_75t_L g3326 ( 
.A(n_2977),
.Y(n_3326)
);

BUFx3_ASAP7_75t_L g3327 ( 
.A(n_3063),
.Y(n_3327)
);

INVx5_ASAP7_75t_L g3328 ( 
.A(n_2976),
.Y(n_3328)
);

BUFx3_ASAP7_75t_L g3329 ( 
.A(n_3167),
.Y(n_3329)
);

NAND2xp5_ASAP7_75t_L g3330 ( 
.A(n_3022),
.B(n_2959),
.Y(n_3330)
);

INVx1_ASAP7_75t_L g3331 ( 
.A(n_3156),
.Y(n_3331)
);

OAI22xp5_ASAP7_75t_L g3332 ( 
.A1(n_3146),
.A2(n_2899),
.B1(n_2520),
.B2(n_2745),
.Y(n_3332)
);

NAND2xp5_ASAP7_75t_L g3333 ( 
.A(n_3025),
.B(n_2811),
.Y(n_3333)
);

AOI22xp5_ASAP7_75t_L g3334 ( 
.A1(n_3138),
.A2(n_2566),
.B1(n_2570),
.B2(n_2614),
.Y(n_3334)
);

INVx3_ASAP7_75t_L g3335 ( 
.A(n_2995),
.Y(n_3335)
);

INVx4_ASAP7_75t_L g3336 ( 
.A(n_2995),
.Y(n_3336)
);

BUFx6f_ASAP7_75t_L g3337 ( 
.A(n_3186),
.Y(n_3337)
);

INVx3_ASAP7_75t_L g3338 ( 
.A(n_2982),
.Y(n_3338)
);

INVx2_ASAP7_75t_L g3339 ( 
.A(n_3158),
.Y(n_3339)
);

INVx3_ASAP7_75t_L g3340 ( 
.A(n_2982),
.Y(n_3340)
);

INVx2_ASAP7_75t_L g3341 ( 
.A(n_3162),
.Y(n_3341)
);

AND2x6_ASAP7_75t_L g3342 ( 
.A(n_3061),
.B(n_2921),
.Y(n_3342)
);

INVx4_ASAP7_75t_L g3343 ( 
.A(n_2976),
.Y(n_3343)
);

AND2x2_ASAP7_75t_SL g3344 ( 
.A(n_3074),
.B(n_3172),
.Y(n_3344)
);

NOR2xp33_ASAP7_75t_SL g3345 ( 
.A(n_3014),
.B(n_2412),
.Y(n_3345)
);

INVx1_ASAP7_75t_L g3346 ( 
.A(n_3171),
.Y(n_3346)
);

INVx1_ASAP7_75t_L g3347 ( 
.A(n_3173),
.Y(n_3347)
);

AND2x4_ASAP7_75t_L g3348 ( 
.A(n_3081),
.B(n_2469),
.Y(n_3348)
);

CKINVDCx6p67_ASAP7_75t_R g3349 ( 
.A(n_3117),
.Y(n_3349)
);

NAND2xp5_ASAP7_75t_L g3350 ( 
.A(n_3049),
.B(n_2823),
.Y(n_3350)
);

INVx1_ASAP7_75t_L g3351 ( 
.A(n_3178),
.Y(n_3351)
);

INVx1_ASAP7_75t_L g3352 ( 
.A(n_3179),
.Y(n_3352)
);

NAND2xp5_ASAP7_75t_L g3353 ( 
.A(n_3086),
.B(n_3088),
.Y(n_3353)
);

OR2x6_ASAP7_75t_L g3354 ( 
.A(n_3175),
.B(n_2843),
.Y(n_3354)
);

INVx4_ASAP7_75t_L g3355 ( 
.A(n_3052),
.Y(n_3355)
);

A2O1A1Ixp33_ASAP7_75t_L g3356 ( 
.A1(n_3067),
.A2(n_2824),
.B(n_2815),
.C(n_2785),
.Y(n_3356)
);

INVx3_ASAP7_75t_L g3357 ( 
.A(n_3052),
.Y(n_3357)
);

INVx1_ASAP7_75t_L g3358 ( 
.A(n_3180),
.Y(n_3358)
);

AOI22xp5_ASAP7_75t_L g3359 ( 
.A1(n_3138),
.A2(n_3073),
.B1(n_3076),
.B2(n_3065),
.Y(n_3359)
);

INVx1_ASAP7_75t_L g3360 ( 
.A(n_3181),
.Y(n_3360)
);

AOI22xp5_ASAP7_75t_L g3361 ( 
.A1(n_3165),
.A2(n_2566),
.B1(n_2570),
.B2(n_2614),
.Y(n_3361)
);

INVx2_ASAP7_75t_L g3362 ( 
.A(n_3184),
.Y(n_3362)
);

INVx1_ASAP7_75t_L g3363 ( 
.A(n_3110),
.Y(n_3363)
);

INVx2_ASAP7_75t_L g3364 ( 
.A(n_3110),
.Y(n_3364)
);

HB1xp67_ASAP7_75t_L g3365 ( 
.A(n_3165),
.Y(n_3365)
);

INVx1_ASAP7_75t_L g3366 ( 
.A(n_3114),
.Y(n_3366)
);

AOI21xp5_ASAP7_75t_L g3367 ( 
.A1(n_3018),
.A2(n_2345),
.B(n_2553),
.Y(n_3367)
);

CKINVDCx16_ASAP7_75t_R g3368 ( 
.A(n_2991),
.Y(n_3368)
);

NOR2xp33_ASAP7_75t_SL g3369 ( 
.A(n_3014),
.B(n_2412),
.Y(n_3369)
);

NAND2xp5_ASAP7_75t_L g3370 ( 
.A(n_3069),
.B(n_2835),
.Y(n_3370)
);

INVxp67_ASAP7_75t_L g3371 ( 
.A(n_3080),
.Y(n_3371)
);

INVx2_ASAP7_75t_L g3372 ( 
.A(n_3114),
.Y(n_3372)
);

BUFx3_ASAP7_75t_L g3373 ( 
.A(n_3079),
.Y(n_3373)
);

INVx2_ASAP7_75t_L g3374 ( 
.A(n_3093),
.Y(n_3374)
);

NOR2xp33_ASAP7_75t_L g3375 ( 
.A(n_2966),
.B(n_2639),
.Y(n_3375)
);

INVx8_ASAP7_75t_L g3376 ( 
.A(n_3103),
.Y(n_3376)
);

AOI22xp5_ASAP7_75t_L g3377 ( 
.A1(n_2973),
.A2(n_2566),
.B1(n_2570),
.B2(n_2614),
.Y(n_3377)
);

INVx1_ASAP7_75t_L g3378 ( 
.A(n_3034),
.Y(n_3378)
);

OR2x6_ASAP7_75t_L g3379 ( 
.A(n_3036),
.B(n_2428),
.Y(n_3379)
);

HB1xp67_ASAP7_75t_L g3380 ( 
.A(n_3029),
.Y(n_3380)
);

INVx3_ASAP7_75t_L g3381 ( 
.A(n_3103),
.Y(n_3381)
);

INVx1_ASAP7_75t_L g3382 ( 
.A(n_3093),
.Y(n_3382)
);

AND2x4_ASAP7_75t_L g3383 ( 
.A(n_2970),
.B(n_2469),
.Y(n_3383)
);

NAND2xp5_ASAP7_75t_L g3384 ( 
.A(n_3043),
.B(n_2840),
.Y(n_3384)
);

AND2x4_ASAP7_75t_L g3385 ( 
.A(n_3070),
.B(n_2470),
.Y(n_3385)
);

OR2x6_ASAP7_75t_L g3386 ( 
.A(n_3013),
.B(n_2428),
.Y(n_3386)
);

INVx1_ASAP7_75t_L g3387 ( 
.A(n_3094),
.Y(n_3387)
);

BUFx3_ASAP7_75t_L g3388 ( 
.A(n_3155),
.Y(n_3388)
);

NAND2xp5_ASAP7_75t_L g3389 ( 
.A(n_3089),
.B(n_2846),
.Y(n_3389)
);

INVx1_ASAP7_75t_L g3390 ( 
.A(n_3094),
.Y(n_3390)
);

NAND2xp5_ASAP7_75t_L g3391 ( 
.A(n_2984),
.B(n_2852),
.Y(n_3391)
);

AND2x6_ASAP7_75t_SL g3392 ( 
.A(n_3127),
.B(n_2607),
.Y(n_3392)
);

INVx2_ASAP7_75t_L g3393 ( 
.A(n_3097),
.Y(n_3393)
);

INVxp67_ASAP7_75t_L g3394 ( 
.A(n_3056),
.Y(n_3394)
);

AND3x1_ASAP7_75t_SL g3395 ( 
.A(n_3082),
.B(n_76),
.C(n_68),
.Y(n_3395)
);

BUFx2_ASAP7_75t_L g3396 ( 
.A(n_3122),
.Y(n_3396)
);

AOI21xp5_ASAP7_75t_L g3397 ( 
.A1(n_3285),
.A2(n_3042),
.B(n_3028),
.Y(n_3397)
);

INVx1_ASAP7_75t_L g3398 ( 
.A(n_3188),
.Y(n_3398)
);

AOI22xp5_ASAP7_75t_L g3399 ( 
.A1(n_3202),
.A2(n_2607),
.B1(n_3053),
.B2(n_3170),
.Y(n_3399)
);

AOI21xp5_ASAP7_75t_L g3400 ( 
.A1(n_3367),
.A2(n_3174),
.B(n_3169),
.Y(n_3400)
);

AOI21xp5_ASAP7_75t_L g3401 ( 
.A1(n_3345),
.A2(n_3174),
.B(n_3169),
.Y(n_3401)
);

INVx1_ASAP7_75t_L g3402 ( 
.A(n_3195),
.Y(n_3402)
);

AOI21xp5_ASAP7_75t_L g3403 ( 
.A1(n_3345),
.A2(n_2785),
.B(n_2345),
.Y(n_3403)
);

NAND2xp5_ASAP7_75t_L g3404 ( 
.A(n_3378),
.B(n_3118),
.Y(n_3404)
);

AOI21xp5_ASAP7_75t_L g3405 ( 
.A1(n_3369),
.A2(n_2553),
.B(n_2502),
.Y(n_3405)
);

NOR2xp33_ASAP7_75t_L g3406 ( 
.A(n_3244),
.B(n_3059),
.Y(n_3406)
);

OAI21xp33_ASAP7_75t_L g3407 ( 
.A1(n_3198),
.A2(n_3159),
.B(n_3054),
.Y(n_3407)
);

AOI21xp5_ASAP7_75t_L g3408 ( 
.A1(n_3369),
.A2(n_2496),
.B(n_3090),
.Y(n_3408)
);

AOI21xp5_ASAP7_75t_L g3409 ( 
.A1(n_3278),
.A2(n_3090),
.B(n_2836),
.Y(n_3409)
);

NAND2xp5_ASAP7_75t_SL g3410 ( 
.A(n_3221),
.B(n_3107),
.Y(n_3410)
);

AOI21xp5_ASAP7_75t_L g3411 ( 
.A1(n_3356),
.A2(n_2839),
.B(n_2812),
.Y(n_3411)
);

OA22x2_ASAP7_75t_L g3412 ( 
.A1(n_3219),
.A2(n_3144),
.B1(n_2607),
.B2(n_3077),
.Y(n_3412)
);

AOI21xp5_ASAP7_75t_L g3413 ( 
.A1(n_3334),
.A2(n_2504),
.B(n_2921),
.Y(n_3413)
);

BUFx8_ASAP7_75t_SL g3414 ( 
.A(n_3209),
.Y(n_3414)
);

NOR2xp33_ASAP7_75t_L g3415 ( 
.A(n_3251),
.B(n_3249),
.Y(n_3415)
);

AOI22xp5_ASAP7_75t_L g3416 ( 
.A1(n_3211),
.A2(n_2607),
.B1(n_3012),
.B2(n_3048),
.Y(n_3416)
);

O2A1O1Ixp33_ASAP7_75t_SL g3417 ( 
.A1(n_3187),
.A2(n_3147),
.B(n_3111),
.C(n_3091),
.Y(n_3417)
);

AOI21xp5_ASAP7_75t_L g3418 ( 
.A1(n_3334),
.A2(n_2954),
.B(n_2929),
.Y(n_3418)
);

AOI21xp5_ASAP7_75t_L g3419 ( 
.A1(n_3264),
.A2(n_2954),
.B(n_2929),
.Y(n_3419)
);

OAI21xp5_ASAP7_75t_L g3420 ( 
.A1(n_3242),
.A2(n_2500),
.B(n_3047),
.Y(n_3420)
);

AOI21xp5_ASAP7_75t_L g3421 ( 
.A1(n_3264),
.A2(n_2790),
.B(n_2767),
.Y(n_3421)
);

INVx2_ASAP7_75t_L g3422 ( 
.A(n_3257),
.Y(n_3422)
);

OAI21xp33_ASAP7_75t_SL g3423 ( 
.A1(n_3361),
.A2(n_3091),
.B(n_2669),
.Y(n_3423)
);

OR2x2_ASAP7_75t_L g3424 ( 
.A(n_3396),
.B(n_3149),
.Y(n_3424)
);

NAND2xp5_ASAP7_75t_L g3425 ( 
.A(n_3227),
.B(n_3144),
.Y(n_3425)
);

INVx4_ASAP7_75t_L g3426 ( 
.A(n_3272),
.Y(n_3426)
);

OAI22xp5_ASAP7_75t_L g3427 ( 
.A1(n_3198),
.A2(n_3142),
.B1(n_3157),
.B2(n_3151),
.Y(n_3427)
);

NAND2xp33_ASAP7_75t_L g3428 ( 
.A(n_3267),
.B(n_2932),
.Y(n_3428)
);

AND2x2_ASAP7_75t_L g3429 ( 
.A(n_3208),
.B(n_3160),
.Y(n_3429)
);

INVx2_ASAP7_75t_L g3430 ( 
.A(n_3269),
.Y(n_3430)
);

HB1xp67_ASAP7_75t_L g3431 ( 
.A(n_3189),
.Y(n_3431)
);

BUFx6f_ASAP7_75t_L g3432 ( 
.A(n_3215),
.Y(n_3432)
);

OR2x6_ASAP7_75t_L g3433 ( 
.A(n_3292),
.B(n_2909),
.Y(n_3433)
);

NOR2x1_ASAP7_75t_L g3434 ( 
.A(n_3388),
.B(n_2917),
.Y(n_3434)
);

NAND3xp33_ASAP7_75t_L g3435 ( 
.A(n_3194),
.B(n_3104),
.C(n_2398),
.Y(n_3435)
);

NAND2xp5_ASAP7_75t_L g3436 ( 
.A(n_3281),
.B(n_3097),
.Y(n_3436)
);

AOI21xp5_ASAP7_75t_L g3437 ( 
.A1(n_3361),
.A2(n_2767),
.B(n_2669),
.Y(n_3437)
);

NAND3xp33_ASAP7_75t_SL g3438 ( 
.A(n_3212),
.B(n_3294),
.C(n_3187),
.Y(n_3438)
);

AOI21xp5_ASAP7_75t_L g3439 ( 
.A1(n_3377),
.A2(n_2809),
.B(n_2520),
.Y(n_3439)
);

NAND2xp5_ASAP7_75t_L g3440 ( 
.A(n_3330),
.B(n_3098),
.Y(n_3440)
);

O2A1O1Ixp33_ASAP7_75t_L g3441 ( 
.A1(n_3332),
.A2(n_3153),
.B(n_3166),
.C(n_3145),
.Y(n_3441)
);

INVx2_ASAP7_75t_SL g3442 ( 
.A(n_3286),
.Y(n_3442)
);

AOI22x1_ASAP7_75t_L g3443 ( 
.A1(n_3293),
.A2(n_2470),
.B1(n_2579),
.B2(n_2847),
.Y(n_3443)
);

NAND2xp5_ASAP7_75t_L g3444 ( 
.A(n_3353),
.B(n_3098),
.Y(n_3444)
);

NOR2xp33_ASAP7_75t_L g3445 ( 
.A(n_3373),
.B(n_2639),
.Y(n_3445)
);

AOI21xp5_ASAP7_75t_L g3446 ( 
.A1(n_3377),
.A2(n_2520),
.B(n_3145),
.Y(n_3446)
);

NAND2xp5_ASAP7_75t_SL g3447 ( 
.A(n_3213),
.B(n_2520),
.Y(n_3447)
);

AOI22xp5_ASAP7_75t_L g3448 ( 
.A1(n_3303),
.A2(n_2476),
.B1(n_3153),
.B2(n_2570),
.Y(n_3448)
);

O2A1O1Ixp33_ASAP7_75t_L g3449 ( 
.A1(n_3332),
.A2(n_3166),
.B(n_3102),
.C(n_3100),
.Y(n_3449)
);

OAI22xp5_ASAP7_75t_SL g3450 ( 
.A1(n_3368),
.A2(n_2962),
.B1(n_2950),
.B2(n_2948),
.Y(n_3450)
);

NAND3xp33_ASAP7_75t_L g3451 ( 
.A(n_3294),
.B(n_3102),
.C(n_3100),
.Y(n_3451)
);

INVx1_ASAP7_75t_SL g3452 ( 
.A(n_3308),
.Y(n_3452)
);

NAND2xp5_ASAP7_75t_L g3453 ( 
.A(n_3289),
.B(n_2854),
.Y(n_3453)
);

OAI21x1_ASAP7_75t_L g3454 ( 
.A1(n_3262),
.A2(n_2426),
.B(n_2421),
.Y(n_3454)
);

AOI22xp33_ASAP7_75t_L g3455 ( 
.A1(n_3344),
.A2(n_2476),
.B1(n_2788),
.B2(n_2779),
.Y(n_3455)
);

AOI22xp33_ASAP7_75t_SL g3456 ( 
.A1(n_3287),
.A2(n_2579),
.B1(n_2476),
.B2(n_2570),
.Y(n_3456)
);

OAI22xp5_ASAP7_75t_L g3457 ( 
.A1(n_3219),
.A2(n_2470),
.B1(n_2868),
.B2(n_2367),
.Y(n_3457)
);

NAND2xp5_ASAP7_75t_SL g3458 ( 
.A(n_3259),
.B(n_3239),
.Y(n_3458)
);

INVx1_ASAP7_75t_L g3459 ( 
.A(n_3196),
.Y(n_3459)
);

INVxp67_ASAP7_75t_L g3460 ( 
.A(n_3204),
.Y(n_3460)
);

OAI22x1_ASAP7_75t_L g3461 ( 
.A1(n_3320),
.A2(n_3177),
.B1(n_2749),
.B2(n_2729),
.Y(n_3461)
);

AOI22xp33_ASAP7_75t_L g3462 ( 
.A1(n_3229),
.A2(n_2476),
.B1(n_2788),
.B2(n_2779),
.Y(n_3462)
);

NAND2xp5_ASAP7_75t_L g3463 ( 
.A(n_3247),
.B(n_2861),
.Y(n_3463)
);

INVx2_ASAP7_75t_SL g3464 ( 
.A(n_3235),
.Y(n_3464)
);

INVx3_ASAP7_75t_L g3465 ( 
.A(n_3290),
.Y(n_3465)
);

AND2x2_ASAP7_75t_SL g3466 ( 
.A(n_3320),
.B(n_2932),
.Y(n_3466)
);

INVx2_ASAP7_75t_L g3467 ( 
.A(n_3282),
.Y(n_3467)
);

OA22x2_ASAP7_75t_L g3468 ( 
.A1(n_3324),
.A2(n_2872),
.B1(n_2869),
.B2(n_2847),
.Y(n_3468)
);

NOR2xp33_ASAP7_75t_R g3469 ( 
.A(n_3230),
.B(n_3190),
.Y(n_3469)
);

AOI221xp5_ASAP7_75t_L g3470 ( 
.A1(n_3324),
.A2(n_3394),
.B1(n_3243),
.B2(n_2579),
.C(n_3371),
.Y(n_3470)
);

OAI21xp33_ASAP7_75t_L g3471 ( 
.A1(n_3359),
.A2(n_2579),
.B(n_2769),
.Y(n_3471)
);

AOI21xp5_ASAP7_75t_L g3472 ( 
.A1(n_3322),
.A2(n_3328),
.B(n_3295),
.Y(n_3472)
);

AND2x2_ASAP7_75t_L g3473 ( 
.A(n_3260),
.B(n_2905),
.Y(n_3473)
);

A2O1A1Ixp33_ASAP7_75t_SL g3474 ( 
.A1(n_3375),
.A2(n_3177),
.B(n_2864),
.C(n_2871),
.Y(n_3474)
);

AOI21xp5_ASAP7_75t_L g3475 ( 
.A1(n_3322),
.A2(n_3328),
.B(n_3232),
.Y(n_3475)
);

NAND2xp5_ASAP7_75t_SL g3476 ( 
.A(n_3259),
.B(n_2422),
.Y(n_3476)
);

A2O1A1Ixp33_ASAP7_75t_SL g3477 ( 
.A1(n_3206),
.A2(n_2882),
.B(n_2888),
.C(n_2862),
.Y(n_3477)
);

AO21x1_ASAP7_75t_L g3478 ( 
.A1(n_3210),
.A2(n_2914),
.B(n_2747),
.Y(n_3478)
);

AOI22xp5_ASAP7_75t_L g3479 ( 
.A1(n_3236),
.A2(n_3287),
.B1(n_3288),
.B2(n_3200),
.Y(n_3479)
);

INVx1_ASAP7_75t_L g3480 ( 
.A(n_3197),
.Y(n_3480)
);

NOR2xp33_ASAP7_75t_L g3481 ( 
.A(n_3205),
.B(n_2932),
.Y(n_3481)
);

O2A1O1Ixp33_ASAP7_75t_L g3482 ( 
.A1(n_3273),
.A2(n_2747),
.B(n_2623),
.C(n_2626),
.Y(n_3482)
);

INVx1_ASAP7_75t_L g3483 ( 
.A(n_3216),
.Y(n_3483)
);

AO32x1_ASAP7_75t_L g3484 ( 
.A1(n_3363),
.A2(n_2778),
.A3(n_2649),
.B1(n_2880),
.B2(n_2454),
.Y(n_3484)
);

BUFx6f_ASAP7_75t_L g3485 ( 
.A(n_3290),
.Y(n_3485)
);

AOI21xp5_ASAP7_75t_L g3486 ( 
.A1(n_3322),
.A2(n_2880),
.B(n_2562),
.Y(n_3486)
);

OAI22xp5_ASAP7_75t_L g3487 ( 
.A1(n_3268),
.A2(n_2374),
.B1(n_2377),
.B2(n_2375),
.Y(n_3487)
);

AOI21xp5_ASAP7_75t_L g3488 ( 
.A1(n_3328),
.A2(n_3231),
.B(n_3391),
.Y(n_3488)
);

BUFx4f_ASAP7_75t_L g3489 ( 
.A(n_3290),
.Y(n_3489)
);

AND2x4_ASAP7_75t_L g3490 ( 
.A(n_3203),
.B(n_2683),
.Y(n_3490)
);

AND2x4_ASAP7_75t_L g3491 ( 
.A(n_3203),
.B(n_2683),
.Y(n_3491)
);

AOI21xp5_ASAP7_75t_L g3492 ( 
.A1(n_3354),
.A2(n_2999),
.B(n_2359),
.Y(n_3492)
);

BUFx12f_ASAP7_75t_L g3493 ( 
.A(n_3228),
.Y(n_3493)
);

BUFx2_ASAP7_75t_L g3494 ( 
.A(n_3365),
.Y(n_3494)
);

INVx1_ASAP7_75t_L g3495 ( 
.A(n_3220),
.Y(n_3495)
);

OR2x2_ASAP7_75t_L g3496 ( 
.A(n_3201),
.B(n_2914),
.Y(n_3496)
);

AO21x2_ASAP7_75t_L g3497 ( 
.A1(n_3359),
.A2(n_2631),
.B(n_2616),
.Y(n_3497)
);

OAI22xp5_ASAP7_75t_L g3498 ( 
.A1(n_3254),
.A2(n_2796),
.B1(n_2392),
.B2(n_2449),
.Y(n_3498)
);

INVx2_ASAP7_75t_L g3499 ( 
.A(n_3297),
.Y(n_3499)
);

O2A1O1Ixp33_ASAP7_75t_L g3500 ( 
.A1(n_3380),
.A2(n_2452),
.B(n_2406),
.C(n_2872),
.Y(n_3500)
);

BUFx2_ASAP7_75t_L g3501 ( 
.A(n_3248),
.Y(n_3501)
);

HB1xp67_ASAP7_75t_L g3502 ( 
.A(n_3261),
.Y(n_3502)
);

AOI21xp5_ASAP7_75t_L g3503 ( 
.A1(n_3354),
.A2(n_2358),
.B(n_2380),
.Y(n_3503)
);

INVx2_ASAP7_75t_L g3504 ( 
.A(n_3299),
.Y(n_3504)
);

OR2x2_ASAP7_75t_L g3505 ( 
.A(n_3214),
.B(n_2860),
.Y(n_3505)
);

AOI21xp5_ASAP7_75t_L g3506 ( 
.A1(n_3354),
.A2(n_2414),
.B(n_2685),
.Y(n_3506)
);

CKINVDCx5p33_ASAP7_75t_R g3507 ( 
.A(n_3316),
.Y(n_3507)
);

AOI21xp5_ASAP7_75t_L g3508 ( 
.A1(n_3222),
.A2(n_2414),
.B(n_2685),
.Y(n_3508)
);

NAND2xp5_ASAP7_75t_L g3509 ( 
.A(n_3313),
.B(n_2908),
.Y(n_3509)
);

NAND2xp5_ASAP7_75t_SL g3510 ( 
.A(n_3217),
.B(n_2422),
.Y(n_3510)
);

CKINVDCx10_ASAP7_75t_R g3511 ( 
.A(n_3368),
.Y(n_3511)
);

O2A1O1Ixp33_ASAP7_75t_L g3512 ( 
.A1(n_3266),
.A2(n_2668),
.B(n_2667),
.C(n_2523),
.Y(n_3512)
);

INVx2_ASAP7_75t_L g3513 ( 
.A(n_3300),
.Y(n_3513)
);

NOR2xp33_ASAP7_75t_L g3514 ( 
.A(n_3275),
.B(n_2936),
.Y(n_3514)
);

INVx3_ASAP7_75t_L g3515 ( 
.A(n_3291),
.Y(n_3515)
);

NAND3xp33_ASAP7_75t_L g3516 ( 
.A(n_3193),
.B(n_2749),
.C(n_2729),
.Y(n_3516)
);

BUFx4f_ASAP7_75t_L g3517 ( 
.A(n_3291),
.Y(n_3517)
);

AO32x2_ASAP7_75t_L g3518 ( 
.A1(n_3392),
.A2(n_2778),
.A3(n_2884),
.B1(n_2920),
.B2(n_2869),
.Y(n_3518)
);

AOI21xp5_ASAP7_75t_L g3519 ( 
.A1(n_3225),
.A2(n_2414),
.B(n_2724),
.Y(n_3519)
);

NOR2xp33_ASAP7_75t_L g3520 ( 
.A(n_3275),
.B(n_2936),
.Y(n_3520)
);

NAND2x1p5_ASAP7_75t_L g3521 ( 
.A(n_3272),
.B(n_2373),
.Y(n_3521)
);

O2A1O1Ixp33_ASAP7_75t_SL g3522 ( 
.A1(n_3255),
.A2(n_3271),
.B(n_3276),
.C(n_3253),
.Y(n_3522)
);

OAI21xp33_ASAP7_75t_L g3523 ( 
.A1(n_3224),
.A2(n_2455),
.B(n_2660),
.Y(n_3523)
);

AOI21xp5_ASAP7_75t_L g3524 ( 
.A1(n_3192),
.A2(n_2724),
.B(n_2860),
.Y(n_3524)
);

NOR2x1_ASAP7_75t_L g3525 ( 
.A(n_3326),
.B(n_2434),
.Y(n_3525)
);

NOR2xp33_ASAP7_75t_L g3526 ( 
.A(n_3301),
.B(n_2936),
.Y(n_3526)
);

NAND2x1_ASAP7_75t_L g3527 ( 
.A(n_3343),
.B(n_2399),
.Y(n_3527)
);

AOI22xp33_ASAP7_75t_SL g3528 ( 
.A1(n_3287),
.A2(n_2476),
.B1(n_2570),
.B2(n_2566),
.Y(n_3528)
);

AND2x4_ASAP7_75t_L g3529 ( 
.A(n_3203),
.B(n_2683),
.Y(n_3529)
);

INVx2_ASAP7_75t_L g3530 ( 
.A(n_3307),
.Y(n_3530)
);

INVx5_ASAP7_75t_L g3531 ( 
.A(n_3272),
.Y(n_3531)
);

NAND2xp5_ASAP7_75t_L g3532 ( 
.A(n_3384),
.B(n_2925),
.Y(n_3532)
);

NOR2xp33_ASAP7_75t_L g3533 ( 
.A(n_3301),
.B(n_2948),
.Y(n_3533)
);

NAND2xp5_ASAP7_75t_L g3534 ( 
.A(n_3350),
.B(n_2937),
.Y(n_3534)
);

AOI21xp5_ASAP7_75t_L g3535 ( 
.A1(n_3192),
.A2(n_2550),
.B(n_2544),
.Y(n_3535)
);

NAND2xp5_ASAP7_75t_L g3536 ( 
.A(n_3364),
.B(n_2945),
.Y(n_3536)
);

NAND2xp5_ASAP7_75t_L g3537 ( 
.A(n_3372),
.B(n_2946),
.Y(n_3537)
);

NAND2xp33_ASAP7_75t_L g3538 ( 
.A(n_3342),
.B(n_2948),
.Y(n_3538)
);

AOI21xp5_ASAP7_75t_L g3539 ( 
.A1(n_3292),
.A2(n_2550),
.B(n_2544),
.Y(n_3539)
);

NOR2xp33_ASAP7_75t_L g3540 ( 
.A(n_3245),
.B(n_2950),
.Y(n_3540)
);

NAND2xp5_ASAP7_75t_L g3541 ( 
.A(n_3374),
.B(n_2722),
.Y(n_3541)
);

AOI221xp5_ASAP7_75t_L g3542 ( 
.A1(n_3274),
.A2(n_2615),
.B1(n_2796),
.B2(n_2834),
.C(n_2826),
.Y(n_3542)
);

NAND2xp5_ASAP7_75t_L g3543 ( 
.A(n_3393),
.B(n_2722),
.Y(n_3543)
);

NOR2x1p5_ASAP7_75t_SL g3544 ( 
.A(n_3366),
.B(n_2435),
.Y(n_3544)
);

NAND2xp33_ASAP7_75t_SL g3545 ( 
.A(n_3291),
.B(n_2950),
.Y(n_3545)
);

INVx2_ASAP7_75t_L g3546 ( 
.A(n_3191),
.Y(n_3546)
);

INVx4_ASAP7_75t_L g3547 ( 
.A(n_3258),
.Y(n_3547)
);

AOI21xp5_ASAP7_75t_L g3548 ( 
.A1(n_3292),
.A2(n_2858),
.B(n_2845),
.Y(n_3548)
);

O2A1O1Ixp33_ASAP7_75t_L g3549 ( 
.A1(n_3379),
.A2(n_2318),
.B(n_2810),
.C(n_2789),
.Y(n_3549)
);

OAI21xp5_ASAP7_75t_L g3550 ( 
.A1(n_3370),
.A2(n_2476),
.B(n_2826),
.Y(n_3550)
);

O2A1O1Ixp33_ASAP7_75t_L g3551 ( 
.A1(n_3379),
.A2(n_2318),
.B(n_2810),
.C(n_2789),
.Y(n_3551)
);

OAI22xp5_ASAP7_75t_SL g3552 ( 
.A1(n_3283),
.A2(n_2920),
.B1(n_2884),
.B2(n_2516),
.Y(n_3552)
);

O2A1O1Ixp33_ASAP7_75t_L g3553 ( 
.A1(n_3379),
.A2(n_2318),
.B(n_2816),
.C(n_2894),
.Y(n_3553)
);

AOI22xp33_ASAP7_75t_L g3554 ( 
.A1(n_3287),
.A2(n_2566),
.B1(n_2834),
.B2(n_2614),
.Y(n_3554)
);

AOI33xp33_ASAP7_75t_L g3555 ( 
.A1(n_3223),
.A2(n_92),
.A3(n_76),
.B1(n_100),
.B2(n_84),
.B3(n_68),
.Y(n_3555)
);

NAND2x1p5_ASAP7_75t_L g3556 ( 
.A(n_3250),
.B(n_2373),
.Y(n_3556)
);

NAND2xp5_ASAP7_75t_L g3557 ( 
.A(n_3382),
.B(n_2722),
.Y(n_3557)
);

NAND2xp5_ASAP7_75t_L g3558 ( 
.A(n_3387),
.B(n_2722),
.Y(n_3558)
);

AOI21xp5_ASAP7_75t_L g3559 ( 
.A1(n_3333),
.A2(n_2858),
.B(n_2845),
.Y(n_3559)
);

BUFx6f_ASAP7_75t_L g3560 ( 
.A(n_3233),
.Y(n_3560)
);

NAND2xp5_ASAP7_75t_L g3561 ( 
.A(n_3390),
.B(n_2800),
.Y(n_3561)
);

AOI21xp5_ASAP7_75t_L g3562 ( 
.A1(n_3343),
.A2(n_2876),
.B(n_2573),
.Y(n_3562)
);

INVx2_ASAP7_75t_L g3563 ( 
.A(n_3199),
.Y(n_3563)
);

NOR2xp33_ASAP7_75t_SL g3564 ( 
.A(n_3250),
.B(n_2444),
.Y(n_3564)
);

OAI22xp5_ASAP7_75t_SL g3565 ( 
.A1(n_3302),
.A2(n_3386),
.B1(n_3329),
.B2(n_3327),
.Y(n_3565)
);

NAND2xp5_ASAP7_75t_SL g3566 ( 
.A(n_3348),
.B(n_2444),
.Y(n_3566)
);

BUFx2_ASAP7_75t_L g3567 ( 
.A(n_3233),
.Y(n_3567)
);

NOR2xp33_ASAP7_75t_L g3568 ( 
.A(n_3348),
.B(n_2444),
.Y(n_3568)
);

OAI21x1_ASAP7_75t_L g3569 ( 
.A1(n_3339),
.A2(n_2426),
.B(n_2421),
.Y(n_3569)
);

NAND2xp5_ASAP7_75t_L g3570 ( 
.A(n_3389),
.B(n_2800),
.Y(n_3570)
);

OAI21xp33_ASAP7_75t_L g3571 ( 
.A1(n_3237),
.A2(n_2515),
.B(n_2816),
.Y(n_3571)
);

NAND2xp5_ASAP7_75t_L g3572 ( 
.A(n_3362),
.B(n_2800),
.Y(n_3572)
);

OAI21x1_ASAP7_75t_L g3573 ( 
.A1(n_3341),
.A2(n_2426),
.B(n_2421),
.Y(n_3573)
);

AOI22xp5_ASAP7_75t_L g3574 ( 
.A1(n_3200),
.A2(n_2566),
.B1(n_2614),
.B2(n_2440),
.Y(n_3574)
);

NAND2xp5_ASAP7_75t_SL g3575 ( 
.A(n_3265),
.B(n_2516),
.Y(n_3575)
);

NAND2xp5_ASAP7_75t_SL g3576 ( 
.A(n_3265),
.B(n_2516),
.Y(n_3576)
);

NAND2xp5_ASAP7_75t_SL g3577 ( 
.A(n_3305),
.B(n_2373),
.Y(n_3577)
);

NAND2xp5_ASAP7_75t_L g3578 ( 
.A(n_3218),
.B(n_3226),
.Y(n_3578)
);

AOI21xp5_ASAP7_75t_L g3579 ( 
.A1(n_3383),
.A2(n_2876),
.B(n_2573),
.Y(n_3579)
);

A2O1A1Ixp33_ASAP7_75t_L g3580 ( 
.A1(n_3263),
.A2(n_2894),
.B(n_2369),
.C(n_2346),
.Y(n_3580)
);

NAND2xp5_ASAP7_75t_L g3581 ( 
.A(n_3234),
.B(n_2800),
.Y(n_3581)
);

AOI22xp5_ASAP7_75t_L g3582 ( 
.A1(n_3395),
.A2(n_2614),
.B1(n_2440),
.B2(n_2399),
.Y(n_3582)
);

NAND2xp5_ASAP7_75t_SL g3583 ( 
.A(n_3305),
.B(n_2373),
.Y(n_3583)
);

NOR2xp33_ASAP7_75t_SL g3584 ( 
.A(n_3263),
.B(n_2895),
.Y(n_3584)
);

INVx1_ASAP7_75t_L g3585 ( 
.A(n_3238),
.Y(n_3585)
);

HB1xp67_ASAP7_75t_L g3586 ( 
.A(n_3240),
.Y(n_3586)
);

AOI21xp5_ASAP7_75t_L g3587 ( 
.A1(n_3383),
.A2(n_3386),
.B(n_3312),
.Y(n_3587)
);

AND2x2_ASAP7_75t_L g3588 ( 
.A(n_3252),
.B(n_2721),
.Y(n_3588)
);

CKINVDCx5p33_ASAP7_75t_R g3589 ( 
.A(n_3317),
.Y(n_3589)
);

INVx4_ASAP7_75t_L g3590 ( 
.A(n_3258),
.Y(n_3590)
);

INVx4_ASAP7_75t_L g3591 ( 
.A(n_3312),
.Y(n_3591)
);

NAND2xp5_ASAP7_75t_L g3592 ( 
.A(n_3256),
.B(n_2439),
.Y(n_3592)
);

BUFx6f_ASAP7_75t_L g3593 ( 
.A(n_3233),
.Y(n_3593)
);

AOI21xp5_ASAP7_75t_L g3594 ( 
.A1(n_3386),
.A2(n_2573),
.B(n_2710),
.Y(n_3594)
);

AOI21xp5_ASAP7_75t_L g3595 ( 
.A1(n_3306),
.A2(n_2453),
.B(n_2435),
.Y(n_3595)
);

AOI21xp5_ASAP7_75t_L g3596 ( 
.A1(n_3306),
.A2(n_3376),
.B(n_3355),
.Y(n_3596)
);

AOI21xp5_ASAP7_75t_L g3597 ( 
.A1(n_3376),
.A2(n_2454),
.B(n_2453),
.Y(n_3597)
);

AOI21xp5_ASAP7_75t_L g3598 ( 
.A1(n_3376),
.A2(n_2459),
.B(n_2443),
.Y(n_3598)
);

AOI21xp5_ASAP7_75t_L g3599 ( 
.A1(n_3355),
.A2(n_2459),
.B(n_2443),
.Y(n_3599)
);

BUFx3_ASAP7_75t_L g3600 ( 
.A(n_3317),
.Y(n_3600)
);

NAND2xp5_ASAP7_75t_L g3601 ( 
.A(n_3311),
.B(n_2439),
.Y(n_3601)
);

NAND2x1_ASAP7_75t_L g3602 ( 
.A(n_3207),
.B(n_2399),
.Y(n_3602)
);

NOR2xp33_ASAP7_75t_L g3603 ( 
.A(n_3349),
.B(n_2696),
.Y(n_3603)
);

NAND2xp5_ASAP7_75t_L g3604 ( 
.A(n_3325),
.B(n_2450),
.Y(n_3604)
);

A2O1A1Ixp33_ASAP7_75t_SL g3605 ( 
.A1(n_3323),
.A2(n_2542),
.B(n_2369),
.C(n_2346),
.Y(n_3605)
);

OAI21x1_ASAP7_75t_L g3606 ( 
.A1(n_3562),
.A2(n_3296),
.B(n_3284),
.Y(n_3606)
);

INVx1_ASAP7_75t_L g3607 ( 
.A(n_3586),
.Y(n_3607)
);

OR2x2_ASAP7_75t_L g3608 ( 
.A(n_3494),
.B(n_3241),
.Y(n_3608)
);

INVx1_ASAP7_75t_L g3609 ( 
.A(n_3502),
.Y(n_3609)
);

OAI21x1_ASAP7_75t_L g3610 ( 
.A1(n_3486),
.A2(n_3304),
.B(n_3298),
.Y(n_3610)
);

A2O1A1Ixp33_ASAP7_75t_L g3611 ( 
.A1(n_3397),
.A2(n_3246),
.B(n_3385),
.C(n_3314),
.Y(n_3611)
);

BUFx2_ASAP7_75t_L g3612 ( 
.A(n_3433),
.Y(n_3612)
);

AOI221x1_ASAP7_75t_L g3613 ( 
.A1(n_3438),
.A2(n_3310),
.B1(n_3319),
.B2(n_3318),
.C(n_3309),
.Y(n_3613)
);

AOI21xp5_ASAP7_75t_L g3614 ( 
.A1(n_3405),
.A2(n_3385),
.B(n_3331),
.Y(n_3614)
);

A2O1A1Ixp33_ASAP7_75t_L g3615 ( 
.A1(n_3415),
.A2(n_3314),
.B(n_3315),
.C(n_3279),
.Y(n_3615)
);

OAI21xp5_ASAP7_75t_L g3616 ( 
.A1(n_3408),
.A2(n_3207),
.B(n_3342),
.Y(n_3616)
);

INVx1_ASAP7_75t_L g3617 ( 
.A(n_3398),
.Y(n_3617)
);

AOI21xp5_ASAP7_75t_L g3618 ( 
.A1(n_3400),
.A2(n_3346),
.B(n_3321),
.Y(n_3618)
);

OAI21x1_ASAP7_75t_L g3619 ( 
.A1(n_3579),
.A2(n_3351),
.B(n_3347),
.Y(n_3619)
);

OAI21x1_ASAP7_75t_L g3620 ( 
.A1(n_3492),
.A2(n_3594),
.B(n_3446),
.Y(n_3620)
);

AOI21xp5_ASAP7_75t_L g3621 ( 
.A1(n_3401),
.A2(n_3358),
.B(n_3352),
.Y(n_3621)
);

INVx4_ASAP7_75t_L g3622 ( 
.A(n_3531),
.Y(n_3622)
);

NAND2xp5_ASAP7_75t_L g3623 ( 
.A(n_3431),
.B(n_3360),
.Y(n_3623)
);

OAI21x1_ASAP7_75t_L g3624 ( 
.A1(n_3419),
.A2(n_3280),
.B(n_3338),
.Y(n_3624)
);

NAND2xp5_ASAP7_75t_L g3625 ( 
.A(n_3460),
.B(n_3392),
.Y(n_3625)
);

OAI21x1_ASAP7_75t_L g3626 ( 
.A1(n_3454),
.A2(n_3340),
.B(n_3338),
.Y(n_3626)
);

NAND2xp5_ASAP7_75t_L g3627 ( 
.A(n_3440),
.B(n_3340),
.Y(n_3627)
);

BUFx6f_ASAP7_75t_L g3628 ( 
.A(n_3432),
.Y(n_3628)
);

INVx2_ASAP7_75t_L g3629 ( 
.A(n_3402),
.Y(n_3629)
);

OR2x6_ASAP7_75t_L g3630 ( 
.A(n_3433),
.B(n_3279),
.Y(n_3630)
);

INVx2_ASAP7_75t_L g3631 ( 
.A(n_3459),
.Y(n_3631)
);

NAND2xp5_ASAP7_75t_L g3632 ( 
.A(n_3424),
.B(n_3357),
.Y(n_3632)
);

AOI21xp5_ASAP7_75t_L g3633 ( 
.A1(n_3522),
.A2(n_3335),
.B(n_3323),
.Y(n_3633)
);

AOI21xp5_ASAP7_75t_L g3634 ( 
.A1(n_3497),
.A2(n_3335),
.B(n_2883),
.Y(n_3634)
);

BUFx2_ASAP7_75t_L g3635 ( 
.A(n_3434),
.Y(n_3635)
);

OR2x2_ASAP7_75t_L g3636 ( 
.A(n_3496),
.B(n_3357),
.Y(n_3636)
);

NAND3xp33_ASAP7_75t_L g3637 ( 
.A(n_3555),
.B(n_3381),
.C(n_3336),
.Y(n_3637)
);

NAND2xp5_ASAP7_75t_L g3638 ( 
.A(n_3436),
.B(n_3381),
.Y(n_3638)
);

NOR2x1_ASAP7_75t_SL g3639 ( 
.A(n_3458),
.B(n_3326),
.Y(n_3639)
);

NAND2xp5_ASAP7_75t_L g3640 ( 
.A(n_3444),
.B(n_3207),
.Y(n_3640)
);

OAI21x1_ASAP7_75t_L g3641 ( 
.A1(n_3539),
.A2(n_3315),
.B(n_2450),
.Y(n_3641)
);

NAND2x1p5_ASAP7_75t_L g3642 ( 
.A(n_3531),
.B(n_3336),
.Y(n_3642)
);

AOI21x1_ASAP7_75t_L g3643 ( 
.A1(n_3476),
.A2(n_2883),
.B(n_2875),
.Y(n_3643)
);

OAI21xp5_ASAP7_75t_L g3644 ( 
.A1(n_3435),
.A2(n_3207),
.B(n_3342),
.Y(n_3644)
);

OAI21x1_ASAP7_75t_SL g3645 ( 
.A1(n_3587),
.A2(n_2875),
.B(n_3342),
.Y(n_3645)
);

OAI21xp5_ASAP7_75t_L g3646 ( 
.A1(n_3488),
.A2(n_2440),
.B(n_2399),
.Y(n_3646)
);

INVx2_ASAP7_75t_L g3647 ( 
.A(n_3480),
.Y(n_3647)
);

HB1xp67_ASAP7_75t_L g3648 ( 
.A(n_3483),
.Y(n_3648)
);

AND2x4_ASAP7_75t_L g3649 ( 
.A(n_3495),
.B(n_3270),
.Y(n_3649)
);

AND2x2_ASAP7_75t_L g3650 ( 
.A(n_3429),
.B(n_3317),
.Y(n_3650)
);

INVx2_ASAP7_75t_L g3651 ( 
.A(n_3585),
.Y(n_3651)
);

OR2x2_ASAP7_75t_L g3652 ( 
.A(n_3425),
.B(n_3270),
.Y(n_3652)
);

OAI21xp5_ASAP7_75t_L g3653 ( 
.A1(n_3399),
.A2(n_2440),
.B(n_2399),
.Y(n_3653)
);

NAND2xp5_ASAP7_75t_L g3654 ( 
.A(n_3404),
.B(n_3270),
.Y(n_3654)
);

NOR2xp33_ASAP7_75t_L g3655 ( 
.A(n_3414),
.B(n_3337),
.Y(n_3655)
);

NAND2x1p5_ASAP7_75t_L g3656 ( 
.A(n_3531),
.B(n_3277),
.Y(n_3656)
);

INVxp67_ASAP7_75t_SL g3657 ( 
.A(n_3549),
.Y(n_3657)
);

INVx2_ASAP7_75t_L g3658 ( 
.A(n_3422),
.Y(n_3658)
);

OAI21x1_ASAP7_75t_L g3659 ( 
.A1(n_3403),
.A2(n_2369),
.B(n_2346),
.Y(n_3659)
);

OAI21x1_ASAP7_75t_L g3660 ( 
.A1(n_3506),
.A2(n_2584),
.B(n_2399),
.Y(n_3660)
);

AO31x2_ASAP7_75t_L g3661 ( 
.A1(n_3478),
.A2(n_3461),
.A3(n_3437),
.B(n_3421),
.Y(n_3661)
);

OA21x2_ASAP7_75t_L g3662 ( 
.A1(n_3420),
.A2(n_2721),
.B(n_2903),
.Y(n_3662)
);

INVx1_ASAP7_75t_L g3663 ( 
.A(n_3430),
.Y(n_3663)
);

OAI22xp5_ASAP7_75t_L g3664 ( 
.A1(n_3582),
.A2(n_3337),
.B1(n_3277),
.B2(n_2904),
.Y(n_3664)
);

OAI21x1_ASAP7_75t_L g3665 ( 
.A1(n_3524),
.A2(n_2440),
.B(n_2696),
.Y(n_3665)
);

AOI21xp5_ASAP7_75t_L g3666 ( 
.A1(n_3497),
.A2(n_2919),
.B(n_2903),
.Y(n_3666)
);

OAI21x1_ASAP7_75t_L g3667 ( 
.A1(n_3548),
.A2(n_2440),
.B(n_2696),
.Y(n_3667)
);

AOI21xp5_ASAP7_75t_L g3668 ( 
.A1(n_3409),
.A2(n_2927),
.B(n_2919),
.Y(n_3668)
);

OAI22xp5_ASAP7_75t_L g3669 ( 
.A1(n_3554),
.A2(n_3528),
.B1(n_3466),
.B2(n_3516),
.Y(n_3669)
);

AOI21xp5_ASAP7_75t_L g3670 ( 
.A1(n_3472),
.A2(n_2927),
.B(n_2904),
.Y(n_3670)
);

INVx2_ASAP7_75t_L g3671 ( 
.A(n_3467),
.Y(n_3671)
);

NAND2xp5_ASAP7_75t_SL g3672 ( 
.A(n_3406),
.B(n_3337),
.Y(n_3672)
);

AOI21xp5_ASAP7_75t_L g3673 ( 
.A1(n_3475),
.A2(n_2904),
.B(n_2895),
.Y(n_3673)
);

CKINVDCx6p67_ASAP7_75t_R g3674 ( 
.A(n_3511),
.Y(n_3674)
);

AO31x2_ASAP7_75t_L g3675 ( 
.A1(n_3413),
.A2(n_2922),
.A3(n_2906),
.B(n_2743),
.Y(n_3675)
);

NAND2xp5_ASAP7_75t_L g3676 ( 
.A(n_3452),
.B(n_3277),
.Y(n_3676)
);

AOI21xp5_ASAP7_75t_L g3677 ( 
.A1(n_3471),
.A2(n_2922),
.B(n_2906),
.Y(n_3677)
);

NOR2xp33_ASAP7_75t_L g3678 ( 
.A(n_3445),
.B(n_148),
.Y(n_3678)
);

AND2x2_ASAP7_75t_L g3679 ( 
.A(n_3473),
.B(n_2714),
.Y(n_3679)
);

NAND2xp5_ASAP7_75t_L g3680 ( 
.A(n_3499),
.B(n_149),
.Y(n_3680)
);

NOR2xp33_ASAP7_75t_L g3681 ( 
.A(n_3481),
.B(n_149),
.Y(n_3681)
);

NAND2xp5_ASAP7_75t_L g3682 ( 
.A(n_3504),
.B(n_150),
.Y(n_3682)
);

CKINVDCx8_ASAP7_75t_R g3683 ( 
.A(n_3507),
.Y(n_3683)
);

OAI21xp5_ASAP7_75t_L g3684 ( 
.A1(n_3411),
.A2(n_69),
.B(n_70),
.Y(n_3684)
);

BUFx2_ASAP7_75t_L g3685 ( 
.A(n_3567),
.Y(n_3685)
);

AOI21xp5_ASAP7_75t_SL g3686 ( 
.A1(n_3512),
.A2(n_3580),
.B(n_3574),
.Y(n_3686)
);

AOI21xp5_ASAP7_75t_L g3687 ( 
.A1(n_3410),
.A2(n_2922),
.B(n_2906),
.Y(n_3687)
);

BUFx3_ASAP7_75t_L g3688 ( 
.A(n_3432),
.Y(n_3688)
);

AOI21xp5_ASAP7_75t_L g3689 ( 
.A1(n_3508),
.A2(n_2743),
.B(n_2714),
.Y(n_3689)
);

CKINVDCx20_ASAP7_75t_R g3690 ( 
.A(n_3469),
.Y(n_3690)
);

AOI21x1_ASAP7_75t_SL g3691 ( 
.A1(n_3557),
.A2(n_152),
.B(n_151),
.Y(n_3691)
);

OAI21x1_ASAP7_75t_L g3692 ( 
.A1(n_3569),
.A2(n_2743),
.B(n_2714),
.Y(n_3692)
);

OAI21x1_ASAP7_75t_SL g3693 ( 
.A1(n_3449),
.A2(n_3553),
.B(n_3443),
.Y(n_3693)
);

NOR2x1_ASAP7_75t_SL g3694 ( 
.A(n_3451),
.B(n_2756),
.Y(n_3694)
);

AOI22xp5_ASAP7_75t_L g3695 ( 
.A1(n_3412),
.A2(n_2757),
.B1(n_2771),
.B2(n_2756),
.Y(n_3695)
);

INVx5_ASAP7_75t_L g3696 ( 
.A(n_3426),
.Y(n_3696)
);

AND2x6_ASAP7_75t_L g3697 ( 
.A(n_3448),
.B(n_2756),
.Y(n_3697)
);

AOI21xp5_ASAP7_75t_L g3698 ( 
.A1(n_3519),
.A2(n_3417),
.B(n_3503),
.Y(n_3698)
);

NAND2xp33_ASAP7_75t_SL g3699 ( 
.A(n_3450),
.B(n_2757),
.Y(n_3699)
);

INVx2_ASAP7_75t_L g3700 ( 
.A(n_3513),
.Y(n_3700)
);

AO31x2_ASAP7_75t_L g3701 ( 
.A1(n_3457),
.A2(n_2771),
.A3(n_2791),
.B(n_2757),
.Y(n_3701)
);

A2O1A1Ixp33_ASAP7_75t_L g3702 ( 
.A1(n_3470),
.A2(n_3423),
.B(n_3407),
.C(n_3456),
.Y(n_3702)
);

NAND2xp5_ASAP7_75t_L g3703 ( 
.A(n_3530),
.B(n_152),
.Y(n_3703)
);

NAND2xp5_ASAP7_75t_L g3704 ( 
.A(n_3546),
.B(n_153),
.Y(n_3704)
);

NAND3xp33_ASAP7_75t_SL g3705 ( 
.A(n_3416),
.B(n_69),
.C(n_71),
.Y(n_3705)
);

BUFx6f_ASAP7_75t_L g3706 ( 
.A(n_3432),
.Y(n_3706)
);

INVx2_ASAP7_75t_SL g3707 ( 
.A(n_3589),
.Y(n_3707)
);

OAI21x1_ASAP7_75t_L g3708 ( 
.A1(n_3573),
.A2(n_2771),
.B(n_2791),
.Y(n_3708)
);

AOI21xp5_ASAP7_75t_L g3709 ( 
.A1(n_3418),
.A2(n_2794),
.B(n_2791),
.Y(n_3709)
);

INVx1_ASAP7_75t_L g3710 ( 
.A(n_3563),
.Y(n_3710)
);

OAI21x1_ASAP7_75t_L g3711 ( 
.A1(n_3439),
.A2(n_2794),
.B(n_2799),
.Y(n_3711)
);

OAI21x1_ASAP7_75t_L g3712 ( 
.A1(n_3551),
.A2(n_2794),
.B(n_2799),
.Y(n_3712)
);

INVx1_ASAP7_75t_L g3713 ( 
.A(n_3578),
.Y(n_3713)
);

INVx1_ASAP7_75t_L g3714 ( 
.A(n_3544),
.Y(n_3714)
);

NAND2xp5_ASAP7_75t_L g3715 ( 
.A(n_3509),
.B(n_3510),
.Y(n_3715)
);

OAI22xp5_ASAP7_75t_L g3716 ( 
.A1(n_3455),
.A2(n_2807),
.B1(n_2799),
.B2(n_2820),
.Y(n_3716)
);

AO31x2_ASAP7_75t_L g3717 ( 
.A1(n_3426),
.A2(n_2820),
.A3(n_2807),
.B(n_72),
.Y(n_3717)
);

AO31x2_ASAP7_75t_L g3718 ( 
.A1(n_3599),
.A2(n_2820),
.A3(n_2807),
.B(n_72),
.Y(n_3718)
);

INVx1_ASAP7_75t_L g3719 ( 
.A(n_3518),
.Y(n_3719)
);

AOI21xp5_ASAP7_75t_L g3720 ( 
.A1(n_3597),
.A2(n_69),
.B(n_71),
.Y(n_3720)
);

OAI21xp5_ASAP7_75t_L g3721 ( 
.A1(n_3523),
.A2(n_79),
.B(n_71),
.Y(n_3721)
);

INVx1_ASAP7_75t_L g3722 ( 
.A(n_3518),
.Y(n_3722)
);

OAI21xp5_ASAP7_75t_L g3723 ( 
.A1(n_3500),
.A2(n_80),
.B(n_72),
.Y(n_3723)
);

AOI21xp5_ASAP7_75t_L g3724 ( 
.A1(n_3598),
.A2(n_73),
.B(n_74),
.Y(n_3724)
);

INVx1_ASAP7_75t_L g3725 ( 
.A(n_3518),
.Y(n_3725)
);

HB1xp67_ASAP7_75t_L g3726 ( 
.A(n_3468),
.Y(n_3726)
);

AOI211x1_ASAP7_75t_L g3727 ( 
.A1(n_3427),
.A2(n_170),
.B(n_180),
.C(n_161),
.Y(n_3727)
);

O2A1O1Ixp33_ASAP7_75t_L g3728 ( 
.A1(n_3474),
.A2(n_75),
.B(n_73),
.C(n_74),
.Y(n_3728)
);

OAI21x1_ASAP7_75t_L g3729 ( 
.A1(n_3482),
.A2(n_3559),
.B(n_3535),
.Y(n_3729)
);

NOR2xp33_ASAP7_75t_L g3730 ( 
.A(n_3514),
.B(n_153),
.Y(n_3730)
);

NAND2xp5_ASAP7_75t_SL g3731 ( 
.A(n_3596),
.B(n_154),
.Y(n_3731)
);

INVx1_ASAP7_75t_L g3732 ( 
.A(n_3453),
.Y(n_3732)
);

NAND2xp5_ASAP7_75t_L g3733 ( 
.A(n_3505),
.B(n_154),
.Y(n_3733)
);

OAI21x1_ASAP7_75t_L g3734 ( 
.A1(n_3550),
.A2(n_73),
.B(n_75),
.Y(n_3734)
);

AND2x2_ASAP7_75t_L g3735 ( 
.A(n_3479),
.B(n_685),
.Y(n_3735)
);

AOI21xp5_ASAP7_75t_L g3736 ( 
.A1(n_3484),
.A2(n_75),
.B(n_76),
.Y(n_3736)
);

OAI21x1_ASAP7_75t_L g3737 ( 
.A1(n_3595),
.A2(n_3602),
.B(n_3527),
.Y(n_3737)
);

OAI21x1_ASAP7_75t_L g3738 ( 
.A1(n_3441),
.A2(n_77),
.B(n_78),
.Y(n_3738)
);

CKINVDCx16_ASAP7_75t_R g3739 ( 
.A(n_3564),
.Y(n_3739)
);

AND2x4_ASAP7_75t_L g3740 ( 
.A(n_3575),
.B(n_77),
.Y(n_3740)
);

OAI21xp5_ASAP7_75t_L g3741 ( 
.A1(n_3498),
.A2(n_3447),
.B(n_3542),
.Y(n_3741)
);

NAND2xp5_ASAP7_75t_L g3742 ( 
.A(n_3463),
.B(n_155),
.Y(n_3742)
);

AND2x2_ASAP7_75t_L g3743 ( 
.A(n_3501),
.B(n_692),
.Y(n_3743)
);

INVx2_ASAP7_75t_L g3744 ( 
.A(n_3588),
.Y(n_3744)
);

OAI21x1_ASAP7_75t_L g3745 ( 
.A1(n_3558),
.A2(n_78),
.B(n_79),
.Y(n_3745)
);

O2A1O1Ixp5_ASAP7_75t_L g3746 ( 
.A1(n_3577),
.A2(n_82),
.B(n_79),
.C(n_81),
.Y(n_3746)
);

A2O1A1Ixp33_ASAP7_75t_L g3747 ( 
.A1(n_3538),
.A2(n_156),
.B(n_157),
.C(n_155),
.Y(n_3747)
);

AO21x1_ASAP7_75t_L g3748 ( 
.A1(n_3545),
.A2(n_81),
.B(n_82),
.Y(n_3748)
);

AOI21xp5_ASAP7_75t_L g3749 ( 
.A1(n_3484),
.A2(n_81),
.B(n_82),
.Y(n_3749)
);

OAI21x1_ASAP7_75t_L g3750 ( 
.A1(n_3561),
.A2(n_83),
.B(n_84),
.Y(n_3750)
);

A2O1A1Ixp33_ASAP7_75t_L g3751 ( 
.A1(n_3489),
.A2(n_157),
.B(n_159),
.C(n_156),
.Y(n_3751)
);

AOI21xp5_ASAP7_75t_L g3752 ( 
.A1(n_3484),
.A2(n_83),
.B(n_84),
.Y(n_3752)
);

OAI21x1_ASAP7_75t_L g3753 ( 
.A1(n_3570),
.A2(n_83),
.B(n_85),
.Y(n_3753)
);

AOI21xp5_ASAP7_75t_L g3754 ( 
.A1(n_3477),
.A2(n_3583),
.B(n_3605),
.Y(n_3754)
);

BUFx2_ASAP7_75t_L g3755 ( 
.A(n_3565),
.Y(n_3755)
);

AND2x2_ASAP7_75t_L g3756 ( 
.A(n_3520),
.B(n_679),
.Y(n_3756)
);

INVx1_ASAP7_75t_L g3757 ( 
.A(n_3536),
.Y(n_3757)
);

NAND2xp5_ASAP7_75t_L g3758 ( 
.A(n_3534),
.B(n_160),
.Y(n_3758)
);

AO31x2_ASAP7_75t_L g3759 ( 
.A1(n_3487),
.A2(n_87),
.A3(n_85),
.B(n_86),
.Y(n_3759)
);

NAND2xp5_ASAP7_75t_L g3760 ( 
.A(n_3532),
.B(n_160),
.Y(n_3760)
);

OAI21xp5_ASAP7_75t_L g3761 ( 
.A1(n_3576),
.A2(n_3566),
.B(n_3462),
.Y(n_3761)
);

AOI21xp5_ASAP7_75t_L g3762 ( 
.A1(n_3584),
.A2(n_3517),
.B(n_3489),
.Y(n_3762)
);

INVx3_ASAP7_75t_L g3763 ( 
.A(n_3485),
.Y(n_3763)
);

OAI22xp5_ASAP7_75t_L g3764 ( 
.A1(n_3464),
.A2(n_88),
.B1(n_85),
.B2(n_87),
.Y(n_3764)
);

AOI21xp5_ASAP7_75t_L g3765 ( 
.A1(n_3517),
.A2(n_88),
.B(n_89),
.Y(n_3765)
);

INVx3_ASAP7_75t_L g3766 ( 
.A(n_3485),
.Y(n_3766)
);

OAI21xp5_ASAP7_75t_L g3767 ( 
.A1(n_3541),
.A2(n_88),
.B(n_89),
.Y(n_3767)
);

NAND2xp5_ASAP7_75t_L g3768 ( 
.A(n_3537),
.B(n_3568),
.Y(n_3768)
);

NAND2xp5_ASAP7_75t_L g3769 ( 
.A(n_3592),
.B(n_161),
.Y(n_3769)
);

NAND2xp5_ASAP7_75t_L g3770 ( 
.A(n_3601),
.B(n_162),
.Y(n_3770)
);

INVx1_ASAP7_75t_L g3771 ( 
.A(n_3604),
.Y(n_3771)
);

NAND2xp5_ASAP7_75t_L g3772 ( 
.A(n_3543),
.B(n_162),
.Y(n_3772)
);

AOI21xp5_ASAP7_75t_L g3773 ( 
.A1(n_3571),
.A2(n_90),
.B(n_91),
.Y(n_3773)
);

INVx4_ASAP7_75t_L g3774 ( 
.A(n_3485),
.Y(n_3774)
);

AO31x2_ASAP7_75t_L g3775 ( 
.A1(n_3547),
.A2(n_92),
.A3(n_90),
.B(n_91),
.Y(n_3775)
);

NAND2xp5_ASAP7_75t_L g3776 ( 
.A(n_3465),
.B(n_164),
.Y(n_3776)
);

NAND2xp5_ASAP7_75t_L g3777 ( 
.A(n_3465),
.B(n_164),
.Y(n_3777)
);

OAI21x1_ASAP7_75t_L g3778 ( 
.A1(n_3572),
.A2(n_90),
.B(n_92),
.Y(n_3778)
);

NAND2xp5_ASAP7_75t_L g3779 ( 
.A(n_3515),
.B(n_165),
.Y(n_3779)
);

NAND2xp5_ASAP7_75t_L g3780 ( 
.A(n_3515),
.B(n_166),
.Y(n_3780)
);

AOI21x1_ASAP7_75t_L g3781 ( 
.A1(n_3581),
.A2(n_3491),
.B(n_3490),
.Y(n_3781)
);

OAI22xp5_ASAP7_75t_L g3782 ( 
.A1(n_3591),
.A2(n_95),
.B1(n_93),
.B2(n_94),
.Y(n_3782)
);

NAND2xp5_ASAP7_75t_SL g3783 ( 
.A(n_3591),
.B(n_167),
.Y(n_3783)
);

AOI21xp5_ASAP7_75t_SL g3784 ( 
.A1(n_3556),
.A2(n_169),
.B(n_168),
.Y(n_3784)
);

AOI21xp5_ASAP7_75t_L g3785 ( 
.A1(n_3521),
.A2(n_93),
.B(n_95),
.Y(n_3785)
);

AOI21x1_ASAP7_75t_L g3786 ( 
.A1(n_3490),
.A2(n_95),
.B(n_96),
.Y(n_3786)
);

INVx1_ASAP7_75t_L g3787 ( 
.A(n_3560),
.Y(n_3787)
);

INVx4_ASAP7_75t_L g3788 ( 
.A(n_3547),
.Y(n_3788)
);

NAND2xp5_ASAP7_75t_L g3789 ( 
.A(n_3526),
.B(n_168),
.Y(n_3789)
);

AOI22xp5_ASAP7_75t_L g3790 ( 
.A1(n_3533),
.A2(n_98),
.B1(n_96),
.B2(n_97),
.Y(n_3790)
);

NAND2xp5_ASAP7_75t_L g3791 ( 
.A(n_3600),
.B(n_3560),
.Y(n_3791)
);

NAND2xp5_ASAP7_75t_L g3792 ( 
.A(n_3560),
.B(n_3593),
.Y(n_3792)
);

AOI21xp33_ASAP7_75t_L g3793 ( 
.A1(n_3603),
.A2(n_97),
.B(n_98),
.Y(n_3793)
);

AO31x2_ASAP7_75t_L g3794 ( 
.A1(n_3590),
.A2(n_3540),
.A3(n_3529),
.B(n_3491),
.Y(n_3794)
);

NAND2xp5_ASAP7_75t_L g3795 ( 
.A(n_3593),
.B(n_170),
.Y(n_3795)
);

NAND2xp5_ASAP7_75t_L g3796 ( 
.A(n_3593),
.B(n_171),
.Y(n_3796)
);

OAI21xp33_ASAP7_75t_L g3797 ( 
.A1(n_3525),
.A2(n_97),
.B(n_98),
.Y(n_3797)
);

AOI21x1_ASAP7_75t_L g3798 ( 
.A1(n_3529),
.A2(n_99),
.B(n_100),
.Y(n_3798)
);

OAI21x1_ASAP7_75t_SL g3799 ( 
.A1(n_3590),
.A2(n_99),
.B(n_100),
.Y(n_3799)
);

OAI21xp5_ASAP7_75t_L g3800 ( 
.A1(n_3428),
.A2(n_101),
.B(n_102),
.Y(n_3800)
);

A2O1A1Ixp33_ASAP7_75t_L g3801 ( 
.A1(n_3442),
.A2(n_175),
.B(n_176),
.C(n_172),
.Y(n_3801)
);

NAND3xp33_ASAP7_75t_L g3802 ( 
.A(n_3552),
.B(n_102),
.C(n_103),
.Y(n_3802)
);

NAND2xp5_ASAP7_75t_L g3803 ( 
.A(n_3493),
.B(n_172),
.Y(n_3803)
);

AOI21xp5_ASAP7_75t_L g3804 ( 
.A1(n_3397),
.A2(n_102),
.B(n_103),
.Y(n_3804)
);

INVx2_ASAP7_75t_L g3805 ( 
.A(n_3398),
.Y(n_3805)
);

A2O1A1Ixp33_ASAP7_75t_L g3806 ( 
.A1(n_3397),
.A2(n_176),
.B(n_177),
.C(n_175),
.Y(n_3806)
);

OAI21xp5_ASAP7_75t_L g3807 ( 
.A1(n_3397),
.A2(n_103),
.B(n_104),
.Y(n_3807)
);

AOI21x1_ASAP7_75t_SL g3808 ( 
.A1(n_3557),
.A2(n_178),
.B(n_177),
.Y(n_3808)
);

AOI22xp5_ASAP7_75t_L g3809 ( 
.A1(n_3438),
.A2(n_106),
.B1(n_104),
.B2(n_105),
.Y(n_3809)
);

OAI21xp5_ASAP7_75t_L g3810 ( 
.A1(n_3397),
.A2(n_104),
.B(n_105),
.Y(n_3810)
);

AOI21x1_ASAP7_75t_L g3811 ( 
.A1(n_3476),
.A2(n_106),
.B(n_178),
.Y(n_3811)
);

AND2x2_ASAP7_75t_L g3812 ( 
.A(n_3429),
.B(n_694),
.Y(n_3812)
);

OAI21x1_ASAP7_75t_SL g3813 ( 
.A1(n_3397),
.A2(n_179),
.B(n_180),
.Y(n_3813)
);

NAND2xp5_ASAP7_75t_L g3814 ( 
.A(n_3431),
.B(n_179),
.Y(n_3814)
);

BUFx12f_ASAP7_75t_L g3815 ( 
.A(n_3507),
.Y(n_3815)
);

OR2x2_ASAP7_75t_L g3816 ( 
.A(n_3494),
.B(n_181),
.Y(n_3816)
);

OAI21x1_ASAP7_75t_L g3817 ( 
.A1(n_3562),
.A2(n_182),
.B(n_183),
.Y(n_3817)
);

OAI21xp5_ASAP7_75t_L g3818 ( 
.A1(n_3397),
.A2(n_183),
.B(n_184),
.Y(n_3818)
);

NAND2xp5_ASAP7_75t_L g3819 ( 
.A(n_3431),
.B(n_185),
.Y(n_3819)
);

BUFx2_ASAP7_75t_L g3820 ( 
.A(n_3494),
.Y(n_3820)
);

NAND3xp33_ASAP7_75t_SL g3821 ( 
.A(n_3555),
.B(n_185),
.C(n_186),
.Y(n_3821)
);

OR2x2_ASAP7_75t_L g3822 ( 
.A(n_3494),
.B(n_187),
.Y(n_3822)
);

OAI21x1_ASAP7_75t_L g3823 ( 
.A1(n_3562),
.A2(n_187),
.B(n_188),
.Y(n_3823)
);

OAI21x1_ASAP7_75t_SL g3824 ( 
.A1(n_3397),
.A2(n_189),
.B(n_190),
.Y(n_3824)
);

OAI21x1_ASAP7_75t_L g3825 ( 
.A1(n_3562),
.A2(n_189),
.B(n_190),
.Y(n_3825)
);

OAI21x1_ASAP7_75t_L g3826 ( 
.A1(n_3562),
.A2(n_191),
.B(n_193),
.Y(n_3826)
);

INVx4_ASAP7_75t_SL g3827 ( 
.A(n_3565),
.Y(n_3827)
);

INVx1_ASAP7_75t_L g3828 ( 
.A(n_3586),
.Y(n_3828)
);

NAND2xp5_ASAP7_75t_L g3829 ( 
.A(n_3431),
.B(n_191),
.Y(n_3829)
);

NAND2xp5_ASAP7_75t_L g3830 ( 
.A(n_3431),
.B(n_193),
.Y(n_3830)
);

AOI21xp5_ASAP7_75t_L g3831 ( 
.A1(n_3397),
.A2(n_195),
.B(n_196),
.Y(n_3831)
);

O2A1O1Ixp33_ASAP7_75t_L g3832 ( 
.A1(n_3806),
.A2(n_198),
.B(n_195),
.C(n_197),
.Y(n_3832)
);

OAI22xp5_ASAP7_75t_L g3833 ( 
.A1(n_3809),
.A2(n_200),
.B1(n_197),
.B2(n_199),
.Y(n_3833)
);

A2O1A1Ixp33_ASAP7_75t_L g3834 ( 
.A1(n_3818),
.A2(n_202),
.B(n_200),
.C(n_201),
.Y(n_3834)
);

CKINVDCx20_ASAP7_75t_R g3835 ( 
.A(n_3690),
.Y(n_3835)
);

INVx3_ASAP7_75t_SL g3836 ( 
.A(n_3674),
.Y(n_3836)
);

NAND2xp5_ASAP7_75t_L g3837 ( 
.A(n_3732),
.B(n_201),
.Y(n_3837)
);

OAI21x1_ASAP7_75t_L g3838 ( 
.A1(n_3698),
.A2(n_202),
.B(n_203),
.Y(n_3838)
);

INVx1_ASAP7_75t_L g3839 ( 
.A(n_3648),
.Y(n_3839)
);

AO32x2_ASAP7_75t_L g3840 ( 
.A1(n_3669),
.A2(n_206),
.A3(n_203),
.B1(n_205),
.B2(n_207),
.Y(n_3840)
);

INVx2_ASAP7_75t_SL g3841 ( 
.A(n_3628),
.Y(n_3841)
);

BUFx6f_ASAP7_75t_L g3842 ( 
.A(n_3628),
.Y(n_3842)
);

CKINVDCx5p33_ASAP7_75t_R g3843 ( 
.A(n_3815),
.Y(n_3843)
);

AOI21xp5_ASAP7_75t_L g3844 ( 
.A1(n_3611),
.A2(n_3686),
.B(n_3807),
.Y(n_3844)
);

NAND2xp5_ASAP7_75t_L g3845 ( 
.A(n_3713),
.B(n_205),
.Y(n_3845)
);

INVx3_ASAP7_75t_L g3846 ( 
.A(n_3628),
.Y(n_3846)
);

CKINVDCx11_ASAP7_75t_R g3847 ( 
.A(n_3683),
.Y(n_3847)
);

INVx2_ASAP7_75t_L g3848 ( 
.A(n_3629),
.Y(n_3848)
);

AOI21xp5_ASAP7_75t_L g3849 ( 
.A1(n_3810),
.A2(n_207),
.B(n_208),
.Y(n_3849)
);

NAND2x1p5_ASAP7_75t_L g3850 ( 
.A(n_3635),
.B(n_208),
.Y(n_3850)
);

O2A1O1Ixp33_ASAP7_75t_L g3851 ( 
.A1(n_3684),
.A2(n_211),
.B(n_209),
.C(n_210),
.Y(n_3851)
);

AOI21xp5_ASAP7_75t_L g3852 ( 
.A1(n_3618),
.A2(n_210),
.B(n_211),
.Y(n_3852)
);

AO22x2_ASAP7_75t_L g3853 ( 
.A1(n_3719),
.A2(n_214),
.B1(n_212),
.B2(n_213),
.Y(n_3853)
);

NOR2xp67_ASAP7_75t_L g3854 ( 
.A(n_3625),
.B(n_212),
.Y(n_3854)
);

OAI21x1_ASAP7_75t_L g3855 ( 
.A1(n_3729),
.A2(n_213),
.B(n_214),
.Y(n_3855)
);

AO31x2_ASAP7_75t_L g3856 ( 
.A1(n_3736),
.A2(n_217),
.A3(n_215),
.B(n_216),
.Y(n_3856)
);

OAI21xp5_ASAP7_75t_L g3857 ( 
.A1(n_3831),
.A2(n_215),
.B(n_216),
.Y(n_3857)
);

BUFx2_ASAP7_75t_L g3858 ( 
.A(n_3820),
.Y(n_3858)
);

OAI21xp5_ASAP7_75t_L g3859 ( 
.A1(n_3804),
.A2(n_217),
.B(n_218),
.Y(n_3859)
);

AND2x2_ASAP7_75t_L g3860 ( 
.A(n_3685),
.B(n_218),
.Y(n_3860)
);

OAI21x1_ASAP7_75t_L g3861 ( 
.A1(n_3620),
.A2(n_219),
.B(n_220),
.Y(n_3861)
);

NAND3xp33_ASAP7_75t_L g3862 ( 
.A(n_3809),
.B(n_219),
.C(n_220),
.Y(n_3862)
);

AOI21xp5_ASAP7_75t_L g3863 ( 
.A1(n_3668),
.A2(n_221),
.B(n_222),
.Y(n_3863)
);

INVx1_ASAP7_75t_SL g3864 ( 
.A(n_3688),
.Y(n_3864)
);

AOI21xp5_ASAP7_75t_L g3865 ( 
.A1(n_3721),
.A2(n_221),
.B(n_222),
.Y(n_3865)
);

NAND2xp5_ASAP7_75t_L g3866 ( 
.A(n_3607),
.B(n_223),
.Y(n_3866)
);

AOI21xp5_ASAP7_75t_L g3867 ( 
.A1(n_3721),
.A2(n_223),
.B(n_224),
.Y(n_3867)
);

AO31x2_ASAP7_75t_L g3868 ( 
.A1(n_3749),
.A2(n_226),
.A3(n_224),
.B(n_225),
.Y(n_3868)
);

INVx1_ASAP7_75t_L g3869 ( 
.A(n_3617),
.Y(n_3869)
);

INVx1_ASAP7_75t_SL g3870 ( 
.A(n_3706),
.Y(n_3870)
);

NOR4xp25_ASAP7_75t_L g3871 ( 
.A(n_3802),
.B(n_3705),
.C(n_3821),
.D(n_3797),
.Y(n_3871)
);

OAI21x1_ASAP7_75t_L g3872 ( 
.A1(n_3660),
.A2(n_225),
.B(n_227),
.Y(n_3872)
);

NAND2xp5_ASAP7_75t_L g3873 ( 
.A(n_3609),
.B(n_228),
.Y(n_3873)
);

AO31x2_ASAP7_75t_L g3874 ( 
.A1(n_3752),
.A2(n_230),
.A3(n_228),
.B(n_229),
.Y(n_3874)
);

INVx1_ASAP7_75t_L g3875 ( 
.A(n_3631),
.Y(n_3875)
);

INVx3_ASAP7_75t_L g3876 ( 
.A(n_3706),
.Y(n_3876)
);

O2A1O1Ixp33_ASAP7_75t_L g3877 ( 
.A1(n_3751),
.A2(n_231),
.B(n_229),
.C(n_230),
.Y(n_3877)
);

INVx3_ASAP7_75t_L g3878 ( 
.A(n_3706),
.Y(n_3878)
);

AO22x2_ASAP7_75t_L g3879 ( 
.A1(n_3722),
.A2(n_233),
.B1(n_231),
.B2(n_232),
.Y(n_3879)
);

AOI21xp5_ASAP7_75t_L g3880 ( 
.A1(n_3702),
.A2(n_232),
.B(n_234),
.Y(n_3880)
);

AND2x2_ASAP7_75t_L g3881 ( 
.A(n_3650),
.B(n_3612),
.Y(n_3881)
);

OR2x6_ASAP7_75t_L g3882 ( 
.A(n_3630),
.B(n_234),
.Y(n_3882)
);

OAI21xp5_ASAP7_75t_L g3883 ( 
.A1(n_3773),
.A2(n_235),
.B(n_236),
.Y(n_3883)
);

INVx1_ASAP7_75t_L g3884 ( 
.A(n_3647),
.Y(n_3884)
);

OAI21x1_ASAP7_75t_L g3885 ( 
.A1(n_3643),
.A2(n_237),
.B(n_238),
.Y(n_3885)
);

AOI21xp5_ASAP7_75t_L g3886 ( 
.A1(n_3723),
.A2(n_237),
.B(n_238),
.Y(n_3886)
);

NOR2xp33_ASAP7_75t_SL g3887 ( 
.A(n_3739),
.B(n_239),
.Y(n_3887)
);

INVxp67_ASAP7_75t_SL g3888 ( 
.A(n_3621),
.Y(n_3888)
);

O2A1O1Ixp33_ASAP7_75t_SL g3889 ( 
.A1(n_3801),
.A2(n_241),
.B(n_239),
.C(n_240),
.Y(n_3889)
);

AOI21xp5_ASAP7_75t_L g3890 ( 
.A1(n_3723),
.A2(n_240),
.B(n_243),
.Y(n_3890)
);

AOI21xp5_ASAP7_75t_L g3891 ( 
.A1(n_3633),
.A2(n_244),
.B(n_246),
.Y(n_3891)
);

OAI22xp33_ASAP7_75t_L g3892 ( 
.A1(n_3802),
.A2(n_248),
.B1(n_244),
.B2(n_247),
.Y(n_3892)
);

AO31x2_ASAP7_75t_L g3893 ( 
.A1(n_3613),
.A2(n_251),
.A3(n_249),
.B(n_250),
.Y(n_3893)
);

OAI21x1_ASAP7_75t_L g3894 ( 
.A1(n_3634),
.A2(n_250),
.B(n_252),
.Y(n_3894)
);

INVx1_ASAP7_75t_L g3895 ( 
.A(n_3651),
.Y(n_3895)
);

O2A1O1Ixp33_ASAP7_75t_L g3896 ( 
.A1(n_3747),
.A2(n_254),
.B(n_252),
.C(n_253),
.Y(n_3896)
);

O2A1O1Ixp33_ASAP7_75t_L g3897 ( 
.A1(n_3800),
.A2(n_255),
.B(n_253),
.C(n_254),
.Y(n_3897)
);

AND2x4_ASAP7_75t_L g3898 ( 
.A(n_3828),
.B(n_255),
.Y(n_3898)
);

OAI21x1_ASAP7_75t_L g3899 ( 
.A1(n_3693),
.A2(n_256),
.B(n_257),
.Y(n_3899)
);

INVx1_ASAP7_75t_L g3900 ( 
.A(n_3805),
.Y(n_3900)
);

NOR2xp33_ASAP7_75t_SL g3901 ( 
.A(n_3739),
.B(n_258),
.Y(n_3901)
);

NOR2xp67_ASAP7_75t_SL g3902 ( 
.A(n_3784),
.B(n_258),
.Y(n_3902)
);

A2O1A1Ixp33_ASAP7_75t_L g3903 ( 
.A1(n_3797),
.A2(n_261),
.B(n_259),
.C(n_260),
.Y(n_3903)
);

NAND3x1_ASAP7_75t_L g3904 ( 
.A(n_3655),
.B(n_3790),
.C(n_3616),
.Y(n_3904)
);

NOR2xp33_ASAP7_75t_L g3905 ( 
.A(n_3678),
.B(n_259),
.Y(n_3905)
);

OAI21x1_ASAP7_75t_L g3906 ( 
.A1(n_3737),
.A2(n_260),
.B(n_261),
.Y(n_3906)
);

CKINVDCx11_ASAP7_75t_R g3907 ( 
.A(n_3827),
.Y(n_3907)
);

AND2x4_ASAP7_75t_L g3908 ( 
.A(n_3794),
.B(n_262),
.Y(n_3908)
);

O2A1O1Ixp33_ASAP7_75t_L g3909 ( 
.A1(n_3765),
.A2(n_265),
.B(n_263),
.C(n_264),
.Y(n_3909)
);

AO31x2_ASAP7_75t_L g3910 ( 
.A1(n_3748),
.A2(n_266),
.A3(n_263),
.B(n_264),
.Y(n_3910)
);

INVx5_ASAP7_75t_L g3911 ( 
.A(n_3622),
.Y(n_3911)
);

O2A1O1Ixp33_ASAP7_75t_L g3912 ( 
.A1(n_3783),
.A2(n_269),
.B(n_267),
.C(n_268),
.Y(n_3912)
);

AND2x2_ASAP7_75t_L g3913 ( 
.A(n_3608),
.B(n_268),
.Y(n_3913)
);

AND2x4_ASAP7_75t_L g3914 ( 
.A(n_3794),
.B(n_269),
.Y(n_3914)
);

OAI21x1_ASAP7_75t_L g3915 ( 
.A1(n_3665),
.A2(n_270),
.B(n_272),
.Y(n_3915)
);

INVx2_ASAP7_75t_L g3916 ( 
.A(n_3663),
.Y(n_3916)
);

O2A1O1Ixp33_ASAP7_75t_SL g3917 ( 
.A1(n_3731),
.A2(n_275),
.B(n_273),
.C(n_274),
.Y(n_3917)
);

AOI221x1_ASAP7_75t_L g3918 ( 
.A1(n_3799),
.A2(n_277),
.B1(n_275),
.B2(n_276),
.C(n_278),
.Y(n_3918)
);

NOR2xp67_ASAP7_75t_L g3919 ( 
.A(n_3696),
.B(n_276),
.Y(n_3919)
);

OAI21x1_ASAP7_75t_L g3920 ( 
.A1(n_3659),
.A2(n_279),
.B(n_281),
.Y(n_3920)
);

AO21x2_ASAP7_75t_L g3921 ( 
.A1(n_3689),
.A2(n_279),
.B(n_281),
.Y(n_3921)
);

AO31x2_ASAP7_75t_L g3922 ( 
.A1(n_3639),
.A2(n_284),
.A3(n_282),
.B(n_283),
.Y(n_3922)
);

AOI21xp5_ASAP7_75t_L g3923 ( 
.A1(n_3646),
.A2(n_282),
.B(n_283),
.Y(n_3923)
);

NAND3xp33_ASAP7_75t_L g3924 ( 
.A(n_3720),
.B(n_285),
.C(n_286),
.Y(n_3924)
);

OAI21x1_ASAP7_75t_L g3925 ( 
.A1(n_3606),
.A2(n_286),
.B(n_287),
.Y(n_3925)
);

BUFx2_ASAP7_75t_L g3926 ( 
.A(n_3794),
.Y(n_3926)
);

INVx2_ASAP7_75t_L g3927 ( 
.A(n_3710),
.Y(n_3927)
);

INVx2_ASAP7_75t_L g3928 ( 
.A(n_3623),
.Y(n_3928)
);

AND2x4_ASAP7_75t_L g3929 ( 
.A(n_3630),
.B(n_287),
.Y(n_3929)
);

NAND2xp5_ASAP7_75t_L g3930 ( 
.A(n_3632),
.B(n_288),
.Y(n_3930)
);

INVx2_ASAP7_75t_L g3931 ( 
.A(n_3658),
.Y(n_3931)
);

AO31x2_ASAP7_75t_L g3932 ( 
.A1(n_3694),
.A2(n_291),
.A3(n_288),
.B(n_289),
.Y(n_3932)
);

NAND2xp33_ASAP7_75t_L g3933 ( 
.A(n_3616),
.B(n_289),
.Y(n_3933)
);

AOI21xp5_ASAP7_75t_L g3934 ( 
.A1(n_3677),
.A2(n_292),
.B(n_293),
.Y(n_3934)
);

INVx4_ASAP7_75t_L g3935 ( 
.A(n_3763),
.Y(n_3935)
);

AO31x2_ASAP7_75t_L g3936 ( 
.A1(n_3714),
.A2(n_295),
.A3(n_292),
.B(n_294),
.Y(n_3936)
);

AO21x1_ASAP7_75t_L g3937 ( 
.A1(n_3672),
.A2(n_3640),
.B(n_3699),
.Y(n_3937)
);

AO31x2_ASAP7_75t_L g3938 ( 
.A1(n_3754),
.A2(n_297),
.A3(n_294),
.B(n_296),
.Y(n_3938)
);

OAI22xp5_ASAP7_75t_L g3939 ( 
.A1(n_3637),
.A2(n_299),
.B1(n_297),
.B2(n_298),
.Y(n_3939)
);

OAI21xp5_ASAP7_75t_L g3940 ( 
.A1(n_3724),
.A2(n_298),
.B(n_299),
.Y(n_3940)
);

O2A1O1Ixp33_ASAP7_75t_SL g3941 ( 
.A1(n_3790),
.A2(n_303),
.B(n_301),
.C(n_302),
.Y(n_3941)
);

OAI21x1_ASAP7_75t_L g3942 ( 
.A1(n_3712),
.A2(n_301),
.B(n_302),
.Y(n_3942)
);

NAND2xp5_ASAP7_75t_L g3943 ( 
.A(n_3715),
.B(n_304),
.Y(n_3943)
);

AOI21xp5_ASAP7_75t_L g3944 ( 
.A1(n_3614),
.A2(n_304),
.B(n_305),
.Y(n_3944)
);

INVx1_ASAP7_75t_L g3945 ( 
.A(n_3619),
.Y(n_3945)
);

A2O1A1Ixp33_ASAP7_75t_L g3946 ( 
.A1(n_3637),
.A2(n_307),
.B(n_305),
.C(n_306),
.Y(n_3946)
);

NOR2xp67_ASAP7_75t_SL g3947 ( 
.A(n_3785),
.B(n_307),
.Y(n_3947)
);

OAI21x1_ASAP7_75t_L g3948 ( 
.A1(n_3817),
.A2(n_308),
.B(n_309),
.Y(n_3948)
);

INVx3_ASAP7_75t_L g3949 ( 
.A(n_3774),
.Y(n_3949)
);

OAI21xp5_ASAP7_75t_L g3950 ( 
.A1(n_3728),
.A2(n_308),
.B(n_310),
.Y(n_3950)
);

NAND2xp5_ASAP7_75t_L g3951 ( 
.A(n_3757),
.B(n_311),
.Y(n_3951)
);

NOR2xp33_ASAP7_75t_L g3952 ( 
.A(n_3768),
.B(n_311),
.Y(n_3952)
);

AO22x2_ASAP7_75t_L g3953 ( 
.A1(n_3725),
.A2(n_314),
.B1(n_312),
.B2(n_313),
.Y(n_3953)
);

BUFx8_ASAP7_75t_SL g3954 ( 
.A(n_3755),
.Y(n_3954)
);

AOI21xp5_ASAP7_75t_L g3955 ( 
.A1(n_3666),
.A2(n_312),
.B(n_314),
.Y(n_3955)
);

NAND2xp5_ASAP7_75t_L g3956 ( 
.A(n_3627),
.B(n_315),
.Y(n_3956)
);

OAI22x1_ASAP7_75t_L g3957 ( 
.A1(n_3695),
.A2(n_318),
.B1(n_316),
.B2(n_317),
.Y(n_3957)
);

AOI21xp5_ASAP7_75t_L g3958 ( 
.A1(n_3657),
.A2(n_316),
.B(n_317),
.Y(n_3958)
);

OAI21xp33_ASAP7_75t_L g3959 ( 
.A1(n_3741),
.A2(n_318),
.B(n_319),
.Y(n_3959)
);

OAI21x1_ASAP7_75t_L g3960 ( 
.A1(n_3823),
.A2(n_320),
.B(n_321),
.Y(n_3960)
);

NOR2xp33_ASAP7_75t_L g3961 ( 
.A(n_3681),
.B(n_320),
.Y(n_3961)
);

OR2x6_ASAP7_75t_L g3962 ( 
.A(n_3630),
.B(n_321),
.Y(n_3962)
);

INVx2_ASAP7_75t_L g3963 ( 
.A(n_3671),
.Y(n_3963)
);

AND2x2_ASAP7_75t_L g3964 ( 
.A(n_3744),
.B(n_3652),
.Y(n_3964)
);

NOR2xp33_ASAP7_75t_L g3965 ( 
.A(n_3789),
.B(n_322),
.Y(n_3965)
);

AO31x2_ASAP7_75t_L g3966 ( 
.A1(n_3622),
.A2(n_324),
.A3(n_322),
.B(n_323),
.Y(n_3966)
);

A2O1A1Ixp33_ASAP7_75t_L g3967 ( 
.A1(n_3644),
.A2(n_327),
.B(n_325),
.C(n_326),
.Y(n_3967)
);

AOI21x1_ASAP7_75t_L g3968 ( 
.A1(n_3811),
.A2(n_325),
.B(n_326),
.Y(n_3968)
);

AOI22xp33_ASAP7_75t_L g3969 ( 
.A1(n_3726),
.A2(n_329),
.B1(n_327),
.B2(n_328),
.Y(n_3969)
);

AOI21xp5_ASAP7_75t_L g3970 ( 
.A1(n_3653),
.A2(n_328),
.B(n_329),
.Y(n_3970)
);

INVx1_ASAP7_75t_L g3971 ( 
.A(n_3700),
.Y(n_3971)
);

INVx1_ASAP7_75t_L g3972 ( 
.A(n_3610),
.Y(n_3972)
);

INVx2_ASAP7_75t_SL g3973 ( 
.A(n_3707),
.Y(n_3973)
);

NAND2xp5_ASAP7_75t_L g3974 ( 
.A(n_3638),
.B(n_330),
.Y(n_3974)
);

OAI21xp5_ASAP7_75t_L g3975 ( 
.A1(n_3738),
.A2(n_3826),
.B(n_3825),
.Y(n_3975)
);

AOI221x1_ASAP7_75t_L g3976 ( 
.A1(n_3813),
.A2(n_333),
.B1(n_330),
.B2(n_331),
.C(n_334),
.Y(n_3976)
);

OAI22x1_ASAP7_75t_L g3977 ( 
.A1(n_3695),
.A2(n_3740),
.B1(n_3735),
.B2(n_3816),
.Y(n_3977)
);

NAND2xp5_ASAP7_75t_L g3978 ( 
.A(n_3771),
.B(n_334),
.Y(n_3978)
);

NAND2xp5_ASAP7_75t_SL g3979 ( 
.A(n_3615),
.B(n_335),
.Y(n_3979)
);

AO31x2_ASAP7_75t_L g3980 ( 
.A1(n_3709),
.A2(n_339),
.A3(n_335),
.B(n_338),
.Y(n_3980)
);

A2O1A1Ixp33_ASAP7_75t_L g3981 ( 
.A1(n_3746),
.A2(n_341),
.B(n_339),
.C(n_340),
.Y(n_3981)
);

BUFx6f_ASAP7_75t_L g3982 ( 
.A(n_3792),
.Y(n_3982)
);

NAND2xp33_ASAP7_75t_L g3983 ( 
.A(n_3642),
.B(n_340),
.Y(n_3983)
);

O2A1O1Ixp33_ASAP7_75t_L g3984 ( 
.A1(n_3824),
.A2(n_344),
.B(n_342),
.C(n_343),
.Y(n_3984)
);

OAI21xp5_ASAP7_75t_L g3985 ( 
.A1(n_3761),
.A2(n_342),
.B(n_344),
.Y(n_3985)
);

NOR2xp33_ASAP7_75t_L g3986 ( 
.A(n_3730),
.B(n_345),
.Y(n_3986)
);

AOI21xp5_ASAP7_75t_L g3987 ( 
.A1(n_3762),
.A2(n_345),
.B(n_346),
.Y(n_3987)
);

NAND2x1p5_ASAP7_75t_L g3988 ( 
.A(n_3696),
.B(n_346),
.Y(n_3988)
);

NAND2xp5_ASAP7_75t_L g3989 ( 
.A(n_3636),
.B(n_347),
.Y(n_3989)
);

OAI21xp5_ASAP7_75t_L g3990 ( 
.A1(n_3767),
.A2(n_347),
.B(n_348),
.Y(n_3990)
);

AOI21xp5_ASAP7_75t_L g3991 ( 
.A1(n_3670),
.A2(n_348),
.B(n_349),
.Y(n_3991)
);

OAI21x1_ASAP7_75t_L g3992 ( 
.A1(n_3667),
.A2(n_349),
.B(n_350),
.Y(n_3992)
);

AOI21xp5_ASAP7_75t_L g3993 ( 
.A1(n_3673),
.A2(n_350),
.B(n_352),
.Y(n_3993)
);

OAI21x1_ASAP7_75t_L g3994 ( 
.A1(n_3624),
.A2(n_352),
.B(n_353),
.Y(n_3994)
);

INVx1_ASAP7_75t_L g3995 ( 
.A(n_3649),
.Y(n_3995)
);

AO31x2_ASAP7_75t_L g3996 ( 
.A1(n_3664),
.A2(n_355),
.A3(n_353),
.B(n_354),
.Y(n_3996)
);

BUFx6f_ASAP7_75t_L g3997 ( 
.A(n_3791),
.Y(n_3997)
);

NOR2xp33_ASAP7_75t_L g3998 ( 
.A(n_3742),
.B(n_354),
.Y(n_3998)
);

NOR2xp67_ASAP7_75t_SL g3999 ( 
.A(n_3696),
.B(n_355),
.Y(n_3999)
);

AO31x2_ASAP7_75t_L g4000 ( 
.A1(n_3788),
.A2(n_358),
.A3(n_356),
.B(n_357),
.Y(n_4000)
);

O2A1O1Ixp33_ASAP7_75t_SL g4001 ( 
.A1(n_3793),
.A2(n_358),
.B(n_356),
.C(n_357),
.Y(n_4001)
);

OAI21xp5_ASAP7_75t_L g4002 ( 
.A1(n_3687),
.A2(n_359),
.B(n_360),
.Y(n_4002)
);

INVx3_ASAP7_75t_SL g4003 ( 
.A(n_3827),
.Y(n_4003)
);

OAI21x1_ASAP7_75t_L g4004 ( 
.A1(n_3711),
.A2(n_359),
.B(n_361),
.Y(n_4004)
);

O2A1O1Ixp33_ASAP7_75t_L g4005 ( 
.A1(n_3782),
.A2(n_363),
.B(n_361),
.C(n_362),
.Y(n_4005)
);

CKINVDCx5p33_ASAP7_75t_R g4006 ( 
.A(n_3676),
.Y(n_4006)
);

BUFx10_ASAP7_75t_L g4007 ( 
.A(n_3740),
.Y(n_4007)
);

INVx1_ASAP7_75t_L g4008 ( 
.A(n_3649),
.Y(n_4008)
);

AOI21xp33_ASAP7_75t_L g4009 ( 
.A1(n_3772),
.A2(n_364),
.B(n_365),
.Y(n_4009)
);

OAI22xp5_ASAP7_75t_L g4010 ( 
.A1(n_3727),
.A2(n_367),
.B1(n_365),
.B2(n_366),
.Y(n_4010)
);

CKINVDCx20_ASAP7_75t_R g4011 ( 
.A(n_3679),
.Y(n_4011)
);

OR2x2_ASAP7_75t_L g4012 ( 
.A(n_3814),
.B(n_366),
.Y(n_4012)
);

AOI22xp33_ASAP7_75t_L g4013 ( 
.A1(n_3844),
.A2(n_3697),
.B1(n_3645),
.B2(n_3803),
.Y(n_4013)
);

NOR2xp67_ASAP7_75t_L g4014 ( 
.A(n_3911),
.B(n_3788),
.Y(n_4014)
);

INVx2_ASAP7_75t_L g4015 ( 
.A(n_3858),
.Y(n_4015)
);

OAI22xp5_ASAP7_75t_L g4016 ( 
.A1(n_3862),
.A2(n_3727),
.B1(n_3716),
.B2(n_3733),
.Y(n_4016)
);

AO31x2_ASAP7_75t_L g4017 ( 
.A1(n_3926),
.A2(n_3774),
.A3(n_3787),
.B(n_3764),
.Y(n_4017)
);

OR2x6_ASAP7_75t_L g4018 ( 
.A(n_3882),
.B(n_3656),
.Y(n_4018)
);

HB1xp67_ASAP7_75t_L g4019 ( 
.A(n_3926),
.Y(n_4019)
);

INVxp33_ASAP7_75t_L g4020 ( 
.A(n_3847),
.Y(n_4020)
);

HB1xp67_ASAP7_75t_L g4021 ( 
.A(n_3858),
.Y(n_4021)
);

AND2x4_ASAP7_75t_L g4022 ( 
.A(n_3995),
.B(n_3781),
.Y(n_4022)
);

AOI22xp33_ASAP7_75t_SL g4023 ( 
.A1(n_3933),
.A2(n_3697),
.B1(n_3734),
.B2(n_3812),
.Y(n_4023)
);

NAND2xp5_ASAP7_75t_SL g4024 ( 
.A(n_3937),
.B(n_3654),
.Y(n_4024)
);

INVx1_ASAP7_75t_L g4025 ( 
.A(n_3869),
.Y(n_4025)
);

AOI21x1_ASAP7_75t_L g4026 ( 
.A1(n_3853),
.A2(n_3798),
.B(n_3786),
.Y(n_4026)
);

BUFx6f_ASAP7_75t_L g4027 ( 
.A(n_3842),
.Y(n_4027)
);

AOI221xp5_ASAP7_75t_L g4028 ( 
.A1(n_3871),
.A2(n_3760),
.B1(n_3758),
.B2(n_3829),
.C(n_3819),
.Y(n_4028)
);

INVx2_ASAP7_75t_L g4029 ( 
.A(n_3916),
.Y(n_4029)
);

AOI221xp5_ASAP7_75t_L g4030 ( 
.A1(n_3892),
.A2(n_3830),
.B1(n_3776),
.B2(n_3780),
.C(n_3779),
.Y(n_4030)
);

AO31x2_ASAP7_75t_L g4031 ( 
.A1(n_3945),
.A2(n_3682),
.A3(n_3703),
.B(n_3680),
.Y(n_4031)
);

OAI21x1_ASAP7_75t_L g4032 ( 
.A1(n_3861),
.A2(n_3626),
.B(n_3692),
.Y(n_4032)
);

INVx2_ASAP7_75t_L g4033 ( 
.A(n_3927),
.Y(n_4033)
);

INVx2_ASAP7_75t_L g4034 ( 
.A(n_3839),
.Y(n_4034)
);

OAI21x1_ASAP7_75t_L g4035 ( 
.A1(n_3855),
.A2(n_3708),
.B(n_3691),
.Y(n_4035)
);

OA21x2_ASAP7_75t_L g4036 ( 
.A1(n_3972),
.A2(n_3753),
.B(n_3750),
.Y(n_4036)
);

HB1xp67_ASAP7_75t_L g4037 ( 
.A(n_3928),
.Y(n_4037)
);

OAI21x1_ASAP7_75t_L g4038 ( 
.A1(n_3975),
.A2(n_3808),
.B(n_3641),
.Y(n_4038)
);

AO21x2_ASAP7_75t_L g4039 ( 
.A1(n_3888),
.A2(n_3873),
.B(n_3866),
.Y(n_4039)
);

NOR2xp33_ASAP7_75t_L g4040 ( 
.A(n_3954),
.B(n_3822),
.Y(n_4040)
);

NAND2xp5_ASAP7_75t_L g4041 ( 
.A(n_3964),
.B(n_3661),
.Y(n_4041)
);

OAI21x1_ASAP7_75t_L g4042 ( 
.A1(n_3872),
.A2(n_3745),
.B(n_3778),
.Y(n_4042)
);

INVx2_ASAP7_75t_L g4043 ( 
.A(n_3848),
.Y(n_4043)
);

AOI221xp5_ASAP7_75t_L g4044 ( 
.A1(n_3941),
.A2(n_3777),
.B1(n_3796),
.B2(n_3795),
.C(n_3769),
.Y(n_4044)
);

INVx1_ASAP7_75t_L g4045 ( 
.A(n_3875),
.Y(n_4045)
);

INVx2_ASAP7_75t_L g4046 ( 
.A(n_3884),
.Y(n_4046)
);

NAND2xp5_ASAP7_75t_L g4047 ( 
.A(n_3971),
.B(n_3661),
.Y(n_4047)
);

BUFx2_ASAP7_75t_R g4048 ( 
.A(n_3836),
.Y(n_4048)
);

INVx2_ASAP7_75t_L g4049 ( 
.A(n_3895),
.Y(n_4049)
);

OAI21x1_ASAP7_75t_L g4050 ( 
.A1(n_3925),
.A2(n_3704),
.B(n_3763),
.Y(n_4050)
);

CKINVDCx11_ASAP7_75t_R g4051 ( 
.A(n_3835),
.Y(n_4051)
);

AND2x4_ASAP7_75t_L g4052 ( 
.A(n_4008),
.B(n_3701),
.Y(n_4052)
);

INVx8_ASAP7_75t_L g4053 ( 
.A(n_3882),
.Y(n_4053)
);

OAI22xp5_ASAP7_75t_L g4054 ( 
.A1(n_3834),
.A2(n_3770),
.B1(n_3766),
.B2(n_3662),
.Y(n_4054)
);

BUFx4f_ASAP7_75t_L g4055 ( 
.A(n_4003),
.Y(n_4055)
);

OAI21xp5_ASAP7_75t_L g4056 ( 
.A1(n_3904),
.A2(n_3756),
.B(n_3743),
.Y(n_4056)
);

INVx1_ASAP7_75t_L g4057 ( 
.A(n_3900),
.Y(n_4057)
);

INVx4_ASAP7_75t_L g4058 ( 
.A(n_3907),
.Y(n_4058)
);

INVx1_ASAP7_75t_L g4059 ( 
.A(n_3931),
.Y(n_4059)
);

NAND2xp5_ASAP7_75t_L g4060 ( 
.A(n_3963),
.B(n_3661),
.Y(n_4060)
);

OAI21x1_ASAP7_75t_L g4061 ( 
.A1(n_3885),
.A2(n_3766),
.B(n_3662),
.Y(n_4061)
);

INVx1_ASAP7_75t_L g4062 ( 
.A(n_3908),
.Y(n_4062)
);

NOR2xp33_ASAP7_75t_SL g4063 ( 
.A(n_3843),
.B(n_3697),
.Y(n_4063)
);

OAI21x1_ASAP7_75t_L g4064 ( 
.A1(n_3994),
.A2(n_3675),
.B(n_3718),
.Y(n_4064)
);

INVx2_ASAP7_75t_L g4065 ( 
.A(n_3982),
.Y(n_4065)
);

OAI21x1_ASAP7_75t_SL g4066 ( 
.A1(n_3886),
.A2(n_3775),
.B(n_3759),
.Y(n_4066)
);

OA21x2_ASAP7_75t_L g4067 ( 
.A1(n_3906),
.A2(n_3775),
.B(n_3759),
.Y(n_4067)
);

NAND2xp5_ASAP7_75t_L g4068 ( 
.A(n_3982),
.B(n_3675),
.Y(n_4068)
);

BUFx2_ASAP7_75t_L g4069 ( 
.A(n_3935),
.Y(n_4069)
);

INVx1_ASAP7_75t_L g4070 ( 
.A(n_3908),
.Y(n_4070)
);

AOI21x1_ASAP7_75t_L g4071 ( 
.A1(n_3853),
.A2(n_3775),
.B(n_3759),
.Y(n_4071)
);

BUFx6f_ASAP7_75t_L g4072 ( 
.A(n_3842),
.Y(n_4072)
);

NAND3xp33_ASAP7_75t_L g4073 ( 
.A(n_3944),
.B(n_3717),
.C(n_3718),
.Y(n_4073)
);

A2O1A1Ixp33_ASAP7_75t_L g4074 ( 
.A1(n_3880),
.A2(n_3717),
.B(n_369),
.C(n_367),
.Y(n_4074)
);

AND2x4_ASAP7_75t_L g4075 ( 
.A(n_3914),
.B(n_3701),
.Y(n_4075)
);

AND2x4_ASAP7_75t_L g4076 ( 
.A(n_3914),
.B(n_3701),
.Y(n_4076)
);

OAI21x1_ASAP7_75t_L g4077 ( 
.A1(n_3894),
.A2(n_3675),
.B(n_3718),
.Y(n_4077)
);

OAI21x1_ASAP7_75t_L g4078 ( 
.A1(n_3920),
.A2(n_3717),
.B(n_3697),
.Y(n_4078)
);

OAI21x1_ASAP7_75t_SL g4079 ( 
.A1(n_3890),
.A2(n_368),
.B(n_369),
.Y(n_4079)
);

HB1xp67_ASAP7_75t_L g4080 ( 
.A(n_3881),
.Y(n_4080)
);

INVx2_ASAP7_75t_L g4081 ( 
.A(n_3997),
.Y(n_4081)
);

INVx4_ASAP7_75t_L g4082 ( 
.A(n_3962),
.Y(n_4082)
);

AND2x4_ASAP7_75t_L g4083 ( 
.A(n_3949),
.B(n_370),
.Y(n_4083)
);

BUFx6f_ASAP7_75t_L g4084 ( 
.A(n_3929),
.Y(n_4084)
);

BUFx3_ASAP7_75t_L g4085 ( 
.A(n_3997),
.Y(n_4085)
);

OAI21x1_ASAP7_75t_L g4086 ( 
.A1(n_3838),
.A2(n_372),
.B(n_373),
.Y(n_4086)
);

NOR2xp33_ASAP7_75t_L g4087 ( 
.A(n_3952),
.B(n_372),
.Y(n_4087)
);

OAI21x1_ASAP7_75t_L g4088 ( 
.A1(n_4004),
.A2(n_373),
.B(n_374),
.Y(n_4088)
);

OA21x2_ASAP7_75t_L g4089 ( 
.A1(n_3899),
.A2(n_3942),
.B(n_3915),
.Y(n_4089)
);

OAI21x1_ASAP7_75t_L g4090 ( 
.A1(n_3992),
.A2(n_375),
.B(n_376),
.Y(n_4090)
);

INVx4_ASAP7_75t_SL g4091 ( 
.A(n_3962),
.Y(n_4091)
);

BUFx3_ASAP7_75t_L g4092 ( 
.A(n_3973),
.Y(n_4092)
);

AOI22xp5_ASAP7_75t_L g4093 ( 
.A1(n_3902),
.A2(n_380),
.B1(n_377),
.B2(n_378),
.Y(n_4093)
);

BUFx2_ASAP7_75t_L g4094 ( 
.A(n_4006),
.Y(n_4094)
);

AOI22x1_ASAP7_75t_L g4095 ( 
.A1(n_3958),
.A2(n_380),
.B1(n_377),
.B2(n_378),
.Y(n_4095)
);

OAI21x1_ASAP7_75t_SL g4096 ( 
.A1(n_3849),
.A2(n_381),
.B(n_382),
.Y(n_4096)
);

OAI21xp5_ASAP7_75t_L g4097 ( 
.A1(n_3863),
.A2(n_381),
.B(n_382),
.Y(n_4097)
);

NAND3xp33_ASAP7_75t_L g4098 ( 
.A(n_3852),
.B(n_383),
.C(n_384),
.Y(n_4098)
);

OAI21x1_ASAP7_75t_L g4099 ( 
.A1(n_3968),
.A2(n_383),
.B(n_384),
.Y(n_4099)
);

INVx1_ASAP7_75t_L g4100 ( 
.A(n_3879),
.Y(n_4100)
);

INVx1_ASAP7_75t_L g4101 ( 
.A(n_3879),
.Y(n_4101)
);

AOI22xp33_ASAP7_75t_SL g4102 ( 
.A1(n_3985),
.A2(n_388),
.B1(n_386),
.B2(n_387),
.Y(n_4102)
);

CKINVDCx20_ASAP7_75t_R g4103 ( 
.A(n_4011),
.Y(n_4103)
);

INVx1_ASAP7_75t_L g4104 ( 
.A(n_3953),
.Y(n_4104)
);

OAI21x1_ASAP7_75t_L g4105 ( 
.A1(n_3968),
.A2(n_386),
.B(n_387),
.Y(n_4105)
);

INVx1_ASAP7_75t_L g4106 ( 
.A(n_3953),
.Y(n_4106)
);

OAI21x1_ASAP7_75t_L g4107 ( 
.A1(n_3955),
.A2(n_3960),
.B(n_3948),
.Y(n_4107)
);

AOI22xp33_ASAP7_75t_L g4108 ( 
.A1(n_3950),
.A2(n_390),
.B1(n_388),
.B2(n_389),
.Y(n_4108)
);

AO31x2_ASAP7_75t_L g4109 ( 
.A1(n_4010),
.A2(n_3957),
.A3(n_3976),
.B(n_3918),
.Y(n_4109)
);

AO31x2_ASAP7_75t_L g4110 ( 
.A1(n_3977),
.A2(n_393),
.A3(n_390),
.B(n_391),
.Y(n_4110)
);

INVx2_ASAP7_75t_L g4111 ( 
.A(n_3841),
.Y(n_4111)
);

OAI22xp33_ASAP7_75t_L g4112 ( 
.A1(n_3887),
.A2(n_394),
.B1(n_391),
.B2(n_393),
.Y(n_4112)
);

CKINVDCx5p33_ASAP7_75t_R g4113 ( 
.A(n_3870),
.Y(n_4113)
);

INVx1_ASAP7_75t_L g4114 ( 
.A(n_3936),
.Y(n_4114)
);

AO21x2_ASAP7_75t_L g4115 ( 
.A1(n_3923),
.A2(n_394),
.B(n_395),
.Y(n_4115)
);

CKINVDCx5p33_ASAP7_75t_R g4116 ( 
.A(n_3846),
.Y(n_4116)
);

OAI21x1_ASAP7_75t_L g4117 ( 
.A1(n_3891),
.A2(n_3934),
.B(n_3993),
.Y(n_4117)
);

AOI21xp5_ASAP7_75t_L g4118 ( 
.A1(n_3851),
.A2(n_396),
.B(n_397),
.Y(n_4118)
);

OR2x2_ASAP7_75t_L g4119 ( 
.A(n_3989),
.B(n_398),
.Y(n_4119)
);

NOR2xp33_ASAP7_75t_R g4120 ( 
.A(n_3901),
.B(n_693),
.Y(n_4120)
);

OAI21x1_ASAP7_75t_L g4121 ( 
.A1(n_3991),
.A2(n_399),
.B(n_400),
.Y(n_4121)
);

OAI22xp5_ASAP7_75t_L g4122 ( 
.A1(n_3967),
.A2(n_401),
.B1(n_399),
.B2(n_400),
.Y(n_4122)
);

NOR2xp33_ASAP7_75t_L g4123 ( 
.A(n_3965),
.B(n_402),
.Y(n_4123)
);

AOI21xp5_ASAP7_75t_L g4124 ( 
.A1(n_3865),
.A2(n_691),
.B(n_402),
.Y(n_4124)
);

OAI22xp33_ASAP7_75t_L g4125 ( 
.A1(n_3970),
.A2(n_406),
.B1(n_403),
.B2(n_405),
.Y(n_4125)
);

OR2x6_ASAP7_75t_L g4126 ( 
.A(n_3929),
.B(n_403),
.Y(n_4126)
);

NAND2x1p5_ASAP7_75t_L g4127 ( 
.A(n_3911),
.B(n_407),
.Y(n_4127)
);

INVx2_ASAP7_75t_L g4128 ( 
.A(n_3876),
.Y(n_4128)
);

AOI21x1_ASAP7_75t_L g4129 ( 
.A1(n_3845),
.A2(n_409),
.B(n_410),
.Y(n_4129)
);

AND2x6_ASAP7_75t_L g4130 ( 
.A(n_3898),
.B(n_409),
.Y(n_4130)
);

OAI21x1_ASAP7_75t_L g4131 ( 
.A1(n_3837),
.A2(n_410),
.B(n_412),
.Y(n_4131)
);

BUFx2_ASAP7_75t_L g4132 ( 
.A(n_3878),
.Y(n_4132)
);

OA21x2_ASAP7_75t_L g4133 ( 
.A1(n_3951),
.A2(n_412),
.B(n_413),
.Y(n_4133)
);

OAI21x1_ASAP7_75t_L g4134 ( 
.A1(n_3978),
.A2(n_413),
.B(n_414),
.Y(n_4134)
);

AOI22xp5_ASAP7_75t_L g4135 ( 
.A1(n_3902),
.A2(n_416),
.B1(n_414),
.B2(n_415),
.Y(n_4135)
);

NAND2xp5_ASAP7_75t_L g4136 ( 
.A(n_3913),
.B(n_690),
.Y(n_4136)
);

OAI21x1_ASAP7_75t_L g4137 ( 
.A1(n_3987),
.A2(n_415),
.B(n_417),
.Y(n_4137)
);

BUFx6f_ASAP7_75t_L g4138 ( 
.A(n_3898),
.Y(n_4138)
);

NAND2xp5_ASAP7_75t_L g4139 ( 
.A(n_3930),
.B(n_689),
.Y(n_4139)
);

NAND2xp5_ASAP7_75t_SL g4140 ( 
.A(n_3911),
.B(n_417),
.Y(n_4140)
);

OR2x6_ASAP7_75t_L g4141 ( 
.A(n_3988),
.B(n_418),
.Y(n_4141)
);

CKINVDCx5p33_ASAP7_75t_R g4142 ( 
.A(n_3864),
.Y(n_4142)
);

OAI21x1_ASAP7_75t_L g4143 ( 
.A1(n_4002),
.A2(n_418),
.B(n_419),
.Y(n_4143)
);

BUFx8_ASAP7_75t_L g4144 ( 
.A(n_3860),
.Y(n_4144)
);

BUFx2_ASAP7_75t_R g4145 ( 
.A(n_3979),
.Y(n_4145)
);

BUFx3_ASAP7_75t_L g4146 ( 
.A(n_4007),
.Y(n_4146)
);

NAND2xp5_ASAP7_75t_L g4147 ( 
.A(n_3956),
.B(n_419),
.Y(n_4147)
);

BUFx3_ASAP7_75t_L g4148 ( 
.A(n_4012),
.Y(n_4148)
);

INVx1_ASAP7_75t_L g4149 ( 
.A(n_3936),
.Y(n_4149)
);

AO21x2_ASAP7_75t_L g4150 ( 
.A1(n_3943),
.A2(n_420),
.B(n_421),
.Y(n_4150)
);

INVx3_ASAP7_75t_L g4151 ( 
.A(n_3922),
.Y(n_4151)
);

INVx1_ASAP7_75t_L g4152 ( 
.A(n_3856),
.Y(n_4152)
);

INVx1_ASAP7_75t_L g4153 ( 
.A(n_3856),
.Y(n_4153)
);

OAI21x1_ASAP7_75t_L g4154 ( 
.A1(n_3857),
.A2(n_3974),
.B(n_3984),
.Y(n_4154)
);

CKINVDCx8_ASAP7_75t_R g4155 ( 
.A(n_3905),
.Y(n_4155)
);

AOI21xp5_ASAP7_75t_SL g4156 ( 
.A1(n_3897),
.A2(n_3903),
.B(n_3946),
.Y(n_4156)
);

OA21x2_ASAP7_75t_L g4157 ( 
.A1(n_3867),
.A2(n_420),
.B(n_421),
.Y(n_4157)
);

OAI21x1_ASAP7_75t_L g4158 ( 
.A1(n_3859),
.A2(n_422),
.B(n_423),
.Y(n_4158)
);

A2O1A1Ixp33_ASAP7_75t_L g4159 ( 
.A1(n_3909),
.A2(n_425),
.B(n_422),
.C(n_424),
.Y(n_4159)
);

INVx1_ASAP7_75t_L g4160 ( 
.A(n_3868),
.Y(n_4160)
);

INVx2_ASAP7_75t_L g4161 ( 
.A(n_3922),
.Y(n_4161)
);

AOI222xp33_ASAP7_75t_L g4162 ( 
.A1(n_3990),
.A2(n_3883),
.B1(n_3959),
.B2(n_3940),
.C1(n_3833),
.C2(n_3939),
.Y(n_4162)
);

OAI21x1_ASAP7_75t_L g4163 ( 
.A1(n_3850),
.A2(n_424),
.B(n_425),
.Y(n_4163)
);

A2O1A1Ixp33_ASAP7_75t_L g4164 ( 
.A1(n_3877),
.A2(n_684),
.B(n_428),
.C(n_426),
.Y(n_4164)
);

NAND2xp5_ASAP7_75t_L g4165 ( 
.A(n_4039),
.B(n_3868),
.Y(n_4165)
);

OAI21x1_ASAP7_75t_L g4166 ( 
.A1(n_4151),
.A2(n_3919),
.B(n_3832),
.Y(n_4166)
);

BUFx2_ASAP7_75t_L g4167 ( 
.A(n_4021),
.Y(n_4167)
);

OAI22xp5_ASAP7_75t_L g4168 ( 
.A1(n_4145),
.A2(n_3854),
.B1(n_3924),
.B2(n_3969),
.Y(n_4168)
);

OAI21x1_ASAP7_75t_L g4169 ( 
.A1(n_4151),
.A2(n_3912),
.B(n_3896),
.Y(n_4169)
);

INVx1_ASAP7_75t_L g4170 ( 
.A(n_4025),
.Y(n_4170)
);

OR2x2_ASAP7_75t_L g4171 ( 
.A(n_4041),
.B(n_3874),
.Y(n_4171)
);

INVx1_ASAP7_75t_L g4172 ( 
.A(n_4025),
.Y(n_4172)
);

AOI21xp5_ASAP7_75t_L g4173 ( 
.A1(n_4156),
.A2(n_3983),
.B(n_3889),
.Y(n_4173)
);

INVx2_ASAP7_75t_L g4174 ( 
.A(n_4022),
.Y(n_4174)
);

INVx1_ASAP7_75t_L g4175 ( 
.A(n_4045),
.Y(n_4175)
);

CKINVDCx20_ASAP7_75t_R g4176 ( 
.A(n_4051),
.Y(n_4176)
);

INVx2_ASAP7_75t_L g4177 ( 
.A(n_4022),
.Y(n_4177)
);

INVx2_ASAP7_75t_L g4178 ( 
.A(n_4062),
.Y(n_4178)
);

NAND2xp5_ASAP7_75t_L g4179 ( 
.A(n_4100),
.B(n_3874),
.Y(n_4179)
);

INVx2_ASAP7_75t_SL g4180 ( 
.A(n_4055),
.Y(n_4180)
);

INVx1_ASAP7_75t_L g4181 ( 
.A(n_4045),
.Y(n_4181)
);

A2O1A1Ixp33_ASAP7_75t_L g4182 ( 
.A1(n_4124),
.A2(n_3961),
.B(n_3986),
.C(n_4005),
.Y(n_4182)
);

AOI21xp33_ASAP7_75t_L g4183 ( 
.A1(n_4162),
.A2(n_3998),
.B(n_3921),
.Y(n_4183)
);

BUFx8_ASAP7_75t_SL g4184 ( 
.A(n_4055),
.Y(n_4184)
);

NAND2xp5_ASAP7_75t_L g4185 ( 
.A(n_4100),
.B(n_3893),
.Y(n_4185)
);

NOR2x1_ASAP7_75t_SL g4186 ( 
.A(n_4024),
.B(n_3999),
.Y(n_4186)
);

BUFx8_ASAP7_75t_SL g4187 ( 
.A(n_4126),
.Y(n_4187)
);

INVx1_ASAP7_75t_L g4188 ( 
.A(n_4057),
.Y(n_4188)
);

NAND2xp5_ASAP7_75t_L g4189 ( 
.A(n_4031),
.B(n_3938),
.Y(n_4189)
);

INVx1_ASAP7_75t_L g4190 ( 
.A(n_4057),
.Y(n_4190)
);

INVx1_ASAP7_75t_L g4191 ( 
.A(n_4046),
.Y(n_4191)
);

INVx3_ASAP7_75t_L g4192 ( 
.A(n_4052),
.Y(n_4192)
);

AOI22xp5_ASAP7_75t_L g4193 ( 
.A1(n_4122),
.A2(n_3947),
.B1(n_4001),
.B2(n_3981),
.Y(n_4193)
);

BUFx4f_ASAP7_75t_L g4194 ( 
.A(n_4127),
.Y(n_4194)
);

NAND2xp5_ASAP7_75t_L g4195 ( 
.A(n_4031),
.B(n_3938),
.Y(n_4195)
);

AOI22xp33_ASAP7_75t_L g4196 ( 
.A1(n_4115),
.A2(n_4009),
.B1(n_3840),
.B2(n_3910),
.Y(n_4196)
);

AOI22xp33_ASAP7_75t_L g4197 ( 
.A1(n_4115),
.A2(n_3840),
.B1(n_3910),
.B2(n_3917),
.Y(n_4197)
);

OAI21x1_ASAP7_75t_L g4198 ( 
.A1(n_4061),
.A2(n_3932),
.B(n_3980),
.Y(n_4198)
);

OA21x2_ASAP7_75t_L g4199 ( 
.A1(n_4047),
.A2(n_3840),
.B(n_3893),
.Y(n_4199)
);

OAI21xp5_ASAP7_75t_L g4200 ( 
.A1(n_4118),
.A2(n_3966),
.B(n_4000),
.Y(n_4200)
);

AND2x2_ASAP7_75t_L g4201 ( 
.A(n_4080),
.B(n_3932),
.Y(n_4201)
);

INVx2_ASAP7_75t_L g4202 ( 
.A(n_4062),
.Y(n_4202)
);

OAI21x1_ASAP7_75t_L g4203 ( 
.A1(n_4060),
.A2(n_4032),
.B(n_4038),
.Y(n_4203)
);

OAI21xp5_ASAP7_75t_L g4204 ( 
.A1(n_4154),
.A2(n_3966),
.B(n_4000),
.Y(n_4204)
);

INVx1_ASAP7_75t_L g4205 ( 
.A(n_4049),
.Y(n_4205)
);

AOI22xp33_ASAP7_75t_L g4206 ( 
.A1(n_4157),
.A2(n_4108),
.B1(n_4102),
.B2(n_4097),
.Y(n_4206)
);

OAI21x1_ASAP7_75t_L g4207 ( 
.A1(n_4064),
.A2(n_3980),
.B(n_3996),
.Y(n_4207)
);

OAI21x1_ASAP7_75t_L g4208 ( 
.A1(n_4077),
.A2(n_3996),
.B(n_427),
.Y(n_4208)
);

OAI21x1_ASAP7_75t_L g4209 ( 
.A1(n_4161),
.A2(n_427),
.B(n_428),
.Y(n_4209)
);

INVx1_ASAP7_75t_L g4210 ( 
.A(n_4059),
.Y(n_4210)
);

AO21x2_ASAP7_75t_L g4211 ( 
.A1(n_4071),
.A2(n_429),
.B(n_430),
.Y(n_4211)
);

AOI21xp5_ASAP7_75t_L g4212 ( 
.A1(n_4164),
.A2(n_681),
.B(n_429),
.Y(n_4212)
);

INVx1_ASAP7_75t_L g4213 ( 
.A(n_4059),
.Y(n_4213)
);

INVx1_ASAP7_75t_SL g4214 ( 
.A(n_4133),
.Y(n_4214)
);

NAND2xp5_ASAP7_75t_L g4215 ( 
.A(n_4101),
.B(n_430),
.Y(n_4215)
);

AOI21xp5_ASAP7_75t_L g4216 ( 
.A1(n_4074),
.A2(n_4098),
.B(n_4159),
.Y(n_4216)
);

INVx3_ASAP7_75t_SL g4217 ( 
.A(n_4058),
.Y(n_4217)
);

INVx1_ASAP7_75t_L g4218 ( 
.A(n_4034),
.Y(n_4218)
);

INVx1_ASAP7_75t_L g4219 ( 
.A(n_4037),
.Y(n_4219)
);

AO21x2_ASAP7_75t_L g4220 ( 
.A1(n_4066),
.A2(n_431),
.B(n_432),
.Y(n_4220)
);

INVx1_ASAP7_75t_L g4221 ( 
.A(n_4029),
.Y(n_4221)
);

NAND2x1p5_ASAP7_75t_L g4222 ( 
.A(n_4069),
.B(n_431),
.Y(n_4222)
);

OAI21x1_ASAP7_75t_L g4223 ( 
.A1(n_4078),
.A2(n_432),
.B(n_433),
.Y(n_4223)
);

INVx2_ASAP7_75t_L g4224 ( 
.A(n_4070),
.Y(n_4224)
);

INVx1_ASAP7_75t_L g4225 ( 
.A(n_4033),
.Y(n_4225)
);

OAI21xp5_ASAP7_75t_L g4226 ( 
.A1(n_4117),
.A2(n_433),
.B(n_434),
.Y(n_4226)
);

NAND2xp5_ASAP7_75t_L g4227 ( 
.A(n_4031),
.B(n_436),
.Y(n_4227)
);

INVx2_ASAP7_75t_L g4228 ( 
.A(n_4070),
.Y(n_4228)
);

AND2x4_ASAP7_75t_L g4229 ( 
.A(n_4075),
.B(n_436),
.Y(n_4229)
);

NOR2xp33_ASAP7_75t_L g4230 ( 
.A(n_4058),
.B(n_438),
.Y(n_4230)
);

NAND2xp5_ASAP7_75t_L g4231 ( 
.A(n_4101),
.B(n_438),
.Y(n_4231)
);

INVx2_ASAP7_75t_SL g4232 ( 
.A(n_4146),
.Y(n_4232)
);

OA21x2_ASAP7_75t_L g4233 ( 
.A1(n_4104),
.A2(n_439),
.B(n_440),
.Y(n_4233)
);

OAI21xp5_ASAP7_75t_L g4234 ( 
.A1(n_4157),
.A2(n_439),
.B(n_440),
.Y(n_4234)
);

AO21x2_ASAP7_75t_L g4235 ( 
.A1(n_4114),
.A2(n_441),
.B(n_442),
.Y(n_4235)
);

NAND2xp5_ASAP7_75t_L g4236 ( 
.A(n_4104),
.B(n_4106),
.Y(n_4236)
);

OR2x2_ASAP7_75t_L g4237 ( 
.A(n_4015),
.B(n_678),
.Y(n_4237)
);

BUFx3_ASAP7_75t_L g4238 ( 
.A(n_4103),
.Y(n_4238)
);

INVx2_ASAP7_75t_SL g4239 ( 
.A(n_4092),
.Y(n_4239)
);

INVx1_ASAP7_75t_L g4240 ( 
.A(n_4043),
.Y(n_4240)
);

OA21x2_ASAP7_75t_L g4241 ( 
.A1(n_4106),
.A2(n_441),
.B(n_443),
.Y(n_4241)
);

NAND2xp5_ASAP7_75t_L g4242 ( 
.A(n_4081),
.B(n_444),
.Y(n_4242)
);

INVx1_ASAP7_75t_L g4243 ( 
.A(n_4114),
.Y(n_4243)
);

INVx2_ASAP7_75t_L g4244 ( 
.A(n_4052),
.Y(n_4244)
);

OR2x6_ASAP7_75t_L g4245 ( 
.A(n_4053),
.B(n_444),
.Y(n_4245)
);

INVx2_ASAP7_75t_L g4246 ( 
.A(n_4138),
.Y(n_4246)
);

AO21x2_ASAP7_75t_L g4247 ( 
.A1(n_4149),
.A2(n_445),
.B(n_446),
.Y(n_4247)
);

INVxp67_ASAP7_75t_L g4248 ( 
.A(n_4150),
.Y(n_4248)
);

AOI22xp33_ASAP7_75t_L g4249 ( 
.A1(n_4095),
.A2(n_677),
.B1(n_447),
.B2(n_445),
.Y(n_4249)
);

OAI21x1_ASAP7_75t_L g4250 ( 
.A1(n_4149),
.A2(n_446),
.B(n_448),
.Y(n_4250)
);

OAI21x1_ASAP7_75t_L g4251 ( 
.A1(n_4050),
.A2(n_449),
.B(n_450),
.Y(n_4251)
);

AOI21xp33_ASAP7_75t_L g4252 ( 
.A1(n_4125),
.A2(n_450),
.B(n_451),
.Y(n_4252)
);

INVx1_ASAP7_75t_L g4253 ( 
.A(n_4152),
.Y(n_4253)
);

AO31x2_ASAP7_75t_L g4254 ( 
.A1(n_4152),
.A2(n_453),
.A3(n_451),
.B(n_452),
.Y(n_4254)
);

NAND2xp5_ASAP7_75t_L g4255 ( 
.A(n_4065),
.B(n_452),
.Y(n_4255)
);

AOI22xp33_ASAP7_75t_SL g4256 ( 
.A1(n_4120),
.A2(n_455),
.B1(n_453),
.B2(n_454),
.Y(n_4256)
);

INVx1_ASAP7_75t_L g4257 ( 
.A(n_4153),
.Y(n_4257)
);

AOI21xp5_ASAP7_75t_L g4258 ( 
.A1(n_4073),
.A2(n_677),
.B(n_455),
.Y(n_4258)
);

INVx1_ASAP7_75t_L g4259 ( 
.A(n_4153),
.Y(n_4259)
);

AOI21xp5_ASAP7_75t_L g4260 ( 
.A1(n_4016),
.A2(n_676),
.B(n_456),
.Y(n_4260)
);

AO21x2_ASAP7_75t_L g4261 ( 
.A1(n_4160),
.A2(n_456),
.B(n_457),
.Y(n_4261)
);

AOI21xp5_ASAP7_75t_L g4262 ( 
.A1(n_4054),
.A2(n_457),
.B(n_458),
.Y(n_4262)
);

AOI21x1_ASAP7_75t_L g4263 ( 
.A1(n_4014),
.A2(n_458),
.B(n_459),
.Y(n_4263)
);

OAI21x1_ASAP7_75t_L g4264 ( 
.A1(n_4160),
.A2(n_459),
.B(n_460),
.Y(n_4264)
);

AO31x2_ASAP7_75t_L g4265 ( 
.A1(n_4068),
.A2(n_462),
.A3(n_460),
.B(n_461),
.Y(n_4265)
);

INVx2_ASAP7_75t_L g4266 ( 
.A(n_4138),
.Y(n_4266)
);

OAI21xp5_ASAP7_75t_L g4267 ( 
.A1(n_4140),
.A2(n_461),
.B(n_463),
.Y(n_4267)
);

INVx2_ASAP7_75t_L g4268 ( 
.A(n_4138),
.Y(n_4268)
);

AOI21xp5_ASAP7_75t_L g4269 ( 
.A1(n_4079),
.A2(n_463),
.B(n_464),
.Y(n_4269)
);

OA21x2_ASAP7_75t_L g4270 ( 
.A1(n_4019),
.A2(n_464),
.B(n_465),
.Y(n_4270)
);

INVx2_ASAP7_75t_L g4271 ( 
.A(n_4075),
.Y(n_4271)
);

INVx1_ASAP7_75t_L g4272 ( 
.A(n_4076),
.Y(n_4272)
);

INVx1_ASAP7_75t_L g4273 ( 
.A(n_4076),
.Y(n_4273)
);

INVx1_ASAP7_75t_L g4274 ( 
.A(n_4067),
.Y(n_4274)
);

NAND2x1p5_ASAP7_75t_L g4275 ( 
.A(n_4094),
.B(n_465),
.Y(n_4275)
);

NAND2x1p5_ASAP7_75t_L g4276 ( 
.A(n_4132),
.B(n_466),
.Y(n_4276)
);

NAND2xp5_ASAP7_75t_L g4277 ( 
.A(n_4036),
.B(n_466),
.Y(n_4277)
);

INVx1_ASAP7_75t_L g4278 ( 
.A(n_4067),
.Y(n_4278)
);

INVx2_ASAP7_75t_L g4279 ( 
.A(n_4111),
.Y(n_4279)
);

OAI21xp5_ASAP7_75t_L g4280 ( 
.A1(n_4143),
.A2(n_468),
.B(n_469),
.Y(n_4280)
);

CKINVDCx20_ASAP7_75t_R g4281 ( 
.A(n_4142),
.Y(n_4281)
);

INVx2_ASAP7_75t_SL g4282 ( 
.A(n_4085),
.Y(n_4282)
);

OR2x6_ASAP7_75t_L g4283 ( 
.A(n_4053),
.B(n_4018),
.Y(n_4283)
);

OR2x2_ASAP7_75t_L g4284 ( 
.A(n_4036),
.B(n_468),
.Y(n_4284)
);

NAND2xp5_ASAP7_75t_L g4285 ( 
.A(n_4028),
.B(n_469),
.Y(n_4285)
);

AOI21xp5_ASAP7_75t_L g4286 ( 
.A1(n_4107),
.A2(n_470),
.B(n_471),
.Y(n_4286)
);

INVx1_ASAP7_75t_L g4287 ( 
.A(n_4017),
.Y(n_4287)
);

OA21x2_ASAP7_75t_L g4288 ( 
.A1(n_4056),
.A2(n_471),
.B(n_472),
.Y(n_4288)
);

OA21x2_ASAP7_75t_L g4289 ( 
.A1(n_4035),
.A2(n_472),
.B(n_473),
.Y(n_4289)
);

NAND2xp5_ASAP7_75t_L g4290 ( 
.A(n_4017),
.B(n_474),
.Y(n_4290)
);

INVx1_ASAP7_75t_L g4291 ( 
.A(n_4017),
.Y(n_4291)
);

INVx1_ASAP7_75t_L g4292 ( 
.A(n_4128),
.Y(n_4292)
);

NAND2xp5_ASAP7_75t_L g4293 ( 
.A(n_4148),
.B(n_474),
.Y(n_4293)
);

BUFx3_ASAP7_75t_L g4294 ( 
.A(n_4113),
.Y(n_4294)
);

INVx4_ASAP7_75t_L g4295 ( 
.A(n_4141),
.Y(n_4295)
);

INVx1_ASAP7_75t_L g4296 ( 
.A(n_4026),
.Y(n_4296)
);

INVx2_ASAP7_75t_L g4297 ( 
.A(n_4084),
.Y(n_4297)
);

AOI22xp33_ASAP7_75t_L g4298 ( 
.A1(n_4095),
.A2(n_676),
.B1(n_477),
.B2(n_475),
.Y(n_4298)
);

OR2x6_ASAP7_75t_L g4299 ( 
.A(n_4018),
.B(n_475),
.Y(n_4299)
);

OAI21x1_ASAP7_75t_L g4300 ( 
.A1(n_4042),
.A2(n_476),
.B(n_477),
.Y(n_4300)
);

OAI211xp5_ASAP7_75t_L g4301 ( 
.A1(n_4093),
.A2(n_479),
.B(n_476),
.C(n_478),
.Y(n_4301)
);

OR2x2_ASAP7_75t_L g4302 ( 
.A(n_4110),
.B(n_675),
.Y(n_4302)
);

NAND2xp5_ASAP7_75t_L g4303 ( 
.A(n_4133),
.B(n_478),
.Y(n_4303)
);

AOI22xp33_ASAP7_75t_L g4304 ( 
.A1(n_4087),
.A2(n_674),
.B1(n_481),
.B2(n_479),
.Y(n_4304)
);

INVx5_ASAP7_75t_L g4305 ( 
.A(n_4141),
.Y(n_4305)
);

OA21x2_ASAP7_75t_L g4306 ( 
.A1(n_4099),
.A2(n_480),
.B(n_481),
.Y(n_4306)
);

AO21x2_ASAP7_75t_L g4307 ( 
.A1(n_4096),
.A2(n_482),
.B(n_483),
.Y(n_4307)
);

OA21x2_ASAP7_75t_L g4308 ( 
.A1(n_4105),
.A2(n_482),
.B(n_484),
.Y(n_4308)
);

OAI21x1_ASAP7_75t_L g4309 ( 
.A1(n_4089),
.A2(n_4013),
.B(n_4086),
.Y(n_4309)
);

INVx1_ASAP7_75t_SL g4310 ( 
.A(n_4091),
.Y(n_4310)
);

AOI21x1_ASAP7_75t_L g4311 ( 
.A1(n_4129),
.A2(n_484),
.B(n_486),
.Y(n_4311)
);

INVx2_ASAP7_75t_L g4312 ( 
.A(n_4084),
.Y(n_4312)
);

OR2x2_ASAP7_75t_L g4313 ( 
.A(n_4110),
.B(n_4119),
.Y(n_4313)
);

OAI22xp5_ASAP7_75t_L g4314 ( 
.A1(n_4206),
.A2(n_4023),
.B1(n_4082),
.B2(n_4135),
.Y(n_4314)
);

BUFx2_ASAP7_75t_L g4315 ( 
.A(n_4283),
.Y(n_4315)
);

INVx1_ASAP7_75t_L g4316 ( 
.A(n_4243),
.Y(n_4316)
);

INVx2_ASAP7_75t_L g4317 ( 
.A(n_4192),
.Y(n_4317)
);

INVx1_ASAP7_75t_L g4318 ( 
.A(n_4170),
.Y(n_4318)
);

AOI22xp33_ASAP7_75t_L g4319 ( 
.A1(n_4183),
.A2(n_4082),
.B1(n_4123),
.B2(n_4130),
.Y(n_4319)
);

AOI22xp33_ASAP7_75t_L g4320 ( 
.A1(n_4183),
.A2(n_4216),
.B1(n_4168),
.B2(n_4260),
.Y(n_4320)
);

OAI21xp33_ASAP7_75t_L g4321 ( 
.A1(n_4196),
.A2(n_4112),
.B(n_4044),
.Y(n_4321)
);

INVx1_ASAP7_75t_L g4322 ( 
.A(n_4172),
.Y(n_4322)
);

AOI22xp33_ASAP7_75t_L g4323 ( 
.A1(n_4168),
.A2(n_4130),
.B1(n_4091),
.B2(n_4084),
.Y(n_4323)
);

INVx1_ASAP7_75t_L g4324 ( 
.A(n_4253),
.Y(n_4324)
);

NAND2xp5_ASAP7_75t_L g4325 ( 
.A(n_4214),
.B(n_4110),
.Y(n_4325)
);

OAI22xp5_ASAP7_75t_SL g4326 ( 
.A1(n_4305),
.A2(n_4155),
.B1(n_4126),
.B2(n_4020),
.Y(n_4326)
);

OAI222xp33_ASAP7_75t_L g4327 ( 
.A1(n_4173),
.A2(n_4136),
.B1(n_4139),
.B2(n_4147),
.C1(n_4083),
.C2(n_4040),
.Y(n_4327)
);

AOI22xp33_ASAP7_75t_L g4328 ( 
.A1(n_4262),
.A2(n_4130),
.B1(n_4158),
.B2(n_4030),
.Y(n_4328)
);

AOI22xp33_ASAP7_75t_L g4329 ( 
.A1(n_4285),
.A2(n_4130),
.B1(n_4137),
.B2(n_4121),
.Y(n_4329)
);

OAI22xp5_ASAP7_75t_L g4330 ( 
.A1(n_4197),
.A2(n_4048),
.B1(n_4089),
.B2(n_4083),
.Y(n_4330)
);

BUFx12f_ASAP7_75t_L g4331 ( 
.A(n_4245),
.Y(n_4331)
);

AOI22xp33_ASAP7_75t_L g4332 ( 
.A1(n_4212),
.A2(n_4144),
.B1(n_4063),
.B2(n_4088),
.Y(n_4332)
);

CKINVDCx14_ASAP7_75t_R g4333 ( 
.A(n_4176),
.Y(n_4333)
);

OR2x2_ASAP7_75t_L g4334 ( 
.A(n_4236),
.B(n_4131),
.Y(n_4334)
);

INVx1_ASAP7_75t_L g4335 ( 
.A(n_4257),
.Y(n_4335)
);

INVx5_ASAP7_75t_SL g4336 ( 
.A(n_4245),
.Y(n_4336)
);

NAND2xp5_ASAP7_75t_L g4337 ( 
.A(n_4214),
.B(n_4134),
.Y(n_4337)
);

INVx1_ASAP7_75t_L g4338 ( 
.A(n_4259),
.Y(n_4338)
);

AOI22xp33_ASAP7_75t_L g4339 ( 
.A1(n_4252),
.A2(n_4144),
.B1(n_4090),
.B2(n_4163),
.Y(n_4339)
);

AOI22xp33_ASAP7_75t_SL g4340 ( 
.A1(n_4186),
.A2(n_4109),
.B1(n_4116),
.B2(n_4072),
.Y(n_4340)
);

BUFx2_ASAP7_75t_L g4341 ( 
.A(n_4283),
.Y(n_4341)
);

AOI22xp33_ASAP7_75t_L g4342 ( 
.A1(n_4252),
.A2(n_4072),
.B1(n_4027),
.B2(n_4109),
.Y(n_4342)
);

AOI22xp33_ASAP7_75t_SL g4343 ( 
.A1(n_4305),
.A2(n_4109),
.B1(n_4072),
.B2(n_4027),
.Y(n_4343)
);

HB1xp67_ASAP7_75t_L g4344 ( 
.A(n_4167),
.Y(n_4344)
);

INVx2_ASAP7_75t_L g4345 ( 
.A(n_4192),
.Y(n_4345)
);

OAI22xp33_ASAP7_75t_L g4346 ( 
.A1(n_4305),
.A2(n_4283),
.B1(n_4193),
.B2(n_4299),
.Y(n_4346)
);

OAI22xp33_ASAP7_75t_L g4347 ( 
.A1(n_4193),
.A2(n_4027),
.B1(n_487),
.B2(n_488),
.Y(n_4347)
);

AOI22xp33_ASAP7_75t_L g4348 ( 
.A1(n_4288),
.A2(n_486),
.B1(n_488),
.B2(n_489),
.Y(n_4348)
);

AOI22xp33_ASAP7_75t_L g4349 ( 
.A1(n_4288),
.A2(n_4226),
.B1(n_4295),
.B2(n_4200),
.Y(n_4349)
);

INVxp67_ASAP7_75t_L g4350 ( 
.A(n_4313),
.Y(n_4350)
);

AOI22xp33_ASAP7_75t_L g4351 ( 
.A1(n_4226),
.A2(n_489),
.B1(n_490),
.B2(n_491),
.Y(n_4351)
);

INVxp67_ASAP7_75t_L g4352 ( 
.A(n_4179),
.Y(n_4352)
);

INVx1_ASAP7_75t_L g4353 ( 
.A(n_4175),
.Y(n_4353)
);

NAND2xp5_ASAP7_75t_L g4354 ( 
.A(n_4248),
.B(n_490),
.Y(n_4354)
);

BUFx12f_ASAP7_75t_L g4355 ( 
.A(n_4245),
.Y(n_4355)
);

AOI22xp33_ASAP7_75t_SL g4356 ( 
.A1(n_4295),
.A2(n_491),
.B1(n_492),
.B2(n_493),
.Y(n_4356)
);

BUFx4f_ASAP7_75t_SL g4357 ( 
.A(n_4281),
.Y(n_4357)
);

AOI22xp5_ASAP7_75t_L g4358 ( 
.A1(n_4310),
.A2(n_493),
.B1(n_494),
.B2(n_495),
.Y(n_4358)
);

AOI22xp33_ASAP7_75t_L g4359 ( 
.A1(n_4200),
.A2(n_494),
.B1(n_496),
.B2(n_497),
.Y(n_4359)
);

OAI22xp5_ASAP7_75t_L g4360 ( 
.A1(n_4310),
.A2(n_4302),
.B1(n_4299),
.B2(n_4194),
.Y(n_4360)
);

OAI21xp5_ASAP7_75t_SL g4361 ( 
.A1(n_4256),
.A2(n_496),
.B(n_498),
.Y(n_4361)
);

AOI22xp33_ASAP7_75t_L g4362 ( 
.A1(n_4204),
.A2(n_498),
.B1(n_499),
.B2(n_500),
.Y(n_4362)
);

OR2x2_ASAP7_75t_L g4363 ( 
.A(n_4179),
.B(n_4185),
.Y(n_4363)
);

HB1xp67_ASAP7_75t_L g4364 ( 
.A(n_4270),
.Y(n_4364)
);

OAI22xp33_ASAP7_75t_SL g4365 ( 
.A1(n_4290),
.A2(n_499),
.B1(n_500),
.B2(n_501),
.Y(n_4365)
);

AOI22xp33_ASAP7_75t_L g4366 ( 
.A1(n_4204),
.A2(n_501),
.B1(n_502),
.B2(n_503),
.Y(n_4366)
);

BUFx5_ASAP7_75t_L g4367 ( 
.A(n_4229),
.Y(n_4367)
);

AOI22xp33_ASAP7_75t_L g4368 ( 
.A1(n_4234),
.A2(n_502),
.B1(n_503),
.B2(n_504),
.Y(n_4368)
);

INVx1_ASAP7_75t_L g4369 ( 
.A(n_4181),
.Y(n_4369)
);

INVx1_ASAP7_75t_L g4370 ( 
.A(n_4188),
.Y(n_4370)
);

AOI222xp33_ASAP7_75t_L g4371 ( 
.A1(n_4182),
.A2(n_504),
.B1(n_505),
.B2(n_506),
.C1(n_507),
.C2(n_508),
.Y(n_4371)
);

AOI22xp33_ASAP7_75t_L g4372 ( 
.A1(n_4234),
.A2(n_505),
.B1(n_506),
.B2(n_507),
.Y(n_4372)
);

AOI22xp33_ASAP7_75t_L g4373 ( 
.A1(n_4258),
.A2(n_509),
.B1(n_510),
.B2(n_511),
.Y(n_4373)
);

AOI22xp33_ASAP7_75t_L g4374 ( 
.A1(n_4220),
.A2(n_509),
.B1(n_510),
.B2(n_511),
.Y(n_4374)
);

INVx2_ASAP7_75t_L g4375 ( 
.A(n_4297),
.Y(n_4375)
);

INVx1_ASAP7_75t_L g4376 ( 
.A(n_4190),
.Y(n_4376)
);

AOI22xp33_ASAP7_75t_L g4377 ( 
.A1(n_4220),
.A2(n_512),
.B1(n_513),
.B2(n_514),
.Y(n_4377)
);

OAI22xp5_ASAP7_75t_L g4378 ( 
.A1(n_4299),
.A2(n_512),
.B1(n_513),
.B2(n_515),
.Y(n_4378)
);

AOI22xp33_ASAP7_75t_L g4379 ( 
.A1(n_4296),
.A2(n_516),
.B1(n_517),
.B2(n_518),
.Y(n_4379)
);

INVx1_ASAP7_75t_L g4380 ( 
.A(n_4284),
.Y(n_4380)
);

AND2x2_ASAP7_75t_L g4381 ( 
.A(n_4246),
.B(n_4266),
.Y(n_4381)
);

NAND2xp5_ASAP7_75t_L g4382 ( 
.A(n_4227),
.B(n_517),
.Y(n_4382)
);

INVx1_ASAP7_75t_L g4383 ( 
.A(n_4210),
.Y(n_4383)
);

OAI22xp5_ASAP7_75t_L g4384 ( 
.A1(n_4194),
.A2(n_518),
.B1(n_519),
.B2(n_520),
.Y(n_4384)
);

BUFx2_ASAP7_75t_L g4385 ( 
.A(n_4217),
.Y(n_4385)
);

AOI222xp33_ASAP7_75t_L g4386 ( 
.A1(n_4267),
.A2(n_519),
.B1(n_520),
.B2(n_521),
.C1(n_522),
.C2(n_523),
.Y(n_4386)
);

AOI22xp33_ASAP7_75t_SL g4387 ( 
.A1(n_4169),
.A2(n_521),
.B1(n_522),
.B2(n_523),
.Y(n_4387)
);

INVx1_ASAP7_75t_L g4388 ( 
.A(n_4213),
.Y(n_4388)
);

BUFx4f_ASAP7_75t_SL g4389 ( 
.A(n_4180),
.Y(n_4389)
);

INVx2_ASAP7_75t_L g4390 ( 
.A(n_4312),
.Y(n_4390)
);

INVx1_ASAP7_75t_L g4391 ( 
.A(n_4178),
.Y(n_4391)
);

CKINVDCx5p33_ASAP7_75t_R g4392 ( 
.A(n_4184),
.Y(n_4392)
);

NAND2xp5_ASAP7_75t_L g4393 ( 
.A(n_4290),
.B(n_524),
.Y(n_4393)
);

AOI222xp33_ASAP7_75t_L g4394 ( 
.A1(n_4267),
.A2(n_524),
.B1(n_525),
.B2(n_526),
.C1(n_528),
.C2(n_529),
.Y(n_4394)
);

AOI22xp33_ASAP7_75t_SL g4395 ( 
.A1(n_4301),
.A2(n_525),
.B1(n_526),
.B2(n_528),
.Y(n_4395)
);

OAI21xp33_ASAP7_75t_L g4396 ( 
.A1(n_4165),
.A2(n_529),
.B(n_531),
.Y(n_4396)
);

INVx1_ASAP7_75t_L g4397 ( 
.A(n_4202),
.Y(n_4397)
);

INVx1_ASAP7_75t_L g4398 ( 
.A(n_4224),
.Y(n_4398)
);

CKINVDCx5p33_ASAP7_75t_R g4399 ( 
.A(n_4238),
.Y(n_4399)
);

INVx1_ASAP7_75t_L g4400 ( 
.A(n_4228),
.Y(n_4400)
);

NAND2x1p5_ASAP7_75t_L g4401 ( 
.A(n_4270),
.B(n_531),
.Y(n_4401)
);

OAI22xp5_ASAP7_75t_L g4402 ( 
.A1(n_4303),
.A2(n_4298),
.B1(n_4249),
.B2(n_4268),
.Y(n_4402)
);

INVx2_ASAP7_75t_SL g4403 ( 
.A(n_4294),
.Y(n_4403)
);

AOI211xp5_ASAP7_75t_SL g4404 ( 
.A1(n_4286),
.A2(n_532),
.B(n_533),
.C(n_534),
.Y(n_4404)
);

OAI21xp5_ASAP7_75t_SL g4405 ( 
.A1(n_4304),
.A2(n_532),
.B(n_533),
.Y(n_4405)
);

BUFx12f_ASAP7_75t_L g4406 ( 
.A(n_4275),
.Y(n_4406)
);

HB1xp67_ASAP7_75t_L g4407 ( 
.A(n_4201),
.Y(n_4407)
);

HB1xp67_ASAP7_75t_L g4408 ( 
.A(n_4289),
.Y(n_4408)
);

OAI222xp33_ASAP7_75t_L g4409 ( 
.A1(n_4303),
.A2(n_4277),
.B1(n_4165),
.B2(n_4185),
.C1(n_4276),
.C2(n_4215),
.Y(n_4409)
);

AOI222xp33_ASAP7_75t_L g4410 ( 
.A1(n_4230),
.A2(n_534),
.B1(n_535),
.B2(n_536),
.C1(n_537),
.C2(n_538),
.Y(n_4410)
);

AOI22xp33_ASAP7_75t_SL g4411 ( 
.A1(n_4166),
.A2(n_535),
.B1(n_537),
.B2(n_540),
.Y(n_4411)
);

OAI22xp5_ASAP7_75t_L g4412 ( 
.A1(n_4277),
.A2(n_540),
.B1(n_541),
.B2(n_542),
.Y(n_4412)
);

AOI22xp33_ASAP7_75t_SL g4413 ( 
.A1(n_4233),
.A2(n_674),
.B1(n_542),
.B2(n_543),
.Y(n_4413)
);

INVx3_ASAP7_75t_L g4414 ( 
.A(n_4229),
.Y(n_4414)
);

BUFx4f_ASAP7_75t_SL g4415 ( 
.A(n_4232),
.Y(n_4415)
);

AOI22xp5_ASAP7_75t_L g4416 ( 
.A1(n_4211),
.A2(n_541),
.B1(n_543),
.B2(n_544),
.Y(n_4416)
);

OAI21xp5_ASAP7_75t_SL g4417 ( 
.A1(n_4280),
.A2(n_544),
.B(n_545),
.Y(n_4417)
);

OAI22xp5_ASAP7_75t_SL g4418 ( 
.A1(n_4222),
.A2(n_546),
.B1(n_548),
.B2(n_549),
.Y(n_4418)
);

INVx2_ASAP7_75t_L g4419 ( 
.A(n_4244),
.Y(n_4419)
);

AOI22xp33_ASAP7_75t_L g4420 ( 
.A1(n_4211),
.A2(n_550),
.B1(n_551),
.B2(n_552),
.Y(n_4420)
);

OAI22xp33_ASAP7_75t_L g4421 ( 
.A1(n_4241),
.A2(n_551),
.B1(n_552),
.B2(n_553),
.Y(n_4421)
);

NAND2xp5_ASAP7_75t_L g4422 ( 
.A(n_4219),
.B(n_553),
.Y(n_4422)
);

AOI22xp33_ASAP7_75t_L g4423 ( 
.A1(n_4280),
.A2(n_555),
.B1(n_556),
.B2(n_557),
.Y(n_4423)
);

INVx2_ASAP7_75t_L g4424 ( 
.A(n_4271),
.Y(n_4424)
);

AOI22xp33_ASAP7_75t_SL g4425 ( 
.A1(n_4241),
.A2(n_556),
.B1(n_558),
.B2(n_559),
.Y(n_4425)
);

INVx2_ASAP7_75t_SL g4426 ( 
.A(n_4239),
.Y(n_4426)
);

AOI22xp33_ASAP7_75t_SL g4427 ( 
.A1(n_4261),
.A2(n_558),
.B1(n_560),
.B2(n_561),
.Y(n_4427)
);

BUFx4f_ASAP7_75t_SL g4428 ( 
.A(n_4282),
.Y(n_4428)
);

OAI21xp33_ASAP7_75t_L g4429 ( 
.A1(n_4189),
.A2(n_561),
.B(n_562),
.Y(n_4429)
);

AOI22xp33_ASAP7_75t_L g4430 ( 
.A1(n_4307),
.A2(n_563),
.B1(n_564),
.B2(n_565),
.Y(n_4430)
);

INVx1_ASAP7_75t_L g4431 ( 
.A(n_4191),
.Y(n_4431)
);

INVx2_ASAP7_75t_L g4432 ( 
.A(n_4174),
.Y(n_4432)
);

OAI21xp5_ASAP7_75t_SL g4433 ( 
.A1(n_4269),
.A2(n_563),
.B(n_564),
.Y(n_4433)
);

BUFx2_ASAP7_75t_L g4434 ( 
.A(n_4187),
.Y(n_4434)
);

AND2x2_ASAP7_75t_L g4435 ( 
.A(n_4177),
.B(n_565),
.Y(n_4435)
);

CKINVDCx5p33_ASAP7_75t_R g4436 ( 
.A(n_4242),
.Y(n_4436)
);

INVx1_ASAP7_75t_L g4437 ( 
.A(n_4205),
.Y(n_4437)
);

AOI22xp33_ASAP7_75t_L g4438 ( 
.A1(n_4307),
.A2(n_566),
.B1(n_567),
.B2(n_568),
.Y(n_4438)
);

CKINVDCx16_ASAP7_75t_R g4439 ( 
.A(n_4237),
.Y(n_4439)
);

AOI22xp33_ASAP7_75t_L g4440 ( 
.A1(n_4289),
.A2(n_569),
.B1(n_570),
.B2(n_571),
.Y(n_4440)
);

INVx1_ASAP7_75t_L g4441 ( 
.A(n_4221),
.Y(n_4441)
);

OAI21xp5_ASAP7_75t_L g4442 ( 
.A1(n_4251),
.A2(n_570),
.B(n_572),
.Y(n_4442)
);

AOI22xp33_ASAP7_75t_L g4443 ( 
.A1(n_4309),
.A2(n_572),
.B1(n_573),
.B2(n_574),
.Y(n_4443)
);

INVx5_ASAP7_75t_L g4444 ( 
.A(n_4254),
.Y(n_4444)
);

OAI22xp5_ASAP7_75t_L g4445 ( 
.A1(n_4215),
.A2(n_574),
.B1(n_575),
.B2(n_576),
.Y(n_4445)
);

CKINVDCx11_ASAP7_75t_R g4446 ( 
.A(n_4279),
.Y(n_4446)
);

HB1xp67_ASAP7_75t_L g4447 ( 
.A(n_4195),
.Y(n_4447)
);

OAI22xp5_ASAP7_75t_SL g4448 ( 
.A1(n_4231),
.A2(n_4293),
.B1(n_4199),
.B2(n_4306),
.Y(n_4448)
);

AND2x2_ASAP7_75t_L g4449 ( 
.A(n_4272),
.B(n_576),
.Y(n_4449)
);

HB1xp67_ASAP7_75t_L g4450 ( 
.A(n_4265),
.Y(n_4450)
);

INVx1_ASAP7_75t_L g4451 ( 
.A(n_4225),
.Y(n_4451)
);

OAI22xp5_ASAP7_75t_L g4452 ( 
.A1(n_4199),
.A2(n_577),
.B1(n_578),
.B2(n_579),
.Y(n_4452)
);

AOI22xp33_ASAP7_75t_L g4453 ( 
.A1(n_4261),
.A2(n_577),
.B1(n_578),
.B2(n_580),
.Y(n_4453)
);

AOI22xp5_ASAP7_75t_L g4454 ( 
.A1(n_4235),
.A2(n_580),
.B1(n_581),
.B2(n_582),
.Y(n_4454)
);

INVx2_ASAP7_75t_L g4455 ( 
.A(n_4273),
.Y(n_4455)
);

INVx6_ASAP7_75t_L g4456 ( 
.A(n_4171),
.Y(n_4456)
);

AOI22xp33_ASAP7_75t_L g4457 ( 
.A1(n_4235),
.A2(n_581),
.B1(n_582),
.B2(n_583),
.Y(n_4457)
);

AOI222xp33_ASAP7_75t_L g4458 ( 
.A1(n_4208),
.A2(n_584),
.B1(n_585),
.B2(n_586),
.C1(n_588),
.C2(n_589),
.Y(n_4458)
);

AOI22xp33_ASAP7_75t_L g4459 ( 
.A1(n_4247),
.A2(n_585),
.B1(n_588),
.B2(n_590),
.Y(n_4459)
);

OAI22xp33_ASAP7_75t_L g4460 ( 
.A1(n_4306),
.A2(n_4308),
.B1(n_4311),
.B2(n_4292),
.Y(n_4460)
);

OAI22xp33_ASAP7_75t_L g4461 ( 
.A1(n_4308),
.A2(n_4255),
.B1(n_4218),
.B2(n_4287),
.Y(n_4461)
);

AOI22xp33_ASAP7_75t_L g4462 ( 
.A1(n_4247),
.A2(n_590),
.B1(n_591),
.B2(n_592),
.Y(n_4462)
);

OAI22xp5_ASAP7_75t_L g4463 ( 
.A1(n_4263),
.A2(n_591),
.B1(n_593),
.B2(n_594),
.Y(n_4463)
);

INVx1_ASAP7_75t_L g4464 ( 
.A(n_4318),
.Y(n_4464)
);

INVx1_ASAP7_75t_L g4465 ( 
.A(n_4322),
.Y(n_4465)
);

NAND2xp5_ASAP7_75t_L g4466 ( 
.A(n_4343),
.B(n_4265),
.Y(n_4466)
);

INVx2_ASAP7_75t_L g4467 ( 
.A(n_4367),
.Y(n_4467)
);

INVx5_ASAP7_75t_L g4468 ( 
.A(n_4331),
.Y(n_4468)
);

BUFx6f_ASAP7_75t_L g4469 ( 
.A(n_4355),
.Y(n_4469)
);

BUFx2_ASAP7_75t_L g4470 ( 
.A(n_4385),
.Y(n_4470)
);

OR2x6_ASAP7_75t_L g4471 ( 
.A(n_4315),
.B(n_4223),
.Y(n_4471)
);

NOR2xp33_ASAP7_75t_L g4472 ( 
.A(n_4434),
.B(n_4240),
.Y(n_4472)
);

HB1xp67_ASAP7_75t_L g4473 ( 
.A(n_4344),
.Y(n_4473)
);

INVx1_ASAP7_75t_L g4474 ( 
.A(n_4353),
.Y(n_4474)
);

INVx1_ASAP7_75t_L g4475 ( 
.A(n_4369),
.Y(n_4475)
);

HB1xp67_ASAP7_75t_L g4476 ( 
.A(n_4444),
.Y(n_4476)
);

AND2x2_ASAP7_75t_L g4477 ( 
.A(n_4341),
.B(n_4291),
.Y(n_4477)
);

INVx1_ASAP7_75t_L g4478 ( 
.A(n_4370),
.Y(n_4478)
);

INVx2_ASAP7_75t_L g4479 ( 
.A(n_4367),
.Y(n_4479)
);

NAND3xp33_ASAP7_75t_L g4480 ( 
.A(n_4320),
.B(n_4278),
.C(n_4274),
.Y(n_4480)
);

INVx2_ASAP7_75t_L g4481 ( 
.A(n_4367),
.Y(n_4481)
);

BUFx2_ASAP7_75t_L g4482 ( 
.A(n_4415),
.Y(n_4482)
);

INVx2_ASAP7_75t_L g4483 ( 
.A(n_4367),
.Y(n_4483)
);

INVx2_ASAP7_75t_SL g4484 ( 
.A(n_4414),
.Y(n_4484)
);

INVx1_ASAP7_75t_L g4485 ( 
.A(n_4376),
.Y(n_4485)
);

AND2x2_ASAP7_75t_L g4486 ( 
.A(n_4317),
.B(n_4203),
.Y(n_4486)
);

AND2x2_ASAP7_75t_L g4487 ( 
.A(n_4345),
.B(n_4198),
.Y(n_4487)
);

AO21x2_ASAP7_75t_L g4488 ( 
.A1(n_4364),
.A2(n_4207),
.B(n_4250),
.Y(n_4488)
);

CKINVDCx20_ASAP7_75t_R g4489 ( 
.A(n_4357),
.Y(n_4489)
);

AND2x2_ASAP7_75t_L g4490 ( 
.A(n_4407),
.B(n_4265),
.Y(n_4490)
);

INVx1_ASAP7_75t_L g4491 ( 
.A(n_4316),
.Y(n_4491)
);

HB1xp67_ASAP7_75t_L g4492 ( 
.A(n_4444),
.Y(n_4492)
);

INVx2_ASAP7_75t_L g4493 ( 
.A(n_4367),
.Y(n_4493)
);

CKINVDCx5p33_ASAP7_75t_R g4494 ( 
.A(n_4333),
.Y(n_4494)
);

OAI21x1_ASAP7_75t_L g4495 ( 
.A1(n_4325),
.A2(n_4300),
.B(n_4209),
.Y(n_4495)
);

HB1xp67_ASAP7_75t_L g4496 ( 
.A(n_4444),
.Y(n_4496)
);

NAND2xp5_ASAP7_75t_L g4497 ( 
.A(n_4342),
.B(n_4254),
.Y(n_4497)
);

OR2x2_ASAP7_75t_L g4498 ( 
.A(n_4380),
.B(n_4254),
.Y(n_4498)
);

AND2x2_ASAP7_75t_L g4499 ( 
.A(n_4432),
.B(n_4264),
.Y(n_4499)
);

INVx1_ASAP7_75t_L g4500 ( 
.A(n_4324),
.Y(n_4500)
);

INVx1_ASAP7_75t_L g4501 ( 
.A(n_4335),
.Y(n_4501)
);

BUFx2_ASAP7_75t_L g4502 ( 
.A(n_4414),
.Y(n_4502)
);

INVx2_ASAP7_75t_L g4503 ( 
.A(n_4444),
.Y(n_4503)
);

INVx2_ASAP7_75t_L g4504 ( 
.A(n_4375),
.Y(n_4504)
);

BUFx6f_ASAP7_75t_L g4505 ( 
.A(n_4392),
.Y(n_4505)
);

OR2x2_ASAP7_75t_L g4506 ( 
.A(n_4334),
.B(n_596),
.Y(n_4506)
);

AO21x2_ASAP7_75t_L g4507 ( 
.A1(n_4408),
.A2(n_596),
.B(n_597),
.Y(n_4507)
);

INVx2_ASAP7_75t_SL g4508 ( 
.A(n_4428),
.Y(n_4508)
);

INVx2_ASAP7_75t_L g4509 ( 
.A(n_4390),
.Y(n_4509)
);

INVx2_ASAP7_75t_L g4510 ( 
.A(n_4381),
.Y(n_4510)
);

OR2x2_ASAP7_75t_L g4511 ( 
.A(n_4337),
.B(n_598),
.Y(n_4511)
);

OAI21x1_ASAP7_75t_L g4512 ( 
.A1(n_4330),
.A2(n_598),
.B(n_599),
.Y(n_4512)
);

OA21x2_ASAP7_75t_L g4513 ( 
.A1(n_4321),
.A2(n_599),
.B(n_600),
.Y(n_4513)
);

INVx3_ASAP7_75t_L g4514 ( 
.A(n_4336),
.Y(n_4514)
);

INVx2_ASAP7_75t_L g4515 ( 
.A(n_4401),
.Y(n_4515)
);

INVx2_ASAP7_75t_L g4516 ( 
.A(n_4401),
.Y(n_4516)
);

INVx3_ASAP7_75t_L g4517 ( 
.A(n_4336),
.Y(n_4517)
);

BUFx3_ASAP7_75t_L g4518 ( 
.A(n_4389),
.Y(n_4518)
);

INVx2_ASAP7_75t_L g4519 ( 
.A(n_4456),
.Y(n_4519)
);

AND2x2_ASAP7_75t_L g4520 ( 
.A(n_4340),
.B(n_602),
.Y(n_4520)
);

INVx1_ASAP7_75t_L g4521 ( 
.A(n_4338),
.Y(n_4521)
);

INVx3_ASAP7_75t_L g4522 ( 
.A(n_4336),
.Y(n_4522)
);

INVx1_ASAP7_75t_L g4523 ( 
.A(n_4383),
.Y(n_4523)
);

AND2x2_ASAP7_75t_L g4524 ( 
.A(n_4419),
.B(n_603),
.Y(n_4524)
);

AOI21x1_ASAP7_75t_L g4525 ( 
.A1(n_4360),
.A2(n_4354),
.B(n_4452),
.Y(n_4525)
);

OA21x2_ASAP7_75t_L g4526 ( 
.A1(n_4349),
.A2(n_603),
.B(n_604),
.Y(n_4526)
);

AND2x2_ASAP7_75t_L g4527 ( 
.A(n_4424),
.B(n_604),
.Y(n_4527)
);

INVx2_ASAP7_75t_L g4528 ( 
.A(n_4456),
.Y(n_4528)
);

OR2x6_ASAP7_75t_L g4529 ( 
.A(n_4326),
.B(n_605),
.Y(n_4529)
);

OAI21x1_ASAP7_75t_L g4530 ( 
.A1(n_4330),
.A2(n_605),
.B(n_606),
.Y(n_4530)
);

HB1xp67_ASAP7_75t_L g4531 ( 
.A(n_4450),
.Y(n_4531)
);

AND2x2_ASAP7_75t_L g4532 ( 
.A(n_4455),
.B(n_606),
.Y(n_4532)
);

BUFx3_ASAP7_75t_L g4533 ( 
.A(n_4406),
.Y(n_4533)
);

INVx3_ASAP7_75t_L g4534 ( 
.A(n_4446),
.Y(n_4534)
);

BUFx6f_ASAP7_75t_L g4535 ( 
.A(n_4435),
.Y(n_4535)
);

NOR2xp33_ASAP7_75t_L g4536 ( 
.A(n_4327),
.B(n_4346),
.Y(n_4536)
);

INVx1_ASAP7_75t_L g4537 ( 
.A(n_4388),
.Y(n_4537)
);

INVxp33_ASAP7_75t_L g4538 ( 
.A(n_4448),
.Y(n_4538)
);

INVx1_ASAP7_75t_L g4539 ( 
.A(n_4431),
.Y(n_4539)
);

BUFx2_ASAP7_75t_L g4540 ( 
.A(n_4426),
.Y(n_4540)
);

AO21x2_ASAP7_75t_L g4541 ( 
.A1(n_4461),
.A2(n_610),
.B(n_612),
.Y(n_4541)
);

AND2x2_ASAP7_75t_L g4542 ( 
.A(n_4350),
.B(n_610),
.Y(n_4542)
);

INVx1_ASAP7_75t_L g4543 ( 
.A(n_4437),
.Y(n_4543)
);

INVx1_ASAP7_75t_L g4544 ( 
.A(n_4441),
.Y(n_4544)
);

INVx2_ASAP7_75t_L g4545 ( 
.A(n_4391),
.Y(n_4545)
);

AND2x2_ASAP7_75t_L g4546 ( 
.A(n_4323),
.B(n_612),
.Y(n_4546)
);

AND2x2_ASAP7_75t_L g4547 ( 
.A(n_4352),
.B(n_613),
.Y(n_4547)
);

AND2x2_ASAP7_75t_L g4548 ( 
.A(n_4397),
.B(n_614),
.Y(n_4548)
);

INVx2_ASAP7_75t_L g4549 ( 
.A(n_4398),
.Y(n_4549)
);

INVx1_ASAP7_75t_L g4550 ( 
.A(n_4451),
.Y(n_4550)
);

INVxp67_ASAP7_75t_L g4551 ( 
.A(n_4363),
.Y(n_4551)
);

INVx2_ASAP7_75t_L g4552 ( 
.A(n_4400),
.Y(n_4552)
);

INVx1_ASAP7_75t_L g4553 ( 
.A(n_4422),
.Y(n_4553)
);

HB1xp67_ASAP7_75t_L g4554 ( 
.A(n_4447),
.Y(n_4554)
);

AO21x2_ASAP7_75t_L g4555 ( 
.A1(n_4393),
.A2(n_614),
.B(n_615),
.Y(n_4555)
);

INVx1_ASAP7_75t_L g4556 ( 
.A(n_4382),
.Y(n_4556)
);

INVx2_ASAP7_75t_L g4557 ( 
.A(n_4439),
.Y(n_4557)
);

BUFx4f_ASAP7_75t_SL g4558 ( 
.A(n_4403),
.Y(n_4558)
);

AO21x2_ASAP7_75t_L g4559 ( 
.A1(n_4421),
.A2(n_615),
.B(n_616),
.Y(n_4559)
);

INVx2_ASAP7_75t_L g4560 ( 
.A(n_4449),
.Y(n_4560)
);

AND2x4_ASAP7_75t_L g4561 ( 
.A(n_4442),
.B(n_616),
.Y(n_4561)
);

AND2x2_ASAP7_75t_L g4562 ( 
.A(n_4319),
.B(n_617),
.Y(n_4562)
);

INVx1_ASAP7_75t_L g4563 ( 
.A(n_4460),
.Y(n_4563)
);

HB1xp67_ASAP7_75t_L g4564 ( 
.A(n_4409),
.Y(n_4564)
);

OA21x2_ASAP7_75t_L g4565 ( 
.A1(n_4443),
.A2(n_620),
.B(n_621),
.Y(n_4565)
);

AND2x2_ASAP7_75t_L g4566 ( 
.A(n_4329),
.B(n_622),
.Y(n_4566)
);

NAND2xp5_ASAP7_75t_L g4567 ( 
.A(n_4314),
.B(n_622),
.Y(n_4567)
);

AND2x2_ASAP7_75t_L g4568 ( 
.A(n_4411),
.B(n_4339),
.Y(n_4568)
);

NAND2xp5_ASAP7_75t_L g4569 ( 
.A(n_4387),
.B(n_623),
.Y(n_4569)
);

INVx1_ASAP7_75t_L g4570 ( 
.A(n_4416),
.Y(n_4570)
);

INVx2_ASAP7_75t_L g4571 ( 
.A(n_4436),
.Y(n_4571)
);

INVx1_ASAP7_75t_L g4572 ( 
.A(n_4402),
.Y(n_4572)
);

INVx1_ASAP7_75t_L g4573 ( 
.A(n_4454),
.Y(n_4573)
);

INVx2_ASAP7_75t_SL g4574 ( 
.A(n_4399),
.Y(n_4574)
);

INVx2_ASAP7_75t_SL g4575 ( 
.A(n_4463),
.Y(n_4575)
);

AND2x4_ASAP7_75t_L g4576 ( 
.A(n_4442),
.B(n_623),
.Y(n_4576)
);

OR2x2_ASAP7_75t_L g4577 ( 
.A(n_4332),
.B(n_4328),
.Y(n_4577)
);

INVx2_ASAP7_75t_L g4578 ( 
.A(n_4463),
.Y(n_4578)
);

INVx1_ASAP7_75t_L g4579 ( 
.A(n_4412),
.Y(n_4579)
);

NOR2xp33_ASAP7_75t_L g4580 ( 
.A(n_4365),
.B(n_4417),
.Y(n_4580)
);

INVx1_ASAP7_75t_L g4581 ( 
.A(n_4413),
.Y(n_4581)
);

HB1xp67_ASAP7_75t_L g4582 ( 
.A(n_4445),
.Y(n_4582)
);

INVx2_ASAP7_75t_SL g4583 ( 
.A(n_4384),
.Y(n_4583)
);

AND2x2_ASAP7_75t_L g4584 ( 
.A(n_4348),
.B(n_624),
.Y(n_4584)
);

BUFx2_ASAP7_75t_L g4585 ( 
.A(n_4418),
.Y(n_4585)
);

AND2x2_ASAP7_75t_L g4586 ( 
.A(n_4425),
.B(n_625),
.Y(n_4586)
);

NOR2x1_ASAP7_75t_SL g4587 ( 
.A(n_4378),
.B(n_626),
.Y(n_4587)
);

AO21x2_ASAP7_75t_L g4588 ( 
.A1(n_4347),
.A2(n_626),
.B(n_627),
.Y(n_4588)
);

AND2x2_ASAP7_75t_L g4589 ( 
.A(n_4440),
.B(n_627),
.Y(n_4589)
);

AOI21x1_ASAP7_75t_L g4590 ( 
.A1(n_4427),
.A2(n_4404),
.B(n_4396),
.Y(n_4590)
);

AO21x2_ASAP7_75t_L g4591 ( 
.A1(n_4358),
.A2(n_628),
.B(n_629),
.Y(n_4591)
);

INVx1_ASAP7_75t_L g4592 ( 
.A(n_4429),
.Y(n_4592)
);

AND2x4_ASAP7_75t_L g4593 ( 
.A(n_4374),
.B(n_630),
.Y(n_4593)
);

INVx1_ASAP7_75t_L g4594 ( 
.A(n_4458),
.Y(n_4594)
);

OR2x2_ASAP7_75t_L g4595 ( 
.A(n_4433),
.B(n_4377),
.Y(n_4595)
);

INVx2_ASAP7_75t_L g4596 ( 
.A(n_4371),
.Y(n_4596)
);

AND2x2_ASAP7_75t_L g4597 ( 
.A(n_4404),
.B(n_631),
.Y(n_4597)
);

INVx1_ASAP7_75t_L g4598 ( 
.A(n_4458),
.Y(n_4598)
);

AND2x4_ASAP7_75t_SL g4599 ( 
.A(n_4420),
.B(n_632),
.Y(n_4599)
);

INVx2_ASAP7_75t_L g4600 ( 
.A(n_4371),
.Y(n_4600)
);

AND2x2_ASAP7_75t_L g4601 ( 
.A(n_4557),
.B(n_4430),
.Y(n_4601)
);

INVx2_ASAP7_75t_L g4602 ( 
.A(n_4470),
.Y(n_4602)
);

INVx1_ASAP7_75t_L g4603 ( 
.A(n_4507),
.Y(n_4603)
);

INVx2_ASAP7_75t_L g4604 ( 
.A(n_4557),
.Y(n_4604)
);

OR2x2_ASAP7_75t_L g4605 ( 
.A(n_4575),
.B(n_4453),
.Y(n_4605)
);

INVx1_ASAP7_75t_L g4606 ( 
.A(n_4507),
.Y(n_4606)
);

INVx2_ASAP7_75t_SL g4607 ( 
.A(n_4534),
.Y(n_4607)
);

INVx2_ASAP7_75t_L g4608 ( 
.A(n_4502),
.Y(n_4608)
);

AND2x2_ASAP7_75t_L g4609 ( 
.A(n_4514),
.B(n_4438),
.Y(n_4609)
);

INVx2_ASAP7_75t_L g4610 ( 
.A(n_4484),
.Y(n_4610)
);

INVx2_ASAP7_75t_L g4611 ( 
.A(n_4484),
.Y(n_4611)
);

NOR2xp67_ASAP7_75t_L g4612 ( 
.A(n_4468),
.B(n_4361),
.Y(n_4612)
);

OR2x2_ASAP7_75t_L g4613 ( 
.A(n_4575),
.B(n_4457),
.Y(n_4613)
);

HB1xp67_ASAP7_75t_L g4614 ( 
.A(n_4473),
.Y(n_4614)
);

NAND2xp5_ASAP7_75t_L g4615 ( 
.A(n_4580),
.B(n_4410),
.Y(n_4615)
);

AND2x2_ASAP7_75t_L g4616 ( 
.A(n_4514),
.B(n_4459),
.Y(n_4616)
);

OAI21xp5_ASAP7_75t_L g4617 ( 
.A1(n_4538),
.A2(n_4405),
.B(n_4395),
.Y(n_4617)
);

INVx2_ASAP7_75t_L g4618 ( 
.A(n_4540),
.Y(n_4618)
);

BUFx2_ASAP7_75t_L g4619 ( 
.A(n_4534),
.Y(n_4619)
);

AND2x2_ASAP7_75t_L g4620 ( 
.A(n_4514),
.B(n_4462),
.Y(n_4620)
);

INVx3_ASAP7_75t_L g4621 ( 
.A(n_4534),
.Y(n_4621)
);

INVxp67_ASAP7_75t_SL g4622 ( 
.A(n_4517),
.Y(n_4622)
);

INVxp67_ASAP7_75t_L g4623 ( 
.A(n_4585),
.Y(n_4623)
);

INVx1_ASAP7_75t_L g4624 ( 
.A(n_4507),
.Y(n_4624)
);

INVx2_ASAP7_75t_L g4625 ( 
.A(n_4535),
.Y(n_4625)
);

BUFx2_ASAP7_75t_L g4626 ( 
.A(n_4541),
.Y(n_4626)
);

INVx1_ASAP7_75t_L g4627 ( 
.A(n_4531),
.Y(n_4627)
);

INVxp67_ASAP7_75t_SL g4628 ( 
.A(n_4517),
.Y(n_4628)
);

INVx2_ASAP7_75t_L g4629 ( 
.A(n_4535),
.Y(n_4629)
);

INVx1_ASAP7_75t_L g4630 ( 
.A(n_4545),
.Y(n_4630)
);

AND2x2_ASAP7_75t_L g4631 ( 
.A(n_4517),
.B(n_4522),
.Y(n_4631)
);

BUFx3_ASAP7_75t_L g4632 ( 
.A(n_4482),
.Y(n_4632)
);

INVx1_ASAP7_75t_L g4633 ( 
.A(n_4545),
.Y(n_4633)
);

OR2x2_ASAP7_75t_L g4634 ( 
.A(n_4578),
.B(n_4368),
.Y(n_4634)
);

AND2x2_ASAP7_75t_L g4635 ( 
.A(n_4522),
.B(n_4356),
.Y(n_4635)
);

HB1xp67_ASAP7_75t_L g4636 ( 
.A(n_4476),
.Y(n_4636)
);

INVx2_ASAP7_75t_L g4637 ( 
.A(n_4535),
.Y(n_4637)
);

BUFx3_ASAP7_75t_L g4638 ( 
.A(n_4518),
.Y(n_4638)
);

AND2x2_ASAP7_75t_L g4639 ( 
.A(n_4522),
.B(n_4515),
.Y(n_4639)
);

AND2x2_ASAP7_75t_L g4640 ( 
.A(n_4515),
.B(n_4516),
.Y(n_4640)
);

INVx2_ASAP7_75t_L g4641 ( 
.A(n_4535),
.Y(n_4641)
);

OAI22xp5_ASAP7_75t_L g4642 ( 
.A1(n_4538),
.A2(n_4359),
.B1(n_4372),
.B2(n_4362),
.Y(n_4642)
);

AND2x2_ASAP7_75t_L g4643 ( 
.A(n_4516),
.B(n_4386),
.Y(n_4643)
);

AND2x2_ASAP7_75t_L g4644 ( 
.A(n_4519),
.B(n_4386),
.Y(n_4644)
);

INVx2_ASAP7_75t_L g4645 ( 
.A(n_4541),
.Y(n_4645)
);

NAND2xp5_ASAP7_75t_L g4646 ( 
.A(n_4580),
.B(n_4410),
.Y(n_4646)
);

AND2x2_ASAP7_75t_L g4647 ( 
.A(n_4519),
.B(n_4394),
.Y(n_4647)
);

AND2x2_ASAP7_75t_L g4648 ( 
.A(n_4528),
.B(n_4394),
.Y(n_4648)
);

OR2x2_ASAP7_75t_L g4649 ( 
.A(n_4578),
.B(n_4351),
.Y(n_4649)
);

AND2x2_ASAP7_75t_L g4650 ( 
.A(n_4528),
.B(n_4423),
.Y(n_4650)
);

INVx2_ASAP7_75t_L g4651 ( 
.A(n_4469),
.Y(n_4651)
);

BUFx2_ASAP7_75t_L g4652 ( 
.A(n_4494),
.Y(n_4652)
);

BUFx8_ASAP7_75t_L g4653 ( 
.A(n_4469),
.Y(n_4653)
);

AND2x2_ASAP7_75t_L g4654 ( 
.A(n_4510),
.B(n_4366),
.Y(n_4654)
);

AND2x4_ASAP7_75t_L g4655 ( 
.A(n_4468),
.B(n_4373),
.Y(n_4655)
);

AND2x2_ASAP7_75t_L g4656 ( 
.A(n_4510),
.B(n_4379),
.Y(n_4656)
);

INVx2_ASAP7_75t_L g4657 ( 
.A(n_4469),
.Y(n_4657)
);

HB1xp67_ASAP7_75t_L g4658 ( 
.A(n_4492),
.Y(n_4658)
);

BUFx3_ASAP7_75t_L g4659 ( 
.A(n_4518),
.Y(n_4659)
);

AND2x2_ASAP7_75t_L g4660 ( 
.A(n_4499),
.B(n_632),
.Y(n_4660)
);

INVx2_ASAP7_75t_L g4661 ( 
.A(n_4469),
.Y(n_4661)
);

INVx2_ASAP7_75t_L g4662 ( 
.A(n_4503),
.Y(n_4662)
);

AND2x2_ASAP7_75t_L g4663 ( 
.A(n_4499),
.B(n_633),
.Y(n_4663)
);

AND2x2_ASAP7_75t_L g4664 ( 
.A(n_4468),
.B(n_633),
.Y(n_4664)
);

INVxp67_ASAP7_75t_L g4665 ( 
.A(n_4529),
.Y(n_4665)
);

AND2x2_ASAP7_75t_L g4666 ( 
.A(n_4468),
.B(n_634),
.Y(n_4666)
);

INVxp67_ASAP7_75t_L g4667 ( 
.A(n_4529),
.Y(n_4667)
);

INVx2_ASAP7_75t_L g4668 ( 
.A(n_4503),
.Y(n_4668)
);

INVx1_ASAP7_75t_L g4669 ( 
.A(n_4549),
.Y(n_4669)
);

AOI21x1_ASAP7_75t_L g4670 ( 
.A1(n_4564),
.A2(n_635),
.B(n_636),
.Y(n_4670)
);

INVx1_ASAP7_75t_L g4671 ( 
.A(n_4549),
.Y(n_4671)
);

INVx2_ASAP7_75t_L g4672 ( 
.A(n_4496),
.Y(n_4672)
);

AND2x4_ASAP7_75t_L g4673 ( 
.A(n_4468),
.B(n_635),
.Y(n_4673)
);

AND2x2_ASAP7_75t_L g4674 ( 
.A(n_4477),
.B(n_636),
.Y(n_4674)
);

INVx2_ASAP7_75t_L g4675 ( 
.A(n_4558),
.Y(n_4675)
);

AND2x2_ASAP7_75t_L g4676 ( 
.A(n_4477),
.B(n_637),
.Y(n_4676)
);

INVx1_ASAP7_75t_L g4677 ( 
.A(n_4552),
.Y(n_4677)
);

NAND2xp5_ASAP7_75t_L g4678 ( 
.A(n_4520),
.B(n_637),
.Y(n_4678)
);

INVx1_ASAP7_75t_L g4679 ( 
.A(n_4552),
.Y(n_4679)
);

INVx2_ASAP7_75t_L g4680 ( 
.A(n_4488),
.Y(n_4680)
);

NAND2xp5_ASAP7_75t_L g4681 ( 
.A(n_4520),
.B(n_638),
.Y(n_4681)
);

AND2x2_ASAP7_75t_L g4682 ( 
.A(n_4563),
.B(n_638),
.Y(n_4682)
);

OR2x2_ASAP7_75t_L g4683 ( 
.A(n_4498),
.B(n_639),
.Y(n_4683)
);

INVx1_ASAP7_75t_L g4684 ( 
.A(n_4464),
.Y(n_4684)
);

INVx3_ASAP7_75t_L g4685 ( 
.A(n_4533),
.Y(n_4685)
);

INVx3_ASAP7_75t_L g4686 ( 
.A(n_4533),
.Y(n_4686)
);

INVx2_ASAP7_75t_L g4687 ( 
.A(n_4488),
.Y(n_4687)
);

INVx2_ASAP7_75t_L g4688 ( 
.A(n_4488),
.Y(n_4688)
);

NAND2x1_ASAP7_75t_L g4689 ( 
.A(n_4471),
.B(n_639),
.Y(n_4689)
);

AND2x2_ASAP7_75t_L g4690 ( 
.A(n_4512),
.B(n_4530),
.Y(n_4690)
);

INVxp67_ASAP7_75t_SL g4691 ( 
.A(n_4587),
.Y(n_4691)
);

AOI22xp33_ASAP7_75t_L g4692 ( 
.A1(n_4596),
.A2(n_673),
.B1(n_641),
.B2(n_643),
.Y(n_4692)
);

INVxp67_ASAP7_75t_SL g4693 ( 
.A(n_4508),
.Y(n_4693)
);

BUFx2_ASAP7_75t_L g4694 ( 
.A(n_4494),
.Y(n_4694)
);

INVx2_ASAP7_75t_SL g4695 ( 
.A(n_4508),
.Y(n_4695)
);

AO21x2_ASAP7_75t_L g4696 ( 
.A1(n_4466),
.A2(n_640),
.B(n_644),
.Y(n_4696)
);

AND2x2_ASAP7_75t_L g4697 ( 
.A(n_4512),
.B(n_4530),
.Y(n_4697)
);

OAI22xp5_ASAP7_75t_L g4698 ( 
.A1(n_4536),
.A2(n_4600),
.B1(n_4596),
.B2(n_4572),
.Y(n_4698)
);

AND2x4_ASAP7_75t_L g4699 ( 
.A(n_4467),
.B(n_640),
.Y(n_4699)
);

BUFx2_ASAP7_75t_SL g4700 ( 
.A(n_4489),
.Y(n_4700)
);

OR2x2_ASAP7_75t_L g4701 ( 
.A(n_4554),
.B(n_644),
.Y(n_4701)
);

INVx1_ASAP7_75t_L g4702 ( 
.A(n_4465),
.Y(n_4702)
);

AND2x4_ASAP7_75t_L g4703 ( 
.A(n_4467),
.B(n_645),
.Y(n_4703)
);

HB1xp67_ASAP7_75t_L g4704 ( 
.A(n_4560),
.Y(n_4704)
);

INVx2_ASAP7_75t_L g4705 ( 
.A(n_4479),
.Y(n_4705)
);

HB1xp67_ASAP7_75t_L g4706 ( 
.A(n_4560),
.Y(n_4706)
);

INVx1_ASAP7_75t_L g4707 ( 
.A(n_4474),
.Y(n_4707)
);

OR2x2_ASAP7_75t_L g4708 ( 
.A(n_4504),
.B(n_647),
.Y(n_4708)
);

NAND2xp5_ASAP7_75t_L g4709 ( 
.A(n_4581),
.B(n_4583),
.Y(n_4709)
);

OAI22xp5_ASAP7_75t_L g4710 ( 
.A1(n_4536),
.A2(n_647),
.B1(n_649),
.B2(n_650),
.Y(n_4710)
);

AND2x2_ASAP7_75t_L g4711 ( 
.A(n_4619),
.B(n_4621),
.Y(n_4711)
);

INVx1_ASAP7_75t_L g4712 ( 
.A(n_4626),
.Y(n_4712)
);

INVx1_ASAP7_75t_L g4713 ( 
.A(n_4626),
.Y(n_4713)
);

AND2x2_ASAP7_75t_L g4714 ( 
.A(n_4619),
.B(n_4631),
.Y(n_4714)
);

INVx2_ASAP7_75t_L g4715 ( 
.A(n_4645),
.Y(n_4715)
);

INVx2_ASAP7_75t_L g4716 ( 
.A(n_4645),
.Y(n_4716)
);

INVx1_ASAP7_75t_L g4717 ( 
.A(n_4614),
.Y(n_4717)
);

AND2x2_ASAP7_75t_L g4718 ( 
.A(n_4621),
.B(n_4529),
.Y(n_4718)
);

INVx2_ASAP7_75t_L g4719 ( 
.A(n_4689),
.Y(n_4719)
);

INVx1_ASAP7_75t_L g4720 ( 
.A(n_4704),
.Y(n_4720)
);

AND2x2_ASAP7_75t_L g4721 ( 
.A(n_4631),
.B(n_4621),
.Y(n_4721)
);

AND2x2_ASAP7_75t_L g4722 ( 
.A(n_4607),
.B(n_4479),
.Y(n_4722)
);

INVx3_ASAP7_75t_L g4723 ( 
.A(n_4689),
.Y(n_4723)
);

OR2x2_ASAP7_75t_L g4724 ( 
.A(n_4605),
.B(n_4497),
.Y(n_4724)
);

AND2x4_ASAP7_75t_SL g4725 ( 
.A(n_4618),
.B(n_4529),
.Y(n_4725)
);

OR2x2_ASAP7_75t_L g4726 ( 
.A(n_4605),
.B(n_4504),
.Y(n_4726)
);

INVx1_ASAP7_75t_L g4727 ( 
.A(n_4706),
.Y(n_4727)
);

HB1xp67_ASAP7_75t_L g4728 ( 
.A(n_4603),
.Y(n_4728)
);

AND2x2_ASAP7_75t_L g4729 ( 
.A(n_4607),
.B(n_4481),
.Y(n_4729)
);

INVx2_ASAP7_75t_L g4730 ( 
.A(n_4680),
.Y(n_4730)
);

INVx2_ASAP7_75t_L g4731 ( 
.A(n_4680),
.Y(n_4731)
);

INVx2_ASAP7_75t_SL g4732 ( 
.A(n_4652),
.Y(n_4732)
);

BUFx3_ASAP7_75t_L g4733 ( 
.A(n_4653),
.Y(n_4733)
);

BUFx3_ASAP7_75t_L g4734 ( 
.A(n_4653),
.Y(n_4734)
);

INVx2_ASAP7_75t_L g4735 ( 
.A(n_4687),
.Y(n_4735)
);

INVx1_ASAP7_75t_SL g4736 ( 
.A(n_4652),
.Y(n_4736)
);

OR2x2_ASAP7_75t_L g4737 ( 
.A(n_4613),
.B(n_4509),
.Y(n_4737)
);

HB1xp67_ASAP7_75t_L g4738 ( 
.A(n_4603),
.Y(n_4738)
);

OR2x2_ASAP7_75t_L g4739 ( 
.A(n_4613),
.B(n_4509),
.Y(n_4739)
);

INVx1_ASAP7_75t_L g4740 ( 
.A(n_4636),
.Y(n_4740)
);

BUFx3_ASAP7_75t_L g4741 ( 
.A(n_4653),
.Y(n_4741)
);

INVx2_ASAP7_75t_SL g4742 ( 
.A(n_4694),
.Y(n_4742)
);

AND2x2_ASAP7_75t_L g4743 ( 
.A(n_4632),
.B(n_4490),
.Y(n_4743)
);

INVx2_ASAP7_75t_L g4744 ( 
.A(n_4687),
.Y(n_4744)
);

INVx3_ASAP7_75t_L g4745 ( 
.A(n_4638),
.Y(n_4745)
);

INVx1_ASAP7_75t_L g4746 ( 
.A(n_4658),
.Y(n_4746)
);

INVx2_ASAP7_75t_L g4747 ( 
.A(n_4688),
.Y(n_4747)
);

INVx4_ASAP7_75t_L g4748 ( 
.A(n_4673),
.Y(n_4748)
);

INVx2_ASAP7_75t_L g4749 ( 
.A(n_4688),
.Y(n_4749)
);

AND2x2_ASAP7_75t_L g4750 ( 
.A(n_4632),
.B(n_4490),
.Y(n_4750)
);

INVx1_ASAP7_75t_L g4751 ( 
.A(n_4708),
.Y(n_4751)
);

INVx2_ASAP7_75t_SL g4752 ( 
.A(n_4694),
.Y(n_4752)
);

INVx2_ASAP7_75t_L g4753 ( 
.A(n_4670),
.Y(n_4753)
);

INVx1_ASAP7_75t_L g4754 ( 
.A(n_4708),
.Y(n_4754)
);

AND2x2_ASAP7_75t_L g4755 ( 
.A(n_4622),
.B(n_4481),
.Y(n_4755)
);

OR2x2_ASAP7_75t_L g4756 ( 
.A(n_4709),
.B(n_4604),
.Y(n_4756)
);

HB1xp67_ASAP7_75t_L g4757 ( 
.A(n_4606),
.Y(n_4757)
);

INVx1_ASAP7_75t_L g4758 ( 
.A(n_4606),
.Y(n_4758)
);

NAND2x1_ASAP7_75t_L g4759 ( 
.A(n_4690),
.B(n_4513),
.Y(n_4759)
);

INVx1_ASAP7_75t_L g4760 ( 
.A(n_4624),
.Y(n_4760)
);

INVxp67_ASAP7_75t_SL g4761 ( 
.A(n_4624),
.Y(n_4761)
);

INVx3_ASAP7_75t_L g4762 ( 
.A(n_4638),
.Y(n_4762)
);

INVx1_ASAP7_75t_L g4763 ( 
.A(n_4627),
.Y(n_4763)
);

AND2x2_ASAP7_75t_L g4764 ( 
.A(n_4693),
.B(n_4471),
.Y(n_4764)
);

INVx3_ASAP7_75t_L g4765 ( 
.A(n_4659),
.Y(n_4765)
);

INVx1_ASAP7_75t_L g4766 ( 
.A(n_4627),
.Y(n_4766)
);

INVx1_ASAP7_75t_L g4767 ( 
.A(n_4630),
.Y(n_4767)
);

INVx2_ASAP7_75t_L g4768 ( 
.A(n_4670),
.Y(n_4768)
);

INVx1_ASAP7_75t_L g4769 ( 
.A(n_4630),
.Y(n_4769)
);

AOI22xp33_ASAP7_75t_L g4770 ( 
.A1(n_4615),
.A2(n_4600),
.B1(n_4598),
.B2(n_4594),
.Y(n_4770)
);

HB1xp67_ASAP7_75t_L g4771 ( 
.A(n_4696),
.Y(n_4771)
);

NOR2x1_ASAP7_75t_SL g4772 ( 
.A(n_4696),
.B(n_4471),
.Y(n_4772)
);

INVx1_ASAP7_75t_L g4773 ( 
.A(n_4633),
.Y(n_4773)
);

AOI22xp33_ASAP7_75t_L g4774 ( 
.A1(n_4646),
.A2(n_4582),
.B1(n_4568),
.B2(n_4570),
.Y(n_4774)
);

INVx2_ASAP7_75t_L g4775 ( 
.A(n_4696),
.Y(n_4775)
);

INVx2_ASAP7_75t_L g4776 ( 
.A(n_4690),
.Y(n_4776)
);

INVx2_ASAP7_75t_L g4777 ( 
.A(n_4697),
.Y(n_4777)
);

OR2x2_ASAP7_75t_L g4778 ( 
.A(n_4736),
.B(n_4604),
.Y(n_4778)
);

OAI22xp5_ASAP7_75t_L g4779 ( 
.A1(n_4774),
.A2(n_4617),
.B1(n_4612),
.B2(n_4691),
.Y(n_4779)
);

INVx1_ASAP7_75t_L g4780 ( 
.A(n_4714),
.Y(n_4780)
);

NAND2xp5_ASAP7_75t_L g4781 ( 
.A(n_4714),
.B(n_4623),
.Y(n_4781)
);

AND2x2_ASAP7_75t_L g4782 ( 
.A(n_4714),
.B(n_4700),
.Y(n_4782)
);

OR2x2_ASAP7_75t_L g4783 ( 
.A(n_4736),
.B(n_4602),
.Y(n_4783)
);

AND2x2_ASAP7_75t_L g4784 ( 
.A(n_4718),
.B(n_4700),
.Y(n_4784)
);

AND2x4_ASAP7_75t_SL g4785 ( 
.A(n_4745),
.B(n_4675),
.Y(n_4785)
);

NAND2xp5_ASAP7_75t_L g4786 ( 
.A(n_4732),
.B(n_4665),
.Y(n_4786)
);

NAND3xp33_ASAP7_75t_L g4787 ( 
.A(n_4770),
.B(n_4698),
.C(n_4617),
.Y(n_4787)
);

AND2x2_ASAP7_75t_L g4788 ( 
.A(n_4718),
.B(n_4685),
.Y(n_4788)
);

INVx1_ASAP7_75t_L g4789 ( 
.A(n_4711),
.Y(n_4789)
);

NAND2xp5_ASAP7_75t_L g4790 ( 
.A(n_4732),
.B(n_4667),
.Y(n_4790)
);

AND2x2_ASAP7_75t_L g4791 ( 
.A(n_4732),
.B(n_4685),
.Y(n_4791)
);

INVx1_ASAP7_75t_L g4792 ( 
.A(n_4711),
.Y(n_4792)
);

NAND2xp5_ASAP7_75t_L g4793 ( 
.A(n_4742),
.B(n_4602),
.Y(n_4793)
);

NOR2x1_ASAP7_75t_L g4794 ( 
.A(n_4723),
.B(n_4659),
.Y(n_4794)
);

AND2x2_ASAP7_75t_L g4795 ( 
.A(n_4742),
.B(n_4685),
.Y(n_4795)
);

AND2x2_ASAP7_75t_L g4796 ( 
.A(n_4742),
.B(n_4686),
.Y(n_4796)
);

AND2x2_ASAP7_75t_L g4797 ( 
.A(n_4752),
.B(n_4686),
.Y(n_4797)
);

INVx1_ASAP7_75t_L g4798 ( 
.A(n_4728),
.Y(n_4798)
);

INVx2_ASAP7_75t_L g4799 ( 
.A(n_4723),
.Y(n_4799)
);

NAND2xp5_ASAP7_75t_SL g4800 ( 
.A(n_4753),
.B(n_4612),
.Y(n_4800)
);

INVx1_ASAP7_75t_L g4801 ( 
.A(n_4728),
.Y(n_4801)
);

NOR2xp33_ASAP7_75t_L g4802 ( 
.A(n_4752),
.B(n_4675),
.Y(n_4802)
);

NAND2xp5_ASAP7_75t_L g4803 ( 
.A(n_4752),
.B(n_4628),
.Y(n_4803)
);

NAND2xp5_ASAP7_75t_L g4804 ( 
.A(n_4745),
.B(n_4618),
.Y(n_4804)
);

NAND2xp5_ASAP7_75t_L g4805 ( 
.A(n_4745),
.B(n_4695),
.Y(n_4805)
);

INVx1_ASAP7_75t_SL g4806 ( 
.A(n_4725),
.Y(n_4806)
);

INVx1_ASAP7_75t_L g4807 ( 
.A(n_4738),
.Y(n_4807)
);

INVx2_ASAP7_75t_L g4808 ( 
.A(n_4723),
.Y(n_4808)
);

HB1xp67_ASAP7_75t_L g4809 ( 
.A(n_4723),
.Y(n_4809)
);

NAND2xp5_ASAP7_75t_L g4810 ( 
.A(n_4745),
.B(n_4695),
.Y(n_4810)
);

INVx1_ASAP7_75t_L g4811 ( 
.A(n_4738),
.Y(n_4811)
);

INVx2_ASAP7_75t_L g4812 ( 
.A(n_4721),
.Y(n_4812)
);

AND2x2_ASAP7_75t_L g4813 ( 
.A(n_4725),
.B(n_4686),
.Y(n_4813)
);

AND2x2_ASAP7_75t_L g4814 ( 
.A(n_4725),
.B(n_4651),
.Y(n_4814)
);

AND2x2_ASAP7_75t_L g4815 ( 
.A(n_4721),
.B(n_4651),
.Y(n_4815)
);

HB1xp67_ASAP7_75t_L g4816 ( 
.A(n_4762),
.Y(n_4816)
);

INVx1_ASAP7_75t_L g4817 ( 
.A(n_4757),
.Y(n_4817)
);

AND2x2_ASAP7_75t_L g4818 ( 
.A(n_4721),
.B(n_4657),
.Y(n_4818)
);

INVx1_ASAP7_75t_L g4819 ( 
.A(n_4757),
.Y(n_4819)
);

INVx1_ASAP7_75t_L g4820 ( 
.A(n_4720),
.Y(n_4820)
);

INVxp67_ASAP7_75t_SL g4821 ( 
.A(n_4762),
.Y(n_4821)
);

INVx1_ASAP7_75t_L g4822 ( 
.A(n_4720),
.Y(n_4822)
);

NAND2xp5_ASAP7_75t_L g4823 ( 
.A(n_4762),
.B(n_4765),
.Y(n_4823)
);

INVx1_ASAP7_75t_L g4824 ( 
.A(n_4727),
.Y(n_4824)
);

NAND2xp5_ASAP7_75t_L g4825 ( 
.A(n_4762),
.B(n_4635),
.Y(n_4825)
);

BUFx3_ASAP7_75t_L g4826 ( 
.A(n_4765),
.Y(n_4826)
);

AOI221xp5_ASAP7_75t_L g4827 ( 
.A1(n_4759),
.A2(n_4642),
.B1(n_4710),
.B2(n_4643),
.C(n_4647),
.Y(n_4827)
);

AND2x2_ASAP7_75t_L g4828 ( 
.A(n_4765),
.B(n_4657),
.Y(n_4828)
);

INVx1_ASAP7_75t_L g4829 ( 
.A(n_4727),
.Y(n_4829)
);

INVx2_ASAP7_75t_L g4830 ( 
.A(n_4765),
.Y(n_4830)
);

INVx2_ASAP7_75t_L g4831 ( 
.A(n_4719),
.Y(n_4831)
);

INVx1_ASAP7_75t_L g4832 ( 
.A(n_4761),
.Y(n_4832)
);

OR2x2_ASAP7_75t_L g4833 ( 
.A(n_4740),
.B(n_4746),
.Y(n_4833)
);

INVx1_ASAP7_75t_L g4834 ( 
.A(n_4761),
.Y(n_4834)
);

AND2x2_ASAP7_75t_L g4835 ( 
.A(n_4782),
.B(n_4661),
.Y(n_4835)
);

NAND2xp5_ASAP7_75t_SL g4836 ( 
.A(n_4782),
.B(n_4697),
.Y(n_4836)
);

NAND2xp5_ASAP7_75t_L g4837 ( 
.A(n_4784),
.B(n_4743),
.Y(n_4837)
);

AND2x2_ASAP7_75t_SL g4838 ( 
.A(n_4784),
.B(n_4655),
.Y(n_4838)
);

BUFx2_ASAP7_75t_L g4839 ( 
.A(n_4809),
.Y(n_4839)
);

INVx1_ASAP7_75t_L g4840 ( 
.A(n_4816),
.Y(n_4840)
);

AND2x2_ASAP7_75t_L g4841 ( 
.A(n_4785),
.B(n_4661),
.Y(n_4841)
);

INVx1_ASAP7_75t_L g4842 ( 
.A(n_4778),
.Y(n_4842)
);

INVx1_ASAP7_75t_L g4843 ( 
.A(n_4812),
.Y(n_4843)
);

AND2x2_ASAP7_75t_L g4844 ( 
.A(n_4785),
.B(n_4764),
.Y(n_4844)
);

AND2x2_ASAP7_75t_L g4845 ( 
.A(n_4815),
.B(n_4818),
.Y(n_4845)
);

INVx2_ASAP7_75t_L g4846 ( 
.A(n_4826),
.Y(n_4846)
);

AND2x2_ASAP7_75t_L g4847 ( 
.A(n_4815),
.B(n_4764),
.Y(n_4847)
);

NAND2x1_ASAP7_75t_L g4848 ( 
.A(n_4794),
.B(n_4719),
.Y(n_4848)
);

AND2x2_ASAP7_75t_L g4849 ( 
.A(n_4818),
.B(n_4743),
.Y(n_4849)
);

NAND2xp5_ASAP7_75t_L g4850 ( 
.A(n_4802),
.B(n_4750),
.Y(n_4850)
);

AND2x4_ASAP7_75t_L g4851 ( 
.A(n_4826),
.B(n_4719),
.Y(n_4851)
);

INVx3_ASAP7_75t_L g4852 ( 
.A(n_4799),
.Y(n_4852)
);

NAND2xp5_ASAP7_75t_L g4853 ( 
.A(n_4802),
.B(n_4750),
.Y(n_4853)
);

NAND2xp5_ASAP7_75t_L g4854 ( 
.A(n_4788),
.B(n_4635),
.Y(n_4854)
);

BUFx2_ASAP7_75t_SL g4855 ( 
.A(n_4830),
.Y(n_4855)
);

INVx1_ASAP7_75t_L g4856 ( 
.A(n_4778),
.Y(n_4856)
);

INVx2_ASAP7_75t_L g4857 ( 
.A(n_4791),
.Y(n_4857)
);

AND2x4_ASAP7_75t_L g4858 ( 
.A(n_4791),
.B(n_4733),
.Y(n_4858)
);

AND2x2_ASAP7_75t_L g4859 ( 
.A(n_4788),
.B(n_4733),
.Y(n_4859)
);

NAND2xp5_ASAP7_75t_L g4860 ( 
.A(n_4795),
.B(n_4796),
.Y(n_4860)
);

NAND2xp5_ASAP7_75t_L g4861 ( 
.A(n_4795),
.B(n_4682),
.Y(n_4861)
);

HB1xp67_ASAP7_75t_L g4862 ( 
.A(n_4796),
.Y(n_4862)
);

AND2x2_ASAP7_75t_L g4863 ( 
.A(n_4813),
.B(n_4733),
.Y(n_4863)
);

INVx2_ASAP7_75t_L g4864 ( 
.A(n_4797),
.Y(n_4864)
);

NAND2xp5_ASAP7_75t_L g4865 ( 
.A(n_4797),
.B(n_4682),
.Y(n_4865)
);

OR2x2_ASAP7_75t_L g4866 ( 
.A(n_4783),
.B(n_4753),
.Y(n_4866)
);

AOI22xp33_ASAP7_75t_L g4867 ( 
.A1(n_4787),
.A2(n_4643),
.B1(n_4647),
.B2(n_4644),
.Y(n_4867)
);

INVx2_ASAP7_75t_L g4868 ( 
.A(n_4799),
.Y(n_4868)
);

AND2x2_ASAP7_75t_L g4869 ( 
.A(n_4813),
.B(n_4814),
.Y(n_4869)
);

AND2x2_ASAP7_75t_L g4870 ( 
.A(n_4814),
.B(n_4734),
.Y(n_4870)
);

AOI22xp33_ASAP7_75t_SL g4871 ( 
.A1(n_4779),
.A2(n_4772),
.B1(n_4648),
.B2(n_4644),
.Y(n_4871)
);

BUFx6f_ASAP7_75t_L g4872 ( 
.A(n_4832),
.Y(n_4872)
);

OR2x2_ASAP7_75t_L g4873 ( 
.A(n_4783),
.B(n_4753),
.Y(n_4873)
);

INVx2_ASAP7_75t_L g4874 ( 
.A(n_4808),
.Y(n_4874)
);

INVx1_ASAP7_75t_L g4875 ( 
.A(n_4812),
.Y(n_4875)
);

INVx1_ASAP7_75t_L g4876 ( 
.A(n_4821),
.Y(n_4876)
);

AND2x2_ASAP7_75t_L g4877 ( 
.A(n_4806),
.B(n_4734),
.Y(n_4877)
);

NOR2xp67_ASAP7_75t_L g4878 ( 
.A(n_4803),
.B(n_4748),
.Y(n_4878)
);

AND2x2_ASAP7_75t_L g4879 ( 
.A(n_4780),
.B(n_4734),
.Y(n_4879)
);

INVx1_ASAP7_75t_L g4880 ( 
.A(n_4834),
.Y(n_4880)
);

AND2x4_ASAP7_75t_L g4881 ( 
.A(n_4808),
.B(n_4741),
.Y(n_4881)
);

AND2x2_ASAP7_75t_L g4882 ( 
.A(n_4828),
.B(n_4741),
.Y(n_4882)
);

INVx2_ASAP7_75t_L g4883 ( 
.A(n_4830),
.Y(n_4883)
);

NAND2xp5_ASAP7_75t_SL g4884 ( 
.A(n_4827),
.B(n_4655),
.Y(n_4884)
);

INVx1_ASAP7_75t_L g4885 ( 
.A(n_4831),
.Y(n_4885)
);

INVx1_ASAP7_75t_L g4886 ( 
.A(n_4831),
.Y(n_4886)
);

AND2x2_ASAP7_75t_L g4887 ( 
.A(n_4869),
.B(n_4741),
.Y(n_4887)
);

OR2x2_ASAP7_75t_L g4888 ( 
.A(n_4854),
.B(n_4781),
.Y(n_4888)
);

INVx1_ASAP7_75t_L g4889 ( 
.A(n_4839),
.Y(n_4889)
);

AND2x4_ASAP7_75t_L g4890 ( 
.A(n_4851),
.B(n_4828),
.Y(n_4890)
);

BUFx3_ASAP7_75t_L g4891 ( 
.A(n_4844),
.Y(n_4891)
);

INVx1_ASAP7_75t_L g4892 ( 
.A(n_4839),
.Y(n_4892)
);

HB1xp67_ASAP7_75t_L g4893 ( 
.A(n_4862),
.Y(n_4893)
);

INVx1_ASAP7_75t_L g4894 ( 
.A(n_4855),
.Y(n_4894)
);

NOR2xp67_ASAP7_75t_L g4895 ( 
.A(n_4842),
.B(n_4748),
.Y(n_4895)
);

HB1xp67_ASAP7_75t_L g4896 ( 
.A(n_4851),
.Y(n_4896)
);

AND2x2_ASAP7_75t_L g4897 ( 
.A(n_4845),
.B(n_4835),
.Y(n_4897)
);

NAND2xp5_ASAP7_75t_L g4898 ( 
.A(n_4838),
.B(n_4789),
.Y(n_4898)
);

AND2x2_ASAP7_75t_L g4899 ( 
.A(n_4845),
.B(n_4792),
.Y(n_4899)
);

AND2x4_ASAP7_75t_L g4900 ( 
.A(n_4851),
.B(n_4748),
.Y(n_4900)
);

AND2x2_ASAP7_75t_L g4901 ( 
.A(n_4835),
.B(n_4639),
.Y(n_4901)
);

AND2x2_ASAP7_75t_L g4902 ( 
.A(n_4869),
.B(n_4639),
.Y(n_4902)
);

AND2x2_ASAP7_75t_L g4903 ( 
.A(n_4859),
.B(n_4601),
.Y(n_4903)
);

INVx2_ASAP7_75t_SL g4904 ( 
.A(n_4848),
.Y(n_4904)
);

INVx1_ASAP7_75t_L g4905 ( 
.A(n_4855),
.Y(n_4905)
);

INVx2_ASAP7_75t_SL g4906 ( 
.A(n_4848),
.Y(n_4906)
);

NAND2xp5_ASAP7_75t_L g4907 ( 
.A(n_4838),
.B(n_4748),
.Y(n_4907)
);

AND2x2_ASAP7_75t_L g4908 ( 
.A(n_4859),
.B(n_4601),
.Y(n_4908)
);

NAND2x1_ASAP7_75t_SL g4909 ( 
.A(n_4844),
.B(n_4771),
.Y(n_4909)
);

INVx2_ASAP7_75t_L g4910 ( 
.A(n_4852),
.Y(n_4910)
);

OR2x2_ASAP7_75t_L g4911 ( 
.A(n_4861),
.B(n_4825),
.Y(n_4911)
);

NAND2xp5_ASAP7_75t_L g4912 ( 
.A(n_4847),
.B(n_4740),
.Y(n_4912)
);

AND2x2_ASAP7_75t_L g4913 ( 
.A(n_4877),
.B(n_4870),
.Y(n_4913)
);

INVx1_ASAP7_75t_L g4914 ( 
.A(n_4852),
.Y(n_4914)
);

AND2x2_ASAP7_75t_L g4915 ( 
.A(n_4847),
.B(n_4625),
.Y(n_4915)
);

INVx1_ASAP7_75t_L g4916 ( 
.A(n_4852),
.Y(n_4916)
);

AND2x4_ASAP7_75t_L g4917 ( 
.A(n_4841),
.B(n_4712),
.Y(n_4917)
);

OR2x2_ASAP7_75t_L g4918 ( 
.A(n_4865),
.B(n_4786),
.Y(n_4918)
);

OR2x2_ASAP7_75t_L g4919 ( 
.A(n_4860),
.B(n_4790),
.Y(n_4919)
);

NAND2x1p5_ASAP7_75t_L g4920 ( 
.A(n_4858),
.B(n_4673),
.Y(n_4920)
);

AND2x4_ASAP7_75t_L g4921 ( 
.A(n_4841),
.B(n_4857),
.Y(n_4921)
);

OR2x2_ASAP7_75t_L g4922 ( 
.A(n_4850),
.B(n_4793),
.Y(n_4922)
);

AND2x2_ASAP7_75t_L g4923 ( 
.A(n_4870),
.B(n_4625),
.Y(n_4923)
);

OR2x2_ASAP7_75t_L g4924 ( 
.A(n_4853),
.B(n_4756),
.Y(n_4924)
);

AND2x2_ASAP7_75t_L g4925 ( 
.A(n_4913),
.B(n_4882),
.Y(n_4925)
);

INVx2_ASAP7_75t_L g4926 ( 
.A(n_4909),
.Y(n_4926)
);

OR2x2_ASAP7_75t_L g4927 ( 
.A(n_4896),
.B(n_4866),
.Y(n_4927)
);

INVx2_ASAP7_75t_L g4928 ( 
.A(n_4896),
.Y(n_4928)
);

NAND2xp5_ASAP7_75t_L g4929 ( 
.A(n_4901),
.B(n_4882),
.Y(n_4929)
);

NAND2xp5_ASAP7_75t_L g4930 ( 
.A(n_4901),
.B(n_4849),
.Y(n_4930)
);

OR2x2_ASAP7_75t_L g4931 ( 
.A(n_4893),
.B(n_4866),
.Y(n_4931)
);

NAND2x1_ASAP7_75t_SL g4932 ( 
.A(n_4890),
.B(n_4771),
.Y(n_4932)
);

INVx1_ASAP7_75t_L g4933 ( 
.A(n_4893),
.Y(n_4933)
);

HB1xp67_ASAP7_75t_L g4934 ( 
.A(n_4890),
.Y(n_4934)
);

AND2x2_ASAP7_75t_L g4935 ( 
.A(n_4902),
.B(n_4849),
.Y(n_4935)
);

AND2x2_ASAP7_75t_L g4936 ( 
.A(n_4902),
.B(n_4897),
.Y(n_4936)
);

INVx2_ASAP7_75t_L g4937 ( 
.A(n_4890),
.Y(n_4937)
);

NAND2xp5_ASAP7_75t_L g4938 ( 
.A(n_4897),
.B(n_4858),
.Y(n_4938)
);

HB1xp67_ASAP7_75t_L g4939 ( 
.A(n_4900),
.Y(n_4939)
);

AND2x2_ASAP7_75t_L g4940 ( 
.A(n_4903),
.B(n_4863),
.Y(n_4940)
);

INVx1_ASAP7_75t_L g4941 ( 
.A(n_4910),
.Y(n_4941)
);

INVx1_ASAP7_75t_L g4942 ( 
.A(n_4910),
.Y(n_4942)
);

OR2x2_ASAP7_75t_L g4943 ( 
.A(n_4889),
.B(n_4873),
.Y(n_4943)
);

AND2x2_ASAP7_75t_L g4944 ( 
.A(n_4908),
.B(n_4863),
.Y(n_4944)
);

INVx1_ASAP7_75t_L g4945 ( 
.A(n_4921),
.Y(n_4945)
);

INVx1_ASAP7_75t_L g4946 ( 
.A(n_4921),
.Y(n_4946)
);

NOR2xp67_ASAP7_75t_L g4947 ( 
.A(n_4904),
.B(n_4842),
.Y(n_4947)
);

INVx2_ASAP7_75t_L g4948 ( 
.A(n_4900),
.Y(n_4948)
);

INVx2_ASAP7_75t_SL g4949 ( 
.A(n_4900),
.Y(n_4949)
);

INVx2_ASAP7_75t_L g4950 ( 
.A(n_4904),
.Y(n_4950)
);

NOR2x1_ASAP7_75t_L g4951 ( 
.A(n_4891),
.B(n_4873),
.Y(n_4951)
);

AND2x2_ASAP7_75t_L g4952 ( 
.A(n_4923),
.B(n_4877),
.Y(n_4952)
);

NOR2xp33_ASAP7_75t_SL g4953 ( 
.A(n_4887),
.B(n_4653),
.Y(n_4953)
);

INVx1_ASAP7_75t_L g4954 ( 
.A(n_4921),
.Y(n_4954)
);

AND2x2_ASAP7_75t_L g4955 ( 
.A(n_4923),
.B(n_4858),
.Y(n_4955)
);

INVx2_ASAP7_75t_L g4956 ( 
.A(n_4906),
.Y(n_4956)
);

INVx1_ASAP7_75t_L g4957 ( 
.A(n_4927),
.Y(n_4957)
);

A2O1A1Ixp33_ASAP7_75t_L g4958 ( 
.A1(n_4932),
.A2(n_4759),
.B(n_4768),
.C(n_4871),
.Y(n_4958)
);

AND2x4_ASAP7_75t_L g4959 ( 
.A(n_4955),
.B(n_4891),
.Y(n_4959)
);

OR2x2_ASAP7_75t_L g4960 ( 
.A(n_4929),
.B(n_4912),
.Y(n_4960)
);

AND2x2_ASAP7_75t_L g4961 ( 
.A(n_4925),
.B(n_4899),
.Y(n_4961)
);

NAND2xp5_ASAP7_75t_L g4962 ( 
.A(n_4952),
.B(n_4915),
.Y(n_4962)
);

NAND2xp5_ASAP7_75t_L g4963 ( 
.A(n_4952),
.B(n_4915),
.Y(n_4963)
);

AND2x2_ASAP7_75t_L g4964 ( 
.A(n_4925),
.B(n_4899),
.Y(n_4964)
);

INVx1_ASAP7_75t_L g4965 ( 
.A(n_4927),
.Y(n_4965)
);

NAND2xp5_ASAP7_75t_L g4966 ( 
.A(n_4955),
.B(n_4857),
.Y(n_4966)
);

AND2x2_ASAP7_75t_L g4967 ( 
.A(n_4940),
.B(n_4879),
.Y(n_4967)
);

AND2x2_ASAP7_75t_L g4968 ( 
.A(n_4940),
.B(n_4879),
.Y(n_4968)
);

NAND2xp5_ASAP7_75t_L g4969 ( 
.A(n_4947),
.B(n_4856),
.Y(n_4969)
);

AND2x2_ASAP7_75t_L g4970 ( 
.A(n_4944),
.B(n_4864),
.Y(n_4970)
);

INVx1_ASAP7_75t_L g4971 ( 
.A(n_4932),
.Y(n_4971)
);

AND2x2_ASAP7_75t_L g4972 ( 
.A(n_4944),
.B(n_4864),
.Y(n_4972)
);

NAND2xp5_ASAP7_75t_L g4973 ( 
.A(n_4951),
.B(n_4856),
.Y(n_4973)
);

INVx1_ASAP7_75t_L g4974 ( 
.A(n_4934),
.Y(n_4974)
);

INVx1_ASAP7_75t_L g4975 ( 
.A(n_4931),
.Y(n_4975)
);

INVx1_ASAP7_75t_L g4976 ( 
.A(n_4931),
.Y(n_4976)
);

OR2x2_ASAP7_75t_L g4977 ( 
.A(n_4938),
.B(n_4804),
.Y(n_4977)
);

INVx1_ASAP7_75t_L g4978 ( 
.A(n_4939),
.Y(n_4978)
);

OR2x2_ASAP7_75t_L g4979 ( 
.A(n_4930),
.B(n_4756),
.Y(n_4979)
);

NAND2xp5_ASAP7_75t_L g4980 ( 
.A(n_4928),
.B(n_4872),
.Y(n_4980)
);

BUFx2_ASAP7_75t_L g4981 ( 
.A(n_4959),
.Y(n_4981)
);

INVx1_ASAP7_75t_L g4982 ( 
.A(n_4961),
.Y(n_4982)
);

OR2x2_ASAP7_75t_L g4983 ( 
.A(n_4962),
.B(n_4837),
.Y(n_4983)
);

INVx2_ASAP7_75t_SL g4984 ( 
.A(n_4959),
.Y(n_4984)
);

NAND2xp5_ASAP7_75t_L g4985 ( 
.A(n_4964),
.B(n_4936),
.Y(n_4985)
);

AND2x2_ASAP7_75t_L g4986 ( 
.A(n_4967),
.B(n_4935),
.Y(n_4986)
);

AOI22xp5_ASAP7_75t_L g4987 ( 
.A1(n_4968),
.A2(n_4884),
.B1(n_4867),
.B2(n_4768),
.Y(n_4987)
);

OR2x2_ASAP7_75t_L g4988 ( 
.A(n_4963),
.B(n_4898),
.Y(n_4988)
);

INVx1_ASAP7_75t_L g4989 ( 
.A(n_4973),
.Y(n_4989)
);

AND2x2_ASAP7_75t_L g4990 ( 
.A(n_4970),
.B(n_4935),
.Y(n_4990)
);

OAI31xp33_ASAP7_75t_L g4991 ( 
.A1(n_4958),
.A2(n_4768),
.A3(n_4712),
.B(n_4713),
.Y(n_4991)
);

INVx2_ASAP7_75t_SL g4992 ( 
.A(n_4972),
.Y(n_4992)
);

AOI22xp5_ASAP7_75t_L g4993 ( 
.A1(n_4973),
.A2(n_4713),
.B1(n_4953),
.B2(n_4906),
.Y(n_4993)
);

INVx1_ASAP7_75t_L g4994 ( 
.A(n_4969),
.Y(n_4994)
);

INVx2_ASAP7_75t_L g4995 ( 
.A(n_4957),
.Y(n_4995)
);

OAI21xp5_ASAP7_75t_L g4996 ( 
.A1(n_4966),
.A2(n_4895),
.B(n_4936),
.Y(n_4996)
);

NAND2xp5_ASAP7_75t_L g4997 ( 
.A(n_4974),
.B(n_4881),
.Y(n_4997)
);

INVx1_ASAP7_75t_L g4998 ( 
.A(n_4969),
.Y(n_4998)
);

HB1xp67_ASAP7_75t_L g4999 ( 
.A(n_4965),
.Y(n_4999)
);

NAND2xp5_ASAP7_75t_L g5000 ( 
.A(n_4978),
.B(n_4881),
.Y(n_5000)
);

OAI31xp33_ASAP7_75t_L g5001 ( 
.A1(n_4981),
.A2(n_4800),
.A3(n_4920),
.B(n_4892),
.Y(n_5001)
);

NAND2x1p5_ASAP7_75t_L g5002 ( 
.A(n_4984),
.B(n_4949),
.Y(n_5002)
);

AOI322xp5_ASAP7_75t_L g5003 ( 
.A1(n_4987),
.A2(n_4836),
.A3(n_4800),
.B1(n_4926),
.B2(n_4717),
.C1(n_4905),
.C2(n_4894),
.Y(n_5003)
);

INVx1_ASAP7_75t_L g5004 ( 
.A(n_4990),
.Y(n_5004)
);

OAI21xp33_ASAP7_75t_SL g5005 ( 
.A1(n_4991),
.A2(n_4716),
.B(n_4715),
.Y(n_5005)
);

INVxp67_ASAP7_75t_SL g5006 ( 
.A(n_4985),
.Y(n_5006)
);

NAND2xp5_ASAP7_75t_L g5007 ( 
.A(n_4986),
.B(n_4881),
.Y(n_5007)
);

INVx2_ASAP7_75t_L g5008 ( 
.A(n_4992),
.Y(n_5008)
);

OAI21xp33_ASAP7_75t_L g5009 ( 
.A1(n_4987),
.A2(n_4888),
.B(n_4810),
.Y(n_5009)
);

AOI22xp5_ASAP7_75t_L g5010 ( 
.A1(n_4982),
.A2(n_4629),
.B1(n_4641),
.B2(n_4637),
.Y(n_5010)
);

NAND2xp5_ASAP7_75t_L g5011 ( 
.A(n_4993),
.B(n_4945),
.Y(n_5011)
);

INVx1_ASAP7_75t_L g5012 ( 
.A(n_4997),
.Y(n_5012)
);

INVx2_ASAP7_75t_L g5013 ( 
.A(n_4995),
.Y(n_5013)
);

OR2x2_ASAP7_75t_L g5014 ( 
.A(n_5000),
.B(n_4920),
.Y(n_5014)
);

INVx1_ASAP7_75t_L g5015 ( 
.A(n_4999),
.Y(n_5015)
);

OAI32xp33_ASAP7_75t_L g5016 ( 
.A1(n_4989),
.A2(n_4926),
.A3(n_4798),
.B1(n_4801),
.B2(n_4811),
.Y(n_5016)
);

AOI22xp5_ASAP7_75t_L g5017 ( 
.A1(n_5004),
.A2(n_4878),
.B1(n_4717),
.B2(n_4629),
.Y(n_5017)
);

INVx1_ASAP7_75t_L g5018 ( 
.A(n_5002),
.Y(n_5018)
);

INVx1_ASAP7_75t_L g5019 ( 
.A(n_5007),
.Y(n_5019)
);

NAND2xp5_ASAP7_75t_L g5020 ( 
.A(n_5003),
.B(n_4949),
.Y(n_5020)
);

INVxp67_ASAP7_75t_SL g5021 ( 
.A(n_5011),
.Y(n_5021)
);

OAI22xp5_ASAP7_75t_L g5022 ( 
.A1(n_5010),
.A2(n_4805),
.B1(n_4716),
.B2(n_4715),
.Y(n_5022)
);

OR2x2_ASAP7_75t_L g5023 ( 
.A(n_5014),
.B(n_4946),
.Y(n_5023)
);

INVxp67_ASAP7_75t_L g5024 ( 
.A(n_5015),
.Y(n_5024)
);

AOI22xp33_ASAP7_75t_L g5025 ( 
.A1(n_5008),
.A2(n_4746),
.B1(n_4777),
.B2(n_4776),
.Y(n_5025)
);

HB1xp67_ASAP7_75t_L g5026 ( 
.A(n_5005),
.Y(n_5026)
);

AOI22xp33_ASAP7_75t_L g5027 ( 
.A1(n_5013),
.A2(n_4776),
.B1(n_4777),
.B2(n_4724),
.Y(n_5027)
);

INVx2_ASAP7_75t_SL g5028 ( 
.A(n_5012),
.Y(n_5028)
);

INVx1_ASAP7_75t_L g5029 ( 
.A(n_5009),
.Y(n_5029)
);

AND2x2_ASAP7_75t_L g5030 ( 
.A(n_5006),
.B(n_4846),
.Y(n_5030)
);

INVx1_ASAP7_75t_L g5031 ( 
.A(n_5016),
.Y(n_5031)
);

OAI221xp5_ASAP7_75t_L g5032 ( 
.A1(n_5001),
.A2(n_4993),
.B1(n_4996),
.B2(n_4907),
.C(n_4975),
.Y(n_5032)
);

OAI22xp5_ASAP7_75t_L g5033 ( 
.A1(n_5016),
.A2(n_4608),
.B1(n_4724),
.B2(n_4641),
.Y(n_5033)
);

INVxp67_ASAP7_75t_L g5034 ( 
.A(n_5007),
.Y(n_5034)
);

AOI22xp5_ASAP7_75t_L g5035 ( 
.A1(n_5004),
.A2(n_4637),
.B1(n_4876),
.B2(n_4846),
.Y(n_5035)
);

AND2x2_ASAP7_75t_L g5036 ( 
.A(n_5002),
.B(n_4954),
.Y(n_5036)
);

OA22x2_ASAP7_75t_L g5037 ( 
.A1(n_5017),
.A2(n_4937),
.B1(n_4840),
.B2(n_4823),
.Y(n_5037)
);

INVx1_ASAP7_75t_L g5038 ( 
.A(n_5036),
.Y(n_5038)
);

NAND2xp5_ASAP7_75t_L g5039 ( 
.A(n_5027),
.B(n_4937),
.Y(n_5039)
);

INVx1_ASAP7_75t_L g5040 ( 
.A(n_5026),
.Y(n_5040)
);

INVx1_ASAP7_75t_L g5041 ( 
.A(n_5033),
.Y(n_5041)
);

OAI22xp5_ASAP7_75t_L g5042 ( 
.A1(n_5035),
.A2(n_4919),
.B1(n_4726),
.B2(n_4739),
.Y(n_5042)
);

INVx1_ASAP7_75t_SL g5043 ( 
.A(n_5030),
.Y(n_5043)
);

OAI22xp33_ASAP7_75t_L g5044 ( 
.A1(n_5020),
.A2(n_4943),
.B1(n_4976),
.B2(n_4872),
.Y(n_5044)
);

NAND2xp5_ASAP7_75t_L g5045 ( 
.A(n_5025),
.B(n_4928),
.Y(n_5045)
);

NAND2xp5_ASAP7_75t_L g5046 ( 
.A(n_5018),
.B(n_4840),
.Y(n_5046)
);

AOI222xp33_ASAP7_75t_L g5047 ( 
.A1(n_5031),
.A2(n_4716),
.B1(n_4715),
.B2(n_4971),
.C1(n_4872),
.C2(n_4933),
.Y(n_5047)
);

INVx1_ASAP7_75t_L g5048 ( 
.A(n_5022),
.Y(n_5048)
);

INVx1_ASAP7_75t_L g5049 ( 
.A(n_5022),
.Y(n_5049)
);

AOI21xp5_ASAP7_75t_L g5050 ( 
.A1(n_5032),
.A2(n_4980),
.B(n_4943),
.Y(n_5050)
);

AOI22xp5_ASAP7_75t_L g5051 ( 
.A1(n_5034),
.A2(n_4917),
.B1(n_4875),
.B2(n_4843),
.Y(n_5051)
);

NAND2xp5_ASAP7_75t_L g5052 ( 
.A(n_5021),
.B(n_4948),
.Y(n_5052)
);

AND2x4_ASAP7_75t_L g5053 ( 
.A(n_5023),
.B(n_4948),
.Y(n_5053)
);

INVx1_ASAP7_75t_L g5054 ( 
.A(n_5019),
.Y(n_5054)
);

OAI21xp33_ASAP7_75t_L g5055 ( 
.A1(n_5029),
.A2(n_4918),
.B(n_4911),
.Y(n_5055)
);

INVx1_ASAP7_75t_L g5056 ( 
.A(n_5024),
.Y(n_5056)
);

INVx1_ASAP7_75t_L g5057 ( 
.A(n_5028),
.Y(n_5057)
);

AOI221xp5_ASAP7_75t_L g5058 ( 
.A1(n_5033),
.A2(n_4872),
.B1(n_4807),
.B2(n_4817),
.C(n_4819),
.Y(n_5058)
);

AOI21xp5_ASAP7_75t_L g5059 ( 
.A1(n_5032),
.A2(n_4980),
.B(n_4979),
.Y(n_5059)
);

INVx1_ASAP7_75t_L g5060 ( 
.A(n_5036),
.Y(n_5060)
);

OR2x2_ASAP7_75t_L g5061 ( 
.A(n_5020),
.B(n_4833),
.Y(n_5061)
);

NAND2xp5_ASAP7_75t_L g5062 ( 
.A(n_5036),
.B(n_4917),
.Y(n_5062)
);

AOI21xp5_ASAP7_75t_L g5063 ( 
.A1(n_5032),
.A2(n_4960),
.B(n_4988),
.Y(n_5063)
);

OAI221xp5_ASAP7_75t_L g5064 ( 
.A1(n_5058),
.A2(n_4922),
.B1(n_4833),
.B2(n_4924),
.C(n_4998),
.Y(n_5064)
);

AOI222xp33_ASAP7_75t_L g5065 ( 
.A1(n_5040),
.A2(n_4872),
.B1(n_4880),
.B2(n_4824),
.C1(n_4829),
.C2(n_4822),
.Y(n_5065)
);

AOI211xp5_ASAP7_75t_L g5066 ( 
.A1(n_5044),
.A2(n_4977),
.B(n_4916),
.C(n_4914),
.Y(n_5066)
);

AOI22xp5_ASAP7_75t_L g5067 ( 
.A1(n_5038),
.A2(n_4917),
.B1(n_4820),
.B2(n_4956),
.Y(n_5067)
);

AOI21xp33_ASAP7_75t_L g5068 ( 
.A1(n_5042),
.A2(n_4983),
.B(n_4994),
.Y(n_5068)
);

NAND2xp5_ASAP7_75t_L g5069 ( 
.A(n_5053),
.B(n_4950),
.Y(n_5069)
);

OAI21xp5_ASAP7_75t_SL g5070 ( 
.A1(n_5051),
.A2(n_4942),
.B(n_4880),
.Y(n_5070)
);

O2A1O1Ixp33_ASAP7_75t_L g5071 ( 
.A1(n_5062),
.A2(n_4956),
.B(n_4950),
.C(n_4941),
.Y(n_5071)
);

NAND3xp33_ASAP7_75t_L g5072 ( 
.A(n_5047),
.B(n_4941),
.C(n_4883),
.Y(n_5072)
);

AOI221x1_ASAP7_75t_L g5073 ( 
.A1(n_5050),
.A2(n_5059),
.B1(n_5055),
.B2(n_5063),
.C(n_5045),
.Y(n_5073)
);

INVx1_ASAP7_75t_L g5074 ( 
.A(n_5037),
.Y(n_5074)
);

NAND2xp5_ASAP7_75t_SL g5075 ( 
.A(n_5060),
.B(n_4883),
.Y(n_5075)
);

AND2x2_ASAP7_75t_L g5076 ( 
.A(n_5043),
.B(n_4751),
.Y(n_5076)
);

NAND2xp5_ASAP7_75t_L g5077 ( 
.A(n_5041),
.B(n_4751),
.Y(n_5077)
);

OAI21xp5_ASAP7_75t_L g5078 ( 
.A1(n_5046),
.A2(n_4886),
.B(n_4885),
.Y(n_5078)
);

INVx1_ASAP7_75t_L g5079 ( 
.A(n_5061),
.Y(n_5079)
);

AOI21xp33_ASAP7_75t_L g5080 ( 
.A1(n_5052),
.A2(n_4886),
.B(n_4885),
.Y(n_5080)
);

AOI22xp33_ASAP7_75t_SL g5081 ( 
.A1(n_5057),
.A2(n_4772),
.B1(n_4874),
.B2(n_4868),
.Y(n_5081)
);

AOI221xp5_ASAP7_75t_SL g5082 ( 
.A1(n_5039),
.A2(n_4874),
.B1(n_4868),
.B2(n_4763),
.C(n_4766),
.Y(n_5082)
);

OAI21xp5_ASAP7_75t_L g5083 ( 
.A1(n_5056),
.A2(n_4766),
.B(n_4763),
.Y(n_5083)
);

AOI21xp5_ASAP7_75t_L g5084 ( 
.A1(n_5054),
.A2(n_4754),
.B(n_4775),
.Y(n_5084)
);

AOI221xp5_ASAP7_75t_L g5085 ( 
.A1(n_5048),
.A2(n_4758),
.B1(n_4760),
.B2(n_4775),
.C(n_4754),
.Y(n_5085)
);

A2O1A1Ixp33_ASAP7_75t_L g5086 ( 
.A1(n_5049),
.A2(n_4775),
.B(n_4758),
.C(n_4760),
.Y(n_5086)
);

OAI32xp33_ASAP7_75t_L g5087 ( 
.A1(n_5061),
.A2(n_4726),
.A3(n_4737),
.B1(n_4739),
.B2(n_4672),
.Y(n_5087)
);

A2O1A1Ixp33_ASAP7_75t_L g5088 ( 
.A1(n_5050),
.A2(n_4777),
.B(n_4776),
.C(n_4672),
.Y(n_5088)
);

NOR2xp33_ASAP7_75t_L g5089 ( 
.A(n_5062),
.B(n_4505),
.Y(n_5089)
);

AOI22xp33_ASAP7_75t_L g5090 ( 
.A1(n_5053),
.A2(n_4729),
.B1(n_4722),
.B2(n_4755),
.Y(n_5090)
);

O2A1O1Ixp33_ASAP7_75t_SL g5091 ( 
.A1(n_5062),
.A2(n_4683),
.B(n_4737),
.C(n_4681),
.Y(n_5091)
);

AOI21xp33_ASAP7_75t_L g5092 ( 
.A1(n_5042),
.A2(n_4731),
.B(n_4730),
.Y(n_5092)
);

AOI221xp5_ASAP7_75t_L g5093 ( 
.A1(n_5044),
.A2(n_4773),
.B1(n_4769),
.B2(n_4767),
.C(n_4731),
.Y(n_5093)
);

NAND2xp5_ASAP7_75t_L g5094 ( 
.A(n_5053),
.B(n_4571),
.Y(n_5094)
);

AOI221xp5_ASAP7_75t_L g5095 ( 
.A1(n_5044),
.A2(n_4773),
.B1(n_4769),
.B2(n_4767),
.C(n_4731),
.Y(n_5095)
);

INVx1_ASAP7_75t_L g5096 ( 
.A(n_5062),
.Y(n_5096)
);

AOI22xp5_ASAP7_75t_L g5097 ( 
.A1(n_5089),
.A2(n_4608),
.B1(n_4755),
.B2(n_4722),
.Y(n_5097)
);

AOI22xp5_ASAP7_75t_L g5098 ( 
.A1(n_5079),
.A2(n_5096),
.B1(n_5094),
.B2(n_5076),
.Y(n_5098)
);

NOR2xp67_ASAP7_75t_L g5099 ( 
.A(n_5072),
.B(n_4664),
.Y(n_5099)
);

NAND2xp5_ASAP7_75t_SL g5100 ( 
.A(n_5090),
.B(n_4673),
.Y(n_5100)
);

OAI211xp5_ASAP7_75t_L g5101 ( 
.A1(n_5067),
.A2(n_4664),
.B(n_4666),
.C(n_4747),
.Y(n_5101)
);

OAI21xp33_ASAP7_75t_SL g5102 ( 
.A1(n_5065),
.A2(n_4729),
.B(n_4722),
.Y(n_5102)
);

AOI32xp33_ASAP7_75t_L g5103 ( 
.A1(n_5081),
.A2(n_4666),
.A3(n_4673),
.B1(n_4747),
.B2(n_4744),
.Y(n_5103)
);

NAND2xp5_ASAP7_75t_L g5104 ( 
.A(n_5088),
.B(n_4571),
.Y(n_5104)
);

AOI21xp5_ASAP7_75t_L g5105 ( 
.A1(n_5071),
.A2(n_4678),
.B(n_4730),
.Y(n_5105)
);

INVx1_ASAP7_75t_L g5106 ( 
.A(n_5069),
.Y(n_5106)
);

O2A1O1Ixp33_ASAP7_75t_SL g5107 ( 
.A1(n_5075),
.A2(n_4683),
.B(n_4749),
.C(n_4747),
.Y(n_5107)
);

OAI221xp5_ASAP7_75t_SL g5108 ( 
.A1(n_5070),
.A2(n_4749),
.B1(n_4744),
.B2(n_4735),
.C(n_4730),
.Y(n_5108)
);

OAI21xp33_ASAP7_75t_L g5109 ( 
.A1(n_5077),
.A2(n_4729),
.B(n_4755),
.Y(n_5109)
);

NAND4xp25_ASAP7_75t_L g5110 ( 
.A(n_5073),
.B(n_4749),
.C(n_4744),
.D(n_4735),
.Y(n_5110)
);

AOI221xp5_ASAP7_75t_L g5111 ( 
.A1(n_5087),
.A2(n_4735),
.B1(n_4668),
.B2(n_4662),
.C(n_4567),
.Y(n_5111)
);

OAI22x1_ASAP7_75t_L g5112 ( 
.A1(n_5074),
.A2(n_4574),
.B1(n_4655),
.B2(n_4610),
.Y(n_5112)
);

INVx2_ASAP7_75t_L g5113 ( 
.A(n_5064),
.Y(n_5113)
);

NAND2xp5_ASAP7_75t_L g5114 ( 
.A(n_5082),
.B(n_4655),
.Y(n_5114)
);

OAI22xp5_ASAP7_75t_L g5115 ( 
.A1(n_5066),
.A2(n_4610),
.B1(n_4611),
.B2(n_4668),
.Y(n_5115)
);

NAND4xp25_ASAP7_75t_L g5116 ( 
.A(n_5068),
.B(n_4692),
.C(n_4662),
.D(n_4648),
.Y(n_5116)
);

NAND2xp5_ASAP7_75t_L g5117 ( 
.A(n_5091),
.B(n_4574),
.Y(n_5117)
);

INVx1_ASAP7_75t_L g5118 ( 
.A(n_5078),
.Y(n_5118)
);

OAI22xp33_ASAP7_75t_L g5119 ( 
.A1(n_5083),
.A2(n_4611),
.B1(n_4701),
.B2(n_4505),
.Y(n_5119)
);

AOI21xp5_ASAP7_75t_L g5120 ( 
.A1(n_5084),
.A2(n_4505),
.B(n_4489),
.Y(n_5120)
);

AOI211xp5_ASAP7_75t_L g5121 ( 
.A1(n_5080),
.A2(n_4701),
.B(n_4505),
.C(n_4640),
.Y(n_5121)
);

NAND2xp33_ASAP7_75t_L g5122 ( 
.A(n_5086),
.B(n_4674),
.Y(n_5122)
);

OAI221xp5_ASAP7_75t_L g5123 ( 
.A1(n_5085),
.A2(n_4707),
.B1(n_4702),
.B2(n_4684),
.C(n_4649),
.Y(n_5123)
);

OAI211xp5_ASAP7_75t_L g5124 ( 
.A1(n_5092),
.A2(n_4705),
.B(n_4707),
.C(n_4702),
.Y(n_5124)
);

NAND3xp33_ASAP7_75t_SL g5125 ( 
.A(n_5120),
.B(n_5095),
.C(n_5093),
.Y(n_5125)
);

AOI221x1_ASAP7_75t_L g5126 ( 
.A1(n_5110),
.A2(n_4705),
.B1(n_4677),
.B2(n_4633),
.C(n_4671),
.Y(n_5126)
);

XNOR2x1_ASAP7_75t_L g5127 ( 
.A(n_5112),
.B(n_4649),
.Y(n_5127)
);

XNOR2x1_ASAP7_75t_L g5128 ( 
.A(n_5113),
.B(n_4634),
.Y(n_5128)
);

NOR2xp33_ASAP7_75t_L g5129 ( 
.A(n_5116),
.B(n_4634),
.Y(n_5129)
);

AO22x2_ASAP7_75t_L g5130 ( 
.A1(n_5106),
.A2(n_4677),
.B1(n_4671),
.B2(n_4669),
.Y(n_5130)
);

OAI221xp5_ASAP7_75t_L g5131 ( 
.A1(n_5103),
.A2(n_4684),
.B1(n_4679),
.B2(n_4669),
.C(n_4583),
.Y(n_5131)
);

INVx1_ASAP7_75t_SL g5132 ( 
.A(n_5117),
.Y(n_5132)
);

OR2x2_ASAP7_75t_L g5133 ( 
.A(n_5114),
.B(n_4640),
.Y(n_5133)
);

NOR2xp67_ASAP7_75t_L g5134 ( 
.A(n_5102),
.B(n_4699),
.Y(n_5134)
);

OAI322xp33_ASAP7_75t_L g5135 ( 
.A1(n_5100),
.A2(n_4679),
.A3(n_4577),
.B1(n_4573),
.B2(n_4511),
.C1(n_4483),
.C2(n_4493),
.Y(n_5135)
);

NAND3xp33_ASAP7_75t_L g5136 ( 
.A(n_5098),
.B(n_4699),
.C(n_4703),
.Y(n_5136)
);

AOI221xp5_ASAP7_75t_L g5137 ( 
.A1(n_5115),
.A2(n_4703),
.B1(n_4699),
.B2(n_4663),
.C(n_4660),
.Y(n_5137)
);

NAND3xp33_ASAP7_75t_L g5138 ( 
.A(n_5099),
.B(n_4699),
.C(n_4703),
.Y(n_5138)
);

AOI211x1_ASAP7_75t_L g5139 ( 
.A1(n_5101),
.A2(n_4663),
.B(n_4660),
.C(n_4674),
.Y(n_5139)
);

NAND2xp5_ASAP7_75t_L g5140 ( 
.A(n_5121),
.B(n_4616),
.Y(n_5140)
);

AOI22xp5_ASAP7_75t_L g5141 ( 
.A1(n_5097),
.A2(n_4703),
.B1(n_4676),
.B2(n_4616),
.Y(n_5141)
);

NAND2xp5_ASAP7_75t_L g5142 ( 
.A(n_5109),
.B(n_4620),
.Y(n_5142)
);

OAI221xp5_ASAP7_75t_L g5143 ( 
.A1(n_5111),
.A2(n_4620),
.B1(n_4609),
.B2(n_4513),
.C(n_4506),
.Y(n_5143)
);

AOI221xp5_ASAP7_75t_L g5144 ( 
.A1(n_5119),
.A2(n_4676),
.B1(n_4609),
.B2(n_4562),
.C(n_4542),
.Y(n_5144)
);

NAND2xp5_ASAP7_75t_L g5145 ( 
.A(n_5139),
.B(n_5105),
.Y(n_5145)
);

INVx2_ASAP7_75t_L g5146 ( 
.A(n_5133),
.Y(n_5146)
);

OR2x2_ASAP7_75t_L g5147 ( 
.A(n_5138),
.B(n_5104),
.Y(n_5147)
);

OAI211xp5_ASAP7_75t_L g5148 ( 
.A1(n_5125),
.A2(n_5118),
.B(n_5124),
.C(n_5107),
.Y(n_5148)
);

OAI21xp33_ASAP7_75t_SL g5149 ( 
.A1(n_5141),
.A2(n_5134),
.B(n_5144),
.Y(n_5149)
);

INVx1_ASAP7_75t_L g5150 ( 
.A(n_5136),
.Y(n_5150)
);

INVx1_ASAP7_75t_L g5151 ( 
.A(n_5142),
.Y(n_5151)
);

NAND2xp5_ASAP7_75t_SL g5152 ( 
.A(n_5140),
.B(n_5122),
.Y(n_5152)
);

AOI21xp5_ASAP7_75t_L g5153 ( 
.A1(n_5129),
.A2(n_5132),
.B(n_5127),
.Y(n_5153)
);

NOR3xp33_ASAP7_75t_L g5154 ( 
.A(n_5131),
.B(n_5108),
.C(n_5123),
.Y(n_5154)
);

NOR2xp67_ASAP7_75t_L g5155 ( 
.A(n_5143),
.B(n_650),
.Y(n_5155)
);

INVx1_ASAP7_75t_L g5156 ( 
.A(n_5130),
.Y(n_5156)
);

NAND2x1p5_ASAP7_75t_SL g5157 ( 
.A(n_5128),
.B(n_4562),
.Y(n_5157)
);

NAND3xp33_ASAP7_75t_L g5158 ( 
.A(n_5137),
.B(n_4542),
.C(n_4513),
.Y(n_5158)
);

NOR3xp33_ASAP7_75t_L g5159 ( 
.A(n_5135),
.B(n_4556),
.C(n_4525),
.Y(n_5159)
);

NOR3xp33_ASAP7_75t_L g5160 ( 
.A(n_5130),
.B(n_4568),
.C(n_4546),
.Y(n_5160)
);

NAND5xp2_ASAP7_75t_L g5161 ( 
.A(n_5126),
.B(n_4597),
.C(n_4546),
.D(n_4590),
.E(n_4566),
.Y(n_5161)
);

NAND4xp25_ASAP7_75t_L g5162 ( 
.A(n_5129),
.B(n_4650),
.C(n_4566),
.D(n_4569),
.Y(n_5162)
);

NOR2xp33_ASAP7_75t_SL g5163 ( 
.A(n_5150),
.B(n_4547),
.Y(n_5163)
);

NOR4xp25_ASAP7_75t_L g5164 ( 
.A(n_5148),
.B(n_4547),
.C(n_4480),
.D(n_4493),
.Y(n_5164)
);

NAND3xp33_ASAP7_75t_SL g5165 ( 
.A(n_5154),
.B(n_4597),
.C(n_4650),
.Y(n_5165)
);

NAND4xp75_ASAP7_75t_L g5166 ( 
.A(n_5149),
.B(n_4526),
.C(n_4656),
.D(n_4548),
.Y(n_5166)
);

OR2x2_ASAP7_75t_L g5167 ( 
.A(n_5161),
.B(n_4483),
.Y(n_5167)
);

NOR4xp25_ASAP7_75t_L g5168 ( 
.A(n_5152),
.B(n_4656),
.C(n_4551),
.D(n_4654),
.Y(n_5168)
);

NAND5xp2_ASAP7_75t_L g5169 ( 
.A(n_5153),
.B(n_4586),
.C(n_4579),
.D(n_4654),
.E(n_4472),
.Y(n_5169)
);

NAND2xp5_ASAP7_75t_SL g5170 ( 
.A(n_5146),
.B(n_4532),
.Y(n_5170)
);

NOR3xp33_ASAP7_75t_L g5171 ( 
.A(n_5145),
.B(n_4595),
.C(n_4553),
.Y(n_5171)
);

O2A1O1Ixp33_ASAP7_75t_L g5172 ( 
.A1(n_5156),
.A2(n_4526),
.B(n_4555),
.C(n_4592),
.Y(n_5172)
);

NOR2x1_ASAP7_75t_L g5173 ( 
.A(n_5147),
.B(n_4555),
.Y(n_5173)
);

NAND4xp25_ASAP7_75t_L g5174 ( 
.A(n_5155),
.B(n_4472),
.C(n_4548),
.D(n_4586),
.Y(n_5174)
);

NOR3xp33_ASAP7_75t_L g5175 ( 
.A(n_5151),
.B(n_4576),
.C(n_4561),
.Y(n_5175)
);

NAND4xp25_ASAP7_75t_L g5176 ( 
.A(n_5160),
.B(n_4532),
.C(n_4576),
.D(n_4561),
.Y(n_5176)
);

NAND3xp33_ASAP7_75t_L g5177 ( 
.A(n_5159),
.B(n_5158),
.C(n_5162),
.Y(n_5177)
);

NAND3xp33_ASAP7_75t_SL g5178 ( 
.A(n_5157),
.B(n_4524),
.C(n_4527),
.Y(n_5178)
);

INVx1_ASAP7_75t_L g5179 ( 
.A(n_5157),
.Y(n_5179)
);

NAND3xp33_ASAP7_75t_L g5180 ( 
.A(n_5154),
.B(n_4526),
.C(n_4524),
.Y(n_5180)
);

NAND3xp33_ASAP7_75t_L g5181 ( 
.A(n_5154),
.B(n_4527),
.C(n_4544),
.Y(n_5181)
);

INVx1_ASAP7_75t_L g5182 ( 
.A(n_5165),
.Y(n_5182)
);

INVxp67_ASAP7_75t_L g5183 ( 
.A(n_5163),
.Y(n_5183)
);

INVx1_ASAP7_75t_L g5184 ( 
.A(n_5167),
.Y(n_5184)
);

AND2x2_ASAP7_75t_L g5185 ( 
.A(n_5175),
.B(n_4486),
.Y(n_5185)
);

INVx2_ASAP7_75t_L g5186 ( 
.A(n_5166),
.Y(n_5186)
);

NOR2xp33_ASAP7_75t_L g5187 ( 
.A(n_5170),
.B(n_4555),
.Y(n_5187)
);

INVx2_ASAP7_75t_L g5188 ( 
.A(n_5179),
.Y(n_5188)
);

INVx2_ASAP7_75t_L g5189 ( 
.A(n_5181),
.Y(n_5189)
);

INVx2_ASAP7_75t_L g5190 ( 
.A(n_5180),
.Y(n_5190)
);

NAND2xp5_ASAP7_75t_L g5191 ( 
.A(n_5164),
.B(n_4539),
.Y(n_5191)
);

INVx1_ASAP7_75t_L g5192 ( 
.A(n_5171),
.Y(n_5192)
);

INVx2_ASAP7_75t_L g5193 ( 
.A(n_5177),
.Y(n_5193)
);

NOR2x1_ASAP7_75t_L g5194 ( 
.A(n_5174),
.B(n_4471),
.Y(n_5194)
);

AO22x2_ASAP7_75t_L g5195 ( 
.A1(n_5178),
.A2(n_4543),
.B1(n_4550),
.B2(n_4475),
.Y(n_5195)
);

AO22x2_ASAP7_75t_L g5196 ( 
.A1(n_5168),
.A2(n_4486),
.B1(n_4478),
.B2(n_4501),
.Y(n_5196)
);

AND2x4_ASAP7_75t_L g5197 ( 
.A(n_5173),
.B(n_4485),
.Y(n_5197)
);

INVxp67_ASAP7_75t_SL g5198 ( 
.A(n_5176),
.Y(n_5198)
);

NOR2x1_ASAP7_75t_L g5199 ( 
.A(n_5169),
.B(n_4591),
.Y(n_5199)
);

NOR3xp33_ASAP7_75t_SL g5200 ( 
.A(n_5182),
.B(n_5172),
.C(n_652),
.Y(n_5200)
);

AND2x4_ASAP7_75t_L g5201 ( 
.A(n_5183),
.B(n_4521),
.Y(n_5201)
);

NOR4xp75_ASAP7_75t_L g5202 ( 
.A(n_5191),
.B(n_4584),
.C(n_4589),
.D(n_4487),
.Y(n_5202)
);

NOR3xp33_ASAP7_75t_SL g5203 ( 
.A(n_5184),
.B(n_651),
.C(n_652),
.Y(n_5203)
);

AND2x4_ASAP7_75t_L g5204 ( 
.A(n_5198),
.B(n_5189),
.Y(n_5204)
);

AND3x2_ASAP7_75t_L g5205 ( 
.A(n_5186),
.B(n_4576),
.C(n_4561),
.Y(n_5205)
);

NAND3xp33_ASAP7_75t_SL g5206 ( 
.A(n_5188),
.B(n_4537),
.C(n_4523),
.Y(n_5206)
);

INVx1_ASAP7_75t_L g5207 ( 
.A(n_5196),
.Y(n_5207)
);

NAND2xp5_ASAP7_75t_L g5208 ( 
.A(n_5199),
.B(n_4500),
.Y(n_5208)
);

INVxp67_ASAP7_75t_L g5209 ( 
.A(n_5190),
.Y(n_5209)
);

NOR3xp33_ASAP7_75t_SL g5210 ( 
.A(n_5192),
.B(n_651),
.C(n_653),
.Y(n_5210)
);

AND2x4_ASAP7_75t_L g5211 ( 
.A(n_5194),
.B(n_4491),
.Y(n_5211)
);

NAND4xp25_ASAP7_75t_L g5212 ( 
.A(n_5209),
.B(n_5193),
.C(n_5204),
.D(n_5201),
.Y(n_5212)
);

HB1xp67_ASAP7_75t_L g5213 ( 
.A(n_5208),
.Y(n_5213)
);

AOI22xp5_ASAP7_75t_L g5214 ( 
.A1(n_5211),
.A2(n_5185),
.B1(n_5187),
.B2(n_5197),
.Y(n_5214)
);

NOR2x1_ASAP7_75t_L g5215 ( 
.A(n_5207),
.B(n_5195),
.Y(n_5215)
);

INVx1_ASAP7_75t_L g5216 ( 
.A(n_5210),
.Y(n_5216)
);

AND2x4_ASAP7_75t_L g5217 ( 
.A(n_5203),
.B(n_5195),
.Y(n_5217)
);

INVx2_ASAP7_75t_L g5218 ( 
.A(n_5205),
.Y(n_5218)
);

INVx2_ASAP7_75t_L g5219 ( 
.A(n_5218),
.Y(n_5219)
);

INVx1_ASAP7_75t_L g5220 ( 
.A(n_5217),
.Y(n_5220)
);

INVx1_ASAP7_75t_L g5221 ( 
.A(n_5215),
.Y(n_5221)
);

INVx1_ASAP7_75t_L g5222 ( 
.A(n_5221),
.Y(n_5222)
);

INVx1_ASAP7_75t_SL g5223 ( 
.A(n_5219),
.Y(n_5223)
);

XNOR2x1_ASAP7_75t_L g5224 ( 
.A(n_5223),
.B(n_5220),
.Y(n_5224)
);

AND2x2_ASAP7_75t_SL g5225 ( 
.A(n_5224),
.B(n_5222),
.Y(n_5225)
);

AOI22x1_ASAP7_75t_L g5226 ( 
.A1(n_5225),
.A2(n_5213),
.B1(n_5216),
.B2(n_5212),
.Y(n_5226)
);

AOI22xp5_ASAP7_75t_L g5227 ( 
.A1(n_5226),
.A2(n_5214),
.B1(n_5200),
.B2(n_5206),
.Y(n_5227)
);

NAND2xp5_ASAP7_75t_L g5228 ( 
.A(n_5227),
.B(n_5202),
.Y(n_5228)
);

OAI22xp5_ASAP7_75t_SL g5229 ( 
.A1(n_5228),
.A2(n_4565),
.B1(n_4593),
.B2(n_655),
.Y(n_5229)
);

AOI21xp33_ASAP7_75t_L g5230 ( 
.A1(n_5229),
.A2(n_653),
.B(n_654),
.Y(n_5230)
);

AND2x2_ASAP7_75t_SL g5231 ( 
.A(n_5230),
.B(n_4599),
.Y(n_5231)
);

NAND3xp33_ASAP7_75t_L g5232 ( 
.A(n_5231),
.B(n_654),
.C(n_655),
.Y(n_5232)
);

INVx1_ASAP7_75t_L g5233 ( 
.A(n_5232),
.Y(n_5233)
);

OR2x6_ASAP7_75t_L g5234 ( 
.A(n_5233),
.B(n_4495),
.Y(n_5234)
);

OAI221xp5_ASAP7_75t_R g5235 ( 
.A1(n_5234),
.A2(n_657),
.B1(n_658),
.B2(n_659),
.C(n_660),
.Y(n_5235)
);

AOI21xp5_ASAP7_75t_L g5236 ( 
.A1(n_5235),
.A2(n_4588),
.B(n_4559),
.Y(n_5236)
);

AOI211xp5_ASAP7_75t_L g5237 ( 
.A1(n_5236),
.A2(n_660),
.B(n_661),
.C(n_663),
.Y(n_5237)
);


endmodule