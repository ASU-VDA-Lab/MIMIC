module fake_jpeg_11263_n_525 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_525);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_525;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx3_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_17),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_12),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_6),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_16),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_17),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_11),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_1),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_15),
.Y(n_34)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_11),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_10),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_4),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_4),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_10),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_2),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_10),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_14),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_5),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_10),
.Y(n_44)
);

CKINVDCx16_ASAP7_75t_R g45 ( 
.A(n_5),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_1),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_15),
.Y(n_47)
);

INVx11_ASAP7_75t_L g48 ( 
.A(n_6),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_13),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_11),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_12),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_13),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_21),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_53),
.Y(n_110)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_27),
.Y(n_54)
);

INVx5_ASAP7_75t_L g159 ( 
.A(n_54),
.Y(n_159)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_29),
.Y(n_55)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_55),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_21),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_56),
.Y(n_121)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_27),
.Y(n_57)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_57),
.Y(n_111)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_29),
.Y(n_58)
);

BUFx12f_ASAP7_75t_L g147 ( 
.A(n_58),
.Y(n_147)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_29),
.Y(n_59)
);

INVx5_ASAP7_75t_L g160 ( 
.A(n_59),
.Y(n_160)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_19),
.Y(n_60)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_60),
.Y(n_108)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_19),
.Y(n_61)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_61),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_27),
.B(n_17),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_62),
.B(n_71),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_21),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_63),
.Y(n_134)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_52),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g149 ( 
.A(n_64),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_21),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g158 ( 
.A(n_65),
.Y(n_158)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_26),
.Y(n_66)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_66),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_24),
.Y(n_67)
);

INVx6_ASAP7_75t_L g129 ( 
.A(n_67),
.Y(n_129)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_27),
.Y(n_68)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_68),
.Y(n_107)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_27),
.Y(n_69)
);

INVx4_ASAP7_75t_L g119 ( 
.A(n_69),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_24),
.Y(n_70)
);

INVx6_ASAP7_75t_L g133 ( 
.A(n_70),
.Y(n_133)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_26),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_30),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_72),
.B(n_74),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_24),
.Y(n_73)
);

INVx6_ASAP7_75t_L g135 ( 
.A(n_73),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_22),
.B(n_0),
.Y(n_74)
);

BUFx3_ASAP7_75t_L g75 ( 
.A(n_18),
.Y(n_75)
);

BUFx3_ASAP7_75t_L g125 ( 
.A(n_75),
.Y(n_125)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_30),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_76),
.B(n_84),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_24),
.Y(n_77)
);

INVx6_ASAP7_75t_L g155 ( 
.A(n_77),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_28),
.Y(n_78)
);

INVx8_ASAP7_75t_L g131 ( 
.A(n_78),
.Y(n_131)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_18),
.Y(n_79)
);

BUFx3_ASAP7_75t_L g126 ( 
.A(n_79),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_28),
.Y(n_80)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_80),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_28),
.Y(n_81)
);

INVx3_ASAP7_75t_L g136 ( 
.A(n_81),
.Y(n_136)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_18),
.Y(n_82)
);

INVx3_ASAP7_75t_L g137 ( 
.A(n_82),
.Y(n_137)
);

BUFx3_ASAP7_75t_L g83 ( 
.A(n_33),
.Y(n_83)
);

INVx4_ASAP7_75t_L g124 ( 
.A(n_83),
.Y(n_124)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_42),
.Y(n_84)
);

BUFx2_ASAP7_75t_L g85 ( 
.A(n_28),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_85),
.Y(n_130)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_33),
.Y(n_86)
);

INVx3_ASAP7_75t_L g143 ( 
.A(n_86),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_39),
.Y(n_87)
);

INVx3_ASAP7_75t_L g144 ( 
.A(n_87),
.Y(n_144)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_33),
.Y(n_88)
);

INVx4_ASAP7_75t_L g156 ( 
.A(n_88),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_39),
.Y(n_89)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_89),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_39),
.Y(n_90)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_90),
.Y(n_113)
);

INVx6_ASAP7_75t_L g91 ( 
.A(n_52),
.Y(n_91)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_91),
.Y(n_115)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_34),
.Y(n_92)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_92),
.Y(n_116)
);

BUFx3_ASAP7_75t_L g93 ( 
.A(n_37),
.Y(n_93)
);

INVx2_ASAP7_75t_SL g153 ( 
.A(n_93),
.Y(n_153)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_34),
.Y(n_94)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_94),
.Y(n_120)
);

INVx8_ASAP7_75t_L g95 ( 
.A(n_32),
.Y(n_95)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_95),
.Y(n_128)
);

INVx8_ASAP7_75t_L g96 ( 
.A(n_32),
.Y(n_96)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_96),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_39),
.Y(n_97)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_97),
.Y(n_146)
);

INVx11_ASAP7_75t_L g98 ( 
.A(n_48),
.Y(n_98)
);

CKINVDCx14_ASAP7_75t_R g132 ( 
.A(n_98),
.Y(n_132)
);

INVx5_ASAP7_75t_L g99 ( 
.A(n_37),
.Y(n_99)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_99),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_40),
.Y(n_100)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_100),
.Y(n_151)
);

AND2x2_ASAP7_75t_L g101 ( 
.A(n_38),
.B(n_0),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_101),
.B(n_102),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_22),
.B(n_1),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_48),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_103),
.B(n_45),
.Y(n_105)
);

NAND3xp33_ASAP7_75t_L g180 ( 
.A(n_105),
.B(n_122),
.C(n_45),
.Y(n_180)
);

OAI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_85),
.A2(n_38),
.B1(n_32),
.B2(n_50),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_106),
.A2(n_139),
.B1(n_100),
.B2(n_90),
.Y(n_171)
);

OR2x2_ASAP7_75t_L g112 ( 
.A(n_55),
.B(n_42),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_112),
.B(n_117),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_101),
.B(n_25),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_114),
.B(n_127),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_95),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_75),
.B(n_25),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_64),
.B(n_23),
.Y(n_127)
);

INVx13_ASAP7_75t_L g138 ( 
.A(n_79),
.Y(n_138)
);

INVx13_ASAP7_75t_L g169 ( 
.A(n_138),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_91),
.A2(n_20),
.B1(n_35),
.B2(n_47),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_58),
.A2(n_20),
.B1(n_35),
.B2(n_37),
.Y(n_145)
);

CKINVDCx16_ASAP7_75t_R g176 ( 
.A(n_145),
.Y(n_176)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_53),
.Y(n_157)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_157),
.Y(n_174)
);

AOI22xp33_ASAP7_75t_L g161 ( 
.A1(n_56),
.A2(n_35),
.B1(n_20),
.B2(n_52),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_161),
.A2(n_47),
.B1(n_40),
.B2(n_50),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_152),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_162),
.B(n_170),
.Y(n_220)
);

OA22x2_ASAP7_75t_L g163 ( 
.A1(n_161),
.A2(n_96),
.B1(n_59),
.B2(n_97),
.Y(n_163)
);

O2A1O1Ixp33_ASAP7_75t_L g254 ( 
.A1(n_163),
.A2(n_173),
.B(n_208),
.C(n_121),
.Y(n_254)
);

BUFx3_ASAP7_75t_L g164 ( 
.A(n_147),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g247 ( 
.A(n_164),
.Y(n_247)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_115),
.Y(n_165)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_165),
.Y(n_233)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_109),
.Y(n_166)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_166),
.Y(n_238)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_113),
.Y(n_167)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_167),
.Y(n_246)
);

INVx1_ASAP7_75t_SL g168 ( 
.A(n_147),
.Y(n_168)
);

AND2x2_ASAP7_75t_L g228 ( 
.A(n_168),
.B(n_171),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_152),
.Y(n_170)
);

AOI22xp33_ASAP7_75t_SL g172 ( 
.A1(n_108),
.A2(n_48),
.B1(n_44),
.B2(n_43),
.Y(n_172)
);

INVxp67_ASAP7_75t_L g243 ( 
.A(n_172),
.Y(n_243)
);

AOI21xp5_ASAP7_75t_L g173 ( 
.A1(n_112),
.A2(n_44),
.B(n_31),
.Y(n_173)
);

INVx3_ASAP7_75t_L g175 ( 
.A(n_128),
.Y(n_175)
);

BUFx2_ASAP7_75t_L g251 ( 
.A(n_175),
.Y(n_251)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_146),
.Y(n_177)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_177),
.Y(n_227)
);

INVx3_ASAP7_75t_SL g178 ( 
.A(n_131),
.Y(n_178)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_178),
.Y(n_232)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_140),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_179),
.B(n_180),
.Y(n_221)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_148),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_181),
.B(n_183),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_154),
.B(n_41),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_182),
.B(n_200),
.Y(n_225)
);

CKINVDCx16_ASAP7_75t_R g183 ( 
.A(n_138),
.Y(n_183)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_151),
.Y(n_184)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_184),
.Y(n_245)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_116),
.Y(n_185)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_185),
.Y(n_253)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_120),
.Y(n_186)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_186),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_141),
.B(n_41),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_187),
.B(n_190),
.Y(n_235)
);

INVx4_ASAP7_75t_L g188 ( 
.A(n_147),
.Y(n_188)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_188),
.Y(n_256)
);

INVx1_ASAP7_75t_SL g189 ( 
.A(n_104),
.Y(n_189)
);

AND2x2_ASAP7_75t_L g231 ( 
.A(n_189),
.B(n_192),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_141),
.B(n_46),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_191),
.A2(n_214),
.B1(n_63),
.B2(n_78),
.Y(n_218)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_123),
.Y(n_192)
);

CKINVDCx16_ASAP7_75t_R g193 ( 
.A(n_132),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_193),
.B(n_197),
.Y(n_239)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_136),
.Y(n_195)
);

AND2x2_ASAP7_75t_L g248 ( 
.A(n_195),
.B(n_198),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_118),
.B(n_93),
.Y(n_196)
);

INVxp67_ASAP7_75t_L g260 ( 
.A(n_196),
.Y(n_260)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_137),
.Y(n_197)
);

INVx2_ASAP7_75t_SL g198 ( 
.A(n_159),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_143),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_199),
.B(n_201),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_154),
.B(n_49),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_142),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_118),
.B(n_83),
.Y(n_202)
);

INVxp67_ASAP7_75t_L g263 ( 
.A(n_202),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_107),
.B(n_46),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_203),
.B(n_205),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_131),
.B(n_36),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_204),
.B(n_51),
.Y(n_249)
);

CKINVDCx14_ASAP7_75t_R g205 ( 
.A(n_153),
.Y(n_205)
);

BUFx6f_ASAP7_75t_L g207 ( 
.A(n_110),
.Y(n_207)
);

AOI22xp33_ASAP7_75t_SL g223 ( 
.A1(n_207),
.A2(n_213),
.B1(n_129),
.B2(n_155),
.Y(n_223)
);

OA22x2_ASAP7_75t_L g208 ( 
.A1(n_106),
.A2(n_89),
.B1(n_87),
.B2(n_81),
.Y(n_208)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_144),
.Y(n_209)
);

AND2x2_ASAP7_75t_L g264 ( 
.A(n_209),
.B(n_210),
.Y(n_264)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_153),
.Y(n_210)
);

CKINVDCx16_ASAP7_75t_R g211 ( 
.A(n_132),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_211),
.B(n_212),
.Y(n_252)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_149),
.Y(n_212)
);

INVx5_ASAP7_75t_L g213 ( 
.A(n_124),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_L g214 ( 
.A1(n_129),
.A2(n_20),
.B1(n_65),
.B2(n_70),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_119),
.B(n_23),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_215),
.B(n_31),
.Y(n_226)
);

INVx4_ASAP7_75t_L g216 ( 
.A(n_160),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_216),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_176),
.A2(n_126),
.B1(n_125),
.B2(n_150),
.Y(n_217)
);

OAI21xp5_ASAP7_75t_SL g292 ( 
.A1(n_217),
.A2(n_234),
.B(n_241),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_L g279 ( 
.A1(n_218),
.A2(n_178),
.B1(n_207),
.B2(n_184),
.Y(n_279)
);

XNOR2x1_ASAP7_75t_SL g219 ( 
.A(n_206),
.B(n_156),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_219),
.B(n_167),
.Y(n_282)
);

INVxp67_ASAP7_75t_L g278 ( 
.A(n_223),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_171),
.A2(n_67),
.B1(n_80),
.B2(n_77),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_224),
.A2(n_236),
.B1(n_237),
.B2(n_240),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_SL g303 ( 
.A(n_226),
.B(n_249),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_182),
.B(n_111),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_229),
.B(n_14),
.C(n_15),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_204),
.A2(n_130),
.B1(n_43),
.B2(n_133),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_208),
.A2(n_73),
.B1(n_149),
.B2(n_155),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_208),
.A2(n_135),
.B1(n_133),
.B2(n_134),
.Y(n_237)
);

OAI22xp33_ASAP7_75t_SL g240 ( 
.A1(n_173),
.A2(n_158),
.B1(n_110),
.B2(n_134),
.Y(n_240)
);

NAND3xp33_ASAP7_75t_SL g241 ( 
.A(n_200),
.B(n_36),
.C(n_49),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_208),
.A2(n_135),
.B1(n_158),
.B2(n_121),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_250),
.A2(n_257),
.B1(n_258),
.B2(n_40),
.Y(n_283)
);

AND2x2_ASAP7_75t_L g297 ( 
.A(n_254),
.B(n_8),
.Y(n_297)
);

OAI22xp33_ASAP7_75t_SL g257 ( 
.A1(n_194),
.A2(n_43),
.B1(n_50),
.B2(n_47),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_163),
.A2(n_52),
.B1(n_50),
.B2(n_47),
.Y(n_258)
);

AOI22xp33_ASAP7_75t_L g259 ( 
.A1(n_163),
.A2(n_212),
.B1(n_185),
.B2(n_186),
.Y(n_259)
);

OA22x2_ASAP7_75t_L g285 ( 
.A1(n_259),
.A2(n_40),
.B1(n_3),
.B2(n_4),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_165),
.B(n_51),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_261),
.B(n_174),
.Y(n_274)
);

A2O1A1Ixp33_ASAP7_75t_L g262 ( 
.A1(n_163),
.A2(n_1),
.B(n_2),
.C(n_3),
.Y(n_262)
);

O2A1O1Ixp33_ASAP7_75t_SL g290 ( 
.A1(n_262),
.A2(n_16),
.B(n_6),
.C(n_7),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_244),
.B(n_210),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_SL g343 ( 
.A(n_265),
.B(n_267),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_244),
.B(n_189),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_264),
.Y(n_268)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_268),
.Y(n_311)
);

AOI21xp33_ASAP7_75t_SL g269 ( 
.A1(n_219),
.A2(n_169),
.B(n_216),
.Y(n_269)
);

OAI21xp5_ASAP7_75t_SL g324 ( 
.A1(n_269),
.A2(n_293),
.B(n_297),
.Y(n_324)
);

FAx1_ASAP7_75t_SL g270 ( 
.A(n_225),
.B(n_169),
.CI(n_175),
.CON(n_270),
.SN(n_270)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_270),
.B(n_271),
.Y(n_334)
);

CKINVDCx14_ASAP7_75t_R g271 ( 
.A(n_230),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_220),
.B(n_213),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_SL g333 ( 
.A(n_272),
.B(n_274),
.Y(n_333)
);

AOI22xp33_ASAP7_75t_L g273 ( 
.A1(n_228),
.A2(n_209),
.B1(n_192),
.B2(n_195),
.Y(n_273)
);

AOI22xp33_ASAP7_75t_SL g344 ( 
.A1(n_273),
.A2(n_280),
.B1(n_287),
.B2(n_295),
.Y(n_344)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_264),
.Y(n_275)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_275),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_229),
.B(n_166),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_276),
.B(n_301),
.Y(n_323)
);

OAI21xp5_ASAP7_75t_L g277 ( 
.A1(n_243),
.A2(n_168),
.B(n_164),
.Y(n_277)
);

OAI21xp5_ASAP7_75t_L g317 ( 
.A1(n_277),
.A2(n_300),
.B(n_269),
.Y(n_317)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_279),
.Y(n_319)
);

AOI22xp33_ASAP7_75t_SL g280 ( 
.A1(n_237),
.A2(n_188),
.B1(n_198),
.B2(n_177),
.Y(n_280)
);

BUFx6f_ASAP7_75t_L g281 ( 
.A(n_247),
.Y(n_281)
);

INVx4_ASAP7_75t_L g309 ( 
.A(n_281),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_SL g310 ( 
.A(n_282),
.B(n_302),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_SL g312 ( 
.A1(n_283),
.A2(n_298),
.B1(n_299),
.B2(n_218),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_264),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_284),
.B(n_290),
.Y(n_340)
);

INVx1_ASAP7_75t_SL g318 ( 
.A(n_285),
.Y(n_318)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_253),
.Y(n_286)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_286),
.Y(n_321)
);

AOI22xp33_ASAP7_75t_SL g287 ( 
.A1(n_250),
.A2(n_2),
.B1(n_5),
.B2(n_6),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_253),
.Y(n_288)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_288),
.Y(n_322)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_233),
.Y(n_289)
);

INVx2_ASAP7_75t_L g308 ( 
.A(n_289),
.Y(n_308)
);

HB1xp67_ASAP7_75t_L g291 ( 
.A(n_233),
.Y(n_291)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_291),
.Y(n_325)
);

OA21x2_ASAP7_75t_L g293 ( 
.A1(n_258),
.A2(n_5),
.B(n_7),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_255),
.Y(n_294)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_294),
.Y(n_331)
);

AOI22xp33_ASAP7_75t_SL g295 ( 
.A1(n_260),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_295)
);

INVxp67_ASAP7_75t_L g296 ( 
.A(n_248),
.Y(n_296)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_296),
.Y(n_338)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_254),
.A2(n_8),
.B1(n_9),
.B2(n_11),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_L g299 ( 
.A1(n_254),
.A2(n_9),
.B1(n_12),
.B2(n_13),
.Y(n_299)
);

AOI22xp33_ASAP7_75t_SL g300 ( 
.A1(n_263),
.A2(n_9),
.B1(n_12),
.B2(n_14),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_259),
.A2(n_16),
.B1(n_14),
.B2(n_15),
.Y(n_301)
);

INVx2_ASAP7_75t_L g304 ( 
.A(n_251),
.Y(n_304)
);

INVx2_ASAP7_75t_L g337 ( 
.A(n_304),
.Y(n_337)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_255),
.Y(n_305)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_305),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_220),
.B(n_16),
.Y(n_306)
);

NAND3xp33_ASAP7_75t_L g328 ( 
.A(n_306),
.B(n_221),
.C(n_226),
.Y(n_328)
);

INVxp67_ASAP7_75t_L g307 ( 
.A(n_248),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_307),
.B(n_231),
.Y(n_332)
);

AOI22xp5_ASAP7_75t_L g357 ( 
.A1(n_312),
.A2(n_315),
.B1(n_320),
.B2(n_336),
.Y(n_357)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_286),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g364 ( 
.A(n_313),
.B(n_327),
.Y(n_364)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_282),
.B(n_225),
.C(n_239),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g347 ( 
.A(n_314),
.B(n_326),
.C(n_329),
.Y(n_347)
);

OAI22xp5_ASAP7_75t_SL g315 ( 
.A1(n_266),
.A2(n_234),
.B1(n_228),
.B2(n_249),
.Y(n_315)
);

INVxp67_ASAP7_75t_L g361 ( 
.A(n_317),
.Y(n_361)
);

OAI22xp5_ASAP7_75t_SL g320 ( 
.A1(n_266),
.A2(n_228),
.B1(n_236),
.B2(n_217),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_276),
.B(n_239),
.C(n_252),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g327 ( 
.A(n_289),
.Y(n_327)
);

INVxp67_ASAP7_75t_L g372 ( 
.A(n_328),
.Y(n_372)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_296),
.B(n_252),
.C(n_230),
.Y(n_329)
);

XOR2xp5_ASAP7_75t_L g330 ( 
.A(n_274),
.B(n_242),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g367 ( 
.A(n_330),
.B(n_342),
.C(n_235),
.Y(n_367)
);

CKINVDCx14_ASAP7_75t_R g370 ( 
.A(n_332),
.Y(n_370)
);

CKINVDCx20_ASAP7_75t_R g335 ( 
.A(n_288),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_335),
.B(n_345),
.Y(n_365)
);

OAI22xp5_ASAP7_75t_SL g336 ( 
.A1(n_283),
.A2(n_262),
.B1(n_224),
.B2(n_261),
.Y(n_336)
);

MAJIxp5_ASAP7_75t_L g339 ( 
.A(n_307),
.B(n_242),
.C(n_256),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_L g350 ( 
.A(n_339),
.B(n_275),
.C(n_268),
.Y(n_350)
);

XOR2xp5_ASAP7_75t_L g342 ( 
.A(n_302),
.B(n_235),
.Y(n_342)
);

OAI22xp5_ASAP7_75t_SL g345 ( 
.A1(n_298),
.A2(n_262),
.B1(n_241),
.B2(n_232),
.Y(n_345)
);

OAI22xp5_ASAP7_75t_SL g346 ( 
.A1(n_299),
.A2(n_232),
.B1(n_222),
.B2(n_221),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_346),
.B(n_285),
.Y(n_366)
);

OAI21xp5_ASAP7_75t_L g348 ( 
.A1(n_334),
.A2(n_297),
.B(n_284),
.Y(n_348)
);

INVxp67_ASAP7_75t_L g389 ( 
.A(n_348),
.Y(n_389)
);

INVx1_ASAP7_75t_SL g349 ( 
.A(n_338),
.Y(n_349)
);

INVx2_ASAP7_75t_L g382 ( 
.A(n_349),
.Y(n_382)
);

MAJIxp5_ASAP7_75t_L g398 ( 
.A(n_350),
.B(n_358),
.C(n_379),
.Y(n_398)
);

NOR2xp33_ASAP7_75t_SL g351 ( 
.A(n_343),
.B(n_303),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_SL g399 ( 
.A(n_351),
.B(n_360),
.Y(n_399)
);

AOI21xp5_ASAP7_75t_L g352 ( 
.A1(n_340),
.A2(n_277),
.B(n_278),
.Y(n_352)
);

AOI21xp5_ASAP7_75t_L g395 ( 
.A1(n_352),
.A2(n_353),
.B(n_324),
.Y(n_395)
);

AOI21xp5_ASAP7_75t_L g353 ( 
.A1(n_317),
.A2(n_278),
.B(n_297),
.Y(n_353)
);

OAI22xp5_ASAP7_75t_SL g354 ( 
.A1(n_318),
.A2(n_293),
.B1(n_270),
.B2(n_285),
.Y(n_354)
);

AOI22xp5_ASAP7_75t_L g393 ( 
.A1(n_354),
.A2(n_355),
.B1(n_368),
.B2(n_377),
.Y(n_393)
);

OAI22xp5_ASAP7_75t_L g355 ( 
.A1(n_318),
.A2(n_270),
.B1(n_293),
.B2(n_285),
.Y(n_355)
);

CKINVDCx20_ASAP7_75t_R g356 ( 
.A(n_335),
.Y(n_356)
);

NOR2xp33_ASAP7_75t_L g392 ( 
.A(n_356),
.B(n_359),
.Y(n_392)
);

XOR2xp5_ASAP7_75t_L g358 ( 
.A(n_310),
.B(n_292),
.Y(n_358)
);

CKINVDCx20_ASAP7_75t_R g359 ( 
.A(n_333),
.Y(n_359)
);

CKINVDCx16_ASAP7_75t_R g360 ( 
.A(n_332),
.Y(n_360)
);

AOI22xp33_ASAP7_75t_SL g362 ( 
.A1(n_319),
.A2(n_281),
.B1(n_290),
.B2(n_292),
.Y(n_362)
);

OAI22xp5_ASAP7_75t_L g383 ( 
.A1(n_362),
.A2(n_344),
.B1(n_338),
.B2(n_316),
.Y(n_383)
);

CKINVDCx20_ASAP7_75t_R g363 ( 
.A(n_327),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_L g396 ( 
.A(n_363),
.B(n_378),
.Y(n_396)
);

HB1xp67_ASAP7_75t_L g381 ( 
.A(n_366),
.Y(n_381)
);

XNOR2xp5_ASAP7_75t_L g404 ( 
.A(n_367),
.B(n_331),
.Y(n_404)
);

OAI22xp5_ASAP7_75t_SL g368 ( 
.A1(n_319),
.A2(n_293),
.B1(n_303),
.B2(n_279),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_323),
.B(n_305),
.Y(n_369)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_369),
.Y(n_385)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_321),
.Y(n_371)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_371),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_323),
.B(n_294),
.Y(n_373)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_373),
.Y(n_387)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_321),
.Y(n_374)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_374),
.Y(n_394)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_322),
.Y(n_375)
);

INVxp67_ASAP7_75t_L g411 ( 
.A(n_375),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_311),
.B(n_304),
.Y(n_376)
);

XOR2x1_ASAP7_75t_L g406 ( 
.A(n_376),
.B(n_380),
.Y(n_406)
);

OAI22xp5_ASAP7_75t_SL g377 ( 
.A1(n_336),
.A2(n_301),
.B1(n_290),
.B2(n_222),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_322),
.Y(n_378)
);

MAJIxp5_ASAP7_75t_L g379 ( 
.A(n_310),
.B(n_256),
.C(n_245),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_311),
.B(n_227),
.Y(n_380)
);

AOI22xp5_ASAP7_75t_L g422 ( 
.A1(n_383),
.A2(n_397),
.B1(n_354),
.B2(n_361),
.Y(n_422)
);

XNOR2xp5_ASAP7_75t_SL g384 ( 
.A(n_358),
.B(n_314),
.Y(n_384)
);

XOR2xp5_ASAP7_75t_L g415 ( 
.A(n_384),
.B(n_386),
.Y(n_415)
);

XOR2xp5_ASAP7_75t_L g386 ( 
.A(n_358),
.B(n_326),
.Y(n_386)
);

XOR2xp5_ASAP7_75t_L g388 ( 
.A(n_347),
.B(n_339),
.Y(n_388)
);

XOR2xp5_ASAP7_75t_L g430 ( 
.A(n_388),
.B(n_402),
.Y(n_430)
);

OAI22xp5_ASAP7_75t_L g390 ( 
.A1(n_359),
.A2(n_312),
.B1(n_316),
.B2(n_345),
.Y(n_390)
);

CKINVDCx16_ASAP7_75t_R g413 ( 
.A(n_390),
.Y(n_413)
);

CKINVDCx20_ASAP7_75t_R g391 ( 
.A(n_380),
.Y(n_391)
);

NOR2xp33_ASAP7_75t_L g436 ( 
.A(n_391),
.B(n_403),
.Y(n_436)
);

OAI21xp5_ASAP7_75t_SL g417 ( 
.A1(n_395),
.A2(n_352),
.B(n_353),
.Y(n_417)
);

OAI22x1_ASAP7_75t_SL g397 ( 
.A1(n_357),
.A2(n_324),
.B1(n_320),
.B2(n_315),
.Y(n_397)
);

AOI22xp5_ASAP7_75t_L g400 ( 
.A1(n_377),
.A2(n_346),
.B1(n_330),
.B2(n_341),
.Y(n_400)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_400),
.Y(n_412)
);

MAJIxp5_ASAP7_75t_L g401 ( 
.A(n_347),
.B(n_329),
.C(n_342),
.Y(n_401)
);

MAJIxp5_ASAP7_75t_L g418 ( 
.A(n_401),
.B(n_379),
.C(n_350),
.Y(n_418)
);

XOR2xp5_ASAP7_75t_L g402 ( 
.A(n_347),
.B(n_341),
.Y(n_402)
);

CKINVDCx20_ASAP7_75t_R g403 ( 
.A(n_364),
.Y(n_403)
);

XNOR2xp5_ASAP7_75t_L g429 ( 
.A(n_404),
.B(n_373),
.Y(n_429)
);

AOI22xp5_ASAP7_75t_L g407 ( 
.A1(n_355),
.A2(n_331),
.B1(n_325),
.B2(n_309),
.Y(n_407)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_407),
.Y(n_421)
);

OAI22xp5_ASAP7_75t_L g408 ( 
.A1(n_357),
.A2(n_325),
.B1(n_309),
.B2(n_337),
.Y(n_408)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_408),
.Y(n_424)
);

NOR2xp33_ASAP7_75t_L g409 ( 
.A(n_351),
.B(n_251),
.Y(n_409)
);

NOR2xp33_ASAP7_75t_SL g423 ( 
.A(n_409),
.B(n_356),
.Y(n_423)
);

AOI22xp5_ASAP7_75t_L g410 ( 
.A1(n_368),
.A2(n_337),
.B1(n_308),
.B2(n_281),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_410),
.B(n_349),
.Y(n_414)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_414),
.Y(n_442)
);

FAx1_ASAP7_75t_SL g416 ( 
.A(n_398),
.B(n_348),
.CI(n_350),
.CON(n_416),
.SN(n_416)
);

FAx1_ASAP7_75t_SL g450 ( 
.A(n_416),
.B(n_395),
.CI(n_370),
.CON(n_450),
.SN(n_450)
);

XOR2xp5_ASAP7_75t_L g438 ( 
.A(n_417),
.B(n_429),
.Y(n_438)
);

MAJIxp5_ASAP7_75t_L g445 ( 
.A(n_418),
.B(n_420),
.C(n_428),
.Y(n_445)
);

INVxp33_ASAP7_75t_L g419 ( 
.A(n_396),
.Y(n_419)
);

INVx1_ASAP7_75t_SL g443 ( 
.A(n_419),
.Y(n_443)
);

MAJIxp5_ASAP7_75t_L g420 ( 
.A(n_402),
.B(n_379),
.C(n_367),
.Y(n_420)
);

OAI22xp5_ASAP7_75t_SL g440 ( 
.A1(n_422),
.A2(n_362),
.B1(n_393),
.B2(n_407),
.Y(n_440)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_423),
.Y(n_448)
);

CKINVDCx20_ASAP7_75t_R g425 ( 
.A(n_392),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_SL g444 ( 
.A(n_425),
.B(n_426),
.Y(n_444)
);

CKINVDCx20_ASAP7_75t_R g426 ( 
.A(n_399),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_411),
.B(n_364),
.Y(n_427)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_427),
.Y(n_457)
);

MAJIxp5_ASAP7_75t_L g428 ( 
.A(n_388),
.B(n_360),
.C(n_349),
.Y(n_428)
);

XOR2xp5_ASAP7_75t_L g431 ( 
.A(n_398),
.B(n_365),
.Y(n_431)
);

XNOR2xp5_ASAP7_75t_SL g451 ( 
.A(n_431),
.B(n_406),
.Y(n_451)
);

MAJIxp5_ASAP7_75t_L g432 ( 
.A(n_401),
.B(n_369),
.C(n_365),
.Y(n_432)
);

MAJIxp5_ASAP7_75t_L g452 ( 
.A(n_432),
.B(n_437),
.C(n_387),
.Y(n_452)
);

CKINVDCx20_ASAP7_75t_R g433 ( 
.A(n_381),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_SL g447 ( 
.A(n_433),
.B(n_435),
.Y(n_447)
);

XNOR2xp5_ASAP7_75t_L g434 ( 
.A(n_404),
.B(n_370),
.Y(n_434)
);

XNOR2xp5_ASAP7_75t_L g449 ( 
.A(n_434),
.B(n_406),
.Y(n_449)
);

CKINVDCx20_ASAP7_75t_R g435 ( 
.A(n_411),
.Y(n_435)
);

MAJIxp5_ASAP7_75t_L g437 ( 
.A(n_386),
.B(n_384),
.C(n_389),
.Y(n_437)
);

AOI22xp5_ASAP7_75t_L g439 ( 
.A1(n_413),
.A2(n_397),
.B1(n_389),
.B2(n_385),
.Y(n_439)
);

OAI22xp5_ASAP7_75t_SL g460 ( 
.A1(n_439),
.A2(n_414),
.B1(n_412),
.B2(n_427),
.Y(n_460)
);

AOI22xp5_ASAP7_75t_SL g459 ( 
.A1(n_440),
.A2(n_442),
.B1(n_424),
.B2(n_457),
.Y(n_459)
);

OAI22xp5_ASAP7_75t_SL g441 ( 
.A1(n_422),
.A2(n_393),
.B1(n_410),
.B2(n_400),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_SL g472 ( 
.A(n_441),
.B(n_446),
.Y(n_472)
);

OAI22xp5_ASAP7_75t_SL g446 ( 
.A1(n_436),
.A2(n_412),
.B1(n_424),
.B2(n_421),
.Y(n_446)
);

XOR2xp5_ASAP7_75t_L g462 ( 
.A(n_449),
.B(n_429),
.Y(n_462)
);

NOR2xp33_ASAP7_75t_L g473 ( 
.A(n_450),
.B(n_454),
.Y(n_473)
);

XNOR2xp5_ASAP7_75t_SL g465 ( 
.A(n_451),
.B(n_434),
.Y(n_465)
);

XNOR2xp5_ASAP7_75t_L g463 ( 
.A(n_452),
.B(n_456),
.Y(n_463)
);

A2O1A1Ixp33_ASAP7_75t_SL g453 ( 
.A1(n_421),
.A2(n_387),
.B(n_385),
.C(n_366),
.Y(n_453)
);

HB1xp67_ASAP7_75t_L g475 ( 
.A(n_453),
.Y(n_475)
);

MAJIxp5_ASAP7_75t_L g454 ( 
.A(n_430),
.B(n_382),
.C(n_363),
.Y(n_454)
);

OAI21xp5_ASAP7_75t_SL g455 ( 
.A1(n_419),
.A2(n_372),
.B(n_382),
.Y(n_455)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_455),
.Y(n_461)
);

MAJIxp5_ASAP7_75t_L g456 ( 
.A(n_430),
.B(n_394),
.C(n_376),
.Y(n_456)
);

XNOR2xp5_ASAP7_75t_L g458 ( 
.A(n_431),
.B(n_405),
.Y(n_458)
);

XNOR2xp5_ASAP7_75t_L g471 ( 
.A(n_458),
.B(n_420),
.Y(n_471)
);

INVxp67_ASAP7_75t_L g479 ( 
.A(n_459),
.Y(n_479)
);

XOR2xp5_ASAP7_75t_L g477 ( 
.A(n_460),
.B(n_474),
.Y(n_477)
);

XNOR2xp5_ASAP7_75t_L g476 ( 
.A(n_462),
.B(n_464),
.Y(n_476)
);

XOR2xp5_ASAP7_75t_L g464 ( 
.A(n_458),
.B(n_437),
.Y(n_464)
);

XNOR2xp5_ASAP7_75t_L g482 ( 
.A(n_465),
.B(n_471),
.Y(n_482)
);

OAI22xp5_ASAP7_75t_SL g466 ( 
.A1(n_448),
.A2(n_432),
.B1(n_394),
.B2(n_428),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_L g490 ( 
.A(n_466),
.B(n_467),
.Y(n_490)
);

CKINVDCx20_ASAP7_75t_R g467 ( 
.A(n_444),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_447),
.Y(n_468)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_468),
.Y(n_487)
);

CKINVDCx20_ASAP7_75t_R g469 ( 
.A(n_454),
.Y(n_469)
);

NOR2xp33_ASAP7_75t_L g478 ( 
.A(n_469),
.B(n_470),
.Y(n_478)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_443),
.Y(n_470)
);

XOR2xp5_ASAP7_75t_L g474 ( 
.A(n_438),
.B(n_415),
.Y(n_474)
);

NOR2xp33_ASAP7_75t_L g480 ( 
.A(n_463),
.B(n_439),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_L g498 ( 
.A(n_480),
.B(n_481),
.Y(n_498)
);

NOR2xp33_ASAP7_75t_L g481 ( 
.A(n_463),
.B(n_443),
.Y(n_481)
);

MAJIxp5_ASAP7_75t_L g483 ( 
.A(n_471),
.B(n_445),
.C(n_452),
.Y(n_483)
);

AOI21xp5_ASAP7_75t_L g493 ( 
.A1(n_483),
.A2(n_485),
.B(n_486),
.Y(n_493)
);

OR2x2_ASAP7_75t_L g484 ( 
.A(n_461),
.B(n_450),
.Y(n_484)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_484),
.Y(n_500)
);

MAJIxp5_ASAP7_75t_L g485 ( 
.A(n_464),
.B(n_445),
.C(n_418),
.Y(n_485)
);

OAI21xp5_ASAP7_75t_SL g486 ( 
.A1(n_473),
.A2(n_459),
.B(n_472),
.Y(n_486)
);

MAJIxp5_ASAP7_75t_L g488 ( 
.A(n_474),
.B(n_456),
.C(n_415),
.Y(n_488)
);

AOI21xp5_ASAP7_75t_L g502 ( 
.A1(n_488),
.A2(n_489),
.B(n_485),
.Y(n_502)
);

MAJIxp5_ASAP7_75t_L g489 ( 
.A(n_462),
.B(n_438),
.C(n_451),
.Y(n_489)
);

AOI22xp5_ASAP7_75t_SL g491 ( 
.A1(n_479),
.A2(n_490),
.B1(n_489),
.B2(n_475),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_L g506 ( 
.A(n_491),
.B(n_492),
.Y(n_506)
);

XNOR2xp5_ASAP7_75t_L g492 ( 
.A(n_476),
.B(n_449),
.Y(n_492)
);

AOI22xp5_ASAP7_75t_SL g494 ( 
.A1(n_479),
.A2(n_460),
.B1(n_416),
.B2(n_450),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_L g507 ( 
.A(n_494),
.B(n_495),
.Y(n_507)
);

AOI22xp5_ASAP7_75t_L g495 ( 
.A1(n_487),
.A2(n_378),
.B1(n_374),
.B2(n_375),
.Y(n_495)
);

OAI21xp5_ASAP7_75t_L g496 ( 
.A1(n_484),
.A2(n_416),
.B(n_417),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_L g509 ( 
.A(n_496),
.B(n_497),
.Y(n_509)
);

INVx3_ASAP7_75t_L g497 ( 
.A(n_478),
.Y(n_497)
);

NOR2xp33_ASAP7_75t_L g499 ( 
.A(n_477),
.B(n_371),
.Y(n_499)
);

OAI21x1_ASAP7_75t_SL g508 ( 
.A1(n_499),
.A2(n_503),
.B(n_453),
.Y(n_508)
);

MAJIxp5_ASAP7_75t_L g501 ( 
.A(n_483),
.B(n_465),
.C(n_453),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_SL g511 ( 
.A(n_501),
.B(n_502),
.Y(n_511)
);

AOI21xp5_ASAP7_75t_L g503 ( 
.A1(n_482),
.A2(n_477),
.B(n_488),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_L g504 ( 
.A(n_497),
.B(n_500),
.Y(n_504)
);

AO21x1_ASAP7_75t_L g514 ( 
.A1(n_504),
.A2(n_508),
.B(n_453),
.Y(n_514)
);

NOR2xp33_ASAP7_75t_L g505 ( 
.A(n_498),
.B(n_308),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_505),
.B(n_510),
.Y(n_515)
);

NOR2xp33_ASAP7_75t_L g510 ( 
.A(n_493),
.B(n_247),
.Y(n_510)
);

NOR2xp33_ASAP7_75t_L g512 ( 
.A(n_511),
.B(n_501),
.Y(n_512)
);

OAI21xp5_ASAP7_75t_SL g517 ( 
.A1(n_512),
.A2(n_513),
.B(n_516),
.Y(n_517)
);

NOR2xp33_ASAP7_75t_L g513 ( 
.A(n_504),
.B(n_499),
.Y(n_513)
);

OAI22xp5_ASAP7_75t_L g518 ( 
.A1(n_514),
.A2(n_507),
.B1(n_506),
.B2(n_251),
.Y(n_518)
);

NOR2xp33_ASAP7_75t_L g516 ( 
.A(n_509),
.B(n_247),
.Y(n_516)
);

OAI321xp33_ASAP7_75t_L g520 ( 
.A1(n_518),
.A2(n_227),
.A3(n_245),
.B1(n_248),
.B2(n_231),
.C(n_246),
.Y(n_520)
);

INVxp67_ASAP7_75t_L g519 ( 
.A(n_515),
.Y(n_519)
);

OAI21xp5_ASAP7_75t_L g521 ( 
.A1(n_519),
.A2(n_231),
.B(n_238),
.Y(n_521)
);

AOI21xp5_ASAP7_75t_L g522 ( 
.A1(n_520),
.A2(n_521),
.B(n_517),
.Y(n_522)
);

BUFx24_ASAP7_75t_SL g523 ( 
.A(n_522),
.Y(n_523)
);

AOI21xp5_ASAP7_75t_L g524 ( 
.A1(n_523),
.A2(n_238),
.B(n_246),
.Y(n_524)
);

BUFx24_ASAP7_75t_SL g525 ( 
.A(n_524),
.Y(n_525)
);


endmodule