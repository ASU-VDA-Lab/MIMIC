module fake_jpeg_22501_n_180 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_180);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_180;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_175;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_118;
wire n_140;
wire n_82;
wire n_128;
wire n_100;
wire n_96;

INVx1_ASAP7_75t_L g15 ( 
.A(n_10),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

BUFx10_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_0),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_13),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_5),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_3),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_12),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_6),
.B(n_8),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_1),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_1),
.Y(n_30)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

CKINVDCx14_ASAP7_75t_R g32 ( 
.A(n_13),
.Y(n_32)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_25),
.Y(n_33)
);

BUFx2_ASAP7_75t_SL g48 ( 
.A(n_33),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_22),
.B(n_0),
.Y(n_34)
);

OR2x2_ASAP7_75t_L g55 ( 
.A(n_34),
.B(n_26),
.Y(n_55)
);

BUFx2_ASAP7_75t_L g35 ( 
.A(n_25),
.Y(n_35)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_35),
.Y(n_52)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_17),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_36),
.B(n_31),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_17),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_37),
.Y(n_60)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_17),
.Y(n_38)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_38),
.A2(n_28),
.B1(n_18),
.B2(n_15),
.Y(n_53)
);

BUFx5_ASAP7_75t_L g39 ( 
.A(n_19),
.Y(n_39)
);

BUFx12_ASAP7_75t_L g47 ( 
.A(n_39),
.Y(n_47)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_19),
.Y(n_40)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_40),
.Y(n_65)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_27),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g56 ( 
.A(n_41),
.B(n_43),
.Y(n_56)
);

INVx5_ASAP7_75t_L g42 ( 
.A(n_19),
.Y(n_42)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_42),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_22),
.B(n_0),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_20),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_44),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_20),
.Y(n_45)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_45),
.Y(n_62)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_46),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g49 ( 
.A1(n_38),
.A2(n_31),
.B1(n_24),
.B2(n_30),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_L g68 ( 
.A1(n_49),
.A2(n_21),
.B1(n_24),
.B2(n_40),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_34),
.B(n_23),
.Y(n_50)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_50),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_37),
.B(n_20),
.Y(n_51)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_51),
.B(n_64),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_53),
.B(n_55),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_42),
.A2(n_16),
.B1(n_15),
.B2(n_29),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_54),
.A2(n_58),
.B1(n_36),
.B2(n_28),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_41),
.B(n_23),
.Y(n_57)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_57),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_38),
.A2(n_16),
.B1(n_30),
.B2(n_29),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_45),
.Y(n_63)
);

INVx5_ASAP7_75t_SL g74 ( 
.A(n_63),
.Y(n_74)
);

NAND2x1_ASAP7_75t_L g64 ( 
.A(n_39),
.B(n_18),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_33),
.B(n_26),
.Y(n_66)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_66),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_68),
.A2(n_88),
.B1(n_61),
.B2(n_60),
.Y(n_108)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_47),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_69),
.B(n_71),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_52),
.B(n_21),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_70),
.B(n_76),
.Y(n_92)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_48),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_51),
.B(n_44),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_73),
.B(n_82),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_52),
.B(n_32),
.Y(n_76)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_47),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_77),
.B(n_78),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_49),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_80),
.A2(n_62),
.B1(n_61),
.B2(n_60),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_55),
.B(n_44),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_56),
.B(n_2),
.Y(n_83)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_83),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_56),
.B(n_2),
.Y(n_84)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_84),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_47),
.B(n_2),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_86),
.B(n_4),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_65),
.B(n_37),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_87),
.B(n_7),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_L g88 ( 
.A1(n_59),
.A2(n_18),
.B1(n_35),
.B2(n_3),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_65),
.B(n_18),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_89),
.Y(n_91)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_64),
.B(n_3),
.Y(n_90)
);

OAI21xp5_ASAP7_75t_SL g102 ( 
.A1(n_90),
.A2(n_4),
.B(n_59),
.Y(n_102)
);

BUFx24_ASAP7_75t_L g95 ( 
.A(n_74),
.Y(n_95)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_95),
.Y(n_112)
);

XNOR2xp5_ASAP7_75t_L g96 ( 
.A(n_75),
.B(n_64),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_96),
.B(n_109),
.Y(n_123)
);

NOR2xp67_ASAP7_75t_L g97 ( 
.A(n_75),
.B(n_7),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_97),
.B(n_103),
.Y(n_116)
);

HAxp5_ASAP7_75t_SL g99 ( 
.A(n_67),
.B(n_35),
.CON(n_99),
.SN(n_99)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_99),
.A2(n_72),
.B1(n_85),
.B2(n_69),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_102),
.A2(n_105),
.B1(n_68),
.B2(n_90),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_SL g103 ( 
.A(n_82),
.B(n_14),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_104),
.B(n_106),
.Y(n_114)
);

BUFx5_ASAP7_75t_L g106 ( 
.A(n_74),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_71),
.B(n_62),
.Y(n_107)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_107),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_108),
.A2(n_80),
.B1(n_87),
.B2(n_73),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_75),
.B(n_63),
.C(n_4),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_110),
.B(n_90),
.Y(n_126)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_101),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_111),
.B(n_113),
.Y(n_137)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_94),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_92),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_115),
.Y(n_136)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_95),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_117),
.B(n_118),
.Y(n_138)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_95),
.Y(n_118)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_95),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_119),
.B(n_124),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_120),
.A2(n_122),
.B1(n_127),
.B2(n_108),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_SL g121 ( 
.A(n_93),
.B(n_79),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_SL g140 ( 
.A(n_121),
.B(n_125),
.Y(n_140)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_106),
.Y(n_124)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_110),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_126),
.B(n_98),
.Y(n_142)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_114),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_129),
.B(n_135),
.Y(n_151)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_120),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_130),
.B(n_103),
.Y(n_145)
);

OA21x2_ASAP7_75t_SL g132 ( 
.A1(n_126),
.A2(n_96),
.B(n_99),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_L g144 ( 
.A1(n_132),
.A2(n_141),
.B(n_142),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_123),
.B(n_98),
.C(n_109),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_133),
.B(n_111),
.C(n_91),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_134),
.B(n_112),
.Y(n_150)
);

INVxp67_ASAP7_75t_L g135 ( 
.A(n_127),
.Y(n_135)
);

INVx2_ASAP7_75t_SL g139 ( 
.A(n_117),
.Y(n_139)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_139),
.Y(n_146)
);

OAI21x1_ASAP7_75t_SL g141 ( 
.A1(n_123),
.A2(n_105),
.B(n_102),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_143),
.B(n_130),
.C(n_134),
.Y(n_155)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_145),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_L g147 ( 
.A(n_133),
.B(n_91),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_L g159 ( 
.A(n_147),
.B(n_129),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_L g148 ( 
.A1(n_135),
.A2(n_142),
.B(n_141),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_148),
.B(n_152),
.Y(n_156)
);

OAI21xp33_ASAP7_75t_L g149 ( 
.A1(n_138),
.A2(n_113),
.B(n_119),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_SL g157 ( 
.A1(n_149),
.A2(n_153),
.B(n_118),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_150),
.A2(n_139),
.B1(n_128),
.B2(n_85),
.Y(n_161)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_137),
.Y(n_152)
);

AND2x4_ASAP7_75t_SL g153 ( 
.A(n_139),
.B(n_112),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_146),
.B(n_131),
.Y(n_154)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_154),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_155),
.B(n_157),
.C(n_151),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_SL g166 ( 
.A(n_159),
.B(n_161),
.Y(n_166)
);

AOI321xp33_ASAP7_75t_L g160 ( 
.A1(n_144),
.A2(n_140),
.A3(n_136),
.B1(n_116),
.B2(n_100),
.C(n_93),
.Y(n_160)
);

AOI21xp33_ASAP7_75t_L g163 ( 
.A1(n_160),
.A2(n_100),
.B(n_79),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_L g171 ( 
.A1(n_162),
.A2(n_163),
.B(n_72),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_155),
.B(n_143),
.C(n_153),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_L g170 ( 
.A(n_165),
.B(n_159),
.Y(n_170)
);

NOR3xp33_ASAP7_75t_L g167 ( 
.A(n_158),
.B(n_153),
.C(n_149),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_167),
.B(n_156),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_168),
.A2(n_81),
.B1(n_11),
.B2(n_14),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_164),
.B(n_147),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_169),
.B(n_81),
.C(n_10),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_170),
.B(n_171),
.C(n_172),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_L g172 ( 
.A(n_166),
.B(n_77),
.Y(n_172)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_173),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_175),
.B(n_168),
.Y(n_176)
);

INVxp67_ASAP7_75t_L g178 ( 
.A(n_176),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_178),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_179),
.B(n_174),
.C(n_177),
.Y(n_180)
);


endmodule