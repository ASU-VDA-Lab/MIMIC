module fake_jpeg_6384_n_337 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_337);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_337;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx4_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_12),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_16),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_10),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_9),
.Y(n_24)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_15),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_16),
.Y(n_27)
);

INVx5_ASAP7_75t_L g28 ( 
.A(n_16),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_0),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_12),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_4),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_15),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_6),
.Y(n_34)
);

INVx11_ASAP7_75t_SL g35 ( 
.A(n_15),
.Y(n_35)
);

BUFx10_ASAP7_75t_L g36 ( 
.A(n_28),
.Y(n_36)
);

CKINVDCx16_ASAP7_75t_R g48 ( 
.A(n_36),
.Y(n_48)
);

INVx5_ASAP7_75t_L g37 ( 
.A(n_28),
.Y(n_37)
);

BUFx2_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_30),
.B(n_0),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_SL g54 ( 
.A(n_38),
.B(n_39),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_30),
.B(n_0),
.Y(n_39)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_26),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_40),
.A2(n_17),
.B1(n_25),
.B2(n_41),
.Y(n_67)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_26),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_41),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_28),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_42),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_20),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_43),
.B(n_44),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_27),
.B(n_7),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_26),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_45),
.B(n_46),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_20),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

BUFx10_ASAP7_75t_L g63 ( 
.A(n_47),
.Y(n_63)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_38),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_49),
.B(n_55),
.Y(n_89)
);

AOI21xp33_ASAP7_75t_L g50 ( 
.A1(n_38),
.A2(n_18),
.B(n_34),
.Y(n_50)
);

AOI21xp33_ASAP7_75t_SL g96 ( 
.A1(n_50),
.A2(n_36),
.B(n_18),
.Y(n_96)
);

OAI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_37),
.A2(n_27),
.B1(n_21),
.B2(n_33),
.Y(n_52)
);

OAI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_52),
.A2(n_46),
.B1(n_43),
.B2(n_21),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_L g53 ( 
.A1(n_37),
.A2(n_27),
.B1(n_17),
.B2(n_25),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_53),
.A2(n_56),
.B1(n_19),
.B2(n_22),
.Y(n_85)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_37),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_L g56 ( 
.A1(n_43),
.A2(n_25),
.B1(n_17),
.B2(n_33),
.Y(n_56)
);

INVx2_ASAP7_75t_SL g58 ( 
.A(n_47),
.Y(n_58)
);

INVx11_ASAP7_75t_L g72 ( 
.A(n_58),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g60 ( 
.A1(n_41),
.A2(n_29),
.B1(n_34),
.B2(n_32),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_60),
.A2(n_24),
.B1(n_20),
.B2(n_21),
.Y(n_88)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_47),
.Y(n_61)
);

INVx6_ASAP7_75t_L g92 ( 
.A(n_61),
.Y(n_92)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_47),
.Y(n_62)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_62),
.Y(n_71)
);

MAJIxp5_ASAP7_75t_L g64 ( 
.A(n_45),
.B(n_30),
.C(n_19),
.Y(n_64)
);

MAJIxp5_ASAP7_75t_L g74 ( 
.A(n_64),
.B(n_66),
.C(n_44),
.Y(n_74)
);

AND2x2_ASAP7_75t_SL g66 ( 
.A(n_36),
.B(n_39),
.Y(n_66)
);

CKINVDCx16_ASAP7_75t_R g87 ( 
.A(n_67),
.Y(n_87)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_39),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_68),
.B(n_22),
.Y(n_93)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_47),
.Y(n_70)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_70),
.Y(n_84)
);

NAND2x1_ASAP7_75t_SL g73 ( 
.A(n_66),
.B(n_35),
.Y(n_73)
);

NAND2xp33_ASAP7_75t_SL g110 ( 
.A(n_73),
.B(n_96),
.Y(n_110)
);

XNOR2xp5_ASAP7_75t_L g123 ( 
.A(n_74),
.B(n_83),
.Y(n_123)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_51),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_75),
.B(n_79),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_L g107 ( 
.A1(n_76),
.A2(n_85),
.B1(n_31),
.B2(n_33),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_L g77 ( 
.A1(n_66),
.A2(n_25),
.B1(n_17),
.B2(n_40),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_77),
.A2(n_80),
.B1(n_88),
.B2(n_81),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_69),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_78),
.B(n_81),
.Y(n_106)
);

BUFx12f_ASAP7_75t_L g79 ( 
.A(n_66),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_L g80 ( 
.A1(n_49),
.A2(n_40),
.B1(n_41),
.B2(n_46),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_69),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_68),
.B(n_45),
.C(n_44),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_82),
.B(n_59),
.C(n_74),
.Y(n_115)
);

XNOR2xp5_ASAP7_75t_L g83 ( 
.A(n_50),
.B(n_36),
.Y(n_83)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_60),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_86),
.B(n_90),
.Y(n_109)
);

INVx6_ASAP7_75t_SL g90 ( 
.A(n_58),
.Y(n_90)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_51),
.Y(n_91)
);

BUFx2_ASAP7_75t_L g113 ( 
.A(n_91),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_93),
.B(n_95),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_48),
.A2(n_40),
.B1(n_31),
.B2(n_23),
.Y(n_94)
);

INVxp67_ASAP7_75t_L g102 ( 
.A(n_94),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_63),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_54),
.B(n_36),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_97),
.B(n_100),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_54),
.A2(n_40),
.B1(n_36),
.B2(n_42),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_98),
.A2(n_87),
.B1(n_94),
.B2(n_73),
.Y(n_114)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_70),
.Y(n_99)
);

INVxp33_ASAP7_75t_L g101 ( 
.A(n_99),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_63),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_87),
.A2(n_55),
.B1(n_48),
.B2(n_62),
.Y(n_104)
);

INVxp67_ASAP7_75t_L g153 ( 
.A(n_104),
.Y(n_153)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_88),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_105),
.B(n_111),
.Y(n_154)
);

AOI22xp33_ASAP7_75t_L g131 ( 
.A1(n_107),
.A2(n_24),
.B1(n_23),
.B2(n_19),
.Y(n_131)
);

OA21x2_ASAP7_75t_L g108 ( 
.A1(n_96),
.A2(n_36),
.B(n_53),
.Y(n_108)
);

HAxp5_ASAP7_75t_SL g133 ( 
.A(n_108),
.B(n_122),
.CON(n_133),
.SN(n_133)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_93),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_86),
.A2(n_59),
.B1(n_61),
.B2(n_62),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_112),
.A2(n_118),
.B1(n_126),
.B2(n_72),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_114),
.A2(n_128),
.B1(n_91),
.B2(n_75),
.Y(n_141)
);

AND2x2_ASAP7_75t_L g147 ( 
.A(n_115),
.B(n_29),
.Y(n_147)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_90),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_116),
.B(n_117),
.Y(n_156)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_89),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_L g118 ( 
.A1(n_73),
.A2(n_70),
.B1(n_31),
.B2(n_24),
.Y(n_118)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_98),
.Y(n_120)
);

CKINVDCx14_ASAP7_75t_R g149 ( 
.A(n_120),
.Y(n_149)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_97),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_121),
.B(n_71),
.Y(n_157)
);

OA21x2_ASAP7_75t_L g122 ( 
.A1(n_85),
.A2(n_36),
.B(n_42),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_79),
.B(n_64),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_124),
.B(n_127),
.Y(n_134)
);

INVxp67_ASAP7_75t_L g125 ( 
.A(n_99),
.Y(n_125)
);

CKINVDCx16_ASAP7_75t_R g148 ( 
.A(n_125),
.Y(n_148)
);

OA22x2_ASAP7_75t_L g126 ( 
.A1(n_83),
.A2(n_42),
.B1(n_65),
.B2(n_51),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_79),
.B(n_32),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_126),
.A2(n_79),
.B1(n_78),
.B2(n_82),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_130),
.A2(n_160),
.B1(n_102),
.B2(n_128),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_131),
.A2(n_141),
.B1(n_155),
.B2(n_158),
.Y(n_172)
);

BUFx2_ASAP7_75t_L g132 ( 
.A(n_113),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_132),
.B(n_138),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_123),
.B(n_100),
.C(n_95),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_135),
.B(n_147),
.C(n_150),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_SL g136 ( 
.A(n_106),
.B(n_23),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_136),
.B(n_143),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_113),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_137),
.Y(n_166)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_106),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_121),
.B(n_119),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_139),
.B(n_151),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_L g140 ( 
.A(n_123),
.B(n_42),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_L g190 ( 
.A(n_140),
.B(n_57),
.Y(n_190)
);

OAI21xp5_ASAP7_75t_SL g142 ( 
.A1(n_126),
.A2(n_71),
.B(n_84),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_SL g191 ( 
.A1(n_142),
.A2(n_146),
.B(n_7),
.Y(n_191)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_103),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_103),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_144),
.B(n_145),
.Y(n_185)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_112),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_L g146 ( 
.A1(n_127),
.A2(n_29),
.B(n_32),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_115),
.B(n_124),
.C(n_129),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_119),
.B(n_84),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_109),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_152),
.B(n_111),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_L g155 ( 
.A1(n_126),
.A2(n_105),
.B1(n_122),
.B2(n_117),
.Y(n_155)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_157),
.Y(n_168)
);

AOI22xp33_ASAP7_75t_L g158 ( 
.A1(n_126),
.A2(n_92),
.B1(n_22),
.B2(n_34),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_114),
.A2(n_58),
.B1(n_92),
.B2(n_72),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_159),
.A2(n_142),
.B1(n_141),
.B2(n_145),
.Y(n_171)
);

CKINVDCx14_ASAP7_75t_R g162 ( 
.A(n_156),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_162),
.B(n_178),
.Y(n_198)
);

AO22x1_ASAP7_75t_SL g163 ( 
.A1(n_133),
.A2(n_122),
.B1(n_108),
.B2(n_110),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_163),
.A2(n_187),
.B1(n_189),
.B2(n_132),
.Y(n_213)
);

BUFx5_ASAP7_75t_L g165 ( 
.A(n_132),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_165),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_L g205 ( 
.A1(n_167),
.A2(n_184),
.B1(n_152),
.B2(n_136),
.Y(n_205)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_169),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_SL g170 ( 
.A(n_130),
.B(n_110),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_170),
.B(n_8),
.C(n_14),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_171),
.A2(n_173),
.B1(n_179),
.B2(n_194),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_L g173 ( 
.A1(n_149),
.A2(n_109),
.B1(n_122),
.B2(n_108),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_SL g174 ( 
.A(n_154),
.B(n_108),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_174),
.B(n_176),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_139),
.B(n_151),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_134),
.B(n_113),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_177),
.B(n_188),
.Y(n_214)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_157),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_149),
.A2(n_159),
.B1(n_138),
.B2(n_154),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_156),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_180),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_153),
.A2(n_116),
.B1(n_18),
.B2(n_26),
.Y(n_181)
);

INVxp67_ASAP7_75t_L g217 ( 
.A(n_181),
.Y(n_217)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_134),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_182),
.B(n_192),
.Y(n_216)
);

AOI22xp33_ASAP7_75t_L g184 ( 
.A1(n_146),
.A2(n_65),
.B1(n_101),
.B2(n_63),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_137),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_186),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_160),
.A2(n_65),
.B1(n_57),
.B2(n_63),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_143),
.B(n_63),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_135),
.A2(n_57),
.B1(n_18),
.B2(n_2),
.Y(n_189)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_190),
.B(n_1),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_SL g206 ( 
.A1(n_191),
.A2(n_147),
.B(n_148),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_SL g192 ( 
.A(n_144),
.B(n_7),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_147),
.Y(n_193)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_193),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_150),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_194)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_161),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_197),
.B(n_199),
.Y(n_248)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_161),
.Y(n_199)
);

INVx1_ASAP7_75t_SL g200 ( 
.A(n_165),
.Y(n_200)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_200),
.Y(n_231)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_176),
.Y(n_201)
);

AOI21xp5_ASAP7_75t_L g235 ( 
.A1(n_201),
.A2(n_206),
.B(n_211),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_205),
.A2(n_213),
.B1(n_221),
.B2(n_172),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_163),
.A2(n_140),
.B1(n_148),
.B2(n_9),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_207),
.A2(n_192),
.B1(n_178),
.B2(n_168),
.Y(n_237)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_208),
.B(n_209),
.Y(n_226)
);

INVx1_ASAP7_75t_SL g210 ( 
.A(n_174),
.Y(n_210)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_210),
.Y(n_236)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_177),
.Y(n_211)
);

AND2x2_ASAP7_75t_L g215 ( 
.A(n_163),
.B(n_1),
.Y(n_215)
);

OAI21xp5_ASAP7_75t_L g249 ( 
.A1(n_215),
.A2(n_3),
.B(n_4),
.Y(n_249)
);

XOR2xp5_ASAP7_75t_L g219 ( 
.A(n_164),
.B(n_14),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_219),
.B(n_220),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_164),
.B(n_2),
.C(n_3),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_L g221 ( 
.A1(n_167),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_221)
);

INVxp67_ASAP7_75t_L g222 ( 
.A(n_175),
.Y(n_222)
);

AOI21xp5_ASAP7_75t_L g243 ( 
.A1(n_222),
.A2(n_186),
.B(n_166),
.Y(n_243)
);

OAI21xp33_ASAP7_75t_L g223 ( 
.A1(n_185),
.A2(n_8),
.B(n_11),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_SL g241 ( 
.A(n_223),
.B(n_11),
.Y(n_241)
);

FAx1_ASAP7_75t_SL g224 ( 
.A(n_202),
.B(n_170),
.CI(n_189),
.CON(n_224),
.SN(n_224)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_224),
.B(n_225),
.Y(n_252)
);

INVxp67_ASAP7_75t_L g225 ( 
.A(n_198),
.Y(n_225)
);

CKINVDCx16_ASAP7_75t_R g227 ( 
.A(n_214),
.Y(n_227)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_227),
.Y(n_250)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_228),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_213),
.A2(n_171),
.B1(n_182),
.B2(n_193),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_229),
.A2(n_233),
.B1(n_228),
.B2(n_234),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_208),
.B(n_190),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_230),
.B(n_240),
.Y(n_253)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_200),
.Y(n_232)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_232),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_215),
.A2(n_194),
.B1(n_191),
.B2(n_187),
.Y(n_233)
);

XOR2x2_ASAP7_75t_L g234 ( 
.A(n_210),
.B(n_169),
.Y(n_234)
);

OAI21xp5_ASAP7_75t_L g263 ( 
.A1(n_234),
.A2(n_249),
.B(n_203),
.Y(n_263)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_237),
.Y(n_266)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_214),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_238),
.B(n_242),
.Y(n_256)
);

OAI21xp5_ASAP7_75t_SL g239 ( 
.A1(n_206),
.A2(n_183),
.B(n_180),
.Y(n_239)
);

OAI21xp5_ASAP7_75t_SL g259 ( 
.A1(n_239),
.A2(n_243),
.B(n_235),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_202),
.B(n_188),
.Y(n_240)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_241),
.Y(n_268)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_216),
.Y(n_242)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_212),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_244),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_219),
.B(n_168),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_246),
.B(n_209),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_L g247 ( 
.A1(n_212),
.A2(n_166),
.B1(n_181),
.B2(n_5),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_247),
.A2(n_249),
.B1(n_241),
.B2(n_195),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_251),
.A2(n_258),
.B1(n_224),
.B2(n_220),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_245),
.B(n_211),
.C(n_207),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_255),
.B(n_226),
.C(n_245),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_229),
.A2(n_233),
.B1(n_236),
.B2(n_201),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_259),
.Y(n_273)
);

HB1xp67_ASAP7_75t_L g260 ( 
.A(n_231),
.Y(n_260)
);

CKINVDCx16_ASAP7_75t_R g277 ( 
.A(n_260),
.Y(n_277)
);

OAI21xp5_ASAP7_75t_SL g262 ( 
.A1(n_248),
.A2(n_195),
.B(n_204),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_262),
.A2(n_265),
.B1(n_222),
.B2(n_217),
.Y(n_274)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_263),
.Y(n_284)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_264),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_225),
.A2(n_215),
.B1(n_199),
.B2(n_197),
.Y(n_265)
);

BUFx3_ASAP7_75t_L g267 ( 
.A(n_246),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_267),
.B(n_253),
.Y(n_276)
);

OAI21xp5_ASAP7_75t_SL g269 ( 
.A1(n_224),
.A2(n_217),
.B(n_218),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_SL g286 ( 
.A1(n_269),
.A2(n_10),
.B1(n_11),
.B2(n_13),
.Y(n_286)
);

XOR2xp5_ASAP7_75t_L g275 ( 
.A(n_270),
.B(n_230),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_271),
.B(n_275),
.C(n_281),
.Y(n_293)
);

BUFx2_ASAP7_75t_L g272 ( 
.A(n_261),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g292 ( 
.A(n_272),
.Y(n_292)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_274),
.Y(n_290)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_276),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_254),
.B(n_196),
.Y(n_278)
);

CKINVDCx16_ASAP7_75t_R g289 ( 
.A(n_278),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_258),
.B(n_240),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_279),
.B(n_282),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_280),
.B(n_283),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_255),
.B(n_226),
.C(n_4),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_SL g282 ( 
.A(n_263),
.B(n_9),
.Y(n_282)
);

BUFx24_ASAP7_75t_SL g283 ( 
.A(n_253),
.Y(n_283)
);

CKINVDCx16_ASAP7_75t_R g285 ( 
.A(n_262),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_285),
.B(n_284),
.Y(n_299)
);

AND2x2_ASAP7_75t_L g294 ( 
.A(n_286),
.B(n_252),
.Y(n_294)
);

NAND4xp25_ASAP7_75t_SL g288 ( 
.A(n_272),
.B(n_250),
.C(n_256),
.D(n_257),
.Y(n_288)
);

HB1xp67_ASAP7_75t_L g307 ( 
.A(n_288),
.Y(n_307)
);

OAI321xp33_ASAP7_75t_L g303 ( 
.A1(n_294),
.A2(n_284),
.A3(n_269),
.B1(n_287),
.B2(n_280),
.C(n_273),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_277),
.B(n_265),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_296),
.B(n_301),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_275),
.B(n_259),
.C(n_252),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_298),
.B(n_297),
.C(n_300),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_L g313 ( 
.A(n_299),
.B(n_5),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_L g300 ( 
.A1(n_287),
.A2(n_251),
.B1(n_266),
.B2(n_256),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_SL g311 ( 
.A1(n_300),
.A2(n_6),
.B1(n_3),
.B2(n_5),
.Y(n_311)
);

INVxp33_ASAP7_75t_L g301 ( 
.A(n_274),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_286),
.B(n_264),
.Y(n_302)
);

OAI21xp5_ASAP7_75t_SL g310 ( 
.A1(n_302),
.A2(n_270),
.B(n_10),
.Y(n_310)
);

AOI21xp5_ASAP7_75t_L g317 ( 
.A1(n_303),
.A2(n_308),
.B(n_310),
.Y(n_317)
);

XOR2xp5_ASAP7_75t_L g304 ( 
.A(n_298),
.B(n_271),
.Y(n_304)
);

XOR2xp5_ASAP7_75t_L g321 ( 
.A(n_304),
.B(n_305),
.Y(n_321)
);

XNOR2x1_ASAP7_75t_L g305 ( 
.A(n_301),
.B(n_273),
.Y(n_305)
);

XOR2xp5_ASAP7_75t_L g306 ( 
.A(n_293),
.B(n_281),
.Y(n_306)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_306),
.Y(n_322)
);

OAI21xp5_ASAP7_75t_L g308 ( 
.A1(n_293),
.A2(n_267),
.B(n_268),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_L g320 ( 
.A1(n_311),
.A2(n_291),
.B1(n_292),
.B2(n_6),
.Y(n_320)
);

OAI21xp5_ASAP7_75t_SL g312 ( 
.A1(n_290),
.A2(n_5),
.B(n_6),
.Y(n_312)
);

OAI21xp5_ASAP7_75t_L g318 ( 
.A1(n_312),
.A2(n_314),
.B(n_288),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_313),
.B(n_294),
.Y(n_319)
);

FAx1_ASAP7_75t_SL g315 ( 
.A(n_305),
.B(n_294),
.CI(n_302),
.CON(n_315),
.SN(n_315)
);

NAND2xp5_ASAP7_75t_SL g327 ( 
.A(n_315),
.B(n_319),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_307),
.B(n_289),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g324 ( 
.A(n_316),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_318),
.B(n_320),
.C(n_323),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_314),
.B(n_295),
.Y(n_323)
);

XOR2xp5_ASAP7_75t_L g326 ( 
.A(n_321),
.B(n_304),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_326),
.B(n_328),
.Y(n_332)
);

HB1xp67_ASAP7_75t_L g328 ( 
.A(n_315),
.Y(n_328)
);

INVxp33_ASAP7_75t_L g329 ( 
.A(n_317),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_329),
.B(n_321),
.Y(n_330)
);

A2O1A1O1Ixp25_ASAP7_75t_L g333 ( 
.A1(n_330),
.A2(n_331),
.B(n_309),
.C(n_318),
.D(n_325),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_324),
.B(n_320),
.Y(n_331)
);

AO221x1_ASAP7_75t_L g334 ( 
.A1(n_333),
.A2(n_329),
.B1(n_332),
.B2(n_306),
.C(n_327),
.Y(n_334)
);

BUFx24_ASAP7_75t_SL g335 ( 
.A(n_334),
.Y(n_335)
);

XNOR2xp5_ASAP7_75t_L g336 ( 
.A(n_335),
.B(n_322),
.Y(n_336)
);

BUFx24_ASAP7_75t_SL g337 ( 
.A(n_336),
.Y(n_337)
);


endmodule