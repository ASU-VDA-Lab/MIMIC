module fake_jpeg_27879_n_153 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_153);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_153;

wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_73;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_150;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_93;
wire n_91;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_135;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_96;

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_34),
.Y(n_39)
);

BUFx16f_ASAP7_75t_L g40 ( 
.A(n_20),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_28),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_4),
.Y(n_42)
);

BUFx5_ASAP7_75t_L g43 ( 
.A(n_17),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_36),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_30),
.Y(n_45)
);

BUFx12_ASAP7_75t_L g46 ( 
.A(n_33),
.Y(n_46)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_6),
.Y(n_47)
);

BUFx5_ASAP7_75t_L g48 ( 
.A(n_6),
.Y(n_48)
);

BUFx5_ASAP7_75t_L g49 ( 
.A(n_2),
.Y(n_49)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_24),
.Y(n_50)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_22),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_26),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_1),
.Y(n_53)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_2),
.Y(n_54)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_29),
.Y(n_55)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_32),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_4),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_21),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_11),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_27),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_38),
.Y(n_61)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_0),
.Y(n_62)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_51),
.Y(n_63)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_63),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_39),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_64),
.B(n_66),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_56),
.Y(n_65)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_65),
.Y(n_70)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_42),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_47),
.B(n_0),
.Y(n_67)
);

AND2x2_ASAP7_75t_L g73 ( 
.A(n_67),
.B(n_47),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_56),
.Y(n_68)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_68),
.Y(n_76)
);

INVx8_ASAP7_75t_L g69 ( 
.A(n_46),
.Y(n_69)
);

INVx5_ASAP7_75t_L g82 ( 
.A(n_69),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_65),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_SL g88 ( 
.A(n_71),
.B(n_39),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_68),
.B(n_57),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_72),
.B(n_73),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_63),
.Y(n_74)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_74),
.Y(n_96)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_69),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_75),
.B(n_78),
.Y(n_91)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_69),
.Y(n_78)
);

INVx2_ASAP7_75t_SL g80 ( 
.A(n_65),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_80),
.B(n_51),
.Y(n_93)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_63),
.Y(n_81)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_81),
.Y(n_92)
);

INVx13_ASAP7_75t_L g83 ( 
.A(n_82),
.Y(n_83)
);

INVx5_ASAP7_75t_L g104 ( 
.A(n_83),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_73),
.B(n_53),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_85),
.B(n_86),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_79),
.B(n_60),
.Y(n_86)
);

AND2x6_ASAP7_75t_L g87 ( 
.A(n_79),
.B(n_31),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_87),
.B(n_89),
.Y(n_102)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_88),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_70),
.B(n_60),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_76),
.A2(n_50),
.B1(n_55),
.B2(n_62),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_90),
.A2(n_54),
.B1(n_45),
.B2(n_58),
.Y(n_99)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_93),
.Y(n_105)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_80),
.Y(n_94)
);

INVx13_ASAP7_75t_L g100 ( 
.A(n_94),
.Y(n_100)
);

CKINVDCx16_ASAP7_75t_R g95 ( 
.A(n_77),
.Y(n_95)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_95),
.Y(n_103)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_74),
.Y(n_97)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_97),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_99),
.A2(n_97),
.B1(n_96),
.B2(n_91),
.Y(n_109)
);

INVx8_ASAP7_75t_L g106 ( 
.A(n_96),
.Y(n_106)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_106),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_109),
.B(n_98),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_102),
.B(n_92),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_110),
.B(n_111),
.Y(n_122)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_106),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_L g112 ( 
.A1(n_105),
.A2(n_84),
.B(n_103),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_L g126 ( 
.A1(n_112),
.A2(n_49),
.B(n_48),
.Y(n_126)
);

INVxp67_ASAP7_75t_L g113 ( 
.A(n_104),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_113),
.B(n_114),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_107),
.B(n_52),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_101),
.B(n_83),
.Y(n_115)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_115),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_100),
.A2(n_87),
.B1(n_61),
.B2(n_59),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_116),
.A2(n_117),
.B1(n_43),
.B2(n_3),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_100),
.A2(n_41),
.B1(n_44),
.B2(n_46),
.Y(n_117)
);

XNOR2xp5_ASAP7_75t_L g119 ( 
.A(n_112),
.B(n_103),
.Y(n_119)
);

XNOR2xp5_ASAP7_75t_SL g136 ( 
.A(n_119),
.B(n_124),
.Y(n_136)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_108),
.Y(n_121)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_121),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_123),
.A2(n_9),
.B1(n_10),
.B2(n_12),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_L g124 ( 
.A(n_113),
.B(n_40),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_114),
.B(n_104),
.Y(n_125)
);

CKINVDCx16_ASAP7_75t_R g137 ( 
.A(n_125),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_SL g133 ( 
.A(n_126),
.B(n_129),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_127),
.A2(n_5),
.B1(n_7),
.B2(n_8),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_L g128 ( 
.A(n_112),
.B(n_19),
.Y(n_128)
);

AOI21xp5_ASAP7_75t_L g138 ( 
.A1(n_128),
.A2(n_130),
.B(n_131),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_114),
.B(n_23),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_SL g130 ( 
.A1(n_110),
.A2(n_18),
.B(n_37),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_115),
.B(n_1),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_112),
.B(n_25),
.C(n_35),
.Y(n_132)
);

OA22x2_ASAP7_75t_L g134 ( 
.A1(n_132),
.A2(n_3),
.B1(n_5),
.B2(n_7),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_134),
.B(n_139),
.Y(n_142)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_140),
.Y(n_143)
);

INVx1_ASAP7_75t_SL g141 ( 
.A(n_133),
.Y(n_141)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_141),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_L g145 ( 
.A(n_144),
.B(n_136),
.Y(n_145)
);

OAI21x1_ASAP7_75t_L g146 ( 
.A1(n_145),
.A2(n_133),
.B(n_138),
.Y(n_146)
);

AND2x2_ASAP7_75t_L g147 ( 
.A(n_146),
.B(n_142),
.Y(n_147)
);

FAx1_ASAP7_75t_SL g148 ( 
.A(n_147),
.B(n_131),
.CI(n_122),
.CON(n_148),
.SN(n_148)
);

XOR2xp5_ASAP7_75t_L g149 ( 
.A(n_148),
.B(n_118),
.Y(n_149)
);

AOI21xp5_ASAP7_75t_L g150 ( 
.A1(n_149),
.A2(n_137),
.B(n_120),
.Y(n_150)
);

AO221x1_ASAP7_75t_L g151 ( 
.A1(n_150),
.A2(n_118),
.B1(n_134),
.B2(n_135),
.C(n_143),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_151),
.A2(n_13),
.B1(n_14),
.B2(n_15),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_152),
.B(n_16),
.Y(n_153)
);


endmodule