module fake_jpeg_19281_n_168 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_168);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_168;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_121;
wire n_99;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_40),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_46),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_9),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_39),
.B(n_15),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_12),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_34),
.Y(n_55)
);

BUFx12f_ASAP7_75t_L g56 ( 
.A(n_21),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_28),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_17),
.Y(n_58)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_16),
.Y(n_59)
);

BUFx4f_ASAP7_75t_L g60 ( 
.A(n_10),
.Y(n_60)
);

INVx11_ASAP7_75t_L g61 ( 
.A(n_48),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_37),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_31),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_19),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_3),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_4),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_1),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_11),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_11),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_13),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_29),
.Y(n_71)
);

BUFx2_ASAP7_75t_L g72 ( 
.A(n_4),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_32),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_3),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_33),
.Y(n_75)
);

BUFx5_ASAP7_75t_L g76 ( 
.A(n_23),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_47),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_2),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_51),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_79),
.Y(n_90)
);

INVx8_ASAP7_75t_L g80 ( 
.A(n_56),
.Y(n_80)
);

INVx6_ASAP7_75t_L g93 ( 
.A(n_80),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_60),
.B(n_24),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_81),
.B(n_69),
.Y(n_88)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_56),
.Y(n_82)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_82),
.Y(n_94)
);

BUFx3_ASAP7_75t_L g83 ( 
.A(n_60),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_83),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_51),
.Y(n_84)
);

BUFx2_ASAP7_75t_L g89 ( 
.A(n_84),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_59),
.A2(n_25),
.B1(n_45),
.B2(n_44),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_85),
.A2(n_53),
.B1(n_66),
.B2(n_74),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_58),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_86),
.B(n_77),
.Y(n_92)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_82),
.Y(n_87)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_87),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_88),
.B(n_81),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_92),
.B(n_54),
.Y(n_102)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_80),
.Y(n_95)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_95),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_85),
.A2(n_59),
.B1(n_61),
.B2(n_50),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_96),
.A2(n_97),
.B1(n_67),
.B2(n_78),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_98),
.B(n_105),
.Y(n_111)
);

BUFx12f_ASAP7_75t_L g100 ( 
.A(n_94),
.Y(n_100)
);

BUFx3_ASAP7_75t_L g123 ( 
.A(n_100),
.Y(n_123)
);

INVx1_ASAP7_75t_SL g101 ( 
.A(n_94),
.Y(n_101)
);

CKINVDCx16_ASAP7_75t_R g113 ( 
.A(n_101),
.Y(n_113)
);

CKINVDCx14_ASAP7_75t_R g116 ( 
.A(n_102),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_93),
.A2(n_84),
.B1(n_79),
.B2(n_75),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_104),
.A2(n_90),
.B1(n_83),
.B2(n_91),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_96),
.A2(n_62),
.B1(n_73),
.B2(n_64),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_106),
.B(n_108),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_90),
.Y(n_107)
);

INVx2_ASAP7_75t_SL g125 ( 
.A(n_107),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_89),
.B(n_68),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_93),
.A2(n_70),
.B1(n_55),
.B2(n_52),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_109),
.B(n_69),
.Y(n_119)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_89),
.Y(n_110)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_110),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_100),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_112),
.B(n_120),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_115),
.A2(n_71),
.B1(n_63),
.B2(n_57),
.Y(n_129)
);

CKINVDCx16_ASAP7_75t_R g118 ( 
.A(n_104),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_118),
.B(n_119),
.Y(n_127)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_100),
.Y(n_120)
);

AOI21xp5_ASAP7_75t_L g121 ( 
.A1(n_101),
.A2(n_91),
.B(n_30),
.Y(n_121)
);

AOI21xp5_ASAP7_75t_L g130 ( 
.A1(n_121),
.A2(n_126),
.B(n_0),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_107),
.B(n_53),
.C(n_71),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_122),
.B(n_0),
.C(n_1),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_103),
.B(n_65),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_124),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_139)
);

OR2x4_ASAP7_75t_L g126 ( 
.A(n_99),
.B(n_72),
.Y(n_126)
);

BUFx3_ASAP7_75t_L g128 ( 
.A(n_123),
.Y(n_128)
);

BUFx3_ASAP7_75t_L g141 ( 
.A(n_128),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_129),
.A2(n_134),
.B1(n_125),
.B2(n_8),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_SL g148 ( 
.A1(n_130),
.A2(n_131),
.B(n_135),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_115),
.A2(n_76),
.B1(n_63),
.B2(n_57),
.Y(n_131)
);

XOR2xp5_ASAP7_75t_L g132 ( 
.A(n_111),
.B(n_72),
.Y(n_132)
);

XOR2xp5_ASAP7_75t_L g140 ( 
.A(n_132),
.B(n_133),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_114),
.A2(n_2),
.B1(n_5),
.B2(n_6),
.Y(n_134)
);

AOI21xp5_ASAP7_75t_L g135 ( 
.A1(n_126),
.A2(n_22),
.B(n_43),
.Y(n_135)
);

AOI21xp5_ASAP7_75t_L g137 ( 
.A1(n_120),
.A2(n_20),
.B(n_42),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_L g146 ( 
.A(n_137),
.B(n_122),
.Y(n_146)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_117),
.Y(n_138)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_138),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_139),
.B(n_121),
.Y(n_145)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_136),
.Y(n_143)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_143),
.Y(n_154)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_128),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_144),
.A2(n_147),
.B1(n_125),
.B2(n_8),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_SL g150 ( 
.A1(n_145),
.A2(n_146),
.B(n_149),
.Y(n_150)
);

CKINVDCx16_ASAP7_75t_R g149 ( 
.A(n_127),
.Y(n_149)
);

OAI22x1_ASAP7_75t_L g151 ( 
.A1(n_148),
.A2(n_131),
.B1(n_132),
.B2(n_123),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_151),
.A2(n_152),
.B1(n_153),
.B2(n_141),
.Y(n_156)
);

NAND2xp33_ASAP7_75t_SL g152 ( 
.A(n_145),
.B(n_113),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_150),
.B(n_140),
.C(n_142),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_L g157 ( 
.A(n_155),
.B(n_156),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_157),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_158),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_159),
.B(n_154),
.C(n_151),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_160),
.B(n_141),
.Y(n_161)
);

BUFx24_ASAP7_75t_SL g162 ( 
.A(n_161),
.Y(n_162)
);

AOI21x1_ASAP7_75t_SL g163 ( 
.A1(n_162),
.A2(n_27),
.B(n_49),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_163),
.B(n_26),
.Y(n_164)
);

AOI321xp33_ASAP7_75t_L g165 ( 
.A1(n_164),
.A2(n_35),
.A3(n_41),
.B1(n_38),
.B2(n_14),
.C(n_18),
.Y(n_165)
);

OA21x2_ASAP7_75t_L g166 ( 
.A1(n_165),
.A2(n_36),
.B(n_116),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_L g167 ( 
.A1(n_166),
.A2(n_7),
.B(n_9),
.Y(n_167)
);

XOR2xp5_ASAP7_75t_L g168 ( 
.A(n_167),
.B(n_10),
.Y(n_168)
);


endmodule