module fake_aes_10820_n_685 (n_44, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_6, n_4, n_40, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_685);
input n_44;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_6;
input n_4;
input n_40;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_685;
wire n_117;
wire n_663;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_672;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_476;
wire n_105;
wire n_227;
wire n_384;
wire n_434;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_360;
wire n_345;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_647;
wire n_367;
wire n_644;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_648;
wire n_613;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_243;
wire n_235;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_77;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_420;
wire n_165;
wire n_195;
wire n_423;
wire n_342;
wire n_446;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_357;
wire n_90;
wire n_653;
wire n_260;
wire n_78;
wire n_539;
wire n_201;
wire n_197;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_522;
wire n_264;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_684;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_618;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_84;
wire n_266;
wire n_683;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_444;
wire n_176;
wire n_521;
wire n_650;
wire n_625;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_261;
wire n_110;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_132;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
CKINVDCx5p33_ASAP7_75t_R g77 ( .A(n_37), .Y(n_77) );
CKINVDCx5p33_ASAP7_75t_R g78 ( .A(n_0), .Y(n_78) );
INVx2_ASAP7_75t_L g79 ( .A(n_18), .Y(n_79) );
INVxp67_ASAP7_75t_L g80 ( .A(n_38), .Y(n_80) );
INVx1_ASAP7_75t_L g81 ( .A(n_45), .Y(n_81) );
INVx1_ASAP7_75t_L g82 ( .A(n_63), .Y(n_82) );
INVxp67_ASAP7_75t_SL g83 ( .A(n_0), .Y(n_83) );
INVx1_ASAP7_75t_L g84 ( .A(n_9), .Y(n_84) );
OR2x2_ASAP7_75t_L g85 ( .A(n_64), .B(n_9), .Y(n_85) );
CKINVDCx5p33_ASAP7_75t_R g86 ( .A(n_16), .Y(n_86) );
INVx1_ASAP7_75t_L g87 ( .A(n_53), .Y(n_87) );
INVxp67_ASAP7_75t_L g88 ( .A(n_27), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_1), .Y(n_89) );
INVxp67_ASAP7_75t_SL g90 ( .A(n_8), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_74), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_34), .Y(n_92) );
INVx1_ASAP7_75t_L g93 ( .A(n_56), .Y(n_93) );
INVx1_ASAP7_75t_L g94 ( .A(n_61), .Y(n_94) );
INVxp33_ASAP7_75t_L g95 ( .A(n_59), .Y(n_95) );
INVxp67_ASAP7_75t_L g96 ( .A(n_23), .Y(n_96) );
CKINVDCx16_ASAP7_75t_R g97 ( .A(n_66), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_2), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_67), .Y(n_99) );
CKINVDCx5p33_ASAP7_75t_R g100 ( .A(n_54), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_71), .Y(n_101) );
BUFx2_ASAP7_75t_L g102 ( .A(n_20), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_10), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_24), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_75), .Y(n_105) );
CKINVDCx5p33_ASAP7_75t_R g106 ( .A(n_52), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_47), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_11), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_41), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_19), .Y(n_110) );
INVx2_ASAP7_75t_L g111 ( .A(n_3), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_51), .Y(n_112) );
HB1xp67_ASAP7_75t_L g113 ( .A(n_5), .Y(n_113) );
INVxp67_ASAP7_75t_SL g114 ( .A(n_35), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_17), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_32), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_49), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_73), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_33), .Y(n_119) );
CKINVDCx14_ASAP7_75t_R g120 ( .A(n_5), .Y(n_120) );
INVxp67_ASAP7_75t_SL g121 ( .A(n_10), .Y(n_121) );
INVxp67_ASAP7_75t_SL g122 ( .A(n_58), .Y(n_122) );
INVxp33_ASAP7_75t_SL g123 ( .A(n_39), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_81), .Y(n_124) );
INVx1_ASAP7_75t_L g125 ( .A(n_81), .Y(n_125) );
INVx3_ASAP7_75t_L g126 ( .A(n_79), .Y(n_126) );
INVx1_ASAP7_75t_L g127 ( .A(n_82), .Y(n_127) );
INVx3_ASAP7_75t_L g128 ( .A(n_79), .Y(n_128) );
BUFx2_ASAP7_75t_L g129 ( .A(n_120), .Y(n_129) );
NAND2xp5_ASAP7_75t_L g130 ( .A(n_102), .B(n_1), .Y(n_130) );
AOI22xp5_ASAP7_75t_L g131 ( .A1(n_97), .A2(n_2), .B1(n_3), .B2(n_4), .Y(n_131) );
NAND2xp5_ASAP7_75t_L g132 ( .A(n_102), .B(n_4), .Y(n_132) );
INVx1_ASAP7_75t_L g133 ( .A(n_82), .Y(n_133) );
NAND2xp5_ASAP7_75t_SL g134 ( .A(n_87), .B(n_6), .Y(n_134) );
INVx2_ASAP7_75t_L g135 ( .A(n_87), .Y(n_135) );
INVx1_ASAP7_75t_L g136 ( .A(n_91), .Y(n_136) );
INVx2_ASAP7_75t_L g137 ( .A(n_91), .Y(n_137) );
INVx1_ASAP7_75t_L g138 ( .A(n_92), .Y(n_138) );
OR2x2_ASAP7_75t_L g139 ( .A(n_113), .B(n_6), .Y(n_139) );
BUFx6f_ASAP7_75t_L g140 ( .A(n_92), .Y(n_140) );
INVx2_ASAP7_75t_L g141 ( .A(n_93), .Y(n_141) );
AND2x2_ASAP7_75t_L g142 ( .A(n_95), .B(n_7), .Y(n_142) );
NAND2xp5_ASAP7_75t_L g143 ( .A(n_98), .B(n_7), .Y(n_143) );
INVx2_ASAP7_75t_L g144 ( .A(n_93), .Y(n_144) );
CKINVDCx20_ASAP7_75t_R g145 ( .A(n_78), .Y(n_145) );
INVx1_ASAP7_75t_L g146 ( .A(n_94), .Y(n_146) );
XNOR2xp5_ASAP7_75t_L g147 ( .A(n_86), .B(n_8), .Y(n_147) );
INVx2_ASAP7_75t_L g148 ( .A(n_94), .Y(n_148) );
INVx1_ASAP7_75t_L g149 ( .A(n_99), .Y(n_149) );
INVx3_ASAP7_75t_L g150 ( .A(n_111), .Y(n_150) );
NOR2xp33_ASAP7_75t_L g151 ( .A(n_101), .B(n_11), .Y(n_151) );
AND2x2_ASAP7_75t_L g152 ( .A(n_111), .B(n_12), .Y(n_152) );
INVx1_ASAP7_75t_L g153 ( .A(n_99), .Y(n_153) );
INVx1_ASAP7_75t_L g154 ( .A(n_105), .Y(n_154) );
AND2x6_ASAP7_75t_L g155 ( .A(n_105), .B(n_40), .Y(n_155) );
INVx1_ASAP7_75t_L g156 ( .A(n_107), .Y(n_156) );
BUFx6f_ASAP7_75t_L g157 ( .A(n_107), .Y(n_157) );
BUFx6f_ASAP7_75t_L g158 ( .A(n_109), .Y(n_158) );
NOR2xp33_ASAP7_75t_L g159 ( .A(n_104), .B(n_12), .Y(n_159) );
XNOR2xp5_ASAP7_75t_L g160 ( .A(n_83), .B(n_13), .Y(n_160) );
INVx1_ASAP7_75t_L g161 ( .A(n_109), .Y(n_161) );
INVx5_ASAP7_75t_L g162 ( .A(n_114), .Y(n_162) );
OA21x2_ASAP7_75t_L g163 ( .A1(n_112), .A2(n_42), .B(n_72), .Y(n_163) );
BUFx6f_ASAP7_75t_L g164 ( .A(n_112), .Y(n_164) );
INVx2_ASAP7_75t_L g165 ( .A(n_116), .Y(n_165) );
NAND2xp5_ASAP7_75t_L g166 ( .A(n_129), .B(n_106), .Y(n_166) );
BUFx6f_ASAP7_75t_L g167 ( .A(n_163), .Y(n_167) );
AND2x2_ASAP7_75t_L g168 ( .A(n_129), .B(n_115), .Y(n_168) );
INVx1_ASAP7_75t_L g169 ( .A(n_140), .Y(n_169) );
INVx2_ASAP7_75t_L g170 ( .A(n_140), .Y(n_170) );
INVx2_ASAP7_75t_L g171 ( .A(n_140), .Y(n_171) );
NAND2xp5_ASAP7_75t_L g172 ( .A(n_124), .B(n_77), .Y(n_172) );
INVx1_ASAP7_75t_L g173 ( .A(n_140), .Y(n_173) );
INVx3_ASAP7_75t_L g174 ( .A(n_140), .Y(n_174) );
BUFx3_ASAP7_75t_L g175 ( .A(n_155), .Y(n_175) );
NOR2xp33_ASAP7_75t_L g176 ( .A(n_124), .B(n_80), .Y(n_176) );
NAND2xp5_ASAP7_75t_SL g177 ( .A(n_162), .B(n_96), .Y(n_177) );
INVx2_ASAP7_75t_L g178 ( .A(n_140), .Y(n_178) );
INVx1_ASAP7_75t_L g179 ( .A(n_157), .Y(n_179) );
INVx1_ASAP7_75t_L g180 ( .A(n_157), .Y(n_180) );
NAND2xp5_ASAP7_75t_L g181 ( .A(n_125), .B(n_100), .Y(n_181) );
AND2x2_ASAP7_75t_L g182 ( .A(n_142), .B(n_84), .Y(n_182) );
INVx3_ASAP7_75t_L g183 ( .A(n_157), .Y(n_183) );
BUFx6f_ASAP7_75t_L g184 ( .A(n_163), .Y(n_184) );
BUFx6f_ASAP7_75t_L g185 ( .A(n_163), .Y(n_185) );
INVx1_ASAP7_75t_L g186 ( .A(n_157), .Y(n_186) );
OAI22xp5_ASAP7_75t_SL g187 ( .A1(n_160), .A2(n_147), .B1(n_145), .B2(n_131), .Y(n_187) );
AND3x4_ASAP7_75t_L g188 ( .A(n_160), .B(n_121), .C(n_90), .Y(n_188) );
NAND2xp5_ASAP7_75t_L g189 ( .A(n_125), .B(n_88), .Y(n_189) );
INVx4_ASAP7_75t_L g190 ( .A(n_155), .Y(n_190) );
BUFx3_ASAP7_75t_L g191 ( .A(n_155), .Y(n_191) );
BUFx3_ASAP7_75t_L g192 ( .A(n_155), .Y(n_192) );
INVx3_ASAP7_75t_L g193 ( .A(n_157), .Y(n_193) );
INVx1_ASAP7_75t_L g194 ( .A(n_157), .Y(n_194) );
INVx3_ASAP7_75t_L g195 ( .A(n_158), .Y(n_195) );
AND2x2_ASAP7_75t_L g196 ( .A(n_142), .B(n_84), .Y(n_196) );
BUFx6f_ASAP7_75t_L g197 ( .A(n_163), .Y(n_197) );
AND2x6_ASAP7_75t_L g198 ( .A(n_152), .B(n_117), .Y(n_198) );
INVx1_ASAP7_75t_L g199 ( .A(n_158), .Y(n_199) );
AND2x2_ASAP7_75t_L g200 ( .A(n_127), .B(n_89), .Y(n_200) );
BUFx6f_ASAP7_75t_L g201 ( .A(n_158), .Y(n_201) );
NAND2xp5_ASAP7_75t_L g202 ( .A(n_127), .B(n_116), .Y(n_202) );
INVx1_ASAP7_75t_L g203 ( .A(n_158), .Y(n_203) );
INVx1_ASAP7_75t_L g204 ( .A(n_158), .Y(n_204) );
BUFx6f_ASAP7_75t_L g205 ( .A(n_158), .Y(n_205) );
AOI22xp33_ASAP7_75t_L g206 ( .A1(n_152), .A2(n_155), .B1(n_139), .B2(n_156), .Y(n_206) );
NAND2x1p5_ASAP7_75t_L g207 ( .A(n_133), .B(n_85), .Y(n_207) );
INVx1_ASAP7_75t_L g208 ( .A(n_164), .Y(n_208) );
AND2x4_ASAP7_75t_L g209 ( .A(n_133), .B(n_136), .Y(n_209) );
INVx1_ASAP7_75t_L g210 ( .A(n_164), .Y(n_210) );
OR2x6_ASAP7_75t_L g211 ( .A(n_139), .B(n_85), .Y(n_211) );
INVx1_ASAP7_75t_L g212 ( .A(n_164), .Y(n_212) );
INVx1_ASAP7_75t_L g213 ( .A(n_164), .Y(n_213) );
AND2x4_ASAP7_75t_L g214 ( .A(n_136), .B(n_89), .Y(n_214) );
AND2x2_ASAP7_75t_L g215 ( .A(n_138), .B(n_103), .Y(n_215) );
AND2x4_ASAP7_75t_L g216 ( .A(n_138), .B(n_103), .Y(n_216) );
NOR2xp33_ASAP7_75t_L g217 ( .A(n_146), .B(n_123), .Y(n_217) );
NAND2xp5_ASAP7_75t_SL g218 ( .A(n_162), .B(n_119), .Y(n_218) );
INVx2_ASAP7_75t_L g219 ( .A(n_164), .Y(n_219) );
NAND2xp5_ASAP7_75t_L g220 ( .A(n_146), .B(n_119), .Y(n_220) );
NAND2x1p5_ASAP7_75t_L g221 ( .A(n_149), .B(n_118), .Y(n_221) );
INVx4_ASAP7_75t_L g222 ( .A(n_155), .Y(n_222) );
INVx1_ASAP7_75t_L g223 ( .A(n_164), .Y(n_223) );
NAND2xp5_ASAP7_75t_SL g224 ( .A(n_162), .B(n_118), .Y(n_224) );
INVx2_ASAP7_75t_L g225 ( .A(n_135), .Y(n_225) );
NOR2xp33_ASAP7_75t_L g226 ( .A(n_149), .B(n_117), .Y(n_226) );
INVx2_ASAP7_75t_L g227 ( .A(n_225), .Y(n_227) );
HB1xp67_ASAP7_75t_L g228 ( .A(n_211), .Y(n_228) );
BUFx2_ASAP7_75t_L g229 ( .A(n_198), .Y(n_229) );
NAND2xp5_ASAP7_75t_SL g230 ( .A(n_190), .B(n_162), .Y(n_230) );
NAND2xp5_ASAP7_75t_L g231 ( .A(n_209), .B(n_153), .Y(n_231) );
AND2x4_ASAP7_75t_L g232 ( .A(n_211), .B(n_130), .Y(n_232) );
HB1xp67_ASAP7_75t_L g233 ( .A(n_211), .Y(n_233) );
INVx1_ASAP7_75t_L g234 ( .A(n_209), .Y(n_234) );
NAND2xp5_ASAP7_75t_L g235 ( .A(n_209), .B(n_156), .Y(n_235) );
INVx1_ASAP7_75t_L g236 ( .A(n_209), .Y(n_236) );
BUFx4f_ASAP7_75t_L g237 ( .A(n_198), .Y(n_237) );
NAND2xp5_ASAP7_75t_SL g238 ( .A(n_190), .B(n_162), .Y(n_238) );
NAND2xp5_ASAP7_75t_L g239 ( .A(n_217), .B(n_153), .Y(n_239) );
INVx1_ASAP7_75t_L g240 ( .A(n_225), .Y(n_240) );
INVx1_ASAP7_75t_L g241 ( .A(n_221), .Y(n_241) );
NAND2xp5_ASAP7_75t_L g242 ( .A(n_172), .B(n_161), .Y(n_242) );
INVx1_ASAP7_75t_L g243 ( .A(n_221), .Y(n_243) );
INVx2_ASAP7_75t_L g244 ( .A(n_201), .Y(n_244) );
INVx1_ASAP7_75t_L g245 ( .A(n_221), .Y(n_245) );
AND2x4_ASAP7_75t_L g246 ( .A(n_211), .B(n_132), .Y(n_246) );
NOR2xp33_ASAP7_75t_L g247 ( .A(n_166), .B(n_162), .Y(n_247) );
NAND2xp5_ASAP7_75t_L g248 ( .A(n_181), .B(n_161), .Y(n_248) );
BUFx2_ASAP7_75t_L g249 ( .A(n_198), .Y(n_249) );
NOR2xp33_ASAP7_75t_R g250 ( .A(n_206), .B(n_147), .Y(n_250) );
INVx2_ASAP7_75t_L g251 ( .A(n_201), .Y(n_251) );
CKINVDCx5p33_ASAP7_75t_R g252 ( .A(n_211), .Y(n_252) );
BUFx4f_ASAP7_75t_L g253 ( .A(n_198), .Y(n_253) );
AND2x4_ASAP7_75t_L g254 ( .A(n_182), .B(n_154), .Y(n_254) );
BUFx3_ASAP7_75t_L g255 ( .A(n_191), .Y(n_255) );
INVx1_ASAP7_75t_L g256 ( .A(n_214), .Y(n_256) );
INVx2_ASAP7_75t_L g257 ( .A(n_201), .Y(n_257) );
AND2x4_ASAP7_75t_SL g258 ( .A(n_190), .B(n_222), .Y(n_258) );
BUFx3_ASAP7_75t_L g259 ( .A(n_191), .Y(n_259) );
AND2x2_ASAP7_75t_L g260 ( .A(n_207), .B(n_154), .Y(n_260) );
AND2x2_ASAP7_75t_L g261 ( .A(n_207), .B(n_165), .Y(n_261) );
BUFx3_ASAP7_75t_L g262 ( .A(n_191), .Y(n_262) );
INVx1_ASAP7_75t_L g263 ( .A(n_214), .Y(n_263) );
INVx2_ASAP7_75t_L g264 ( .A(n_201), .Y(n_264) );
NOR2xp33_ASAP7_75t_L g265 ( .A(n_168), .B(n_143), .Y(n_265) );
NAND2xp5_ASAP7_75t_L g266 ( .A(n_189), .B(n_159), .Y(n_266) );
AOI21xp33_ASAP7_75t_L g267 ( .A1(n_182), .A2(n_151), .B(n_134), .Y(n_267) );
CKINVDCx5p33_ASAP7_75t_R g268 ( .A(n_187), .Y(n_268) );
INVx3_ASAP7_75t_L g269 ( .A(n_214), .Y(n_269) );
BUFx6f_ASAP7_75t_L g270 ( .A(n_175), .Y(n_270) );
BUFx2_ASAP7_75t_L g271 ( .A(n_198), .Y(n_271) );
NAND2xp5_ASAP7_75t_L g272 ( .A(n_196), .B(n_165), .Y(n_272) );
INVx1_ASAP7_75t_L g273 ( .A(n_214), .Y(n_273) );
INVx1_ASAP7_75t_L g274 ( .A(n_216), .Y(n_274) );
INVx2_ASAP7_75t_L g275 ( .A(n_201), .Y(n_275) );
INVx2_ASAP7_75t_L g276 ( .A(n_205), .Y(n_276) );
NAND2xp5_ASAP7_75t_L g277 ( .A(n_196), .B(n_165), .Y(n_277) );
INVxp67_ASAP7_75t_L g278 ( .A(n_168), .Y(n_278) );
NAND2xp5_ASAP7_75t_L g279 ( .A(n_198), .B(n_135), .Y(n_279) );
INVx1_ASAP7_75t_L g280 ( .A(n_216), .Y(n_280) );
NAND2xp5_ASAP7_75t_L g281 ( .A(n_198), .B(n_135), .Y(n_281) );
AOI22xp33_ASAP7_75t_L g282 ( .A1(n_216), .A2(n_155), .B1(n_137), .B2(n_148), .Y(n_282) );
OAI21xp5_ASAP7_75t_L g283 ( .A1(n_176), .A2(n_155), .B(n_148), .Y(n_283) );
INVx5_ASAP7_75t_L g284 ( .A(n_190), .Y(n_284) );
AND2x6_ASAP7_75t_SL g285 ( .A(n_188), .B(n_108), .Y(n_285) );
INVx3_ASAP7_75t_L g286 ( .A(n_216), .Y(n_286) );
OAI21x1_ASAP7_75t_L g287 ( .A1(n_202), .A2(n_137), .B(n_148), .Y(n_287) );
INVx1_ASAP7_75t_L g288 ( .A(n_200), .Y(n_288) );
NAND2xp5_ASAP7_75t_L g289 ( .A(n_207), .B(n_137), .Y(n_289) );
INVx1_ASAP7_75t_L g290 ( .A(n_200), .Y(n_290) );
INVx1_ASAP7_75t_SL g291 ( .A(n_261), .Y(n_291) );
INVx3_ASAP7_75t_L g292 ( .A(n_286), .Y(n_292) );
AND2x4_ASAP7_75t_L g293 ( .A(n_254), .B(n_215), .Y(n_293) );
BUFx3_ASAP7_75t_L g294 ( .A(n_237), .Y(n_294) );
NOR2xp33_ASAP7_75t_L g295 ( .A(n_232), .B(n_222), .Y(n_295) );
NAND2xp5_ASAP7_75t_L g296 ( .A(n_260), .B(n_215), .Y(n_296) );
BUFx2_ASAP7_75t_L g297 ( .A(n_252), .Y(n_297) );
AND2x6_ASAP7_75t_L g298 ( .A(n_241), .B(n_175), .Y(n_298) );
AND2x2_ASAP7_75t_SL g299 ( .A(n_237), .B(n_222), .Y(n_299) );
INVx4_ASAP7_75t_L g300 ( .A(n_237), .Y(n_300) );
O2A1O1Ixp33_ASAP7_75t_L g301 ( .A1(n_278), .A2(n_220), .B(n_226), .C(n_224), .Y(n_301) );
NAND2xp5_ASAP7_75t_L g302 ( .A(n_260), .B(n_222), .Y(n_302) );
BUFx3_ASAP7_75t_L g303 ( .A(n_253), .Y(n_303) );
INVx5_ASAP7_75t_L g304 ( .A(n_229), .Y(n_304) );
INVx1_ASAP7_75t_L g305 ( .A(n_256), .Y(n_305) );
AOI221xp5_ASAP7_75t_L g306 ( .A1(n_265), .A2(n_187), .B1(n_188), .B2(n_115), .C(n_108), .Y(n_306) );
INVx1_ASAP7_75t_L g307 ( .A(n_256), .Y(n_307) );
HB1xp67_ASAP7_75t_L g308 ( .A(n_241), .Y(n_308) );
BUFx6f_ASAP7_75t_L g309 ( .A(n_255), .Y(n_309) );
OR2x6_ASAP7_75t_L g310 ( .A(n_228), .B(n_188), .Y(n_310) );
INVx2_ASAP7_75t_L g311 ( .A(n_286), .Y(n_311) );
INVx1_ASAP7_75t_L g312 ( .A(n_263), .Y(n_312) );
NAND2xp5_ASAP7_75t_L g313 ( .A(n_261), .B(n_192), .Y(n_313) );
INVx4_ASAP7_75t_L g314 ( .A(n_253), .Y(n_314) );
INVx3_ASAP7_75t_L g315 ( .A(n_286), .Y(n_315) );
BUFx5_ASAP7_75t_L g316 ( .A(n_243), .Y(n_316) );
NOR2x1_ASAP7_75t_L g317 ( .A(n_232), .B(n_177), .Y(n_317) );
O2A1O1Ixp33_ASAP7_75t_L g318 ( .A1(n_288), .A2(n_218), .B(n_141), .C(n_144), .Y(n_318) );
INVx2_ASAP7_75t_SL g319 ( .A(n_254), .Y(n_319) );
NAND2xp5_ASAP7_75t_L g320 ( .A(n_254), .B(n_192), .Y(n_320) );
BUFx6f_ASAP7_75t_L g321 ( .A(n_255), .Y(n_321) );
OAI22xp5_ASAP7_75t_L g322 ( .A1(n_243), .A2(n_141), .B1(n_144), .B2(n_185), .Y(n_322) );
INVx2_ASAP7_75t_L g323 ( .A(n_227), .Y(n_323) );
INVxp67_ASAP7_75t_L g324 ( .A(n_233), .Y(n_324) );
OR2x2_ASAP7_75t_L g325 ( .A(n_268), .B(n_126), .Y(n_325) );
AOI22xp5_ASAP7_75t_SL g326 ( .A1(n_252), .A2(n_122), .B1(n_110), .B2(n_126), .Y(n_326) );
AOI222xp33_ASAP7_75t_L g327 ( .A1(n_268), .A2(n_110), .B1(n_126), .B2(n_150), .C1(n_128), .C2(n_144), .Y(n_327) );
HB1xp67_ASAP7_75t_L g328 ( .A(n_245), .Y(n_328) );
AOI21xp5_ASAP7_75t_L g329 ( .A1(n_283), .A2(n_242), .B(n_248), .Y(n_329) );
INVx2_ASAP7_75t_L g330 ( .A(n_227), .Y(n_330) );
BUFx2_ASAP7_75t_L g331 ( .A(n_285), .Y(n_331) );
AOI22xp33_ASAP7_75t_L g332 ( .A1(n_288), .A2(n_141), .B1(n_197), .B2(n_167), .Y(n_332) );
INVx1_ASAP7_75t_L g333 ( .A(n_263), .Y(n_333) );
OAI22xp33_ASAP7_75t_L g334 ( .A1(n_253), .A2(n_126), .B1(n_150), .B2(n_128), .Y(n_334) );
INVx1_ASAP7_75t_SL g335 ( .A(n_254), .Y(n_335) );
INVx1_ASAP7_75t_L g336 ( .A(n_273), .Y(n_336) );
BUFx2_ASAP7_75t_SL g337 ( .A(n_245), .Y(n_337) );
AOI21xp5_ASAP7_75t_L g338 ( .A1(n_230), .A2(n_167), .B(n_184), .Y(n_338) );
CKINVDCx11_ASAP7_75t_R g339 ( .A(n_285), .Y(n_339) );
INVx1_ASAP7_75t_L g340 ( .A(n_273), .Y(n_340) );
NAND2xp5_ASAP7_75t_L g341 ( .A(n_296), .B(n_291), .Y(n_341) );
NOR2xp67_ASAP7_75t_L g342 ( .A(n_308), .B(n_286), .Y(n_342) );
INVxp67_ASAP7_75t_SL g343 ( .A(n_308), .Y(n_343) );
INVx3_ASAP7_75t_L g344 ( .A(n_316), .Y(n_344) );
INVx2_ASAP7_75t_L g345 ( .A(n_323), .Y(n_345) );
INVx2_ASAP7_75t_L g346 ( .A(n_323), .Y(n_346) );
INVx3_ASAP7_75t_SL g347 ( .A(n_316), .Y(n_347) );
AOI22xp33_ASAP7_75t_L g348 ( .A1(n_306), .A2(n_310), .B1(n_250), .B2(n_232), .Y(n_348) );
OAI22xp5_ASAP7_75t_L g349 ( .A1(n_337), .A2(n_246), .B1(n_232), .B2(n_289), .Y(n_349) );
NOR2xp33_ASAP7_75t_L g350 ( .A(n_310), .B(n_297), .Y(n_350) );
AOI22xp5_ASAP7_75t_L g351 ( .A1(n_310), .A2(n_246), .B1(n_290), .B2(n_274), .Y(n_351) );
AOI21xp5_ASAP7_75t_L g352 ( .A1(n_338), .A2(n_238), .B(n_239), .Y(n_352) );
INVx2_ASAP7_75t_L g353 ( .A(n_330), .Y(n_353) );
NAND2xp5_ASAP7_75t_L g354 ( .A(n_293), .B(n_246), .Y(n_354) );
AOI22xp33_ASAP7_75t_L g355 ( .A1(n_331), .A2(n_246), .B1(n_229), .B2(n_249), .Y(n_355) );
AOI22xp5_ASAP7_75t_L g356 ( .A1(n_335), .A2(n_290), .B1(n_280), .B2(n_274), .Y(n_356) );
INVx2_ASAP7_75t_SL g357 ( .A(n_316), .Y(n_357) );
OAI22xp5_ASAP7_75t_SL g358 ( .A1(n_325), .A2(n_266), .B1(n_272), .B2(n_277), .Y(n_358) );
AOI22xp33_ASAP7_75t_L g359 ( .A1(n_293), .A2(n_249), .B1(n_271), .B2(n_269), .Y(n_359) );
INVx1_ASAP7_75t_L g360 ( .A(n_305), .Y(n_360) );
CKINVDCx20_ASAP7_75t_R g361 ( .A(n_339), .Y(n_361) );
OAI22xp5_ASAP7_75t_L g362 ( .A1(n_328), .A2(n_271), .B1(n_235), .B2(n_231), .Y(n_362) );
AOI22xp33_ASAP7_75t_L g363 ( .A1(n_319), .A2(n_269), .B1(n_236), .B2(n_234), .Y(n_363) );
INVxp67_ASAP7_75t_L g364 ( .A(n_328), .Y(n_364) );
AND2x4_ASAP7_75t_L g365 ( .A(n_300), .B(n_234), .Y(n_365) );
INVx2_ASAP7_75t_L g366 ( .A(n_330), .Y(n_366) );
OAI22xp5_ASAP7_75t_L g367 ( .A1(n_334), .A2(n_280), .B1(n_269), .B2(n_236), .Y(n_367) );
OAI22xp33_ASAP7_75t_L g368 ( .A1(n_324), .A2(n_279), .B1(n_281), .B2(n_267), .Y(n_368) );
OAI22xp5_ASAP7_75t_L g369 ( .A1(n_334), .A2(n_282), .B1(n_240), .B2(n_259), .Y(n_369) );
INVx1_ASAP7_75t_L g370 ( .A(n_307), .Y(n_370) );
NAND2xp5_ASAP7_75t_L g371 ( .A(n_324), .B(n_240), .Y(n_371) );
OR2x2_ASAP7_75t_L g372 ( .A(n_341), .B(n_287), .Y(n_372) );
NAND2xp5_ASAP7_75t_L g373 ( .A(n_360), .B(n_329), .Y(n_373) );
AO31x2_ASAP7_75t_L g374 ( .A1(n_369), .A2(n_322), .A3(n_336), .B(n_333), .Y(n_374) );
INVx1_ASAP7_75t_L g375 ( .A(n_360), .Y(n_375) );
CKINVDCx5p33_ASAP7_75t_R g376 ( .A(n_361), .Y(n_376) );
OAI211xp5_ASAP7_75t_L g377 ( .A1(n_348), .A2(n_327), .B(n_339), .C(n_301), .Y(n_377) );
INVxp67_ASAP7_75t_L g378 ( .A(n_343), .Y(n_378) );
AOI22xp33_ASAP7_75t_L g379 ( .A1(n_358), .A2(n_295), .B1(n_317), .B2(n_340), .Y(n_379) );
AND2x2_ASAP7_75t_L g380 ( .A(n_345), .B(n_316), .Y(n_380) );
AOI22xp33_ASAP7_75t_L g381 ( .A1(n_351), .A2(n_295), .B1(n_312), .B2(n_292), .Y(n_381) );
AOI22xp33_ASAP7_75t_SL g382 ( .A1(n_350), .A2(n_326), .B1(n_316), .B2(n_304), .Y(n_382) );
INVx1_ASAP7_75t_L g383 ( .A(n_370), .Y(n_383) );
CKINVDCx5p33_ASAP7_75t_R g384 ( .A(n_361), .Y(n_384) );
HB1xp67_ASAP7_75t_L g385 ( .A(n_364), .Y(n_385) );
AOI22xp33_ASAP7_75t_L g386 ( .A1(n_351), .A2(n_292), .B1(n_315), .B2(n_311), .Y(n_386) );
AOI222xp33_ASAP7_75t_L g387 ( .A1(n_370), .A2(n_128), .B1(n_150), .B2(n_320), .C1(n_302), .C2(n_315), .Y(n_387) );
AOI21xp33_ASAP7_75t_L g388 ( .A1(n_368), .A2(n_318), .B(n_287), .Y(n_388) );
OAI22xp5_ASAP7_75t_L g389 ( .A1(n_356), .A2(n_332), .B1(n_313), .B2(n_304), .Y(n_389) );
OAI22xp5_ASAP7_75t_L g390 ( .A1(n_356), .A2(n_332), .B1(n_304), .B2(n_299), .Y(n_390) );
AND2x2_ASAP7_75t_L g391 ( .A(n_345), .B(n_316), .Y(n_391) );
OAI21x1_ASAP7_75t_L g392 ( .A1(n_352), .A2(n_344), .B(n_366), .Y(n_392) );
A2O1A1Ixp33_ASAP7_75t_L g393 ( .A1(n_342), .A2(n_247), .B(n_299), .C(n_294), .Y(n_393) );
AOI22xp33_ASAP7_75t_L g394 ( .A1(n_349), .A2(n_304), .B1(n_300), .B2(n_314), .Y(n_394) );
AND2x2_ASAP7_75t_L g395 ( .A(n_346), .B(n_309), .Y(n_395) );
AOI22xp33_ASAP7_75t_L g396 ( .A1(n_354), .A2(n_314), .B1(n_303), .B2(n_294), .Y(n_396) );
INVx1_ASAP7_75t_L g397 ( .A(n_346), .Y(n_397) );
OAI211xp5_ASAP7_75t_SL g398 ( .A1(n_355), .A2(n_128), .B(n_150), .C(n_199), .Y(n_398) );
OAI332xp33_ASAP7_75t_SL g399 ( .A1(n_375), .A2(n_367), .A3(n_362), .B1(n_15), .B2(n_16), .B3(n_13), .C1(n_18), .C2(n_19), .Y(n_399) );
INVx2_ASAP7_75t_L g400 ( .A(n_397), .Y(n_400) );
NAND3xp33_ASAP7_75t_L g401 ( .A(n_379), .B(n_342), .C(n_366), .Y(n_401) );
INVx1_ASAP7_75t_L g402 ( .A(n_375), .Y(n_402) );
INVxp67_ASAP7_75t_L g403 ( .A(n_385), .Y(n_403) );
NOR4xp25_ASAP7_75t_L g404 ( .A(n_377), .B(n_371), .C(n_353), .D(n_344), .Y(n_404) );
AOI22xp33_ASAP7_75t_L g405 ( .A1(n_387), .A2(n_365), .B1(n_347), .B2(n_363), .Y(n_405) );
AND2x2_ASAP7_75t_L g406 ( .A(n_397), .B(n_353), .Y(n_406) );
INVx2_ASAP7_75t_L g407 ( .A(n_392), .Y(n_407) );
INVx1_ASAP7_75t_L g408 ( .A(n_383), .Y(n_408) );
INVx1_ASAP7_75t_L g409 ( .A(n_383), .Y(n_409) );
INVx2_ASAP7_75t_L g410 ( .A(n_392), .Y(n_410) );
NAND2xp5_ASAP7_75t_SL g411 ( .A(n_378), .B(n_347), .Y(n_411) );
OAI21x1_ASAP7_75t_L g412 ( .A1(n_373), .A2(n_344), .B(n_171), .Y(n_412) );
AND2x2_ASAP7_75t_L g413 ( .A(n_380), .B(n_357), .Y(n_413) );
INVx1_ASAP7_75t_L g414 ( .A(n_372), .Y(n_414) );
AOI22xp33_ASAP7_75t_L g415 ( .A1(n_387), .A2(n_365), .B1(n_347), .B2(n_359), .Y(n_415) );
AOI221xp5_ASAP7_75t_L g416 ( .A1(n_381), .A2(n_365), .B1(n_357), .B2(n_197), .C(n_167), .Y(n_416) );
OAI211xp5_ASAP7_75t_L g417 ( .A1(n_382), .A2(n_376), .B(n_384), .C(n_386), .Y(n_417) );
INVx1_ASAP7_75t_L g418 ( .A(n_372), .Y(n_418) );
HB1xp67_ASAP7_75t_L g419 ( .A(n_380), .Y(n_419) );
AOI221xp5_ASAP7_75t_L g420 ( .A1(n_373), .A2(n_167), .B1(n_184), .B2(n_185), .C(n_197), .Y(n_420) );
OAI22xp5_ASAP7_75t_L g421 ( .A1(n_390), .A2(n_309), .B1(n_321), .B2(n_167), .Y(n_421) );
AOI22xp33_ASAP7_75t_L g422 ( .A1(n_398), .A2(n_321), .B1(n_309), .B2(n_298), .Y(n_422) );
AND2x4_ASAP7_75t_L g423 ( .A(n_391), .B(n_309), .Y(n_423) );
AOI22xp33_ASAP7_75t_L g424 ( .A1(n_390), .A2(n_321), .B1(n_298), .B2(n_303), .Y(n_424) );
NAND3xp33_ASAP7_75t_L g425 ( .A(n_388), .B(n_197), .C(n_185), .Y(n_425) );
INVx1_ASAP7_75t_SL g426 ( .A(n_391), .Y(n_426) );
AOI221xp5_ASAP7_75t_L g427 ( .A1(n_388), .A2(n_184), .B1(n_185), .B2(n_197), .C(n_213), .Y(n_427) );
AOI322xp5_ASAP7_75t_L g428 ( .A1(n_394), .A2(n_14), .A3(n_15), .B1(n_17), .B2(n_185), .C1(n_184), .C2(n_179), .Y(n_428) );
INVx2_ASAP7_75t_L g429 ( .A(n_374), .Y(n_429) );
AOI22xp33_ASAP7_75t_L g430 ( .A1(n_389), .A2(n_321), .B1(n_298), .B2(n_184), .Y(n_430) );
AND2x2_ASAP7_75t_L g431 ( .A(n_395), .B(n_14), .Y(n_431) );
AND2x2_ASAP7_75t_L g432 ( .A(n_395), .B(n_21), .Y(n_432) );
OR2x2_ASAP7_75t_L g433 ( .A(n_374), .B(n_180), .Y(n_433) );
OAI33xp33_ASAP7_75t_L g434 ( .A1(n_403), .A2(n_389), .A3(n_186), .B1(n_208), .B2(n_169), .B3(n_179), .Y(n_434) );
AND2x2_ASAP7_75t_L g435 ( .A(n_400), .B(n_374), .Y(n_435) );
HB1xp67_ASAP7_75t_L g436 ( .A(n_400), .Y(n_436) );
OR2x2_ASAP7_75t_L g437 ( .A(n_414), .B(n_374), .Y(n_437) );
OAI221xp5_ASAP7_75t_SL g438 ( .A1(n_404), .A2(n_396), .B1(n_393), .B2(n_186), .C(n_210), .Y(n_438) );
INVx2_ASAP7_75t_L g439 ( .A(n_400), .Y(n_439) );
OAI221xp5_ASAP7_75t_L g440 ( .A1(n_417), .A2(n_180), .B1(n_173), .B2(n_204), .C(n_199), .Y(n_440) );
INVx1_ASAP7_75t_SL g441 ( .A(n_431), .Y(n_441) );
INVx4_ASAP7_75t_L g442 ( .A(n_423), .Y(n_442) );
INVx3_ASAP7_75t_L g443 ( .A(n_407), .Y(n_443) );
AO21x2_ASAP7_75t_L g444 ( .A1(n_425), .A2(n_374), .B(n_223), .Y(n_444) );
AND2x2_ASAP7_75t_L g445 ( .A(n_414), .B(n_374), .Y(n_445) );
AND2x2_ASAP7_75t_L g446 ( .A(n_418), .B(n_22), .Y(n_446) );
INVx1_ASAP7_75t_L g447 ( .A(n_402), .Y(n_447) );
NAND2xp5_ASAP7_75t_L g448 ( .A(n_402), .B(n_208), .Y(n_448) );
INVx2_ASAP7_75t_L g449 ( .A(n_408), .Y(n_449) );
NAND4xp25_ASAP7_75t_L g450 ( .A(n_428), .B(n_212), .C(n_173), .D(n_169), .Y(n_450) );
AND2x2_ASAP7_75t_L g451 ( .A(n_418), .B(n_25), .Y(n_451) );
NAND2xp5_ASAP7_75t_L g452 ( .A(n_408), .B(n_212), .Y(n_452) );
NOR3xp33_ASAP7_75t_L g453 ( .A(n_411), .B(n_194), .C(n_203), .Y(n_453) );
INVx1_ASAP7_75t_L g454 ( .A(n_409), .Y(n_454) );
NAND3xp33_ASAP7_75t_L g455 ( .A(n_428), .B(n_205), .C(n_203), .Y(n_455) );
AOI22xp5_ASAP7_75t_L g456 ( .A1(n_415), .A2(n_298), .B1(n_223), .B2(n_213), .Y(n_456) );
OAI22xp5_ASAP7_75t_L g457 ( .A1(n_405), .A2(n_298), .B1(n_284), .B2(n_262), .Y(n_457) );
AO21x2_ASAP7_75t_L g458 ( .A1(n_425), .A2(n_194), .B(n_204), .Y(n_458) );
OAI21xp33_ASAP7_75t_L g459 ( .A1(n_404), .A2(n_210), .B(n_171), .Y(n_459) );
AND2x2_ASAP7_75t_L g460 ( .A(n_406), .B(n_26), .Y(n_460) );
AND2x2_ASAP7_75t_L g461 ( .A(n_406), .B(n_28), .Y(n_461) );
NAND2xp5_ASAP7_75t_L g462 ( .A(n_409), .B(n_170), .Y(n_462) );
HB1xp67_ASAP7_75t_L g463 ( .A(n_419), .Y(n_463) );
INVx1_ASAP7_75t_L g464 ( .A(n_429), .Y(n_464) );
OR2x2_ASAP7_75t_L g465 ( .A(n_426), .B(n_170), .Y(n_465) );
AND2x2_ASAP7_75t_L g466 ( .A(n_426), .B(n_29), .Y(n_466) );
INVx1_ASAP7_75t_L g467 ( .A(n_429), .Y(n_467) );
AND2x2_ASAP7_75t_L g468 ( .A(n_413), .B(n_30), .Y(n_468) );
INVx1_ASAP7_75t_L g469 ( .A(n_429), .Y(n_469) );
INVx2_ASAP7_75t_SL g470 ( .A(n_423), .Y(n_470) );
NOR3xp33_ASAP7_75t_L g471 ( .A(n_401), .B(n_174), .C(n_183), .Y(n_471) );
AO21x2_ASAP7_75t_L g472 ( .A1(n_407), .A2(n_178), .B(n_219), .Y(n_472) );
AND2x2_ASAP7_75t_L g473 ( .A(n_413), .B(n_31), .Y(n_473) );
AO21x2_ASAP7_75t_L g474 ( .A1(n_407), .A2(n_219), .B(n_178), .Y(n_474) );
OAI31xp33_ASAP7_75t_L g475 ( .A1(n_421), .A2(n_258), .A3(n_174), .B(n_193), .Y(n_475) );
AND2x2_ASAP7_75t_L g476 ( .A(n_431), .B(n_36), .Y(n_476) );
NOR3xp33_ASAP7_75t_L g477 ( .A(n_401), .B(n_183), .C(n_193), .Y(n_477) );
OR2x6_ASAP7_75t_SL g478 ( .A(n_421), .B(n_43), .Y(n_478) );
AND2x2_ASAP7_75t_L g479 ( .A(n_423), .B(n_44), .Y(n_479) );
INVx1_ASAP7_75t_L g480 ( .A(n_433), .Y(n_480) );
OR2x6_ASAP7_75t_L g481 ( .A(n_412), .B(n_205), .Y(n_481) );
BUFx3_ASAP7_75t_L g482 ( .A(n_423), .Y(n_482) );
OAI22xp5_ASAP7_75t_L g483 ( .A1(n_424), .A2(n_284), .B1(n_262), .B2(n_259), .Y(n_483) );
NAND2xp5_ASAP7_75t_L g484 ( .A(n_463), .B(n_433), .Y(n_484) );
OR2x2_ASAP7_75t_L g485 ( .A(n_480), .B(n_410), .Y(n_485) );
INVx2_ASAP7_75t_L g486 ( .A(n_439), .Y(n_486) );
INVx2_ASAP7_75t_L g487 ( .A(n_439), .Y(n_487) );
OAI221xp5_ASAP7_75t_L g488 ( .A1(n_438), .A2(n_430), .B1(n_416), .B2(n_422), .C(n_399), .Y(n_488) );
NAND2x1_ASAP7_75t_L g489 ( .A(n_481), .B(n_410), .Y(n_489) );
HB1xp67_ASAP7_75t_L g490 ( .A(n_436), .Y(n_490) );
INVx1_ASAP7_75t_L g491 ( .A(n_447), .Y(n_491) );
INVx1_ASAP7_75t_L g492 ( .A(n_447), .Y(n_492) );
INVx1_ASAP7_75t_L g493 ( .A(n_454), .Y(n_493) );
INVx1_ASAP7_75t_L g494 ( .A(n_454), .Y(n_494) );
INVx2_ASAP7_75t_L g495 ( .A(n_464), .Y(n_495) );
HB1xp67_ASAP7_75t_L g496 ( .A(n_441), .Y(n_496) );
INVx1_ASAP7_75t_L g497 ( .A(n_449), .Y(n_497) );
AND2x2_ASAP7_75t_L g498 ( .A(n_445), .B(n_410), .Y(n_498) );
AND2x2_ASAP7_75t_SL g499 ( .A(n_476), .B(n_416), .Y(n_499) );
NOR3xp33_ASAP7_75t_SL g500 ( .A(n_450), .B(n_427), .C(n_420), .Y(n_500) );
INVx1_ASAP7_75t_L g501 ( .A(n_449), .Y(n_501) );
HB1xp67_ASAP7_75t_L g502 ( .A(n_480), .Y(n_502) );
INVx1_ASAP7_75t_L g503 ( .A(n_464), .Y(n_503) );
AND4x1_ASAP7_75t_L g504 ( .A(n_475), .B(n_432), .C(n_420), .D(n_427), .Y(n_504) );
NOR2xp67_ASAP7_75t_L g505 ( .A(n_450), .B(n_432), .Y(n_505) );
AND2x2_ASAP7_75t_L g506 ( .A(n_445), .B(n_412), .Y(n_506) );
OR2x2_ASAP7_75t_L g507 ( .A(n_437), .B(n_205), .Y(n_507) );
INVx1_ASAP7_75t_L g508 ( .A(n_467), .Y(n_508) );
INVx1_ASAP7_75t_SL g509 ( .A(n_466), .Y(n_509) );
INVx1_ASAP7_75t_L g510 ( .A(n_467), .Y(n_510) );
OR2x2_ASAP7_75t_L g511 ( .A(n_437), .B(n_205), .Y(n_511) );
AOI211xp5_ASAP7_75t_L g512 ( .A1(n_476), .A2(n_193), .B(n_183), .C(n_195), .Y(n_512) );
AND2x2_ASAP7_75t_L g513 ( .A(n_435), .B(n_46), .Y(n_513) );
AND2x2_ASAP7_75t_L g514 ( .A(n_435), .B(n_48), .Y(n_514) );
OR2x2_ASAP7_75t_L g515 ( .A(n_469), .B(n_195), .Y(n_515) );
AND2x2_ASAP7_75t_L g516 ( .A(n_469), .B(n_50), .Y(n_516) );
INVx1_ASAP7_75t_L g517 ( .A(n_446), .Y(n_517) );
NAND2xp5_ASAP7_75t_L g518 ( .A(n_468), .B(n_55), .Y(n_518) );
INVxp67_ASAP7_75t_L g519 ( .A(n_478), .Y(n_519) );
INVx2_ASAP7_75t_L g520 ( .A(n_443), .Y(n_520) );
NAND2xp5_ASAP7_75t_L g521 ( .A(n_468), .B(n_57), .Y(n_521) );
AOI31xp33_ASAP7_75t_L g522 ( .A1(n_473), .A2(n_60), .A3(n_62), .B(n_65), .Y(n_522) );
INVx1_ASAP7_75t_L g523 ( .A(n_443), .Y(n_523) );
INVx1_ASAP7_75t_L g524 ( .A(n_443), .Y(n_524) );
AND2x2_ASAP7_75t_L g525 ( .A(n_482), .B(n_68), .Y(n_525) );
INVx1_ASAP7_75t_SL g526 ( .A(n_466), .Y(n_526) );
OR2x2_ASAP7_75t_L g527 ( .A(n_482), .B(n_442), .Y(n_527) );
NAND2xp5_ASAP7_75t_L g528 ( .A(n_473), .B(n_69), .Y(n_528) );
NAND2xp5_ASAP7_75t_L g529 ( .A(n_470), .B(n_70), .Y(n_529) );
OR2x2_ASAP7_75t_L g530 ( .A(n_482), .B(n_174), .Y(n_530) );
INVx1_ASAP7_75t_L g531 ( .A(n_443), .Y(n_531) );
OR2x2_ASAP7_75t_L g532 ( .A(n_442), .B(n_195), .Y(n_532) );
INVx2_ASAP7_75t_L g533 ( .A(n_472), .Y(n_533) );
INVx2_ASAP7_75t_L g534 ( .A(n_472), .Y(n_534) );
AND2x2_ASAP7_75t_L g535 ( .A(n_442), .B(n_76), .Y(n_535) );
INVx1_ASAP7_75t_L g536 ( .A(n_446), .Y(n_536) );
INVx1_ASAP7_75t_L g537 ( .A(n_451), .Y(n_537) );
AND2x2_ASAP7_75t_L g538 ( .A(n_442), .B(n_244), .Y(n_538) );
AOI221x1_ASAP7_75t_L g539 ( .A1(n_459), .A2(n_244), .B1(n_251), .B2(n_276), .C(n_257), .Y(n_539) );
AND2x2_ASAP7_75t_L g540 ( .A(n_470), .B(n_251), .Y(n_540) );
INVx2_ASAP7_75t_SL g541 ( .A(n_481), .Y(n_541) );
NOR2xp33_ASAP7_75t_L g542 ( .A(n_519), .B(n_434), .Y(n_542) );
AND2x2_ASAP7_75t_L g543 ( .A(n_498), .B(n_444), .Y(n_543) );
INVx1_ASAP7_75t_L g544 ( .A(n_502), .Y(n_544) );
INVx2_ASAP7_75t_L g545 ( .A(n_495), .Y(n_545) );
OR2x2_ASAP7_75t_L g546 ( .A(n_484), .B(n_461), .Y(n_546) );
INVxp67_ASAP7_75t_L g547 ( .A(n_490), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g548 ( .A(n_496), .B(n_478), .Y(n_548) );
INVx1_ASAP7_75t_L g549 ( .A(n_491), .Y(n_549) );
NAND4xp25_ASAP7_75t_L g550 ( .A(n_505), .B(n_456), .C(n_455), .D(n_459), .Y(n_550) );
AND2x2_ASAP7_75t_L g551 ( .A(n_509), .B(n_479), .Y(n_551) );
OR2x2_ASAP7_75t_L g552 ( .A(n_498), .B(n_460), .Y(n_552) );
INVx2_ASAP7_75t_L g553 ( .A(n_495), .Y(n_553) );
NOR2xp33_ASAP7_75t_L g554 ( .A(n_499), .B(n_456), .Y(n_554) );
INVx1_ASAP7_75t_L g555 ( .A(n_492), .Y(n_555) );
INVx1_ASAP7_75t_L g556 ( .A(n_493), .Y(n_556) );
OR2x2_ASAP7_75t_L g557 ( .A(n_527), .B(n_460), .Y(n_557) );
INVx2_ASAP7_75t_SL g558 ( .A(n_527), .Y(n_558) );
NAND2xp5_ASAP7_75t_L g559 ( .A(n_494), .B(n_451), .Y(n_559) );
OAI21xp33_ASAP7_75t_L g560 ( .A1(n_522), .A2(n_455), .B(n_461), .Y(n_560) );
NAND2xp5_ASAP7_75t_L g561 ( .A(n_517), .B(n_479), .Y(n_561) );
NOR2xp33_ASAP7_75t_L g562 ( .A(n_499), .B(n_457), .Y(n_562) );
INVx1_ASAP7_75t_L g563 ( .A(n_501), .Y(n_563) );
AOI211x1_ASAP7_75t_SL g564 ( .A1(n_518), .A2(n_448), .B(n_452), .C(n_462), .Y(n_564) );
INVx3_ASAP7_75t_L g565 ( .A(n_489), .Y(n_565) );
AND2x2_ASAP7_75t_L g566 ( .A(n_526), .B(n_481), .Y(n_566) );
OR2x2_ASAP7_75t_L g567 ( .A(n_485), .B(n_465), .Y(n_567) );
NAND2xp5_ASAP7_75t_L g568 ( .A(n_536), .B(n_444), .Y(n_568) );
AND2x2_ASAP7_75t_L g569 ( .A(n_513), .B(n_481), .Y(n_569) );
AND2x2_ASAP7_75t_L g570 ( .A(n_513), .B(n_514), .Y(n_570) );
NAND2xp5_ASAP7_75t_L g571 ( .A(n_537), .B(n_444), .Y(n_571) );
AOI32xp33_ASAP7_75t_L g572 ( .A1(n_512), .A2(n_477), .A3(n_471), .B1(n_453), .B2(n_440), .Y(n_572) );
INVx1_ASAP7_75t_L g573 ( .A(n_501), .Y(n_573) );
INVx1_ASAP7_75t_L g574 ( .A(n_503), .Y(n_574) );
NOR2x1_ASAP7_75t_L g575 ( .A(n_535), .B(n_481), .Y(n_575) );
AOI21xp5_ASAP7_75t_L g576 ( .A1(n_489), .A2(n_475), .B(n_458), .Y(n_576) );
INVx1_ASAP7_75t_L g577 ( .A(n_503), .Y(n_577) );
OR2x2_ASAP7_75t_L g578 ( .A(n_485), .B(n_465), .Y(n_578) );
AND2x2_ASAP7_75t_L g579 ( .A(n_514), .B(n_474), .Y(n_579) );
INVxp67_ASAP7_75t_L g580 ( .A(n_508), .Y(n_580) );
AND2x2_ASAP7_75t_L g581 ( .A(n_506), .B(n_474), .Y(n_581) );
BUFx2_ASAP7_75t_L g582 ( .A(n_535), .Y(n_582) );
INVx2_ASAP7_75t_L g583 ( .A(n_508), .Y(n_583) );
INVx1_ASAP7_75t_L g584 ( .A(n_497), .Y(n_584) );
NAND3xp33_ASAP7_75t_L g585 ( .A(n_500), .B(n_483), .C(n_257), .Y(n_585) );
INVx2_ASAP7_75t_SL g586 ( .A(n_541), .Y(n_586) );
OAI321xp33_ASAP7_75t_L g587 ( .A1(n_541), .A2(n_458), .A3(n_275), .B1(n_276), .B2(n_264), .C(n_474), .Y(n_587) );
INVxp67_ASAP7_75t_L g588 ( .A(n_523), .Y(n_588) );
NAND2xp5_ASAP7_75t_L g589 ( .A(n_510), .B(n_472), .Y(n_589) );
NAND2xp5_ASAP7_75t_L g590 ( .A(n_506), .B(n_458), .Y(n_590) );
NAND2xp5_ASAP7_75t_L g591 ( .A(n_486), .B(n_264), .Y(n_591) );
INVx1_ASAP7_75t_L g592 ( .A(n_486), .Y(n_592) );
AND2x2_ASAP7_75t_L g593 ( .A(n_543), .B(n_524), .Y(n_593) );
AND2x4_ASAP7_75t_L g594 ( .A(n_575), .B(n_524), .Y(n_594) );
XNOR2xp5_ASAP7_75t_L g595 ( .A(n_570), .B(n_504), .Y(n_595) );
INVx2_ASAP7_75t_L g596 ( .A(n_545), .Y(n_596) );
O2A1O1Ixp5_ASAP7_75t_L g597 ( .A1(n_542), .A2(n_521), .B(n_528), .C(n_525), .Y(n_597) );
INVx1_ASAP7_75t_L g598 ( .A(n_544), .Y(n_598) );
OAI211xp5_ASAP7_75t_L g599 ( .A1(n_560), .A2(n_488), .B(n_525), .C(n_529), .Y(n_599) );
AND2x2_ASAP7_75t_L g600 ( .A(n_543), .B(n_523), .Y(n_600) );
OR2x2_ASAP7_75t_L g601 ( .A(n_558), .B(n_511), .Y(n_601) );
INVx2_ASAP7_75t_L g602 ( .A(n_545), .Y(n_602) );
NAND2xp5_ASAP7_75t_SL g603 ( .A(n_565), .B(n_487), .Y(n_603) );
AND2x2_ASAP7_75t_L g604 ( .A(n_558), .B(n_531), .Y(n_604) );
NAND2xp5_ASAP7_75t_L g605 ( .A(n_547), .B(n_531), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g606 ( .A(n_547), .B(n_487), .Y(n_606) );
AOI21xp33_ASAP7_75t_SL g607 ( .A1(n_548), .A2(n_532), .B(n_516), .Y(n_607) );
NAND2xp5_ASAP7_75t_L g608 ( .A(n_580), .B(n_507), .Y(n_608) );
NAND2x1_ASAP7_75t_L g609 ( .A(n_582), .B(n_516), .Y(n_609) );
INVx1_ASAP7_75t_L g610 ( .A(n_580), .Y(n_610) );
NAND2xp5_ASAP7_75t_L g611 ( .A(n_542), .B(n_511), .Y(n_611) );
NOR2xp33_ASAP7_75t_L g612 ( .A(n_554), .B(n_562), .Y(n_612) );
INVx1_ASAP7_75t_L g613 ( .A(n_549), .Y(n_613) );
INVx1_ASAP7_75t_L g614 ( .A(n_555), .Y(n_614) );
INVxp67_ASAP7_75t_L g615 ( .A(n_586), .Y(n_615) );
NOR2xp33_ASAP7_75t_L g616 ( .A(n_554), .B(n_532), .Y(n_616) );
NAND2xp5_ASAP7_75t_L g617 ( .A(n_556), .B(n_507), .Y(n_617) );
AND2x4_ASAP7_75t_L g618 ( .A(n_565), .B(n_586), .Y(n_618) );
NOR2x1p5_ASAP7_75t_L g619 ( .A(n_550), .B(n_530), .Y(n_619) );
INVxp67_ASAP7_75t_L g620 ( .A(n_551), .Y(n_620) );
OR2x2_ASAP7_75t_L g621 ( .A(n_567), .B(n_520), .Y(n_621) );
INVx2_ASAP7_75t_L g622 ( .A(n_553), .Y(n_622) );
INVx1_ASAP7_75t_L g623 ( .A(n_574), .Y(n_623) );
NAND2xp5_ASAP7_75t_SL g624 ( .A(n_565), .B(n_520), .Y(n_624) );
OR2x2_ASAP7_75t_L g625 ( .A(n_578), .B(n_534), .Y(n_625) );
NOR2x1_ASAP7_75t_L g626 ( .A(n_576), .B(n_515), .Y(n_626) );
INVx1_ASAP7_75t_L g627 ( .A(n_577), .Y(n_627) );
INVx1_ASAP7_75t_L g628 ( .A(n_584), .Y(n_628) );
INVx1_ASAP7_75t_L g629 ( .A(n_583), .Y(n_629) );
INVx1_ASAP7_75t_L g630 ( .A(n_583), .Y(n_630) );
AOI221xp5_ASAP7_75t_L g631 ( .A1(n_562), .A2(n_540), .B1(n_538), .B2(n_534), .C(n_533), .Y(n_631) );
CKINVDCx14_ASAP7_75t_R g632 ( .A(n_552), .Y(n_632) );
INVx1_ASAP7_75t_L g633 ( .A(n_563), .Y(n_633) );
INVx2_ASAP7_75t_L g634 ( .A(n_553), .Y(n_634) );
NOR3xp33_ASAP7_75t_L g635 ( .A(n_585), .B(n_530), .C(n_538), .Y(n_635) );
AOI21xp33_ASAP7_75t_SL g636 ( .A1(n_572), .A2(n_515), .B(n_533), .Y(n_636) );
AOI221xp5_ASAP7_75t_L g637 ( .A1(n_588), .A2(n_540), .B1(n_275), .B2(n_539), .C(n_270), .Y(n_637) );
AOI221xp5_ASAP7_75t_L g638 ( .A1(n_561), .A2(n_539), .B1(n_270), .B2(n_259), .C(n_262), .Y(n_638) );
NOR2x1_ASAP7_75t_L g639 ( .A(n_573), .B(n_255), .Y(n_639) );
NOR3xp33_ASAP7_75t_L g640 ( .A(n_587), .B(n_258), .C(n_284), .Y(n_640) );
INVx1_ASAP7_75t_L g641 ( .A(n_592), .Y(n_641) );
INVx1_ASAP7_75t_L g642 ( .A(n_588), .Y(n_642) );
XNOR2x1_ASAP7_75t_L g643 ( .A(n_546), .B(n_270), .Y(n_643) );
OAI21xp33_ASAP7_75t_SL g644 ( .A1(n_569), .A2(n_284), .B(n_270), .Y(n_644) );
NAND2xp5_ASAP7_75t_L g645 ( .A(n_568), .B(n_270), .Y(n_645) );
INVx1_ASAP7_75t_L g646 ( .A(n_589), .Y(n_646) );
INVx1_ASAP7_75t_L g647 ( .A(n_557), .Y(n_647) );
OAI22xp5_ASAP7_75t_L g648 ( .A1(n_559), .A2(n_284), .B1(n_590), .B2(n_579), .Y(n_648) );
OAI21xp33_ASAP7_75t_SL g649 ( .A1(n_566), .A2(n_284), .B(n_581), .Y(n_649) );
INVx2_ASAP7_75t_SL g650 ( .A(n_591), .Y(n_650) );
INVx2_ASAP7_75t_SL g651 ( .A(n_601), .Y(n_651) );
OAI211xp5_ASAP7_75t_L g652 ( .A1(n_636), .A2(n_599), .B(n_611), .C(n_649), .Y(n_652) );
AO22x1_ASAP7_75t_L g653 ( .A1(n_635), .A2(n_626), .B1(n_618), .B2(n_612), .Y(n_653) );
NAND2x1_ASAP7_75t_SL g654 ( .A(n_618), .B(n_594), .Y(n_654) );
BUFx2_ASAP7_75t_L g655 ( .A(n_632), .Y(n_655) );
NAND4xp25_ASAP7_75t_L g656 ( .A(n_597), .B(n_612), .C(n_564), .D(n_631), .Y(n_656) );
AOI22xp5_ASAP7_75t_L g657 ( .A1(n_619), .A2(n_616), .B1(n_595), .B2(n_643), .Y(n_657) );
AOI31xp33_ASAP7_75t_L g658 ( .A1(n_644), .A2(n_607), .A3(n_615), .B(n_618), .Y(n_658) );
AOI211x1_ASAP7_75t_SL g659 ( .A1(n_648), .A2(n_605), .B(n_606), .C(n_603), .Y(n_659) );
OAI22xp33_ASAP7_75t_L g660 ( .A1(n_609), .A2(n_620), .B1(n_648), .B2(n_647), .Y(n_660) );
AOI21xp33_ASAP7_75t_L g661 ( .A1(n_616), .A2(n_598), .B(n_646), .Y(n_661) );
OAI31xp33_ASAP7_75t_L g662 ( .A1(n_594), .A2(n_610), .A3(n_642), .B(n_604), .Y(n_662) );
OA22x2_ASAP7_75t_L g663 ( .A1(n_594), .A2(n_614), .B1(n_613), .B2(n_603), .Y(n_663) );
OAI211xp5_ASAP7_75t_L g664 ( .A1(n_657), .A2(n_624), .B(n_638), .C(n_608), .Y(n_664) );
CKINVDCx20_ASAP7_75t_R g665 ( .A(n_655), .Y(n_665) );
OAI332xp33_ASAP7_75t_L g666 ( .A1(n_660), .A2(n_628), .A3(n_650), .B1(n_621), .B2(n_625), .B3(n_627), .C1(n_623), .C2(n_633), .Y(n_666) );
OA22x2_ASAP7_75t_L g667 ( .A1(n_657), .A2(n_593), .B1(n_600), .B2(n_624), .Y(n_667) );
OAI211xp5_ASAP7_75t_SL g668 ( .A1(n_659), .A2(n_638), .B(n_637), .C(n_639), .Y(n_668) );
OAI322xp33_ASAP7_75t_L g669 ( .A1(n_663), .A2(n_617), .A3(n_641), .B1(n_630), .B2(n_629), .C1(n_571), .C2(n_602), .Y(n_669) );
AOI21xp5_ASAP7_75t_L g670 ( .A1(n_658), .A2(n_622), .B(n_596), .Y(n_670) );
XNOR2xp5_ASAP7_75t_L g671 ( .A(n_653), .B(n_593), .Y(n_671) );
NAND2xp5_ASAP7_75t_L g672 ( .A(n_664), .B(n_656), .Y(n_672) );
INVx1_ASAP7_75t_SL g673 ( .A(n_665), .Y(n_673) );
OAI21xp33_ASAP7_75t_SL g674 ( .A1(n_667), .A2(n_654), .B(n_662), .Y(n_674) );
NAND4xp75_ASAP7_75t_L g675 ( .A(n_670), .B(n_661), .C(n_652), .D(n_651), .Y(n_675) );
NOR3xp33_ASAP7_75t_L g676 ( .A(n_675), .B(n_666), .C(n_668), .Y(n_676) );
OAI22x1_ASAP7_75t_L g677 ( .A1(n_672), .A2(n_671), .B1(n_669), .B2(n_602), .Y(n_677) );
HB1xp67_ASAP7_75t_L g678 ( .A(n_673), .Y(n_678) );
NOR3xp33_ASAP7_75t_L g679 ( .A(n_678), .B(n_676), .C(n_674), .Y(n_679) );
BUFx2_ASAP7_75t_L g680 ( .A(n_677), .Y(n_680) );
NAND2xp5_ASAP7_75t_L g681 ( .A(n_679), .B(n_600), .Y(n_681) );
INVx1_ASAP7_75t_SL g682 ( .A(n_680), .Y(n_682) );
AOI21xp5_ASAP7_75t_L g683 ( .A1(n_682), .A2(n_645), .B(n_640), .Y(n_683) );
AO21x2_ASAP7_75t_L g684 ( .A1(n_683), .A2(n_681), .B(n_645), .Y(n_684) );
AOI221xp5_ASAP7_75t_L g685 ( .A1(n_684), .A2(n_596), .B1(n_622), .B2(n_634), .C(n_679), .Y(n_685) );
endmodule