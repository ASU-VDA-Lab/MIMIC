module fake_aes_9009_n_15 (n_1, n_2, n_4, n_3, n_0, n_15);
input n_1;
input n_2;
input n_4;
input n_3;
input n_0;
output n_15;
wire n_11;
wire n_13;
wire n_12;
wire n_6;
wire n_9;
wire n_5;
wire n_14;
wire n_8;
wire n_10;
wire n_7;
NAND2xp5_ASAP7_75t_L g5 ( .A(n_1), .B(n_0), .Y(n_5) );
INVx1_ASAP7_75t_L g6 ( .A(n_2), .Y(n_6) );
NAND2xp5_ASAP7_75t_L g7 ( .A(n_0), .B(n_4), .Y(n_7) );
BUFx3_ASAP7_75t_L g8 ( .A(n_3), .Y(n_8) );
OA21x2_ASAP7_75t_L g9 ( .A1(n_6), .A2(n_0), .B(n_1), .Y(n_9) );
BUFx2_ASAP7_75t_L g10 ( .A(n_8), .Y(n_10) );
BUFx3_ASAP7_75t_L g11 ( .A(n_8), .Y(n_11) );
OAI211xp5_ASAP7_75t_L g12 ( .A1(n_10), .A2(n_5), .B(n_7), .C(n_6), .Y(n_12) );
INVxp67_ASAP7_75t_L g13 ( .A(n_12), .Y(n_13) );
AND2x2_ASAP7_75t_L g14 ( .A(n_13), .B(n_9), .Y(n_14) );
NAND2xp5_ASAP7_75t_L g15 ( .A(n_14), .B(n_11), .Y(n_15) );
endmodule