module real_jpeg_6715_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_271;
wire n_47;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_425;
wire n_50;
wire n_409;
wire n_186;
wire n_137;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_366;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_417;
wire n_428;
wire n_216;
wire n_128;
wire n_202;
wire n_367;
wire n_127;
wire n_365;
wire n_356;
wire n_423;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_83;
wire n_288;
wire n_78;
wire n_221;
wire n_393;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_200;
wire n_432;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_338;
wire n_175;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_372;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_286;
wire n_215;
wire n_166;
wire n_176;
wire n_323;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_18;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_299;
wire n_243;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

INVx8_ASAP7_75t_L g54 ( 
.A(n_0),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_1),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_1),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_2),
.A2(n_107),
.B1(n_109),
.B2(n_110),
.Y(n_106)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_2),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_SL g170 ( 
.A1(n_2),
.A2(n_109),
.B1(n_171),
.B2(n_172),
.Y(n_170)
);

OAI22xp33_ASAP7_75t_L g225 ( 
.A1(n_2),
.A2(n_109),
.B1(n_226),
.B2(n_227),
.Y(n_225)
);

AOI22xp33_ASAP7_75t_L g376 ( 
.A1(n_2),
.A2(n_109),
.B1(n_179),
.B2(n_377),
.Y(n_376)
);

INVx6_ASAP7_75t_L g93 ( 
.A(n_3),
.Y(n_93)
);

INVx8_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_4),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g164 ( 
.A(n_4),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g185 ( 
.A(n_4),
.Y(n_185)
);

BUFx6f_ASAP7_75t_L g264 ( 
.A(n_4),
.Y(n_264)
);

INVx2_ASAP7_75t_L g402 ( 
.A(n_4),
.Y(n_402)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_5),
.A2(n_50),
.B1(n_81),
.B2(n_82),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_5),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_L g177 ( 
.A1(n_5),
.A2(n_81),
.B1(n_178),
.B2(n_180),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_5),
.A2(n_81),
.B1(n_206),
.B2(n_207),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_6),
.A2(n_127),
.B1(n_138),
.B2(n_189),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_6),
.Y(n_189)
);

AOI22xp33_ASAP7_75t_L g314 ( 
.A1(n_6),
.A2(n_189),
.B1(n_315),
.B2(n_316),
.Y(n_314)
);

OAI22xp5_ASAP7_75t_L g337 ( 
.A1(n_6),
.A2(n_189),
.B1(n_338),
.B2(n_341),
.Y(n_337)
);

AOI22xp33_ASAP7_75t_SL g395 ( 
.A1(n_6),
.A2(n_110),
.B1(n_189),
.B2(n_396),
.Y(n_395)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_7),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_7),
.Y(n_130)
);

INVx8_ASAP7_75t_L g96 ( 
.A(n_8),
.Y(n_96)
);

OAI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_9),
.A2(n_49),
.B1(n_55),
.B2(n_56),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_9),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_9),
.A2(n_55),
.B1(n_115),
.B2(n_117),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g260 ( 
.A1(n_9),
.A2(n_28),
.B1(n_55),
.B2(n_261),
.Y(n_260)
);

INVx6_ASAP7_75t_L g127 ( 
.A(n_10),
.Y(n_127)
);

BUFx5_ASAP7_75t_L g128 ( 
.A(n_10),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g138 ( 
.A(n_10),
.Y(n_138)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_10),
.Y(n_142)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_10),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g226 ( 
.A(n_10),
.Y(n_226)
);

OAI22xp33_ASAP7_75t_SL g31 ( 
.A1(n_11),
.A2(n_28),
.B1(n_32),
.B2(n_35),
.Y(n_31)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_11),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_11),
.A2(n_35),
.B1(n_155),
.B2(n_158),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_12),
.A2(n_137),
.B1(n_139),
.B2(n_140),
.Y(n_136)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_12),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_L g268 ( 
.A1(n_12),
.A2(n_139),
.B1(n_269),
.B2(n_271),
.Y(n_268)
);

OAI22xp33_ASAP7_75t_SL g299 ( 
.A1(n_12),
.A2(n_41),
.B1(n_139),
.B2(n_300),
.Y(n_299)
);

AOI22xp33_ASAP7_75t_SL g364 ( 
.A1(n_12),
.A2(n_139),
.B1(n_365),
.B2(n_367),
.Y(n_364)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_13),
.Y(n_256)
);

AOI22xp33_ASAP7_75t_SL g284 ( 
.A1(n_13),
.A2(n_172),
.B1(n_256),
.B2(n_285),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_13),
.B(n_294),
.C(n_295),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_SL g320 ( 
.A(n_13),
.B(n_101),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_13),
.B(n_332),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_13),
.B(n_84),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_L g372 ( 
.A(n_13),
.B(n_195),
.Y(n_372)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_14),
.Y(n_68)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_14),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g294 ( 
.A(n_14),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_15),
.A2(n_145),
.B1(n_146),
.B2(n_147),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_15),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_15),
.A2(n_115),
.B1(n_145),
.B2(n_194),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_15),
.A2(n_145),
.B1(n_156),
.B2(n_288),
.Y(n_287)
);

AOI22xp33_ASAP7_75t_L g306 ( 
.A1(n_15),
.A2(n_145),
.B1(n_307),
.B2(n_308),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_L g39 ( 
.A1(n_16),
.A2(n_40),
.B1(n_41),
.B2(n_44),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_16),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_SL g214 ( 
.A1(n_16),
.A2(n_40),
.B1(n_215),
.B2(n_216),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_230),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_229),
.Y(n_18)
);

OR2x2_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_197),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_20),
.B(n_197),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_151),
.C(n_166),
.Y(n_20)
);

FAx1_ASAP7_75t_SL g274 ( 
.A(n_21),
.B(n_151),
.CI(n_166),
.CON(n_274),
.SN(n_274)
);

XNOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_85),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_22),
.B(n_86),
.C(n_120),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_47),
.Y(n_22)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_23),
.B(n_47),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_31),
.B1(n_36),
.B2(n_39),
.Y(n_23)
);

OAI21xp5_ASAP7_75t_SL g161 ( 
.A1(n_24),
.A2(n_39),
.B(n_162),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_24),
.A2(n_259),
.B1(n_262),
.B2(n_265),
.Y(n_258)
);

AOI21xp5_ASAP7_75t_L g298 ( 
.A1(n_24),
.A2(n_299),
.B(n_303),
.Y(n_298)
);

AOI21xp5_ASAP7_75t_L g334 ( 
.A1(n_24),
.A2(n_256),
.B(n_303),
.Y(n_334)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_25),
.A2(n_177),
.B1(n_183),
.B2(n_184),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g346 ( 
.A(n_25),
.B(n_306),
.Y(n_346)
);

OAI22xp5_ASAP7_75t_SL g350 ( 
.A1(n_25),
.A2(n_351),
.B1(n_352),
.B2(n_353),
.Y(n_350)
);

OAI22xp5_ASAP7_75t_SL g401 ( 
.A1(n_25),
.A2(n_260),
.B1(n_376),
.B2(n_402),
.Y(n_401)
);

OR2x2_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_28),
.Y(n_25)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVx2_ASAP7_75t_L g305 ( 
.A(n_27),
.Y(n_305)
);

BUFx6f_ASAP7_75t_L g333 ( 
.A(n_27),
.Y(n_333)
);

INVx2_ASAP7_75t_L g345 ( 
.A(n_27),
.Y(n_345)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

BUFx2_ASAP7_75t_L g261 ( 
.A(n_29),
.Y(n_261)
);

BUFx8_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g46 ( 
.A(n_30),
.Y(n_46)
);

INVx2_ASAP7_75t_L g330 ( 
.A(n_30),
.Y(n_330)
);

BUFx3_ASAP7_75t_L g340 ( 
.A(n_30),
.Y(n_340)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_31),
.Y(n_183)
);

INVx4_ASAP7_75t_L g307 ( 
.A(n_32),
.Y(n_307)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

HB1xp67_ASAP7_75t_L g296 ( 
.A(n_33),
.Y(n_296)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_34),
.Y(n_77)
);

BUFx3_ASAP7_75t_L g182 ( 
.A(n_34),
.Y(n_182)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_43),
.Y(n_78)
);

BUFx5_ASAP7_75t_L g342 ( 
.A(n_43),
.Y(n_342)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

BUFx2_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_L g47 ( 
.A1(n_48),
.A2(n_61),
.B1(n_80),
.B2(n_84),
.Y(n_47)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_48),
.Y(n_175)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx4_ASAP7_75t_SL g51 ( 
.A(n_52),
.Y(n_51)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g292 ( 
.A(n_53),
.Y(n_292)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx11_ASAP7_75t_L g60 ( 
.A(n_54),
.Y(n_60)
);

BUFx5_ASAP7_75t_L g83 ( 
.A(n_54),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g289 ( 
.A(n_54),
.Y(n_289)
);

INVx2_ASAP7_75t_L g317 ( 
.A(n_54),
.Y(n_317)
);

INVx3_ASAP7_75t_L g383 ( 
.A(n_54),
.Y(n_383)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_59),
.Y(n_285)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_60),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_60),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g157 ( 
.A(n_60),
.Y(n_157)
);

INVx5_ASAP7_75t_L g160 ( 
.A(n_60),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_61),
.A2(n_80),
.B1(n_84),
.B2(n_154),
.Y(n_153)
);

INVx2_ASAP7_75t_SL g169 ( 
.A(n_61),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_61),
.A2(n_84),
.B1(n_154),
.B2(n_213),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_61),
.B(n_287),
.Y(n_318)
);

AND2x2_ASAP7_75t_L g61 ( 
.A(n_62),
.B(n_73),
.Y(n_61)
);

OAI22xp33_ASAP7_75t_L g62 ( 
.A1(n_63),
.A2(n_66),
.B1(n_69),
.B2(n_72),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx5_ASAP7_75t_L g216 ( 
.A(n_65),
.Y(n_216)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_68),
.Y(n_74)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_71),
.Y(n_79)
);

AO22x2_ASAP7_75t_L g101 ( 
.A1(n_72),
.A2(n_83),
.B1(n_102),
.B2(n_104),
.Y(n_101)
);

INVx11_ASAP7_75t_L g315 ( 
.A(n_72),
.Y(n_315)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_73),
.Y(n_84)
);

OAI21xp5_ASAP7_75t_SL g313 ( 
.A1(n_73),
.A2(n_314),
.B(n_318),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_74),
.A2(n_75),
.B1(n_78),
.B2(n_79),
.Y(n_73)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g179 ( 
.A(n_76),
.Y(n_179)
);

INVx5_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx2_ASAP7_75t_L g310 ( 
.A(n_77),
.Y(n_310)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_82),
.Y(n_171)
);

INVx5_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_84),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g286 ( 
.A(n_84),
.B(n_287),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g85 ( 
.A(n_86),
.B(n_120),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_87),
.A2(n_106),
.B1(n_113),
.B2(n_114),
.Y(n_86)
);

INVx3_ASAP7_75t_SL g191 ( 
.A(n_87),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g423 ( 
.A1(n_87),
.A2(n_113),
.B1(n_268),
.B2(n_395),
.Y(n_423)
);

OR2x2_ASAP7_75t_L g87 ( 
.A(n_88),
.B(n_101),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_L g88 ( 
.A1(n_89),
.A2(n_94),
.B1(n_97),
.B2(n_98),
.Y(n_88)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_91),
.Y(n_97)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g380 ( 
.A(n_92),
.Y(n_380)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

BUFx3_ASAP7_75t_L g103 ( 
.A(n_93),
.Y(n_103)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_93),
.Y(n_105)
);

INVx3_ASAP7_75t_L g195 ( 
.A(n_94),
.Y(n_195)
);

INVx5_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_95),
.Y(n_210)
);

BUFx5_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_96),
.Y(n_100)
);

INVx6_ASAP7_75t_L g108 ( 
.A(n_96),
.Y(n_108)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_96),
.Y(n_116)
);

INVx3_ASAP7_75t_L g134 ( 
.A(n_96),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g246 ( 
.A(n_96),
.Y(n_246)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

BUFx2_ASAP7_75t_L g206 ( 
.A(n_99),
.Y(n_206)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_100),
.Y(n_270)
);

INVx3_ASAP7_75t_L g397 ( 
.A(n_100),
.Y(n_397)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_101),
.Y(n_113)
);

AOI22x1_ASAP7_75t_L g190 ( 
.A1(n_101),
.A2(n_191),
.B1(n_192),
.B2(n_196),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_101),
.A2(n_191),
.B1(n_204),
.B2(n_205),
.Y(n_203)
);

INVx6_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx4_ASAP7_75t_L g384 ( 
.A(n_104),
.Y(n_384)
);

INVx6_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_106),
.Y(n_196)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_108),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_108),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_108),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g254 ( 
.A(n_108),
.Y(n_254)
);

BUFx6f_ASAP7_75t_L g272 ( 
.A(n_108),
.Y(n_272)
);

AOI32xp33_ASAP7_75t_L g378 ( 
.A1(n_110),
.A2(n_289),
.A3(n_372),
.B1(n_379),
.B2(n_381),
.Y(n_378)
);

INVx6_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVx6_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_113),
.B(n_193),
.Y(n_273)
);

OAI21xp5_ASAP7_75t_SL g394 ( 
.A1(n_113),
.A2(n_395),
.B(n_398),
.Y(n_394)
);

INVxp67_ASAP7_75t_L g204 ( 
.A(n_114),
.Y(n_204)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

OAI21xp33_ASAP7_75t_SL g370 ( 
.A1(n_117),
.A2(n_256),
.B(n_371),
.Y(n_370)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_SL g120 ( 
.A1(n_121),
.A2(n_136),
.B(n_143),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_121),
.A2(n_131),
.B1(n_136),
.B2(n_188),
.Y(n_187)
);

INVx1_ASAP7_75t_SL g121 ( 
.A(n_122),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_122),
.B(n_144),
.Y(n_228)
);

AOI21xp5_ASAP7_75t_L g416 ( 
.A1(n_122),
.A2(n_417),
.B(n_421),
.Y(n_416)
);

AND2x2_ASAP7_75t_L g122 ( 
.A(n_123),
.B(n_131),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_124),
.A2(n_127),
.B1(n_128),
.B2(n_129),
.Y(n_123)
);

INVx6_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVx5_ASAP7_75t_L g250 ( 
.A(n_126),
.Y(n_250)
);

INVx8_ASAP7_75t_L g146 ( 
.A(n_127),
.Y(n_146)
);

INVx3_ASAP7_75t_L g247 ( 
.A(n_128),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_128),
.B(n_256),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_129),
.A2(n_132),
.B1(n_133),
.B2(n_135),
.Y(n_131)
);

INVx4_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_130),
.Y(n_132)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_131),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g400 ( 
.A(n_131),
.B(n_256),
.Y(n_400)
);

INVx4_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

INVx4_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

INVx2_ASAP7_75t_L g420 ( 
.A(n_142),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_143),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_150),
.Y(n_143)
);

INVx5_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

INVx3_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_150),
.B(n_225),
.Y(n_224)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_150),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_152),
.A2(n_153),
.B1(n_161),
.B2(n_165),
.Y(n_151)
);

INVxp67_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_153),
.B(n_161),
.Y(n_220)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

INVx4_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_157),
.Y(n_173)
);

INVx3_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

INVx4_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

BUFx2_ASAP7_75t_L g215 ( 
.A(n_160),
.Y(n_215)
);

INVx5_ASAP7_75t_L g366 ( 
.A(n_160),
.Y(n_366)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_161),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_161),
.A2(n_165),
.B1(n_222),
.B2(n_223),
.Y(n_221)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_167),
.B(n_186),
.C(n_190),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_L g235 ( 
.A(n_167),
.B(n_236),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_168),
.B(n_176),
.Y(n_167)
);

XOR2xp5_ASAP7_75t_L g436 ( 
.A(n_168),
.B(n_176),
.Y(n_436)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_169),
.A2(n_170),
.B1(n_174),
.B2(n_175),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_SL g283 ( 
.A1(n_169),
.A2(n_284),
.B(n_286),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_SL g363 ( 
.A1(n_169),
.A2(n_174),
.B1(n_314),
.B2(n_364),
.Y(n_363)
);

OAI21xp5_ASAP7_75t_SL g391 ( 
.A1(n_169),
.A2(n_286),
.B(n_364),
.Y(n_391)
);

OAI21xp5_ASAP7_75t_SL g424 ( 
.A1(n_170),
.A2(n_174),
.B(n_318),
.Y(n_424)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

INVxp67_ASAP7_75t_L g265 ( 
.A(n_177),
.Y(n_265)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

BUFx3_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

BUFx6f_ASAP7_75t_L g302 ( 
.A(n_182),
.Y(n_302)
);

INVx4_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_186),
.A2(n_187),
.B1(n_190),
.B2(n_237),
.Y(n_236)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_L g241 ( 
.A1(n_188),
.A2(n_228),
.B(n_242),
.Y(n_241)
);

INVx1_ASAP7_75t_SL g237 ( 
.A(n_190),
.Y(n_237)
);

AOI21xp5_ASAP7_75t_L g266 ( 
.A1(n_191),
.A2(n_267),
.B(n_273),
.Y(n_266)
);

AOI21xp5_ASAP7_75t_L g369 ( 
.A1(n_191),
.A2(n_273),
.B(n_370),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_191),
.B(n_192),
.Y(n_398)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

INVx4_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_199),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_200),
.A2(n_201),
.B1(n_218),
.B2(n_219),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

AOI21xp5_ASAP7_75t_L g201 ( 
.A1(n_202),
.A2(n_211),
.B(n_217),
.Y(n_201)
);

INVxp67_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

AND2x2_ASAP7_75t_L g217 ( 
.A(n_203),
.B(n_212),
.Y(n_217)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

INVx3_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

INVxp67_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_220),
.B(n_221),
.Y(n_219)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_224),
.B(n_228),
.Y(n_223)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_226),
.Y(n_227)
);

OAI21xp5_ASAP7_75t_L g230 ( 
.A1(n_231),
.A2(n_275),
.B(n_449),
.Y(n_230)
);

INVxp67_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_233),
.B(n_274),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g450 ( 
.A(n_233),
.B(n_274),
.Y(n_450)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_234),
.B(n_238),
.C(n_239),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_SL g439 ( 
.A1(n_234),
.A2(n_235),
.B1(n_238),
.B2(n_440),
.Y(n_439)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_238),
.Y(n_440)
);

XNOR2xp5_ASAP7_75t_L g438 ( 
.A(n_239),
.B(n_439),
.Y(n_438)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_240),
.B(n_243),
.C(n_266),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g433 ( 
.A1(n_240),
.A2(n_241),
.B1(n_266),
.B2(n_434),
.Y(n_433)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g432 ( 
.A(n_243),
.B(n_433),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_244),
.B(n_257),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_L g409 ( 
.A1(n_244),
.A2(n_257),
.B1(n_258),
.B2(n_410),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_244),
.Y(n_410)
);

OAI32xp33_ASAP7_75t_L g244 ( 
.A1(n_245),
.A2(n_247),
.A3(n_248),
.B1(n_251),
.B2(n_255),
.Y(n_244)
);

INVx4_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_249),
.B(n_252),
.Y(n_251)
);

INVx6_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

BUFx6f_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

OAI21xp33_ASAP7_75t_SL g417 ( 
.A1(n_255),
.A2(n_256),
.B(n_418),
.Y(n_417)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

INVxp67_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

INVx3_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_266),
.Y(n_434)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

INVx3_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

BUFx12f_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

BUFx24_ASAP7_75t_SL g451 ( 
.A(n_274),
.Y(n_451)
);

AOI21xp5_ASAP7_75t_L g275 ( 
.A1(n_276),
.A2(n_427),
.B(n_446),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

AOI21xp5_ASAP7_75t_SL g277 ( 
.A1(n_278),
.A2(n_405),
.B(n_426),
.Y(n_277)
);

AO21x1_ASAP7_75t_SL g278 ( 
.A1(n_279),
.A2(n_386),
.B(n_404),
.Y(n_278)
);

OAI21xp5_ASAP7_75t_SL g279 ( 
.A1(n_280),
.A2(n_358),
.B(n_385),
.Y(n_279)
);

AOI21xp5_ASAP7_75t_L g280 ( 
.A1(n_281),
.A2(n_321),
.B(n_357),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_282),
.B(n_297),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g357 ( 
.A(n_282),
.B(n_297),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_SL g282 ( 
.A(n_283),
.B(n_290),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_SL g354 ( 
.A1(n_283),
.A2(n_290),
.B1(n_291),
.B2(n_355),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_283),
.Y(n_355)
);

INVx5_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_292),
.B(n_293),
.Y(n_291)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_298),
.B(n_311),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g359 ( 
.A(n_298),
.B(n_312),
.C(n_320),
.Y(n_359)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_299),
.Y(n_352)
);

INVx6_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

INVx4_ASAP7_75t_L g301 ( 
.A(n_302),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_304),
.B(n_306),
.Y(n_303)
);

INVx4_ASAP7_75t_L g304 ( 
.A(n_305),
.Y(n_304)
);

INVx2_ASAP7_75t_L g377 ( 
.A(n_308),
.Y(n_377)
);

INVx4_ASAP7_75t_SL g308 ( 
.A(n_309),
.Y(n_308)
);

INVx4_ASAP7_75t_L g309 ( 
.A(n_310),
.Y(n_309)
);

AOI22xp5_ASAP7_75t_SL g311 ( 
.A1(n_312),
.A2(n_313),
.B1(n_319),
.B2(n_320),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_313),
.Y(n_312)
);

INVx2_ASAP7_75t_L g367 ( 
.A(n_315),
.Y(n_367)
);

BUFx3_ASAP7_75t_L g316 ( 
.A(n_317),
.Y(n_316)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

OAI21xp5_ASAP7_75t_L g321 ( 
.A1(n_322),
.A2(n_349),
.B(n_356),
.Y(n_321)
);

AOI21xp5_ASAP7_75t_L g322 ( 
.A1(n_323),
.A2(n_335),
.B(n_348),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_324),
.B(n_334),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_325),
.B(n_331),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_326),
.Y(n_325)
);

INVx1_ASAP7_75t_SL g326 ( 
.A(n_327),
.Y(n_326)
);

INVx2_ASAP7_75t_L g327 ( 
.A(n_328),
.Y(n_327)
);

INVx2_ASAP7_75t_L g328 ( 
.A(n_329),
.Y(n_328)
);

INVx2_ASAP7_75t_L g329 ( 
.A(n_330),
.Y(n_329)
);

INVx2_ASAP7_75t_L g353 ( 
.A(n_332),
.Y(n_353)
);

INVx8_ASAP7_75t_L g332 ( 
.A(n_333),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_SL g335 ( 
.A(n_336),
.B(n_347),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g348 ( 
.A(n_336),
.B(n_347),
.Y(n_348)
);

AOI21xp5_ASAP7_75t_L g336 ( 
.A1(n_337),
.A2(n_343),
.B(n_346),
.Y(n_336)
);

INVxp67_ASAP7_75t_L g351 ( 
.A(n_337),
.Y(n_351)
);

INVx2_ASAP7_75t_L g338 ( 
.A(n_339),
.Y(n_338)
);

INVx5_ASAP7_75t_L g339 ( 
.A(n_340),
.Y(n_339)
);

INVx5_ASAP7_75t_L g341 ( 
.A(n_342),
.Y(n_341)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_344),
.Y(n_343)
);

INVx3_ASAP7_75t_L g344 ( 
.A(n_345),
.Y(n_344)
);

AOI21xp5_ASAP7_75t_L g374 ( 
.A1(n_345),
.A2(n_346),
.B(n_375),
.Y(n_374)
);

NOR2xp33_ASAP7_75t_L g349 ( 
.A(n_350),
.B(n_354),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_350),
.B(n_354),
.Y(n_356)
);

NOR2xp33_ASAP7_75t_L g358 ( 
.A(n_359),
.B(n_360),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_359),
.B(n_360),
.Y(n_385)
);

XNOR2xp5_ASAP7_75t_L g360 ( 
.A(n_361),
.B(n_373),
.Y(n_360)
);

AOI22xp5_ASAP7_75t_L g361 ( 
.A1(n_362),
.A2(n_363),
.B1(n_368),
.B2(n_369),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_363),
.Y(n_362)
);

MAJIxp5_ASAP7_75t_L g387 ( 
.A(n_363),
.B(n_368),
.C(n_373),
.Y(n_387)
);

INVx2_ASAP7_75t_L g365 ( 
.A(n_366),
.Y(n_365)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_369),
.Y(n_368)
);

INVxp33_ASAP7_75t_L g371 ( 
.A(n_372),
.Y(n_371)
);

XOR2xp5_ASAP7_75t_L g373 ( 
.A(n_374),
.B(n_378),
.Y(n_373)
);

NOR2xp33_ASAP7_75t_L g392 ( 
.A(n_374),
.B(n_378),
.Y(n_392)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_376),
.Y(n_375)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_380),
.Y(n_379)
);

NAND2xp33_ASAP7_75t_SL g381 ( 
.A(n_382),
.B(n_384),
.Y(n_381)
);

BUFx6f_ASAP7_75t_L g382 ( 
.A(n_383),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_387),
.B(n_388),
.Y(n_386)
);

NOR2xp33_ASAP7_75t_SL g404 ( 
.A(n_387),
.B(n_388),
.Y(n_404)
);

AOI22xp5_ASAP7_75t_L g388 ( 
.A1(n_389),
.A2(n_390),
.B1(n_393),
.B2(n_403),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_390),
.Y(n_389)
);

XNOR2xp5_ASAP7_75t_SL g390 ( 
.A(n_391),
.B(n_392),
.Y(n_390)
);

MAJIxp5_ASAP7_75t_L g406 ( 
.A(n_391),
.B(n_392),
.C(n_403),
.Y(n_406)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_393),
.Y(n_403)
);

XNOR2xp5_ASAP7_75t_SL g393 ( 
.A(n_394),
.B(n_399),
.Y(n_393)
);

MAJIxp5_ASAP7_75t_L g411 ( 
.A(n_394),
.B(n_400),
.C(n_401),
.Y(n_411)
);

INVx2_ASAP7_75t_L g396 ( 
.A(n_397),
.Y(n_396)
);

XOR2xp5_ASAP7_75t_L g399 ( 
.A(n_400),
.B(n_401),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_406),
.B(n_407),
.Y(n_405)
);

NOR2xp33_ASAP7_75t_SL g426 ( 
.A(n_406),
.B(n_407),
.Y(n_426)
);

XNOR2xp5_ASAP7_75t_L g407 ( 
.A(n_408),
.B(n_414),
.Y(n_407)
);

AOI22xp5_ASAP7_75t_L g408 ( 
.A1(n_409),
.A2(n_411),
.B1(n_412),
.B2(n_413),
.Y(n_408)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_409),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_411),
.Y(n_413)
);

MAJIxp5_ASAP7_75t_L g442 ( 
.A(n_411),
.B(n_412),
.C(n_414),
.Y(n_442)
);

AOI22xp5_ASAP7_75t_L g414 ( 
.A1(n_415),
.A2(n_416),
.B1(n_422),
.B2(n_425),
.Y(n_414)
);

MAJIxp5_ASAP7_75t_L g437 ( 
.A(n_415),
.B(n_423),
.C(n_424),
.Y(n_437)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_416),
.Y(n_415)
);

INVx3_ASAP7_75t_L g418 ( 
.A(n_419),
.Y(n_418)
);

INVx4_ASAP7_75t_L g419 ( 
.A(n_420),
.Y(n_419)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_422),
.Y(n_425)
);

XNOR2xp5_ASAP7_75t_SL g422 ( 
.A(n_423),
.B(n_424),
.Y(n_422)
);

INVxp67_ASAP7_75t_L g427 ( 
.A(n_428),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_SL g428 ( 
.A(n_429),
.B(n_441),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_430),
.Y(n_429)
);

OAI21xp5_ASAP7_75t_L g446 ( 
.A1(n_430),
.A2(n_447),
.B(n_448),
.Y(n_446)
);

NOR2x1_ASAP7_75t_L g430 ( 
.A(n_431),
.B(n_438),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_431),
.B(n_438),
.Y(n_448)
);

MAJIxp5_ASAP7_75t_L g431 ( 
.A(n_432),
.B(n_435),
.C(n_437),
.Y(n_431)
);

XOR2xp5_ASAP7_75t_L g443 ( 
.A(n_432),
.B(n_444),
.Y(n_443)
);

AOI22xp5_ASAP7_75t_L g444 ( 
.A1(n_435),
.A2(n_436),
.B1(n_437),
.B2(n_445),
.Y(n_444)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_436),
.Y(n_435)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_437),
.Y(n_445)
);

OR2x2_ASAP7_75t_L g441 ( 
.A(n_442),
.B(n_443),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_442),
.B(n_443),
.Y(n_447)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_450),
.Y(n_449)
);


endmodule