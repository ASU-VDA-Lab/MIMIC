module fake_jpeg_18253_n_254 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_254);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_254;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_11;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_12;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_96;

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_1),
.Y(n_11)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_6),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_2),
.Y(n_13)
);

BUFx5_ASAP7_75t_L g14 ( 
.A(n_9),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_5),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

INVx11_ASAP7_75t_SL g17 ( 
.A(n_3),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_10),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

INVx6_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_24),
.Y(n_37)
);

INVx11_ASAP7_75t_L g25 ( 
.A(n_17),
.Y(n_25)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_25),
.Y(n_36)
);

INVx8_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_26),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_15),
.B(n_22),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_27),
.B(n_29),
.Y(n_39)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_17),
.Y(n_28)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_28),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_12),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_SL g30 ( 
.A(n_19),
.B(n_10),
.Y(n_30)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_30),
.Y(n_34)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_21),
.Y(n_31)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_31),
.Y(n_41)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_21),
.Y(n_32)
);

BUFx16f_ASAP7_75t_L g40 ( 
.A(n_32),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_19),
.B(n_8),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_L g42 ( 
.A1(n_33),
.A2(n_11),
.B1(n_13),
.B2(n_12),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_42),
.B(n_30),
.Y(n_44)
);

INVx1_ASAP7_75t_SL g43 ( 
.A(n_41),
.Y(n_43)
);

INVx1_ASAP7_75t_SL g60 ( 
.A(n_43),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_L g76 ( 
.A1(n_44),
.A2(n_33),
.B1(n_29),
.B2(n_16),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_L g45 ( 
.A1(n_39),
.A2(n_32),
.B1(n_31),
.B2(n_26),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_45),
.A2(n_59),
.B1(n_26),
.B2(n_35),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g46 ( 
.A(n_39),
.B(n_27),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_46),
.B(n_48),
.Y(n_65)
);

BUFx2_ASAP7_75t_L g47 ( 
.A(n_38),
.Y(n_47)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_47),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_39),
.B(n_27),
.Y(n_48)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_38),
.Y(n_49)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_49),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_41),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_50),
.B(n_52),
.Y(n_72)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_35),
.Y(n_51)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_51),
.Y(n_70)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

BUFx2_ASAP7_75t_L g53 ( 
.A(n_38),
.Y(n_53)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_53),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_37),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_54),
.B(n_37),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_34),
.B(n_27),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_55),
.B(n_56),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_34),
.B(n_29),
.Y(n_56)
);

INVx2_ASAP7_75t_SL g57 ( 
.A(n_37),
.Y(n_57)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_57),
.Y(n_71)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_42),
.Y(n_58)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_58),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g59 ( 
.A1(n_35),
.A2(n_31),
.B1(n_32),
.B2(n_26),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_56),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_63),
.B(n_40),
.Y(n_92)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_57),
.Y(n_64)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_64),
.Y(n_90)
);

AND2x4_ASAP7_75t_L g68 ( 
.A(n_45),
.B(n_31),
.Y(n_68)
);

AND2x2_ASAP7_75t_L g94 ( 
.A(n_68),
.B(n_40),
.Y(n_94)
);

OAI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_58),
.A2(n_29),
.B1(n_32),
.B2(n_31),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_69),
.A2(n_73),
.B1(n_74),
.B2(n_26),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_48),
.A2(n_32),
.B1(n_26),
.B2(n_24),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_43),
.A2(n_24),
.B1(n_23),
.B2(n_25),
.Y(n_75)
);

INVxp67_ASAP7_75t_L g83 ( 
.A(n_75),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_76),
.B(n_44),
.Y(n_81)
);

CKINVDCx16_ASAP7_75t_R g93 ( 
.A(n_78),
.Y(n_93)
);

BUFx5_ASAP7_75t_L g79 ( 
.A(n_64),
.Y(n_79)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_79),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_80),
.A2(n_81),
.B1(n_71),
.B2(n_70),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_77),
.A2(n_24),
.B1(n_43),
.B2(n_57),
.Y(n_82)
);

INVxp67_ASAP7_75t_L g97 ( 
.A(n_82),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_77),
.A2(n_46),
.B1(n_55),
.B2(n_50),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_84),
.A2(n_65),
.B1(n_66),
.B2(n_63),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_68),
.A2(n_59),
.B1(n_51),
.B2(n_24),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_85),
.A2(n_73),
.B1(n_68),
.B2(n_74),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_78),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_86),
.B(n_92),
.Y(n_96)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_61),
.Y(n_87)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_87),
.Y(n_110)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_61),
.Y(n_88)
);

CKINVDCx16_ASAP7_75t_R g113 ( 
.A(n_88),
.Y(n_113)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_72),
.Y(n_89)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_89),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_65),
.B(n_40),
.C(n_51),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_91),
.B(n_37),
.C(n_40),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_94),
.B(n_37),
.Y(n_99)
);

CKINVDCx16_ASAP7_75t_R g95 ( 
.A(n_72),
.Y(n_95)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_95),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_98),
.B(n_100),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_SL g122 ( 
.A1(n_99),
.A2(n_107),
.B(n_67),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_89),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_L g101 ( 
.A1(n_83),
.A2(n_81),
.B(n_86),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_L g140 ( 
.A1(n_101),
.A2(n_115),
.B(n_13),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_102),
.A2(n_109),
.B1(n_93),
.B2(n_84),
.Y(n_117)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_79),
.Y(n_106)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_106),
.Y(n_118)
);

AND2x2_ASAP7_75t_L g107 ( 
.A(n_94),
.B(n_68),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_80),
.A2(n_68),
.B1(n_66),
.B2(n_60),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_108),
.A2(n_112),
.B1(n_83),
.B2(n_91),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_85),
.A2(n_60),
.B1(n_67),
.B2(n_62),
.Y(n_109)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_90),
.Y(n_111)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_111),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_95),
.B(n_71),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_114),
.B(n_53),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_94),
.A2(n_23),
.B1(n_16),
.B2(n_70),
.Y(n_115)
);

XNOR2xp5_ASAP7_75t_L g133 ( 
.A(n_116),
.B(n_40),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_117),
.A2(n_132),
.B1(n_143),
.B2(n_25),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_119),
.A2(n_125),
.B1(n_127),
.B2(n_136),
.Y(n_155)
);

AND2x2_ASAP7_75t_L g120 ( 
.A(n_104),
.B(n_88),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_SL g146 ( 
.A1(n_120),
.A2(n_113),
.B(n_99),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_101),
.A2(n_90),
.B1(n_87),
.B2(n_23),
.Y(n_121)
);

INVxp67_ASAP7_75t_L g158 ( 
.A(n_121),
.Y(n_158)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_122),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_114),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_123),
.B(n_128),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_108),
.A2(n_62),
.B1(n_52),
.B2(n_49),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_97),
.A2(n_54),
.B1(n_36),
.B2(n_28),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_104),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_110),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_129),
.B(n_135),
.Y(n_162)
);

XOR2xp5_ASAP7_75t_L g130 ( 
.A(n_98),
.B(n_33),
.Y(n_130)
);

XOR2xp5_ASAP7_75t_L g164 ( 
.A(n_130),
.B(n_137),
.Y(n_164)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_131),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_102),
.A2(n_36),
.B1(n_28),
.B2(n_57),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_L g147 ( 
.A(n_133),
.B(n_138),
.Y(n_147)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_111),
.Y(n_134)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_134),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_105),
.B(n_30),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_97),
.A2(n_36),
.B1(n_28),
.B2(n_53),
.Y(n_136)
);

XOR2xp5_ASAP7_75t_L g137 ( 
.A(n_96),
.B(n_14),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_L g138 ( 
.A(n_96),
.B(n_30),
.Y(n_138)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_105),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_139),
.Y(n_148)
);

XNOR2xp5_ASAP7_75t_L g150 ( 
.A(n_140),
.B(n_115),
.Y(n_150)
);

XOR2xp5_ASAP7_75t_L g141 ( 
.A(n_116),
.B(n_20),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_SL g151 ( 
.A(n_141),
.B(n_107),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_107),
.A2(n_28),
.B1(n_47),
.B2(n_25),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_142),
.A2(n_136),
.B1(n_127),
.B2(n_125),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_109),
.A2(n_11),
.B1(n_47),
.B2(n_22),
.Y(n_143)
);

OA21x2_ASAP7_75t_L g144 ( 
.A1(n_126),
.A2(n_121),
.B(n_117),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_144),
.B(n_165),
.Y(n_181)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_146),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_150),
.B(n_140),
.Y(n_169)
);

XOR2xp5_ASAP7_75t_L g170 ( 
.A(n_151),
.B(n_153),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_120),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_152),
.B(n_154),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_L g153 ( 
.A(n_137),
.B(n_103),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_120),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_133),
.B(n_106),
.C(n_103),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_156),
.B(n_18),
.C(n_14),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g157 ( 
.A(n_119),
.B(n_20),
.Y(n_157)
);

XOR2xp5_ASAP7_75t_L g174 ( 
.A(n_157),
.B(n_161),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_124),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_159),
.B(n_148),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_160),
.A2(n_143),
.B1(n_25),
.B2(n_2),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_SL g161 ( 
.A(n_130),
.B(n_20),
.Y(n_161)
);

INVxp33_ASAP7_75t_L g165 ( 
.A(n_142),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_166),
.A2(n_22),
.B1(n_15),
.B2(n_18),
.Y(n_183)
);

XOR2xp5_ASAP7_75t_L g193 ( 
.A(n_169),
.B(n_164),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_156),
.B(n_141),
.C(n_118),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_171),
.B(n_185),
.C(n_151),
.Y(n_195)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_145),
.Y(n_172)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_172),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_175),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_147),
.B(n_138),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_L g191 ( 
.A(n_176),
.B(n_178),
.Y(n_191)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_167),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_177),
.B(n_179),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_L g178 ( 
.A(n_147),
.B(n_132),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_158),
.A2(n_18),
.B1(n_22),
.B2(n_15),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_180),
.A2(n_183),
.B1(n_155),
.B2(n_1),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_162),
.B(n_0),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_182),
.B(n_184),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_SL g184 ( 
.A(n_149),
.B(n_0),
.Y(n_184)
);

BUFx24_ASAP7_75t_SL g186 ( 
.A(n_176),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_186),
.B(n_189),
.Y(n_208)
);

CKINVDCx16_ASAP7_75t_R g189 ( 
.A(n_173),
.Y(n_189)
);

AOI21xp5_ASAP7_75t_L g190 ( 
.A1(n_168),
.A2(n_163),
.B(n_158),
.Y(n_190)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_190),
.Y(n_212)
);

INVxp33_ASAP7_75t_L g192 ( 
.A(n_181),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_192),
.B(n_194),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_193),
.B(n_198),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g194 ( 
.A(n_171),
.B(n_153),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g209 ( 
.A(n_195),
.B(n_174),
.Y(n_209)
);

OAI21xp5_ASAP7_75t_L g197 ( 
.A1(n_185),
.A2(n_144),
.B(n_150),
.Y(n_197)
);

AOI21xp5_ASAP7_75t_L g211 ( 
.A1(n_197),
.A2(n_0),
.B(n_1),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g198 ( 
.A(n_170),
.B(n_164),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_178),
.B(n_157),
.C(n_161),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_199),
.B(n_174),
.C(n_170),
.Y(n_204)
);

CKINVDCx16_ASAP7_75t_R g202 ( 
.A(n_201),
.Y(n_202)
);

CKINVDCx16_ASAP7_75t_R g203 ( 
.A(n_187),
.Y(n_203)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_203),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_L g218 ( 
.A(n_204),
.B(n_209),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_200),
.A2(n_188),
.B1(n_169),
.B2(n_192),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_207),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_224)
);

AOI21xp33_ASAP7_75t_L g210 ( 
.A1(n_195),
.A2(n_165),
.B(n_144),
.Y(n_210)
);

AOI21xp5_ASAP7_75t_L g217 ( 
.A1(n_210),
.A2(n_191),
.B(n_2),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_211),
.B(n_213),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_198),
.B(n_0),
.Y(n_213)
);

BUFx6f_ASAP7_75t_L g214 ( 
.A(n_196),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_214),
.B(n_2),
.C(n_3),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_L g216 ( 
.A1(n_202),
.A2(n_199),
.B1(n_193),
.B2(n_191),
.Y(n_216)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_216),
.Y(n_228)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_217),
.Y(n_231)
);

NOR2x1_ASAP7_75t_L g220 ( 
.A(n_212),
.B(n_1),
.Y(n_220)
);

NAND2x1p5_ASAP7_75t_L g225 ( 
.A(n_220),
.B(n_4),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_221),
.B(n_223),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_205),
.A2(n_209),
.B1(n_214),
.B2(n_208),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_L g232 ( 
.A1(n_222),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_213),
.B(n_3),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_224),
.B(n_4),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_225),
.B(n_229),
.Y(n_237)
);

AOI21x1_ASAP7_75t_L g226 ( 
.A1(n_215),
.A2(n_204),
.B(n_206),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g235 ( 
.A(n_226),
.B(n_232),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_218),
.B(n_206),
.Y(n_230)
);

OR2x2_ASAP7_75t_L g238 ( 
.A(n_230),
.B(n_233),
.Y(n_238)
);

INVx6_ASAP7_75t_L g233 ( 
.A(n_220),
.Y(n_233)
);

NOR3xp33_ASAP7_75t_SL g234 ( 
.A(n_225),
.B(n_218),
.C(n_219),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_234),
.B(n_236),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_L g236 ( 
.A1(n_228),
.A2(n_231),
.B1(n_233),
.B2(n_227),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_230),
.B(n_219),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_239),
.B(n_241),
.Y(n_243)
);

OAI21xp5_ASAP7_75t_L g240 ( 
.A1(n_228),
.A2(n_221),
.B(n_223),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_SL g246 ( 
.A(n_240),
.B(n_7),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g241 ( 
.A(n_226),
.B(n_7),
.Y(n_241)
);

BUFx6f_ASAP7_75t_L g244 ( 
.A(n_238),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_244),
.B(n_245),
.Y(n_247)
);

OAI21xp5_ASAP7_75t_SL g245 ( 
.A1(n_235),
.A2(n_7),
.B(n_8),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_246),
.B(n_237),
.Y(n_248)
);

INVxp33_ASAP7_75t_L g249 ( 
.A(n_248),
.Y(n_249)
);

AOI21xp5_ASAP7_75t_SL g250 ( 
.A1(n_247),
.A2(n_242),
.B(n_243),
.Y(n_250)
);

AO21x1_ASAP7_75t_L g251 ( 
.A1(n_250),
.A2(n_237),
.B(n_7),
.Y(n_251)
);

BUFx24_ASAP7_75t_SL g252 ( 
.A(n_251),
.Y(n_252)
);

BUFx24_ASAP7_75t_SL g253 ( 
.A(n_252),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_253),
.B(n_249),
.Y(n_254)
);


endmodule