module fake_jpeg_29687_n_253 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_253);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_253;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_122;
wire n_75;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx4f_ASAP7_75t_L g18 ( 
.A(n_16),
.Y(n_18)
);

BUFx24_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

INVx8_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_15),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_8),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_11),
.Y(n_27)
);

INVx11_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_3),
.B(n_4),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

INVx5_ASAP7_75t_L g34 ( 
.A(n_13),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_4),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_1),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_5),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_0),
.Y(n_38)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_15),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_9),
.Y(n_40)
);

BUFx5_ASAP7_75t_L g41 ( 
.A(n_37),
.Y(n_41)
);

BUFx2_ASAP7_75t_L g71 ( 
.A(n_41),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_31),
.B(n_17),
.Y(n_42)
);

AND2x2_ASAP7_75t_L g74 ( 
.A(n_42),
.B(n_59),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g43 ( 
.A(n_23),
.B(n_0),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_43),
.B(n_46),
.Y(n_80)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_19),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g85 ( 
.A(n_44),
.Y(n_85)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_32),
.Y(n_45)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_45),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_32),
.B(n_0),
.Y(n_46)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_19),
.Y(n_47)
);

BUFx10_ASAP7_75t_L g79 ( 
.A(n_47),
.Y(n_79)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_35),
.Y(n_48)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_48),
.Y(n_70)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_49),
.Y(n_82)
);

INVx5_ASAP7_75t_L g50 ( 
.A(n_28),
.Y(n_50)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_50),
.Y(n_75)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_24),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_51),
.Y(n_81)
);

BUFx5_ASAP7_75t_L g52 ( 
.A(n_37),
.Y(n_52)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_52),
.Y(n_73)
);

BUFx5_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

INVx6_ASAP7_75t_L g89 ( 
.A(n_53),
.Y(n_89)
);

OR2x2_ASAP7_75t_L g54 ( 
.A(n_23),
.B(n_2),
.Y(n_54)
);

OR2x2_ASAP7_75t_L g86 ( 
.A(n_54),
.B(n_60),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_28),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_55),
.Y(n_101)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_24),
.Y(n_56)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_56),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_29),
.Y(n_57)
);

INVx6_ASAP7_75t_L g102 ( 
.A(n_57),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_SL g58 ( 
.A(n_22),
.B(n_17),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_58),
.B(n_62),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_22),
.B(n_16),
.Y(n_59)
);

OR2x2_ASAP7_75t_L g60 ( 
.A(n_40),
.B(n_2),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_40),
.B(n_3),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_61),
.B(n_66),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_27),
.B(n_12),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_SL g63 ( 
.A(n_27),
.B(n_12),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_63),
.B(n_14),
.Y(n_87)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_29),
.Y(n_64)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_64),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_36),
.Y(n_65)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_65),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_25),
.B(n_5),
.Y(n_66)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_20),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_67),
.Y(n_96)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_36),
.Y(n_68)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_68),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_51),
.A2(n_39),
.B1(n_38),
.B2(n_18),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_72),
.A2(n_94),
.B1(n_100),
.B2(n_65),
.Y(n_105)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_45),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_77),
.B(n_78),
.Y(n_104)
);

INVxp67_ASAP7_75t_L g78 ( 
.A(n_44),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_SL g83 ( 
.A(n_46),
.B(n_33),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_SL g126 ( 
.A(n_83),
.B(n_87),
.Y(n_126)
);

BUFx12_ASAP7_75t_L g90 ( 
.A(n_50),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_90),
.B(n_99),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_54),
.B(n_33),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g127 ( 
.A(n_91),
.B(n_98),
.Y(n_127)
);

OAI22xp33_ASAP7_75t_L g94 ( 
.A1(n_64),
.A2(n_38),
.B1(n_18),
.B2(n_39),
.Y(n_94)
);

BUFx16f_ASAP7_75t_L g95 ( 
.A(n_44),
.Y(n_95)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_95),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_60),
.B(n_25),
.Y(n_98)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_48),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_56),
.A2(n_18),
.B1(n_34),
.B2(n_30),
.Y(n_100)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_69),
.Y(n_103)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_103),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_105),
.A2(n_114),
.B1(n_6),
.B2(n_8),
.Y(n_147)
);

AO22x1_ASAP7_75t_SL g107 ( 
.A1(n_70),
.A2(n_49),
.B1(n_68),
.B2(n_57),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_107),
.A2(n_116),
.B1(n_128),
.B2(n_85),
.Y(n_148)
);

AND2x2_ASAP7_75t_L g108 ( 
.A(n_80),
.B(n_53),
.Y(n_108)
);

XNOR2xp5_ASAP7_75t_L g155 ( 
.A(n_108),
.B(n_115),
.Y(n_155)
);

CKINVDCx16_ASAP7_75t_R g109 ( 
.A(n_95),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_109),
.B(n_129),
.Y(n_141)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_76),
.Y(n_111)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_111),
.Y(n_150)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_92),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_112),
.B(n_119),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_84),
.B(n_26),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_SL g145 ( 
.A(n_113),
.B(n_131),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_88),
.A2(n_67),
.B1(n_55),
.B2(n_20),
.Y(n_114)
);

AND2x2_ASAP7_75t_L g115 ( 
.A(n_82),
.B(n_52),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_L g116 ( 
.A1(n_94),
.A2(n_37),
.B1(n_21),
.B2(n_30),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_86),
.B(n_26),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_117),
.B(n_132),
.Y(n_144)
);

AND2x2_ASAP7_75t_SL g118 ( 
.A(n_93),
.B(n_41),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_118),
.B(n_85),
.C(n_90),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_79),
.Y(n_119)
);

INVx1_ASAP7_75t_SL g120 ( 
.A(n_78),
.Y(n_120)
);

INVxp67_ASAP7_75t_L g143 ( 
.A(n_120),
.Y(n_143)
);

INVx6_ASAP7_75t_L g121 ( 
.A(n_102),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_121),
.Y(n_140)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_97),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_122),
.B(n_130),
.Y(n_157)
);

OR2x4_ASAP7_75t_L g123 ( 
.A(n_86),
.B(n_19),
.Y(n_123)
);

O2A1O1Ixp33_ASAP7_75t_L g153 ( 
.A1(n_123),
.A2(n_125),
.B(n_10),
.C(n_117),
.Y(n_153)
);

INVx8_ASAP7_75t_L g124 ( 
.A(n_73),
.Y(n_124)
);

INVx4_ASAP7_75t_L g134 ( 
.A(n_124),
.Y(n_134)
);

OR2x4_ASAP7_75t_L g125 ( 
.A(n_74),
.B(n_21),
.Y(n_125)
);

AO22x1_ASAP7_75t_SL g128 ( 
.A1(n_81),
.A2(n_47),
.B1(n_34),
.B2(n_7),
.Y(n_128)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_79),
.Y(n_129)
);

A2O1A1Ixp33_ASAP7_75t_L g130 ( 
.A1(n_74),
.A2(n_47),
.B(n_14),
.C(n_7),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_96),
.B(n_5),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_81),
.B(n_6),
.Y(n_132)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_75),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_133),
.B(n_111),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_104),
.Y(n_136)
);

OR2x2_ASAP7_75t_L g160 ( 
.A(n_136),
.B(n_137),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_106),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_108),
.A2(n_102),
.B1(n_101),
.B2(n_73),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_138),
.A2(n_142),
.B1(n_158),
.B2(n_118),
.Y(n_171)
);

AOI32xp33_ASAP7_75t_L g139 ( 
.A1(n_123),
.A2(n_89),
.A3(n_71),
.B1(n_90),
.B2(n_79),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_139),
.B(n_151),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_108),
.A2(n_101),
.B1(n_89),
.B2(n_71),
.Y(n_142)
);

XNOR2x1_ASAP7_75t_L g166 ( 
.A(n_146),
.B(n_118),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_147),
.A2(n_149),
.B1(n_128),
.B2(n_130),
.Y(n_170)
);

CKINVDCx16_ASAP7_75t_R g162 ( 
.A(n_148),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_105),
.A2(n_8),
.B1(n_10),
.B2(n_85),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_115),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_127),
.B(n_10),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_152),
.B(n_153),
.Y(n_167)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_154),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_132),
.B(n_114),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_156),
.B(n_107),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_107),
.A2(n_128),
.B1(n_112),
.B2(n_122),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_161),
.B(n_169),
.Y(n_183)
);

BUFx12_ASAP7_75t_L g165 ( 
.A(n_159),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_165),
.B(n_177),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_SL g198 ( 
.A1(n_166),
.A2(n_181),
.B(n_140),
.Y(n_198)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_150),
.Y(n_168)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_168),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_144),
.B(n_103),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_170),
.B(n_171),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_144),
.B(n_115),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_172),
.B(n_174),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_SL g173 ( 
.A(n_157),
.B(n_126),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_SL g189 ( 
.A(n_173),
.B(n_141),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_156),
.B(n_133),
.Y(n_174)
);

AND2x6_ASAP7_75t_L g175 ( 
.A(n_153),
.B(n_125),
.Y(n_175)
);

NOR3xp33_ASAP7_75t_L g182 ( 
.A(n_175),
.B(n_137),
.C(n_136),
.Y(n_182)
);

INVx4_ASAP7_75t_L g176 ( 
.A(n_134),
.Y(n_176)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_176),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_155),
.B(n_120),
.C(n_124),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_147),
.A2(n_121),
.B1(n_129),
.B2(n_110),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_L g199 ( 
.A1(n_178),
.A2(n_140),
.B1(n_162),
.B2(n_161),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_145),
.B(n_110),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_179),
.B(n_180),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_135),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_SL g181 ( 
.A1(n_146),
.A2(n_154),
.B(n_155),
.Y(n_181)
);

INVxp67_ASAP7_75t_L g211 ( 
.A(n_182),
.Y(n_211)
);

OAI21xp5_ASAP7_75t_L g185 ( 
.A1(n_164),
.A2(n_151),
.B(n_149),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_L g213 ( 
.A1(n_185),
.A2(n_174),
.B(n_172),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_162),
.A2(n_158),
.B1(n_148),
.B2(n_150),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_187),
.A2(n_199),
.B1(n_171),
.B2(n_178),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_189),
.B(n_196),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_160),
.B(n_143),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_190),
.B(n_193),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_160),
.B(n_143),
.Y(n_193)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_168),
.Y(n_195)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_195),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_160),
.B(n_134),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_180),
.B(n_159),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_197),
.B(n_165),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_SL g207 ( 
.A(n_198),
.B(n_181),
.Y(n_207)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_202),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_183),
.B(n_163),
.Y(n_203)
);

OAI21x1_ASAP7_75t_L g224 ( 
.A1(n_203),
.A2(n_208),
.B(n_209),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_186),
.Y(n_204)
);

AOI21xp5_ASAP7_75t_L g221 ( 
.A1(n_204),
.A2(n_205),
.B(n_167),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_186),
.Y(n_205)
);

CKINVDCx16_ASAP7_75t_R g206 ( 
.A(n_191),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_L g220 ( 
.A1(n_206),
.A2(n_212),
.B1(n_213),
.B2(n_214),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_SL g225 ( 
.A(n_207),
.B(n_185),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_183),
.B(n_163),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_189),
.B(n_173),
.Y(n_209)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_191),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_207),
.B(n_198),
.C(n_184),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_215),
.B(n_218),
.C(n_222),
.Y(n_229)
);

A2O1A1Ixp33_ASAP7_75t_L g216 ( 
.A1(n_211),
.A2(n_192),
.B(n_193),
.C(n_190),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_216),
.B(n_219),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_213),
.B(n_177),
.Y(n_217)
);

XOR2xp5_ASAP7_75t_L g227 ( 
.A(n_217),
.B(n_200),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_203),
.B(n_166),
.C(n_188),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_204),
.A2(n_199),
.B1(n_187),
.B2(n_170),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_221),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_208),
.B(n_188),
.C(n_192),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_SL g228 ( 
.A(n_225),
.B(n_200),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g235 ( 
.A(n_227),
.B(n_228),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_222),
.A2(n_214),
.B1(n_211),
.B2(n_205),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_230),
.A2(n_220),
.B1(n_217),
.B2(n_216),
.Y(n_236)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_224),
.Y(n_232)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_232),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_223),
.B(n_201),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_233),
.B(n_169),
.Y(n_239)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_236),
.B(n_228),
.Y(n_242)
);

AOI21xp5_ASAP7_75t_SL g237 ( 
.A1(n_232),
.A2(n_225),
.B(n_210),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_237),
.B(n_238),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_231),
.A2(n_226),
.B1(n_230),
.B2(n_206),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_239),
.B(n_194),
.Y(n_244)
);

AOI21xp5_ASAP7_75t_L g240 ( 
.A1(n_229),
.A2(n_215),
.B(n_212),
.Y(n_240)
);

AOI21xp5_ASAP7_75t_L g245 ( 
.A1(n_240),
.A2(n_218),
.B(n_194),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_242),
.B(n_245),
.Y(n_247)
);

AOI322xp5_ASAP7_75t_L g243 ( 
.A1(n_234),
.A2(n_175),
.A3(n_237),
.B1(n_210),
.B2(n_229),
.C1(n_227),
.C2(n_195),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_243),
.B(n_244),
.Y(n_246)
);

AOI21xp5_ASAP7_75t_L g248 ( 
.A1(n_241),
.A2(n_235),
.B(n_176),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_SL g249 ( 
.A(n_248),
.B(n_242),
.Y(n_249)
);

NOR3xp33_ASAP7_75t_SL g251 ( 
.A(n_249),
.B(n_250),
.C(n_247),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_246),
.B(n_165),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g252 ( 
.A(n_251),
.B(n_235),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_252),
.B(n_165),
.Y(n_253)
);


endmodule