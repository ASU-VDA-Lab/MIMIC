module real_jpeg_15987_n_19 (n_17, n_8, n_0, n_2, n_132, n_139, n_10, n_137, n_9, n_129, n_12, n_135, n_130, n_134, n_6, n_136, n_128, n_133, n_11, n_14, n_131, n_138, n_7, n_18, n_3, n_5, n_4, n_1, n_16, n_15, n_13, n_19);

input n_17;
input n_8;
input n_0;
input n_2;
input n_132;
input n_139;
input n_10;
input n_137;
input n_9;
input n_129;
input n_12;
input n_135;
input n_130;
input n_134;
input n_6;
input n_136;
input n_128;
input n_133;
input n_11;
input n_14;
input n_131;
input n_138;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;

output n_19;

wire n_108;
wire n_54;
wire n_37;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_78;
wire n_83;
wire n_104;
wire n_64;
wire n_47;
wire n_22;
wire n_87;
wire n_40;
wire n_105;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_126;
wire n_113;
wire n_120;
wire n_93;
wire n_95;
wire n_33;
wire n_65;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_66;
wire n_28;
wire n_44;
wire n_62;
wire n_121;
wire n_106;
wire n_45;
wire n_112;
wire n_42;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_118;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_69;
wire n_31;
wire n_72;
wire n_100;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_117;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_30;
wire n_103;
wire n_43;
wire n_57;
wire n_84;
wire n_82;
wire n_111;
wire n_125;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_25;
wire n_53;
wire n_119;
wire n_36;
wire n_102;
wire n_81;
wire n_85;
wire n_101;
wire n_96;
wire n_89;

NOR2xp33_ASAP7_75t_SL g110 ( 
.A(n_0),
.B(n_111),
.Y(n_110)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_0),
.Y(n_115)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_1),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_1),
.B(n_43),
.Y(n_105)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

NOR2xp67_ASAP7_75t_L g62 ( 
.A(n_3),
.B(n_63),
.Y(n_62)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_3),
.Y(n_108)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

AND2x2_ASAP7_75t_L g78 ( 
.A(n_5),
.B(n_79),
.Y(n_78)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_6),
.Y(n_91)
);

AOI21x1_ASAP7_75t_L g75 ( 
.A1(n_7),
.A2(n_76),
.B(n_85),
.Y(n_75)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_7),
.Y(n_87)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_8),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_SL g86 ( 
.A(n_8),
.B(n_78),
.C(n_83),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_9),
.B(n_50),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_9),
.B(n_50),
.Y(n_101)
);

MAJx2_ASAP7_75t_L g73 ( 
.A(n_10),
.B(n_74),
.C(n_96),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_SL g120 ( 
.A(n_11),
.B(n_121),
.Y(n_120)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_11),
.Y(n_125)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_12),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_12),
.B(n_57),
.Y(n_102)
);

XOR2xp5_ASAP7_75t_L g20 ( 
.A(n_13),
.B(n_21),
.Y(n_20)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_14),
.Y(n_112)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_15),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_16),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_16),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_16),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_16),
.Y(n_65)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_17),
.Y(n_68)
);

AOI322xp5_ASAP7_75t_SL g103 ( 
.A1(n_17),
.A2(n_54),
.A3(n_67),
.B1(n_70),
.B2(n_104),
.C1(n_106),
.C2(n_139),
.Y(n_103)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_18),
.Y(n_36)
);

XOR2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_26),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_23),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_24),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

AOI21xp5_ASAP7_75t_SL g26 ( 
.A1(n_27),
.A2(n_119),
.B(n_124),
.Y(n_26)
);

OAI21xp5_ASAP7_75t_L g27 ( 
.A1(n_28),
.A2(n_37),
.B(n_117),
.Y(n_27)
);

INVxp67_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_SL g29 ( 
.A(n_30),
.B(n_36),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_30),
.B(n_36),
.Y(n_118)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_32),
.B(n_33),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

NOR2x1_ASAP7_75t_L g83 ( 
.A(n_34),
.B(n_84),
.Y(n_83)
);

BUFx4f_ASAP7_75t_SL g34 ( 
.A(n_35),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_35),
.Y(n_52)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_35),
.Y(n_59)
);

BUFx5_ASAP7_75t_L g95 ( 
.A(n_35),
.Y(n_95)
);

AOI21xp5_ASAP7_75t_SL g37 ( 
.A1(n_38),
.A2(n_109),
.B(n_114),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

AOI31xp67_ASAP7_75t_L g39 ( 
.A1(n_40),
.A2(n_48),
.A3(n_73),
.B(n_100),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_41),
.B(n_42),
.Y(n_40)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_44),
.B(n_45),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_SL g89 ( 
.A(n_45),
.B(n_90),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

NOR3xp33_ASAP7_75t_SL g48 ( 
.A(n_49),
.B(n_53),
.C(n_60),
.Y(n_48)
);

NOR3xp33_ASAP7_75t_L g104 ( 
.A(n_49),
.B(n_62),
.C(n_105),
.Y(n_104)
);

NOR2x1_ASAP7_75t_L g50 ( 
.A(n_51),
.B(n_52),
.Y(n_50)
);

BUFx2_ASAP7_75t_L g99 ( 
.A(n_52),
.Y(n_99)
);

OAI321xp33_ASAP7_75t_L g100 ( 
.A1(n_53),
.A2(n_60),
.A3(n_101),
.B1(n_102),
.B2(n_103),
.C(n_138),
.Y(n_100)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_55),
.B(n_56),
.Y(n_54)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_58),
.B(n_59),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_61),
.B(n_67),
.Y(n_60)
);

INVxp67_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_63),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_SL g63 ( 
.A(n_64),
.B(n_66),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

BUFx12f_ASAP7_75t_L g71 ( 
.A(n_65),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_65),
.B(n_80),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_68),
.B(n_69),
.Y(n_67)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g70 ( 
.A(n_71),
.B(n_72),
.Y(n_70)
);

BUFx3_ASAP7_75t_L g123 ( 
.A(n_71),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g74 ( 
.A(n_75),
.B(n_91),
.C(n_92),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_L g76 ( 
.A(n_77),
.B(n_81),
.C(n_82),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

AOI21xp5_ASAP7_75t_L g85 ( 
.A1(n_86),
.A2(n_87),
.B(n_88),
.Y(n_85)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_95),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_98),
.Y(n_96)
);

BUFx3_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g106 ( 
.A(n_107),
.B(n_108),
.Y(n_106)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_111),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_112),
.B(n_113),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_115),
.B(n_116),
.Y(n_114)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_121),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_122),
.B(n_123),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_125),
.B(n_126),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_128),
.Y(n_44)
);

CKINVDCx16_ASAP7_75t_R g51 ( 
.A(n_129),
.Y(n_51)
);

INVxp67_ASAP7_75t_L g58 ( 
.A(n_130),
.Y(n_58)
);

INVxp67_ASAP7_75t_L g66 ( 
.A(n_131),
.Y(n_66)
);

INVxp67_ASAP7_75t_L g72 ( 
.A(n_132),
.Y(n_72)
);

INVxp67_ASAP7_75t_L g80 ( 
.A(n_133),
.Y(n_80)
);

CKINVDCx16_ASAP7_75t_R g84 ( 
.A(n_134),
.Y(n_84)
);

CKINVDCx16_ASAP7_75t_R g90 ( 
.A(n_135),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_136),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_137),
.Y(n_97)
);


endmodule