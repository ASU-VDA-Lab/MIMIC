module fake_jpeg_17078_n_343 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_343);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_343;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx3_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

INVx2_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

BUFx16f_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_4),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

INVx1_ASAP7_75t_SL g23 ( 
.A(n_8),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

INVxp33_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

CKINVDCx16_ASAP7_75t_R g27 ( 
.A(n_3),
.Y(n_27)
);

BUFx16f_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

INVx1_ASAP7_75t_SL g30 ( 
.A(n_12),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_0),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_4),
.Y(n_34)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_2),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_18),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_36),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_19),
.Y(n_37)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_37),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_17),
.B(n_0),
.Y(n_38)
);

AND2x2_ASAP7_75t_L g52 ( 
.A(n_38),
.B(n_40),
.Y(n_52)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_17),
.Y(n_39)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_39),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_23),
.B(n_0),
.Y(n_40)
);

INVx5_ASAP7_75t_SL g41 ( 
.A(n_19),
.Y(n_41)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_41),
.A2(n_30),
.B1(n_35),
.B2(n_33),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_23),
.B(n_1),
.Y(n_42)
);

AND2x2_ASAP7_75t_L g64 ( 
.A(n_42),
.B(n_48),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_18),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_43),
.Y(n_69)
);

BUFx6f_ASAP7_75t_SL g44 ( 
.A(n_19),
.Y(n_44)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_44),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_SL g45 ( 
.A(n_26),
.B(n_14),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_45),
.B(n_30),
.Y(n_50)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_16),
.Y(n_46)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_46),
.Y(n_59)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_33),
.Y(n_47)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_47),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_24),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_50),
.B(n_48),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_46),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_51),
.B(n_53),
.Y(n_79)
);

HB1xp67_ASAP7_75t_L g53 ( 
.A(n_46),
.Y(n_53)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_47),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g77 ( 
.A(n_56),
.Y(n_77)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_39),
.Y(n_58)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_58),
.Y(n_91)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_39),
.Y(n_60)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_60),
.Y(n_101)
);

AOI21xp33_ASAP7_75t_L g61 ( 
.A1(n_45),
.A2(n_28),
.B(n_34),
.Y(n_61)
);

AND2x2_ASAP7_75t_L g87 ( 
.A(n_61),
.B(n_68),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_45),
.B(n_30),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_62),
.B(n_66),
.Y(n_103)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_47),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g106 ( 
.A(n_63),
.Y(n_106)
);

CKINVDCx14_ASAP7_75t_R g85 ( 
.A(n_65),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_40),
.B(n_31),
.Y(n_66)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_39),
.Y(n_67)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_67),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_48),
.A2(n_35),
.B1(n_28),
.B2(n_27),
.Y(n_68)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_47),
.Y(n_70)
);

INVx11_ASAP7_75t_L g96 ( 
.A(n_70),
.Y(n_96)
);

OAI22xp33_ASAP7_75t_L g71 ( 
.A1(n_47),
.A2(n_19),
.B1(n_28),
.B2(n_18),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_71),
.A2(n_41),
.B1(n_44),
.B2(n_42),
.Y(n_78)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_36),
.Y(n_72)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_72),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_38),
.B(n_34),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_73),
.B(n_38),
.Y(n_83)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_44),
.Y(n_74)
);

HB1xp67_ASAP7_75t_L g89 ( 
.A(n_74),
.Y(n_89)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_58),
.Y(n_76)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_76),
.Y(n_126)
);

OAI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_78),
.A2(n_108),
.B1(n_63),
.B2(n_56),
.Y(n_129)
);

INVxp67_ASAP7_75t_L g80 ( 
.A(n_59),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_80),
.B(n_82),
.Y(n_117)
);

AND2x4_ASAP7_75t_L g81 ( 
.A(n_64),
.B(n_44),
.Y(n_81)
);

AND2x2_ASAP7_75t_L g114 ( 
.A(n_81),
.B(n_43),
.Y(n_114)
);

INVx5_ASAP7_75t_L g82 ( 
.A(n_55),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_83),
.B(n_24),
.Y(n_118)
);

INVx13_ASAP7_75t_L g84 ( 
.A(n_75),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_84),
.B(n_88),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_52),
.B(n_38),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_86),
.B(n_98),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_75),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_90),
.B(n_93),
.Y(n_125)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_59),
.Y(n_92)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_92),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_73),
.B(n_42),
.Y(n_93)
);

CKINVDCx14_ASAP7_75t_R g94 ( 
.A(n_68),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_94),
.B(n_95),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_57),
.Y(n_95)
);

INVx4_ASAP7_75t_L g97 ( 
.A(n_57),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_97),
.B(n_104),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_52),
.B(n_42),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_52),
.A2(n_40),
.B1(n_28),
.B2(n_43),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_99),
.A2(n_105),
.B1(n_86),
.B2(n_98),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_64),
.B(n_37),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_100),
.B(n_110),
.Y(n_138)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_49),
.Y(n_102)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_102),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_64),
.B(n_31),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_49),
.A2(n_43),
.B1(n_36),
.B2(n_41),
.Y(n_105)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_69),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_107),
.B(n_22),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_L g108 ( 
.A1(n_60),
.A2(n_67),
.B1(n_54),
.B2(n_70),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_54),
.B(n_37),
.Y(n_110)
);

A2O1A1Ixp33_ASAP7_75t_SL g111 ( 
.A1(n_71),
.A2(n_41),
.B(n_43),
.C(n_36),
.Y(n_111)
);

AOI21xp5_ASAP7_75t_L g115 ( 
.A1(n_111),
.A2(n_55),
.B(n_74),
.Y(n_115)
);

MAJx2_ASAP7_75t_L g113 ( 
.A(n_81),
.B(n_41),
.C(n_37),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_113),
.B(n_132),
.C(n_16),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_L g147 ( 
.A1(n_114),
.A2(n_134),
.B(n_141),
.Y(n_147)
);

O2A1O1Ixp33_ASAP7_75t_L g168 ( 
.A1(n_115),
.A2(n_77),
.B(n_21),
.C(n_22),
.Y(n_168)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_110),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_116),
.B(n_123),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_118),
.B(n_20),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_101),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_119),
.B(n_121),
.Y(n_165)
);

CKINVDCx16_ASAP7_75t_R g121 ( 
.A(n_79),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_122),
.A2(n_129),
.B1(n_130),
.B2(n_133),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_101),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_83),
.B(n_25),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_127),
.B(n_139),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_85),
.A2(n_81),
.B1(n_100),
.B2(n_87),
.Y(n_130)
);

MAJx2_ASAP7_75t_L g132 ( 
.A(n_81),
.B(n_87),
.C(n_99),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_81),
.A2(n_72),
.B1(n_36),
.B2(n_69),
.Y(n_133)
);

AND2x2_ASAP7_75t_L g134 ( 
.A(n_78),
.B(n_1),
.Y(n_134)
);

INVxp67_ASAP7_75t_L g135 ( 
.A(n_102),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_135),
.B(n_106),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_87),
.B(n_37),
.Y(n_139)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_140),
.Y(n_151)
);

AND2x2_ASAP7_75t_L g141 ( 
.A(n_105),
.B(n_1),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_90),
.B(n_25),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_142),
.B(n_96),
.Y(n_157)
);

A2O1A1O1Ixp25_ASAP7_75t_L g144 ( 
.A1(n_132),
.A2(n_103),
.B(n_111),
.C(n_80),
.D(n_92),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_SL g182 ( 
.A1(n_144),
.A2(n_152),
.B(n_168),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_137),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_146),
.B(n_150),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_134),
.A2(n_111),
.B1(n_91),
.B2(n_76),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g204 ( 
.A1(n_148),
.A2(n_149),
.B1(n_153),
.B2(n_160),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_134),
.A2(n_111),
.B1(n_91),
.B2(n_109),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_137),
.Y(n_150)
);

AOI21xp5_ASAP7_75t_L g152 ( 
.A1(n_128),
.A2(n_111),
.B(n_82),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_134),
.A2(n_109),
.B1(n_112),
.B2(n_95),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_131),
.Y(n_154)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_154),
.Y(n_185)
);

CKINVDCx14_ASAP7_75t_R g155 ( 
.A(n_120),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_155),
.B(n_156),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_131),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_157),
.B(n_158),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_124),
.B(n_112),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_124),
.B(n_96),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_159),
.B(n_170),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_114),
.A2(n_107),
.B1(n_97),
.B2(n_84),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_115),
.A2(n_20),
.B1(n_21),
.B2(n_22),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_161),
.A2(n_169),
.B1(n_176),
.B2(n_27),
.Y(n_181)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_117),
.Y(n_162)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_162),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_164),
.B(n_167),
.Y(n_178)
);

AO22x1_ASAP7_75t_L g166 ( 
.A1(n_115),
.A2(n_89),
.B1(n_106),
.B2(n_77),
.Y(n_166)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_166),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_114),
.A2(n_11),
.B1(n_15),
.B2(n_14),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_125),
.B(n_118),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_171),
.B(n_130),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_139),
.A2(n_21),
.B1(n_29),
.B2(n_32),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_172),
.A2(n_141),
.B1(n_133),
.B2(n_140),
.Y(n_183)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_117),
.Y(n_173)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_173),
.Y(n_201)
);

BUFx6f_ASAP7_75t_L g174 ( 
.A(n_126),
.Y(n_174)
);

INVx4_ASAP7_75t_L g180 ( 
.A(n_174),
.Y(n_180)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_126),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_175),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_114),
.A2(n_11),
.B1(n_15),
.B2(n_14),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_SL g213 ( 
.A1(n_179),
.A2(n_184),
.B(n_191),
.Y(n_213)
);

AOI22xp33_ASAP7_75t_L g218 ( 
.A1(n_181),
.A2(n_183),
.B1(n_200),
.B2(n_172),
.Y(n_218)
);

OAI21xp5_ASAP7_75t_SL g184 ( 
.A1(n_152),
.A2(n_149),
.B(n_148),
.Y(n_184)
);

INVxp67_ASAP7_75t_L g186 ( 
.A(n_160),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_186),
.B(n_199),
.Y(n_212)
);

NOR2x1_ASAP7_75t_L g189 ( 
.A(n_144),
.B(n_128),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_SL g232 ( 
.A(n_189),
.B(n_210),
.Y(n_232)
);

OAI21xp5_ASAP7_75t_SL g191 ( 
.A1(n_166),
.A2(n_132),
.B(n_113),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_SL g192 ( 
.A1(n_166),
.A2(n_113),
.B(n_138),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_SL g214 ( 
.A1(n_192),
.A2(n_206),
.B(n_169),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_143),
.A2(n_122),
.B1(n_141),
.B2(n_138),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g211 ( 
.A1(n_193),
.A2(n_205),
.B1(n_153),
.B2(n_176),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g195 ( 
.A(n_171),
.B(n_127),
.Y(n_195)
);

AOI21xp5_ASAP7_75t_L g223 ( 
.A1(n_195),
.A2(n_196),
.B(n_203),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_145),
.B(n_125),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_162),
.A2(n_141),
.B1(n_121),
.B2(n_129),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_L g230 ( 
.A1(n_198),
.A2(n_190),
.B(n_194),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_165),
.B(n_142),
.Y(n_199)
);

AOI22xp33_ASAP7_75t_L g200 ( 
.A1(n_168),
.A2(n_120),
.B1(n_136),
.B2(n_123),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_154),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_202),
.B(n_174),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g203 ( 
.A(n_145),
.B(n_136),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_143),
.A2(n_119),
.B1(n_32),
.B2(n_29),
.Y(n_205)
);

AOI32xp33_ASAP7_75t_L g206 ( 
.A1(n_147),
.A2(n_25),
.A3(n_16),
.B1(n_32),
.B2(n_29),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_159),
.B(n_25),
.C(n_13),
.Y(n_207)
);

INVxp67_ASAP7_75t_L g236 ( 
.A(n_207),
.Y(n_236)
);

AO22x1_ASAP7_75t_SL g209 ( 
.A1(n_161),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_209)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_209),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g210 ( 
.A(n_147),
.B(n_13),
.Y(n_210)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_210),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_211),
.A2(n_216),
.B1(n_227),
.B2(n_180),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_214),
.B(n_182),
.Y(n_245)
);

INVx1_ASAP7_75t_SL g215 ( 
.A(n_198),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_215),
.B(n_217),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_L g216 ( 
.A1(n_208),
.A2(n_173),
.B1(n_163),
.B2(n_165),
.Y(n_216)
);

INVx1_ASAP7_75t_SL g217 ( 
.A(n_188),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_218),
.A2(n_205),
.B1(n_201),
.B2(n_207),
.Y(n_239)
);

CKINVDCx16_ASAP7_75t_R g219 ( 
.A(n_177),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_219),
.B(n_220),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_185),
.Y(n_220)
);

AOI22xp33_ASAP7_75t_SL g221 ( 
.A1(n_208),
.A2(n_156),
.B1(n_151),
.B2(n_146),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_L g246 ( 
.A1(n_221),
.A2(n_222),
.B1(n_225),
.B2(n_209),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_204),
.A2(n_158),
.B1(n_157),
.B2(n_151),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_186),
.A2(n_189),
.B1(n_184),
.B2(n_193),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_185),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_226),
.B(n_234),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_L g227 ( 
.A1(n_183),
.A2(n_150),
.B1(n_175),
.B2(n_170),
.Y(n_227)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_229),
.Y(n_244)
);

OAI21xp5_ASAP7_75t_L g243 ( 
.A1(n_230),
.A2(n_232),
.B(n_187),
.Y(n_243)
);

HB1xp67_ASAP7_75t_L g231 ( 
.A(n_190),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_231),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_SL g233 ( 
.A(n_197),
.B(n_164),
.Y(n_233)
);

CKINVDCx14_ASAP7_75t_R g242 ( 
.A(n_233),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_SL g234 ( 
.A(n_197),
.B(n_174),
.Y(n_234)
);

CKINVDCx16_ASAP7_75t_R g235 ( 
.A(n_178),
.Y(n_235)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_235),
.Y(n_250)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_201),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_237),
.B(n_238),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_187),
.Y(n_238)
);

AOI22xp33_ASAP7_75t_L g281 ( 
.A1(n_239),
.A2(n_246),
.B1(n_252),
.B2(n_254),
.Y(n_281)
);

AO22x1_ASAP7_75t_L g240 ( 
.A1(n_215),
.A2(n_182),
.B1(n_192),
.B2(n_191),
.Y(n_240)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_240),
.Y(n_264)
);

NAND3xp33_ASAP7_75t_L g241 ( 
.A(n_217),
.B(n_212),
.C(n_238),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_241),
.B(n_261),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g265 ( 
.A(n_243),
.B(n_227),
.Y(n_265)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_245),
.B(n_263),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_L g247 ( 
.A1(n_225),
.A2(n_209),
.B1(n_181),
.B2(n_179),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_247),
.A2(n_258),
.B1(n_236),
.B2(n_219),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_223),
.B(n_195),
.C(n_213),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_249),
.B(n_251),
.C(n_256),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_223),
.B(n_196),
.C(n_203),
.Y(n_251)
);

OAI21xp5_ASAP7_75t_L g252 ( 
.A1(n_230),
.A2(n_212),
.B(n_232),
.Y(n_252)
);

OAI21xp5_ASAP7_75t_L g254 ( 
.A1(n_224),
.A2(n_180),
.B(n_11),
.Y(n_254)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_255),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_213),
.B(n_2),
.C(n_3),
.Y(n_256)
);

NAND2x1_ASAP7_75t_SL g257 ( 
.A(n_234),
.B(n_3),
.Y(n_257)
);

CKINVDCx16_ASAP7_75t_R g268 ( 
.A(n_257),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_L g258 ( 
.A1(n_222),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_216),
.B(n_5),
.Y(n_261)
);

XOR2xp5_ASAP7_75t_L g263 ( 
.A(n_214),
.B(n_5),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_L g288 ( 
.A(n_265),
.B(n_263),
.Y(n_288)
);

INVxp33_ASAP7_75t_SL g266 ( 
.A(n_260),
.Y(n_266)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_266),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_253),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_270),
.B(n_271),
.Y(n_291)
);

INVxp67_ASAP7_75t_L g271 ( 
.A(n_259),
.Y(n_271)
);

NOR2x1_ASAP7_75t_L g272 ( 
.A(n_242),
.B(n_224),
.Y(n_272)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_272),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_251),
.B(n_228),
.C(n_211),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_275),
.B(n_276),
.C(n_278),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_249),
.B(n_228),
.C(n_226),
.Y(n_276)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_277),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_253),
.B(n_220),
.C(n_233),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_245),
.B(n_229),
.C(n_235),
.Y(n_279)
);

HB1xp67_ASAP7_75t_L g295 ( 
.A(n_279),
.Y(n_295)
);

HB1xp67_ASAP7_75t_L g280 ( 
.A(n_244),
.Y(n_280)
);

BUFx2_ASAP7_75t_L g297 ( 
.A(n_280),
.Y(n_297)
);

AND2x2_ASAP7_75t_L g282 ( 
.A(n_244),
.B(n_231),
.Y(n_282)
);

INVxp67_ASAP7_75t_L g286 ( 
.A(n_282),
.Y(n_286)
);

INVxp67_ASAP7_75t_L g283 ( 
.A(n_255),
.Y(n_283)
);

OAI22xp33_ASAP7_75t_SL g292 ( 
.A1(n_283),
.A2(n_262),
.B1(n_254),
.B2(n_257),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_283),
.A2(n_267),
.B1(n_264),
.B2(n_282),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_285),
.A2(n_268),
.B1(n_248),
.B2(n_273),
.Y(n_307)
);

XOR2xp5_ASAP7_75t_L g309 ( 
.A(n_288),
.B(n_293),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_278),
.B(n_250),
.Y(n_289)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_289),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_292),
.B(n_296),
.Y(n_301)
);

XOR2xp5_ASAP7_75t_L g293 ( 
.A(n_274),
.B(n_243),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_L g294 ( 
.A(n_275),
.B(n_252),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_294),
.B(n_269),
.C(n_256),
.Y(n_302)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_272),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_271),
.B(n_250),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_298),
.B(n_262),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_299),
.B(n_276),
.C(n_279),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_SL g323 ( 
.A(n_300),
.B(n_307),
.Y(n_323)
);

XNOR2xp5_ASAP7_75t_L g321 ( 
.A(n_302),
.B(n_313),
.Y(n_321)
);

XNOR2x1_ASAP7_75t_L g303 ( 
.A(n_286),
.B(n_281),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_SL g318 ( 
.A(n_303),
.B(n_305),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_299),
.B(n_294),
.C(n_269),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_304),
.B(n_240),
.Y(n_316)
);

MAJx2_ASAP7_75t_L g305 ( 
.A(n_293),
.B(n_274),
.C(n_240),
.Y(n_305)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_306),
.Y(n_315)
);

AOI21xp5_ASAP7_75t_SL g308 ( 
.A1(n_287),
.A2(n_290),
.B(n_291),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_L g319 ( 
.A1(n_308),
.A2(n_257),
.B1(n_297),
.B2(n_7),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_288),
.B(n_239),
.C(n_261),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_310),
.B(n_6),
.Y(n_322)
);

XOR2xp5_ASAP7_75t_L g311 ( 
.A(n_285),
.B(n_248),
.Y(n_311)
);

XOR2xp5_ASAP7_75t_L g320 ( 
.A(n_311),
.B(n_5),
.Y(n_320)
);

HB1xp67_ASAP7_75t_L g313 ( 
.A(n_284),
.Y(n_313)
);

AND2x2_ASAP7_75t_L g314 ( 
.A(n_303),
.B(n_286),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_SL g327 ( 
.A(n_314),
.B(n_319),
.Y(n_327)
);

AOI21xp5_ASAP7_75t_L g330 ( 
.A1(n_316),
.A2(n_322),
.B(n_6),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_L g317 ( 
.A1(n_301),
.A2(n_295),
.B1(n_237),
.B2(n_297),
.Y(n_317)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_317),
.Y(n_328)
);

XNOR2xp5_ASAP7_75t_L g329 ( 
.A(n_320),
.B(n_309),
.Y(n_329)
);

AOI21xp5_ASAP7_75t_SL g324 ( 
.A1(n_323),
.A2(n_308),
.B(n_312),
.Y(n_324)
);

OAI21xp5_ASAP7_75t_SL g336 ( 
.A1(n_324),
.A2(n_318),
.B(n_9),
.Y(n_336)
);

AOI22xp5_ASAP7_75t_SL g325 ( 
.A1(n_315),
.A2(n_305),
.B1(n_300),
.B2(n_309),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_325),
.B(n_330),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_321),
.B(n_311),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_SL g333 ( 
.A(n_326),
.B(n_329),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_320),
.B(n_6),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_SL g335 ( 
.A(n_331),
.B(n_7),
.Y(n_335)
);

AOI21xp5_ASAP7_75t_L g334 ( 
.A1(n_328),
.A2(n_314),
.B(n_318),
.Y(n_334)
);

MAJx2_ASAP7_75t_L g337 ( 
.A(n_334),
.B(n_336),
.C(n_327),
.Y(n_337)
);

AOI22xp33_ASAP7_75t_SL g338 ( 
.A1(n_335),
.A2(n_327),
.B1(n_9),
.B2(n_10),
.Y(n_338)
);

OAI21xp5_ASAP7_75t_L g339 ( 
.A1(n_337),
.A2(n_338),
.B(n_332),
.Y(n_339)
);

CKINVDCx20_ASAP7_75t_R g340 ( 
.A(n_339),
.Y(n_340)
);

OAI21xp5_ASAP7_75t_L g341 ( 
.A1(n_340),
.A2(n_333),
.B(n_7),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_L g342 ( 
.A(n_341),
.B(n_7),
.Y(n_342)
);

NAND3xp33_ASAP7_75t_SL g343 ( 
.A(n_342),
.B(n_10),
.C(n_339),
.Y(n_343)
);


endmodule