module real_jpeg_16501_n_10 (n_5, n_4, n_8, n_0, n_1, n_2, n_6, n_7, n_3, n_9, n_10);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_2;
input n_6;
input n_7;
input n_3;
input n_9;

output n_10;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_247;
wire n_146;
wire n_78;
wire n_83;
wire n_249;
wire n_166;
wire n_176;
wire n_215;
wire n_221;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_11;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_243;
wire n_255;
wire n_115;
wire n_98;
wire n_27;
wire n_184;
wire n_56;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_13;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_141;
wire n_95;
wire n_242;
wire n_65;
wire n_33;
wire n_188;
wire n_139;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_172;
wire n_160;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_262;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_205;
wire n_258;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_241;
wire n_103;
wire n_259;
wire n_225;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_185;
wire n_240;
wire n_209;
wire n_55;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_12;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_167;
wire n_216;
wire n_128;
wire n_179;
wire n_202;
wire n_213;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_256;
wire n_182;
wire n_253;
wire n_96;
wire n_89;
wire n_16;

OAI32xp33_ASAP7_75t_L g16 ( 
.A1(n_0),
.A2(n_17),
.A3(n_20),
.B1(n_23),
.B2(n_29),
.Y(n_16)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_L g37 ( 
.A1(n_0),
.A2(n_38),
.B1(n_39),
.B2(n_41),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_0),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_0),
.A2(n_74),
.B1(n_76),
.B2(n_77),
.Y(n_73)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_0),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_0),
.B(n_132),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_0),
.B(n_167),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_0),
.B(n_197),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_0),
.A2(n_176),
.B1(n_224),
.B2(n_227),
.Y(n_223)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_1),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_L g80 ( 
.A1(n_2),
.A2(n_81),
.B1(n_84),
.B2(n_85),
.Y(n_80)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_2),
.Y(n_84)
);

OAI22xp33_ASAP7_75t_L g111 ( 
.A1(n_2),
.A2(n_84),
.B1(n_112),
.B2(n_115),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_2),
.A2(n_84),
.B1(n_125),
.B2(n_127),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_2),
.A2(n_84),
.B1(n_232),
.B2(n_241),
.Y(n_240)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_3),
.Y(n_102)
);

BUFx5_ASAP7_75t_L g103 ( 
.A(n_3),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_3),
.Y(n_110)
);

BUFx5_ASAP7_75t_L g147 ( 
.A(n_3),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g150 ( 
.A(n_3),
.Y(n_150)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_4),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_4),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g68 ( 
.A(n_5),
.Y(n_68)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_5),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_5),
.Y(n_100)
);

BUFx3_ASAP7_75t_L g105 ( 
.A(n_5),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g201 ( 
.A(n_6),
.Y(n_201)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_6),
.Y(n_204)
);

INVx6_ASAP7_75t_L g235 ( 
.A(n_6),
.Y(n_235)
);

BUFx5_ASAP7_75t_L g238 ( 
.A(n_6),
.Y(n_238)
);

BUFx6f_ASAP7_75t_L g251 ( 
.A(n_6),
.Y(n_251)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_7),
.Y(n_66)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_8),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_8),
.Y(n_43)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_8),
.Y(n_108)
);

BUFx3_ASAP7_75t_L g226 ( 
.A(n_9),
.Y(n_226)
);

BUFx8_ASAP7_75t_L g229 ( 
.A(n_9),
.Y(n_229)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_9),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g10 ( 
.A(n_11),
.B(n_209),
.Y(n_10)
);

AOI21x1_ASAP7_75t_L g11 ( 
.A1(n_12),
.A2(n_185),
.B(n_208),
.Y(n_11)
);

OAI21x1_ASAP7_75t_L g12 ( 
.A1(n_13),
.A2(n_133),
.B(n_184),
.Y(n_12)
);

NOR2xp67_ASAP7_75t_SL g13 ( 
.A(n_14),
.B(n_119),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_14),
.B(n_119),
.Y(n_184)
);

XOR2x2_ASAP7_75t_SL g14 ( 
.A(n_15),
.B(n_56),
.Y(n_14)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_15),
.B(n_88),
.C(n_117),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_35),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_16),
.B(n_35),
.Y(n_188)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_18),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_19),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_19),
.Y(n_87)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

INVx4_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_SL g23 ( 
.A(n_24),
.B(n_28),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_27),
.Y(n_92)
);

BUFx3_ASAP7_75t_L g95 ( 
.A(n_27),
.Y(n_95)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_27),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_28),
.B(n_94),
.Y(n_93)
);

BUFx2_ASAP7_75t_L g176 ( 
.A(n_28),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_29),
.B(n_60),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_30),
.B(n_33),
.Y(n_29)
);

OA22x2_ASAP7_75t_L g67 ( 
.A1(n_30),
.A2(n_68),
.B1(n_69),
.B2(n_71),
.Y(n_67)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_34),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_36),
.B(n_44),
.Y(n_35)
);

OA22x2_ASAP7_75t_L g122 ( 
.A1(n_36),
.A2(n_123),
.B1(n_124),
.B2(n_129),
.Y(n_122)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_37),
.B(n_45),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_L g89 ( 
.A1(n_38),
.A2(n_90),
.B(n_93),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

AO22x2_ASAP7_75t_L g106 ( 
.A1(n_40),
.A2(n_102),
.B1(n_107),
.B2(n_109),
.Y(n_106)
);

BUFx3_ASAP7_75t_L g126 ( 
.A(n_40),
.Y(n_126)
);

INVx4_ASAP7_75t_L g128 ( 
.A(n_40),
.Y(n_128)
);

INVx3_ASAP7_75t_L g165 ( 
.A(n_40),
.Y(n_165)
);

HB1xp67_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_43),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g153 ( 
.A(n_43),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_SL g44 ( 
.A(n_45),
.B(n_51),
.Y(n_44)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_45),
.Y(n_123)
);

AND2x2_ASAP7_75t_L g45 ( 
.A(n_46),
.B(n_49),
.Y(n_45)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_47),
.Y(n_130)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_48),
.Y(n_170)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_49),
.Y(n_142)
);

INVx5_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

OA21x2_ASAP7_75t_L g171 ( 
.A1(n_52),
.A2(n_124),
.B(n_172),
.Y(n_171)
);

INVx5_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_SL g56 ( 
.A1(n_57),
.A2(n_88),
.B1(n_117),
.B2(n_118),
.Y(n_56)
);

INVx2_ASAP7_75t_SL g117 ( 
.A(n_57),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g215 ( 
.A1(n_57),
.A2(n_117),
.B1(n_216),
.B2(n_217),
.Y(n_215)
);

OA22x2_ASAP7_75t_L g57 ( 
.A1(n_58),
.A2(n_67),
.B1(n_73),
.B2(n_80),
.Y(n_57)
);

OA22x2_ASAP7_75t_L g192 ( 
.A1(n_58),
.A2(n_67),
.B1(n_73),
.B2(n_80),
.Y(n_192)
);

NAND2x1p5_ASAP7_75t_L g58 ( 
.A(n_59),
.B(n_67),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_61),
.B(n_64),
.Y(n_60)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_63),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g202 ( 
.A(n_65),
.Y(n_202)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

BUFx5_ASAP7_75t_L g79 ( 
.A(n_66),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_66),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g199 ( 
.A(n_66),
.Y(n_199)
);

BUFx6f_ASAP7_75t_L g257 ( 
.A(n_66),
.Y(n_257)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_67),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_70),
.Y(n_114)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx2_ASAP7_75t_SL g78 ( 
.A(n_79),
.Y(n_78)
);

BUFx2_ASAP7_75t_SL g81 ( 
.A(n_82),
.Y(n_81)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx6_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx6_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g262 ( 
.A(n_87),
.Y(n_262)
);

INVx1_ASAP7_75t_SL g118 ( 
.A(n_88),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_88),
.B(n_136),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_88),
.A2(n_118),
.B1(n_136),
.B2(n_181),
.Y(n_180)
);

AO22x2_ASAP7_75t_L g88 ( 
.A1(n_89),
.A2(n_96),
.B1(n_106),
.B2(n_111),
.Y(n_88)
);

AO22x1_ASAP7_75t_L g121 ( 
.A1(n_89),
.A2(n_96),
.B1(n_106),
.B2(n_111),
.Y(n_121)
);

INVxp67_ASAP7_75t_L g220 ( 
.A(n_89),
.Y(n_220)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVx5_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

OAI32xp33_ASAP7_75t_L g136 ( 
.A1(n_93),
.A2(n_137),
.A3(n_141),
.B1(n_143),
.B2(n_148),
.Y(n_136)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_96),
.Y(n_218)
);

NOR2x1p5_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_106),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_98),
.A2(n_101),
.B1(n_103),
.B2(n_104),
.Y(n_97)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVx6_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_100),
.Y(n_140)
);

INVx8_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx5_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_106),
.B(n_175),
.Y(n_174)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_106),
.Y(n_219)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx6_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_120),
.B(n_122),
.C(n_131),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_120),
.A2(n_121),
.B1(n_188),
.B2(n_189),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_120),
.B(n_188),
.C(n_190),
.Y(n_212)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

XNOR2xp5_ASAP7_75t_L g157 ( 
.A(n_121),
.B(n_131),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_122),
.A2(n_155),
.B1(n_156),
.B2(n_157),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_122),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_122),
.B(n_174),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_122),
.B(n_174),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_L g246 ( 
.A1(n_122),
.A2(n_155),
.B1(n_247),
.B2(n_248),
.Y(n_246)
);

INVx3_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

AOI21x1_ASAP7_75t_L g133 ( 
.A1(n_134),
.A2(n_158),
.B(n_183),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_135),
.B(n_154),
.Y(n_134)
);

NOR2xp67_ASAP7_75t_SL g183 ( 
.A(n_135),
.B(n_154),
.Y(n_183)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_136),
.Y(n_181)
);

INVx4_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

INVx5_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

INVx1_ASAP7_75t_SL g143 ( 
.A(n_144),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_151),
.Y(n_148)
);

INVx6_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

BUFx3_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

OAI21x1_ASAP7_75t_L g158 ( 
.A1(n_159),
.A2(n_178),
.B(n_182),
.Y(n_158)
);

AOI21xp5_ASAP7_75t_SL g159 ( 
.A1(n_160),
.A2(n_173),
.B(n_177),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_161),
.B(n_171),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_162),
.B(n_166),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

INVx3_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_171),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_171),
.A2(n_179),
.B1(n_195),
.B2(n_196),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_171),
.B(n_192),
.C(n_196),
.Y(n_245)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g258 ( 
.A(n_176),
.B(n_259),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_180),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_179),
.B(n_180),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_186),
.B(n_207),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_186),
.B(n_207),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_187),
.A2(n_190),
.B1(n_191),
.B2(n_206),
.Y(n_186)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_187),
.Y(n_206)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_188),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_192),
.A2(n_193),
.B1(n_194),
.B2(n_205),
.Y(n_191)
);

INVx1_ASAP7_75t_SL g205 ( 
.A(n_192),
.Y(n_205)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

INVxp67_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

OA22x2_ASAP7_75t_L g222 ( 
.A1(n_198),
.A2(n_223),
.B1(n_230),
.B2(n_240),
.Y(n_222)
);

OAI21x1_ASAP7_75t_L g230 ( 
.A1(n_198),
.A2(n_231),
.B(n_236),
.Y(n_230)
);

OA22x2_ASAP7_75t_L g198 ( 
.A1(n_199),
.A2(n_200),
.B1(n_202),
.B2(n_203),
.Y(n_198)
);

INVx6_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_210),
.B(n_263),
.Y(n_209)
);

INVxp67_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_212),
.B(n_213),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_212),
.B(n_213),
.Y(n_263)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_214),
.B(n_244),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_SL g214 ( 
.A(n_215),
.B(n_221),
.Y(n_214)
);

INVxp67_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

AOI21xp5_ASAP7_75t_L g217 ( 
.A1(n_218),
.A2(n_219),
.B(n_220),
.Y(n_217)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

INVx3_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

BUFx6f_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

BUFx12f_ASAP7_75t_L g232 ( 
.A(n_226),
.Y(n_232)
);

BUFx6f_ASAP7_75t_L g239 ( 
.A(n_226),
.Y(n_239)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

INVx3_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

INVxp67_ASAP7_75t_L g261 ( 
.A(n_231),
.Y(n_261)
);

AND2x2_ASAP7_75t_L g231 ( 
.A(n_232),
.B(n_233),
.Y(n_231)
);

INVx3_ASAP7_75t_L g260 ( 
.A(n_232),
.Y(n_260)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

INVx3_ASAP7_75t_SL g234 ( 
.A(n_235),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_237),
.B(n_239),
.Y(n_236)
);

INVx4_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

HB1xp67_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

BUFx6f_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_SL g244 ( 
.A(n_245),
.B(n_246),
.Y(n_244)
);

INVx1_ASAP7_75t_SL g247 ( 
.A(n_248),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_249),
.A2(n_258),
.B1(n_261),
.B2(n_262),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_250),
.B(n_252),
.Y(n_249)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

INVx1_ASAP7_75t_SL g252 ( 
.A(n_253),
.Y(n_252)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

INVx3_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);


endmodule