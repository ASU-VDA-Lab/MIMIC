module fake_jpeg_12731_n_433 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_433);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_433;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_430;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_9),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

BUFx12_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_9),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

BUFx12_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_8),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

INVx13_ASAP7_75t_L g32 ( 
.A(n_16),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_4),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_13),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_10),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_11),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_11),
.Y(n_37)
);

INVx5_ASAP7_75t_L g38 ( 
.A(n_4),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_0),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_7),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_16),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_14),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_7),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_8),
.Y(n_44)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_3),
.Y(n_45)
);

BUFx16f_ASAP7_75t_L g46 ( 
.A(n_16),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_4),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_2),
.Y(n_48)
);

BUFx2_ASAP7_75t_L g49 ( 
.A(n_15),
.Y(n_49)
);

BUFx5_ASAP7_75t_L g50 ( 
.A(n_2),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_8),
.Y(n_51)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_14),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_5),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_18),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_54),
.Y(n_113)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_22),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g122 ( 
.A(n_55),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_18),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_56),
.Y(n_131)
);

BUFx5_ASAP7_75t_L g57 ( 
.A(n_22),
.Y(n_57)
);

BUFx5_ASAP7_75t_L g139 ( 
.A(n_57),
.Y(n_139)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_50),
.Y(n_58)
);

INVx5_ASAP7_75t_L g170 ( 
.A(n_58),
.Y(n_170)
);

INVx5_ASAP7_75t_L g59 ( 
.A(n_23),
.Y(n_59)
);

INVx3_ASAP7_75t_L g164 ( 
.A(n_59),
.Y(n_164)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_46),
.Y(n_60)
);

INVx4_ASAP7_75t_L g116 ( 
.A(n_60),
.Y(n_116)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_20),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_61),
.Y(n_132)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_52),
.Y(n_62)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_62),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_18),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g138 ( 
.A(n_63),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_31),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_64),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_17),
.B(n_15),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g171 ( 
.A(n_65),
.B(n_88),
.Y(n_171)
);

INVx8_ASAP7_75t_L g66 ( 
.A(n_50),
.Y(n_66)
);

INVx5_ASAP7_75t_L g175 ( 
.A(n_66),
.Y(n_175)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_49),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_67),
.A2(n_53),
.B1(n_48),
.B2(n_39),
.Y(n_118)
);

HB1xp67_ASAP7_75t_L g68 ( 
.A(n_38),
.Y(n_68)
);

CKINVDCx16_ASAP7_75t_R g153 ( 
.A(n_68),
.Y(n_153)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_52),
.Y(n_69)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_69),
.Y(n_133)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_31),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g147 ( 
.A(n_70),
.Y(n_147)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_23),
.Y(n_71)
);

BUFx3_ASAP7_75t_L g143 ( 
.A(n_71),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_31),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g149 ( 
.A(n_72),
.Y(n_149)
);

INVx11_ASAP7_75t_L g73 ( 
.A(n_32),
.Y(n_73)
);

INVx11_ASAP7_75t_L g167 ( 
.A(n_73),
.Y(n_167)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_23),
.Y(n_74)
);

INVx4_ASAP7_75t_L g146 ( 
.A(n_74),
.Y(n_146)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_49),
.Y(n_75)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_75),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_33),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g161 ( 
.A(n_76),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_33),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g165 ( 
.A(n_77),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_33),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g172 ( 
.A(n_78),
.Y(n_172)
);

INVx3_ASAP7_75t_SL g79 ( 
.A(n_45),
.Y(n_79)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_79),
.Y(n_140)
);

INVx13_ASAP7_75t_L g80 ( 
.A(n_32),
.Y(n_80)
);

INVx13_ASAP7_75t_L g128 ( 
.A(n_80),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_45),
.Y(n_81)
);

INVx8_ASAP7_75t_L g126 ( 
.A(n_81),
.Y(n_126)
);

BUFx12f_ASAP7_75t_L g82 ( 
.A(n_51),
.Y(n_82)
);

BUFx3_ASAP7_75t_L g154 ( 
.A(n_82),
.Y(n_154)
);

INVx8_ASAP7_75t_L g83 ( 
.A(n_20),
.Y(n_83)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_83),
.Y(n_119)
);

BUFx2_ASAP7_75t_L g84 ( 
.A(n_38),
.Y(n_84)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_84),
.Y(n_156)
);

BUFx3_ASAP7_75t_L g85 ( 
.A(n_23),
.Y(n_85)
);

BUFx12f_ASAP7_75t_L g114 ( 
.A(n_85),
.Y(n_114)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_46),
.Y(n_86)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_86),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_45),
.Y(n_87)
);

INVx8_ASAP7_75t_L g155 ( 
.A(n_87),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_17),
.B(n_15),
.Y(n_88)
);

CKINVDCx16_ASAP7_75t_R g89 ( 
.A(n_32),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_89),
.B(n_101),
.Y(n_112)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_27),
.Y(n_90)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_90),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_20),
.Y(n_91)
);

BUFx12f_ASAP7_75t_L g150 ( 
.A(n_91),
.Y(n_150)
);

BUFx12f_ASAP7_75t_L g92 ( 
.A(n_51),
.Y(n_92)
);

BUFx4f_ASAP7_75t_SL g111 ( 
.A(n_92),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_29),
.Y(n_93)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_93),
.Y(n_176)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_46),
.Y(n_94)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_94),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_26),
.B(n_14),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_95),
.B(n_107),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_29),
.Y(n_96)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_96),
.Y(n_163)
);

INVx8_ASAP7_75t_L g97 ( 
.A(n_29),
.Y(n_97)
);

BUFx4f_ASAP7_75t_SL g159 ( 
.A(n_97),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_26),
.B(n_10),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_98),
.B(n_100),
.Y(n_127)
);

AND2x2_ASAP7_75t_L g99 ( 
.A(n_49),
.B(n_41),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g174 ( 
.A(n_99),
.B(n_102),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_34),
.B(n_10),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_34),
.B(n_0),
.Y(n_101)
);

BUFx5_ASAP7_75t_L g102 ( 
.A(n_19),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_24),
.Y(n_103)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_103),
.Y(n_168)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_24),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_104),
.B(n_106),
.Y(n_115)
);

INVx8_ASAP7_75t_L g105 ( 
.A(n_25),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_105),
.B(n_47),
.Y(n_152)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_27),
.Y(n_106)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_19),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_24),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_108),
.B(n_41),
.Y(n_125)
);

INVx11_ASAP7_75t_L g109 ( 
.A(n_25),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_109),
.Y(n_166)
);

INVx5_ASAP7_75t_L g110 ( 
.A(n_24),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_110),
.B(n_41),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_118),
.A2(n_80),
.B1(n_63),
.B2(n_78),
.Y(n_189)
);

OA22x2_ASAP7_75t_L g120 ( 
.A1(n_81),
.A2(n_53),
.B1(n_48),
.B2(n_39),
.Y(n_120)
);

OA22x2_ASAP7_75t_L g206 ( 
.A1(n_120),
.A2(n_28),
.B1(n_6),
.B2(n_8),
.Y(n_206)
);

INVxp67_ASAP7_75t_L g179 ( 
.A(n_121),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_65),
.B(n_37),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_SL g203 ( 
.A(n_123),
.B(n_141),
.Y(n_203)
);

AND2x2_ASAP7_75t_L g225 ( 
.A(n_125),
.B(n_152),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_88),
.B(n_37),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_130),
.B(n_148),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_98),
.A2(n_21),
.B1(n_35),
.B2(n_36),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_135),
.A2(n_151),
.B1(n_177),
.B2(n_79),
.Y(n_181)
);

AOI22xp33_ASAP7_75t_L g136 ( 
.A1(n_91),
.A2(n_47),
.B1(n_44),
.B2(n_43),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g215 ( 
.A1(n_136),
.A2(n_162),
.B1(n_157),
.B2(n_119),
.Y(n_215)
);

AOI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_58),
.A2(n_66),
.B1(n_84),
.B2(n_21),
.Y(n_137)
);

AOI21xp5_ASAP7_75t_L g184 ( 
.A1(n_137),
.A2(n_145),
.B(n_157),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_100),
.B(n_36),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_SL g145 ( 
.A1(n_68),
.A2(n_41),
.B1(n_44),
.B2(n_43),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_82),
.B(n_35),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_67),
.A2(n_42),
.B1(n_30),
.B2(n_40),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_SL g157 ( 
.A1(n_55),
.A2(n_40),
.B1(n_42),
.B2(n_30),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_99),
.B(n_0),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_160),
.B(n_5),
.Y(n_194)
);

AOI22xp33_ASAP7_75t_SL g162 ( 
.A1(n_70),
.A2(n_1),
.B1(n_3),
.B2(n_5),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_92),
.B(n_1),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_169),
.B(n_173),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_105),
.B(n_3),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_93),
.A2(n_28),
.B1(n_25),
.B2(n_7),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_103),
.B(n_5),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_178),
.B(n_6),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_115),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_180),
.B(n_187),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_L g259 ( 
.A1(n_181),
.A2(n_189),
.B1(n_212),
.B2(n_138),
.Y(n_259)
);

INVxp67_ASAP7_75t_L g182 ( 
.A(n_167),
.Y(n_182)
);

HB1xp67_ASAP7_75t_L g273 ( 
.A(n_182),
.Y(n_273)
);

INVx4_ASAP7_75t_L g183 ( 
.A(n_150),
.Y(n_183)
);

INVx3_ASAP7_75t_L g263 ( 
.A(n_183),
.Y(n_263)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_140),
.Y(n_185)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_185),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_124),
.B(n_108),
.C(n_87),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_186),
.B(n_205),
.Y(n_251)
);

INVxp67_ASAP7_75t_L g187 ( 
.A(n_167),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_117),
.Y(n_188)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_188),
.Y(n_246)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_142),
.Y(n_190)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_190),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_163),
.A2(n_96),
.B1(n_54),
.B2(n_56),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_191),
.A2(n_192),
.B1(n_144),
.B2(n_149),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_120),
.A2(n_77),
.B1(n_76),
.B2(n_72),
.Y(n_192)
);

AOI22xp33_ASAP7_75t_SL g193 ( 
.A1(n_170),
.A2(n_64),
.B1(n_25),
.B2(n_28),
.Y(n_193)
);

INVxp67_ASAP7_75t_L g250 ( 
.A(n_193),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_SL g244 ( 
.A(n_194),
.B(n_208),
.Y(n_244)
);

BUFx6f_ASAP7_75t_L g195 ( 
.A(n_113),
.Y(n_195)
);

BUFx6f_ASAP7_75t_L g241 ( 
.A(n_195),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_127),
.B(n_6),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_196),
.B(n_217),
.Y(n_240)
);

AOI22xp33_ASAP7_75t_SL g197 ( 
.A1(n_170),
.A2(n_175),
.B1(n_156),
.B2(n_137),
.Y(n_197)
);

AOI22xp33_ASAP7_75t_SL g236 ( 
.A1(n_197),
.A2(n_211),
.B1(n_143),
.B2(n_126),
.Y(n_236)
);

INVxp33_ASAP7_75t_L g198 ( 
.A(n_128),
.Y(n_198)
);

NAND2xp33_ASAP7_75t_SL g239 ( 
.A(n_198),
.B(n_223),
.Y(n_239)
);

BUFx3_ASAP7_75t_L g199 ( 
.A(n_114),
.Y(n_199)
);

INVx1_ASAP7_75t_SL g267 ( 
.A(n_199),
.Y(n_267)
);

BUFx6f_ASAP7_75t_L g200 ( 
.A(n_113),
.Y(n_200)
);

INVx6_ASAP7_75t_L g270 ( 
.A(n_200),
.Y(n_270)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_168),
.Y(n_202)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_202),
.Y(n_276)
);

INVx8_ASAP7_75t_L g204 ( 
.A(n_147),
.Y(n_204)
);

INVx3_ASAP7_75t_SL g278 ( 
.A(n_204),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_174),
.B(n_28),
.C(n_7),
.Y(n_205)
);

AND2x2_ASAP7_75t_L g242 ( 
.A(n_206),
.B(n_221),
.Y(n_242)
);

INVx4_ASAP7_75t_L g207 ( 
.A(n_150),
.Y(n_207)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_207),
.Y(n_245)
);

INVx6_ASAP7_75t_L g210 ( 
.A(n_131),
.Y(n_210)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_210),
.Y(n_248)
);

AOI22xp33_ASAP7_75t_SL g211 ( 
.A1(n_175),
.A2(n_122),
.B1(n_154),
.B2(n_145),
.Y(n_211)
);

AOI22xp33_ASAP7_75t_L g212 ( 
.A1(n_120),
.A2(n_174),
.B1(n_136),
.B2(n_153),
.Y(n_212)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_176),
.Y(n_213)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_213),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_128),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_214),
.B(n_216),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_215),
.A2(n_222),
.B1(n_149),
.B2(n_131),
.Y(n_238)
);

CKINVDCx16_ASAP7_75t_R g216 ( 
.A(n_111),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_129),
.B(n_133),
.Y(n_217)
);

CKINVDCx16_ASAP7_75t_R g218 ( 
.A(n_111),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_218),
.B(n_226),
.Y(n_256)
);

O2A1O1Ixp33_ASAP7_75t_L g219 ( 
.A1(n_119),
.A2(n_112),
.B(n_162),
.C(n_159),
.Y(n_219)
);

A2O1A1Ixp33_ASAP7_75t_L g271 ( 
.A1(n_219),
.A2(n_205),
.B(n_179),
.C(n_220),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_171),
.A2(n_143),
.B1(n_122),
.B2(n_154),
.Y(n_220)
);

AOI21xp5_ASAP7_75t_L g274 ( 
.A1(n_220),
.A2(n_223),
.B(n_229),
.Y(n_274)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_134),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_L g222 ( 
.A1(n_132),
.A2(n_172),
.B1(n_165),
.B2(n_161),
.Y(n_222)
);

INVx1_ASAP7_75t_SL g223 ( 
.A(n_114),
.Y(n_223)
);

INVx3_ASAP7_75t_L g224 ( 
.A(n_150),
.Y(n_224)
);

CKINVDCx16_ASAP7_75t_R g279 ( 
.A(n_224),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_116),
.Y(n_226)
);

INVx3_ASAP7_75t_L g227 ( 
.A(n_147),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_227),
.B(n_229),
.Y(n_258)
);

INVx13_ASAP7_75t_L g228 ( 
.A(n_111),
.Y(n_228)
);

NAND2xp33_ASAP7_75t_SL g257 ( 
.A(n_228),
.B(n_231),
.Y(n_257)
);

INVxp67_ASAP7_75t_L g229 ( 
.A(n_126),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_116),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_230),
.Y(n_252)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_132),
.Y(n_231)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_146),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_232),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_166),
.B(n_158),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_233),
.B(n_234),
.Y(n_261)
);

CKINVDCx14_ASAP7_75t_R g234 ( 
.A(n_159),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_146),
.B(n_164),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_235),
.B(n_198),
.Y(n_266)
);

OAI22x1_ASAP7_75t_L g309 ( 
.A1(n_236),
.A2(n_271),
.B1(n_274),
.B2(n_278),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_L g289 ( 
.A1(n_238),
.A2(n_262),
.B1(n_269),
.B2(n_272),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_SL g243 ( 
.A(n_225),
.B(n_139),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g303 ( 
.A(n_243),
.B(n_255),
.Y(n_303)
);

OA22x2_ASAP7_75t_L g247 ( 
.A1(n_192),
.A2(n_155),
.B1(n_138),
.B2(n_144),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_247),
.B(n_264),
.Y(n_283)
);

MAJx2_ASAP7_75t_L g255 ( 
.A(n_225),
.B(n_114),
.C(n_155),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g312 ( 
.A1(n_259),
.A2(n_265),
.B1(n_242),
.B2(n_260),
.Y(n_312)
);

AOI22xp33_ASAP7_75t_L g313 ( 
.A1(n_260),
.A2(n_247),
.B1(n_248),
.B2(n_264),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_181),
.A2(n_161),
.B1(n_165),
.B2(n_172),
.Y(n_262)
);

OA22x2_ASAP7_75t_L g264 ( 
.A1(n_184),
.A2(n_206),
.B1(n_189),
.B2(n_191),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_184),
.A2(n_186),
.B1(n_206),
.B2(n_201),
.Y(n_265)
);

CKINVDCx16_ASAP7_75t_R g306 ( 
.A(n_266),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_225),
.A2(n_219),
.B1(n_206),
.B2(n_217),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_179),
.A2(n_194),
.B1(n_196),
.B2(n_221),
.Y(n_272)
);

AND2x2_ASAP7_75t_SL g275 ( 
.A(n_185),
.B(n_202),
.Y(n_275)
);

INVx1_ASAP7_75t_SL g293 ( 
.A(n_275),
.Y(n_293)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_276),
.Y(n_280)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_280),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_261),
.B(n_203),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_SL g323 ( 
.A(n_281),
.B(n_290),
.Y(n_323)
);

AOI22xp33_ASAP7_75t_SL g282 ( 
.A1(n_250),
.A2(n_204),
.B1(n_227),
.B2(n_199),
.Y(n_282)
);

AOI22xp33_ASAP7_75t_SL g319 ( 
.A1(n_282),
.A2(n_305),
.B1(n_307),
.B2(n_309),
.Y(n_319)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_276),
.Y(n_284)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_284),
.Y(n_325)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_248),
.Y(n_285)
);

BUFx2_ASAP7_75t_L g335 ( 
.A(n_285),
.Y(n_335)
);

OAI22xp5_ASAP7_75t_SL g286 ( 
.A1(n_269),
.A2(n_231),
.B1(n_209),
.B2(n_213),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g326 ( 
.A1(n_286),
.A2(n_292),
.B1(n_300),
.B2(n_289),
.Y(n_326)
);

XOR2xp5_ASAP7_75t_L g287 ( 
.A(n_251),
.B(n_182),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_287),
.B(n_303),
.C(n_296),
.Y(n_321)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_253),
.Y(n_288)
);

INVx2_ASAP7_75t_SL g329 ( 
.A(n_288),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_261),
.B(n_232),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_240),
.B(n_210),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_291),
.B(n_296),
.Y(n_315)
);

OAI22xp33_ASAP7_75t_SL g292 ( 
.A1(n_238),
.A2(n_195),
.B1(n_200),
.B2(n_224),
.Y(n_292)
);

AOI21xp33_ASAP7_75t_L g294 ( 
.A1(n_250),
.A2(n_187),
.B(n_228),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_SL g317 ( 
.A(n_294),
.B(n_298),
.Y(n_317)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_253),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_SL g333 ( 
.A(n_295),
.B(n_297),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_240),
.B(n_251),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_237),
.B(n_183),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_265),
.B(n_207),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g299 ( 
.A(n_249),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_SL g324 ( 
.A(n_299),
.B(n_301),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_L g300 ( 
.A1(n_262),
.A2(n_264),
.B1(n_272),
.B2(n_242),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_SL g301 ( 
.A(n_244),
.B(n_275),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g302 ( 
.A(n_275),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g327 ( 
.A(n_302),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_252),
.B(n_242),
.Y(n_304)
);

XOR2xp5_ASAP7_75t_SL g314 ( 
.A(n_304),
.B(n_255),
.Y(n_314)
);

BUFx6f_ASAP7_75t_L g305 ( 
.A(n_241),
.Y(n_305)
);

BUFx6f_ASAP7_75t_L g307 ( 
.A(n_241),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_256),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g328 ( 
.A(n_308),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_246),
.B(n_268),
.Y(n_310)
);

CKINVDCx16_ASAP7_75t_R g330 ( 
.A(n_310),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_266),
.B(n_279),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g331 ( 
.A(n_311),
.Y(n_331)
);

OAI22xp5_ASAP7_75t_L g316 ( 
.A1(n_312),
.A2(n_313),
.B1(n_264),
.B2(n_274),
.Y(n_316)
);

XOR2xp5_ASAP7_75t_L g347 ( 
.A(n_314),
.B(n_286),
.Y(n_347)
);

AOI22xp5_ASAP7_75t_L g353 ( 
.A1(n_316),
.A2(n_320),
.B1(n_338),
.B2(n_277),
.Y(n_353)
);

OAI22xp5_ASAP7_75t_L g320 ( 
.A1(n_312),
.A2(n_247),
.B1(n_271),
.B2(n_243),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g343 ( 
.A(n_321),
.B(n_303),
.C(n_301),
.Y(n_343)
);

AO21x1_ASAP7_75t_L g322 ( 
.A1(n_298),
.A2(n_283),
.B(n_300),
.Y(n_322)
);

INVxp67_ASAP7_75t_L g359 ( 
.A(n_322),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_326),
.B(n_339),
.Y(n_356)
);

AOI22xp5_ASAP7_75t_L g332 ( 
.A1(n_289),
.A2(n_247),
.B1(n_278),
.B2(n_270),
.Y(n_332)
);

OAI22xp5_ASAP7_75t_SL g351 ( 
.A1(n_332),
.A2(n_295),
.B1(n_288),
.B2(n_285),
.Y(n_351)
);

AND2x6_ASAP7_75t_L g334 ( 
.A(n_287),
.B(n_257),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g354 ( 
.A(n_334),
.B(n_337),
.Y(n_354)
);

OAI21xp5_ASAP7_75t_L g336 ( 
.A1(n_304),
.A2(n_239),
.B(n_258),
.Y(n_336)
);

OAI21xp5_ASAP7_75t_SL g357 ( 
.A1(n_336),
.A2(n_267),
.B(n_245),
.Y(n_357)
);

AND2x6_ASAP7_75t_L g337 ( 
.A(n_309),
.B(n_254),
.Y(n_337)
);

OAI22xp5_ASAP7_75t_SL g338 ( 
.A1(n_283),
.A2(n_291),
.B1(n_306),
.B2(n_293),
.Y(n_338)
);

CKINVDCx20_ASAP7_75t_R g339 ( 
.A(n_280),
.Y(n_339)
);

CKINVDCx16_ASAP7_75t_R g340 ( 
.A(n_324),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_SL g369 ( 
.A(n_340),
.B(n_355),
.Y(n_369)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_329),
.Y(n_341)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_341),
.Y(n_376)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_329),
.Y(n_342)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_342),
.Y(n_378)
);

MAJIxp5_ASAP7_75t_L g365 ( 
.A(n_343),
.B(n_349),
.C(n_350),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_SL g344 ( 
.A(n_328),
.B(n_299),
.Y(n_344)
);

CKINVDCx14_ASAP7_75t_R g364 ( 
.A(n_344),
.Y(n_364)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_329),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_345),
.B(n_346),
.Y(n_375)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_318),
.Y(n_346)
);

XNOR2xp5_ASAP7_75t_SL g367 ( 
.A(n_347),
.B(n_334),
.Y(n_367)
);

OAI22xp5_ASAP7_75t_L g348 ( 
.A1(n_326),
.A2(n_306),
.B1(n_302),
.B2(n_293),
.Y(n_348)
);

OAI22xp5_ASAP7_75t_SL g368 ( 
.A1(n_348),
.A2(n_353),
.B1(n_322),
.B2(n_327),
.Y(n_368)
);

XNOR2xp5_ASAP7_75t_L g349 ( 
.A(n_321),
.B(n_315),
.Y(n_349)
);

MAJIxp5_ASAP7_75t_L g350 ( 
.A(n_314),
.B(n_308),
.C(n_284),
.Y(n_350)
);

AND2x4_ASAP7_75t_L g374 ( 
.A(n_351),
.B(n_325),
.Y(n_374)
);

XOR2xp5_ASAP7_75t_L g352 ( 
.A(n_315),
.B(n_273),
.Y(n_352)
);

MAJIxp5_ASAP7_75t_L g371 ( 
.A(n_352),
.B(n_333),
.C(n_331),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_SL g355 ( 
.A(n_328),
.B(n_277),
.Y(n_355)
);

OAI21xp33_ASAP7_75t_L g363 ( 
.A1(n_357),
.A2(n_327),
.B(n_336),
.Y(n_363)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_318),
.Y(n_358)
);

NOR2xp33_ASAP7_75t_L g370 ( 
.A(n_358),
.B(n_360),
.Y(n_370)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_325),
.Y(n_360)
);

CKINVDCx16_ASAP7_75t_R g361 ( 
.A(n_355),
.Y(n_361)
);

NOR2xp33_ASAP7_75t_L g382 ( 
.A(n_361),
.B(n_377),
.Y(n_382)
);

XOR2xp5_ASAP7_75t_L g362 ( 
.A(n_349),
.B(n_338),
.Y(n_362)
);

XOR2xp5_ASAP7_75t_L g387 ( 
.A(n_362),
.B(n_366),
.Y(n_387)
);

AOI22xp33_ASAP7_75t_SL g389 ( 
.A1(n_363),
.A2(n_317),
.B1(n_351),
.B2(n_337),
.Y(n_389)
);

XNOR2xp5_ASAP7_75t_L g366 ( 
.A(n_343),
.B(n_320),
.Y(n_366)
);

XNOR2xp5_ASAP7_75t_SL g380 ( 
.A(n_367),
.B(n_347),
.Y(n_380)
);

AOI22xp5_ASAP7_75t_SL g392 ( 
.A1(n_368),
.A2(n_345),
.B1(n_341),
.B2(n_339),
.Y(n_392)
);

MAJIxp5_ASAP7_75t_L g383 ( 
.A(n_371),
.B(n_373),
.C(n_357),
.Y(n_383)
);

NOR2xp33_ASAP7_75t_L g372 ( 
.A(n_352),
.B(n_324),
.Y(n_372)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_372),
.Y(n_388)
);

MAJIxp5_ASAP7_75t_L g373 ( 
.A(n_350),
.B(n_322),
.C(n_331),
.Y(n_373)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_374),
.Y(n_379)
);

CKINVDCx20_ASAP7_75t_R g377 ( 
.A(n_348),
.Y(n_377)
);

XOR2xp5_ASAP7_75t_L g394 ( 
.A(n_380),
.B(n_362),
.Y(n_394)
);

OAI21xp5_ASAP7_75t_L g381 ( 
.A1(n_368),
.A2(n_359),
.B(n_354),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_381),
.B(n_384),
.Y(n_397)
);

MAJx2_ASAP7_75t_L g395 ( 
.A(n_383),
.B(n_365),
.C(n_367),
.Y(n_395)
);

OAI22xp5_ASAP7_75t_L g384 ( 
.A1(n_364),
.A2(n_332),
.B1(n_323),
.B2(n_356),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_370),
.Y(n_385)
);

OAI22xp5_ASAP7_75t_L g400 ( 
.A1(n_385),
.A2(n_389),
.B1(n_391),
.B2(n_369),
.Y(n_400)
);

OAI22xp5_ASAP7_75t_SL g386 ( 
.A1(n_373),
.A2(n_353),
.B1(n_359),
.B2(n_356),
.Y(n_386)
);

AOI22xp5_ASAP7_75t_L g402 ( 
.A1(n_386),
.A2(n_390),
.B1(n_374),
.B2(n_381),
.Y(n_402)
);

OAI22xp5_ASAP7_75t_SL g390 ( 
.A1(n_371),
.A2(n_319),
.B1(n_317),
.B2(n_342),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_375),
.Y(n_391)
);

OAI22xp5_ASAP7_75t_SL g401 ( 
.A1(n_392),
.A2(n_374),
.B1(n_360),
.B2(n_358),
.Y(n_401)
);

MAJIxp5_ASAP7_75t_L g393 ( 
.A(n_387),
.B(n_365),
.C(n_366),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_393),
.B(n_398),
.Y(n_404)
);

XNOR2xp5_ASAP7_75t_L g406 ( 
.A(n_394),
.B(n_395),
.Y(n_406)
);

OA21x2_ASAP7_75t_L g396 ( 
.A1(n_379),
.A2(n_375),
.B(n_374),
.Y(n_396)
);

INVxp67_ASAP7_75t_L g405 ( 
.A(n_396),
.Y(n_405)
);

MAJIxp5_ASAP7_75t_L g398 ( 
.A(n_387),
.B(n_378),
.C(n_376),
.Y(n_398)
);

MAJIxp5_ASAP7_75t_L g399 ( 
.A(n_383),
.B(n_378),
.C(n_376),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_SL g408 ( 
.A(n_399),
.B(n_402),
.Y(n_408)
);

AOI22xp5_ASAP7_75t_L g410 ( 
.A1(n_400),
.A2(n_403),
.B1(n_390),
.B2(n_386),
.Y(n_410)
);

INVxp67_ASAP7_75t_L g412 ( 
.A(n_401),
.Y(n_412)
);

OAI22xp5_ASAP7_75t_SL g403 ( 
.A1(n_392),
.A2(n_330),
.B1(n_346),
.B2(n_305),
.Y(n_403)
);

XNOR2xp5_ASAP7_75t_L g407 ( 
.A(n_393),
.B(n_382),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g417 ( 
.A(n_407),
.B(n_409),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_SL g409 ( 
.A(n_399),
.B(n_388),
.Y(n_409)
);

HB1xp67_ASAP7_75t_L g418 ( 
.A(n_410),
.Y(n_418)
);

MAJIxp5_ASAP7_75t_L g411 ( 
.A(n_398),
.B(n_391),
.C(n_379),
.Y(n_411)
);

AND2x2_ASAP7_75t_L g414 ( 
.A(n_411),
.B(n_408),
.Y(n_414)
);

OAI21xp5_ASAP7_75t_L g413 ( 
.A1(n_404),
.A2(n_397),
.B(n_403),
.Y(n_413)
);

NOR2xp33_ASAP7_75t_SL g423 ( 
.A(n_413),
.B(n_415),
.Y(n_423)
);

CKINVDCx20_ASAP7_75t_R g424 ( 
.A(n_414),
.Y(n_424)
);

NOR2xp33_ASAP7_75t_L g415 ( 
.A(n_411),
.B(n_385),
.Y(n_415)
);

NOR2xp33_ASAP7_75t_L g416 ( 
.A(n_412),
.B(n_402),
.Y(n_416)
);

AOI322xp5_ASAP7_75t_L g420 ( 
.A1(n_416),
.A2(n_419),
.A3(n_405),
.B1(n_418),
.B2(n_396),
.C1(n_417),
.C2(n_395),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_SL g419 ( 
.A(n_412),
.B(n_401),
.Y(n_419)
);

OR2x2_ASAP7_75t_L g427 ( 
.A(n_420),
.B(n_421),
.Y(n_427)
);

MAJIxp5_ASAP7_75t_L g421 ( 
.A(n_419),
.B(n_406),
.C(n_405),
.Y(n_421)
);

AOI322xp5_ASAP7_75t_L g422 ( 
.A1(n_415),
.A2(n_396),
.A3(n_380),
.B1(n_307),
.B2(n_305),
.C1(n_394),
.C2(n_335),
.Y(n_422)
);

MAJIxp5_ASAP7_75t_L g426 ( 
.A(n_422),
.B(n_335),
.C(n_267),
.Y(n_426)
);

OAI21xp5_ASAP7_75t_L g425 ( 
.A1(n_424),
.A2(n_335),
.B(n_307),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_425),
.B(n_426),
.Y(n_428)
);

XOR2x2_ASAP7_75t_L g429 ( 
.A(n_427),
.B(n_421),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_429),
.B(n_423),
.Y(n_430)
);

NOR2xp33_ASAP7_75t_SL g431 ( 
.A(n_430),
.B(n_428),
.Y(n_431)
);

OAI21xp5_ASAP7_75t_SL g432 ( 
.A1(n_431),
.A2(n_245),
.B(n_270),
.Y(n_432)
);

XNOR2xp5_ASAP7_75t_L g433 ( 
.A(n_432),
.B(n_263),
.Y(n_433)
);


endmodule