module fake_jpeg_21518_n_187 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_187);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_187;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_175;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_121;
wire n_102;
wire n_130;
wire n_99;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_5),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_12),
.Y(n_14)
);

INVx4_ASAP7_75t_L g15 ( 
.A(n_7),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_5),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

INVx3_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

INVxp67_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

BUFx10_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

BUFx4f_ASAP7_75t_SL g28 ( 
.A(n_0),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_27),
.B(n_0),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_30),
.B(n_34),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_24),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_31),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_26),
.Y(n_32)
);

INVx5_ASAP7_75t_L g58 ( 
.A(n_32),
.Y(n_58)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_17),
.Y(n_33)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_33),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_27),
.B(n_1),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_17),
.Y(n_35)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_35),
.Y(n_54)
);

INVx2_ASAP7_75t_R g36 ( 
.A(n_28),
.Y(n_36)
);

AND2x2_ASAP7_75t_L g49 ( 
.A(n_36),
.B(n_27),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_24),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_37),
.Y(n_55)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_26),
.Y(n_38)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_38),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_24),
.Y(n_39)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_39),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_27),
.B(n_2),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_40),
.B(n_16),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_26),
.Y(n_41)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_41),
.Y(n_50)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_18),
.Y(n_42)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_42),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_26),
.Y(n_43)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_43),
.Y(n_52)
);

HB1xp67_ASAP7_75t_L g44 ( 
.A(n_28),
.Y(n_44)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_44),
.Y(n_62)
);

CKINVDCx12_ASAP7_75t_R g47 ( 
.A(n_36),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_47),
.B(n_28),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_49),
.A2(n_61),
.B1(n_44),
.B2(n_19),
.Y(n_82)
);

INVxp67_ASAP7_75t_L g56 ( 
.A(n_36),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_56),
.B(n_43),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_38),
.A2(n_15),
.B1(n_21),
.B2(n_16),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_57),
.A2(n_64),
.B1(n_13),
.B2(n_29),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g93 ( 
.A(n_59),
.B(n_2),
.Y(n_93)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_32),
.Y(n_60)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_60),
.Y(n_66)
);

MAJIxp5_ASAP7_75t_L g61 ( 
.A(n_32),
.B(n_27),
.C(n_15),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g64 ( 
.A1(n_30),
.A2(n_21),
.B1(n_13),
.B2(n_14),
.Y(n_64)
);

OAI21xp5_ASAP7_75t_L g65 ( 
.A1(n_49),
.A2(n_34),
.B(n_40),
.Y(n_65)
);

AOI21xp5_ASAP7_75t_SL g106 ( 
.A1(n_65),
.A2(n_83),
.B(n_41),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_51),
.B(n_42),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_67),
.B(n_79),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_L g68 ( 
.A1(n_54),
.A2(n_33),
.B1(n_35),
.B2(n_37),
.Y(n_68)
);

OAI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_68),
.A2(n_69),
.B1(n_3),
.B2(n_4),
.Y(n_114)
);

AOI21xp33_ASAP7_75t_L g70 ( 
.A1(n_48),
.A2(n_20),
.B(n_22),
.Y(n_70)
);

NOR2x1_ASAP7_75t_L g104 ( 
.A(n_70),
.B(n_19),
.Y(n_104)
);

CKINVDCx16_ASAP7_75t_R g113 ( 
.A(n_71),
.Y(n_113)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_62),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_72),
.Y(n_108)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_62),
.Y(n_73)
);

INVx6_ASAP7_75t_L g111 ( 
.A(n_73),
.Y(n_111)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_63),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_74),
.B(n_75),
.Y(n_102)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_50),
.Y(n_75)
);

AOI32xp33_ASAP7_75t_L g76 ( 
.A1(n_56),
.A2(n_25),
.A3(n_20),
.B1(n_22),
.B2(n_14),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_76),
.B(n_77),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_61),
.B(n_28),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_45),
.Y(n_78)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_78),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_49),
.B(n_39),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_46),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_80),
.B(n_84),
.Y(n_105)
);

HB1xp67_ASAP7_75t_L g81 ( 
.A(n_46),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_81),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_82),
.B(n_41),
.C(n_60),
.Y(n_94)
);

AND2x4_ASAP7_75t_L g83 ( 
.A(n_53),
.B(n_32),
.Y(n_83)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_50),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_53),
.A2(n_18),
.B1(n_29),
.B2(n_23),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_85),
.A2(n_88),
.B1(n_55),
.B2(n_31),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_45),
.B(n_39),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_86),
.B(n_93),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_58),
.B(n_23),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_87),
.B(n_89),
.Y(n_107)
);

OA22x2_ASAP7_75t_L g88 ( 
.A1(n_52),
.A2(n_37),
.B1(n_31),
.B2(n_43),
.Y(n_88)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_52),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_90),
.B(n_91),
.Y(n_109)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_55),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_58),
.B(n_11),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_92),
.Y(n_99)
);

XNOR2xp5_ASAP7_75t_L g129 ( 
.A(n_94),
.B(n_106),
.Y(n_129)
);

CKINVDCx14_ASAP7_75t_R g126 ( 
.A(n_100),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_67),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_101),
.B(n_104),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_82),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_110),
.A2(n_72),
.B1(n_90),
.B2(n_75),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_86),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_112),
.B(n_84),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_114),
.B(n_88),
.Y(n_118)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_88),
.Y(n_115)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_115),
.Y(n_116)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_105),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_117),
.B(n_119),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_118),
.A2(n_131),
.B1(n_115),
.B2(n_126),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_101),
.B(n_79),
.Y(n_119)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_109),
.Y(n_121)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_121),
.Y(n_134)
);

INVx4_ASAP7_75t_L g122 ( 
.A(n_111),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_122),
.B(n_127),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_95),
.B(n_65),
.C(n_83),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_123),
.B(n_103),
.C(n_107),
.Y(n_140)
);

NAND2xp67_ASAP7_75t_L g124 ( 
.A(n_106),
.B(n_83),
.Y(n_124)
);

XNOR2xp5_ASAP7_75t_L g143 ( 
.A(n_124),
.B(n_110),
.Y(n_143)
);

AOI21xp5_ASAP7_75t_L g125 ( 
.A1(n_100),
.A2(n_83),
.B(n_73),
.Y(n_125)
);

AOI21xp5_ASAP7_75t_L g138 ( 
.A1(n_125),
.A2(n_95),
.B(n_94),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_102),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_112),
.B(n_88),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_128),
.B(n_130),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_132),
.B(n_143),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_121),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_135),
.B(n_137),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_130),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_L g148 ( 
.A1(n_138),
.A2(n_123),
.B(n_120),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_140),
.B(n_141),
.C(n_142),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_129),
.B(n_113),
.C(n_96),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_129),
.B(n_113),
.C(n_96),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_125),
.A2(n_104),
.B1(n_97),
.B2(n_98),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_144),
.B(n_145),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_116),
.A2(n_128),
.B1(n_118),
.B2(n_124),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_133),
.B(n_127),
.Y(n_146)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_146),
.Y(n_163)
);

XNOR2x1_ASAP7_75t_L g161 ( 
.A(n_148),
.B(n_122),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_136),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_149),
.B(n_150),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_134),
.Y(n_150)
);

AND2x6_ASAP7_75t_L g153 ( 
.A(n_144),
.B(n_120),
.Y(n_153)
);

INVxp67_ASAP7_75t_L g162 ( 
.A(n_153),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_139),
.B(n_119),
.Y(n_154)
);

CKINVDCx16_ASAP7_75t_R g165 ( 
.A(n_154),
.Y(n_165)
);

AOI322xp5_ASAP7_75t_L g155 ( 
.A1(n_138),
.A2(n_116),
.A3(n_131),
.B1(n_99),
.B2(n_98),
.C1(n_97),
.C2(n_111),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_155),
.B(n_140),
.C(n_143),
.Y(n_160)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_145),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_157),
.A2(n_132),
.B1(n_142),
.B2(n_141),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_SL g158 ( 
.A(n_156),
.B(n_99),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_158),
.B(n_159),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_160),
.A2(n_147),
.B1(n_148),
.B2(n_153),
.Y(n_167)
);

XOR2xp5_ASAP7_75t_L g171 ( 
.A(n_161),
.B(n_108),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_147),
.B(n_108),
.C(n_66),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_L g172 ( 
.A(n_164),
.B(n_108),
.Y(n_172)
);

XOR2xp5_ASAP7_75t_L g176 ( 
.A(n_167),
.B(n_168),
.Y(n_176)
);

OAI322xp33_ASAP7_75t_L g168 ( 
.A1(n_163),
.A2(n_150),
.A3(n_154),
.B1(n_157),
.B2(n_151),
.C1(n_152),
.C2(n_5),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_162),
.A2(n_152),
.B1(n_151),
.B2(n_66),
.Y(n_170)
);

XOR2xp5_ASAP7_75t_L g175 ( 
.A(n_170),
.B(n_171),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_172),
.B(n_164),
.C(n_161),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_L g173 ( 
.A1(n_162),
.A2(n_6),
.B(n_8),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_L g178 ( 
.A1(n_173),
.A2(n_6),
.B(n_8),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_174),
.B(n_177),
.C(n_172),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_169),
.B(n_166),
.C(n_165),
.Y(n_177)
);

AOI21xp5_ASAP7_75t_SL g179 ( 
.A1(n_178),
.A2(n_173),
.B(n_170),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_179),
.B(n_180),
.Y(n_182)
);

AOI322xp5_ASAP7_75t_L g181 ( 
.A1(n_176),
.A2(n_175),
.A3(n_171),
.B1(n_78),
.B2(n_10),
.C1(n_9),
.C2(n_6),
.Y(n_181)
);

OR2x2_ASAP7_75t_L g183 ( 
.A(n_181),
.B(n_175),
.Y(n_183)
);

AOI21xp5_ASAP7_75t_SL g184 ( 
.A1(n_183),
.A2(n_10),
.B(n_182),
.Y(n_184)
);

INVxp67_ASAP7_75t_L g185 ( 
.A(n_184),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_185),
.B(n_10),
.Y(n_186)
);

BUFx24_ASAP7_75t_SL g187 ( 
.A(n_186),
.Y(n_187)
);


endmodule