module fake_ibex_1777_n_37 (n_4, n_2, n_7, n_5, n_11, n_6, n_8, n_10, n_0, n_9, n_3, n_1, n_37);

input n_4;
input n_2;
input n_7;
input n_5;
input n_11;
input n_6;
input n_8;
input n_10;
input n_0;
input n_9;
input n_3;
input n_1;

output n_37;

wire n_20;
wire n_17;
wire n_25;
wire n_36;
wire n_18;
wire n_22;
wire n_28;
wire n_32;
wire n_33;
wire n_30;
wire n_29;
wire n_13;
wire n_26;
wire n_35;
wire n_14;
wire n_34;
wire n_12;
wire n_15;
wire n_24;
wire n_31;
wire n_23;
wire n_21;
wire n_27;
wire n_19;
wire n_16;

INVx1_ASAP7_75t_L g12 ( 
.A(n_2),
.Y(n_12)
);

BUFx3_ASAP7_75t_L g13 ( 
.A(n_7),
.Y(n_13)
);

AND2x6_ASAP7_75t_L g14 ( 
.A(n_5),
.B(n_8),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_0),
.Y(n_15)
);

INVx2_ASAP7_75t_L g16 ( 
.A(n_11),
.Y(n_16)
);

BUFx10_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

HB1xp67_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

AOI21xp5_ASAP7_75t_L g23 ( 
.A1(n_16),
.A2(n_4),
.B(n_6),
.Y(n_23)
);

OAI21x1_ASAP7_75t_L g24 ( 
.A1(n_20),
.A2(n_22),
.B(n_18),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_19),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

INVx2_ASAP7_75t_SL g27 ( 
.A(n_17),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_21),
.Y(n_28)
);

AOI22xp33_ASAP7_75t_L g29 ( 
.A1(n_25),
.A2(n_12),
.B1(n_15),
.B2(n_14),
.Y(n_29)
);

AND2x2_ASAP7_75t_L g30 ( 
.A(n_27),
.B(n_14),
.Y(n_30)
);

AO21x2_ASAP7_75t_L g31 ( 
.A1(n_24),
.A2(n_14),
.B(n_1),
.Y(n_31)
);

AOI22xp33_ASAP7_75t_L g32 ( 
.A1(n_24),
.A2(n_1),
.B1(n_28),
.B2(n_26),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_30),
.B(n_27),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_31),
.Y(n_34)
);

AOI221xp5_ASAP7_75t_L g35 ( 
.A1(n_33),
.A2(n_29),
.B1(n_32),
.B2(n_26),
.C(n_31),
.Y(n_35)
);

AOI31xp33_ASAP7_75t_L g36 ( 
.A1(n_35),
.A2(n_34),
.A3(n_23),
.B(n_26),
.Y(n_36)
);

XNOR2xp5_ASAP7_75t_L g37 ( 
.A(n_36),
.B(n_26),
.Y(n_37)
);


endmodule