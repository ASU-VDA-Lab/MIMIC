module real_jpeg_4647_n_15 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_6, n_7, n_3, n_10, n_9, n_15);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_15;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_201;
wire n_114;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_78;
wire n_83;
wire n_249;
wire n_215;
wire n_176;
wire n_166;
wire n_221;
wire n_300;
wire n_286;
wire n_288;
wire n_292;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_301;
wire n_280;
wire n_64;
wire n_177;
wire n_291;
wire n_236;
wire n_47;
wire n_131;
wire n_281;
wire n_271;
wire n_276;
wire n_163;
wire n_22;
wire n_287;
wire n_174;
wire n_237;
wire n_87;
wire n_255;
wire n_105;
wire n_40;
wire n_197;
wire n_173;
wire n_299;
wire n_115;
wire n_243;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_275;
wire n_293;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_120;
wire n_155;
wire n_113;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_139;
wire n_33;
wire n_65;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_282;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_44;
wire n_28;
wire n_267;
wire n_305;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_290;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_285;
wire n_304;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_302;
wire n_26;
wire n_148;
wire n_222;
wire n_19;
wire n_262;
wire n_118;
wire n_220;
wire n_294;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_137;
wire n_31;
wire n_298;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_296;
wire n_134;
wire n_270;
wire n_223;
wire n_159;
wire n_72;
wire n_303;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_205;
wire n_195;
wire n_258;
wire n_289;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_278;
wire n_130;
wire n_241;
wire n_225;
wire n_103;
wire n_259;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_284;
wire n_226;
wire n_277;
wire n_125;
wire n_297;
wire n_185;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_240;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_97;
wire n_187;
wire n_75;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_279;
wire n_216;
wire n_244;
wire n_295;
wire n_128;
wire n_167;
wire n_179;
wire n_133;
wire n_213;
wire n_202;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_102;
wire n_81;
wire n_85;
wire n_181;
wire n_283;
wire n_101;
wire n_256;
wire n_274;
wire n_182;
wire n_253;
wire n_96;
wire n_273;
wire n_269;
wire n_89;
wire n_16;

INVx8_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_1),
.A2(n_96),
.B1(n_97),
.B2(n_101),
.Y(n_95)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_1),
.Y(n_101)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_2),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_2),
.Y(n_94)
);

BUFx3_ASAP7_75t_L g161 ( 
.A(n_2),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_SL g34 ( 
.A1(n_3),
.A2(n_35),
.B1(n_39),
.B2(n_43),
.Y(n_34)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_3),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_L g260 ( 
.A1(n_3),
.A2(n_43),
.B1(n_129),
.B2(n_148),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_L g275 ( 
.A1(n_3),
.A2(n_43),
.B1(n_159),
.B2(n_250),
.Y(n_275)
);

AOI22xp33_ASAP7_75t_L g79 ( 
.A1(n_4),
.A2(n_80),
.B1(n_86),
.B2(n_87),
.Y(n_79)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_4),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g221 ( 
.A1(n_4),
.A2(n_86),
.B1(n_109),
.B2(n_222),
.Y(n_221)
);

INVx6_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

INVx8_ASAP7_75t_L g91 ( 
.A(n_6),
.Y(n_91)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_6),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g156 ( 
.A(n_6),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g256 ( 
.A(n_6),
.Y(n_256)
);

AOI22xp33_ASAP7_75t_L g185 ( 
.A1(n_7),
.A2(n_159),
.B1(n_186),
.B2(n_187),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_7),
.Y(n_186)
);

BUFx5_ASAP7_75t_L g71 ( 
.A(n_8),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_8),
.Y(n_77)
);

INVx3_ASAP7_75t_L g173 ( 
.A(n_8),
.Y(n_173)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_9),
.Y(n_38)
);

BUFx5_ASAP7_75t_L g169 ( 
.A(n_10),
.Y(n_169)
);

BUFx5_ASAP7_75t_L g179 ( 
.A(n_10),
.Y(n_179)
);

BUFx6f_ASAP7_75t_L g199 ( 
.A(n_10),
.Y(n_199)
);

BUFx6f_ASAP7_75t_L g201 ( 
.A(n_10),
.Y(n_201)
);

BUFx6f_ASAP7_75t_L g207 ( 
.A(n_10),
.Y(n_207)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_10),
.Y(n_211)
);

AOI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_11),
.A2(n_129),
.B1(n_130),
.B2(n_133),
.Y(n_128)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_11),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_L g215 ( 
.A1(n_11),
.A2(n_133),
.B1(n_216),
.B2(n_218),
.Y(n_215)
);

OAI22xp33_ASAP7_75t_SL g249 ( 
.A1(n_11),
.A2(n_80),
.B1(n_133),
.B2(n_250),
.Y(n_249)
);

BUFx3_ASAP7_75t_L g113 ( 
.A(n_12),
.Y(n_113)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_12),
.Y(n_117)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_12),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g46 ( 
.A1(n_13),
.A2(n_47),
.B1(n_51),
.B2(n_52),
.Y(n_46)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_13),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_13),
.A2(n_51),
.B1(n_136),
.B2(n_137),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_L g158 ( 
.A1(n_13),
.A2(n_51),
.B1(n_87),
.B2(n_159),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g204 ( 
.A1(n_13),
.A2(n_51),
.B1(n_205),
.B2(n_208),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_14),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_14),
.B(n_144),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_SL g233 ( 
.A1(n_14),
.A2(n_69),
.B1(n_129),
.B2(n_234),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_14),
.B(n_241),
.C(n_244),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_SL g262 ( 
.A(n_14),
.B(n_23),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_14),
.B(n_256),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_14),
.B(n_139),
.Y(n_277)
);

XOR2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_227),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_225),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_162),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_SL g226 ( 
.A(n_18),
.B(n_162),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_105),
.C(n_140),
.Y(n_18)
);

AOI22xp5_ASAP7_75t_L g302 ( 
.A1(n_19),
.A2(n_20),
.B1(n_303),
.B2(n_304),
.Y(n_302)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

XNOR2xp5_ASAP7_75t_SL g20 ( 
.A(n_21),
.B(n_67),
.Y(n_20)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_21),
.B(n_68),
.C(n_78),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_SL g21 ( 
.A1(n_22),
.A2(n_34),
.B(n_44),
.Y(n_21)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_22),
.A2(n_34),
.B1(n_56),
.B2(n_215),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_22),
.B(n_46),
.Y(n_297)
);

INVx1_ASAP7_75t_SL g22 ( 
.A(n_23),
.Y(n_22)
);

OR2x2_ASAP7_75t_L g56 ( 
.A(n_23),
.B(n_57),
.Y(n_56)
);

AO22x2_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_27),
.B1(n_29),
.B2(n_31),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_25),
.Y(n_64)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_26),
.Y(n_33)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVx11_ASAP7_75t_L g30 ( 
.A(n_28),
.Y(n_30)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_28),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_28),
.Y(n_129)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_28),
.Y(n_132)
);

INVx3_ASAP7_75t_L g138 ( 
.A(n_28),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx5_ASAP7_75t_L g119 ( 
.A(n_30),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g222 ( 
.A(n_30),
.Y(n_222)
);

INVx6_ASAP7_75t_L g237 ( 
.A(n_30),
.Y(n_237)
);

AOI32xp33_ASAP7_75t_L g141 ( 
.A1(n_31),
.A2(n_129),
.A3(n_142),
.B1(n_143),
.B2(n_147),
.Y(n_141)
);

INVx5_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

BUFx2_ASAP7_75t_L g151 ( 
.A(n_32),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_33),
.Y(n_60)
);

INVx5_ASAP7_75t_L g218 ( 
.A(n_35),
.Y(n_218)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_37),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

BUFx5_ASAP7_75t_L g42 ( 
.A(n_38),
.Y(n_42)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_38),
.Y(n_75)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx6_ASAP7_75t_L g146 ( 
.A(n_42),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_45),
.B(n_55),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

BUFx5_ASAP7_75t_L g61 ( 
.A(n_50),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_50),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g167 ( 
.A(n_50),
.Y(n_167)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

AOI21xp5_ASAP7_75t_L g294 ( 
.A1(n_55),
.A2(n_295),
.B(n_297),
.Y(n_294)
);

INVx3_ASAP7_75t_SL g55 ( 
.A(n_56),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_L g57 ( 
.A1(n_58),
.A2(n_61),
.B1(n_62),
.B2(n_65),
.Y(n_57)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_65),
.B(n_175),
.Y(n_174)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

OAI21xp33_ASAP7_75t_SL g295 ( 
.A1(n_66),
.A2(n_69),
.B(n_296),
.Y(n_295)
);

XOR2xp5_ASAP7_75t_L g67 ( 
.A(n_68),
.B(n_78),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_69),
.B(n_70),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_69),
.B(n_177),
.Y(n_176)
);

OAI21xp33_ASAP7_75t_SL g200 ( 
.A1(n_69),
.A2(n_176),
.B(n_201),
.Y(n_200)
);

AOI21xp5_ASAP7_75t_L g272 ( 
.A1(n_69),
.A2(n_182),
.B(n_254),
.Y(n_272)
);

AND2x2_ASAP7_75t_L g195 ( 
.A(n_70),
.B(n_196),
.Y(n_195)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_70),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_71),
.A2(n_72),
.B1(n_74),
.B2(n_76),
.Y(n_70)
);

INVx6_ASAP7_75t_L g217 ( 
.A(n_72),
.Y(n_217)
);

INVx5_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx6_ASAP7_75t_SL g142 ( 
.A(n_75),
.Y(n_142)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_79),
.A2(n_89),
.B1(n_95),
.B2(n_102),
.Y(n_78)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_79),
.Y(n_153)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx4_ASAP7_75t_SL g81 ( 
.A(n_82),
.Y(n_81)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx5_ASAP7_75t_L g88 ( 
.A(n_84),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g253 ( 
.A(n_84),
.Y(n_253)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_85),
.Y(n_100)
);

BUFx3_ASAP7_75t_L g125 ( 
.A(n_85),
.Y(n_125)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_87),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx3_ASAP7_75t_L g246 ( 
.A(n_88),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_89),
.B(n_158),
.Y(n_157)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_89),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_89),
.A2(n_155),
.B1(n_281),
.B2(n_282),
.Y(n_280)
);

OR2x2_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_92),
.Y(n_89)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVxp67_ASAP7_75t_L g183 ( 
.A(n_95),
.Y(n_183)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVx8_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx4_ASAP7_75t_L g126 ( 
.A(n_100),
.Y(n_126)
);

INVx5_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

XNOR2xp5_ASAP7_75t_SL g304 ( 
.A(n_105),
.B(n_140),
.Y(n_304)
);

OAI21xp5_ASAP7_75t_SL g105 ( 
.A1(n_106),
.A2(n_128),
.B(n_134),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_SL g232 ( 
.A1(n_106),
.A2(n_134),
.B(n_233),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_106),
.A2(n_128),
.B1(n_220),
.B2(n_260),
.Y(n_292)
);

INVx1_ASAP7_75t_SL g106 ( 
.A(n_107),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_107),
.B(n_135),
.Y(n_223)
);

AND2x2_ASAP7_75t_L g107 ( 
.A(n_108),
.B(n_120),
.Y(n_107)
);

OAI22xp33_ASAP7_75t_L g108 ( 
.A1(n_109),
.A2(n_111),
.B1(n_114),
.B2(n_118),
.Y(n_108)
);

INVx4_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVx4_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

BUFx3_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

BUFx5_ASAP7_75t_L g127 ( 
.A(n_117),
.Y(n_127)
);

INVx4_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_120),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_SL g259 ( 
.A1(n_120),
.A2(n_223),
.B(n_260),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_121),
.A2(n_123),
.B1(n_126),
.B2(n_127),
.Y(n_120)
);

INVx5_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVx4_ASAP7_75t_L g243 ( 
.A(n_122),
.Y(n_243)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g270 ( 
.A(n_125),
.Y(n_270)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

INVx4_ASAP7_75t_L g136 ( 
.A(n_131),
.Y(n_136)
);

INVx4_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_135),
.B(n_139),
.Y(n_134)
);

INVx4_ASAP7_75t_SL g150 ( 
.A(n_137),
.Y(n_150)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_139),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_141),
.B(n_152),
.Y(n_140)
);

XOR2xp5_ASAP7_75t_L g298 ( 
.A(n_141),
.B(n_152),
.Y(n_298)
);

INVxp33_ASAP7_75t_L g296 ( 
.A(n_143),
.Y(n_296)
);

INVx3_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

BUFx2_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

NAND2xp33_ASAP7_75t_SL g147 ( 
.A(n_148),
.B(n_151),
.Y(n_147)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

AOI21xp5_ASAP7_75t_L g152 ( 
.A1(n_153),
.A2(n_154),
.B(n_157),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_154),
.A2(n_182),
.B1(n_183),
.B2(n_184),
.Y(n_181)
);

INVx4_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

INVx4_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

AOI21xp5_ASAP7_75t_L g274 ( 
.A1(n_157),
.A2(n_275),
.B(n_276),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_158),
.B(n_255),
.Y(n_254)
);

INVx8_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

BUFx8_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_161),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_192),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_164),
.A2(n_189),
.B1(n_190),
.B2(n_191),
.Y(n_163)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_164),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_165),
.A2(n_166),
.B1(n_180),
.B2(n_181),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

OAI32xp33_ASAP7_75t_L g166 ( 
.A1(n_167),
.A2(n_168),
.A3(n_170),
.B1(n_174),
.B2(n_176),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_168),
.A2(n_171),
.B1(n_197),
.B2(n_199),
.Y(n_196)
);

INVx8_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

INVx6_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

INVx3_ASAP7_75t_L g175 ( 
.A(n_172),
.Y(n_175)
);

INVx5_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g198 ( 
.A(n_173),
.Y(n_198)
);

INVx4_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

INVx3_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

AOI21xp5_ASAP7_75t_L g248 ( 
.A1(n_182),
.A2(n_249),
.B(n_254),
.Y(n_248)
);

INVxp67_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_189),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_193),
.A2(n_194),
.B1(n_213),
.B2(n_224),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

AOI21xp5_ASAP7_75t_L g194 ( 
.A1(n_195),
.A2(n_200),
.B(n_202),
.Y(n_194)
);

INVx4_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_204),
.B(n_212),
.Y(n_203)
);

INVx3_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

INVx4_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

INVx4_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

BUFx6f_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_213),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_SL g213 ( 
.A(n_214),
.B(n_219),
.Y(n_213)
);

INVx3_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_SL g219 ( 
.A1(n_220),
.A2(n_221),
.B(n_223),
.Y(n_219)
);

INVxp67_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

AO21x1_ASAP7_75t_L g227 ( 
.A1(n_228),
.A2(n_300),
.B(n_305),
.Y(n_227)
);

OAI21xp5_ASAP7_75t_SL g228 ( 
.A1(n_229),
.A2(n_287),
.B(n_299),
.Y(n_228)
);

AOI21xp5_ASAP7_75t_L g229 ( 
.A1(n_230),
.A2(n_263),
.B(n_286),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_231),
.B(n_247),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_231),
.B(n_247),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_232),
.B(n_238),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_232),
.A2(n_238),
.B1(n_239),
.B2(n_284),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_232),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_234),
.B(n_240),
.Y(n_239)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

INVx3_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

INVx4_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

HB1xp67_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_248),
.B(n_257),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_248),
.B(n_258),
.C(n_262),
.Y(n_288)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_249),
.Y(n_282)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

INVx6_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_255),
.Y(n_276)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_258),
.A2(n_259),
.B1(n_261),
.B2(n_262),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

OAI21xp5_ASAP7_75t_L g263 ( 
.A1(n_264),
.A2(n_279),
.B(n_285),
.Y(n_263)
);

AOI21xp5_ASAP7_75t_L g264 ( 
.A1(n_265),
.A2(n_273),
.B(n_278),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_266),
.B(n_272),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_267),
.B(n_271),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

INVx6_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

INVx4_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_SL g273 ( 
.A(n_274),
.B(n_277),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_274),
.B(n_277),
.Y(n_278)
);

INVxp67_ASAP7_75t_L g281 ( 
.A(n_275),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_280),
.B(n_283),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_280),
.B(n_283),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_288),
.B(n_289),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_288),
.B(n_289),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_L g289 ( 
.A(n_290),
.B(n_298),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_291),
.A2(n_292),
.B1(n_293),
.B2(n_294),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_292),
.B(n_293),
.C(n_298),
.Y(n_301)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_301),
.B(n_302),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_SL g305 ( 
.A(n_301),
.B(n_302),
.Y(n_305)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_304),
.Y(n_303)
);


endmodule