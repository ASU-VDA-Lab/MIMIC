module fake_jpeg_4618_n_332 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_332);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_332;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx4f_ASAP7_75t_SL g17 ( 
.A(n_11),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_15),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_4),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_7),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_8),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_10),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_35),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_36),
.B(n_41),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_17),
.Y(n_37)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_37),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_17),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_38),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_29),
.B(n_7),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_SL g51 ( 
.A(n_39),
.B(n_44),
.Y(n_51)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_35),
.Y(n_40)
);

INVx5_ASAP7_75t_L g67 ( 
.A(n_40),
.Y(n_67)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_35),
.Y(n_41)
);

INVx5_ASAP7_75t_L g42 ( 
.A(n_17),
.Y(n_42)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_42),
.Y(n_53)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_18),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_43),
.B(n_45),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_19),
.B(n_7),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_19),
.B(n_9),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g46 ( 
.A(n_20),
.B(n_0),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_46),
.B(n_0),
.Y(n_56)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_46),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_49),
.B(n_54),
.Y(n_71)
);

BUFx4f_ASAP7_75t_SL g50 ( 
.A(n_42),
.Y(n_50)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_50),
.Y(n_82)
);

AND2x2_ASAP7_75t_SL g52 ( 
.A(n_42),
.B(n_30),
.Y(n_52)
);

AND2x2_ASAP7_75t_L g99 ( 
.A(n_52),
.B(n_61),
.Y(n_99)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_42),
.Y(n_54)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_55),
.B(n_57),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_SL g91 ( 
.A(n_56),
.B(n_59),
.Y(n_91)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_46),
.Y(n_57)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_40),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_58),
.B(n_60),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_44),
.B(n_22),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_45),
.B(n_22),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_39),
.B(n_31),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_39),
.B(n_24),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_62),
.B(n_68),
.Y(n_87)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_43),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_63),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_43),
.A2(n_26),
.B1(n_29),
.B2(n_28),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_64),
.A2(n_17),
.B1(n_25),
.B2(n_33),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_37),
.B(n_24),
.Y(n_68)
);

CKINVDCx12_ASAP7_75t_R g69 ( 
.A(n_43),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_69),
.B(n_70),
.Y(n_94)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_41),
.Y(n_70)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_47),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_72),
.B(n_74),
.Y(n_101)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_47),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_52),
.A2(n_49),
.B1(n_57),
.B2(n_41),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_75),
.A2(n_77),
.B1(n_84),
.B2(n_53),
.Y(n_113)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_68),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_76),
.B(n_83),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_52),
.A2(n_28),
.B1(n_26),
.B2(n_36),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_L g78 ( 
.A1(n_52),
.A2(n_29),
.B1(n_26),
.B2(n_17),
.Y(n_78)
);

OAI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_78),
.A2(n_65),
.B1(n_25),
.B2(n_21),
.Y(n_107)
);

INVx6_ASAP7_75t_L g79 ( 
.A(n_67),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_79),
.A2(n_90),
.B1(n_65),
.B2(n_55),
.Y(n_117)
);

AND2x4_ASAP7_75t_L g81 ( 
.A(n_50),
.B(n_30),
.Y(n_81)
);

MAJx2_ASAP7_75t_L g119 ( 
.A(n_81),
.B(n_21),
.C(n_23),
.Y(n_119)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_67),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_48),
.A2(n_36),
.B1(n_70),
.B2(n_54),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_56),
.B(n_20),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_85),
.B(n_60),
.Y(n_111)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_48),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_88),
.B(n_89),
.Y(n_124)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_61),
.Y(n_89)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_50),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_92),
.B(n_93),
.Y(n_127)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_50),
.Y(n_93)
);

AOI21xp5_ASAP7_75t_L g95 ( 
.A1(n_51),
.A2(n_30),
.B(n_21),
.Y(n_95)
);

XNOR2xp5_ASAP7_75t_L g104 ( 
.A(n_95),
.B(n_25),
.Y(n_104)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_62),
.Y(n_96)
);

INVx13_ASAP7_75t_L g112 ( 
.A(n_96),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_55),
.Y(n_97)
);

INVx6_ASAP7_75t_L g109 ( 
.A(n_97),
.Y(n_109)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_59),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_98),
.B(n_58),
.Y(n_118)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_80),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_100),
.B(n_102),
.Y(n_136)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_80),
.Y(n_102)
);

CKINVDCx16_ASAP7_75t_R g103 ( 
.A(n_94),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_103),
.B(n_105),
.Y(n_144)
);

AND2x2_ASAP7_75t_L g128 ( 
.A(n_104),
.B(n_113),
.Y(n_128)
);

CKINVDCx16_ASAP7_75t_R g105 ( 
.A(n_94),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_86),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_106),
.B(n_118),
.Y(n_146)
);

CKINVDCx16_ASAP7_75t_R g152 ( 
.A(n_107),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_75),
.B(n_69),
.C(n_53),
.Y(n_108)
);

XNOR2xp5_ASAP7_75t_L g142 ( 
.A(n_108),
.B(n_37),
.Y(n_142)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_81),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_110),
.B(n_115),
.Y(n_149)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_111),
.Y(n_147)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_81),
.Y(n_114)
);

INVx3_ASAP7_75t_L g137 ( 
.A(n_114),
.Y(n_137)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_97),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g135 ( 
.A1(n_117),
.A2(n_121),
.B1(n_79),
.B2(n_76),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_SL g156 ( 
.A1(n_119),
.A2(n_31),
.B(n_27),
.Y(n_156)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_81),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_120),
.B(n_126),
.Y(n_150)
);

AOI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_81),
.A2(n_88),
.B1(n_89),
.B2(n_96),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_99),
.A2(n_58),
.B1(n_65),
.B2(n_51),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_122),
.A2(n_123),
.B1(n_84),
.B2(n_87),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_99),
.A2(n_33),
.B1(n_23),
.B2(n_27),
.Y(n_123)
);

INVxp67_ASAP7_75t_SL g125 ( 
.A(n_79),
.Y(n_125)
);

INVx2_ASAP7_75t_R g158 ( 
.A(n_125),
.Y(n_158)
);

INVx1_ASAP7_75t_SL g126 ( 
.A(n_91),
.Y(n_126)
);

OR2x4_ASAP7_75t_L g129 ( 
.A(n_110),
.B(n_99),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_SL g159 ( 
.A1(n_129),
.A2(n_132),
.B(n_133),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_106),
.B(n_100),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_130),
.B(n_134),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_120),
.A2(n_95),
.B1(n_74),
.B2(n_72),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_131),
.A2(n_140),
.B1(n_145),
.B2(n_118),
.Y(n_166)
);

AOI21xp5_ASAP7_75t_L g132 ( 
.A1(n_108),
.A2(n_77),
.B(n_71),
.Y(n_132)
);

AOI21xp5_ASAP7_75t_L g133 ( 
.A1(n_113),
.A2(n_71),
.B(n_99),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_102),
.B(n_86),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g188 ( 
.A1(n_135),
.A2(n_138),
.B1(n_34),
.B2(n_109),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_122),
.B(n_87),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_139),
.B(n_143),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_104),
.A2(n_83),
.B1(n_98),
.B2(n_91),
.Y(n_140)
);

OAI211xp5_ASAP7_75t_L g141 ( 
.A1(n_119),
.A2(n_85),
.B(n_33),
.C(n_23),
.Y(n_141)
);

FAx1_ASAP7_75t_SL g179 ( 
.A(n_141),
.B(n_154),
.CI(n_156),
.CON(n_179),
.SN(n_179)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_142),
.B(n_155),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_126),
.B(n_92),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_124),
.A2(n_73),
.B1(n_93),
.B2(n_82),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_127),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_148),
.B(n_151),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_127),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_112),
.B(n_97),
.Y(n_153)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_153),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_124),
.B(n_73),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_L g155 ( 
.A(n_123),
.B(n_37),
.Y(n_155)
);

INVx5_ASAP7_75t_L g157 ( 
.A(n_115),
.Y(n_157)
);

INVxp67_ASAP7_75t_SL g168 ( 
.A(n_157),
.Y(n_168)
);

INVx13_ASAP7_75t_L g160 ( 
.A(n_158),
.Y(n_160)
);

INVx13_ASAP7_75t_L g200 ( 
.A(n_160),
.Y(n_200)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_130),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_162),
.B(n_171),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_129),
.B(n_119),
.C(n_103),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_163),
.B(n_180),
.C(n_184),
.Y(n_195)
);

INVx13_ASAP7_75t_L g165 ( 
.A(n_158),
.Y(n_165)
);

CKINVDCx16_ASAP7_75t_R g207 ( 
.A(n_165),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_L g215 ( 
.A1(n_166),
.A2(n_172),
.B1(n_32),
.B2(n_18),
.Y(n_215)
);

OAI21xp33_ASAP7_75t_L g167 ( 
.A1(n_139),
.A2(n_105),
.B(n_112),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_167),
.B(n_18),
.Y(n_208)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_157),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_170),
.Y(n_219)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_146),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_128),
.A2(n_101),
.B1(n_111),
.B2(n_116),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_SL g173 ( 
.A(n_136),
.B(n_101),
.Y(n_173)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_173),
.Y(n_206)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_146),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_175),
.B(n_176),
.Y(n_216)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_134),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_153),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_177),
.B(n_191),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_133),
.B(n_132),
.C(n_142),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_148),
.B(n_112),
.Y(n_181)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_181),
.Y(n_218)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_158),
.Y(n_182)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_182),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_138),
.A2(n_116),
.B1(n_82),
.B2(n_109),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_183),
.A2(n_188),
.B1(n_189),
.B2(n_152),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_128),
.B(n_63),
.C(n_38),
.Y(n_184)
);

INVxp67_ASAP7_75t_SL g185 ( 
.A(n_145),
.Y(n_185)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_185),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_151),
.B(n_109),
.Y(n_186)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_186),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_136),
.B(n_147),
.Y(n_187)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_187),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_152),
.A2(n_34),
.B1(n_38),
.B2(n_66),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_147),
.B(n_11),
.Y(n_190)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_190),
.Y(n_213)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_143),
.Y(n_191)
);

XOR2xp5_ASAP7_75t_L g192 ( 
.A(n_180),
.B(n_131),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_192),
.B(n_203),
.Y(n_241)
);

AOI21xp33_ASAP7_75t_L g193 ( 
.A1(n_159),
.A2(n_150),
.B(n_156),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_L g222 ( 
.A1(n_193),
.A2(n_205),
.B(n_209),
.Y(n_222)
);

AND2x2_ASAP7_75t_L g194 ( 
.A(n_163),
.B(n_155),
.Y(n_194)
);

AOI21xp5_ASAP7_75t_L g234 ( 
.A1(n_194),
.A2(n_198),
.B(n_202),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_L g224 ( 
.A1(n_196),
.A2(n_166),
.B1(n_172),
.B2(n_171),
.Y(n_224)
);

OAI21xp5_ASAP7_75t_L g198 ( 
.A1(n_159),
.A2(n_149),
.B(n_128),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_183),
.A2(n_140),
.B1(n_137),
.B2(n_144),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_201),
.A2(n_175),
.B1(n_184),
.B2(n_191),
.Y(n_227)
);

OAI21xp5_ASAP7_75t_SL g202 ( 
.A1(n_174),
.A2(n_144),
.B(n_154),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_L g203 ( 
.A1(n_174),
.A2(n_137),
.B(n_18),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_SL g205 ( 
.A1(n_161),
.A2(n_63),
.B(n_38),
.Y(n_205)
);

AND2x2_ASAP7_75t_L g235 ( 
.A(n_208),
.B(n_169),
.Y(n_235)
);

OAI21xp5_ASAP7_75t_SL g209 ( 
.A1(n_161),
.A2(n_63),
.B(n_66),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_L g212 ( 
.A(n_169),
.B(n_18),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_212),
.B(n_189),
.Y(n_243)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_178),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_SL g225 ( 
.A(n_214),
.B(n_220),
.Y(n_225)
);

NOR3xp33_ASAP7_75t_L g232 ( 
.A(n_215),
.B(n_164),
.C(n_177),
.Y(n_232)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_168),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_217),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_221),
.B(n_226),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_217),
.B(n_162),
.Y(n_223)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_223),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_224),
.A2(n_227),
.B1(n_233),
.B2(n_235),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_219),
.Y(n_226)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_204),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_SL g267 ( 
.A(n_228),
.B(n_230),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_204),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_229),
.Y(n_250)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_216),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_216),
.Y(n_231)
);

OAI21xp5_ASAP7_75t_SL g253 ( 
.A1(n_231),
.A2(n_238),
.B(n_240),
.Y(n_253)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_232),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_L g233 ( 
.A1(n_199),
.A2(n_176),
.B1(n_182),
.B2(n_179),
.Y(n_233)
);

CKINVDCx16_ASAP7_75t_R g236 ( 
.A(n_209),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_SL g261 ( 
.A(n_236),
.B(n_237),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_SL g237 ( 
.A(n_206),
.B(n_179),
.Y(n_237)
);

INVxp67_ASAP7_75t_L g238 ( 
.A(n_205),
.Y(n_238)
);

OAI21xp5_ASAP7_75t_L g239 ( 
.A1(n_202),
.A2(n_179),
.B(n_165),
.Y(n_239)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_239),
.B(n_242),
.Y(n_255)
);

AND2x6_ASAP7_75t_L g240 ( 
.A(n_198),
.B(n_160),
.Y(n_240)
);

OAI21xp5_ASAP7_75t_L g242 ( 
.A1(n_199),
.A2(n_201),
.B(n_207),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_243),
.B(n_227),
.Y(n_262)
);

INVxp67_ASAP7_75t_SL g244 ( 
.A(n_220),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_L g254 ( 
.A1(n_244),
.A2(n_197),
.B1(n_210),
.B2(n_196),
.Y(n_254)
);

NOR2x1_ASAP7_75t_L g245 ( 
.A(n_211),
.B(n_66),
.Y(n_245)
);

OAI21xp5_ASAP7_75t_L g256 ( 
.A1(n_245),
.A2(n_213),
.B(n_197),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_203),
.A2(n_170),
.B1(n_32),
.B2(n_2),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_246),
.A2(n_214),
.B1(n_211),
.B2(n_218),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_241),
.B(n_195),
.C(n_192),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_247),
.B(n_248),
.C(n_251),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_241),
.B(n_195),
.C(n_194),
.Y(n_248)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_249),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_234),
.B(n_235),
.C(n_221),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_254),
.B(n_225),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_256),
.B(n_0),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_234),
.B(n_235),
.C(n_230),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_257),
.B(n_259),
.C(n_266),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_238),
.A2(n_194),
.B1(n_210),
.B2(n_208),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_258),
.A2(n_264),
.B1(n_32),
.B2(n_1),
.Y(n_276)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_240),
.B(n_212),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_262),
.B(n_245),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_242),
.A2(n_200),
.B1(n_213),
.B2(n_32),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_239),
.B(n_200),
.Y(n_266)
);

OAI21xp5_ASAP7_75t_L g268 ( 
.A1(n_253),
.A2(n_231),
.B(n_223),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_268),
.A2(n_272),
.B1(n_276),
.B2(n_281),
.Y(n_296)
);

OA21x2_ASAP7_75t_SL g271 ( 
.A1(n_262),
.A2(n_222),
.B(n_243),
.Y(n_271)
);

OAI21xp33_ASAP7_75t_L g297 ( 
.A1(n_271),
.A2(n_249),
.B(n_13),
.Y(n_297)
);

OAI21xp5_ASAP7_75t_L g272 ( 
.A1(n_253),
.A2(n_246),
.B(n_222),
.Y(n_272)
);

OAI21xp5_ASAP7_75t_L g291 ( 
.A1(n_274),
.A2(n_265),
.B(n_273),
.Y(n_291)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_275),
.B(n_278),
.Y(n_288)
);

A2O1A1Ixp33_ASAP7_75t_SL g277 ( 
.A1(n_263),
.A2(n_0),
.B(n_1),
.C(n_2),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_277),
.A2(n_280),
.B1(n_264),
.B2(n_250),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_251),
.B(n_9),
.Y(n_278)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_279),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_257),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_252),
.A2(n_10),
.B1(n_15),
.B2(n_14),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_260),
.B(n_9),
.Y(n_282)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_282),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_261),
.B(n_11),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_SL g293 ( 
.A(n_283),
.B(n_256),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_248),
.B(n_2),
.C(n_3),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_284),
.B(n_280),
.C(n_272),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_270),
.A2(n_252),
.B1(n_258),
.B2(n_259),
.Y(n_285)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_285),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_286),
.B(n_290),
.C(n_294),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_287),
.B(n_275),
.Y(n_300)
);

XOR2xp5_ASAP7_75t_L g289 ( 
.A(n_273),
.B(n_247),
.Y(n_289)
);

XOR2xp5_ASAP7_75t_L g304 ( 
.A(n_289),
.B(n_277),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_269),
.B(n_255),
.C(n_267),
.Y(n_290)
);

AOI21xp5_ASAP7_75t_L g310 ( 
.A1(n_291),
.A2(n_15),
.B(n_16),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_SL g299 ( 
.A(n_293),
.B(n_278),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_269),
.B(n_255),
.C(n_266),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_L g307 ( 
.A(n_297),
.B(n_14),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_268),
.B(n_3),
.C(n_4),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_298),
.B(n_3),
.C(n_5),
.Y(n_305)
);

OAI21xp5_ASAP7_75t_SL g319 ( 
.A1(n_299),
.A2(n_306),
.B(n_309),
.Y(n_319)
);

AOI21xp5_ASAP7_75t_L g317 ( 
.A1(n_300),
.A2(n_302),
.B(n_305),
.Y(n_317)
);

OAI21xp5_ASAP7_75t_L g302 ( 
.A1(n_296),
.A2(n_284),
.B(n_277),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_SL g303 ( 
.A1(n_296),
.A2(n_277),
.B1(n_5),
.B2(n_6),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_303),
.B(n_307),
.Y(n_314)
);

XOR2xp5_ASAP7_75t_L g312 ( 
.A(n_304),
.B(n_310),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_295),
.B(n_13),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_292),
.B(n_5),
.Y(n_309)
);

AOI21x1_ASAP7_75t_L g311 ( 
.A1(n_304),
.A2(n_302),
.B(n_285),
.Y(n_311)
);

OAI31xp33_ASAP7_75t_L g323 ( 
.A1(n_311),
.A2(n_315),
.A3(n_288),
.B(n_16),
.Y(n_323)
);

XNOR2xp5_ASAP7_75t_L g313 ( 
.A(n_301),
.B(n_290),
.Y(n_313)
);

XOR2xp5_ASAP7_75t_L g325 ( 
.A(n_313),
.B(n_6),
.Y(n_325)
);

AO21x1_ASAP7_75t_L g315 ( 
.A1(n_308),
.A2(n_291),
.B(n_286),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_307),
.B(n_298),
.Y(n_316)
);

OAI21xp5_ASAP7_75t_L g321 ( 
.A1(n_316),
.A2(n_318),
.B(n_305),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_303),
.B(n_288),
.Y(n_318)
);

NAND4xp25_ASAP7_75t_L g320 ( 
.A(n_315),
.B(n_301),
.C(n_289),
.D(n_294),
.Y(n_320)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_320),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_321),
.B(n_325),
.Y(n_327)
);

INVxp67_ASAP7_75t_L g322 ( 
.A(n_317),
.Y(n_322)
);

OAI22xp33_ASAP7_75t_L g326 ( 
.A1(n_322),
.A2(n_323),
.B1(n_324),
.B2(n_314),
.Y(n_326)
);

NOR2xp67_ASAP7_75t_L g324 ( 
.A(n_313),
.B(n_16),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_326),
.B(n_322),
.Y(n_329)
);

OAI22xp5_ASAP7_75t_L g330 ( 
.A1(n_329),
.A2(n_328),
.B1(n_327),
.B2(n_312),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_330),
.B(n_312),
.C(n_319),
.Y(n_331)
);

XNOR2xp5_ASAP7_75t_L g332 ( 
.A(n_331),
.B(n_6),
.Y(n_332)
);


endmodule