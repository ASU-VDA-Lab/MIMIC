module fake_netlist_6_1734_n_868 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_161, n_68, n_166, n_28, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_178, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_180, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_181, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_175, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_104, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_173, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_171, n_31, n_57, n_169, n_53, n_51, n_44, n_56, n_868);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_161;
input n_68;
input n_166;
input n_28;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_178;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_181;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_175;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_104;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_173;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_171;
input n_31;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_868;

wire n_591;
wire n_435;
wire n_793;
wire n_326;
wire n_801;
wire n_256;
wire n_853;
wire n_440;
wire n_587;
wire n_695;
wire n_507;
wire n_580;
wire n_762;
wire n_209;
wire n_367;
wire n_465;
wire n_680;
wire n_741;
wire n_760;
wire n_590;
wire n_625;
wire n_661;
wire n_223;
wire n_278;
wire n_341;
wire n_362;
wire n_226;
wire n_828;
wire n_208;
wire n_462;
wire n_607;
wire n_671;
wire n_726;
wire n_316;
wire n_419;
wire n_304;
wire n_212;
wire n_700;
wire n_694;
wire n_740;
wire n_578;
wire n_703;
wire n_365;
wire n_384;
wire n_297;
wire n_627;
wire n_595;
wire n_524;
wire n_342;
wire n_820;
wire n_783;
wire n_725;
wire n_358;
wire n_751;
wire n_449;
wire n_749;
wire n_798;
wire n_188;
wire n_310;
wire n_509;
wire n_186;
wire n_245;
wire n_368;
wire n_575;
wire n_677;
wire n_805;
wire n_396;
wire n_495;
wire n_815;
wire n_350;
wire n_585;
wire n_732;
wire n_568;
wire n_392;
wire n_840;
wire n_442;
wire n_480;
wire n_724;
wire n_382;
wire n_673;
wire n_628;
wire n_557;
wire n_823;
wire n_349;
wire n_643;
wire n_233;
wire n_617;
wire n_698;
wire n_845;
wire n_255;
wire n_807;
wire n_739;
wire n_284;
wire n_400;
wire n_337;
wire n_865;
wire n_214;
wire n_485;
wire n_443;
wire n_246;
wire n_768;
wire n_471;
wire n_289;
wire n_421;
wire n_781;
wire n_424;
wire n_789;
wire n_615;
wire n_182;
wire n_238;
wire n_573;
wire n_769;
wire n_202;
wire n_320;
wire n_639;
wire n_676;
wire n_327;
wire n_794;
wire n_727;
wire n_369;
wire n_597;
wire n_685;
wire n_280;
wire n_287;
wire n_832;
wire n_353;
wire n_610;
wire n_555;
wire n_389;
wire n_814;
wire n_415;
wire n_830;
wire n_230;
wire n_605;
wire n_461;
wire n_383;
wire n_826;
wire n_669;
wire n_200;
wire n_447;
wire n_198;
wire n_300;
wire n_222;
wire n_248;
wire n_517;
wire n_718;
wire n_747;
wire n_852;
wire n_667;
wire n_229;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_621;
wire n_305;
wire n_721;
wire n_750;
wire n_532;
wire n_742;
wire n_535;
wire n_691;
wire n_250;
wire n_372;
wire n_468;
wire n_544;
wire n_504;
wire n_314;
wire n_378;
wire n_413;
wire n_377;
wire n_791;
wire n_183;
wire n_510;
wire n_837;
wire n_836;
wire n_863;
wire n_375;
wire n_601;
wire n_338;
wire n_522;
wire n_466;
wire n_704;
wire n_748;
wire n_506;
wire n_763;
wire n_360;
wire n_603;
wire n_235;
wire n_536;
wire n_866;
wire n_622;
wire n_191;
wire n_340;
wire n_710;
wire n_387;
wire n_452;
wire n_616;
wire n_658;
wire n_744;
wire n_344;
wire n_581;
wire n_428;
wire n_785;
wire n_761;
wire n_746;
wire n_609;
wire n_765;
wire n_432;
wire n_641;
wire n_822;
wire n_693;
wire n_631;
wire n_516;
wire n_758;
wire n_525;
wire n_720;
wire n_842;
wire n_611;
wire n_491;
wire n_656;
wire n_772;
wire n_843;
wire n_797;
wire n_666;
wire n_371;
wire n_795;
wire n_770;
wire n_567;
wire n_189;
wire n_738;
wire n_405;
wire n_213;
wire n_538;
wire n_294;
wire n_302;
wire n_499;
wire n_380;
wire n_838;
wire n_705;
wire n_647;
wire n_197;
wire n_343;
wire n_844;
wire n_448;
wire n_494;
wire n_539;
wire n_493;
wire n_397;
wire n_614;
wire n_529;
wire n_445;
wire n_425;
wire n_684;
wire n_454;
wire n_218;
wire n_638;
wire n_234;
wire n_486;
wire n_381;
wire n_236;
wire n_653;
wire n_752;
wire n_713;
wire n_648;
wire n_657;
wire n_576;
wire n_472;
wire n_270;
wire n_239;
wire n_414;
wire n_563;
wire n_782;
wire n_490;
wire n_803;
wire n_290;
wire n_220;
wire n_809;
wire n_224;
wire n_839;
wire n_734;
wire n_708;
wire n_196;
wire n_402;
wire n_352;
wire n_668;
wire n_478;
wire n_626;
wire n_574;
wire n_779;
wire n_800;
wire n_460;
wire n_854;
wire n_417;
wire n_446;
wire n_498;
wire n_662;
wire n_374;
wire n_659;
wire n_709;
wire n_366;
wire n_777;
wire n_407;
wire n_450;
wire n_808;
wire n_867;
wire n_272;
wire n_526;
wire n_185;
wire n_712;
wire n_348;
wire n_711;
wire n_579;
wire n_376;
wire n_390;
wire n_473;
wire n_293;
wire n_334;
wire n_559;
wire n_370;
wire n_458;
wire n_232;
wire n_650;
wire n_717;
wire n_330;
wire n_771;
wire n_470;
wire n_475;
wire n_298;
wire n_492;
wire n_281;
wire n_258;
wire n_551;
wire n_699;
wire n_456;
wire n_564;
wire n_265;
wire n_260;
wire n_313;
wire n_451;
wire n_624;
wire n_824;
wire n_279;
wire n_686;
wire n_796;
wire n_252;
wire n_757;
wire n_228;
wire n_565;
wire n_594;
wire n_719;
wire n_356;
wire n_577;
wire n_184;
wire n_552;
wire n_619;
wire n_216;
wire n_455;
wire n_521;
wire n_363;
wire n_572;
wire n_395;
wire n_813;
wire n_592;
wire n_745;
wire n_654;
wire n_323;
wire n_829;
wire n_606;
wire n_393;
wire n_818;
wire n_411;
wire n_503;
wire n_716;
wire n_623;
wire n_599;
wire n_513;
wire n_855;
wire n_776;
wire n_321;
wire n_645;
wire n_331;
wire n_227;
wire n_570;
wire n_731;
wire n_859;
wire n_406;
wire n_483;
wire n_735;
wire n_204;
wire n_482;
wire n_755;
wire n_474;
wire n_527;
wire n_261;
wire n_608;
wire n_620;
wire n_420;
wire n_683;
wire n_630;
wire n_312;
wire n_394;
wire n_519;
wire n_541;
wire n_512;
wire n_292;
wire n_307;
wire n_469;
wire n_433;
wire n_500;
wire n_792;
wire n_476;
wire n_714;
wire n_291;
wire n_219;
wire n_543;
wire n_357;
wire n_264;
wire n_263;
wire n_589;
wire n_860;
wire n_481;
wire n_788;
wire n_819;
wire n_821;
wire n_325;
wire n_767;
wire n_804;
wire n_329;
wire n_464;
wire n_600;
wire n_831;
wire n_802;
wire n_561;
wire n_477;
wire n_549;
wire n_533;
wire n_408;
wire n_806;
wire n_864;
wire n_237;
wire n_584;
wire n_244;
wire n_399;
wire n_243;
wire n_548;
wire n_282;
wire n_436;
wire n_833;
wire n_211;
wire n_523;
wire n_322;
wire n_707;
wire n_345;
wire n_409;
wire n_231;
wire n_354;
wire n_689;
wire n_799;
wire n_505;
wire n_240;
wire n_756;
wire n_319;
wire n_547;
wire n_537;
wire n_273;
wire n_558;
wire n_810;
wire n_635;
wire n_787;
wire n_311;
wire n_403;
wire n_723;
wire n_253;
wire n_634;
wire n_583;
wire n_596;
wire n_546;
wire n_562;
wire n_249;
wire n_201;
wire n_386;
wire n_764;
wire n_556;
wire n_692;
wire n_733;
wire n_754;
wire n_487;
wire n_550;
wire n_241;
wire n_275;
wire n_553;
wire n_652;
wire n_849;
wire n_560;
wire n_753;
wire n_642;
wire n_276;
wire n_569;
wire n_441;
wire n_221;
wire n_811;
wire n_444;
wire n_586;
wire n_423;
wire n_737;
wire n_318;
wire n_303;
wire n_511;
wire n_715;
wire n_467;
wire n_306;
wire n_193;
wire n_269;
wire n_359;
wire n_346;
wire n_416;
wire n_530;
wire n_277;
wire n_520;
wire n_418;
wire n_618;
wire n_790;
wire n_582;
wire n_199;
wire n_266;
wire n_296;
wire n_861;
wire n_674;
wire n_857;
wire n_775;
wire n_571;
wire n_268;
wire n_404;
wire n_271;
wire n_651;
wire n_439;
wire n_217;
wire n_210;
wire n_299;
wire n_518;
wire n_206;
wire n_679;
wire n_453;
wire n_612;
wire n_633;
wire n_665;
wire n_333;
wire n_588;
wire n_215;
wire n_247;
wire n_225;
wire n_308;
wire n_309;
wire n_759;
wire n_355;
wire n_426;
wire n_317;
wire n_632;
wire n_702;
wire n_431;
wire n_347;
wire n_812;
wire n_459;
wire n_502;
wire n_328;
wire n_672;
wire n_534;
wire n_488;
wire n_429;
wire n_373;
wire n_195;
wire n_285;
wire n_497;
wire n_780;
wire n_773;
wire n_675;
wire n_257;
wire n_730;
wire n_655;
wire n_706;
wire n_786;
wire n_670;
wire n_203;
wire n_286;
wire n_254;
wire n_207;
wire n_834;
wire n_242;
wire n_835;
wire n_690;
wire n_850;
wire n_401;
wire n_324;
wire n_766;
wire n_743;
wire n_816;
wire n_335;
wire n_430;
wire n_463;
wire n_545;
wire n_489;
wire n_205;
wire n_604;
wire n_848;
wire n_251;
wire n_301;
wire n_274;
wire n_636;
wire n_825;
wire n_728;
wire n_681;
wire n_729;
wire n_774;
wire n_412;
wire n_640;
wire n_660;
wire n_267;
wire n_438;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_515;
wire n_288;
wire n_427;
wire n_479;
wire n_496;
wire n_598;
wire n_422;
wire n_696;
wire n_688;
wire n_722;
wire n_862;
wire n_351;
wire n_437;
wire n_259;
wire n_540;
wire n_593;
wire n_514;
wire n_646;
wire n_528;
wire n_391;
wire n_457;
wire n_697;
wire n_687;
wire n_364;
wire n_637;
wire n_295;
wire n_385;
wire n_701;
wire n_817;
wire n_629;
wire n_388;
wire n_190;
wire n_858;
wire n_262;
wire n_484;
wire n_613;
wire n_736;
wire n_187;
wire n_846;
wire n_501;
wire n_841;
wire n_531;
wire n_827;
wire n_361;
wire n_508;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_332;
wire n_336;
wire n_398;
wire n_410;
wire n_566;
wire n_554;
wire n_602;
wire n_194;
wire n_664;
wire n_678;
wire n_192;
wire n_649;
wire n_283;

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_132),
.Y(n_182)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_168),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_91),
.Y(n_184)
);

INVxp33_ASAP7_75t_L g185 ( 
.A(n_73),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_118),
.B(n_105),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_124),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_167),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_61),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_71),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_153),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_150),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_100),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_62),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_130),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_48),
.Y(n_196)
);

HB1xp67_ASAP7_75t_L g197 ( 
.A(n_126),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_31),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_135),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_46),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_9),
.Y(n_201)
);

HB1xp67_ASAP7_75t_L g202 ( 
.A(n_159),
.Y(n_202)
);

BUFx10_ASAP7_75t_L g203 ( 
.A(n_55),
.Y(n_203)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_87),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_154),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_161),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_121),
.Y(n_207)
);

INVx1_ASAP7_75t_SL g208 ( 
.A(n_165),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_25),
.Y(n_209)
);

INVx2_ASAP7_75t_SL g210 ( 
.A(n_96),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_14),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_157),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_156),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_15),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_32),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_173),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_175),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_111),
.Y(n_218)
);

INVx1_ASAP7_75t_SL g219 ( 
.A(n_30),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_60),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_37),
.Y(n_221)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_178),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_14),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_131),
.Y(n_224)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_74),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_70),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_149),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_108),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_58),
.Y(n_229)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_57),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_64),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_164),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_5),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_11),
.Y(n_234)
);

BUFx3_ASAP7_75t_L g235 ( 
.A(n_117),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_125),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_53),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_13),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_170),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_177),
.Y(n_240)
);

BUFx2_ASAP7_75t_L g241 ( 
.A(n_16),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_176),
.Y(n_242)
);

INVxp67_ASAP7_75t_L g243 ( 
.A(n_20),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_113),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_63),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_76),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_54),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_49),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_102),
.Y(n_249)
);

BUFx6f_ASAP7_75t_L g250 ( 
.A(n_109),
.Y(n_250)
);

INVx1_ASAP7_75t_SL g251 ( 
.A(n_110),
.Y(n_251)
);

AND2x2_ASAP7_75t_L g252 ( 
.A(n_241),
.B(n_0),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_211),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_214),
.Y(n_254)
);

BUFx6f_ASAP7_75t_L g255 ( 
.A(n_250),
.Y(n_255)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_233),
.Y(n_256)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_234),
.Y(n_257)
);

OA21x2_ASAP7_75t_L g258 ( 
.A1(n_183),
.A2(n_0),
.B(n_1),
.Y(n_258)
);

OA21x2_ASAP7_75t_L g259 ( 
.A1(n_183),
.A2(n_1),
.B(n_2),
.Y(n_259)
);

NOR2x1_ASAP7_75t_L g260 ( 
.A(n_235),
.B(n_23),
.Y(n_260)
);

BUFx6f_ASAP7_75t_L g261 ( 
.A(n_250),
.Y(n_261)
);

BUFx3_ASAP7_75t_L g262 ( 
.A(n_235),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_210),
.B(n_2),
.Y(n_263)
);

BUFx2_ASAP7_75t_L g264 ( 
.A(n_223),
.Y(n_264)
);

BUFx2_ASAP7_75t_L g265 ( 
.A(n_238),
.Y(n_265)
);

INVx5_ASAP7_75t_L g266 ( 
.A(n_250),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_204),
.Y(n_267)
);

INVx4_ASAP7_75t_L g268 ( 
.A(n_250),
.Y(n_268)
);

OA21x2_ASAP7_75t_L g269 ( 
.A1(n_204),
.A2(n_3),
.B(n_4),
.Y(n_269)
);

BUFx6f_ASAP7_75t_L g270 ( 
.A(n_222),
.Y(n_270)
);

BUFx2_ASAP7_75t_L g271 ( 
.A(n_201),
.Y(n_271)
);

AND2x6_ASAP7_75t_L g272 ( 
.A(n_222),
.B(n_24),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_225),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_187),
.Y(n_274)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_225),
.Y(n_275)
);

AND2x4_ASAP7_75t_L g276 ( 
.A(n_230),
.B(n_26),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_230),
.Y(n_277)
);

INVx3_ASAP7_75t_L g278 ( 
.A(n_203),
.Y(n_278)
);

BUFx6f_ASAP7_75t_L g279 ( 
.A(n_189),
.Y(n_279)
);

INVx4_ASAP7_75t_L g280 ( 
.A(n_203),
.Y(n_280)
);

OAI21x1_ASAP7_75t_L g281 ( 
.A1(n_191),
.A2(n_3),
.B(n_4),
.Y(n_281)
);

CKINVDCx16_ASAP7_75t_R g282 ( 
.A(n_242),
.Y(n_282)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_192),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_185),
.B(n_5),
.Y(n_284)
);

OA21x2_ASAP7_75t_L g285 ( 
.A1(n_243),
.A2(n_6),
.B(n_7),
.Y(n_285)
);

BUFx3_ASAP7_75t_L g286 ( 
.A(n_203),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_196),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_199),
.Y(n_288)
);

BUFx8_ASAP7_75t_SL g289 ( 
.A(n_201),
.Y(n_289)
);

BUFx12f_ASAP7_75t_L g290 ( 
.A(n_188),
.Y(n_290)
);

NAND2xp33_ASAP7_75t_L g291 ( 
.A(n_185),
.B(n_6),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_197),
.B(n_7),
.Y(n_292)
);

BUFx2_ASAP7_75t_L g293 ( 
.A(n_242),
.Y(n_293)
);

BUFx6f_ASAP7_75t_L g294 ( 
.A(n_200),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_212),
.Y(n_295)
);

BUFx6f_ASAP7_75t_L g296 ( 
.A(n_217),
.Y(n_296)
);

INVx2_ASAP7_75t_L g297 ( 
.A(n_220),
.Y(n_297)
);

BUFx6f_ASAP7_75t_L g298 ( 
.A(n_224),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_202),
.B(n_8),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_188),
.Y(n_300)
);

OAI21x1_ASAP7_75t_L g301 ( 
.A1(n_232),
.A2(n_240),
.B(n_237),
.Y(n_301)
);

INVx3_ASAP7_75t_L g302 ( 
.A(n_244),
.Y(n_302)
);

AO21x2_ASAP7_75t_L g303 ( 
.A1(n_281),
.A2(n_248),
.B(n_247),
.Y(n_303)
);

INVxp33_ASAP7_75t_SL g304 ( 
.A(n_300),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_SL g305 ( 
.A(n_280),
.B(n_245),
.Y(n_305)
);

BUFx10_ASAP7_75t_L g306 ( 
.A(n_284),
.Y(n_306)
);

AO21x2_ASAP7_75t_L g307 ( 
.A1(n_281),
.A2(n_249),
.B(n_186),
.Y(n_307)
);

INVx2_ASAP7_75t_L g308 ( 
.A(n_270),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_SL g309 ( 
.A(n_280),
.B(n_245),
.Y(n_309)
);

BUFx6f_ASAP7_75t_SL g310 ( 
.A(n_286),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_280),
.B(n_208),
.Y(n_311)
);

INVx5_ASAP7_75t_L g312 ( 
.A(n_272),
.Y(n_312)
);

INVx2_ASAP7_75t_L g313 ( 
.A(n_270),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_SL g314 ( 
.A(n_278),
.B(n_246),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_278),
.B(n_300),
.Y(n_315)
);

OR2x6_ASAP7_75t_L g316 ( 
.A(n_290),
.B(n_246),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_283),
.Y(n_317)
);

INVx2_ASAP7_75t_L g318 ( 
.A(n_270),
.Y(n_318)
);

INVx2_ASAP7_75t_L g319 ( 
.A(n_270),
.Y(n_319)
);

INVx2_ASAP7_75t_L g320 ( 
.A(n_270),
.Y(n_320)
);

OR2x6_ASAP7_75t_L g321 ( 
.A(n_290),
.B(n_182),
.Y(n_321)
);

INVx2_ASAP7_75t_L g322 ( 
.A(n_255),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_289),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_SL g324 ( 
.A(n_278),
.B(n_219),
.Y(n_324)
);

BUFx10_ASAP7_75t_L g325 ( 
.A(n_276),
.Y(n_325)
);

INVx8_ASAP7_75t_L g326 ( 
.A(n_266),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_SL g327 ( 
.A(n_276),
.B(n_251),
.Y(n_327)
);

NOR2x1p5_ASAP7_75t_L g328 ( 
.A(n_286),
.B(n_184),
.Y(n_328)
);

INVx2_ASAP7_75t_SL g329 ( 
.A(n_264),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_283),
.Y(n_330)
);

INVx2_ASAP7_75t_L g331 ( 
.A(n_255),
.Y(n_331)
);

INVx1_ASAP7_75t_SL g332 ( 
.A(n_293),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_262),
.B(n_239),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_SL g334 ( 
.A(n_276),
.B(n_190),
.Y(n_334)
);

INVx2_ASAP7_75t_L g335 ( 
.A(n_255),
.Y(n_335)
);

INVx2_ASAP7_75t_L g336 ( 
.A(n_255),
.Y(n_336)
);

INVx2_ASAP7_75t_L g337 ( 
.A(n_255),
.Y(n_337)
);

AND2x2_ASAP7_75t_L g338 ( 
.A(n_264),
.B(n_193),
.Y(n_338)
);

INVx2_ASAP7_75t_SL g339 ( 
.A(n_265),
.Y(n_339)
);

NAND2xp33_ASAP7_75t_SL g340 ( 
.A(n_252),
.B(n_194),
.Y(n_340)
);

INVx2_ASAP7_75t_L g341 ( 
.A(n_261),
.Y(n_341)
);

INVx2_ASAP7_75t_SL g342 ( 
.A(n_265),
.Y(n_342)
);

INVx2_ASAP7_75t_L g343 ( 
.A(n_261),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_297),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_262),
.B(n_236),
.Y(n_345)
);

AOI21x1_ASAP7_75t_L g346 ( 
.A1(n_275),
.A2(n_198),
.B(n_195),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_297),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_275),
.Y(n_348)
);

INVx2_ASAP7_75t_L g349 ( 
.A(n_261),
.Y(n_349)
);

INVx2_ASAP7_75t_L g350 ( 
.A(n_261),
.Y(n_350)
);

INVx2_ASAP7_75t_L g351 ( 
.A(n_261),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_268),
.B(n_205),
.Y(n_352)
);

INVx2_ASAP7_75t_L g353 ( 
.A(n_267),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_274),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_SL g355 ( 
.A(n_311),
.B(n_252),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_354),
.Y(n_356)
);

NAND2xp33_ASAP7_75t_L g357 ( 
.A(n_327),
.B(n_292),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_308),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_325),
.B(n_268),
.Y(n_359)
);

BUFx3_ASAP7_75t_L g360 ( 
.A(n_333),
.Y(n_360)
);

AND2x4_ASAP7_75t_L g361 ( 
.A(n_328),
.B(n_254),
.Y(n_361)
);

NAND2xp33_ASAP7_75t_L g362 ( 
.A(n_327),
.B(n_345),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_SL g363 ( 
.A(n_315),
.B(n_299),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_325),
.B(n_268),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_L g365 ( 
.A(n_314),
.B(n_263),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_325),
.B(n_266),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_308),
.Y(n_367)
);

OR2x2_ASAP7_75t_L g368 ( 
.A(n_332),
.B(n_282),
.Y(n_368)
);

NAND3xp33_ASAP7_75t_L g369 ( 
.A(n_334),
.B(n_291),
.C(n_285),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_313),
.Y(n_370)
);

NOR2xp33_ASAP7_75t_L g371 ( 
.A(n_314),
.B(n_293),
.Y(n_371)
);

AO221x1_ASAP7_75t_L g372 ( 
.A1(n_307),
.A2(n_302),
.B1(n_285),
.B2(n_291),
.C(n_296),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_352),
.B(n_266),
.Y(n_373)
);

AND2x2_ASAP7_75t_L g374 ( 
.A(n_329),
.B(n_287),
.Y(n_374)
);

INVx2_ASAP7_75t_L g375 ( 
.A(n_313),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_334),
.B(n_266),
.Y(n_376)
);

INVx8_ASAP7_75t_L g377 ( 
.A(n_321),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_324),
.B(n_288),
.Y(n_378)
);

INVxp67_ASAP7_75t_L g379 ( 
.A(n_339),
.Y(n_379)
);

BUFx6f_ASAP7_75t_SL g380 ( 
.A(n_316),
.Y(n_380)
);

INVxp67_ASAP7_75t_L g381 ( 
.A(n_342),
.Y(n_381)
);

NOR2xp33_ASAP7_75t_L g382 ( 
.A(n_305),
.B(n_295),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_318),
.B(n_302),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_318),
.B(n_302),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_319),
.Y(n_385)
);

NOR2xp33_ASAP7_75t_L g386 ( 
.A(n_305),
.B(n_279),
.Y(n_386)
);

AND2x6_ASAP7_75t_L g387 ( 
.A(n_338),
.B(n_260),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_320),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_320),
.B(n_279),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_322),
.B(n_279),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_322),
.B(n_279),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_348),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_331),
.B(n_294),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_331),
.B(n_294),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_335),
.B(n_336),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_317),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_330),
.Y(n_397)
);

INVx3_ASAP7_75t_L g398 ( 
.A(n_335),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g399 ( 
.A(n_336),
.B(n_294),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_SL g400 ( 
.A(n_306),
.B(n_206),
.Y(n_400)
);

NAND2xp33_ASAP7_75t_L g401 ( 
.A(n_340),
.B(n_272),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_337),
.B(n_294),
.Y(n_402)
);

NOR2xp33_ASAP7_75t_SL g403 ( 
.A(n_304),
.B(n_272),
.Y(n_403)
);

NOR2xp33_ASAP7_75t_L g404 ( 
.A(n_309),
.B(n_294),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_341),
.B(n_296),
.Y(n_405)
);

NOR2xp33_ASAP7_75t_L g406 ( 
.A(n_309),
.B(n_296),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_341),
.B(n_296),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_343),
.B(n_298),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_343),
.B(n_298),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_349),
.B(n_298),
.Y(n_410)
);

INVx8_ASAP7_75t_L g411 ( 
.A(n_321),
.Y(n_411)
);

NAND2xp33_ASAP7_75t_L g412 ( 
.A(n_340),
.B(n_272),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_344),
.Y(n_413)
);

INVx2_ASAP7_75t_SL g414 ( 
.A(n_306),
.Y(n_414)
);

NOR2xp67_ASAP7_75t_L g415 ( 
.A(n_312),
.B(n_207),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_349),
.B(n_298),
.Y(n_416)
);

BUFx6f_ASAP7_75t_L g417 ( 
.A(n_350),
.Y(n_417)
);

INVx2_ASAP7_75t_L g418 ( 
.A(n_350),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_351),
.B(n_298),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_347),
.Y(n_420)
);

BUFx8_ASAP7_75t_L g421 ( 
.A(n_310),
.Y(n_421)
);

INVx2_ASAP7_75t_L g422 ( 
.A(n_351),
.Y(n_422)
);

NOR2xp67_ASAP7_75t_L g423 ( 
.A(n_312),
.B(n_209),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_365),
.B(n_360),
.Y(n_424)
);

AO21x1_ASAP7_75t_L g425 ( 
.A1(n_357),
.A2(n_301),
.B(n_346),
.Y(n_425)
);

HB1xp67_ASAP7_75t_SL g426 ( 
.A(n_421),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_356),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_386),
.B(n_306),
.Y(n_428)
);

OAI21xp33_ASAP7_75t_L g429 ( 
.A1(n_371),
.A2(n_304),
.B(n_253),
.Y(n_429)
);

A2O1A1Ixp33_ASAP7_75t_L g430 ( 
.A1(n_382),
.A2(n_301),
.B(n_353),
.C(n_267),
.Y(n_430)
);

AOI21xp5_ASAP7_75t_L g431 ( 
.A1(n_362),
.A2(n_364),
.B(n_359),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_404),
.B(n_307),
.Y(n_432)
);

AOI21xp5_ASAP7_75t_L g433 ( 
.A1(n_366),
.A2(n_326),
.B(n_401),
.Y(n_433)
);

NOR2xp33_ASAP7_75t_L g434 ( 
.A(n_379),
.B(n_381),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_406),
.B(n_353),
.Y(n_435)
);

HB1xp67_ASAP7_75t_L g436 ( 
.A(n_374),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_SL g437 ( 
.A(n_355),
.B(n_312),
.Y(n_437)
);

NOR2xp33_ASAP7_75t_L g438 ( 
.A(n_363),
.B(n_271),
.Y(n_438)
);

INVx2_ASAP7_75t_L g439 ( 
.A(n_392),
.Y(n_439)
);

AOI21xp33_ASAP7_75t_L g440 ( 
.A1(n_369),
.A2(n_316),
.B(n_321),
.Y(n_440)
);

NOR2xp33_ASAP7_75t_L g441 ( 
.A(n_400),
.B(n_271),
.Y(n_441)
);

AO21x1_ASAP7_75t_L g442 ( 
.A1(n_412),
.A2(n_277),
.B(n_273),
.Y(n_442)
);

AOI21xp5_ASAP7_75t_L g443 ( 
.A1(n_373),
.A2(n_326),
.B(n_312),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_396),
.Y(n_444)
);

OAI21xp5_ASAP7_75t_L g445 ( 
.A1(n_369),
.A2(n_378),
.B(n_376),
.Y(n_445)
);

INVx3_ASAP7_75t_L g446 ( 
.A(n_417),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_387),
.B(n_397),
.Y(n_447)
);

AOI21xp5_ASAP7_75t_L g448 ( 
.A1(n_395),
.A2(n_326),
.B(n_303),
.Y(n_448)
);

NOR2xp33_ASAP7_75t_L g449 ( 
.A(n_414),
.B(n_316),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_387),
.B(n_303),
.Y(n_450)
);

AO21x1_ASAP7_75t_L g451 ( 
.A1(n_403),
.A2(n_277),
.B(n_273),
.Y(n_451)
);

AND2x4_ASAP7_75t_L g452 ( 
.A(n_361),
.B(n_256),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_387),
.B(n_285),
.Y(n_453)
);

AO21x1_ASAP7_75t_L g454 ( 
.A1(n_372),
.A2(n_285),
.B(n_253),
.Y(n_454)
);

OR2x2_ASAP7_75t_L g455 ( 
.A(n_368),
.B(n_316),
.Y(n_455)
);

OAI21xp5_ASAP7_75t_L g456 ( 
.A1(n_383),
.A2(n_259),
.B(n_258),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_L g457 ( 
.A(n_413),
.B(n_420),
.Y(n_457)
);

AOI21xp5_ASAP7_75t_L g458 ( 
.A1(n_389),
.A2(n_259),
.B(n_258),
.Y(n_458)
);

AND2x4_ASAP7_75t_L g459 ( 
.A(n_361),
.B(n_256),
.Y(n_459)
);

AOI21xp5_ASAP7_75t_L g460 ( 
.A1(n_390),
.A2(n_259),
.B(n_258),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g461 ( 
.A(n_417),
.B(n_259),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_384),
.Y(n_462)
);

INVx2_ASAP7_75t_L g463 ( 
.A(n_375),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_L g464 ( 
.A(n_417),
.B(n_269),
.Y(n_464)
);

O2A1O1Ixp5_ASAP7_75t_L g465 ( 
.A1(n_418),
.A2(n_257),
.B(n_269),
.C(n_272),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_358),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_L g467 ( 
.A(n_398),
.B(n_269),
.Y(n_467)
);

O2A1O1Ixp33_ASAP7_75t_L g468 ( 
.A1(n_391),
.A2(n_257),
.B(n_269),
.C(n_321),
.Y(n_468)
);

INVx2_ASAP7_75t_L g469 ( 
.A(n_422),
.Y(n_469)
);

NAND2xp33_ASAP7_75t_L g470 ( 
.A(n_367),
.B(n_272),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_370),
.Y(n_471)
);

INVx3_ASAP7_75t_L g472 ( 
.A(n_385),
.Y(n_472)
);

AOI21xp5_ASAP7_75t_L g473 ( 
.A1(n_393),
.A2(n_399),
.B(n_394),
.Y(n_473)
);

BUFx2_ASAP7_75t_L g474 ( 
.A(n_421),
.Y(n_474)
);

AOI21xp5_ASAP7_75t_L g475 ( 
.A1(n_402),
.A2(n_215),
.B(n_213),
.Y(n_475)
);

INVx3_ASAP7_75t_L g476 ( 
.A(n_388),
.Y(n_476)
);

AOI21xp5_ASAP7_75t_L g477 ( 
.A1(n_405),
.A2(n_216),
.B(n_218),
.Y(n_477)
);

OAI21xp5_ASAP7_75t_L g478 ( 
.A1(n_415),
.A2(n_228),
.B(n_226),
.Y(n_478)
);

CKINVDCx20_ASAP7_75t_R g479 ( 
.A(n_377),
.Y(n_479)
);

AND2x2_ASAP7_75t_SL g480 ( 
.A(n_380),
.B(n_310),
.Y(n_480)
);

CKINVDCx8_ASAP7_75t_R g481 ( 
.A(n_377),
.Y(n_481)
);

OAI21xp5_ASAP7_75t_L g482 ( 
.A1(n_423),
.A2(n_231),
.B(n_229),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_407),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_L g484 ( 
.A(n_408),
.B(n_221),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_L g485 ( 
.A(n_409),
.B(n_227),
.Y(n_485)
);

AND2x4_ASAP7_75t_L g486 ( 
.A(n_410),
.B(n_27),
.Y(n_486)
);

OAI21xp33_ASAP7_75t_L g487 ( 
.A1(n_416),
.A2(n_323),
.B(n_9),
.Y(n_487)
);

AOI21xp5_ASAP7_75t_L g488 ( 
.A1(n_419),
.A2(n_411),
.B(n_377),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_411),
.Y(n_489)
);

OAI21xp33_ASAP7_75t_L g490 ( 
.A1(n_411),
.A2(n_8),
.B(n_10),
.Y(n_490)
);

AOI21x1_ASAP7_75t_L g491 ( 
.A1(n_380),
.A2(n_90),
.B(n_180),
.Y(n_491)
);

OAI22xp5_ASAP7_75t_L g492 ( 
.A1(n_365),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_492)
);

HB1xp67_ASAP7_75t_L g493 ( 
.A(n_379),
.Y(n_493)
);

OAI22xp5_ASAP7_75t_L g494 ( 
.A1(n_424),
.A2(n_12),
.B1(n_13),
.B2(n_15),
.Y(n_494)
);

OAI21x1_ASAP7_75t_L g495 ( 
.A1(n_473),
.A2(n_93),
.B(n_179),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_L g496 ( 
.A(n_428),
.B(n_16),
.Y(n_496)
);

INVx2_ASAP7_75t_L g497 ( 
.A(n_444),
.Y(n_497)
);

AOI21xp5_ASAP7_75t_L g498 ( 
.A1(n_461),
.A2(n_92),
.B(n_174),
.Y(n_498)
);

OAI21xp5_ASAP7_75t_L g499 ( 
.A1(n_432),
.A2(n_465),
.B(n_460),
.Y(n_499)
);

INVx2_ASAP7_75t_L g500 ( 
.A(n_472),
.Y(n_500)
);

AND2x2_ASAP7_75t_L g501 ( 
.A(n_436),
.B(n_17),
.Y(n_501)
);

AOI21xp5_ASAP7_75t_L g502 ( 
.A1(n_464),
.A2(n_89),
.B(n_172),
.Y(n_502)
);

AOI21x1_ASAP7_75t_L g503 ( 
.A1(n_448),
.A2(n_88),
.B(n_171),
.Y(n_503)
);

OAI21x1_ASAP7_75t_L g504 ( 
.A1(n_458),
.A2(n_181),
.B(n_86),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_427),
.Y(n_505)
);

INVxp67_ASAP7_75t_L g506 ( 
.A(n_434),
.Y(n_506)
);

OAI21x1_ASAP7_75t_L g507 ( 
.A1(n_433),
.A2(n_169),
.B(n_85),
.Y(n_507)
);

HB1xp67_ASAP7_75t_L g508 ( 
.A(n_493),
.Y(n_508)
);

INVxp67_ASAP7_75t_L g509 ( 
.A(n_438),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_466),
.Y(n_510)
);

OAI21x1_ASAP7_75t_L g511 ( 
.A1(n_456),
.A2(n_166),
.B(n_84),
.Y(n_511)
);

A2O1A1Ixp33_ASAP7_75t_L g512 ( 
.A1(n_445),
.A2(n_17),
.B(n_18),
.C(n_19),
.Y(n_512)
);

A2O1A1Ixp33_ASAP7_75t_L g513 ( 
.A1(n_445),
.A2(n_18),
.B(n_19),
.C(n_20),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_L g514 ( 
.A(n_462),
.B(n_21),
.Y(n_514)
);

OR2x2_ASAP7_75t_L g515 ( 
.A(n_455),
.B(n_21),
.Y(n_515)
);

BUFx2_ASAP7_75t_L g516 ( 
.A(n_452),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_471),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_L g518 ( 
.A(n_483),
.B(n_22),
.Y(n_518)
);

BUFx4_ASAP7_75t_SL g519 ( 
.A(n_479),
.Y(n_519)
);

NAND2xp33_ASAP7_75t_L g520 ( 
.A(n_450),
.B(n_28),
.Y(n_520)
);

AOI21xp5_ASAP7_75t_L g521 ( 
.A1(n_431),
.A2(n_97),
.B(n_29),
.Y(n_521)
);

AOI21xp5_ASAP7_75t_L g522 ( 
.A1(n_467),
.A2(n_98),
.B(n_33),
.Y(n_522)
);

AOI21x1_ASAP7_75t_L g523 ( 
.A1(n_435),
.A2(n_99),
.B(n_34),
.Y(n_523)
);

AOI21xp33_ASAP7_75t_L g524 ( 
.A1(n_441),
.A2(n_22),
.B(n_35),
.Y(n_524)
);

OR2x6_ASAP7_75t_L g525 ( 
.A(n_474),
.B(n_36),
.Y(n_525)
);

OAI21xp5_ASAP7_75t_L g526 ( 
.A1(n_456),
.A2(n_38),
.B(n_39),
.Y(n_526)
);

INVx4_ASAP7_75t_L g527 ( 
.A(n_446),
.Y(n_527)
);

BUFx2_ASAP7_75t_L g528 ( 
.A(n_452),
.Y(n_528)
);

NAND3xp33_ASAP7_75t_L g529 ( 
.A(n_447),
.B(n_40),
.C(n_41),
.Y(n_529)
);

AOI21xp33_ASAP7_75t_L g530 ( 
.A1(n_453),
.A2(n_42),
.B(n_43),
.Y(n_530)
);

OAI22x1_ASAP7_75t_L g531 ( 
.A1(n_449),
.A2(n_44),
.B1(n_45),
.B2(n_47),
.Y(n_531)
);

NOR2xp33_ASAP7_75t_SL g532 ( 
.A(n_481),
.B(n_50),
.Y(n_532)
);

OAI21x1_ASAP7_75t_L g533 ( 
.A1(n_472),
.A2(n_51),
.B(n_52),
.Y(n_533)
);

CKINVDCx5p33_ASAP7_75t_R g534 ( 
.A(n_426),
.Y(n_534)
);

OAI21x1_ASAP7_75t_L g535 ( 
.A1(n_476),
.A2(n_56),
.B(n_59),
.Y(n_535)
);

AND2x2_ASAP7_75t_L g536 ( 
.A(n_429),
.B(n_65),
.Y(n_536)
);

OAI21x1_ASAP7_75t_L g537 ( 
.A1(n_476),
.A2(n_163),
.B(n_67),
.Y(n_537)
);

INVx3_ASAP7_75t_L g538 ( 
.A(n_446),
.Y(n_538)
);

OAI21xp5_ASAP7_75t_L g539 ( 
.A1(n_430),
.A2(n_66),
.B(n_68),
.Y(n_539)
);

AND3x4_ASAP7_75t_L g540 ( 
.A(n_459),
.B(n_69),
.C(n_72),
.Y(n_540)
);

AOI21xp33_ASAP7_75t_L g541 ( 
.A1(n_440),
.A2(n_75),
.B(n_77),
.Y(n_541)
);

OAI21xp5_ASAP7_75t_L g542 ( 
.A1(n_468),
.A2(n_78),
.B(n_79),
.Y(n_542)
);

OAI21x1_ASAP7_75t_L g543 ( 
.A1(n_488),
.A2(n_162),
.B(n_81),
.Y(n_543)
);

INVxp67_ASAP7_75t_L g544 ( 
.A(n_459),
.Y(n_544)
);

OAI21x1_ASAP7_75t_L g545 ( 
.A1(n_425),
.A2(n_160),
.B(n_82),
.Y(n_545)
);

A2O1A1Ixp33_ASAP7_75t_L g546 ( 
.A1(n_487),
.A2(n_80),
.B(n_83),
.C(n_94),
.Y(n_546)
);

OAI21xp33_ASAP7_75t_L g547 ( 
.A1(n_490),
.A2(n_95),
.B(n_101),
.Y(n_547)
);

INVx2_ASAP7_75t_L g548 ( 
.A(n_439),
.Y(n_548)
);

OR2x2_ASAP7_75t_L g549 ( 
.A(n_457),
.B(n_103),
.Y(n_549)
);

O2A1O1Ixp5_ASAP7_75t_L g550 ( 
.A1(n_442),
.A2(n_104),
.B(n_106),
.C(n_107),
.Y(n_550)
);

OA21x2_ASAP7_75t_L g551 ( 
.A1(n_499),
.A2(n_454),
.B(n_451),
.Y(n_551)
);

AOI22xp5_ASAP7_75t_L g552 ( 
.A1(n_547),
.A2(n_492),
.B1(n_437),
.B2(n_486),
.Y(n_552)
);

AND2x4_ASAP7_75t_L g553 ( 
.A(n_544),
.B(n_489),
.Y(n_553)
);

INVx5_ASAP7_75t_L g554 ( 
.A(n_527),
.Y(n_554)
);

OAI21x1_ASAP7_75t_SL g555 ( 
.A1(n_526),
.A2(n_491),
.B(n_492),
.Y(n_555)
);

BUFx6f_ASAP7_75t_L g556 ( 
.A(n_516),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_505),
.Y(n_557)
);

BUFx12f_ASAP7_75t_L g558 ( 
.A(n_534),
.Y(n_558)
);

OAI21x1_ASAP7_75t_L g559 ( 
.A1(n_504),
.A2(n_463),
.B(n_469),
.Y(n_559)
);

OAI21x1_ASAP7_75t_L g560 ( 
.A1(n_507),
.A2(n_485),
.B(n_484),
.Y(n_560)
);

OAI21x1_ASAP7_75t_L g561 ( 
.A1(n_495),
.A2(n_443),
.B(n_482),
.Y(n_561)
);

INVx2_ASAP7_75t_SL g562 ( 
.A(n_508),
.Y(n_562)
);

NOR2xp33_ASAP7_75t_L g563 ( 
.A(n_509),
.B(n_480),
.Y(n_563)
);

OAI21x1_ASAP7_75t_L g564 ( 
.A1(n_499),
.A2(n_478),
.B(n_477),
.Y(n_564)
);

BUFx4f_ASAP7_75t_L g565 ( 
.A(n_540),
.Y(n_565)
);

AO21x2_ASAP7_75t_L g566 ( 
.A1(n_542),
.A2(n_470),
.B(n_486),
.Y(n_566)
);

OAI21x1_ASAP7_75t_L g567 ( 
.A1(n_511),
.A2(n_475),
.B(n_114),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_L g568 ( 
.A(n_506),
.B(n_500),
.Y(n_568)
);

AO21x2_ASAP7_75t_L g569 ( 
.A1(n_542),
.A2(n_112),
.B(n_115),
.Y(n_569)
);

AOI22xp33_ASAP7_75t_L g570 ( 
.A1(n_524),
.A2(n_116),
.B1(n_119),
.B2(n_120),
.Y(n_570)
);

OA21x2_ASAP7_75t_L g571 ( 
.A1(n_539),
.A2(n_122),
.B(n_123),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_510),
.Y(n_572)
);

OAI21x1_ASAP7_75t_L g573 ( 
.A1(n_543),
.A2(n_127),
.B(n_128),
.Y(n_573)
);

AO21x2_ASAP7_75t_L g574 ( 
.A1(n_539),
.A2(n_129),
.B(n_133),
.Y(n_574)
);

OAI21x1_ASAP7_75t_L g575 ( 
.A1(n_503),
.A2(n_134),
.B(n_136),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_L g576 ( 
.A(n_496),
.B(n_137),
.Y(n_576)
);

INVx3_ASAP7_75t_L g577 ( 
.A(n_527),
.Y(n_577)
);

OAI21x1_ASAP7_75t_L g578 ( 
.A1(n_533),
.A2(n_138),
.B(n_139),
.Y(n_578)
);

NOR2xp33_ASAP7_75t_L g579 ( 
.A(n_514),
.B(n_158),
.Y(n_579)
);

OAI21xp5_ASAP7_75t_L g580 ( 
.A1(n_526),
.A2(n_140),
.B(n_141),
.Y(n_580)
);

OAI21x1_ASAP7_75t_L g581 ( 
.A1(n_535),
.A2(n_142),
.B(n_143),
.Y(n_581)
);

OR2x2_ASAP7_75t_L g582 ( 
.A(n_528),
.B(n_144),
.Y(n_582)
);

OAI21xp5_ASAP7_75t_L g583 ( 
.A1(n_518),
.A2(n_155),
.B(n_146),
.Y(n_583)
);

OA21x2_ASAP7_75t_L g584 ( 
.A1(n_545),
.A2(n_145),
.B(n_147),
.Y(n_584)
);

AOI21x1_ASAP7_75t_L g585 ( 
.A1(n_521),
.A2(n_148),
.B(n_151),
.Y(n_585)
);

OAI21x1_ASAP7_75t_L g586 ( 
.A1(n_537),
.A2(n_152),
.B(n_538),
.Y(n_586)
);

INVx3_ASAP7_75t_L g587 ( 
.A(n_538),
.Y(n_587)
);

OA21x2_ASAP7_75t_L g588 ( 
.A1(n_530),
.A2(n_550),
.B(n_541),
.Y(n_588)
);

INVx1_ASAP7_75t_SL g589 ( 
.A(n_515),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_L g590 ( 
.A(n_497),
.B(n_536),
.Y(n_590)
);

INVx1_ASAP7_75t_SL g591 ( 
.A(n_501),
.Y(n_591)
);

INVx5_ASAP7_75t_L g592 ( 
.A(n_525),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_L g593 ( 
.A(n_517),
.B(n_549),
.Y(n_593)
);

INVx6_ASAP7_75t_L g594 ( 
.A(n_525),
.Y(n_594)
);

OAI21x1_ASAP7_75t_L g595 ( 
.A1(n_522),
.A2(n_498),
.B(n_502),
.Y(n_595)
);

INVx2_ASAP7_75t_L g596 ( 
.A(n_548),
.Y(n_596)
);

OAI21x1_ASAP7_75t_L g597 ( 
.A1(n_523),
.A2(n_529),
.B(n_494),
.Y(n_597)
);

AOI21x1_ASAP7_75t_L g598 ( 
.A1(n_531),
.A2(n_529),
.B(n_494),
.Y(n_598)
);

BUFx6f_ASAP7_75t_L g599 ( 
.A(n_525),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_557),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_572),
.Y(n_601)
);

INVx2_ASAP7_75t_L g602 ( 
.A(n_587),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_596),
.Y(n_603)
);

OAI22xp5_ASAP7_75t_L g604 ( 
.A1(n_590),
.A2(n_546),
.B1(n_513),
.B2(n_512),
.Y(n_604)
);

BUFx3_ASAP7_75t_L g605 ( 
.A(n_556),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_587),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_593),
.Y(n_607)
);

AND2x4_ASAP7_75t_L g608 ( 
.A(n_592),
.B(n_519),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_593),
.Y(n_609)
);

INVx4_ASAP7_75t_L g610 ( 
.A(n_554),
.Y(n_610)
);

INVx2_ASAP7_75t_L g611 ( 
.A(n_551),
.Y(n_611)
);

HB1xp67_ASAP7_75t_L g612 ( 
.A(n_562),
.Y(n_612)
);

INVx2_ASAP7_75t_L g613 ( 
.A(n_551),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_590),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_568),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_568),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_577),
.Y(n_617)
);

NAND2x1p5_ASAP7_75t_L g618 ( 
.A(n_554),
.B(n_520),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_577),
.Y(n_619)
);

OAI21x1_ASAP7_75t_L g620 ( 
.A1(n_586),
.A2(n_530),
.B(n_532),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_552),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_552),
.Y(n_622)
);

BUFx2_ASAP7_75t_L g623 ( 
.A(n_556),
.Y(n_623)
);

AND2x2_ASAP7_75t_L g624 ( 
.A(n_565),
.B(n_532),
.Y(n_624)
);

INVx2_ASAP7_75t_L g625 ( 
.A(n_559),
.Y(n_625)
);

OAI21x1_ASAP7_75t_L g626 ( 
.A1(n_567),
.A2(n_578),
.B(n_581),
.Y(n_626)
);

OR2x2_ASAP7_75t_L g627 ( 
.A(n_589),
.B(n_591),
.Y(n_627)
);

INVx2_ASAP7_75t_L g628 ( 
.A(n_554),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_554),
.Y(n_629)
);

HB1xp67_ASAP7_75t_L g630 ( 
.A(n_556),
.Y(n_630)
);

INVx2_ASAP7_75t_L g631 ( 
.A(n_597),
.Y(n_631)
);

OAI22xp5_ASAP7_75t_L g632 ( 
.A1(n_591),
.A2(n_565),
.B1(n_563),
.B2(n_592),
.Y(n_632)
);

INVx4_ASAP7_75t_L g633 ( 
.A(n_592),
.Y(n_633)
);

HB1xp67_ASAP7_75t_L g634 ( 
.A(n_589),
.Y(n_634)
);

AND2x2_ASAP7_75t_L g635 ( 
.A(n_579),
.B(n_580),
.Y(n_635)
);

INVx2_ASAP7_75t_L g636 ( 
.A(n_573),
.Y(n_636)
);

INVx2_ASAP7_75t_L g637 ( 
.A(n_585),
.Y(n_637)
);

AND2x2_ASAP7_75t_L g638 ( 
.A(n_579),
.B(n_580),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_553),
.Y(n_639)
);

BUFx2_ASAP7_75t_L g640 ( 
.A(n_553),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_598),
.Y(n_641)
);

INVx2_ASAP7_75t_L g642 ( 
.A(n_575),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_571),
.Y(n_643)
);

HB1xp67_ASAP7_75t_L g644 ( 
.A(n_582),
.Y(n_644)
);

AOI22xp33_ASAP7_75t_L g645 ( 
.A1(n_555),
.A2(n_563),
.B1(n_574),
.B2(n_592),
.Y(n_645)
);

INVx2_ASAP7_75t_SL g646 ( 
.A(n_605),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_L g647 ( 
.A(n_607),
.B(n_599),
.Y(n_647)
);

OR2x2_ASAP7_75t_L g648 ( 
.A(n_621),
.B(n_576),
.Y(n_648)
);

INVx2_ASAP7_75t_L g649 ( 
.A(n_600),
.Y(n_649)
);

BUFx6f_ASAP7_75t_L g650 ( 
.A(n_610),
.Y(n_650)
);

INVx2_ASAP7_75t_L g651 ( 
.A(n_600),
.Y(n_651)
);

INVx2_ASAP7_75t_L g652 ( 
.A(n_601),
.Y(n_652)
);

INVxp67_ASAP7_75t_SL g653 ( 
.A(n_634),
.Y(n_653)
);

INVx4_ASAP7_75t_L g654 ( 
.A(n_610),
.Y(n_654)
);

HB1xp67_ASAP7_75t_L g655 ( 
.A(n_627),
.Y(n_655)
);

AND2x2_ASAP7_75t_L g656 ( 
.A(n_614),
.B(n_583),
.Y(n_656)
);

INVx2_ASAP7_75t_L g657 ( 
.A(n_601),
.Y(n_657)
);

INVxp67_ASAP7_75t_SL g658 ( 
.A(n_627),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_L g659 ( 
.A(n_607),
.B(n_599),
.Y(n_659)
);

HB1xp67_ASAP7_75t_L g660 ( 
.A(n_612),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_603),
.Y(n_661)
);

INVx2_ASAP7_75t_L g662 ( 
.A(n_611),
.Y(n_662)
);

AND2x4_ASAP7_75t_L g663 ( 
.A(n_633),
.B(n_599),
.Y(n_663)
);

HB1xp67_ASAP7_75t_L g664 ( 
.A(n_640),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_611),
.Y(n_665)
);

AND2x4_ASAP7_75t_L g666 ( 
.A(n_633),
.B(n_583),
.Y(n_666)
);

HB1xp67_ASAP7_75t_L g667 ( 
.A(n_640),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_613),
.Y(n_668)
);

AND2x2_ASAP7_75t_L g669 ( 
.A(n_614),
.B(n_574),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_603),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_615),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_615),
.Y(n_672)
);

AND2x2_ASAP7_75t_L g673 ( 
.A(n_609),
.B(n_576),
.Y(n_673)
);

AND2x2_ASAP7_75t_L g674 ( 
.A(n_609),
.B(n_571),
.Y(n_674)
);

BUFx5_ASAP7_75t_L g675 ( 
.A(n_643),
.Y(n_675)
);

INVx3_ASAP7_75t_L g676 ( 
.A(n_610),
.Y(n_676)
);

BUFx2_ASAP7_75t_L g677 ( 
.A(n_641),
.Y(n_677)
);

AND2x2_ASAP7_75t_L g678 ( 
.A(n_616),
.B(n_570),
.Y(n_678)
);

AND2x4_ASAP7_75t_L g679 ( 
.A(n_633),
.B(n_569),
.Y(n_679)
);

AND2x2_ASAP7_75t_L g680 ( 
.A(n_616),
.B(n_570),
.Y(n_680)
);

AND2x2_ASAP7_75t_L g681 ( 
.A(n_621),
.B(n_569),
.Y(n_681)
);

INVx2_ASAP7_75t_SL g682 ( 
.A(n_605),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_639),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_641),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_606),
.Y(n_685)
);

AOI22xp5_ASAP7_75t_L g686 ( 
.A1(n_635),
.A2(n_594),
.B1(n_558),
.B2(n_566),
.Y(n_686)
);

AND2x2_ASAP7_75t_L g687 ( 
.A(n_622),
.B(n_584),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_L g688 ( 
.A(n_644),
.B(n_594),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_L g689 ( 
.A(n_622),
.B(n_638),
.Y(n_689)
);

AND2x2_ASAP7_75t_L g690 ( 
.A(n_635),
.B(n_584),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_631),
.Y(n_691)
);

AND2x2_ASAP7_75t_L g692 ( 
.A(n_638),
.B(n_566),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_606),
.Y(n_693)
);

AND2x2_ASAP7_75t_L g694 ( 
.A(n_602),
.B(n_564),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_631),
.Y(n_695)
);

INVx2_ASAP7_75t_SL g696 ( 
.A(n_623),
.Y(n_696)
);

NOR2xp33_ASAP7_75t_L g697 ( 
.A(n_624),
.B(n_588),
.Y(n_697)
);

OAI22xp5_ASAP7_75t_L g698 ( 
.A1(n_645),
.A2(n_595),
.B1(n_561),
.B2(n_560),
.Y(n_698)
);

AND2x4_ASAP7_75t_L g699 ( 
.A(n_649),
.B(n_628),
.Y(n_699)
);

INVx2_ASAP7_75t_L g700 ( 
.A(n_675),
.Y(n_700)
);

AND2x2_ASAP7_75t_L g701 ( 
.A(n_692),
.B(n_602),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_649),
.Y(n_702)
);

NOR2x1_ASAP7_75t_SL g703 ( 
.A(n_671),
.B(n_637),
.Y(n_703)
);

OR2x2_ASAP7_75t_L g704 ( 
.A(n_692),
.B(n_632),
.Y(n_704)
);

AOI22xp33_ASAP7_75t_L g705 ( 
.A1(n_697),
.A2(n_624),
.B1(n_608),
.B2(n_604),
.Y(n_705)
);

AND2x2_ASAP7_75t_L g706 ( 
.A(n_681),
.B(n_623),
.Y(n_706)
);

AOI22xp33_ASAP7_75t_L g707 ( 
.A1(n_666),
.A2(n_608),
.B1(n_630),
.B2(n_619),
.Y(n_707)
);

AOI22xp33_ASAP7_75t_L g708 ( 
.A1(n_666),
.A2(n_608),
.B1(n_617),
.B2(n_619),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_651),
.Y(n_709)
);

AND2x2_ASAP7_75t_L g710 ( 
.A(n_681),
.B(n_689),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_651),
.Y(n_711)
);

OR2x2_ASAP7_75t_L g712 ( 
.A(n_658),
.B(n_677),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_L g713 ( 
.A(n_655),
.B(n_617),
.Y(n_713)
);

AOI22xp33_ASAP7_75t_L g714 ( 
.A1(n_666),
.A2(n_618),
.B1(n_637),
.B2(n_629),
.Y(n_714)
);

AND2x4_ASAP7_75t_L g715 ( 
.A(n_652),
.B(n_657),
.Y(n_715)
);

OAI22xp5_ASAP7_75t_SL g716 ( 
.A1(n_688),
.A2(n_629),
.B1(n_618),
.B2(n_628),
.Y(n_716)
);

OR2x2_ASAP7_75t_L g717 ( 
.A(n_677),
.B(n_625),
.Y(n_717)
);

BUFx2_ASAP7_75t_L g718 ( 
.A(n_675),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_652),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_657),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_684),
.Y(n_721)
);

OR2x2_ASAP7_75t_L g722 ( 
.A(n_648),
.B(n_625),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_684),
.Y(n_723)
);

INVx2_ASAP7_75t_SL g724 ( 
.A(n_696),
.Y(n_724)
);

AND2x2_ASAP7_75t_L g725 ( 
.A(n_669),
.B(n_620),
.Y(n_725)
);

AND2x2_ASAP7_75t_L g726 ( 
.A(n_669),
.B(n_620),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_672),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_661),
.Y(n_728)
);

BUFx3_ASAP7_75t_L g729 ( 
.A(n_663),
.Y(n_729)
);

AOI22xp5_ASAP7_75t_L g730 ( 
.A1(n_686),
.A2(n_618),
.B1(n_636),
.B2(n_642),
.Y(n_730)
);

INVx2_ASAP7_75t_L g731 ( 
.A(n_675),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_670),
.Y(n_732)
);

AND2x2_ASAP7_75t_L g733 ( 
.A(n_678),
.B(n_636),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_685),
.Y(n_734)
);

HB1xp67_ASAP7_75t_L g735 ( 
.A(n_664),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_693),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_L g737 ( 
.A(n_673),
.B(n_642),
.Y(n_737)
);

AND2x2_ASAP7_75t_L g738 ( 
.A(n_678),
.B(n_626),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_665),
.Y(n_739)
);

OR2x2_ASAP7_75t_L g740 ( 
.A(n_648),
.B(n_626),
.Y(n_740)
);

AOI22xp33_ASAP7_75t_L g741 ( 
.A1(n_680),
.A2(n_656),
.B1(n_673),
.B2(n_667),
.Y(n_741)
);

INVx2_ASAP7_75t_L g742 ( 
.A(n_675),
.Y(n_742)
);

INVx2_ASAP7_75t_L g743 ( 
.A(n_675),
.Y(n_743)
);

AND2x2_ASAP7_75t_L g744 ( 
.A(n_710),
.B(n_690),
.Y(n_744)
);

AND2x4_ASAP7_75t_L g745 ( 
.A(n_715),
.B(n_679),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_721),
.Y(n_746)
);

AND2x4_ASAP7_75t_L g747 ( 
.A(n_715),
.B(n_679),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_723),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_728),
.Y(n_749)
);

AND2x2_ASAP7_75t_L g750 ( 
.A(n_710),
.B(n_690),
.Y(n_750)
);

INVx2_ASAP7_75t_L g751 ( 
.A(n_715),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_L g752 ( 
.A(n_735),
.B(n_653),
.Y(n_752)
);

AND2x2_ASAP7_75t_L g753 ( 
.A(n_738),
.B(n_694),
.Y(n_753)
);

INVx2_ASAP7_75t_L g754 ( 
.A(n_727),
.Y(n_754)
);

INVx2_ASAP7_75t_L g755 ( 
.A(n_702),
.Y(n_755)
);

NOR2x1p5_ASAP7_75t_L g756 ( 
.A(n_729),
.B(n_647),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_L g757 ( 
.A(n_701),
.B(n_656),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_SL g758 ( 
.A(n_705),
.B(n_680),
.Y(n_758)
);

NOR2x1_ASAP7_75t_L g759 ( 
.A(n_713),
.B(n_659),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_L g760 ( 
.A(n_701),
.B(n_706),
.Y(n_760)
);

AND2x2_ASAP7_75t_L g761 ( 
.A(n_738),
.B(n_694),
.Y(n_761)
);

NAND2x1_ASAP7_75t_L g762 ( 
.A(n_718),
.B(n_679),
.Y(n_762)
);

NAND2xp33_ASAP7_75t_SL g763 ( 
.A(n_716),
.B(n_650),
.Y(n_763)
);

INVx2_ASAP7_75t_L g764 ( 
.A(n_709),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_732),
.Y(n_765)
);

AOI221xp5_ASAP7_75t_L g766 ( 
.A1(n_741),
.A2(n_660),
.B1(n_683),
.B2(n_696),
.C(n_698),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_734),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_736),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_712),
.Y(n_769)
);

AND2x2_ASAP7_75t_L g770 ( 
.A(n_706),
.B(n_675),
.Y(n_770)
);

INVx2_ASAP7_75t_L g771 ( 
.A(n_711),
.Y(n_771)
);

AND2x4_ASAP7_75t_L g772 ( 
.A(n_700),
.B(n_695),
.Y(n_772)
);

NAND3xp33_ASAP7_75t_L g773 ( 
.A(n_707),
.B(n_663),
.C(n_674),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_L g774 ( 
.A(n_733),
.B(n_674),
.Y(n_774)
);

AND2x2_ASAP7_75t_L g775 ( 
.A(n_725),
.B(n_675),
.Y(n_775)
);

AND2x2_ASAP7_75t_L g776 ( 
.A(n_725),
.B(n_675),
.Y(n_776)
);

BUFx2_ASAP7_75t_L g777 ( 
.A(n_718),
.Y(n_777)
);

AND2x2_ASAP7_75t_L g778 ( 
.A(n_726),
.B(n_733),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_754),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_754),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_749),
.Y(n_781)
);

INVx2_ASAP7_75t_L g782 ( 
.A(n_755),
.Y(n_782)
);

NOR2x1p5_ASAP7_75t_SL g783 ( 
.A(n_755),
.B(n_740),
.Y(n_783)
);

AND3x2_ASAP7_75t_L g784 ( 
.A(n_766),
.B(n_663),
.C(n_699),
.Y(n_784)
);

OAI222xp33_ASAP7_75t_L g785 ( 
.A1(n_758),
.A2(n_704),
.B1(n_730),
.B2(n_708),
.C1(n_712),
.C2(n_714),
.Y(n_785)
);

INVx2_ASAP7_75t_L g786 ( 
.A(n_764),
.Y(n_786)
);

OR2x2_ASAP7_75t_L g787 ( 
.A(n_778),
.B(n_726),
.Y(n_787)
);

INVx3_ASAP7_75t_L g788 ( 
.A(n_762),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_L g789 ( 
.A(n_752),
.B(n_704),
.Y(n_789)
);

AND2x2_ASAP7_75t_L g790 ( 
.A(n_778),
.B(n_700),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_765),
.Y(n_791)
);

OR2x2_ASAP7_75t_L g792 ( 
.A(n_769),
.B(n_740),
.Y(n_792)
);

AND2x2_ASAP7_75t_L g793 ( 
.A(n_775),
.B(n_743),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_767),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_768),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_746),
.Y(n_796)
);

NOR2x1_ASAP7_75t_L g797 ( 
.A(n_759),
.B(n_699),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_L g798 ( 
.A(n_744),
.B(n_719),
.Y(n_798)
);

AND2x2_ASAP7_75t_L g799 ( 
.A(n_775),
.B(n_743),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_L g800 ( 
.A(n_744),
.B(n_750),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_L g801 ( 
.A(n_750),
.B(n_720),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_748),
.Y(n_802)
);

NAND4xp25_ASAP7_75t_L g803 ( 
.A(n_789),
.B(n_773),
.C(n_763),
.D(n_758),
.Y(n_803)
);

AOI22xp33_ASAP7_75t_SL g804 ( 
.A1(n_785),
.A2(n_784),
.B1(n_763),
.B2(n_770),
.Y(n_804)
);

AND2x2_ASAP7_75t_L g805 ( 
.A(n_793),
.B(n_776),
.Y(n_805)
);

NAND2x1p5_ASAP7_75t_L g806 ( 
.A(n_797),
.B(n_762),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_779),
.Y(n_807)
);

NOR2xp33_ASAP7_75t_L g808 ( 
.A(n_800),
.B(n_760),
.Y(n_808)
);

INVx2_ASAP7_75t_L g809 ( 
.A(n_782),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_780),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_796),
.Y(n_811)
);

AND2x2_ASAP7_75t_L g812 ( 
.A(n_793),
.B(n_776),
.Y(n_812)
);

AOI33xp33_ASAP7_75t_L g813 ( 
.A1(n_784),
.A2(n_764),
.A3(n_771),
.B1(n_770),
.B2(n_724),
.B3(n_751),
.Y(n_813)
);

OAI222xp33_ASAP7_75t_L g814 ( 
.A1(n_804),
.A2(n_787),
.B1(n_801),
.B2(n_798),
.C1(n_757),
.C2(n_792),
.Y(n_814)
);

OAI22xp5_ASAP7_75t_L g815 ( 
.A1(n_804),
.A2(n_808),
.B1(n_806),
.B2(n_756),
.Y(n_815)
);

OAI211xp5_ASAP7_75t_SL g816 ( 
.A1(n_813),
.A2(n_795),
.B(n_794),
.C(n_791),
.Y(n_816)
);

OAI21xp33_ASAP7_75t_L g817 ( 
.A1(n_803),
.A2(n_783),
.B(n_781),
.Y(n_817)
);

NAND2xp33_ASAP7_75t_SL g818 ( 
.A(n_805),
.B(n_788),
.Y(n_818)
);

AOI22xp5_ASAP7_75t_L g819 ( 
.A1(n_808),
.A2(n_745),
.B1(n_747),
.B2(n_811),
.Y(n_819)
);

AOI22xp33_ASAP7_75t_L g820 ( 
.A1(n_806),
.A2(n_745),
.B1(n_747),
.B2(n_729),
.Y(n_820)
);

NAND4xp25_ASAP7_75t_L g821 ( 
.A(n_815),
.B(n_802),
.C(n_810),
.D(n_807),
.Y(n_821)
);

OAI21xp33_ASAP7_75t_L g822 ( 
.A1(n_817),
.A2(n_792),
.B(n_799),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_L g823 ( 
.A(n_819),
.B(n_812),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_816),
.Y(n_824)
);

AOI22xp33_ASAP7_75t_SL g825 ( 
.A1(n_814),
.A2(n_788),
.B1(n_745),
.B2(n_747),
.Y(n_825)
);

AOI221xp5_ASAP7_75t_L g826 ( 
.A1(n_818),
.A2(n_799),
.B1(n_809),
.B2(n_790),
.C(n_786),
.Y(n_826)
);

AOI21xp33_ASAP7_75t_SL g827 ( 
.A1(n_820),
.A2(n_788),
.B(n_646),
.Y(n_827)
);

OAI321xp33_ASAP7_75t_L g828 ( 
.A1(n_824),
.A2(n_751),
.A3(n_777),
.B1(n_771),
.B2(n_724),
.C(n_737),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_SL g829 ( 
.A(n_825),
.B(n_790),
.Y(n_829)
);

INVx2_ASAP7_75t_L g830 ( 
.A(n_823),
.Y(n_830)
);

AOI211xp5_ASAP7_75t_SL g831 ( 
.A1(n_822),
.A2(n_739),
.B(n_699),
.C(n_774),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_L g832 ( 
.A(n_830),
.B(n_821),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_L g833 ( 
.A(n_831),
.B(n_826),
.Y(n_833)
);

NOR3xp33_ASAP7_75t_L g834 ( 
.A(n_829),
.B(n_827),
.C(n_646),
.Y(n_834)
);

NOR3x1_ASAP7_75t_L g835 ( 
.A(n_832),
.B(n_828),
.C(n_682),
.Y(n_835)
);

NOR3xp33_ASAP7_75t_L g836 ( 
.A(n_833),
.B(n_682),
.C(n_654),
.Y(n_836)
);

NOR3xp33_ASAP7_75t_L g837 ( 
.A(n_834),
.B(n_654),
.C(n_676),
.Y(n_837)
);

NOR2xp33_ASAP7_75t_L g838 ( 
.A(n_832),
.B(n_786),
.Y(n_838)
);

NAND2xp33_ASAP7_75t_L g839 ( 
.A(n_836),
.B(n_782),
.Y(n_839)
);

XOR2x1_ASAP7_75t_L g840 ( 
.A(n_835),
.B(n_772),
.Y(n_840)
);

XOR2xp5_ASAP7_75t_L g841 ( 
.A(n_837),
.B(n_703),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_L g842 ( 
.A(n_838),
.B(n_761),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_L g843 ( 
.A(n_836),
.B(n_761),
.Y(n_843)
);

AND3x4_ASAP7_75t_L g844 ( 
.A(n_840),
.B(n_772),
.C(n_731),
.Y(n_844)
);

AOI21xp5_ASAP7_75t_L g845 ( 
.A1(n_839),
.A2(n_703),
.B(n_654),
.Y(n_845)
);

NOR4xp25_ASAP7_75t_L g846 ( 
.A(n_843),
.B(n_676),
.C(n_742),
.D(n_731),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_842),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_SL g848 ( 
.A(n_841),
.B(n_650),
.Y(n_848)
);

XNOR2xp5_ASAP7_75t_L g849 ( 
.A(n_847),
.B(n_753),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_844),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_L g851 ( 
.A(n_846),
.B(n_753),
.Y(n_851)
);

AOI22xp5_ASAP7_75t_L g852 ( 
.A1(n_848),
.A2(n_845),
.B1(n_777),
.B2(n_772),
.Y(n_852)
);

OAI22xp5_ASAP7_75t_L g853 ( 
.A1(n_850),
.A2(n_852),
.B1(n_851),
.B2(n_849),
.Y(n_853)
);

INVx2_ASAP7_75t_L g854 ( 
.A(n_850),
.Y(n_854)
);

INVx2_ASAP7_75t_SL g855 ( 
.A(n_850),
.Y(n_855)
);

INVx2_ASAP7_75t_L g856 ( 
.A(n_850),
.Y(n_856)
);

OAI22xp5_ASAP7_75t_L g857 ( 
.A1(n_850),
.A2(n_742),
.B1(n_722),
.B2(n_717),
.Y(n_857)
);

AOI22xp33_ASAP7_75t_L g858 ( 
.A1(n_855),
.A2(n_650),
.B1(n_676),
.B2(n_687),
.Y(n_858)
);

AOI22xp5_ASAP7_75t_L g859 ( 
.A1(n_854),
.A2(n_650),
.B1(n_687),
.B2(n_691),
.Y(n_859)
);

INVx2_ASAP7_75t_L g860 ( 
.A(n_856),
.Y(n_860)
);

INVx1_ASAP7_75t_L g861 ( 
.A(n_853),
.Y(n_861)
);

AOI21xp5_ASAP7_75t_L g862 ( 
.A1(n_861),
.A2(n_857),
.B(n_650),
.Y(n_862)
);

OAI21xp5_ASAP7_75t_L g863 ( 
.A1(n_860),
.A2(n_722),
.B(n_717),
.Y(n_863)
);

NAND2x1_ASAP7_75t_L g864 ( 
.A(n_858),
.B(n_691),
.Y(n_864)
);

OAI22xp5_ASAP7_75t_L g865 ( 
.A1(n_862),
.A2(n_859),
.B1(n_695),
.B2(n_668),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_L g866 ( 
.A(n_865),
.B(n_863),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_SL g867 ( 
.A(n_866),
.B(n_864),
.Y(n_867)
);

AOI22xp33_ASAP7_75t_L g868 ( 
.A1(n_867),
.A2(n_665),
.B1(n_668),
.B2(n_662),
.Y(n_868)
);


endmodule