module fake_netlist_5_16_n_1491 (n_137, n_294, n_318, n_82, n_194, n_316, n_248, n_124, n_86, n_136, n_146, n_315, n_268, n_61, n_127, n_75, n_235, n_226, n_74, n_57, n_111, n_155, n_43, n_116, n_22, n_284, n_46, n_245, n_21, n_139, n_38, n_105, n_280, n_4, n_17, n_254, n_33, n_23, n_302, n_265, n_293, n_244, n_47, n_173, n_198, n_247, n_314, n_8, n_321, n_292, n_100, n_212, n_119, n_275, n_252, n_26, n_295, n_133, n_330, n_2, n_6, n_39, n_147, n_67, n_307, n_87, n_150, n_106, n_209, n_259, n_301, n_68, n_93, n_186, n_134, n_191, n_51, n_63, n_171, n_153, n_204, n_250, n_260, n_298, n_320, n_286, n_122, n_282, n_331, n_10, n_24, n_325, n_132, n_90, n_101, n_281, n_240, n_189, n_220, n_291, n_231, n_257, n_31, n_13, n_152, n_317, n_9, n_323, n_195, n_42, n_227, n_45, n_271, n_94, n_123, n_167, n_234, n_308, n_267, n_297, n_156, n_5, n_225, n_219, n_157, n_131, n_192, n_223, n_158, n_138, n_264, n_109, n_163, n_276, n_95, n_183, n_185, n_243, n_169, n_59, n_255, n_215, n_196, n_211, n_218, n_181, n_3, n_290, n_221, n_178, n_287, n_72, n_104, n_41, n_56, n_141, n_15, n_145, n_48, n_50, n_313, n_88, n_216, n_168, n_164, n_311, n_208, n_142, n_214, n_328, n_140, n_299, n_303, n_296, n_241, n_184, n_65, n_78, n_144, n_114, n_96, n_165, n_213, n_129, n_98, n_197, n_107, n_69, n_236, n_1, n_249, n_304, n_329, n_203, n_274, n_80, n_35, n_73, n_277, n_92, n_19, n_149, n_309, n_30, n_14, n_84, n_130, n_322, n_258, n_29, n_79, n_151, n_25, n_306, n_288, n_188, n_190, n_201, n_263, n_44, n_224, n_40, n_34, n_228, n_283, n_112, n_85, n_239, n_55, n_49, n_310, n_54, n_12, n_76, n_170, n_27, n_77, n_102, n_161, n_273, n_270, n_230, n_81, n_118, n_279, n_70, n_253, n_261, n_174, n_289, n_172, n_206, n_217, n_312, n_210, n_91, n_176, n_182, n_143, n_83, n_237, n_180, n_207, n_37, n_229, n_108, n_66, n_177, n_60, n_16, n_0, n_58, n_18, n_117, n_326, n_233, n_205, n_113, n_246, n_179, n_125, n_269, n_128, n_285, n_120, n_232, n_327, n_135, n_126, n_202, n_266, n_272, n_193, n_251, n_53, n_160, n_154, n_62, n_148, n_71, n_300, n_159, n_175, n_262, n_238, n_99, n_319, n_20, n_121, n_242, n_36, n_200, n_162, n_64, n_222, n_28, n_89, n_115, n_324, n_199, n_187, n_32, n_103, n_97, n_166, n_11, n_7, n_256, n_305, n_52, n_278, n_110, n_1491);

input n_137;
input n_294;
input n_318;
input n_82;
input n_194;
input n_316;
input n_248;
input n_124;
input n_86;
input n_136;
input n_146;
input n_315;
input n_268;
input n_61;
input n_127;
input n_75;
input n_235;
input n_226;
input n_74;
input n_57;
input n_111;
input n_155;
input n_43;
input n_116;
input n_22;
input n_284;
input n_46;
input n_245;
input n_21;
input n_139;
input n_38;
input n_105;
input n_280;
input n_4;
input n_17;
input n_254;
input n_33;
input n_23;
input n_302;
input n_265;
input n_293;
input n_244;
input n_47;
input n_173;
input n_198;
input n_247;
input n_314;
input n_8;
input n_321;
input n_292;
input n_100;
input n_212;
input n_119;
input n_275;
input n_252;
input n_26;
input n_295;
input n_133;
input n_330;
input n_2;
input n_6;
input n_39;
input n_147;
input n_67;
input n_307;
input n_87;
input n_150;
input n_106;
input n_209;
input n_259;
input n_301;
input n_68;
input n_93;
input n_186;
input n_134;
input n_191;
input n_51;
input n_63;
input n_171;
input n_153;
input n_204;
input n_250;
input n_260;
input n_298;
input n_320;
input n_286;
input n_122;
input n_282;
input n_331;
input n_10;
input n_24;
input n_325;
input n_132;
input n_90;
input n_101;
input n_281;
input n_240;
input n_189;
input n_220;
input n_291;
input n_231;
input n_257;
input n_31;
input n_13;
input n_152;
input n_317;
input n_9;
input n_323;
input n_195;
input n_42;
input n_227;
input n_45;
input n_271;
input n_94;
input n_123;
input n_167;
input n_234;
input n_308;
input n_267;
input n_297;
input n_156;
input n_5;
input n_225;
input n_219;
input n_157;
input n_131;
input n_192;
input n_223;
input n_158;
input n_138;
input n_264;
input n_109;
input n_163;
input n_276;
input n_95;
input n_183;
input n_185;
input n_243;
input n_169;
input n_59;
input n_255;
input n_215;
input n_196;
input n_211;
input n_218;
input n_181;
input n_3;
input n_290;
input n_221;
input n_178;
input n_287;
input n_72;
input n_104;
input n_41;
input n_56;
input n_141;
input n_15;
input n_145;
input n_48;
input n_50;
input n_313;
input n_88;
input n_216;
input n_168;
input n_164;
input n_311;
input n_208;
input n_142;
input n_214;
input n_328;
input n_140;
input n_299;
input n_303;
input n_296;
input n_241;
input n_184;
input n_65;
input n_78;
input n_144;
input n_114;
input n_96;
input n_165;
input n_213;
input n_129;
input n_98;
input n_197;
input n_107;
input n_69;
input n_236;
input n_1;
input n_249;
input n_304;
input n_329;
input n_203;
input n_274;
input n_80;
input n_35;
input n_73;
input n_277;
input n_92;
input n_19;
input n_149;
input n_309;
input n_30;
input n_14;
input n_84;
input n_130;
input n_322;
input n_258;
input n_29;
input n_79;
input n_151;
input n_25;
input n_306;
input n_288;
input n_188;
input n_190;
input n_201;
input n_263;
input n_44;
input n_224;
input n_40;
input n_34;
input n_228;
input n_283;
input n_112;
input n_85;
input n_239;
input n_55;
input n_49;
input n_310;
input n_54;
input n_12;
input n_76;
input n_170;
input n_27;
input n_77;
input n_102;
input n_161;
input n_273;
input n_270;
input n_230;
input n_81;
input n_118;
input n_279;
input n_70;
input n_253;
input n_261;
input n_174;
input n_289;
input n_172;
input n_206;
input n_217;
input n_312;
input n_210;
input n_91;
input n_176;
input n_182;
input n_143;
input n_83;
input n_237;
input n_180;
input n_207;
input n_37;
input n_229;
input n_108;
input n_66;
input n_177;
input n_60;
input n_16;
input n_0;
input n_58;
input n_18;
input n_117;
input n_326;
input n_233;
input n_205;
input n_113;
input n_246;
input n_179;
input n_125;
input n_269;
input n_128;
input n_285;
input n_120;
input n_232;
input n_327;
input n_135;
input n_126;
input n_202;
input n_266;
input n_272;
input n_193;
input n_251;
input n_53;
input n_160;
input n_154;
input n_62;
input n_148;
input n_71;
input n_300;
input n_159;
input n_175;
input n_262;
input n_238;
input n_99;
input n_319;
input n_20;
input n_121;
input n_242;
input n_36;
input n_200;
input n_162;
input n_64;
input n_222;
input n_28;
input n_89;
input n_115;
input n_324;
input n_199;
input n_187;
input n_32;
input n_103;
input n_97;
input n_166;
input n_11;
input n_7;
input n_256;
input n_305;
input n_52;
input n_278;
input n_110;

output n_1491;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1166;
wire n_469;
wire n_785;
wire n_549;
wire n_532;
wire n_1161;
wire n_1150;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_880;
wire n_544;
wire n_1007;
wire n_552;
wire n_1370;
wire n_1292;
wire n_1198;
wire n_1360;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1021;
wire n_551;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1353;
wire n_800;
wire n_1347;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_915;
wire n_864;
wire n_859;
wire n_951;
wire n_1264;
wire n_447;
wire n_625;
wire n_854;
wire n_1462;
wire n_674;
wire n_417;
wire n_516;
wire n_933;
wire n_1152;
wire n_497;
wire n_606;
wire n_877;
wire n_755;
wire n_1118;
wire n_947;
wire n_1285;
wire n_373;
wire n_1359;
wire n_530;
wire n_1107;
wire n_556;
wire n_1230;
wire n_668;
wire n_375;
wire n_929;
wire n_1124;
wire n_902;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1257;
wire n_1182;
wire n_579;
wire n_1261;
wire n_938;
wire n_1098;
wire n_1154;
wire n_1242;
wire n_1135;
wire n_406;
wire n_519;
wire n_1016;
wire n_1243;
wire n_546;
wire n_1280;
wire n_731;
wire n_371;
wire n_1483;
wire n_1314;
wire n_709;
wire n_1490;
wire n_1236;
wire n_569;
wire n_920;
wire n_1289;
wire n_335;
wire n_370;
wire n_976;
wire n_343;
wire n_1449;
wire n_1078;
wire n_775;
wire n_600;
wire n_1484;
wire n_1374;
wire n_1328;
wire n_955;
wire n_339;
wire n_1146;
wire n_882;
wire n_1097;
wire n_1036;
wire n_347;
wire n_550;
wire n_696;
wire n_897;
wire n_798;
wire n_350;
wire n_646;
wire n_1428;
wire n_436;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_580;
wire n_1040;
wire n_578;
wire n_926;
wire n_344;
wire n_1218;
wire n_422;
wire n_475;
wire n_777;
wire n_1070;
wire n_1030;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_496;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_521;
wire n_663;
wire n_845;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_680;
wire n_1473;
wire n_395;
wire n_553;
wire n_901;
wire n_813;
wire n_1284;
wire n_675;
wire n_888;
wire n_1167;
wire n_637;
wire n_1384;
wire n_446;
wire n_1064;
wire n_858;
wire n_923;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_468;
wire n_342;
wire n_464;
wire n_363;
wire n_1069;
wire n_1075;
wire n_1450;
wire n_1322;
wire n_1471;
wire n_1459;
wire n_460;
wire n_889;
wire n_973;
wire n_477;
wire n_571;
wire n_461;
wire n_1211;
wire n_1197;
wire n_907;
wire n_1447;
wire n_1377;
wire n_989;
wire n_1039;
wire n_1403;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_1002;
wire n_1463;
wire n_593;
wire n_748;
wire n_586;
wire n_1058;
wire n_838;
wire n_332;
wire n_1053;
wire n_1224;
wire n_349;
wire n_1248;
wire n_1331;
wire n_953;
wire n_1014;
wire n_1241;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_440;
wire n_793;
wire n_478;
wire n_476;
wire n_534;
wire n_884;
wire n_345;
wire n_944;
wire n_647;
wire n_407;
wire n_1072;
wire n_832;
wire n_857;
wire n_561;
wire n_1319;
wire n_1387;
wire n_1027;
wire n_971;
wire n_1156;
wire n_794;
wire n_404;
wire n_686;
wire n_847;
wire n_1393;
wire n_596;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_728;
wire n_1162;
wire n_1199;
wire n_352;
wire n_1038;
wire n_520;
wire n_1369;
wire n_409;
wire n_887;
wire n_809;
wire n_870;
wire n_931;
wire n_599;
wire n_1481;
wire n_434;
wire n_868;
wire n_639;
wire n_914;
wire n_411;
wire n_414;
wire n_1293;
wire n_965;
wire n_935;
wire n_1175;
wire n_817;
wire n_360;
wire n_1479;
wire n_759;
wire n_806;
wire n_1477;
wire n_1189;
wire n_1259;
wire n_706;
wire n_746;
wire n_747;
wire n_784;
wire n_1244;
wire n_431;
wire n_1194;
wire n_615;
wire n_851;
wire n_843;
wire n_523;
wire n_913;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_776;
wire n_1415;
wire n_367;
wire n_452;
wire n_525;
wire n_1260;
wire n_1464;
wire n_649;
wire n_547;
wire n_1444;
wire n_1191;
wire n_1128;
wire n_744;
wire n_629;
wire n_590;
wire n_1308;
wire n_1233;
wire n_526;
wire n_372;
wire n_677;
wire n_1333;
wire n_1121;
wire n_433;
wire n_368;
wire n_604;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1001;
wire n_498;
wire n_1468;
wire n_689;
wire n_738;
wire n_640;
wire n_624;
wire n_1380;
wire n_1010;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_1195;
wire n_610;
wire n_936;
wire n_568;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_448;
wire n_758;
wire n_999;
wire n_1158;
wire n_563;
wire n_1145;
wire n_878;
wire n_524;
wire n_394;
wire n_1049;
wire n_1153;
wire n_741;
wire n_1306;
wire n_1068;
wire n_906;
wire n_1163;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_658;
wire n_1362;
wire n_456;
wire n_959;
wire n_535;
wire n_940;
wire n_1445;
wire n_592;
wire n_1169;
wire n_1017;
wire n_978;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1269;
wire n_1095;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_603;
wire n_1431;
wire n_484;
wire n_1033;
wire n_442;
wire n_636;
wire n_660;
wire n_1009;
wire n_1148;
wire n_742;
wire n_750;
wire n_995;
wire n_454;
wire n_374;
wire n_396;
wire n_1383;
wire n_1073;
wire n_662;
wire n_459;
wire n_962;
wire n_1215;
wire n_1171;
wire n_723;
wire n_1065;
wire n_1336;
wire n_473;
wire n_1309;
wire n_1426;
wire n_1043;
wire n_355;
wire n_486;
wire n_614;
wire n_337;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_743;
wire n_613;
wire n_1119;
wire n_1240;
wire n_829;
wire n_1416;
wire n_361;
wire n_1237;
wire n_700;
wire n_573;
wire n_1420;
wire n_1132;
wire n_388;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_761;
wire n_1006;
wire n_1270;
wire n_1486;
wire n_582;
wire n_1332;
wire n_1390;
wire n_512;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1349;
wire n_1093;
wire n_1031;
wire n_609;
wire n_1041;
wire n_1265;
wire n_383;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_630;
wire n_504;
wire n_511;
wire n_874;
wire n_358;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_1304;
wire n_1324;
wire n_987;
wire n_1455;
wire n_767;
wire n_993;
wire n_1407;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_429;
wire n_948;
wire n_1217;
wire n_628;
wire n_365;
wire n_729;
wire n_1131;
wire n_1084;
wire n_970;
wire n_911;
wire n_1430;
wire n_513;
wire n_1094;
wire n_1354;
wire n_560;
wire n_340;
wire n_1351;
wire n_1044;
wire n_1205;
wire n_346;
wire n_1209;
wire n_495;
wire n_602;
wire n_574;
wire n_1435;
wire n_879;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_490;
wire n_1327;
wire n_996;
wire n_921;
wire n_572;
wire n_366;
wire n_815;
wire n_1381;
wire n_1037;
wire n_1080;
wire n_1274;
wire n_1316;
wire n_426;
wire n_1438;
wire n_1082;
wire n_589;
wire n_716;
wire n_562;
wire n_1436;
wire n_952;
wire n_1229;
wire n_391;
wire n_701;
wire n_1437;
wire n_1023;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_531;
wire n_890;
wire n_764;
wire n_1056;
wire n_1424;
wire n_960;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_634;
wire n_1252;
wire n_348;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_1311;
wire n_950;
wire n_380;
wire n_419;
wire n_1346;
wire n_444;
wire n_1299;
wire n_1060;
wire n_1141;
wire n_389;
wire n_418;
wire n_912;
wire n_968;
wire n_451;
wire n_619;
wire n_408;
wire n_1386;
wire n_376;
wire n_967;
wire n_1442;
wire n_1139;
wire n_515;
wire n_351;
wire n_885;
wire n_397;
wire n_1432;
wire n_1357;
wire n_483;
wire n_683;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_983;
wire n_1305;
wire n_873;
wire n_378;
wire n_1112;
wire n_762;
wire n_1283;
wire n_690;
wire n_583;
wire n_1343;
wire n_1203;
wire n_821;
wire n_1179;
wire n_621;
wire n_753;
wire n_455;
wire n_1048;
wire n_1288;
wire n_385;
wire n_507;
wire n_1228;
wire n_972;
wire n_692;
wire n_820;
wire n_1200;
wire n_1301;
wire n_1363;
wire n_1185;
wire n_991;
wire n_828;
wire n_779;
wire n_576;
wire n_1143;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_537;
wire n_945;
wire n_492;
wire n_943;
wire n_341;
wire n_992;
wire n_543;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_883;
wire n_470;
wire n_449;
wire n_1214;
wire n_1342;
wire n_1400;
wire n_900;
wire n_856;
wire n_918;
wire n_942;
wire n_1147;
wire n_1077;
wire n_1422;
wire n_540;
wire n_618;
wire n_896;
wire n_356;
wire n_894;
wire n_831;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1470;
wire n_1096;
wire n_833;
wire n_1307;
wire n_988;
wire n_814;
wire n_1201;
wire n_1114;
wire n_655;
wire n_1446;
wire n_669;
wire n_472;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_387;
wire n_1149;
wire n_398;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_1219;
wire n_1204;
wire n_1035;
wire n_783;
wire n_555;
wire n_1188;
wire n_661;
wire n_849;
wire n_336;
wire n_681;
wire n_584;
wire n_430;
wire n_510;
wire n_830;
wire n_1296;
wire n_1413;
wire n_801;
wire n_875;
wire n_357;
wire n_1110;
wire n_445;
wire n_749;
wire n_1134;
wire n_1358;
wire n_717;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_1338;
wire n_577;
wire n_1419;
wire n_338;
wire n_693;
wire n_836;
wire n_990;
wire n_1389;
wire n_975;
wire n_1256;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_458;
wire n_770;
wire n_1375;
wire n_1102;
wire n_711;
wire n_1187;
wire n_1441;
wire n_1392;
wire n_1164;
wire n_489;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_876;
wire n_1190;
wire n_601;
wire n_917;
wire n_966;
wire n_1116;
wire n_1212;
wire n_726;
wire n_982;
wire n_1453;
wire n_818;
wire n_861;
wire n_1183;
wire n_899;
wire n_1253;
wire n_774;
wire n_1335;
wire n_1059;
wire n_1345;
wire n_1133;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_527;
wire n_1168;
wire n_707;
wire n_937;
wire n_1427;
wire n_393;
wire n_487;
wire n_665;
wire n_1440;
wire n_421;
wire n_1356;
wire n_910;
wire n_768;
wire n_1475;
wire n_1302;
wire n_1136;
wire n_1313;
wire n_754;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_735;
wire n_1109;
wire n_895;
wire n_1310;
wire n_427;
wire n_1399;
wire n_791;
wire n_732;
wire n_808;
wire n_797;
wire n_1025;
wire n_500;
wire n_1067;
wire n_435;
wire n_766;
wire n_1457;
wire n_541;
wire n_538;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_594;
wire n_1291;
wire n_1297;
wire n_1155;
wire n_1418;
wire n_1485;
wire n_1011;
wire n_1184;
wire n_985;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_1352;
wire n_626;
wire n_1144;
wire n_1137;
wire n_1170;
wire n_676;
wire n_653;
wire n_642;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_664;
wire n_503;
wire n_1372;
wire n_605;
wire n_1273;
wire n_353;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_1282;
wire n_1318;
wire n_780;
wire n_998;
wire n_1454;
wire n_467;
wire n_1227;
wire n_840;
wire n_1334;
wire n_501;
wire n_823;
wire n_725;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_672;
wire n_581;
wire n_382;
wire n_554;
wire n_898;
wire n_1013;
wire n_1452;
wire n_718;
wire n_1120;
wire n_719;
wire n_443;
wire n_714;
wire n_909;
wire n_997;
wire n_932;
wire n_612;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_508;
wire n_506;
wire n_1320;
wire n_737;
wire n_986;
wire n_509;
wire n_1317;
wire n_1281;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_733;
wire n_1489;
wire n_1376;
wire n_941;
wire n_981;
wire n_867;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_518;
wire n_505;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_381;
wire n_390;
wire n_1330;
wire n_481;
wire n_769;
wire n_1046;
wire n_934;
wire n_826;
wire n_886;
wire n_1221;
wire n_654;
wire n_1172;
wire n_379;
wire n_428;
wire n_1341;
wire n_570;
wire n_1361;
wire n_853;
wire n_377;
wire n_751;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_392;
wire n_704;
wire n_787;
wire n_961;
wire n_771;
wire n_1225;
wire n_522;
wire n_1287;
wire n_1262;
wire n_400;
wire n_930;
wire n_1411;
wire n_622;
wire n_1087;
wire n_386;
wire n_994;
wire n_848;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1247;
wire n_922;
wire n_816;
wire n_591;
wire n_1344;
wire n_631;
wire n_479;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_432;
wire n_839;
wire n_1210;
wire n_1364;
wire n_1250;
wire n_369;
wire n_871;
wire n_598;
wire n_685;
wire n_928;
wire n_608;
wire n_1367;
wire n_1460;
wire n_772;
wire n_499;
wire n_517;
wire n_402;
wire n_413;
wire n_1086;
wire n_796;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_903;
wire n_740;
wire n_384;
wire n_1404;
wire n_1315;
wire n_1061;
wire n_333;
wire n_1298;
wire n_462;
wire n_1193;
wire n_1255;
wire n_1113;
wire n_1226;
wire n_722;
wire n_1277;
wire n_844;
wire n_471;
wire n_852;
wire n_1487;
wire n_1028;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_1337;
wire n_632;
wire n_699;
wire n_979;
wire n_1245;
wire n_846;
wire n_465;
wire n_362;
wire n_1321;
wire n_585;
wire n_616;
wire n_745;
wire n_1103;
wire n_648;
wire n_1379;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_494;
wire n_641;
wire n_730;
wire n_1325;
wire n_354;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_695;
wire n_656;
wire n_1220;
wire n_437;
wire n_403;
wire n_453;
wire n_1130;
wire n_720;
wire n_863;
wire n_805;
wire n_1275;
wire n_712;
wire n_1042;
wire n_1402;
wire n_412;
wire n_657;
wire n_644;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_566;
wire n_565;
wire n_1448;
wire n_1398;
wire n_597;
wire n_1181;
wire n_1196;
wire n_651;
wire n_1340;
wire n_334;
wire n_811;
wire n_807;
wire n_835;
wire n_666;
wire n_1433;
wire n_1254;
wire n_1026;
wire n_1234;
wire n_364;
wire n_1138;
wire n_927;
wire n_1089;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_1018;
wire n_438;
wire n_713;
wire n_904;
wire n_1180;
wire n_1271;
wire n_533;
wire n_1251;

INVx2_ASAP7_75t_L g332 ( 
.A(n_34),
.Y(n_332)
);

CKINVDCx14_ASAP7_75t_R g333 ( 
.A(n_65),
.Y(n_333)
);

BUFx2_ASAP7_75t_L g334 ( 
.A(n_18),
.Y(n_334)
);

CKINVDCx20_ASAP7_75t_R g335 ( 
.A(n_176),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_97),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_259),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_105),
.Y(n_338)
);

BUFx3_ASAP7_75t_L g339 ( 
.A(n_167),
.Y(n_339)
);

INVx3_ASAP7_75t_L g340 ( 
.A(n_135),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_69),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_28),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_115),
.Y(n_343)
);

INVxp67_ASAP7_75t_SL g344 ( 
.A(n_227),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_213),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_36),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_11),
.Y(n_347)
);

INVx1_ASAP7_75t_SL g348 ( 
.A(n_256),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_29),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_161),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_255),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_303),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_314),
.Y(n_353)
);

CKINVDCx16_ASAP7_75t_R g354 ( 
.A(n_254),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_111),
.Y(n_355)
);

INVx3_ASAP7_75t_L g356 ( 
.A(n_191),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_249),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_162),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_117),
.Y(n_359)
);

INVx2_ASAP7_75t_L g360 ( 
.A(n_204),
.Y(n_360)
);

NOR2xp67_ASAP7_75t_L g361 ( 
.A(n_235),
.B(n_312),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_218),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_126),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_129),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_220),
.Y(n_365)
);

BUFx10_ASAP7_75t_L g366 ( 
.A(n_121),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_246),
.Y(n_367)
);

CKINVDCx20_ASAP7_75t_R g368 ( 
.A(n_300),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_132),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_206),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_79),
.Y(n_371)
);

INVx1_ASAP7_75t_SL g372 ( 
.A(n_2),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_221),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_107),
.Y(n_374)
);

CKINVDCx20_ASAP7_75t_R g375 ( 
.A(n_110),
.Y(n_375)
);

NOR2xp67_ASAP7_75t_L g376 ( 
.A(n_118),
.B(n_258),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_41),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_208),
.Y(n_378)
);

INVx2_ASAP7_75t_L g379 ( 
.A(n_120),
.Y(n_379)
);

HB1xp67_ASAP7_75t_L g380 ( 
.A(n_138),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_139),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_243),
.Y(n_382)
);

CKINVDCx20_ASAP7_75t_R g383 ( 
.A(n_287),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_37),
.Y(n_384)
);

INVxp67_ASAP7_75t_SL g385 ( 
.A(n_269),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_77),
.Y(n_386)
);

INVx2_ASAP7_75t_L g387 ( 
.A(n_301),
.Y(n_387)
);

INVx1_ASAP7_75t_SL g388 ( 
.A(n_252),
.Y(n_388)
);

BUFx6f_ASAP7_75t_L g389 ( 
.A(n_101),
.Y(n_389)
);

HB1xp67_ASAP7_75t_SL g390 ( 
.A(n_71),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_322),
.Y(n_391)
);

BUFx10_ASAP7_75t_L g392 ( 
.A(n_305),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_88),
.Y(n_393)
);

INVx2_ASAP7_75t_L g394 ( 
.A(n_284),
.Y(n_394)
);

BUFx6f_ASAP7_75t_L g395 ( 
.A(n_56),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_151),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_207),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_116),
.Y(n_398)
);

BUFx6f_ASAP7_75t_L g399 ( 
.A(n_123),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_33),
.Y(n_400)
);

CKINVDCx16_ASAP7_75t_R g401 ( 
.A(n_247),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_38),
.Y(n_402)
);

INVx1_ASAP7_75t_SL g403 ( 
.A(n_124),
.Y(n_403)
);

INVx2_ASAP7_75t_L g404 ( 
.A(n_328),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_152),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_229),
.Y(n_406)
);

INVx2_ASAP7_75t_L g407 ( 
.A(n_224),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_104),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_122),
.Y(n_409)
);

BUFx5_ASAP7_75t_L g410 ( 
.A(n_80),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_309),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_282),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_62),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_310),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_197),
.Y(n_415)
);

INVx2_ASAP7_75t_L g416 ( 
.A(n_302),
.Y(n_416)
);

NOR2xp67_ASAP7_75t_L g417 ( 
.A(n_299),
.B(n_146),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_127),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_327),
.Y(n_419)
);

BUFx3_ASAP7_75t_L g420 ( 
.A(n_196),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_145),
.Y(n_421)
);

INVx2_ASAP7_75t_L g422 ( 
.A(n_263),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_268),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_211),
.Y(n_424)
);

INVx2_ASAP7_75t_L g425 ( 
.A(n_200),
.Y(n_425)
);

BUFx6f_ASAP7_75t_L g426 ( 
.A(n_140),
.Y(n_426)
);

BUFx3_ASAP7_75t_L g427 ( 
.A(n_103),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_223),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_53),
.Y(n_429)
);

CKINVDCx14_ASAP7_75t_R g430 ( 
.A(n_306),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_264),
.Y(n_431)
);

CKINVDCx20_ASAP7_75t_R g432 ( 
.A(n_157),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_141),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_147),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_21),
.Y(n_435)
);

INVx1_ASAP7_75t_SL g436 ( 
.A(n_153),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_82),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_158),
.Y(n_438)
);

BUFx10_ASAP7_75t_L g439 ( 
.A(n_202),
.Y(n_439)
);

INVx2_ASAP7_75t_L g440 ( 
.A(n_78),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_50),
.Y(n_441)
);

CKINVDCx5p33_ASAP7_75t_R g442 ( 
.A(n_81),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_236),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_144),
.Y(n_444)
);

CKINVDCx5p33_ASAP7_75t_R g445 ( 
.A(n_37),
.Y(n_445)
);

CKINVDCx5p33_ASAP7_75t_R g446 ( 
.A(n_137),
.Y(n_446)
);

INVx2_ASAP7_75t_SL g447 ( 
.A(n_320),
.Y(n_447)
);

CKINVDCx5p33_ASAP7_75t_R g448 ( 
.A(n_185),
.Y(n_448)
);

CKINVDCx5p33_ASAP7_75t_R g449 ( 
.A(n_114),
.Y(n_449)
);

CKINVDCx5p33_ASAP7_75t_R g450 ( 
.A(n_251),
.Y(n_450)
);

BUFx5_ASAP7_75t_L g451 ( 
.A(n_325),
.Y(n_451)
);

BUFx2_ASAP7_75t_L g452 ( 
.A(n_248),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_240),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_143),
.Y(n_454)
);

CKINVDCx5p33_ASAP7_75t_R g455 ( 
.A(n_257),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_46),
.Y(n_456)
);

BUFx3_ASAP7_75t_L g457 ( 
.A(n_163),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_298),
.Y(n_458)
);

CKINVDCx5p33_ASAP7_75t_R g459 ( 
.A(n_34),
.Y(n_459)
);

CKINVDCx20_ASAP7_75t_R g460 ( 
.A(n_89),
.Y(n_460)
);

BUFx6f_ASAP7_75t_L g461 ( 
.A(n_20),
.Y(n_461)
);

INVx1_ASAP7_75t_SL g462 ( 
.A(n_273),
.Y(n_462)
);

BUFx3_ASAP7_75t_L g463 ( 
.A(n_27),
.Y(n_463)
);

BUFx5_ASAP7_75t_L g464 ( 
.A(n_199),
.Y(n_464)
);

CKINVDCx5p33_ASAP7_75t_R g465 ( 
.A(n_297),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_166),
.Y(n_466)
);

INVx1_ASAP7_75t_SL g467 ( 
.A(n_29),
.Y(n_467)
);

CKINVDCx5p33_ASAP7_75t_R g468 ( 
.A(n_296),
.Y(n_468)
);

CKINVDCx5p33_ASAP7_75t_R g469 ( 
.A(n_192),
.Y(n_469)
);

BUFx10_ASAP7_75t_L g470 ( 
.A(n_61),
.Y(n_470)
);

BUFx6f_ASAP7_75t_L g471 ( 
.A(n_20),
.Y(n_471)
);

CKINVDCx5p33_ASAP7_75t_R g472 ( 
.A(n_319),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_1),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_98),
.Y(n_474)
);

CKINVDCx5p33_ASAP7_75t_R g475 ( 
.A(n_154),
.Y(n_475)
);

CKINVDCx5p33_ASAP7_75t_R g476 ( 
.A(n_317),
.Y(n_476)
);

CKINVDCx5p33_ASAP7_75t_R g477 ( 
.A(n_96),
.Y(n_477)
);

CKINVDCx5p33_ASAP7_75t_R g478 ( 
.A(n_286),
.Y(n_478)
);

CKINVDCx5p33_ASAP7_75t_R g479 ( 
.A(n_9),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_186),
.Y(n_480)
);

CKINVDCx5p33_ASAP7_75t_R g481 ( 
.A(n_133),
.Y(n_481)
);

CKINVDCx20_ASAP7_75t_R g482 ( 
.A(n_1),
.Y(n_482)
);

CKINVDCx5p33_ASAP7_75t_R g483 ( 
.A(n_238),
.Y(n_483)
);

CKINVDCx5p33_ASAP7_75t_R g484 ( 
.A(n_233),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_311),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_136),
.Y(n_486)
);

CKINVDCx5p33_ASAP7_75t_R g487 ( 
.A(n_54),
.Y(n_487)
);

CKINVDCx5p33_ASAP7_75t_R g488 ( 
.A(n_265),
.Y(n_488)
);

CKINVDCx5p33_ASAP7_75t_R g489 ( 
.A(n_281),
.Y(n_489)
);

INVxp67_ASAP7_75t_L g490 ( 
.A(n_45),
.Y(n_490)
);

BUFx2_ASAP7_75t_L g491 ( 
.A(n_84),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_212),
.Y(n_492)
);

CKINVDCx5p33_ASAP7_75t_R g493 ( 
.A(n_178),
.Y(n_493)
);

CKINVDCx5p33_ASAP7_75t_R g494 ( 
.A(n_179),
.Y(n_494)
);

INVx2_ASAP7_75t_L g495 ( 
.A(n_275),
.Y(n_495)
);

INVx2_ASAP7_75t_L g496 ( 
.A(n_274),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_315),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_316),
.Y(n_498)
);

INVx1_ASAP7_75t_SL g499 ( 
.A(n_290),
.Y(n_499)
);

CKINVDCx16_ASAP7_75t_R g500 ( 
.A(n_142),
.Y(n_500)
);

CKINVDCx5p33_ASAP7_75t_R g501 ( 
.A(n_324),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_175),
.Y(n_502)
);

BUFx10_ASAP7_75t_L g503 ( 
.A(n_6),
.Y(n_503)
);

CKINVDCx5p33_ASAP7_75t_R g504 ( 
.A(n_45),
.Y(n_504)
);

CKINVDCx5p33_ASAP7_75t_R g505 ( 
.A(n_134),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_63),
.Y(n_506)
);

CKINVDCx5p33_ASAP7_75t_R g507 ( 
.A(n_250),
.Y(n_507)
);

CKINVDCx5p33_ASAP7_75t_R g508 ( 
.A(n_271),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_23),
.Y(n_509)
);

CKINVDCx5p33_ASAP7_75t_R g510 ( 
.A(n_261),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_222),
.Y(n_511)
);

BUFx3_ASAP7_75t_L g512 ( 
.A(n_27),
.Y(n_512)
);

CKINVDCx5p33_ASAP7_75t_R g513 ( 
.A(n_308),
.Y(n_513)
);

CKINVDCx5p33_ASAP7_75t_R g514 ( 
.A(n_168),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_11),
.Y(n_515)
);

CKINVDCx5p33_ASAP7_75t_R g516 ( 
.A(n_285),
.Y(n_516)
);

CKINVDCx5p33_ASAP7_75t_R g517 ( 
.A(n_326),
.Y(n_517)
);

INVx3_ASAP7_75t_L g518 ( 
.A(n_50),
.Y(n_518)
);

CKINVDCx20_ASAP7_75t_R g519 ( 
.A(n_323),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_278),
.Y(n_520)
);

CKINVDCx5p33_ASAP7_75t_R g521 ( 
.A(n_216),
.Y(n_521)
);

BUFx6f_ASAP7_75t_L g522 ( 
.A(n_289),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_188),
.Y(n_523)
);

BUFx6f_ASAP7_75t_L g524 ( 
.A(n_174),
.Y(n_524)
);

CKINVDCx5p33_ASAP7_75t_R g525 ( 
.A(n_64),
.Y(n_525)
);

BUFx6f_ASAP7_75t_L g526 ( 
.A(n_183),
.Y(n_526)
);

CKINVDCx5p33_ASAP7_75t_R g527 ( 
.A(n_93),
.Y(n_527)
);

CKINVDCx16_ASAP7_75t_R g528 ( 
.A(n_75),
.Y(n_528)
);

CKINVDCx20_ASAP7_75t_R g529 ( 
.A(n_321),
.Y(n_529)
);

CKINVDCx5p33_ASAP7_75t_R g530 ( 
.A(n_205),
.Y(n_530)
);

CKINVDCx5p33_ASAP7_75t_R g531 ( 
.A(n_231),
.Y(n_531)
);

CKINVDCx5p33_ASAP7_75t_R g532 ( 
.A(n_187),
.Y(n_532)
);

BUFx2_ASAP7_75t_L g533 ( 
.A(n_6),
.Y(n_533)
);

NOR2xp67_ASAP7_75t_L g534 ( 
.A(n_219),
.B(n_288),
.Y(n_534)
);

CKINVDCx5p33_ASAP7_75t_R g535 ( 
.A(n_232),
.Y(n_535)
);

BUFx8_ASAP7_75t_SL g536 ( 
.A(n_272),
.Y(n_536)
);

CKINVDCx5p33_ASAP7_75t_R g537 ( 
.A(n_184),
.Y(n_537)
);

CKINVDCx20_ASAP7_75t_R g538 ( 
.A(n_51),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_193),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_59),
.Y(n_540)
);

CKINVDCx5p33_ASAP7_75t_R g541 ( 
.A(n_24),
.Y(n_541)
);

CKINVDCx5p33_ASAP7_75t_R g542 ( 
.A(n_24),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_177),
.Y(n_543)
);

CKINVDCx5p33_ASAP7_75t_R g544 ( 
.A(n_214),
.Y(n_544)
);

CKINVDCx5p33_ASAP7_75t_R g545 ( 
.A(n_226),
.Y(n_545)
);

BUFx10_ASAP7_75t_L g546 ( 
.A(n_267),
.Y(n_546)
);

INVx1_ASAP7_75t_SL g547 ( 
.A(n_13),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_109),
.Y(n_548)
);

NOR2xp67_ASAP7_75t_L g549 ( 
.A(n_67),
.B(n_19),
.Y(n_549)
);

CKINVDCx5p33_ASAP7_75t_R g550 ( 
.A(n_85),
.Y(n_550)
);

CKINVDCx5p33_ASAP7_75t_R g551 ( 
.A(n_295),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_119),
.Y(n_552)
);

BUFx3_ASAP7_75t_L g553 ( 
.A(n_18),
.Y(n_553)
);

BUFx10_ASAP7_75t_L g554 ( 
.A(n_48),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_329),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_244),
.Y(n_556)
);

CKINVDCx5p33_ASAP7_75t_R g557 ( 
.A(n_19),
.Y(n_557)
);

INVx2_ASAP7_75t_L g558 ( 
.A(n_283),
.Y(n_558)
);

CKINVDCx5p33_ASAP7_75t_R g559 ( 
.A(n_47),
.Y(n_559)
);

CKINVDCx5p33_ASAP7_75t_R g560 ( 
.A(n_156),
.Y(n_560)
);

BUFx6f_ASAP7_75t_L g561 ( 
.A(n_25),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_155),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_209),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_461),
.Y(n_564)
);

AND2x4_ASAP7_75t_L g565 ( 
.A(n_339),
.B(n_0),
.Y(n_565)
);

AND2x2_ASAP7_75t_L g566 ( 
.A(n_334),
.B(n_0),
.Y(n_566)
);

BUFx6f_ASAP7_75t_L g567 ( 
.A(n_389),
.Y(n_567)
);

BUFx3_ASAP7_75t_L g568 ( 
.A(n_366),
.Y(n_568)
);

BUFx3_ASAP7_75t_L g569 ( 
.A(n_366),
.Y(n_569)
);

BUFx6f_ASAP7_75t_L g570 ( 
.A(n_389),
.Y(n_570)
);

BUFx12f_ASAP7_75t_L g571 ( 
.A(n_503),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_461),
.Y(n_572)
);

INVx2_ASAP7_75t_L g573 ( 
.A(n_461),
.Y(n_573)
);

AND2x6_ASAP7_75t_L g574 ( 
.A(n_340),
.B(n_52),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_L g575 ( 
.A(n_340),
.B(n_2),
.Y(n_575)
);

INVx2_ASAP7_75t_L g576 ( 
.A(n_471),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_471),
.Y(n_577)
);

AND2x4_ASAP7_75t_L g578 ( 
.A(n_420),
.B(n_427),
.Y(n_578)
);

INVx2_ASAP7_75t_L g579 ( 
.A(n_471),
.Y(n_579)
);

INVx2_ASAP7_75t_SL g580 ( 
.A(n_503),
.Y(n_580)
);

HB1xp67_ASAP7_75t_L g581 ( 
.A(n_533),
.Y(n_581)
);

BUFx6f_ASAP7_75t_L g582 ( 
.A(n_389),
.Y(n_582)
);

BUFx6f_ASAP7_75t_L g583 ( 
.A(n_395),
.Y(n_583)
);

AND2x4_ASAP7_75t_L g584 ( 
.A(n_457),
.B(n_3),
.Y(n_584)
);

BUFx3_ASAP7_75t_L g585 ( 
.A(n_392),
.Y(n_585)
);

BUFx6f_ASAP7_75t_L g586 ( 
.A(n_395),
.Y(n_586)
);

INVx2_ASAP7_75t_L g587 ( 
.A(n_561),
.Y(n_587)
);

HB1xp67_ASAP7_75t_L g588 ( 
.A(n_463),
.Y(n_588)
);

AND2x4_ASAP7_75t_L g589 ( 
.A(n_356),
.B(n_3),
.Y(n_589)
);

BUFx6f_ASAP7_75t_L g590 ( 
.A(n_395),
.Y(n_590)
);

OAI22x1_ASAP7_75t_R g591 ( 
.A1(n_482),
.A2(n_4),
.B1(n_5),
.B2(n_7),
.Y(n_591)
);

INVx5_ASAP7_75t_L g592 ( 
.A(n_399),
.Y(n_592)
);

INVx2_ASAP7_75t_L g593 ( 
.A(n_561),
.Y(n_593)
);

OAI21x1_ASAP7_75t_L g594 ( 
.A1(n_356),
.A2(n_57),
.B(n_55),
.Y(n_594)
);

BUFx6f_ASAP7_75t_L g595 ( 
.A(n_399),
.Y(n_595)
);

BUFx6f_ASAP7_75t_L g596 ( 
.A(n_399),
.Y(n_596)
);

HB1xp67_ASAP7_75t_L g597 ( 
.A(n_512),
.Y(n_597)
);

BUFx6f_ASAP7_75t_SL g598 ( 
.A(n_554),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_561),
.Y(n_599)
);

HB1xp67_ASAP7_75t_L g600 ( 
.A(n_553),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_518),
.Y(n_601)
);

OAI22xp5_ASAP7_75t_SL g602 ( 
.A1(n_372),
.A2(n_4),
.B1(n_5),
.B2(n_7),
.Y(n_602)
);

HB1xp67_ASAP7_75t_L g603 ( 
.A(n_346),
.Y(n_603)
);

BUFx2_ASAP7_75t_L g604 ( 
.A(n_347),
.Y(n_604)
);

AND2x2_ASAP7_75t_L g605 ( 
.A(n_452),
.B(n_8),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_L g606 ( 
.A(n_491),
.B(n_447),
.Y(n_606)
);

OAI22xp5_ASAP7_75t_L g607 ( 
.A1(n_333),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_607)
);

BUFx6f_ASAP7_75t_L g608 ( 
.A(n_426),
.Y(n_608)
);

INVx2_ASAP7_75t_L g609 ( 
.A(n_410),
.Y(n_609)
);

INVx5_ASAP7_75t_L g610 ( 
.A(n_426),
.Y(n_610)
);

BUFx12f_ASAP7_75t_L g611 ( 
.A(n_554),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_518),
.Y(n_612)
);

BUFx6f_ASAP7_75t_L g613 ( 
.A(n_426),
.Y(n_613)
);

OA21x2_ASAP7_75t_L g614 ( 
.A1(n_338),
.A2(n_10),
.B(n_12),
.Y(n_614)
);

INVx5_ASAP7_75t_L g615 ( 
.A(n_522),
.Y(n_615)
);

CKINVDCx16_ASAP7_75t_R g616 ( 
.A(n_354),
.Y(n_616)
);

INVx1_ASAP7_75t_SL g617 ( 
.A(n_467),
.Y(n_617)
);

BUFx6f_ASAP7_75t_L g618 ( 
.A(n_522),
.Y(n_618)
);

INVx2_ASAP7_75t_L g619 ( 
.A(n_410),
.Y(n_619)
);

HB1xp67_ASAP7_75t_L g620 ( 
.A(n_377),
.Y(n_620)
);

INVx2_ASAP7_75t_SL g621 ( 
.A(n_392),
.Y(n_621)
);

INVx5_ASAP7_75t_L g622 ( 
.A(n_522),
.Y(n_622)
);

INVx2_ASAP7_75t_L g623 ( 
.A(n_410),
.Y(n_623)
);

NOR2xp33_ASAP7_75t_L g624 ( 
.A(n_380),
.B(n_12),
.Y(n_624)
);

INVx2_ASAP7_75t_L g625 ( 
.A(n_410),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_332),
.Y(n_626)
);

AND2x4_ASAP7_75t_L g627 ( 
.A(n_360),
.B(n_14),
.Y(n_627)
);

BUFx8_ASAP7_75t_SL g628 ( 
.A(n_536),
.Y(n_628)
);

INVxp33_ASAP7_75t_SL g629 ( 
.A(n_384),
.Y(n_629)
);

HB1xp67_ASAP7_75t_L g630 ( 
.A(n_400),
.Y(n_630)
);

BUFx12f_ASAP7_75t_L g631 ( 
.A(n_439),
.Y(n_631)
);

CKINVDCx5p33_ASAP7_75t_R g632 ( 
.A(n_336),
.Y(n_632)
);

INVx2_ASAP7_75t_L g633 ( 
.A(n_410),
.Y(n_633)
);

BUFx6f_ASAP7_75t_L g634 ( 
.A(n_524),
.Y(n_634)
);

INVx2_ASAP7_75t_L g635 ( 
.A(n_451),
.Y(n_635)
);

BUFx6f_ASAP7_75t_L g636 ( 
.A(n_524),
.Y(n_636)
);

BUFx6f_ASAP7_75t_L g637 ( 
.A(n_524),
.Y(n_637)
);

HB1xp67_ASAP7_75t_L g638 ( 
.A(n_435),
.Y(n_638)
);

OAI22xp5_ASAP7_75t_L g639 ( 
.A1(n_430),
.A2(n_14),
.B1(n_15),
.B2(n_16),
.Y(n_639)
);

OAI21x1_ASAP7_75t_L g640 ( 
.A1(n_379),
.A2(n_60),
.B(n_58),
.Y(n_640)
);

INVx2_ASAP7_75t_L g641 ( 
.A(n_451),
.Y(n_641)
);

BUFx6f_ASAP7_75t_L g642 ( 
.A(n_526),
.Y(n_642)
);

BUFx6f_ASAP7_75t_L g643 ( 
.A(n_526),
.Y(n_643)
);

INVx2_ASAP7_75t_L g644 ( 
.A(n_451),
.Y(n_644)
);

BUFx6f_ASAP7_75t_L g645 ( 
.A(n_526),
.Y(n_645)
);

BUFx2_ASAP7_75t_L g646 ( 
.A(n_445),
.Y(n_646)
);

CKINVDCx5p33_ASAP7_75t_R g647 ( 
.A(n_337),
.Y(n_647)
);

BUFx8_ASAP7_75t_L g648 ( 
.A(n_342),
.Y(n_648)
);

BUFx12f_ASAP7_75t_L g649 ( 
.A(n_439),
.Y(n_649)
);

INVx2_ASAP7_75t_L g650 ( 
.A(n_451),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_349),
.Y(n_651)
);

BUFx2_ASAP7_75t_L g652 ( 
.A(n_459),
.Y(n_652)
);

BUFx12f_ASAP7_75t_L g653 ( 
.A(n_470),
.Y(n_653)
);

BUFx2_ASAP7_75t_L g654 ( 
.A(n_479),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_L g655 ( 
.A(n_387),
.B(n_15),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_402),
.Y(n_656)
);

INVx3_ASAP7_75t_L g657 ( 
.A(n_470),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_L g658 ( 
.A(n_394),
.B(n_16),
.Y(n_658)
);

OA21x2_ASAP7_75t_L g659 ( 
.A1(n_341),
.A2(n_17),
.B(n_21),
.Y(n_659)
);

OA21x2_ASAP7_75t_L g660 ( 
.A1(n_345),
.A2(n_357),
.B(n_355),
.Y(n_660)
);

XNOR2xp5_ASAP7_75t_L g661 ( 
.A(n_504),
.B(n_17),
.Y(n_661)
);

OA21x2_ASAP7_75t_L g662 ( 
.A1(n_359),
.A2(n_22),
.B(n_23),
.Y(n_662)
);

INVx5_ASAP7_75t_L g663 ( 
.A(n_546),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_441),
.Y(n_664)
);

AND2x4_ASAP7_75t_L g665 ( 
.A(n_404),
.B(n_22),
.Y(n_665)
);

INVx5_ASAP7_75t_L g666 ( 
.A(n_546),
.Y(n_666)
);

INVx2_ASAP7_75t_L g667 ( 
.A(n_451),
.Y(n_667)
);

BUFx6f_ASAP7_75t_L g668 ( 
.A(n_407),
.Y(n_668)
);

CKINVDCx16_ASAP7_75t_R g669 ( 
.A(n_401),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_L g670 ( 
.A(n_416),
.B(n_25),
.Y(n_670)
);

CKINVDCx5p33_ASAP7_75t_R g671 ( 
.A(n_343),
.Y(n_671)
);

OAI21x1_ASAP7_75t_L g672 ( 
.A1(n_422),
.A2(n_68),
.B(n_66),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_L g673 ( 
.A(n_425),
.B(n_26),
.Y(n_673)
);

BUFx3_ASAP7_75t_L g674 ( 
.A(n_350),
.Y(n_674)
);

INVx2_ASAP7_75t_L g675 ( 
.A(n_464),
.Y(n_675)
);

AOI22x1_ASAP7_75t_SL g676 ( 
.A1(n_541),
.A2(n_26),
.B1(n_28),
.B2(n_30),
.Y(n_676)
);

AND2x2_ASAP7_75t_L g677 ( 
.A(n_500),
.B(n_31),
.Y(n_677)
);

INVx2_ASAP7_75t_L g678 ( 
.A(n_464),
.Y(n_678)
);

OA21x2_ASAP7_75t_L g679 ( 
.A1(n_363),
.A2(n_31),
.B(n_32),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_456),
.Y(n_680)
);

NOR2xp33_ASAP7_75t_L g681 ( 
.A(n_348),
.B(n_32),
.Y(n_681)
);

BUFx3_ASAP7_75t_L g682 ( 
.A(n_351),
.Y(n_682)
);

INVx2_ASAP7_75t_L g683 ( 
.A(n_464),
.Y(n_683)
);

OA21x2_ASAP7_75t_L g684 ( 
.A1(n_364),
.A2(n_33),
.B(n_35),
.Y(n_684)
);

NOR2x1_ASAP7_75t_L g685 ( 
.A(n_361),
.B(n_70),
.Y(n_685)
);

CKINVDCx5p33_ASAP7_75t_R g686 ( 
.A(n_352),
.Y(n_686)
);

BUFx6f_ASAP7_75t_L g687 ( 
.A(n_440),
.Y(n_687)
);

AND2x2_ASAP7_75t_L g688 ( 
.A(n_528),
.B(n_35),
.Y(n_688)
);

BUFx2_ASAP7_75t_L g689 ( 
.A(n_542),
.Y(n_689)
);

HB1xp67_ASAP7_75t_L g690 ( 
.A(n_557),
.Y(n_690)
);

BUFx2_ASAP7_75t_L g691 ( 
.A(n_559),
.Y(n_691)
);

CKINVDCx5p33_ASAP7_75t_R g692 ( 
.A(n_353),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_L g693 ( 
.A(n_495),
.B(n_496),
.Y(n_693)
);

OAI22x1_ASAP7_75t_L g694 ( 
.A1(n_473),
.A2(n_36),
.B1(n_38),
.B2(n_39),
.Y(n_694)
);

NOR2x1_ASAP7_75t_L g695 ( 
.A(n_376),
.B(n_72),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_L g696 ( 
.A(n_558),
.B(n_39),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_L g697 ( 
.A(n_369),
.B(n_40),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_L g698 ( 
.A(n_374),
.B(n_40),
.Y(n_698)
);

INVx2_ASAP7_75t_L g699 ( 
.A(n_464),
.Y(n_699)
);

OAI22x1_ASAP7_75t_R g700 ( 
.A1(n_509),
.A2(n_41),
.B1(n_42),
.B2(n_43),
.Y(n_700)
);

INVx5_ASAP7_75t_L g701 ( 
.A(n_464),
.Y(n_701)
);

NOR2xp33_ASAP7_75t_L g702 ( 
.A(n_388),
.B(n_42),
.Y(n_702)
);

AND2x4_ASAP7_75t_L g703 ( 
.A(n_386),
.B(n_43),
.Y(n_703)
);

BUFx3_ASAP7_75t_L g704 ( 
.A(n_358),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_515),
.Y(n_705)
);

BUFx2_ASAP7_75t_L g706 ( 
.A(n_490),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_391),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_393),
.Y(n_708)
);

BUFx12f_ASAP7_75t_L g709 ( 
.A(n_362),
.Y(n_709)
);

HB1xp67_ASAP7_75t_L g710 ( 
.A(n_547),
.Y(n_710)
);

BUFx6f_ASAP7_75t_L g711 ( 
.A(n_396),
.Y(n_711)
);

BUFx3_ASAP7_75t_L g712 ( 
.A(n_365),
.Y(n_712)
);

BUFx12f_ASAP7_75t_L g713 ( 
.A(n_367),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_406),
.Y(n_714)
);

INVx2_ASAP7_75t_L g715 ( 
.A(n_418),
.Y(n_715)
);

OAI21x1_ASAP7_75t_L g716 ( 
.A1(n_563),
.A2(n_74),
.B(n_73),
.Y(n_716)
);

BUFx12f_ASAP7_75t_L g717 ( 
.A(n_370),
.Y(n_717)
);

INVx2_ASAP7_75t_L g718 ( 
.A(n_421),
.Y(n_718)
);

BUFx2_ASAP7_75t_L g719 ( 
.A(n_335),
.Y(n_719)
);

OA21x2_ASAP7_75t_L g720 ( 
.A1(n_424),
.A2(n_44),
.B(n_46),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_L g721 ( 
.A(n_433),
.B(n_44),
.Y(n_721)
);

INVx4_ASAP7_75t_L g722 ( 
.A(n_371),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_573),
.Y(n_723)
);

CKINVDCx5p33_ASAP7_75t_R g724 ( 
.A(n_628),
.Y(n_724)
);

HB1xp67_ASAP7_75t_L g725 ( 
.A(n_617),
.Y(n_725)
);

CKINVDCx5p33_ASAP7_75t_R g726 ( 
.A(n_632),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_576),
.Y(n_727)
);

CKINVDCx5p33_ASAP7_75t_R g728 ( 
.A(n_647),
.Y(n_728)
);

CKINVDCx5p33_ASAP7_75t_R g729 ( 
.A(n_671),
.Y(n_729)
);

CKINVDCx5p33_ASAP7_75t_R g730 ( 
.A(n_686),
.Y(n_730)
);

CKINVDCx5p33_ASAP7_75t_R g731 ( 
.A(n_692),
.Y(n_731)
);

CKINVDCx5p33_ASAP7_75t_R g732 ( 
.A(n_709),
.Y(n_732)
);

NOR2xp33_ASAP7_75t_R g733 ( 
.A(n_616),
.B(n_669),
.Y(n_733)
);

XOR2xp5_ASAP7_75t_L g734 ( 
.A(n_719),
.B(n_368),
.Y(n_734)
);

CKINVDCx5p33_ASAP7_75t_R g735 ( 
.A(n_713),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_579),
.Y(n_736)
);

INVx2_ASAP7_75t_L g737 ( 
.A(n_587),
.Y(n_737)
);

CKINVDCx5p33_ASAP7_75t_R g738 ( 
.A(n_717),
.Y(n_738)
);

NOR2xp33_ASAP7_75t_R g739 ( 
.A(n_657),
.B(n_375),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_593),
.Y(n_740)
);

CKINVDCx5p33_ASAP7_75t_R g741 ( 
.A(n_674),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_567),
.Y(n_742)
);

CKINVDCx5p33_ASAP7_75t_R g743 ( 
.A(n_682),
.Y(n_743)
);

NOR2xp33_ASAP7_75t_L g744 ( 
.A(n_606),
.B(n_403),
.Y(n_744)
);

CKINVDCx5p33_ASAP7_75t_R g745 ( 
.A(n_704),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_567),
.Y(n_746)
);

NOR2xp33_ASAP7_75t_R g747 ( 
.A(n_657),
.B(n_383),
.Y(n_747)
);

CKINVDCx20_ASAP7_75t_R g748 ( 
.A(n_712),
.Y(n_748)
);

INVx2_ASAP7_75t_L g749 ( 
.A(n_567),
.Y(n_749)
);

CKINVDCx5p33_ASAP7_75t_R g750 ( 
.A(n_629),
.Y(n_750)
);

CKINVDCx5p33_ASAP7_75t_R g751 ( 
.A(n_631),
.Y(n_751)
);

CKINVDCx20_ASAP7_75t_R g752 ( 
.A(n_604),
.Y(n_752)
);

AND2x2_ASAP7_75t_L g753 ( 
.A(n_603),
.B(n_436),
.Y(n_753)
);

CKINVDCx5p33_ASAP7_75t_R g754 ( 
.A(n_649),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_570),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_570),
.Y(n_756)
);

CKINVDCx5p33_ASAP7_75t_R g757 ( 
.A(n_653),
.Y(n_757)
);

NOR2xp33_ASAP7_75t_R g758 ( 
.A(n_571),
.B(n_432),
.Y(n_758)
);

CKINVDCx20_ASAP7_75t_R g759 ( 
.A(n_646),
.Y(n_759)
);

CKINVDCx5p33_ASAP7_75t_R g760 ( 
.A(n_722),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_570),
.Y(n_761)
);

CKINVDCx5p33_ASAP7_75t_R g762 ( 
.A(n_722),
.Y(n_762)
);

INVx2_ASAP7_75t_L g763 ( 
.A(n_582),
.Y(n_763)
);

CKINVDCx5p33_ASAP7_75t_R g764 ( 
.A(n_611),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_582),
.Y(n_765)
);

HB1xp67_ASAP7_75t_L g766 ( 
.A(n_710),
.Y(n_766)
);

NOR2xp33_ASAP7_75t_L g767 ( 
.A(n_605),
.B(n_462),
.Y(n_767)
);

CKINVDCx5p33_ASAP7_75t_R g768 ( 
.A(n_598),
.Y(n_768)
);

CKINVDCx5p33_ASAP7_75t_R g769 ( 
.A(n_598),
.Y(n_769)
);

BUFx6f_ASAP7_75t_L g770 ( 
.A(n_582),
.Y(n_770)
);

CKINVDCx20_ASAP7_75t_R g771 ( 
.A(n_652),
.Y(n_771)
);

AND2x6_ASAP7_75t_L g772 ( 
.A(n_589),
.B(n_434),
.Y(n_772)
);

CKINVDCx5p33_ASAP7_75t_R g773 ( 
.A(n_654),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_583),
.Y(n_774)
);

INVx2_ASAP7_75t_L g775 ( 
.A(n_583),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_583),
.Y(n_776)
);

CKINVDCx5p33_ASAP7_75t_R g777 ( 
.A(n_689),
.Y(n_777)
);

CKINVDCx5p33_ASAP7_75t_R g778 ( 
.A(n_691),
.Y(n_778)
);

CKINVDCx5p33_ASAP7_75t_R g779 ( 
.A(n_568),
.Y(n_779)
);

CKINVDCx5p33_ASAP7_75t_R g780 ( 
.A(n_569),
.Y(n_780)
);

HB1xp67_ASAP7_75t_L g781 ( 
.A(n_588),
.Y(n_781)
);

INVx1_ASAP7_75t_L g782 ( 
.A(n_586),
.Y(n_782)
);

AO22x2_ASAP7_75t_L g783 ( 
.A1(n_589),
.A2(n_453),
.B1(n_454),
.B2(n_437),
.Y(n_783)
);

CKINVDCx5p33_ASAP7_75t_R g784 ( 
.A(n_585),
.Y(n_784)
);

INVx1_ASAP7_75t_L g785 ( 
.A(n_586),
.Y(n_785)
);

CKINVDCx16_ASAP7_75t_R g786 ( 
.A(n_581),
.Y(n_786)
);

NAND2xp33_ASAP7_75t_R g787 ( 
.A(n_706),
.B(n_373),
.Y(n_787)
);

NOR2xp33_ASAP7_75t_R g788 ( 
.A(n_621),
.B(n_460),
.Y(n_788)
);

NAND2xp33_ASAP7_75t_R g789 ( 
.A(n_614),
.B(n_378),
.Y(n_789)
);

NOR2xp33_ASAP7_75t_R g790 ( 
.A(n_574),
.B(n_519),
.Y(n_790)
);

HB1xp67_ASAP7_75t_L g791 ( 
.A(n_597),
.Y(n_791)
);

CKINVDCx5p33_ASAP7_75t_R g792 ( 
.A(n_663),
.Y(n_792)
);

CKINVDCx5p33_ASAP7_75t_R g793 ( 
.A(n_663),
.Y(n_793)
);

NOR2xp33_ASAP7_75t_R g794 ( 
.A(n_574),
.B(n_529),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_586),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_L g796 ( 
.A(n_578),
.B(n_458),
.Y(n_796)
);

NOR2xp33_ASAP7_75t_R g797 ( 
.A(n_574),
.B(n_538),
.Y(n_797)
);

CKINVDCx5p33_ASAP7_75t_R g798 ( 
.A(n_666),
.Y(n_798)
);

CKINVDCx20_ASAP7_75t_R g799 ( 
.A(n_620),
.Y(n_799)
);

CKINVDCx5p33_ASAP7_75t_R g800 ( 
.A(n_666),
.Y(n_800)
);

INVx2_ASAP7_75t_L g801 ( 
.A(n_590),
.Y(n_801)
);

AND2x2_ASAP7_75t_L g802 ( 
.A(n_630),
.B(n_499),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_590),
.Y(n_803)
);

AND3x2_ASAP7_75t_L g804 ( 
.A(n_677),
.B(n_385),
.C(n_344),
.Y(n_804)
);

CKINVDCx16_ASAP7_75t_R g805 ( 
.A(n_638),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_595),
.Y(n_806)
);

CKINVDCx5p33_ASAP7_75t_R g807 ( 
.A(n_666),
.Y(n_807)
);

CKINVDCx5p33_ASAP7_75t_R g808 ( 
.A(n_690),
.Y(n_808)
);

CKINVDCx5p33_ASAP7_75t_R g809 ( 
.A(n_578),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_595),
.Y(n_810)
);

INVx2_ASAP7_75t_L g811 ( 
.A(n_595),
.Y(n_811)
);

CKINVDCx5p33_ASAP7_75t_R g812 ( 
.A(n_648),
.Y(n_812)
);

CKINVDCx16_ASAP7_75t_R g813 ( 
.A(n_688),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_596),
.Y(n_814)
);

CKINVDCx20_ASAP7_75t_R g815 ( 
.A(n_648),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_596),
.Y(n_816)
);

CKINVDCx5p33_ASAP7_75t_R g817 ( 
.A(n_600),
.Y(n_817)
);

NOR2xp33_ASAP7_75t_R g818 ( 
.A(n_574),
.B(n_381),
.Y(n_818)
);

CKINVDCx5p33_ASAP7_75t_R g819 ( 
.A(n_580),
.Y(n_819)
);

INVx2_ASAP7_75t_L g820 ( 
.A(n_608),
.Y(n_820)
);

CKINVDCx5p33_ASAP7_75t_R g821 ( 
.A(n_668),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_608),
.Y(n_822)
);

HB1xp67_ASAP7_75t_L g823 ( 
.A(n_661),
.Y(n_823)
);

CKINVDCx5p33_ASAP7_75t_R g824 ( 
.A(n_668),
.Y(n_824)
);

BUFx6f_ASAP7_75t_L g825 ( 
.A(n_770),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_L g826 ( 
.A(n_767),
.B(n_592),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_SL g827 ( 
.A(n_744),
.B(n_566),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_L g828 ( 
.A(n_821),
.B(n_592),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_SL g829 ( 
.A(n_725),
.B(n_681),
.Y(n_829)
);

NAND2xp33_ASAP7_75t_L g830 ( 
.A(n_790),
.B(n_575),
.Y(n_830)
);

INVxp33_ASAP7_75t_L g831 ( 
.A(n_725),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_749),
.Y(n_832)
);

BUFx6f_ASAP7_75t_L g833 ( 
.A(n_770),
.Y(n_833)
);

NOR2xp33_ASAP7_75t_L g834 ( 
.A(n_824),
.B(n_702),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_SL g835 ( 
.A(n_813),
.B(n_565),
.Y(n_835)
);

BUFx6f_ASAP7_75t_SL g836 ( 
.A(n_723),
.Y(n_836)
);

NOR2xp33_ASAP7_75t_L g837 ( 
.A(n_760),
.B(n_624),
.Y(n_837)
);

INVx5_ASAP7_75t_L g838 ( 
.A(n_770),
.Y(n_838)
);

BUFx6f_ASAP7_75t_L g839 ( 
.A(n_770),
.Y(n_839)
);

NOR2xp33_ASAP7_75t_L g840 ( 
.A(n_762),
.B(n_697),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_L g841 ( 
.A(n_772),
.B(n_592),
.Y(n_841)
);

INVx2_ASAP7_75t_L g842 ( 
.A(n_763),
.Y(n_842)
);

INVx2_ASAP7_75t_L g843 ( 
.A(n_775),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_L g844 ( 
.A(n_772),
.B(n_610),
.Y(n_844)
);

NOR2xp33_ASAP7_75t_L g845 ( 
.A(n_809),
.B(n_698),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_SL g846 ( 
.A(n_753),
.B(n_565),
.Y(n_846)
);

OR2x6_ASAP7_75t_L g847 ( 
.A(n_766),
.B(n_694),
.Y(n_847)
);

NOR2x1p5_ASAP7_75t_L g848 ( 
.A(n_768),
.B(n_721),
.Y(n_848)
);

INVxp33_ASAP7_75t_L g849 ( 
.A(n_766),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_L g850 ( 
.A(n_772),
.B(n_610),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_L g851 ( 
.A(n_772),
.B(n_610),
.Y(n_851)
);

INVx3_ASAP7_75t_L g852 ( 
.A(n_801),
.Y(n_852)
);

INVx2_ASAP7_75t_L g853 ( 
.A(n_811),
.Y(n_853)
);

CKINVDCx5p33_ASAP7_75t_R g854 ( 
.A(n_726),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_820),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_L g856 ( 
.A(n_772),
.B(n_615),
.Y(n_856)
);

NAND3xp33_ASAP7_75t_L g857 ( 
.A(n_796),
.B(n_658),
.C(n_655),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_SL g858 ( 
.A(n_802),
.B(n_584),
.Y(n_858)
);

BUFx6f_ASAP7_75t_L g859 ( 
.A(n_742),
.Y(n_859)
);

NOR3xp33_ASAP7_75t_L g860 ( 
.A(n_786),
.B(n_639),
.C(n_607),
.Y(n_860)
);

INVx4_ASAP7_75t_L g861 ( 
.A(n_741),
.Y(n_861)
);

AOI221xp5_ASAP7_75t_L g862 ( 
.A1(n_823),
.A2(n_602),
.B1(n_665),
.B2(n_627),
.C(n_703),
.Y(n_862)
);

NOR2xp33_ASAP7_75t_L g863 ( 
.A(n_728),
.B(n_729),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_SL g864 ( 
.A(n_739),
.B(n_584),
.Y(n_864)
);

INVxp33_ASAP7_75t_L g865 ( 
.A(n_781),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_L g866 ( 
.A(n_783),
.B(n_615),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_L g867 ( 
.A(n_783),
.B(n_615),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_L g868 ( 
.A(n_783),
.B(n_622),
.Y(n_868)
);

INVxp67_ASAP7_75t_L g869 ( 
.A(n_787),
.Y(n_869)
);

BUFx6f_ASAP7_75t_L g870 ( 
.A(n_746),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_SL g871 ( 
.A(n_747),
.B(n_627),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_755),
.Y(n_872)
);

NAND3xp33_ASAP7_75t_L g873 ( 
.A(n_781),
.B(n_791),
.C(n_808),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_SL g874 ( 
.A(n_819),
.B(n_665),
.Y(n_874)
);

INVx2_ASAP7_75t_L g875 ( 
.A(n_737),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_SL g876 ( 
.A(n_788),
.B(n_703),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_756),
.Y(n_877)
);

NOR2xp33_ASAP7_75t_L g878 ( 
.A(n_730),
.B(n_693),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_761),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_765),
.Y(n_880)
);

INVxp67_ASAP7_75t_L g881 ( 
.A(n_791),
.Y(n_881)
);

NOR2xp33_ASAP7_75t_L g882 ( 
.A(n_731),
.B(n_714),
.Y(n_882)
);

INVx2_ASAP7_75t_L g883 ( 
.A(n_774),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_776),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_782),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_785),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_795),
.Y(n_887)
);

INVx2_ASAP7_75t_L g888 ( 
.A(n_803),
.Y(n_888)
);

INVx2_ASAP7_75t_L g889 ( 
.A(n_806),
.Y(n_889)
);

NOR2xp33_ASAP7_75t_L g890 ( 
.A(n_743),
.B(n_745),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_SL g891 ( 
.A(n_817),
.B(n_382),
.Y(n_891)
);

INVxp67_ASAP7_75t_L g892 ( 
.A(n_734),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_SL g893 ( 
.A(n_779),
.B(n_780),
.Y(n_893)
);

NOR2xp33_ASAP7_75t_L g894 ( 
.A(n_784),
.B(n_670),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_SL g895 ( 
.A(n_773),
.B(n_397),
.Y(n_895)
);

INVx1_ASAP7_75t_L g896 ( 
.A(n_810),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_SL g897 ( 
.A(n_777),
.B(n_398),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_L g898 ( 
.A(n_814),
.B(n_622),
.Y(n_898)
);

INVx2_ASAP7_75t_L g899 ( 
.A(n_816),
.Y(n_899)
);

INVx1_ASAP7_75t_SL g900 ( 
.A(n_752),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_L g901 ( 
.A(n_822),
.B(n_622),
.Y(n_901)
);

INVx1_ASAP7_75t_L g902 ( 
.A(n_727),
.Y(n_902)
);

BUFx6f_ASAP7_75t_L g903 ( 
.A(n_736),
.Y(n_903)
);

INVx2_ASAP7_75t_SL g904 ( 
.A(n_778),
.Y(n_904)
);

NOR2xp67_ASAP7_75t_L g905 ( 
.A(n_750),
.B(n_701),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_740),
.Y(n_906)
);

CKINVDCx20_ASAP7_75t_R g907 ( 
.A(n_748),
.Y(n_907)
);

NOR2xp33_ASAP7_75t_L g908 ( 
.A(n_804),
.B(n_673),
.Y(n_908)
);

NOR3xp33_ASAP7_75t_L g909 ( 
.A(n_805),
.B(n_696),
.C(n_549),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_SL g910 ( 
.A(n_794),
.B(n_405),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_804),
.Y(n_911)
);

INVx2_ASAP7_75t_L g912 ( 
.A(n_792),
.Y(n_912)
);

NOR2xp33_ASAP7_75t_L g913 ( 
.A(n_793),
.B(n_715),
.Y(n_913)
);

NAND2xp33_ASAP7_75t_L g914 ( 
.A(n_797),
.B(n_685),
.Y(n_914)
);

AND2x4_ASAP7_75t_L g915 ( 
.A(n_798),
.B(n_601),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_SL g916 ( 
.A(n_800),
.B(n_408),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_807),
.Y(n_917)
);

NOR2xp33_ASAP7_75t_L g918 ( 
.A(n_769),
.B(n_718),
.Y(n_918)
);

NAND2xp5_ASAP7_75t_L g919 ( 
.A(n_818),
.B(n_660),
.Y(n_919)
);

HB1xp67_ASAP7_75t_L g920 ( 
.A(n_831),
.Y(n_920)
);

NAND3xp33_ASAP7_75t_L g921 ( 
.A(n_827),
.B(n_789),
.C(n_708),
.Y(n_921)
);

INVx1_ASAP7_75t_L g922 ( 
.A(n_875),
.Y(n_922)
);

NAND2xp5_ASAP7_75t_L g923 ( 
.A(n_878),
.B(n_660),
.Y(n_923)
);

AOI22xp5_ASAP7_75t_L g924 ( 
.A1(n_908),
.A2(n_759),
.B1(n_771),
.B2(n_799),
.Y(n_924)
);

NAND3xp33_ASAP7_75t_L g925 ( 
.A(n_862),
.B(n_708),
.C(n_707),
.Y(n_925)
);

CKINVDCx5p33_ASAP7_75t_R g926 ( 
.A(n_854),
.Y(n_926)
);

OAI22xp5_ASAP7_75t_L g927 ( 
.A1(n_919),
.A2(n_390),
.B1(n_474),
.B2(n_466),
.Y(n_927)
);

NAND2x1p5_ASAP7_75t_L g928 ( 
.A(n_861),
.B(n_594),
.Y(n_928)
);

INVxp67_ASAP7_75t_L g929 ( 
.A(n_882),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_SL g930 ( 
.A(n_869),
.B(n_733),
.Y(n_930)
);

BUFx2_ASAP7_75t_L g931 ( 
.A(n_907),
.Y(n_931)
);

AND2x4_ASAP7_75t_L g932 ( 
.A(n_902),
.B(n_664),
.Y(n_932)
);

NOR2xp33_ASAP7_75t_L g933 ( 
.A(n_840),
.B(n_812),
.Y(n_933)
);

BUFx3_ASAP7_75t_L g934 ( 
.A(n_903),
.Y(n_934)
);

NAND2xp5_ASAP7_75t_L g935 ( 
.A(n_894),
.B(n_668),
.Y(n_935)
);

OAI22x1_ASAP7_75t_SL g936 ( 
.A1(n_900),
.A2(n_591),
.B1(n_724),
.B2(n_815),
.Y(n_936)
);

BUFx2_ASAP7_75t_L g937 ( 
.A(n_911),
.Y(n_937)
);

NAND2xp5_ASAP7_75t_L g938 ( 
.A(n_837),
.B(n_687),
.Y(n_938)
);

INVx2_ASAP7_75t_L g939 ( 
.A(n_906),
.Y(n_939)
);

INVx2_ASAP7_75t_L g940 ( 
.A(n_842),
.Y(n_940)
);

INVx1_ASAP7_75t_L g941 ( 
.A(n_843),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_L g942 ( 
.A(n_845),
.B(n_687),
.Y(n_942)
);

NOR2xp33_ASAP7_75t_L g943 ( 
.A(n_865),
.B(n_732),
.Y(n_943)
);

AOI22xp5_ASAP7_75t_L g944 ( 
.A1(n_830),
.A2(n_695),
.B1(n_411),
.B2(n_412),
.Y(n_944)
);

AND2x2_ASAP7_75t_SL g945 ( 
.A(n_860),
.B(n_909),
.Y(n_945)
);

NOR2xp33_ASAP7_75t_L g946 ( 
.A(n_849),
.B(n_735),
.Y(n_946)
);

INVx1_ASAP7_75t_L g947 ( 
.A(n_853),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_L g948 ( 
.A(n_834),
.B(n_687),
.Y(n_948)
);

NOR2xp33_ASAP7_75t_L g949 ( 
.A(n_871),
.B(n_738),
.Y(n_949)
);

INVx1_ASAP7_75t_L g950 ( 
.A(n_832),
.Y(n_950)
);

AND2x2_ASAP7_75t_SL g951 ( 
.A(n_863),
.B(n_614),
.Y(n_951)
);

BUFx4f_ASAP7_75t_L g952 ( 
.A(n_904),
.Y(n_952)
);

BUFx3_ASAP7_75t_L g953 ( 
.A(n_903),
.Y(n_953)
);

NOR2xp33_ASAP7_75t_L g954 ( 
.A(n_829),
.B(n_751),
.Y(n_954)
);

BUFx2_ASAP7_75t_L g955 ( 
.A(n_881),
.Y(n_955)
);

INVx2_ASAP7_75t_L g956 ( 
.A(n_903),
.Y(n_956)
);

AOI21xp5_ASAP7_75t_L g957 ( 
.A1(n_914),
.A2(n_844),
.B(n_841),
.Y(n_957)
);

AOI22xp5_ASAP7_75t_L g958 ( 
.A1(n_846),
.A2(n_413),
.B1(n_414),
.B2(n_409),
.Y(n_958)
);

NAND2xp5_ASAP7_75t_SL g959 ( 
.A(n_858),
.B(n_758),
.Y(n_959)
);

NAND2xp5_ASAP7_75t_SL g960 ( 
.A(n_905),
.B(n_864),
.Y(n_960)
);

NAND2xp5_ASAP7_75t_SL g961 ( 
.A(n_861),
.B(n_754),
.Y(n_961)
);

INVx2_ASAP7_75t_L g962 ( 
.A(n_852),
.Y(n_962)
);

INVx2_ASAP7_75t_L g963 ( 
.A(n_852),
.Y(n_963)
);

NAND2xp5_ASAP7_75t_L g964 ( 
.A(n_826),
.B(n_480),
.Y(n_964)
);

INVx1_ASAP7_75t_L g965 ( 
.A(n_855),
.Y(n_965)
);

INVx1_ASAP7_75t_L g966 ( 
.A(n_872),
.Y(n_966)
);

NAND2x1_ASAP7_75t_L g967 ( 
.A(n_825),
.B(n_659),
.Y(n_967)
);

HB1xp67_ASAP7_75t_L g968 ( 
.A(n_835),
.Y(n_968)
);

INVx2_ASAP7_75t_SL g969 ( 
.A(n_915),
.Y(n_969)
);

BUFx6f_ASAP7_75t_L g970 ( 
.A(n_825),
.Y(n_970)
);

AND2x2_ASAP7_75t_L g971 ( 
.A(n_890),
.B(n_757),
.Y(n_971)
);

NOR2xp33_ASAP7_75t_L g972 ( 
.A(n_876),
.B(n_764),
.Y(n_972)
);

NAND2xp5_ASAP7_75t_L g973 ( 
.A(n_857),
.B(n_859),
.Y(n_973)
);

INVxp67_ASAP7_75t_L g974 ( 
.A(n_874),
.Y(n_974)
);

AND2x2_ASAP7_75t_L g975 ( 
.A(n_915),
.B(n_651),
.Y(n_975)
);

NOR2xp33_ASAP7_75t_L g976 ( 
.A(n_873),
.B(n_895),
.Y(n_976)
);

AND2x4_ASAP7_75t_L g977 ( 
.A(n_883),
.B(n_651),
.Y(n_977)
);

INVx2_ASAP7_75t_SL g978 ( 
.A(n_888),
.Y(n_978)
);

AND2x4_ASAP7_75t_L g979 ( 
.A(n_889),
.B(n_656),
.Y(n_979)
);

INVx1_ASAP7_75t_L g980 ( 
.A(n_877),
.Y(n_980)
);

BUFx3_ASAP7_75t_L g981 ( 
.A(n_859),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_L g982 ( 
.A(n_859),
.B(n_870),
.Y(n_982)
);

NOR2xp33_ASAP7_75t_L g983 ( 
.A(n_897),
.B(n_415),
.Y(n_983)
);

INVx3_ASAP7_75t_L g984 ( 
.A(n_899),
.Y(n_984)
);

NAND2xp5_ASAP7_75t_L g985 ( 
.A(n_870),
.B(n_485),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_SL g986 ( 
.A(n_866),
.B(n_419),
.Y(n_986)
);

NAND2xp5_ASAP7_75t_L g987 ( 
.A(n_870),
.B(n_486),
.Y(n_987)
);

INVx1_ASAP7_75t_L g988 ( 
.A(n_879),
.Y(n_988)
);

NAND2xp5_ASAP7_75t_SL g989 ( 
.A(n_867),
.B(n_423),
.Y(n_989)
);

AOI22xp5_ASAP7_75t_L g990 ( 
.A1(n_910),
.A2(n_428),
.B1(n_431),
.B2(n_429),
.Y(n_990)
);

INVx4_ASAP7_75t_L g991 ( 
.A(n_825),
.Y(n_991)
);

INVx1_ASAP7_75t_L g992 ( 
.A(n_880),
.Y(n_992)
);

BUFx8_ASAP7_75t_L g993 ( 
.A(n_836),
.Y(n_993)
);

NOR3xp33_ASAP7_75t_SL g994 ( 
.A(n_891),
.B(n_700),
.C(n_442),
.Y(n_994)
);

NOR2xp33_ASAP7_75t_R g995 ( 
.A(n_917),
.B(n_438),
.Y(n_995)
);

INVx2_ASAP7_75t_SL g996 ( 
.A(n_884),
.Y(n_996)
);

NAND2xp5_ASAP7_75t_L g997 ( 
.A(n_913),
.B(n_492),
.Y(n_997)
);

AND2x2_ASAP7_75t_L g998 ( 
.A(n_918),
.B(n_656),
.Y(n_998)
);

NAND2xp5_ASAP7_75t_SL g999 ( 
.A(n_868),
.B(n_912),
.Y(n_999)
);

INVx1_ASAP7_75t_L g1000 ( 
.A(n_885),
.Y(n_1000)
);

INVx1_ASAP7_75t_L g1001 ( 
.A(n_886),
.Y(n_1001)
);

INVx1_ASAP7_75t_L g1002 ( 
.A(n_887),
.Y(n_1002)
);

INVxp67_ASAP7_75t_L g1003 ( 
.A(n_847),
.Y(n_1003)
);

NAND2xp33_ASAP7_75t_SL g1004 ( 
.A(n_848),
.B(n_443),
.Y(n_1004)
);

AOI22xp33_ASAP7_75t_SL g1005 ( 
.A1(n_847),
.A2(n_676),
.B1(n_662),
.B2(n_659),
.Y(n_1005)
);

NAND2xp5_ASAP7_75t_L g1006 ( 
.A(n_896),
.B(n_497),
.Y(n_1006)
);

INVx5_ASAP7_75t_L g1007 ( 
.A(n_833),
.Y(n_1007)
);

INVx3_ASAP7_75t_L g1008 ( 
.A(n_833),
.Y(n_1008)
);

BUFx6f_ASAP7_75t_L g1009 ( 
.A(n_833),
.Y(n_1009)
);

INVxp67_ASAP7_75t_L g1010 ( 
.A(n_836),
.Y(n_1010)
);

AOI22xp33_ASAP7_75t_L g1011 ( 
.A1(n_850),
.A2(n_679),
.B1(n_684),
.B2(n_662),
.Y(n_1011)
);

INVx1_ASAP7_75t_L g1012 ( 
.A(n_898),
.Y(n_1012)
);

INVx1_ASAP7_75t_L g1013 ( 
.A(n_901),
.Y(n_1013)
);

NOR2xp33_ASAP7_75t_L g1014 ( 
.A(n_893),
.B(n_444),
.Y(n_1014)
);

INVx5_ASAP7_75t_L g1015 ( 
.A(n_839),
.Y(n_1015)
);

NAND2xp5_ASAP7_75t_SL g1016 ( 
.A(n_828),
.B(n_446),
.Y(n_1016)
);

INVx1_ASAP7_75t_L g1017 ( 
.A(n_839),
.Y(n_1017)
);

AND2x2_ASAP7_75t_L g1018 ( 
.A(n_916),
.B(n_680),
.Y(n_1018)
);

INVxp67_ASAP7_75t_L g1019 ( 
.A(n_892),
.Y(n_1019)
);

INVx1_ASAP7_75t_SL g1020 ( 
.A(n_839),
.Y(n_1020)
);

AOI22xp33_ASAP7_75t_SL g1021 ( 
.A1(n_851),
.A2(n_676),
.B1(n_684),
.B2(n_679),
.Y(n_1021)
);

AOI21xp5_ASAP7_75t_L g1022 ( 
.A1(n_923),
.A2(n_856),
.B(n_716),
.Y(n_1022)
);

AOI21xp5_ASAP7_75t_L g1023 ( 
.A1(n_957),
.A2(n_838),
.B(n_672),
.Y(n_1023)
);

INVx2_ASAP7_75t_L g1024 ( 
.A(n_1002),
.Y(n_1024)
);

NAND2xp5_ASAP7_75t_L g1025 ( 
.A(n_929),
.B(n_498),
.Y(n_1025)
);

A2O1A1Ixp33_ASAP7_75t_L g1026 ( 
.A1(n_921),
.A2(n_534),
.B(n_417),
.C(n_506),
.Y(n_1026)
);

AND2x4_ASAP7_75t_L g1027 ( 
.A(n_969),
.B(n_680),
.Y(n_1027)
);

A2O1A1Ixp33_ASAP7_75t_L g1028 ( 
.A1(n_976),
.A2(n_511),
.B(n_520),
.C(n_502),
.Y(n_1028)
);

NOR2xp33_ASAP7_75t_R g1029 ( 
.A(n_926),
.B(n_448),
.Y(n_1029)
);

NAND2xp5_ASAP7_75t_L g1030 ( 
.A(n_938),
.B(n_523),
.Y(n_1030)
);

OAI22xp5_ASAP7_75t_L g1031 ( 
.A1(n_951),
.A2(n_540),
.B1(n_543),
.B2(n_539),
.Y(n_1031)
);

O2A1O1Ixp5_ASAP7_75t_L g1032 ( 
.A1(n_967),
.A2(n_552),
.B(n_555),
.C(n_548),
.Y(n_1032)
);

AOI21xp5_ASAP7_75t_L g1033 ( 
.A1(n_982),
.A2(n_838),
.B(n_640),
.Y(n_1033)
);

HB1xp67_ASAP7_75t_L g1034 ( 
.A(n_920),
.Y(n_1034)
);

AND2x4_ASAP7_75t_L g1035 ( 
.A(n_932),
.B(n_705),
.Y(n_1035)
);

OAI22xp5_ASAP7_75t_L g1036 ( 
.A1(n_973),
.A2(n_562),
.B1(n_556),
.B2(n_720),
.Y(n_1036)
);

NAND2xp5_ASAP7_75t_L g1037 ( 
.A(n_998),
.B(n_720),
.Y(n_1037)
);

NOR2xp33_ASAP7_75t_L g1038 ( 
.A(n_933),
.B(n_955),
.Y(n_1038)
);

AND2x4_ASAP7_75t_L g1039 ( 
.A(n_932),
.B(n_705),
.Y(n_1039)
);

NAND2xp33_ASAP7_75t_SL g1040 ( 
.A(n_995),
.B(n_449),
.Y(n_1040)
);

AOI21xp5_ASAP7_75t_L g1041 ( 
.A1(n_1011),
.A2(n_838),
.B(n_618),
.Y(n_1041)
);

OR2x6_ASAP7_75t_L g1042 ( 
.A(n_931),
.B(n_626),
.Y(n_1042)
);

NOR2xp33_ASAP7_75t_L g1043 ( 
.A(n_974),
.B(n_450),
.Y(n_1043)
);

A2O1A1Ixp33_ASAP7_75t_SL g1044 ( 
.A1(n_983),
.A2(n_1014),
.B(n_1012),
.C(n_1013),
.Y(n_1044)
);

INVx1_ASAP7_75t_L g1045 ( 
.A(n_977),
.Y(n_1045)
);

NAND2xp5_ASAP7_75t_L g1046 ( 
.A(n_948),
.B(n_455),
.Y(n_1046)
);

BUFx2_ASAP7_75t_L g1047 ( 
.A(n_1003),
.Y(n_1047)
);

O2A1O1Ixp33_ASAP7_75t_L g1048 ( 
.A1(n_927),
.A2(n_707),
.B(n_612),
.C(n_601),
.Y(n_1048)
);

INVx1_ASAP7_75t_L g1049 ( 
.A(n_977),
.Y(n_1049)
);

AOI21xp5_ASAP7_75t_L g1050 ( 
.A1(n_1007),
.A2(n_618),
.B(n_613),
.Y(n_1050)
);

AOI22xp33_ASAP7_75t_L g1051 ( 
.A1(n_1021),
.A2(n_619),
.B1(n_623),
.B2(n_609),
.Y(n_1051)
);

INVx1_ASAP7_75t_L g1052 ( 
.A(n_979),
.Y(n_1052)
);

AOI21xp5_ASAP7_75t_L g1053 ( 
.A1(n_1007),
.A2(n_1015),
.B(n_935),
.Y(n_1053)
);

AOI21xp5_ASAP7_75t_L g1054 ( 
.A1(n_1007),
.A2(n_618),
.B(n_613),
.Y(n_1054)
);

NAND2xp5_ASAP7_75t_L g1055 ( 
.A(n_942),
.B(n_465),
.Y(n_1055)
);

AOI21xp5_ASAP7_75t_L g1056 ( 
.A1(n_1015),
.A2(n_634),
.B(n_613),
.Y(n_1056)
);

BUFx2_ASAP7_75t_L g1057 ( 
.A(n_937),
.Y(n_1057)
);

NAND2xp5_ASAP7_75t_SL g1058 ( 
.A(n_952),
.B(n_468),
.Y(n_1058)
);

INVxp67_ASAP7_75t_L g1059 ( 
.A(n_975),
.Y(n_1059)
);

BUFx3_ASAP7_75t_L g1060 ( 
.A(n_952),
.Y(n_1060)
);

BUFx4f_ASAP7_75t_L g1061 ( 
.A(n_945),
.Y(n_1061)
);

NOR2xp33_ASAP7_75t_L g1062 ( 
.A(n_968),
.B(n_469),
.Y(n_1062)
);

NAND2xp5_ASAP7_75t_SL g1063 ( 
.A(n_934),
.B(n_472),
.Y(n_1063)
);

CKINVDCx16_ASAP7_75t_R g1064 ( 
.A(n_924),
.Y(n_1064)
);

O2A1O1Ixp33_ASAP7_75t_L g1065 ( 
.A1(n_999),
.A2(n_989),
.B(n_986),
.C(n_997),
.Y(n_1065)
);

NAND2xp5_ASAP7_75t_L g1066 ( 
.A(n_1018),
.B(n_475),
.Y(n_1066)
);

INVx1_ASAP7_75t_L g1067 ( 
.A(n_979),
.Y(n_1067)
);

INVx3_ASAP7_75t_L g1068 ( 
.A(n_1008),
.Y(n_1068)
);

OAI21xp33_ASAP7_75t_L g1069 ( 
.A1(n_925),
.A2(n_626),
.B(n_612),
.Y(n_1069)
);

NAND2xp5_ASAP7_75t_L g1070 ( 
.A(n_956),
.B(n_476),
.Y(n_1070)
);

CKINVDCx5p33_ASAP7_75t_R g1071 ( 
.A(n_971),
.Y(n_1071)
);

INVx2_ASAP7_75t_L g1072 ( 
.A(n_922),
.Y(n_1072)
);

INVx1_ASAP7_75t_L g1073 ( 
.A(n_966),
.Y(n_1073)
);

A2O1A1Ixp33_ASAP7_75t_L g1074 ( 
.A1(n_949),
.A2(n_625),
.B(n_633),
.C(n_699),
.Y(n_1074)
);

CKINVDCx11_ASAP7_75t_R g1075 ( 
.A(n_936),
.Y(n_1075)
);

NAND2xp5_ASAP7_75t_L g1076 ( 
.A(n_964),
.B(n_477),
.Y(n_1076)
);

AOI21xp5_ASAP7_75t_L g1077 ( 
.A1(n_1015),
.A2(n_636),
.B(n_634),
.Y(n_1077)
);

OAI21xp5_ASAP7_75t_L g1078 ( 
.A1(n_928),
.A2(n_641),
.B(n_635),
.Y(n_1078)
);

A2O1A1Ixp33_ASAP7_75t_L g1079 ( 
.A1(n_972),
.A2(n_644),
.B(n_650),
.C(n_683),
.Y(n_1079)
);

INVx1_ASAP7_75t_L g1080 ( 
.A(n_980),
.Y(n_1080)
);

O2A1O1Ixp5_ASAP7_75t_L g1081 ( 
.A1(n_939),
.A2(n_678),
.B(n_675),
.C(n_667),
.Y(n_1081)
);

AOI21xp5_ASAP7_75t_L g1082 ( 
.A1(n_991),
.A2(n_636),
.B(n_634),
.Y(n_1082)
);

AOI22xp5_ASAP7_75t_L g1083 ( 
.A1(n_988),
.A2(n_527),
.B1(n_481),
.B2(n_483),
.Y(n_1083)
);

INVx2_ASAP7_75t_L g1084 ( 
.A(n_940),
.Y(n_1084)
);

A2O1A1Ixp33_ASAP7_75t_L g1085 ( 
.A1(n_992),
.A2(n_530),
.B(n_484),
.C(n_487),
.Y(n_1085)
);

OAI22xp5_ASAP7_75t_L g1086 ( 
.A1(n_1005),
.A2(n_531),
.B1(n_488),
.B2(n_489),
.Y(n_1086)
);

HB1xp67_ASAP7_75t_L g1087 ( 
.A(n_1020),
.Y(n_1087)
);

OAI22xp5_ASAP7_75t_L g1088 ( 
.A1(n_1000),
.A2(n_535),
.B1(n_493),
.B2(n_494),
.Y(n_1088)
);

OAI22xp5_ASAP7_75t_L g1089 ( 
.A1(n_1001),
.A2(n_537),
.B1(n_501),
.B2(n_505),
.Y(n_1089)
);

OAI22xp5_ASAP7_75t_L g1090 ( 
.A1(n_960),
.A2(n_545),
.B1(n_507),
.B2(n_508),
.Y(n_1090)
);

NAND2xp5_ASAP7_75t_L g1091 ( 
.A(n_953),
.B(n_478),
.Y(n_1091)
);

INVx4_ASAP7_75t_L g1092 ( 
.A(n_970),
.Y(n_1092)
);

NOR2xp33_ASAP7_75t_L g1093 ( 
.A(n_1019),
.B(n_510),
.Y(n_1093)
);

NAND2xp5_ASAP7_75t_L g1094 ( 
.A(n_996),
.B(n_941),
.Y(n_1094)
);

HB1xp67_ASAP7_75t_L g1095 ( 
.A(n_978),
.Y(n_1095)
);

NAND2xp5_ASAP7_75t_L g1096 ( 
.A(n_947),
.B(n_513),
.Y(n_1096)
);

INVx3_ASAP7_75t_SL g1097 ( 
.A(n_930),
.Y(n_1097)
);

BUFx2_ASAP7_75t_L g1098 ( 
.A(n_1010),
.Y(n_1098)
);

A2O1A1Ixp33_ASAP7_75t_L g1099 ( 
.A1(n_954),
.A2(n_560),
.B(n_516),
.C(n_517),
.Y(n_1099)
);

A2O1A1Ixp33_ASAP7_75t_L g1100 ( 
.A1(n_950),
.A2(n_514),
.B(n_521),
.C(n_525),
.Y(n_1100)
);

CKINVDCx5p33_ASAP7_75t_R g1101 ( 
.A(n_993),
.Y(n_1101)
);

AOI21xp5_ASAP7_75t_L g1102 ( 
.A1(n_991),
.A2(n_1009),
.B(n_970),
.Y(n_1102)
);

AOI21xp5_ASAP7_75t_L g1103 ( 
.A1(n_970),
.A2(n_637),
.B(n_636),
.Y(n_1103)
);

BUFx6f_ASAP7_75t_L g1104 ( 
.A(n_1092),
.Y(n_1104)
);

BUFx2_ASAP7_75t_SL g1105 ( 
.A(n_1060),
.Y(n_1105)
);

OAI21x1_ASAP7_75t_L g1106 ( 
.A1(n_1023),
.A2(n_1008),
.B(n_1017),
.Y(n_1106)
);

INVx2_ASAP7_75t_L g1107 ( 
.A(n_1024),
.Y(n_1107)
);

HB1xp67_ASAP7_75t_L g1108 ( 
.A(n_1034),
.Y(n_1108)
);

INVx4_ASAP7_75t_L g1109 ( 
.A(n_1092),
.Y(n_1109)
);

OA21x2_ASAP7_75t_L g1110 ( 
.A1(n_1022),
.A2(n_987),
.B(n_985),
.Y(n_1110)
);

AO21x2_ASAP7_75t_L g1111 ( 
.A1(n_1078),
.A2(n_944),
.B(n_1006),
.Y(n_1111)
);

AND2x4_ASAP7_75t_L g1112 ( 
.A(n_1059),
.B(n_965),
.Y(n_1112)
);

AOI22x1_ASAP7_75t_L g1113 ( 
.A1(n_1033),
.A2(n_963),
.B1(n_962),
.B2(n_984),
.Y(n_1113)
);

CKINVDCx5p33_ASAP7_75t_R g1114 ( 
.A(n_1071),
.Y(n_1114)
);

NOR2xp33_ASAP7_75t_L g1115 ( 
.A(n_1038),
.B(n_959),
.Y(n_1115)
);

INVx1_ASAP7_75t_L g1116 ( 
.A(n_1073),
.Y(n_1116)
);

NAND2x1p5_ASAP7_75t_L g1117 ( 
.A(n_1068),
.B(n_981),
.Y(n_1117)
);

BUFx6f_ASAP7_75t_L g1118 ( 
.A(n_1068),
.Y(n_1118)
);

NAND2x1p5_ASAP7_75t_L g1119 ( 
.A(n_1080),
.B(n_1009),
.Y(n_1119)
);

INVx1_ASAP7_75t_L g1120 ( 
.A(n_1072),
.Y(n_1120)
);

BUFx2_ASAP7_75t_L g1121 ( 
.A(n_1042),
.Y(n_1121)
);

INVx1_ASAP7_75t_L g1122 ( 
.A(n_1027),
.Y(n_1122)
);

OA21x2_ASAP7_75t_L g1123 ( 
.A1(n_1032),
.A2(n_1016),
.B(n_572),
.Y(n_1123)
);

AND2x2_ASAP7_75t_L g1124 ( 
.A(n_1027),
.B(n_943),
.Y(n_1124)
);

AO21x2_ASAP7_75t_L g1125 ( 
.A1(n_1044),
.A2(n_990),
.B(n_958),
.Y(n_1125)
);

HB1xp67_ASAP7_75t_L g1126 ( 
.A(n_1087),
.Y(n_1126)
);

INVx1_ASAP7_75t_SL g1127 ( 
.A(n_1057),
.Y(n_1127)
);

AND2x4_ASAP7_75t_L g1128 ( 
.A(n_1045),
.B(n_984),
.Y(n_1128)
);

BUFx10_ASAP7_75t_L g1129 ( 
.A(n_1093),
.Y(n_1129)
);

OAI21xp5_ASAP7_75t_L g1130 ( 
.A1(n_1037),
.A2(n_1004),
.B(n_994),
.Y(n_1130)
);

INVx2_ASAP7_75t_L g1131 ( 
.A(n_1084),
.Y(n_1131)
);

OAI21x1_ASAP7_75t_L g1132 ( 
.A1(n_1041),
.A2(n_572),
.B(n_564),
.Y(n_1132)
);

BUFx6f_ASAP7_75t_L g1133 ( 
.A(n_1035),
.Y(n_1133)
);

AND2x4_ASAP7_75t_L g1134 ( 
.A(n_1049),
.B(n_961),
.Y(n_1134)
);

OAI21x1_ASAP7_75t_L g1135 ( 
.A1(n_1102),
.A2(n_577),
.B(n_564),
.Y(n_1135)
);

INVx1_ASAP7_75t_L g1136 ( 
.A(n_1052),
.Y(n_1136)
);

AO21x2_ASAP7_75t_L g1137 ( 
.A1(n_1031),
.A2(n_599),
.B(n_577),
.Y(n_1137)
);

INVx4_ASAP7_75t_L g1138 ( 
.A(n_1097),
.Y(n_1138)
);

HB1xp67_ASAP7_75t_L g1139 ( 
.A(n_1035),
.Y(n_1139)
);

BUFx10_ASAP7_75t_L g1140 ( 
.A(n_1062),
.Y(n_1140)
);

INVx1_ASAP7_75t_L g1141 ( 
.A(n_1067),
.Y(n_1141)
);

INVx3_ASAP7_75t_L g1142 ( 
.A(n_1039),
.Y(n_1142)
);

AO21x2_ASAP7_75t_L g1143 ( 
.A1(n_1036),
.A2(n_599),
.B(n_946),
.Y(n_1143)
);

INVx1_ASAP7_75t_L g1144 ( 
.A(n_1094),
.Y(n_1144)
);

AND2x4_ASAP7_75t_L g1145 ( 
.A(n_1095),
.B(n_1009),
.Y(n_1145)
);

INVx4_ASAP7_75t_L g1146 ( 
.A(n_1042),
.Y(n_1146)
);

INVx1_ASAP7_75t_L g1147 ( 
.A(n_1069),
.Y(n_1147)
);

AND2x2_ASAP7_75t_L g1148 ( 
.A(n_1043),
.B(n_711),
.Y(n_1148)
);

INVx2_ASAP7_75t_L g1149 ( 
.A(n_1081),
.Y(n_1149)
);

NOR2xp67_ASAP7_75t_L g1150 ( 
.A(n_1066),
.B(n_76),
.Y(n_1150)
);

INVx8_ASAP7_75t_L g1151 ( 
.A(n_1042),
.Y(n_1151)
);

INVx3_ASAP7_75t_SL g1152 ( 
.A(n_1101),
.Y(n_1152)
);

AOI22xp33_ASAP7_75t_L g1153 ( 
.A1(n_1051),
.A2(n_1061),
.B1(n_1086),
.B2(n_1025),
.Y(n_1153)
);

OAI21x1_ASAP7_75t_L g1154 ( 
.A1(n_1053),
.A2(n_86),
.B(n_83),
.Y(n_1154)
);

INVx1_ASAP7_75t_L g1155 ( 
.A(n_1070),
.Y(n_1155)
);

BUFx2_ASAP7_75t_R g1156 ( 
.A(n_1098),
.Y(n_1156)
);

INVx3_ASAP7_75t_SL g1157 ( 
.A(n_1064),
.Y(n_1157)
);

AOI22xp33_ASAP7_75t_L g1158 ( 
.A1(n_1061),
.A2(n_711),
.B1(n_532),
.B2(n_544),
.Y(n_1158)
);

BUFx6f_ASAP7_75t_L g1159 ( 
.A(n_1047),
.Y(n_1159)
);

NAND2xp5_ASAP7_75t_SL g1160 ( 
.A(n_1065),
.B(n_550),
.Y(n_1160)
);

INVx5_ASAP7_75t_L g1161 ( 
.A(n_1028),
.Y(n_1161)
);

OAI21x1_ASAP7_75t_L g1162 ( 
.A1(n_1030),
.A2(n_90),
.B(n_87),
.Y(n_1162)
);

INVx1_ASAP7_75t_SL g1163 ( 
.A(n_1091),
.Y(n_1163)
);

INVx2_ASAP7_75t_L g1164 ( 
.A(n_1096),
.Y(n_1164)
);

OAI21x1_ASAP7_75t_L g1165 ( 
.A1(n_1103),
.A2(n_237),
.B(n_331),
.Y(n_1165)
);

AND2x4_ASAP7_75t_L g1166 ( 
.A(n_1063),
.B(n_91),
.Y(n_1166)
);

AND2x2_ASAP7_75t_L g1167 ( 
.A(n_1029),
.B(n_711),
.Y(n_1167)
);

INVx5_ASAP7_75t_SL g1168 ( 
.A(n_1075),
.Y(n_1168)
);

INVx2_ASAP7_75t_L g1169 ( 
.A(n_1055),
.Y(n_1169)
);

OR2x6_ASAP7_75t_L g1170 ( 
.A(n_1048),
.B(n_993),
.Y(n_1170)
);

INVx2_ASAP7_75t_L g1171 ( 
.A(n_1046),
.Y(n_1171)
);

INVx1_ASAP7_75t_L g1172 ( 
.A(n_1074),
.Y(n_1172)
);

AO21x2_ASAP7_75t_L g1173 ( 
.A1(n_1143),
.A2(n_1026),
.B(n_1079),
.Y(n_1173)
);

NAND2x1p5_ASAP7_75t_L g1174 ( 
.A(n_1104),
.B(n_1058),
.Y(n_1174)
);

AOI22xp5_ASAP7_75t_L g1175 ( 
.A1(n_1115),
.A2(n_1040),
.B1(n_1088),
.B2(n_1089),
.Y(n_1175)
);

INVx1_ASAP7_75t_L g1176 ( 
.A(n_1116),
.Y(n_1176)
);

INVx8_ASAP7_75t_L g1177 ( 
.A(n_1151),
.Y(n_1177)
);

INVx2_ASAP7_75t_L g1178 ( 
.A(n_1107),
.Y(n_1178)
);

INVx1_ASAP7_75t_L g1179 ( 
.A(n_1120),
.Y(n_1179)
);

INVx2_ASAP7_75t_L g1180 ( 
.A(n_1131),
.Y(n_1180)
);

NAND2xp5_ASAP7_75t_L g1181 ( 
.A(n_1169),
.B(n_1076),
.Y(n_1181)
);

NAND2xp5_ASAP7_75t_L g1182 ( 
.A(n_1171),
.B(n_1099),
.Y(n_1182)
);

INVx2_ASAP7_75t_L g1183 ( 
.A(n_1136),
.Y(n_1183)
);

OAI21xp5_ASAP7_75t_L g1184 ( 
.A1(n_1172),
.A2(n_1085),
.B(n_1100),
.Y(n_1184)
);

INVx3_ASAP7_75t_L g1185 ( 
.A(n_1118),
.Y(n_1185)
);

BUFx6f_ASAP7_75t_L g1186 ( 
.A(n_1104),
.Y(n_1186)
);

AOI22xp33_ASAP7_75t_L g1187 ( 
.A1(n_1115),
.A2(n_1090),
.B1(n_1083),
.B2(n_551),
.Y(n_1187)
);

AO21x1_ASAP7_75t_SL g1188 ( 
.A1(n_1153),
.A2(n_47),
.B(n_48),
.Y(n_1188)
);

INVx1_ASAP7_75t_L g1189 ( 
.A(n_1141),
.Y(n_1189)
);

INVx2_ASAP7_75t_SL g1190 ( 
.A(n_1159),
.Y(n_1190)
);

INVx1_ASAP7_75t_L g1191 ( 
.A(n_1122),
.Y(n_1191)
);

AOI22xp33_ASAP7_75t_L g1192 ( 
.A1(n_1153),
.A2(n_1082),
.B1(n_701),
.B2(n_1056),
.Y(n_1192)
);

NAND2xp5_ASAP7_75t_L g1193 ( 
.A(n_1144),
.B(n_1050),
.Y(n_1193)
);

INVx1_ASAP7_75t_L g1194 ( 
.A(n_1112),
.Y(n_1194)
);

INVx2_ASAP7_75t_L g1195 ( 
.A(n_1112),
.Y(n_1195)
);

INVx1_ASAP7_75t_L g1196 ( 
.A(n_1147),
.Y(n_1196)
);

INVx1_ASAP7_75t_L g1197 ( 
.A(n_1128),
.Y(n_1197)
);

HB1xp67_ASAP7_75t_L g1198 ( 
.A(n_1108),
.Y(n_1198)
);

HB1xp67_ASAP7_75t_L g1199 ( 
.A(n_1126),
.Y(n_1199)
);

AO21x1_ASAP7_75t_L g1200 ( 
.A1(n_1160),
.A2(n_1077),
.B(n_1054),
.Y(n_1200)
);

BUFx6f_ASAP7_75t_L g1201 ( 
.A(n_1104),
.Y(n_1201)
);

AOI22xp33_ASAP7_75t_L g1202 ( 
.A1(n_1124),
.A2(n_1139),
.B1(n_1142),
.B2(n_1158),
.Y(n_1202)
);

OAI21xp33_ASAP7_75t_L g1203 ( 
.A1(n_1158),
.A2(n_645),
.B(n_643),
.Y(n_1203)
);

NAND2x1p5_ASAP7_75t_L g1204 ( 
.A(n_1109),
.B(n_637),
.Y(n_1204)
);

AO21x2_ASAP7_75t_L g1205 ( 
.A1(n_1143),
.A2(n_701),
.B(n_92),
.Y(n_1205)
);

OAI22xp33_ASAP7_75t_L g1206 ( 
.A1(n_1157),
.A2(n_645),
.B1(n_643),
.B2(n_642),
.Y(n_1206)
);

INVx6_ASAP7_75t_L g1207 ( 
.A(n_1138),
.Y(n_1207)
);

BUFx3_ASAP7_75t_L g1208 ( 
.A(n_1159),
.Y(n_1208)
);

NAND2xp5_ASAP7_75t_L g1209 ( 
.A(n_1164),
.B(n_49),
.Y(n_1209)
);

CKINVDCx5p33_ASAP7_75t_R g1210 ( 
.A(n_1114),
.Y(n_1210)
);

AO21x1_ASAP7_75t_L g1211 ( 
.A1(n_1160),
.A2(n_49),
.B(n_94),
.Y(n_1211)
);

INVx6_ASAP7_75t_L g1212 ( 
.A(n_1138),
.Y(n_1212)
);

NAND2x1p5_ASAP7_75t_L g1213 ( 
.A(n_1109),
.B(n_637),
.Y(n_1213)
);

OAI21x1_ASAP7_75t_L g1214 ( 
.A1(n_1106),
.A2(n_95),
.B(n_99),
.Y(n_1214)
);

OAI21x1_ASAP7_75t_L g1215 ( 
.A1(n_1113),
.A2(n_100),
.B(n_102),
.Y(n_1215)
);

INVx1_ASAP7_75t_L g1216 ( 
.A(n_1142),
.Y(n_1216)
);

OAI21xp5_ASAP7_75t_L g1217 ( 
.A1(n_1130),
.A2(n_106),
.B(n_108),
.Y(n_1217)
);

INVx1_ASAP7_75t_L g1218 ( 
.A(n_1119),
.Y(n_1218)
);

INVx1_ASAP7_75t_L g1219 ( 
.A(n_1126),
.Y(n_1219)
);

OR2x6_ASAP7_75t_L g1220 ( 
.A(n_1151),
.B(n_642),
.Y(n_1220)
);

AND2x2_ASAP7_75t_L g1221 ( 
.A(n_1157),
.B(n_643),
.Y(n_1221)
);

INVx1_ASAP7_75t_L g1222 ( 
.A(n_1117),
.Y(n_1222)
);

CKINVDCx20_ASAP7_75t_R g1223 ( 
.A(n_1152),
.Y(n_1223)
);

HB1xp67_ASAP7_75t_L g1224 ( 
.A(n_1127),
.Y(n_1224)
);

AND2x2_ASAP7_75t_L g1225 ( 
.A(n_1167),
.B(n_645),
.Y(n_1225)
);

INVx1_ASAP7_75t_L g1226 ( 
.A(n_1117),
.Y(n_1226)
);

OAI21x1_ASAP7_75t_L g1227 ( 
.A1(n_1132),
.A2(n_112),
.B(n_113),
.Y(n_1227)
);

INVx1_ASAP7_75t_L g1228 ( 
.A(n_1145),
.Y(n_1228)
);

INVx2_ASAP7_75t_L g1229 ( 
.A(n_1135),
.Y(n_1229)
);

NAND2xp33_ASAP7_75t_R g1230 ( 
.A(n_1210),
.B(n_1121),
.Y(n_1230)
);

AND2x2_ASAP7_75t_L g1231 ( 
.A(n_1195),
.B(n_1194),
.Y(n_1231)
);

HB1xp67_ASAP7_75t_L g1232 ( 
.A(n_1224),
.Y(n_1232)
);

BUFx3_ASAP7_75t_L g1233 ( 
.A(n_1208),
.Y(n_1233)
);

OA21x2_ASAP7_75t_L g1234 ( 
.A1(n_1215),
.A2(n_1162),
.B(n_1154),
.Y(n_1234)
);

CKINVDCx5p33_ASAP7_75t_R g1235 ( 
.A(n_1223),
.Y(n_1235)
);

INVx1_ASAP7_75t_L g1236 ( 
.A(n_1176),
.Y(n_1236)
);

AO32x2_ASAP7_75t_L g1237 ( 
.A1(n_1188),
.A2(n_1146),
.A3(n_1125),
.B1(n_1170),
.B2(n_1137),
.Y(n_1237)
);

A2O1A1Ixp33_ASAP7_75t_L g1238 ( 
.A1(n_1175),
.A2(n_1150),
.B(n_1155),
.C(n_1163),
.Y(n_1238)
);

CKINVDCx5p33_ASAP7_75t_R g1239 ( 
.A(n_1224),
.Y(n_1239)
);

NAND2xp33_ASAP7_75t_R g1240 ( 
.A(n_1221),
.B(n_1166),
.Y(n_1240)
);

HB1xp67_ASAP7_75t_L g1241 ( 
.A(n_1199),
.Y(n_1241)
);

INVx4_ASAP7_75t_L g1242 ( 
.A(n_1186),
.Y(n_1242)
);

NAND2xp5_ASAP7_75t_L g1243 ( 
.A(n_1196),
.B(n_1148),
.Y(n_1243)
);

INVx1_ASAP7_75t_L g1244 ( 
.A(n_1189),
.Y(n_1244)
);

INVx2_ASAP7_75t_L g1245 ( 
.A(n_1178),
.Y(n_1245)
);

INVx1_ASAP7_75t_L g1246 ( 
.A(n_1183),
.Y(n_1246)
);

BUFx3_ASAP7_75t_L g1247 ( 
.A(n_1207),
.Y(n_1247)
);

HB1xp67_ASAP7_75t_L g1248 ( 
.A(n_1198),
.Y(n_1248)
);

NAND2xp5_ASAP7_75t_L g1249 ( 
.A(n_1181),
.B(n_1150),
.Y(n_1249)
);

INVx1_ASAP7_75t_L g1250 ( 
.A(n_1179),
.Y(n_1250)
);

NAND2xp33_ASAP7_75t_R g1251 ( 
.A(n_1228),
.B(n_1166),
.Y(n_1251)
);

AND2x2_ASAP7_75t_L g1252 ( 
.A(n_1225),
.B(n_1133),
.Y(n_1252)
);

AOI22xp33_ASAP7_75t_L g1253 ( 
.A1(n_1217),
.A2(n_1134),
.B1(n_1140),
.B2(n_1161),
.Y(n_1253)
);

NAND2xp33_ASAP7_75t_R g1254 ( 
.A(n_1182),
.B(n_1134),
.Y(n_1254)
);

INVx2_ASAP7_75t_SL g1255 ( 
.A(n_1212),
.Y(n_1255)
);

CKINVDCx5p33_ASAP7_75t_R g1256 ( 
.A(n_1212),
.Y(n_1256)
);

AOI22xp33_ASAP7_75t_L g1257 ( 
.A1(n_1217),
.A2(n_1140),
.B1(n_1161),
.B2(n_1146),
.Y(n_1257)
);

CKINVDCx5p33_ASAP7_75t_R g1258 ( 
.A(n_1190),
.Y(n_1258)
);

INVx1_ASAP7_75t_L g1259 ( 
.A(n_1191),
.Y(n_1259)
);

NAND2xp5_ASAP7_75t_L g1260 ( 
.A(n_1181),
.B(n_1161),
.Y(n_1260)
);

BUFx3_ASAP7_75t_L g1261 ( 
.A(n_1219),
.Y(n_1261)
);

NAND2xp5_ASAP7_75t_L g1262 ( 
.A(n_1182),
.B(n_1161),
.Y(n_1262)
);

BUFx6f_ASAP7_75t_L g1263 ( 
.A(n_1186),
.Y(n_1263)
);

NAND2xp33_ASAP7_75t_SL g1264 ( 
.A(n_1186),
.B(n_1105),
.Y(n_1264)
);

AND2x2_ASAP7_75t_L g1265 ( 
.A(n_1202),
.B(n_1129),
.Y(n_1265)
);

BUFx3_ASAP7_75t_L g1266 ( 
.A(n_1177),
.Y(n_1266)
);

NOR3xp33_ASAP7_75t_SL g1267 ( 
.A(n_1206),
.B(n_1170),
.C(n_1156),
.Y(n_1267)
);

NOR2x1p5_ASAP7_75t_L g1268 ( 
.A(n_1209),
.B(n_1156),
.Y(n_1268)
);

CKINVDCx20_ASAP7_75t_R g1269 ( 
.A(n_1177),
.Y(n_1269)
);

NAND2xp33_ASAP7_75t_R g1270 ( 
.A(n_1197),
.B(n_1170),
.Y(n_1270)
);

INVx2_ASAP7_75t_L g1271 ( 
.A(n_1180),
.Y(n_1271)
);

CKINVDCx5p33_ASAP7_75t_R g1272 ( 
.A(n_1177),
.Y(n_1272)
);

OAI22xp5_ASAP7_75t_L g1273 ( 
.A1(n_1203),
.A2(n_1149),
.B1(n_1123),
.B2(n_1110),
.Y(n_1273)
);

OAI222xp33_ASAP7_75t_L g1274 ( 
.A1(n_1175),
.A2(n_1125),
.B1(n_1137),
.B2(n_1111),
.C1(n_1168),
.C2(n_1165),
.Y(n_1274)
);

HB1xp67_ASAP7_75t_L g1275 ( 
.A(n_1173),
.Y(n_1275)
);

CKINVDCx5p33_ASAP7_75t_R g1276 ( 
.A(n_1201),
.Y(n_1276)
);

AOI22xp33_ASAP7_75t_L g1277 ( 
.A1(n_1187),
.A2(n_1111),
.B1(n_1123),
.B2(n_1110),
.Y(n_1277)
);

OR2x2_ASAP7_75t_SL g1278 ( 
.A(n_1209),
.B(n_1168),
.Y(n_1278)
);

CKINVDCx20_ASAP7_75t_R g1279 ( 
.A(n_1201),
.Y(n_1279)
);

INVx1_ASAP7_75t_L g1280 ( 
.A(n_1216),
.Y(n_1280)
);

AND2x4_ASAP7_75t_L g1281 ( 
.A(n_1185),
.B(n_125),
.Y(n_1281)
);

NAND2xp33_ASAP7_75t_SL g1282 ( 
.A(n_1201),
.B(n_128),
.Y(n_1282)
);

NAND2xp5_ASAP7_75t_L g1283 ( 
.A(n_1203),
.B(n_330),
.Y(n_1283)
);

BUFx12f_ASAP7_75t_L g1284 ( 
.A(n_1220),
.Y(n_1284)
);

INVx1_ASAP7_75t_L g1285 ( 
.A(n_1236),
.Y(n_1285)
);

INVx1_ASAP7_75t_L g1286 ( 
.A(n_1244),
.Y(n_1286)
);

INVx2_ASAP7_75t_L g1287 ( 
.A(n_1250),
.Y(n_1287)
);

AOI22xp33_ASAP7_75t_L g1288 ( 
.A1(n_1253),
.A2(n_1265),
.B1(n_1257),
.B2(n_1268),
.Y(n_1288)
);

INVx2_ASAP7_75t_SL g1289 ( 
.A(n_1232),
.Y(n_1289)
);

AND2x4_ASAP7_75t_L g1290 ( 
.A(n_1259),
.B(n_1280),
.Y(n_1290)
);

BUFx2_ASAP7_75t_L g1291 ( 
.A(n_1239),
.Y(n_1291)
);

OR2x2_ASAP7_75t_L g1292 ( 
.A(n_1241),
.B(n_1173),
.Y(n_1292)
);

NAND2xp5_ASAP7_75t_L g1293 ( 
.A(n_1249),
.B(n_1260),
.Y(n_1293)
);

NAND2xp5_ASAP7_75t_L g1294 ( 
.A(n_1249),
.B(n_1174),
.Y(n_1294)
);

INVx2_ASAP7_75t_L g1295 ( 
.A(n_1246),
.Y(n_1295)
);

BUFx6f_ASAP7_75t_L g1296 ( 
.A(n_1263),
.Y(n_1296)
);

AND2x2_ASAP7_75t_L g1297 ( 
.A(n_1231),
.B(n_1222),
.Y(n_1297)
);

INVxp67_ASAP7_75t_L g1298 ( 
.A(n_1248),
.Y(n_1298)
);

INVxp67_ASAP7_75t_SL g1299 ( 
.A(n_1275),
.Y(n_1299)
);

AND2x4_ASAP7_75t_L g1300 ( 
.A(n_1281),
.B(n_1226),
.Y(n_1300)
);

INVx2_ASAP7_75t_L g1301 ( 
.A(n_1275),
.Y(n_1301)
);

INVx2_ASAP7_75t_L g1302 ( 
.A(n_1245),
.Y(n_1302)
);

NAND2xp5_ASAP7_75t_L g1303 ( 
.A(n_1243),
.B(n_1193),
.Y(n_1303)
);

OAI22xp5_ASAP7_75t_L g1304 ( 
.A1(n_1267),
.A2(n_1220),
.B1(n_1218),
.B2(n_1192),
.Y(n_1304)
);

NAND3xp33_ASAP7_75t_L g1305 ( 
.A(n_1238),
.B(n_1184),
.C(n_1220),
.Y(n_1305)
);

AND2x2_ASAP7_75t_L g1306 ( 
.A(n_1252),
.B(n_1184),
.Y(n_1306)
);

INVx2_ASAP7_75t_L g1307 ( 
.A(n_1271),
.Y(n_1307)
);

AND2x2_ASAP7_75t_L g1308 ( 
.A(n_1261),
.B(n_1211),
.Y(n_1308)
);

INVx3_ASAP7_75t_L g1309 ( 
.A(n_1263),
.Y(n_1309)
);

INVx2_ASAP7_75t_L g1310 ( 
.A(n_1262),
.Y(n_1310)
);

AND2x4_ASAP7_75t_L g1311 ( 
.A(n_1281),
.B(n_1214),
.Y(n_1311)
);

BUFx3_ASAP7_75t_L g1312 ( 
.A(n_1247),
.Y(n_1312)
);

OR2x2_ASAP7_75t_L g1313 ( 
.A(n_1262),
.B(n_1205),
.Y(n_1313)
);

INVx1_ASAP7_75t_L g1314 ( 
.A(n_1243),
.Y(n_1314)
);

INVx2_ASAP7_75t_SL g1315 ( 
.A(n_1263),
.Y(n_1315)
);

INVx2_ASAP7_75t_SL g1316 ( 
.A(n_1266),
.Y(n_1316)
);

AND2x2_ASAP7_75t_L g1317 ( 
.A(n_1242),
.B(n_1205),
.Y(n_1317)
);

INVx2_ASAP7_75t_L g1318 ( 
.A(n_1234),
.Y(n_1318)
);

CKINVDCx6p67_ASAP7_75t_R g1319 ( 
.A(n_1279),
.Y(n_1319)
);

INVx2_ASAP7_75t_SL g1320 ( 
.A(n_1276),
.Y(n_1320)
);

INVx1_ASAP7_75t_L g1321 ( 
.A(n_1237),
.Y(n_1321)
);

AO21x2_ASAP7_75t_L g1322 ( 
.A1(n_1274),
.A2(n_1229),
.B(n_1200),
.Y(n_1322)
);

INVx1_ASAP7_75t_L g1323 ( 
.A(n_1237),
.Y(n_1323)
);

AND2x2_ASAP7_75t_L g1324 ( 
.A(n_1242),
.B(n_1204),
.Y(n_1324)
);

INVx1_ASAP7_75t_L g1325 ( 
.A(n_1237),
.Y(n_1325)
);

INVx2_ASAP7_75t_L g1326 ( 
.A(n_1234),
.Y(n_1326)
);

OAI21x1_ASAP7_75t_L g1327 ( 
.A1(n_1273),
.A2(n_1227),
.B(n_1213),
.Y(n_1327)
);

INVx1_ASAP7_75t_L g1328 ( 
.A(n_1283),
.Y(n_1328)
);

NAND2x1p5_ASAP7_75t_L g1329 ( 
.A(n_1255),
.B(n_1204),
.Y(n_1329)
);

CKINVDCx5p33_ASAP7_75t_R g1330 ( 
.A(n_1230),
.Y(n_1330)
);

INVx2_ASAP7_75t_SL g1331 ( 
.A(n_1233),
.Y(n_1331)
);

OR2x2_ASAP7_75t_L g1332 ( 
.A(n_1278),
.B(n_1213),
.Y(n_1332)
);

NAND2xp5_ASAP7_75t_L g1333 ( 
.A(n_1235),
.B(n_130),
.Y(n_1333)
);

AND2x4_ASAP7_75t_L g1334 ( 
.A(n_1269),
.B(n_1272),
.Y(n_1334)
);

INVx1_ASAP7_75t_L g1335 ( 
.A(n_1273),
.Y(n_1335)
);

INVx2_ASAP7_75t_L g1336 ( 
.A(n_1258),
.Y(n_1336)
);

INVx2_ASAP7_75t_L g1337 ( 
.A(n_1284),
.Y(n_1337)
);

INVx1_ASAP7_75t_L g1338 ( 
.A(n_1287),
.Y(n_1338)
);

INVx2_ASAP7_75t_L g1339 ( 
.A(n_1287),
.Y(n_1339)
);

AND2x4_ASAP7_75t_L g1340 ( 
.A(n_1290),
.B(n_1277),
.Y(n_1340)
);

INVx1_ASAP7_75t_L g1341 ( 
.A(n_1285),
.Y(n_1341)
);

OAI221xp5_ASAP7_75t_L g1342 ( 
.A1(n_1288),
.A2(n_1240),
.B1(n_1251),
.B2(n_1305),
.C(n_1332),
.Y(n_1342)
);

INVx1_ASAP7_75t_L g1343 ( 
.A(n_1286),
.Y(n_1343)
);

NOR2xp33_ASAP7_75t_L g1344 ( 
.A(n_1294),
.B(n_1274),
.Y(n_1344)
);

INVx2_ASAP7_75t_SL g1345 ( 
.A(n_1290),
.Y(n_1345)
);

NAND2xp5_ASAP7_75t_L g1346 ( 
.A(n_1293),
.B(n_1256),
.Y(n_1346)
);

INVx2_ASAP7_75t_L g1347 ( 
.A(n_1310),
.Y(n_1347)
);

AND2x2_ASAP7_75t_L g1348 ( 
.A(n_1306),
.B(n_1254),
.Y(n_1348)
);

NAND2xp5_ASAP7_75t_L g1349 ( 
.A(n_1310),
.B(n_1264),
.Y(n_1349)
);

AND2x4_ASAP7_75t_L g1350 ( 
.A(n_1290),
.B(n_1270),
.Y(n_1350)
);

INVx1_ASAP7_75t_L g1351 ( 
.A(n_1295),
.Y(n_1351)
);

INVx2_ASAP7_75t_L g1352 ( 
.A(n_1318),
.Y(n_1352)
);

OR2x2_ASAP7_75t_L g1353 ( 
.A(n_1292),
.B(n_1282),
.Y(n_1353)
);

NAND2xp5_ASAP7_75t_L g1354 ( 
.A(n_1314),
.B(n_1303),
.Y(n_1354)
);

INVx1_ASAP7_75t_L g1355 ( 
.A(n_1295),
.Y(n_1355)
);

INVx2_ASAP7_75t_L g1356 ( 
.A(n_1318),
.Y(n_1356)
);

HB1xp67_ASAP7_75t_L g1357 ( 
.A(n_1301),
.Y(n_1357)
);

INVx2_ASAP7_75t_L g1358 ( 
.A(n_1326),
.Y(n_1358)
);

AND2x4_ASAP7_75t_L g1359 ( 
.A(n_1301),
.B(n_131),
.Y(n_1359)
);

INVx2_ASAP7_75t_L g1360 ( 
.A(n_1326),
.Y(n_1360)
);

INVx1_ASAP7_75t_L g1361 ( 
.A(n_1298),
.Y(n_1361)
);

INVx1_ASAP7_75t_L g1362 ( 
.A(n_1289),
.Y(n_1362)
);

INVx1_ASAP7_75t_L g1363 ( 
.A(n_1299),
.Y(n_1363)
);

HB1xp67_ASAP7_75t_L g1364 ( 
.A(n_1299),
.Y(n_1364)
);

NOR2xp33_ASAP7_75t_SL g1365 ( 
.A(n_1330),
.B(n_148),
.Y(n_1365)
);

NOR3xp33_ASAP7_75t_L g1366 ( 
.A(n_1304),
.B(n_149),
.C(n_150),
.Y(n_1366)
);

INVx2_ASAP7_75t_L g1367 ( 
.A(n_1302),
.Y(n_1367)
);

NAND2xp5_ASAP7_75t_L g1368 ( 
.A(n_1328),
.B(n_159),
.Y(n_1368)
);

HB1xp67_ASAP7_75t_L g1369 ( 
.A(n_1335),
.Y(n_1369)
);

AND2x2_ASAP7_75t_L g1370 ( 
.A(n_1321),
.B(n_160),
.Y(n_1370)
);

NAND2xp5_ASAP7_75t_SL g1371 ( 
.A(n_1288),
.B(n_164),
.Y(n_1371)
);

INVx2_ASAP7_75t_L g1372 ( 
.A(n_1307),
.Y(n_1372)
);

OR2x2_ASAP7_75t_L g1373 ( 
.A(n_1313),
.B(n_165),
.Y(n_1373)
);

OAI22xp5_ASAP7_75t_L g1374 ( 
.A1(n_1330),
.A2(n_169),
.B1(n_170),
.B2(n_171),
.Y(n_1374)
);

INVx1_ASAP7_75t_L g1375 ( 
.A(n_1323),
.Y(n_1375)
);

BUFx2_ASAP7_75t_L g1376 ( 
.A(n_1350),
.Y(n_1376)
);

NAND2xp5_ASAP7_75t_L g1377 ( 
.A(n_1354),
.B(n_1308),
.Y(n_1377)
);

AND2x2_ASAP7_75t_L g1378 ( 
.A(n_1345),
.B(n_1325),
.Y(n_1378)
);

OR2x2_ASAP7_75t_L g1379 ( 
.A(n_1357),
.B(n_1322),
.Y(n_1379)
);

INVx1_ASAP7_75t_L g1380 ( 
.A(n_1341),
.Y(n_1380)
);

NAND2xp5_ASAP7_75t_L g1381 ( 
.A(n_1361),
.B(n_1297),
.Y(n_1381)
);

AND2x2_ASAP7_75t_L g1382 ( 
.A(n_1375),
.B(n_1317),
.Y(n_1382)
);

INVx1_ASAP7_75t_L g1383 ( 
.A(n_1343),
.Y(n_1383)
);

AND2x2_ASAP7_75t_L g1384 ( 
.A(n_1348),
.B(n_1327),
.Y(n_1384)
);

INVx2_ASAP7_75t_L g1385 ( 
.A(n_1352),
.Y(n_1385)
);

INVx4_ASAP7_75t_L g1386 ( 
.A(n_1359),
.Y(n_1386)
);

INVx2_ASAP7_75t_L g1387 ( 
.A(n_1352),
.Y(n_1387)
);

OR2x2_ASAP7_75t_L g1388 ( 
.A(n_1364),
.B(n_1291),
.Y(n_1388)
);

HB1xp67_ASAP7_75t_L g1389 ( 
.A(n_1369),
.Y(n_1389)
);

HB1xp67_ASAP7_75t_L g1390 ( 
.A(n_1369),
.Y(n_1390)
);

HB1xp67_ASAP7_75t_L g1391 ( 
.A(n_1363),
.Y(n_1391)
);

HB1xp67_ASAP7_75t_L g1392 ( 
.A(n_1362),
.Y(n_1392)
);

NOR2xp33_ASAP7_75t_L g1393 ( 
.A(n_1342),
.B(n_1331),
.Y(n_1393)
);

HB1xp67_ASAP7_75t_L g1394 ( 
.A(n_1347),
.Y(n_1394)
);

INVx1_ASAP7_75t_L g1395 ( 
.A(n_1339),
.Y(n_1395)
);

INVx3_ASAP7_75t_L g1396 ( 
.A(n_1356),
.Y(n_1396)
);

INVx1_ASAP7_75t_L g1397 ( 
.A(n_1338),
.Y(n_1397)
);

AND2x2_ASAP7_75t_L g1398 ( 
.A(n_1340),
.B(n_1337),
.Y(n_1398)
);

NOR2xp33_ASAP7_75t_R g1399 ( 
.A(n_1365),
.B(n_1319),
.Y(n_1399)
);

INVx2_ASAP7_75t_L g1400 ( 
.A(n_1356),
.Y(n_1400)
);

AOI22xp5_ASAP7_75t_L g1401 ( 
.A1(n_1393),
.A2(n_1371),
.B1(n_1366),
.B2(n_1344),
.Y(n_1401)
);

NOR2xp33_ASAP7_75t_L g1402 ( 
.A(n_1393),
.B(n_1346),
.Y(n_1402)
);

INVx2_ASAP7_75t_SL g1403 ( 
.A(n_1388),
.Y(n_1403)
);

HB1xp67_ASAP7_75t_L g1404 ( 
.A(n_1389),
.Y(n_1404)
);

OAI22xp33_ASAP7_75t_L g1405 ( 
.A1(n_1386),
.A2(n_1371),
.B1(n_1353),
.B2(n_1344),
.Y(n_1405)
);

OAI22xp33_ASAP7_75t_L g1406 ( 
.A1(n_1386),
.A2(n_1349),
.B1(n_1373),
.B2(n_1350),
.Y(n_1406)
);

OR2x2_ASAP7_75t_L g1407 ( 
.A(n_1384),
.B(n_1358),
.Y(n_1407)
);

OAI32xp33_ASAP7_75t_L g1408 ( 
.A1(n_1377),
.A2(n_1379),
.A3(n_1390),
.B1(n_1381),
.B2(n_1392),
.Y(n_1408)
);

AND2x4_ASAP7_75t_L g1409 ( 
.A(n_1376),
.B(n_1340),
.Y(n_1409)
);

NAND2xp5_ASAP7_75t_L g1410 ( 
.A(n_1398),
.B(n_1351),
.Y(n_1410)
);

INVx2_ASAP7_75t_L g1411 ( 
.A(n_1396),
.Y(n_1411)
);

INVx1_ASAP7_75t_L g1412 ( 
.A(n_1380),
.Y(n_1412)
);

AND2x4_ASAP7_75t_L g1413 ( 
.A(n_1398),
.B(n_1340),
.Y(n_1413)
);

INVx1_ASAP7_75t_L g1414 ( 
.A(n_1383),
.Y(n_1414)
);

OAI22xp33_ASAP7_75t_L g1415 ( 
.A1(n_1386),
.A2(n_1368),
.B1(n_1319),
.B2(n_1374),
.Y(n_1415)
);

INVx1_ASAP7_75t_L g1416 ( 
.A(n_1391),
.Y(n_1416)
);

INVxp67_ASAP7_75t_SL g1417 ( 
.A(n_1394),
.Y(n_1417)
);

AOI22xp5_ASAP7_75t_L g1418 ( 
.A1(n_1401),
.A2(n_1405),
.B1(n_1402),
.B2(n_1415),
.Y(n_1418)
);

INVx1_ASAP7_75t_L g1419 ( 
.A(n_1412),
.Y(n_1419)
);

INVx1_ASAP7_75t_L g1420 ( 
.A(n_1414),
.Y(n_1420)
);

INVxp67_ASAP7_75t_SL g1421 ( 
.A(n_1404),
.Y(n_1421)
);

INVx2_ASAP7_75t_L g1422 ( 
.A(n_1411),
.Y(n_1422)
);

INVx1_ASAP7_75t_L g1423 ( 
.A(n_1416),
.Y(n_1423)
);

XNOR2xp5_ASAP7_75t_L g1424 ( 
.A(n_1406),
.B(n_1334),
.Y(n_1424)
);

OAI22xp33_ASAP7_75t_L g1425 ( 
.A1(n_1403),
.A2(n_1397),
.B1(n_1359),
.B2(n_1370),
.Y(n_1425)
);

AOI22xp5_ASAP7_75t_L g1426 ( 
.A1(n_1409),
.A2(n_1413),
.B1(n_1410),
.B2(n_1300),
.Y(n_1426)
);

AOI21xp33_ASAP7_75t_L g1427 ( 
.A1(n_1408),
.A2(n_1417),
.B(n_1333),
.Y(n_1427)
);

OAI22xp33_ASAP7_75t_L g1428 ( 
.A1(n_1407),
.A2(n_1370),
.B1(n_1355),
.B2(n_1395),
.Y(n_1428)
);

OAI21xp33_ASAP7_75t_L g1429 ( 
.A1(n_1418),
.A2(n_1382),
.B(n_1399),
.Y(n_1429)
);

INVx1_ASAP7_75t_L g1430 ( 
.A(n_1419),
.Y(n_1430)
);

AO32x1_ASAP7_75t_L g1431 ( 
.A1(n_1424),
.A2(n_1320),
.A3(n_1316),
.B1(n_1336),
.B2(n_1315),
.Y(n_1431)
);

INVx1_ASAP7_75t_L g1432 ( 
.A(n_1420),
.Y(n_1432)
);

AOI21xp5_ASAP7_75t_L g1433 ( 
.A1(n_1427),
.A2(n_1334),
.B(n_1316),
.Y(n_1433)
);

NAND2x1_ASAP7_75t_SL g1434 ( 
.A(n_1426),
.B(n_1378),
.Y(n_1434)
);

AOI22xp5_ASAP7_75t_L g1435 ( 
.A1(n_1423),
.A2(n_1300),
.B1(n_1324),
.B2(n_1311),
.Y(n_1435)
);

NAND2xp5_ASAP7_75t_L g1436 ( 
.A(n_1421),
.B(n_1385),
.Y(n_1436)
);

INVx1_ASAP7_75t_L g1437 ( 
.A(n_1422),
.Y(n_1437)
);

NAND2xp5_ASAP7_75t_L g1438 ( 
.A(n_1428),
.B(n_1387),
.Y(n_1438)
);

OR2x2_ASAP7_75t_L g1439 ( 
.A(n_1425),
.B(n_1400),
.Y(n_1439)
);

INVxp67_ASAP7_75t_L g1440 ( 
.A(n_1421),
.Y(n_1440)
);

NAND2xp5_ASAP7_75t_L g1441 ( 
.A(n_1440),
.B(n_1312),
.Y(n_1441)
);

XOR2x2_ASAP7_75t_L g1442 ( 
.A(n_1433),
.B(n_1329),
.Y(n_1442)
);

NAND3xp33_ASAP7_75t_L g1443 ( 
.A(n_1429),
.B(n_1372),
.C(n_1367),
.Y(n_1443)
);

NOR2x1_ASAP7_75t_L g1444 ( 
.A(n_1430),
.B(n_1432),
.Y(n_1444)
);

INVx1_ASAP7_75t_L g1445 ( 
.A(n_1437),
.Y(n_1445)
);

INVxp67_ASAP7_75t_SL g1446 ( 
.A(n_1434),
.Y(n_1446)
);

AND2x2_ASAP7_75t_L g1447 ( 
.A(n_1446),
.B(n_1435),
.Y(n_1447)
);

NOR2x1_ASAP7_75t_L g1448 ( 
.A(n_1444),
.B(n_1439),
.Y(n_1448)
);

INVx1_ASAP7_75t_L g1449 ( 
.A(n_1445),
.Y(n_1449)
);

OAI22xp5_ASAP7_75t_SL g1450 ( 
.A1(n_1441),
.A2(n_1431),
.B1(n_1438),
.B2(n_1436),
.Y(n_1450)
);

AOI21xp5_ASAP7_75t_L g1451 ( 
.A1(n_1442),
.A2(n_1315),
.B(n_1367),
.Y(n_1451)
);

NOR3xp33_ASAP7_75t_L g1452 ( 
.A(n_1443),
.B(n_1309),
.C(n_1358),
.Y(n_1452)
);

OAI22xp5_ASAP7_75t_L g1453 ( 
.A1(n_1448),
.A2(n_1296),
.B1(n_1360),
.B2(n_180),
.Y(n_1453)
);

AOI21xp5_ASAP7_75t_L g1454 ( 
.A1(n_1450),
.A2(n_1360),
.B(n_1296),
.Y(n_1454)
);

NOR4xp25_ASAP7_75t_L g1455 ( 
.A(n_1449),
.B(n_172),
.C(n_173),
.D(n_181),
.Y(n_1455)
);

NAND3xp33_ASAP7_75t_L g1456 ( 
.A(n_1447),
.B(n_1296),
.C(n_189),
.Y(n_1456)
);

AOI221xp5_ASAP7_75t_L g1457 ( 
.A1(n_1452),
.A2(n_182),
.B1(n_190),
.B2(n_194),
.C(n_195),
.Y(n_1457)
);

INVx1_ASAP7_75t_SL g1458 ( 
.A(n_1451),
.Y(n_1458)
);

INVxp67_ASAP7_75t_SL g1459 ( 
.A(n_1453),
.Y(n_1459)
);

INVx1_ASAP7_75t_L g1460 ( 
.A(n_1458),
.Y(n_1460)
);

INVx2_ASAP7_75t_L g1461 ( 
.A(n_1456),
.Y(n_1461)
);

INVx1_ASAP7_75t_L g1462 ( 
.A(n_1454),
.Y(n_1462)
);

AOI22xp5_ASAP7_75t_L g1463 ( 
.A1(n_1455),
.A2(n_198),
.B1(n_201),
.B2(n_203),
.Y(n_1463)
);

AND2x4_ASAP7_75t_L g1464 ( 
.A(n_1457),
.B(n_210),
.Y(n_1464)
);

NAND4xp75_ASAP7_75t_L g1465 ( 
.A(n_1460),
.B(n_215),
.C(n_217),
.D(n_225),
.Y(n_1465)
);

AOI22xp5_ASAP7_75t_L g1466 ( 
.A1(n_1464),
.A2(n_228),
.B1(n_230),
.B2(n_234),
.Y(n_1466)
);

XOR2xp5_ASAP7_75t_L g1467 ( 
.A(n_1459),
.B(n_239),
.Y(n_1467)
);

NOR2xp33_ASAP7_75t_L g1468 ( 
.A(n_1461),
.B(n_241),
.Y(n_1468)
);

CKINVDCx5p33_ASAP7_75t_R g1469 ( 
.A(n_1467),
.Y(n_1469)
);

CKINVDCx5p33_ASAP7_75t_R g1470 ( 
.A(n_1468),
.Y(n_1470)
);

NAND2xp5_ASAP7_75t_SL g1471 ( 
.A(n_1466),
.B(n_1462),
.Y(n_1471)
);

OR2x2_ASAP7_75t_L g1472 ( 
.A(n_1465),
.B(n_1463),
.Y(n_1472)
);

INVx1_ASAP7_75t_L g1473 ( 
.A(n_1469),
.Y(n_1473)
);

XOR2x1_ASAP7_75t_L g1474 ( 
.A(n_1472),
.B(n_242),
.Y(n_1474)
);

XOR2xp5_ASAP7_75t_L g1475 ( 
.A(n_1471),
.B(n_245),
.Y(n_1475)
);

HB1xp67_ASAP7_75t_L g1476 ( 
.A(n_1469),
.Y(n_1476)
);

INVx2_ASAP7_75t_L g1477 ( 
.A(n_1470),
.Y(n_1477)
);

INVx1_ASAP7_75t_L g1478 ( 
.A(n_1476),
.Y(n_1478)
);

OR2x2_ASAP7_75t_L g1479 ( 
.A(n_1473),
.B(n_253),
.Y(n_1479)
);

NOR2xp33_ASAP7_75t_L g1480 ( 
.A(n_1474),
.B(n_260),
.Y(n_1480)
);

INVx1_ASAP7_75t_L g1481 ( 
.A(n_1475),
.Y(n_1481)
);

NOR2xp33_ASAP7_75t_L g1482 ( 
.A(n_1477),
.B(n_262),
.Y(n_1482)
);

INVx1_ASAP7_75t_L g1483 ( 
.A(n_1478),
.Y(n_1483)
);

OAI21xp5_ASAP7_75t_L g1484 ( 
.A1(n_1481),
.A2(n_1480),
.B(n_1482),
.Y(n_1484)
);

CKINVDCx20_ASAP7_75t_R g1485 ( 
.A(n_1479),
.Y(n_1485)
);

AOI22xp33_ASAP7_75t_R g1486 ( 
.A1(n_1483),
.A2(n_266),
.B1(n_270),
.B2(n_276),
.Y(n_1486)
);

OAI211xp5_ASAP7_75t_SL g1487 ( 
.A1(n_1484),
.A2(n_277),
.B(n_279),
.C(n_280),
.Y(n_1487)
);

OAI22xp5_ASAP7_75t_L g1488 ( 
.A1(n_1486),
.A2(n_1485),
.B1(n_1487),
.B2(n_291),
.Y(n_1488)
);

AOI22xp5_ASAP7_75t_SL g1489 ( 
.A1(n_1488),
.A2(n_292),
.B1(n_293),
.B2(n_294),
.Y(n_1489)
);

OR2x6_ASAP7_75t_L g1490 ( 
.A(n_1489),
.B(n_304),
.Y(n_1490)
);

OAI22xp33_ASAP7_75t_L g1491 ( 
.A1(n_1490),
.A2(n_307),
.B1(n_313),
.B2(n_318),
.Y(n_1491)
);


endmodule