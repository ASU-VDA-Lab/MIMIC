module real_aes_17269_n_101 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_101);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_101;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_830;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_838;
wire n_485;
wire n_822;
wire n_846;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_841;
wire n_318;
wire n_718;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_555;
wire n_421;
wire n_329;
wire n_852;
wire n_766;
wire n_132;
wire n_857;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_556;
wire n_545;
wire n_341;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_865;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_594;
wire n_856;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_564;
wire n_519;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_824;
wire n_467;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_559;
wire n_466;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_840;
wire n_570;
wire n_675;
wire n_530;
wire n_835;
wire n_104;
wire n_535;
wire n_732;
wire n_834;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_755;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_746;
wire n_178;
wire n_409;
wire n_781;
wire n_748;
wire n_860;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_455;
wire n_310;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_102;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_812;
wire n_817;
wire n_565;
wire n_443;
wire n_782;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_417;
wire n_363;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_617;
wire n_402;
wire n_552;
wire n_602;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_807;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_832;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_859;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_848;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_569;
wire n_303;
wire n_563;
wire n_785;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_853;
wire n_810;
wire n_843;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_851;
wire n_133;
wire n_494;
wire n_711;
wire n_864;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_845;
wire n_850;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_847;
wire n_779;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_765;
wire n_826;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_831;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_866;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_858;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_456;
wire n_359;
wire n_717;
wire n_312;
wire n_266;
wire n_183;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_861;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_839;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_863;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_836;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_837;
wire n_474;
wire n_829;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_241;
wire n_175;
wire n_687;
wire n_729;
wire n_844;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_854;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_802;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_842;
wire n_259;
wire n_143;
wire n_849;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_855;
wire n_798;
wire n_237;
wire n_668;
wire n_797;
wire n_862;
CKINVDCx5p33_ASAP7_75t_R g621 ( .A(n_0), .Y(n_621) );
AND2x4_ASAP7_75t_L g105 ( .A(n_1), .B(n_106), .Y(n_105) );
AOI22xp5_ASAP7_75t_L g172 ( .A1(n_2), .A2(n_4), .B1(n_173), .B2(n_174), .Y(n_172) );
AOI22xp33_ASAP7_75t_L g141 ( .A1(n_3), .A2(n_20), .B1(n_142), .B2(n_144), .Y(n_141) );
AOI22xp33_ASAP7_75t_L g240 ( .A1(n_5), .A2(n_52), .B1(n_232), .B2(n_241), .Y(n_240) );
BUFx3_ASAP7_75t_L g560 ( .A(n_6), .Y(n_560) );
AOI22xp5_ASAP7_75t_L g295 ( .A1(n_7), .A2(n_13), .B1(n_149), .B2(n_224), .Y(n_295) );
INVx1_ASAP7_75t_L g106 ( .A(n_8), .Y(n_106) );
CKINVDCx5p33_ASAP7_75t_R g195 ( .A(n_9), .Y(n_195) );
NAND2xp5_ASAP7_75t_L g545 ( .A(n_10), .B(n_171), .Y(n_545) );
BUFx2_ASAP7_75t_L g113 ( .A(n_11), .Y(n_113) );
OR2x2_ASAP7_75t_L g124 ( .A(n_11), .B(n_29), .Y(n_124) );
BUFx6f_ASAP7_75t_L g143 ( .A(n_12), .Y(n_143) );
INVx5_ASAP7_75t_SL g865 ( .A(n_14), .Y(n_865) );
NAND2xp5_ASAP7_75t_SL g570 ( .A(n_15), .B(n_247), .Y(n_570) );
NAND2xp5_ASAP7_75t_L g571 ( .A(n_16), .B(n_252), .Y(n_571) );
AOI22xp33_ASAP7_75t_L g592 ( .A1(n_17), .A2(n_86), .B1(n_142), .B2(n_247), .Y(n_592) );
OAI21x1_ASAP7_75t_L g157 ( .A1(n_18), .A2(n_47), .B(n_158), .Y(n_157) );
CKINVDCx5p33_ASAP7_75t_R g163 ( .A(n_19), .Y(n_163) );
NAND2xp5_ASAP7_75t_L g566 ( .A(n_21), .B(n_144), .Y(n_566) );
INVx4_ASAP7_75t_R g260 ( .A(n_22), .Y(n_260) );
NAND2xp5_ASAP7_75t_L g202 ( .A(n_23), .B(n_147), .Y(n_202) );
AO32x1_ASAP7_75t_L g589 ( .A1(n_24), .A2(n_155), .A3(n_156), .B1(n_585), .B2(n_590), .Y(n_589) );
AO32x2_ASAP7_75t_L g624 ( .A1(n_24), .A2(n_155), .A3(n_156), .B1(n_585), .B2(n_590), .Y(n_624) );
INVx1_ASAP7_75t_L g181 ( .A(n_25), .Y(n_181) );
NAND2xp5_ASAP7_75t_SL g210 ( .A(n_26), .B(n_144), .Y(n_210) );
A2O1A1Ixp33_ASAP7_75t_SL g193 ( .A1(n_27), .A2(n_146), .B(n_149), .C(n_194), .Y(n_193) );
AOI22xp33_ASAP7_75t_L g148 ( .A1(n_28), .A2(n_43), .B1(n_149), .B2(n_150), .Y(n_148) );
HB1xp67_ASAP7_75t_L g111 ( .A(n_29), .Y(n_111) );
CKINVDCx5p33_ASAP7_75t_R g190 ( .A(n_30), .Y(n_190) );
AOI22xp33_ASAP7_75t_L g597 ( .A1(n_31), .A2(n_51), .B1(n_144), .B2(n_261), .Y(n_597) );
NAND2xp5_ASAP7_75t_L g580 ( .A(n_32), .B(n_547), .Y(n_580) );
AOI22xp5_ASAP7_75t_L g591 ( .A1(n_33), .A2(n_91), .B1(n_142), .B2(n_150), .Y(n_591) );
NAND2xp5_ASAP7_75t_SL g582 ( .A(n_34), .B(n_531), .Y(n_582) );
INVx1_ASAP7_75t_L g207 ( .A(n_35), .Y(n_207) );
NAND2xp5_ASAP7_75t_L g209 ( .A(n_36), .B(n_149), .Y(n_209) );
AOI22xp33_ASAP7_75t_L g595 ( .A1(n_37), .A2(n_68), .B1(n_150), .B2(n_596), .Y(n_595) );
CKINVDCx5p33_ASAP7_75t_R g225 ( .A(n_38), .Y(n_225) );
OAI22x1_ASAP7_75t_SL g129 ( .A1(n_39), .A2(n_54), .B1(n_130), .B2(n_131), .Y(n_129) );
INVx1_ASAP7_75t_L g131 ( .A(n_39), .Y(n_131) );
INVx2_ASAP7_75t_L g505 ( .A(n_40), .Y(n_505) );
BUFx3_ASAP7_75t_L g109 ( .A(n_41), .Y(n_109) );
INVx1_ASAP7_75t_L g122 ( .A(n_41), .Y(n_122) );
OAI22x1_ASAP7_75t_L g513 ( .A1(n_42), .A2(n_78), .B1(n_514), .B2(n_515), .Y(n_513) );
INVx1_ASAP7_75t_L g515 ( .A(n_42), .Y(n_515) );
NAND2xp5_ASAP7_75t_L g583 ( .A(n_44), .B(n_584), .Y(n_583) );
AOI22xp33_ASAP7_75t_L g296 ( .A1(n_45), .A2(n_85), .B1(n_149), .B2(n_150), .Y(n_296) );
CKINVDCx5p33_ASAP7_75t_R g262 ( .A(n_46), .Y(n_262) );
CKINVDCx5p33_ASAP7_75t_R g617 ( .A(n_48), .Y(n_617) );
CKINVDCx5p33_ASAP7_75t_R g856 ( .A(n_49), .Y(n_856) );
CKINVDCx5p33_ASAP7_75t_R g535 ( .A(n_50), .Y(n_535) );
AOI22xp5_ASAP7_75t_L g530 ( .A1(n_53), .A2(n_79), .B1(n_204), .B2(n_531), .Y(n_530) );
INVx1_ASAP7_75t_L g130 ( .A(n_54), .Y(n_130) );
CKINVDCx5p33_ASAP7_75t_R g299 ( .A(n_55), .Y(n_299) );
AOI22xp33_ASAP7_75t_L g556 ( .A1(n_56), .A2(n_83), .B1(n_142), .B2(n_247), .Y(n_556) );
INVx1_ASAP7_75t_L g158 ( .A(n_57), .Y(n_158) );
AND2x4_ASAP7_75t_L g160 ( .A(n_58), .B(n_161), .Y(n_160) );
INVx1_ASAP7_75t_L g116 ( .A(n_59), .Y(n_116) );
AOI22xp33_ASAP7_75t_L g169 ( .A1(n_60), .A2(n_90), .B1(n_150), .B2(n_170), .Y(n_169) );
AO22x1_ASAP7_75t_L g245 ( .A1(n_61), .A2(n_73), .B1(n_203), .B2(n_246), .Y(n_245) );
NAND2xp5_ASAP7_75t_L g544 ( .A(n_62), .B(n_142), .Y(n_544) );
INVx1_ASAP7_75t_L g161 ( .A(n_63), .Y(n_161) );
AND2x2_ASAP7_75t_L g197 ( .A(n_64), .B(n_155), .Y(n_197) );
NAND2xp5_ASAP7_75t_L g551 ( .A(n_65), .B(n_155), .Y(n_551) );
A2O1A1Ixp33_ASAP7_75t_L g619 ( .A1(n_66), .A2(n_152), .B(n_232), .C(n_620), .Y(n_619) );
NAND3xp33_ASAP7_75t_L g550 ( .A(n_67), .B(n_142), .C(n_549), .Y(n_550) );
CKINVDCx5p33_ASAP7_75t_R g188 ( .A(n_69), .Y(n_188) );
NAND2xp5_ASAP7_75t_L g231 ( .A(n_70), .B(n_232), .Y(n_231) );
AND2x2_ASAP7_75t_L g622 ( .A(n_71), .B(n_266), .Y(n_622) );
CKINVDCx5p33_ASAP7_75t_R g599 ( .A(n_72), .Y(n_599) );
NAND2xp5_ASAP7_75t_L g226 ( .A(n_74), .B(n_144), .Y(n_226) );
AOI22xp33_ASAP7_75t_L g533 ( .A1(n_75), .A2(n_96), .B1(n_204), .B2(n_247), .Y(n_533) );
INVx2_ASAP7_75t_L g147 ( .A(n_76), .Y(n_147) );
NAND2xp5_ASAP7_75t_L g568 ( .A(n_77), .B(n_227), .Y(n_568) );
INVx1_ASAP7_75t_L g514 ( .A(n_78), .Y(n_514) );
NAND2xp5_ASAP7_75t_L g199 ( .A(n_80), .B(n_155), .Y(n_199) );
CKINVDCx5p33_ASAP7_75t_R g257 ( .A(n_81), .Y(n_257) );
CKINVDCx5p33_ASAP7_75t_R g616 ( .A(n_82), .Y(n_616) );
NAND2xp5_ASAP7_75t_L g243 ( .A(n_84), .B(n_165), .Y(n_243) );
NAND2xp5_ASAP7_75t_L g548 ( .A(n_87), .B(n_549), .Y(n_548) );
AOI22xp33_ASAP7_75t_L g557 ( .A1(n_88), .A2(n_100), .B1(n_150), .B2(n_261), .Y(n_557) );
NAND2xp5_ASAP7_75t_SL g579 ( .A(n_89), .B(n_531), .Y(n_579) );
NAND2xp5_ASAP7_75t_SL g221 ( .A(n_92), .B(n_155), .Y(n_221) );
INVx1_ASAP7_75t_L g108 ( .A(n_93), .Y(n_108) );
NOR2xp33_ASAP7_75t_L g120 ( .A(n_93), .B(n_121), .Y(n_120) );
NAND2xp5_ASAP7_75t_L g586 ( .A(n_94), .B(n_252), .Y(n_586) );
A2O1A1Ixp33_ASAP7_75t_L g255 ( .A1(n_95), .A2(n_177), .B(n_232), .C(n_256), .Y(n_255) );
AND2x2_ASAP7_75t_L g265 ( .A(n_97), .B(n_266), .Y(n_265) );
NAND2xp33_ASAP7_75t_L g230 ( .A(n_98), .B(n_171), .Y(n_230) );
CKINVDCx5p33_ASAP7_75t_R g565 ( .A(n_99), .Y(n_565) );
AOI21xp5_ASAP7_75t_L g101 ( .A1(n_102), .A2(n_114), .B(n_864), .Y(n_101) );
AND2x6_ASAP7_75t_L g102 ( .A(n_103), .B(n_110), .Y(n_102) );
AND2x2_ASAP7_75t_SL g866 ( .A(n_103), .B(n_110), .Y(n_866) );
NOR3x1_ASAP7_75t_L g103 ( .A(n_104), .B(n_107), .C(n_109), .Y(n_103) );
INVx2_ASAP7_75t_SL g104 ( .A(n_105), .Y(n_104) );
BUFx6f_ASAP7_75t_L g853 ( .A(n_107), .Y(n_853) );
BUFx2_ASAP7_75t_L g107 ( .A(n_108), .Y(n_107) );
INVx2_ASAP7_75t_L g851 ( .A(n_108), .Y(n_851) );
INVx1_ASAP7_75t_L g511 ( .A(n_109), .Y(n_511) );
NOR2x1_ASAP7_75t_L g863 ( .A(n_109), .B(n_124), .Y(n_863) );
NOR2x1p5_ASAP7_75t_L g110 ( .A(n_111), .B(n_112), .Y(n_110) );
INVx1_ASAP7_75t_L g112 ( .A(n_113), .Y(n_112) );
OR2x6_ASAP7_75t_L g114 ( .A(n_115), .B(n_125), .Y(n_114) );
NOR2xp67_ASAP7_75t_L g126 ( .A(n_115), .B(n_127), .Y(n_126) );
NOR2x1_ASAP7_75t_L g115 ( .A(n_116), .B(n_117), .Y(n_115) );
BUFx2_ASAP7_75t_SL g117 ( .A(n_118), .Y(n_117) );
INVx5_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
CKINVDCx8_ASAP7_75t_R g500 ( .A(n_119), .Y(n_500) );
AND2x6_ASAP7_75t_SL g119 ( .A(n_120), .B(n_123), .Y(n_119) );
INVx1_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
NAND2xp5_ASAP7_75t_L g510 ( .A(n_123), .B(n_511), .Y(n_510) );
INVx1_ASAP7_75t_L g123 ( .A(n_124), .Y(n_123) );
OAI21xp5_ASAP7_75t_L g125 ( .A1(n_126), .A2(n_501), .B(n_506), .Y(n_125) );
AND2x2_ASAP7_75t_L g127 ( .A(n_128), .B(n_497), .Y(n_127) );
XNOR2x1_ASAP7_75t_L g128 ( .A(n_129), .B(n_132), .Y(n_128) );
OA22x2_ASAP7_75t_L g517 ( .A1(n_132), .A2(n_518), .B1(n_850), .B2(n_852), .Y(n_517) );
AND2x4_ASAP7_75t_L g132 ( .A(n_133), .B(n_389), .Y(n_132) );
NOR2xp67_ASAP7_75t_L g133 ( .A(n_134), .B(n_331), .Y(n_133) );
NAND3xp33_ASAP7_75t_SL g134 ( .A(n_135), .B(n_267), .C(n_313), .Y(n_134) );
OAI21xp5_ASAP7_75t_L g135 ( .A1(n_136), .A2(n_212), .B(n_235), .Y(n_135) );
AOI22xp5_ASAP7_75t_L g267 ( .A1(n_136), .A2(n_268), .B1(n_287), .B2(n_300), .Y(n_267) );
AOI22x1_ASAP7_75t_L g393 ( .A1(n_136), .A2(n_394), .B1(n_398), .B2(n_399), .Y(n_393) );
INVx2_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
OR2x2_ASAP7_75t_L g137 ( .A(n_138), .B(n_182), .Y(n_137) );
OR2x2_ASAP7_75t_L g354 ( .A(n_138), .B(n_355), .Y(n_354) );
NAND2xp5_ASAP7_75t_L g138 ( .A(n_139), .B(n_166), .Y(n_138) );
OR2x2_ASAP7_75t_L g217 ( .A(n_139), .B(n_166), .Y(n_217) );
AND2x2_ASAP7_75t_L g271 ( .A(n_139), .B(n_272), .Y(n_271) );
INVx2_ASAP7_75t_SL g279 ( .A(n_139), .Y(n_279) );
BUFx2_ASAP7_75t_L g330 ( .A(n_139), .Y(n_330) );
AO31x2_ASAP7_75t_L g139 ( .A1(n_140), .A2(n_154), .A3(n_159), .B(n_162), .Y(n_139) );
OAI22xp5_ASAP7_75t_L g140 ( .A1(n_141), .A2(n_145), .B1(n_148), .B2(n_151), .Y(n_140) );
NOR2xp33_ASAP7_75t_L g194 ( .A(n_142), .B(n_195), .Y(n_194) );
INVx2_ASAP7_75t_SL g531 ( .A(n_142), .Y(n_531) );
INVx2_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
BUFx6f_ASAP7_75t_L g144 ( .A(n_143), .Y(n_144) );
INVx3_ASAP7_75t_L g149 ( .A(n_143), .Y(n_149) );
BUFx6f_ASAP7_75t_L g150 ( .A(n_143), .Y(n_150) );
BUFx6f_ASAP7_75t_L g171 ( .A(n_143), .Y(n_171) );
INVx1_ASAP7_75t_L g175 ( .A(n_143), .Y(n_175) );
INVx1_ASAP7_75t_L g204 ( .A(n_143), .Y(n_204) );
INVx1_ASAP7_75t_L g232 ( .A(n_143), .Y(n_232) );
INVx1_ASAP7_75t_L g242 ( .A(n_143), .Y(n_242) );
BUFx6f_ASAP7_75t_L g247 ( .A(n_143), .Y(n_247) );
INVx1_ASAP7_75t_L g261 ( .A(n_143), .Y(n_261) );
NOR2xp33_ASAP7_75t_L g187 ( .A(n_144), .B(n_188), .Y(n_187) );
INVx2_ASAP7_75t_L g596 ( .A(n_144), .Y(n_596) );
OAI22xp5_ASAP7_75t_L g615 ( .A1(n_144), .A2(n_261), .B1(n_616), .B2(n_617), .Y(n_615) );
OAI22xp5_ASAP7_75t_L g168 ( .A1(n_145), .A2(n_169), .B1(n_172), .B2(n_176), .Y(n_168) );
OAI22x1_ASAP7_75t_L g294 ( .A1(n_145), .A2(n_176), .B1(n_295), .B2(n_296), .Y(n_294) );
OAI22xp5_ASAP7_75t_L g529 ( .A1(n_145), .A2(n_530), .B1(n_532), .B2(n_533), .Y(n_529) );
OAI22xp5_ASAP7_75t_L g555 ( .A1(n_145), .A2(n_146), .B1(n_556), .B2(n_557), .Y(n_555) );
AOI21xp5_ASAP7_75t_L g581 ( .A1(n_145), .A2(n_582), .B(n_583), .Y(n_581) );
OAI22xp5_ASAP7_75t_L g594 ( .A1(n_145), .A2(n_151), .B1(n_595), .B2(n_597), .Y(n_594) );
INVx6_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
AOI21xp5_ASAP7_75t_L g229 ( .A1(n_146), .A2(n_230), .B(n_231), .Y(n_229) );
NAND2xp5_ASAP7_75t_L g244 ( .A(n_146), .B(n_245), .Y(n_244) );
A2O1A1Ixp33_ASAP7_75t_L g310 ( .A1(n_146), .A2(n_239), .B(n_245), .C(n_249), .Y(n_310) );
AOI21xp5_ASAP7_75t_L g543 ( .A1(n_146), .A2(n_544), .B(n_545), .Y(n_543) );
OAI22xp5_ASAP7_75t_L g590 ( .A1(n_146), .A2(n_191), .B1(n_591), .B2(n_592), .Y(n_590) );
BUFx8_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
INVx2_ASAP7_75t_L g153 ( .A(n_147), .Y(n_153) );
INVx1_ASAP7_75t_L g177 ( .A(n_147), .Y(n_177) );
INVx1_ASAP7_75t_L g192 ( .A(n_147), .Y(n_192) );
INVx4_ASAP7_75t_L g224 ( .A(n_149), .Y(n_224) );
INVx2_ASAP7_75t_L g173 ( .A(n_150), .Y(n_173) );
NAND2xp5_ASAP7_75t_L g205 ( .A(n_150), .B(n_206), .Y(n_205) );
INVx2_ASAP7_75t_L g547 ( .A(n_150), .Y(n_547) );
AOI21xp5_ASAP7_75t_L g208 ( .A1(n_151), .A2(n_209), .B(n_210), .Y(n_208) );
OAI21x1_ASAP7_75t_L g239 ( .A1(n_151), .A2(n_240), .B(n_243), .Y(n_239) );
AOI21x1_ASAP7_75t_L g578 ( .A1(n_151), .A2(n_579), .B(n_580), .Y(n_578) );
INVx2_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
BUFx3_ASAP7_75t_L g152 ( .A(n_153), .Y(n_152) );
INVx2_ASAP7_75t_L g228 ( .A(n_153), .Y(n_228) );
AOI31xp67_ASAP7_75t_L g554 ( .A1(n_154), .A2(n_159), .A3(n_555), .B(n_558), .Y(n_554) );
INVx2_ASAP7_75t_L g154 ( .A(n_155), .Y(n_154) );
NOR2x1_ASAP7_75t_L g233 ( .A(n_155), .B(n_234), .Y(n_233) );
INVx4_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
AND2x2_ASAP7_75t_L g211 ( .A(n_156), .B(n_159), .Y(n_211) );
BUFx3_ASAP7_75t_L g528 ( .A(n_156), .Y(n_528) );
NOR2xp33_ASAP7_75t_L g558 ( .A(n_156), .B(n_559), .Y(n_558) );
INVx2_ASAP7_75t_L g562 ( .A(n_156), .Y(n_562) );
INVx2_ASAP7_75t_SL g576 ( .A(n_156), .Y(n_576) );
NOR2xp33_ASAP7_75t_L g598 ( .A(n_156), .B(n_599), .Y(n_598) );
BUFx6f_ASAP7_75t_L g156 ( .A(n_157), .Y(n_156) );
INVx2_ASAP7_75t_L g165 ( .A(n_157), .Y(n_165) );
INVx1_ASAP7_75t_L g234 ( .A(n_159), .Y(n_234) );
OAI21x1_ASAP7_75t_L g542 ( .A1(n_159), .A2(n_543), .B(n_546), .Y(n_542) );
OAI21x1_ASAP7_75t_L g563 ( .A1(n_159), .A2(n_564), .B(n_567), .Y(n_563) );
BUFx10_ASAP7_75t_L g159 ( .A(n_160), .Y(n_159) );
INVx1_ASAP7_75t_L g179 ( .A(n_160), .Y(n_179) );
INVx1_ASAP7_75t_L g196 ( .A(n_160), .Y(n_196) );
BUFx10_ASAP7_75t_L g264 ( .A(n_160), .Y(n_264) );
AO31x2_ASAP7_75t_L g593 ( .A1(n_160), .A2(n_528), .A3(n_594), .B(n_598), .Y(n_593) );
NOR2xp33_ASAP7_75t_L g162 ( .A(n_163), .B(n_164), .Y(n_162) );
BUFx2_ASAP7_75t_L g167 ( .A(n_164), .Y(n_167) );
NOR2xp33_ASAP7_75t_L g180 ( .A(n_164), .B(n_181), .Y(n_180) );
INVx2_ASAP7_75t_L g266 ( .A(n_164), .Y(n_266) );
NOR2xp33_ASAP7_75t_L g298 ( .A(n_164), .B(n_299), .Y(n_298) );
NOR2xp33_ASAP7_75t_L g534 ( .A(n_164), .B(n_535), .Y(n_534) );
INVx2_ASAP7_75t_L g164 ( .A(n_165), .Y(n_164) );
OAI21xp33_ASAP7_75t_L g249 ( .A1(n_165), .A2(n_196), .B(n_243), .Y(n_249) );
INVx2_ASAP7_75t_L g253 ( .A(n_165), .Y(n_253) );
INVx2_ASAP7_75t_L g297 ( .A(n_165), .Y(n_297) );
AND2x2_ASAP7_75t_L g274 ( .A(n_166), .B(n_198), .Y(n_274) );
INVx1_ASAP7_75t_L g281 ( .A(n_166), .Y(n_281) );
INVx1_ASAP7_75t_L g286 ( .A(n_166), .Y(n_286) );
NAND2xp5_ASAP7_75t_L g349 ( .A(n_166), .B(n_279), .Y(n_349) );
INVx1_ASAP7_75t_L g370 ( .A(n_166), .Y(n_370) );
NOR2xp33_ASAP7_75t_L g440 ( .A(n_166), .B(n_272), .Y(n_440) );
AO31x2_ASAP7_75t_L g166 ( .A1(n_167), .A2(n_168), .A3(n_178), .B(n_180), .Y(n_166) );
AOI21x1_ASAP7_75t_L g184 ( .A1(n_167), .A2(n_185), .B(n_197), .Y(n_184) );
INVx2_ASAP7_75t_L g170 ( .A(n_171), .Y(n_170) );
OAI22xp33_ASAP7_75t_L g259 ( .A1(n_171), .A2(n_260), .B1(n_261), .B2(n_262), .Y(n_259) );
O2A1O1Ixp5_ASAP7_75t_L g564 ( .A1(n_174), .A2(n_191), .B(n_565), .C(n_566), .Y(n_564) );
INVx2_ASAP7_75t_L g174 ( .A(n_175), .Y(n_174) );
NOR2xp33_ASAP7_75t_L g189 ( .A(n_175), .B(n_190), .Y(n_189) );
NAND2xp5_ASAP7_75t_SL g258 ( .A(n_176), .B(n_259), .Y(n_258) );
INVx1_ASAP7_75t_L g176 ( .A(n_177), .Y(n_176) );
INVx1_ASAP7_75t_SL g532 ( .A(n_177), .Y(n_532) );
INVx1_ASAP7_75t_L g618 ( .A(n_177), .Y(n_618) );
AO31x2_ASAP7_75t_L g527 ( .A1(n_178), .A2(n_528), .A3(n_529), .B(n_534), .Y(n_527) );
INVx2_ASAP7_75t_SL g178 ( .A(n_179), .Y(n_178) );
INVx2_ASAP7_75t_SL g585 ( .A(n_179), .Y(n_585) );
INVx1_ASAP7_75t_L g333 ( .A(n_182), .Y(n_333) );
OR2x2_ASAP7_75t_L g385 ( .A(n_182), .B(n_349), .Y(n_385) );
NAND2xp5_ASAP7_75t_L g182 ( .A(n_183), .B(n_198), .Y(n_182) );
AND2x2_ASAP7_75t_L g218 ( .A(n_183), .B(n_219), .Y(n_218) );
OR2x2_ASAP7_75t_L g277 ( .A(n_183), .B(n_278), .Y(n_277) );
INVxp67_ASAP7_75t_L g283 ( .A(n_183), .Y(n_283) );
NAND2xp5_ASAP7_75t_L g361 ( .A(n_183), .B(n_215), .Y(n_361) );
INVx1_ASAP7_75t_L g183 ( .A(n_184), .Y(n_183) );
INVx2_ASAP7_75t_L g272 ( .A(n_184), .Y(n_272) );
AOI21xp5_ASAP7_75t_L g185 ( .A1(n_186), .A2(n_193), .B(n_196), .Y(n_185) );
OAI21xp5_ASAP7_75t_L g186 ( .A1(n_187), .A2(n_189), .B(n_191), .Y(n_186) );
BUFx4f_ASAP7_75t_L g191 ( .A(n_192), .Y(n_191) );
NOR2xp33_ASAP7_75t_L g206 ( .A(n_192), .B(n_207), .Y(n_206) );
INVx1_ASAP7_75t_L g549 ( .A(n_192), .Y(n_549) );
AOI21xp5_ASAP7_75t_L g613 ( .A1(n_196), .A2(n_614), .B(n_619), .Y(n_613) );
INVx3_ASAP7_75t_L g215 ( .A(n_198), .Y(n_215) );
INVx1_ASAP7_75t_L g327 ( .A(n_198), .Y(n_327) );
AND2x2_ASAP7_75t_L g329 ( .A(n_198), .B(n_330), .Y(n_329) );
AND2x2_ASAP7_75t_L g347 ( .A(n_198), .B(n_348), .Y(n_347) );
OR2x2_ASAP7_75t_L g369 ( .A(n_198), .B(n_370), .Y(n_369) );
NAND2x1p5_ASAP7_75t_SL g380 ( .A(n_198), .B(n_356), .Y(n_380) );
NAND2xp5_ASAP7_75t_L g470 ( .A(n_198), .B(n_286), .Y(n_470) );
AND2x4_ASAP7_75t_L g198 ( .A(n_199), .B(n_200), .Y(n_198) );
OAI21xp5_ASAP7_75t_L g200 ( .A1(n_201), .A2(n_208), .B(n_211), .Y(n_200) );
OAI21xp33_ASAP7_75t_SL g201 ( .A1(n_202), .A2(n_203), .B(n_205), .Y(n_201) );
INVx1_ASAP7_75t_L g203 ( .A(n_204), .Y(n_203) );
NOR2xp33_ASAP7_75t_L g620 ( .A(n_204), .B(n_621), .Y(n_620) );
AND2x2_ASAP7_75t_L g212 ( .A(n_213), .B(n_218), .Y(n_212) );
AOI22xp5_ASAP7_75t_L g408 ( .A1(n_213), .A2(n_409), .B1(n_410), .B2(n_412), .Y(n_408) );
AND2x2_ASAP7_75t_L g213 ( .A(n_214), .B(n_216), .Y(n_213) );
NAND2xp5_ASAP7_75t_L g343 ( .A(n_214), .B(n_344), .Y(n_343) );
NAND2xp5_ASAP7_75t_L g464 ( .A(n_214), .B(n_465), .Y(n_464) );
OR2x2_ASAP7_75t_L g487 ( .A(n_214), .B(n_345), .Y(n_487) );
INVx2_ASAP7_75t_L g214 ( .A(n_215), .Y(n_214) );
AND2x4_ASAP7_75t_L g285 ( .A(n_215), .B(n_286), .Y(n_285) );
NAND2xp5_ASAP7_75t_L g355 ( .A(n_215), .B(n_356), .Y(n_355) );
OR2x2_ASAP7_75t_L g375 ( .A(n_215), .B(n_376), .Y(n_375) );
AND2x4_ASAP7_75t_L g326 ( .A(n_216), .B(n_327), .Y(n_326) );
INVx2_ASAP7_75t_L g216 ( .A(n_217), .Y(n_216) );
INVx2_ASAP7_75t_L g416 ( .A(n_217), .Y(n_416) );
OR2x2_ASAP7_75t_L g490 ( .A(n_217), .B(n_417), .Y(n_490) );
INVx1_ASAP7_75t_L g321 ( .A(n_218), .Y(n_321) );
INVx3_ASAP7_75t_L g325 ( .A(n_219), .Y(n_325) );
BUFx2_ASAP7_75t_L g336 ( .A(n_219), .Y(n_336) );
BUFx3_ASAP7_75t_L g219 ( .A(n_220), .Y(n_219) );
AND2x2_ASAP7_75t_L g306 ( .A(n_220), .B(n_250), .Y(n_306) );
INVx2_ASAP7_75t_L g352 ( .A(n_220), .Y(n_352) );
INVx1_ASAP7_75t_L g384 ( .A(n_220), .Y(n_384) );
AND2x2_ASAP7_75t_L g397 ( .A(n_220), .B(n_293), .Y(n_397) );
AND2x2_ASAP7_75t_L g419 ( .A(n_220), .B(n_318), .Y(n_419) );
NAND2x1p5_ASAP7_75t_L g220 ( .A(n_221), .B(n_222), .Y(n_220) );
OAI21x1_ASAP7_75t_L g222 ( .A1(n_223), .A2(n_229), .B(n_233), .Y(n_222) );
O2A1O1Ixp33_ASAP7_75t_L g223 ( .A1(n_224), .A2(n_225), .B(n_226), .C(n_227), .Y(n_223) );
INVx2_ASAP7_75t_SL g227 ( .A(n_228), .Y(n_227) );
OAI22xp5_ASAP7_75t_L g567 ( .A1(n_228), .A2(n_568), .B1(n_569), .B2(n_570), .Y(n_567) );
HB1xp67_ASAP7_75t_L g235 ( .A(n_236), .Y(n_235) );
AND2x2_ASAP7_75t_L g410 ( .A(n_236), .B(n_411), .Y(n_410) );
NAND2xp5_ASAP7_75t_L g418 ( .A(n_236), .B(n_419), .Y(n_418) );
AND2x2_ASAP7_75t_L g435 ( .A(n_236), .B(n_303), .Y(n_435) );
NAND2xp5_ASAP7_75t_L g436 ( .A(n_236), .B(n_437), .Y(n_436) );
AND2x4_ASAP7_75t_L g236 ( .A(n_237), .B(n_250), .Y(n_236) );
INVx2_ASAP7_75t_L g291 ( .A(n_237), .Y(n_291) );
AND2x2_ASAP7_75t_L g319 ( .A(n_237), .B(n_320), .Y(n_319) );
AOI21x1_ASAP7_75t_L g237 ( .A1(n_238), .A2(n_244), .B(n_248), .Y(n_237) );
INVx1_ASAP7_75t_L g238 ( .A(n_239), .Y(n_238) );
INVx2_ASAP7_75t_L g241 ( .A(n_242), .Y(n_241) );
NOR2xp33_ASAP7_75t_L g256 ( .A(n_242), .B(n_257), .Y(n_256) );
INVxp67_ASAP7_75t_SL g246 ( .A(n_247), .Y(n_246) );
INVx3_ASAP7_75t_L g584 ( .A(n_247), .Y(n_584) );
INVx1_ASAP7_75t_L g248 ( .A(n_249), .Y(n_248) );
AND2x2_ASAP7_75t_L g292 ( .A(n_250), .B(n_293), .Y(n_292) );
INVx1_ASAP7_75t_L g312 ( .A(n_250), .Y(n_312) );
INVx2_ASAP7_75t_L g320 ( .A(n_250), .Y(n_320) );
OR2x2_ASAP7_75t_L g340 ( .A(n_250), .B(n_293), .Y(n_340) );
AND2x2_ASAP7_75t_L g351 ( .A(n_250), .B(n_352), .Y(n_351) );
AO21x2_ASAP7_75t_L g250 ( .A1(n_251), .A2(n_254), .B(n_265), .Y(n_250) );
AOI21x1_ASAP7_75t_L g612 ( .A1(n_251), .A2(n_613), .B(n_622), .Y(n_612) );
INVx2_ASAP7_75t_L g251 ( .A(n_252), .Y(n_251) );
INVx2_ASAP7_75t_L g252 ( .A(n_253), .Y(n_252) );
AOI21xp5_ASAP7_75t_L g254 ( .A1(n_255), .A2(n_258), .B(n_263), .Y(n_254) );
INVx1_ASAP7_75t_L g569 ( .A(n_261), .Y(n_569) );
INVx2_ASAP7_75t_L g263 ( .A(n_264), .Y(n_263) );
AO31x2_ASAP7_75t_L g293 ( .A1(n_264), .A2(n_294), .A3(n_297), .B(n_298), .Y(n_293) );
OAI221xp5_ASAP7_75t_L g268 ( .A1(n_269), .A2(n_273), .B1(n_275), .B2(n_280), .C(n_282), .Y(n_268) );
INVx1_ASAP7_75t_L g269 ( .A(n_270), .Y(n_269) );
OAI32xp33_ASAP7_75t_L g381 ( .A1(n_270), .A2(n_284), .A3(n_382), .B1(n_385), .B2(n_386), .Y(n_381) );
HB1xp67_ASAP7_75t_L g270 ( .A(n_271), .Y(n_270) );
INVx1_ASAP7_75t_L g371 ( .A(n_271), .Y(n_371) );
AND2x2_ASAP7_75t_L g407 ( .A(n_271), .B(n_285), .Y(n_407) );
INVx1_ASAP7_75t_L g471 ( .A(n_271), .Y(n_471) );
OR2x2_ASAP7_75t_L g345 ( .A(n_272), .B(n_279), .Y(n_345) );
INVx2_ASAP7_75t_L g356 ( .A(n_272), .Y(n_356) );
BUFx2_ASAP7_75t_SL g273 ( .A(n_274), .Y(n_273) );
AND2x2_ASAP7_75t_L g495 ( .A(n_274), .B(n_496), .Y(n_495) );
INVx1_ASAP7_75t_L g275 ( .A(n_276), .Y(n_275) );
INVx1_ASAP7_75t_L g276 ( .A(n_277), .Y(n_276) );
INVxp67_ASAP7_75t_L g482 ( .A(n_277), .Y(n_482) );
INVx1_ASAP7_75t_L g496 ( .A(n_277), .Y(n_496) );
OR2x2_ASAP7_75t_L g376 ( .A(n_278), .B(n_356), .Y(n_376) );
INVx1_ASAP7_75t_L g278 ( .A(n_279), .Y(n_278) );
NOR2xp33_ASAP7_75t_L g398 ( .A(n_280), .B(n_376), .Y(n_398) );
INVx1_ASAP7_75t_L g429 ( .A(n_280), .Y(n_429) );
BUFx3_ASAP7_75t_L g280 ( .A(n_281), .Y(n_280) );
INVx1_ASAP7_75t_L g463 ( .A(n_281), .Y(n_463) );
OR2x2_ASAP7_75t_L g282 ( .A(n_283), .B(n_284), .Y(n_282) );
NAND2x1_ASAP7_75t_L g432 ( .A(n_283), .B(n_433), .Y(n_432) );
OAI21xp5_ASAP7_75t_SL g454 ( .A1(n_284), .A2(n_455), .B(n_460), .Y(n_454) );
INVx2_ASAP7_75t_L g284 ( .A(n_285), .Y(n_284) );
INVx2_ASAP7_75t_SL g287 ( .A(n_288), .Y(n_287) );
NAND2xp5_ASAP7_75t_L g288 ( .A(n_289), .B(n_292), .Y(n_288) );
AND2x2_ASAP7_75t_L g364 ( .A(n_289), .B(n_306), .Y(n_364) );
INVxp67_ASAP7_75t_SL g494 ( .A(n_289), .Y(n_494) );
INVx1_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
INVx2_ASAP7_75t_L g396 ( .A(n_290), .Y(n_396) );
INVx1_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
AND2x2_ASAP7_75t_L g378 ( .A(n_291), .B(n_352), .Y(n_378) );
AND2x2_ASAP7_75t_L g449 ( .A(n_291), .B(n_320), .Y(n_449) );
NAND2xp5_ASAP7_75t_L g324 ( .A(n_292), .B(n_325), .Y(n_324) );
AND2x2_ASAP7_75t_L g377 ( .A(n_292), .B(n_378), .Y(n_377) );
AND2x2_ASAP7_75t_L g456 ( .A(n_292), .B(n_457), .Y(n_456) );
INVx2_ASAP7_75t_L g305 ( .A(n_293), .Y(n_305) );
INVx2_ASAP7_75t_L g318 ( .A(n_293), .Y(n_318) );
NAND2xp5_ASAP7_75t_L g366 ( .A(n_293), .B(n_309), .Y(n_366) );
AND2x2_ASAP7_75t_L g426 ( .A(n_293), .B(n_320), .Y(n_426) );
INVx2_ASAP7_75t_L g541 ( .A(n_297), .Y(n_541) );
NAND2xp33_ASAP7_75t_SL g300 ( .A(n_301), .B(n_307), .Y(n_300) );
INVx2_ASAP7_75t_SL g301 ( .A(n_302), .Y(n_301) );
AND2x2_ASAP7_75t_L g302 ( .A(n_303), .B(n_306), .Y(n_302) );
INVx1_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
INVx1_ASAP7_75t_L g401 ( .A(n_304), .Y(n_401) );
NAND2xp5_ASAP7_75t_L g476 ( .A(n_304), .B(n_384), .Y(n_476) );
INVx1_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
OR2x2_ASAP7_75t_L g308 ( .A(n_305), .B(n_309), .Y(n_308) );
AND2x2_ASAP7_75t_L g437 ( .A(n_305), .B(n_352), .Y(n_437) );
OR2x2_ASAP7_75t_L g307 ( .A(n_308), .B(n_311), .Y(n_307) );
OR2x2_ASAP7_75t_L g382 ( .A(n_308), .B(n_383), .Y(n_382) );
INVx2_ASAP7_75t_L g339 ( .A(n_309), .Y(n_339) );
INVx1_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
INVx1_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
OR2x2_ASAP7_75t_L g365 ( .A(n_312), .B(n_366), .Y(n_365) );
AOI22xp5_ASAP7_75t_L g313 ( .A1(n_314), .A2(n_326), .B1(n_328), .B2(n_329), .Y(n_313) );
OAI21xp33_ASAP7_75t_L g314 ( .A1(n_315), .A2(n_321), .B(n_322), .Y(n_314) );
INVx1_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
AND2x2_ASAP7_75t_L g328 ( .A(n_316), .B(n_325), .Y(n_328) );
BUFx2_ASAP7_75t_L g346 ( .A(n_316), .Y(n_346) );
AND2x2_ASAP7_75t_L g316 ( .A(n_317), .B(n_319), .Y(n_316) );
INVx1_ASAP7_75t_L g357 ( .A(n_317), .Y(n_357) );
INVx1_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
AND2x2_ASAP7_75t_L g372 ( .A(n_319), .B(n_336), .Y(n_372) );
INVx2_ASAP7_75t_L g388 ( .A(n_319), .Y(n_388) );
AND2x2_ASAP7_75t_L g430 ( .A(n_319), .B(n_352), .Y(n_430) );
INVx1_ASAP7_75t_L g322 ( .A(n_323), .Y(n_322) );
INVx1_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
AND2x2_ASAP7_75t_L g405 ( .A(n_325), .B(n_406), .Y(n_405) );
AND2x2_ASAP7_75t_L g452 ( .A(n_326), .B(n_453), .Y(n_452) );
INVx1_ASAP7_75t_L g483 ( .A(n_327), .Y(n_483) );
INVx2_ASAP7_75t_L g422 ( .A(n_330), .Y(n_422) );
NAND4xp25_ASAP7_75t_L g331 ( .A(n_332), .B(n_341), .C(n_358), .D(n_373), .Y(n_331) );
NAND2xp33_ASAP7_75t_SL g332 ( .A(n_333), .B(n_334), .Y(n_332) );
AOI221xp5_ASAP7_75t_L g427 ( .A1(n_334), .A2(n_412), .B1(n_428), .B2(n_430), .C(n_431), .Y(n_427) );
INVx2_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
NAND2x1_ASAP7_75t_L g335 ( .A(n_336), .B(n_337), .Y(n_335) );
INVx2_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
INVx1_ASAP7_75t_L g409 ( .A(n_338), .Y(n_409) );
OR2x2_ASAP7_75t_L g338 ( .A(n_339), .B(n_340), .Y(n_338) );
INVx2_ASAP7_75t_L g402 ( .A(n_339), .Y(n_402) );
INVx2_ASAP7_75t_L g474 ( .A(n_340), .Y(n_474) );
AOI222xp33_ASAP7_75t_L g341 ( .A1(n_342), .A2(n_346), .B1(n_347), .B2(n_350), .C1(n_353), .C2(n_357), .Y(n_341) );
INVx1_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
AND2x2_ASAP7_75t_L g428 ( .A(n_344), .B(n_429), .Y(n_428) );
AOI21xp5_ASAP7_75t_L g455 ( .A1(n_344), .A2(n_456), .B(n_458), .Y(n_455) );
INVx1_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
OR2x2_ASAP7_75t_L g467 ( .A(n_345), .B(n_411), .Y(n_467) );
OAI21xp33_ASAP7_75t_SL g441 ( .A1(n_346), .A2(n_367), .B(n_442), .Y(n_441) );
INVx1_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
OR2x2_ASAP7_75t_L g360 ( .A(n_349), .B(n_361), .Y(n_360) );
INVxp67_ASAP7_75t_SL g412 ( .A(n_349), .Y(n_412) );
HB1xp67_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
BUFx2_ASAP7_75t_L g411 ( .A(n_352), .Y(n_411) );
INVx1_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
INVx1_ASAP7_75t_L g417 ( .A(n_356), .Y(n_417) );
AOI22xp33_ASAP7_75t_SL g358 ( .A1(n_359), .A2(n_362), .B1(n_367), .B2(n_372), .Y(n_358) );
INVx1_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
NAND2xp5_ASAP7_75t_L g362 ( .A(n_363), .B(n_365), .Y(n_362) );
INVx2_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
AOI221xp5_ASAP7_75t_L g373 ( .A1(n_364), .A2(n_374), .B1(n_377), .B2(n_379), .C(n_381), .Y(n_373) );
INVx3_ASAP7_75t_R g488 ( .A(n_365), .Y(n_488) );
INVx1_ASAP7_75t_L g406 ( .A(n_366), .Y(n_406) );
INVx2_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
OR2x2_ASAP7_75t_L g368 ( .A(n_369), .B(n_371), .Y(n_368) );
INVxp67_ASAP7_75t_SL g423 ( .A(n_369), .Y(n_423) );
INVx1_ASAP7_75t_L g433 ( .A(n_369), .Y(n_433) );
INVx1_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
NAND2xp5_ASAP7_75t_L g424 ( .A(n_378), .B(n_425), .Y(n_424) );
INVx1_ASAP7_75t_L g451 ( .A(n_378), .Y(n_451) );
AND2x2_ASAP7_75t_L g479 ( .A(n_378), .B(n_426), .Y(n_479) );
INVx2_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
AND2x2_ASAP7_75t_L g473 ( .A(n_383), .B(n_474), .Y(n_473) );
INVx2_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
INVx1_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
INVx3_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
NOR2x1_ASAP7_75t_L g389 ( .A(n_390), .B(n_445), .Y(n_389) );
NAND3xp33_ASAP7_75t_L g390 ( .A(n_391), .B(n_427), .C(n_441), .Y(n_390) );
NOR3xp33_ASAP7_75t_L g391 ( .A(n_392), .B(n_403), .C(n_413), .Y(n_391) );
INVx1_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
OAI21xp33_ASAP7_75t_L g404 ( .A1(n_394), .A2(n_405), .B(n_407), .Y(n_404) );
INVx1_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
NAND2xp5_ASAP7_75t_L g395 ( .A(n_396), .B(n_397), .Y(n_395) );
INVx1_ASAP7_75t_L g444 ( .A(n_396), .Y(n_444) );
AND2x2_ASAP7_75t_L g485 ( .A(n_396), .B(n_474), .Y(n_485) );
NAND2x1_ASAP7_75t_L g443 ( .A(n_397), .B(n_444), .Y(n_443) );
INVx1_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
NAND2xp5_ASAP7_75t_L g400 ( .A(n_401), .B(n_402), .Y(n_400) );
INVx1_ASAP7_75t_L g465 ( .A(n_402), .Y(n_465) );
NAND2xp5_ASAP7_75t_L g403 ( .A(n_404), .B(n_408), .Y(n_403) );
INVx1_ASAP7_75t_L g457 ( .A(n_411), .Y(n_457) );
OAI22xp33_ASAP7_75t_L g413 ( .A1(n_414), .A2(n_418), .B1(n_420), .B2(n_424), .Y(n_413) );
HB1xp67_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
NAND2xp5_ASAP7_75t_L g415 ( .A(n_416), .B(n_417), .Y(n_415) );
INVx1_ASAP7_75t_L g453 ( .A(n_417), .Y(n_453) );
NAND2xp5_ASAP7_75t_L g459 ( .A(n_419), .B(n_449), .Y(n_459) );
NAND2xp5_ASAP7_75t_L g420 ( .A(n_421), .B(n_423), .Y(n_420) );
INVx2_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
INVx1_ASAP7_75t_L g492 ( .A(n_425), .Y(n_492) );
INVx2_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
OAI22xp33_ASAP7_75t_SL g431 ( .A1(n_432), .A2(n_434), .B1(n_436), .B2(n_438), .Y(n_431) );
INVx1_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
INVx1_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
HB1xp67_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
INVx2_ASAP7_75t_SL g442 ( .A(n_443), .Y(n_442) );
NAND2xp5_ASAP7_75t_L g445 ( .A(n_446), .B(n_472), .Y(n_445) );
O2A1O1Ixp33_ASAP7_75t_L g446 ( .A1(n_447), .A2(n_450), .B(n_452), .C(n_454), .Y(n_446) );
INVx1_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
OAI21xp33_ASAP7_75t_L g461 ( .A1(n_448), .A2(n_462), .B(n_464), .Y(n_461) );
INVx2_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
INVx1_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
O2A1O1Ixp5_ASAP7_75t_SL g472 ( .A1(n_452), .A2(n_473), .B(n_475), .C(n_477), .Y(n_472) );
AOI22xp33_ASAP7_75t_L g460 ( .A1(n_456), .A2(n_461), .B1(n_466), .B2(n_468), .Y(n_460) );
INVx1_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
INVx1_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
INVx1_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
INVx1_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
OR2x2_ASAP7_75t_L g469 ( .A(n_470), .B(n_471), .Y(n_469) );
INVx2_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
OAI211xp5_ASAP7_75t_L g477 ( .A1(n_478), .A2(n_480), .B(n_484), .C(n_491), .Y(n_477) );
INVx1_ASAP7_75t_L g478 ( .A(n_479), .Y(n_478) );
INVx2_ASAP7_75t_L g480 ( .A(n_481), .Y(n_480) );
AND2x2_ASAP7_75t_L g481 ( .A(n_482), .B(n_483), .Y(n_481) );
AOI22xp5_ASAP7_75t_L g484 ( .A1(n_485), .A2(n_486), .B1(n_488), .B2(n_489), .Y(n_484) );
INVx2_ASAP7_75t_L g486 ( .A(n_487), .Y(n_486) );
INVx2_ASAP7_75t_L g489 ( .A(n_490), .Y(n_489) );
OAI21xp5_ASAP7_75t_SL g491 ( .A1(n_492), .A2(n_493), .B(n_495), .Y(n_491) );
INVx1_ASAP7_75t_L g493 ( .A(n_494), .Y(n_493) );
BUFx6f_ASAP7_75t_L g497 ( .A(n_498), .Y(n_497) );
INVx3_ASAP7_75t_L g498 ( .A(n_499), .Y(n_498) );
INVx3_ASAP7_75t_L g499 ( .A(n_500), .Y(n_499) );
INVx1_ASAP7_75t_L g501 ( .A(n_502), .Y(n_501) );
BUFx2_ASAP7_75t_L g502 ( .A(n_503), .Y(n_502) );
INVx2_ASAP7_75t_L g503 ( .A(n_504), .Y(n_503) );
INVx3_ASAP7_75t_L g504 ( .A(n_505), .Y(n_504) );
INVx1_ASAP7_75t_L g509 ( .A(n_505), .Y(n_509) );
NOR2xp33_ASAP7_75t_L g860 ( .A(n_505), .B(n_861), .Y(n_860) );
AOI21xp5_ASAP7_75t_L g506 ( .A1(n_507), .A2(n_512), .B(n_855), .Y(n_506) );
BUFx12f_ASAP7_75t_L g507 ( .A(n_508), .Y(n_507) );
AND2x6_ASAP7_75t_SL g508 ( .A(n_509), .B(n_510), .Y(n_508) );
OAI22xp5_ASAP7_75t_L g512 ( .A1(n_513), .A2(n_516), .B1(n_517), .B2(n_854), .Y(n_512) );
INVx1_ASAP7_75t_L g854 ( .A(n_513), .Y(n_854) );
INVx2_ASAP7_75t_L g516 ( .A(n_517), .Y(n_516) );
INVx1_ASAP7_75t_L g518 ( .A(n_519), .Y(n_518) );
OR2x2_ASAP7_75t_L g519 ( .A(n_520), .B(n_738), .Y(n_519) );
NAND4xp25_ASAP7_75t_L g520 ( .A(n_521), .B(n_670), .C(n_697), .D(n_728), .Y(n_520) );
NOR2xp33_ASAP7_75t_L g521 ( .A(n_522), .B(n_636), .Y(n_521) );
OAI21xp33_ASAP7_75t_L g522 ( .A1(n_523), .A2(n_572), .B(n_600), .Y(n_522) );
OR2x2_ASAP7_75t_L g523 ( .A(n_524), .B(n_536), .Y(n_523) );
INVx2_ASAP7_75t_L g524 ( .A(n_525), .Y(n_524) );
OR2x2_ASAP7_75t_L g758 ( .A(n_525), .B(n_647), .Y(n_758) );
AND2x2_ASAP7_75t_L g765 ( .A(n_525), .B(n_766), .Y(n_765) );
INVx2_ASAP7_75t_SL g525 ( .A(n_526), .Y(n_525) );
OR2x2_ASAP7_75t_L g674 ( .A(n_526), .B(n_675), .Y(n_674) );
INVx2_ASAP7_75t_L g526 ( .A(n_527), .Y(n_526) );
AND2x2_ASAP7_75t_L g607 ( .A(n_527), .B(n_553), .Y(n_607) );
AND2x2_ASAP7_75t_L g631 ( .A(n_527), .B(n_632), .Y(n_631) );
INVx1_ASAP7_75t_L g640 ( .A(n_527), .Y(n_640) );
OR2x2_ASAP7_75t_L g648 ( .A(n_527), .B(n_604), .Y(n_648) );
OR2x2_ASAP7_75t_L g669 ( .A(n_527), .B(n_632), .Y(n_669) );
AND2x2_ASAP7_75t_L g678 ( .A(n_527), .B(n_561), .Y(n_678) );
INVx1_ASAP7_75t_L g751 ( .A(n_527), .Y(n_751) );
AND2x2_ASAP7_75t_L g754 ( .A(n_527), .B(n_755), .Y(n_754) );
NAND2xp5_ASAP7_75t_L g536 ( .A(n_537), .B(n_552), .Y(n_536) );
INVx2_ASAP7_75t_L g667 ( .A(n_537), .Y(n_667) );
INVx2_ASAP7_75t_L g537 ( .A(n_538), .Y(n_537) );
INVx1_ASAP7_75t_L g775 ( .A(n_538), .Y(n_775) );
INVx1_ASAP7_75t_L g538 ( .A(n_539), .Y(n_538) );
INVx1_ASAP7_75t_L g720 ( .A(n_539), .Y(n_720) );
INVx2_ASAP7_75t_L g539 ( .A(n_540), .Y(n_539) );
OR2x2_ASAP7_75t_L g647 ( .A(n_540), .B(n_633), .Y(n_647) );
OAI21x1_ASAP7_75t_L g540 ( .A1(n_541), .A2(n_542), .B(n_551), .Y(n_540) );
OAI21xp5_ASAP7_75t_L g605 ( .A1(n_541), .A2(n_542), .B(n_551), .Y(n_605) );
OAI21xp5_ASAP7_75t_L g546 ( .A1(n_547), .A2(n_548), .B(n_550), .Y(n_546) );
HB1xp67_ASAP7_75t_L g829 ( .A(n_552), .Y(n_829) );
AND2x2_ASAP7_75t_L g552 ( .A(n_553), .B(n_561), .Y(n_552) );
INVx2_ASAP7_75t_L g641 ( .A(n_553), .Y(n_641) );
AND2x2_ASAP7_75t_L g679 ( .A(n_553), .B(n_605), .Y(n_679) );
INVx2_ASAP7_75t_L g553 ( .A(n_554), .Y(n_553) );
INVx1_ASAP7_75t_L g633 ( .A(n_554), .Y(n_633) );
CKINVDCx5p33_ASAP7_75t_R g559 ( .A(n_560), .Y(n_559) );
AND2x2_ASAP7_75t_L g635 ( .A(n_561), .B(n_605), .Y(n_635) );
INVx1_ASAP7_75t_L g721 ( .A(n_561), .Y(n_721) );
OA21x2_ASAP7_75t_L g561 ( .A1(n_562), .A2(n_563), .B(n_571), .Y(n_561) );
OA21x2_ASAP7_75t_L g604 ( .A1(n_562), .A2(n_563), .B(n_571), .Y(n_604) );
O2A1O1Ixp33_ASAP7_75t_SL g779 ( .A1(n_572), .A2(n_780), .B(n_781), .C(n_783), .Y(n_779) );
OR2x2_ASAP7_75t_L g572 ( .A(n_573), .B(n_587), .Y(n_572) );
OR2x2_ASAP7_75t_L g727 ( .A(n_573), .B(n_711), .Y(n_727) );
INVxp67_ASAP7_75t_SL g789 ( .A(n_573), .Y(n_789) );
INVx2_ASAP7_75t_L g573 ( .A(n_574), .Y(n_573) );
AND2x2_ASAP7_75t_L g623 ( .A(n_574), .B(n_624), .Y(n_623) );
OR2x2_ASAP7_75t_L g655 ( .A(n_574), .B(n_627), .Y(n_655) );
INVx3_ASAP7_75t_L g657 ( .A(n_574), .Y(n_657) );
INVxp67_ASAP7_75t_L g665 ( .A(n_574), .Y(n_665) );
INVx1_ASAP7_75t_L g675 ( .A(n_574), .Y(n_675) );
BUFx2_ASAP7_75t_L g701 ( .A(n_574), .Y(n_701) );
OR2x2_ASAP7_75t_L g724 ( .A(n_574), .B(n_725), .Y(n_724) );
AND2x2_ASAP7_75t_L g763 ( .A(n_574), .B(n_725), .Y(n_763) );
NAND2xp5_ASAP7_75t_L g811 ( .A(n_574), .B(n_593), .Y(n_811) );
INVx1_ASAP7_75t_L g837 ( .A(n_574), .Y(n_837) );
BUFx6f_ASAP7_75t_L g574 ( .A(n_575), .Y(n_574) );
OAI21x1_ASAP7_75t_L g575 ( .A1(n_576), .A2(n_577), .B(n_586), .Y(n_575) );
OAI21x1_ASAP7_75t_L g577 ( .A1(n_578), .A2(n_581), .B(n_585), .Y(n_577) );
NOR2xp33_ASAP7_75t_L g816 ( .A(n_587), .B(n_655), .Y(n_816) );
INVx2_ASAP7_75t_SL g587 ( .A(n_588), .Y(n_587) );
AND2x2_ASAP7_75t_L g656 ( .A(n_588), .B(n_657), .Y(n_656) );
AND2x2_ASAP7_75t_L g742 ( .A(n_588), .B(n_689), .Y(n_742) );
AND2x2_ASAP7_75t_L g759 ( .A(n_588), .B(n_688), .Y(n_759) );
AND2x2_ASAP7_75t_L g588 ( .A(n_589), .B(n_593), .Y(n_588) );
OR2x2_ASAP7_75t_L g711 ( .A(n_589), .B(n_593), .Y(n_711) );
INVx1_ASAP7_75t_L g778 ( .A(n_589), .Y(n_778) );
INVx1_ASAP7_75t_L g791 ( .A(n_589), .Y(n_791) );
INVx3_ASAP7_75t_L g626 ( .A(n_593), .Y(n_626) );
AND2x2_ASAP7_75t_L g681 ( .A(n_593), .B(n_611), .Y(n_681) );
AND2x2_ASAP7_75t_L g702 ( .A(n_593), .B(n_703), .Y(n_702) );
AOI22xp5_ASAP7_75t_L g600 ( .A1(n_601), .A2(n_608), .B1(n_625), .B2(n_628), .Y(n_600) );
AOI22xp5_ASAP7_75t_L g838 ( .A1(n_601), .A2(n_736), .B1(n_839), .B2(n_841), .Y(n_838) );
INVx3_ASAP7_75t_L g601 ( .A(n_602), .Y(n_601) );
OR2x2_ASAP7_75t_L g602 ( .A(n_603), .B(n_606), .Y(n_602) );
OR2x2_ASAP7_75t_L g750 ( .A(n_603), .B(n_751), .Y(n_750) );
INVx1_ASAP7_75t_L g784 ( .A(n_603), .Y(n_784) );
OR2x2_ASAP7_75t_L g603 ( .A(n_604), .B(n_605), .Y(n_603) );
BUFx2_ASAP7_75t_L g660 ( .A(n_604), .Y(n_660) );
INVx2_ASAP7_75t_SL g684 ( .A(n_604), .Y(n_684) );
AND2x2_ASAP7_75t_L g704 ( .A(n_604), .B(n_640), .Y(n_704) );
INVx1_ASAP7_75t_L g755 ( .A(n_604), .Y(n_755) );
INVx1_ASAP7_75t_L g744 ( .A(n_606), .Y(n_744) );
INVx2_ASAP7_75t_L g606 ( .A(n_607), .Y(n_606) );
AND2x4_ASAP7_75t_L g736 ( .A(n_607), .B(n_718), .Y(n_736) );
AO22x1_ASAP7_75t_L g824 ( .A1(n_608), .A2(n_677), .B1(n_825), .B2(n_826), .Y(n_824) );
AND2x2_ASAP7_75t_L g608 ( .A(n_609), .B(n_623), .Y(n_608) );
INVx1_ASAP7_75t_L g609 ( .A(n_610), .Y(n_609) );
HB1xp67_ASAP7_75t_L g610 ( .A(n_611), .Y(n_610) );
INVx1_ASAP7_75t_L g643 ( .A(n_611), .Y(n_643) );
INVx1_ASAP7_75t_L g652 ( .A(n_611), .Y(n_652) );
INVx1_ASAP7_75t_L g703 ( .A(n_611), .Y(n_703) );
INVx2_ASAP7_75t_L g611 ( .A(n_612), .Y(n_611) );
INVx1_ASAP7_75t_L g627 ( .A(n_612), .Y(n_627) );
NAND2xp5_ASAP7_75t_SL g614 ( .A(n_615), .B(n_618), .Y(n_614) );
AND2x2_ASAP7_75t_L g823 ( .A(n_623), .B(n_733), .Y(n_823) );
AND2x4_ASAP7_75t_L g690 ( .A(n_624), .B(n_626), .Y(n_690) );
INVx1_ASAP7_75t_L g725 ( .A(n_624), .Y(n_725) );
INVx1_ASAP7_75t_L g799 ( .A(n_624), .Y(n_799) );
NAND2xp5_ASAP7_75t_L g664 ( .A(n_625), .B(n_665), .Y(n_664) );
NAND2xp5_ASAP7_75t_L g842 ( .A(n_625), .B(n_843), .Y(n_842) );
AND2x2_ASAP7_75t_L g625 ( .A(n_626), .B(n_627), .Y(n_625) );
AND2x4_ASAP7_75t_L g651 ( .A(n_626), .B(n_652), .Y(n_651) );
INVx1_ASAP7_75t_L g770 ( .A(n_626), .Y(n_770) );
INVx1_ASAP7_75t_L g689 ( .A(n_627), .Y(n_689) );
INVx1_ASAP7_75t_L g709 ( .A(n_627), .Y(n_709) );
OR2x2_ASAP7_75t_L g790 ( .A(n_627), .B(n_791), .Y(n_790) );
INVx2_ASAP7_75t_L g628 ( .A(n_629), .Y(n_628) );
OR2x2_ASAP7_75t_L g629 ( .A(n_630), .B(n_634), .Y(n_629) );
INVx1_ASAP7_75t_L g630 ( .A(n_631), .Y(n_630) );
AND2x2_ASAP7_75t_L g817 ( .A(n_631), .B(n_660), .Y(n_817) );
AND2x2_ASAP7_75t_L g825 ( .A(n_631), .B(n_667), .Y(n_825) );
INVx1_ASAP7_75t_L g632 ( .A(n_633), .Y(n_632) );
OR2x2_ASAP7_75t_L g767 ( .A(n_634), .B(n_717), .Y(n_767) );
INVx1_ASAP7_75t_L g634 ( .A(n_635), .Y(n_634) );
AND2x2_ASAP7_75t_L g638 ( .A(n_635), .B(n_639), .Y(n_638) );
INVx1_ASAP7_75t_SL g745 ( .A(n_635), .Y(n_745) );
OAI211xp5_ASAP7_75t_L g636 ( .A1(n_637), .A2(n_642), .B(n_644), .C(n_662), .Y(n_636) );
OAI322xp33_ASAP7_75t_L g682 ( .A1(n_637), .A2(n_674), .A3(n_683), .B1(n_686), .B2(n_691), .C1(n_694), .C2(n_696), .Y(n_682) );
INVx2_ASAP7_75t_L g637 ( .A(n_638), .Y(n_637) );
AND2x2_ASAP7_75t_L g692 ( .A(n_639), .B(n_693), .Y(n_692) );
INVx2_ASAP7_75t_L g748 ( .A(n_639), .Y(n_748) );
AND2x2_ASAP7_75t_L g639 ( .A(n_640), .B(n_641), .Y(n_639) );
INVx1_ASAP7_75t_L g717 ( .A(n_641), .Y(n_717) );
AND2x2_ASAP7_75t_L g756 ( .A(n_641), .B(n_720), .Y(n_756) );
INVx1_ASAP7_75t_L g849 ( .A(n_641), .Y(n_849) );
INVx1_ASAP7_75t_L g827 ( .A(n_642), .Y(n_827) );
OAI211xp5_ASAP7_75t_L g847 ( .A1(n_642), .A2(n_726), .B(n_769), .C(n_848), .Y(n_847) );
INVx1_ASAP7_75t_L g642 ( .A(n_643), .Y(n_642) );
AOI22xp5_ASAP7_75t_L g644 ( .A1(n_645), .A2(n_649), .B1(n_656), .B2(n_658), .Y(n_644) );
OAI21xp5_ASAP7_75t_L g722 ( .A1(n_645), .A2(n_723), .B(n_726), .Y(n_722) );
INVx1_ASAP7_75t_L g645 ( .A(n_646), .Y(n_645) );
OR2x2_ASAP7_75t_L g646 ( .A(n_647), .B(n_648), .Y(n_646) );
INVx2_ASAP7_75t_L g661 ( .A(n_647), .Y(n_661) );
INVx1_ASAP7_75t_L g685 ( .A(n_647), .Y(n_685) );
INVx1_ASAP7_75t_L g766 ( .A(n_647), .Y(n_766) );
INVx1_ASAP7_75t_L g795 ( .A(n_648), .Y(n_795) );
NAND2xp5_ASAP7_75t_L g649 ( .A(n_650), .B(n_653), .Y(n_649) );
HB1xp67_ASAP7_75t_L g846 ( .A(n_650), .Y(n_846) );
INVx2_ASAP7_75t_L g650 ( .A(n_651), .Y(n_650) );
NAND2x1p5_ASAP7_75t_L g782 ( .A(n_651), .B(n_763), .Y(n_782) );
INVx1_ASAP7_75t_L g733 ( .A(n_652), .Y(n_733) );
INVx1_ASAP7_75t_L g653 ( .A(n_654), .Y(n_653) );
NAND2x1_ASAP7_75t_SL g694 ( .A(n_654), .B(n_695), .Y(n_694) );
INVx3_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
NOR2xp33_ASAP7_75t_L g714 ( .A(n_655), .B(n_690), .Y(n_714) );
AND2x2_ASAP7_75t_L g777 ( .A(n_657), .B(n_778), .Y(n_777) );
AND2x2_ASAP7_75t_L g658 ( .A(n_659), .B(n_661), .Y(n_658) );
INVx1_ASAP7_75t_L g659 ( .A(n_660), .Y(n_659) );
AND2x2_ASAP7_75t_L g676 ( .A(n_660), .B(n_661), .Y(n_676) );
NAND2xp5_ASAP7_75t_L g662 ( .A(n_663), .B(n_666), .Y(n_662) );
INVx1_ASAP7_75t_L g663 ( .A(n_664), .Y(n_663) );
AND2x2_ASAP7_75t_L g830 ( .A(n_665), .B(n_687), .Y(n_830) );
INVx1_ASAP7_75t_L g843 ( .A(n_665), .Y(n_843) );
AND2x2_ASAP7_75t_L g666 ( .A(n_667), .B(n_668), .Y(n_666) );
INVx1_ASAP7_75t_L g747 ( .A(n_667), .Y(n_747) );
NAND2xp5_ASAP7_75t_L g737 ( .A(n_668), .B(n_693), .Y(n_737) );
INVx1_ASAP7_75t_L g780 ( .A(n_668), .Y(n_780) );
INVx1_ASAP7_75t_L g668 ( .A(n_669), .Y(n_668) );
INVx1_ASAP7_75t_L g707 ( .A(n_669), .Y(n_707) );
OR2x2_ASAP7_75t_L g836 ( .A(n_669), .B(n_837), .Y(n_836) );
O2A1O1Ixp5_ASAP7_75t_L g670 ( .A1(n_671), .A2(n_677), .B(n_680), .C(n_682), .Y(n_670) );
INVxp67_ASAP7_75t_SL g671 ( .A(n_672), .Y(n_671) );
NAND2xp5_ASAP7_75t_SL g672 ( .A(n_673), .B(n_676), .Y(n_672) );
INVx1_ASAP7_75t_L g673 ( .A(n_674), .Y(n_673) );
AND2x2_ASAP7_75t_L g769 ( .A(n_675), .B(n_770), .Y(n_769) );
INVx2_ASAP7_75t_L g814 ( .A(n_676), .Y(n_814) );
INVx2_ASAP7_75t_L g807 ( .A(n_677), .Y(n_807) );
AND2x2_ASAP7_75t_L g677 ( .A(n_678), .B(n_679), .Y(n_677) );
AOI21xp5_ASAP7_75t_L g728 ( .A1(n_678), .A2(n_729), .B(n_734), .Y(n_728) );
AND2x2_ASAP7_75t_L g794 ( .A(n_679), .B(n_795), .Y(n_794) );
BUFx2_ASAP7_75t_L g680 ( .A(n_681), .Y(n_680) );
AND2x2_ASAP7_75t_L g762 ( .A(n_681), .B(n_763), .Y(n_762) );
AND2x4_ASAP7_75t_L g776 ( .A(n_681), .B(n_777), .Y(n_776) );
NAND2xp5_ASAP7_75t_L g803 ( .A(n_681), .B(n_804), .Y(n_803) );
NAND2xp5_ASAP7_75t_L g683 ( .A(n_684), .B(n_685), .Y(n_683) );
INVx2_ASAP7_75t_L g693 ( .A(n_684), .Y(n_693) );
NAND2xp5_ASAP7_75t_L g706 ( .A(n_684), .B(n_707), .Y(n_706) );
HB1xp67_ASAP7_75t_L g832 ( .A(n_684), .Y(n_832) );
AOI21xp33_ASAP7_75t_L g734 ( .A1(n_686), .A2(n_735), .B(n_737), .Y(n_734) );
INVx2_ASAP7_75t_L g686 ( .A(n_687), .Y(n_686) );
AND2x2_ASAP7_75t_L g687 ( .A(n_688), .B(n_690), .Y(n_687) );
INVx1_ASAP7_75t_L g688 ( .A(n_689), .Y(n_688) );
INVx3_ASAP7_75t_L g696 ( .A(n_690), .Y(n_696) );
AND2x4_ASAP7_75t_L g821 ( .A(n_690), .B(n_709), .Y(n_821) );
INVx2_ASAP7_75t_SL g691 ( .A(n_692), .Y(n_691) );
INVx2_ASAP7_75t_L g695 ( .A(n_696), .Y(n_695) );
AOI221xp5_ASAP7_75t_L g697 ( .A1(n_698), .A2(n_704), .B1(n_705), .B2(n_708), .C(n_712), .Y(n_697) );
INVx1_ASAP7_75t_L g698 ( .A(n_699), .Y(n_698) );
HB1xp67_ASAP7_75t_L g699 ( .A(n_700), .Y(n_699) );
INVx1_ASAP7_75t_L g818 ( .A(n_700), .Y(n_818) );
NAND2xp5_ASAP7_75t_L g700 ( .A(n_701), .B(n_702), .Y(n_700) );
BUFx2_ASAP7_75t_L g731 ( .A(n_701), .Y(n_731) );
INVx1_ASAP7_75t_L g705 ( .A(n_706), .Y(n_705) );
AND2x2_ASAP7_75t_L g708 ( .A(n_709), .B(n_710), .Y(n_708) );
OR2x2_ASAP7_75t_L g840 ( .A(n_709), .B(n_724), .Y(n_840) );
AND2x4_ASAP7_75t_L g732 ( .A(n_710), .B(n_733), .Y(n_732) );
INVx2_ASAP7_75t_L g710 ( .A(n_711), .Y(n_710) );
OAI21xp5_ASAP7_75t_SL g712 ( .A1(n_713), .A2(n_715), .B(n_722), .Y(n_712) );
INVxp67_ASAP7_75t_L g713 ( .A(n_714), .Y(n_713) );
INVx1_ASAP7_75t_L g715 ( .A(n_716), .Y(n_715) );
AND2x2_ASAP7_75t_L g716 ( .A(n_717), .B(n_718), .Y(n_716) );
AND2x2_ASAP7_75t_L g801 ( .A(n_718), .B(n_751), .Y(n_801) );
INVx2_ASAP7_75t_L g718 ( .A(n_719), .Y(n_718) );
NAND2x1p5_ASAP7_75t_L g719 ( .A(n_720), .B(n_721), .Y(n_719) );
INVx2_ASAP7_75t_L g723 ( .A(n_724), .Y(n_723) );
INVx2_ASAP7_75t_L g726 ( .A(n_727), .Y(n_726) );
INVx1_ASAP7_75t_L g729 ( .A(n_730), .Y(n_729) );
NAND2xp5_ASAP7_75t_L g730 ( .A(n_731), .B(n_732), .Y(n_730) );
INVx1_ASAP7_75t_L g813 ( .A(n_732), .Y(n_813) );
INVx1_ASAP7_75t_L g735 ( .A(n_736), .Y(n_735) );
NAND2xp5_ASAP7_75t_L g822 ( .A(n_736), .B(n_823), .Y(n_822) );
NAND3xp33_ASAP7_75t_SL g738 ( .A(n_739), .B(n_785), .C(n_828), .Y(n_738) );
NOR3xp33_ASAP7_75t_L g739 ( .A(n_740), .B(n_760), .C(n_779), .Y(n_739) );
OAI21xp5_ASAP7_75t_SL g740 ( .A1(n_741), .A2(n_743), .B(n_752), .Y(n_740) );
INVx2_ASAP7_75t_L g741 ( .A(n_742), .Y(n_741) );
AOI211x1_ASAP7_75t_SL g743 ( .A1(n_744), .A2(n_745), .B(n_746), .C(n_749), .Y(n_743) );
OAI322xp33_ASAP7_75t_L g786 ( .A1(n_744), .A2(n_787), .A3(n_792), .B1(n_793), .B2(n_796), .C1(n_800), .C2(n_802), .Y(n_786) );
NOR2xp67_ASAP7_75t_L g746 ( .A(n_747), .B(n_748), .Y(n_746) );
O2A1O1Ixp5_ASAP7_75t_SL g844 ( .A1(n_747), .A2(n_845), .B(n_846), .C(n_847), .Y(n_844) );
INVx3_ASAP7_75t_L g749 ( .A(n_750), .Y(n_749) );
NAND2xp5_ASAP7_75t_L g774 ( .A(n_751), .B(n_775), .Y(n_774) );
OAI21xp5_ASAP7_75t_L g752 ( .A1(n_753), .A2(n_757), .B(n_759), .Y(n_752) );
AOI22xp5_ASAP7_75t_L g815 ( .A1(n_753), .A2(n_816), .B1(n_817), .B2(n_818), .Y(n_815) );
AND2x4_ASAP7_75t_L g753 ( .A(n_754), .B(n_756), .Y(n_753) );
INVx1_ASAP7_75t_L g757 ( .A(n_758), .Y(n_757) );
OAI221xp5_ASAP7_75t_L g760 ( .A1(n_761), .A2(n_764), .B1(n_767), .B2(n_768), .C(n_771), .Y(n_760) );
INVx1_ASAP7_75t_L g761 ( .A(n_762), .Y(n_761) );
INVx1_ASAP7_75t_L g764 ( .A(n_765), .Y(n_764) );
INVx1_ASAP7_75t_L g768 ( .A(n_769), .Y(n_768) );
NAND2xp5_ASAP7_75t_L g771 ( .A(n_772), .B(n_776), .Y(n_771) );
INVx1_ASAP7_75t_L g772 ( .A(n_773), .Y(n_772) );
HB1xp67_ASAP7_75t_L g773 ( .A(n_774), .Y(n_773) );
INVx2_ASAP7_75t_L g805 ( .A(n_778), .Y(n_805) );
INVx1_ASAP7_75t_L g812 ( .A(n_778), .Y(n_812) );
HB1xp67_ASAP7_75t_L g781 ( .A(n_782), .Y(n_781) );
INVx1_ASAP7_75t_L g783 ( .A(n_784), .Y(n_783) );
INVx1_ASAP7_75t_L g792 ( .A(n_784), .Y(n_792) );
NOR4xp25_ASAP7_75t_L g785 ( .A(n_786), .B(n_806), .C(n_819), .D(n_824), .Y(n_785) );
INVx1_ASAP7_75t_L g787 ( .A(n_788), .Y(n_787) );
NOR2x1p5_ASAP7_75t_L g788 ( .A(n_789), .B(n_790), .Y(n_788) );
INVx2_ASAP7_75t_L g793 ( .A(n_794), .Y(n_793) );
INVx1_ASAP7_75t_L g796 ( .A(n_797), .Y(n_796) );
INVx2_ASAP7_75t_L g797 ( .A(n_798), .Y(n_797) );
INVx1_ASAP7_75t_L g798 ( .A(n_799), .Y(n_798) );
INVx2_ASAP7_75t_L g800 ( .A(n_801), .Y(n_800) );
HB1xp67_ASAP7_75t_L g802 ( .A(n_803), .Y(n_802) );
INVx2_ASAP7_75t_L g804 ( .A(n_805), .Y(n_804) );
NOR2xp33_ASAP7_75t_L g826 ( .A(n_805), .B(n_827), .Y(n_826) );
OAI221xp5_ASAP7_75t_L g806 ( .A1(n_807), .A2(n_808), .B1(n_813), .B2(n_814), .C(n_815), .Y(n_806) );
OAI21xp33_ASAP7_75t_L g819 ( .A1(n_807), .A2(n_820), .B(n_822), .Y(n_819) );
INVxp67_ASAP7_75t_L g808 ( .A(n_809), .Y(n_808) );
INVx2_ASAP7_75t_L g809 ( .A(n_810), .Y(n_809) );
OR2x2_ASAP7_75t_L g810 ( .A(n_811), .B(n_812), .Y(n_810) );
INVx1_ASAP7_75t_L g820 ( .A(n_821), .Y(n_820) );
INVx1_ASAP7_75t_L g835 ( .A(n_827), .Y(n_835) );
AOI211xp5_ASAP7_75t_L g828 ( .A1(n_829), .A2(n_830), .B(n_831), .C(n_844), .Y(n_828) );
OAI21xp5_ASAP7_75t_SL g831 ( .A1(n_832), .A2(n_833), .B(n_838), .Y(n_831) );
INVx1_ASAP7_75t_L g833 ( .A(n_834), .Y(n_833) );
NOR2x1_ASAP7_75t_L g834 ( .A(n_835), .B(n_836), .Y(n_834) );
HB1xp67_ASAP7_75t_L g845 ( .A(n_836), .Y(n_845) );
INVx1_ASAP7_75t_L g839 ( .A(n_840), .Y(n_839) );
INVx1_ASAP7_75t_L g841 ( .A(n_842), .Y(n_841) );
INVx1_ASAP7_75t_L g848 ( .A(n_849), .Y(n_848) );
CKINVDCx5p33_ASAP7_75t_R g850 ( .A(n_851), .Y(n_850) );
AND2x2_ASAP7_75t_L g862 ( .A(n_851), .B(n_863), .Y(n_862) );
CKINVDCx5p33_ASAP7_75t_R g852 ( .A(n_853), .Y(n_852) );
NOR2xp33_ASAP7_75t_L g855 ( .A(n_856), .B(n_857), .Y(n_855) );
BUFx6f_ASAP7_75t_L g857 ( .A(n_858), .Y(n_857) );
INVx2_ASAP7_75t_L g858 ( .A(n_859), .Y(n_858) );
BUFx10_ASAP7_75t_L g859 ( .A(n_860), .Y(n_859) );
INVx1_ASAP7_75t_L g861 ( .A(n_862), .Y(n_861) );
NOR2xp33_ASAP7_75t_SL g864 ( .A(n_865), .B(n_866), .Y(n_864) );
endmodule