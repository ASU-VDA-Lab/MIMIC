module fake_jpeg_22079_n_178 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_178);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_178;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_175;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_143;
wire n_17;
wire n_25;
wire n_122;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

INVx3_ASAP7_75t_L g15 ( 
.A(n_10),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_12),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_4),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_8),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_2),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_8),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_4),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

INVx1_ASAP7_75t_SL g30 ( 
.A(n_13),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

CKINVDCx16_ASAP7_75t_R g33 ( 
.A(n_18),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_33),
.B(n_35),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_21),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_34),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_30),
.B(n_0),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_21),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_36),
.B(n_38),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_17),
.B(n_0),
.Y(n_37)
);

AND2x2_ASAP7_75t_L g59 ( 
.A(n_37),
.B(n_42),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g38 ( 
.A(n_23),
.B(n_29),
.Y(n_38)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_31),
.Y(n_39)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_39),
.Y(n_58)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_21),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_40),
.B(n_23),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_18),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_41),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_R g42 ( 
.A(n_30),
.B(n_1),
.Y(n_42)
);

INVx5_ASAP7_75t_L g43 ( 
.A(n_16),
.Y(n_43)
);

BUFx2_ASAP7_75t_L g48 ( 
.A(n_43),
.Y(n_48)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_31),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_44),
.A2(n_15),
.B1(n_24),
.B2(n_27),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_16),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_45),
.Y(n_61)
);

MAJIxp5_ASAP7_75t_L g46 ( 
.A(n_36),
.B(n_37),
.C(n_30),
.Y(n_46)
);

AND2x2_ASAP7_75t_L g78 ( 
.A(n_46),
.B(n_60),
.Y(n_78)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_45),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_47),
.B(n_51),
.Y(n_69)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_45),
.Y(n_51)
);

INVxp67_ASAP7_75t_L g70 ( 
.A(n_52),
.Y(n_70)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_42),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_54),
.B(n_55),
.Y(n_87)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_43),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_39),
.A2(n_15),
.B1(n_24),
.B2(n_27),
.Y(n_56)
);

INVxp67_ASAP7_75t_L g77 ( 
.A(n_56),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_44),
.A2(n_15),
.B1(n_24),
.B2(n_40),
.Y(n_57)
);

INVxp67_ASAP7_75t_L g80 ( 
.A(n_57),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_L g60 ( 
.A(n_34),
.B(n_17),
.C(n_20),
.Y(n_60)
);

INVx13_ASAP7_75t_L g62 ( 
.A(n_41),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_62),
.B(n_3),
.Y(n_85)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_64),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_34),
.Y(n_65)
);

INVx1_ASAP7_75t_SL g90 ( 
.A(n_65),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_41),
.B(n_22),
.Y(n_66)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_66),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_L g67 ( 
.A1(n_44),
.A2(n_25),
.B1(n_19),
.B2(n_28),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_67),
.A2(n_20),
.B1(n_32),
.B2(n_29),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_68),
.A2(n_81),
.B1(n_62),
.B2(n_58),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_59),
.B(n_31),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_71),
.B(n_73),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_L g72 ( 
.A1(n_59),
.A2(n_28),
.B1(n_25),
.B2(n_19),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_72),
.A2(n_50),
.B1(n_14),
.B2(n_9),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_59),
.B(n_16),
.Y(n_73)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_63),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_74),
.B(n_79),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_54),
.A2(n_32),
.B1(n_26),
.B2(n_22),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_76),
.A2(n_55),
.B1(n_51),
.B2(n_47),
.Y(n_92)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_63),
.Y(n_79)
);

O2A1O1Ixp33_ASAP7_75t_L g81 ( 
.A1(n_48),
.A2(n_26),
.B(n_3),
.C(n_4),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_46),
.B(n_1),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_82),
.B(n_83),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_48),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_85),
.B(n_5),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_SL g86 ( 
.A(n_53),
.B(n_7),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_86),
.B(n_13),
.Y(n_101)
);

AND2x2_ASAP7_75t_SL g88 ( 
.A(n_48),
.B(n_5),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_88),
.B(n_50),
.C(n_6),
.Y(n_105)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_60),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_89),
.B(n_91),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_49),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_92),
.B(n_102),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_L g116 ( 
.A1(n_93),
.A2(n_99),
.B1(n_90),
.B2(n_102),
.Y(n_116)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_74),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_95),
.B(n_97),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_71),
.A2(n_58),
.B1(n_61),
.B2(n_63),
.Y(n_96)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_96),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_69),
.Y(n_97)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_68),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_99),
.B(n_101),
.Y(n_125)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_79),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_100),
.B(n_103),
.Y(n_117)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_76),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_81),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_105),
.B(n_106),
.C(n_88),
.Y(n_120)
);

XOR2xp5_ASAP7_75t_L g106 ( 
.A(n_73),
.B(n_82),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_107),
.B(n_9),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_83),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_108),
.B(n_109),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_108),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_111),
.Y(n_128)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_94),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_112),
.B(n_100),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_SL g113 ( 
.A(n_106),
.B(n_89),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_113),
.B(n_122),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_116),
.A2(n_127),
.B1(n_93),
.B2(n_105),
.Y(n_138)
);

AOI21xp5_ASAP7_75t_L g118 ( 
.A1(n_104),
.A2(n_77),
.B(n_70),
.Y(n_118)
);

INVxp67_ASAP7_75t_L g133 ( 
.A(n_118),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_L g131 ( 
.A(n_120),
.B(n_124),
.Y(n_131)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_96),
.Y(n_122)
);

AND2x2_ASAP7_75t_SL g123 ( 
.A(n_104),
.B(n_78),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_123),
.B(n_78),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_SL g124 ( 
.A1(n_98),
.A2(n_87),
.B(n_77),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_97),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_126),
.B(n_84),
.Y(n_136)
);

NOR3xp33_ASAP7_75t_SL g129 ( 
.A(n_126),
.B(n_110),
.C(n_91),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_129),
.B(n_130),
.Y(n_144)
);

INVx5_ASAP7_75t_L g130 ( 
.A(n_115),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_132),
.B(n_137),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_114),
.A2(n_70),
.B1(n_80),
.B2(n_103),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_134),
.A2(n_138),
.B1(n_124),
.B2(n_122),
.Y(n_148)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_136),
.Y(n_145)
);

INVxp67_ASAP7_75t_L g137 ( 
.A(n_117),
.Y(n_137)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_119),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_139),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_114),
.A2(n_80),
.B1(n_78),
.B2(n_92),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_140),
.A2(n_121),
.B1(n_127),
.B2(n_112),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_141),
.B(n_120),
.C(n_123),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_L g154 ( 
.A(n_143),
.B(n_147),
.Y(n_154)
);

XNOR2x1_ASAP7_75t_L g146 ( 
.A(n_133),
.B(n_113),
.Y(n_146)
);

AOI21xp5_ASAP7_75t_L g155 ( 
.A1(n_146),
.A2(n_131),
.B(n_137),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_141),
.B(n_123),
.C(n_118),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_148),
.B(n_149),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_135),
.B(n_123),
.C(n_111),
.Y(n_149)
);

A2O1A1Ixp33_ASAP7_75t_L g152 ( 
.A1(n_151),
.A2(n_134),
.B(n_133),
.C(n_140),
.Y(n_152)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_152),
.Y(n_163)
);

XOR2xp5_ASAP7_75t_L g160 ( 
.A(n_155),
.B(n_147),
.Y(n_160)
);

OA21x2_ASAP7_75t_SL g156 ( 
.A1(n_146),
.A2(n_131),
.B(n_129),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_156),
.B(n_157),
.Y(n_161)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_150),
.Y(n_157)
);

AOI21xp5_ASAP7_75t_SL g158 ( 
.A1(n_144),
.A2(n_128),
.B(n_130),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_158),
.B(n_159),
.Y(n_165)
);

NOR3xp33_ASAP7_75t_SL g159 ( 
.A(n_151),
.B(n_125),
.C(n_121),
.Y(n_159)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_160),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_154),
.B(n_143),
.C(n_149),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_162),
.B(n_75),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_153),
.A2(n_142),
.B1(n_145),
.B2(n_90),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_164),
.A2(n_163),
.B1(n_165),
.B2(n_161),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_166),
.B(n_168),
.Y(n_173)
);

A2O1A1Ixp33_ASAP7_75t_L g167 ( 
.A1(n_160),
.A2(n_159),
.B(n_158),
.C(n_152),
.Y(n_167)
);

AOI21xp5_ASAP7_75t_SL g172 ( 
.A1(n_167),
.A2(n_88),
.B(n_12),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_162),
.B(n_95),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_170),
.B(n_84),
.C(n_75),
.Y(n_171)
);

AND2x2_ASAP7_75t_L g174 ( 
.A(n_171),
.B(n_14),
.Y(n_174)
);

AOI21xp5_ASAP7_75t_L g175 ( 
.A1(n_172),
.A2(n_168),
.B(n_169),
.Y(n_175)
);

AOI21xp5_ASAP7_75t_L g176 ( 
.A1(n_174),
.A2(n_175),
.B(n_173),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_176),
.B(n_65),
.C(n_6),
.Y(n_177)
);

XOR2xp5_ASAP7_75t_L g178 ( 
.A(n_177),
.B(n_5),
.Y(n_178)
);


endmodule