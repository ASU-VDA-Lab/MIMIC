module fake_aes_1569_n_17 (n_1, n_2, n_0, n_17);
input n_1;
input n_2;
input n_0;
output n_17;
wire n_11;
wire n_13;
wire n_16;
wire n_12;
wire n_6;
wire n_4;
wire n_3;
wire n_9;
wire n_5;
wire n_14;
wire n_7;
wire n_15;
wire n_10;
wire n_8;
INVx2_ASAP7_75t_L g3 ( .A(n_2), .Y(n_3) );
INVx2_ASAP7_75t_L g4 ( .A(n_2), .Y(n_4) );
INVx2_ASAP7_75t_L g5 ( .A(n_2), .Y(n_5) );
O2A1O1Ixp33_ASAP7_75t_L g6 ( .A1(n_3), .A2(n_0), .B(n_1), .C(n_2), .Y(n_6) );
NAND2xp5_ASAP7_75t_L g7 ( .A(n_4), .B(n_0), .Y(n_7) );
INVx1_ASAP7_75t_L g8 ( .A(n_7), .Y(n_8) );
INVx2_ASAP7_75t_L g9 ( .A(n_6), .Y(n_9) );
INVx1_ASAP7_75t_L g10 ( .A(n_8), .Y(n_10) );
OR2x2_ASAP7_75t_L g11 ( .A(n_9), .B(n_1), .Y(n_11) );
AOI21xp5_ASAP7_75t_L g12 ( .A1(n_10), .A2(n_9), .B(n_5), .Y(n_12) );
AOI21xp5_ASAP7_75t_L g13 ( .A1(n_11), .A2(n_0), .B(n_1), .Y(n_13) );
NAND3xp33_ASAP7_75t_L g14 ( .A(n_13), .B(n_11), .C(n_1), .Y(n_14) );
HB1xp67_ASAP7_75t_L g15 ( .A(n_12), .Y(n_15) );
AO22x2_ASAP7_75t_L g16 ( .A1(n_14), .A2(n_0), .B1(n_11), .B2(n_13), .Y(n_16) );
NAND2xp5_ASAP7_75t_L g17 ( .A(n_16), .B(n_15), .Y(n_17) );
endmodule