module fake_jpeg_6345_n_158 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_158);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_158;

wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_15;
wire n_124;
wire n_141;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_125;
wire n_80;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_121;
wire n_99;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx11_ASAP7_75t_SL g14 ( 
.A(n_9),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_7),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

INVxp67_ASAP7_75t_L g17 ( 
.A(n_12),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_8),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_8),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_2),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_10),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

INVx13_ASAP7_75t_L g62 ( 
.A(n_30),
.Y(n_62)
);

INVx5_ASAP7_75t_L g31 ( 
.A(n_28),
.Y(n_31)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_31),
.Y(n_70)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_23),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_32),
.B(n_33),
.Y(n_44)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_28),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_15),
.B(n_0),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_34),
.B(n_37),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_23),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_35),
.B(n_39),
.Y(n_47)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_23),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_36),
.B(n_38),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_15),
.B(n_1),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_16),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_23),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_17),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_40),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_16),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_41),
.B(n_29),
.Y(n_50)
);

INVx11_ASAP7_75t_L g42 ( 
.A(n_19),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_42),
.B(n_43),
.Y(n_57)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_19),
.Y(n_43)
);

INVx4_ASAP7_75t_SL g45 ( 
.A(n_31),
.Y(n_45)
);

INVx3_ASAP7_75t_SL g88 ( 
.A(n_45),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g49 ( 
.A1(n_33),
.A2(n_29),
.B1(n_22),
.B2(n_25),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_49),
.B(n_52),
.Y(n_73)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_50),
.Y(n_76)
);

INVx1_ASAP7_75t_SL g51 ( 
.A(n_30),
.Y(n_51)
);

HB1xp67_ASAP7_75t_L g89 ( 
.A(n_51),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_L g52 ( 
.A1(n_42),
.A2(n_22),
.B1(n_25),
.B2(n_26),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_41),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_53),
.B(n_68),
.Y(n_95)
);

INVx1_ASAP7_75t_SL g54 ( 
.A(n_30),
.Y(n_54)
);

OR2x2_ASAP7_75t_L g78 ( 
.A(n_54),
.B(n_5),
.Y(n_78)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_30),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_55),
.B(n_56),
.Y(n_74)
);

AOI21xp5_ASAP7_75t_L g56 ( 
.A1(n_39),
.A2(n_20),
.B(n_18),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_38),
.B(n_43),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_58),
.B(n_4),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_36),
.B(n_20),
.Y(n_60)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_60),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_SL g61 ( 
.A(n_32),
.B(n_26),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_61),
.B(n_69),
.Y(n_91)
);

A2O1A1Ixp33_ASAP7_75t_L g63 ( 
.A1(n_40),
.A2(n_18),
.B(n_24),
.C(n_21),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_SL g87 ( 
.A(n_63),
.B(n_72),
.Y(n_87)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_41),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_64),
.B(n_65),
.Y(n_94)
);

O2A1O1Ixp33_ASAP7_75t_L g65 ( 
.A1(n_40),
.A2(n_27),
.B(n_24),
.C(n_21),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_40),
.A2(n_27),
.B1(n_2),
.B2(n_3),
.Y(n_66)
);

INVxp67_ASAP7_75t_L g75 ( 
.A(n_66),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_35),
.B(n_1),
.Y(n_67)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_67),
.Y(n_81)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_34),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_34),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_L g71 ( 
.A1(n_33),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_71)
);

INVxp67_ASAP7_75t_L g84 ( 
.A(n_71),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_33),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_72)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_77),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_78),
.B(n_79),
.Y(n_99)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_45),
.Y(n_79)
);

INVx8_ASAP7_75t_L g82 ( 
.A(n_45),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_82),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_58),
.B(n_6),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_83),
.B(n_90),
.Y(n_104)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_64),
.Y(n_85)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_85),
.Y(n_113)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_61),
.Y(n_86)
);

INVx13_ASAP7_75t_L g101 ( 
.A(n_86),
.Y(n_101)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_53),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_63),
.B(n_10),
.Y(n_92)
);

NOR3xp33_ASAP7_75t_L g110 ( 
.A(n_92),
.B(n_12),
.C(n_13),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_56),
.B(n_11),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_93),
.B(n_13),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_74),
.B(n_48),
.C(n_47),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_96),
.B(n_97),
.C(n_108),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_SL g97 ( 
.A1(n_93),
.A2(n_57),
.B(n_46),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_87),
.A2(n_49),
.B1(n_70),
.B2(n_44),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_100),
.A2(n_102),
.B1(n_105),
.B2(n_106),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_73),
.A2(n_70),
.B1(n_44),
.B2(n_57),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_84),
.A2(n_70),
.B1(n_46),
.B2(n_69),
.Y(n_105)
);

OA22x2_ASAP7_75t_L g106 ( 
.A1(n_88),
.A2(n_65),
.B1(n_62),
.B2(n_51),
.Y(n_106)
);

OR2x2_ASAP7_75t_L g107 ( 
.A(n_88),
.B(n_48),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_107),
.B(n_110),
.Y(n_118)
);

XOR2xp5_ASAP7_75t_L g108 ( 
.A(n_77),
.B(n_59),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_SL g109 ( 
.A1(n_94),
.A2(n_59),
.B(n_68),
.Y(n_109)
);

XNOR2xp5_ASAP7_75t_L g123 ( 
.A(n_109),
.B(n_88),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_111),
.B(n_83),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_87),
.A2(n_55),
.B1(n_54),
.B2(n_62),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_112),
.A2(n_114),
.B1(n_75),
.B2(n_78),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_84),
.A2(n_75),
.B1(n_86),
.B2(n_91),
.Y(n_114)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_104),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_115),
.B(n_116),
.Y(n_129)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_106),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_117),
.A2(n_123),
.B1(n_111),
.B2(n_98),
.Y(n_135)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_104),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_121),
.B(n_122),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_103),
.Y(n_124)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_124),
.Y(n_130)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_102),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_125),
.B(n_126),
.Y(n_127)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_100),
.Y(n_126)
);

NOR2xp67_ASAP7_75t_SL g128 ( 
.A(n_123),
.B(n_96),
.Y(n_128)
);

AOI221xp5_ASAP7_75t_L g145 ( 
.A1(n_128),
.A2(n_135),
.B1(n_81),
.B2(n_80),
.C(n_76),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_121),
.B(n_119),
.Y(n_131)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_131),
.Y(n_144)
);

NAND4xp25_ASAP7_75t_SL g133 ( 
.A(n_116),
.B(n_106),
.C(n_89),
.D(n_85),
.Y(n_133)
);

AO221x1_ASAP7_75t_L g142 ( 
.A1(n_133),
.A2(n_136),
.B1(n_79),
.B2(n_82),
.C(n_113),
.Y(n_142)
);

AOI322xp5_ASAP7_75t_SL g134 ( 
.A1(n_118),
.A2(n_109),
.A3(n_97),
.B1(n_106),
.B2(n_108),
.C1(n_114),
.C2(n_81),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_SL g137 ( 
.A(n_134),
.B(n_119),
.Y(n_137)
);

INVxp67_ASAP7_75t_L g136 ( 
.A(n_120),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_137),
.B(n_138),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_SL g138 ( 
.A(n_132),
.B(n_98),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_131),
.B(n_126),
.C(n_120),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_139),
.B(n_145),
.C(n_129),
.Y(n_149)
);

OR2x2_ASAP7_75t_L g140 ( 
.A(n_133),
.B(n_125),
.Y(n_140)
);

AND2x2_ASAP7_75t_L g148 ( 
.A(n_140),
.B(n_127),
.Y(n_148)
);

A2O1A1O1Ixp25_ASAP7_75t_L g141 ( 
.A1(n_127),
.A2(n_99),
.B(n_107),
.C(n_101),
.D(n_95),
.Y(n_141)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_142),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_136),
.A2(n_101),
.B1(n_80),
.B2(n_76),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_143),
.B(n_130),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_SL g152 ( 
.A(n_148),
.B(n_141),
.Y(n_152)
);

INVxp67_ASAP7_75t_L g151 ( 
.A(n_150),
.Y(n_151)
);

OAI31xp33_ASAP7_75t_L g154 ( 
.A1(n_152),
.A2(n_148),
.A3(n_140),
.B(n_146),
.Y(n_154)
);

NOR2xp67_ASAP7_75t_SL g153 ( 
.A(n_151),
.B(n_149),
.Y(n_153)
);

INVxp67_ASAP7_75t_L g156 ( 
.A(n_153),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_154),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_155),
.B(n_147),
.Y(n_157)
);

AOI21xp5_ASAP7_75t_SL g158 ( 
.A1(n_157),
.A2(n_156),
.B(n_144),
.Y(n_158)
);


endmodule