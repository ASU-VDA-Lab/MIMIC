module fake_jpeg_13648_n_472 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_472);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_472;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx3_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_8),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_11),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_9),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

BUFx8_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

BUFx4f_ASAP7_75t_SL g29 ( 
.A(n_9),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_0),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

INVx5_ASAP7_75t_L g34 ( 
.A(n_4),
.Y(n_34)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_10),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_6),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_7),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_4),
.Y(n_38)
);

BUFx5_ASAP7_75t_L g39 ( 
.A(n_12),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_11),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_0),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_13),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_1),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_12),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_6),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_1),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_8),
.Y(n_47)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_14),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_17),
.B(n_6),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_SL g107 ( 
.A(n_49),
.B(n_75),
.Y(n_107)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_24),
.Y(n_50)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_50),
.Y(n_100)
);

BUFx5_ASAP7_75t_L g51 ( 
.A(n_20),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g111 ( 
.A(n_51),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_29),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_52),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_29),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_53),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_29),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_54),
.Y(n_132)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_23),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g106 ( 
.A(n_55),
.Y(n_106)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_20),
.Y(n_56)
);

BUFx2_ASAP7_75t_L g152 ( 
.A(n_56),
.Y(n_152)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_28),
.Y(n_57)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_57),
.Y(n_102)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_28),
.Y(n_58)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_58),
.Y(n_105)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_39),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g130 ( 
.A(n_59),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_29),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_60),
.Y(n_134)
);

BUFx5_ASAP7_75t_L g61 ( 
.A(n_39),
.Y(n_61)
);

BUFx12f_ASAP7_75t_L g120 ( 
.A(n_61),
.Y(n_120)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_48),
.Y(n_62)
);

INVx4_ASAP7_75t_L g149 ( 
.A(n_62),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_30),
.Y(n_63)
);

INVx6_ASAP7_75t_L g113 ( 
.A(n_63),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_30),
.Y(n_64)
);

INVx8_ASAP7_75t_L g103 ( 
.A(n_64),
.Y(n_103)
);

BUFx8_ASAP7_75t_L g65 ( 
.A(n_23),
.Y(n_65)
);

BUFx12f_ASAP7_75t_L g139 ( 
.A(n_65),
.Y(n_139)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_33),
.Y(n_66)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_66),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_30),
.Y(n_67)
);

INVx5_ASAP7_75t_L g143 ( 
.A(n_67),
.Y(n_143)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_33),
.Y(n_68)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_68),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_17),
.B(n_15),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_69),
.B(n_73),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_31),
.Y(n_70)
);

INVx5_ASAP7_75t_L g153 ( 
.A(n_70),
.Y(n_153)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_48),
.Y(n_71)
);

INVx4_ASAP7_75t_L g150 ( 
.A(n_71),
.Y(n_150)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_23),
.Y(n_72)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_72),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_43),
.B(n_6),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_31),
.Y(n_74)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_74),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_18),
.B(n_7),
.Y(n_75)
);

HB1xp67_ASAP7_75t_L g76 ( 
.A(n_41),
.Y(n_76)
);

CKINVDCx16_ASAP7_75t_R g137 ( 
.A(n_76),
.Y(n_137)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_23),
.B(n_7),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_77),
.B(n_95),
.Y(n_108)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_16),
.Y(n_78)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_78),
.Y(n_114)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_16),
.Y(n_79)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_79),
.Y(n_115)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_35),
.Y(n_80)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_80),
.Y(n_119)
);

INVx6_ASAP7_75t_L g81 ( 
.A(n_31),
.Y(n_81)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_81),
.Y(n_121)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_35),
.Y(n_82)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_82),
.Y(n_122)
);

INVx5_ASAP7_75t_L g83 ( 
.A(n_34),
.Y(n_83)
);

INVx3_ASAP7_75t_L g125 ( 
.A(n_83),
.Y(n_125)
);

INVx8_ASAP7_75t_L g84 ( 
.A(n_37),
.Y(n_84)
);

INVx3_ASAP7_75t_L g138 ( 
.A(n_84),
.Y(n_138)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_47),
.Y(n_85)
);

INVx3_ASAP7_75t_L g145 ( 
.A(n_85),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_37),
.Y(n_86)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_86),
.Y(n_101)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_19),
.Y(n_87)
);

INVx4_ASAP7_75t_L g136 ( 
.A(n_87),
.Y(n_136)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_47),
.Y(n_88)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_88),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_37),
.Y(n_89)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_89),
.Y(n_148)
);

INVx6_ASAP7_75t_L g90 ( 
.A(n_44),
.Y(n_90)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_90),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_44),
.Y(n_91)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_91),
.Y(n_133)
);

INVx8_ASAP7_75t_L g92 ( 
.A(n_44),
.Y(n_92)
);

INVx1_ASAP7_75t_SL g123 ( 
.A(n_92),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_41),
.Y(n_93)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_93),
.Y(n_144)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_19),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_94),
.B(n_96),
.Y(n_141)
);

BUFx3_ASAP7_75t_L g95 ( 
.A(n_19),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_18),
.B(n_7),
.Y(n_96)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_24),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_97),
.B(n_27),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_56),
.A2(n_41),
.B1(n_34),
.B2(n_22),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g162 ( 
.A1(n_112),
.A2(n_126),
.B1(n_54),
.B2(n_52),
.Y(n_162)
);

AOI22xp33_ASAP7_75t_L g116 ( 
.A1(n_63),
.A2(n_32),
.B1(n_43),
.B2(n_46),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_116),
.A2(n_117),
.B1(n_147),
.B2(n_25),
.Y(n_156)
);

AOI22xp33_ASAP7_75t_L g117 ( 
.A1(n_64),
.A2(n_32),
.B1(n_46),
.B2(n_42),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_55),
.A2(n_19),
.B1(n_22),
.B2(n_38),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_127),
.B(n_129),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_96),
.B(n_45),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_49),
.B(n_45),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_135),
.B(n_140),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_75),
.B(n_21),
.Y(n_140)
);

OA22x2_ASAP7_75t_L g142 ( 
.A1(n_77),
.A2(n_21),
.B1(n_40),
.B2(n_42),
.Y(n_142)
);

OA22x2_ASAP7_75t_SL g178 ( 
.A1(n_142),
.A2(n_38),
.B1(n_36),
.B2(n_22),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_76),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_146),
.B(n_151),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_67),
.A2(n_40),
.B1(n_27),
.B2(n_26),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_73),
.B(n_26),
.Y(n_151)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_148),
.Y(n_154)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_154),
.Y(n_221)
);

CKINVDCx16_ASAP7_75t_R g155 ( 
.A(n_116),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_155),
.B(n_157),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_156),
.A2(n_173),
.B1(n_113),
.B2(n_101),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_100),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_144),
.Y(n_158)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_158),
.Y(n_209)
);

CKINVDCx16_ASAP7_75t_R g159 ( 
.A(n_126),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_159),
.B(n_163),
.Y(n_236)
);

AO22x1_ASAP7_75t_SL g160 ( 
.A1(n_102),
.A2(n_84),
.B1(n_93),
.B2(n_65),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_160),
.B(n_168),
.Y(n_215)
);

HB1xp67_ASAP7_75t_L g161 ( 
.A(n_128),
.Y(n_161)
);

CKINVDCx16_ASAP7_75t_R g219 ( 
.A(n_161),
.Y(n_219)
);

INVxp67_ASAP7_75t_L g229 ( 
.A(n_162),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_117),
.Y(n_163)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_121),
.Y(n_164)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_164),
.Y(n_232)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_133),
.Y(n_165)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_165),
.Y(n_237)
);

INVx3_ASAP7_75t_SL g166 ( 
.A(n_103),
.Y(n_166)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_166),
.Y(n_211)
);

AOI22xp33_ASAP7_75t_SL g167 ( 
.A1(n_152),
.A2(n_25),
.B1(n_60),
.B2(n_53),
.Y(n_167)
);

INVxp67_ASAP7_75t_L g242 ( 
.A(n_167),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_104),
.B(n_0),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_108),
.B(n_91),
.C(n_89),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_169),
.B(n_170),
.C(n_174),
.Y(n_205)
);

AND2x2_ASAP7_75t_L g170 ( 
.A(n_105),
.B(n_38),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_124),
.Y(n_171)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_171),
.Y(n_213)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_114),
.Y(n_172)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_172),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_141),
.A2(n_86),
.B1(n_74),
.B2(n_70),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_107),
.A2(n_38),
.B1(n_36),
.B2(n_22),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_109),
.Y(n_175)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_175),
.Y(n_223)
);

BUFx4f_ASAP7_75t_SL g176 ( 
.A(n_139),
.Y(n_176)
);

BUFx8_ASAP7_75t_L g235 ( 
.A(n_176),
.Y(n_235)
);

AOI21xp33_ASAP7_75t_L g208 ( 
.A1(n_178),
.A2(n_181),
.B(n_199),
.Y(n_208)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_110),
.Y(n_179)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_179),
.Y(n_228)
);

INVx4_ASAP7_75t_L g180 ( 
.A(n_139),
.Y(n_180)
);

INVx4_ASAP7_75t_L g206 ( 
.A(n_180),
.Y(n_206)
);

AOI32xp33_ASAP7_75t_L g181 ( 
.A1(n_111),
.A2(n_36),
.A3(n_8),
.B1(n_2),
.B2(n_3),
.Y(n_181)
);

BUFx2_ASAP7_75t_L g182 ( 
.A(n_118),
.Y(n_182)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_182),
.Y(n_238)
);

AOI22xp33_ASAP7_75t_L g183 ( 
.A1(n_115),
.A2(n_36),
.B1(n_5),
.B2(n_2),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_L g214 ( 
.A1(n_183),
.A2(n_195),
.B1(n_106),
.B2(n_130),
.Y(n_214)
);

INVx11_ASAP7_75t_L g184 ( 
.A(n_139),
.Y(n_184)
);

INVxp33_ASAP7_75t_L g207 ( 
.A(n_184),
.Y(n_207)
);

BUFx2_ASAP7_75t_L g187 ( 
.A(n_118),
.Y(n_187)
);

INVx8_ASAP7_75t_L g204 ( 
.A(n_187),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_142),
.B(n_0),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_188),
.B(n_200),
.Y(n_217)
);

INVx8_ASAP7_75t_L g189 ( 
.A(n_131),
.Y(n_189)
);

INVx5_ASAP7_75t_L g234 ( 
.A(n_189),
.Y(n_234)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_98),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_190),
.B(n_192),
.Y(n_243)
);

INVx4_ASAP7_75t_L g191 ( 
.A(n_131),
.Y(n_191)
);

INVx6_ASAP7_75t_L g230 ( 
.A(n_191),
.Y(n_230)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_98),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_137),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_193),
.Y(n_210)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_119),
.Y(n_194)
);

NAND3xp33_ASAP7_75t_L g241 ( 
.A(n_194),
.B(n_196),
.C(n_197),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_142),
.A2(n_130),
.B1(n_152),
.B2(n_122),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_145),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_99),
.Y(n_197)
);

INVx3_ASAP7_75t_L g198 ( 
.A(n_132),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_198),
.Y(n_222)
);

INVxp67_ASAP7_75t_L g199 ( 
.A(n_112),
.Y(n_199)
);

AND2x2_ASAP7_75t_L g200 ( 
.A(n_149),
.B(n_0),
.Y(n_200)
);

HB1xp67_ASAP7_75t_L g201 ( 
.A(n_136),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_201),
.Y(n_233)
);

INVx5_ASAP7_75t_L g202 ( 
.A(n_132),
.Y(n_202)
);

INVx8_ASAP7_75t_L g240 ( 
.A(n_202),
.Y(n_240)
);

BUFx5_ASAP7_75t_L g203 ( 
.A(n_134),
.Y(n_203)
);

OAI22xp33_ASAP7_75t_L g224 ( 
.A1(n_203),
.A2(n_184),
.B1(n_180),
.B2(n_106),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_L g244 ( 
.A1(n_212),
.A2(n_226),
.B1(n_227),
.B2(n_166),
.Y(n_244)
);

AND2x2_ASAP7_75t_L g246 ( 
.A(n_214),
.B(n_160),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_188),
.A2(n_113),
.B1(n_101),
.B2(n_138),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_220),
.A2(n_225),
.B1(n_231),
.B2(n_202),
.Y(n_258)
);

HB1xp67_ASAP7_75t_L g245 ( 
.A(n_224),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_195),
.A2(n_103),
.B1(n_153),
.B2(n_143),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_156),
.A2(n_123),
.B1(n_125),
.B2(n_150),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_173),
.A2(n_136),
.B1(n_134),
.B2(n_120),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_199),
.A2(n_111),
.B1(n_120),
.B2(n_1),
.Y(n_231)
);

FAx1_ASAP7_75t_SL g239 ( 
.A(n_168),
.B(n_120),
.CI(n_111),
.CON(n_239),
.SN(n_239)
);

NOR2xp33_ASAP7_75t_SL g260 ( 
.A(n_239),
.B(n_200),
.Y(n_260)
);

AND2x2_ASAP7_75t_L g291 ( 
.A(n_244),
.B(n_250),
.Y(n_291)
);

AOI22xp33_ASAP7_75t_L g311 ( 
.A1(n_246),
.A2(n_240),
.B1(n_230),
.B2(n_232),
.Y(n_311)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_209),
.Y(n_247)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_247),
.Y(n_284)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_223),
.Y(n_248)
);

INVx2_ASAP7_75t_L g307 ( 
.A(n_248),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_241),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_249),
.B(n_262),
.Y(n_281)
);

OAI21xp33_ASAP7_75t_L g250 ( 
.A1(n_217),
.A2(n_186),
.B(n_185),
.Y(n_250)
);

AOI32xp33_ASAP7_75t_L g251 ( 
.A1(n_217),
.A2(n_178),
.A3(n_174),
.B1(n_177),
.B2(n_169),
.Y(n_251)
);

OAI21xp5_ASAP7_75t_L g293 ( 
.A1(n_251),
.A2(n_254),
.B(n_274),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_215),
.A2(n_178),
.B1(n_160),
.B2(n_175),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_252),
.A2(n_270),
.B1(n_273),
.B2(n_224),
.Y(n_283)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_209),
.Y(n_253)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_253),
.Y(n_289)
);

OR2x2_ASAP7_75t_L g254 ( 
.A(n_239),
.B(n_158),
.Y(n_254)
);

AOI22xp33_ASAP7_75t_SL g255 ( 
.A1(n_242),
.A2(n_187),
.B1(n_182),
.B2(n_189),
.Y(n_255)
);

AOI22xp33_ASAP7_75t_SL g280 ( 
.A1(n_255),
.A2(n_271),
.B1(n_204),
.B2(n_206),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_205),
.B(n_170),
.C(n_179),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_256),
.B(n_257),
.C(n_228),
.Y(n_292)
);

XOR2xp5_ASAP7_75t_L g257 ( 
.A(n_205),
.B(n_170),
.Y(n_257)
);

BUFx2_ASAP7_75t_L g282 ( 
.A(n_258),
.Y(n_282)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_213),
.Y(n_259)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_259),
.Y(n_294)
);

INVxp67_ASAP7_75t_L g298 ( 
.A(n_260),
.Y(n_298)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_213),
.Y(n_261)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_261),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_239),
.B(n_200),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_215),
.B(n_210),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_263),
.B(n_264),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_210),
.B(n_171),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_233),
.B(n_165),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_265),
.B(n_266),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_216),
.B(n_164),
.Y(n_266)
);

INVx2_ASAP7_75t_SL g267 ( 
.A(n_238),
.Y(n_267)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_267),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_SL g268 ( 
.A(n_236),
.B(n_208),
.Y(n_268)
);

CKINVDCx16_ASAP7_75t_R g297 ( 
.A(n_268),
.Y(n_297)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_223),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_269),
.B(n_272),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_212),
.A2(n_154),
.B1(n_198),
.B2(n_191),
.Y(n_270)
);

BUFx2_ASAP7_75t_L g271 ( 
.A(n_204),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_SL g272 ( 
.A(n_220),
.B(n_243),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_L g273 ( 
.A1(n_229),
.A2(n_192),
.B1(n_190),
.B2(n_203),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_233),
.B(n_176),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_229),
.A2(n_242),
.B1(n_225),
.B2(n_231),
.Y(n_275)
);

OAI21xp5_ASAP7_75t_L g296 ( 
.A1(n_275),
.A2(n_277),
.B(n_207),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_219),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g299 ( 
.A(n_276),
.Y(n_299)
);

CKINVDCx14_ASAP7_75t_R g277 ( 
.A(n_235),
.Y(n_277)
);

INVxp67_ASAP7_75t_L g278 ( 
.A(n_228),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_278),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_226),
.A2(n_176),
.B1(n_2),
.B2(n_3),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_L g306 ( 
.A1(n_279),
.A2(n_234),
.B1(n_237),
.B2(n_230),
.Y(n_306)
);

INVxp67_ASAP7_75t_L g329 ( 
.A(n_280),
.Y(n_329)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_283),
.Y(n_314)
);

OAI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_263),
.A2(n_227),
.B1(n_222),
.B2(n_211),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g336 ( 
.A1(n_285),
.A2(n_290),
.B1(n_301),
.B2(n_306),
.Y(n_336)
);

OAI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_254),
.A2(n_222),
.B1(n_211),
.B2(n_218),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g343 ( 
.A(n_292),
.B(n_300),
.C(n_302),
.Y(n_343)
);

INVxp67_ASAP7_75t_L g339 ( 
.A(n_296),
.Y(n_339)
);

XOR2xp5_ASAP7_75t_L g300 ( 
.A(n_257),
.B(n_218),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_254),
.A2(n_262),
.B1(n_275),
.B2(n_272),
.Y(n_301)
);

XOR2xp5_ASAP7_75t_L g302 ( 
.A(n_256),
.B(n_238),
.Y(n_302)
);

AOI21xp5_ASAP7_75t_L g303 ( 
.A1(n_260),
.A2(n_206),
.B(n_235),
.Y(n_303)
);

OAI21xp5_ASAP7_75t_SL g338 ( 
.A1(n_303),
.A2(n_305),
.B(n_310),
.Y(n_338)
);

OAI21xp33_ASAP7_75t_SL g305 ( 
.A1(n_266),
.A2(n_234),
.B(n_237),
.Y(n_305)
);

AOI22xp33_ASAP7_75t_SL g309 ( 
.A1(n_245),
.A2(n_271),
.B1(n_270),
.B2(n_268),
.Y(n_309)
);

INVxp67_ASAP7_75t_L g341 ( 
.A(n_309),
.Y(n_341)
);

AOI21xp5_ASAP7_75t_L g310 ( 
.A1(n_274),
.A2(n_235),
.B(n_232),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_SL g333 ( 
.A1(n_311),
.A2(n_267),
.B1(n_271),
.B2(n_240),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_264),
.B(n_269),
.C(n_261),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_L g334 ( 
.A(n_312),
.B(n_267),
.Y(n_334)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_265),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_313),
.B(n_276),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_L g315 ( 
.A1(n_282),
.A2(n_251),
.B1(n_258),
.B2(n_252),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_L g352 ( 
.A1(n_315),
.A2(n_325),
.B1(n_291),
.B2(n_285),
.Y(n_352)
);

HB1xp67_ASAP7_75t_L g316 ( 
.A(n_312),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g348 ( 
.A(n_316),
.Y(n_348)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_284),
.Y(n_317)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_317),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_286),
.B(n_259),
.Y(n_318)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_318),
.Y(n_363)
);

CKINVDCx20_ASAP7_75t_R g319 ( 
.A(n_287),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_319),
.B(n_320),
.Y(n_350)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_287),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_SL g345 ( 
.A(n_321),
.B(n_323),
.Y(n_345)
);

INVx4_ASAP7_75t_L g322 ( 
.A(n_307),
.Y(n_322)
);

BUFx2_ASAP7_75t_L g347 ( 
.A(n_322),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_299),
.B(n_249),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_SL g324 ( 
.A(n_286),
.B(n_253),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_SL g361 ( 
.A(n_324),
.B(n_331),
.Y(n_361)
);

OAI22xp5_ASAP7_75t_L g325 ( 
.A1(n_282),
.A2(n_246),
.B1(n_279),
.B2(n_244),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_284),
.Y(n_326)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_326),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_313),
.B(n_288),
.Y(n_327)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_327),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_288),
.B(n_247),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_328),
.B(n_332),
.Y(n_354)
);

XOR2xp5_ASAP7_75t_L g330 ( 
.A(n_302),
.B(n_246),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g353 ( 
.A(n_330),
.B(n_334),
.C(n_300),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_SL g331 ( 
.A(n_290),
.B(n_248),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_308),
.B(n_299),
.Y(n_332)
);

AOI22xp33_ASAP7_75t_SL g351 ( 
.A1(n_333),
.A2(n_282),
.B1(n_329),
.B2(n_341),
.Y(n_351)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_289),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_335),
.B(n_340),
.Y(n_356)
);

NOR2xp33_ASAP7_75t_L g337 ( 
.A(n_308),
.B(n_277),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_SL g367 ( 
.A(n_337),
.B(n_323),
.Y(n_367)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_289),
.Y(n_340)
);

CKINVDCx20_ASAP7_75t_R g342 ( 
.A(n_306),
.Y(n_342)
);

CKINVDCx20_ASAP7_75t_R g359 ( 
.A(n_342),
.Y(n_359)
);

XOR2xp5_ASAP7_75t_L g344 ( 
.A(n_343),
.B(n_292),
.Y(n_344)
);

MAJIxp5_ASAP7_75t_L g374 ( 
.A(n_344),
.B(n_353),
.C(n_358),
.Y(n_374)
);

AND2x2_ASAP7_75t_L g349 ( 
.A(n_332),
.B(n_296),
.Y(n_349)
);

INVxp67_ASAP7_75t_L g390 ( 
.A(n_349),
.Y(n_390)
);

OAI22xp5_ASAP7_75t_L g377 ( 
.A1(n_351),
.A2(n_352),
.B1(n_360),
.B2(n_314),
.Y(n_377)
);

OAI21xp5_ASAP7_75t_SL g355 ( 
.A1(n_339),
.A2(n_291),
.B(n_297),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_SL g378 ( 
.A(n_355),
.B(n_319),
.Y(n_378)
);

OAI21xp5_ASAP7_75t_L g357 ( 
.A1(n_338),
.A2(n_293),
.B(n_301),
.Y(n_357)
);

NOR2xp33_ASAP7_75t_L g388 ( 
.A(n_357),
.B(n_362),
.Y(n_388)
);

MAJIxp5_ASAP7_75t_L g358 ( 
.A(n_343),
.B(n_293),
.C(n_298),
.Y(n_358)
);

OAI22xp5_ASAP7_75t_L g360 ( 
.A1(n_314),
.A2(n_283),
.B1(n_281),
.B2(n_297),
.Y(n_360)
);

AOI21xp5_ASAP7_75t_L g362 ( 
.A1(n_338),
.A2(n_291),
.B(n_310),
.Y(n_362)
);

OAI21xp5_ASAP7_75t_L g364 ( 
.A1(n_327),
.A2(n_303),
.B(n_281),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_364),
.B(n_368),
.Y(n_373)
);

AOI22xp5_ASAP7_75t_L g366 ( 
.A1(n_315),
.A2(n_305),
.B1(n_294),
.B2(n_295),
.Y(n_366)
);

OAI22xp5_ASAP7_75t_SL g384 ( 
.A1(n_366),
.A2(n_336),
.B1(n_331),
.B2(n_342),
.Y(n_384)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_367),
.Y(n_371)
);

INVxp67_ASAP7_75t_L g368 ( 
.A(n_337),
.Y(n_368)
);

MAJIxp5_ASAP7_75t_L g370 ( 
.A(n_330),
.B(n_295),
.C(n_294),
.Y(n_370)
);

MAJIxp5_ASAP7_75t_L g380 ( 
.A(n_370),
.B(n_324),
.C(n_340),
.Y(n_380)
);

NOR2xp33_ASAP7_75t_SL g372 ( 
.A(n_345),
.B(n_321),
.Y(n_372)
);

NOR2x1_ASAP7_75t_L g411 ( 
.A(n_372),
.B(n_379),
.Y(n_411)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_354),
.Y(n_375)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_375),
.Y(n_395)
);

XOR2xp5_ASAP7_75t_L g376 ( 
.A(n_344),
.B(n_334),
.Y(n_376)
);

XOR2xp5_ASAP7_75t_L g409 ( 
.A(n_376),
.B(n_364),
.Y(n_409)
);

AOI22xp5_ASAP7_75t_L g396 ( 
.A1(n_377),
.A2(n_384),
.B1(n_360),
.B2(n_325),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g399 ( 
.A(n_378),
.B(n_381),
.Y(n_399)
);

NOR2xp33_ASAP7_75t_SL g379 ( 
.A(n_345),
.B(n_320),
.Y(n_379)
);

XNOR2xp5_ASAP7_75t_L g397 ( 
.A(n_380),
.B(n_370),
.Y(n_397)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_354),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_369),
.B(n_318),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_382),
.B(n_385),
.Y(n_400)
);

MAJIxp5_ASAP7_75t_L g383 ( 
.A(n_344),
.B(n_336),
.C(n_328),
.Y(n_383)
);

MAJIxp5_ASAP7_75t_L g405 ( 
.A(n_383),
.B(n_386),
.C(n_362),
.Y(n_405)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_356),
.Y(n_385)
);

MAJIxp5_ASAP7_75t_SL g386 ( 
.A(n_349),
.B(n_358),
.C(n_357),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_356),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_387),
.B(n_389),
.Y(n_406)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_350),
.Y(n_389)
);

OAI22xp5_ASAP7_75t_L g391 ( 
.A1(n_352),
.A2(n_351),
.B1(n_366),
.B2(n_369),
.Y(n_391)
);

HB1xp67_ASAP7_75t_L g404 ( 
.A(n_391),
.Y(n_404)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_350),
.Y(n_392)
);

OAI22xp5_ASAP7_75t_L g407 ( 
.A1(n_392),
.A2(n_393),
.B1(n_365),
.B2(n_346),
.Y(n_407)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_346),
.Y(n_393)
);

OAI22xp5_ASAP7_75t_SL g394 ( 
.A1(n_379),
.A2(n_363),
.B1(n_361),
.B2(n_367),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_SL g420 ( 
.A(n_394),
.B(n_397),
.Y(n_420)
);

OAI22xp33_ASAP7_75t_L g419 ( 
.A1(n_396),
.A2(n_402),
.B1(n_392),
.B2(n_385),
.Y(n_419)
);

XNOR2xp5_ASAP7_75t_L g398 ( 
.A(n_374),
.B(n_353),
.Y(n_398)
);

XNOR2xp5_ASAP7_75t_L g426 ( 
.A(n_398),
.B(n_403),
.Y(n_426)
);

NOR2xp33_ASAP7_75t_L g401 ( 
.A(n_380),
.B(n_348),
.Y(n_401)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_401),
.Y(n_414)
);

AOI22xp5_ASAP7_75t_L g402 ( 
.A1(n_384),
.A2(n_349),
.B1(n_359),
.B2(n_363),
.Y(n_402)
);

XNOR2xp5_ASAP7_75t_L g403 ( 
.A(n_374),
.B(n_355),
.Y(n_403)
);

MAJIxp5_ASAP7_75t_L g412 ( 
.A(n_405),
.B(n_410),
.C(n_383),
.Y(n_412)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_407),
.Y(n_422)
);

NOR2xp33_ASAP7_75t_L g408 ( 
.A(n_372),
.B(n_348),
.Y(n_408)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_408),
.Y(n_424)
);

XOR2xp5_ASAP7_75t_L g423 ( 
.A(n_409),
.B(n_382),
.Y(n_423)
);

MAJIxp5_ASAP7_75t_L g410 ( 
.A(n_376),
.B(n_349),
.C(n_361),
.Y(n_410)
);

MAJx2_ASAP7_75t_L g428 ( 
.A(n_412),
.B(n_405),
.C(n_403),
.Y(n_428)
);

AOI21xp5_ASAP7_75t_L g413 ( 
.A1(n_411),
.A2(n_373),
.B(n_388),
.Y(n_413)
);

AOI21xp5_ASAP7_75t_L g429 ( 
.A1(n_413),
.A2(n_416),
.B(n_406),
.Y(n_429)
);

NOR2xp33_ASAP7_75t_L g415 ( 
.A(n_411),
.B(n_371),
.Y(n_415)
);

NOR2xp33_ASAP7_75t_SL g431 ( 
.A(n_415),
.B(n_418),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_399),
.B(n_389),
.Y(n_416)
);

MAJIxp5_ASAP7_75t_L g417 ( 
.A(n_397),
.B(n_386),
.C(n_390),
.Y(n_417)
);

MAJIxp5_ASAP7_75t_L g427 ( 
.A(n_417),
.B(n_409),
.C(n_398),
.Y(n_427)
);

NOR2xp33_ASAP7_75t_L g418 ( 
.A(n_410),
.B(n_371),
.Y(n_418)
);

XOR2xp5_ASAP7_75t_L g438 ( 
.A(n_419),
.B(n_423),
.Y(n_438)
);

AOI22xp5_ASAP7_75t_SL g421 ( 
.A1(n_404),
.A2(n_390),
.B1(n_373),
.B2(n_387),
.Y(n_421)
);

OAI22xp5_ASAP7_75t_SL g437 ( 
.A1(n_421),
.A2(n_359),
.B1(n_347),
.B2(n_365),
.Y(n_437)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_400),
.Y(n_425)
);

AOI22xp33_ASAP7_75t_SL g430 ( 
.A1(n_425),
.A2(n_395),
.B1(n_393),
.B2(n_347),
.Y(n_430)
);

AOI21xp5_ASAP7_75t_L g440 ( 
.A1(n_427),
.A2(n_428),
.B(n_429),
.Y(n_440)
);

AOI21xp5_ASAP7_75t_L g444 ( 
.A1(n_430),
.A2(n_417),
.B(n_423),
.Y(n_444)
);

AO21x1_ASAP7_75t_L g432 ( 
.A1(n_416),
.A2(n_402),
.B(n_381),
.Y(n_432)
);

AOI21xp5_ASAP7_75t_SL g447 ( 
.A1(n_432),
.A2(n_426),
.B(n_304),
.Y(n_447)
);

XNOR2xp5_ASAP7_75t_L g433 ( 
.A(n_412),
.B(n_426),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g441 ( 
.A(n_433),
.B(n_435),
.Y(n_441)
);

NOR2xp33_ASAP7_75t_SL g434 ( 
.A(n_424),
.B(n_375),
.Y(n_434)
);

NOR2xp33_ASAP7_75t_SL g442 ( 
.A(n_434),
.B(n_436),
.Y(n_442)
);

NOR2xp33_ASAP7_75t_L g435 ( 
.A(n_414),
.B(n_396),
.Y(n_435)
);

NOR2xp33_ASAP7_75t_SL g436 ( 
.A(n_413),
.B(n_326),
.Y(n_436)
);

AOI22xp5_ASAP7_75t_L g443 ( 
.A1(n_437),
.A2(n_439),
.B1(n_422),
.B2(n_419),
.Y(n_443)
);

OAI22xp5_ASAP7_75t_SL g439 ( 
.A1(n_421),
.A2(n_317),
.B1(n_335),
.B2(n_347),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_443),
.B(n_444),
.Y(n_454)
);

BUFx24_ASAP7_75t_SL g445 ( 
.A(n_433),
.Y(n_445)
);

NOR2xp33_ASAP7_75t_L g452 ( 
.A(n_445),
.B(n_447),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_L g446 ( 
.A(n_437),
.B(n_420),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_L g455 ( 
.A(n_446),
.B(n_448),
.Y(n_455)
);

OAI22xp5_ASAP7_75t_L g448 ( 
.A1(n_432),
.A2(n_322),
.B1(n_304),
.B2(n_307),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_438),
.B(n_322),
.Y(n_449)
);

AOI21xp5_ASAP7_75t_L g451 ( 
.A1(n_449),
.A2(n_450),
.B(n_438),
.Y(n_451)
);

AOI21xp5_ASAP7_75t_L g450 ( 
.A1(n_431),
.A2(n_333),
.B(n_273),
.Y(n_450)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_451),
.Y(n_460)
);

OAI21xp5_ASAP7_75t_SL g453 ( 
.A1(n_440),
.A2(n_427),
.B(n_428),
.Y(n_453)
);

OAI21xp5_ASAP7_75t_L g462 ( 
.A1(n_453),
.A2(n_456),
.B(n_3),
.Y(n_462)
);

MAJIxp5_ASAP7_75t_L g456 ( 
.A(n_441),
.B(n_439),
.C(n_221),
.Y(n_456)
);

AOI21xp5_ASAP7_75t_L g457 ( 
.A1(n_442),
.A2(n_221),
.B(n_235),
.Y(n_457)
);

OAI21x1_ASAP7_75t_L g463 ( 
.A1(n_457),
.A2(n_458),
.B(n_3),
.Y(n_463)
);

AOI21xp5_ASAP7_75t_L g458 ( 
.A1(n_447),
.A2(n_5),
.B(n_2),
.Y(n_458)
);

INVxp67_ASAP7_75t_L g459 ( 
.A(n_452),
.Y(n_459)
);

MAJIxp5_ASAP7_75t_L g466 ( 
.A(n_459),
.B(n_461),
.C(n_10),
.Y(n_466)
);

INVxp67_ASAP7_75t_L g461 ( 
.A(n_455),
.Y(n_461)
);

MAJIxp5_ASAP7_75t_L g465 ( 
.A(n_462),
.B(n_454),
.C(n_4),
.Y(n_465)
);

INVx2_ASAP7_75t_SL g464 ( 
.A(n_463),
.Y(n_464)
);

MAJIxp5_ASAP7_75t_L g467 ( 
.A(n_465),
.B(n_466),
.C(n_460),
.Y(n_467)
);

OAI321xp33_ASAP7_75t_L g469 ( 
.A1(n_467),
.A2(n_468),
.A3(n_1),
.B1(n_14),
.B2(n_15),
.C(n_332),
.Y(n_469)
);

MAJIxp5_ASAP7_75t_L g468 ( 
.A(n_464),
.B(n_10),
.C(n_11),
.Y(n_468)
);

BUFx24_ASAP7_75t_SL g470 ( 
.A(n_469),
.Y(n_470)
);

OAI21xp5_ASAP7_75t_SL g471 ( 
.A1(n_470),
.A2(n_14),
.B(n_15),
.Y(n_471)
);

MAJIxp5_ASAP7_75t_L g472 ( 
.A(n_471),
.B(n_14),
.C(n_15),
.Y(n_472)
);


endmodule