module fake_jpeg_16848_n_60 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_60);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_60;

wire n_57;
wire n_21;
wire n_53;
wire n_33;
wire n_54;
wire n_45;
wire n_23;
wire n_27;
wire n_55;
wire n_22;
wire n_47;
wire n_51;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_59;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_25;
wire n_31;
wire n_56;
wire n_37;
wire n_43;
wire n_50;
wire n_29;
wire n_32;

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_13),
.B(n_3),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_17),
.Y(n_19)
);

INVx3_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_16),
.Y(n_21)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

INVx8_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

BUFx16f_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_2),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_3),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_8),
.B(n_6),
.Y(n_31)
);

CKINVDCx16_ASAP7_75t_R g32 ( 
.A(n_27),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_32),
.B(n_33),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_27),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_25),
.B(n_0),
.Y(n_34)
);

MAJIxp5_ASAP7_75t_L g42 ( 
.A(n_34),
.B(n_35),
.C(n_36),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_30),
.B(n_1),
.Y(n_35)
);

MAJIxp5_ASAP7_75t_L g36 ( 
.A(n_31),
.B(n_1),
.C(n_4),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_26),
.Y(n_37)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_37),
.Y(n_44)
);

INVx5_ASAP7_75t_L g38 ( 
.A(n_27),
.Y(n_38)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_38),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_24),
.Y(n_39)
);

CKINVDCx14_ASAP7_75t_R g40 ( 
.A(n_18),
.Y(n_40)
);

AND2x2_ASAP7_75t_L g41 ( 
.A(n_28),
.B(n_5),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_L g46 ( 
.A1(n_45),
.A2(n_20),
.B1(n_23),
.B2(n_22),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_46),
.A2(n_47),
.B1(n_45),
.B2(n_35),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g47 ( 
.A1(n_42),
.A2(n_22),
.B1(n_20),
.B2(n_23),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_44),
.B(n_34),
.Y(n_48)
);

XNOR2xp5_ASAP7_75t_L g49 ( 
.A(n_48),
.B(n_42),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_49),
.B(n_50),
.Y(n_51)
);

AO22x1_ASAP7_75t_L g52 ( 
.A1(n_49),
.A2(n_46),
.B1(n_39),
.B2(n_24),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_52),
.B(n_41),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g55 ( 
.A1(n_53),
.A2(n_54),
.B1(n_41),
.B2(n_52),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_SL g54 ( 
.A(n_51),
.B(n_44),
.Y(n_54)
);

AOI21xp5_ASAP7_75t_L g57 ( 
.A1(n_55),
.A2(n_56),
.B(n_43),
.Y(n_57)
);

HB1xp67_ASAP7_75t_L g56 ( 
.A(n_54),
.Y(n_56)
);

AOI21xp5_ASAP7_75t_L g58 ( 
.A1(n_57),
.A2(n_40),
.B(n_29),
.Y(n_58)
);

A2O1A1O1Ixp25_ASAP7_75t_L g59 ( 
.A1(n_58),
.A2(n_10),
.B(n_14),
.C(n_15),
.D(n_19),
.Y(n_59)
);

XNOR2xp5_ASAP7_75t_L g60 ( 
.A(n_59),
.B(n_21),
.Y(n_60)
);


endmodule