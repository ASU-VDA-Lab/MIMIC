module fake_jpeg_31367_n_471 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_471);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_471;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_393;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_15),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_1),
.Y(n_18)
);

CKINVDCx11_ASAP7_75t_R g19 ( 
.A(n_6),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_4),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_9),
.Y(n_28)
);

INVxp67_ASAP7_75t_L g29 ( 
.A(n_15),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_3),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_10),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_3),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_2),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_12),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_10),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_7),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_2),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_11),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_12),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_12),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_3),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_2),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_1),
.Y(n_45)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_13),
.Y(n_46)
);

CKINVDCx14_ASAP7_75t_R g47 ( 
.A(n_0),
.Y(n_47)
);

INVx11_ASAP7_75t_SL g48 ( 
.A(n_11),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_20),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_49),
.Y(n_101)
);

INVx11_ASAP7_75t_L g50 ( 
.A(n_48),
.Y(n_50)
);

INVx5_ASAP7_75t_L g117 ( 
.A(n_50),
.Y(n_117)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_23),
.Y(n_51)
);

INVx2_ASAP7_75t_SL g108 ( 
.A(n_51),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_20),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_52),
.Y(n_110)
);

BUFx24_ASAP7_75t_L g53 ( 
.A(n_48),
.Y(n_53)
);

INVx5_ASAP7_75t_SL g119 ( 
.A(n_53),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_20),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_54),
.Y(n_125)
);

BUFx5_ASAP7_75t_L g55 ( 
.A(n_24),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g114 ( 
.A(n_55),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_29),
.B(n_15),
.Y(n_56)
);

AND2x2_ASAP7_75t_L g107 ( 
.A(n_56),
.B(n_63),
.Y(n_107)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_23),
.Y(n_57)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_57),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_20),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_58),
.Y(n_129)
);

INVx11_ASAP7_75t_L g59 ( 
.A(n_32),
.Y(n_59)
);

INVx5_ASAP7_75t_L g131 ( 
.A(n_59),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_21),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_60),
.Y(n_132)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_46),
.Y(n_61)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_61),
.Y(n_123)
);

INVx2_ASAP7_75t_SL g62 ( 
.A(n_19),
.Y(n_62)
);

INVx1_ASAP7_75t_SL g98 ( 
.A(n_62),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_17),
.B(n_14),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_21),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g148 ( 
.A(n_64),
.Y(n_148)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_23),
.Y(n_65)
);

INVx11_ASAP7_75t_L g105 ( 
.A(n_65),
.Y(n_105)
);

CKINVDCx9p33_ASAP7_75t_R g66 ( 
.A(n_19),
.Y(n_66)
);

INVx8_ASAP7_75t_L g128 ( 
.A(n_66),
.Y(n_128)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_25),
.Y(n_67)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_67),
.Y(n_106)
);

INVx8_ASAP7_75t_L g68 ( 
.A(n_25),
.Y(n_68)
);

INVx8_ASAP7_75t_L g143 ( 
.A(n_68),
.Y(n_143)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_25),
.Y(n_69)
);

INVx3_ASAP7_75t_L g144 ( 
.A(n_69),
.Y(n_144)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_31),
.Y(n_70)
);

INVx6_ASAP7_75t_L g142 ( 
.A(n_70),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_21),
.Y(n_71)
);

INVx4_ASAP7_75t_L g141 ( 
.A(n_71),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g72 ( 
.A1(n_34),
.A2(n_14),
.B1(n_1),
.B2(n_2),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_72),
.A2(n_90),
.B1(n_47),
.B2(n_30),
.Y(n_111)
);

INVx8_ASAP7_75t_L g73 ( 
.A(n_31),
.Y(n_73)
);

BUFx3_ASAP7_75t_L g133 ( 
.A(n_73),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_17),
.B(n_14),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_74),
.B(n_77),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_18),
.B(n_0),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_75),
.B(n_78),
.Y(n_100)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_31),
.Y(n_76)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_76),
.Y(n_138)
);

AOI21xp33_ASAP7_75t_L g77 ( 
.A1(n_16),
.A2(n_1),
.B(n_3),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_18),
.B(n_39),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_21),
.Y(n_79)
);

BUFx12f_ASAP7_75t_L g99 ( 
.A(n_79),
.Y(n_99)
);

INVx6_ASAP7_75t_SL g80 ( 
.A(n_26),
.Y(n_80)
);

INVx6_ASAP7_75t_SL g147 ( 
.A(n_80),
.Y(n_147)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_46),
.Y(n_81)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_81),
.Y(n_113)
);

INVx5_ASAP7_75t_L g82 ( 
.A(n_32),
.Y(n_82)
);

BUFx12f_ASAP7_75t_L g104 ( 
.A(n_82),
.Y(n_104)
);

INVx8_ASAP7_75t_L g83 ( 
.A(n_32),
.Y(n_83)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_83),
.Y(n_121)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_26),
.Y(n_84)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_84),
.Y(n_146)
);

INVx8_ASAP7_75t_L g85 ( 
.A(n_34),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_85),
.B(n_86),
.Y(n_115)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_26),
.Y(n_86)
);

BUFx12f_ASAP7_75t_L g87 ( 
.A(n_26),
.Y(n_87)
);

BUFx12f_ASAP7_75t_L g135 ( 
.A(n_87),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_41),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_88),
.B(n_91),
.Y(n_140)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_16),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_89),
.B(n_94),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_34),
.A2(n_4),
.B1(n_5),
.B2(n_7),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_41),
.Y(n_91)
);

BUFx3_ASAP7_75t_L g92 ( 
.A(n_41),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_92),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_41),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_93),
.B(n_44),
.Y(n_145)
);

BUFx12f_ASAP7_75t_L g94 ( 
.A(n_44),
.Y(n_94)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_24),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_95),
.B(n_24),
.Y(n_118)
);

XOR2xp5_ASAP7_75t_L g97 ( 
.A(n_62),
.B(n_33),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_97),
.B(n_35),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_49),
.A2(n_46),
.B1(n_36),
.B2(n_42),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_102),
.A2(n_103),
.B1(n_111),
.B2(n_122),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_85),
.A2(n_47),
.B1(n_42),
.B2(n_36),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_52),
.A2(n_36),
.B1(n_42),
.B2(n_44),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_112),
.A2(n_120),
.B1(n_134),
.B2(n_91),
.Y(n_153)
);

AND2x2_ASAP7_75t_L g160 ( 
.A(n_118),
.B(n_145),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_54),
.A2(n_58),
.B1(n_71),
.B2(n_93),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_60),
.A2(n_28),
.B1(n_43),
.B2(n_40),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_64),
.A2(n_28),
.B1(n_43),
.B2(n_40),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_L g195 ( 
.A1(n_126),
.A2(n_130),
.B1(n_5),
.B2(n_8),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_57),
.B(n_27),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_SL g187 ( 
.A(n_127),
.B(n_136),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_79),
.A2(n_27),
.B1(n_39),
.B2(n_30),
.Y(n_130)
);

OAI22xp33_ASAP7_75t_L g134 ( 
.A1(n_88),
.A2(n_44),
.B1(n_45),
.B2(n_22),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_76),
.B(n_22),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_95),
.B(n_45),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_SL g193 ( 
.A(n_137),
.B(n_139),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_92),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_116),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_149),
.B(n_150),
.Y(n_206)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_146),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_100),
.B(n_35),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_151),
.B(n_154),
.Y(n_210)
);

OA22x2_ASAP7_75t_L g152 ( 
.A1(n_111),
.A2(n_86),
.B1(n_84),
.B2(n_73),
.Y(n_152)
);

AND2x2_ASAP7_75t_L g214 ( 
.A(n_152),
.B(n_175),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_153),
.A2(n_174),
.B1(n_188),
.B2(n_197),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_107),
.B(n_37),
.Y(n_154)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_113),
.Y(n_155)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_155),
.Y(n_220)
);

AOI22xp33_ASAP7_75t_SL g156 ( 
.A1(n_128),
.A2(n_83),
.B1(n_82),
.B2(n_65),
.Y(n_156)
);

INVxp67_ASAP7_75t_L g204 ( 
.A(n_156),
.Y(n_204)
);

INVxp67_ASAP7_75t_L g157 ( 
.A(n_119),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_157),
.B(n_161),
.Y(n_215)
);

INVx3_ASAP7_75t_L g158 ( 
.A(n_119),
.Y(n_158)
);

INVx1_ASAP7_75t_SL g205 ( 
.A(n_158),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_SL g230 ( 
.A(n_159),
.B(n_105),
.Y(n_230)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_113),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g162 ( 
.A(n_101),
.Y(n_162)
);

BUFx3_ASAP7_75t_L g226 ( 
.A(n_162),
.Y(n_226)
);

AND2x2_ASAP7_75t_SL g163 ( 
.A(n_97),
.B(n_68),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_163),
.B(n_108),
.C(n_120),
.Y(n_203)
);

INVx4_ASAP7_75t_L g164 ( 
.A(n_96),
.Y(n_164)
);

INVx1_ASAP7_75t_SL g213 ( 
.A(n_164),
.Y(n_213)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_138),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_165),
.B(n_169),
.Y(n_235)
);

INVx6_ASAP7_75t_L g166 ( 
.A(n_101),
.Y(n_166)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_166),
.Y(n_222)
);

BUFx6f_ASAP7_75t_L g167 ( 
.A(n_110),
.Y(n_167)
);

HB1xp67_ASAP7_75t_L g236 ( 
.A(n_167),
.Y(n_236)
);

INVx3_ASAP7_75t_L g168 ( 
.A(n_117),
.Y(n_168)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_168),
.Y(n_207)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_123),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_107),
.B(n_33),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_170),
.B(n_179),
.Y(n_201)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_96),
.Y(n_171)
);

CKINVDCx14_ASAP7_75t_R g211 ( 
.A(n_171),
.Y(n_211)
);

CKINVDCx16_ASAP7_75t_R g173 ( 
.A(n_121),
.Y(n_173)
);

BUFx4f_ASAP7_75t_SL g221 ( 
.A(n_173),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_109),
.A2(n_59),
.B1(n_87),
.B2(n_94),
.Y(n_174)
);

OAI21xp33_ASAP7_75t_L g175 ( 
.A1(n_140),
.A2(n_38),
.B(n_37),
.Y(n_175)
);

CKINVDCx16_ASAP7_75t_R g176 ( 
.A(n_115),
.Y(n_176)
);

INVxp67_ASAP7_75t_L g217 ( 
.A(n_176),
.Y(n_217)
);

BUFx4f_ASAP7_75t_L g177 ( 
.A(n_99),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_177),
.Y(n_225)
);

CKINVDCx16_ASAP7_75t_R g178 ( 
.A(n_147),
.Y(n_178)
);

INVxp67_ASAP7_75t_L g219 ( 
.A(n_178),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_98),
.B(n_38),
.Y(n_179)
);

INVx4_ASAP7_75t_L g180 ( 
.A(n_117),
.Y(n_180)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_180),
.Y(n_208)
);

OA22x2_ASAP7_75t_L g181 ( 
.A1(n_112),
.A2(n_70),
.B1(n_87),
.B2(n_94),
.Y(n_181)
);

AND2x2_ASAP7_75t_L g228 ( 
.A(n_181),
.B(n_196),
.Y(n_228)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_106),
.Y(n_182)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_182),
.Y(n_218)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_141),
.Y(n_183)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_183),
.Y(n_233)
);

HB1xp67_ASAP7_75t_L g184 ( 
.A(n_106),
.Y(n_184)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_184),
.Y(n_240)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_141),
.Y(n_185)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_185),
.Y(n_241)
);

AOI22xp33_ASAP7_75t_SL g186 ( 
.A1(n_128),
.A2(n_24),
.B1(n_53),
.B2(n_50),
.Y(n_186)
);

INVxp67_ASAP7_75t_L g227 ( 
.A(n_186),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_103),
.A2(n_24),
.B1(n_53),
.B2(n_7),
.Y(n_188)
);

O2A1O1Ixp33_ASAP7_75t_L g189 ( 
.A1(n_134),
.A2(n_4),
.B(n_5),
.C(n_7),
.Y(n_189)
);

OAI22xp33_ASAP7_75t_L g234 ( 
.A1(n_189),
.A2(n_131),
.B1(n_133),
.B2(n_105),
.Y(n_234)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_144),
.Y(n_190)
);

INVxp67_ASAP7_75t_L g238 ( 
.A(n_190),
.Y(n_238)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_144),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_191),
.Y(n_231)
);

AOI22xp33_ASAP7_75t_SL g192 ( 
.A1(n_98),
.A2(n_4),
.B1(n_5),
.B2(n_8),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_L g229 ( 
.A1(n_192),
.A2(n_114),
.B1(n_142),
.B2(n_143),
.Y(n_229)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_110),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_194),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_195),
.A2(n_108),
.B1(n_148),
.B2(n_132),
.Y(n_200)
);

INVx3_ASAP7_75t_L g196 ( 
.A(n_99),
.Y(n_196)
);

AND2x2_ASAP7_75t_L g197 ( 
.A(n_147),
.B(n_8),
.Y(n_197)
);

AND2x2_ASAP7_75t_L g242 ( 
.A(n_197),
.B(n_198),
.Y(n_242)
);

HB1xp67_ASAP7_75t_L g198 ( 
.A(n_142),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_SL g199 ( 
.A(n_187),
.B(n_124),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_SL g249 ( 
.A(n_199),
.B(n_223),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_200),
.A2(n_202),
.B1(n_224),
.B2(n_229),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_172),
.A2(n_152),
.B1(n_153),
.B2(n_163),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_203),
.B(n_183),
.C(n_114),
.Y(n_267)
);

AND2x2_ASAP7_75t_L g253 ( 
.A(n_209),
.B(n_188),
.Y(n_253)
);

AOI22xp33_ASAP7_75t_L g212 ( 
.A1(n_152),
.A2(n_148),
.B1(n_125),
.B2(n_129),
.Y(n_212)
);

AOI22xp33_ASAP7_75t_L g268 ( 
.A1(n_212),
.A2(n_166),
.B1(n_162),
.B2(n_167),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_163),
.B(n_125),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_216),
.B(n_232),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_SL g223 ( 
.A(n_193),
.B(n_143),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_152),
.A2(n_129),
.B1(n_132),
.B2(n_99),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_SL g245 ( 
.A(n_230),
.B(n_160),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_160),
.B(n_197),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_234),
.A2(n_237),
.B1(n_177),
.B2(n_180),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_160),
.A2(n_131),
.B1(n_104),
.B2(n_133),
.Y(n_237)
);

CKINVDCx16_ASAP7_75t_R g243 ( 
.A(n_215),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_243),
.B(n_247),
.Y(n_282)
);

HB1xp67_ASAP7_75t_L g244 ( 
.A(n_208),
.Y(n_244)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_244),
.Y(n_283)
);

XNOR2x1_ASAP7_75t_L g315 ( 
.A(n_245),
.B(n_267),
.Y(n_315)
);

INVxp33_ASAP7_75t_L g247 ( 
.A(n_215),
.Y(n_247)
);

OA21x2_ASAP7_75t_L g248 ( 
.A1(n_214),
.A2(n_228),
.B(n_202),
.Y(n_248)
);

AND2x2_ASAP7_75t_L g294 ( 
.A(n_248),
.B(n_253),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_SL g250 ( 
.A(n_216),
.B(n_174),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_250),
.B(n_251),
.Y(n_285)
);

OR2x2_ASAP7_75t_L g251 ( 
.A(n_214),
.B(n_189),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_218),
.Y(n_252)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_252),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_232),
.B(n_155),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_255),
.B(n_256),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_214),
.B(n_175),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_203),
.B(n_191),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_257),
.B(n_260),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_199),
.B(n_158),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_258),
.B(n_263),
.Y(n_284)
);

INVx4_ASAP7_75t_L g259 ( 
.A(n_226),
.Y(n_259)
);

INVx2_ASAP7_75t_L g303 ( 
.A(n_259),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_230),
.B(n_157),
.Y(n_260)
);

O2A1O1Ixp33_ASAP7_75t_L g261 ( 
.A1(n_204),
.A2(n_181),
.B(n_177),
.C(n_171),
.Y(n_261)
);

O2A1O1Ixp33_ASAP7_75t_L g302 ( 
.A1(n_261),
.A2(n_219),
.B(n_238),
.C(n_225),
.Y(n_302)
);

OAI21xp5_ASAP7_75t_L g262 ( 
.A1(n_242),
.A2(n_228),
.B(n_227),
.Y(n_262)
);

OAI21xp5_ASAP7_75t_L g309 ( 
.A1(n_262),
.A2(n_213),
.B(n_207),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_223),
.B(n_206),
.Y(n_263)
);

AND2x2_ASAP7_75t_SL g264 ( 
.A(n_201),
.B(n_164),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_264),
.B(n_275),
.Y(n_301)
);

AND2x2_ASAP7_75t_L g265 ( 
.A(n_242),
.B(n_181),
.Y(n_265)
);

OAI21xp5_ASAP7_75t_SL g304 ( 
.A1(n_265),
.A2(n_266),
.B(n_281),
.Y(n_304)
);

AND2x2_ASAP7_75t_L g266 ( 
.A(n_242),
.B(n_181),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_SL g314 ( 
.A1(n_268),
.A2(n_271),
.B1(n_273),
.B2(n_213),
.Y(n_314)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_218),
.Y(n_269)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_269),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_206),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_270),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_217),
.B(n_168),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_272),
.B(n_221),
.Y(n_291)
);

AOI22xp33_ASAP7_75t_L g273 ( 
.A1(n_209),
.A2(n_104),
.B1(n_196),
.B2(n_135),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_233),
.Y(n_274)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_274),
.Y(n_308)
);

AO22x2_ASAP7_75t_L g275 ( 
.A1(n_224),
.A2(n_104),
.B1(n_135),
.B2(n_11),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_SL g276 ( 
.A(n_201),
.B(n_9),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_SL g286 ( 
.A(n_276),
.B(n_205),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_SL g277 ( 
.A(n_210),
.B(n_9),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_277),
.B(n_280),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_235),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_278),
.Y(n_287)
);

HB1xp67_ASAP7_75t_L g279 ( 
.A(n_208),
.Y(n_279)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_279),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_SL g280 ( 
.A(n_210),
.B(n_10),
.Y(n_280)
);

AOI22xp33_ASAP7_75t_SL g281 ( 
.A1(n_205),
.A2(n_13),
.B1(n_135),
.B2(n_240),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_SL g332 ( 
.A(n_286),
.B(n_292),
.Y(n_332)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_291),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_270),
.B(n_221),
.Y(n_292)
);

XOR2xp5_ASAP7_75t_L g293 ( 
.A(n_245),
.B(n_237),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_293),
.B(n_300),
.C(n_267),
.Y(n_318)
);

OAI21xp33_ASAP7_75t_SL g295 ( 
.A1(n_256),
.A2(n_228),
.B(n_229),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g325 ( 
.A1(n_295),
.A2(n_305),
.B1(n_314),
.B2(n_266),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g296 ( 
.A(n_264),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_296),
.Y(n_320)
);

NOR2x1_ASAP7_75t_L g297 ( 
.A(n_265),
.B(n_200),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_297),
.B(n_302),
.Y(n_346)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_257),
.B(n_240),
.C(n_207),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_L g305 ( 
.A1(n_253),
.A2(n_236),
.B1(n_235),
.B2(n_222),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_249),
.B(n_221),
.Y(n_306)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_306),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_249),
.B(n_221),
.Y(n_307)
);

CKINVDCx16_ASAP7_75t_R g319 ( 
.A(n_307),
.Y(n_319)
);

INVxp67_ASAP7_75t_L g334 ( 
.A(n_309),
.Y(n_334)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_252),
.Y(n_311)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_311),
.Y(n_322)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_269),
.Y(n_312)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_312),
.Y(n_340)
);

NAND3xp33_ASAP7_75t_L g313 ( 
.A(n_277),
.B(n_225),
.C(n_211),
.Y(n_313)
);

NAND3xp33_ASAP7_75t_L g333 ( 
.A(n_313),
.B(n_280),
.C(n_243),
.Y(n_333)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_274),
.Y(n_317)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_317),
.Y(n_348)
);

XNOR2xp5_ASAP7_75t_SL g359 ( 
.A(n_318),
.B(n_344),
.Y(n_359)
);

HB1xp67_ASAP7_75t_L g321 ( 
.A(n_303),
.Y(n_321)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_321),
.Y(n_353)
);

XOR2xp5_ASAP7_75t_L g323 ( 
.A(n_315),
.B(n_260),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g351 ( 
.A(n_323),
.B(n_331),
.C(n_342),
.Y(n_351)
);

INVx1_ASAP7_75t_SL g324 ( 
.A(n_294),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_324),
.B(n_339),
.Y(n_352)
);

OAI22xp5_ASAP7_75t_L g354 ( 
.A1(n_325),
.A2(n_338),
.B1(n_341),
.B2(n_301),
.Y(n_354)
);

CKINVDCx20_ASAP7_75t_R g327 ( 
.A(n_282),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g349 ( 
.A(n_327),
.B(n_333),
.Y(n_349)
);

AOI21xp5_ASAP7_75t_L g328 ( 
.A1(n_294),
.A2(n_262),
.B(n_266),
.Y(n_328)
);

AOI21xp5_ASAP7_75t_L g360 ( 
.A1(n_328),
.A2(n_330),
.B(n_336),
.Y(n_360)
);

A2O1A1O1Ixp25_ASAP7_75t_L g329 ( 
.A1(n_285),
.A2(n_246),
.B(n_255),
.C(n_248),
.D(n_250),
.Y(n_329)
);

A2O1A1O1Ixp25_ASAP7_75t_L g372 ( 
.A1(n_329),
.A2(n_316),
.B(n_311),
.C(n_298),
.D(n_288),
.Y(n_372)
);

OAI21xp5_ASAP7_75t_SL g330 ( 
.A1(n_294),
.A2(n_251),
.B(n_265),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_315),
.B(n_246),
.C(n_264),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g335 ( 
.A(n_282),
.Y(n_335)
);

NAND3xp33_ASAP7_75t_L g373 ( 
.A(n_335),
.B(n_345),
.C(n_275),
.Y(n_373)
);

AOI21xp5_ASAP7_75t_L g336 ( 
.A1(n_304),
.A2(n_251),
.B(n_253),
.Y(n_336)
);

OAI22xp5_ASAP7_75t_L g337 ( 
.A1(n_287),
.A2(n_254),
.B1(n_278),
.B2(n_271),
.Y(n_337)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_337),
.Y(n_357)
);

AOI22xp5_ASAP7_75t_L g338 ( 
.A1(n_297),
.A2(n_305),
.B1(n_314),
.B2(n_293),
.Y(n_338)
);

INVxp67_ASAP7_75t_L g339 ( 
.A(n_309),
.Y(n_339)
);

AOI22xp5_ASAP7_75t_L g341 ( 
.A1(n_297),
.A2(n_254),
.B1(n_248),
.B2(n_264),
.Y(n_341)
);

XOR2xp5_ASAP7_75t_L g342 ( 
.A(n_290),
.B(n_248),
.Y(n_342)
);

XNOR2xp5_ASAP7_75t_SL g344 ( 
.A(n_290),
.B(n_276),
.Y(n_344)
);

OAI21xp33_ASAP7_75t_L g345 ( 
.A1(n_287),
.A2(n_275),
.B(n_261),
.Y(n_345)
);

INVx2_ASAP7_75t_L g347 ( 
.A(n_303),
.Y(n_347)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_347),
.Y(n_365)
);

AOI22xp5_ASAP7_75t_L g350 ( 
.A1(n_342),
.A2(n_296),
.B1(n_301),
.B2(n_284),
.Y(n_350)
);

AOI22xp5_ASAP7_75t_L g386 ( 
.A1(n_350),
.A2(n_354),
.B1(n_362),
.B2(n_375),
.Y(n_386)
);

MAJIxp5_ASAP7_75t_L g355 ( 
.A(n_318),
.B(n_300),
.C(n_289),
.Y(n_355)
);

MAJIxp5_ASAP7_75t_L g378 ( 
.A(n_355),
.B(n_364),
.C(n_371),
.Y(n_378)
);

OAI22xp5_ASAP7_75t_L g356 ( 
.A1(n_319),
.A2(n_284),
.B1(n_299),
.B2(n_285),
.Y(n_356)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_356),
.Y(n_376)
);

OR2x2_ASAP7_75t_L g358 ( 
.A(n_320),
.B(n_299),
.Y(n_358)
);

CKINVDCx20_ASAP7_75t_R g392 ( 
.A(n_358),
.Y(n_392)
);

CKINVDCx20_ASAP7_75t_R g361 ( 
.A(n_332),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_361),
.B(n_369),
.Y(n_382)
);

AOI22xp5_ASAP7_75t_L g362 ( 
.A1(n_334),
.A2(n_304),
.B1(n_302),
.B2(n_275),
.Y(n_362)
);

XNOR2xp5_ASAP7_75t_L g363 ( 
.A(n_323),
.B(n_289),
.Y(n_363)
);

XNOR2xp5_ASAP7_75t_L g379 ( 
.A(n_363),
.B(n_374),
.Y(n_379)
);

MAJIxp5_ASAP7_75t_L g364 ( 
.A(n_331),
.B(n_283),
.C(n_310),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_343),
.Y(n_366)
);

CKINVDCx14_ASAP7_75t_R g388 ( 
.A(n_366),
.Y(n_388)
);

OAI22xp5_ASAP7_75t_L g367 ( 
.A1(n_326),
.A2(n_286),
.B1(n_316),
.B2(n_312),
.Y(n_367)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_367),
.Y(n_380)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_322),
.Y(n_368)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_368),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_346),
.B(n_317),
.Y(n_369)
);

INVxp67_ASAP7_75t_L g370 ( 
.A(n_341),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_370),
.B(n_373),
.Y(n_383)
);

MAJIxp5_ASAP7_75t_L g371 ( 
.A(n_334),
.B(n_310),
.C(n_283),
.Y(n_371)
);

XOR2xp5_ASAP7_75t_L g381 ( 
.A(n_372),
.B(n_329),
.Y(n_381)
);

XNOR2xp5_ASAP7_75t_L g374 ( 
.A(n_344),
.B(n_298),
.Y(n_374)
);

AOI22xp5_ASAP7_75t_L g375 ( 
.A1(n_339),
.A2(n_275),
.B1(n_288),
.B2(n_308),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_L g377 ( 
.A(n_366),
.B(n_231),
.Y(n_377)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_377),
.Y(n_404)
);

XNOR2xp5_ASAP7_75t_SL g399 ( 
.A(n_381),
.B(n_350),
.Y(n_399)
);

MAJIxp5_ASAP7_75t_L g384 ( 
.A(n_364),
.B(n_338),
.C(n_324),
.Y(n_384)
);

MAJIxp5_ASAP7_75t_L g401 ( 
.A(n_384),
.B(n_391),
.C(n_393),
.Y(n_401)
);

XNOR2xp5_ASAP7_75t_L g387 ( 
.A(n_351),
.B(n_328),
.Y(n_387)
);

XNOR2xp5_ASAP7_75t_L g405 ( 
.A(n_387),
.B(n_389),
.Y(n_405)
);

XNOR2xp5_ASAP7_75t_L g389 ( 
.A(n_351),
.B(n_336),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_358),
.B(n_348),
.Y(n_390)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_390),
.Y(n_411)
);

MAJIxp5_ASAP7_75t_L g391 ( 
.A(n_355),
.B(n_325),
.C(n_330),
.Y(n_391)
);

MAJIxp5_ASAP7_75t_L g393 ( 
.A(n_359),
.B(n_346),
.C(n_348),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_SL g394 ( 
.A(n_349),
.B(n_340),
.Y(n_394)
);

XNOR2xp5_ASAP7_75t_L g408 ( 
.A(n_394),
.B(n_395),
.Y(n_408)
);

XNOR2xp5_ASAP7_75t_L g395 ( 
.A(n_359),
.B(n_340),
.Y(n_395)
);

NOR2xp33_ASAP7_75t_L g396 ( 
.A(n_371),
.B(n_374),
.Y(n_396)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_396),
.Y(n_416)
);

AO21x1_ASAP7_75t_L g397 ( 
.A1(n_369),
.A2(n_322),
.B(n_308),
.Y(n_397)
);

XNOR2xp5_ASAP7_75t_L g410 ( 
.A(n_397),
.B(n_352),
.Y(n_410)
);

MAJIxp5_ASAP7_75t_L g398 ( 
.A(n_363),
.B(n_347),
.C(n_231),
.Y(n_398)
);

MAJIxp5_ASAP7_75t_L g414 ( 
.A(n_398),
.B(n_211),
.C(n_241),
.Y(n_414)
);

XNOR2xp5_ASAP7_75t_L g420 ( 
.A(n_399),
.B(n_400),
.Y(n_420)
);

XOR2xp5_ASAP7_75t_L g400 ( 
.A(n_387),
.B(n_360),
.Y(n_400)
);

NOR2xp67_ASAP7_75t_SL g402 ( 
.A(n_389),
.B(n_360),
.Y(n_402)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_402),
.Y(n_419)
);

AOI22xp5_ASAP7_75t_L g403 ( 
.A1(n_380),
.A2(n_357),
.B1(n_370),
.B2(n_353),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_SL g421 ( 
.A(n_403),
.B(n_409),
.Y(n_421)
);

AOI22xp5_ASAP7_75t_SL g406 ( 
.A1(n_376),
.A2(n_362),
.B1(n_372),
.B2(n_375),
.Y(n_406)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_406),
.Y(n_422)
);

HB1xp67_ASAP7_75t_L g407 ( 
.A(n_382),
.Y(n_407)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_407),
.Y(n_424)
);

CKINVDCx20_ASAP7_75t_R g409 ( 
.A(n_392),
.Y(n_409)
);

NOR2xp33_ASAP7_75t_L g428 ( 
.A(n_410),
.B(n_413),
.Y(n_428)
);

MAJx2_ASAP7_75t_L g412 ( 
.A(n_393),
.B(n_352),
.C(n_365),
.Y(n_412)
);

MAJIxp5_ASAP7_75t_L g429 ( 
.A(n_412),
.B(n_414),
.C(n_398),
.Y(n_429)
);

AOI22xp5_ASAP7_75t_L g413 ( 
.A1(n_388),
.A2(n_259),
.B1(n_236),
.B2(n_239),
.Y(n_413)
);

NOR2xp33_ASAP7_75t_SL g415 ( 
.A(n_378),
.B(n_239),
.Y(n_415)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_415),
.Y(n_426)
);

NAND4xp25_ASAP7_75t_L g417 ( 
.A(n_411),
.B(n_386),
.C(n_383),
.D(n_381),
.Y(n_417)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_417),
.Y(n_432)
);

OAI21xp5_ASAP7_75t_SL g418 ( 
.A1(n_406),
.A2(n_391),
.B(n_384),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_SL g439 ( 
.A(n_418),
.B(n_427),
.Y(n_439)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_404),
.Y(n_423)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_423),
.Y(n_435)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_412),
.Y(n_425)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_425),
.Y(n_436)
);

AOI21xp5_ASAP7_75t_L g427 ( 
.A1(n_400),
.A2(n_386),
.B(n_397),
.Y(n_427)
);

XNOR2xp5_ASAP7_75t_L g434 ( 
.A(n_429),
.B(n_401),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_414),
.B(n_385),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g441 ( 
.A(n_430),
.B(n_379),
.Y(n_441)
);

AOI21x1_ASAP7_75t_L g431 ( 
.A1(n_421),
.A2(n_399),
.B(n_408),
.Y(n_431)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_431),
.Y(n_444)
);

MAJIxp5_ASAP7_75t_L g433 ( 
.A(n_429),
.B(n_378),
.C(n_401),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_SL g453 ( 
.A(n_433),
.B(n_434),
.Y(n_453)
);

OR2x2_ASAP7_75t_L g437 ( 
.A(n_428),
.B(n_416),
.Y(n_437)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_437),
.Y(n_450)
);

AOI22xp5_ASAP7_75t_SL g438 ( 
.A1(n_422),
.A2(n_405),
.B1(n_395),
.B2(n_379),
.Y(n_438)
);

XNOR2xp5_ASAP7_75t_L g445 ( 
.A(n_438),
.B(n_418),
.Y(n_445)
);

XOR2xp5_ASAP7_75t_L g440 ( 
.A(n_420),
.B(n_405),
.Y(n_440)
);

XOR2xp5_ASAP7_75t_L g451 ( 
.A(n_440),
.B(n_442),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_441),
.B(n_443),
.Y(n_447)
);

XOR2xp5_ASAP7_75t_L g442 ( 
.A(n_420),
.B(n_241),
.Y(n_442)
);

NOR2xp33_ASAP7_75t_SL g443 ( 
.A(n_423),
.B(n_233),
.Y(n_443)
);

NOR2xp33_ASAP7_75t_L g457 ( 
.A(n_445),
.B(n_13),
.Y(n_457)
);

OAI22xp5_ASAP7_75t_L g446 ( 
.A1(n_432),
.A2(n_425),
.B1(n_426),
.B2(n_422),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_446),
.B(n_448),
.Y(n_460)
);

OAI22xp5_ASAP7_75t_SL g448 ( 
.A1(n_439),
.A2(n_436),
.B1(n_419),
.B2(n_417),
.Y(n_448)
);

OAI21xp5_ASAP7_75t_SL g449 ( 
.A1(n_437),
.A2(n_427),
.B(n_430),
.Y(n_449)
);

AOI21xp5_ASAP7_75t_L g456 ( 
.A1(n_449),
.A2(n_440),
.B(n_220),
.Y(n_456)
);

AOI322xp5_ASAP7_75t_L g452 ( 
.A1(n_435),
.A2(n_13),
.A3(n_220),
.B1(n_222),
.B2(n_226),
.C1(n_424),
.C2(n_438),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_L g461 ( 
.A(n_452),
.B(n_448),
.Y(n_461)
);

NOR2xp67_ASAP7_75t_SL g454 ( 
.A(n_433),
.B(n_226),
.Y(n_454)
);

NOR2xp33_ASAP7_75t_SL g455 ( 
.A(n_454),
.B(n_442),
.Y(n_455)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_455),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_456),
.B(n_457),
.Y(n_462)
);

NOR2xp33_ASAP7_75t_L g458 ( 
.A(n_447),
.B(n_450),
.Y(n_458)
);

XNOR2xp5_ASAP7_75t_L g463 ( 
.A(n_458),
.B(n_459),
.Y(n_463)
);

OAI21x1_ASAP7_75t_L g459 ( 
.A1(n_453),
.A2(n_444),
.B(n_449),
.Y(n_459)
);

INVxp67_ASAP7_75t_L g464 ( 
.A(n_461),
.Y(n_464)
);

INVxp33_ASAP7_75t_L g466 ( 
.A(n_464),
.Y(n_466)
);

OAI31xp33_ASAP7_75t_L g469 ( 
.A1(n_466),
.A2(n_467),
.A3(n_468),
.B(n_456),
.Y(n_469)
);

XOR2xp5_ASAP7_75t_L g467 ( 
.A(n_463),
.B(n_445),
.Y(n_467)
);

XNOR2xp5_ASAP7_75t_L g468 ( 
.A(n_465),
.B(n_460),
.Y(n_468)
);

OAI21xp5_ASAP7_75t_SL g470 ( 
.A1(n_469),
.A2(n_462),
.B(n_451),
.Y(n_470)
);

XOR2xp5_ASAP7_75t_L g471 ( 
.A(n_470),
.B(n_451),
.Y(n_471)
);


endmodule