module fake_jpeg_1210_n_679 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_679);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_679;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_657;
wire n_27;
wire n_664;
wire n_365;
wire n_179;
wire n_620;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_678;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_417;
wire n_362;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_635;
wire n_517;
wire n_629;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_643;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_647;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_641;
wire n_48;
wire n_465;
wire n_638;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_623;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_637;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_672;
wire n_309;
wire n_624;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_596;
wire n_569;
wire n_400;
wire n_646;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_663;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_634;
wire n_23;
wire n_69;
wire n_658;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_666;
wire n_639;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_645;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_622;
wire n_463;
wire n_667;
wire n_92;
wire n_332;
wire n_640;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_653;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_626;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_668;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_642;
wire n_101;
wire n_226;
wire n_509;
wire n_644;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_656;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_649;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_615;
wire n_598;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_662;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_676;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_648;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_670;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_631;
wire n_433;
wire n_636;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_650;
wire n_218;
wire n_63;
wire n_652;
wire n_599;
wire n_239;
wire n_674;
wire n_243;
wire n_481;
wire n_628;
wire n_619;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_655;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_625;
wire n_147;
wire n_449;
wire n_627;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_659;
wire n_125;
wire n_661;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_673;
wire n_58;
wire n_41;
wire n_613;
wire n_630;
wire n_266;
wire n_548;
wire n_665;
wire n_72;
wire n_512;
wire n_654;
wire n_445;
wire n_443;
wire n_677;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_671;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_669;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_660;
wire n_373;
wire n_633;
wire n_112;
wire n_632;
wire n_616;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_651;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_675;
wire n_335;
wire n_120;
wire n_621;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_18),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_18),
.Y(n_22)
);

CKINVDCx16_ASAP7_75t_R g23 ( 
.A(n_4),
.Y(n_23)
);

INVx6_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_18),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_18),
.Y(n_28)
);

CKINVDCx14_ASAP7_75t_R g29 ( 
.A(n_9),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

BUFx12_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

INVx1_ASAP7_75t_SL g33 ( 
.A(n_0),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_4),
.Y(n_34)
);

BUFx2_ASAP7_75t_L g35 ( 
.A(n_8),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_6),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_6),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_1),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_13),
.Y(n_39)
);

INVx11_ASAP7_75t_L g40 ( 
.A(n_14),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_2),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_7),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_4),
.Y(n_43)
);

BUFx5_ASAP7_75t_L g44 ( 
.A(n_9),
.Y(n_44)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_1),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_6),
.Y(n_46)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_2),
.Y(n_47)
);

BUFx8_ASAP7_75t_L g48 ( 
.A(n_2),
.Y(n_48)
);

BUFx2_ASAP7_75t_L g49 ( 
.A(n_13),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_14),
.Y(n_50)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_9),
.Y(n_51)
);

BUFx5_ASAP7_75t_L g52 ( 
.A(n_8),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_2),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_4),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_13),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_9),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_0),
.Y(n_57)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_12),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_5),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_28),
.B(n_55),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_60),
.B(n_82),
.Y(n_139)
);

BUFx2_ASAP7_75t_L g61 ( 
.A(n_35),
.Y(n_61)
);

INVx2_ASAP7_75t_SL g217 ( 
.A(n_61),
.Y(n_217)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_50),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_62),
.Y(n_134)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_34),
.Y(n_63)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_63),
.Y(n_136)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_34),
.Y(n_64)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_64),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_50),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g150 ( 
.A(n_65),
.Y(n_150)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_50),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g173 ( 
.A(n_66),
.Y(n_173)
);

BUFx4f_ASAP7_75t_L g67 ( 
.A(n_48),
.Y(n_67)
);

INVx1_ASAP7_75t_SL g185 ( 
.A(n_67),
.Y(n_185)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_50),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g183 ( 
.A(n_68),
.Y(n_183)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_34),
.Y(n_69)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_69),
.Y(n_143)
);

CKINVDCx9p33_ASAP7_75t_R g70 ( 
.A(n_48),
.Y(n_70)
);

INVx4_ASAP7_75t_SL g155 ( 
.A(n_70),
.Y(n_155)
);

CKINVDCx6p67_ASAP7_75t_R g71 ( 
.A(n_48),
.Y(n_71)
);

INVx1_ASAP7_75t_SL g188 ( 
.A(n_71),
.Y(n_188)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_51),
.Y(n_72)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_72),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_31),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g192 ( 
.A(n_73),
.Y(n_192)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_31),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g195 ( 
.A(n_74),
.Y(n_195)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_49),
.Y(n_75)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_75),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_31),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g208 ( 
.A(n_76),
.Y(n_208)
);

INVx5_ASAP7_75t_L g77 ( 
.A(n_53),
.Y(n_77)
);

BUFx3_ASAP7_75t_L g135 ( 
.A(n_77),
.Y(n_135)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_51),
.Y(n_78)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_78),
.Y(n_163)
);

BUFx5_ASAP7_75t_L g79 ( 
.A(n_48),
.Y(n_79)
);

INVx4_ASAP7_75t_L g141 ( 
.A(n_79),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_31),
.Y(n_80)
);

INVx6_ASAP7_75t_L g170 ( 
.A(n_80),
.Y(n_170)
);

INVx6_ASAP7_75t_L g81 ( 
.A(n_42),
.Y(n_81)
);

BUFx2_ASAP7_75t_L g148 ( 
.A(n_81),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_28),
.B(n_19),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_55),
.B(n_19),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_83),
.B(n_96),
.Y(n_147)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_45),
.Y(n_84)
);

INVx3_ASAP7_75t_L g137 ( 
.A(n_84),
.Y(n_137)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_49),
.Y(n_85)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_85),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_59),
.Y(n_86)
);

INVx8_ASAP7_75t_L g158 ( 
.A(n_86),
.Y(n_158)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_45),
.Y(n_87)
);

INVx3_ASAP7_75t_L g138 ( 
.A(n_87),
.Y(n_138)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_49),
.Y(n_88)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_88),
.Y(n_161)
);

BUFx3_ASAP7_75t_L g89 ( 
.A(n_21),
.Y(n_89)
);

INVx5_ASAP7_75t_L g153 ( 
.A(n_89),
.Y(n_153)
);

BUFx12f_ASAP7_75t_L g90 ( 
.A(n_48),
.Y(n_90)
);

INVx5_ASAP7_75t_L g146 ( 
.A(n_90),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_SL g91 ( 
.A(n_36),
.B(n_19),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_91),
.B(n_95),
.Y(n_159)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_45),
.Y(n_92)
);

INVx3_ASAP7_75t_L g144 ( 
.A(n_92),
.Y(n_144)
);

INVx6_ASAP7_75t_L g93 ( 
.A(n_42),
.Y(n_93)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_93),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_59),
.Y(n_94)
);

INVx5_ASAP7_75t_L g174 ( 
.A(n_94),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_SL g95 ( 
.A(n_36),
.B(n_19),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_37),
.B(n_17),
.Y(n_96)
);

BUFx12f_ASAP7_75t_L g97 ( 
.A(n_32),
.Y(n_97)
);

INVx5_ASAP7_75t_L g179 ( 
.A(n_97),
.Y(n_179)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_53),
.Y(n_98)
);

INVx3_ASAP7_75t_L g151 ( 
.A(n_98),
.Y(n_151)
);

INVx6_ASAP7_75t_L g99 ( 
.A(n_42),
.Y(n_99)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_99),
.Y(n_169)
);

INVx4_ASAP7_75t_SL g100 ( 
.A(n_58),
.Y(n_100)
);

INVx6_ASAP7_75t_SL g224 ( 
.A(n_100),
.Y(n_224)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_42),
.Y(n_101)
);

INVx5_ASAP7_75t_L g197 ( 
.A(n_101),
.Y(n_197)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_59),
.Y(n_102)
);

INVx4_ASAP7_75t_L g149 ( 
.A(n_102),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_23),
.B(n_17),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_103),
.B(n_111),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_59),
.Y(n_104)
);

INVx4_ASAP7_75t_L g162 ( 
.A(n_104),
.Y(n_162)
);

BUFx4f_ASAP7_75t_SL g105 ( 
.A(n_58),
.Y(n_105)
);

BUFx12_ASAP7_75t_L g156 ( 
.A(n_105),
.Y(n_156)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_51),
.Y(n_106)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_106),
.Y(n_178)
);

INVx2_ASAP7_75t_SL g107 ( 
.A(n_35),
.Y(n_107)
);

INVx4_ASAP7_75t_L g181 ( 
.A(n_107),
.Y(n_181)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_35),
.Y(n_108)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_108),
.Y(n_191)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_35),
.Y(n_109)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_109),
.Y(n_199)
);

CKINVDCx16_ASAP7_75t_R g110 ( 
.A(n_49),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_110),
.B(n_129),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_23),
.B(n_17),
.Y(n_111)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_24),
.Y(n_112)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_112),
.Y(n_172)
);

BUFx5_ASAP7_75t_L g113 ( 
.A(n_44),
.Y(n_113)
);

INVx4_ASAP7_75t_L g200 ( 
.A(n_113),
.Y(n_200)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_47),
.Y(n_114)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_114),
.Y(n_202)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_57),
.Y(n_115)
);

INVx4_ASAP7_75t_L g204 ( 
.A(n_115),
.Y(n_204)
);

INVx5_ASAP7_75t_L g116 ( 
.A(n_53),
.Y(n_116)
);

INVx4_ASAP7_75t_L g205 ( 
.A(n_116),
.Y(n_205)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_47),
.Y(n_117)
);

INVx3_ASAP7_75t_L g194 ( 
.A(n_117),
.Y(n_194)
);

BUFx12_ASAP7_75t_L g118 ( 
.A(n_58),
.Y(n_118)
);

BUFx12_ASAP7_75t_L g207 ( 
.A(n_118),
.Y(n_207)
);

INVx4_ASAP7_75t_L g119 ( 
.A(n_44),
.Y(n_119)
);

INVx3_ASAP7_75t_L g196 ( 
.A(n_119),
.Y(n_196)
);

BUFx5_ASAP7_75t_L g120 ( 
.A(n_44),
.Y(n_120)
);

INVx4_ASAP7_75t_L g211 ( 
.A(n_120),
.Y(n_211)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_47),
.Y(n_121)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_121),
.Y(n_215)
);

INVx11_ASAP7_75t_L g122 ( 
.A(n_47),
.Y(n_122)
);

INVx11_ASAP7_75t_L g164 ( 
.A(n_122),
.Y(n_164)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_21),
.Y(n_123)
);

INVx3_ASAP7_75t_L g212 ( 
.A(n_123),
.Y(n_212)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_57),
.Y(n_124)
);

INVx4_ASAP7_75t_L g218 ( 
.A(n_124),
.Y(n_218)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_47),
.Y(n_125)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_125),
.Y(n_220)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_21),
.Y(n_126)
);

INVx3_ASAP7_75t_L g226 ( 
.A(n_126),
.Y(n_226)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_57),
.Y(n_127)
);

INVx4_ASAP7_75t_L g225 ( 
.A(n_127),
.Y(n_225)
);

INVx3_ASAP7_75t_L g128 ( 
.A(n_47),
.Y(n_128)
);

HB1xp67_ASAP7_75t_L g152 ( 
.A(n_128),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_SL g129 ( 
.A(n_37),
.B(n_17),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_57),
.Y(n_130)
);

INVx4_ASAP7_75t_L g222 ( 
.A(n_130),
.Y(n_222)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_24),
.Y(n_131)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_131),
.Y(n_177)
);

AOI21xp33_ASAP7_75t_L g132 ( 
.A1(n_71),
.A2(n_22),
.B(n_39),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_SL g270 ( 
.A(n_132),
.B(n_175),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_84),
.B(n_33),
.C(n_22),
.Y(n_133)
);

AND2x2_ASAP7_75t_L g230 ( 
.A(n_133),
.B(n_184),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_66),
.A2(n_24),
.B1(n_46),
.B2(n_43),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g253 ( 
.A1(n_165),
.A2(n_166),
.B1(n_167),
.B2(n_171),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_62),
.A2(n_22),
.B1(n_26),
.B2(n_39),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_81),
.A2(n_24),
.B1(n_46),
.B2(n_43),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_93),
.A2(n_46),
.B1(n_43),
.B2(n_58),
.Y(n_171)
);

AND2x2_ASAP7_75t_L g175 ( 
.A(n_107),
.B(n_33),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_97),
.B(n_33),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_SL g275 ( 
.A(n_176),
.B(n_180),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_97),
.B(n_58),
.Y(n_180)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_61),
.Y(n_182)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_182),
.Y(n_237)
);

NAND2xp33_ASAP7_75t_SL g184 ( 
.A(n_71),
.B(n_29),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_92),
.B(n_29),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_186),
.B(n_193),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_105),
.B(n_58),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_187),
.B(n_190),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_65),
.A2(n_26),
.B1(n_39),
.B2(n_38),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_L g280 ( 
.A1(n_189),
.A2(n_198),
.B1(n_214),
.B2(n_221),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_99),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_87),
.B(n_26),
.Y(n_193)
);

AOI22xp33_ASAP7_75t_L g198 ( 
.A1(n_73),
.A2(n_40),
.B1(n_54),
.B2(n_30),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_100),
.B(n_30),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_201),
.B(n_210),
.Y(n_260)
);

AOI22xp33_ASAP7_75t_SL g203 ( 
.A1(n_67),
.A2(n_40),
.B1(n_54),
.B2(n_20),
.Y(n_203)
);

OA22x2_ASAP7_75t_L g297 ( 
.A1(n_203),
.A2(n_32),
.B1(n_3),
.B2(n_5),
.Y(n_297)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_117),
.Y(n_206)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_206),
.Y(n_246)
);

OAI22xp33_ASAP7_75t_SL g209 ( 
.A1(n_74),
.A2(n_40),
.B1(n_56),
.B2(n_38),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_209),
.A2(n_213),
.B1(n_32),
.B2(n_2),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_89),
.B(n_56),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_68),
.A2(n_56),
.B1(n_54),
.B2(n_25),
.Y(n_213)
);

AOI22xp33_ASAP7_75t_L g214 ( 
.A1(n_76),
.A2(n_41),
.B1(n_38),
.B2(n_30),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_77),
.B(n_20),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_216),
.B(n_90),
.Y(n_229)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_116),
.Y(n_219)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_219),
.Y(n_256)
);

AOI22xp33_ASAP7_75t_L g221 ( 
.A1(n_80),
.A2(n_41),
.B1(n_27),
.B2(n_25),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_90),
.B(n_20),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_223),
.B(n_16),
.Y(n_276)
);

INVx4_ASAP7_75t_L g227 ( 
.A(n_217),
.Y(n_227)
);

INVx4_ASAP7_75t_L g347 ( 
.A(n_227),
.Y(n_347)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_168),
.Y(n_228)
);

INVx2_ASAP7_75t_L g313 ( 
.A(n_228),
.Y(n_313)
);

AND2x2_ASAP7_75t_L g342 ( 
.A(n_229),
.B(n_282),
.Y(n_342)
);

INVx3_ASAP7_75t_L g232 ( 
.A(n_181),
.Y(n_232)
);

INVx3_ASAP7_75t_L g351 ( 
.A(n_232),
.Y(n_351)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_169),
.Y(n_233)
);

INVx2_ASAP7_75t_L g314 ( 
.A(n_233),
.Y(n_314)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_224),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_SL g322 ( 
.A(n_234),
.B(n_249),
.Y(n_322)
);

AND2x2_ASAP7_75t_L g235 ( 
.A(n_175),
.B(n_181),
.Y(n_235)
);

CKINVDCx14_ASAP7_75t_R g357 ( 
.A(n_235),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_147),
.B(n_25),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_236),
.B(n_254),
.Y(n_330)
);

INVx8_ASAP7_75t_L g238 ( 
.A(n_192),
.Y(n_238)
);

INVx5_ASAP7_75t_L g358 ( 
.A(n_238),
.Y(n_358)
);

BUFx2_ASAP7_75t_L g239 ( 
.A(n_217),
.Y(n_239)
);

HB1xp67_ASAP7_75t_L g335 ( 
.A(n_239),
.Y(n_335)
);

BUFx8_ASAP7_75t_L g240 ( 
.A(n_155),
.Y(n_240)
);

INVxp67_ASAP7_75t_L g318 ( 
.A(n_240),
.Y(n_318)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_172),
.Y(n_241)
);

INVx2_ASAP7_75t_L g315 ( 
.A(n_241),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_198),
.A2(n_130),
.B1(n_127),
.B2(n_124),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g326 ( 
.A1(n_242),
.A2(n_290),
.B1(n_195),
.B2(n_192),
.Y(n_326)
);

INVx3_ASAP7_75t_L g243 ( 
.A(n_185),
.Y(n_243)
);

INVx2_ASAP7_75t_L g320 ( 
.A(n_243),
.Y(n_320)
);

AOI22xp33_ASAP7_75t_SL g245 ( 
.A1(n_188),
.A2(n_119),
.B1(n_27),
.B2(n_41),
.Y(n_245)
);

INVxp67_ASAP7_75t_L g362 ( 
.A(n_245),
.Y(n_362)
);

AOI22xp33_ASAP7_75t_SL g247 ( 
.A1(n_188),
.A2(n_27),
.B1(n_122),
.B2(n_115),
.Y(n_247)
);

INVxp67_ASAP7_75t_L g367 ( 
.A(n_247),
.Y(n_367)
);

AOI22xp33_ASAP7_75t_SL g248 ( 
.A1(n_155),
.A2(n_94),
.B1(n_104),
.B2(n_102),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_L g340 ( 
.A1(n_248),
.A2(n_289),
.B1(n_292),
.B2(n_306),
.Y(n_340)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_152),
.Y(n_249)
);

INVx4_ASAP7_75t_L g250 ( 
.A(n_146),
.Y(n_250)
);

INVx2_ASAP7_75t_L g323 ( 
.A(n_250),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_152),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_SL g327 ( 
.A(n_251),
.B(n_262),
.Y(n_327)
);

INVx3_ASAP7_75t_L g252 ( 
.A(n_185),
.Y(n_252)
);

INVx2_ASAP7_75t_L g332 ( 
.A(n_252),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_160),
.B(n_136),
.Y(n_254)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_177),
.Y(n_255)
);

INVx2_ASAP7_75t_L g343 ( 
.A(n_255),
.Y(n_343)
);

BUFx2_ASAP7_75t_SL g257 ( 
.A(n_141),
.Y(n_257)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_257),
.Y(n_311)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_140),
.Y(n_258)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_258),
.Y(n_316)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_143),
.Y(n_259)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_259),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_154),
.B(n_101),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_261),
.B(n_281),
.Y(n_338)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_148),
.Y(n_262)
);

HB1xp67_ASAP7_75t_L g263 ( 
.A(n_194),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g355 ( 
.A(n_263),
.Y(n_355)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_148),
.Y(n_264)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_264),
.Y(n_321)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_142),
.Y(n_265)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_265),
.Y(n_334)
);

AO22x1_ASAP7_75t_L g266 ( 
.A1(n_164),
.A2(n_86),
.B1(n_118),
.B2(n_52),
.Y(n_266)
);

OAI21xp5_ASAP7_75t_L g324 ( 
.A1(n_266),
.A2(n_301),
.B(n_305),
.Y(n_324)
);

INVx3_ASAP7_75t_L g267 ( 
.A(n_205),
.Y(n_267)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_267),
.Y(n_336)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_145),
.Y(n_268)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_268),
.Y(n_339)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_151),
.Y(n_269)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_269),
.Y(n_350)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_202),
.Y(n_271)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_271),
.Y(n_356)
);

AOI21xp5_ASAP7_75t_L g272 ( 
.A1(n_209),
.A2(n_118),
.B(n_52),
.Y(n_272)
);

AOI21xp5_ASAP7_75t_L g312 ( 
.A1(n_272),
.A2(n_211),
.B(n_200),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_174),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_SL g344 ( 
.A(n_273),
.B(n_293),
.Y(n_344)
);

INVx6_ASAP7_75t_L g274 ( 
.A(n_134),
.Y(n_274)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_274),
.Y(n_368)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_276),
.B(n_284),
.Y(n_308)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_161),
.Y(n_277)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_277),
.Y(n_369)
);

INVx11_ASAP7_75t_L g278 ( 
.A(n_164),
.Y(n_278)
);

INVx6_ASAP7_75t_L g348 ( 
.A(n_278),
.Y(n_348)
);

BUFx16f_ASAP7_75t_L g279 ( 
.A(n_156),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g317 ( 
.A(n_279),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_215),
.B(n_0),
.Y(n_281)
);

INVx3_ASAP7_75t_L g282 ( 
.A(n_205),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_220),
.B(n_0),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_283),
.B(n_288),
.Y(n_353)
);

INVx6_ASAP7_75t_L g284 ( 
.A(n_134),
.Y(n_284)
);

BUFx2_ASAP7_75t_L g285 ( 
.A(n_153),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_285),
.B(n_286),
.Y(n_331)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_191),
.Y(n_286)
);

OAI22xp33_ASAP7_75t_SL g287 ( 
.A1(n_214),
.A2(n_52),
.B1(n_32),
.B2(n_16),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_SL g329 ( 
.A1(n_287),
.A2(n_296),
.B1(n_297),
.B2(n_302),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_199),
.B(n_1),
.Y(n_288)
);

AOI22xp33_ASAP7_75t_L g289 ( 
.A1(n_157),
.A2(n_178),
.B1(n_163),
.B2(n_221),
.Y(n_289)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_212),
.Y(n_291)
);

OR2x2_ASAP7_75t_L g363 ( 
.A(n_291),
.B(n_295),
.Y(n_363)
);

AOI22xp33_ASAP7_75t_SL g292 ( 
.A1(n_141),
.A2(n_32),
.B1(n_16),
.B2(n_15),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_139),
.B(n_16),
.Y(n_293)
);

AND2x2_ASAP7_75t_L g294 ( 
.A(n_138),
.B(n_1),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g359 ( 
.A(n_294),
.B(n_300),
.C(n_303),
.Y(n_359)
);

INVx4_ASAP7_75t_L g295 ( 
.A(n_153),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_159),
.B(n_15),
.Y(n_296)
);

INVx3_ASAP7_75t_L g298 ( 
.A(n_135),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_298),
.B(n_299),
.Y(n_364)
);

HB1xp67_ASAP7_75t_L g299 ( 
.A(n_226),
.Y(n_299)
);

AND2x2_ASAP7_75t_L g300 ( 
.A(n_137),
.B(n_1),
.Y(n_300)
);

A2O1A1Ixp33_ASAP7_75t_L g301 ( 
.A1(n_156),
.A2(n_15),
.B(n_14),
.C(n_13),
.Y(n_301)
);

INVx3_ASAP7_75t_L g302 ( 
.A(n_135),
.Y(n_302)
);

AND2x2_ASAP7_75t_L g303 ( 
.A(n_144),
.B(n_3),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_196),
.B(n_3),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_L g361 ( 
.A(n_304),
.B(n_7),
.Y(n_361)
);

HB1xp67_ASAP7_75t_L g305 ( 
.A(n_179),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_L g306 ( 
.A1(n_173),
.A2(n_15),
.B1(n_14),
.B2(n_12),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_149),
.Y(n_307)
);

AOI22xp33_ASAP7_75t_L g325 ( 
.A1(n_307),
.A2(n_197),
.B1(n_222),
.B2(n_218),
.Y(n_325)
);

AO21x2_ASAP7_75t_SL g309 ( 
.A1(n_272),
.A2(n_203),
.B(n_156),
.Y(n_309)
);

INVx5_ASAP7_75t_L g395 ( 
.A(n_309),
.Y(n_395)
);

OAI22xp5_ASAP7_75t_SL g310 ( 
.A1(n_290),
.A2(n_173),
.B1(n_170),
.B2(n_225),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_L g379 ( 
.A1(n_310),
.A2(n_326),
.B1(n_333),
.B2(n_337),
.Y(n_379)
);

OAI21xp33_ASAP7_75t_SL g410 ( 
.A1(n_312),
.A2(n_279),
.B(n_252),
.Y(n_410)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_325),
.Y(n_377)
);

MAJx2_ASAP7_75t_L g328 ( 
.A(n_270),
.B(n_211),
.C(n_200),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g371 ( 
.A(n_328),
.B(n_366),
.C(n_301),
.Y(n_371)
);

OAI22xp33_ASAP7_75t_L g333 ( 
.A1(n_280),
.A2(n_170),
.B1(n_222),
.B2(n_218),
.Y(n_333)
);

OAI22xp33_ASAP7_75t_SL g337 ( 
.A1(n_260),
.A2(n_225),
.B1(n_204),
.B2(n_162),
.Y(n_337)
);

OAI22xp5_ASAP7_75t_L g341 ( 
.A1(n_231),
.A2(n_208),
.B1(n_195),
.B2(n_183),
.Y(n_341)
);

AOI22xp5_ASAP7_75t_L g404 ( 
.A1(n_341),
.A2(n_345),
.B1(n_346),
.B2(n_354),
.Y(n_404)
);

OAI22xp5_ASAP7_75t_L g345 ( 
.A1(n_261),
.A2(n_208),
.B1(n_183),
.B2(n_150),
.Y(n_345)
);

OAI22xp5_ASAP7_75t_SL g346 ( 
.A1(n_230),
.A2(n_204),
.B1(n_162),
.B2(n_149),
.Y(n_346)
);

AOI22xp5_ASAP7_75t_L g349 ( 
.A1(n_253),
.A2(n_150),
.B1(n_158),
.B2(n_207),
.Y(n_349)
);

OAI22xp5_ASAP7_75t_L g400 ( 
.A1(n_349),
.A2(n_278),
.B1(n_238),
.B2(n_264),
.Y(n_400)
);

AOI22xp33_ASAP7_75t_L g352 ( 
.A1(n_242),
.A2(n_158),
.B1(n_6),
.B2(n_7),
.Y(n_352)
);

OAI22xp33_ASAP7_75t_SL g373 ( 
.A1(n_352),
.A2(n_360),
.B1(n_306),
.B2(n_240),
.Y(n_373)
);

OAI22xp5_ASAP7_75t_SL g354 ( 
.A1(n_230),
.A2(n_207),
.B1(n_6),
.B2(n_7),
.Y(n_354)
);

AOI22xp33_ASAP7_75t_L g360 ( 
.A1(n_236),
.A2(n_5),
.B1(n_7),
.B2(n_8),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_SL g382 ( 
.A(n_361),
.B(n_294),
.Y(n_382)
);

MAJIxp5_ASAP7_75t_L g365 ( 
.A(n_230),
.B(n_207),
.C(n_12),
.Y(n_365)
);

MAJIxp5_ASAP7_75t_L g380 ( 
.A(n_365),
.B(n_235),
.C(n_303),
.Y(n_380)
);

XNOR2xp5_ASAP7_75t_L g366 ( 
.A(n_254),
.B(n_8),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_338),
.B(n_304),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_370),
.B(n_376),
.Y(n_421)
);

XNOR2xp5_ASAP7_75t_L g432 ( 
.A(n_371),
.B(n_380),
.Y(n_432)
);

CKINVDCx16_ASAP7_75t_R g372 ( 
.A(n_363),
.Y(n_372)
);

NOR2xp33_ASAP7_75t_L g435 ( 
.A(n_372),
.B(n_374),
.Y(n_435)
);

INVxp67_ASAP7_75t_L g420 ( 
.A(n_373),
.Y(n_420)
);

CKINVDCx20_ASAP7_75t_R g374 ( 
.A(n_322),
.Y(n_374)
);

INVx2_ASAP7_75t_L g375 ( 
.A(n_368),
.Y(n_375)
);

INVx2_ASAP7_75t_SL g450 ( 
.A(n_375),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_338),
.B(n_288),
.Y(n_376)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_364),
.Y(n_378)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_378),
.Y(n_443)
);

OAI22xp5_ASAP7_75t_SL g381 ( 
.A1(n_349),
.A2(n_229),
.B1(n_244),
.B2(n_281),
.Y(n_381)
);

AOI22xp5_ASAP7_75t_L g425 ( 
.A1(n_381),
.A2(n_387),
.B1(n_388),
.B2(n_392),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_382),
.B(n_343),
.Y(n_459)
);

MAJIxp5_ASAP7_75t_L g383 ( 
.A(n_328),
.B(n_235),
.C(n_246),
.Y(n_383)
);

MAJIxp5_ASAP7_75t_L g426 ( 
.A(n_383),
.B(n_365),
.C(n_359),
.Y(n_426)
);

AOI22xp33_ASAP7_75t_SL g384 ( 
.A1(n_367),
.A2(n_297),
.B1(n_266),
.B2(n_298),
.Y(n_384)
);

AOI22xp33_ASAP7_75t_SL g453 ( 
.A1(n_384),
.A2(n_408),
.B1(n_416),
.B2(n_347),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_353),
.B(n_283),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_385),
.B(n_386),
.Y(n_422)
);

CKINVDCx14_ASAP7_75t_R g386 ( 
.A(n_363),
.Y(n_386)
);

OAI22xp5_ASAP7_75t_SL g387 ( 
.A1(n_326),
.A2(n_303),
.B1(n_300),
.B2(n_294),
.Y(n_387)
);

OAI22xp5_ASAP7_75t_SL g388 ( 
.A1(n_329),
.A2(n_300),
.B1(n_297),
.B2(n_284),
.Y(n_388)
);

BUFx24_ASAP7_75t_SL g389 ( 
.A(n_344),
.Y(n_389)
);

INVxp67_ASAP7_75t_L g441 ( 
.A(n_389),
.Y(n_441)
);

OAI21xp5_ASAP7_75t_SL g390 ( 
.A1(n_312),
.A2(n_275),
.B(n_240),
.Y(n_390)
);

OAI21xp5_ASAP7_75t_SL g433 ( 
.A1(n_390),
.A2(n_396),
.B(n_417),
.Y(n_433)
);

CKINVDCx20_ASAP7_75t_R g391 ( 
.A(n_327),
.Y(n_391)
);

CKINVDCx14_ASAP7_75t_R g428 ( 
.A(n_391),
.Y(n_428)
);

OAI22xp5_ASAP7_75t_SL g392 ( 
.A1(n_329),
.A2(n_297),
.B1(n_274),
.B2(n_233),
.Y(n_392)
);

OAI22xp5_ASAP7_75t_SL g393 ( 
.A1(n_309),
.A2(n_228),
.B1(n_258),
.B2(n_259),
.Y(n_393)
);

AOI22xp5_ASAP7_75t_L g430 ( 
.A1(n_393),
.A2(n_398),
.B1(n_400),
.B2(n_318),
.Y(n_430)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_364),
.Y(n_394)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_394),
.Y(n_446)
);

OAI21xp5_ASAP7_75t_L g396 ( 
.A1(n_324),
.A2(n_266),
.B(n_255),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_334),
.Y(n_397)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_397),
.Y(n_451)
);

OAI22xp5_ASAP7_75t_SL g398 ( 
.A1(n_309),
.A2(n_269),
.B1(n_307),
.B2(n_271),
.Y(n_398)
);

INVxp67_ASAP7_75t_L g399 ( 
.A(n_331),
.Y(n_399)
);

INVxp67_ASAP7_75t_L g452 ( 
.A(n_399),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_353),
.B(n_286),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_401),
.B(n_402),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_330),
.B(n_241),
.Y(n_402)
);

NOR2xp33_ASAP7_75t_L g403 ( 
.A(n_355),
.B(n_237),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g438 ( 
.A(n_403),
.B(n_414),
.Y(n_438)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_334),
.Y(n_405)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_405),
.Y(n_454)
);

AOI22xp5_ASAP7_75t_L g406 ( 
.A1(n_324),
.A2(n_267),
.B1(n_282),
.B2(n_256),
.Y(n_406)
);

OAI22xp5_ASAP7_75t_L g439 ( 
.A1(n_406),
.A2(n_407),
.B1(n_415),
.B2(n_311),
.Y(n_439)
);

AOI22xp5_ASAP7_75t_L g407 ( 
.A1(n_333),
.A2(n_232),
.B1(n_302),
.B2(n_285),
.Y(n_407)
);

AOI22xp33_ASAP7_75t_SL g408 ( 
.A1(n_367),
.A2(n_362),
.B1(n_309),
.B2(n_340),
.Y(n_408)
);

AOI21xp5_ASAP7_75t_L g409 ( 
.A1(n_362),
.A2(n_279),
.B(n_250),
.Y(n_409)
);

OAI21xp5_ASAP7_75t_L g447 ( 
.A1(n_409),
.A2(n_418),
.B(n_317),
.Y(n_447)
);

OR2x2_ASAP7_75t_L g419 ( 
.A(n_410),
.B(n_396),
.Y(n_419)
);

INVxp67_ASAP7_75t_L g411 ( 
.A(n_342),
.Y(n_411)
);

CKINVDCx20_ASAP7_75t_R g423 ( 
.A(n_411),
.Y(n_423)
);

MAJx2_ASAP7_75t_L g412 ( 
.A(n_330),
.B(n_239),
.C(n_295),
.Y(n_412)
);

MAJIxp5_ASAP7_75t_L g437 ( 
.A(n_412),
.B(n_318),
.C(n_311),
.Y(n_437)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_339),
.Y(n_413)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_413),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_361),
.B(n_227),
.Y(n_414)
);

AOI22xp5_ASAP7_75t_L g415 ( 
.A1(n_310),
.A2(n_243),
.B1(n_9),
.B2(n_10),
.Y(n_415)
);

AOI22xp33_ASAP7_75t_SL g416 ( 
.A1(n_346),
.A2(n_8),
.B1(n_10),
.B2(n_11),
.Y(n_416)
);

A2O1A1O1Ixp25_ASAP7_75t_L g417 ( 
.A1(n_359),
.A2(n_10),
.B(n_11),
.C(n_342),
.D(n_357),
.Y(n_417)
);

OAI21xp5_ASAP7_75t_SL g418 ( 
.A1(n_342),
.A2(n_10),
.B(n_11),
.Y(n_418)
);

AOI21xp5_ASAP7_75t_L g472 ( 
.A1(n_419),
.A2(n_371),
.B(n_417),
.Y(n_472)
);

OAI22xp5_ASAP7_75t_SL g424 ( 
.A1(n_395),
.A2(n_308),
.B1(n_339),
.B2(n_369),
.Y(n_424)
);

AOI22xp5_ASAP7_75t_L g465 ( 
.A1(n_424),
.A2(n_427),
.B1(n_429),
.B2(n_431),
.Y(n_465)
);

MAJIxp5_ASAP7_75t_L g466 ( 
.A(n_426),
.B(n_448),
.C(n_456),
.Y(n_466)
);

OAI22xp5_ASAP7_75t_SL g427 ( 
.A1(n_395),
.A2(n_369),
.B1(n_368),
.B2(n_355),
.Y(n_427)
);

OAI22xp5_ASAP7_75t_SL g429 ( 
.A1(n_395),
.A2(n_354),
.B1(n_358),
.B2(n_356),
.Y(n_429)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_430),
.Y(n_464)
);

OAI22xp5_ASAP7_75t_SL g431 ( 
.A1(n_408),
.A2(n_358),
.B1(n_316),
.B2(n_356),
.Y(n_431)
);

XNOR2xp5_ASAP7_75t_L g436 ( 
.A(n_376),
.B(n_366),
.Y(n_436)
);

XNOR2xp5_ASAP7_75t_SL g495 ( 
.A(n_436),
.B(n_437),
.Y(n_495)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_439),
.Y(n_471)
);

OAI22xp5_ASAP7_75t_SL g440 ( 
.A1(n_378),
.A2(n_319),
.B1(n_316),
.B2(n_350),
.Y(n_440)
);

AOI22xp5_ASAP7_75t_L g494 ( 
.A1(n_440),
.A2(n_442),
.B1(n_375),
.B2(n_315),
.Y(n_494)
);

OAI22xp5_ASAP7_75t_SL g442 ( 
.A1(n_394),
.A2(n_319),
.B1(n_350),
.B2(n_336),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_L g444 ( 
.A(n_385),
.B(n_321),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g483 ( 
.A(n_444),
.B(n_455),
.Y(n_483)
);

CKINVDCx20_ASAP7_75t_R g445 ( 
.A(n_403),
.Y(n_445)
);

NOR2xp33_ASAP7_75t_L g460 ( 
.A(n_445),
.B(n_374),
.Y(n_460)
);

INVxp67_ASAP7_75t_L g490 ( 
.A(n_447),
.Y(n_490)
);

MAJIxp5_ASAP7_75t_L g448 ( 
.A(n_383),
.B(n_336),
.C(n_321),
.Y(n_448)
);

AOI22xp5_ASAP7_75t_L g449 ( 
.A1(n_388),
.A2(n_323),
.B1(n_351),
.B2(n_315),
.Y(n_449)
);

OAI22xp5_ASAP7_75t_SL g461 ( 
.A1(n_449),
.A2(n_379),
.B1(n_407),
.B2(n_404),
.Y(n_461)
);

INVxp67_ASAP7_75t_L g491 ( 
.A(n_453),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_L g455 ( 
.A(n_370),
.B(n_343),
.Y(n_455)
);

MAJIxp5_ASAP7_75t_L g456 ( 
.A(n_383),
.B(n_313),
.C(n_314),
.Y(n_456)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_397),
.Y(n_458)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_458),
.Y(n_485)
);

XNOR2xp5_ASAP7_75t_L g480 ( 
.A(n_459),
.B(n_418),
.Y(n_480)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_460),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_L g506 ( 
.A(n_461),
.B(n_463),
.Y(n_506)
);

OAI22xp5_ASAP7_75t_L g462 ( 
.A1(n_425),
.A2(n_384),
.B1(n_404),
.B2(n_379),
.Y(n_462)
);

OAI22xp5_ASAP7_75t_L g502 ( 
.A1(n_462),
.A2(n_467),
.B1(n_446),
.B2(n_428),
.Y(n_502)
);

INVx2_ASAP7_75t_SL g463 ( 
.A(n_450),
.Y(n_463)
);

OAI22xp5_ASAP7_75t_L g467 ( 
.A1(n_425),
.A2(n_401),
.B1(n_402),
.B2(n_406),
.Y(n_467)
);

OAI21xp5_ASAP7_75t_L g468 ( 
.A1(n_419),
.A2(n_390),
.B(n_410),
.Y(n_468)
);

OAI21xp5_ASAP7_75t_SL g499 ( 
.A1(n_468),
.A2(n_470),
.B(n_472),
.Y(n_499)
);

OAI22xp5_ASAP7_75t_SL g469 ( 
.A1(n_420),
.A2(n_392),
.B1(n_398),
.B2(n_393),
.Y(n_469)
);

AOI22xp5_ASAP7_75t_L g534 ( 
.A1(n_469),
.A2(n_481),
.B1(n_486),
.B2(n_450),
.Y(n_534)
);

OAI21xp5_ASAP7_75t_L g470 ( 
.A1(n_419),
.A2(n_386),
.B(n_409),
.Y(n_470)
);

XOR2xp5_ASAP7_75t_L g473 ( 
.A(n_432),
.B(n_412),
.Y(n_473)
);

MAJIxp5_ASAP7_75t_L g504 ( 
.A(n_473),
.B(n_482),
.C(n_487),
.Y(n_504)
);

OAI22xp5_ASAP7_75t_SL g474 ( 
.A1(n_453),
.A2(n_391),
.B1(n_412),
.B2(n_372),
.Y(n_474)
);

AOI22xp5_ASAP7_75t_L g509 ( 
.A1(n_474),
.A2(n_437),
.B1(n_447),
.B2(n_431),
.Y(n_509)
);

INVx2_ASAP7_75t_L g475 ( 
.A(n_450),
.Y(n_475)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_475),
.Y(n_505)
);

OA21x2_ASAP7_75t_L g476 ( 
.A1(n_427),
.A2(n_400),
.B(n_377),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_L g521 ( 
.A(n_476),
.B(n_479),
.Y(n_521)
);

NOR2xp33_ASAP7_75t_L g477 ( 
.A(n_445),
.B(n_413),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_SL g501 ( 
.A(n_477),
.B(n_493),
.Y(n_501)
);

CKINVDCx16_ASAP7_75t_R g478 ( 
.A(n_442),
.Y(n_478)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_478),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_SL g479 ( 
.A(n_428),
.B(n_381),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_L g523 ( 
.A(n_480),
.B(n_497),
.Y(n_523)
);

OAI22xp5_ASAP7_75t_SL g481 ( 
.A1(n_443),
.A2(n_415),
.B1(n_387),
.B2(n_377),
.Y(n_481)
);

MAJIxp5_ASAP7_75t_L g482 ( 
.A(n_432),
.B(n_380),
.C(n_414),
.Y(n_482)
);

OAI21xp5_ASAP7_75t_L g484 ( 
.A1(n_433),
.A2(n_417),
.B(n_405),
.Y(n_484)
);

OAI21xp5_ASAP7_75t_SL g510 ( 
.A1(n_484),
.A2(n_435),
.B(n_444),
.Y(n_510)
);

OAI22xp5_ASAP7_75t_SL g486 ( 
.A1(n_443),
.A2(n_446),
.B1(n_430),
.B2(n_434),
.Y(n_486)
);

XOR2xp5_ASAP7_75t_L g487 ( 
.A(n_426),
.B(n_380),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_451),
.Y(n_488)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_488),
.Y(n_517)
);

XNOR2xp5_ASAP7_75t_L g489 ( 
.A(n_426),
.B(n_382),
.Y(n_489)
);

XOR2xp5_ASAP7_75t_L g500 ( 
.A(n_489),
.B(n_448),
.Y(n_500)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_451),
.Y(n_492)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_492),
.Y(n_522)
);

INVxp67_ASAP7_75t_L g493 ( 
.A(n_433),
.Y(n_493)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_494),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_L g496 ( 
.A(n_421),
.B(n_373),
.Y(n_496)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_496),
.Y(n_529)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_454),
.Y(n_497)
);

XNOR2xp5_ASAP7_75t_L g498 ( 
.A(n_487),
.B(n_448),
.Y(n_498)
);

XOR2xp5_ASAP7_75t_L g550 ( 
.A(n_498),
.B(n_507),
.Y(n_550)
);

MAJIxp5_ASAP7_75t_L g543 ( 
.A(n_500),
.B(n_518),
.C(n_530),
.Y(n_543)
);

AOI22xp5_ASAP7_75t_L g548 ( 
.A1(n_502),
.A2(n_503),
.B1(n_481),
.B2(n_465),
.Y(n_548)
);

OAI22xp5_ASAP7_75t_SL g503 ( 
.A1(n_471),
.A2(n_434),
.B1(n_422),
.B2(n_421),
.Y(n_503)
);

XOR2xp5_ASAP7_75t_L g507 ( 
.A(n_489),
.B(n_495),
.Y(n_507)
);

OAI22xp5_ASAP7_75t_L g508 ( 
.A1(n_460),
.A2(n_435),
.B1(n_422),
.B2(n_449),
.Y(n_508)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_508),
.Y(n_538)
);

OAI22xp5_ASAP7_75t_SL g544 ( 
.A1(n_509),
.A2(n_513),
.B1(n_519),
.B2(n_534),
.Y(n_544)
);

OAI21xp5_ASAP7_75t_SL g558 ( 
.A1(n_510),
.A2(n_485),
.B(n_476),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_SL g511 ( 
.A(n_466),
.B(n_452),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_SL g547 ( 
.A(n_511),
.B(n_497),
.Y(n_547)
);

AOI22xp5_ASAP7_75t_L g513 ( 
.A1(n_462),
.A2(n_424),
.B1(n_429),
.B2(n_439),
.Y(n_513)
);

OAI22xp5_ASAP7_75t_L g514 ( 
.A1(n_471),
.A2(n_455),
.B1(n_423),
.B2(n_438),
.Y(n_514)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_514),
.Y(n_540)
);

XNOR2xp5_ASAP7_75t_L g515 ( 
.A(n_482),
.B(n_456),
.Y(n_515)
);

XOR2xp5_ASAP7_75t_L g551 ( 
.A(n_515),
.B(n_527),
.Y(n_551)
);

CKINVDCx20_ASAP7_75t_R g516 ( 
.A(n_477),
.Y(n_516)
);

CKINVDCx20_ASAP7_75t_R g559 ( 
.A(n_516),
.Y(n_559)
);

MAJIxp5_ASAP7_75t_L g518 ( 
.A(n_466),
.B(n_456),
.C(n_438),
.Y(n_518)
);

AOI22xp5_ASAP7_75t_L g519 ( 
.A1(n_464),
.A2(n_423),
.B1(n_459),
.B2(n_440),
.Y(n_519)
);

CKINVDCx20_ASAP7_75t_R g520 ( 
.A(n_483),
.Y(n_520)
);

CKINVDCx20_ASAP7_75t_R g562 ( 
.A(n_520),
.Y(n_562)
);

OAI22xp5_ASAP7_75t_L g524 ( 
.A1(n_496),
.A2(n_458),
.B1(n_457),
.B2(n_454),
.Y(n_524)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_524),
.Y(n_542)
);

XNOR2xp5_ASAP7_75t_SL g526 ( 
.A(n_495),
.B(n_436),
.Y(n_526)
);

XNOR2xp5_ASAP7_75t_SL g535 ( 
.A(n_526),
.B(n_484),
.Y(n_535)
);

XNOR2xp5_ASAP7_75t_L g527 ( 
.A(n_495),
.B(n_457),
.Y(n_527)
);

XNOR2xp5_ASAP7_75t_L g530 ( 
.A(n_473),
.B(n_313),
.Y(n_530)
);

MAJIxp5_ASAP7_75t_L g531 ( 
.A(n_472),
.B(n_323),
.C(n_351),
.Y(n_531)
);

MAJIxp5_ASAP7_75t_L g553 ( 
.A(n_531),
.B(n_533),
.C(n_494),
.Y(n_553)
);

HB1xp67_ASAP7_75t_L g532 ( 
.A(n_467),
.Y(n_532)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_532),
.Y(n_555)
);

MAJIxp5_ASAP7_75t_L g533 ( 
.A(n_480),
.B(n_450),
.C(n_314),
.Y(n_533)
);

XNOR2xp5_ASAP7_75t_SL g580 ( 
.A(n_535),
.B(n_563),
.Y(n_580)
);

OAI21xp5_ASAP7_75t_L g536 ( 
.A1(n_521),
.A2(n_490),
.B(n_468),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_L g588 ( 
.A(n_536),
.B(n_549),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_L g537 ( 
.A(n_503),
.B(n_486),
.Y(n_537)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_537),
.Y(n_574)
);

FAx1_ASAP7_75t_SL g539 ( 
.A(n_499),
.B(n_470),
.CI(n_474),
.CON(n_539),
.SN(n_539)
);

XNOR2x2_ASAP7_75t_SL g587 ( 
.A(n_539),
.B(n_522),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_L g541 ( 
.A(n_525),
.B(n_483),
.Y(n_541)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_541),
.Y(n_590)
);

AOI21xp5_ASAP7_75t_L g545 ( 
.A1(n_499),
.A2(n_491),
.B(n_464),
.Y(n_545)
);

NOR2xp33_ASAP7_75t_L g571 ( 
.A(n_545),
.B(n_557),
.Y(n_571)
);

OAI22xp5_ASAP7_75t_SL g546 ( 
.A1(n_529),
.A2(n_465),
.B1(n_478),
.B2(n_479),
.Y(n_546)
);

AOI22xp5_ASAP7_75t_L g575 ( 
.A1(n_546),
.A2(n_512),
.B1(n_506),
.B2(n_513),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_SL g579 ( 
.A(n_547),
.B(n_559),
.Y(n_579)
);

OAI22xp5_ASAP7_75t_L g569 ( 
.A1(n_548),
.A2(n_554),
.B1(n_561),
.B2(n_564),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_L g549 ( 
.A(n_529),
.B(n_463),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_L g552 ( 
.A(n_528),
.B(n_463),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_L g589 ( 
.A(n_552),
.B(n_556),
.Y(n_589)
);

XNOR2xp5_ASAP7_75t_L g573 ( 
.A(n_553),
.B(n_558),
.Y(n_573)
);

OAI22xp5_ASAP7_75t_L g554 ( 
.A1(n_534),
.A2(n_476),
.B1(n_488),
.B2(n_492),
.Y(n_554)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_517),
.Y(n_556)
);

AOI21xp5_ASAP7_75t_L g557 ( 
.A1(n_509),
.A2(n_469),
.B(n_485),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_L g560 ( 
.A(n_528),
.B(n_475),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_L g592 ( 
.A(n_560),
.B(n_565),
.Y(n_592)
);

AOI22xp5_ASAP7_75t_L g561 ( 
.A1(n_506),
.A2(n_461),
.B1(n_476),
.B2(n_416),
.Y(n_561)
);

XNOR2xp5_ASAP7_75t_SL g563 ( 
.A(n_507),
.B(n_320),
.Y(n_563)
);

AOI21xp5_ASAP7_75t_L g564 ( 
.A1(n_521),
.A2(n_348),
.B(n_320),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_517),
.Y(n_565)
);

XNOR2xp5_ASAP7_75t_SL g566 ( 
.A(n_526),
.B(n_332),
.Y(n_566)
);

XNOR2xp5_ASAP7_75t_L g578 ( 
.A(n_566),
.B(n_530),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_SL g567 ( 
.A(n_510),
.B(n_348),
.Y(n_567)
);

CKINVDCx16_ASAP7_75t_R g577 ( 
.A(n_567),
.Y(n_577)
);

MAJIxp5_ASAP7_75t_L g568 ( 
.A(n_543),
.B(n_504),
.C(n_515),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_L g595 ( 
.A(n_568),
.B(n_570),
.Y(n_595)
);

CKINVDCx20_ASAP7_75t_R g570 ( 
.A(n_541),
.Y(n_570)
);

MAJIxp5_ASAP7_75t_L g572 ( 
.A(n_543),
.B(n_504),
.C(n_518),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_L g610 ( 
.A(n_572),
.B(n_579),
.Y(n_610)
);

OAI22xp5_ASAP7_75t_SL g596 ( 
.A1(n_575),
.A2(n_576),
.B1(n_585),
.B2(n_564),
.Y(n_596)
);

AOI22xp5_ASAP7_75t_L g576 ( 
.A1(n_544),
.A2(n_512),
.B1(n_501),
.B2(n_519),
.Y(n_576)
);

XNOR2xp5_ASAP7_75t_L g599 ( 
.A(n_578),
.B(n_586),
.Y(n_599)
);

NOR2xp33_ASAP7_75t_SL g581 ( 
.A(n_559),
.B(n_441),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_L g613 ( 
.A(n_581),
.B(n_582),
.Y(n_613)
);

NOR2xp33_ASAP7_75t_SL g582 ( 
.A(n_547),
.B(n_498),
.Y(n_582)
);

MAJIxp5_ASAP7_75t_L g583 ( 
.A(n_550),
.B(n_500),
.C(n_533),
.Y(n_583)
);

MAJIxp5_ASAP7_75t_L g598 ( 
.A(n_583),
.B(n_584),
.C(n_593),
.Y(n_598)
);

MAJIxp5_ASAP7_75t_L g584 ( 
.A(n_550),
.B(n_527),
.C(n_531),
.Y(n_584)
);

AOI22xp5_ASAP7_75t_L g585 ( 
.A1(n_544),
.A2(n_523),
.B1(n_522),
.B2(n_505),
.Y(n_585)
);

XNOR2xp5_ASAP7_75t_L g586 ( 
.A(n_551),
.B(n_523),
.Y(n_586)
);

XNOR2xp5_ASAP7_75t_L g603 ( 
.A(n_587),
.B(n_536),
.Y(n_603)
);

OAI22xp5_ASAP7_75t_SL g591 ( 
.A1(n_538),
.A2(n_548),
.B1(n_557),
.B2(n_540),
.Y(n_591)
);

AOI22xp5_ASAP7_75t_L g602 ( 
.A1(n_591),
.A2(n_561),
.B1(n_554),
.B2(n_540),
.Y(n_602)
);

MAJIxp5_ASAP7_75t_L g593 ( 
.A(n_551),
.B(n_505),
.C(n_332),
.Y(n_593)
);

CKINVDCx16_ASAP7_75t_R g594 ( 
.A(n_588),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_L g633 ( 
.A(n_594),
.B(n_601),
.Y(n_633)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_596),
.Y(n_625)
);

XOR2xp5_ASAP7_75t_L g597 ( 
.A(n_584),
.B(n_563),
.Y(n_597)
);

XNOR2xp5_ASAP7_75t_L g623 ( 
.A(n_597),
.B(n_600),
.Y(n_623)
);

XOR2xp5_ASAP7_75t_L g600 ( 
.A(n_573),
.B(n_563),
.Y(n_600)
);

MAJIxp5_ASAP7_75t_L g601 ( 
.A(n_568),
.B(n_553),
.C(n_538),
.Y(n_601)
);

OAI22xp5_ASAP7_75t_SL g624 ( 
.A1(n_602),
.A2(n_609),
.B1(n_575),
.B2(n_589),
.Y(n_624)
);

XNOR2xp5_ASAP7_75t_L g630 ( 
.A(n_603),
.B(n_608),
.Y(n_630)
);

AOI21xp5_ASAP7_75t_L g604 ( 
.A1(n_573),
.A2(n_558),
.B(n_545),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_SL g629 ( 
.A(n_604),
.B(n_607),
.Y(n_629)
);

NOR2xp33_ASAP7_75t_L g605 ( 
.A(n_591),
.B(n_572),
.Y(n_605)
);

CKINVDCx14_ASAP7_75t_R g619 ( 
.A(n_605),
.Y(n_619)
);

NOR2xp33_ASAP7_75t_L g606 ( 
.A(n_593),
.B(n_542),
.Y(n_606)
);

NOR2xp33_ASAP7_75t_SL g627 ( 
.A(n_606),
.B(n_615),
.Y(n_627)
);

MAJIxp5_ASAP7_75t_L g607 ( 
.A(n_583),
.B(n_542),
.C(n_567),
.Y(n_607)
);

XNOR2xp5_ASAP7_75t_L g608 ( 
.A(n_586),
.B(n_555),
.Y(n_608)
);

AOI22xp5_ASAP7_75t_L g609 ( 
.A1(n_569),
.A2(n_555),
.B1(n_546),
.B2(n_562),
.Y(n_609)
);

XNOR2xp5_ASAP7_75t_L g611 ( 
.A(n_587),
.B(n_566),
.Y(n_611)
);

NOR2xp33_ASAP7_75t_L g618 ( 
.A(n_611),
.B(n_580),
.Y(n_618)
);

XOR2xp5_ASAP7_75t_L g612 ( 
.A(n_585),
.B(n_566),
.Y(n_612)
);

XOR2xp5_ASAP7_75t_L g622 ( 
.A(n_612),
.B(n_608),
.Y(n_622)
);

MAJIxp5_ASAP7_75t_L g614 ( 
.A(n_578),
.B(n_552),
.C(n_560),
.Y(n_614)
);

MAJIxp5_ASAP7_75t_L g620 ( 
.A(n_614),
.B(n_574),
.C(n_592),
.Y(n_620)
);

NOR2xp33_ASAP7_75t_L g615 ( 
.A(n_590),
.B(n_562),
.Y(n_615)
);

A2O1A1Ixp33_ASAP7_75t_L g616 ( 
.A1(n_603),
.A2(n_588),
.B(n_590),
.C(n_574),
.Y(n_616)
);

AOI22xp5_ASAP7_75t_L g636 ( 
.A1(n_616),
.A2(n_624),
.B1(n_628),
.B2(n_596),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_L g617 ( 
.A(n_595),
.B(n_589),
.Y(n_617)
);

OR2x2_ASAP7_75t_L g638 ( 
.A(n_617),
.B(n_618),
.Y(n_638)
);

XNOR2xp5_ASAP7_75t_L g645 ( 
.A(n_620),
.B(n_622),
.Y(n_645)
);

MAJIxp5_ASAP7_75t_L g621 ( 
.A(n_601),
.B(n_571),
.C(n_576),
.Y(n_621)
);

MAJIxp5_ASAP7_75t_L g635 ( 
.A(n_621),
.B(n_598),
.C(n_607),
.Y(n_635)
);

CKINVDCx20_ASAP7_75t_R g626 ( 
.A(n_613),
.Y(n_626)
);

NOR2xp33_ASAP7_75t_SL g643 ( 
.A(n_626),
.B(n_599),
.Y(n_643)
);

OAI22xp33_ASAP7_75t_L g628 ( 
.A1(n_609),
.A2(n_577),
.B1(n_592),
.B2(n_549),
.Y(n_628)
);

BUFx24_ASAP7_75t_SL g631 ( 
.A(n_610),
.Y(n_631)
);

NOR2xp33_ASAP7_75t_L g637 ( 
.A(n_631),
.B(n_632),
.Y(n_637)
);

NOR2xp33_ASAP7_75t_SL g632 ( 
.A(n_598),
.B(n_565),
.Y(n_632)
);

XOR2xp5_ASAP7_75t_L g634 ( 
.A(n_597),
.B(n_580),
.Y(n_634)
);

NOR2xp33_ASAP7_75t_L g640 ( 
.A(n_634),
.B(n_599),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_SL g653 ( 
.A(n_635),
.B(n_642),
.Y(n_653)
);

OR2x2_ASAP7_75t_L g657 ( 
.A(n_636),
.B(n_641),
.Y(n_657)
);

OR2x2_ASAP7_75t_L g639 ( 
.A(n_625),
.B(n_539),
.Y(n_639)
);

O2A1O1Ixp33_ASAP7_75t_SL g660 ( 
.A1(n_639),
.A2(n_644),
.B(n_535),
.C(n_600),
.Y(n_660)
);

XNOR2xp5_ASAP7_75t_L g652 ( 
.A(n_640),
.B(n_649),
.Y(n_652)
);

AOI22xp5_ASAP7_75t_SL g641 ( 
.A1(n_624),
.A2(n_537),
.B1(n_602),
.B2(n_539),
.Y(n_641)
);

NOR2xp33_ASAP7_75t_L g642 ( 
.A(n_627),
.B(n_621),
.Y(n_642)
);

AOI21xp33_ASAP7_75t_L g658 ( 
.A1(n_643),
.A2(n_646),
.B(n_647),
.Y(n_658)
);

OR2x2_ASAP7_75t_L g644 ( 
.A(n_617),
.B(n_539),
.Y(n_644)
);

OAI21xp5_ASAP7_75t_SL g646 ( 
.A1(n_629),
.A2(n_611),
.B(n_612),
.Y(n_646)
);

AND2x2_ASAP7_75t_L g647 ( 
.A(n_628),
.B(n_614),
.Y(n_647)
);

INVxp33_ASAP7_75t_L g654 ( 
.A(n_647),
.Y(n_654)
);

INVx6_ASAP7_75t_L g648 ( 
.A(n_619),
.Y(n_648)
);

NOR2xp33_ASAP7_75t_L g651 ( 
.A(n_648),
.B(n_620),
.Y(n_651)
);

NOR2xp33_ASAP7_75t_L g649 ( 
.A(n_633),
.B(n_556),
.Y(n_649)
);

INVxp67_ASAP7_75t_L g650 ( 
.A(n_643),
.Y(n_650)
);

AO21x1_ASAP7_75t_L g667 ( 
.A1(n_650),
.A2(n_646),
.B(n_639),
.Y(n_667)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_651),
.Y(n_662)
);

XNOR2xp5_ASAP7_75t_L g655 ( 
.A(n_645),
.B(n_622),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_L g664 ( 
.A(n_655),
.B(n_656),
.Y(n_664)
);

NOR2xp33_ASAP7_75t_L g656 ( 
.A(n_648),
.B(n_630),
.Y(n_656)
);

AOI21xp5_ASAP7_75t_L g665 ( 
.A1(n_658),
.A2(n_659),
.B(n_638),
.Y(n_665)
);

A2O1A1Ixp33_ASAP7_75t_L g659 ( 
.A1(n_647),
.A2(n_616),
.B(n_630),
.C(n_535),
.Y(n_659)
);

OAI21xp5_ASAP7_75t_L g663 ( 
.A1(n_660),
.A2(n_644),
.B(n_639),
.Y(n_663)
);

NOR2xp33_ASAP7_75t_L g661 ( 
.A(n_652),
.B(n_645),
.Y(n_661)
);

AOI21xp5_ASAP7_75t_L g672 ( 
.A1(n_661),
.A2(n_666),
.B(n_668),
.Y(n_672)
);

AO21x1_ASAP7_75t_L g671 ( 
.A1(n_663),
.A2(n_665),
.B(n_667),
.Y(n_671)
);

AOI21xp5_ASAP7_75t_L g666 ( 
.A1(n_653),
.A2(n_635),
.B(n_638),
.Y(n_666)
);

AOI21x1_ASAP7_75t_SL g668 ( 
.A1(n_654),
.A2(n_637),
.B(n_636),
.Y(n_668)
);

AND2x2_ASAP7_75t_L g669 ( 
.A(n_662),
.B(n_654),
.Y(n_669)
);

NAND3xp33_ASAP7_75t_L g675 ( 
.A(n_669),
.B(n_670),
.C(n_673),
.Y(n_675)
);

NOR2xp33_ASAP7_75t_L g670 ( 
.A(n_664),
.B(n_657),
.Y(n_670)
);

AOI21xp5_ASAP7_75t_L g673 ( 
.A1(n_665),
.A2(n_657),
.B(n_623),
.Y(n_673)
);

MAJIxp5_ASAP7_75t_L g674 ( 
.A(n_672),
.B(n_641),
.C(n_623),
.Y(n_674)
);

AOI21xp5_ASAP7_75t_L g676 ( 
.A1(n_674),
.A2(n_671),
.B(n_660),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_SL g677 ( 
.A(n_676),
.B(n_675),
.Y(n_677)
);

O2A1O1Ixp33_ASAP7_75t_SL g678 ( 
.A1(n_677),
.A2(n_634),
.B(n_347),
.C(n_335),
.Y(n_678)
);

AOI21xp5_ASAP7_75t_L g679 ( 
.A1(n_678),
.A2(n_10),
.B(n_11),
.Y(n_679)
);


endmodule