module real_jpeg_31545_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_626, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_626;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_598;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_95;
wire n_541;
wire n_441;
wire n_557;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_553;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_574;
wire n_595;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_562;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_366;
wire n_620;
wire n_456;
wire n_578;
wire n_259;
wire n_556;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_560;
wire n_538;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_565;
wire n_466;
wire n_623;
wire n_353;
wire n_453;
wire n_551;
wire n_230;
wire n_417;
wire n_428;
wire n_216;
wire n_128;
wire n_202;
wire n_605;
wire n_483;
wire n_367;
wire n_127;
wire n_365;
wire n_356;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_550;
wire n_233;
wire n_73;
wire n_621;
wire n_532;
wire n_348;
wire n_516;
wire n_473;
wire n_252;
wire n_601;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_288;
wire n_83;
wire n_525;
wire n_221;
wire n_393;
wire n_489;
wire n_611;
wire n_104;
wire n_153;
wire n_443;
wire n_599;
wire n_337;
wire n_544;
wire n_131;
wire n_439;
wire n_607;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_561;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_569;
wire n_335;
wire n_214;
wire n_113;
wire n_566;
wire n_543;
wire n_251;
wire n_459;
wire n_576;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_577;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_564;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_593;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_590;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_612;
wire n_110;
wire n_195;
wire n_592;
wire n_533;
wire n_289;
wire n_117;
wire n_614;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_559;
wire n_232;
wire n_582;
wire n_448;
wire n_615;
wire n_212;
wire n_284;
wire n_579;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_583;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_589;
wire n_25;
wire n_542;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_515;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_323;
wire n_166;
wire n_176;
wire n_215;
wire n_286;
wire n_596;
wire n_312;
wire n_617;
wire n_325;
wire n_307;
wire n_316;
wire n_594;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_604;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_572;
wire n_155;
wire n_405;
wire n_412;
wire n_586;
wire n_548;
wire n_319;
wire n_493;
wire n_93;
wire n_242;
wire n_487;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_613;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_531;
wire n_546;
wire n_112;
wire n_554;
wire n_508;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_616;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_536;
wire n_148;
wire n_373;
wire n_563;
wire n_558;
wire n_510;
wire n_396;
wire n_501;
wire n_600;
wire n_392;
wire n_575;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_584;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_622;
wire n_183;
wire n_248;
wire n_192;
wire n_624;
wire n_318;
wire n_537;
wire n_603;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_475;
wire n_74;
wire n_404;
wire n_204;
wire n_158;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_585;
wire n_494;
wire n_539;
wire n_512;
wire n_75;
wire n_581;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_534;
wire n_256;
wire n_520;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_545;
wire n_484;
wire n_587;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_608;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_299;
wire n_243;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_602;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_571;
wire n_610;
wire n_573;
wire n_379;
wire n_141;
wire n_555;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_570;
wire n_28;
wire n_606;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_313;
wire n_42;
wire n_268;
wire n_597;
wire n_618;
wire n_609;
wire n_94;
wire n_547;
wire n_309;
wire n_294;
wire n_619;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_588;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_540;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_567;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_530;
wire n_361;
wire n_324;
wire n_86;
wire n_261;
wire n_549;
wire n_70;
wire n_568;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_580;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_468;
wire n_133;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_552;
wire n_408;
wire n_85;
wire n_591;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_0),
.Y(n_212)
);

BUFx12f_ASAP7_75t_L g321 ( 
.A(n_0),
.Y(n_321)
);

AOI22xp5_ASAP7_75t_L g46 ( 
.A1(n_1),
.A2(n_47),
.B1(n_51),
.B2(n_52),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_1),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_1),
.A2(n_51),
.B1(n_185),
.B2(n_186),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g313 ( 
.A1(n_1),
.A2(n_51),
.B1(n_314),
.B2(n_317),
.Y(n_313)
);

AOI22xp33_ASAP7_75t_L g80 ( 
.A1(n_2),
.A2(n_81),
.B1(n_85),
.B2(n_86),
.Y(n_80)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_2),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_2),
.A2(n_85),
.B1(n_216),
.B2(n_219),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_2),
.A2(n_85),
.B1(n_254),
.B2(n_258),
.Y(n_253)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_3),
.Y(n_99)
);

BUFx3_ASAP7_75t_L g105 ( 
.A(n_3),
.Y(n_105)
);

BUFx3_ASAP7_75t_L g240 ( 
.A(n_3),
.Y(n_240)
);

BUFx6f_ASAP7_75t_L g172 ( 
.A(n_4),
.Y(n_172)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_5),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_5),
.Y(n_71)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_5),
.Y(n_440)
);

AO22x1_ASAP7_75t_SL g36 ( 
.A1(n_6),
.A2(n_37),
.B1(n_41),
.B2(n_44),
.Y(n_36)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_6),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_6),
.A2(n_44),
.B1(n_147),
.B2(n_149),
.Y(n_146)
);

NOR2xp67_ASAP7_75t_SL g380 ( 
.A(n_7),
.B(n_381),
.Y(n_380)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_7),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_7),
.B(n_139),
.Y(n_443)
);

OAI32xp33_ASAP7_75t_L g470 ( 
.A1(n_7),
.A2(n_52),
.A3(n_471),
.B1(n_475),
.B2(n_482),
.Y(n_470)
);

AOI22xp33_ASAP7_75t_L g514 ( 
.A1(n_7),
.A2(n_414),
.B1(n_515),
.B2(n_517),
.Y(n_514)
);

OAI32xp33_ASAP7_75t_L g522 ( 
.A1(n_7),
.A2(n_52),
.A3(n_471),
.B1(n_475),
.B2(n_482),
.Y(n_522)
);

OAI21xp33_ASAP7_75t_L g582 ( 
.A1(n_7),
.A2(n_214),
.B(n_583),
.Y(n_582)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_8),
.A2(n_131),
.B1(n_132),
.B2(n_135),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_8),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_8),
.A2(n_131),
.B1(n_225),
.B2(n_228),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_SL g323 ( 
.A1(n_8),
.A2(n_131),
.B1(n_324),
.B2(n_329),
.Y(n_323)
);

AOI22xp5_ASAP7_75t_SL g436 ( 
.A1(n_8),
.A2(n_131),
.B1(n_437),
.B2(n_441),
.Y(n_436)
);

OAI22xp5_ASAP7_75t_L g235 ( 
.A1(n_9),
.A2(n_236),
.B1(n_237),
.B2(n_241),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_9),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g348 ( 
.A1(n_9),
.A2(n_236),
.B1(n_349),
.B2(n_353),
.Y(n_348)
);

AOI22xp33_ASAP7_75t_SL g465 ( 
.A1(n_9),
.A2(n_236),
.B1(n_405),
.B2(n_466),
.Y(n_465)
);

AOI22xp33_ASAP7_75t_SL g539 ( 
.A1(n_9),
.A2(n_236),
.B1(n_540),
.B2(n_542),
.Y(n_539)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_10),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_10),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_10),
.Y(n_67)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_10),
.Y(n_203)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_11),
.Y(n_102)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_11),
.Y(n_109)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_12),
.Y(n_61)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_12),
.Y(n_64)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_12),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_13),
.A2(n_154),
.B1(n_159),
.B2(n_160),
.Y(n_153)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_13),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_13),
.A2(n_159),
.B1(n_199),
.B2(n_204),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_13),
.A2(n_159),
.B1(n_241),
.B2(n_248),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g360 ( 
.A1(n_13),
.A2(n_159),
.B1(n_361),
.B2(n_363),
.Y(n_360)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_14),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_14),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g158 ( 
.A(n_14),
.Y(n_158)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_14),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g302 ( 
.A1(n_15),
.A2(n_303),
.B1(n_304),
.B2(n_307),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_15),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_SL g417 ( 
.A1(n_15),
.A2(n_303),
.B1(n_418),
.B2(n_422),
.Y(n_417)
);

AOI22xp33_ASAP7_75t_SL g505 ( 
.A1(n_15),
.A2(n_303),
.B1(n_506),
.B2(n_510),
.Y(n_505)
);

AOI22xp33_ASAP7_75t_SL g529 ( 
.A1(n_15),
.A2(n_303),
.B1(n_530),
.B2(n_533),
.Y(n_529)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_16),
.A2(n_123),
.B1(n_125),
.B2(n_126),
.Y(n_122)
);

INVx1_ASAP7_75t_SL g125 ( 
.A(n_16),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g294 ( 
.A1(n_16),
.A2(n_116),
.B1(n_125),
.B2(n_295),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_SL g403 ( 
.A1(n_16),
.A2(n_125),
.B1(n_404),
.B2(n_405),
.Y(n_403)
);

OAI22xp33_ASAP7_75t_SL g492 ( 
.A1(n_16),
.A2(n_125),
.B1(n_217),
.B2(n_493),
.Y(n_492)
);

XNOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_271),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_SL g18 ( 
.A(n_19),
.B(n_270),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_242),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_21),
.B(n_242),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_140),
.C(n_193),
.Y(n_21)
);

HB1xp67_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_23),
.B(n_141),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_91),
.Y(n_23)
);

OAI21xp33_ASAP7_75t_SL g265 ( 
.A1(n_24),
.A2(n_266),
.B(n_267),
.Y(n_265)
);

AND2x2_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_45),
.Y(n_24)
);

XOR2xp5_ASAP7_75t_L g91 ( 
.A(n_25),
.B(n_92),
.Y(n_91)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_25),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_SL g286 ( 
.A1(n_25),
.A2(n_266),
.B1(n_287),
.B2(n_288),
.Y(n_286)
);

OA21x2_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_33),
.B(n_36),
.Y(n_25)
);

INVx1_ASAP7_75t_SL g214 ( 
.A(n_26),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g358 ( 
.A1(n_26),
.A2(n_313),
.B1(n_359),
.B2(n_365),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g491 ( 
.A(n_26),
.B(n_492),
.Y(n_491)
);

AOI22xp33_ASAP7_75t_L g527 ( 
.A1(n_26),
.A2(n_528),
.B1(n_536),
.B2(n_538),
.Y(n_527)
);

AND2x2_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_30),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_28),
.Y(n_362)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_28),
.Y(n_535)
);

HB1xp67_ASAP7_75t_L g565 ( 
.A(n_28),
.Y(n_565)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_29),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g316 ( 
.A(n_29),
.Y(n_316)
);

INVx3_ASAP7_75t_L g547 ( 
.A(n_29),
.Y(n_547)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_32),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g367 ( 
.A(n_32),
.Y(n_367)
);

INVx2_ASAP7_75t_L g588 ( 
.A(n_32),
.Y(n_588)
);

INVx3_ASAP7_75t_SL g33 ( 
.A(n_34),
.Y(n_33)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_36),
.Y(n_213)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

BUFx2_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx2_ASAP7_75t_L g364 ( 
.A(n_42),
.Y(n_364)
);

BUFx2_ASAP7_75t_SL g532 ( 
.A(n_42),
.Y(n_532)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_43),
.Y(n_77)
);

INVx2_ASAP7_75t_L g495 ( 
.A(n_43),
.Y(n_495)
);

INVxp67_ASAP7_75t_SL g288 ( 
.A(n_45),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_L g45 ( 
.A1(n_46),
.A2(n_56),
.B1(n_80),
.B2(n_89),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_46),
.A2(n_56),
.B1(n_89),
.B2(n_198),
.Y(n_197)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx2_ASAP7_75t_SL g49 ( 
.A(n_50),
.Y(n_49)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_50),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g331 ( 
.A(n_50),
.Y(n_331)
);

INVx1_ASAP7_75t_SL g52 ( 
.A(n_53),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx4_ASAP7_75t_L g558 ( 
.A(n_54),
.Y(n_558)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_55),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g148 ( 
.A(n_55),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g169 ( 
.A(n_55),
.Y(n_169)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_55),
.Y(n_207)
);

BUFx6f_ASAP7_75t_L g509 ( 
.A(n_55),
.Y(n_509)
);

BUFx6f_ASAP7_75t_L g576 ( 
.A(n_55),
.Y(n_576)
);

INVx2_ASAP7_75t_SL g145 ( 
.A(n_56),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g322 ( 
.A1(n_56),
.A2(n_89),
.B1(n_198),
.B2(n_323),
.Y(n_322)
);

OAI21xp33_ASAP7_75t_SL g464 ( 
.A1(n_56),
.A2(n_465),
.B(n_468),
.Y(n_464)
);

OAI22xp5_ASAP7_75t_SL g504 ( 
.A1(n_56),
.A2(n_89),
.B1(n_465),
.B2(n_505),
.Y(n_504)
);

OR2x2_ASAP7_75t_L g56 ( 
.A(n_57),
.B(n_68),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_L g57 ( 
.A1(n_58),
.A2(n_60),
.B1(n_62),
.B2(n_65),
.Y(n_57)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

HB1xp67_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx2_ASAP7_75t_L g568 ( 
.A(n_61),
.Y(n_568)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_64),
.Y(n_79)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_66),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_67),
.Y(n_84)
);

BUFx3_ASAP7_75t_L g90 ( 
.A(n_68),
.Y(n_90)
);

OAI22x1_ASAP7_75t_L g68 ( 
.A1(n_69),
.A2(n_72),
.B1(n_76),
.B2(n_78),
.Y(n_68)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g218 ( 
.A(n_71),
.Y(n_218)
);

INVx6_ASAP7_75t_L g221 ( 
.A(n_71),
.Y(n_221)
);

BUFx6f_ASAP7_75t_L g554 ( 
.A(n_71),
.Y(n_554)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_79),
.Y(n_560)
);

INVxp67_ASAP7_75t_L g144 ( 
.A(n_80),
.Y(n_144)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g511 ( 
.A(n_84),
.Y(n_511)
);

BUFx2_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx3_ASAP7_75t_SL g87 ( 
.A(n_88),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_SL g579 ( 
.A(n_89),
.B(n_414),
.Y(n_579)
);

INVx2_ASAP7_75t_SL g89 ( 
.A(n_90),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_90),
.A2(n_144),
.B1(n_145),
.B2(n_146),
.Y(n_143)
);

OA21x2_ASAP7_75t_L g251 ( 
.A1(n_90),
.A2(n_145),
.B(n_146),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_SL g402 ( 
.A1(n_90),
.A2(n_145),
.B1(n_403),
.B2(n_407),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g468 ( 
.A(n_90),
.B(n_403),
.Y(n_468)
);

AO22x1_ASAP7_75t_L g608 ( 
.A1(n_90),
.A2(n_145),
.B1(n_403),
.B2(n_609),
.Y(n_608)
);

HB1xp67_ASAP7_75t_L g267 ( 
.A(n_92),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_93),
.B(n_129),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_93),
.B(n_344),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_122),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_94),
.B(n_235),
.Y(n_234)
);

BUFx2_ASAP7_75t_L g245 ( 
.A(n_94),
.Y(n_245)
);

AO22x2_ASAP7_75t_SL g301 ( 
.A1(n_94),
.A2(n_139),
.B1(n_235),
.B2(n_302),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_SL g409 ( 
.A(n_94),
.B(n_410),
.Y(n_409)
);

AND2x2_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_110),
.Y(n_94)
);

OAI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_96),
.A2(n_100),
.B1(n_103),
.B2(n_106),
.Y(n_95)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVx2_ASAP7_75t_L g306 ( 
.A(n_98),
.Y(n_306)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_99),
.Y(n_124)
);

INVx6_ASAP7_75t_L g128 ( 
.A(n_99),
.Y(n_128)
);

BUFx3_ASAP7_75t_L g134 ( 
.A(n_99),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g249 ( 
.A(n_99),
.Y(n_249)
);

BUFx3_ASAP7_75t_L g309 ( 
.A(n_99),
.Y(n_309)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_102),
.Y(n_112)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_102),
.Y(n_121)
);

INVx2_ASAP7_75t_L g374 ( 
.A(n_102),
.Y(n_374)
);

BUFx3_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g138 ( 
.A(n_105),
.Y(n_138)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_109),
.Y(n_390)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_110),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_111),
.A2(n_113),
.B1(n_116),
.B2(n_119),
.Y(n_110)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g516 ( 
.A(n_114),
.Y(n_516)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g188 ( 
.A(n_115),
.Y(n_188)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_115),
.Y(n_227)
);

BUFx6f_ASAP7_75t_L g298 ( 
.A(n_115),
.Y(n_298)
);

BUFx12f_ASAP7_75t_L g352 ( 
.A(n_115),
.Y(n_352)
);

BUFx6f_ASAP7_75t_L g387 ( 
.A(n_115),
.Y(n_387)
);

INVx5_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

BUFx2_ASAP7_75t_L g354 ( 
.A(n_117),
.Y(n_354)
);

INVx8_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g185 ( 
.A(n_118),
.Y(n_185)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_122),
.B(n_139),
.Y(n_233)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_123),
.Y(n_241)
);

BUFx4f_ASAP7_75t_SL g123 ( 
.A(n_124),
.Y(n_123)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVx3_ASAP7_75t_L g379 ( 
.A(n_128),
.Y(n_379)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_128),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_139),
.Y(n_129)
);

AOI22x1_ASAP7_75t_SL g244 ( 
.A1(n_130),
.A2(n_245),
.B1(n_246),
.B2(n_247),
.Y(n_244)
);

INVx2_ASAP7_75t_SL g132 ( 
.A(n_133),
.Y(n_132)
);

INVx3_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

HB1xp67_ASAP7_75t_L g246 ( 
.A(n_139),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_139),
.B(n_302),
.Y(n_344)
);

HB1xp67_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_192),
.Y(n_141)
);

OR2x2_ASAP7_75t_L g142 ( 
.A(n_143),
.B(n_152),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_143),
.B(n_152),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g571 ( 
.A(n_145),
.B(n_572),
.Y(n_571)
);

BUFx6f_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_148),
.A2(n_168),
.B1(n_170),
.B2(n_173),
.Y(n_167)
);

INVx1_ASAP7_75t_SL g149 ( 
.A(n_150),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

BUFx2_ASAP7_75t_L g467 ( 
.A(n_151),
.Y(n_467)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_153),
.A2(n_166),
.B1(n_184),
.B2(n_189),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_153),
.A2(n_166),
.B1(n_191),
.B2(n_224),
.Y(n_223)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

INVx8_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

INVx3_ASAP7_75t_L g371 ( 
.A(n_158),
.Y(n_371)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_161),
.A2(n_176),
.B1(n_178),
.B2(n_181),
.Y(n_175)
);

INVx3_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

INVx4_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_164),
.Y(n_177)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_164),
.Y(n_423)
);

BUFx6f_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g231 ( 
.A(n_165),
.Y(n_231)
);

BUFx5_ASAP7_75t_L g257 ( 
.A(n_165),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_166),
.A2(n_184),
.B1(n_189),
.B2(n_253),
.Y(n_252)
);

INVx2_ASAP7_75t_L g299 ( 
.A(n_166),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g416 ( 
.A1(n_166),
.A2(n_417),
.B1(n_424),
.B2(n_425),
.Y(n_416)
);

AO22x1_ASAP7_75t_SL g434 ( 
.A1(n_166),
.A2(n_191),
.B1(n_294),
.B2(n_417),
.Y(n_434)
);

AND2x4_ASAP7_75t_L g166 ( 
.A(n_167),
.B(n_175),
.Y(n_166)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_167),
.Y(n_191)
);

INVxp67_ASAP7_75t_SL g356 ( 
.A(n_167),
.Y(n_356)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

INVx3_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

BUFx3_ASAP7_75t_L g174 ( 
.A(n_172),
.Y(n_174)
);

BUFx6f_ASAP7_75t_L g180 ( 
.A(n_172),
.Y(n_180)
);

BUFx6f_ASAP7_75t_L g183 ( 
.A(n_172),
.Y(n_183)
);

BUFx3_ASAP7_75t_L g481 ( 
.A(n_172),
.Y(n_481)
);

INVx5_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

INVx4_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

INVx5_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

BUFx6f_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

BUFx4f_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

INVx2_ASAP7_75t_SL g187 ( 
.A(n_188),
.Y(n_187)
);

INVx4_ASAP7_75t_L g519 ( 
.A(n_188),
.Y(n_519)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

OAI22x1_ASAP7_75t_L g292 ( 
.A1(n_190),
.A2(n_293),
.B1(n_299),
.B2(n_300),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_SL g611 ( 
.A(n_190),
.B(n_414),
.Y(n_611)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

HB1xp67_ASAP7_75t_L g264 ( 
.A(n_192),
.Y(n_264)
);

INVxp33_ASAP7_75t_SL g193 ( 
.A(n_194),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_194),
.B(n_278),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_195),
.B(n_222),
.C(n_232),
.Y(n_194)
);

INVxp67_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_196),
.B(n_283),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_197),
.B(n_208),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g340 ( 
.A(n_197),
.B(n_208),
.Y(n_340)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

HB1xp67_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

BUFx6f_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

BUFx5_ASAP7_75t_L g328 ( 
.A(n_203),
.Y(n_328)
);

BUFx3_ASAP7_75t_L g487 ( 
.A(n_203),
.Y(n_487)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

INVx3_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

INVx3_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

OAI22xp33_ASAP7_75t_SL g208 ( 
.A1(n_209),
.A2(n_213),
.B1(n_214),
.B2(n_215),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

BUFx2_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_212),
.Y(n_594)
);

OAI22xp5_ASAP7_75t_SL g311 ( 
.A1(n_214),
.A2(n_215),
.B1(n_312),
.B2(n_318),
.Y(n_311)
);

OAI22xp5_ASAP7_75t_L g435 ( 
.A1(n_214),
.A2(n_318),
.B1(n_360),
.B2(n_436),
.Y(n_435)
);

OAI21xp5_ASAP7_75t_L g605 ( 
.A1(n_214),
.A2(n_539),
.B(n_583),
.Y(n_605)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

HB1xp67_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_218),
.Y(n_317)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

BUFx2_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

INVx2_ASAP7_75t_L g598 ( 
.A(n_221),
.Y(n_598)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_222),
.A2(n_223),
.B1(n_232),
.B2(n_284),
.Y(n_283)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_224),
.Y(n_300)
);

HB1xp67_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

HB1xp67_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_231),
.Y(n_260)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_231),
.Y(n_421)
);

INVx2_ASAP7_75t_L g477 ( 
.A(n_231),
.Y(n_477)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_232),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_233),
.B(n_234),
.Y(n_232)
);

AND2x2_ASAP7_75t_L g408 ( 
.A(n_233),
.B(n_409),
.Y(n_408)
);

HB1xp67_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_243),
.B(n_263),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_244),
.B(n_250),
.Y(n_243)
);

BUFx6f_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_251),
.A2(n_252),
.B1(n_261),
.B2(n_262),
.Y(n_250)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_251),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_252),
.Y(n_262)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

INVx3_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

HB1xp67_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_L g263 ( 
.A1(n_264),
.A2(n_265),
.B1(n_268),
.B2(n_269),
.Y(n_263)
);

INVxp67_ASAP7_75t_SL g269 ( 
.A(n_264),
.Y(n_269)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_265),
.Y(n_268)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

NAND2x1_ASAP7_75t_L g272 ( 
.A(n_273),
.B(n_451),
.Y(n_272)
);

AOI21xp5_ASAP7_75t_L g273 ( 
.A1(n_274),
.A2(n_391),
.B(n_447),
.Y(n_273)
);

INVxp67_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g621 ( 
.A(n_275),
.B(n_622),
.Y(n_621)
);

OAI21xp5_ASAP7_75t_SL g275 ( 
.A1(n_276),
.A2(n_279),
.B(n_332),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_276),
.B(n_279),
.Y(n_450)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

AND2x2_ASAP7_75t_L g449 ( 
.A(n_277),
.B(n_280),
.Y(n_449)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_281),
.B(n_285),
.C(n_289),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g333 ( 
.A(n_281),
.B(n_334),
.Y(n_333)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

INVxp67_ASAP7_75t_SL g285 ( 
.A(n_286),
.Y(n_285)
);

XOR2xp5_ASAP7_75t_L g334 ( 
.A(n_286),
.B(n_290),
.Y(n_334)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

INVxp33_ASAP7_75t_SL g289 ( 
.A(n_290),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_291),
.B(n_301),
.C(n_310),
.Y(n_290)
);

HB1xp67_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_L g338 ( 
.A(n_292),
.B(n_301),
.Y(n_338)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_294),
.B(n_356),
.Y(n_355)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

INVx2_ASAP7_75t_L g296 ( 
.A(n_297),
.Y(n_296)
);

INVx2_ASAP7_75t_L g474 ( 
.A(n_297),
.Y(n_474)
);

INVx2_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

OAI21xp5_ASAP7_75t_L g347 ( 
.A1(n_299),
.A2(n_348),
.B(n_355),
.Y(n_347)
);

OAI21xp5_ASAP7_75t_L g513 ( 
.A1(n_299),
.A2(n_355),
.B(n_514),
.Y(n_513)
);

INVx3_ASAP7_75t_L g304 ( 
.A(n_305),
.Y(n_304)
);

INVx4_ASAP7_75t_L g305 ( 
.A(n_306),
.Y(n_305)
);

BUFx3_ASAP7_75t_L g307 ( 
.A(n_308),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_309),
.Y(n_308)
);

BUFx6f_ASAP7_75t_L g413 ( 
.A(n_309),
.Y(n_413)
);

XNOR2xp5_ASAP7_75t_L g337 ( 
.A(n_310),
.B(n_338),
.Y(n_337)
);

AND2x2_ASAP7_75t_L g310 ( 
.A(n_311),
.B(n_322),
.Y(n_310)
);

XNOR2x2_ASAP7_75t_L g400 ( 
.A(n_311),
.B(n_322),
.Y(n_400)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_313),
.Y(n_312)
);

BUFx3_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

INVx6_ASAP7_75t_L g315 ( 
.A(n_316),
.Y(n_315)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_317),
.Y(n_441)
);

OAI21xp5_ASAP7_75t_SL g580 ( 
.A1(n_318),
.A2(n_491),
.B(n_529),
.Y(n_580)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_319),
.Y(n_318)
);

INVx5_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

BUFx3_ASAP7_75t_L g537 ( 
.A(n_320),
.Y(n_537)
);

INVx8_ASAP7_75t_L g320 ( 
.A(n_321),
.Y(n_320)
);

INVx8_ASAP7_75t_L g490 ( 
.A(n_321),
.Y(n_490)
);

INVxp67_ASAP7_75t_SL g407 ( 
.A(n_323),
.Y(n_407)
);

INVx2_ASAP7_75t_L g324 ( 
.A(n_325),
.Y(n_324)
);

INVx3_ASAP7_75t_L g325 ( 
.A(n_326),
.Y(n_325)
);

INVx2_ASAP7_75t_L g326 ( 
.A(n_327),
.Y(n_326)
);

INVx4_ASAP7_75t_L g327 ( 
.A(n_328),
.Y(n_327)
);

INVx4_ASAP7_75t_L g329 ( 
.A(n_330),
.Y(n_329)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_330),
.Y(n_404)
);

INVx4_ASAP7_75t_L g330 ( 
.A(n_331),
.Y(n_330)
);

BUFx6f_ASAP7_75t_L g406 ( 
.A(n_331),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_333),
.B(n_335),
.Y(n_332)
);

OR2x2_ASAP7_75t_L g448 ( 
.A(n_333),
.B(n_335),
.Y(n_448)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_336),
.B(n_339),
.C(n_341),
.Y(n_335)
);

HB1xp67_ASAP7_75t_L g336 ( 
.A(n_337),
.Y(n_336)
);

XOR2xp5_ASAP7_75t_L g394 ( 
.A(n_337),
.B(n_340),
.Y(n_394)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_340),
.Y(n_339)
);

XNOR2x1_ASAP7_75t_L g393 ( 
.A(n_341),
.B(n_394),
.Y(n_393)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_342),
.B(n_345),
.C(n_357),
.Y(n_341)
);

OAI22xp5_ASAP7_75t_L g398 ( 
.A1(n_342),
.A2(n_343),
.B1(n_346),
.B2(n_347),
.Y(n_398)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_343),
.Y(n_342)
);

HB1xp67_ASAP7_75t_L g345 ( 
.A(n_346),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_347),
.Y(n_346)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_348),
.Y(n_424)
);

INVx2_ASAP7_75t_L g349 ( 
.A(n_350),
.Y(n_349)
);

INVx3_ASAP7_75t_L g350 ( 
.A(n_351),
.Y(n_350)
);

INVx2_ASAP7_75t_L g351 ( 
.A(n_352),
.Y(n_351)
);

INVx1_ASAP7_75t_SL g353 ( 
.A(n_354),
.Y(n_353)
);

BUFx2_ASAP7_75t_L g425 ( 
.A(n_356),
.Y(n_425)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_357),
.Y(n_399)
);

OR2x2_ASAP7_75t_L g357 ( 
.A(n_358),
.B(n_368),
.Y(n_357)
);

XOR2xp5_ASAP7_75t_SL g430 ( 
.A(n_358),
.B(n_431),
.Y(n_430)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_360),
.Y(n_359)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_362),
.Y(n_361)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_364),
.Y(n_363)
);

INVx3_ASAP7_75t_L g365 ( 
.A(n_366),
.Y(n_365)
);

INVx3_ASAP7_75t_L g366 ( 
.A(n_367),
.Y(n_366)
);

AOI32xp33_ASAP7_75t_L g368 ( 
.A1(n_369),
.A2(n_372),
.A3(n_375),
.B1(n_380),
.B2(n_383),
.Y(n_368)
);

AOI32xp33_ASAP7_75t_L g431 ( 
.A1(n_369),
.A2(n_372),
.A3(n_375),
.B1(n_380),
.B2(n_383),
.Y(n_431)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_370),
.Y(n_369)
);

INVx2_ASAP7_75t_L g370 ( 
.A(n_371),
.Y(n_370)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_373),
.Y(n_372)
);

INVx2_ASAP7_75t_L g373 ( 
.A(n_374),
.Y(n_373)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_376),
.Y(n_375)
);

INVx2_ASAP7_75t_L g376 ( 
.A(n_377),
.Y(n_376)
);

INVx2_ASAP7_75t_L g377 ( 
.A(n_378),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_379),
.Y(n_378)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_380),
.Y(n_415)
);

INVx3_ASAP7_75t_L g381 ( 
.A(n_382),
.Y(n_381)
);

NAND2xp33_ASAP7_75t_L g383 ( 
.A(n_384),
.B(n_388),
.Y(n_383)
);

BUFx2_ASAP7_75t_L g384 ( 
.A(n_385),
.Y(n_384)
);

INVx2_ASAP7_75t_L g385 ( 
.A(n_386),
.Y(n_385)
);

INVx2_ASAP7_75t_L g386 ( 
.A(n_387),
.Y(n_386)
);

INVx3_ASAP7_75t_L g388 ( 
.A(n_389),
.Y(n_388)
);

INVx3_ASAP7_75t_L g389 ( 
.A(n_390),
.Y(n_389)
);

MAJIxp5_ASAP7_75t_L g391 ( 
.A(n_392),
.B(n_395),
.C(n_426),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_393),
.Y(n_392)
);

OAI21xp33_ASAP7_75t_L g622 ( 
.A1(n_393),
.A2(n_623),
.B(n_624),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_395),
.Y(n_623)
);

MAJx2_ASAP7_75t_L g395 ( 
.A(n_396),
.B(n_400),
.C(n_401),
.Y(n_395)
);

AOI22xp5_ASAP7_75t_SL g444 ( 
.A1(n_396),
.A2(n_397),
.B1(n_445),
.B2(n_446),
.Y(n_444)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_397),
.Y(n_396)
);

XNOR2xp5_ASAP7_75t_L g397 ( 
.A(n_398),
.B(n_399),
.Y(n_397)
);

XNOR2x1_ASAP7_75t_L g445 ( 
.A(n_400),
.B(n_401),
.Y(n_445)
);

MAJx2_ASAP7_75t_L g401 ( 
.A(n_402),
.B(n_408),
.C(n_416),
.Y(n_401)
);

XNOR2xp5_ASAP7_75t_L g429 ( 
.A(n_402),
.B(n_416),
.Y(n_429)
);

INVx3_ASAP7_75t_L g405 ( 
.A(n_406),
.Y(n_405)
);

XOR2xp5_ASAP7_75t_L g428 ( 
.A(n_408),
.B(n_429),
.Y(n_428)
);

OAI21xp5_ASAP7_75t_SL g410 ( 
.A1(n_411),
.A2(n_414),
.B(n_415),
.Y(n_410)
);

INVx3_ASAP7_75t_L g411 ( 
.A(n_412),
.Y(n_411)
);

INVx8_ASAP7_75t_L g412 ( 
.A(n_413),
.Y(n_412)
);

NOR2xp33_ASAP7_75t_L g482 ( 
.A(n_414),
.B(n_483),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_SL g569 ( 
.A(n_414),
.B(n_486),
.Y(n_569)
);

OAI21xp33_ASAP7_75t_SL g572 ( 
.A1(n_414),
.A2(n_569),
.B(n_573),
.Y(n_572)
);

NOR2xp33_ASAP7_75t_L g590 ( 
.A(n_414),
.B(n_591),
.Y(n_590)
);

INVx2_ASAP7_75t_L g418 ( 
.A(n_419),
.Y(n_418)
);

HB1xp67_ASAP7_75t_L g419 ( 
.A(n_420),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_421),
.Y(n_420)
);

INVx1_ASAP7_75t_SL g422 ( 
.A(n_423),
.Y(n_422)
);

OR2x2_ASAP7_75t_L g426 ( 
.A(n_427),
.B(n_444),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_SL g624 ( 
.A(n_427),
.B(n_444),
.Y(n_624)
);

MAJIxp5_ASAP7_75t_L g427 ( 
.A(n_428),
.B(n_430),
.C(n_432),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_SL g454 ( 
.A(n_428),
.B(n_455),
.Y(n_454)
);

OR2x2_ASAP7_75t_L g457 ( 
.A(n_428),
.B(n_455),
.Y(n_457)
);

OAI22xp5_ASAP7_75t_SL g455 ( 
.A1(n_430),
.A2(n_432),
.B1(n_433),
.B2(n_456),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_430),
.Y(n_456)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_433),
.Y(n_432)
);

MAJIxp5_ASAP7_75t_L g433 ( 
.A(n_434),
.B(n_435),
.C(n_442),
.Y(n_433)
);

XNOR2xp5_ASAP7_75t_SL g460 ( 
.A(n_434),
.B(n_461),
.Y(n_460)
);

AOI22xp5_ASAP7_75t_L g461 ( 
.A1(n_435),
.A2(n_442),
.B1(n_443),
.B2(n_462),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_435),
.Y(n_462)
);

OAI21xp5_ASAP7_75t_L g488 ( 
.A1(n_436),
.A2(n_489),
.B(n_491),
.Y(n_488)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_438),
.Y(n_437)
);

BUFx2_ASAP7_75t_L g438 ( 
.A(n_439),
.Y(n_438)
);

INVx2_ASAP7_75t_L g439 ( 
.A(n_440),
.Y(n_439)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_443),
.Y(n_442)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_445),
.Y(n_446)
);

OAI21xp5_ASAP7_75t_L g447 ( 
.A1(n_448),
.A2(n_449),
.B(n_450),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_452),
.B(n_621),
.Y(n_451)
);

OAI21x1_ASAP7_75t_L g452 ( 
.A1(n_453),
.A2(n_496),
.B(n_620),
.Y(n_452)
);

AOI21xp5_ASAP7_75t_L g453 ( 
.A1(n_454),
.A2(n_457),
.B(n_458),
.Y(n_453)
);

NAND3xp33_ASAP7_75t_L g620 ( 
.A(n_454),
.B(n_457),
.C(n_458),
.Y(n_620)
);

MAJIxp5_ASAP7_75t_L g458 ( 
.A(n_459),
.B(n_463),
.C(n_469),
.Y(n_458)
);

INVxp67_ASAP7_75t_L g459 ( 
.A(n_460),
.Y(n_459)
);

XNOR2xp5_ASAP7_75t_L g498 ( 
.A(n_460),
.B(n_499),
.Y(n_498)
);

OAI22xp5_ASAP7_75t_L g499 ( 
.A1(n_463),
.A2(n_464),
.B1(n_469),
.B2(n_500),
.Y(n_499)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_464),
.Y(n_463)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_467),
.Y(n_466)
);

AND2x2_ASAP7_75t_L g570 ( 
.A(n_468),
.B(n_571),
.Y(n_570)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_469),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_470),
.B(n_488),
.Y(n_469)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_472),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_473),
.Y(n_472)
);

INVx2_ASAP7_75t_L g473 ( 
.A(n_474),
.Y(n_473)
);

NAND2xp67_ASAP7_75t_SL g475 ( 
.A(n_476),
.B(n_478),
.Y(n_475)
);

BUFx3_ASAP7_75t_L g476 ( 
.A(n_477),
.Y(n_476)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_479),
.Y(n_478)
);

HB1xp67_ASAP7_75t_L g479 ( 
.A(n_480),
.Y(n_479)
);

BUFx3_ASAP7_75t_L g480 ( 
.A(n_481),
.Y(n_480)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_484),
.Y(n_483)
);

INVx2_ASAP7_75t_L g484 ( 
.A(n_485),
.Y(n_484)
);

INVx2_ASAP7_75t_L g485 ( 
.A(n_486),
.Y(n_485)
);

INVx5_ASAP7_75t_L g486 ( 
.A(n_487),
.Y(n_486)
);

XOR2xp5_ASAP7_75t_L g521 ( 
.A(n_488),
.B(n_522),
.Y(n_521)
);

BUFx2_ASAP7_75t_L g489 ( 
.A(n_490),
.Y(n_489)
);

NAND2xp33_ASAP7_75t_SL g583 ( 
.A(n_492),
.B(n_584),
.Y(n_583)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_493),
.Y(n_541)
);

INVx4_ASAP7_75t_L g493 ( 
.A(n_494),
.Y(n_493)
);

INVx4_ASAP7_75t_L g494 ( 
.A(n_495),
.Y(n_494)
);

AOI21x1_ASAP7_75t_L g496 ( 
.A1(n_497),
.A2(n_524),
.B(n_619),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_SL g497 ( 
.A(n_498),
.B(n_501),
.Y(n_497)
);

NOR2xp67_ASAP7_75t_SL g619 ( 
.A(n_498),
.B(n_501),
.Y(n_619)
);

OAI21xp5_ASAP7_75t_L g501 ( 
.A1(n_502),
.A2(n_520),
.B(n_523),
.Y(n_501)
);

NOR2xp33_ASAP7_75t_L g502 ( 
.A(n_503),
.B(n_512),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_SL g523 ( 
.A(n_503),
.B(n_512),
.Y(n_523)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_504),
.Y(n_503)
);

XNOR2xp5_ASAP7_75t_L g603 ( 
.A(n_504),
.B(n_513),
.Y(n_603)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_505),
.Y(n_609)
);

INVx1_ASAP7_75t_SL g506 ( 
.A(n_507),
.Y(n_506)
);

INVx2_ASAP7_75t_L g507 ( 
.A(n_508),
.Y(n_507)
);

INVx2_ASAP7_75t_SL g508 ( 
.A(n_509),
.Y(n_508)
);

BUFx2_ASAP7_75t_L g510 ( 
.A(n_511),
.Y(n_510)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_513),
.Y(n_512)
);

INVx2_ASAP7_75t_L g515 ( 
.A(n_516),
.Y(n_515)
);

BUFx3_ASAP7_75t_L g517 ( 
.A(n_518),
.Y(n_517)
);

INVx3_ASAP7_75t_L g518 ( 
.A(n_519),
.Y(n_518)
);

HB1xp67_ASAP7_75t_L g520 ( 
.A(n_521),
.Y(n_520)
);

XOR2xp5_ASAP7_75t_L g602 ( 
.A(n_521),
.B(n_603),
.Y(n_602)
);

OAI321xp33_ASAP7_75t_L g524 ( 
.A1(n_525),
.A2(n_601),
.A3(n_612),
.B1(n_617),
.B2(n_618),
.C(n_626),
.Y(n_524)
);

AOI21xp5_ASAP7_75t_L g525 ( 
.A1(n_526),
.A2(n_577),
.B(n_600),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_L g526 ( 
.A(n_527),
.B(n_548),
.Y(n_526)
);

NOR2xp33_ASAP7_75t_L g600 ( 
.A(n_527),
.B(n_548),
.Y(n_600)
);

INVxp67_ASAP7_75t_L g528 ( 
.A(n_529),
.Y(n_528)
);

BUFx3_ASAP7_75t_L g530 ( 
.A(n_531),
.Y(n_530)
);

INVx2_ASAP7_75t_L g531 ( 
.A(n_532),
.Y(n_531)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_534),
.Y(n_533)
);

INVx2_ASAP7_75t_L g534 ( 
.A(n_535),
.Y(n_534)
);

INVx1_ASAP7_75t_SL g536 ( 
.A(n_537),
.Y(n_536)
);

INVxp67_ASAP7_75t_L g538 ( 
.A(n_539),
.Y(n_538)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_541),
.Y(n_540)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_543),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_544),
.Y(n_543)
);

BUFx3_ASAP7_75t_L g544 ( 
.A(n_545),
.Y(n_544)
);

INVx2_ASAP7_75t_L g545 ( 
.A(n_546),
.Y(n_545)
);

INVx2_ASAP7_75t_L g546 ( 
.A(n_547),
.Y(n_546)
);

XNOR2xp5_ASAP7_75t_L g548 ( 
.A(n_549),
.B(n_570),
.Y(n_548)
);

NOR2xp33_ASAP7_75t_L g613 ( 
.A(n_549),
.B(n_570),
.Y(n_613)
);

AOI21xp33_ASAP7_75t_L g549 ( 
.A1(n_550),
.A2(n_555),
.B(n_561),
.Y(n_549)
);

INVx1_ASAP7_75t_SL g550 ( 
.A(n_551),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_552),
.Y(n_551)
);

HB1xp67_ASAP7_75t_L g552 ( 
.A(n_553),
.Y(n_552)
);

INVx3_ASAP7_75t_L g553 ( 
.A(n_554),
.Y(n_553)
);

NOR2xp33_ASAP7_75t_L g555 ( 
.A(n_556),
.B(n_559),
.Y(n_555)
);

INVx2_ASAP7_75t_L g556 ( 
.A(n_557),
.Y(n_556)
);

INVx2_ASAP7_75t_L g557 ( 
.A(n_558),
.Y(n_557)
);

HB1xp67_ASAP7_75t_L g559 ( 
.A(n_560),
.Y(n_559)
);

AOI21xp5_ASAP7_75t_L g561 ( 
.A1(n_562),
.A2(n_566),
.B(n_569),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_563),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_564),
.Y(n_563)
);

INVx2_ASAP7_75t_L g564 ( 
.A(n_565),
.Y(n_564)
);

INVx2_ASAP7_75t_SL g566 ( 
.A(n_567),
.Y(n_566)
);

INVx3_ASAP7_75t_L g567 ( 
.A(n_568),
.Y(n_567)
);

INVx2_ASAP7_75t_SL g573 ( 
.A(n_574),
.Y(n_573)
);

BUFx6f_ASAP7_75t_L g574 ( 
.A(n_575),
.Y(n_574)
);

INVx4_ASAP7_75t_L g575 ( 
.A(n_576),
.Y(n_575)
);

OAI21xp5_ASAP7_75t_SL g577 ( 
.A1(n_578),
.A2(n_581),
.B(n_599),
.Y(n_577)
);

NOR2xp33_ASAP7_75t_L g578 ( 
.A(n_579),
.B(n_580),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_SL g599 ( 
.A(n_579),
.B(n_580),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_SL g581 ( 
.A(n_582),
.B(n_589),
.Y(n_581)
);

INVx2_ASAP7_75t_L g584 ( 
.A(n_585),
.Y(n_584)
);

INVx3_ASAP7_75t_SL g585 ( 
.A(n_586),
.Y(n_585)
);

BUFx6f_ASAP7_75t_L g586 ( 
.A(n_587),
.Y(n_586)
);

INVx3_ASAP7_75t_L g587 ( 
.A(n_588),
.Y(n_587)
);

NOR2xp33_ASAP7_75t_SL g589 ( 
.A(n_590),
.B(n_595),
.Y(n_589)
);

INVx2_ASAP7_75t_L g591 ( 
.A(n_592),
.Y(n_591)
);

INVx4_ASAP7_75t_L g592 ( 
.A(n_593),
.Y(n_592)
);

INVx2_ASAP7_75t_SL g593 ( 
.A(n_594),
.Y(n_593)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_596),
.Y(n_595)
);

INVx3_ASAP7_75t_L g596 ( 
.A(n_597),
.Y(n_596)
);

INVx2_ASAP7_75t_L g597 ( 
.A(n_598),
.Y(n_597)
);

AND2x2_ASAP7_75t_L g601 ( 
.A(n_602),
.B(n_604),
.Y(n_601)
);

OR2x2_ASAP7_75t_L g618 ( 
.A(n_602),
.B(n_604),
.Y(n_618)
);

MAJIxp5_ASAP7_75t_L g604 ( 
.A(n_605),
.B(n_606),
.C(n_610),
.Y(n_604)
);

XNOR2xp5_ASAP7_75t_L g614 ( 
.A(n_605),
.B(n_615),
.Y(n_614)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_607),
.Y(n_606)
);

OAI22xp5_ASAP7_75t_L g615 ( 
.A1(n_607),
.A2(n_608),
.B1(n_611),
.B2(n_616),
.Y(n_615)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_608),
.Y(n_607)
);

HB1xp67_ASAP7_75t_L g610 ( 
.A(n_611),
.Y(n_610)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_611),
.Y(n_616)
);

NOR2xp33_ASAP7_75t_L g612 ( 
.A(n_613),
.B(n_614),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_L g617 ( 
.A(n_613),
.B(n_614),
.Y(n_617)
);


endmodule