module fake_jpeg_10657_n_311 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_311);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_311;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_12),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_14),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_15),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_16),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_5),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_12),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_2),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_6),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_16),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_0),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_3),
.Y(n_32)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_4),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

BUFx6f_ASAP7_75t_SL g35 ( 
.A(n_1),
.Y(n_35)
);

INVx5_ASAP7_75t_L g36 ( 
.A(n_35),
.Y(n_36)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_36),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_35),
.Y(n_37)
);

OR2x2_ASAP7_75t_L g63 ( 
.A(n_37),
.B(n_38),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_35),
.Y(n_38)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_25),
.Y(n_39)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_39),
.Y(n_52)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_25),
.Y(n_40)
);

AND2x2_ASAP7_75t_L g57 ( 
.A(n_40),
.B(n_22),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_25),
.Y(n_41)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_41),
.Y(n_66)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_21),
.Y(n_42)
);

BUFx2_ASAP7_75t_L g62 ( 
.A(n_42),
.Y(n_62)
);

INVx6_ASAP7_75t_SL g43 ( 
.A(n_34),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_43),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_20),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_44),
.B(n_18),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_43),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_47),
.B(n_56),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_48),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_36),
.A2(n_33),
.B1(n_18),
.B2(n_19),
.Y(n_49)
);

AOI21xp5_ASAP7_75t_L g91 ( 
.A1(n_49),
.A2(n_60),
.B(n_58),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_37),
.A2(n_33),
.B1(n_30),
.B2(n_20),
.Y(n_50)
);

OAI21xp5_ASAP7_75t_L g87 ( 
.A1(n_50),
.A2(n_31),
.B(n_24),
.Y(n_87)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_51),
.B(n_61),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_43),
.Y(n_53)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_53),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_44),
.B(n_30),
.Y(n_54)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_54),
.Y(n_98)
);

AND2x2_ASAP7_75t_SL g55 ( 
.A(n_40),
.B(n_18),
.Y(n_55)
);

AND2x2_ASAP7_75t_L g88 ( 
.A(n_55),
.B(n_57),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_SL g56 ( 
.A(n_44),
.B(n_20),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_37),
.A2(n_33),
.B1(n_19),
.B2(n_22),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_L g71 ( 
.A1(n_58),
.A2(n_59),
.B1(n_29),
.B2(n_26),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_37),
.A2(n_26),
.B1(n_19),
.B2(n_22),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_36),
.A2(n_26),
.B1(n_29),
.B2(n_30),
.Y(n_60)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_36),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_43),
.Y(n_64)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_64),
.Y(n_67)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_42),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_65),
.B(n_38),
.Y(n_82)
);

OR2x2_ASAP7_75t_SL g68 ( 
.A(n_57),
.B(n_29),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_68),
.B(n_63),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_55),
.B(n_44),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_69),
.B(n_92),
.Y(n_104)
);

HB1xp67_ASAP7_75t_L g70 ( 
.A(n_46),
.Y(n_70)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_70),
.Y(n_114)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_71),
.Y(n_105)
);

INVx13_ASAP7_75t_L g72 ( 
.A(n_45),
.Y(n_72)
);

INVx11_ASAP7_75t_L g103 ( 
.A(n_72),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_L g74 ( 
.A1(n_48),
.A2(n_38),
.B1(n_39),
.B2(n_23),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_74),
.A2(n_100),
.B1(n_27),
.B2(n_28),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_62),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_75),
.B(n_78),
.Y(n_107)
);

CKINVDCx16_ASAP7_75t_R g78 ( 
.A(n_45),
.Y(n_78)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_45),
.Y(n_79)
);

INVx11_ASAP7_75t_L g130 ( 
.A(n_79),
.Y(n_130)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_62),
.Y(n_80)
);

CKINVDCx10_ASAP7_75t_R g126 ( 
.A(n_80),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_50),
.A2(n_38),
.B1(n_32),
.B2(n_23),
.Y(n_81)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_81),
.Y(n_120)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_82),
.Y(n_112)
);

AND2x2_ASAP7_75t_SL g83 ( 
.A(n_55),
.B(n_57),
.Y(n_83)
);

AND2x2_ASAP7_75t_L g111 ( 
.A(n_83),
.B(n_40),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_45),
.Y(n_84)
);

BUFx2_ASAP7_75t_L g109 ( 
.A(n_84),
.Y(n_109)
);

INVx8_ASAP7_75t_L g85 ( 
.A(n_46),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_85),
.A2(n_91),
.B1(n_95),
.B2(n_99),
.Y(n_106)
);

XNOR2x2_ASAP7_75t_L g86 ( 
.A(n_55),
.B(n_42),
.Y(n_86)
);

AOI21xp5_ASAP7_75t_L g128 ( 
.A1(n_86),
.A2(n_87),
.B(n_27),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_62),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_89),
.B(n_90),
.Y(n_123)
);

INVx13_ASAP7_75t_L g90 ( 
.A(n_53),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_56),
.B(n_17),
.Y(n_92)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_65),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_93),
.B(n_96),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_66),
.Y(n_94)
);

INVx13_ASAP7_75t_L g122 ( 
.A(n_94),
.Y(n_122)
);

AOI32xp33_ASAP7_75t_L g95 ( 
.A1(n_47),
.A2(n_52),
.A3(n_39),
.B1(n_66),
.B2(n_21),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_52),
.B(n_32),
.Y(n_96)
);

HB1xp67_ASAP7_75t_L g97 ( 
.A(n_51),
.Y(n_97)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_97),
.Y(n_116)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_53),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_L g100 ( 
.A1(n_61),
.A2(n_39),
.B1(n_28),
.B2(n_24),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_59),
.Y(n_101)
);

INVx13_ASAP7_75t_L g127 ( 
.A(n_101),
.Y(n_127)
);

CKINVDCx12_ASAP7_75t_R g108 ( 
.A(n_72),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_108),
.B(n_79),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_69),
.B(n_83),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_110),
.B(n_111),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_73),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_113),
.B(n_115),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_101),
.A2(n_52),
.B1(n_39),
.B2(n_40),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_117),
.A2(n_85),
.B1(n_99),
.B2(n_102),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_SL g135 ( 
.A(n_118),
.B(n_68),
.Y(n_135)
);

AND2x2_ASAP7_75t_L g119 ( 
.A(n_86),
.B(n_63),
.Y(n_119)
);

AOI21xp5_ASAP7_75t_L g143 ( 
.A1(n_119),
.A2(n_88),
.B(n_92),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_83),
.B(n_63),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_121),
.B(n_125),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_88),
.B(n_64),
.Y(n_125)
);

XOR2xp5_ASAP7_75t_L g147 ( 
.A(n_128),
.B(n_87),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_81),
.A2(n_39),
.B1(n_42),
.B2(n_31),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_129),
.A2(n_120),
.B1(n_105),
.B2(n_115),
.Y(n_152)
);

AND2x2_ASAP7_75t_SL g131 ( 
.A(n_125),
.B(n_77),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_L g166 ( 
.A1(n_131),
.A2(n_143),
.B(n_121),
.Y(n_166)
);

CKINVDCx16_ASAP7_75t_R g132 ( 
.A(n_123),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_132),
.B(n_135),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_133),
.A2(n_159),
.B1(n_114),
.B2(n_122),
.Y(n_178)
);

CKINVDCx14_ASAP7_75t_R g167 ( 
.A(n_134),
.Y(n_167)
);

CKINVDCx16_ASAP7_75t_R g138 ( 
.A(n_123),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_138),
.B(n_139),
.Y(n_171)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_107),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_SL g140 ( 
.A(n_118),
.B(n_77),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_140),
.B(n_146),
.Y(n_162)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_107),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_141),
.B(n_145),
.Y(n_183)
);

INVxp67_ASAP7_75t_L g144 ( 
.A(n_126),
.Y(n_144)
);

HB1xp67_ASAP7_75t_L g174 ( 
.A(n_144),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_112),
.B(n_76),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_104),
.B(n_88),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_SL g190 ( 
.A1(n_147),
.A2(n_155),
.B(n_21),
.Y(n_190)
);

INVx1_ASAP7_75t_SL g148 ( 
.A(n_126),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_148),
.B(n_149),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_109),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_124),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_150),
.B(n_151),
.Y(n_164)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_124),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_152),
.A2(n_105),
.B1(n_127),
.B2(n_128),
.Y(n_168)
);

HB1xp67_ASAP7_75t_L g153 ( 
.A(n_122),
.Y(n_153)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_153),
.Y(n_163)
);

OA22x2_ASAP7_75t_L g154 ( 
.A1(n_117),
.A2(n_91),
.B1(n_102),
.B2(n_67),
.Y(n_154)
);

OA22x2_ASAP7_75t_L g172 ( 
.A1(n_154),
.A2(n_127),
.B1(n_103),
.B2(n_111),
.Y(n_172)
);

INVxp67_ASAP7_75t_L g155 ( 
.A(n_106),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_112),
.B(n_98),
.Y(n_156)
);

CKINVDCx16_ASAP7_75t_R g187 ( 
.A(n_156),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_130),
.B(n_113),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_157),
.Y(n_189)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_129),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_158),
.B(n_111),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_127),
.A2(n_67),
.B1(n_90),
.B2(n_42),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_110),
.B(n_64),
.C(n_84),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_160),
.B(n_104),
.C(n_116),
.Y(n_170)
);

CKINVDCx16_ASAP7_75t_R g161 ( 
.A(n_109),
.Y(n_161)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_161),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_SL g205 ( 
.A1(n_166),
.A2(n_169),
.B(n_178),
.Y(n_205)
);

OAI32xp33_ASAP7_75t_L g211 ( 
.A1(n_168),
.A2(n_140),
.A3(n_135),
.B1(n_144),
.B2(n_148),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_170),
.B(n_176),
.C(n_138),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_172),
.A2(n_186),
.B1(n_188),
.B2(n_191),
.Y(n_214)
);

OAI21xp5_ASAP7_75t_L g173 ( 
.A1(n_143),
.A2(n_119),
.B(n_116),
.Y(n_173)
);

AOI21xp5_ASAP7_75t_L g207 ( 
.A1(n_173),
.A2(n_182),
.B(n_190),
.Y(n_207)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_159),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_175),
.B(n_177),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_136),
.B(n_119),
.C(n_114),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_133),
.Y(n_177)
);

BUFx2_ASAP7_75t_L g179 ( 
.A(n_161),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_179),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_137),
.B(n_93),
.Y(n_180)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_180),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_L g182 ( 
.A1(n_155),
.A2(n_34),
.B(n_17),
.Y(n_182)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_131),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_185),
.B(n_192),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_158),
.A2(n_122),
.B1(n_130),
.B2(n_103),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_154),
.A2(n_94),
.B1(n_41),
.B2(n_17),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_154),
.A2(n_41),
.B1(n_17),
.B2(n_80),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_131),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_154),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_193),
.B(n_152),
.Y(n_202)
);

NOR2x1_ASAP7_75t_L g195 ( 
.A(n_181),
.B(n_142),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_195),
.B(n_218),
.Y(n_237)
);

XOR2xp5_ASAP7_75t_L g198 ( 
.A(n_173),
.B(n_170),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_198),
.B(n_199),
.C(n_210),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_176),
.B(n_160),
.Y(n_199)
);

A2O1A1O1Ixp25_ASAP7_75t_L g200 ( 
.A1(n_166),
.A2(n_147),
.B(n_136),
.C(n_137),
.D(n_146),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_200),
.B(n_201),
.Y(n_223)
);

INVx13_ASAP7_75t_L g201 ( 
.A(n_179),
.Y(n_201)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_202),
.Y(n_222)
);

AOI21xp5_ASAP7_75t_SL g203 ( 
.A1(n_169),
.A2(n_139),
.B(n_141),
.Y(n_203)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_203),
.Y(n_235)
);

INVxp67_ASAP7_75t_L g206 ( 
.A(n_184),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_206),
.B(n_208),
.Y(n_231)
);

INVxp67_ASAP7_75t_L g208 ( 
.A(n_186),
.Y(n_208)
);

NAND3xp33_ASAP7_75t_L g209 ( 
.A(n_164),
.B(n_151),
.C(n_150),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_SL g229 ( 
.A(n_209),
.B(n_217),
.Y(n_229)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_211),
.Y(n_238)
);

XOR2xp5_ASAP7_75t_L g212 ( 
.A(n_190),
.B(n_108),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_212),
.B(n_215),
.C(n_219),
.Y(n_225)
);

AOI21xp5_ASAP7_75t_L g213 ( 
.A1(n_193),
.A2(n_149),
.B(n_109),
.Y(n_213)
);

AOI21xp5_ASAP7_75t_L g226 ( 
.A1(n_213),
.A2(n_220),
.B(n_192),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g215 ( 
.A(n_162),
.B(n_41),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_188),
.A2(n_41),
.B1(n_34),
.B2(n_15),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_216),
.A2(n_178),
.B1(n_189),
.B2(n_167),
.Y(n_240)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_164),
.Y(n_217)
);

OR2x2_ASAP7_75t_L g218 ( 
.A(n_171),
.B(n_0),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g219 ( 
.A(n_162),
.B(n_41),
.Y(n_219)
);

AOI21xp5_ASAP7_75t_L g220 ( 
.A1(n_185),
.A2(n_0),
.B(n_1),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_197),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_221),
.B(n_239),
.Y(n_248)
);

OAI21xp5_ASAP7_75t_SL g257 ( 
.A1(n_226),
.A2(n_220),
.B(n_214),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_199),
.B(n_180),
.C(n_182),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_227),
.B(n_230),
.C(n_232),
.Y(n_243)
);

HB1xp67_ASAP7_75t_L g228 ( 
.A(n_201),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_228),
.B(n_241),
.Y(n_247)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_198),
.B(n_191),
.Y(n_230)
);

XOR2xp5_ASAP7_75t_L g232 ( 
.A(n_212),
.B(n_183),
.Y(n_232)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_210),
.B(n_172),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_233),
.B(n_234),
.C(n_236),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_205),
.B(n_172),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_215),
.B(n_189),
.C(n_175),
.Y(n_236)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_203),
.Y(n_239)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_240),
.Y(n_244)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_194),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_219),
.B(n_172),
.C(n_163),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_242),
.B(n_207),
.C(n_214),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_222),
.B(n_196),
.Y(n_245)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_245),
.Y(n_264)
);

NOR2xp67_ASAP7_75t_SL g246 ( 
.A(n_226),
.B(n_195),
.Y(n_246)
);

CKINVDCx14_ASAP7_75t_R g268 ( 
.A(n_246),
.Y(n_268)
);

AO221x1_ASAP7_75t_L g249 ( 
.A1(n_231),
.A2(n_204),
.B1(n_163),
.B2(n_174),
.C(n_165),
.Y(n_249)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_249),
.Y(n_267)
);

A2O1A1O1Ixp25_ASAP7_75t_L g250 ( 
.A1(n_223),
.A2(n_238),
.B(n_234),
.C(n_200),
.D(n_230),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g262 ( 
.A(n_250),
.B(n_253),
.Y(n_262)
);

AOI21xp5_ASAP7_75t_L g252 ( 
.A1(n_235),
.A2(n_208),
.B(n_206),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_L g265 ( 
.A1(n_252),
.A2(n_258),
.B1(n_259),
.B2(n_225),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_225),
.B(n_224),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_254),
.B(n_260),
.C(n_242),
.Y(n_261)
);

NAND3xp33_ASAP7_75t_L g255 ( 
.A(n_237),
.B(n_211),
.C(n_187),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_255),
.B(n_256),
.Y(n_272)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_229),
.Y(n_256)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_257),
.Y(n_274)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_240),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_L g259 ( 
.A1(n_237),
.A2(n_216),
.B1(n_165),
.B2(n_218),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_236),
.B(n_1),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_261),
.B(n_263),
.C(n_251),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_253),
.B(n_224),
.C(n_227),
.Y(n_263)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_265),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_244),
.A2(n_233),
.B1(n_232),
.B2(n_4),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_L g282 ( 
.A1(n_266),
.A2(n_270),
.B1(n_6),
.B2(n_7),
.Y(n_282)
);

NOR2xp67_ASAP7_75t_L g269 ( 
.A(n_248),
.B(n_2),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_269),
.B(n_257),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_252),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_243),
.B(n_3),
.C(n_5),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_271),
.B(n_273),
.C(n_8),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_243),
.B(n_6),
.C(n_7),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_275),
.B(n_277),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_276),
.B(n_278),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_SL g277 ( 
.A(n_266),
.B(n_250),
.Y(n_277)
);

AOI21xp5_ASAP7_75t_SL g278 ( 
.A1(n_274),
.A2(n_245),
.B(n_260),
.Y(n_278)
);

INVxp67_ASAP7_75t_L g279 ( 
.A(n_270),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_279),
.B(n_280),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_261),
.B(n_254),
.C(n_251),
.Y(n_280)
);

XOR2xp5_ASAP7_75t_L g281 ( 
.A(n_262),
.B(n_247),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_281),
.B(n_282),
.Y(n_294)
);

XOR2xp5_ASAP7_75t_L g283 ( 
.A(n_263),
.B(n_8),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_283),
.B(n_284),
.Y(n_291)
);

XOR2xp5_ASAP7_75t_L g284 ( 
.A(n_262),
.B(n_273),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_286),
.B(n_9),
.Y(n_293)
);

BUFx24_ASAP7_75t_SL g287 ( 
.A(n_285),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_287),
.B(n_293),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_279),
.A2(n_268),
.B1(n_264),
.B2(n_267),
.Y(n_289)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_289),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_278),
.B(n_272),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_295),
.B(n_9),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_294),
.B(n_281),
.Y(n_296)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_296),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_292),
.B(n_271),
.Y(n_297)
);

XOR2x2_ASAP7_75t_L g306 ( 
.A(n_297),
.B(n_296),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_SL g298 ( 
.A(n_290),
.B(n_277),
.Y(n_298)
);

AOI322xp5_ASAP7_75t_L g305 ( 
.A1(n_298),
.A2(n_291),
.A3(n_292),
.B1(n_13),
.B2(n_14),
.C1(n_10),
.C2(n_11),
.Y(n_305)
);

AOI21xp5_ASAP7_75t_L g303 ( 
.A1(n_301),
.A2(n_302),
.B(n_10),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_288),
.B(n_9),
.Y(n_302)
);

NAND4xp25_ASAP7_75t_SL g308 ( 
.A(n_303),
.B(n_11),
.C(n_13),
.D(n_300),
.Y(n_308)
);

AOI21xp5_ASAP7_75t_L g307 ( 
.A1(n_305),
.A2(n_306),
.B(n_299),
.Y(n_307)
);

AOI21xp5_ASAP7_75t_L g309 ( 
.A1(n_307),
.A2(n_308),
.B(n_304),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_309),
.B(n_11),
.Y(n_310)
);

XOR2xp5_ASAP7_75t_L g311 ( 
.A(n_310),
.B(n_13),
.Y(n_311)
);


endmodule