module fake_jpeg_17096_n_143 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_143);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_143;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_93;
wire n_91;
wire n_138;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_39),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_13),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_17),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_6),
.Y(n_46)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_9),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_7),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_33),
.Y(n_49)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_35),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_8),
.Y(n_51)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_28),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_4),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_4),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_3),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_21),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_2),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_14),
.Y(n_58)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_3),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_18),
.Y(n_60)
);

INVx11_ASAP7_75t_L g61 ( 
.A(n_52),
.Y(n_61)
);

INVx5_ASAP7_75t_L g83 ( 
.A(n_61),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_44),
.Y(n_62)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_62),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_44),
.Y(n_63)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_63),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_59),
.B(n_49),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_64),
.B(n_49),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_51),
.Y(n_65)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_65),
.Y(n_84)
);

INVx11_ASAP7_75t_L g66 ( 
.A(n_52),
.Y(n_66)
);

BUFx10_ASAP7_75t_L g74 ( 
.A(n_66),
.Y(n_74)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_49),
.Y(n_67)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_67),
.Y(n_80)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_54),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_68),
.B(n_53),
.Y(n_75)
);

INVx13_ASAP7_75t_L g70 ( 
.A(n_67),
.Y(n_70)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_70),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_SL g71 ( 
.A(n_68),
.B(n_57),
.Y(n_71)
);

AND2x2_ASAP7_75t_L g96 ( 
.A(n_71),
.B(n_73),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_64),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_75),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_66),
.B(n_48),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_76),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_61),
.B(n_46),
.Y(n_77)
);

AND2x4_ASAP7_75t_L g95 ( 
.A(n_77),
.B(n_78),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_65),
.B(n_55),
.Y(n_78)
);

INVx6_ASAP7_75t_SL g79 ( 
.A(n_62),
.Y(n_79)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_79),
.Y(n_91)
);

XOR2xp5_ASAP7_75t_L g86 ( 
.A(n_81),
.B(n_50),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_63),
.A2(n_50),
.B1(n_47),
.B2(n_51),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_82),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_97)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_69),
.Y(n_85)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_85),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_86),
.B(n_74),
.Y(n_110)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_72),
.Y(n_87)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_87),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_82),
.A2(n_60),
.B1(n_58),
.B2(n_56),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_89),
.A2(n_90),
.B1(n_92),
.B2(n_98),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_84),
.A2(n_45),
.B1(n_43),
.B2(n_26),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_83),
.A2(n_24),
.B1(n_41),
.B2(n_40),
.Y(n_92)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_83),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_93),
.B(n_94),
.Y(n_109)
);

HB1xp67_ASAP7_75t_L g94 ( 
.A(n_74),
.Y(n_94)
);

OA22x2_ASAP7_75t_L g106 ( 
.A1(n_97),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_80),
.A2(n_0),
.B1(n_1),
.B2(n_5),
.Y(n_98)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_80),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_99),
.Y(n_108)
);

CKINVDCx14_ASAP7_75t_R g103 ( 
.A(n_90),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_103),
.B(n_111),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_88),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_104),
.B(n_110),
.Y(n_113)
);

AOI21x1_ASAP7_75t_L g105 ( 
.A1(n_95),
.A2(n_70),
.B(n_74),
.Y(n_105)
);

MAJx2_ASAP7_75t_L g116 ( 
.A(n_105),
.B(n_101),
.C(n_100),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_106),
.A2(n_95),
.B1(n_92),
.B2(n_91),
.Y(n_115)
);

BUFx3_ASAP7_75t_L g111 ( 
.A(n_94),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_103),
.B(n_96),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_114),
.B(n_115),
.Y(n_121)
);

AOI21xp5_ASAP7_75t_SL g122 ( 
.A1(n_116),
.A2(n_118),
.B(n_109),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_102),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_117),
.B(n_112),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_119),
.B(n_16),
.Y(n_128)
);

AOI21xp5_ASAP7_75t_L g120 ( 
.A1(n_118),
.A2(n_113),
.B(n_109),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_120),
.A2(n_10),
.B1(n_11),
.B2(n_15),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_122),
.A2(n_121),
.B1(n_106),
.B2(n_12),
.Y(n_124)
);

XOR2xp5_ASAP7_75t_L g123 ( 
.A(n_113),
.B(n_107),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_123),
.B(n_106),
.C(n_108),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_124),
.B(n_127),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_119),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_125),
.B(n_126),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_128),
.B(n_19),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_SL g132 ( 
.A(n_131),
.B(n_128),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_L g134 ( 
.A(n_132),
.B(n_133),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_129),
.A2(n_20),
.B1(n_22),
.B2(n_23),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_134),
.B(n_130),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_135),
.B(n_42),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_136),
.B(n_25),
.C(n_27),
.Y(n_137)
);

NAND3xp33_ASAP7_75t_L g138 ( 
.A(n_137),
.B(n_29),
.C(n_30),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_138),
.B(n_31),
.C(n_32),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_139),
.Y(n_140)
);

OAI21x1_ASAP7_75t_L g141 ( 
.A1(n_140),
.A2(n_34),
.B(n_36),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_141),
.B(n_37),
.Y(n_142)
);

XNOR2xp5_ASAP7_75t_L g143 ( 
.A(n_142),
.B(n_38),
.Y(n_143)
);


endmodule