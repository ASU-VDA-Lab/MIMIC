module fake_jpeg_13184_n_480 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_480);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_480;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx10_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_2),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

BUFx12_ASAP7_75t_L g21 ( 
.A(n_16),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_9),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_0),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_14),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_8),
.Y(n_26)
);

BUFx4f_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

BUFx24_ASAP7_75t_L g29 ( 
.A(n_15),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_16),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_13),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_8),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_11),
.Y(n_33)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_8),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_17),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_15),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_0),
.Y(n_37)
);

BUFx5_ASAP7_75t_L g38 ( 
.A(n_10),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_10),
.Y(n_39)
);

BUFx12_ASAP7_75t_L g40 ( 
.A(n_10),
.Y(n_40)
);

BUFx16f_ASAP7_75t_L g41 ( 
.A(n_2),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_1),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_10),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_0),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_17),
.Y(n_45)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_1),
.Y(n_46)
);

INVx11_ASAP7_75t_L g47 ( 
.A(n_3),
.Y(n_47)
);

BUFx5_ASAP7_75t_L g48 ( 
.A(n_4),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_14),
.Y(n_49)
);

CKINVDCx16_ASAP7_75t_R g50 ( 
.A(n_15),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_14),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_9),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_5),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_5),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_3),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_7),
.Y(n_56)
);

CKINVDCx16_ASAP7_75t_R g57 ( 
.A(n_29),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_57),
.B(n_77),
.Y(n_121)
);

INVx6_ASAP7_75t_SL g58 ( 
.A(n_29),
.Y(n_58)
);

BUFx12f_ASAP7_75t_L g156 ( 
.A(n_58),
.Y(n_156)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_45),
.Y(n_59)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_59),
.Y(n_131)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_45),
.Y(n_60)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_60),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_25),
.B(n_17),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_61),
.B(n_63),
.Y(n_128)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_22),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g148 ( 
.A(n_62),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_25),
.B(n_16),
.Y(n_63)
);

INVx5_ASAP7_75t_L g64 ( 
.A(n_29),
.Y(n_64)
);

INVx2_ASAP7_75t_SL g129 ( 
.A(n_64),
.Y(n_129)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_32),
.Y(n_65)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_65),
.Y(n_170)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_33),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_66),
.Y(n_118)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_20),
.Y(n_67)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_67),
.Y(n_160)
);

INVx8_ASAP7_75t_L g68 ( 
.A(n_29),
.Y(n_68)
);

INVx5_ASAP7_75t_L g124 ( 
.A(n_68),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_33),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_69),
.Y(n_119)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_28),
.Y(n_70)
);

INVx5_ASAP7_75t_L g138 ( 
.A(n_70),
.Y(n_138)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_41),
.Y(n_71)
);

INVx3_ASAP7_75t_L g137 ( 
.A(n_71),
.Y(n_137)
);

BUFx12f_ASAP7_75t_L g72 ( 
.A(n_28),
.Y(n_72)
);

INVx5_ASAP7_75t_L g163 ( 
.A(n_72),
.Y(n_163)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_22),
.Y(n_73)
);

INVx3_ASAP7_75t_L g157 ( 
.A(n_73),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_33),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_74),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_53),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_75),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_30),
.B(n_13),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_76),
.B(n_79),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_21),
.Y(n_77)
);

HB1xp67_ASAP7_75t_L g78 ( 
.A(n_20),
.Y(n_78)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_78),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_30),
.B(n_13),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_53),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g165 ( 
.A(n_80),
.Y(n_165)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_22),
.Y(n_81)
);

INVx3_ASAP7_75t_L g172 ( 
.A(n_81),
.Y(n_172)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_32),
.Y(n_82)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_82),
.Y(n_177)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_53),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g185 ( 
.A(n_83),
.Y(n_185)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_56),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g188 ( 
.A(n_84),
.Y(n_188)
);

INVx6_ASAP7_75t_L g85 ( 
.A(n_56),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g189 ( 
.A(n_85),
.Y(n_189)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_27),
.Y(n_86)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_86),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_21),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_87),
.B(n_88),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_21),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_21),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_89),
.B(n_93),
.Y(n_126)
);

BUFx3_ASAP7_75t_L g90 ( 
.A(n_22),
.Y(n_90)
);

INVx4_ASAP7_75t_L g132 ( 
.A(n_90),
.Y(n_132)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_27),
.Y(n_91)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_91),
.Y(n_173)
);

INVx11_ASAP7_75t_L g92 ( 
.A(n_47),
.Y(n_92)
);

BUFx10_ASAP7_75t_L g125 ( 
.A(n_92),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_40),
.Y(n_93)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_27),
.Y(n_94)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_94),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_31),
.B(n_0),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_95),
.B(n_106),
.Y(n_152)
);

INVx6_ASAP7_75t_L g96 ( 
.A(n_56),
.Y(n_96)
);

INVx6_ASAP7_75t_L g123 ( 
.A(n_96),
.Y(n_123)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_37),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_97),
.B(n_98),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_40),
.Y(n_98)
);

INVx4_ASAP7_75t_SL g99 ( 
.A(n_18),
.Y(n_99)
);

INVx4_ASAP7_75t_L g144 ( 
.A(n_99),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_27),
.Y(n_100)
);

INVx8_ASAP7_75t_L g143 ( 
.A(n_100),
.Y(n_143)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_41),
.Y(n_101)
);

INVx3_ASAP7_75t_L g179 ( 
.A(n_101),
.Y(n_179)
);

HAxp5_ASAP7_75t_SL g102 ( 
.A(n_18),
.B(n_1),
.CON(n_102),
.SN(n_102)
);

AND2x2_ASAP7_75t_L g176 ( 
.A(n_102),
.B(n_103),
.Y(n_176)
);

AND2x2_ASAP7_75t_L g103 ( 
.A(n_34),
.B(n_1),
.Y(n_103)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_41),
.Y(n_104)
);

INVx2_ASAP7_75t_SL g130 ( 
.A(n_104),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_46),
.Y(n_105)
);

INVx4_ASAP7_75t_L g139 ( 
.A(n_105),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_31),
.B(n_2),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_46),
.Y(n_107)
);

INVx4_ASAP7_75t_L g146 ( 
.A(n_107),
.Y(n_146)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_37),
.Y(n_108)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_108),
.Y(n_181)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_34),
.Y(n_109)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_109),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_36),
.B(n_50),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_110),
.B(n_113),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_36),
.B(n_2),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_111),
.B(n_117),
.Y(n_159)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_42),
.Y(n_112)
);

INVx4_ASAP7_75t_L g151 ( 
.A(n_112),
.Y(n_151)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_43),
.Y(n_113)
);

INVx8_ASAP7_75t_L g114 ( 
.A(n_38),
.Y(n_114)
);

INVx4_ASAP7_75t_L g174 ( 
.A(n_114),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_50),
.B(n_3),
.Y(n_115)
);

AND2x2_ASAP7_75t_L g178 ( 
.A(n_115),
.B(n_4),
.Y(n_178)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_46),
.Y(n_116)
);

INVx4_ASAP7_75t_L g190 ( 
.A(n_116),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_40),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_67),
.A2(n_35),
.B1(n_51),
.B2(n_49),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_134),
.A2(n_171),
.B1(n_129),
.B2(n_163),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_85),
.A2(n_49),
.B1(n_35),
.B2(n_51),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g220 ( 
.A1(n_135),
.A2(n_136),
.B1(n_140),
.B2(n_141),
.Y(n_220)
);

AOI22xp33_ASAP7_75t_SL g136 ( 
.A1(n_58),
.A2(n_55),
.B1(n_39),
.B2(n_18),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_103),
.A2(n_49),
.B1(n_35),
.B2(n_51),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_96),
.A2(n_26),
.B1(n_52),
.B2(n_24),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_109),
.A2(n_26),
.B1(n_52),
.B2(n_24),
.Y(n_142)
);

OAI22xp33_ASAP7_75t_L g194 ( 
.A1(n_142),
.A2(n_145),
.B1(n_153),
.B2(n_158),
.Y(n_194)
);

AOI22xp33_ASAP7_75t_L g145 ( 
.A1(n_66),
.A2(n_18),
.B1(n_54),
.B2(n_44),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_92),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_147),
.B(n_149),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_71),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_101),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_150),
.B(n_186),
.Y(n_207)
);

AOI22xp33_ASAP7_75t_L g153 ( 
.A1(n_69),
.A2(n_18),
.B1(n_54),
.B2(n_44),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_SL g154 ( 
.A1(n_68),
.A2(n_55),
.B1(n_39),
.B2(n_47),
.Y(n_154)
);

AOI22xp33_ASAP7_75t_SL g193 ( 
.A1(n_154),
.A2(n_175),
.B1(n_187),
.B2(n_72),
.Y(n_193)
);

AOI22xp33_ASAP7_75t_L g158 ( 
.A1(n_74),
.A2(n_43),
.B1(n_19),
.B2(n_23),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_86),
.B(n_23),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_161),
.B(n_167),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_75),
.A2(n_19),
.B1(n_42),
.B2(n_38),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_166),
.B(n_129),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_91),
.B(n_42),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_80),
.A2(n_42),
.B1(n_48),
.B2(n_40),
.Y(n_171)
);

AOI22xp33_ASAP7_75t_SL g175 ( 
.A1(n_70),
.A2(n_48),
.B1(n_5),
.B2(n_6),
.Y(n_175)
);

AOI21xp33_ASAP7_75t_L g234 ( 
.A1(n_178),
.A2(n_12),
.B(n_121),
.Y(n_234)
);

INVx4_ASAP7_75t_L g182 ( 
.A(n_99),
.Y(n_182)
);

HB1xp67_ASAP7_75t_L g213 ( 
.A(n_182),
.Y(n_213)
);

BUFx10_ASAP7_75t_L g183 ( 
.A(n_64),
.Y(n_183)
);

CKINVDCx6p67_ASAP7_75t_R g251 ( 
.A(n_183),
.Y(n_251)
);

NOR2x1_ASAP7_75t_L g186 ( 
.A(n_73),
.B(n_4),
.Y(n_186)
);

AOI22xp33_ASAP7_75t_SL g187 ( 
.A1(n_114),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_187)
);

NAND3xp33_ASAP7_75t_L g191 ( 
.A(n_152),
.B(n_104),
.C(n_102),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_191),
.B(n_211),
.Y(n_253)
);

AOI22xp33_ASAP7_75t_SL g255 ( 
.A1(n_193),
.A2(n_198),
.B1(n_214),
.B2(n_246),
.Y(n_255)
);

AOI22xp33_ASAP7_75t_SL g195 ( 
.A1(n_174),
.A2(n_116),
.B1(n_107),
.B2(n_105),
.Y(n_195)
);

INVxp67_ASAP7_75t_L g288 ( 
.A(n_195),
.Y(n_288)
);

BUFx3_ASAP7_75t_L g196 ( 
.A(n_156),
.Y(n_196)
);

INVx5_ASAP7_75t_L g277 ( 
.A(n_196),
.Y(n_277)
);

AOI22xp33_ASAP7_75t_SL g197 ( 
.A1(n_174),
.A2(n_81),
.B1(n_112),
.B2(n_72),
.Y(n_197)
);

INVxp67_ASAP7_75t_L g298 ( 
.A(n_197),
.Y(n_298)
);

AOI22xp33_ASAP7_75t_SL g198 ( 
.A1(n_170),
.A2(n_62),
.B1(n_90),
.B2(n_94),
.Y(n_198)
);

INVx1_ASAP7_75t_SL g200 ( 
.A(n_156),
.Y(n_200)
);

AND2x2_ASAP7_75t_L g267 ( 
.A(n_200),
.B(n_206),
.Y(n_267)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_131),
.Y(n_201)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_201),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_155),
.B(n_6),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_SL g263 ( 
.A(n_202),
.B(n_205),
.Y(n_263)
);

INVx5_ASAP7_75t_L g203 ( 
.A(n_156),
.Y(n_203)
);

INVx3_ASAP7_75t_L g258 ( 
.A(n_203),
.Y(n_258)
);

INVx3_ASAP7_75t_L g204 ( 
.A(n_139),
.Y(n_204)
);

INVx3_ASAP7_75t_L g275 ( 
.A(n_204),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_128),
.B(n_6),
.Y(n_205)
);

INVx1_ASAP7_75t_SL g206 ( 
.A(n_183),
.Y(n_206)
);

INVx6_ASAP7_75t_L g208 ( 
.A(n_118),
.Y(n_208)
);

INVx3_ASAP7_75t_L g286 ( 
.A(n_208),
.Y(n_286)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_169),
.Y(n_209)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_209),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_162),
.B(n_100),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_SL g269 ( 
.A(n_210),
.B(n_212),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_127),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_159),
.B(n_7),
.Y(n_212)
);

AOI22xp33_ASAP7_75t_SL g214 ( 
.A1(n_177),
.A2(n_83),
.B1(n_84),
.B2(n_11),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_164),
.Y(n_215)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_215),
.Y(n_260)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_173),
.Y(n_216)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_216),
.Y(n_261)
);

AND2x2_ASAP7_75t_L g217 ( 
.A(n_176),
.B(n_7),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_217),
.B(n_223),
.C(n_241),
.Y(n_272)
);

BUFx2_ASAP7_75t_SL g218 ( 
.A(n_183),
.Y(n_218)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_218),
.Y(n_299)
);

INVx4_ASAP7_75t_L g219 ( 
.A(n_132),
.Y(n_219)
);

INVx2_ASAP7_75t_L g287 ( 
.A(n_219),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_126),
.B(n_7),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_221),
.B(n_228),
.Y(n_279)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_180),
.Y(n_222)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_222),
.Y(n_271)
);

AND2x2_ASAP7_75t_L g223 ( 
.A(n_176),
.B(n_8),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_181),
.Y(n_224)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_224),
.Y(n_283)
);

AOI22xp33_ASAP7_75t_L g225 ( 
.A1(n_158),
.A2(n_12),
.B1(n_145),
.B2(n_153),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_L g266 ( 
.A1(n_225),
.A2(n_243),
.B1(n_244),
.B2(n_248),
.Y(n_266)
);

BUFx6f_ASAP7_75t_L g226 ( 
.A(n_118),
.Y(n_226)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_226),
.Y(n_264)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_160),
.Y(n_227)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_227),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_122),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_184),
.Y(n_229)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_229),
.Y(n_292)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_123),
.Y(n_230)
);

AND2x2_ASAP7_75t_L g289 ( 
.A(n_230),
.B(n_233),
.Y(n_289)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_130),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_231),
.B(n_232),
.Y(n_280)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_130),
.Y(n_232)
);

INVx3_ASAP7_75t_L g233 ( 
.A(n_139),
.Y(n_233)
);

OR2x6_ASAP7_75t_L g285 ( 
.A(n_234),
.B(n_125),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_178),
.B(n_12),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_235),
.B(n_238),
.Y(n_268)
);

BUFx2_ASAP7_75t_L g236 ( 
.A(n_124),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_236),
.B(n_240),
.Y(n_284)
);

INVx13_ASAP7_75t_L g237 ( 
.A(n_144),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_237),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_186),
.B(n_12),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_168),
.B(n_123),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_239),
.B(n_247),
.Y(n_276)
);

INVx3_ASAP7_75t_L g240 ( 
.A(n_146),
.Y(n_240)
);

AND2x2_ASAP7_75t_SL g241 ( 
.A(n_157),
.B(n_172),
.Y(n_241)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_151),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_242),
.Y(n_278)
);

OR2x2_ASAP7_75t_L g244 ( 
.A(n_136),
.B(n_179),
.Y(n_244)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_189),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g296 ( 
.A(n_245),
.Y(n_296)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_137),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_143),
.Y(n_247)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_189),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_249),
.B(n_250),
.Y(n_281)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_143),
.Y(n_250)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_119),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_252),
.B(n_120),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_243),
.A2(n_154),
.B1(n_175),
.B2(n_187),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_254),
.A2(n_274),
.B1(n_295),
.B2(n_241),
.Y(n_307)
);

AND2x4_ASAP7_75t_SL g256 ( 
.A(n_199),
.B(n_148),
.Y(n_256)
);

AND2x2_ASAP7_75t_L g304 ( 
.A(n_256),
.B(n_241),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_220),
.A2(n_146),
.B1(n_190),
.B2(n_119),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_L g301 ( 
.A1(n_270),
.A2(n_291),
.B1(n_297),
.B2(n_252),
.Y(n_301)
);

AOI21xp5_ASAP7_75t_L g273 ( 
.A1(n_244),
.A2(n_138),
.B(n_125),
.Y(n_273)
);

OAI21xp5_ASAP7_75t_L g311 ( 
.A1(n_273),
.A2(n_285),
.B(n_236),
.Y(n_311)
);

OAI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_194),
.A2(n_190),
.B1(n_120),
.B2(n_133),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_SL g282 ( 
.A(n_217),
.B(n_125),
.C(n_148),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_282),
.B(n_206),
.C(n_213),
.Y(n_314)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_290),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_L g291 ( 
.A1(n_194),
.A2(n_239),
.B1(n_238),
.B2(n_217),
.Y(n_291)
);

NOR2x1_ASAP7_75t_SL g293 ( 
.A(n_207),
.B(n_133),
.Y(n_293)
);

OR2x4_ASAP7_75t_L g321 ( 
.A(n_293),
.B(n_251),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_235),
.B(n_165),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_294),
.B(n_196),
.Y(n_317)
);

OAI22xp5_ASAP7_75t_SL g295 ( 
.A1(n_192),
.A2(n_230),
.B1(n_185),
.B2(n_188),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g297 ( 
.A1(n_223),
.A2(n_165),
.B1(n_185),
.B2(n_188),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_L g338 ( 
.A1(n_301),
.A2(n_306),
.B1(n_318),
.B2(n_329),
.Y(n_338)
);

CKINVDCx20_ASAP7_75t_R g302 ( 
.A(n_281),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_302),
.B(n_308),
.Y(n_341)
);

BUFx3_ASAP7_75t_L g303 ( 
.A(n_258),
.Y(n_303)
);

BUFx3_ASAP7_75t_L g343 ( 
.A(n_303),
.Y(n_343)
);

OAI21xp5_ASAP7_75t_SL g363 ( 
.A1(n_304),
.A2(n_311),
.B(n_314),
.Y(n_363)
);

INVxp67_ASAP7_75t_L g305 ( 
.A(n_267),
.Y(n_305)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_305),
.Y(n_344)
);

OAI22xp5_ASAP7_75t_SL g306 ( 
.A1(n_291),
.A2(n_249),
.B1(n_245),
.B2(n_208),
.Y(n_306)
);

AND2x2_ASAP7_75t_L g337 ( 
.A(n_307),
.B(n_331),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_SL g308 ( 
.A(n_276),
.B(n_223),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_L g309 ( 
.A1(n_266),
.A2(n_227),
.B1(n_233),
.B2(n_240),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_L g340 ( 
.A1(n_309),
.A2(n_310),
.B1(n_312),
.B2(n_315),
.Y(n_340)
);

AOI22xp5_ASAP7_75t_L g310 ( 
.A1(n_274),
.A2(n_204),
.B1(n_209),
.B2(n_222),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_L g312 ( 
.A1(n_254),
.A2(n_216),
.B1(n_226),
.B2(n_242),
.Y(n_312)
);

INVx5_ASAP7_75t_L g313 ( 
.A(n_258),
.Y(n_313)
);

BUFx2_ASAP7_75t_L g342 ( 
.A(n_313),
.Y(n_342)
);

AOI22xp5_ASAP7_75t_L g315 ( 
.A1(n_276),
.A2(n_219),
.B1(n_251),
.B2(n_203),
.Y(n_315)
);

BUFx5_ASAP7_75t_L g316 ( 
.A(n_299),
.Y(n_316)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_316),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_317),
.B(n_324),
.Y(n_352)
);

OAI22xp5_ASAP7_75t_SL g318 ( 
.A1(n_270),
.A2(n_251),
.B1(n_200),
.B2(n_237),
.Y(n_318)
);

INVxp67_ASAP7_75t_L g319 ( 
.A(n_267),
.Y(n_319)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_319),
.Y(n_353)
);

AOI22xp5_ASAP7_75t_L g320 ( 
.A1(n_288),
.A2(n_251),
.B1(n_295),
.B2(n_268),
.Y(n_320)
);

OAI22xp5_ASAP7_75t_L g346 ( 
.A1(n_320),
.A2(n_326),
.B1(n_328),
.B2(n_282),
.Y(n_346)
);

CKINVDCx14_ASAP7_75t_R g358 ( 
.A(n_321),
.Y(n_358)
);

OAI21xp5_ASAP7_75t_L g322 ( 
.A1(n_285),
.A2(n_273),
.B(n_298),
.Y(n_322)
);

OAI21xp5_ASAP7_75t_L g339 ( 
.A1(n_322),
.A2(n_323),
.B(n_336),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_SL g323 ( 
.A(n_253),
.B(n_268),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_294),
.B(n_256),
.Y(n_324)
);

INVxp33_ASAP7_75t_SL g325 ( 
.A(n_284),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_325),
.B(n_330),
.Y(n_355)
);

AOI22xp5_ASAP7_75t_L g326 ( 
.A1(n_288),
.A2(n_256),
.B1(n_272),
.B2(n_298),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_279),
.B(n_269),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g361 ( 
.A(n_327),
.Y(n_361)
);

AOI22xp5_ASAP7_75t_L g328 ( 
.A1(n_272),
.A2(n_293),
.B1(n_285),
.B2(n_290),
.Y(n_328)
);

OAI22xp5_ASAP7_75t_L g329 ( 
.A1(n_255),
.A2(n_285),
.B1(n_297),
.B2(n_281),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_280),
.B(n_285),
.Y(n_330)
);

AND2x2_ASAP7_75t_L g331 ( 
.A(n_289),
.B(n_267),
.Y(n_331)
);

XOR2xp5_ASAP7_75t_L g332 ( 
.A(n_259),
.B(n_260),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_L g345 ( 
.A(n_332),
.B(n_271),
.C(n_283),
.Y(n_345)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_292),
.Y(n_333)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_333),
.Y(n_354)
);

OAI22xp33_ASAP7_75t_SL g334 ( 
.A1(n_292),
.A2(n_286),
.B1(n_275),
.B2(n_264),
.Y(n_334)
);

AOI22xp5_ASAP7_75t_L g351 ( 
.A1(n_334),
.A2(n_265),
.B1(n_299),
.B2(n_275),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_278),
.B(n_296),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_335),
.B(n_257),
.Y(n_357)
);

NOR2xp33_ASAP7_75t_SL g336 ( 
.A(n_263),
.B(n_262),
.Y(n_336)
);

XOR2xp5_ASAP7_75t_L g381 ( 
.A(n_345),
.B(n_363),
.Y(n_381)
);

INVxp67_ASAP7_75t_L g378 ( 
.A(n_346),
.Y(n_378)
);

XOR2xp5_ASAP7_75t_L g347 ( 
.A(n_328),
.B(n_289),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_L g386 ( 
.A(n_347),
.B(n_349),
.C(n_356),
.Y(n_386)
);

OAI22xp5_ASAP7_75t_SL g348 ( 
.A1(n_307),
.A2(n_264),
.B1(n_286),
.B2(n_265),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_348),
.B(n_357),
.Y(n_387)
);

XOR2xp5_ASAP7_75t_L g349 ( 
.A(n_324),
.B(n_289),
.Y(n_349)
);

AND2x2_ASAP7_75t_L g368 ( 
.A(n_351),
.B(n_318),
.Y(n_368)
);

MAJIxp5_ASAP7_75t_L g356 ( 
.A(n_330),
.B(n_257),
.C(n_261),
.Y(n_356)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_335),
.Y(n_359)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_359),
.Y(n_367)
);

OAI22xp5_ASAP7_75t_SL g360 ( 
.A1(n_302),
.A2(n_261),
.B1(n_287),
.B2(n_277),
.Y(n_360)
);

AOI22xp5_ASAP7_75t_SL g372 ( 
.A1(n_360),
.A2(n_365),
.B1(n_306),
.B2(n_305),
.Y(n_372)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_333),
.Y(n_362)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_362),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_300),
.B(n_287),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_SL g377 ( 
.A(n_364),
.B(n_332),
.Y(n_377)
);

OAI22xp5_ASAP7_75t_L g365 ( 
.A1(n_312),
.A2(n_277),
.B1(n_320),
.B2(n_300),
.Y(n_365)
);

CKINVDCx20_ASAP7_75t_R g366 ( 
.A(n_357),
.Y(n_366)
);

NOR2xp33_ASAP7_75t_L g403 ( 
.A(n_366),
.B(n_371),
.Y(n_403)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_368),
.Y(n_400)
);

AOI22x1_ASAP7_75t_L g369 ( 
.A1(n_337),
.A2(n_329),
.B1(n_321),
.B2(n_301),
.Y(n_369)
);

OAI22xp33_ASAP7_75t_SL g394 ( 
.A1(n_369),
.A2(n_372),
.B1(n_337),
.B2(n_365),
.Y(n_394)
);

OAI22xp5_ASAP7_75t_L g370 ( 
.A1(n_338),
.A2(n_326),
.B1(n_309),
.B2(n_311),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_370),
.B(n_373),
.Y(n_391)
);

CKINVDCx20_ASAP7_75t_R g371 ( 
.A(n_364),
.Y(n_371)
);

OAI22xp5_ASAP7_75t_SL g373 ( 
.A1(n_338),
.A2(n_322),
.B1(n_317),
.B2(n_310),
.Y(n_373)
);

INVx2_ASAP7_75t_L g374 ( 
.A(n_354),
.Y(n_374)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_374),
.Y(n_406)
);

NOR2xp33_ASAP7_75t_L g375 ( 
.A(n_361),
.B(n_336),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_L g410 ( 
.A(n_375),
.B(n_380),
.Y(n_410)
);

OAI22xp5_ASAP7_75t_L g376 ( 
.A1(n_359),
.A2(n_315),
.B1(n_323),
.B2(n_319),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_376),
.B(n_377),
.Y(n_396)
);

AOI21xp5_ASAP7_75t_L g379 ( 
.A1(n_337),
.A2(n_358),
.B(n_347),
.Y(n_379)
);

OAI21xp5_ASAP7_75t_L g401 ( 
.A1(n_379),
.A2(n_353),
.B(n_344),
.Y(n_401)
);

INVxp67_ASAP7_75t_L g380 ( 
.A(n_339),
.Y(n_380)
);

MAJIxp5_ASAP7_75t_L g393 ( 
.A(n_381),
.B(n_388),
.C(n_356),
.Y(n_393)
);

CKINVDCx20_ASAP7_75t_R g382 ( 
.A(n_360),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_382),
.B(n_383),
.Y(n_402)
);

OR2x2_ASAP7_75t_L g383 ( 
.A(n_355),
.B(n_304),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_SL g384 ( 
.A(n_341),
.B(n_308),
.Y(n_384)
);

XOR2xp5_ASAP7_75t_L g398 ( 
.A(n_384),
.B(n_385),
.Y(n_398)
);

OAI32xp33_ASAP7_75t_L g385 ( 
.A1(n_358),
.A2(n_304),
.A3(n_331),
.B1(n_314),
.B2(n_313),
.Y(n_385)
);

MAJIxp5_ASAP7_75t_L g388 ( 
.A(n_363),
.B(n_331),
.C(n_303),
.Y(n_388)
);

XNOR2x1_ASAP7_75t_L g390 ( 
.A(n_386),
.B(n_337),
.Y(n_390)
);

XNOR2x1_ASAP7_75t_L g417 ( 
.A(n_390),
.B(n_392),
.Y(n_417)
);

OA21x2_ASAP7_75t_SL g392 ( 
.A1(n_383),
.A2(n_355),
.B(n_352),
.Y(n_392)
);

MAJIxp5_ASAP7_75t_L g411 ( 
.A(n_393),
.B(n_395),
.C(n_397),
.Y(n_411)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_394),
.Y(n_415)
);

MAJIxp5_ASAP7_75t_L g395 ( 
.A(n_381),
.B(n_349),
.C(n_346),
.Y(n_395)
);

MAJIxp5_ASAP7_75t_L g397 ( 
.A(n_386),
.B(n_388),
.C(n_349),
.Y(n_397)
);

OAI22xp5_ASAP7_75t_SL g399 ( 
.A1(n_378),
.A2(n_352),
.B1(n_341),
.B2(n_339),
.Y(n_399)
);

OAI22xp5_ASAP7_75t_SL g416 ( 
.A1(n_399),
.A2(n_405),
.B1(n_408),
.B2(n_409),
.Y(n_416)
);

XOR2xp5_ASAP7_75t_L g427 ( 
.A(n_401),
.B(n_402),
.Y(n_427)
);

MAJIxp5_ASAP7_75t_L g404 ( 
.A(n_379),
.B(n_345),
.C(n_353),
.Y(n_404)
);

MAJIxp5_ASAP7_75t_L g419 ( 
.A(n_404),
.B(n_407),
.C(n_383),
.Y(n_419)
);

OAI22xp5_ASAP7_75t_L g405 ( 
.A1(n_366),
.A2(n_351),
.B1(n_348),
.B2(n_344),
.Y(n_405)
);

MAJIxp5_ASAP7_75t_L g407 ( 
.A(n_377),
.B(n_362),
.C(n_354),
.Y(n_407)
);

OAI22xp5_ASAP7_75t_SL g408 ( 
.A1(n_372),
.A2(n_340),
.B1(n_361),
.B2(n_350),
.Y(n_408)
);

OAI22xp5_ASAP7_75t_L g409 ( 
.A1(n_371),
.A2(n_340),
.B1(n_350),
.B2(n_342),
.Y(n_409)
);

NOR2xp33_ASAP7_75t_L g412 ( 
.A(n_410),
.B(n_376),
.Y(n_412)
);

NOR2xp33_ASAP7_75t_SL g433 ( 
.A(n_412),
.B(n_413),
.Y(n_433)
);

NOR2xp33_ASAP7_75t_L g413 ( 
.A(n_410),
.B(n_384),
.Y(n_413)
);

NOR2xp33_ASAP7_75t_L g414 ( 
.A(n_407),
.B(n_367),
.Y(n_414)
);

CKINVDCx20_ASAP7_75t_R g432 ( 
.A(n_414),
.Y(n_432)
);

CKINVDCx20_ASAP7_75t_R g418 ( 
.A(n_403),
.Y(n_418)
);

NOR3xp33_ASAP7_75t_L g440 ( 
.A(n_418),
.B(n_420),
.C(n_424),
.Y(n_440)
);

MAJIxp5_ASAP7_75t_L g435 ( 
.A(n_419),
.B(n_421),
.C(n_423),
.Y(n_435)
);

NOR2xp33_ASAP7_75t_L g420 ( 
.A(n_399),
.B(n_367),
.Y(n_420)
);

MAJIxp5_ASAP7_75t_L g421 ( 
.A(n_397),
.B(n_370),
.C(n_369),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_403),
.Y(n_422)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_422),
.Y(n_429)
);

MAJIxp5_ASAP7_75t_L g423 ( 
.A(n_393),
.B(n_369),
.C(n_373),
.Y(n_423)
);

CKINVDCx20_ASAP7_75t_R g424 ( 
.A(n_402),
.Y(n_424)
);

MAJIxp5_ASAP7_75t_L g425 ( 
.A(n_395),
.B(n_385),
.C(n_387),
.Y(n_425)
);

MAJIxp5_ASAP7_75t_L g436 ( 
.A(n_425),
.B(n_426),
.C(n_404),
.Y(n_436)
);

MAJIxp5_ASAP7_75t_L g426 ( 
.A(n_390),
.B(n_387),
.C(n_389),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_427),
.B(n_401),
.Y(n_430)
);

CKINVDCx20_ASAP7_75t_R g428 ( 
.A(n_427),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_428),
.B(n_438),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_430),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_416),
.B(n_406),
.Y(n_431)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_431),
.Y(n_446)
);

OAI21xp33_ASAP7_75t_L g434 ( 
.A1(n_417),
.A2(n_396),
.B(n_391),
.Y(n_434)
);

XOR2xp5_ASAP7_75t_L g445 ( 
.A(n_434),
.B(n_436),
.Y(n_445)
);

NOR3xp33_ASAP7_75t_SL g437 ( 
.A(n_415),
.B(n_392),
.C(n_396),
.Y(n_437)
);

NOR2xp33_ASAP7_75t_SL g443 ( 
.A(n_437),
.B(n_408),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g438 ( 
.A(n_416),
.B(n_406),
.Y(n_438)
);

AOI21xp5_ASAP7_75t_L g439 ( 
.A1(n_415),
.A2(n_398),
.B(n_400),
.Y(n_439)
);

NOR2xp33_ASAP7_75t_L g441 ( 
.A(n_439),
.B(n_398),
.Y(n_441)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_441),
.Y(n_457)
);

NOR2xp33_ASAP7_75t_L g442 ( 
.A(n_432),
.B(n_419),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_L g455 ( 
.A(n_442),
.B(n_444),
.Y(n_455)
);

OR2x2_ASAP7_75t_L g451 ( 
.A(n_443),
.B(n_447),
.Y(n_451)
);

AOI22xp5_ASAP7_75t_L g444 ( 
.A1(n_431),
.A2(n_391),
.B1(n_421),
.B2(n_400),
.Y(n_444)
);

OAI22xp5_ASAP7_75t_SL g447 ( 
.A1(n_439),
.A2(n_423),
.B1(n_425),
.B2(n_426),
.Y(n_447)
);

MAJIxp5_ASAP7_75t_L g448 ( 
.A(n_435),
.B(n_411),
.C(n_390),
.Y(n_448)
);

XOR2xp5_ASAP7_75t_L g454 ( 
.A(n_448),
.B(n_411),
.Y(n_454)
);

OAI21xp5_ASAP7_75t_L g452 ( 
.A1(n_448),
.A2(n_436),
.B(n_435),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_L g466 ( 
.A(n_452),
.B(n_453),
.Y(n_466)
);

AOI22xp33_ASAP7_75t_SL g453 ( 
.A1(n_446),
.A2(n_429),
.B1(n_438),
.B2(n_433),
.Y(n_453)
);

NOR2xp67_ASAP7_75t_SL g465 ( 
.A(n_454),
.B(n_389),
.Y(n_465)
);

AOI22xp33_ASAP7_75t_SL g456 ( 
.A1(n_449),
.A2(n_429),
.B1(n_440),
.B2(n_382),
.Y(n_456)
);

NOR2xp33_ASAP7_75t_L g464 ( 
.A(n_456),
.B(n_445),
.Y(n_464)
);

NOR2xp33_ASAP7_75t_L g458 ( 
.A(n_444),
.B(n_428),
.Y(n_458)
);

NOR2xp33_ASAP7_75t_SL g461 ( 
.A(n_458),
.B(n_450),
.Y(n_461)
);

XOR2xp5_ASAP7_75t_L g459 ( 
.A(n_447),
.B(n_417),
.Y(n_459)
);

XNOR2xp5_ASAP7_75t_L g460 ( 
.A(n_459),
.B(n_445),
.Y(n_460)
);

INVxp67_ASAP7_75t_L g467 ( 
.A(n_460),
.Y(n_467)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_461),
.Y(n_470)
);

OAI21xp5_ASAP7_75t_SL g462 ( 
.A1(n_451),
.A2(n_449),
.B(n_450),
.Y(n_462)
);

AOI21xp33_ASAP7_75t_L g469 ( 
.A1(n_462),
.A2(n_464),
.B(n_465),
.Y(n_469)
);

OAI21xp33_ASAP7_75t_L g463 ( 
.A1(n_457),
.A2(n_430),
.B(n_437),
.Y(n_463)
);

AOI22xp5_ASAP7_75t_L g468 ( 
.A1(n_463),
.A2(n_459),
.B1(n_455),
.B2(n_456),
.Y(n_468)
);

INVxp67_ASAP7_75t_L g473 ( 
.A(n_468),
.Y(n_473)
);

NOR3xp33_ASAP7_75t_SL g471 ( 
.A(n_466),
.B(n_451),
.C(n_453),
.Y(n_471)
);

AOI21xp5_ASAP7_75t_SL g474 ( 
.A1(n_471),
.A2(n_368),
.B(n_405),
.Y(n_474)
);

MAJx2_ASAP7_75t_L g472 ( 
.A(n_470),
.B(n_463),
.C(n_409),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_472),
.B(n_342),
.Y(n_476)
);

OAI311xp33_ASAP7_75t_L g475 ( 
.A1(n_474),
.A2(n_469),
.A3(n_467),
.B1(n_368),
.C1(n_374),
.Y(n_475)
);

AOI21xp5_ASAP7_75t_L g477 ( 
.A1(n_475),
.A2(n_476),
.B(n_473),
.Y(n_477)
);

OAI21xp5_ASAP7_75t_L g478 ( 
.A1(n_477),
.A2(n_342),
.B(n_343),
.Y(n_478)
);

XOR2xp5_ASAP7_75t_L g479 ( 
.A(n_478),
.B(n_343),
.Y(n_479)
);

OAI21xp5_ASAP7_75t_SL g480 ( 
.A1(n_479),
.A2(n_343),
.B(n_316),
.Y(n_480)
);


endmodule