module real_jpeg_31401_n_8 (n_5, n_4, n_0, n_1, n_2, n_6, n_7, n_3, n_8);

input n_5;
input n_4;
input n_0;
input n_1;
input n_2;
input n_6;
input n_7;
input n_3;

output n_8;

wire n_17;
wire n_43;
wire n_54;
wire n_37;
wire n_21;
wire n_35;
wire n_38;
wire n_50;
wire n_33;
wire n_29;
wire n_49;
wire n_10;
wire n_31;
wire n_9;
wire n_52;
wire n_12;
wire n_24;
wire n_34;
wire n_44;
wire n_28;
wire n_46;
wire n_23;
wire n_47;
wire n_14;
wire n_11;
wire n_51;
wire n_45;
wire n_25;
wire n_42;
wire n_22;
wire n_18;
wire n_53;
wire n_40;
wire n_36;
wire n_39;
wire n_41;
wire n_27;
wire n_26;
wire n_20;
wire n_19;
wire n_32;
wire n_48;
wire n_30;
wire n_16;
wire n_15;
wire n_13;

AND2x2_ASAP7_75t_L g18 ( 
.A(n_0),
.B(n_1),
.Y(n_18)
);

AND2x2_ASAP7_75t_L g40 ( 
.A(n_0),
.B(n_41),
.Y(n_40)
);

CKINVDCx5p33_ASAP7_75t_R g49 ( 
.A(n_0),
.Y(n_49)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_1),
.Y(n_41)
);

BUFx2_ASAP7_75t_R g13 ( 
.A(n_2),
.Y(n_13)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

NAND2x1p5_ASAP7_75t_L g26 ( 
.A(n_2),
.B(n_27),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_2),
.B(n_35),
.Y(n_34)
);

AOI322xp5_ASAP7_75t_L g42 ( 
.A1(n_3),
.A2(n_43),
.A3(n_44),
.B1(n_45),
.B2(n_47),
.C1(n_50),
.C2(n_54),
.Y(n_42)
);

INVx4_ASAP7_75t_L g11 ( 
.A(n_4),
.Y(n_11)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_4),
.B(n_23),
.Y(n_29)
);

AND2x2_ASAP7_75t_L g30 ( 
.A(n_4),
.B(n_31),
.Y(n_30)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

AND2x2_ASAP7_75t_L g24 ( 
.A(n_7),
.B(n_25),
.Y(n_24)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

OAI221xp5_ASAP7_75t_L g8 ( 
.A1(n_9),
.A2(n_14),
.B1(n_28),
.B2(n_38),
.C(n_42),
.Y(n_8)
);

INVx1_ASAP7_75t_L g9 ( 
.A(n_10),
.Y(n_9)
);

NAND2xp5_ASAP7_75t_SL g10 ( 
.A(n_11),
.B(n_12),
.Y(n_10)
);

OR2x2_ASAP7_75t_L g21 ( 
.A(n_11),
.B(n_22),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_SL g43 ( 
.A(n_11),
.B(n_22),
.Y(n_43)
);

OR2x2_ASAP7_75t_L g44 ( 
.A(n_11),
.B(n_12),
.Y(n_44)
);

OR2x2_ASAP7_75t_L g52 ( 
.A(n_11),
.B(n_23),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_11),
.B(n_31),
.Y(n_53)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_13),
.Y(n_12)
);

INVxp67_ASAP7_75t_L g14 ( 
.A(n_15),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_20),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_17),
.Y(n_16)
);

AND2x2_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_19),
.Y(n_17)
);

AND2x4_ASAP7_75t_L g54 ( 
.A(n_18),
.B(n_46),
.Y(n_54)
);

AND2x2_ASAP7_75t_SL g39 ( 
.A(n_19),
.B(n_40),
.Y(n_39)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_19),
.Y(n_46)
);

CKINVDCx16_ASAP7_75t_R g20 ( 
.A(n_21),
.Y(n_20)
);

OA21x2_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_24),
.B(n_26),
.Y(n_22)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_23),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_25),
.B(n_27),
.Y(n_37)
);

INVx1_ASAP7_75t_SL g35 ( 
.A(n_27),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_30),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_32),
.Y(n_31)
);

OA21x2_ASAP7_75t_L g32 ( 
.A1(n_33),
.A2(n_34),
.B(n_36),
.Y(n_32)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_39),
.Y(n_38)
);

AND2x4_ASAP7_75t_L g45 ( 
.A(n_40),
.B(n_46),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

BUFx12f_ASAP7_75t_SL g48 ( 
.A(n_49),
.Y(n_48)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_52),
.B(n_53),
.Y(n_51)
);


endmodule