module fake_netlist_6_1555_n_1611 (n_52, n_16, n_1, n_91, n_119, n_46, n_18, n_21, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_138, n_22, n_68, n_28, n_50, n_49, n_7, n_83, n_5, n_101, n_127, n_125, n_77, n_106, n_92, n_42, n_133, n_96, n_8, n_90, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_75, n_109, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_1611);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_18;
input n_21;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_138;
input n_22;
input n_68;
input n_28;
input n_50;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_127;
input n_125;
input n_77;
input n_106;
input n_92;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_75;
input n_109;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1611;

wire n_992;
wire n_801;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_168;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_783;
wire n_798;
wire n_188;
wire n_1575;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_805;
wire n_1151;
wire n_396;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1009;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_424;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_200;
wire n_447;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1078;
wire n_250;
wire n_544;
wire n_1140;
wire n_1444;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1572;
wire n_658;
wire n_616;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_494;
wire n_539;
wire n_493;
wire n_155;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_407;
wire n_913;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_163;
wire n_1558;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_577;
wire n_166;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_243;
wire n_979;
wire n_905;
wire n_175;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_692;
wire n_733;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_318;
wire n_1111;
wire n_715;
wire n_1251;
wire n_1265;
wire n_530;
wire n_1563;
wire n_277;
wire n_618;
wire n_1297;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_210;
wire n_1069;
wire n_612;
wire n_178;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_429;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1504;
wire n_286;
wire n_254;
wire n_242;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_816;
wire n_1157;
wire n_1462;
wire n_1188;
wire n_877;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_170;
wire n_891;
wire n_1412;
wire n_949;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_148;
wire n_161;
wire n_462;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_297;
wire n_627;
wire n_595;
wire n_524;
wire n_1465;
wire n_342;
wire n_1044;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_353;
wire n_605;
wire n_1514;
wire n_826;
wire n_872;
wire n_1139;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_173;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_622;
wire n_147;
wire n_1469;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_631;
wire n_720;
wire n_153;
wire n_842;
wire n_1432;
wire n_156;
wire n_145;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1246;
wire n_899;
wire n_189;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1474;
wire n_1571;
wire n_1577;
wire n_1181;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1505;
wire n_803;
wire n_290;
wire n_926;
wire n_927;
wire n_919;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_154;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1507;
wire n_184;
wire n_552;
wire n_1358;
wire n_1388;
wire n_216;
wire n_912;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1395;
wire n_731;
wire n_1502;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_527;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_150;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_211;
wire n_1483;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_319;
wire n_1339;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1220;
wire n_556;
wire n_162;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_146;
wire n_1252;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1053;
wire n_416;
wire n_520;
wire n_418;
wire n_1093;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_914;
wire n_759;
wire n_426;
wire n_317;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1224;
wire n_1459;
wire n_1135;
wire n_1179;
wire n_1169;
wire n_401;
wire n_324;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1580;
wire n_1425;
wire n_1267;
wire n_1281;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1419;
wire n_351;
wire n_259;
wire n_177;
wire n_1437;
wire n_385;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1594;
wire n_664;
wire n_171;
wire n_169;
wire n_1429;
wire n_1610;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1079;
wire n_341;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_144;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_160;
wire n_186;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1024;
wire n_198;
wire n_179;
wire n_248;
wire n_517;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_183;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1182;
wire n_1298;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_167;
wire n_1356;
wire n_1589;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1586;
wire n_302;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_397;
wire n_1262;
wire n_218;
wire n_1213;
wire n_1350;
wire n_172;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_352;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1361;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_450;
wire n_921;
wire n_1346;
wire n_711;
wire n_579;
wire n_1352;
wire n_937;
wire n_370;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_152;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_227;
wire n_204;
wire n_482;
wire n_934;
wire n_1407;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1489;
wire n_164;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_282;
wire n_833;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_159;
wire n_1086;
wire n_1066;
wire n_157;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1484;
wire n_1321;
wire n_1241;
wire n_569;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_786;
wire n_1236;
wire n_1559;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1325;
wire n_1002;
wire n_545;
wire n_489;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_151;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_187;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1562;
wire n_398;
wire n_1191;
wire n_566;
wire n_1023;
wire n_1118;
wire n_1076;
wire n_194;
wire n_1007;
wire n_1378;
wire n_855;
wire n_1592;
wire n_591;
wire n_1377;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_661;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_310;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_180;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_181;
wire n_182;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_555;
wire n_389;
wire n_814;
wire n_669;
wire n_176;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_763;
wire n_1147;
wire n_360;
wire n_1506;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_174;
wire n_1173;
wire n_525;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1219;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1109;
wire n_185;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1525;
wire n_455;
wire n_1585;
wire n_363;
wire n_1090;
wire n_592;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_503;
wire n_1450;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1574;
wire n_240;
wire n_756;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1479;
wire n_1055;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_404;
wire n_271;
wire n_158;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1010;
wire n_149;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_534;
wire n_1578;
wire n_1006;
wire n_373;
wire n_257;
wire n_1557;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_207;
wire n_1089;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_1576;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_165;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_1259;
wire n_192;
wire n_1538;
wire n_649;
wire n_1240;

INVx1_ASAP7_75t_L g144 ( 
.A(n_85),
.Y(n_144)
);

BUFx3_ASAP7_75t_L g145 ( 
.A(n_116),
.Y(n_145)
);

INVx1_ASAP7_75t_SL g146 ( 
.A(n_108),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_83),
.Y(n_147)
);

CKINVDCx5p33_ASAP7_75t_R g148 ( 
.A(n_31),
.Y(n_148)
);

INVx2_ASAP7_75t_SL g149 ( 
.A(n_0),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_47),
.Y(n_150)
);

INVx2_ASAP7_75t_SL g151 ( 
.A(n_101),
.Y(n_151)
);

CKINVDCx5p33_ASAP7_75t_R g152 ( 
.A(n_93),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_132),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g154 ( 
.A(n_9),
.Y(n_154)
);

BUFx10_ASAP7_75t_L g155 ( 
.A(n_82),
.Y(n_155)
);

CKINVDCx5p33_ASAP7_75t_R g156 ( 
.A(n_121),
.Y(n_156)
);

CKINVDCx5p33_ASAP7_75t_R g157 ( 
.A(n_65),
.Y(n_157)
);

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_26),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_12),
.Y(n_159)
);

CKINVDCx5p33_ASAP7_75t_R g160 ( 
.A(n_7),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_3),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_127),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_3),
.Y(n_163)
);

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_77),
.Y(n_164)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_6),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_115),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_53),
.Y(n_167)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_7),
.Y(n_168)
);

BUFx10_ASAP7_75t_L g169 ( 
.A(n_4),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g170 ( 
.A(n_56),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_84),
.Y(n_171)
);

BUFx6f_ASAP7_75t_L g172 ( 
.A(n_28),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_73),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_91),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_78),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_124),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_29),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_55),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_11),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_129),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_97),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_137),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_14),
.Y(n_183)
);

BUFx3_ASAP7_75t_L g184 ( 
.A(n_5),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_9),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_27),
.Y(n_186)
);

CKINVDCx16_ASAP7_75t_R g187 ( 
.A(n_45),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_45),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_27),
.Y(n_189)
);

INVx1_ASAP7_75t_SL g190 ( 
.A(n_48),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_46),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_46),
.Y(n_192)
);

BUFx6f_ASAP7_75t_L g193 ( 
.A(n_98),
.Y(n_193)
);

BUFx3_ASAP7_75t_L g194 ( 
.A(n_89),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_35),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_2),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_64),
.Y(n_197)
);

INVx1_ASAP7_75t_SL g198 ( 
.A(n_2),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_41),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_18),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_118),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_36),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_30),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_102),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_16),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_94),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_16),
.Y(n_207)
);

BUFx8_ASAP7_75t_SL g208 ( 
.A(n_15),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_25),
.Y(n_209)
);

INVx1_ASAP7_75t_SL g210 ( 
.A(n_122),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_23),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_69),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_18),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_59),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_139),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_104),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_51),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_5),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_95),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_33),
.Y(n_220)
);

BUFx6f_ASAP7_75t_L g221 ( 
.A(n_6),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_112),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_128),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_103),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_96),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_48),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_61),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_29),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_142),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_22),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_87),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_36),
.Y(n_232)
);

INVxp67_ASAP7_75t_L g233 ( 
.A(n_28),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_111),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_39),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_90),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_26),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_50),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_100),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_133),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_32),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_109),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_123),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_106),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_113),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_11),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_41),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_58),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_42),
.Y(n_249)
);

CKINVDCx11_ASAP7_75t_R g250 ( 
.A(n_130),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_79),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_17),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_117),
.Y(n_253)
);

BUFx6f_ASAP7_75t_L g254 ( 
.A(n_136),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_4),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_99),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_126),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_134),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_19),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_107),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_31),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_60),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_57),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_66),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_43),
.Y(n_265)
);

BUFx5_ASAP7_75t_L g266 ( 
.A(n_37),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_15),
.Y(n_267)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_72),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_71),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_70),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_141),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_47),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_30),
.Y(n_273)
);

BUFx6f_ASAP7_75t_L g274 ( 
.A(n_62),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_33),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_14),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_143),
.Y(n_277)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_67),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_63),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_42),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_8),
.Y(n_281)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_140),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_173),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_208),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_266),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_173),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_227),
.Y(n_287)
);

INVxp67_ASAP7_75t_SL g288 ( 
.A(n_145),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g289 ( 
.A(n_227),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_266),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_262),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_250),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_266),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_262),
.Y(n_294)
);

BUFx3_ASAP7_75t_L g295 ( 
.A(n_145),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_266),
.Y(n_296)
);

BUFx3_ASAP7_75t_L g297 ( 
.A(n_194),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_266),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_266),
.Y(n_299)
);

HB1xp67_ASAP7_75t_L g300 ( 
.A(n_187),
.Y(n_300)
);

INVxp67_ASAP7_75t_SL g301 ( 
.A(n_194),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_175),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g303 ( 
.A(n_176),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_266),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_154),
.Y(n_305)
);

INVx1_ASAP7_75t_SL g306 ( 
.A(n_169),
.Y(n_306)
);

INVxp67_ASAP7_75t_L g307 ( 
.A(n_169),
.Y(n_307)
);

INVx2_ASAP7_75t_L g308 ( 
.A(n_154),
.Y(n_308)
);

INVxp67_ASAP7_75t_SL g309 ( 
.A(n_154),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_178),
.Y(n_310)
);

BUFx6f_ASAP7_75t_L g311 ( 
.A(n_170),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_182),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_151),
.B(n_1),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_154),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_172),
.Y(n_315)
);

CKINVDCx16_ASAP7_75t_R g316 ( 
.A(n_169),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_172),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_172),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_151),
.B(n_1),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_201),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_172),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_204),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_206),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_212),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_221),
.Y(n_325)
);

OR2x2_ASAP7_75t_L g326 ( 
.A(n_150),
.B(n_8),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_221),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_221),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_215),
.Y(n_329)
);

CKINVDCx20_ASAP7_75t_R g330 ( 
.A(n_217),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_222),
.Y(n_331)
);

AND2x2_ASAP7_75t_L g332 ( 
.A(n_184),
.B(n_10),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_223),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_221),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_165),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_165),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_225),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_168),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_168),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_229),
.Y(n_340)
);

HB1xp67_ASAP7_75t_L g341 ( 
.A(n_158),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_231),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_184),
.Y(n_343)
);

BUFx3_ASAP7_75t_L g344 ( 
.A(n_155),
.Y(n_344)
);

CKINVDCx20_ASAP7_75t_R g345 ( 
.A(n_234),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_236),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_159),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_238),
.Y(n_348)
);

INVxp33_ASAP7_75t_L g349 ( 
.A(n_183),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_188),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_305),
.Y(n_351)
);

INVx3_ASAP7_75t_L g352 ( 
.A(n_311),
.Y(n_352)
);

INVx3_ASAP7_75t_L g353 ( 
.A(n_311),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_309),
.B(n_152),
.Y(n_354)
);

AND2x2_ASAP7_75t_L g355 ( 
.A(n_332),
.B(n_268),
.Y(n_355)
);

INVx2_ASAP7_75t_L g356 ( 
.A(n_304),
.Y(n_356)
);

INVx2_ASAP7_75t_L g357 ( 
.A(n_285),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_308),
.B(n_152),
.Y(n_358)
);

HB1xp67_ASAP7_75t_L g359 ( 
.A(n_300),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_305),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_314),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_314),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_315),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_315),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_308),
.B(n_156),
.Y(n_365)
);

BUFx2_ASAP7_75t_L g366 ( 
.A(n_307),
.Y(n_366)
);

HB1xp67_ASAP7_75t_L g367 ( 
.A(n_341),
.Y(n_367)
);

CKINVDCx20_ASAP7_75t_R g368 ( 
.A(n_283),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_317),
.Y(n_369)
);

BUFx2_ASAP7_75t_L g370 ( 
.A(n_344),
.Y(n_370)
);

INVx1_ASAP7_75t_SL g371 ( 
.A(n_306),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_317),
.Y(n_372)
);

INVx3_ASAP7_75t_L g373 ( 
.A(n_311),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_302),
.Y(n_374)
);

INVxp33_ASAP7_75t_SL g375 ( 
.A(n_292),
.Y(n_375)
);

BUFx3_ASAP7_75t_L g376 ( 
.A(n_295),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_318),
.Y(n_377)
);

CKINVDCx20_ASAP7_75t_R g378 ( 
.A(n_286),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_318),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_310),
.Y(n_380)
);

INVxp67_ASAP7_75t_L g381 ( 
.A(n_295),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_321),
.Y(n_382)
);

INVxp67_ASAP7_75t_L g383 ( 
.A(n_297),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_321),
.Y(n_384)
);

CKINVDCx16_ASAP7_75t_R g385 ( 
.A(n_316),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_312),
.Y(n_386)
);

BUFx6f_ASAP7_75t_L g387 ( 
.A(n_311),
.Y(n_387)
);

CKINVDCx16_ASAP7_75t_R g388 ( 
.A(n_287),
.Y(n_388)
);

INVx2_ASAP7_75t_L g389 ( 
.A(n_285),
.Y(n_389)
);

CKINVDCx20_ASAP7_75t_R g390 ( 
.A(n_289),
.Y(n_390)
);

INVx3_ASAP7_75t_L g391 ( 
.A(n_311),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_320),
.Y(n_392)
);

INVx2_ASAP7_75t_L g393 ( 
.A(n_290),
.Y(n_393)
);

CKINVDCx20_ASAP7_75t_R g394 ( 
.A(n_291),
.Y(n_394)
);

INVx2_ASAP7_75t_L g395 ( 
.A(n_290),
.Y(n_395)
);

INVx2_ASAP7_75t_L g396 ( 
.A(n_293),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_322),
.Y(n_397)
);

INVx2_ASAP7_75t_L g398 ( 
.A(n_293),
.Y(n_398)
);

INVx3_ASAP7_75t_L g399 ( 
.A(n_296),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_325),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_323),
.Y(n_401)
);

INVx2_ASAP7_75t_L g402 ( 
.A(n_296),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_288),
.B(n_156),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_325),
.Y(n_404)
);

BUFx6f_ASAP7_75t_L g405 ( 
.A(n_298),
.Y(n_405)
);

BUFx3_ASAP7_75t_L g406 ( 
.A(n_297),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_327),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_324),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_329),
.Y(n_409)
);

BUFx6f_ASAP7_75t_L g410 ( 
.A(n_298),
.Y(n_410)
);

CKINVDCx20_ASAP7_75t_R g411 ( 
.A(n_294),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_301),
.B(n_327),
.Y(n_412)
);

BUFx3_ASAP7_75t_L g413 ( 
.A(n_328),
.Y(n_413)
);

BUFx8_ASAP7_75t_L g414 ( 
.A(n_332),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_328),
.Y(n_415)
);

AND2x4_ASAP7_75t_L g416 ( 
.A(n_299),
.B(n_268),
.Y(n_416)
);

BUFx2_ASAP7_75t_L g417 ( 
.A(n_344),
.Y(n_417)
);

INVx2_ASAP7_75t_L g418 ( 
.A(n_299),
.Y(n_418)
);

INVx2_ASAP7_75t_L g419 ( 
.A(n_334),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_331),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_413),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_413),
.Y(n_422)
);

NOR2xp33_ASAP7_75t_L g423 ( 
.A(n_403),
.B(n_333),
.Y(n_423)
);

INVx2_ASAP7_75t_L g424 ( 
.A(n_419),
.Y(n_424)
);

NOR2xp33_ASAP7_75t_L g425 ( 
.A(n_403),
.B(n_337),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_SL g426 ( 
.A(n_414),
.B(n_278),
.Y(n_426)
);

BUFx4f_ASAP7_75t_L g427 ( 
.A(n_370),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_355),
.B(n_340),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_356),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_356),
.Y(n_430)
);

BUFx3_ASAP7_75t_L g431 ( 
.A(n_376),
.Y(n_431)
);

INVx4_ASAP7_75t_L g432 ( 
.A(n_405),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_355),
.B(n_342),
.Y(n_433)
);

BUFx6f_ASAP7_75t_L g434 ( 
.A(n_387),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_356),
.Y(n_435)
);

INVx1_ASAP7_75t_SL g436 ( 
.A(n_371),
.Y(n_436)
);

INVx4_ASAP7_75t_L g437 ( 
.A(n_405),
.Y(n_437)
);

INVx4_ASAP7_75t_L g438 ( 
.A(n_405),
.Y(n_438)
);

AND2x2_ASAP7_75t_L g439 ( 
.A(n_371),
.B(n_346),
.Y(n_439)
);

INVxp67_ASAP7_75t_SL g440 ( 
.A(n_412),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_SL g441 ( 
.A(n_414),
.B(n_278),
.Y(n_441)
);

NOR2xp33_ASAP7_75t_L g442 ( 
.A(n_354),
.B(n_348),
.Y(n_442)
);

BUFx2_ASAP7_75t_L g443 ( 
.A(n_381),
.Y(n_443)
);

NAND3xp33_ASAP7_75t_L g444 ( 
.A(n_381),
.B(n_319),
.C(n_313),
.Y(n_444)
);

INVx2_ASAP7_75t_SL g445 ( 
.A(n_370),
.Y(n_445)
);

INVx2_ASAP7_75t_SL g446 ( 
.A(n_417),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_399),
.Y(n_447)
);

OR2x2_ASAP7_75t_L g448 ( 
.A(n_354),
.B(n_343),
.Y(n_448)
);

OAI22xp5_ASAP7_75t_L g449 ( 
.A1(n_383),
.A2(n_303),
.B1(n_345),
.B2(n_330),
.Y(n_449)
);

HB1xp67_ASAP7_75t_L g450 ( 
.A(n_359),
.Y(n_450)
);

INVx5_ASAP7_75t_L g451 ( 
.A(n_387),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_399),
.Y(n_452)
);

INVx3_ASAP7_75t_L g453 ( 
.A(n_387),
.Y(n_453)
);

INVx1_ASAP7_75t_SL g454 ( 
.A(n_368),
.Y(n_454)
);

AND2x2_ASAP7_75t_L g455 ( 
.A(n_417),
.B(n_349),
.Y(n_455)
);

AND2x2_ASAP7_75t_L g456 ( 
.A(n_383),
.B(n_343),
.Y(n_456)
);

BUFx4f_ASAP7_75t_L g457 ( 
.A(n_416),
.Y(n_457)
);

INVx2_ASAP7_75t_L g458 ( 
.A(n_419),
.Y(n_458)
);

AOI22xp33_ASAP7_75t_L g459 ( 
.A1(n_355),
.A2(n_326),
.B1(n_149),
.B2(n_282),
.Y(n_459)
);

BUFx6f_ASAP7_75t_L g460 ( 
.A(n_387),
.Y(n_460)
);

NOR2xp33_ASAP7_75t_L g461 ( 
.A(n_358),
.B(n_334),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_399),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_357),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_357),
.Y(n_464)
);

INVx4_ASAP7_75t_L g465 ( 
.A(n_405),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_357),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_L g467 ( 
.A(n_376),
.B(n_146),
.Y(n_467)
);

NOR2xp33_ASAP7_75t_L g468 ( 
.A(n_358),
.B(n_347),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_SL g469 ( 
.A(n_414),
.B(n_282),
.Y(n_469)
);

BUFx10_ASAP7_75t_L g470 ( 
.A(n_374),
.Y(n_470)
);

BUFx6f_ASAP7_75t_L g471 ( 
.A(n_387),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_SL g472 ( 
.A(n_414),
.B(n_170),
.Y(n_472)
);

BUFx6f_ASAP7_75t_L g473 ( 
.A(n_387),
.Y(n_473)
);

INVx4_ASAP7_75t_SL g474 ( 
.A(n_416),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_SL g475 ( 
.A(n_414),
.B(n_170),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_389),
.Y(n_476)
);

INVx4_ASAP7_75t_L g477 ( 
.A(n_405),
.Y(n_477)
);

INVx2_ASAP7_75t_L g478 ( 
.A(n_352),
.Y(n_478)
);

NOR2xp33_ASAP7_75t_L g479 ( 
.A(n_365),
.B(n_347),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_SL g480 ( 
.A(n_416),
.B(n_170),
.Y(n_480)
);

AND2x6_ASAP7_75t_L g481 ( 
.A(n_416),
.B(n_193),
.Y(n_481)
);

BUFx3_ASAP7_75t_L g482 ( 
.A(n_376),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_389),
.Y(n_483)
);

INVx2_ASAP7_75t_L g484 ( 
.A(n_352),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_389),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_393),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_393),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_SL g488 ( 
.A(n_416),
.B(n_193),
.Y(n_488)
);

BUFx3_ASAP7_75t_L g489 ( 
.A(n_406),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_L g490 ( 
.A(n_406),
.B(n_210),
.Y(n_490)
);

NOR2xp33_ASAP7_75t_L g491 ( 
.A(n_365),
.B(n_406),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_L g492 ( 
.A(n_412),
.B(n_239),
.Y(n_492)
);

NAND2x1p5_ASAP7_75t_L g493 ( 
.A(n_405),
.B(n_144),
.Y(n_493)
);

BUFx10_ASAP7_75t_L g494 ( 
.A(n_380),
.Y(n_494)
);

NAND2x1p5_ASAP7_75t_L g495 ( 
.A(n_405),
.B(n_147),
.Y(n_495)
);

INVx2_ASAP7_75t_L g496 ( 
.A(n_352),
.Y(n_496)
);

AND2x2_ASAP7_75t_SL g497 ( 
.A(n_366),
.B(n_193),
.Y(n_497)
);

INVx4_ASAP7_75t_L g498 ( 
.A(n_410),
.Y(n_498)
);

NOR2xp33_ASAP7_75t_L g499 ( 
.A(n_366),
.B(n_350),
.Y(n_499)
);

AND2x6_ASAP7_75t_L g500 ( 
.A(n_395),
.B(n_193),
.Y(n_500)
);

NOR2xp33_ASAP7_75t_L g501 ( 
.A(n_351),
.B(n_350),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_395),
.Y(n_502)
);

BUFx3_ASAP7_75t_L g503 ( 
.A(n_410),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_L g504 ( 
.A(n_396),
.B(n_242),
.Y(n_504)
);

INVx4_ASAP7_75t_L g505 ( 
.A(n_410),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_SL g506 ( 
.A(n_386),
.B(n_254),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_L g507 ( 
.A(n_396),
.B(n_245),
.Y(n_507)
);

BUFx6f_ASAP7_75t_L g508 ( 
.A(n_410),
.Y(n_508)
);

NOR2x1p5_ASAP7_75t_L g509 ( 
.A(n_392),
.B(n_284),
.Y(n_509)
);

BUFx10_ASAP7_75t_L g510 ( 
.A(n_397),
.Y(n_510)
);

BUFx6f_ASAP7_75t_L g511 ( 
.A(n_410),
.Y(n_511)
);

AND2x6_ASAP7_75t_L g512 ( 
.A(n_398),
.B(n_254),
.Y(n_512)
);

AOI22xp33_ASAP7_75t_L g513 ( 
.A1(n_398),
.A2(n_326),
.B1(n_149),
.B2(n_280),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_L g514 ( 
.A(n_402),
.B(n_248),
.Y(n_514)
);

INVx1_ASAP7_75t_SL g515 ( 
.A(n_368),
.Y(n_515)
);

INVx2_ASAP7_75t_L g516 ( 
.A(n_353),
.Y(n_516)
);

BUFx6f_ASAP7_75t_L g517 ( 
.A(n_410),
.Y(n_517)
);

XNOR2x2_ASAP7_75t_L g518 ( 
.A(n_388),
.B(n_190),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_402),
.Y(n_519)
);

AND2x4_ASAP7_75t_L g520 ( 
.A(n_351),
.B(n_335),
.Y(n_520)
);

CKINVDCx5p33_ASAP7_75t_R g521 ( 
.A(n_401),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_SL g522 ( 
.A(n_408),
.B(n_254),
.Y(n_522)
);

INVx4_ASAP7_75t_L g523 ( 
.A(n_410),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_402),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_418),
.Y(n_525)
);

INVx3_ASAP7_75t_L g526 ( 
.A(n_353),
.Y(n_526)
);

AOI22xp33_ASAP7_75t_L g527 ( 
.A1(n_418),
.A2(n_196),
.B1(n_275),
.B2(n_189),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_418),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_L g529 ( 
.A(n_353),
.B(n_253),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_SL g530 ( 
.A(n_409),
.B(n_254),
.Y(n_530)
);

INVxp33_ASAP7_75t_L g531 ( 
.A(n_359),
.Y(n_531)
);

INVx5_ASAP7_75t_L g532 ( 
.A(n_353),
.Y(n_532)
);

OR2x2_ASAP7_75t_L g533 ( 
.A(n_367),
.B(n_198),
.Y(n_533)
);

OR2x2_ASAP7_75t_L g534 ( 
.A(n_367),
.B(n_335),
.Y(n_534)
);

INVx3_ASAP7_75t_L g535 ( 
.A(n_353),
.Y(n_535)
);

AND2x6_ASAP7_75t_L g536 ( 
.A(n_360),
.B(n_274),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_L g537 ( 
.A(n_373),
.B(n_256),
.Y(n_537)
);

INVx2_ASAP7_75t_L g538 ( 
.A(n_373),
.Y(n_538)
);

CKINVDCx5p33_ASAP7_75t_R g539 ( 
.A(n_420),
.Y(n_539)
);

NOR2xp33_ASAP7_75t_L g540 ( 
.A(n_361),
.B(n_233),
.Y(n_540)
);

HB1xp67_ASAP7_75t_L g541 ( 
.A(n_361),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_SL g542 ( 
.A(n_385),
.B(n_274),
.Y(n_542)
);

INVx2_ASAP7_75t_L g543 ( 
.A(n_373),
.Y(n_543)
);

AND2x2_ASAP7_75t_L g544 ( 
.A(n_385),
.B(n_336),
.Y(n_544)
);

AND2x6_ASAP7_75t_L g545 ( 
.A(n_362),
.B(n_274),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_362),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_363),
.Y(n_547)
);

INVx4_ASAP7_75t_L g548 ( 
.A(n_373),
.Y(n_548)
);

NOR2xp33_ASAP7_75t_L g549 ( 
.A(n_363),
.B(n_157),
.Y(n_549)
);

BUFx10_ASAP7_75t_L g550 ( 
.A(n_375),
.Y(n_550)
);

AND2x2_ASAP7_75t_L g551 ( 
.A(n_364),
.B(n_336),
.Y(n_551)
);

INVx1_ASAP7_75t_SL g552 ( 
.A(n_378),
.Y(n_552)
);

AOI22xp33_ASAP7_75t_L g553 ( 
.A1(n_364),
.A2(n_191),
.B1(n_200),
.B2(n_203),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_L g554 ( 
.A(n_391),
.B(n_257),
.Y(n_554)
);

OR2x2_ASAP7_75t_L g555 ( 
.A(n_388),
.B(n_338),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_SL g556 ( 
.A(n_497),
.B(n_274),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_L g557 ( 
.A(n_440),
.B(n_369),
.Y(n_557)
);

NOR2xp33_ASAP7_75t_L g558 ( 
.A(n_440),
.B(n_428),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_L g559 ( 
.A(n_491),
.B(n_369),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_L g560 ( 
.A(n_491),
.B(n_372),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_SL g561 ( 
.A(n_497),
.B(n_153),
.Y(n_561)
);

INVx2_ASAP7_75t_L g562 ( 
.A(n_424),
.Y(n_562)
);

INVx4_ASAP7_75t_L g563 ( 
.A(n_431),
.Y(n_563)
);

AND2x2_ASAP7_75t_L g564 ( 
.A(n_436),
.B(n_338),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_L g565 ( 
.A(n_442),
.B(n_372),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_L g566 ( 
.A(n_442),
.B(n_377),
.Y(n_566)
);

NOR2xp33_ASAP7_75t_L g567 ( 
.A(n_433),
.B(n_157),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_L g568 ( 
.A(n_423),
.B(n_377),
.Y(n_568)
);

INVx2_ASAP7_75t_L g569 ( 
.A(n_424),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_421),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_422),
.Y(n_571)
);

INVx8_ASAP7_75t_L g572 ( 
.A(n_521),
.Y(n_572)
);

AOI22xp5_ASAP7_75t_L g573 ( 
.A1(n_423),
.A2(n_425),
.B1(n_441),
.B2(n_426),
.Y(n_573)
);

AOI21x1_ASAP7_75t_L g574 ( 
.A1(n_529),
.A2(n_382),
.B(n_379),
.Y(n_574)
);

INVxp67_ASAP7_75t_L g575 ( 
.A(n_455),
.Y(n_575)
);

INVx2_ASAP7_75t_L g576 ( 
.A(n_458),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_L g577 ( 
.A(n_425),
.B(n_379),
.Y(n_577)
);

INVx2_ASAP7_75t_L g578 ( 
.A(n_458),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_L g579 ( 
.A(n_461),
.B(n_382),
.Y(n_579)
);

AND2x6_ASAP7_75t_SL g580 ( 
.A(n_439),
.B(n_207),
.Y(n_580)
);

AOI22xp5_ASAP7_75t_L g581 ( 
.A1(n_426),
.A2(n_264),
.B1(n_269),
.B2(n_270),
.Y(n_581)
);

AND2x6_ASAP7_75t_SL g582 ( 
.A(n_499),
.B(n_211),
.Y(n_582)
);

NOR2xp33_ASAP7_75t_L g583 ( 
.A(n_443),
.B(n_162),
.Y(n_583)
);

NOR2xp33_ASAP7_75t_L g584 ( 
.A(n_499),
.B(n_162),
.Y(n_584)
);

NOR2xp33_ASAP7_75t_L g585 ( 
.A(n_448),
.B(n_164),
.Y(n_585)
);

INVx2_ASAP7_75t_L g586 ( 
.A(n_429),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_L g587 ( 
.A(n_461),
.B(n_384),
.Y(n_587)
);

NOR2xp33_ASAP7_75t_L g588 ( 
.A(n_492),
.B(n_544),
.Y(n_588)
);

NAND3xp33_ASAP7_75t_SL g589 ( 
.A(n_459),
.B(n_533),
.C(n_531),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_L g590 ( 
.A(n_468),
.B(n_384),
.Y(n_590)
);

INVx3_ASAP7_75t_L g591 ( 
.A(n_520),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_541),
.Y(n_592)
);

INVx3_ASAP7_75t_L g593 ( 
.A(n_520),
.Y(n_593)
);

INVx2_ASAP7_75t_L g594 ( 
.A(n_430),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_541),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_551),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_L g597 ( 
.A(n_468),
.B(n_479),
.Y(n_597)
);

BUFx4f_ASAP7_75t_L g598 ( 
.A(n_555),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_546),
.Y(n_599)
);

NAND3xp33_ASAP7_75t_L g600 ( 
.A(n_459),
.B(n_192),
.C(n_213),
.Y(n_600)
);

NOR2xp33_ASAP7_75t_L g601 ( 
.A(n_444),
.B(n_534),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_L g602 ( 
.A(n_479),
.B(n_400),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_L g603 ( 
.A(n_504),
.B(n_404),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_L g604 ( 
.A(n_507),
.B(n_404),
.Y(n_604)
);

INVx2_ASAP7_75t_SL g605 ( 
.A(n_456),
.Y(n_605)
);

BUFx8_ASAP7_75t_L g606 ( 
.A(n_445),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_L g607 ( 
.A(n_514),
.B(n_407),
.Y(n_607)
);

NOR2xp33_ASAP7_75t_L g608 ( 
.A(n_467),
.B(n_164),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_547),
.Y(n_609)
);

BUFx8_ASAP7_75t_L g610 ( 
.A(n_446),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_L g611 ( 
.A(n_447),
.B(n_415),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_452),
.Y(n_612)
);

INVx2_ASAP7_75t_L g613 ( 
.A(n_463),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_SL g614 ( 
.A(n_457),
.B(n_167),
.Y(n_614)
);

AOI22xp33_ASAP7_75t_L g615 ( 
.A1(n_513),
.A2(n_237),
.B1(n_255),
.B2(n_218),
.Y(n_615)
);

AND2x6_ASAP7_75t_SL g616 ( 
.A(n_540),
.B(n_226),
.Y(n_616)
);

HB1xp67_ASAP7_75t_L g617 ( 
.A(n_450),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_L g618 ( 
.A(n_462),
.B(n_391),
.Y(n_618)
);

OAI21xp33_ASAP7_75t_L g619 ( 
.A1(n_540),
.A2(n_246),
.B(n_265),
.Y(n_619)
);

INVx2_ASAP7_75t_L g620 ( 
.A(n_435),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_482),
.Y(n_621)
);

INVx2_ASAP7_75t_L g622 ( 
.A(n_464),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_482),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_489),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_SL g625 ( 
.A(n_474),
.B(n_171),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_L g626 ( 
.A(n_549),
.B(n_419),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_L g627 ( 
.A(n_490),
.B(n_174),
.Y(n_627)
);

NOR2xp33_ASAP7_75t_L g628 ( 
.A(n_542),
.B(n_166),
.Y(n_628)
);

AOI22xp33_ASAP7_75t_L g629 ( 
.A1(n_513),
.A2(n_272),
.B1(n_163),
.B2(n_230),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_489),
.Y(n_630)
);

INVxp67_ASAP7_75t_SL g631 ( 
.A(n_508),
.Y(n_631)
);

INVx2_ASAP7_75t_L g632 ( 
.A(n_466),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_SL g633 ( 
.A(n_474),
.B(n_180),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_SL g634 ( 
.A(n_427),
.B(n_181),
.Y(n_634)
);

NOR2xp33_ASAP7_75t_L g635 ( 
.A(n_542),
.B(n_166),
.Y(n_635)
);

INVx2_ASAP7_75t_L g636 ( 
.A(n_476),
.Y(n_636)
);

AND2x6_ASAP7_75t_SL g637 ( 
.A(n_518),
.B(n_163),
.Y(n_637)
);

HB1xp67_ASAP7_75t_L g638 ( 
.A(n_454),
.Y(n_638)
);

INVx2_ASAP7_75t_L g639 ( 
.A(n_483),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_SL g640 ( 
.A(n_427),
.B(n_197),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_L g641 ( 
.A(n_526),
.B(n_535),
.Y(n_641)
);

INVx2_ASAP7_75t_L g642 ( 
.A(n_485),
.Y(n_642)
);

NOR2xp33_ASAP7_75t_L g643 ( 
.A(n_506),
.B(n_258),
.Y(n_643)
);

BUFx3_ASAP7_75t_L g644 ( 
.A(n_470),
.Y(n_644)
);

A2O1A1Ixp33_ASAP7_75t_L g645 ( 
.A1(n_501),
.A2(n_214),
.B(n_244),
.C(n_243),
.Y(n_645)
);

INVx2_ASAP7_75t_L g646 ( 
.A(n_486),
.Y(n_646)
);

AOI22xp5_ASAP7_75t_L g647 ( 
.A1(n_441),
.A2(n_263),
.B1(n_271),
.B2(n_260),
.Y(n_647)
);

NOR2xp33_ASAP7_75t_L g648 ( 
.A(n_506),
.B(n_522),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_501),
.Y(n_649)
);

INVx2_ASAP7_75t_L g650 ( 
.A(n_487),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_L g651 ( 
.A(n_537),
.B(n_216),
.Y(n_651)
);

AOI21xp5_ASAP7_75t_L g652 ( 
.A1(n_554),
.A2(n_224),
.B(n_219),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_SL g653 ( 
.A(n_469),
.B(n_240),
.Y(n_653)
);

NOR2xp33_ASAP7_75t_L g654 ( 
.A(n_522),
.B(n_258),
.Y(n_654)
);

INVx2_ASAP7_75t_L g655 ( 
.A(n_502),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_L g656 ( 
.A(n_503),
.B(n_251),
.Y(n_656)
);

NOR2xp33_ASAP7_75t_L g657 ( 
.A(n_530),
.B(n_260),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_SL g658 ( 
.A(n_469),
.B(n_277),
.Y(n_658)
);

HB1xp67_ASAP7_75t_L g659 ( 
.A(n_515),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_L g660 ( 
.A(n_503),
.B(n_277),
.Y(n_660)
);

NOR2xp33_ASAP7_75t_L g661 ( 
.A(n_530),
.B(n_279),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_L g662 ( 
.A(n_519),
.B(n_279),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_L g663 ( 
.A(n_524),
.B(n_148),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_L g664 ( 
.A(n_525),
.B(n_177),
.Y(n_664)
);

AOI22xp5_ASAP7_75t_L g665 ( 
.A1(n_472),
.A2(n_186),
.B1(n_230),
.B2(n_241),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_SL g666 ( 
.A(n_472),
.B(n_155),
.Y(n_666)
);

BUFx3_ASAP7_75t_L g667 ( 
.A(n_470),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_L g668 ( 
.A(n_528),
.B(n_548),
.Y(n_668)
);

NOR2xp67_ASAP7_75t_SL g669 ( 
.A(n_475),
.B(n_160),
.Y(n_669)
);

AOI22xp5_ASAP7_75t_L g670 ( 
.A1(n_475),
.A2(n_488),
.B1(n_480),
.B2(n_509),
.Y(n_670)
);

NAND2x1p5_ASAP7_75t_L g671 ( 
.A(n_480),
.B(n_339),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_SL g672 ( 
.A(n_478),
.B(n_155),
.Y(n_672)
);

INVx2_ASAP7_75t_L g673 ( 
.A(n_484),
.Y(n_673)
);

BUFx2_ASAP7_75t_L g674 ( 
.A(n_552),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_SL g675 ( 
.A(n_496),
.B(n_179),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_SL g676 ( 
.A(n_516),
.B(n_538),
.Y(n_676)
);

AND2x6_ASAP7_75t_L g677 ( 
.A(n_508),
.B(n_49),
.Y(n_677)
);

INVx4_ASAP7_75t_L g678 ( 
.A(n_508),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_L g679 ( 
.A(n_453),
.B(n_195),
.Y(n_679)
);

A2O1A1Ixp33_ASAP7_75t_L g680 ( 
.A1(n_527),
.A2(n_160),
.B(n_161),
.C(n_185),
.Y(n_680)
);

AOI22xp5_ASAP7_75t_L g681 ( 
.A1(n_488),
.A2(n_241),
.B1(n_259),
.B2(n_186),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_SL g682 ( 
.A(n_543),
.B(n_199),
.Y(n_682)
);

INVx5_ASAP7_75t_L g683 ( 
.A(n_481),
.Y(n_683)
);

INVx2_ASAP7_75t_SL g684 ( 
.A(n_494),
.Y(n_684)
);

NOR2xp33_ASAP7_75t_L g685 ( 
.A(n_432),
.B(n_202),
.Y(n_685)
);

NOR2xp33_ASAP7_75t_L g686 ( 
.A(n_432),
.B(n_281),
.Y(n_686)
);

NOR2xp33_ASAP7_75t_L g687 ( 
.A(n_437),
.B(n_205),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_L g688 ( 
.A(n_511),
.B(n_517),
.Y(n_688)
);

NOR2xp33_ASAP7_75t_L g689 ( 
.A(n_437),
.B(n_235),
.Y(n_689)
);

O2A1O1Ixp33_ASAP7_75t_L g690 ( 
.A1(n_527),
.A2(n_259),
.B(n_261),
.C(n_394),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_493),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_SL g692 ( 
.A(n_517),
.B(n_249),
.Y(n_692)
);

INVxp67_ASAP7_75t_L g693 ( 
.A(n_550),
.Y(n_693)
);

AOI22xp33_ASAP7_75t_L g694 ( 
.A1(n_553),
.A2(n_261),
.B1(n_185),
.B2(n_161),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_493),
.Y(n_695)
);

AOI21xp5_ASAP7_75t_L g696 ( 
.A1(n_688),
.A2(n_465),
.B(n_498),
.Y(n_696)
);

NOR2xp33_ASAP7_75t_L g697 ( 
.A(n_597),
.B(n_539),
.Y(n_697)
);

BUFx3_ASAP7_75t_L g698 ( 
.A(n_572),
.Y(n_698)
);

OR2x2_ASAP7_75t_L g699 ( 
.A(n_617),
.B(n_553),
.Y(n_699)
);

AOI21xp5_ASAP7_75t_L g700 ( 
.A1(n_668),
.A2(n_465),
.B(n_438),
.Y(n_700)
);

OAI321xp33_ASAP7_75t_L g701 ( 
.A1(n_573),
.A2(n_495),
.A3(n_276),
.B1(n_228),
.B2(n_232),
.C(n_247),
.Y(n_701)
);

INVx1_ASAP7_75t_SL g702 ( 
.A(n_674),
.Y(n_702)
);

AOI21xp5_ASAP7_75t_L g703 ( 
.A1(n_557),
.A2(n_477),
.B(n_438),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_SL g704 ( 
.A(n_558),
.B(n_588),
.Y(n_704)
);

O2A1O1Ixp33_ASAP7_75t_L g705 ( 
.A1(n_558),
.A2(n_495),
.B(n_411),
.C(n_390),
.Y(n_705)
);

OAI21xp5_ASAP7_75t_L g706 ( 
.A1(n_588),
.A2(n_477),
.B(n_505),
.Y(n_706)
);

A2O1A1Ixp33_ASAP7_75t_L g707 ( 
.A1(n_648),
.A2(n_209),
.B(n_273),
.C(n_252),
.Y(n_707)
);

BUFx8_ASAP7_75t_L g708 ( 
.A(n_684),
.Y(n_708)
);

INVx3_ASAP7_75t_L g709 ( 
.A(n_591),
.Y(n_709)
);

OAI22xp5_ASAP7_75t_L g710 ( 
.A1(n_649),
.A2(n_276),
.B1(n_267),
.B2(n_220),
.Y(n_710)
);

INVx2_ASAP7_75t_L g711 ( 
.A(n_569),
.Y(n_711)
);

NOR2xp33_ASAP7_75t_L g712 ( 
.A(n_575),
.B(n_390),
.Y(n_712)
);

OAI22xp5_ASAP7_75t_L g713 ( 
.A1(n_665),
.A2(n_411),
.B1(n_517),
.B2(n_471),
.Y(n_713)
);

OAI21xp5_ASAP7_75t_L g714 ( 
.A1(n_559),
.A2(n_523),
.B(n_505),
.Y(n_714)
);

AOI21xp5_ASAP7_75t_L g715 ( 
.A1(n_641),
.A2(n_498),
.B(n_523),
.Y(n_715)
);

AND2x2_ASAP7_75t_L g716 ( 
.A(n_584),
.B(n_510),
.Y(n_716)
);

INVx2_ASAP7_75t_L g717 ( 
.A(n_569),
.Y(n_717)
);

O2A1O1Ixp33_ASAP7_75t_L g718 ( 
.A1(n_556),
.A2(n_481),
.B(n_13),
.C(n_17),
.Y(n_718)
);

AOI21x1_ASAP7_75t_L g719 ( 
.A1(n_676),
.A2(n_434),
.B(n_460),
.Y(n_719)
);

AO21x1_ASAP7_75t_L g720 ( 
.A1(n_653),
.A2(n_556),
.B(n_658),
.Y(n_720)
);

AND2x2_ASAP7_75t_L g721 ( 
.A(n_584),
.B(n_10),
.Y(n_721)
);

AND2x2_ASAP7_75t_L g722 ( 
.A(n_585),
.B(n_13),
.Y(n_722)
);

OR2x6_ASAP7_75t_L g723 ( 
.A(n_572),
.B(n_434),
.Y(n_723)
);

AOI21xp5_ASAP7_75t_L g724 ( 
.A1(n_603),
.A2(n_434),
.B(n_460),
.Y(n_724)
);

BUFx2_ASAP7_75t_L g725 ( 
.A(n_638),
.Y(n_725)
);

OAI21xp5_ASAP7_75t_L g726 ( 
.A1(n_560),
.A2(n_481),
.B(n_500),
.Y(n_726)
);

INVx4_ASAP7_75t_L g727 ( 
.A(n_563),
.Y(n_727)
);

BUFx3_ASAP7_75t_L g728 ( 
.A(n_572),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_L g729 ( 
.A(n_565),
.B(n_434),
.Y(n_729)
);

AOI21xp5_ASAP7_75t_L g730 ( 
.A1(n_604),
.A2(n_460),
.B(n_471),
.Y(n_730)
);

AOI22xp5_ASAP7_75t_L g731 ( 
.A1(n_601),
.A2(n_481),
.B1(n_460),
.B2(n_471),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_L g732 ( 
.A(n_566),
.B(n_473),
.Y(n_732)
);

A2O1A1Ixp33_ASAP7_75t_L g733 ( 
.A1(n_628),
.A2(n_473),
.B(n_532),
.C(n_451),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_599),
.Y(n_734)
);

AOI21xp5_ASAP7_75t_L g735 ( 
.A1(n_607),
.A2(n_631),
.B(n_678),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_L g736 ( 
.A(n_568),
.B(n_473),
.Y(n_736)
);

CKINVDCx10_ASAP7_75t_R g737 ( 
.A(n_637),
.Y(n_737)
);

AOI21x1_ASAP7_75t_L g738 ( 
.A1(n_676),
.A2(n_532),
.B(n_451),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_L g739 ( 
.A(n_577),
.B(n_532),
.Y(n_739)
);

INVx5_ASAP7_75t_L g740 ( 
.A(n_677),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_609),
.Y(n_741)
);

O2A1O1Ixp5_ASAP7_75t_L g742 ( 
.A1(n_614),
.A2(n_545),
.B(n_536),
.C(n_512),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_612),
.Y(n_743)
);

INVx1_ASAP7_75t_SL g744 ( 
.A(n_659),
.Y(n_744)
);

BUFx6f_ASAP7_75t_L g745 ( 
.A(n_563),
.Y(n_745)
);

OAI21xp5_ASAP7_75t_L g746 ( 
.A1(n_626),
.A2(n_512),
.B(n_500),
.Y(n_746)
);

NOR2xp33_ASAP7_75t_L g747 ( 
.A(n_567),
.B(n_19),
.Y(n_747)
);

AOI21xp5_ASAP7_75t_L g748 ( 
.A1(n_691),
.A2(n_536),
.B(n_545),
.Y(n_748)
);

AOI21xp5_ASAP7_75t_L g749 ( 
.A1(n_695),
.A2(n_536),
.B(n_545),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_L g750 ( 
.A(n_590),
.B(n_545),
.Y(n_750)
);

A2O1A1Ixp33_ASAP7_75t_L g751 ( 
.A1(n_628),
.A2(n_20),
.B(n_21),
.C(n_22),
.Y(n_751)
);

BUFx6f_ASAP7_75t_L g752 ( 
.A(n_677),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_L g753 ( 
.A(n_602),
.B(n_545),
.Y(n_753)
);

OAI21xp33_ASAP7_75t_L g754 ( 
.A1(n_694),
.A2(n_20),
.B(n_21),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_SL g755 ( 
.A(n_593),
.B(n_536),
.Y(n_755)
);

AOI21xp5_ASAP7_75t_L g756 ( 
.A1(n_614),
.A2(n_536),
.B(n_80),
.Y(n_756)
);

A2O1A1Ixp33_ASAP7_75t_L g757 ( 
.A1(n_635),
.A2(n_23),
.B(n_24),
.C(n_25),
.Y(n_757)
);

OAI22xp5_ASAP7_75t_L g758 ( 
.A1(n_629),
.A2(n_24),
.B1(n_34),
.B2(n_37),
.Y(n_758)
);

AOI21xp5_ASAP7_75t_L g759 ( 
.A1(n_679),
.A2(n_86),
.B(n_135),
.Y(n_759)
);

A2O1A1Ixp33_ASAP7_75t_L g760 ( 
.A1(n_635),
.A2(n_34),
.B(n_38),
.C(n_39),
.Y(n_760)
);

A2O1A1Ixp33_ASAP7_75t_L g761 ( 
.A1(n_643),
.A2(n_38),
.B(n_40),
.C(n_44),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_L g762 ( 
.A(n_608),
.B(n_44),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_L g763 ( 
.A(n_608),
.B(n_52),
.Y(n_763)
);

NOR2xp67_ASAP7_75t_L g764 ( 
.A(n_693),
.B(n_54),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_613),
.Y(n_765)
);

INVx2_ASAP7_75t_L g766 ( 
.A(n_632),
.Y(n_766)
);

AOI21x1_ASAP7_75t_L g767 ( 
.A1(n_656),
.A2(n_68),
.B(n_74),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_L g768 ( 
.A(n_585),
.B(n_75),
.Y(n_768)
);

OAI21x1_ASAP7_75t_L g769 ( 
.A1(n_611),
.A2(n_76),
.B(n_81),
.Y(n_769)
);

BUFx6f_ASAP7_75t_L g770 ( 
.A(n_677),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_L g771 ( 
.A(n_567),
.B(n_88),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_L g772 ( 
.A(n_579),
.B(n_92),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_SL g773 ( 
.A(n_605),
.B(n_105),
.Y(n_773)
);

OAI21xp5_ASAP7_75t_L g774 ( 
.A1(n_601),
.A2(n_110),
.B(n_114),
.Y(n_774)
);

OAI22xp5_ASAP7_75t_L g775 ( 
.A1(n_629),
.A2(n_119),
.B1(n_120),
.B2(n_125),
.Y(n_775)
);

A2O1A1Ixp33_ASAP7_75t_L g776 ( 
.A1(n_643),
.A2(n_131),
.B(n_138),
.C(n_654),
.Y(n_776)
);

AND2x2_ASAP7_75t_L g777 ( 
.A(n_583),
.B(n_592),
.Y(n_777)
);

AOI21xp5_ASAP7_75t_L g778 ( 
.A1(n_651),
.A2(n_660),
.B(n_587),
.Y(n_778)
);

BUFx4f_ASAP7_75t_L g779 ( 
.A(n_677),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_L g780 ( 
.A(n_627),
.B(n_596),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_L g781 ( 
.A(n_570),
.B(n_571),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_SL g782 ( 
.A(n_598),
.B(n_654),
.Y(n_782)
);

A2O1A1Ixp33_ASAP7_75t_L g783 ( 
.A1(n_657),
.A2(n_661),
.B(n_670),
.C(n_561),
.Y(n_783)
);

AOI21xp5_ASAP7_75t_L g784 ( 
.A1(n_625),
.A2(n_633),
.B(n_683),
.Y(n_784)
);

HB1xp67_ASAP7_75t_L g785 ( 
.A(n_595),
.Y(n_785)
);

NOR2xp33_ASAP7_75t_L g786 ( 
.A(n_589),
.B(n_583),
.Y(n_786)
);

NOR2xp33_ASAP7_75t_L g787 ( 
.A(n_598),
.B(n_681),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_SL g788 ( 
.A(n_657),
.B(n_661),
.Y(n_788)
);

BUFx6f_ASAP7_75t_L g789 ( 
.A(n_677),
.Y(n_789)
);

AOI22xp5_ASAP7_75t_L g790 ( 
.A1(n_666),
.A2(n_692),
.B1(n_561),
.B2(n_689),
.Y(n_790)
);

AO22x1_ASAP7_75t_L g791 ( 
.A1(n_606),
.A2(n_610),
.B1(n_621),
.B2(n_624),
.Y(n_791)
);

NOR2xp33_ASAP7_75t_L g792 ( 
.A(n_623),
.B(n_630),
.Y(n_792)
);

AOI22xp33_ASAP7_75t_L g793 ( 
.A1(n_669),
.A2(n_620),
.B1(n_594),
.B2(n_586),
.Y(n_793)
);

AO21x1_ASAP7_75t_L g794 ( 
.A1(n_692),
.A2(n_634),
.B(n_640),
.Y(n_794)
);

NOR2xp33_ASAP7_75t_L g795 ( 
.A(n_634),
.B(n_640),
.Y(n_795)
);

BUFx6f_ASAP7_75t_L g796 ( 
.A(n_644),
.Y(n_796)
);

O2A1O1Ixp33_ASAP7_75t_L g797 ( 
.A1(n_680),
.A2(n_645),
.B(n_675),
.C(n_682),
.Y(n_797)
);

OAI21xp5_ASAP7_75t_L g798 ( 
.A1(n_562),
.A2(n_576),
.B(n_578),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_622),
.Y(n_799)
);

INVx3_ASAP7_75t_L g800 ( 
.A(n_673),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_L g801 ( 
.A(n_685),
.B(n_686),
.Y(n_801)
);

AOI21xp5_ASAP7_75t_L g802 ( 
.A1(n_636),
.A2(n_646),
.B(n_650),
.Y(n_802)
);

NOR3xp33_ASAP7_75t_L g803 ( 
.A(n_690),
.B(n_600),
.C(n_672),
.Y(n_803)
);

OAI21xp5_ASAP7_75t_L g804 ( 
.A1(n_652),
.A2(n_680),
.B(n_645),
.Y(n_804)
);

NAND3xp33_ASAP7_75t_L g805 ( 
.A(n_694),
.B(n_615),
.C(n_647),
.Y(n_805)
);

AOI21xp5_ASAP7_75t_L g806 ( 
.A1(n_639),
.A2(n_642),
.B(n_655),
.Y(n_806)
);

AOI21xp5_ASAP7_75t_L g807 ( 
.A1(n_685),
.A2(n_689),
.B(n_687),
.Y(n_807)
);

AOI21xp5_ASAP7_75t_L g808 ( 
.A1(n_686),
.A2(n_687),
.B(n_664),
.Y(n_808)
);

AOI22xp5_ASAP7_75t_L g809 ( 
.A1(n_675),
.A2(n_682),
.B1(n_663),
.B2(n_662),
.Y(n_809)
);

AOI21xp5_ASAP7_75t_L g810 ( 
.A1(n_672),
.A2(n_671),
.B(n_619),
.Y(n_810)
);

AOI21xp5_ASAP7_75t_L g811 ( 
.A1(n_671),
.A2(n_581),
.B(n_615),
.Y(n_811)
);

NAND2x1p5_ASAP7_75t_L g812 ( 
.A(n_644),
.B(n_667),
.Y(n_812)
);

INVx3_ASAP7_75t_L g813 ( 
.A(n_667),
.Y(n_813)
);

NOR3xp33_ASAP7_75t_L g814 ( 
.A(n_580),
.B(n_616),
.C(n_582),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_L g815 ( 
.A(n_606),
.B(n_610),
.Y(n_815)
);

NOR2xp33_ASAP7_75t_L g816 ( 
.A(n_597),
.B(n_436),
.Y(n_816)
);

BUFx4f_ASAP7_75t_L g817 ( 
.A(n_572),
.Y(n_817)
);

AOI22xp33_ASAP7_75t_L g818 ( 
.A1(n_597),
.A2(n_573),
.B1(n_558),
.B2(n_653),
.Y(n_818)
);

INVx2_ASAP7_75t_L g819 ( 
.A(n_569),
.Y(n_819)
);

CKINVDCx5p33_ASAP7_75t_R g820 ( 
.A(n_572),
.Y(n_820)
);

OAI22xp5_ASAP7_75t_L g821 ( 
.A1(n_597),
.A2(n_573),
.B1(n_459),
.B2(n_558),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_L g822 ( 
.A(n_597),
.B(n_558),
.Y(n_822)
);

BUFx2_ASAP7_75t_L g823 ( 
.A(n_674),
.Y(n_823)
);

AOI21xp5_ASAP7_75t_L g824 ( 
.A1(n_688),
.A2(n_457),
.B(n_668),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_L g825 ( 
.A(n_597),
.B(n_558),
.Y(n_825)
);

AOI21xp5_ASAP7_75t_L g826 ( 
.A1(n_688),
.A2(n_457),
.B(n_668),
.Y(n_826)
);

OAI21xp5_ASAP7_75t_L g827 ( 
.A1(n_597),
.A2(n_558),
.B(n_573),
.Y(n_827)
);

AOI21xp5_ASAP7_75t_L g828 ( 
.A1(n_688),
.A2(n_457),
.B(n_668),
.Y(n_828)
);

AOI21x1_ASAP7_75t_L g829 ( 
.A1(n_676),
.A2(n_574),
.B(n_688),
.Y(n_829)
);

BUFx6f_ASAP7_75t_L g830 ( 
.A(n_563),
.Y(n_830)
);

INVx2_ASAP7_75t_L g831 ( 
.A(n_569),
.Y(n_831)
);

AND2x2_ASAP7_75t_L g832 ( 
.A(n_564),
.B(n_436),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_L g833 ( 
.A(n_597),
.B(n_558),
.Y(n_833)
);

INVx2_ASAP7_75t_L g834 ( 
.A(n_569),
.Y(n_834)
);

OAI21xp5_ASAP7_75t_L g835 ( 
.A1(n_597),
.A2(n_558),
.B(n_573),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_L g836 ( 
.A(n_597),
.B(n_558),
.Y(n_836)
);

AOI21x1_ASAP7_75t_L g837 ( 
.A1(n_676),
.A2(n_574),
.B(n_688),
.Y(n_837)
);

NOR2xp33_ASAP7_75t_L g838 ( 
.A(n_597),
.B(n_436),
.Y(n_838)
);

NOR2xp33_ASAP7_75t_L g839 ( 
.A(n_597),
.B(n_436),
.Y(n_839)
);

OAI22xp5_ASAP7_75t_L g840 ( 
.A1(n_597),
.A2(n_573),
.B1(n_459),
.B2(n_558),
.Y(n_840)
);

AOI21xp5_ASAP7_75t_L g841 ( 
.A1(n_688),
.A2(n_457),
.B(n_668),
.Y(n_841)
);

AOI21x1_ASAP7_75t_L g842 ( 
.A1(n_676),
.A2(n_574),
.B(n_688),
.Y(n_842)
);

BUFx2_ASAP7_75t_L g843 ( 
.A(n_674),
.Y(n_843)
);

OAI21x1_ASAP7_75t_L g844 ( 
.A1(n_574),
.A2(n_641),
.B(n_618),
.Y(n_844)
);

AOI21xp5_ASAP7_75t_L g845 ( 
.A1(n_688),
.A2(n_457),
.B(n_668),
.Y(n_845)
);

NOR2xp33_ASAP7_75t_L g846 ( 
.A(n_597),
.B(n_436),
.Y(n_846)
);

OAI21xp5_ASAP7_75t_L g847 ( 
.A1(n_597),
.A2(n_558),
.B(n_573),
.Y(n_847)
);

NOR3xp33_ASAP7_75t_L g848 ( 
.A(n_589),
.B(n_449),
.C(n_388),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_L g849 ( 
.A(n_597),
.B(n_558),
.Y(n_849)
);

INVxp67_ASAP7_75t_SL g850 ( 
.A(n_591),
.Y(n_850)
);

AO21x1_ASAP7_75t_L g851 ( 
.A1(n_573),
.A2(n_597),
.B(n_653),
.Y(n_851)
);

OR2x6_ASAP7_75t_L g852 ( 
.A(n_572),
.B(n_644),
.Y(n_852)
);

BUFx2_ASAP7_75t_L g853 ( 
.A(n_823),
.Y(n_853)
);

O2A1O1Ixp33_ASAP7_75t_L g854 ( 
.A1(n_821),
.A2(n_840),
.B(n_783),
.C(n_825),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_L g855 ( 
.A(n_822),
.B(n_833),
.Y(n_855)
);

AOI21xp5_ASAP7_75t_L g856 ( 
.A1(n_807),
.A2(n_801),
.B(n_827),
.Y(n_856)
);

INVx1_ASAP7_75t_L g857 ( 
.A(n_734),
.Y(n_857)
);

OAI21xp5_ASAP7_75t_L g858 ( 
.A1(n_827),
.A2(n_847),
.B(n_835),
.Y(n_858)
);

HB1xp67_ASAP7_75t_L g859 ( 
.A(n_702),
.Y(n_859)
);

INVx5_ASAP7_75t_L g860 ( 
.A(n_752),
.Y(n_860)
);

BUFx12f_ASAP7_75t_L g861 ( 
.A(n_820),
.Y(n_861)
);

AOI21xp5_ASAP7_75t_L g862 ( 
.A1(n_835),
.A2(n_847),
.B(n_836),
.Y(n_862)
);

OAI21x1_ASAP7_75t_L g863 ( 
.A1(n_738),
.A2(n_842),
.B(n_837),
.Y(n_863)
);

AOI21xp5_ASAP7_75t_L g864 ( 
.A1(n_849),
.A2(n_778),
.B(n_714),
.Y(n_864)
);

OAI21x1_ASAP7_75t_L g865 ( 
.A1(n_844),
.A2(n_696),
.B(n_715),
.Y(n_865)
);

AND2x2_ASAP7_75t_L g866 ( 
.A(n_832),
.B(n_816),
.Y(n_866)
);

AOI21xp5_ASAP7_75t_L g867 ( 
.A1(n_714),
.A2(n_704),
.B(n_808),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_741),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_L g869 ( 
.A(n_821),
.B(n_840),
.Y(n_869)
);

NOR2xp33_ASAP7_75t_L g870 ( 
.A(n_697),
.B(n_838),
.Y(n_870)
);

AOI21xp5_ASAP7_75t_L g871 ( 
.A1(n_772),
.A2(n_732),
.B(n_729),
.Y(n_871)
);

NAND3xp33_ASAP7_75t_SL g872 ( 
.A(n_705),
.B(n_747),
.C(n_716),
.Y(n_872)
);

AO31x2_ASAP7_75t_L g873 ( 
.A1(n_851),
.A2(n_794),
.A3(n_720),
.B(n_733),
.Y(n_873)
);

CKINVDCx20_ASAP7_75t_R g874 ( 
.A(n_698),
.Y(n_874)
);

OAI21x1_ASAP7_75t_L g875 ( 
.A1(n_824),
.A2(n_828),
.B(n_826),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_L g876 ( 
.A(n_839),
.B(n_846),
.Y(n_876)
);

OAI21xp5_ASAP7_75t_L g877 ( 
.A1(n_818),
.A2(n_811),
.B(n_788),
.Y(n_877)
);

AOI21xp5_ASAP7_75t_L g878 ( 
.A1(n_736),
.A2(n_706),
.B(n_841),
.Y(n_878)
);

AOI21xp5_ASAP7_75t_L g879 ( 
.A1(n_706),
.A2(n_845),
.B(n_735),
.Y(n_879)
);

AOI21x1_ASAP7_75t_L g880 ( 
.A1(n_771),
.A2(n_768),
.B(n_763),
.Y(n_880)
);

INVx5_ASAP7_75t_L g881 ( 
.A(n_752),
.Y(n_881)
);

NAND3xp33_ASAP7_75t_L g882 ( 
.A(n_805),
.B(n_787),
.C(n_848),
.Y(n_882)
);

INVx2_ASAP7_75t_L g883 ( 
.A(n_711),
.Y(n_883)
);

NAND3x1_ASAP7_75t_L g884 ( 
.A(n_814),
.B(n_815),
.C(n_712),
.Y(n_884)
);

A2O1A1Ixp33_ASAP7_75t_L g885 ( 
.A1(n_795),
.A2(n_721),
.B(n_722),
.C(n_797),
.Y(n_885)
);

INVx2_ASAP7_75t_L g886 ( 
.A(n_717),
.Y(n_886)
);

AND2x2_ASAP7_75t_L g887 ( 
.A(n_777),
.B(n_744),
.Y(n_887)
);

HB1xp67_ASAP7_75t_L g888 ( 
.A(n_702),
.Y(n_888)
);

OAI21xp5_ASAP7_75t_L g889 ( 
.A1(n_790),
.A2(n_750),
.B(n_753),
.Y(n_889)
);

OAI21x1_ASAP7_75t_L g890 ( 
.A1(n_798),
.A2(n_700),
.B(n_724),
.Y(n_890)
);

AND2x2_ASAP7_75t_L g891 ( 
.A(n_744),
.B(n_725),
.Y(n_891)
);

OAI21x1_ASAP7_75t_L g892 ( 
.A1(n_798),
.A2(n_730),
.B(n_703),
.Y(n_892)
);

BUFx6f_ASAP7_75t_L g893 ( 
.A(n_745),
.Y(n_893)
);

AOI21xp5_ASAP7_75t_L g894 ( 
.A1(n_739),
.A2(n_810),
.B(n_780),
.Y(n_894)
);

AND2x2_ASAP7_75t_L g895 ( 
.A(n_843),
.B(n_785),
.Y(n_895)
);

NOR2x1_ASAP7_75t_L g896 ( 
.A(n_728),
.B(n_852),
.Y(n_896)
);

INVx1_ASAP7_75t_L g897 ( 
.A(n_765),
.Y(n_897)
);

OAI21xp5_ASAP7_75t_L g898 ( 
.A1(n_809),
.A2(n_726),
.B(n_804),
.Y(n_898)
);

NOR2xp33_ASAP7_75t_L g899 ( 
.A(n_782),
.B(n_699),
.Y(n_899)
);

INVx2_ASAP7_75t_L g900 ( 
.A(n_819),
.Y(n_900)
);

AOI21xp5_ASAP7_75t_L g901 ( 
.A1(n_779),
.A2(n_726),
.B(n_802),
.Y(n_901)
);

O2A1O1Ixp5_ASAP7_75t_L g902 ( 
.A1(n_762),
.A2(n_804),
.B(n_774),
.C(n_746),
.Y(n_902)
);

BUFx6f_ASAP7_75t_L g903 ( 
.A(n_745),
.Y(n_903)
);

A2O1A1Ixp33_ASAP7_75t_L g904 ( 
.A1(n_803),
.A2(n_707),
.B(n_701),
.C(n_792),
.Y(n_904)
);

AOI21xp5_ASAP7_75t_L g905 ( 
.A1(n_779),
.A2(n_806),
.B(n_781),
.Y(n_905)
);

NOR2xp33_ASAP7_75t_SL g906 ( 
.A(n_817),
.B(n_852),
.Y(n_906)
);

BUFx3_ASAP7_75t_L g907 ( 
.A(n_796),
.Y(n_907)
);

INVx2_ASAP7_75t_L g908 ( 
.A(n_831),
.Y(n_908)
);

NAND2x1p5_ASAP7_75t_L g909 ( 
.A(n_740),
.B(n_752),
.Y(n_909)
);

AO31x2_ASAP7_75t_L g910 ( 
.A1(n_776),
.A2(n_757),
.A3(n_751),
.B(n_760),
.Y(n_910)
);

AOI21xp5_ASAP7_75t_L g911 ( 
.A1(n_850),
.A2(n_784),
.B(n_740),
.Y(n_911)
);

AND2x2_ASAP7_75t_L g912 ( 
.A(n_813),
.B(n_796),
.Y(n_912)
);

OAI22xp5_ASAP7_75t_L g913 ( 
.A1(n_740),
.A2(n_709),
.B1(n_731),
.B2(n_830),
.Y(n_913)
);

NAND2x1p5_ASAP7_75t_L g914 ( 
.A(n_740),
.B(n_789),
.Y(n_914)
);

BUFx6f_ASAP7_75t_L g915 ( 
.A(n_745),
.Y(n_915)
);

AOI21xp5_ASAP7_75t_L g916 ( 
.A1(n_793),
.A2(n_766),
.B(n_799),
.Y(n_916)
);

AOI21xp5_ASAP7_75t_L g917 ( 
.A1(n_773),
.A2(n_834),
.B(n_709),
.Y(n_917)
);

O2A1O1Ixp5_ASAP7_75t_L g918 ( 
.A1(n_755),
.A2(n_742),
.B(n_767),
.C(n_775),
.Y(n_918)
);

OAI21x1_ASAP7_75t_L g919 ( 
.A1(n_769),
.A2(n_749),
.B(n_748),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_L g920 ( 
.A(n_743),
.B(n_800),
.Y(n_920)
);

AOI21xp5_ASAP7_75t_L g921 ( 
.A1(n_759),
.A2(n_775),
.B(n_756),
.Y(n_921)
);

NAND2x1p5_ASAP7_75t_L g922 ( 
.A(n_770),
.B(n_789),
.Y(n_922)
);

NAND2xp5_ASAP7_75t_SL g923 ( 
.A(n_830),
.B(n_713),
.Y(n_923)
);

OAI21xp5_ASAP7_75t_L g924 ( 
.A1(n_701),
.A2(n_718),
.B(n_713),
.Y(n_924)
);

AOI21xp5_ASAP7_75t_L g925 ( 
.A1(n_800),
.A2(n_770),
.B(n_789),
.Y(n_925)
);

AOI21x1_ASAP7_75t_L g926 ( 
.A1(n_764),
.A2(n_723),
.B(n_758),
.Y(n_926)
);

A2O1A1Ixp33_ASAP7_75t_L g927 ( 
.A1(n_758),
.A2(n_761),
.B(n_817),
.C(n_813),
.Y(n_927)
);

AOI21xp5_ASAP7_75t_L g928 ( 
.A1(n_770),
.A2(n_830),
.B(n_723),
.Y(n_928)
);

AOI21x1_ASAP7_75t_L g929 ( 
.A1(n_723),
.A2(n_710),
.B(n_791),
.Y(n_929)
);

OAI21xp5_ASAP7_75t_L g930 ( 
.A1(n_710),
.A2(n_727),
.B(n_812),
.Y(n_930)
);

AOI21xp5_ASAP7_75t_L g931 ( 
.A1(n_727),
.A2(n_852),
.B(n_796),
.Y(n_931)
);

AOI21xp5_ASAP7_75t_L g932 ( 
.A1(n_708),
.A2(n_807),
.B(n_801),
.Y(n_932)
);

OAI22xp5_ASAP7_75t_L g933 ( 
.A1(n_708),
.A2(n_597),
.B1(n_822),
.B2(n_825),
.Y(n_933)
);

AOI21xp5_ASAP7_75t_L g934 ( 
.A1(n_737),
.A2(n_807),
.B(n_801),
.Y(n_934)
);

INVx1_ASAP7_75t_L g935 ( 
.A(n_734),
.Y(n_935)
);

OAI21x1_ASAP7_75t_L g936 ( 
.A1(n_719),
.A2(n_738),
.B(n_829),
.Y(n_936)
);

AND2x2_ASAP7_75t_L g937 ( 
.A(n_832),
.B(n_816),
.Y(n_937)
);

AND2x4_ASAP7_75t_L g938 ( 
.A(n_813),
.B(n_723),
.Y(n_938)
);

OAI21x1_ASAP7_75t_L g939 ( 
.A1(n_719),
.A2(n_738),
.B(n_829),
.Y(n_939)
);

AND2x4_ASAP7_75t_L g940 ( 
.A(n_813),
.B(n_723),
.Y(n_940)
);

AOI22xp33_ASAP7_75t_L g941 ( 
.A1(n_805),
.A2(n_747),
.B1(n_786),
.B2(n_721),
.Y(n_941)
);

AND2x2_ASAP7_75t_L g942 ( 
.A(n_832),
.B(n_816),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_L g943 ( 
.A(n_822),
.B(n_825),
.Y(n_943)
);

AOI21xp5_ASAP7_75t_L g944 ( 
.A1(n_807),
.A2(n_801),
.B(n_827),
.Y(n_944)
);

AO31x2_ASAP7_75t_L g945 ( 
.A1(n_851),
.A2(n_794),
.A3(n_720),
.B(n_783),
.Y(n_945)
);

AND2x2_ASAP7_75t_L g946 ( 
.A(n_832),
.B(n_816),
.Y(n_946)
);

NAND2xp5_ASAP7_75t_L g947 ( 
.A(n_822),
.B(n_825),
.Y(n_947)
);

OAI21x1_ASAP7_75t_L g948 ( 
.A1(n_719),
.A2(n_738),
.B(n_829),
.Y(n_948)
);

AO21x1_ASAP7_75t_L g949 ( 
.A1(n_821),
.A2(n_840),
.B(n_835),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_L g950 ( 
.A(n_822),
.B(n_825),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_L g951 ( 
.A(n_822),
.B(n_825),
.Y(n_951)
);

CKINVDCx5p33_ASAP7_75t_R g952 ( 
.A(n_820),
.Y(n_952)
);

OAI21xp5_ASAP7_75t_L g953 ( 
.A1(n_807),
.A2(n_801),
.B(n_783),
.Y(n_953)
);

OAI21xp5_ASAP7_75t_L g954 ( 
.A1(n_807),
.A2(n_801),
.B(n_783),
.Y(n_954)
);

OAI21xp5_ASAP7_75t_L g955 ( 
.A1(n_807),
.A2(n_801),
.B(n_783),
.Y(n_955)
);

INVx1_ASAP7_75t_L g956 ( 
.A(n_734),
.Y(n_956)
);

NOR2xp33_ASAP7_75t_L g957 ( 
.A(n_697),
.B(n_816),
.Y(n_957)
);

NAND2xp5_ASAP7_75t_L g958 ( 
.A(n_822),
.B(n_825),
.Y(n_958)
);

OAI21x1_ASAP7_75t_L g959 ( 
.A1(n_719),
.A2(n_738),
.B(n_829),
.Y(n_959)
);

AOI21xp5_ASAP7_75t_L g960 ( 
.A1(n_807),
.A2(n_801),
.B(n_827),
.Y(n_960)
);

INVx3_ASAP7_75t_L g961 ( 
.A(n_752),
.Y(n_961)
);

A2O1A1Ixp33_ASAP7_75t_L g962 ( 
.A1(n_827),
.A2(n_847),
.B(n_835),
.C(n_573),
.Y(n_962)
);

AND2x4_ASAP7_75t_L g963 ( 
.A(n_813),
.B(n_723),
.Y(n_963)
);

AOI21xp5_ASAP7_75t_SL g964 ( 
.A1(n_783),
.A2(n_835),
.B(n_827),
.Y(n_964)
);

NOR2x1_ASAP7_75t_SL g965 ( 
.A(n_740),
.B(n_752),
.Y(n_965)
);

OAI22xp5_ASAP7_75t_L g966 ( 
.A1(n_822),
.A2(n_597),
.B1(n_833),
.B2(n_825),
.Y(n_966)
);

INVx1_ASAP7_75t_L g967 ( 
.A(n_734),
.Y(n_967)
);

AND2x2_ASAP7_75t_L g968 ( 
.A(n_832),
.B(n_816),
.Y(n_968)
);

AO21x1_ASAP7_75t_L g969 ( 
.A1(n_821),
.A2(n_840),
.B(n_835),
.Y(n_969)
);

OAI21x1_ASAP7_75t_L g970 ( 
.A1(n_719),
.A2(n_738),
.B(n_829),
.Y(n_970)
);

OAI21x1_ASAP7_75t_L g971 ( 
.A1(n_719),
.A2(n_738),
.B(n_829),
.Y(n_971)
);

AOI21xp5_ASAP7_75t_L g972 ( 
.A1(n_807),
.A2(n_801),
.B(n_827),
.Y(n_972)
);

AOI21xp5_ASAP7_75t_L g973 ( 
.A1(n_807),
.A2(n_801),
.B(n_827),
.Y(n_973)
);

INVx5_ASAP7_75t_L g974 ( 
.A(n_752),
.Y(n_974)
);

NAND2xp5_ASAP7_75t_L g975 ( 
.A(n_822),
.B(n_825),
.Y(n_975)
);

NAND2xp5_ASAP7_75t_L g976 ( 
.A(n_822),
.B(n_825),
.Y(n_976)
);

INVx4_ASAP7_75t_L g977 ( 
.A(n_745),
.Y(n_977)
);

OAI21x1_ASAP7_75t_L g978 ( 
.A1(n_719),
.A2(n_738),
.B(n_829),
.Y(n_978)
);

AND2x2_ASAP7_75t_L g979 ( 
.A(n_832),
.B(n_816),
.Y(n_979)
);

OAI22xp5_ASAP7_75t_L g980 ( 
.A1(n_822),
.A2(n_597),
.B1(n_833),
.B2(n_825),
.Y(n_980)
);

OAI21x1_ASAP7_75t_L g981 ( 
.A1(n_719),
.A2(n_738),
.B(n_829),
.Y(n_981)
);

INVxp67_ASAP7_75t_L g982 ( 
.A(n_832),
.Y(n_982)
);

OAI21x1_ASAP7_75t_L g983 ( 
.A1(n_719),
.A2(n_738),
.B(n_829),
.Y(n_983)
);

A2O1A1Ixp33_ASAP7_75t_L g984 ( 
.A1(n_827),
.A2(n_847),
.B(n_835),
.C(n_573),
.Y(n_984)
);

AO21x1_ASAP7_75t_L g985 ( 
.A1(n_821),
.A2(n_840),
.B(n_835),
.Y(n_985)
);

OAI21x1_ASAP7_75t_L g986 ( 
.A1(n_719),
.A2(n_738),
.B(n_829),
.Y(n_986)
);

AND2x4_ASAP7_75t_L g987 ( 
.A(n_912),
.B(n_896),
.Y(n_987)
);

OR2x6_ASAP7_75t_SL g988 ( 
.A(n_952),
.B(n_933),
.Y(n_988)
);

OAI22xp5_ASAP7_75t_L g989 ( 
.A1(n_855),
.A2(n_951),
.B1(n_958),
.B2(n_950),
.Y(n_989)
);

OAI21xp5_ASAP7_75t_L g990 ( 
.A1(n_962),
.A2(n_984),
.B(n_902),
.Y(n_990)
);

NOR2xp33_ASAP7_75t_R g991 ( 
.A(n_874),
.B(n_872),
.Y(n_991)
);

INVxp67_ASAP7_75t_SL g992 ( 
.A(n_855),
.Y(n_992)
);

AOI221x1_ASAP7_75t_L g993 ( 
.A1(n_964),
.A2(n_955),
.B1(n_954),
.B2(n_953),
.C(n_924),
.Y(n_993)
);

AND2x2_ASAP7_75t_L g994 ( 
.A(n_866),
.B(n_937),
.Y(n_994)
);

AND2x4_ASAP7_75t_L g995 ( 
.A(n_938),
.B(n_940),
.Y(n_995)
);

AND2x2_ASAP7_75t_L g996 ( 
.A(n_942),
.B(n_946),
.Y(n_996)
);

CKINVDCx5p33_ASAP7_75t_R g997 ( 
.A(n_861),
.Y(n_997)
);

NOR2xp33_ASAP7_75t_L g998 ( 
.A(n_870),
.B(n_957),
.Y(n_998)
);

NAND2x1p5_ASAP7_75t_L g999 ( 
.A(n_860),
.B(n_881),
.Y(n_999)
);

CKINVDCx5p33_ASAP7_75t_R g1000 ( 
.A(n_853),
.Y(n_1000)
);

INVx3_ASAP7_75t_L g1001 ( 
.A(n_909),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_L g1002 ( 
.A(n_943),
.B(n_947),
.Y(n_1002)
);

A2O1A1Ixp33_ASAP7_75t_L g1003 ( 
.A1(n_885),
.A2(n_898),
.B(n_941),
.C(n_854),
.Y(n_1003)
);

NOR2xp33_ASAP7_75t_L g1004 ( 
.A(n_876),
.B(n_968),
.Y(n_1004)
);

AND2x4_ASAP7_75t_L g1005 ( 
.A(n_938),
.B(n_940),
.Y(n_1005)
);

OAI22xp5_ASAP7_75t_SL g1006 ( 
.A1(n_876),
.A2(n_982),
.B1(n_882),
.B2(n_899),
.Y(n_1006)
);

AND2x4_ASAP7_75t_L g1007 ( 
.A(n_963),
.B(n_907),
.Y(n_1007)
);

BUFx3_ASAP7_75t_L g1008 ( 
.A(n_891),
.Y(n_1008)
);

HB1xp67_ASAP7_75t_L g1009 ( 
.A(n_859),
.Y(n_1009)
);

NAND2xp5_ASAP7_75t_L g1010 ( 
.A(n_943),
.B(n_947),
.Y(n_1010)
);

OR2x6_ASAP7_75t_L g1011 ( 
.A(n_931),
.B(n_928),
.Y(n_1011)
);

NAND2xp5_ASAP7_75t_L g1012 ( 
.A(n_950),
.B(n_951),
.Y(n_1012)
);

OR2x2_ASAP7_75t_L g1013 ( 
.A(n_979),
.B(n_887),
.Y(n_1013)
);

INVx3_ASAP7_75t_L g1014 ( 
.A(n_909),
.Y(n_1014)
);

AO22x1_ASAP7_75t_SL g1015 ( 
.A1(n_963),
.A2(n_935),
.B1(n_868),
.B2(n_956),
.Y(n_1015)
);

CKINVDCx5p33_ASAP7_75t_R g1016 ( 
.A(n_888),
.Y(n_1016)
);

HB1xp67_ASAP7_75t_L g1017 ( 
.A(n_895),
.Y(n_1017)
);

BUFx12f_ASAP7_75t_L g1018 ( 
.A(n_893),
.Y(n_1018)
);

INVx1_ASAP7_75t_L g1019 ( 
.A(n_967),
.Y(n_1019)
);

NOR2xp33_ASAP7_75t_R g1020 ( 
.A(n_906),
.B(n_929),
.Y(n_1020)
);

BUFx4_ASAP7_75t_R g1021 ( 
.A(n_965),
.Y(n_1021)
);

AND2x4_ASAP7_75t_L g1022 ( 
.A(n_931),
.B(n_977),
.Y(n_1022)
);

BUFx12f_ASAP7_75t_L g1023 ( 
.A(n_893),
.Y(n_1023)
);

O2A1O1Ixp5_ASAP7_75t_L g1024 ( 
.A1(n_880),
.A2(n_921),
.B(n_985),
.C(n_949),
.Y(n_1024)
);

BUFx3_ASAP7_75t_L g1025 ( 
.A(n_893),
.Y(n_1025)
);

INVx4_ASAP7_75t_L g1026 ( 
.A(n_903),
.Y(n_1026)
);

INVx1_ASAP7_75t_L g1027 ( 
.A(n_897),
.Y(n_1027)
);

INVx3_ASAP7_75t_L g1028 ( 
.A(n_914),
.Y(n_1028)
);

NAND2xp5_ASAP7_75t_L g1029 ( 
.A(n_958),
.B(n_975),
.Y(n_1029)
);

INVx1_ASAP7_75t_SL g1030 ( 
.A(n_884),
.Y(n_1030)
);

O2A1O1Ixp33_ASAP7_75t_L g1031 ( 
.A1(n_904),
.A2(n_966),
.B(n_980),
.C(n_975),
.Y(n_1031)
);

INVx3_ASAP7_75t_SL g1032 ( 
.A(n_903),
.Y(n_1032)
);

NAND2xp5_ASAP7_75t_L g1033 ( 
.A(n_976),
.B(n_862),
.Y(n_1033)
);

BUFx2_ASAP7_75t_L g1034 ( 
.A(n_903),
.Y(n_1034)
);

INVx2_ASAP7_75t_L g1035 ( 
.A(n_883),
.Y(n_1035)
);

INVx2_ASAP7_75t_L g1036 ( 
.A(n_886),
.Y(n_1036)
);

BUFx6f_ASAP7_75t_L g1037 ( 
.A(n_915),
.Y(n_1037)
);

NAND2xp33_ASAP7_75t_L g1038 ( 
.A(n_976),
.B(n_915),
.Y(n_1038)
);

INVxp67_ASAP7_75t_L g1039 ( 
.A(n_920),
.Y(n_1039)
);

AOI21xp5_ASAP7_75t_L g1040 ( 
.A1(n_864),
.A2(n_879),
.B(n_856),
.Y(n_1040)
);

O2A1O1Ixp5_ASAP7_75t_L g1041 ( 
.A1(n_921),
.A2(n_969),
.B(n_858),
.C(n_877),
.Y(n_1041)
);

AND2x2_ASAP7_75t_L g1042 ( 
.A(n_934),
.B(n_920),
.Y(n_1042)
);

AND2x2_ASAP7_75t_L g1043 ( 
.A(n_900),
.B(n_908),
.Y(n_1043)
);

BUFx6f_ASAP7_75t_L g1044 ( 
.A(n_915),
.Y(n_1044)
);

AOI21xp5_ASAP7_75t_L g1045 ( 
.A1(n_864),
.A2(n_879),
.B(n_856),
.Y(n_1045)
);

INVx3_ASAP7_75t_L g1046 ( 
.A(n_914),
.Y(n_1046)
);

AOI22xp33_ASAP7_75t_L g1047 ( 
.A1(n_869),
.A2(n_923),
.B1(n_973),
.B2(n_944),
.Y(n_1047)
);

INVx2_ASAP7_75t_SL g1048 ( 
.A(n_961),
.Y(n_1048)
);

AOI21xp5_ASAP7_75t_L g1049 ( 
.A1(n_944),
.A2(n_973),
.B(n_960),
.Y(n_1049)
);

NAND2xp5_ASAP7_75t_L g1050 ( 
.A(n_862),
.B(n_854),
.Y(n_1050)
);

NOR2xp67_ASAP7_75t_SL g1051 ( 
.A(n_860),
.B(n_881),
.Y(n_1051)
);

BUFx12f_ASAP7_75t_L g1052 ( 
.A(n_922),
.Y(n_1052)
);

INVx3_ASAP7_75t_SL g1053 ( 
.A(n_860),
.Y(n_1053)
);

OR2x6_ASAP7_75t_L g1054 ( 
.A(n_928),
.B(n_922),
.Y(n_1054)
);

OR2x6_ASAP7_75t_L g1055 ( 
.A(n_932),
.B(n_925),
.Y(n_1055)
);

BUFx12f_ASAP7_75t_L g1056 ( 
.A(n_860),
.Y(n_1056)
);

INVx2_ASAP7_75t_SL g1057 ( 
.A(n_881),
.Y(n_1057)
);

INVx3_ASAP7_75t_L g1058 ( 
.A(n_881),
.Y(n_1058)
);

OR2x2_ASAP7_75t_L g1059 ( 
.A(n_932),
.B(n_930),
.Y(n_1059)
);

NOR2xp33_ASAP7_75t_SL g1060 ( 
.A(n_974),
.B(n_927),
.Y(n_1060)
);

NAND2x1p5_ASAP7_75t_L g1061 ( 
.A(n_974),
.B(n_925),
.Y(n_1061)
);

AOI21xp5_ASAP7_75t_L g1062 ( 
.A1(n_972),
.A2(n_867),
.B(n_894),
.Y(n_1062)
);

AOI21xp5_ASAP7_75t_L g1063 ( 
.A1(n_867),
.A2(n_894),
.B(n_878),
.Y(n_1063)
);

BUFx6f_ASAP7_75t_L g1064 ( 
.A(n_974),
.Y(n_1064)
);

AND2x2_ASAP7_75t_L g1065 ( 
.A(n_910),
.B(n_974),
.Y(n_1065)
);

AND2x2_ASAP7_75t_L g1066 ( 
.A(n_910),
.B(n_945),
.Y(n_1066)
);

INVx1_ASAP7_75t_SL g1067 ( 
.A(n_916),
.Y(n_1067)
);

AND2x2_ASAP7_75t_L g1068 ( 
.A(n_910),
.B(n_945),
.Y(n_1068)
);

NAND2xp5_ASAP7_75t_L g1069 ( 
.A(n_916),
.B(n_889),
.Y(n_1069)
);

NAND3xp33_ASAP7_75t_L g1070 ( 
.A(n_905),
.B(n_901),
.C(n_878),
.Y(n_1070)
);

OR2x6_ASAP7_75t_L g1071 ( 
.A(n_913),
.B(n_905),
.Y(n_1071)
);

BUFx6f_ASAP7_75t_L g1072 ( 
.A(n_926),
.Y(n_1072)
);

BUFx6f_ASAP7_75t_L g1073 ( 
.A(n_919),
.Y(n_1073)
);

AND2x2_ASAP7_75t_L g1074 ( 
.A(n_873),
.B(n_917),
.Y(n_1074)
);

AOI21xp5_ASAP7_75t_L g1075 ( 
.A1(n_871),
.A2(n_901),
.B(n_875),
.Y(n_1075)
);

O2A1O1Ixp33_ASAP7_75t_L g1076 ( 
.A1(n_871),
.A2(n_918),
.B(n_917),
.C(n_911),
.Y(n_1076)
);

NAND2xp5_ASAP7_75t_L g1077 ( 
.A(n_873),
.B(n_911),
.Y(n_1077)
);

NAND2xp5_ASAP7_75t_L g1078 ( 
.A(n_873),
.B(n_863),
.Y(n_1078)
);

NAND2xp5_ASAP7_75t_L g1079 ( 
.A(n_892),
.B(n_890),
.Y(n_1079)
);

INVxp67_ASAP7_75t_L g1080 ( 
.A(n_936),
.Y(n_1080)
);

NAND2xp5_ASAP7_75t_L g1081 ( 
.A(n_939),
.B(n_970),
.Y(n_1081)
);

NOR2xp33_ASAP7_75t_L g1082 ( 
.A(n_948),
.B(n_986),
.Y(n_1082)
);

INVx1_ASAP7_75t_L g1083 ( 
.A(n_959),
.Y(n_1083)
);

AND2x4_ASAP7_75t_L g1084 ( 
.A(n_971),
.B(n_978),
.Y(n_1084)
);

NAND3xp33_ASAP7_75t_SL g1085 ( 
.A(n_865),
.B(n_981),
.C(n_983),
.Y(n_1085)
);

INVx3_ASAP7_75t_L g1086 ( 
.A(n_909),
.Y(n_1086)
);

OR2x2_ASAP7_75t_L g1087 ( 
.A(n_866),
.B(n_436),
.Y(n_1087)
);

INVx2_ASAP7_75t_L g1088 ( 
.A(n_857),
.Y(n_1088)
);

BUFx3_ASAP7_75t_L g1089 ( 
.A(n_853),
.Y(n_1089)
);

CKINVDCx5p33_ASAP7_75t_R g1090 ( 
.A(n_952),
.Y(n_1090)
);

NAND2xp5_ASAP7_75t_L g1091 ( 
.A(n_855),
.B(n_943),
.Y(n_1091)
);

NAND2xp5_ASAP7_75t_L g1092 ( 
.A(n_855),
.B(n_943),
.Y(n_1092)
);

INVx1_ASAP7_75t_SL g1093 ( 
.A(n_891),
.Y(n_1093)
);

NAND2xp5_ASAP7_75t_L g1094 ( 
.A(n_855),
.B(n_943),
.Y(n_1094)
);

OAI21x1_ASAP7_75t_L g1095 ( 
.A1(n_936),
.A2(n_948),
.B(n_939),
.Y(n_1095)
);

HB1xp67_ASAP7_75t_L g1096 ( 
.A(n_859),
.Y(n_1096)
);

NAND2x1p5_ASAP7_75t_L g1097 ( 
.A(n_860),
.B(n_881),
.Y(n_1097)
);

INVx2_ASAP7_75t_L g1098 ( 
.A(n_857),
.Y(n_1098)
);

OAI21xp5_ASAP7_75t_L g1099 ( 
.A1(n_962),
.A2(n_984),
.B(n_902),
.Y(n_1099)
);

INVx2_ASAP7_75t_L g1100 ( 
.A(n_857),
.Y(n_1100)
);

AND2x2_ASAP7_75t_L g1101 ( 
.A(n_866),
.B(n_937),
.Y(n_1101)
);

INVx3_ASAP7_75t_L g1102 ( 
.A(n_909),
.Y(n_1102)
);

INVx3_ASAP7_75t_L g1103 ( 
.A(n_909),
.Y(n_1103)
);

OA21x2_ASAP7_75t_L g1104 ( 
.A1(n_877),
.A2(n_898),
.B(n_864),
.Y(n_1104)
);

INVx3_ASAP7_75t_L g1105 ( 
.A(n_909),
.Y(n_1105)
);

BUFx3_ASAP7_75t_L g1106 ( 
.A(n_853),
.Y(n_1106)
);

INVx1_ASAP7_75t_L g1107 ( 
.A(n_857),
.Y(n_1107)
);

NAND2xp5_ASAP7_75t_L g1108 ( 
.A(n_855),
.B(n_943),
.Y(n_1108)
);

AND2x2_ASAP7_75t_L g1109 ( 
.A(n_866),
.B(n_937),
.Y(n_1109)
);

INVx2_ASAP7_75t_SL g1110 ( 
.A(n_891),
.Y(n_1110)
);

INVx1_ASAP7_75t_L g1111 ( 
.A(n_857),
.Y(n_1111)
);

INVx2_ASAP7_75t_L g1112 ( 
.A(n_857),
.Y(n_1112)
);

INVx1_ASAP7_75t_L g1113 ( 
.A(n_857),
.Y(n_1113)
);

AOI22xp5_ASAP7_75t_L g1114 ( 
.A1(n_870),
.A2(n_957),
.B1(n_697),
.B2(n_712),
.Y(n_1114)
);

INVx4_ASAP7_75t_L g1115 ( 
.A(n_893),
.Y(n_1115)
);

OAI22xp5_ASAP7_75t_L g1116 ( 
.A1(n_855),
.A2(n_597),
.B1(n_825),
.B2(n_822),
.Y(n_1116)
);

BUFx12f_ASAP7_75t_L g1117 ( 
.A(n_861),
.Y(n_1117)
);

AND2x2_ASAP7_75t_L g1118 ( 
.A(n_866),
.B(n_937),
.Y(n_1118)
);

INVx4_ASAP7_75t_L g1119 ( 
.A(n_1053),
.Y(n_1119)
);

AOI22xp33_ASAP7_75t_L g1120 ( 
.A1(n_998),
.A2(n_1114),
.B1(n_1042),
.B2(n_1006),
.Y(n_1120)
);

CKINVDCx20_ASAP7_75t_R g1121 ( 
.A(n_1090),
.Y(n_1121)
);

INVx1_ASAP7_75t_L g1122 ( 
.A(n_1088),
.Y(n_1122)
);

OAI22xp5_ASAP7_75t_L g1123 ( 
.A1(n_1002),
.A2(n_1092),
.B1(n_1012),
.B2(n_1108),
.Y(n_1123)
);

AND2x2_ASAP7_75t_L g1124 ( 
.A(n_992),
.B(n_1002),
.Y(n_1124)
);

INVx1_ASAP7_75t_L g1125 ( 
.A(n_1098),
.Y(n_1125)
);

BUFx12f_ASAP7_75t_L g1126 ( 
.A(n_997),
.Y(n_1126)
);

BUFx2_ASAP7_75t_L g1127 ( 
.A(n_1065),
.Y(n_1127)
);

INVx1_ASAP7_75t_L g1128 ( 
.A(n_1100),
.Y(n_1128)
);

INVx1_ASAP7_75t_L g1129 ( 
.A(n_1112),
.Y(n_1129)
);

HB1xp67_ASAP7_75t_L g1130 ( 
.A(n_1017),
.Y(n_1130)
);

AOI222xp33_ASAP7_75t_L g1131 ( 
.A1(n_1004),
.A2(n_1118),
.B1(n_1109),
.B2(n_1101),
.C1(n_996),
.C2(n_994),
.Y(n_1131)
);

INVx3_ASAP7_75t_L g1132 ( 
.A(n_1072),
.Y(n_1132)
);

INVx1_ASAP7_75t_L g1133 ( 
.A(n_1019),
.Y(n_1133)
);

BUFx8_ASAP7_75t_SL g1134 ( 
.A(n_1117),
.Y(n_1134)
);

INVx2_ASAP7_75t_SL g1135 ( 
.A(n_1037),
.Y(n_1135)
);

CKINVDCx20_ASAP7_75t_R g1136 ( 
.A(n_1000),
.Y(n_1136)
);

AOI22xp33_ASAP7_75t_SL g1137 ( 
.A1(n_991),
.A2(n_1060),
.B1(n_1030),
.B2(n_1020),
.Y(n_1137)
);

OAI22xp33_ASAP7_75t_L g1138 ( 
.A1(n_1010),
.A2(n_1108),
.B1(n_1091),
.B2(n_1012),
.Y(n_1138)
);

INVx1_ASAP7_75t_L g1139 ( 
.A(n_1066),
.Y(n_1139)
);

AND2x2_ASAP7_75t_L g1140 ( 
.A(n_992),
.B(n_1010),
.Y(n_1140)
);

INVx1_ASAP7_75t_L g1141 ( 
.A(n_1107),
.Y(n_1141)
);

INVx1_ASAP7_75t_L g1142 ( 
.A(n_1111),
.Y(n_1142)
);

INVx3_ASAP7_75t_L g1143 ( 
.A(n_1072),
.Y(n_1143)
);

INVx1_ASAP7_75t_L g1144 ( 
.A(n_1113),
.Y(n_1144)
);

AOI21x1_ASAP7_75t_L g1145 ( 
.A1(n_1075),
.A2(n_1079),
.B(n_1045),
.Y(n_1145)
);

INVx1_ASAP7_75t_L g1146 ( 
.A(n_1027),
.Y(n_1146)
);

AOI22xp33_ASAP7_75t_SL g1147 ( 
.A1(n_1116),
.A2(n_989),
.B1(n_1008),
.B2(n_1029),
.Y(n_1147)
);

INVx1_ASAP7_75t_L g1148 ( 
.A(n_1068),
.Y(n_1148)
);

INVx1_ASAP7_75t_L g1149 ( 
.A(n_1083),
.Y(n_1149)
);

NAND2x1p5_ASAP7_75t_L g1150 ( 
.A(n_1072),
.B(n_1059),
.Y(n_1150)
);

BUFx2_ASAP7_75t_L g1151 ( 
.A(n_1009),
.Y(n_1151)
);

AND2x2_ASAP7_75t_L g1152 ( 
.A(n_1029),
.B(n_1091),
.Y(n_1152)
);

AOI21x1_ASAP7_75t_L g1153 ( 
.A1(n_1079),
.A2(n_1045),
.B(n_1040),
.Y(n_1153)
);

BUFx3_ASAP7_75t_L g1154 ( 
.A(n_1018),
.Y(n_1154)
);

INVx2_ASAP7_75t_L g1155 ( 
.A(n_1067),
.Y(n_1155)
);

OA21x2_ASAP7_75t_L g1156 ( 
.A1(n_993),
.A2(n_1024),
.B(n_1063),
.Y(n_1156)
);

AND2x2_ASAP7_75t_L g1157 ( 
.A(n_1092),
.B(n_1094),
.Y(n_1157)
);

INVxp67_ASAP7_75t_SL g1158 ( 
.A(n_1051),
.Y(n_1158)
);

INVx1_ASAP7_75t_L g1159 ( 
.A(n_1043),
.Y(n_1159)
);

BUFx12f_ASAP7_75t_L g1160 ( 
.A(n_1016),
.Y(n_1160)
);

AOI22xp33_ASAP7_75t_L g1161 ( 
.A1(n_990),
.A2(n_1099),
.B1(n_1013),
.B2(n_1110),
.Y(n_1161)
);

INVx1_ASAP7_75t_L g1162 ( 
.A(n_1035),
.Y(n_1162)
);

OAI21x1_ASAP7_75t_L g1163 ( 
.A1(n_1095),
.A2(n_1063),
.B(n_1062),
.Y(n_1163)
);

INVx1_ASAP7_75t_L g1164 ( 
.A(n_1036),
.Y(n_1164)
);

INVx6_ASAP7_75t_L g1165 ( 
.A(n_1056),
.Y(n_1165)
);

NAND2x1p5_ASAP7_75t_L g1166 ( 
.A(n_1022),
.B(n_1074),
.Y(n_1166)
);

INVx1_ASAP7_75t_SL g1167 ( 
.A(n_1093),
.Y(n_1167)
);

BUFx12f_ASAP7_75t_L g1168 ( 
.A(n_1023),
.Y(n_1168)
);

BUFx3_ASAP7_75t_L g1169 ( 
.A(n_1089),
.Y(n_1169)
);

OAI22xp5_ASAP7_75t_L g1170 ( 
.A1(n_1094),
.A2(n_1087),
.B1(n_1116),
.B2(n_1003),
.Y(n_1170)
);

CKINVDCx5p33_ASAP7_75t_R g1171 ( 
.A(n_1106),
.Y(n_1171)
);

INVx1_ASAP7_75t_L g1172 ( 
.A(n_1078),
.Y(n_1172)
);

OAI22x1_ASAP7_75t_L g1173 ( 
.A1(n_1050),
.A2(n_1033),
.B1(n_1039),
.B2(n_1080),
.Y(n_1173)
);

AOI22xp33_ASAP7_75t_L g1174 ( 
.A1(n_990),
.A2(n_1071),
.B1(n_1050),
.B2(n_1038),
.Y(n_1174)
);

CKINVDCx11_ASAP7_75t_R g1175 ( 
.A(n_988),
.Y(n_1175)
);

NAND2xp5_ASAP7_75t_L g1176 ( 
.A(n_1039),
.B(n_1033),
.Y(n_1176)
);

NAND2x1p5_ASAP7_75t_L g1177 ( 
.A(n_1022),
.B(n_1104),
.Y(n_1177)
);

BUFx12f_ASAP7_75t_L g1178 ( 
.A(n_1007),
.Y(n_1178)
);

OAI22xp5_ASAP7_75t_L g1179 ( 
.A1(n_1031),
.A2(n_1096),
.B1(n_1071),
.B2(n_987),
.Y(n_1179)
);

CKINVDCx11_ASAP7_75t_R g1180 ( 
.A(n_1032),
.Y(n_1180)
);

INVx1_ASAP7_75t_L g1181 ( 
.A(n_1015),
.Y(n_1181)
);

AND2x2_ASAP7_75t_L g1182 ( 
.A(n_1031),
.B(n_1047),
.Y(n_1182)
);

INVx4_ASAP7_75t_L g1183 ( 
.A(n_1064),
.Y(n_1183)
);

BUFx2_ASAP7_75t_L g1184 ( 
.A(n_1011),
.Y(n_1184)
);

INVx2_ASAP7_75t_L g1185 ( 
.A(n_1077),
.Y(n_1185)
);

AND2x2_ASAP7_75t_L g1186 ( 
.A(n_995),
.B(n_1005),
.Y(n_1186)
);

AO21x2_ASAP7_75t_L g1187 ( 
.A1(n_1049),
.A2(n_1085),
.B(n_1070),
.Y(n_1187)
);

OAI22xp33_ASAP7_75t_L g1188 ( 
.A1(n_1011),
.A2(n_1071),
.B1(n_1054),
.B2(n_1069),
.Y(n_1188)
);

INVx1_ASAP7_75t_L g1189 ( 
.A(n_1048),
.Y(n_1189)
);

BUFx2_ASAP7_75t_L g1190 ( 
.A(n_1011),
.Y(n_1190)
);

INVx1_ASAP7_75t_L g1191 ( 
.A(n_1077),
.Y(n_1191)
);

CKINVDCx5p33_ASAP7_75t_R g1192 ( 
.A(n_1032),
.Y(n_1192)
);

AOI22xp5_ASAP7_75t_L g1193 ( 
.A1(n_995),
.A2(n_1005),
.B1(n_1054),
.B2(n_1055),
.Y(n_1193)
);

BUFx2_ASAP7_75t_L g1194 ( 
.A(n_1055),
.Y(n_1194)
);

AOI22xp33_ASAP7_75t_SL g1195 ( 
.A1(n_1054),
.A2(n_1055),
.B1(n_1052),
.B2(n_1061),
.Y(n_1195)
);

INVx1_ASAP7_75t_L g1196 ( 
.A(n_1037),
.Y(n_1196)
);

INVx1_ASAP7_75t_L g1197 ( 
.A(n_1037),
.Y(n_1197)
);

INVx4_ASAP7_75t_SL g1198 ( 
.A(n_1064),
.Y(n_1198)
);

AOI21x1_ASAP7_75t_L g1199 ( 
.A1(n_1081),
.A2(n_1084),
.B(n_1085),
.Y(n_1199)
);

OAI21x1_ASAP7_75t_L g1200 ( 
.A1(n_1076),
.A2(n_1041),
.B(n_1082),
.Y(n_1200)
);

INVx1_ASAP7_75t_L g1201 ( 
.A(n_1080),
.Y(n_1201)
);

OAI22xp5_ASAP7_75t_L g1202 ( 
.A1(n_1061),
.A2(n_1034),
.B1(n_999),
.B2(n_1097),
.Y(n_1202)
);

HB1xp67_ASAP7_75t_L g1203 ( 
.A(n_1025),
.Y(n_1203)
);

INVx1_ASAP7_75t_L g1204 ( 
.A(n_1044),
.Y(n_1204)
);

INVx1_ASAP7_75t_L g1205 ( 
.A(n_1044),
.Y(n_1205)
);

OAI21x1_ASAP7_75t_L g1206 ( 
.A1(n_999),
.A2(n_1097),
.B(n_1058),
.Y(n_1206)
);

BUFx6f_ASAP7_75t_L g1207 ( 
.A(n_1058),
.Y(n_1207)
);

CKINVDCx20_ASAP7_75t_R g1208 ( 
.A(n_1044),
.Y(n_1208)
);

BUFx2_ASAP7_75t_L g1209 ( 
.A(n_1026),
.Y(n_1209)
);

INVx3_ASAP7_75t_L g1210 ( 
.A(n_1001),
.Y(n_1210)
);

BUFx3_ASAP7_75t_L g1211 ( 
.A(n_1115),
.Y(n_1211)
);

OA21x2_ASAP7_75t_L g1212 ( 
.A1(n_1073),
.A2(n_1057),
.B(n_1021),
.Y(n_1212)
);

HB1xp67_ASAP7_75t_L g1213 ( 
.A(n_1115),
.Y(n_1213)
);

AOI22xp33_ASAP7_75t_L g1214 ( 
.A1(n_1014),
.A2(n_1086),
.B1(n_1028),
.B2(n_1046),
.Y(n_1214)
);

NAND2xp5_ASAP7_75t_L g1215 ( 
.A(n_1014),
.B(n_1086),
.Y(n_1215)
);

CKINVDCx6p67_ASAP7_75t_R g1216 ( 
.A(n_1073),
.Y(n_1216)
);

AOI22xp33_ASAP7_75t_L g1217 ( 
.A1(n_1028),
.A2(n_1046),
.B1(n_1102),
.B2(n_1103),
.Y(n_1217)
);

AOI22xp33_ASAP7_75t_L g1218 ( 
.A1(n_1103),
.A2(n_998),
.B1(n_870),
.B2(n_957),
.Y(n_1218)
);

INVx3_ASAP7_75t_L g1219 ( 
.A(n_1105),
.Y(n_1219)
);

AO21x2_ASAP7_75t_L g1220 ( 
.A1(n_1040),
.A2(n_1045),
.B(n_1075),
.Y(n_1220)
);

AOI222xp33_ASAP7_75t_L g1221 ( 
.A1(n_998),
.A2(n_758),
.B1(n_754),
.B2(n_805),
.C1(n_957),
.C2(n_870),
.Y(n_1221)
);

OAI22xp33_ASAP7_75t_SL g1222 ( 
.A1(n_1114),
.A2(n_870),
.B1(n_957),
.B2(n_998),
.Y(n_1222)
);

BUFx2_ASAP7_75t_R g1223 ( 
.A(n_1090),
.Y(n_1223)
);

AOI22xp33_ASAP7_75t_L g1224 ( 
.A1(n_998),
.A2(n_870),
.B1(n_957),
.B2(n_747),
.Y(n_1224)
);

OAI21x1_ASAP7_75t_L g1225 ( 
.A1(n_1145),
.A2(n_1163),
.B(n_1153),
.Y(n_1225)
);

AND2x2_ASAP7_75t_L g1226 ( 
.A(n_1139),
.B(n_1148),
.Y(n_1226)
);

INVx2_ASAP7_75t_L g1227 ( 
.A(n_1149),
.Y(n_1227)
);

AND2x2_ASAP7_75t_L g1228 ( 
.A(n_1185),
.B(n_1191),
.Y(n_1228)
);

INVx3_ASAP7_75t_L g1229 ( 
.A(n_1177),
.Y(n_1229)
);

OR2x2_ASAP7_75t_SL g1230 ( 
.A(n_1212),
.B(n_1181),
.Y(n_1230)
);

INVx1_ASAP7_75t_L g1231 ( 
.A(n_1201),
.Y(n_1231)
);

AND2x2_ASAP7_75t_L g1232 ( 
.A(n_1172),
.B(n_1127),
.Y(n_1232)
);

NAND2xp5_ASAP7_75t_L g1233 ( 
.A(n_1124),
.B(n_1140),
.Y(n_1233)
);

INVx2_ASAP7_75t_SL g1234 ( 
.A(n_1184),
.Y(n_1234)
);

AND2x2_ASAP7_75t_L g1235 ( 
.A(n_1127),
.B(n_1156),
.Y(n_1235)
);

AND2x2_ASAP7_75t_L g1236 ( 
.A(n_1156),
.B(n_1182),
.Y(n_1236)
);

INVx1_ASAP7_75t_L g1237 ( 
.A(n_1173),
.Y(n_1237)
);

AND2x2_ASAP7_75t_L g1238 ( 
.A(n_1156),
.B(n_1182),
.Y(n_1238)
);

AND2x2_ASAP7_75t_L g1239 ( 
.A(n_1177),
.B(n_1200),
.Y(n_1239)
);

NAND2xp5_ASAP7_75t_L g1240 ( 
.A(n_1124),
.B(n_1140),
.Y(n_1240)
);

HB1xp67_ASAP7_75t_L g1241 ( 
.A(n_1150),
.Y(n_1241)
);

BUFx6f_ASAP7_75t_L g1242 ( 
.A(n_1194),
.Y(n_1242)
);

AOI22xp33_ASAP7_75t_L g1243 ( 
.A1(n_1224),
.A2(n_1222),
.B1(n_1221),
.B2(n_1120),
.Y(n_1243)
);

NAND2xp5_ASAP7_75t_L g1244 ( 
.A(n_1152),
.B(n_1157),
.Y(n_1244)
);

BUFx3_ASAP7_75t_L g1245 ( 
.A(n_1212),
.Y(n_1245)
);

AND2x2_ASAP7_75t_L g1246 ( 
.A(n_1166),
.B(n_1194),
.Y(n_1246)
);

AND2x4_ASAP7_75t_L g1247 ( 
.A(n_1184),
.B(n_1190),
.Y(n_1247)
);

OR2x2_ASAP7_75t_L g1248 ( 
.A(n_1220),
.B(n_1187),
.Y(n_1248)
);

OA21x2_ASAP7_75t_L g1249 ( 
.A1(n_1174),
.A2(n_1199),
.B(n_1176),
.Y(n_1249)
);

AND2x2_ASAP7_75t_L g1250 ( 
.A(n_1166),
.B(n_1152),
.Y(n_1250)
);

INVx2_ASAP7_75t_SL g1251 ( 
.A(n_1190),
.Y(n_1251)
);

HB1xp67_ASAP7_75t_L g1252 ( 
.A(n_1155),
.Y(n_1252)
);

BUFx6f_ASAP7_75t_L g1253 ( 
.A(n_1199),
.Y(n_1253)
);

OR2x6_ASAP7_75t_L g1254 ( 
.A(n_1179),
.B(n_1155),
.Y(n_1254)
);

BUFx6f_ASAP7_75t_L g1255 ( 
.A(n_1216),
.Y(n_1255)
);

BUFx3_ASAP7_75t_L g1256 ( 
.A(n_1212),
.Y(n_1256)
);

AND2x2_ASAP7_75t_L g1257 ( 
.A(n_1157),
.B(n_1187),
.Y(n_1257)
);

BUFx3_ASAP7_75t_L g1258 ( 
.A(n_1216),
.Y(n_1258)
);

NAND2xp5_ASAP7_75t_L g1259 ( 
.A(n_1138),
.B(n_1123),
.Y(n_1259)
);

BUFx2_ASAP7_75t_L g1260 ( 
.A(n_1151),
.Y(n_1260)
);

HB1xp67_ASAP7_75t_L g1261 ( 
.A(n_1151),
.Y(n_1261)
);

AND2x4_ASAP7_75t_L g1262 ( 
.A(n_1193),
.B(n_1132),
.Y(n_1262)
);

OA21x2_ASAP7_75t_L g1263 ( 
.A1(n_1161),
.A2(n_1170),
.B(n_1146),
.Y(n_1263)
);

HB1xp67_ASAP7_75t_L g1264 ( 
.A(n_1130),
.Y(n_1264)
);

INVx1_ASAP7_75t_L g1265 ( 
.A(n_1133),
.Y(n_1265)
);

INVx1_ASAP7_75t_L g1266 ( 
.A(n_1141),
.Y(n_1266)
);

AO21x2_ASAP7_75t_L g1267 ( 
.A1(n_1188),
.A2(n_1142),
.B(n_1144),
.Y(n_1267)
);

AND2x2_ASAP7_75t_L g1268 ( 
.A(n_1147),
.B(n_1143),
.Y(n_1268)
);

OAI21x1_ASAP7_75t_L g1269 ( 
.A1(n_1143),
.A2(n_1206),
.B(n_1210),
.Y(n_1269)
);

INVx1_ASAP7_75t_L g1270 ( 
.A(n_1122),
.Y(n_1270)
);

INVx1_ASAP7_75t_L g1271 ( 
.A(n_1125),
.Y(n_1271)
);

AO21x2_ASAP7_75t_L g1272 ( 
.A1(n_1128),
.A2(n_1129),
.B(n_1206),
.Y(n_1272)
);

BUFx3_ASAP7_75t_L g1273 ( 
.A(n_1165),
.Y(n_1273)
);

AND2x2_ASAP7_75t_L g1274 ( 
.A(n_1159),
.B(n_1131),
.Y(n_1274)
);

INVx1_ASAP7_75t_L g1275 ( 
.A(n_1162),
.Y(n_1275)
);

INVx1_ASAP7_75t_L g1276 ( 
.A(n_1164),
.Y(n_1276)
);

AND2x2_ASAP7_75t_L g1277 ( 
.A(n_1250),
.B(n_1195),
.Y(n_1277)
);

INVx2_ASAP7_75t_SL g1278 ( 
.A(n_1261),
.Y(n_1278)
);

OAI33xp33_ASAP7_75t_L g1279 ( 
.A1(n_1259),
.A2(n_1189),
.A3(n_1196),
.B1(n_1197),
.B2(n_1204),
.B3(n_1205),
.Y(n_1279)
);

INVx2_ASAP7_75t_L g1280 ( 
.A(n_1227),
.Y(n_1280)
);

BUFx6f_ASAP7_75t_L g1281 ( 
.A(n_1253),
.Y(n_1281)
);

NAND2xp5_ASAP7_75t_L g1282 ( 
.A(n_1244),
.B(n_1218),
.Y(n_1282)
);

OR2x2_ASAP7_75t_L g1283 ( 
.A(n_1257),
.B(n_1167),
.Y(n_1283)
);

AND2x2_ASAP7_75t_L g1284 ( 
.A(n_1257),
.B(n_1219),
.Y(n_1284)
);

OR2x2_ASAP7_75t_L g1285 ( 
.A(n_1257),
.B(n_1203),
.Y(n_1285)
);

NAND2xp5_ASAP7_75t_L g1286 ( 
.A(n_1244),
.B(n_1137),
.Y(n_1286)
);

AND2x2_ASAP7_75t_L g1287 ( 
.A(n_1236),
.B(n_1219),
.Y(n_1287)
);

HB1xp67_ASAP7_75t_L g1288 ( 
.A(n_1261),
.Y(n_1288)
);

AOI222xp33_ASAP7_75t_L g1289 ( 
.A1(n_1243),
.A2(n_1175),
.B1(n_1186),
.B2(n_1160),
.C1(n_1178),
.C2(n_1180),
.Y(n_1289)
);

INVx1_ASAP7_75t_SL g1290 ( 
.A(n_1260),
.Y(n_1290)
);

INVx5_ASAP7_75t_SL g1291 ( 
.A(n_1254),
.Y(n_1291)
);

AND2x2_ASAP7_75t_L g1292 ( 
.A(n_1236),
.B(n_1219),
.Y(n_1292)
);

AOI22xp33_ASAP7_75t_L g1293 ( 
.A1(n_1243),
.A2(n_1175),
.B1(n_1160),
.B2(n_1186),
.Y(n_1293)
);

NOR4xp25_ASAP7_75t_SL g1294 ( 
.A(n_1237),
.B(n_1158),
.C(n_1192),
.D(n_1209),
.Y(n_1294)
);

INVxp67_ASAP7_75t_L g1295 ( 
.A(n_1264),
.Y(n_1295)
);

AND2x2_ASAP7_75t_L g1296 ( 
.A(n_1236),
.B(n_1207),
.Y(n_1296)
);

AND2x2_ASAP7_75t_L g1297 ( 
.A(n_1238),
.B(n_1207),
.Y(n_1297)
);

AND2x2_ASAP7_75t_L g1298 ( 
.A(n_1238),
.B(n_1207),
.Y(n_1298)
);

OR2x2_ASAP7_75t_L g1299 ( 
.A(n_1235),
.B(n_1169),
.Y(n_1299)
);

HB1xp67_ASAP7_75t_L g1300 ( 
.A(n_1260),
.Y(n_1300)
);

AND2x2_ASAP7_75t_L g1301 ( 
.A(n_1238),
.B(n_1207),
.Y(n_1301)
);

OAI221xp5_ASAP7_75t_L g1302 ( 
.A1(n_1259),
.A2(n_1214),
.B1(n_1217),
.B2(n_1169),
.C(n_1165),
.Y(n_1302)
);

AND2x2_ASAP7_75t_L g1303 ( 
.A(n_1235),
.B(n_1215),
.Y(n_1303)
);

AO21x2_ASAP7_75t_L g1304 ( 
.A1(n_1225),
.A2(n_1202),
.B(n_1213),
.Y(n_1304)
);

NAND2xp5_ASAP7_75t_L g1305 ( 
.A(n_1264),
.B(n_1171),
.Y(n_1305)
);

NAND2xp5_ASAP7_75t_L g1306 ( 
.A(n_1233),
.B(n_1171),
.Y(n_1306)
);

INVx1_ASAP7_75t_L g1307 ( 
.A(n_1231),
.Y(n_1307)
);

OAI211xp5_ASAP7_75t_L g1308 ( 
.A1(n_1263),
.A2(n_1180),
.B(n_1192),
.C(n_1154),
.Y(n_1308)
);

INVx1_ASAP7_75t_L g1309 ( 
.A(n_1231),
.Y(n_1309)
);

INVx3_ASAP7_75t_L g1310 ( 
.A(n_1269),
.Y(n_1310)
);

OR2x2_ASAP7_75t_L g1311 ( 
.A(n_1235),
.B(n_1237),
.Y(n_1311)
);

OR2x2_ASAP7_75t_L g1312 ( 
.A(n_1240),
.B(n_1119),
.Y(n_1312)
);

AND2x2_ASAP7_75t_L g1313 ( 
.A(n_1232),
.B(n_1135),
.Y(n_1313)
);

HB1xp67_ASAP7_75t_L g1314 ( 
.A(n_1252),
.Y(n_1314)
);

AND2x2_ASAP7_75t_L g1315 ( 
.A(n_1232),
.B(n_1135),
.Y(n_1315)
);

INVx2_ASAP7_75t_SL g1316 ( 
.A(n_1242),
.Y(n_1316)
);

AND2x2_ASAP7_75t_L g1317 ( 
.A(n_1232),
.B(n_1183),
.Y(n_1317)
);

AND2x2_ASAP7_75t_L g1318 ( 
.A(n_1226),
.B(n_1183),
.Y(n_1318)
);

HB1xp67_ASAP7_75t_L g1319 ( 
.A(n_1252),
.Y(n_1319)
);

AND2x4_ASAP7_75t_L g1320 ( 
.A(n_1229),
.B(n_1198),
.Y(n_1320)
);

OR2x2_ASAP7_75t_L g1321 ( 
.A(n_1240),
.B(n_1119),
.Y(n_1321)
);

BUFx3_ASAP7_75t_L g1322 ( 
.A(n_1245),
.Y(n_1322)
);

AND2x2_ASAP7_75t_L g1323 ( 
.A(n_1296),
.B(n_1245),
.Y(n_1323)
);

NAND2xp5_ASAP7_75t_L g1324 ( 
.A(n_1283),
.B(n_1267),
.Y(n_1324)
);

AND2x6_ASAP7_75t_L g1325 ( 
.A(n_1291),
.B(n_1255),
.Y(n_1325)
);

OAI221xp5_ASAP7_75t_L g1326 ( 
.A1(n_1293),
.A2(n_1274),
.B1(n_1251),
.B2(n_1234),
.C(n_1273),
.Y(n_1326)
);

NAND2xp5_ASAP7_75t_L g1327 ( 
.A(n_1303),
.B(n_1267),
.Y(n_1327)
);

NAND2xp5_ASAP7_75t_L g1328 ( 
.A(n_1303),
.B(n_1267),
.Y(n_1328)
);

OA211x2_ASAP7_75t_L g1329 ( 
.A1(n_1295),
.A2(n_1230),
.B(n_1255),
.C(n_1258),
.Y(n_1329)
);

OAI21xp5_ASAP7_75t_SL g1330 ( 
.A1(n_1289),
.A2(n_1308),
.B(n_1302),
.Y(n_1330)
);

NAND2xp5_ASAP7_75t_L g1331 ( 
.A(n_1290),
.B(n_1267),
.Y(n_1331)
);

NAND2xp5_ASAP7_75t_L g1332 ( 
.A(n_1312),
.B(n_1247),
.Y(n_1332)
);

NAND2xp5_ASAP7_75t_L g1333 ( 
.A(n_1312),
.B(n_1247),
.Y(n_1333)
);

NAND4xp25_ASAP7_75t_L g1334 ( 
.A(n_1282),
.B(n_1274),
.C(n_1268),
.D(n_1265),
.Y(n_1334)
);

OAI221xp5_ASAP7_75t_SL g1335 ( 
.A1(n_1286),
.A2(n_1274),
.B1(n_1254),
.B2(n_1268),
.C(n_1248),
.Y(n_1335)
);

INVx2_ASAP7_75t_L g1336 ( 
.A(n_1280),
.Y(n_1336)
);

NAND2xp5_ASAP7_75t_L g1337 ( 
.A(n_1321),
.B(n_1247),
.Y(n_1337)
);

AOI211xp5_ASAP7_75t_SL g1338 ( 
.A1(n_1285),
.A2(n_1268),
.B(n_1239),
.C(n_1229),
.Y(n_1338)
);

OAI22xp5_ASAP7_75t_L g1339 ( 
.A1(n_1291),
.A2(n_1230),
.B1(n_1305),
.B2(n_1306),
.Y(n_1339)
);

NAND2xp5_ASAP7_75t_SL g1340 ( 
.A(n_1291),
.B(n_1242),
.Y(n_1340)
);

AND2x2_ASAP7_75t_L g1341 ( 
.A(n_1297),
.B(n_1256),
.Y(n_1341)
);

NAND3xp33_ASAP7_75t_L g1342 ( 
.A(n_1294),
.B(n_1263),
.C(n_1248),
.Y(n_1342)
);

NAND2xp5_ASAP7_75t_L g1343 ( 
.A(n_1288),
.B(n_1247),
.Y(n_1343)
);

NAND2xp5_ASAP7_75t_L g1344 ( 
.A(n_1300),
.B(n_1265),
.Y(n_1344)
);

NOR2xp33_ASAP7_75t_SL g1345 ( 
.A(n_1279),
.B(n_1223),
.Y(n_1345)
);

AND2x2_ASAP7_75t_L g1346 ( 
.A(n_1297),
.B(n_1256),
.Y(n_1346)
);

NAND2xp5_ASAP7_75t_L g1347 ( 
.A(n_1285),
.B(n_1266),
.Y(n_1347)
);

OAI221xp5_ASAP7_75t_L g1348 ( 
.A1(n_1299),
.A2(n_1251),
.B1(n_1234),
.B2(n_1273),
.C(n_1165),
.Y(n_1348)
);

OAI21xp33_ASAP7_75t_L g1349 ( 
.A1(n_1277),
.A2(n_1254),
.B(n_1234),
.Y(n_1349)
);

NOR2x1_ASAP7_75t_L g1350 ( 
.A(n_1304),
.B(n_1272),
.Y(n_1350)
);

NOR2xp33_ASAP7_75t_L g1351 ( 
.A(n_1299),
.B(n_1273),
.Y(n_1351)
);

AND2x2_ASAP7_75t_L g1352 ( 
.A(n_1298),
.B(n_1246),
.Y(n_1352)
);

OR2x2_ASAP7_75t_L g1353 ( 
.A(n_1311),
.B(n_1251),
.Y(n_1353)
);

NAND2xp5_ASAP7_75t_SL g1354 ( 
.A(n_1291),
.B(n_1242),
.Y(n_1354)
);

NAND2xp5_ASAP7_75t_L g1355 ( 
.A(n_1313),
.B(n_1266),
.Y(n_1355)
);

NAND2xp5_ASAP7_75t_L g1356 ( 
.A(n_1313),
.B(n_1246),
.Y(n_1356)
);

AND2x2_ASAP7_75t_L g1357 ( 
.A(n_1301),
.B(n_1246),
.Y(n_1357)
);

NAND2xp5_ASAP7_75t_L g1358 ( 
.A(n_1315),
.B(n_1241),
.Y(n_1358)
);

NAND3xp33_ASAP7_75t_L g1359 ( 
.A(n_1294),
.B(n_1263),
.C(n_1248),
.Y(n_1359)
);

NAND3xp33_ASAP7_75t_L g1360 ( 
.A(n_1278),
.B(n_1263),
.C(n_1241),
.Y(n_1360)
);

NAND2xp5_ASAP7_75t_SL g1361 ( 
.A(n_1291),
.B(n_1242),
.Y(n_1361)
);

NAND2xp5_ASAP7_75t_L g1362 ( 
.A(n_1315),
.B(n_1228),
.Y(n_1362)
);

NAND3xp33_ASAP7_75t_L g1363 ( 
.A(n_1278),
.B(n_1263),
.C(n_1242),
.Y(n_1363)
);

AND2x2_ASAP7_75t_L g1364 ( 
.A(n_1284),
.B(n_1239),
.Y(n_1364)
);

AOI221xp5_ASAP7_75t_L g1365 ( 
.A1(n_1277),
.A2(n_1270),
.B1(n_1271),
.B2(n_1276),
.C(n_1275),
.Y(n_1365)
);

AOI21xp5_ASAP7_75t_SL g1366 ( 
.A1(n_1320),
.A2(n_1249),
.B(n_1258),
.Y(n_1366)
);

OAI22xp5_ASAP7_75t_L g1367 ( 
.A1(n_1311),
.A2(n_1230),
.B1(n_1254),
.B2(n_1262),
.Y(n_1367)
);

AND2x4_ASAP7_75t_L g1368 ( 
.A(n_1340),
.B(n_1322),
.Y(n_1368)
);

INVx2_ASAP7_75t_L g1369 ( 
.A(n_1336),
.Y(n_1369)
);

AND2x4_ASAP7_75t_L g1370 ( 
.A(n_1340),
.B(n_1310),
.Y(n_1370)
);

INVx1_ASAP7_75t_SL g1371 ( 
.A(n_1353),
.Y(n_1371)
);

AND2x2_ASAP7_75t_L g1372 ( 
.A(n_1364),
.B(n_1287),
.Y(n_1372)
);

AND2x2_ASAP7_75t_L g1373 ( 
.A(n_1323),
.B(n_1292),
.Y(n_1373)
);

BUFx3_ASAP7_75t_L g1374 ( 
.A(n_1325),
.Y(n_1374)
);

INVx1_ASAP7_75t_L g1375 ( 
.A(n_1344),
.Y(n_1375)
);

INVx1_ASAP7_75t_L g1376 ( 
.A(n_1347),
.Y(n_1376)
);

AND2x4_ASAP7_75t_L g1377 ( 
.A(n_1354),
.B(n_1310),
.Y(n_1377)
);

INVx2_ASAP7_75t_L g1378 ( 
.A(n_1327),
.Y(n_1378)
);

OR2x2_ASAP7_75t_L g1379 ( 
.A(n_1328),
.B(n_1324),
.Y(n_1379)
);

NOR2xp33_ASAP7_75t_L g1380 ( 
.A(n_1345),
.B(n_1121),
.Y(n_1380)
);

NAND2xp5_ASAP7_75t_L g1381 ( 
.A(n_1331),
.B(n_1314),
.Y(n_1381)
);

INVx1_ASAP7_75t_L g1382 ( 
.A(n_1355),
.Y(n_1382)
);

INVx2_ASAP7_75t_L g1383 ( 
.A(n_1350),
.Y(n_1383)
);

INVx1_ASAP7_75t_L g1384 ( 
.A(n_1362),
.Y(n_1384)
);

INVx1_ASAP7_75t_L g1385 ( 
.A(n_1343),
.Y(n_1385)
);

NAND2xp5_ASAP7_75t_L g1386 ( 
.A(n_1358),
.B(n_1319),
.Y(n_1386)
);

INVx1_ASAP7_75t_SL g1387 ( 
.A(n_1341),
.Y(n_1387)
);

NAND2xp5_ASAP7_75t_L g1388 ( 
.A(n_1332),
.B(n_1333),
.Y(n_1388)
);

OR2x2_ASAP7_75t_L g1389 ( 
.A(n_1337),
.B(n_1356),
.Y(n_1389)
);

INVx2_ASAP7_75t_L g1390 ( 
.A(n_1346),
.Y(n_1390)
);

AND2x4_ASAP7_75t_SL g1391 ( 
.A(n_1346),
.B(n_1320),
.Y(n_1391)
);

NOR2xp33_ASAP7_75t_L g1392 ( 
.A(n_1330),
.B(n_1121),
.Y(n_1392)
);

INVx2_ASAP7_75t_L g1393 ( 
.A(n_1352),
.Y(n_1393)
);

NAND2xp5_ASAP7_75t_L g1394 ( 
.A(n_1365),
.B(n_1307),
.Y(n_1394)
);

OR2x2_ASAP7_75t_L g1395 ( 
.A(n_1363),
.B(n_1316),
.Y(n_1395)
);

AND2x2_ASAP7_75t_L g1396 ( 
.A(n_1352),
.B(n_1281),
.Y(n_1396)
);

OR2x2_ASAP7_75t_L g1397 ( 
.A(n_1360),
.B(n_1280),
.Y(n_1397)
);

INVx1_ASAP7_75t_L g1398 ( 
.A(n_1357),
.Y(n_1398)
);

INVx1_ASAP7_75t_L g1399 ( 
.A(n_1357),
.Y(n_1399)
);

NOR2xp67_ASAP7_75t_L g1400 ( 
.A(n_1395),
.B(n_1339),
.Y(n_1400)
);

NAND2xp5_ASAP7_75t_L g1401 ( 
.A(n_1375),
.B(n_1351),
.Y(n_1401)
);

HB1xp67_ASAP7_75t_L g1402 ( 
.A(n_1381),
.Y(n_1402)
);

INVx2_ASAP7_75t_L g1403 ( 
.A(n_1369),
.Y(n_1403)
);

NAND2xp5_ASAP7_75t_L g1404 ( 
.A(n_1375),
.B(n_1334),
.Y(n_1404)
);

NOR4xp75_ASAP7_75t_L g1405 ( 
.A(n_1394),
.B(n_1348),
.C(n_1326),
.D(n_1361),
.Y(n_1405)
);

OR2x2_ASAP7_75t_L g1406 ( 
.A(n_1379),
.B(n_1366),
.Y(n_1406)
);

NAND2xp5_ASAP7_75t_L g1407 ( 
.A(n_1376),
.B(n_1317),
.Y(n_1407)
);

INVx1_ASAP7_75t_L g1408 ( 
.A(n_1369),
.Y(n_1408)
);

NAND2xp5_ASAP7_75t_L g1409 ( 
.A(n_1376),
.B(n_1317),
.Y(n_1409)
);

AND2x2_ASAP7_75t_L g1410 ( 
.A(n_1391),
.B(n_1338),
.Y(n_1410)
);

INVx1_ASAP7_75t_L g1411 ( 
.A(n_1369),
.Y(n_1411)
);

INVx1_ASAP7_75t_L g1412 ( 
.A(n_1381),
.Y(n_1412)
);

INVx2_ASAP7_75t_SL g1413 ( 
.A(n_1391),
.Y(n_1413)
);

INVx2_ASAP7_75t_SL g1414 ( 
.A(n_1391),
.Y(n_1414)
);

AND2x2_ASAP7_75t_L g1415 ( 
.A(n_1396),
.B(n_1361),
.Y(n_1415)
);

AND2x2_ASAP7_75t_L g1416 ( 
.A(n_1396),
.B(n_1367),
.Y(n_1416)
);

INVx1_ASAP7_75t_L g1417 ( 
.A(n_1397),
.Y(n_1417)
);

INVx2_ASAP7_75t_L g1418 ( 
.A(n_1397),
.Y(n_1418)
);

INVx1_ASAP7_75t_L g1419 ( 
.A(n_1398),
.Y(n_1419)
);

INVx1_ASAP7_75t_L g1420 ( 
.A(n_1398),
.Y(n_1420)
);

AND2x2_ASAP7_75t_L g1421 ( 
.A(n_1393),
.B(n_1349),
.Y(n_1421)
);

NAND2xp5_ASAP7_75t_L g1422 ( 
.A(n_1385),
.B(n_1318),
.Y(n_1422)
);

OR2x2_ASAP7_75t_L g1423 ( 
.A(n_1379),
.B(n_1342),
.Y(n_1423)
);

INVx2_ASAP7_75t_L g1424 ( 
.A(n_1383),
.Y(n_1424)
);

OR2x2_ASAP7_75t_L g1425 ( 
.A(n_1378),
.B(n_1359),
.Y(n_1425)
);

AND2x2_ASAP7_75t_L g1426 ( 
.A(n_1393),
.B(n_1390),
.Y(n_1426)
);

NOR2xp33_ASAP7_75t_L g1427 ( 
.A(n_1392),
.B(n_1126),
.Y(n_1427)
);

INVx1_ASAP7_75t_L g1428 ( 
.A(n_1399),
.Y(n_1428)
);

INVx1_ASAP7_75t_L g1429 ( 
.A(n_1399),
.Y(n_1429)
);

INVx1_ASAP7_75t_L g1430 ( 
.A(n_1382),
.Y(n_1430)
);

INVx1_ASAP7_75t_L g1431 ( 
.A(n_1382),
.Y(n_1431)
);

INVx1_ASAP7_75t_L g1432 ( 
.A(n_1394),
.Y(n_1432)
);

NAND2xp5_ASAP7_75t_L g1433 ( 
.A(n_1384),
.B(n_1307),
.Y(n_1433)
);

NAND2xp5_ASAP7_75t_L g1434 ( 
.A(n_1384),
.B(n_1309),
.Y(n_1434)
);

NAND2xp5_ASAP7_75t_L g1435 ( 
.A(n_1432),
.B(n_1378),
.Y(n_1435)
);

INVx2_ASAP7_75t_L g1436 ( 
.A(n_1403),
.Y(n_1436)
);

OR2x2_ASAP7_75t_L g1437 ( 
.A(n_1423),
.B(n_1378),
.Y(n_1437)
);

NOR2x2_ASAP7_75t_L g1438 ( 
.A(n_1418),
.B(n_1383),
.Y(n_1438)
);

OR2x2_ASAP7_75t_L g1439 ( 
.A(n_1423),
.B(n_1425),
.Y(n_1439)
);

INVx2_ASAP7_75t_L g1440 ( 
.A(n_1403),
.Y(n_1440)
);

INVx2_ASAP7_75t_L g1441 ( 
.A(n_1424),
.Y(n_1441)
);

NAND2x1_ASAP7_75t_L g1442 ( 
.A(n_1410),
.B(n_1368),
.Y(n_1442)
);

INVx1_ASAP7_75t_L g1443 ( 
.A(n_1430),
.Y(n_1443)
);

INVx1_ASAP7_75t_L g1444 ( 
.A(n_1430),
.Y(n_1444)
);

INVx1_ASAP7_75t_L g1445 ( 
.A(n_1431),
.Y(n_1445)
);

INVx1_ASAP7_75t_L g1446 ( 
.A(n_1419),
.Y(n_1446)
);

INVx2_ASAP7_75t_L g1447 ( 
.A(n_1424),
.Y(n_1447)
);

NAND2xp5_ASAP7_75t_L g1448 ( 
.A(n_1432),
.B(n_1371),
.Y(n_1448)
);

OR2x2_ASAP7_75t_L g1449 ( 
.A(n_1425),
.B(n_1395),
.Y(n_1449)
);

CKINVDCx16_ASAP7_75t_R g1450 ( 
.A(n_1427),
.Y(n_1450)
);

INVx2_ASAP7_75t_L g1451 ( 
.A(n_1408),
.Y(n_1451)
);

INVx1_ASAP7_75t_L g1452 ( 
.A(n_1431),
.Y(n_1452)
);

AOI22xp33_ASAP7_75t_L g1453 ( 
.A1(n_1404),
.A2(n_1380),
.B1(n_1374),
.B2(n_1368),
.Y(n_1453)
);

AND2x4_ASAP7_75t_L g1454 ( 
.A(n_1413),
.B(n_1374),
.Y(n_1454)
);

NAND2xp5_ASAP7_75t_L g1455 ( 
.A(n_1402),
.B(n_1371),
.Y(n_1455)
);

NAND2xp5_ASAP7_75t_L g1456 ( 
.A(n_1412),
.B(n_1373),
.Y(n_1456)
);

INVxp67_ASAP7_75t_L g1457 ( 
.A(n_1401),
.Y(n_1457)
);

INVx1_ASAP7_75t_L g1458 ( 
.A(n_1419),
.Y(n_1458)
);

OR2x2_ASAP7_75t_L g1459 ( 
.A(n_1418),
.B(n_1417),
.Y(n_1459)
);

NOR2x1p5_ASAP7_75t_SL g1460 ( 
.A(n_1406),
.B(n_1383),
.Y(n_1460)
);

AOI21xp5_ASAP7_75t_L g1461 ( 
.A1(n_1400),
.A2(n_1335),
.B(n_1374),
.Y(n_1461)
);

AOI21xp33_ASAP7_75t_L g1462 ( 
.A1(n_1406),
.A2(n_1377),
.B(n_1370),
.Y(n_1462)
);

OAI21xp5_ASAP7_75t_L g1463 ( 
.A1(n_1412),
.A2(n_1368),
.B(n_1370),
.Y(n_1463)
);

AND2x2_ASAP7_75t_L g1464 ( 
.A(n_1410),
.B(n_1387),
.Y(n_1464)
);

OR2x2_ASAP7_75t_L g1465 ( 
.A(n_1417),
.B(n_1389),
.Y(n_1465)
);

NAND2xp5_ASAP7_75t_L g1466 ( 
.A(n_1421),
.B(n_1373),
.Y(n_1466)
);

INVx2_ASAP7_75t_L g1467 ( 
.A(n_1408),
.Y(n_1467)
);

INVx2_ASAP7_75t_L g1468 ( 
.A(n_1411),
.Y(n_1468)
);

INVx1_ASAP7_75t_L g1469 ( 
.A(n_1420),
.Y(n_1469)
);

NAND2xp5_ASAP7_75t_L g1470 ( 
.A(n_1421),
.B(n_1390),
.Y(n_1470)
);

OAI211xp5_ASAP7_75t_L g1471 ( 
.A1(n_1405),
.A2(n_1386),
.B(n_1387),
.C(n_1388),
.Y(n_1471)
);

INVx1_ASAP7_75t_L g1472 ( 
.A(n_1420),
.Y(n_1472)
);

INVx1_ASAP7_75t_L g1473 ( 
.A(n_1428),
.Y(n_1473)
);

AND2x2_ASAP7_75t_L g1474 ( 
.A(n_1413),
.B(n_1372),
.Y(n_1474)
);

INVx1_ASAP7_75t_L g1475 ( 
.A(n_1428),
.Y(n_1475)
);

AOI21xp33_ASAP7_75t_L g1476 ( 
.A1(n_1429),
.A2(n_1377),
.B(n_1370),
.Y(n_1476)
);

AND2x2_ASAP7_75t_L g1477 ( 
.A(n_1414),
.B(n_1415),
.Y(n_1477)
);

NAND2xp5_ASAP7_75t_SL g1478 ( 
.A(n_1450),
.B(n_1414),
.Y(n_1478)
);

NAND2xp5_ASAP7_75t_L g1479 ( 
.A(n_1457),
.B(n_1415),
.Y(n_1479)
);

INVx1_ASAP7_75t_SL g1480 ( 
.A(n_1439),
.Y(n_1480)
);

AND2x2_ASAP7_75t_L g1481 ( 
.A(n_1477),
.B(n_1416),
.Y(n_1481)
);

BUFx3_ASAP7_75t_L g1482 ( 
.A(n_1442),
.Y(n_1482)
);

OAI22xp5_ASAP7_75t_L g1483 ( 
.A1(n_1471),
.A2(n_1329),
.B1(n_1368),
.B2(n_1416),
.Y(n_1483)
);

HB1xp67_ASAP7_75t_L g1484 ( 
.A(n_1439),
.Y(n_1484)
);

INVx1_ASAP7_75t_L g1485 ( 
.A(n_1446),
.Y(n_1485)
);

AND2x2_ASAP7_75t_L g1486 ( 
.A(n_1477),
.B(n_1426),
.Y(n_1486)
);

OR2x2_ASAP7_75t_L g1487 ( 
.A(n_1449),
.B(n_1429),
.Y(n_1487)
);

INVx1_ASAP7_75t_L g1488 ( 
.A(n_1446),
.Y(n_1488)
);

INVx2_ASAP7_75t_L g1489 ( 
.A(n_1438),
.Y(n_1489)
);

AND2x4_ASAP7_75t_L g1490 ( 
.A(n_1454),
.B(n_1460),
.Y(n_1490)
);

AND2x2_ASAP7_75t_L g1491 ( 
.A(n_1464),
.B(n_1454),
.Y(n_1491)
);

INVx1_ASAP7_75t_SL g1492 ( 
.A(n_1438),
.Y(n_1492)
);

INVx2_ASAP7_75t_L g1493 ( 
.A(n_1459),
.Y(n_1493)
);

INVx1_ASAP7_75t_SL g1494 ( 
.A(n_1454),
.Y(n_1494)
);

INVxp67_ASAP7_75t_L g1495 ( 
.A(n_1449),
.Y(n_1495)
);

OR2x2_ASAP7_75t_L g1496 ( 
.A(n_1465),
.B(n_1433),
.Y(n_1496)
);

OR2x2_ASAP7_75t_L g1497 ( 
.A(n_1465),
.B(n_1459),
.Y(n_1497)
);

NAND2xp5_ASAP7_75t_L g1498 ( 
.A(n_1461),
.B(n_1407),
.Y(n_1498)
);

INVx1_ASAP7_75t_L g1499 ( 
.A(n_1458),
.Y(n_1499)
);

BUFx3_ASAP7_75t_L g1500 ( 
.A(n_1442),
.Y(n_1500)
);

INVx2_ASAP7_75t_L g1501 ( 
.A(n_1451),
.Y(n_1501)
);

INVx1_ASAP7_75t_L g1502 ( 
.A(n_1469),
.Y(n_1502)
);

HB1xp67_ASAP7_75t_L g1503 ( 
.A(n_1464),
.Y(n_1503)
);

INVx1_ASAP7_75t_L g1504 ( 
.A(n_1472),
.Y(n_1504)
);

OR2x2_ASAP7_75t_L g1505 ( 
.A(n_1437),
.B(n_1434),
.Y(n_1505)
);

NAND2x1p5_ASAP7_75t_L g1506 ( 
.A(n_1437),
.B(n_1258),
.Y(n_1506)
);

INVx1_ASAP7_75t_L g1507 ( 
.A(n_1473),
.Y(n_1507)
);

INVx1_ASAP7_75t_SL g1508 ( 
.A(n_1455),
.Y(n_1508)
);

INVx1_ASAP7_75t_SL g1509 ( 
.A(n_1448),
.Y(n_1509)
);

INVx2_ASAP7_75t_L g1510 ( 
.A(n_1451),
.Y(n_1510)
);

INVx1_ASAP7_75t_SL g1511 ( 
.A(n_1474),
.Y(n_1511)
);

INVx3_ASAP7_75t_SL g1512 ( 
.A(n_1474),
.Y(n_1512)
);

AND2x2_ASAP7_75t_L g1513 ( 
.A(n_1463),
.B(n_1426),
.Y(n_1513)
);

INVx1_ASAP7_75t_L g1514 ( 
.A(n_1484),
.Y(n_1514)
);

AND2x2_ASAP7_75t_L g1515 ( 
.A(n_1491),
.B(n_1453),
.Y(n_1515)
);

INVxp67_ASAP7_75t_L g1516 ( 
.A(n_1503),
.Y(n_1516)
);

AO221x1_ASAP7_75t_L g1517 ( 
.A1(n_1483),
.A2(n_1475),
.B1(n_1443),
.B2(n_1452),
.C(n_1445),
.Y(n_1517)
);

NOR2xp67_ASAP7_75t_L g1518 ( 
.A(n_1490),
.B(n_1466),
.Y(n_1518)
);

NOR3xp33_ASAP7_75t_L g1519 ( 
.A(n_1478),
.B(n_1462),
.C(n_1476),
.Y(n_1519)
);

AND2x2_ASAP7_75t_L g1520 ( 
.A(n_1491),
.B(n_1512),
.Y(n_1520)
);

NAND3xp33_ASAP7_75t_L g1521 ( 
.A(n_1495),
.B(n_1444),
.C(n_1435),
.Y(n_1521)
);

NAND3x2_ASAP7_75t_L g1522 ( 
.A(n_1490),
.B(n_1460),
.C(n_1377),
.Y(n_1522)
);

NAND2xp5_ASAP7_75t_L g1523 ( 
.A(n_1480),
.B(n_1456),
.Y(n_1523)
);

NOR2xp33_ASAP7_75t_L g1524 ( 
.A(n_1508),
.B(n_1134),
.Y(n_1524)
);

INVx2_ASAP7_75t_L g1525 ( 
.A(n_1490),
.Y(n_1525)
);

INVx2_ASAP7_75t_L g1526 ( 
.A(n_1490),
.Y(n_1526)
);

NAND3xp33_ASAP7_75t_L g1527 ( 
.A(n_1498),
.B(n_1447),
.C(n_1441),
.Y(n_1527)
);

INVx1_ASAP7_75t_L g1528 ( 
.A(n_1485),
.Y(n_1528)
);

INVx2_ASAP7_75t_L g1529 ( 
.A(n_1512),
.Y(n_1529)
);

NAND2xp5_ASAP7_75t_L g1530 ( 
.A(n_1509),
.B(n_1470),
.Y(n_1530)
);

INVx1_ASAP7_75t_L g1531 ( 
.A(n_1485),
.Y(n_1531)
);

INVx3_ASAP7_75t_L g1532 ( 
.A(n_1482),
.Y(n_1532)
);

OAI221xp5_ASAP7_75t_L g1533 ( 
.A1(n_1492),
.A2(n_1447),
.B1(n_1441),
.B2(n_1440),
.C(n_1436),
.Y(n_1533)
);

OR2x2_ASAP7_75t_L g1534 ( 
.A(n_1479),
.B(n_1422),
.Y(n_1534)
);

NAND2xp5_ASAP7_75t_L g1535 ( 
.A(n_1509),
.B(n_1409),
.Y(n_1535)
);

INVx1_ASAP7_75t_L g1536 ( 
.A(n_1488),
.Y(n_1536)
);

OAI221xp5_ASAP7_75t_L g1537 ( 
.A1(n_1492),
.A2(n_1440),
.B1(n_1436),
.B2(n_1468),
.C(n_1467),
.Y(n_1537)
);

OR2x2_ASAP7_75t_L g1538 ( 
.A(n_1497),
.B(n_1467),
.Y(n_1538)
);

NAND2xp5_ASAP7_75t_SL g1539 ( 
.A(n_1518),
.B(n_1482),
.Y(n_1539)
);

AND2x2_ASAP7_75t_L g1540 ( 
.A(n_1520),
.B(n_1512),
.Y(n_1540)
);

AOI22xp33_ASAP7_75t_L g1541 ( 
.A1(n_1517),
.A2(n_1489),
.B1(n_1494),
.B2(n_1511),
.Y(n_1541)
);

INVxp67_ASAP7_75t_L g1542 ( 
.A(n_1520),
.Y(n_1542)
);

BUFx2_ASAP7_75t_L g1543 ( 
.A(n_1532),
.Y(n_1543)
);

INVx1_ASAP7_75t_L g1544 ( 
.A(n_1528),
.Y(n_1544)
);

NOR2xp33_ASAP7_75t_L g1545 ( 
.A(n_1524),
.B(n_1482),
.Y(n_1545)
);

NAND2xp5_ASAP7_75t_L g1546 ( 
.A(n_1529),
.B(n_1516),
.Y(n_1546)
);

XOR2xp5_ASAP7_75t_L g1547 ( 
.A(n_1515),
.B(n_1136),
.Y(n_1547)
);

NAND2xp5_ASAP7_75t_L g1548 ( 
.A(n_1529),
.B(n_1481),
.Y(n_1548)
);

OR2x2_ASAP7_75t_L g1549 ( 
.A(n_1514),
.B(n_1497),
.Y(n_1549)
);

INVx1_ASAP7_75t_L g1550 ( 
.A(n_1531),
.Y(n_1550)
);

NOR2xp33_ASAP7_75t_L g1551 ( 
.A(n_1524),
.B(n_1515),
.Y(n_1551)
);

NAND2xp5_ASAP7_75t_L g1552 ( 
.A(n_1525),
.B(n_1481),
.Y(n_1552)
);

INVx1_ASAP7_75t_L g1553 ( 
.A(n_1536),
.Y(n_1553)
);

NAND2xp5_ASAP7_75t_L g1554 ( 
.A(n_1525),
.B(n_1489),
.Y(n_1554)
);

INVx2_ASAP7_75t_L g1555 ( 
.A(n_1532),
.Y(n_1555)
);

INVx1_ASAP7_75t_L g1556 ( 
.A(n_1538),
.Y(n_1556)
);

OR2x2_ASAP7_75t_L g1557 ( 
.A(n_1530),
.B(n_1493),
.Y(n_1557)
);

O2A1O1Ixp33_ASAP7_75t_L g1558 ( 
.A1(n_1539),
.A2(n_1519),
.B(n_1537),
.C(n_1533),
.Y(n_1558)
);

AOI22xp5_ASAP7_75t_L g1559 ( 
.A1(n_1545),
.A2(n_1522),
.B1(n_1523),
.B2(n_1526),
.Y(n_1559)
);

AO21x1_ASAP7_75t_L g1560 ( 
.A1(n_1539),
.A2(n_1526),
.B(n_1489),
.Y(n_1560)
);

NAND3xp33_ASAP7_75t_L g1561 ( 
.A(n_1541),
.B(n_1527),
.C(n_1532),
.Y(n_1561)
);

NAND2xp5_ASAP7_75t_SL g1562 ( 
.A(n_1551),
.B(n_1545),
.Y(n_1562)
);

NAND2xp5_ASAP7_75t_L g1563 ( 
.A(n_1542),
.B(n_1486),
.Y(n_1563)
);

OAI211xp5_ASAP7_75t_SL g1564 ( 
.A1(n_1551),
.A2(n_1535),
.B(n_1521),
.C(n_1534),
.Y(n_1564)
);

INVx1_ASAP7_75t_L g1565 ( 
.A(n_1543),
.Y(n_1565)
);

AO21x1_ASAP7_75t_L g1566 ( 
.A1(n_1555),
.A2(n_1506),
.B(n_1488),
.Y(n_1566)
);

AOI21xp5_ASAP7_75t_L g1567 ( 
.A1(n_1547),
.A2(n_1493),
.B(n_1538),
.Y(n_1567)
);

NOR2xp33_ASAP7_75t_L g1568 ( 
.A(n_1546),
.B(n_1134),
.Y(n_1568)
);

NAND3xp33_ASAP7_75t_SL g1569 ( 
.A(n_1558),
.B(n_1541),
.C(n_1540),
.Y(n_1569)
);

NAND2xp5_ASAP7_75t_L g1570 ( 
.A(n_1565),
.B(n_1562),
.Y(n_1570)
);

INVxp67_ASAP7_75t_L g1571 ( 
.A(n_1568),
.Y(n_1571)
);

INVx1_ASAP7_75t_L g1572 ( 
.A(n_1563),
.Y(n_1572)
);

NOR2x1_ASAP7_75t_L g1573 ( 
.A(n_1561),
.B(n_1554),
.Y(n_1573)
);

INVx1_ASAP7_75t_L g1574 ( 
.A(n_1560),
.Y(n_1574)
);

AND2x2_ASAP7_75t_L g1575 ( 
.A(n_1559),
.B(n_1548),
.Y(n_1575)
);

NOR3xp33_ASAP7_75t_L g1576 ( 
.A(n_1564),
.B(n_1552),
.C(n_1549),
.Y(n_1576)
);

NAND3xp33_ASAP7_75t_SL g1577 ( 
.A(n_1566),
.B(n_1557),
.C(n_1556),
.Y(n_1577)
);

NAND2xp5_ASAP7_75t_L g1578 ( 
.A(n_1567),
.B(n_1544),
.Y(n_1578)
);

NAND2xp5_ASAP7_75t_SL g1579 ( 
.A(n_1573),
.B(n_1500),
.Y(n_1579)
);

AOI31xp33_ASAP7_75t_L g1580 ( 
.A1(n_1577),
.A2(n_1553),
.A3(n_1550),
.B(n_1506),
.Y(n_1580)
);

AOI22xp5_ASAP7_75t_L g1581 ( 
.A1(n_1569),
.A2(n_1500),
.B1(n_1493),
.B2(n_1499),
.Y(n_1581)
);

AOI211xp5_ASAP7_75t_L g1582 ( 
.A1(n_1576),
.A2(n_1500),
.B(n_1513),
.C(n_1499),
.Y(n_1582)
);

NOR2xp33_ASAP7_75t_SL g1583 ( 
.A(n_1570),
.B(n_1126),
.Y(n_1583)
);

NOR3x1_ASAP7_75t_L g1584 ( 
.A(n_1578),
.B(n_1504),
.C(n_1502),
.Y(n_1584)
);

INVx1_ASAP7_75t_L g1585 ( 
.A(n_1584),
.Y(n_1585)
);

AOI22xp5_ASAP7_75t_L g1586 ( 
.A1(n_1583),
.A2(n_1574),
.B1(n_1575),
.B2(n_1571),
.Y(n_1586)
);

OAI22xp33_ASAP7_75t_L g1587 ( 
.A1(n_1580),
.A2(n_1506),
.B1(n_1572),
.B2(n_1502),
.Y(n_1587)
);

INVx1_ASAP7_75t_L g1588 ( 
.A(n_1579),
.Y(n_1588)
);

INVx1_ASAP7_75t_L g1589 ( 
.A(n_1581),
.Y(n_1589)
);

AOI22xp5_ASAP7_75t_L g1590 ( 
.A1(n_1582),
.A2(n_1504),
.B1(n_1507),
.B2(n_1513),
.Y(n_1590)
);

INVx1_ASAP7_75t_L g1591 ( 
.A(n_1584),
.Y(n_1591)
);

INVx2_ASAP7_75t_L g1592 ( 
.A(n_1588),
.Y(n_1592)
);

CKINVDCx5p33_ASAP7_75t_R g1593 ( 
.A(n_1586),
.Y(n_1593)
);

NOR3xp33_ASAP7_75t_SL g1594 ( 
.A(n_1589),
.B(n_1507),
.C(n_1168),
.Y(n_1594)
);

NAND3xp33_ASAP7_75t_SL g1595 ( 
.A(n_1585),
.B(n_1136),
.C(n_1487),
.Y(n_1595)
);

INVx1_ASAP7_75t_L g1596 ( 
.A(n_1591),
.Y(n_1596)
);

XNOR2x2_ASAP7_75t_SL g1597 ( 
.A(n_1596),
.B(n_1590),
.Y(n_1597)
);

OR2x2_ASAP7_75t_L g1598 ( 
.A(n_1592),
.B(n_1587),
.Y(n_1598)
);

XNOR2x1_ASAP7_75t_SL g1599 ( 
.A(n_1593),
.B(n_1168),
.Y(n_1599)
);

INVx2_ASAP7_75t_L g1600 ( 
.A(n_1598),
.Y(n_1600)
);

NAND5xp2_ASAP7_75t_L g1601 ( 
.A(n_1600),
.B(n_1594),
.C(n_1599),
.D(n_1597),
.E(n_1595),
.Y(n_1601)
);

NAND2xp5_ASAP7_75t_L g1602 ( 
.A(n_1601),
.B(n_1592),
.Y(n_1602)
);

INVx1_ASAP7_75t_L g1603 ( 
.A(n_1601),
.Y(n_1603)
);

XOR2xp5_ASAP7_75t_L g1604 ( 
.A(n_1603),
.B(n_1602),
.Y(n_1604)
);

OAI21xp5_ASAP7_75t_L g1605 ( 
.A1(n_1602),
.A2(n_1510),
.B(n_1501),
.Y(n_1605)
);

NAND2xp5_ASAP7_75t_L g1606 ( 
.A(n_1604),
.B(n_1501),
.Y(n_1606)
);

AO21x1_ASAP7_75t_L g1607 ( 
.A1(n_1605),
.A2(n_1510),
.B(n_1501),
.Y(n_1607)
);

NAND3xp33_ASAP7_75t_L g1608 ( 
.A(n_1606),
.B(n_1154),
.C(n_1510),
.Y(n_1608)
);

AOI222xp33_ASAP7_75t_L g1609 ( 
.A1(n_1608),
.A2(n_1607),
.B1(n_1486),
.B2(n_1468),
.C1(n_1165),
.C2(n_1411),
.Y(n_1609)
);

OAI221xp5_ASAP7_75t_R g1610 ( 
.A1(n_1609),
.A2(n_1487),
.B1(n_1208),
.B2(n_1505),
.C(n_1496),
.Y(n_1610)
);

AOI211xp5_ASAP7_75t_L g1611 ( 
.A1(n_1610),
.A2(n_1505),
.B(n_1496),
.C(n_1211),
.Y(n_1611)
);


endmodule