module fake_ariane_1157_n_1138 (n_83, n_8, n_56, n_60, n_170, n_190, n_160, n_64, n_179, n_180, n_119, n_124, n_167, n_90, n_195, n_38, n_213, n_47, n_110, n_153, n_18, n_197, n_221, n_86, n_75, n_89, n_67, n_176, n_149, n_34, n_158, n_172, n_69, n_95, n_175, n_92, n_143, n_183, n_203, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_181, n_152, n_120, n_169, n_106, n_12, n_53, n_173, n_111, n_21, n_115, n_133, n_66, n_205, n_71, n_24, n_7, n_109, n_208, n_96, n_156, n_209, n_49, n_20, n_174, n_100, n_17, n_50, n_187, n_132, n_62, n_210, n_147, n_204, n_200, n_51, n_166, n_76, n_218, n_103, n_79, n_26, n_3, n_46, n_220, n_0, n_84, n_36, n_199, n_91, n_159, n_107, n_189, n_72, n_105, n_128, n_217, n_44, n_30, n_82, n_178, n_31, n_42, n_57, n_131, n_201, n_70, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_6, n_214, n_48, n_94, n_101, n_4, n_134, n_188, n_185, n_2, n_32, n_37, n_58, n_65, n_123, n_212, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_198, n_148, n_164, n_52, n_157, n_184, n_177, n_135, n_73, n_77, n_171, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_182, n_196, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_206, n_13, n_27, n_207, n_29, n_41, n_219, n_140, n_55, n_191, n_151, n_136, n_192, n_28, n_80, n_146, n_211, n_194, n_97, n_154, n_215, n_142, n_161, n_14, n_163, n_88, n_186, n_141, n_68, n_116, n_104, n_202, n_145, n_78, n_193, n_39, n_59, n_63, n_99, n_216, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_1138);

input n_83;
input n_8;
input n_56;
input n_60;
input n_170;
input n_190;
input n_160;
input n_64;
input n_179;
input n_180;
input n_119;
input n_124;
input n_167;
input n_90;
input n_195;
input n_38;
input n_213;
input n_47;
input n_110;
input n_153;
input n_18;
input n_197;
input n_221;
input n_86;
input n_75;
input n_89;
input n_67;
input n_176;
input n_149;
input n_34;
input n_158;
input n_172;
input n_69;
input n_95;
input n_175;
input n_92;
input n_143;
input n_183;
input n_203;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_181;
input n_152;
input n_120;
input n_169;
input n_106;
input n_12;
input n_53;
input n_173;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_205;
input n_71;
input n_24;
input n_7;
input n_109;
input n_208;
input n_96;
input n_156;
input n_209;
input n_49;
input n_20;
input n_174;
input n_100;
input n_17;
input n_50;
input n_187;
input n_132;
input n_62;
input n_210;
input n_147;
input n_204;
input n_200;
input n_51;
input n_166;
input n_76;
input n_218;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_220;
input n_0;
input n_84;
input n_36;
input n_199;
input n_91;
input n_159;
input n_107;
input n_189;
input n_72;
input n_105;
input n_128;
input n_217;
input n_44;
input n_30;
input n_82;
input n_178;
input n_31;
input n_42;
input n_57;
input n_131;
input n_201;
input n_70;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_6;
input n_214;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_188;
input n_185;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_212;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_198;
input n_148;
input n_164;
input n_52;
input n_157;
input n_184;
input n_177;
input n_135;
input n_73;
input n_77;
input n_171;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_182;
input n_196;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_206;
input n_13;
input n_27;
input n_207;
input n_29;
input n_41;
input n_219;
input n_140;
input n_55;
input n_191;
input n_151;
input n_136;
input n_192;
input n_28;
input n_80;
input n_146;
input n_211;
input n_194;
input n_97;
input n_154;
input n_215;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_186;
input n_141;
input n_68;
input n_116;
input n_104;
input n_202;
input n_145;
input n_78;
input n_193;
input n_39;
input n_59;
input n_63;
input n_99;
input n_216;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_1138;

wire n_295;
wire n_356;
wire n_556;
wire n_698;
wire n_1127;
wire n_1072;
wire n_695;
wire n_913;
wire n_730;
wire n_386;
wire n_307;
wire n_516;
wire n_589;
wire n_332;
wire n_1008;
wire n_581;
wire n_294;
wire n_1020;
wire n_1137;
wire n_646;
wire n_640;
wire n_463;
wire n_1024;
wire n_830;
wire n_691;
wire n_404;
wire n_943;
wire n_1118;
wire n_678;
wire n_1058;
wire n_651;
wire n_987;
wire n_936;
wire n_347;
wire n_423;
wire n_1042;
wire n_961;
wire n_469;
wire n_1046;
wire n_479;
wire n_726;
wire n_603;
wire n_1123;
wire n_878;
wire n_373;
wire n_299;
wire n_836;
wire n_541;
wire n_499;
wire n_789;
wire n_788;
wire n_850;
wire n_908;
wire n_771;
wire n_1036;
wire n_564;
wire n_610;
wire n_752;
wire n_341;
wire n_1029;
wire n_985;
wire n_421;
wire n_245;
wire n_549;
wire n_522;
wire n_319;
wire n_591;
wire n_760;
wire n_690;
wire n_906;
wire n_416;
wire n_969;
wire n_283;
wire n_1109;
wire n_919;
wire n_525;
wire n_806;
wire n_367;
wire n_1111;
wire n_970;
wire n_713;
wire n_649;
wire n_598;
wire n_374;
wire n_345;
wire n_318;
wire n_817;
wire n_244;
wire n_643;
wire n_679;
wire n_226;
wire n_924;
wire n_927;
wire n_781;
wire n_261;
wire n_1095;
wire n_682;
wire n_663;
wire n_370;
wire n_706;
wire n_717;
wire n_819;
wire n_286;
wire n_443;
wire n_586;
wire n_864;
wire n_952;
wire n_1096;
wire n_686;
wire n_605;
wire n_776;
wire n_424;
wire n_584;
wire n_528;
wire n_387;
wire n_406;
wire n_826;
wire n_1130;
wire n_524;
wire n_634;
wire n_391;
wire n_349;
wire n_466;
wire n_756;
wire n_940;
wire n_346;
wire n_1016;
wire n_764;
wire n_979;
wire n_348;
wire n_552;
wire n_1077;
wire n_462;
wire n_607;
wire n_670;
wire n_897;
wire n_956;
wire n_949;
wire n_410;
wire n_445;
wire n_379;
wire n_515;
wire n_807;
wire n_765;
wire n_1131;
wire n_264;
wire n_891;
wire n_737;
wire n_885;
wire n_232;
wire n_441;
wire n_568;
wire n_1032;
wire n_385;
wire n_637;
wire n_917;
wire n_327;
wire n_1088;
wire n_766;
wire n_372;
wire n_377;
wire n_396;
wire n_802;
wire n_631;
wire n_399;
wire n_554;
wire n_960;
wire n_520;
wire n_980;
wire n_870;
wire n_714;
wire n_279;
wire n_945;
wire n_702;
wire n_958;
wire n_905;
wire n_790;
wire n_857;
wire n_898;
wire n_363;
wire n_720;
wire n_1067;
wire n_968;
wire n_354;
wire n_813;
wire n_926;
wire n_725;
wire n_419;
wire n_1009;
wire n_230;
wire n_270;
wire n_1064;
wire n_633;
wire n_900;
wire n_1133;
wire n_883;
wire n_338;
wire n_995;
wire n_285;
wire n_1093;
wire n_473;
wire n_801;
wire n_733;
wire n_761;
wire n_818;
wire n_500;
wire n_665;
wire n_731;
wire n_336;
wire n_754;
wire n_779;
wire n_903;
wire n_315;
wire n_871;
wire n_1073;
wire n_594;
wire n_311;
wire n_239;
wire n_402;
wire n_1052;
wire n_1068;
wire n_272;
wire n_829;
wire n_1062;
wire n_668;
wire n_339;
wire n_738;
wire n_758;
wire n_833;
wire n_672;
wire n_487;
wire n_740;
wire n_879;
wire n_1117;
wire n_422;
wire n_1106;
wire n_648;
wire n_784;
wire n_269;
wire n_597;
wire n_816;
wire n_1018;
wire n_855;
wire n_1047;
wire n_259;
wire n_835;
wire n_808;
wire n_953;
wire n_446;
wire n_553;
wire n_1076;
wire n_753;
wire n_1050;
wire n_566;
wire n_814;
wire n_578;
wire n_701;
wire n_1003;
wire n_1125;
wire n_625;
wire n_405;
wire n_557;
wire n_1107;
wire n_858;
wire n_242;
wire n_645;
wire n_989;
wire n_309;
wire n_320;
wire n_331;
wire n_559;
wire n_1134;
wire n_485;
wire n_401;
wire n_267;
wire n_495;
wire n_504;
wire n_647;
wire n_483;
wire n_335;
wire n_435;
wire n_1035;
wire n_350;
wire n_291;
wire n_822;
wire n_381;
wire n_344;
wire n_795;
wire n_426;
wire n_433;
wire n_481;
wire n_600;
wire n_721;
wire n_840;
wire n_1053;
wire n_1084;
wire n_398;
wire n_1090;
wire n_529;
wire n_502;
wire n_253;
wire n_561;
wire n_770;
wire n_839;
wire n_821;
wire n_928;
wire n_1099;
wire n_271;
wire n_507;
wire n_486;
wire n_465;
wire n_901;
wire n_759;
wire n_247;
wire n_569;
wire n_567;
wire n_825;
wire n_732;
wire n_1103;
wire n_971;
wire n_240;
wire n_369;
wire n_224;
wire n_787;
wire n_894;
wire n_1105;
wire n_547;
wire n_420;
wire n_562;
wire n_518;
wire n_439;
wire n_604;
wire n_614;
wire n_677;
wire n_222;
wire n_478;
wire n_703;
wire n_748;
wire n_786;
wire n_510;
wire n_1061;
wire n_1045;
wire n_831;
wire n_256;
wire n_868;
wire n_326;
wire n_681;
wire n_778;
wire n_227;
wire n_874;
wire n_323;
wire n_550;
wire n_1023;
wire n_988;
wire n_635;
wire n_707;
wire n_997;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_694;
wire n_884;
wire n_1116;
wire n_983;
wire n_282;
wire n_328;
wire n_368;
wire n_1113;
wire n_1034;
wire n_590;
wire n_727;
wire n_699;
wire n_277;
wire n_248;
wire n_301;
wire n_467;
wire n_1085;
wire n_432;
wire n_545;
wire n_1015;
wire n_536;
wire n_644;
wire n_293;
wire n_823;
wire n_921;
wire n_620;
wire n_228;
wire n_325;
wire n_276;
wire n_688;
wire n_1074;
wire n_859;
wire n_636;
wire n_427;
wire n_587;
wire n_497;
wire n_1098;
wire n_693;
wire n_863;
wire n_303;
wire n_671;
wire n_442;
wire n_777;
wire n_929;
wire n_352;
wire n_538;
wire n_899;
wire n_920;
wire n_576;
wire n_843;
wire n_1080;
wire n_511;
wire n_1086;
wire n_611;
wire n_1092;
wire n_238;
wire n_365;
wire n_429;
wire n_455;
wire n_654;
wire n_588;
wire n_1013;
wire n_986;
wire n_1104;
wire n_638;
wire n_334;
wire n_1128;
wire n_729;
wire n_887;
wire n_661;
wire n_488;
wire n_1048;
wire n_775;
wire n_667;
wire n_1122;
wire n_1049;
wire n_300;
wire n_533;
wire n_904;
wire n_505;
wire n_869;
wire n_846;
wire n_1132;
wire n_390;
wire n_498;
wire n_501;
wire n_438;
wire n_1059;
wire n_314;
wire n_684;
wire n_1120;
wire n_440;
wire n_627;
wire n_1039;
wire n_273;
wire n_305;
wire n_539;
wire n_312;
wire n_233;
wire n_728;
wire n_388;
wire n_333;
wire n_612;
wire n_449;
wire n_413;
wire n_392;
wire n_376;
wire n_977;
wire n_957;
wire n_512;
wire n_715;
wire n_889;
wire n_1066;
wire n_935;
wire n_579;
wire n_844;
wire n_1012;
wire n_459;
wire n_685;
wire n_321;
wire n_911;
wire n_1136;
wire n_361;
wire n_458;
wire n_383;
wire n_623;
wire n_838;
wire n_237;
wire n_780;
wire n_861;
wire n_950;
wire n_1017;
wire n_711;
wire n_877;
wire n_1021;
wire n_1065;
wire n_453;
wire n_1119;
wire n_734;
wire n_491;
wire n_810;
wire n_723;
wire n_617;
wire n_616;
wire n_658;
wire n_630;
wire n_705;
wire n_570;
wire n_1055;
wire n_260;
wire n_362;
wire n_543;
wire n_942;
wire n_310;
wire n_709;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_1089;
wire n_281;
wire n_628;
wire n_809;
wire n_461;
wire n_1121;
wire n_490;
wire n_262;
wire n_743;
wire n_225;
wire n_907;
wire n_235;
wire n_1006;
wire n_881;
wire n_660;
wire n_464;
wire n_735;
wire n_575;
wire n_546;
wire n_1019;
wire n_297;
wire n_962;
wire n_662;
wire n_641;
wire n_1005;
wire n_503;
wire n_941;
wire n_1112;
wire n_700;
wire n_910;
wire n_290;
wire n_527;
wire n_741;
wire n_772;
wire n_747;
wire n_847;
wire n_939;
wire n_371;
wire n_845;
wire n_888;
wire n_1135;
wire n_918;
wire n_639;
wire n_452;
wire n_673;
wire n_1114;
wire n_676;
wire n_551;
wire n_308;
wire n_708;
wire n_417;
wire n_1038;
wire n_572;
wire n_343;
wire n_865;
wire n_1041;
wire n_414;
wire n_571;
wire n_680;
wire n_287;
wire n_302;
wire n_993;
wire n_380;
wire n_948;
wire n_582;
wire n_284;
wire n_922;
wire n_1004;
wire n_448;
wire n_593;
wire n_755;
wire n_1097;
wire n_710;
wire n_860;
wire n_249;
wire n_534;
wire n_1108;
wire n_355;
wire n_444;
wire n_609;
wire n_278;
wire n_851;
wire n_1043;
wire n_255;
wire n_560;
wire n_450;
wire n_890;
wire n_257;
wire n_842;
wire n_652;
wire n_451;
wire n_613;
wire n_745;
wire n_475;
wire n_1022;
wire n_1033;
wire n_896;
wire n_409;
wire n_947;
wire n_930;
wire n_519;
wire n_902;
wire n_384;
wire n_1031;
wire n_468;
wire n_1056;
wire n_853;
wire n_526;
wire n_716;
wire n_742;
wire n_696;
wire n_1040;
wire n_674;
wire n_1081;
wire n_482;
wire n_316;
wire n_798;
wire n_769;
wire n_820;
wire n_577;
wire n_407;
wire n_774;
wire n_872;
wire n_933;
wire n_916;
wire n_254;
wire n_596;
wire n_954;
wire n_912;
wire n_476;
wire n_460;
wire n_832;
wire n_535;
wire n_231;
wire n_366;
wire n_744;
wire n_762;
wire n_656;
wire n_555;
wire n_234;
wire n_492;
wire n_574;
wire n_848;
wire n_804;
wire n_280;
wire n_982;
wire n_915;
wire n_252;
wire n_664;
wire n_629;
wire n_1075;
wire n_454;
wire n_992;
wire n_966;
wire n_298;
wire n_955;
wire n_532;
wire n_415;
wire n_794;
wire n_763;
wire n_655;
wire n_544;
wire n_540;
wire n_692;
wire n_599;
wire n_768;
wire n_1091;
wire n_514;
wire n_418;
wire n_984;
wire n_537;
wire n_1063;
wire n_223;
wire n_403;
wire n_750;
wire n_834;
wire n_991;
wire n_389;
wire n_1007;
wire n_800;
wire n_657;
wire n_513;
wire n_837;
wire n_288;
wire n_812;
wire n_1126;
wire n_395;
wire n_621;
wire n_606;
wire n_1026;
wire n_951;
wire n_938;
wire n_862;
wire n_304;
wire n_895;
wire n_659;
wire n_583;
wire n_509;
wire n_1014;
wire n_724;
wire n_306;
wire n_666;
wire n_1000;
wire n_313;
wire n_430;
wire n_626;
wire n_493;
wire n_722;
wire n_378;
wire n_436;
wire n_946;
wire n_757;
wire n_375;
wire n_324;
wire n_1030;
wire n_1100;
wire n_585;
wire n_875;
wire n_669;
wire n_785;
wire n_827;
wire n_931;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_622;
wire n_697;
wire n_967;
wire n_999;
wire n_998;
wire n_1083;
wire n_472;
wire n_937;
wire n_296;
wire n_265;
wire n_746;
wire n_456;
wire n_292;
wire n_880;
wire n_793;
wire n_852;
wire n_1079;
wire n_275;
wire n_704;
wire n_1060;
wire n_1044;
wire n_751;
wire n_615;
wire n_1027;
wire n_1070;
wire n_996;
wire n_521;
wire n_963;
wire n_873;
wire n_1082;
wire n_496;
wire n_739;
wire n_1028;
wire n_342;
wire n_866;
wire n_246;
wire n_517;
wire n_925;
wire n_530;
wire n_1094;
wire n_792;
wire n_1001;
wire n_1115;
wire n_824;
wire n_428;
wire n_1002;
wire n_358;
wire n_580;
wire n_892;
wire n_608;
wire n_959;
wire n_494;
wire n_1051;
wire n_719;
wire n_263;
wire n_434;
wire n_360;
wire n_1102;
wire n_975;
wire n_1101;
wire n_1129;
wire n_563;
wire n_229;
wire n_394;
wire n_923;
wire n_1124;
wire n_250;
wire n_932;
wire n_773;
wire n_1037;
wire n_981;
wire n_1010;
wire n_882;
wire n_990;
wire n_1110;
wire n_317;
wire n_867;
wire n_243;
wire n_803;
wire n_329;
wire n_718;
wire n_340;
wire n_944;
wire n_749;
wire n_994;
wire n_289;
wire n_548;
wire n_542;
wire n_815;
wire n_973;
wire n_523;
wire n_1078;
wire n_268;
wire n_972;
wire n_266;
wire n_470;
wire n_457;
wire n_1087;
wire n_632;
wire n_477;
wire n_364;
wire n_258;
wire n_650;
wire n_782;
wire n_856;
wire n_425;
wire n_431;
wire n_811;
wire n_1054;
wire n_508;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1071;
wire n_411;
wire n_484;
wire n_712;
wire n_849;
wire n_976;
wire n_909;
wire n_353;
wire n_736;
wire n_767;
wire n_1025;
wire n_241;
wire n_357;
wire n_412;
wire n_687;
wire n_447;
wire n_964;
wire n_1057;
wire n_382;
wire n_797;
wire n_489;
wire n_480;
wire n_1011;
wire n_642;
wire n_978;
wire n_408;
wire n_828;
wire n_595;
wire n_322;
wire n_251;
wire n_974;
wire n_506;
wire n_893;
wire n_602;
wire n_799;
wire n_558;
wire n_592;
wire n_397;
wire n_854;
wire n_841;
wire n_471;
wire n_351;
wire n_886;
wire n_965;
wire n_393;
wire n_1069;
wire n_474;
wire n_653;
wire n_359;
wire n_573;
wire n_796;
wire n_805;
wire n_531;
wire n_934;
wire n_783;
wire n_675;

INVx1_ASAP7_75t_L g222 ( 
.A(n_56),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_45),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_195),
.Y(n_224)
);

INVxp67_ASAP7_75t_L g225 ( 
.A(n_35),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_202),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_132),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_16),
.Y(n_228)
);

BUFx2_ASAP7_75t_L g229 ( 
.A(n_162),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_22),
.Y(n_230)
);

INVx1_ASAP7_75t_SL g231 ( 
.A(n_70),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_168),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_129),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_16),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_159),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_63),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_115),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_185),
.Y(n_238)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_201),
.Y(n_239)
);

BUFx6f_ASAP7_75t_L g240 ( 
.A(n_57),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_172),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_104),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_100),
.Y(n_243)
);

BUFx10_ASAP7_75t_L g244 ( 
.A(n_126),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_33),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_137),
.Y(n_246)
);

INVx1_ASAP7_75t_SL g247 ( 
.A(n_171),
.Y(n_247)
);

BUFx3_ASAP7_75t_L g248 ( 
.A(n_80),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_37),
.Y(n_249)
);

INVx2_ASAP7_75t_SL g250 ( 
.A(n_53),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_204),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_140),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_174),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_31),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_196),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_175),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_143),
.Y(n_257)
);

BUFx6f_ASAP7_75t_L g258 ( 
.A(n_122),
.Y(n_258)
);

BUFx3_ASAP7_75t_L g259 ( 
.A(n_19),
.Y(n_259)
);

CKINVDCx14_ASAP7_75t_R g260 ( 
.A(n_123),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_153),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_189),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_71),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_6),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_149),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_81),
.Y(n_266)
);

INVxp67_ASAP7_75t_L g267 ( 
.A(n_216),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_221),
.Y(n_268)
);

INVxp67_ASAP7_75t_SL g269 ( 
.A(n_15),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_208),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_148),
.Y(n_271)
);

BUFx3_ASAP7_75t_L g272 ( 
.A(n_40),
.Y(n_272)
);

BUFx3_ASAP7_75t_L g273 ( 
.A(n_107),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_178),
.Y(n_274)
);

BUFx10_ASAP7_75t_L g275 ( 
.A(n_2),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_89),
.Y(n_276)
);

BUFx2_ASAP7_75t_L g277 ( 
.A(n_173),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_4),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_69),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_151),
.Y(n_280)
);

INVx2_ASAP7_75t_L g281 ( 
.A(n_29),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_212),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_94),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_19),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_211),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_82),
.Y(n_286)
);

INVx1_ASAP7_75t_SL g287 ( 
.A(n_6),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_43),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_219),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_77),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_229),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_259),
.Y(n_292)
);

INVxp67_ASAP7_75t_SL g293 ( 
.A(n_259),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_230),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_264),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_277),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_244),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g298 ( 
.A(n_275),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_244),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g300 ( 
.A(n_275),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_244),
.Y(n_301)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_248),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_236),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_260),
.Y(n_304)
);

INVx2_ASAP7_75t_L g305 ( 
.A(n_248),
.Y(n_305)
);

INVx2_ASAP7_75t_L g306 ( 
.A(n_272),
.Y(n_306)
);

INVxp33_ASAP7_75t_SL g307 ( 
.A(n_228),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_275),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_260),
.Y(n_309)
);

BUFx2_ASAP7_75t_L g310 ( 
.A(n_234),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_269),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_222),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_253),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_223),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_232),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_265),
.Y(n_316)
);

INVxp67_ASAP7_75t_SL g317 ( 
.A(n_272),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_235),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_237),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_241),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_254),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_255),
.Y(n_322)
);

INVxp67_ASAP7_75t_L g323 ( 
.A(n_278),
.Y(n_323)
);

INVxp67_ASAP7_75t_L g324 ( 
.A(n_284),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_268),
.Y(n_325)
);

INVxp67_ASAP7_75t_SL g326 ( 
.A(n_273),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_262),
.Y(n_327)
);

BUFx2_ASAP7_75t_L g328 ( 
.A(n_287),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_286),
.Y(n_329)
);

BUFx3_ASAP7_75t_L g330 ( 
.A(n_273),
.Y(n_330)
);

INVxp67_ASAP7_75t_SL g331 ( 
.A(n_239),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_270),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_283),
.Y(n_333)
);

INVxp67_ASAP7_75t_L g334 ( 
.A(n_285),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_224),
.Y(n_335)
);

INVx2_ASAP7_75t_L g336 ( 
.A(n_239),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_281),
.Y(n_337)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_226),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_281),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_250),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_317),
.B(n_326),
.Y(n_341)
);

OAI22xp5_ASAP7_75t_SL g342 ( 
.A1(n_298),
.A2(n_231),
.B1(n_247),
.B2(n_225),
.Y(n_342)
);

AND2x4_ASAP7_75t_L g343 ( 
.A(n_330),
.B(n_267),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_294),
.Y(n_344)
);

BUFx8_ASAP7_75t_L g345 ( 
.A(n_328),
.Y(n_345)
);

AND2x2_ASAP7_75t_L g346 ( 
.A(n_293),
.B(n_227),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_297),
.B(n_233),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_299),
.B(n_238),
.Y(n_348)
);

CKINVDCx20_ASAP7_75t_R g349 ( 
.A(n_316),
.Y(n_349)
);

INVx2_ASAP7_75t_L g350 ( 
.A(n_336),
.Y(n_350)
);

HB1xp67_ASAP7_75t_L g351 ( 
.A(n_291),
.Y(n_351)
);

BUFx12f_ASAP7_75t_L g352 ( 
.A(n_304),
.Y(n_352)
);

AND2x4_ASAP7_75t_L g353 ( 
.A(n_330),
.B(n_240),
.Y(n_353)
);

AOI22xp5_ASAP7_75t_L g354 ( 
.A1(n_291),
.A2(n_290),
.B1(n_289),
.B2(n_288),
.Y(n_354)
);

NAND2xp33_ASAP7_75t_L g355 ( 
.A(n_312),
.B(n_240),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_295),
.Y(n_356)
);

BUFx12f_ASAP7_75t_L g357 ( 
.A(n_304),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_292),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_336),
.Y(n_359)
);

INVx3_ASAP7_75t_L g360 ( 
.A(n_302),
.Y(n_360)
);

OAI22xp5_ASAP7_75t_SL g361 ( 
.A1(n_298),
.A2(n_282),
.B1(n_280),
.B2(n_279),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_337),
.Y(n_362)
);

BUFx3_ASAP7_75t_L g363 ( 
.A(n_302),
.Y(n_363)
);

BUFx6f_ASAP7_75t_L g364 ( 
.A(n_305),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_301),
.B(n_242),
.Y(n_365)
);

AND2x4_ASAP7_75t_L g366 ( 
.A(n_334),
.B(n_240),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_309),
.B(n_243),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_339),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_309),
.B(n_245),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_305),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_306),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_306),
.Y(n_372)
);

INVx3_ASAP7_75t_L g373 ( 
.A(n_314),
.Y(n_373)
);

HB1xp67_ASAP7_75t_L g374 ( 
.A(n_310),
.Y(n_374)
);

AOI22x1_ASAP7_75t_SL g375 ( 
.A1(n_316),
.A2(n_276),
.B1(n_274),
.B2(n_271),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_315),
.Y(n_376)
);

OAI22xp5_ASAP7_75t_SL g377 ( 
.A1(n_300),
.A2(n_325),
.B1(n_329),
.B2(n_313),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_SL g378 ( 
.A(n_335),
.B(n_266),
.Y(n_378)
);

INVx2_ASAP7_75t_SL g379 ( 
.A(n_335),
.Y(n_379)
);

HB1xp67_ASAP7_75t_L g380 ( 
.A(n_323),
.Y(n_380)
);

INVx4_ASAP7_75t_L g381 ( 
.A(n_308),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_303),
.Y(n_382)
);

AOI22xp5_ASAP7_75t_L g383 ( 
.A1(n_338),
.A2(n_263),
.B1(n_261),
.B2(n_246),
.Y(n_383)
);

INVx2_ASAP7_75t_L g384 ( 
.A(n_318),
.Y(n_384)
);

OAI21x1_ASAP7_75t_L g385 ( 
.A1(n_319),
.A2(n_258),
.B(n_240),
.Y(n_385)
);

INVxp67_ASAP7_75t_L g386 ( 
.A(n_296),
.Y(n_386)
);

INVx3_ASAP7_75t_L g387 ( 
.A(n_320),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_331),
.B(n_249),
.Y(n_388)
);

INVx3_ASAP7_75t_L g389 ( 
.A(n_321),
.Y(n_389)
);

BUFx6f_ASAP7_75t_L g390 ( 
.A(n_322),
.Y(n_390)
);

AND2x2_ASAP7_75t_L g391 ( 
.A(n_324),
.B(n_251),
.Y(n_391)
);

INVx2_ASAP7_75t_L g392 ( 
.A(n_327),
.Y(n_392)
);

XNOR2x2_ASAP7_75t_R g393 ( 
.A(n_300),
.B(n_0),
.Y(n_393)
);

AND2x4_ASAP7_75t_L g394 ( 
.A(n_340),
.B(n_258),
.Y(n_394)
);

HB1xp67_ASAP7_75t_L g395 ( 
.A(n_338),
.Y(n_395)
);

NOR2xp33_ASAP7_75t_L g396 ( 
.A(n_341),
.B(n_307),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_350),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_350),
.Y(n_398)
);

BUFx6f_ASAP7_75t_L g399 ( 
.A(n_364),
.Y(n_399)
);

INVx2_ASAP7_75t_SL g400 ( 
.A(n_380),
.Y(n_400)
);

INVx2_ASAP7_75t_L g401 ( 
.A(n_364),
.Y(n_401)
);

INVx2_ASAP7_75t_L g402 ( 
.A(n_364),
.Y(n_402)
);

INVx2_ASAP7_75t_L g403 ( 
.A(n_364),
.Y(n_403)
);

INVx2_ASAP7_75t_L g404 ( 
.A(n_359),
.Y(n_404)
);

OR2x2_ASAP7_75t_L g405 ( 
.A(n_351),
.B(n_313),
.Y(n_405)
);

INVx2_ASAP7_75t_L g406 ( 
.A(n_363),
.Y(n_406)
);

INVx2_ASAP7_75t_L g407 ( 
.A(n_385),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_346),
.B(n_332),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_370),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_371),
.Y(n_410)
);

INVx2_ASAP7_75t_L g411 ( 
.A(n_363),
.Y(n_411)
);

INVx2_ASAP7_75t_L g412 ( 
.A(n_372),
.Y(n_412)
);

INVx2_ASAP7_75t_L g413 ( 
.A(n_390),
.Y(n_413)
);

INVx2_ASAP7_75t_L g414 ( 
.A(n_390),
.Y(n_414)
);

INVx2_ASAP7_75t_L g415 ( 
.A(n_390),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_SL g416 ( 
.A(n_354),
.B(n_307),
.Y(n_416)
);

INVx3_ASAP7_75t_L g417 ( 
.A(n_390),
.Y(n_417)
);

INVx2_ASAP7_75t_SL g418 ( 
.A(n_380),
.Y(n_418)
);

INVx2_ASAP7_75t_L g419 ( 
.A(n_360),
.Y(n_419)
);

AND2x2_ASAP7_75t_L g420 ( 
.A(n_373),
.B(n_333),
.Y(n_420)
);

AND2x2_ASAP7_75t_L g421 ( 
.A(n_373),
.B(n_311),
.Y(n_421)
);

INVx2_ASAP7_75t_SL g422 ( 
.A(n_343),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_384),
.Y(n_423)
);

INVx2_ASAP7_75t_L g424 ( 
.A(n_360),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_384),
.Y(n_425)
);

AO21x2_ASAP7_75t_L g426 ( 
.A1(n_378),
.A2(n_348),
.B(n_347),
.Y(n_426)
);

BUFx3_ASAP7_75t_L g427 ( 
.A(n_353),
.Y(n_427)
);

INVx2_ASAP7_75t_L g428 ( 
.A(n_362),
.Y(n_428)
);

INVx2_ASAP7_75t_SL g429 ( 
.A(n_343),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_392),
.Y(n_430)
);

INVx2_ASAP7_75t_L g431 ( 
.A(n_368),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_392),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_376),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_SL g434 ( 
.A(n_379),
.B(n_325),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_388),
.B(n_252),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_387),
.Y(n_436)
);

INVx3_ASAP7_75t_L g437 ( 
.A(n_353),
.Y(n_437)
);

AO21x2_ASAP7_75t_L g438 ( 
.A1(n_378),
.A2(n_257),
.B(n_256),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_387),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_SL g440 ( 
.A(n_383),
.B(n_329),
.Y(n_440)
);

INVx2_ASAP7_75t_L g441 ( 
.A(n_389),
.Y(n_441)
);

NOR2xp33_ASAP7_75t_L g442 ( 
.A(n_381),
.B(n_258),
.Y(n_442)
);

INVx2_ASAP7_75t_L g443 ( 
.A(n_389),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_358),
.Y(n_444)
);

INVx2_ASAP7_75t_L g445 ( 
.A(n_344),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_L g446 ( 
.A(n_353),
.B(n_366),
.Y(n_446)
);

NAND3xp33_ASAP7_75t_L g447 ( 
.A(n_356),
.B(n_258),
.C(n_0),
.Y(n_447)
);

INVx2_ASAP7_75t_L g448 ( 
.A(n_394),
.Y(n_448)
);

AOI21x1_ASAP7_75t_L g449 ( 
.A1(n_394),
.A2(n_220),
.B(n_30),
.Y(n_449)
);

AND2x2_ASAP7_75t_L g450 ( 
.A(n_366),
.B(n_1),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_SL g451 ( 
.A(n_391),
.B(n_1),
.Y(n_451)
);

NOR2x1p5_ASAP7_75t_L g452 ( 
.A(n_352),
.B(n_2),
.Y(n_452)
);

INVx3_ASAP7_75t_L g453 ( 
.A(n_394),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_366),
.B(n_3),
.Y(n_454)
);

INVx2_ASAP7_75t_L g455 ( 
.A(n_381),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_355),
.Y(n_456)
);

INVx2_ASAP7_75t_L g457 ( 
.A(n_343),
.Y(n_457)
);

INVx3_ASAP7_75t_L g458 ( 
.A(n_365),
.Y(n_458)
);

CKINVDCx5p33_ASAP7_75t_R g459 ( 
.A(n_382),
.Y(n_459)
);

INVx2_ASAP7_75t_L g460 ( 
.A(n_386),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_SL g461 ( 
.A(n_367),
.B(n_3),
.Y(n_461)
);

INVx2_ASAP7_75t_SL g462 ( 
.A(n_374),
.Y(n_462)
);

INVx2_ASAP7_75t_L g463 ( 
.A(n_369),
.Y(n_463)
);

INVx2_ASAP7_75t_L g464 ( 
.A(n_374),
.Y(n_464)
);

INVx2_ASAP7_75t_L g465 ( 
.A(n_355),
.Y(n_465)
);

CKINVDCx5p33_ASAP7_75t_R g466 ( 
.A(n_382),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_351),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_342),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_352),
.Y(n_469)
);

AND2x2_ASAP7_75t_L g470 ( 
.A(n_357),
.B(n_4),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_437),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_437),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_437),
.Y(n_473)
);

OR2x6_ASAP7_75t_L g474 ( 
.A(n_469),
.B(n_377),
.Y(n_474)
);

XOR2xp5_ASAP7_75t_L g475 ( 
.A(n_459),
.B(n_349),
.Y(n_475)
);

AND2x4_ASAP7_75t_L g476 ( 
.A(n_422),
.B(n_395),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_437),
.Y(n_477)
);

AND2x4_ASAP7_75t_L g478 ( 
.A(n_422),
.B(n_429),
.Y(n_478)
);

AND2x2_ASAP7_75t_L g479 ( 
.A(n_400),
.B(n_357),
.Y(n_479)
);

NOR2xp33_ASAP7_75t_L g480 ( 
.A(n_463),
.B(n_361),
.Y(n_480)
);

OAI21xp5_ASAP7_75t_L g481 ( 
.A1(n_407),
.A2(n_395),
.B(n_375),
.Y(n_481)
);

AND2x2_ASAP7_75t_L g482 ( 
.A(n_400),
.B(n_349),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_419),
.Y(n_483)
);

NOR2xp33_ASAP7_75t_L g484 ( 
.A(n_463),
.B(n_345),
.Y(n_484)
);

BUFx8_ASAP7_75t_L g485 ( 
.A(n_469),
.Y(n_485)
);

XOR2xp5_ASAP7_75t_L g486 ( 
.A(n_466),
.B(n_345),
.Y(n_486)
);

AND2x2_ASAP7_75t_L g487 ( 
.A(n_418),
.B(n_345),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_424),
.Y(n_488)
);

INVx2_ASAP7_75t_L g489 ( 
.A(n_411),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_424),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_424),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_436),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_L g493 ( 
.A(n_463),
.B(n_5),
.Y(n_493)
);

OAI21xp5_ASAP7_75t_L g494 ( 
.A1(n_407),
.A2(n_5),
.B(n_7),
.Y(n_494)
);

OR2x2_ASAP7_75t_L g495 ( 
.A(n_462),
.B(n_393),
.Y(n_495)
);

NOR2xp33_ASAP7_75t_L g496 ( 
.A(n_396),
.B(n_7),
.Y(n_496)
);

XOR2xp5_ASAP7_75t_L g497 ( 
.A(n_405),
.B(n_28),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_436),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_439),
.Y(n_499)
);

XOR2x2_ASAP7_75t_L g500 ( 
.A(n_468),
.B(n_8),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_439),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_444),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_444),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_433),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_433),
.Y(n_505)
);

NOR2xp33_ASAP7_75t_SL g506 ( 
.A(n_468),
.B(n_8),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_423),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_423),
.Y(n_508)
);

BUFx6f_ASAP7_75t_L g509 ( 
.A(n_399),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_425),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_425),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_430),
.Y(n_512)
);

NOR2xp67_ASAP7_75t_L g513 ( 
.A(n_458),
.B(n_32),
.Y(n_513)
);

INVx2_ASAP7_75t_L g514 ( 
.A(n_411),
.Y(n_514)
);

OAI21xp5_ASAP7_75t_L g515 ( 
.A1(n_407),
.A2(n_9),
.B(n_10),
.Y(n_515)
);

INVxp67_ASAP7_75t_SL g516 ( 
.A(n_427),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_430),
.Y(n_517)
);

AND2x2_ASAP7_75t_L g518 ( 
.A(n_418),
.B(n_9),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_432),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_432),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_397),
.Y(n_521)
);

CKINVDCx20_ASAP7_75t_R g522 ( 
.A(n_462),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_397),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_398),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_398),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_441),
.Y(n_526)
);

CKINVDCx5p33_ASAP7_75t_R g527 ( 
.A(n_405),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_441),
.Y(n_528)
);

CKINVDCx5p33_ASAP7_75t_R g529 ( 
.A(n_464),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_443),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_443),
.Y(n_531)
);

CKINVDCx5p33_ASAP7_75t_R g532 ( 
.A(n_464),
.Y(n_532)
);

INVx2_ASAP7_75t_SL g533 ( 
.A(n_464),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_445),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_445),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_L g536 ( 
.A(n_458),
.B(n_10),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_409),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_409),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_410),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_410),
.Y(n_540)
);

XNOR2xp5_ASAP7_75t_L g541 ( 
.A(n_440),
.B(n_11),
.Y(n_541)
);

NOR2xp33_ASAP7_75t_L g542 ( 
.A(n_458),
.B(n_11),
.Y(n_542)
);

INVx4_ASAP7_75t_SL g543 ( 
.A(n_470),
.Y(n_543)
);

INVx4_ASAP7_75t_L g544 ( 
.A(n_427),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_428),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_L g546 ( 
.A(n_458),
.B(n_12),
.Y(n_546)
);

NOR2xp33_ASAP7_75t_L g547 ( 
.A(n_416),
.B(n_12),
.Y(n_547)
);

AND2x2_ASAP7_75t_L g548 ( 
.A(n_467),
.B(n_13),
.Y(n_548)
);

INVxp33_ASAP7_75t_L g549 ( 
.A(n_467),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_428),
.Y(n_550)
);

AND2x2_ASAP7_75t_L g551 ( 
.A(n_460),
.B(n_13),
.Y(n_551)
);

CKINVDCx16_ASAP7_75t_R g552 ( 
.A(n_470),
.Y(n_552)
);

INVx2_ASAP7_75t_L g553 ( 
.A(n_411),
.Y(n_553)
);

XOR2xp5_ASAP7_75t_L g554 ( 
.A(n_434),
.B(n_34),
.Y(n_554)
);

AND2x6_ASAP7_75t_SL g555 ( 
.A(n_474),
.B(n_454),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_SL g556 ( 
.A(n_480),
.B(n_429),
.Y(n_556)
);

NOR2x1p5_ASAP7_75t_L g557 ( 
.A(n_527),
.B(n_460),
.Y(n_557)
);

NOR2xp33_ASAP7_75t_L g558 ( 
.A(n_484),
.B(n_460),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_545),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_502),
.Y(n_560)
);

AOI22xp5_ASAP7_75t_L g561 ( 
.A1(n_496),
.A2(n_457),
.B1(n_408),
.B2(n_438),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_503),
.Y(n_562)
);

NAND3xp33_ASAP7_75t_L g563 ( 
.A(n_547),
.B(n_451),
.C(n_461),
.Y(n_563)
);

INVx2_ASAP7_75t_L g564 ( 
.A(n_471),
.Y(n_564)
);

OR2x6_ASAP7_75t_L g565 ( 
.A(n_487),
.B(n_457),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_L g566 ( 
.A(n_478),
.B(n_420),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_L g567 ( 
.A(n_478),
.B(n_420),
.Y(n_567)
);

AND2x2_ASAP7_75t_SL g568 ( 
.A(n_506),
.B(n_450),
.Y(n_568)
);

INVx2_ASAP7_75t_L g569 ( 
.A(n_472),
.Y(n_569)
);

BUFx6f_ASAP7_75t_L g570 ( 
.A(n_509),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_L g571 ( 
.A(n_533),
.B(n_421),
.Y(n_571)
);

CKINVDCx5p33_ASAP7_75t_R g572 ( 
.A(n_522),
.Y(n_572)
);

AOI22xp33_ASAP7_75t_L g573 ( 
.A1(n_506),
.A2(n_438),
.B1(n_448),
.B2(n_427),
.Y(n_573)
);

AOI21xp5_ASAP7_75t_L g574 ( 
.A1(n_492),
.A2(n_426),
.B(n_435),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_L g575 ( 
.A(n_529),
.B(n_421),
.Y(n_575)
);

INVx2_ASAP7_75t_SL g576 ( 
.A(n_479),
.Y(n_576)
);

BUFx6f_ASAP7_75t_L g577 ( 
.A(n_509),
.Y(n_577)
);

INVx2_ASAP7_75t_L g578 ( 
.A(n_473),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_SL g579 ( 
.A(n_544),
.B(n_455),
.Y(n_579)
);

NOR2x2_ASAP7_75t_L g580 ( 
.A(n_474),
.B(n_455),
.Y(n_580)
);

INVxp67_ASAP7_75t_SL g581 ( 
.A(n_516),
.Y(n_581)
);

AOI22xp5_ASAP7_75t_L g582 ( 
.A1(n_532),
.A2(n_438),
.B1(n_426),
.B2(n_450),
.Y(n_582)
);

BUFx6f_ASAP7_75t_L g583 ( 
.A(n_509),
.Y(n_583)
);

INVx2_ASAP7_75t_SL g584 ( 
.A(n_482),
.Y(n_584)
);

NAND2xp5_ASAP7_75t_L g585 ( 
.A(n_551),
.B(n_453),
.Y(n_585)
);

INVx2_ASAP7_75t_L g586 ( 
.A(n_477),
.Y(n_586)
);

AOI22xp5_ASAP7_75t_L g587 ( 
.A1(n_542),
.A2(n_426),
.B1(n_453),
.B2(n_446),
.Y(n_587)
);

INVx2_ASAP7_75t_L g588 ( 
.A(n_489),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_SL g589 ( 
.A(n_544),
.B(n_453),
.Y(n_589)
);

AOI22xp5_ASAP7_75t_L g590 ( 
.A1(n_476),
.A2(n_453),
.B1(n_417),
.B2(n_448),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_L g591 ( 
.A(n_504),
.B(n_428),
.Y(n_591)
);

OR2x2_ASAP7_75t_L g592 ( 
.A(n_475),
.B(n_431),
.Y(n_592)
);

BUFx6f_ASAP7_75t_L g593 ( 
.A(n_514),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_L g594 ( 
.A(n_505),
.B(n_431),
.Y(n_594)
);

NOR2xp33_ASAP7_75t_L g595 ( 
.A(n_549),
.B(n_476),
.Y(n_595)
);

INVx8_ASAP7_75t_L g596 ( 
.A(n_474),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_537),
.Y(n_597)
);

INVx3_ASAP7_75t_L g598 ( 
.A(n_553),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_538),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_L g600 ( 
.A(n_518),
.B(n_431),
.Y(n_600)
);

INVxp67_ASAP7_75t_L g601 ( 
.A(n_495),
.Y(n_601)
);

INVx2_ASAP7_75t_SL g602 ( 
.A(n_485),
.Y(n_602)
);

INVxp67_ASAP7_75t_L g603 ( 
.A(n_548),
.Y(n_603)
);

NOR3xp33_ASAP7_75t_L g604 ( 
.A(n_481),
.B(n_447),
.C(n_417),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_L g605 ( 
.A(n_539),
.B(n_406),
.Y(n_605)
);

INVx8_ASAP7_75t_L g606 ( 
.A(n_486),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_SL g607 ( 
.A(n_481),
.B(n_442),
.Y(n_607)
);

NAND2xp33_ASAP7_75t_L g608 ( 
.A(n_536),
.B(n_399),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_L g609 ( 
.A(n_540),
.B(n_406),
.Y(n_609)
);

NOR2xp33_ASAP7_75t_L g610 ( 
.A(n_552),
.B(n_417),
.Y(n_610)
);

NAND2xp33_ASAP7_75t_L g611 ( 
.A(n_536),
.B(n_546),
.Y(n_611)
);

AOI22xp33_ASAP7_75t_SL g612 ( 
.A1(n_485),
.A2(n_447),
.B1(n_452),
.B2(n_456),
.Y(n_612)
);

A2O1A1Ixp33_ASAP7_75t_SL g613 ( 
.A1(n_494),
.A2(n_417),
.B(n_413),
.C(n_414),
.Y(n_613)
);

AND2x6_ASAP7_75t_SL g614 ( 
.A(n_500),
.B(n_493),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_L g615 ( 
.A(n_534),
.B(n_412),
.Y(n_615)
);

AND2x6_ASAP7_75t_SL g616 ( 
.A(n_493),
.B(n_452),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_535),
.Y(n_617)
);

INVx8_ASAP7_75t_L g618 ( 
.A(n_543),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_L g619 ( 
.A(n_498),
.B(n_412),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_499),
.Y(n_620)
);

NOR2xp67_ASAP7_75t_L g621 ( 
.A(n_541),
.B(n_404),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_560),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_562),
.Y(n_623)
);

AND2x4_ASAP7_75t_L g624 ( 
.A(n_557),
.B(n_543),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_L g625 ( 
.A(n_558),
.B(n_550),
.Y(n_625)
);

AOI22xp5_ASAP7_75t_L g626 ( 
.A1(n_568),
.A2(n_497),
.B1(n_554),
.B2(n_513),
.Y(n_626)
);

AND2x2_ASAP7_75t_L g627 ( 
.A(n_595),
.B(n_404),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_L g628 ( 
.A(n_597),
.B(n_507),
.Y(n_628)
);

INVx3_ASAP7_75t_L g629 ( 
.A(n_570),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_SL g630 ( 
.A(n_576),
.B(n_513),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_599),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_620),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_L g633 ( 
.A(n_559),
.B(n_508),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_617),
.Y(n_634)
);

BUFx6f_ASAP7_75t_L g635 ( 
.A(n_618),
.Y(n_635)
);

BUFx2_ASAP7_75t_L g636 ( 
.A(n_572),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_L g637 ( 
.A(n_559),
.B(n_510),
.Y(n_637)
);

INVx3_ASAP7_75t_L g638 ( 
.A(n_570),
.Y(n_638)
);

AND2x2_ASAP7_75t_L g639 ( 
.A(n_575),
.B(n_494),
.Y(n_639)
);

BUFx3_ASAP7_75t_L g640 ( 
.A(n_618),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_619),
.Y(n_641)
);

NAND2xp33_ASAP7_75t_R g642 ( 
.A(n_592),
.B(n_610),
.Y(n_642)
);

BUFx3_ASAP7_75t_L g643 ( 
.A(n_606),
.Y(n_643)
);

A2O1A1Ixp33_ASAP7_75t_L g644 ( 
.A1(n_563),
.A2(n_515),
.B(n_512),
.C(n_511),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_SL g645 ( 
.A(n_584),
.B(n_566),
.Y(n_645)
);

INVx3_ASAP7_75t_L g646 ( 
.A(n_570),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_L g647 ( 
.A(n_567),
.B(n_517),
.Y(n_647)
);

INVx2_ASAP7_75t_L g648 ( 
.A(n_564),
.Y(n_648)
);

NAND2x1p5_ASAP7_75t_L g649 ( 
.A(n_577),
.B(n_519),
.Y(n_649)
);

CKINVDCx5p33_ASAP7_75t_R g650 ( 
.A(n_606),
.Y(n_650)
);

INVx2_ASAP7_75t_L g651 ( 
.A(n_569),
.Y(n_651)
);

NOR3xp33_ASAP7_75t_SL g652 ( 
.A(n_607),
.B(n_515),
.C(n_501),
.Y(n_652)
);

INVx2_ASAP7_75t_L g653 ( 
.A(n_578),
.Y(n_653)
);

INVx2_ASAP7_75t_L g654 ( 
.A(n_586),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_L g655 ( 
.A(n_591),
.B(n_594),
.Y(n_655)
);

HB1xp67_ASAP7_75t_L g656 ( 
.A(n_571),
.Y(n_656)
);

INVx2_ASAP7_75t_L g657 ( 
.A(n_588),
.Y(n_657)
);

NOR2xp33_ASAP7_75t_L g658 ( 
.A(n_601),
.B(n_526),
.Y(n_658)
);

HB1xp67_ASAP7_75t_L g659 ( 
.A(n_581),
.Y(n_659)
);

NOR2xp33_ASAP7_75t_L g660 ( 
.A(n_556),
.B(n_528),
.Y(n_660)
);

NOR2xp33_ASAP7_75t_L g661 ( 
.A(n_565),
.B(n_530),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_605),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_609),
.Y(n_663)
);

INVx2_ASAP7_75t_SL g664 ( 
.A(n_596),
.Y(n_664)
);

OA22x2_ASAP7_75t_L g665 ( 
.A1(n_565),
.A2(n_520),
.B1(n_525),
.B2(n_524),
.Y(n_665)
);

NOR2xp33_ASAP7_75t_L g666 ( 
.A(n_603),
.B(n_531),
.Y(n_666)
);

BUFx6f_ASAP7_75t_L g667 ( 
.A(n_577),
.Y(n_667)
);

BUFx3_ASAP7_75t_L g668 ( 
.A(n_602),
.Y(n_668)
);

BUFx12f_ASAP7_75t_L g669 ( 
.A(n_555),
.Y(n_669)
);

NOR3xp33_ASAP7_75t_SL g670 ( 
.A(n_589),
.B(n_523),
.C(n_521),
.Y(n_670)
);

NOR3xp33_ASAP7_75t_SL g671 ( 
.A(n_600),
.B(n_488),
.C(n_483),
.Y(n_671)
);

BUFx12f_ASAP7_75t_L g672 ( 
.A(n_616),
.Y(n_672)
);

AND2x2_ASAP7_75t_L g673 ( 
.A(n_621),
.B(n_413),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_615),
.Y(n_674)
);

INVx5_ASAP7_75t_L g675 ( 
.A(n_577),
.Y(n_675)
);

BUFx6f_ASAP7_75t_L g676 ( 
.A(n_583),
.Y(n_676)
);

BUFx3_ASAP7_75t_L g677 ( 
.A(n_596),
.Y(n_677)
);

AND2x6_ASAP7_75t_L g678 ( 
.A(n_583),
.B(n_456),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_598),
.Y(n_679)
);

BUFx2_ASAP7_75t_L g680 ( 
.A(n_580),
.Y(n_680)
);

NOR3xp33_ASAP7_75t_SL g681 ( 
.A(n_574),
.B(n_491),
.C(n_490),
.Y(n_681)
);

NAND3xp33_ASAP7_75t_L g682 ( 
.A(n_604),
.B(n_414),
.C(n_413),
.Y(n_682)
);

NOR3xp33_ASAP7_75t_SL g683 ( 
.A(n_579),
.B(n_14),
.C(n_15),
.Y(n_683)
);

AOI21xp5_ASAP7_75t_L g684 ( 
.A1(n_611),
.A2(n_608),
.B(n_613),
.Y(n_684)
);

INVx3_ASAP7_75t_L g685 ( 
.A(n_675),
.Y(n_685)
);

AND2x2_ASAP7_75t_L g686 ( 
.A(n_626),
.B(n_612),
.Y(n_686)
);

AND2x2_ASAP7_75t_L g687 ( 
.A(n_627),
.B(n_573),
.Y(n_687)
);

NAND3xp33_ASAP7_75t_L g688 ( 
.A(n_652),
.B(n_561),
.C(n_582),
.Y(n_688)
);

AOI21xp5_ASAP7_75t_L g689 ( 
.A1(n_655),
.A2(n_585),
.B(n_587),
.Y(n_689)
);

BUFx6f_ASAP7_75t_L g690 ( 
.A(n_635),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_L g691 ( 
.A(n_656),
.B(n_614),
.Y(n_691)
);

AND2x4_ASAP7_75t_L g692 ( 
.A(n_624),
.B(n_590),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_L g693 ( 
.A(n_656),
.B(n_598),
.Y(n_693)
);

AOI21x1_ASAP7_75t_L g694 ( 
.A1(n_684),
.A2(n_449),
.B(n_414),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_SL g695 ( 
.A(n_659),
.B(n_583),
.Y(n_695)
);

OAI21xp5_ASAP7_75t_L g696 ( 
.A1(n_652),
.A2(n_415),
.B(n_402),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_L g697 ( 
.A(n_641),
.B(n_662),
.Y(n_697)
);

NAND3xp33_ASAP7_75t_L g698 ( 
.A(n_683),
.B(n_415),
.C(n_593),
.Y(n_698)
);

OAI21x1_ASAP7_75t_L g699 ( 
.A1(n_684),
.A2(n_449),
.B(n_402),
.Y(n_699)
);

OAI22xp5_ASAP7_75t_L g700 ( 
.A1(n_639),
.A2(n_593),
.B1(n_403),
.B2(n_401),
.Y(n_700)
);

AOI21xp5_ASAP7_75t_L g701 ( 
.A1(n_655),
.A2(n_593),
.B(n_399),
.Y(n_701)
);

OAI21x1_ASAP7_75t_L g702 ( 
.A1(n_665),
.A2(n_682),
.B(n_649),
.Y(n_702)
);

OAI21xp5_ASAP7_75t_L g703 ( 
.A1(n_644),
.A2(n_403),
.B(n_401),
.Y(n_703)
);

AND2x2_ASAP7_75t_L g704 ( 
.A(n_658),
.B(n_465),
.Y(n_704)
);

A2O1A1Ixp33_ASAP7_75t_L g705 ( 
.A1(n_671),
.A2(n_465),
.B(n_399),
.C(n_18),
.Y(n_705)
);

AOI21xp5_ASAP7_75t_L g706 ( 
.A1(n_625),
.A2(n_399),
.B(n_38),
.Y(n_706)
);

AND2x4_ASAP7_75t_L g707 ( 
.A(n_624),
.B(n_399),
.Y(n_707)
);

OAI21x1_ASAP7_75t_L g708 ( 
.A1(n_665),
.A2(n_39),
.B(n_36),
.Y(n_708)
);

AOI21x1_ASAP7_75t_L g709 ( 
.A1(n_625),
.A2(n_42),
.B(n_41),
.Y(n_709)
);

O2A1O1Ixp5_ASAP7_75t_L g710 ( 
.A1(n_630),
.A2(n_14),
.B(n_17),
.C(n_18),
.Y(n_710)
);

AOI21xp5_ASAP7_75t_L g711 ( 
.A1(n_633),
.A2(n_46),
.B(n_44),
.Y(n_711)
);

NOR2xp33_ASAP7_75t_SL g712 ( 
.A(n_669),
.B(n_17),
.Y(n_712)
);

OAI21x1_ASAP7_75t_L g713 ( 
.A1(n_649),
.A2(n_48),
.B(n_47),
.Y(n_713)
);

OAI21x1_ASAP7_75t_L g714 ( 
.A1(n_633),
.A2(n_50),
.B(n_49),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_L g715 ( 
.A(n_663),
.B(n_20),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_L g716 ( 
.A(n_659),
.B(n_20),
.Y(n_716)
);

INVx2_ASAP7_75t_L g717 ( 
.A(n_648),
.Y(n_717)
);

AO31x2_ASAP7_75t_L g718 ( 
.A1(n_637),
.A2(n_127),
.A3(n_217),
.B(n_215),
.Y(n_718)
);

OAI21x1_ASAP7_75t_L g719 ( 
.A1(n_637),
.A2(n_124),
.B(n_214),
.Y(n_719)
);

AOI21xp5_ASAP7_75t_L g720 ( 
.A1(n_628),
.A2(n_647),
.B(n_674),
.Y(n_720)
);

OR2x6_ASAP7_75t_L g721 ( 
.A(n_664),
.B(n_21),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_L g722 ( 
.A(n_628),
.B(n_647),
.Y(n_722)
);

AOI21xp5_ASAP7_75t_L g723 ( 
.A1(n_622),
.A2(n_121),
.B(n_213),
.Y(n_723)
);

O2A1O1Ixp5_ASAP7_75t_L g724 ( 
.A1(n_666),
.A2(n_21),
.B(n_22),
.C(n_23),
.Y(n_724)
);

OAI21x1_ASAP7_75t_L g725 ( 
.A1(n_629),
.A2(n_125),
.B(n_210),
.Y(n_725)
);

INVx2_ASAP7_75t_L g726 ( 
.A(n_651),
.Y(n_726)
);

BUFx3_ASAP7_75t_L g727 ( 
.A(n_643),
.Y(n_727)
);

A2O1A1Ixp33_ASAP7_75t_L g728 ( 
.A1(n_671),
.A2(n_23),
.B(n_24),
.C(n_25),
.Y(n_728)
);

AOI21xp5_ASAP7_75t_L g729 ( 
.A1(n_623),
.A2(n_128),
.B(n_209),
.Y(n_729)
);

BUFx8_ASAP7_75t_L g730 ( 
.A(n_636),
.Y(n_730)
);

A2O1A1Ixp33_ASAP7_75t_L g731 ( 
.A1(n_660),
.A2(n_24),
.B(n_25),
.C(n_26),
.Y(n_731)
);

AOI21xp5_ASAP7_75t_L g732 ( 
.A1(n_631),
.A2(n_130),
.B(n_207),
.Y(n_732)
);

INVxp67_ASAP7_75t_L g733 ( 
.A(n_642),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_634),
.Y(n_734)
);

INVx2_ASAP7_75t_SL g735 ( 
.A(n_635),
.Y(n_735)
);

OAI21x1_ASAP7_75t_L g736 ( 
.A1(n_629),
.A2(n_646),
.B(n_638),
.Y(n_736)
);

INVx4_ASAP7_75t_L g737 ( 
.A(n_675),
.Y(n_737)
);

AOI21xp33_ASAP7_75t_L g738 ( 
.A1(n_673),
.A2(n_26),
.B(n_27),
.Y(n_738)
);

BUFx3_ASAP7_75t_L g739 ( 
.A(n_640),
.Y(n_739)
);

OAI21x1_ASAP7_75t_L g740 ( 
.A1(n_638),
.A2(n_120),
.B(n_51),
.Y(n_740)
);

HB1xp67_ASAP7_75t_L g741 ( 
.A(n_632),
.Y(n_741)
);

CKINVDCx6p67_ASAP7_75t_R g742 ( 
.A(n_672),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_L g743 ( 
.A(n_661),
.B(n_27),
.Y(n_743)
);

AO31x2_ASAP7_75t_L g744 ( 
.A1(n_681),
.A2(n_52),
.A3(n_54),
.B(n_55),
.Y(n_744)
);

INVxp67_ASAP7_75t_SL g745 ( 
.A(n_667),
.Y(n_745)
);

AO31x2_ASAP7_75t_L g746 ( 
.A1(n_689),
.A2(n_657),
.A3(n_654),
.B(n_653),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_SL g747 ( 
.A(n_722),
.B(n_670),
.Y(n_747)
);

AO31x2_ASAP7_75t_L g748 ( 
.A1(n_720),
.A2(n_679),
.A3(n_681),
.B(n_680),
.Y(n_748)
);

AO22x2_ASAP7_75t_L g749 ( 
.A1(n_688),
.A2(n_645),
.B1(n_677),
.B2(n_668),
.Y(n_749)
);

AOI21xp5_ASAP7_75t_L g750 ( 
.A1(n_688),
.A2(n_706),
.B(n_701),
.Y(n_750)
);

OR2x6_ASAP7_75t_L g751 ( 
.A(n_727),
.B(n_635),
.Y(n_751)
);

NOR4xp25_ASAP7_75t_L g752 ( 
.A(n_731),
.B(n_683),
.C(n_646),
.D(n_670),
.Y(n_752)
);

A2O1A1Ixp33_ASAP7_75t_L g753 ( 
.A1(n_686),
.A2(n_675),
.B(n_676),
.C(n_667),
.Y(n_753)
);

AOI22xp5_ASAP7_75t_L g754 ( 
.A1(n_712),
.A2(n_650),
.B1(n_678),
.B2(n_675),
.Y(n_754)
);

AO31x2_ASAP7_75t_L g755 ( 
.A1(n_700),
.A2(n_678),
.A3(n_676),
.B(n_667),
.Y(n_755)
);

NOR2xp33_ASAP7_75t_L g756 ( 
.A(n_691),
.B(n_743),
.Y(n_756)
);

AOI21xp5_ASAP7_75t_L g757 ( 
.A1(n_703),
.A2(n_676),
.B(n_678),
.Y(n_757)
);

A2O1A1Ixp33_ASAP7_75t_L g758 ( 
.A1(n_705),
.A2(n_678),
.B(n_59),
.C(n_60),
.Y(n_758)
);

BUFx2_ASAP7_75t_L g759 ( 
.A(n_730),
.Y(n_759)
);

BUFx6f_ASAP7_75t_L g760 ( 
.A(n_739),
.Y(n_760)
);

AOI21xp5_ASAP7_75t_L g761 ( 
.A1(n_711),
.A2(n_696),
.B(n_697),
.Y(n_761)
);

OAI22xp5_ASAP7_75t_L g762 ( 
.A1(n_728),
.A2(n_678),
.B1(n_61),
.B2(n_62),
.Y(n_762)
);

OA21x2_ASAP7_75t_L g763 ( 
.A1(n_699),
.A2(n_702),
.B(n_694),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_741),
.Y(n_764)
);

AO31x2_ASAP7_75t_L g765 ( 
.A1(n_734),
.A2(n_58),
.A3(n_64),
.B(n_65),
.Y(n_765)
);

AOI21xp5_ASAP7_75t_L g766 ( 
.A1(n_696),
.A2(n_66),
.B(n_67),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_L g767 ( 
.A(n_704),
.B(n_693),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_734),
.Y(n_768)
);

BUFx3_ASAP7_75t_L g769 ( 
.A(n_730),
.Y(n_769)
);

OAI21x1_ASAP7_75t_L g770 ( 
.A1(n_714),
.A2(n_68),
.B(n_72),
.Y(n_770)
);

AO32x2_ASAP7_75t_L g771 ( 
.A1(n_737),
.A2(n_73),
.A3(n_74),
.B1(n_75),
.B2(n_76),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_717),
.Y(n_772)
);

OAI21x1_ASAP7_75t_L g773 ( 
.A1(n_719),
.A2(n_78),
.B(n_79),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_L g774 ( 
.A(n_716),
.B(n_83),
.Y(n_774)
);

O2A1O1Ixp33_ASAP7_75t_SL g775 ( 
.A1(n_715),
.A2(n_84),
.B(n_85),
.C(n_86),
.Y(n_775)
);

AO31x2_ASAP7_75t_L g776 ( 
.A1(n_726),
.A2(n_87),
.A3(n_88),
.B(n_90),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_L g777 ( 
.A(n_733),
.B(n_218),
.Y(n_777)
);

INVx2_ASAP7_75t_L g778 ( 
.A(n_736),
.Y(n_778)
);

AOI21xp5_ASAP7_75t_L g779 ( 
.A1(n_723),
.A2(n_91),
.B(n_92),
.Y(n_779)
);

AOI21xp5_ASAP7_75t_L g780 ( 
.A1(n_729),
.A2(n_93),
.B(n_95),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_695),
.Y(n_781)
);

OR2x2_ASAP7_75t_L g782 ( 
.A(n_687),
.B(n_96),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_745),
.Y(n_783)
);

AOI21xp5_ASAP7_75t_L g784 ( 
.A1(n_732),
.A2(n_206),
.B(n_98),
.Y(n_784)
);

OA21x2_ASAP7_75t_L g785 ( 
.A1(n_708),
.A2(n_97),
.B(n_99),
.Y(n_785)
);

INVxp67_ASAP7_75t_SL g786 ( 
.A(n_685),
.Y(n_786)
);

CKINVDCx8_ASAP7_75t_R g787 ( 
.A(n_690),
.Y(n_787)
);

BUFx3_ASAP7_75t_L g788 ( 
.A(n_690),
.Y(n_788)
);

INVx2_ASAP7_75t_L g789 ( 
.A(n_707),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_L g790 ( 
.A(n_692),
.B(n_205),
.Y(n_790)
);

AOI21xp5_ASAP7_75t_L g791 ( 
.A1(n_698),
.A2(n_101),
.B(n_102),
.Y(n_791)
);

AOI21xp5_ASAP7_75t_L g792 ( 
.A1(n_698),
.A2(n_103),
.B(n_105),
.Y(n_792)
);

A2O1A1Ixp33_ASAP7_75t_L g793 ( 
.A1(n_724),
.A2(n_106),
.B(n_108),
.C(n_109),
.Y(n_793)
);

A2O1A1Ixp33_ASAP7_75t_L g794 ( 
.A1(n_710),
.A2(n_738),
.B(n_692),
.C(n_712),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_718),
.Y(n_795)
);

AOI21x1_ASAP7_75t_L g796 ( 
.A1(n_709),
.A2(n_110),
.B(n_111),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_718),
.Y(n_797)
);

INVx2_ASAP7_75t_L g798 ( 
.A(n_718),
.Y(n_798)
);

NOR2xp33_ASAP7_75t_L g799 ( 
.A(n_721),
.B(n_112),
.Y(n_799)
);

OR2x2_ASAP7_75t_L g800 ( 
.A(n_721),
.B(n_113),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_L g801 ( 
.A(n_690),
.B(n_203),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_L g802 ( 
.A(n_721),
.B(n_735),
.Y(n_802)
);

AOI21xp5_ASAP7_75t_L g803 ( 
.A1(n_713),
.A2(n_114),
.B(n_116),
.Y(n_803)
);

A2O1A1Ixp33_ASAP7_75t_L g804 ( 
.A1(n_725),
.A2(n_117),
.B(n_118),
.C(n_119),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_L g805 ( 
.A(n_685),
.B(n_200),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_L g806 ( 
.A(n_737),
.B(n_131),
.Y(n_806)
);

AND2x6_ASAP7_75t_L g807 ( 
.A(n_744),
.B(n_740),
.Y(n_807)
);

INVx2_ASAP7_75t_SL g808 ( 
.A(n_742),
.Y(n_808)
);

OR2x2_ASAP7_75t_L g809 ( 
.A(n_744),
.B(n_133),
.Y(n_809)
);

AOI22xp33_ASAP7_75t_SL g810 ( 
.A1(n_749),
.A2(n_744),
.B1(n_135),
.B2(n_136),
.Y(n_810)
);

BUFx2_ASAP7_75t_SL g811 ( 
.A(n_760),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_768),
.Y(n_812)
);

INVx2_ASAP7_75t_L g813 ( 
.A(n_772),
.Y(n_813)
);

OAI22xp33_ASAP7_75t_L g814 ( 
.A1(n_754),
.A2(n_134),
.B1(n_138),
.B2(n_139),
.Y(n_814)
);

OAI22xp33_ASAP7_75t_L g815 ( 
.A1(n_800),
.A2(n_141),
.B1(n_142),
.B2(n_144),
.Y(n_815)
);

OAI21xp5_ASAP7_75t_L g816 ( 
.A1(n_747),
.A2(n_761),
.B(n_758),
.Y(n_816)
);

AOI22xp33_ASAP7_75t_L g817 ( 
.A1(n_756),
.A2(n_145),
.B1(n_146),
.B2(n_147),
.Y(n_817)
);

AOI22xp33_ASAP7_75t_SL g818 ( 
.A1(n_749),
.A2(n_150),
.B1(n_152),
.B2(n_154),
.Y(n_818)
);

AND2x2_ASAP7_75t_L g819 ( 
.A(n_764),
.B(n_155),
.Y(n_819)
);

INVx1_ASAP7_75t_SL g820 ( 
.A(n_783),
.Y(n_820)
);

OAI22xp5_ASAP7_75t_L g821 ( 
.A1(n_794),
.A2(n_156),
.B1(n_157),
.B2(n_158),
.Y(n_821)
);

BUFx10_ASAP7_75t_L g822 ( 
.A(n_760),
.Y(n_822)
);

AND2x2_ASAP7_75t_L g823 ( 
.A(n_767),
.B(n_160),
.Y(n_823)
);

AOI22xp5_ASAP7_75t_L g824 ( 
.A1(n_799),
.A2(n_161),
.B1(n_163),
.B2(n_164),
.Y(n_824)
);

INVx5_ASAP7_75t_L g825 ( 
.A(n_807),
.Y(n_825)
);

INVx3_ASAP7_75t_SL g826 ( 
.A(n_751),
.Y(n_826)
);

OAI22xp5_ASAP7_75t_L g827 ( 
.A1(n_762),
.A2(n_165),
.B1(n_166),
.B2(n_167),
.Y(n_827)
);

BUFx6f_ASAP7_75t_SL g828 ( 
.A(n_769),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_L g829 ( 
.A(n_781),
.B(n_169),
.Y(n_829)
);

AND2x2_ASAP7_75t_L g830 ( 
.A(n_786),
.B(n_170),
.Y(n_830)
);

CKINVDCx5p33_ASAP7_75t_R g831 ( 
.A(n_759),
.Y(n_831)
);

OAI22xp5_ASAP7_75t_L g832 ( 
.A1(n_793),
.A2(n_176),
.B1(n_177),
.B2(n_179),
.Y(n_832)
);

INVx1_ASAP7_75t_SL g833 ( 
.A(n_802),
.Y(n_833)
);

INVx6_ASAP7_75t_L g834 ( 
.A(n_751),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_SL g835 ( 
.A(n_753),
.B(n_180),
.Y(n_835)
);

CKINVDCx6p67_ASAP7_75t_R g836 ( 
.A(n_788),
.Y(n_836)
);

AOI22xp33_ASAP7_75t_L g837 ( 
.A1(n_782),
.A2(n_181),
.B1(n_182),
.B2(n_183),
.Y(n_837)
);

OAI22xp5_ASAP7_75t_L g838 ( 
.A1(n_774),
.A2(n_184),
.B1(n_186),
.B2(n_187),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_746),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_746),
.Y(n_840)
);

BUFx6f_ASAP7_75t_L g841 ( 
.A(n_787),
.Y(n_841)
);

CKINVDCx20_ASAP7_75t_R g842 ( 
.A(n_808),
.Y(n_842)
);

AOI22xp33_ASAP7_75t_SL g843 ( 
.A1(n_809),
.A2(n_188),
.B1(n_190),
.B2(n_191),
.Y(n_843)
);

AOI22xp33_ASAP7_75t_L g844 ( 
.A1(n_777),
.A2(n_192),
.B1(n_193),
.B2(n_194),
.Y(n_844)
);

AOI22xp33_ASAP7_75t_L g845 ( 
.A1(n_789),
.A2(n_197),
.B1(n_198),
.B2(n_199),
.Y(n_845)
);

INVx2_ASAP7_75t_L g846 ( 
.A(n_748),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_748),
.Y(n_847)
);

AOI22xp33_ASAP7_75t_L g848 ( 
.A1(n_790),
.A2(n_797),
.B1(n_795),
.B2(n_798),
.Y(n_848)
);

CKINVDCx20_ASAP7_75t_R g849 ( 
.A(n_801),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_778),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_755),
.Y(n_851)
);

AOI22xp33_ASAP7_75t_SL g852 ( 
.A1(n_807),
.A2(n_785),
.B1(n_766),
.B2(n_771),
.Y(n_852)
);

INVx1_ASAP7_75t_L g853 ( 
.A(n_755),
.Y(n_853)
);

INVx3_ASAP7_75t_L g854 ( 
.A(n_763),
.Y(n_854)
);

AOI22xp33_ASAP7_75t_L g855 ( 
.A1(n_807),
.A2(n_750),
.B1(n_757),
.B2(n_779),
.Y(n_855)
);

OAI22xp33_ASAP7_75t_L g856 ( 
.A1(n_806),
.A2(n_792),
.B1(n_791),
.B2(n_780),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_L g857 ( 
.A(n_752),
.B(n_805),
.Y(n_857)
);

BUFx12f_ASAP7_75t_L g858 ( 
.A(n_771),
.Y(n_858)
);

INVx3_ASAP7_75t_L g859 ( 
.A(n_765),
.Y(n_859)
);

INVx6_ASAP7_75t_L g860 ( 
.A(n_775),
.Y(n_860)
);

BUFx2_ASAP7_75t_L g861 ( 
.A(n_765),
.Y(n_861)
);

AOI22xp33_ASAP7_75t_L g862 ( 
.A1(n_784),
.A2(n_803),
.B1(n_773),
.B2(n_770),
.Y(n_862)
);

CKINVDCx11_ASAP7_75t_R g863 ( 
.A(n_776),
.Y(n_863)
);

BUFx3_ASAP7_75t_L g864 ( 
.A(n_776),
.Y(n_864)
);

BUFx8_ASAP7_75t_L g865 ( 
.A(n_804),
.Y(n_865)
);

BUFx12f_ASAP7_75t_L g866 ( 
.A(n_796),
.Y(n_866)
);

BUFx6f_ASAP7_75t_L g867 ( 
.A(n_787),
.Y(n_867)
);

INVx2_ASAP7_75t_L g868 ( 
.A(n_850),
.Y(n_868)
);

INVx3_ASAP7_75t_L g869 ( 
.A(n_854),
.Y(n_869)
);

AND2x4_ASAP7_75t_L g870 ( 
.A(n_825),
.B(n_851),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_812),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_847),
.Y(n_872)
);

INVx2_ASAP7_75t_L g873 ( 
.A(n_854),
.Y(n_873)
);

BUFx6f_ASAP7_75t_L g874 ( 
.A(n_825),
.Y(n_874)
);

AO21x2_ASAP7_75t_L g875 ( 
.A1(n_846),
.A2(n_839),
.B(n_840),
.Y(n_875)
);

INVx2_ASAP7_75t_L g876 ( 
.A(n_813),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_853),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_861),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_820),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_820),
.Y(n_880)
);

INVx2_ASAP7_75t_L g881 ( 
.A(n_859),
.Y(n_881)
);

BUFx3_ASAP7_75t_L g882 ( 
.A(n_825),
.Y(n_882)
);

BUFx6f_ASAP7_75t_L g883 ( 
.A(n_866),
.Y(n_883)
);

INVx2_ASAP7_75t_L g884 ( 
.A(n_859),
.Y(n_884)
);

BUFx3_ASAP7_75t_L g885 ( 
.A(n_841),
.Y(n_885)
);

INVx2_ASAP7_75t_L g886 ( 
.A(n_864),
.Y(n_886)
);

INVx3_ASAP7_75t_L g887 ( 
.A(n_858),
.Y(n_887)
);

AND2x2_ASAP7_75t_L g888 ( 
.A(n_833),
.B(n_816),
.Y(n_888)
);

OA21x2_ASAP7_75t_L g889 ( 
.A1(n_816),
.A2(n_855),
.B(n_848),
.Y(n_889)
);

INVx2_ASAP7_75t_L g890 ( 
.A(n_863),
.Y(n_890)
);

HB1xp67_ASAP7_75t_L g891 ( 
.A(n_833),
.Y(n_891)
);

AOI22xp33_ASAP7_75t_L g892 ( 
.A1(n_857),
.A2(n_865),
.B1(n_818),
.B2(n_810),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_819),
.Y(n_893)
);

INVx1_ASAP7_75t_L g894 ( 
.A(n_829),
.Y(n_894)
);

AND2x2_ASAP7_75t_L g895 ( 
.A(n_852),
.B(n_823),
.Y(n_895)
);

INVx1_ASAP7_75t_SL g896 ( 
.A(n_826),
.Y(n_896)
);

INVx1_ASAP7_75t_L g897 ( 
.A(n_860),
.Y(n_897)
);

INVx2_ASAP7_75t_L g898 ( 
.A(n_860),
.Y(n_898)
);

INVx2_ASAP7_75t_L g899 ( 
.A(n_830),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_L g900 ( 
.A(n_836),
.B(n_867),
.Y(n_900)
);

INVx2_ASAP7_75t_SL g901 ( 
.A(n_822),
.Y(n_901)
);

INVxp67_ASAP7_75t_L g902 ( 
.A(n_811),
.Y(n_902)
);

INVx3_ASAP7_75t_L g903 ( 
.A(n_865),
.Y(n_903)
);

OAI22xp5_ASAP7_75t_L g904 ( 
.A1(n_824),
.A2(n_843),
.B1(n_821),
.B2(n_827),
.Y(n_904)
);

INVx2_ASAP7_75t_L g905 ( 
.A(n_834),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_835),
.Y(n_906)
);

OAI21x1_ASAP7_75t_L g907 ( 
.A1(n_862),
.A2(n_832),
.B(n_838),
.Y(n_907)
);

INVx2_ASAP7_75t_L g908 ( 
.A(n_834),
.Y(n_908)
);

AND2x2_ASAP7_75t_L g909 ( 
.A(n_822),
.B(n_824),
.Y(n_909)
);

BUFx3_ASAP7_75t_L g910 ( 
.A(n_841),
.Y(n_910)
);

OAI21x1_ASAP7_75t_L g911 ( 
.A1(n_838),
.A2(n_845),
.B(n_844),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_841),
.Y(n_912)
);

OR2x2_ASAP7_75t_L g913 ( 
.A(n_867),
.B(n_831),
.Y(n_913)
);

NAND2x1p5_ASAP7_75t_L g914 ( 
.A(n_903),
.B(n_867),
.Y(n_914)
);

BUFx3_ASAP7_75t_L g915 ( 
.A(n_885),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_871),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_871),
.Y(n_917)
);

INVx2_ASAP7_75t_L g918 ( 
.A(n_877),
.Y(n_918)
);

AND2x2_ASAP7_75t_L g919 ( 
.A(n_888),
.B(n_899),
.Y(n_919)
);

INVx1_ASAP7_75t_L g920 ( 
.A(n_879),
.Y(n_920)
);

HB1xp67_ASAP7_75t_L g921 ( 
.A(n_879),
.Y(n_921)
);

AND2x2_ASAP7_75t_L g922 ( 
.A(n_888),
.B(n_849),
.Y(n_922)
);

INVx2_ASAP7_75t_L g923 ( 
.A(n_877),
.Y(n_923)
);

CKINVDCx20_ASAP7_75t_R g924 ( 
.A(n_896),
.Y(n_924)
);

INVx2_ASAP7_75t_L g925 ( 
.A(n_872),
.Y(n_925)
);

INVx1_ASAP7_75t_L g926 ( 
.A(n_880),
.Y(n_926)
);

INVxp67_ASAP7_75t_L g927 ( 
.A(n_891),
.Y(n_927)
);

AND2x2_ASAP7_75t_L g928 ( 
.A(n_899),
.B(n_842),
.Y(n_928)
);

BUFx2_ASAP7_75t_L g929 ( 
.A(n_869),
.Y(n_929)
);

INVx1_ASAP7_75t_L g930 ( 
.A(n_880),
.Y(n_930)
);

OA21x2_ASAP7_75t_L g931 ( 
.A1(n_881),
.A2(n_817),
.B(n_837),
.Y(n_931)
);

BUFx2_ASAP7_75t_L g932 ( 
.A(n_869),
.Y(n_932)
);

NOR2xp33_ASAP7_75t_L g933 ( 
.A(n_896),
.B(n_828),
.Y(n_933)
);

INVx1_ASAP7_75t_L g934 ( 
.A(n_872),
.Y(n_934)
);

AOI21xp5_ASAP7_75t_L g935 ( 
.A1(n_904),
.A2(n_856),
.B(n_814),
.Y(n_935)
);

NOR2xp33_ASAP7_75t_L g936 ( 
.A(n_913),
.B(n_828),
.Y(n_936)
);

OR2x2_ASAP7_75t_L g937 ( 
.A(n_878),
.B(n_876),
.Y(n_937)
);

INVx1_ASAP7_75t_L g938 ( 
.A(n_868),
.Y(n_938)
);

AO21x2_ASAP7_75t_L g939 ( 
.A1(n_875),
.A2(n_815),
.B(n_886),
.Y(n_939)
);

INVx3_ASAP7_75t_L g940 ( 
.A(n_869),
.Y(n_940)
);

OA21x2_ASAP7_75t_L g941 ( 
.A1(n_881),
.A2(n_884),
.B(n_907),
.Y(n_941)
);

INVx1_ASAP7_75t_L g942 ( 
.A(n_868),
.Y(n_942)
);

BUFx2_ASAP7_75t_L g943 ( 
.A(n_869),
.Y(n_943)
);

HB1xp67_ASAP7_75t_L g944 ( 
.A(n_894),
.Y(n_944)
);

AND2x4_ASAP7_75t_L g945 ( 
.A(n_882),
.B(n_874),
.Y(n_945)
);

INVx1_ASAP7_75t_L g946 ( 
.A(n_868),
.Y(n_946)
);

INVx2_ASAP7_75t_L g947 ( 
.A(n_937),
.Y(n_947)
);

INVx3_ASAP7_75t_L g948 ( 
.A(n_940),
.Y(n_948)
);

AND2x2_ASAP7_75t_L g949 ( 
.A(n_919),
.B(n_873),
.Y(n_949)
);

INVx1_ASAP7_75t_L g950 ( 
.A(n_918),
.Y(n_950)
);

AND2x2_ASAP7_75t_L g951 ( 
.A(n_919),
.B(n_873),
.Y(n_951)
);

AND2x2_ASAP7_75t_L g952 ( 
.A(n_922),
.B(n_873),
.Y(n_952)
);

AND2x2_ASAP7_75t_L g953 ( 
.A(n_922),
.B(n_887),
.Y(n_953)
);

HB1xp67_ASAP7_75t_L g954 ( 
.A(n_921),
.Y(n_954)
);

NAND2xp5_ASAP7_75t_L g955 ( 
.A(n_944),
.B(n_894),
.Y(n_955)
);

HB1xp67_ASAP7_75t_L g956 ( 
.A(n_927),
.Y(n_956)
);

INVx2_ASAP7_75t_SL g957 ( 
.A(n_915),
.Y(n_957)
);

OAI22xp5_ASAP7_75t_L g958 ( 
.A1(n_935),
.A2(n_892),
.B1(n_904),
.B2(n_903),
.Y(n_958)
);

BUFx3_ASAP7_75t_L g959 ( 
.A(n_924),
.Y(n_959)
);

AND2x2_ASAP7_75t_L g960 ( 
.A(n_928),
.B(n_887),
.Y(n_960)
);

INVx1_ASAP7_75t_L g961 ( 
.A(n_918),
.Y(n_961)
);

AND2x4_ASAP7_75t_L g962 ( 
.A(n_945),
.B(n_882),
.Y(n_962)
);

INVx1_ASAP7_75t_L g963 ( 
.A(n_923),
.Y(n_963)
);

INVx2_ASAP7_75t_L g964 ( 
.A(n_937),
.Y(n_964)
);

AND2x4_ASAP7_75t_L g965 ( 
.A(n_945),
.B(n_882),
.Y(n_965)
);

INVx1_ASAP7_75t_L g966 ( 
.A(n_923),
.Y(n_966)
);

AND2x2_ASAP7_75t_L g967 ( 
.A(n_928),
.B(n_887),
.Y(n_967)
);

INVx1_ASAP7_75t_L g968 ( 
.A(n_925),
.Y(n_968)
);

HB1xp67_ASAP7_75t_L g969 ( 
.A(n_954),
.Y(n_969)
);

INVxp67_ASAP7_75t_SL g970 ( 
.A(n_955),
.Y(n_970)
);

BUFx2_ASAP7_75t_L g971 ( 
.A(n_959),
.Y(n_971)
);

INVx1_ASAP7_75t_L g972 ( 
.A(n_956),
.Y(n_972)
);

INVx1_ASAP7_75t_SL g973 ( 
.A(n_959),
.Y(n_973)
);

INVx1_ASAP7_75t_L g974 ( 
.A(n_950),
.Y(n_974)
);

INVx2_ASAP7_75t_L g975 ( 
.A(n_950),
.Y(n_975)
);

AND2x2_ASAP7_75t_L g976 ( 
.A(n_953),
.B(n_915),
.Y(n_976)
);

NAND3xp33_ASAP7_75t_L g977 ( 
.A(n_958),
.B(n_926),
.C(n_920),
.Y(n_977)
);

INVx2_ASAP7_75t_L g978 ( 
.A(n_961),
.Y(n_978)
);

BUFx3_ASAP7_75t_L g979 ( 
.A(n_959),
.Y(n_979)
);

AND2x2_ASAP7_75t_L g980 ( 
.A(n_953),
.B(n_932),
.Y(n_980)
);

INVxp67_ASAP7_75t_L g981 ( 
.A(n_960),
.Y(n_981)
);

BUFx2_ASAP7_75t_L g982 ( 
.A(n_962),
.Y(n_982)
);

INVx2_ASAP7_75t_L g983 ( 
.A(n_961),
.Y(n_983)
);

OR2x2_ASAP7_75t_L g984 ( 
.A(n_972),
.B(n_947),
.Y(n_984)
);

NAND2xp5_ASAP7_75t_L g985 ( 
.A(n_970),
.B(n_920),
.Y(n_985)
);

INVx1_ASAP7_75t_L g986 ( 
.A(n_969),
.Y(n_986)
);

NOR2x1p5_ASAP7_75t_L g987 ( 
.A(n_979),
.B(n_903),
.Y(n_987)
);

NAND2xp5_ASAP7_75t_L g988 ( 
.A(n_974),
.B(n_926),
.Y(n_988)
);

INVx2_ASAP7_75t_L g989 ( 
.A(n_975),
.Y(n_989)
);

AND2x2_ASAP7_75t_L g990 ( 
.A(n_971),
.B(n_960),
.Y(n_990)
);

INVx1_ASAP7_75t_L g991 ( 
.A(n_971),
.Y(n_991)
);

INVx2_ASAP7_75t_L g992 ( 
.A(n_975),
.Y(n_992)
);

AND2x4_ASAP7_75t_L g993 ( 
.A(n_979),
.B(n_982),
.Y(n_993)
);

AND2x2_ASAP7_75t_L g994 ( 
.A(n_976),
.B(n_982),
.Y(n_994)
);

AND2x2_ASAP7_75t_L g995 ( 
.A(n_976),
.B(n_967),
.Y(n_995)
);

INVx1_ASAP7_75t_L g996 ( 
.A(n_986),
.Y(n_996)
);

INVx1_ASAP7_75t_L g997 ( 
.A(n_991),
.Y(n_997)
);

BUFx3_ASAP7_75t_L g998 ( 
.A(n_993),
.Y(n_998)
);

NAND3xp33_ASAP7_75t_L g999 ( 
.A(n_993),
.B(n_977),
.C(n_985),
.Y(n_999)
);

INVx1_ASAP7_75t_L g1000 ( 
.A(n_984),
.Y(n_1000)
);

BUFx2_ASAP7_75t_L g1001 ( 
.A(n_990),
.Y(n_1001)
);

AND2x2_ASAP7_75t_L g1002 ( 
.A(n_994),
.B(n_981),
.Y(n_1002)
);

INVxp67_ASAP7_75t_SL g1003 ( 
.A(n_985),
.Y(n_1003)
);

OR2x2_ASAP7_75t_L g1004 ( 
.A(n_988),
.B(n_973),
.Y(n_1004)
);

AO221x1_ASAP7_75t_L g1005 ( 
.A1(n_1001),
.A2(n_903),
.B1(n_948),
.B2(n_887),
.C(n_987),
.Y(n_1005)
);

OAI221xp5_ASAP7_75t_L g1006 ( 
.A1(n_1003),
.A2(n_999),
.B1(n_1000),
.B2(n_1004),
.C(n_998),
.Y(n_1006)
);

CKINVDCx20_ASAP7_75t_R g1007 ( 
.A(n_998),
.Y(n_1007)
);

OAI221xp5_ASAP7_75t_L g1008 ( 
.A1(n_1003),
.A2(n_992),
.B1(n_989),
.B2(n_895),
.C(n_890),
.Y(n_1008)
);

NAND2xp5_ASAP7_75t_L g1009 ( 
.A(n_1002),
.B(n_995),
.Y(n_1009)
);

NAND2xp5_ASAP7_75t_L g1010 ( 
.A(n_1002),
.B(n_988),
.Y(n_1010)
);

INVx2_ASAP7_75t_SL g1011 ( 
.A(n_996),
.Y(n_1011)
);

AND2x2_ASAP7_75t_L g1012 ( 
.A(n_1007),
.B(n_997),
.Y(n_1012)
);

INVx2_ASAP7_75t_L g1013 ( 
.A(n_1009),
.Y(n_1013)
);

INVx1_ASAP7_75t_L g1014 ( 
.A(n_1010),
.Y(n_1014)
);

HB1xp67_ASAP7_75t_L g1015 ( 
.A(n_1006),
.Y(n_1015)
);

INVx1_ASAP7_75t_L g1016 ( 
.A(n_1011),
.Y(n_1016)
);

INVx1_ASAP7_75t_L g1017 ( 
.A(n_1008),
.Y(n_1017)
);

OR2x2_ASAP7_75t_L g1018 ( 
.A(n_1005),
.B(n_989),
.Y(n_1018)
);

INVx1_ASAP7_75t_L g1019 ( 
.A(n_1010),
.Y(n_1019)
);

AND2x2_ASAP7_75t_L g1020 ( 
.A(n_1007),
.B(n_980),
.Y(n_1020)
);

INVx1_ASAP7_75t_L g1021 ( 
.A(n_1010),
.Y(n_1021)
);

NAND2xp33_ASAP7_75t_SL g1022 ( 
.A(n_1020),
.B(n_980),
.Y(n_1022)
);

INVx1_ASAP7_75t_L g1023 ( 
.A(n_1013),
.Y(n_1023)
);

INVx2_ASAP7_75t_L g1024 ( 
.A(n_1012),
.Y(n_1024)
);

INVx2_ASAP7_75t_L g1025 ( 
.A(n_1018),
.Y(n_1025)
);

INVx1_ASAP7_75t_L g1026 ( 
.A(n_1013),
.Y(n_1026)
);

NOR2xp67_ASAP7_75t_L g1027 ( 
.A(n_1016),
.B(n_933),
.Y(n_1027)
);

INVxp67_ASAP7_75t_SL g1028 ( 
.A(n_1015),
.Y(n_1028)
);

AOI22xp5_ASAP7_75t_L g1029 ( 
.A1(n_1015),
.A2(n_895),
.B1(n_992),
.B2(n_890),
.Y(n_1029)
);

AOI21xp5_ASAP7_75t_L g1030 ( 
.A1(n_1014),
.A2(n_936),
.B(n_900),
.Y(n_1030)
);

NOR3xp33_ASAP7_75t_SL g1031 ( 
.A(n_1028),
.B(n_1021),
.C(n_1019),
.Y(n_1031)
);

AND2x2_ASAP7_75t_L g1032 ( 
.A(n_1024),
.B(n_1017),
.Y(n_1032)
);

OAI21xp5_ASAP7_75t_L g1033 ( 
.A1(n_1027),
.A2(n_907),
.B(n_911),
.Y(n_1033)
);

INVx1_ASAP7_75t_L g1034 ( 
.A(n_1023),
.Y(n_1034)
);

AND2x2_ASAP7_75t_L g1035 ( 
.A(n_1025),
.B(n_967),
.Y(n_1035)
);

AOI21xp5_ASAP7_75t_L g1036 ( 
.A1(n_1022),
.A2(n_913),
.B(n_978),
.Y(n_1036)
);

NAND2xp5_ASAP7_75t_L g1037 ( 
.A(n_1026),
.B(n_952),
.Y(n_1037)
);

NAND2xp5_ASAP7_75t_L g1038 ( 
.A(n_1029),
.B(n_952),
.Y(n_1038)
);

AOI221xp5_ASAP7_75t_L g1039 ( 
.A1(n_1030),
.A2(n_890),
.B1(n_906),
.B2(n_983),
.C(n_978),
.Y(n_1039)
);

OAI222xp33_ASAP7_75t_L g1040 ( 
.A1(n_1035),
.A2(n_1030),
.B1(n_902),
.B2(n_909),
.C1(n_897),
.C2(n_906),
.Y(n_1040)
);

OAI21xp5_ASAP7_75t_L g1041 ( 
.A1(n_1031),
.A2(n_911),
.B(n_909),
.Y(n_1041)
);

NAND2xp5_ASAP7_75t_L g1042 ( 
.A(n_1032),
.B(n_1034),
.Y(n_1042)
);

INVx1_ASAP7_75t_L g1043 ( 
.A(n_1037),
.Y(n_1043)
);

INVx1_ASAP7_75t_L g1044 ( 
.A(n_1038),
.Y(n_1044)
);

AOI21xp5_ASAP7_75t_L g1045 ( 
.A1(n_1033),
.A2(n_901),
.B(n_957),
.Y(n_1045)
);

INVx2_ASAP7_75t_L g1046 ( 
.A(n_1039),
.Y(n_1046)
);

INVx2_ASAP7_75t_L g1047 ( 
.A(n_1042),
.Y(n_1047)
);

INVx2_ASAP7_75t_L g1048 ( 
.A(n_1043),
.Y(n_1048)
);

HB1xp67_ASAP7_75t_L g1049 ( 
.A(n_1044),
.Y(n_1049)
);

INVx1_ASAP7_75t_L g1050 ( 
.A(n_1046),
.Y(n_1050)
);

INVx1_ASAP7_75t_L g1051 ( 
.A(n_1041),
.Y(n_1051)
);

INVx1_ASAP7_75t_L g1052 ( 
.A(n_1045),
.Y(n_1052)
);

INVx2_ASAP7_75t_L g1053 ( 
.A(n_1040),
.Y(n_1053)
);

INVx1_ASAP7_75t_L g1054 ( 
.A(n_1042),
.Y(n_1054)
);

INVxp67_ASAP7_75t_L g1055 ( 
.A(n_1042),
.Y(n_1055)
);

HB1xp67_ASAP7_75t_L g1056 ( 
.A(n_1042),
.Y(n_1056)
);

INVx2_ASAP7_75t_L g1057 ( 
.A(n_1042),
.Y(n_1057)
);

NAND2xp5_ASAP7_75t_L g1058 ( 
.A(n_1056),
.B(n_1036),
.Y(n_1058)
);

AND5x1_ASAP7_75t_L g1059 ( 
.A(n_1053),
.B(n_901),
.C(n_914),
.D(n_885),
.E(n_910),
.Y(n_1059)
);

XNOR2x2_ASAP7_75t_L g1060 ( 
.A(n_1054),
.B(n_897),
.Y(n_1060)
);

NAND2xp5_ASAP7_75t_L g1061 ( 
.A(n_1047),
.B(n_983),
.Y(n_1061)
);

CKINVDCx20_ASAP7_75t_R g1062 ( 
.A(n_1049),
.Y(n_1062)
);

NAND2xp5_ASAP7_75t_L g1063 ( 
.A(n_1057),
.B(n_957),
.Y(n_1063)
);

INVx1_ASAP7_75t_L g1064 ( 
.A(n_1055),
.Y(n_1064)
);

OA22x2_ASAP7_75t_L g1065 ( 
.A1(n_1051),
.A2(n_948),
.B1(n_965),
.B2(n_962),
.Y(n_1065)
);

NOR2xp67_ASAP7_75t_L g1066 ( 
.A(n_1048),
.B(n_1052),
.Y(n_1066)
);

XNOR2x2_ASAP7_75t_L g1067 ( 
.A(n_1050),
.B(n_912),
.Y(n_1067)
);

INVx1_ASAP7_75t_L g1068 ( 
.A(n_1052),
.Y(n_1068)
);

OAI321xp33_ASAP7_75t_L g1069 ( 
.A1(n_1058),
.A2(n_883),
.A3(n_912),
.B1(n_914),
.B2(n_898),
.C(n_878),
.Y(n_1069)
);

NAND5xp2_ASAP7_75t_L g1070 ( 
.A(n_1064),
.B(n_914),
.C(n_893),
.D(n_883),
.E(n_951),
.Y(n_1070)
);

NOR3xp33_ASAP7_75t_L g1071 ( 
.A(n_1066),
.B(n_898),
.C(n_910),
.Y(n_1071)
);

NAND2xp5_ASAP7_75t_L g1072 ( 
.A(n_1062),
.B(n_930),
.Y(n_1072)
);

NAND2xp5_ASAP7_75t_L g1073 ( 
.A(n_1068),
.B(n_930),
.Y(n_1073)
);

NOR2x1_ASAP7_75t_L g1074 ( 
.A(n_1063),
.B(n_948),
.Y(n_1074)
);

OAI21xp5_ASAP7_75t_SL g1075 ( 
.A1(n_1061),
.A2(n_1060),
.B(n_1059),
.Y(n_1075)
);

NAND4xp25_ASAP7_75t_SL g1076 ( 
.A(n_1065),
.B(n_1067),
.C(n_898),
.D(n_951),
.Y(n_1076)
);

NAND2xp5_ASAP7_75t_L g1077 ( 
.A(n_1075),
.B(n_968),
.Y(n_1077)
);

NOR2x1p5_ASAP7_75t_L g1078 ( 
.A(n_1072),
.B(n_948),
.Y(n_1078)
);

NOR2xp67_ASAP7_75t_L g1079 ( 
.A(n_1076),
.B(n_965),
.Y(n_1079)
);

NOR3xp33_ASAP7_75t_L g1080 ( 
.A(n_1071),
.B(n_910),
.C(n_885),
.Y(n_1080)
);

NAND4xp25_ASAP7_75t_L g1081 ( 
.A(n_1074),
.B(n_962),
.C(n_965),
.D(n_945),
.Y(n_1081)
);

INVx1_ASAP7_75t_L g1082 ( 
.A(n_1073),
.Y(n_1082)
);

NOR2x1_ASAP7_75t_L g1083 ( 
.A(n_1070),
.B(n_962),
.Y(n_1083)
);

AND3x1_ASAP7_75t_L g1084 ( 
.A(n_1069),
.B(n_940),
.C(n_916),
.Y(n_1084)
);

NOR2x1_ASAP7_75t_L g1085 ( 
.A(n_1076),
.B(n_965),
.Y(n_1085)
);

AOI22xp33_ASAP7_75t_L g1086 ( 
.A1(n_1077),
.A2(n_883),
.B1(n_939),
.B2(n_889),
.Y(n_1086)
);

NOR2xp33_ASAP7_75t_L g1087 ( 
.A(n_1082),
.B(n_883),
.Y(n_1087)
);

NOR2xp33_ASAP7_75t_L g1088 ( 
.A(n_1085),
.B(n_883),
.Y(n_1088)
);

INVxp33_ASAP7_75t_SL g1089 ( 
.A(n_1083),
.Y(n_1089)
);

NOR4xp75_ASAP7_75t_L g1090 ( 
.A(n_1079),
.B(n_940),
.C(n_949),
.D(n_883),
.Y(n_1090)
);

NOR2xp33_ASAP7_75t_L g1091 ( 
.A(n_1081),
.B(n_964),
.Y(n_1091)
);

NOR2x1p5_ASAP7_75t_L g1092 ( 
.A(n_1084),
.B(n_945),
.Y(n_1092)
);

AND2x4_ASAP7_75t_L g1093 ( 
.A(n_1078),
.B(n_964),
.Y(n_1093)
);

BUFx2_ASAP7_75t_L g1094 ( 
.A(n_1080),
.Y(n_1094)
);

OR2x2_ASAP7_75t_L g1095 ( 
.A(n_1093),
.B(n_947),
.Y(n_1095)
);

NAND4xp75_ASAP7_75t_L g1096 ( 
.A(n_1087),
.B(n_889),
.C(n_941),
.D(n_893),
.Y(n_1096)
);

NAND2xp5_ASAP7_75t_L g1097 ( 
.A(n_1089),
.B(n_968),
.Y(n_1097)
);

INVxp67_ASAP7_75t_SL g1098 ( 
.A(n_1094),
.Y(n_1098)
);

NAND4xp75_ASAP7_75t_L g1099 ( 
.A(n_1088),
.B(n_889),
.C(n_941),
.D(n_949),
.Y(n_1099)
);

NOR2x1_ASAP7_75t_L g1100 ( 
.A(n_1092),
.B(n_943),
.Y(n_1100)
);

INVx2_ASAP7_75t_L g1101 ( 
.A(n_1093),
.Y(n_1101)
);

NAND2xp33_ASAP7_75t_SL g1102 ( 
.A(n_1086),
.B(n_1090),
.Y(n_1102)
);

NOR2xp33_ASAP7_75t_L g1103 ( 
.A(n_1091),
.B(n_966),
.Y(n_1103)
);

AND4x1_ASAP7_75t_L g1104 ( 
.A(n_1087),
.B(n_917),
.C(n_916),
.D(n_934),
.Y(n_1104)
);

INVx1_ASAP7_75t_L g1105 ( 
.A(n_1089),
.Y(n_1105)
);

NAND2xp5_ASAP7_75t_L g1106 ( 
.A(n_1089),
.B(n_963),
.Y(n_1106)
);

XNOR2x1_ASAP7_75t_L g1107 ( 
.A(n_1090),
.B(n_908),
.Y(n_1107)
);

AOI21xp5_ASAP7_75t_L g1108 ( 
.A1(n_1105),
.A2(n_1098),
.B(n_1102),
.Y(n_1108)
);

INVx1_ASAP7_75t_L g1109 ( 
.A(n_1101),
.Y(n_1109)
);

OAI21xp5_ASAP7_75t_L g1110 ( 
.A1(n_1097),
.A2(n_966),
.B(n_963),
.Y(n_1110)
);

NOR3xp33_ASAP7_75t_L g1111 ( 
.A(n_1106),
.B(n_908),
.C(n_905),
.Y(n_1111)
);

INVx1_ASAP7_75t_L g1112 ( 
.A(n_1100),
.Y(n_1112)
);

NAND2xp5_ASAP7_75t_L g1113 ( 
.A(n_1107),
.B(n_939),
.Y(n_1113)
);

INVx2_ASAP7_75t_L g1114 ( 
.A(n_1095),
.Y(n_1114)
);

NAND2xp5_ASAP7_75t_L g1115 ( 
.A(n_1103),
.B(n_1104),
.Y(n_1115)
);

AOI22xp5_ASAP7_75t_L g1116 ( 
.A1(n_1099),
.A2(n_889),
.B1(n_939),
.B2(n_917),
.Y(n_1116)
);

INVx1_ASAP7_75t_L g1117 ( 
.A(n_1109),
.Y(n_1117)
);

AOI22xp5_ASAP7_75t_L g1118 ( 
.A1(n_1112),
.A2(n_1096),
.B1(n_899),
.B2(n_941),
.Y(n_1118)
);

INVx1_ASAP7_75t_SL g1119 ( 
.A(n_1114),
.Y(n_1119)
);

AOI22xp5_ASAP7_75t_L g1120 ( 
.A1(n_1108),
.A2(n_941),
.B1(n_934),
.B2(n_931),
.Y(n_1120)
);

AOI22xp5_ASAP7_75t_L g1121 ( 
.A1(n_1115),
.A2(n_931),
.B1(n_874),
.B2(n_905),
.Y(n_1121)
);

HB1xp67_ASAP7_75t_L g1122 ( 
.A(n_1113),
.Y(n_1122)
);

OAI22xp5_ASAP7_75t_L g1123 ( 
.A1(n_1119),
.A2(n_1117),
.B1(n_1118),
.B2(n_1122),
.Y(n_1123)
);

INVx2_ASAP7_75t_L g1124 ( 
.A(n_1121),
.Y(n_1124)
);

OAI22x1_ASAP7_75t_L g1125 ( 
.A1(n_1120),
.A2(n_1116),
.B1(n_1111),
.B2(n_1110),
.Y(n_1125)
);

OAI21xp5_ASAP7_75t_L g1126 ( 
.A1(n_1123),
.A2(n_905),
.B(n_908),
.Y(n_1126)
);

INVx1_ASAP7_75t_L g1127 ( 
.A(n_1126),
.Y(n_1127)
);

OAI21xp5_ASAP7_75t_L g1128 ( 
.A1(n_1127),
.A2(n_1124),
.B(n_1125),
.Y(n_1128)
);

OAI22xp5_ASAP7_75t_L g1129 ( 
.A1(n_1128),
.A2(n_943),
.B1(n_932),
.B2(n_929),
.Y(n_1129)
);

OAI22xp33_ASAP7_75t_L g1130 ( 
.A1(n_1128),
.A2(n_874),
.B1(n_929),
.B2(n_925),
.Y(n_1130)
);

AOI22xp5_ASAP7_75t_L g1131 ( 
.A1(n_1128),
.A2(n_874),
.B1(n_931),
.B2(n_870),
.Y(n_1131)
);

AOI21xp5_ASAP7_75t_L g1132 ( 
.A1(n_1130),
.A2(n_874),
.B(n_931),
.Y(n_1132)
);

AOI21xp5_ASAP7_75t_L g1133 ( 
.A1(n_1129),
.A2(n_874),
.B(n_870),
.Y(n_1133)
);

OAI21xp5_ASAP7_75t_L g1134 ( 
.A1(n_1131),
.A2(n_870),
.B(n_942),
.Y(n_1134)
);

OA21x2_ASAP7_75t_L g1135 ( 
.A1(n_1132),
.A2(n_946),
.B(n_942),
.Y(n_1135)
);

AO21x2_ASAP7_75t_L g1136 ( 
.A1(n_1133),
.A2(n_1134),
.B(n_870),
.Y(n_1136)
);

AOI221xp5_ASAP7_75t_L g1137 ( 
.A1(n_1136),
.A2(n_946),
.B1(n_938),
.B2(n_886),
.C(n_884),
.Y(n_1137)
);

AOI211xp5_ASAP7_75t_L g1138 ( 
.A1(n_1137),
.A2(n_1135),
.B(n_886),
.C(n_938),
.Y(n_1138)
);


endmodule