module fake_jpeg_14056_n_565 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_565);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_565;

wire n_529;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_547;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_419;
wire n_378;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_10),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

CKINVDCx14_ASAP7_75t_R g24 ( 
.A(n_16),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_4),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_2),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_18),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_1),
.Y(n_33)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_18),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_17),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_0),
.Y(n_36)
);

INVx11_ASAP7_75t_L g37 ( 
.A(n_1),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_14),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_15),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_16),
.Y(n_40)
);

BUFx16f_ASAP7_75t_L g41 ( 
.A(n_0),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_12),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_7),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_15),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_4),
.Y(n_45)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_14),
.Y(n_46)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_10),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_16),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_12),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_8),
.Y(n_50)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_2),
.Y(n_51)
);

INVxp67_ASAP7_75t_L g52 ( 
.A(n_6),
.Y(n_52)
);

BUFx8_ASAP7_75t_L g53 ( 
.A(n_17),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_20),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g141 ( 
.A(n_54),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g55 ( 
.A(n_21),
.B(n_18),
.C(n_17),
.Y(n_55)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_55),
.B(n_48),
.C(n_35),
.Y(n_115)
);

BUFx5_ASAP7_75t_L g56 ( 
.A(n_37),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g134 ( 
.A(n_56),
.Y(n_134)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_32),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g164 ( 
.A(n_57),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_20),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_58),
.Y(n_145)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_20),
.Y(n_59)
);

INVx5_ASAP7_75t_L g111 ( 
.A(n_59),
.Y(n_111)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_21),
.Y(n_60)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_60),
.Y(n_125)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_26),
.Y(n_61)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_61),
.Y(n_146)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_26),
.Y(n_62)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_62),
.Y(n_148)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_53),
.Y(n_63)
);

INVx5_ASAP7_75t_L g132 ( 
.A(n_63),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_37),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_64),
.B(n_67),
.Y(n_121)
);

INVx8_ASAP7_75t_L g65 ( 
.A(n_43),
.Y(n_65)
);

INVx5_ASAP7_75t_L g144 ( 
.A(n_65),
.Y(n_144)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_51),
.Y(n_66)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_66),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_37),
.Y(n_67)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_53),
.Y(n_68)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_68),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_43),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g152 ( 
.A(n_69),
.Y(n_152)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_23),
.Y(n_70)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_70),
.Y(n_110)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_23),
.Y(n_71)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_71),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_43),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g176 ( 
.A(n_72),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_47),
.Y(n_73)
);

INVx6_ASAP7_75t_L g159 ( 
.A(n_73),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_47),
.Y(n_74)
);

INVx6_ASAP7_75t_L g168 ( 
.A(n_74),
.Y(n_168)
);

INVx6_ASAP7_75t_L g75 ( 
.A(n_47),
.Y(n_75)
);

INVx6_ASAP7_75t_L g171 ( 
.A(n_75),
.Y(n_171)
);

BUFx3_ASAP7_75t_L g76 ( 
.A(n_32),
.Y(n_76)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_76),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_28),
.Y(n_77)
);

INVx8_ASAP7_75t_L g142 ( 
.A(n_77),
.Y(n_142)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_32),
.Y(n_78)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_78),
.Y(n_118)
);

INVx11_ASAP7_75t_L g79 ( 
.A(n_41),
.Y(n_79)
);

INVx11_ASAP7_75t_L g129 ( 
.A(n_79),
.Y(n_129)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_32),
.Y(n_80)
);

INVx4_ASAP7_75t_L g119 ( 
.A(n_80),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_28),
.Y(n_81)
);

BUFx2_ASAP7_75t_L g167 ( 
.A(n_81),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_31),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_82),
.B(n_84),
.Y(n_135)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_32),
.Y(n_83)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_83),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_31),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_28),
.Y(n_85)
);

INVx4_ASAP7_75t_L g163 ( 
.A(n_85),
.Y(n_163)
);

INVx6_ASAP7_75t_L g86 ( 
.A(n_39),
.Y(n_86)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_86),
.Y(n_158)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_53),
.Y(n_87)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_87),
.Y(n_124)
);

INVx6_ASAP7_75t_L g88 ( 
.A(n_39),
.Y(n_88)
);

INVx3_ASAP7_75t_L g157 ( 
.A(n_88),
.Y(n_157)
);

BUFx12f_ASAP7_75t_L g89 ( 
.A(n_53),
.Y(n_89)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_89),
.Y(n_126)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_51),
.Y(n_90)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_90),
.Y(n_114)
);

INVx11_ASAP7_75t_L g91 ( 
.A(n_41),
.Y(n_91)
);

INVx11_ASAP7_75t_L g139 ( 
.A(n_91),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_39),
.Y(n_92)
);

INVx3_ASAP7_75t_L g177 ( 
.A(n_92),
.Y(n_177)
);

BUFx5_ASAP7_75t_L g93 ( 
.A(n_34),
.Y(n_93)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_93),
.Y(n_127)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_40),
.Y(n_94)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_94),
.Y(n_128)
);

INVx2_ASAP7_75t_R g95 ( 
.A(n_24),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_95),
.B(n_102),
.Y(n_153)
);

BUFx3_ASAP7_75t_L g96 ( 
.A(n_49),
.Y(n_96)
);

INVx3_ASAP7_75t_L g130 ( 
.A(n_96),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_40),
.Y(n_97)
);

INVx3_ASAP7_75t_L g131 ( 
.A(n_97),
.Y(n_131)
);

INVx8_ASAP7_75t_L g98 ( 
.A(n_34),
.Y(n_98)
);

INVx3_ASAP7_75t_L g137 ( 
.A(n_98),
.Y(n_137)
);

INVx11_ASAP7_75t_L g99 ( 
.A(n_41),
.Y(n_99)
);

INVx11_ASAP7_75t_L g161 ( 
.A(n_99),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_40),
.Y(n_100)
);

INVx3_ASAP7_75t_L g154 ( 
.A(n_100),
.Y(n_154)
);

INVx6_ASAP7_75t_L g101 ( 
.A(n_34),
.Y(n_101)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_101),
.Y(n_136)
);

AND2x2_ASAP7_75t_L g102 ( 
.A(n_40),
.B(n_0),
.Y(n_102)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_35),
.Y(n_103)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_103),
.Y(n_149)
);

INVx8_ASAP7_75t_L g104 ( 
.A(n_41),
.Y(n_104)
);

INVx11_ASAP7_75t_L g172 ( 
.A(n_104),
.Y(n_172)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_40),
.Y(n_105)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_105),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_38),
.B(n_0),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_106),
.B(n_3),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_49),
.Y(n_107)
);

INVx4_ASAP7_75t_SL g123 ( 
.A(n_107),
.Y(n_123)
);

INVx6_ASAP7_75t_SL g108 ( 
.A(n_52),
.Y(n_108)
);

INVx6_ASAP7_75t_SL g117 ( 
.A(n_108),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_38),
.B(n_2),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_109),
.B(n_22),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_115),
.B(n_33),
.C(n_29),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_120),
.B(n_170),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_79),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_133),
.B(n_156),
.Y(n_200)
);

AO22x1_ASAP7_75t_SL g138 ( 
.A1(n_102),
.A2(n_48),
.B1(n_50),
.B2(n_27),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_138),
.A2(n_87),
.B1(n_42),
.B2(n_36),
.Y(n_181)
);

BUFx12_ASAP7_75t_L g140 ( 
.A(n_91),
.Y(n_140)
);

INVx13_ASAP7_75t_L g206 ( 
.A(n_140),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_55),
.A2(n_46),
.B1(n_44),
.B2(n_24),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_143),
.A2(n_92),
.B1(n_65),
.B2(n_58),
.Y(n_239)
);

INVx13_ASAP7_75t_L g147 ( 
.A(n_99),
.Y(n_147)
);

INVx13_ASAP7_75t_L g236 ( 
.A(n_147),
.Y(n_236)
);

INVx6_ASAP7_75t_SL g155 ( 
.A(n_104),
.Y(n_155)
);

CKINVDCx9p33_ASAP7_75t_R g197 ( 
.A(n_155),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_78),
.Y(n_156)
);

AND2x2_ASAP7_75t_L g193 ( 
.A(n_160),
.B(n_89),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_95),
.B(n_22),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_162),
.B(n_166),
.Y(n_185)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_105),
.Y(n_165)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_165),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_83),
.B(n_45),
.Y(n_166)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_68),
.Y(n_169)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_169),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_63),
.B(n_36),
.Y(n_170)
);

HAxp5_ASAP7_75t_SL g173 ( 
.A(n_63),
.B(n_42),
.CON(n_173),
.SN(n_173)
);

OR2x2_ASAP7_75t_L g203 ( 
.A(n_173),
.B(n_46),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_98),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_174),
.B(n_175),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_59),
.Y(n_175)
);

INVx4_ASAP7_75t_L g178 ( 
.A(n_123),
.Y(n_178)
);

BUFx2_ASAP7_75t_L g256 ( 
.A(n_178),
.Y(n_256)
);

INVx3_ASAP7_75t_L g180 ( 
.A(n_111),
.Y(n_180)
);

INVx3_ASAP7_75t_L g273 ( 
.A(n_180),
.Y(n_273)
);

NAND2xp33_ASAP7_75t_SL g245 ( 
.A(n_181),
.B(n_203),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_135),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_182),
.B(n_213),
.Y(n_244)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_158),
.Y(n_183)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_183),
.Y(n_242)
);

CKINVDCx12_ASAP7_75t_R g184 ( 
.A(n_117),
.Y(n_184)
);

CKINVDCx16_ASAP7_75t_R g248 ( 
.A(n_184),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_153),
.B(n_30),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g251 ( 
.A(n_186),
.B(n_190),
.Y(n_251)
);

AOI22xp33_ASAP7_75t_SL g187 ( 
.A1(n_173),
.A2(n_89),
.B1(n_75),
.B2(n_46),
.Y(n_187)
);

AOI22xp33_ASAP7_75t_SL g282 ( 
.A1(n_187),
.A2(n_235),
.B1(n_238),
.B2(n_241),
.Y(n_282)
);

CKINVDCx12_ASAP7_75t_R g188 ( 
.A(n_172),
.Y(n_188)
);

BUFx12f_ASAP7_75t_L g286 ( 
.A(n_188),
.Y(n_286)
);

INVx3_ASAP7_75t_L g189 ( 
.A(n_111),
.Y(n_189)
);

INVx3_ASAP7_75t_L g281 ( 
.A(n_189),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_110),
.B(n_45),
.Y(n_190)
);

INVx2_ASAP7_75t_SL g191 ( 
.A(n_129),
.Y(n_191)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_191),
.Y(n_261)
);

INVx5_ASAP7_75t_L g192 ( 
.A(n_132),
.Y(n_192)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_192),
.Y(n_247)
);

OAI21xp33_ASAP7_75t_L g278 ( 
.A1(n_193),
.A2(n_215),
.B(n_218),
.Y(n_278)
);

INVx5_ASAP7_75t_L g194 ( 
.A(n_132),
.Y(n_194)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_194),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_195),
.B(n_208),
.C(n_237),
.Y(n_280)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_136),
.Y(n_196)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_196),
.Y(n_263)
);

BUFx6f_ASAP7_75t_L g198 ( 
.A(n_141),
.Y(n_198)
);

BUFx6f_ASAP7_75t_L g284 ( 
.A(n_198),
.Y(n_284)
);

INVx5_ASAP7_75t_L g199 ( 
.A(n_172),
.Y(n_199)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_199),
.Y(n_270)
);

BUFx16f_ASAP7_75t_L g201 ( 
.A(n_129),
.Y(n_201)
);

BUFx3_ASAP7_75t_L g255 ( 
.A(n_201),
.Y(n_255)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_128),
.Y(n_202)
);

INVx2_ASAP7_75t_L g291 ( 
.A(n_202),
.Y(n_291)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_112),
.Y(n_204)
);

INVx1_ASAP7_75t_SL g260 ( 
.A(n_204),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_114),
.A2(n_101),
.B1(n_86),
.B2(n_88),
.Y(n_205)
);

AOI22xp33_ASAP7_75t_L g243 ( 
.A1(n_205),
.A2(n_167),
.B1(n_176),
.B2(n_145),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_149),
.B(n_148),
.C(n_125),
.Y(n_208)
);

INVx8_ASAP7_75t_L g209 ( 
.A(n_159),
.Y(n_209)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_209),
.Y(n_268)
);

AND2x4_ASAP7_75t_L g210 ( 
.A(n_146),
.B(n_57),
.Y(n_210)
);

AND2x2_ASAP7_75t_L g275 ( 
.A(n_210),
.B(n_232),
.Y(n_275)
);

CKINVDCx12_ASAP7_75t_R g211 ( 
.A(n_147),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_211),
.Y(n_249)
);

INVxp67_ASAP7_75t_L g213 ( 
.A(n_139),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_121),
.B(n_44),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_214),
.B(n_221),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_138),
.B(n_29),
.Y(n_215)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_150),
.Y(n_217)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_217),
.Y(n_257)
);

AND2x2_ASAP7_75t_L g218 ( 
.A(n_151),
.B(n_80),
.Y(n_218)
);

INVx3_ASAP7_75t_L g219 ( 
.A(n_144),
.Y(n_219)
);

BUFx3_ASAP7_75t_L g276 ( 
.A(n_219),
.Y(n_276)
);

INVx4_ASAP7_75t_L g220 ( 
.A(n_123),
.Y(n_220)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_220),
.Y(n_289)
);

BUFx12f_ASAP7_75t_L g221 ( 
.A(n_164),
.Y(n_221)
);

INVx4_ASAP7_75t_L g222 ( 
.A(n_139),
.Y(n_222)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_222),
.Y(n_293)
);

BUFx6f_ASAP7_75t_L g223 ( 
.A(n_141),
.Y(n_223)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_223),
.Y(n_269)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_118),
.Y(n_224)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_224),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_140),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_225),
.B(n_227),
.Y(n_254)
);

NAND2x1p5_ASAP7_75t_L g226 ( 
.A(n_161),
.B(n_100),
.Y(n_226)
);

OAI21xp5_ASAP7_75t_L g277 ( 
.A1(n_226),
.A2(n_167),
.B(n_76),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_116),
.B(n_44),
.Y(n_227)
);

CKINVDCx16_ASAP7_75t_R g228 ( 
.A(n_161),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_228),
.B(n_229),
.Y(n_266)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_157),
.Y(n_229)
);

OR2x2_ASAP7_75t_L g230 ( 
.A(n_124),
.B(n_50),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_230),
.B(n_231),
.Y(n_274)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_122),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_113),
.B(n_19),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_157),
.B(n_33),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_233),
.B(n_30),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_L g234 ( 
.A1(n_171),
.A2(n_85),
.B1(n_77),
.B2(n_81),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_L g296 ( 
.A1(n_234),
.A2(n_239),
.B1(n_197),
.B2(n_223),
.Y(n_296)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_131),
.Y(n_235)
);

AND2x2_ASAP7_75t_SL g237 ( 
.A(n_113),
.B(n_96),
.Y(n_237)
);

BUFx2_ASAP7_75t_L g238 ( 
.A(n_144),
.Y(n_238)
);

INVx4_ASAP7_75t_L g240 ( 
.A(n_126),
.Y(n_240)
);

AOI22xp33_ASAP7_75t_SL g297 ( 
.A1(n_240),
.A2(n_49),
.B1(n_5),
.B2(n_6),
.Y(n_297)
);

INVx3_ASAP7_75t_L g241 ( 
.A(n_154),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_L g299 ( 
.A1(n_243),
.A2(n_191),
.B1(n_198),
.B2(n_220),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_239),
.A2(n_171),
.B1(n_69),
.B2(n_54),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_250),
.A2(n_253),
.B1(n_265),
.B2(n_272),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_SL g319 ( 
.A(n_252),
.B(n_178),
.Y(n_319)
);

OAI22xp33_ASAP7_75t_SL g253 ( 
.A1(n_203),
.A2(n_137),
.B1(n_177),
.B2(n_163),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_185),
.B(n_19),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_258),
.B(n_264),
.Y(n_303)
);

OAI21xp5_ASAP7_75t_SL g262 ( 
.A1(n_230),
.A2(n_27),
.B(n_25),
.Y(n_262)
);

OR2x2_ASAP7_75t_L g324 ( 
.A(n_262),
.B(n_236),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_208),
.B(n_25),
.Y(n_264)
);

OAI22xp33_ASAP7_75t_L g265 ( 
.A1(n_187),
.A2(n_168),
.B1(n_159),
.B2(n_163),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_200),
.B(n_119),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_267),
.B(n_279),
.Y(n_312)
);

OAI22xp33_ASAP7_75t_L g272 ( 
.A1(n_226),
.A2(n_168),
.B1(n_74),
.B2(n_73),
.Y(n_272)
);

AND2x2_ASAP7_75t_L g315 ( 
.A(n_277),
.B(n_237),
.Y(n_315)
);

A2O1A1Ixp33_ASAP7_75t_L g279 ( 
.A1(n_195),
.A2(n_140),
.B(n_119),
.C(n_130),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_179),
.B(n_142),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_283),
.B(n_285),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_212),
.B(n_142),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_205),
.A2(n_72),
.B1(n_177),
.B2(n_176),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_287),
.A2(n_292),
.B1(n_294),
.B2(n_295),
.Y(n_305)
);

AOI22xp33_ASAP7_75t_SL g288 ( 
.A1(n_238),
.A2(n_164),
.B1(n_134),
.B2(n_127),
.Y(n_288)
);

AOI22xp33_ASAP7_75t_SL g335 ( 
.A1(n_288),
.A2(n_297),
.B1(n_221),
.B2(n_201),
.Y(n_335)
);

AOI21xp5_ASAP7_75t_SL g290 ( 
.A1(n_193),
.A2(n_134),
.B(n_4),
.Y(n_290)
);

OAI21xp5_ASAP7_75t_L g337 ( 
.A1(n_290),
.A2(n_3),
.B(n_5),
.Y(n_337)
);

OAI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_209),
.A2(n_152),
.B1(n_145),
.B2(n_210),
.Y(n_292)
);

OAI22xp33_ASAP7_75t_SL g294 ( 
.A1(n_197),
.A2(n_152),
.B1(n_97),
.B2(n_107),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_SL g295 ( 
.A1(n_210),
.A2(n_49),
.B1(n_93),
.B2(n_56),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_296),
.A2(n_250),
.B1(n_287),
.B2(n_292),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_267),
.B(n_216),
.Y(n_298)
);

CKINVDCx14_ASAP7_75t_R g374 ( 
.A(n_298),
.Y(n_374)
);

INVxp67_ASAP7_75t_SL g384 ( 
.A(n_299),
.Y(n_384)
);

INVx3_ASAP7_75t_L g300 ( 
.A(n_276),
.Y(n_300)
);

INVx2_ASAP7_75t_SL g381 ( 
.A(n_300),
.Y(n_381)
);

AO22x1_ASAP7_75t_L g301 ( 
.A1(n_272),
.A2(n_210),
.B1(n_213),
.B2(n_222),
.Y(n_301)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_301),
.Y(n_350)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_261),
.Y(n_302)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_302),
.Y(n_356)
);

INVx5_ASAP7_75t_L g306 ( 
.A(n_286),
.Y(n_306)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_306),
.Y(n_372)
);

OAI22xp5_ASAP7_75t_L g348 ( 
.A1(n_307),
.A2(n_335),
.B1(n_344),
.B2(n_282),
.Y(n_348)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_257),
.Y(n_308)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_308),
.Y(n_377)
);

INVx8_ASAP7_75t_L g309 ( 
.A(n_284),
.Y(n_309)
);

INVx3_ASAP7_75t_SL g367 ( 
.A(n_309),
.Y(n_367)
);

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_285),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g365 ( 
.A(n_310),
.B(n_318),
.Y(n_365)
);

OAI22xp5_ASAP7_75t_SL g311 ( 
.A1(n_280),
.A2(n_241),
.B1(n_189),
.B2(n_180),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_L g376 ( 
.A1(n_311),
.A2(n_332),
.B1(n_336),
.B2(n_256),
.Y(n_376)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_280),
.B(n_218),
.C(n_237),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g368 ( 
.A(n_313),
.B(n_317),
.C(n_329),
.Y(n_368)
);

BUFx2_ASAP7_75t_L g314 ( 
.A(n_268),
.Y(n_314)
);

INVxp67_ASAP7_75t_L g357 ( 
.A(n_314),
.Y(n_357)
);

AND2x2_ASAP7_75t_L g347 ( 
.A(n_315),
.B(n_325),
.Y(n_347)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_261),
.Y(n_316)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_316),
.Y(n_378)
);

XNOR2xp5_ASAP7_75t_L g317 ( 
.A(n_264),
.B(n_207),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_SL g318 ( 
.A(n_251),
.B(n_240),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g385 ( 
.A(n_319),
.B(n_320),
.Y(n_385)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_283),
.B(n_192),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_291),
.Y(n_321)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_321),
.Y(n_380)
);

CKINVDCx16_ASAP7_75t_R g322 ( 
.A(n_244),
.Y(n_322)
);

CKINVDCx16_ASAP7_75t_R g370 ( 
.A(n_322),
.Y(n_370)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_249),
.B(n_194),
.Y(n_323)
);

INVxp67_ASAP7_75t_L g366 ( 
.A(n_323),
.Y(n_366)
);

INVxp67_ASAP7_75t_L g386 ( 
.A(n_324),
.Y(n_386)
);

INVx8_ASAP7_75t_L g325 ( 
.A(n_284),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_SL g326 ( 
.A(n_248),
.B(n_49),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g352 ( 
.A(n_326),
.Y(n_352)
);

INVx6_ASAP7_75t_L g327 ( 
.A(n_273),
.Y(n_327)
);

AND2x2_ASAP7_75t_L g353 ( 
.A(n_327),
.B(n_328),
.Y(n_353)
);

AND2x2_ASAP7_75t_L g328 ( 
.A(n_275),
.B(n_219),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_275),
.B(n_254),
.C(n_245),
.Y(n_329)
);

INVx2_ASAP7_75t_L g331 ( 
.A(n_273),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_331),
.B(n_334),
.Y(n_354)
);

OAI22xp5_ASAP7_75t_L g332 ( 
.A1(n_252),
.A2(n_199),
.B1(n_236),
.B2(n_206),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_275),
.B(n_206),
.C(n_221),
.Y(n_333)
);

XNOR2xp5_ASAP7_75t_L g371 ( 
.A(n_333),
.B(n_259),
.Y(n_371)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_271),
.Y(n_334)
);

OAI22xp5_ASAP7_75t_SL g336 ( 
.A1(n_277),
.A2(n_201),
.B1(n_5),
.B2(n_6),
.Y(n_336)
);

OAI21xp5_ASAP7_75t_L g351 ( 
.A1(n_337),
.A2(n_339),
.B(n_343),
.Y(n_351)
);

INVx5_ASAP7_75t_L g338 ( 
.A(n_286),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_338),
.B(n_340),
.Y(n_359)
);

OAI21xp5_ASAP7_75t_L g339 ( 
.A1(n_274),
.A2(n_13),
.B(n_6),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_271),
.Y(n_340)
);

INVx2_ASAP7_75t_L g341 ( 
.A(n_281),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_341),
.B(n_345),
.Y(n_369)
);

CKINVDCx12_ASAP7_75t_R g342 ( 
.A(n_286),
.Y(n_342)
);

CKINVDCx20_ASAP7_75t_R g358 ( 
.A(n_342),
.Y(n_358)
);

AOI32xp33_ASAP7_75t_L g343 ( 
.A1(n_279),
.A2(n_278),
.A3(n_258),
.B1(n_290),
.B2(n_246),
.Y(n_343)
);

AOI22xp33_ASAP7_75t_SL g344 ( 
.A1(n_295),
.A2(n_3),
.B1(n_7),
.B2(n_8),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_291),
.Y(n_345)
);

XOR2xp5_ASAP7_75t_L g346 ( 
.A(n_317),
.B(n_266),
.Y(n_346)
);

MAJIxp5_ASAP7_75t_L g405 ( 
.A(n_346),
.B(n_364),
.C(n_345),
.Y(n_405)
);

AOI22xp5_ASAP7_75t_SL g410 ( 
.A1(n_348),
.A2(n_300),
.B1(n_306),
.B2(n_338),
.Y(n_410)
);

OAI22xp5_ASAP7_75t_SL g349 ( 
.A1(n_312),
.A2(n_265),
.B1(n_268),
.B2(n_269),
.Y(n_349)
);

AOI22xp5_ASAP7_75t_L g412 ( 
.A1(n_349),
.A2(n_363),
.B1(n_263),
.B2(n_255),
.Y(n_412)
);

XNOR2xp5_ASAP7_75t_SL g355 ( 
.A(n_329),
.B(n_262),
.Y(n_355)
);

XOR2xp5_ASAP7_75t_L g399 ( 
.A(n_355),
.B(n_371),
.Y(n_399)
);

AOI22xp5_ASAP7_75t_SL g360 ( 
.A1(n_312),
.A2(n_281),
.B1(n_276),
.B2(n_286),
.Y(n_360)
);

OAI21xp5_ASAP7_75t_SL g394 ( 
.A1(n_360),
.A2(n_301),
.B(n_328),
.Y(n_394)
);

CKINVDCx20_ASAP7_75t_R g361 ( 
.A(n_330),
.Y(n_361)
);

NOR2xp33_ASAP7_75t_L g388 ( 
.A(n_361),
.B(n_362),
.Y(n_388)
);

CKINVDCx20_ASAP7_75t_R g362 ( 
.A(n_330),
.Y(n_362)
);

OAI22xp5_ASAP7_75t_SL g363 ( 
.A1(n_307),
.A2(n_269),
.B1(n_289),
.B2(n_293),
.Y(n_363)
);

XOR2xp5_ASAP7_75t_L g364 ( 
.A(n_313),
.B(n_260),
.Y(n_364)
);

OAI22xp5_ASAP7_75t_L g373 ( 
.A1(n_304),
.A2(n_259),
.B1(n_247),
.B2(n_270),
.Y(n_373)
);

OAI22xp5_ASAP7_75t_L g391 ( 
.A1(n_373),
.A2(n_376),
.B1(n_379),
.B2(n_305),
.Y(n_391)
);

AOI21xp5_ASAP7_75t_L g375 ( 
.A1(n_315),
.A2(n_256),
.B(n_270),
.Y(n_375)
);

AOI21xp5_ASAP7_75t_L g395 ( 
.A1(n_375),
.A2(n_315),
.B(n_328),
.Y(n_395)
);

AOI22xp5_ASAP7_75t_L g379 ( 
.A1(n_311),
.A2(n_247),
.B1(n_260),
.B2(n_242),
.Y(n_379)
);

CKINVDCx20_ASAP7_75t_R g382 ( 
.A(n_324),
.Y(n_382)
);

NOR2xp33_ASAP7_75t_L g402 ( 
.A(n_382),
.B(n_339),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_303),
.B(n_242),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_383),
.B(n_316),
.Y(n_398)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_356),
.Y(n_387)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_387),
.Y(n_426)
);

BUFx12_ASAP7_75t_L g389 ( 
.A(n_358),
.Y(n_389)
);

CKINVDCx20_ASAP7_75t_R g437 ( 
.A(n_389),
.Y(n_437)
);

INVx8_ASAP7_75t_L g390 ( 
.A(n_370),
.Y(n_390)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_390),
.Y(n_435)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_391),
.Y(n_454)
);

AOI22xp33_ASAP7_75t_L g392 ( 
.A1(n_384),
.A2(n_336),
.B1(n_304),
.B2(n_301),
.Y(n_392)
);

OAI22xp5_ASAP7_75t_L g445 ( 
.A1(n_392),
.A2(n_410),
.B1(n_412),
.B2(n_418),
.Y(n_445)
);

CKINVDCx20_ASAP7_75t_R g393 ( 
.A(n_354),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_393),
.B(n_397),
.Y(n_430)
);

AND2x2_ASAP7_75t_L g425 ( 
.A(n_394),
.B(n_347),
.Y(n_425)
);

OAI21xp5_ASAP7_75t_SL g444 ( 
.A1(n_395),
.A2(n_401),
.B(n_403),
.Y(n_444)
);

XNOR2xp5_ASAP7_75t_L g396 ( 
.A(n_364),
.B(n_303),
.Y(n_396)
);

MAJIxp5_ASAP7_75t_L g429 ( 
.A(n_396),
.B(n_405),
.C(n_421),
.Y(n_429)
);

CKINVDCx20_ASAP7_75t_R g397 ( 
.A(n_354),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_398),
.B(n_416),
.Y(n_434)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_356),
.Y(n_400)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_400),
.Y(n_446)
);

NOR2x1_ASAP7_75t_L g401 ( 
.A(n_347),
.B(n_333),
.Y(n_401)
);

CKINVDCx14_ASAP7_75t_R g441 ( 
.A(n_402),
.Y(n_441)
);

OAI21xp5_ASAP7_75t_SL g403 ( 
.A1(n_386),
.A2(n_305),
.B(n_302),
.Y(n_403)
);

OAI21xp5_ASAP7_75t_SL g404 ( 
.A1(n_386),
.A2(n_341),
.B(n_331),
.Y(n_404)
);

O2A1O1Ixp33_ASAP7_75t_L g428 ( 
.A1(n_404),
.A2(n_406),
.B(n_419),
.C(n_353),
.Y(n_428)
);

OAI21xp5_ASAP7_75t_SL g406 ( 
.A1(n_382),
.A2(n_337),
.B(n_321),
.Y(n_406)
);

OAI21xp33_ASAP7_75t_L g407 ( 
.A1(n_360),
.A2(n_361),
.B(n_362),
.Y(n_407)
);

AOI21xp33_ASAP7_75t_L g436 ( 
.A1(n_407),
.A2(n_347),
.B(n_366),
.Y(n_436)
);

OAI22xp5_ASAP7_75t_SL g408 ( 
.A1(n_350),
.A2(n_314),
.B1(n_327),
.B2(n_325),
.Y(n_408)
);

AOI22xp5_ASAP7_75t_L g427 ( 
.A1(n_408),
.A2(n_367),
.B1(n_363),
.B2(n_381),
.Y(n_427)
);

CKINVDCx16_ASAP7_75t_R g409 ( 
.A(n_359),
.Y(n_409)
);

INVxp67_ASAP7_75t_SL g433 ( 
.A(n_409),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_383),
.B(n_309),
.Y(n_411)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_411),
.Y(n_451)
);

OA22x2_ASAP7_75t_L g413 ( 
.A1(n_350),
.A2(n_263),
.B1(n_255),
.B2(n_8),
.Y(n_413)
);

INVx2_ASAP7_75t_SL g431 ( 
.A(n_413),
.Y(n_431)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_378),
.Y(n_414)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_414),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_365),
.B(n_3),
.Y(n_415)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_415),
.Y(n_453)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_378),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_377),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_417),
.B(n_420),
.Y(n_443)
);

AOI22xp5_ASAP7_75t_L g418 ( 
.A1(n_349),
.A2(n_13),
.B1(n_8),
.B2(n_9),
.Y(n_418)
);

AO21x1_ASAP7_75t_L g419 ( 
.A1(n_351),
.A2(n_7),
.B(n_9),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_385),
.B(n_366),
.Y(n_420)
);

XOR2xp5_ASAP7_75t_L g421 ( 
.A(n_368),
.B(n_7),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_377),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_422),
.B(n_380),
.Y(n_448)
);

XOR2xp5_ASAP7_75t_L g423 ( 
.A(n_399),
.B(n_368),
.Y(n_423)
);

XOR2xp5_ASAP7_75t_L g462 ( 
.A(n_423),
.B(n_401),
.Y(n_462)
);

NOR2xp33_ASAP7_75t_SL g424 ( 
.A(n_420),
.B(n_352),
.Y(n_424)
);

NOR2xp33_ASAP7_75t_SL g467 ( 
.A(n_424),
.B(n_415),
.Y(n_467)
);

AOI21xp5_ASAP7_75t_L g479 ( 
.A1(n_425),
.A2(n_436),
.B(n_416),
.Y(n_479)
);

OAI22xp5_ASAP7_75t_L g460 ( 
.A1(n_427),
.A2(n_438),
.B1(n_412),
.B2(n_410),
.Y(n_460)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_428),
.Y(n_463)
);

OAI22xp5_ASAP7_75t_SL g432 ( 
.A1(n_388),
.A2(n_376),
.B1(n_351),
.B2(n_379),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_L g455 ( 
.A(n_432),
.B(n_449),
.Y(n_455)
);

AOI22xp5_ASAP7_75t_L g438 ( 
.A1(n_393),
.A2(n_353),
.B1(n_374),
.B2(n_381),
.Y(n_438)
);

AO22x1_ASAP7_75t_SL g439 ( 
.A1(n_403),
.A2(n_380),
.B1(n_372),
.B2(n_353),
.Y(n_439)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_439),
.Y(n_464)
);

MAJIxp5_ASAP7_75t_L g440 ( 
.A(n_405),
.B(n_371),
.C(n_355),
.Y(n_440)
);

MAJIxp5_ASAP7_75t_L g457 ( 
.A(n_440),
.B(n_447),
.C(n_450),
.Y(n_457)
);

CKINVDCx20_ASAP7_75t_R g442 ( 
.A(n_389),
.Y(n_442)
);

NOR2xp33_ASAP7_75t_L g461 ( 
.A(n_442),
.B(n_372),
.Y(n_461)
);

MAJIxp5_ASAP7_75t_L g447 ( 
.A(n_399),
.B(n_346),
.C(n_375),
.Y(n_447)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_448),
.Y(n_459)
);

OAI22xp5_ASAP7_75t_SL g449 ( 
.A1(n_397),
.A2(n_369),
.B1(n_359),
.B2(n_367),
.Y(n_449)
);

MAJIxp5_ASAP7_75t_L g450 ( 
.A(n_396),
.B(n_369),
.C(n_357),
.Y(n_450)
);

INVxp67_ASAP7_75t_SL g456 ( 
.A(n_443),
.Y(n_456)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_456),
.Y(n_484)
);

MAJIxp5_ASAP7_75t_L g458 ( 
.A(n_423),
.B(n_421),
.C(n_395),
.Y(n_458)
);

MAJIxp5_ASAP7_75t_L g483 ( 
.A(n_458),
.B(n_466),
.C(n_474),
.Y(n_483)
);

AOI22xp5_ASAP7_75t_L g491 ( 
.A1(n_460),
.A2(n_445),
.B1(n_454),
.B2(n_431),
.Y(n_491)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_461),
.Y(n_487)
);

XOR2xp5_ASAP7_75t_L g500 ( 
.A(n_462),
.B(n_465),
.Y(n_500)
);

XOR2xp5_ASAP7_75t_L g465 ( 
.A(n_447),
.B(n_398),
.Y(n_465)
);

MAJIxp5_ASAP7_75t_L g466 ( 
.A(n_440),
.B(n_429),
.C(n_450),
.Y(n_466)
);

NOR2xp33_ASAP7_75t_SL g501 ( 
.A(n_467),
.B(n_453),
.Y(n_501)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_443),
.Y(n_468)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_468),
.Y(n_499)
);

OAI22xp5_ASAP7_75t_L g469 ( 
.A1(n_441),
.A2(n_419),
.B1(n_418),
.B2(n_411),
.Y(n_469)
);

HB1xp67_ASAP7_75t_L g494 ( 
.A(n_469),
.Y(n_494)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_434),
.Y(n_470)
);

OAI22xp5_ASAP7_75t_L g502 ( 
.A1(n_470),
.A2(n_471),
.B1(n_472),
.B2(n_452),
.Y(n_502)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_434),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_433),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_L g473 ( 
.A(n_448),
.B(n_413),
.Y(n_473)
);

CKINVDCx20_ASAP7_75t_R g496 ( 
.A(n_473),
.Y(n_496)
);

MAJIxp5_ASAP7_75t_L g474 ( 
.A(n_429),
.B(n_394),
.C(n_406),
.Y(n_474)
);

XNOR2xp5_ASAP7_75t_L g475 ( 
.A(n_432),
.B(n_404),
.Y(n_475)
);

XNOR2xp5_ASAP7_75t_L g493 ( 
.A(n_475),
.B(n_476),
.Y(n_493)
);

XOR2xp5_ASAP7_75t_L g476 ( 
.A(n_444),
.B(n_408),
.Y(n_476)
);

XOR2xp5_ASAP7_75t_L g477 ( 
.A(n_444),
.B(n_387),
.Y(n_477)
);

MAJIxp5_ASAP7_75t_L g486 ( 
.A(n_477),
.B(n_481),
.C(n_451),
.Y(n_486)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_426),
.Y(n_478)
);

NOR2xp33_ASAP7_75t_L g495 ( 
.A(n_478),
.B(n_480),
.Y(n_495)
);

AOI21xp5_ASAP7_75t_L g482 ( 
.A1(n_479),
.A2(n_425),
.B(n_438),
.Y(n_482)
);

CKINVDCx14_ASAP7_75t_R g480 ( 
.A(n_430),
.Y(n_480)
);

MAJIxp5_ASAP7_75t_L g481 ( 
.A(n_425),
.B(n_414),
.C(n_400),
.Y(n_481)
);

A2O1A1Ixp33_ASAP7_75t_SL g506 ( 
.A1(n_482),
.A2(n_479),
.B(n_463),
.C(n_464),
.Y(n_506)
);

OAI22xp5_ASAP7_75t_SL g485 ( 
.A1(n_455),
.A2(n_454),
.B1(n_431),
.B2(n_430),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_L g512 ( 
.A(n_485),
.B(n_488),
.Y(n_512)
);

XNOR2xp5_ASAP7_75t_L g509 ( 
.A(n_486),
.B(n_477),
.Y(n_509)
);

MAJIxp5_ASAP7_75t_L g488 ( 
.A(n_466),
.B(n_457),
.C(n_465),
.Y(n_488)
);

MAJIxp5_ASAP7_75t_L g489 ( 
.A(n_457),
.B(n_437),
.C(n_439),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_L g514 ( 
.A(n_489),
.B(n_490),
.Y(n_514)
);

MAJIxp5_ASAP7_75t_L g490 ( 
.A(n_462),
.B(n_439),
.C(n_451),
.Y(n_490)
);

OAI22xp5_ASAP7_75t_SL g507 ( 
.A1(n_491),
.A2(n_498),
.B1(n_464),
.B2(n_471),
.Y(n_507)
);

MAJIxp5_ASAP7_75t_L g492 ( 
.A(n_474),
.B(n_449),
.C(n_435),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_L g518 ( 
.A(n_492),
.B(n_497),
.Y(n_518)
);

OAI22xp5_ASAP7_75t_SL g497 ( 
.A1(n_455),
.A2(n_431),
.B1(n_427),
.B2(n_428),
.Y(n_497)
);

AOI22xp5_ASAP7_75t_L g498 ( 
.A1(n_459),
.A2(n_453),
.B1(n_452),
.B2(n_446),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_SL g516 ( 
.A(n_501),
.B(n_435),
.Y(n_516)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_502),
.Y(n_508)
);

AOI21xp33_ASAP7_75t_L g503 ( 
.A1(n_463),
.A2(n_446),
.B(n_426),
.Y(n_503)
);

MAJIxp5_ASAP7_75t_SL g505 ( 
.A(n_503),
.B(n_473),
.C(n_470),
.Y(n_505)
);

MAJIxp5_ASAP7_75t_L g504 ( 
.A(n_488),
.B(n_481),
.C(n_458),
.Y(n_504)
);

MAJIxp5_ASAP7_75t_L g536 ( 
.A(n_504),
.B(n_521),
.C(n_413),
.Y(n_536)
);

AOI21xp5_ASAP7_75t_L g533 ( 
.A1(n_505),
.A2(n_482),
.B(n_499),
.Y(n_533)
);

OR2x2_ASAP7_75t_L g534 ( 
.A(n_506),
.B(n_500),
.Y(n_534)
);

AOI22xp5_ASAP7_75t_SL g531 ( 
.A1(n_507),
.A2(n_485),
.B1(n_490),
.B2(n_496),
.Y(n_531)
);

XNOR2xp5_ASAP7_75t_L g532 ( 
.A(n_509),
.B(n_520),
.Y(n_532)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_495),
.Y(n_510)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_510),
.Y(n_523)
);

CKINVDCx20_ASAP7_75t_R g511 ( 
.A(n_498),
.Y(n_511)
);

AOI22xp5_ASAP7_75t_L g530 ( 
.A1(n_511),
.A2(n_515),
.B1(n_517),
.B2(n_497),
.Y(n_530)
);

NOR2xp33_ASAP7_75t_L g513 ( 
.A(n_486),
.B(n_390),
.Y(n_513)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_513),
.Y(n_525)
);

OAI22xp5_ASAP7_75t_SL g515 ( 
.A1(n_494),
.A2(n_475),
.B1(n_476),
.B2(n_472),
.Y(n_515)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_516),
.Y(n_527)
);

OAI22xp5_ASAP7_75t_SL g517 ( 
.A1(n_491),
.A2(n_422),
.B1(n_417),
.B2(n_413),
.Y(n_517)
);

INVx13_ASAP7_75t_L g519 ( 
.A(n_484),
.Y(n_519)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_519),
.Y(n_528)
);

XNOR2xp5_ASAP7_75t_L g520 ( 
.A(n_493),
.B(n_381),
.Y(n_520)
);

XOR2xp5_ASAP7_75t_L g521 ( 
.A(n_493),
.B(n_357),
.Y(n_521)
);

BUFx24_ASAP7_75t_SL g522 ( 
.A(n_512),
.Y(n_522)
);

NOR2xp33_ASAP7_75t_L g537 ( 
.A(n_522),
.B(n_529),
.Y(n_537)
);

INVxp67_ASAP7_75t_L g524 ( 
.A(n_518),
.Y(n_524)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_524),
.Y(n_538)
);

OAI21xp5_ASAP7_75t_SL g526 ( 
.A1(n_514),
.A2(n_483),
.B(n_489),
.Y(n_526)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_526),
.Y(n_544)
);

OAI21xp5_ASAP7_75t_SL g529 ( 
.A1(n_504),
.A2(n_483),
.B(n_492),
.Y(n_529)
);

XNOR2xp5_ASAP7_75t_L g542 ( 
.A(n_530),
.B(n_531),
.Y(n_542)
);

OAI21x1_ASAP7_75t_SL g547 ( 
.A1(n_533),
.A2(n_534),
.B(n_535),
.Y(n_547)
);

OAI21x1_ASAP7_75t_SL g535 ( 
.A1(n_508),
.A2(n_487),
.B(n_500),
.Y(n_535)
);

NOR2xp33_ASAP7_75t_L g540 ( 
.A(n_536),
.B(n_520),
.Y(n_540)
);

NOR2x1_ASAP7_75t_L g539 ( 
.A(n_527),
.B(n_507),
.Y(n_539)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_539),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_SL g550 ( 
.A(n_540),
.B(n_545),
.Y(n_550)
);

MAJIxp5_ASAP7_75t_L g541 ( 
.A(n_532),
.B(n_509),
.C(n_521),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_L g549 ( 
.A(n_541),
.B(n_543),
.Y(n_549)
);

AOI22xp5_ASAP7_75t_L g543 ( 
.A1(n_524),
.A2(n_515),
.B1(n_517),
.B2(n_506),
.Y(n_543)
);

INVx2_ASAP7_75t_L g545 ( 
.A(n_525),
.Y(n_545)
);

OAI221xp5_ASAP7_75t_L g546 ( 
.A1(n_523),
.A2(n_519),
.B1(n_506),
.B2(n_389),
.C(n_367),
.Y(n_546)
);

OAI21xp5_ASAP7_75t_L g553 ( 
.A1(n_546),
.A2(n_534),
.B(n_531),
.Y(n_553)
);

NOR2xp33_ASAP7_75t_SL g551 ( 
.A(n_537),
.B(n_528),
.Y(n_551)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_551),
.Y(n_555)
);

XOR2xp5_ASAP7_75t_L g552 ( 
.A(n_541),
.B(n_532),
.Y(n_552)
);

NOR2xp33_ASAP7_75t_SL g557 ( 
.A(n_552),
.B(n_542),
.Y(n_557)
);

OAI22xp5_ASAP7_75t_SL g556 ( 
.A1(n_553),
.A2(n_543),
.B1(n_536),
.B2(n_547),
.Y(n_556)
);

A2O1A1Ixp33_ASAP7_75t_L g554 ( 
.A1(n_548),
.A2(n_544),
.B(n_538),
.C(n_506),
.Y(n_554)
);

AOI21xp5_ASAP7_75t_L g559 ( 
.A1(n_554),
.A2(n_539),
.B(n_542),
.Y(n_559)
);

NOR2xp33_ASAP7_75t_L g558 ( 
.A(n_556),
.B(n_557),
.Y(n_558)
);

AOI322xp5_ASAP7_75t_L g560 ( 
.A1(n_559),
.A2(n_550),
.A3(n_554),
.B1(n_555),
.B2(n_549),
.C1(n_389),
.C2(n_552),
.Y(n_560)
);

MAJIxp5_ASAP7_75t_L g561 ( 
.A(n_560),
.B(n_558),
.C(n_10),
.Y(n_561)
);

OAI21xp5_ASAP7_75t_L g562 ( 
.A1(n_561),
.A2(n_9),
.B(n_11),
.Y(n_562)
);

AOI221xp5_ASAP7_75t_L g563 ( 
.A1(n_562),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.C(n_197),
.Y(n_563)
);

MAJIxp5_ASAP7_75t_L g564 ( 
.A(n_563),
.B(n_11),
.C(n_12),
.Y(n_564)
);

NOR2xp33_ASAP7_75t_L g565 ( 
.A(n_564),
.B(n_11),
.Y(n_565)
);


endmodule