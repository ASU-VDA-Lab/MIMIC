module fake_jpeg_30013_n_351 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_351);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_351;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_137;
wire n_74;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_122;
wire n_75;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_347;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVxp67_ASAP7_75t_L g15 ( 
.A(n_2),
.Y(n_15)
);

INVx3_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

INVx3_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_12),
.Y(n_26)
);

INVx5_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

BUFx16f_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_3),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_8),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_9),
.Y(n_36)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_3),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_7),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_8),
.Y(n_39)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_17),
.Y(n_40)
);

INVx11_ASAP7_75t_L g84 ( 
.A(n_40),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_17),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_41),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_17),
.Y(n_42)
);

INVx6_ASAP7_75t_L g75 ( 
.A(n_42),
.Y(n_75)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_17),
.Y(n_43)
);

INVx5_ASAP7_75t_L g61 ( 
.A(n_43),
.Y(n_61)
);

HB1xp67_ASAP7_75t_L g44 ( 
.A(n_32),
.Y(n_44)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_44),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_22),
.Y(n_45)
);

INVx6_ASAP7_75t_L g85 ( 
.A(n_45),
.Y(n_85)
);

INVx13_ASAP7_75t_L g46 ( 
.A(n_32),
.Y(n_46)
);

BUFx24_ASAP7_75t_L g62 ( 
.A(n_46),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_22),
.Y(n_47)
);

INVx5_ASAP7_75t_L g63 ( 
.A(n_47),
.Y(n_63)
);

BUFx5_ASAP7_75t_L g48 ( 
.A(n_32),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g74 ( 
.A(n_48),
.Y(n_74)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_27),
.Y(n_49)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_49),
.Y(n_92)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_27),
.Y(n_50)
);

BUFx5_ASAP7_75t_L g66 ( 
.A(n_50),
.Y(n_66)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_24),
.Y(n_51)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_51),
.Y(n_77)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_22),
.Y(n_52)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_52),
.Y(n_81)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_16),
.Y(n_53)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_53),
.Y(n_64)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_32),
.Y(n_54)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_54),
.Y(n_91)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_32),
.Y(n_55)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_55),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_26),
.B(n_13),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_56),
.B(n_57),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_26),
.B(n_13),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_22),
.Y(n_58)
);

BUFx12f_ASAP7_75t_L g94 ( 
.A(n_58),
.Y(n_94)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_16),
.Y(n_59)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_59),
.Y(n_72)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_16),
.Y(n_60)
);

INVx4_ASAP7_75t_SL g80 ( 
.A(n_60),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_51),
.A2(n_15),
.B1(n_25),
.B2(n_38),
.Y(n_67)
);

AND2x2_ASAP7_75t_L g107 ( 
.A(n_67),
.B(n_70),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_53),
.A2(n_37),
.B1(n_19),
.B2(n_27),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_68),
.A2(n_88),
.B1(n_21),
.B2(n_35),
.Y(n_122)
);

CKINVDCx16_ASAP7_75t_R g69 ( 
.A(n_46),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_69),
.B(n_73),
.Y(n_135)
);

AND2x2_ASAP7_75t_L g70 ( 
.A(n_59),
.B(n_19),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_41),
.B(n_31),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_71),
.B(n_78),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_49),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_41),
.B(n_31),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_60),
.A2(n_25),
.B1(n_34),
.B2(n_38),
.Y(n_79)
);

AND2x2_ASAP7_75t_L g112 ( 
.A(n_79),
.B(n_99),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_54),
.B(n_33),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_83),
.B(n_89),
.Y(n_114)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_55),
.Y(n_86)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_86),
.Y(n_113)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_40),
.Y(n_87)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_87),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_40),
.A2(n_19),
.B1(n_37),
.B2(n_28),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_54),
.B(n_24),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_42),
.B(n_36),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_90),
.B(n_93),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_54),
.B(n_33),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_48),
.B(n_39),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_95),
.B(n_98),
.Y(n_126)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_43),
.Y(n_96)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_96),
.Y(n_121)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_42),
.Y(n_97)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_97),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_46),
.B(n_39),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_45),
.B(n_18),
.Y(n_99)
);

A2O1A1Ixp33_ASAP7_75t_L g100 ( 
.A1(n_50),
.A2(n_25),
.B(n_20),
.C(n_18),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_100),
.B(n_102),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_43),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_62),
.Y(n_103)
);

CKINVDCx14_ASAP7_75t_R g143 ( 
.A(n_103),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_70),
.A2(n_20),
.B1(n_30),
.B2(n_37),
.Y(n_104)
);

AND2x2_ASAP7_75t_L g166 ( 
.A(n_104),
.B(n_122),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_76),
.Y(n_106)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_106),
.Y(n_144)
);

INVx8_ASAP7_75t_L g108 ( 
.A(n_81),
.Y(n_108)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_108),
.Y(n_148)
);

CKINVDCx16_ASAP7_75t_R g109 ( 
.A(n_62),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_109),
.B(n_127),
.Y(n_149)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_86),
.Y(n_110)
);

HB1xp67_ASAP7_75t_L g151 ( 
.A(n_110),
.Y(n_151)
);

INVx4_ASAP7_75t_L g111 ( 
.A(n_101),
.Y(n_111)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_111),
.Y(n_150)
);

INVx6_ASAP7_75t_L g115 ( 
.A(n_76),
.Y(n_115)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_115),
.Y(n_156)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_62),
.Y(n_120)
);

CKINVDCx14_ASAP7_75t_R g152 ( 
.A(n_120),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_71),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_123),
.B(n_124),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_78),
.Y(n_124)
);

OAI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_100),
.A2(n_58),
.B1(n_47),
.B2(n_45),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_125),
.A2(n_138),
.B1(n_80),
.B2(n_104),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_99),
.Y(n_127)
);

INVx3_ASAP7_75t_L g128 ( 
.A(n_94),
.Y(n_128)
);

INVxp67_ASAP7_75t_L g158 ( 
.A(n_128),
.Y(n_158)
);

AO22x1_ASAP7_75t_SL g129 ( 
.A1(n_64),
.A2(n_58),
.B1(n_47),
.B2(n_52),
.Y(n_129)
);

AO22x1_ASAP7_75t_SL g171 ( 
.A1(n_129),
.A2(n_131),
.B1(n_63),
.B2(n_61),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_82),
.B(n_36),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_SL g147 ( 
.A(n_130),
.B(n_126),
.Y(n_147)
);

AO22x2_ASAP7_75t_L g131 ( 
.A1(n_75),
.A2(n_52),
.B1(n_28),
.B2(n_29),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_77),
.Y(n_132)
);

CKINVDCx16_ASAP7_75t_R g162 ( 
.A(n_132),
.Y(n_162)
);

INVx3_ASAP7_75t_L g133 ( 
.A(n_94),
.Y(n_133)
);

INVxp67_ASAP7_75t_L g169 ( 
.A(n_133),
.Y(n_169)
);

INVx3_ASAP7_75t_L g134 ( 
.A(n_94),
.Y(n_134)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_134),
.Y(n_161)
);

OA21x2_ASAP7_75t_L g136 ( 
.A1(n_67),
.A2(n_35),
.B(n_23),
.Y(n_136)
);

AND2x2_ASAP7_75t_L g168 ( 
.A(n_136),
.B(n_140),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_75),
.Y(n_137)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_137),
.Y(n_165)
);

AOI22xp33_ASAP7_75t_SL g138 ( 
.A1(n_80),
.A2(n_30),
.B1(n_29),
.B2(n_28),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_85),
.Y(n_139)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_139),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_70),
.A2(n_34),
.B1(n_35),
.B2(n_23),
.Y(n_140)
);

OAI32xp33_ASAP7_75t_L g141 ( 
.A1(n_105),
.A2(n_116),
.A3(n_112),
.B1(n_107),
.B2(n_119),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_141),
.B(n_147),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_L g142 ( 
.A1(n_107),
.A2(n_79),
.B(n_65),
.Y(n_142)
);

OR2x2_ASAP7_75t_L g184 ( 
.A(n_142),
.B(n_164),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_112),
.A2(n_97),
.B1(n_64),
.B2(n_72),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_145),
.A2(n_146),
.B1(n_154),
.B2(n_171),
.Y(n_180)
);

FAx1_ASAP7_75t_SL g153 ( 
.A(n_112),
.B(n_72),
.CI(n_101),
.CON(n_153),
.SN(n_153)
);

NOR2xp33_ASAP7_75t_SL g202 ( 
.A(n_153),
.B(n_157),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_107),
.A2(n_136),
.B1(n_140),
.B2(n_131),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_136),
.B(n_85),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_155),
.B(n_157),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_114),
.B(n_21),
.Y(n_157)
);

AOI21xp5_ASAP7_75t_L g159 ( 
.A1(n_103),
.A2(n_92),
.B(n_74),
.Y(n_159)
);

OA21x2_ASAP7_75t_L g203 ( 
.A1(n_159),
.A2(n_0),
.B(n_2),
.Y(n_203)
);

OAI32xp33_ASAP7_75t_L g160 ( 
.A1(n_131),
.A2(n_81),
.A3(n_21),
.B1(n_23),
.B2(n_91),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_160),
.B(n_174),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_L g164 ( 
.A1(n_135),
.A2(n_91),
.B(n_84),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_117),
.B(n_63),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_170),
.B(n_0),
.Y(n_204)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_118),
.Y(n_172)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_172),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_121),
.B(n_92),
.C(n_74),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_173),
.B(n_134),
.C(n_133),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_111),
.B(n_120),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_131),
.A2(n_84),
.B1(n_61),
.B2(n_29),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_175),
.A2(n_66),
.B1(n_28),
.B2(n_3),
.Y(n_194)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_118),
.Y(n_176)
);

CKINVDCx16_ASAP7_75t_R g195 ( 
.A(n_176),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_110),
.B(n_113),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_177),
.B(n_128),
.Y(n_186)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_113),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_178),
.B(n_108),
.Y(n_179)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_179),
.Y(n_223)
);

INVx5_ASAP7_75t_L g181 ( 
.A(n_144),
.Y(n_181)
);

BUFx2_ASAP7_75t_L g236 ( 
.A(n_181),
.Y(n_236)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_182),
.B(n_156),
.Y(n_240)
);

CKINVDCx14_ASAP7_75t_R g238 ( 
.A(n_186),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_155),
.A2(n_129),
.B1(n_139),
.B2(n_137),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_187),
.A2(n_197),
.B1(n_198),
.B2(n_200),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_149),
.B(n_29),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_188),
.B(n_191),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_168),
.B(n_129),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_189),
.B(n_196),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_163),
.B(n_115),
.C(n_106),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_190),
.B(n_192),
.C(n_207),
.Y(n_217)
);

INVxp33_ASAP7_75t_L g191 ( 
.A(n_159),
.Y(n_191)
);

MAJx2_ASAP7_75t_L g192 ( 
.A(n_168),
.B(n_66),
.C(n_12),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_194),
.A2(n_206),
.B1(n_184),
.B2(n_213),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_168),
.B(n_12),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_166),
.A2(n_142),
.B1(n_154),
.B2(n_141),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g198 ( 
.A1(n_166),
.A2(n_11),
.B1(n_10),
.B2(n_3),
.Y(n_198)
);

INVx11_ASAP7_75t_L g199 ( 
.A(n_158),
.Y(n_199)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_199),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_L g200 ( 
.A1(n_166),
.A2(n_10),
.B1(n_11),
.B2(n_5),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_170),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_201),
.B(n_202),
.Y(n_222)
);

AND2x2_ASAP7_75t_L g239 ( 
.A(n_203),
.B(n_144),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_SL g242 ( 
.A(n_204),
.B(n_205),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_153),
.B(n_0),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_L g206 ( 
.A1(n_171),
.A2(n_160),
.B1(n_175),
.B2(n_153),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_145),
.B(n_11),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_147),
.B(n_0),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_208),
.B(n_209),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_162),
.Y(n_209)
);

AOI22xp33_ASAP7_75t_SL g210 ( 
.A1(n_143),
.A2(n_2),
.B1(n_5),
.B2(n_6),
.Y(n_210)
);

OAI22x1_ASAP7_75t_L g241 ( 
.A1(n_210),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_241)
);

INVxp67_ASAP7_75t_L g211 ( 
.A(n_164),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_211),
.B(n_213),
.Y(n_233)
);

OR2x2_ASAP7_75t_L g213 ( 
.A(n_171),
.B(n_5),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_SL g214 ( 
.A(n_173),
.B(n_5),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_SL g219 ( 
.A(n_214),
.B(n_6),
.Y(n_219)
);

INVx13_ASAP7_75t_L g215 ( 
.A(n_152),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_215),
.Y(n_224)
);

O2A1O1Ixp33_ASAP7_75t_SL g216 ( 
.A1(n_183),
.A2(n_158),
.B(n_169),
.C(n_148),
.Y(n_216)
);

AOI21xp5_ASAP7_75t_L g264 ( 
.A1(n_216),
.A2(n_179),
.B(n_185),
.Y(n_264)
);

AOI21xp5_ASAP7_75t_L g218 ( 
.A1(n_184),
.A2(n_148),
.B(n_169),
.Y(n_218)
);

OAI21xp5_ASAP7_75t_SL g267 ( 
.A1(n_218),
.A2(n_229),
.B(n_235),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_SL g249 ( 
.A(n_219),
.B(n_231),
.Y(n_249)
);

OAI21xp5_ASAP7_75t_L g221 ( 
.A1(n_184),
.A2(n_150),
.B(n_151),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_L g259 ( 
.A1(n_221),
.A2(n_203),
.B(n_214),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_197),
.B(n_150),
.C(n_178),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_225),
.B(n_240),
.C(n_182),
.Y(n_248)
);

AOI21xp5_ASAP7_75t_SL g229 ( 
.A1(n_203),
.A2(n_161),
.B(n_172),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_SL g231 ( 
.A(n_193),
.B(n_161),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_209),
.B(n_176),
.Y(n_232)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_232),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_234),
.A2(n_198),
.B1(n_187),
.B2(n_180),
.Y(n_262)
);

AOI21xp5_ASAP7_75t_L g235 ( 
.A1(n_206),
.A2(n_167),
.B(n_165),
.Y(n_235)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_212),
.Y(n_237)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_237),
.Y(n_265)
);

AND2x2_ASAP7_75t_L g260 ( 
.A(n_239),
.B(n_194),
.Y(n_260)
);

OAI22x1_ASAP7_75t_L g247 ( 
.A1(n_241),
.A2(n_203),
.B1(n_192),
.B2(n_200),
.Y(n_247)
);

BUFx24_ASAP7_75t_SL g243 ( 
.A(n_193),
.Y(n_243)
);

BUFx24_ASAP7_75t_SL g251 ( 
.A(n_243),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_SL g244 ( 
.A(n_196),
.B(n_156),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_244),
.B(n_202),
.Y(n_250)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_237),
.Y(n_245)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_245),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_236),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_246),
.B(n_253),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_247),
.A2(n_216),
.B1(n_233),
.B2(n_220),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_SL g284 ( 
.A(n_248),
.B(n_242),
.Y(n_284)
);

CKINVDCx14_ASAP7_75t_R g270 ( 
.A(n_250),
.Y(n_270)
);

INVxp67_ASAP7_75t_L g252 ( 
.A(n_218),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_252),
.B(n_256),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_231),
.B(n_190),
.Y(n_253)
);

AOI21x1_ASAP7_75t_L g254 ( 
.A1(n_221),
.A2(n_189),
.B(n_205),
.Y(n_254)
);

AOI21xp5_ASAP7_75t_L g273 ( 
.A1(n_254),
.A2(n_259),
.B(n_260),
.Y(n_273)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_223),
.Y(n_255)
);

INVx1_ASAP7_75t_SL g288 ( 
.A(n_255),
.Y(n_288)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_223),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_240),
.B(n_201),
.C(n_180),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_257),
.B(n_217),
.C(n_228),
.Y(n_274)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_227),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_SL g280 ( 
.A(n_258),
.B(n_264),
.Y(n_280)
);

OA21x2_ASAP7_75t_L g261 ( 
.A1(n_233),
.A2(n_213),
.B(n_185),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_261),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_262),
.A2(n_266),
.B1(n_230),
.B2(n_225),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_235),
.A2(n_234),
.B1(n_239),
.B2(n_216),
.Y(n_266)
);

AOI21xp5_ASAP7_75t_L g268 ( 
.A1(n_239),
.A2(n_215),
.B(n_192),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_L g289 ( 
.A1(n_268),
.A2(n_241),
.B1(n_204),
.B2(n_219),
.Y(n_289)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_227),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_SL g286 ( 
.A(n_269),
.B(n_224),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g301 ( 
.A1(n_271),
.A2(n_281),
.B1(n_282),
.B2(n_285),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_274),
.B(n_278),
.C(n_284),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_L g303 ( 
.A1(n_275),
.A2(n_279),
.B1(n_249),
.B2(n_263),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_248),
.B(n_217),
.C(n_222),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_260),
.A2(n_222),
.B1(n_220),
.B2(n_238),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_262),
.A2(n_230),
.B1(n_228),
.B2(n_229),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_266),
.A2(n_229),
.B1(n_242),
.B2(n_226),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_247),
.A2(n_226),
.B1(n_224),
.B2(n_241),
.Y(n_285)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_286),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_257),
.B(n_195),
.C(n_244),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_287),
.B(n_252),
.C(n_259),
.Y(n_302)
);

AOI21xp5_ASAP7_75t_L g290 ( 
.A1(n_289),
.A2(n_260),
.B(n_264),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g312 ( 
.A1(n_290),
.A2(n_303),
.B1(n_289),
.B2(n_282),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_286),
.B(n_256),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_291),
.B(n_295),
.Y(n_317)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_274),
.B(n_254),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g314 ( 
.A(n_292),
.B(n_293),
.Y(n_314)
);

XOR2xp5_ASAP7_75t_L g293 ( 
.A(n_278),
.B(n_268),
.Y(n_293)
);

XOR2xp5_ASAP7_75t_L g311 ( 
.A(n_293),
.B(n_294),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_SL g294 ( 
.A(n_284),
.B(n_250),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_SL g295 ( 
.A(n_270),
.B(n_251),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_288),
.B(n_255),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_296),
.B(n_298),
.Y(n_318)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_288),
.Y(n_298)
);

XOR2xp5_ASAP7_75t_L g299 ( 
.A(n_287),
.B(n_273),
.Y(n_299)
);

XOR2xp5_ASAP7_75t_L g313 ( 
.A(n_299),
.B(n_272),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_302),
.B(n_273),
.C(n_277),
.Y(n_308)
);

OAI21xp5_ASAP7_75t_L g304 ( 
.A1(n_280),
.A2(n_261),
.B(n_267),
.Y(n_304)
);

AOI21xp5_ASAP7_75t_L g309 ( 
.A1(n_304),
.A2(n_267),
.B(n_275),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_276),
.B(n_272),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_305),
.B(n_276),
.Y(n_306)
);

OR2x2_ASAP7_75t_L g325 ( 
.A(n_306),
.B(n_291),
.Y(n_325)
);

AOI22xp5_ASAP7_75t_SL g307 ( 
.A1(n_297),
.A2(n_285),
.B1(n_271),
.B2(n_281),
.Y(n_307)
);

XOR2xp5_ASAP7_75t_L g324 ( 
.A(n_307),
.B(n_309),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_308),
.B(n_316),
.C(n_294),
.Y(n_327)
);

AOI21xp5_ASAP7_75t_L g310 ( 
.A1(n_304),
.A2(n_280),
.B(n_279),
.Y(n_310)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_310),
.Y(n_320)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_312),
.Y(n_322)
);

XNOR2xp5_ASAP7_75t_L g321 ( 
.A(n_313),
.B(n_314),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_290),
.B(n_261),
.Y(n_315)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_315),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_300),
.B(n_269),
.C(n_258),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_SL g319 ( 
.A(n_317),
.B(n_300),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_319),
.B(n_325),
.Y(n_336)
);

XNOR2xp5_ASAP7_75t_L g326 ( 
.A(n_316),
.B(n_302),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_SL g330 ( 
.A(n_326),
.B(n_314),
.Y(n_330)
);

AOI21xp5_ASAP7_75t_L g335 ( 
.A1(n_327),
.A2(n_328),
.B(n_311),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_313),
.B(n_292),
.C(n_299),
.Y(n_328)
);

OAI21xp5_ASAP7_75t_SL g329 ( 
.A1(n_320),
.A2(n_308),
.B(n_318),
.Y(n_329)
);

AOI21xp5_ASAP7_75t_L g340 ( 
.A1(n_329),
.A2(n_333),
.B(n_212),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_SL g339 ( 
.A(n_330),
.B(n_334),
.Y(n_339)
);

AOI22xp5_ASAP7_75t_L g331 ( 
.A1(n_322),
.A2(n_283),
.B1(n_245),
.B2(n_307),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_331),
.B(n_332),
.Y(n_341)
);

AOI22xp5_ASAP7_75t_L g332 ( 
.A1(n_323),
.A2(n_301),
.B1(n_311),
.B2(n_305),
.Y(n_332)
);

OAI21xp5_ASAP7_75t_SL g333 ( 
.A1(n_327),
.A2(n_296),
.B(n_283),
.Y(n_333)
);

BUFx24_ASAP7_75t_SL g334 ( 
.A(n_324),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_SL g342 ( 
.A(n_335),
.B(n_207),
.Y(n_342)
);

AOI322xp5_ASAP7_75t_L g337 ( 
.A1(n_336),
.A2(n_325),
.A3(n_324),
.B1(n_332),
.B2(n_265),
.C1(n_301),
.C2(n_328),
.Y(n_337)
);

AOI21xp33_ASAP7_75t_L g343 ( 
.A1(n_337),
.A2(n_215),
.B(n_236),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_335),
.B(n_321),
.C(n_195),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_338),
.B(n_340),
.Y(n_344)
);

OAI21xp5_ASAP7_75t_L g345 ( 
.A1(n_342),
.A2(n_199),
.B(n_167),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_343),
.B(n_236),
.Y(n_346)
);

INVxp67_ASAP7_75t_L g347 ( 
.A(n_345),
.Y(n_347)
);

MAJx2_ASAP7_75t_L g348 ( 
.A(n_346),
.B(n_344),
.C(n_341),
.Y(n_348)
);

A2O1A1O1Ixp25_ASAP7_75t_L g349 ( 
.A1(n_348),
.A2(n_339),
.B(n_347),
.C(n_165),
.D(n_181),
.Y(n_349)
);

NOR3xp33_ASAP7_75t_L g350 ( 
.A(n_349),
.B(n_6),
.C(n_7),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_350),
.B(n_9),
.Y(n_351)
);


endmodule