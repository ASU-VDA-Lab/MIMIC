module fake_jpeg_28272_n_130 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_130);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_130;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

BUFx12_ASAP7_75t_L g13 ( 
.A(n_3),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_0),
.Y(n_14)
);

BUFx12f_ASAP7_75t_L g15 ( 
.A(n_5),
.Y(n_15)
);

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

INVx6_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_6),
.Y(n_20)
);

INVx11_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

INVx11_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

BUFx24_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_1),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_12),
.Y(n_27)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

INVx5_ASAP7_75t_SL g45 ( 
.A(n_28),
.Y(n_45)
);

CKINVDCx16_ASAP7_75t_R g29 ( 
.A(n_23),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_29),
.B(n_36),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_23),
.Y(n_30)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_30),
.Y(n_55)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_20),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_SL g48 ( 
.A(n_31),
.B(n_33),
.Y(n_48)
);

INVx11_ASAP7_75t_L g32 ( 
.A(n_25),
.Y(n_32)
);

INVx5_ASAP7_75t_L g49 ( 
.A(n_32),
.Y(n_49)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_20),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_23),
.B(n_0),
.Y(n_34)
);

AND2x2_ASAP7_75t_L g43 ( 
.A(n_34),
.B(n_0),
.Y(n_43)
);

INVx5_ASAP7_75t_L g35 ( 
.A(n_25),
.Y(n_35)
);

BUFx2_ASAP7_75t_L g53 ( 
.A(n_35),
.Y(n_53)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_27),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_15),
.Y(n_37)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_37),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_23),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_38),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_34),
.B(n_25),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_40),
.B(n_47),
.Y(n_67)
);

CKINVDCx14_ASAP7_75t_R g41 ( 
.A(n_31),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_41),
.B(n_43),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_SL g44 ( 
.A1(n_28),
.A2(n_17),
.B1(n_24),
.B2(n_14),
.Y(n_44)
);

INVxp67_ASAP7_75t_L g64 ( 
.A(n_44),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_37),
.B(n_25),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_33),
.B(n_27),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_SL g56 ( 
.A(n_50),
.B(n_36),
.Y(n_56)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_29),
.Y(n_51)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_51),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g52 ( 
.A1(n_35),
.A2(n_17),
.B1(n_22),
.B2(n_21),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_52),
.A2(n_16),
.B1(n_15),
.B2(n_13),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_L g54 ( 
.A1(n_32),
.A2(n_22),
.B1(n_21),
.B2(n_26),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g59 ( 
.A1(n_54),
.A2(n_14),
.B1(n_24),
.B2(n_18),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_SL g81 ( 
.A(n_56),
.B(n_66),
.Y(n_81)
);

AND2x2_ASAP7_75t_L g57 ( 
.A(n_40),
.B(n_37),
.Y(n_57)
);

OAI21xp5_ASAP7_75t_L g86 ( 
.A1(n_57),
.A2(n_69),
.B(n_64),
.Y(n_86)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_55),
.Y(n_58)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_58),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_59),
.A2(n_60),
.B1(n_61),
.B2(n_70),
.Y(n_73)
);

OAI32xp33_ASAP7_75t_L g60 ( 
.A1(n_47),
.A2(n_18),
.A3(n_19),
.B1(n_16),
.B2(n_15),
.Y(n_60)
);

AO22x2_ASAP7_75t_SL g61 ( 
.A1(n_44),
.A2(n_52),
.B1(n_42),
.B2(n_38),
.Y(n_61)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_39),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_63),
.B(n_65),
.Y(n_76)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_48),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g66 ( 
.A(n_43),
.B(n_19),
.Y(n_66)
);

NOR2xp67_ASAP7_75t_L g68 ( 
.A(n_43),
.B(n_38),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_68),
.B(n_71),
.Y(n_79)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_53),
.Y(n_71)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_46),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_72),
.A2(n_55),
.B1(n_49),
.B2(n_46),
.Y(n_78)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_60),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_74),
.B(n_83),
.Y(n_94)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_67),
.B(n_37),
.Y(n_75)
);

OAI21xp5_ASAP7_75t_SL g88 ( 
.A1(n_75),
.A2(n_80),
.B(n_57),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_67),
.B(n_51),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_77),
.B(n_82),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_78),
.A2(n_61),
.B1(n_45),
.B2(n_85),
.Y(n_90)
);

AND2x2_ASAP7_75t_L g80 ( 
.A(n_62),
.B(n_30),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_69),
.B(n_42),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_58),
.Y(n_83)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_61),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_85),
.B(n_30),
.Y(n_93)
);

OAI21xp5_ASAP7_75t_L g89 ( 
.A1(n_86),
.A2(n_64),
.B(n_57),
.Y(n_89)
);

AOI21xp5_ASAP7_75t_L g106 ( 
.A1(n_88),
.A2(n_3),
.B(n_4),
.Y(n_106)
);

XNOR2xp5_ASAP7_75t_SL g104 ( 
.A(n_89),
.B(n_98),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_90),
.A2(n_91),
.B1(n_92),
.B2(n_75),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_74),
.A2(n_70),
.B1(n_45),
.B2(n_72),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_73),
.A2(n_45),
.B1(n_49),
.B2(n_16),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_93),
.B(n_95),
.Y(n_99)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_82),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_77),
.B(n_16),
.C(n_13),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_96),
.B(n_84),
.C(n_76),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_75),
.B(n_2),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_97),
.B(n_80),
.Y(n_102)
);

A2O1A1O1Ixp25_ASAP7_75t_L g98 ( 
.A1(n_86),
.A2(n_13),
.B(n_53),
.C(n_4),
.D(n_2),
.Y(n_98)
);

OAI21xp5_ASAP7_75t_SL g114 ( 
.A1(n_100),
.A2(n_101),
.B(n_105),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_91),
.A2(n_79),
.B1(n_73),
.B2(n_80),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_102),
.B(n_103),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_94),
.A2(n_81),
.B1(n_53),
.B2(n_3),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_L g110 ( 
.A1(n_106),
.A2(n_97),
.B(n_89),
.Y(n_110)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_87),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_107),
.B(n_87),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_99),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_108),
.B(n_109),
.Y(n_119)
);

XOR2xp5_ASAP7_75t_L g118 ( 
.A(n_110),
.B(n_88),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_105),
.B(n_96),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_112),
.B(n_113),
.Y(n_116)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_101),
.Y(n_113)
);

NAND4xp25_ASAP7_75t_L g115 ( 
.A(n_110),
.B(n_98),
.C(n_104),
.D(n_100),
.Y(n_115)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_115),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_111),
.B(n_103),
.C(n_104),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_117),
.B(n_116),
.C(n_119),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_118),
.A2(n_114),
.B1(n_9),
.B2(n_10),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_121),
.B(n_11),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_L g122 ( 
.A1(n_116),
.A2(n_114),
.B(n_8),
.Y(n_122)
);

AO21x1_ASAP7_75t_L g124 ( 
.A1(n_122),
.A2(n_7),
.B(n_9),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_123),
.B(n_7),
.Y(n_125)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_124),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_125),
.A2(n_126),
.B1(n_120),
.B2(n_122),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_128),
.B(n_121),
.C(n_11),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_L g130 ( 
.A(n_129),
.B(n_127),
.Y(n_130)
);


endmodule