module real_jpeg_12096_n_18 (n_17, n_8, n_0, n_2, n_331, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_3, n_5, n_4, n_1, n_16, n_15, n_13, n_18);

input n_17;
input n_8;
input n_0;
input n_2;
input n_331;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;

output n_18;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

BUFx16f_ASAP7_75t_L g46 ( 
.A(n_1),
.Y(n_46)
);

BUFx12_ASAP7_75t_L g62 ( 
.A(n_2),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_3),
.A2(n_60),
.B1(n_61),
.B2(n_120),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_3),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_SL g180 ( 
.A1(n_3),
.A2(n_41),
.B1(n_43),
.B2(n_120),
.Y(n_180)
);

AOI22xp33_ASAP7_75t_SL g201 ( 
.A1(n_3),
.A2(n_55),
.B1(n_58),
.B2(n_120),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_3),
.A2(n_30),
.B1(n_36),
.B2(n_120),
.Y(n_231)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_4),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_L g49 ( 
.A1(n_5),
.A2(n_41),
.B1(n_43),
.B2(n_50),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_5),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_L g92 ( 
.A1(n_5),
.A2(n_50),
.B1(n_55),
.B2(n_58),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_L g110 ( 
.A1(n_5),
.A2(n_30),
.B1(n_36),
.B2(n_50),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g317 ( 
.A1(n_5),
.A2(n_50),
.B1(n_60),
.B2(n_61),
.Y(n_317)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_6),
.A2(n_60),
.B1(n_61),
.B2(n_66),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_6),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_6),
.A2(n_55),
.B1(n_58),
.B2(n_66),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_6),
.A2(n_41),
.B1(n_43),
.B2(n_66),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_6),
.A2(n_30),
.B1(n_36),
.B2(n_66),
.Y(n_176)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_7),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_8),
.A2(n_55),
.B1(n_58),
.B2(n_72),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_8),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_8),
.A2(n_60),
.B1(n_61),
.B2(n_72),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_L g114 ( 
.A1(n_8),
.A2(n_41),
.B1(n_43),
.B2(n_72),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g177 ( 
.A1(n_8),
.A2(n_30),
.B1(n_36),
.B2(n_72),
.Y(n_177)
);

AOI22xp33_ASAP7_75t_SL g168 ( 
.A1(n_9),
.A2(n_55),
.B1(n_58),
.B2(n_169),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_9),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_L g198 ( 
.A1(n_9),
.A2(n_60),
.B1(n_61),
.B2(n_169),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_L g222 ( 
.A1(n_9),
.A2(n_41),
.B1(n_43),
.B2(n_169),
.Y(n_222)
);

OAI22xp33_ASAP7_75t_SL g243 ( 
.A1(n_9),
.A2(n_30),
.B1(n_36),
.B2(n_169),
.Y(n_243)
);

BUFx12_ASAP7_75t_L g75 ( 
.A(n_10),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_11),
.B(n_174),
.Y(n_173)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_11),
.Y(n_187)
);

AOI21xp33_ASAP7_75t_L g195 ( 
.A1(n_11),
.A2(n_60),
.B(n_196),
.Y(n_195)
);

OAI22xp33_ASAP7_75t_L g221 ( 
.A1(n_11),
.A2(n_41),
.B1(n_43),
.B2(n_187),
.Y(n_221)
);

O2A1O1Ixp33_ASAP7_75t_L g223 ( 
.A1(n_11),
.A2(n_43),
.B(n_46),
.C(n_224),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_11),
.B(n_79),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_11),
.B(n_33),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_11),
.B(n_51),
.Y(n_248)
);

A2O1A1Ixp33_ASAP7_75t_L g257 ( 
.A1(n_11),
.A2(n_58),
.B(n_73),
.C(n_258),
.Y(n_257)
);

BUFx8_ASAP7_75t_L g57 ( 
.A(n_12),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g39 ( 
.A1(n_13),
.A2(n_40),
.B1(n_41),
.B2(n_43),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_13),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_13),
.A2(n_40),
.B1(n_55),
.B2(n_58),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_13),
.A2(n_40),
.B1(n_60),
.B2(n_61),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_13),
.A2(n_30),
.B1(n_36),
.B2(n_40),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g34 ( 
.A1(n_14),
.A2(n_30),
.B1(n_35),
.B2(n_36),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_14),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_14),
.A2(n_35),
.B1(n_41),
.B2(n_43),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_14),
.A2(n_35),
.B1(n_55),
.B2(n_58),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g326 ( 
.A1(n_14),
.A2(n_35),
.B1(n_60),
.B2(n_61),
.Y(n_326)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_15),
.A2(n_60),
.B1(n_61),
.B2(n_64),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_15),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g153 ( 
.A1(n_15),
.A2(n_55),
.B1(n_58),
.B2(n_64),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_15),
.A2(n_41),
.B1(n_43),
.B2(n_64),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_15),
.A2(n_30),
.B1(n_36),
.B2(n_64),
.Y(n_190)
);

AOI22xp33_ASAP7_75t_SL g155 ( 
.A1(n_16),
.A2(n_60),
.B1(n_61),
.B2(n_156),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_16),
.Y(n_156)
);

AOI22xp33_ASAP7_75t_SL g171 ( 
.A1(n_16),
.A2(n_55),
.B1(n_58),
.B2(n_156),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_L g229 ( 
.A1(n_16),
.A2(n_41),
.B1(n_43),
.B2(n_156),
.Y(n_229)
);

OAI22xp33_ASAP7_75t_SL g236 ( 
.A1(n_16),
.A2(n_30),
.B1(n_36),
.B2(n_156),
.Y(n_236)
);

INVx11_ASAP7_75t_L g31 ( 
.A(n_17),
.Y(n_31)
);

XOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_322),
.Y(n_18)
);

AOI21xp5_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_309),
.B(n_321),
.Y(n_19)
);

AO21x1_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_134),
.B(n_306),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_121),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_SL g22 ( 
.A(n_23),
.B(n_96),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_23),
.B(n_96),
.Y(n_307)
);

XOR2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_67),
.Y(n_23)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_24),
.B(n_82),
.C(n_94),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_28),
.B(n_52),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_25),
.A2(n_26),
.B1(n_99),
.B2(n_100),
.Y(n_98)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_37),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_27),
.A2(n_28),
.B1(n_52),
.B2(n_101),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_27),
.A2(n_28),
.B1(n_37),
.B2(n_38),
.Y(n_140)
);

CKINVDCx16_ASAP7_75t_R g27 ( 
.A(n_28),
.Y(n_27)
);

OAI21xp5_ASAP7_75t_SL g28 ( 
.A1(n_29),
.A2(n_33),
.B(n_34),
.Y(n_28)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_29),
.A2(n_33),
.B1(n_34),
.B2(n_109),
.Y(n_108)
);

CKINVDCx16_ASAP7_75t_R g145 ( 
.A(n_29),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_29),
.A2(n_33),
.B1(n_176),
.B2(n_177),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_29),
.A2(n_33),
.B1(n_176),
.B2(n_190),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_29),
.A2(n_33),
.B1(n_147),
.B2(n_177),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_29),
.A2(n_33),
.B1(n_190),
.B2(n_231),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_29),
.A2(n_33),
.B1(n_187),
.B2(n_243),
.Y(n_242)
);

AOI22xp33_ASAP7_75t_L g247 ( 
.A1(n_29),
.A2(n_33),
.B1(n_236),
.B2(n_243),
.Y(n_247)
);

AND2x2_ASAP7_75t_L g29 ( 
.A(n_30),
.B(n_32),
.Y(n_29)
);

INVx3_ASAP7_75t_SL g36 ( 
.A(n_30),
.Y(n_36)
);

OA22x2_ASAP7_75t_L g48 ( 
.A1(n_30),
.A2(n_36),
.B1(n_46),
.B2(n_47),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_SL g244 ( 
.A(n_30),
.B(n_245),
.Y(n_244)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_32),
.A2(n_110),
.B1(n_145),
.B2(n_146),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_32),
.A2(n_145),
.B1(n_235),
.B2(n_237),
.Y(n_234)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

OAI21xp33_ASAP7_75t_L g224 ( 
.A1(n_36),
.A2(n_47),
.B(n_187),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_38),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_L g38 ( 
.A1(n_39),
.A2(n_44),
.B1(n_49),
.B2(n_51),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_39),
.A2(n_44),
.B1(n_51),
.B2(n_113),
.Y(n_112)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_41),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_L g45 ( 
.A1(n_41),
.A2(n_43),
.B1(n_46),
.B2(n_47),
.Y(n_45)
);

OA22x2_ASAP7_75t_L g77 ( 
.A1(n_41),
.A2(n_43),
.B1(n_75),
.B2(n_76),
.Y(n_77)
);

OAI32xp33_ASAP7_75t_L g185 ( 
.A1(n_41),
.A2(n_58),
.A3(n_75),
.B1(n_186),
.B2(n_188),
.Y(n_185)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_43),
.B(n_76),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_44),
.A2(n_49),
.B1(n_51),
.B2(n_81),
.Y(n_80)
);

OAI21xp5_ASAP7_75t_L g88 ( 
.A1(n_44),
.A2(n_51),
.B(n_81),
.Y(n_88)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_44),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_44),
.A2(n_51),
.B1(n_179),
.B2(n_181),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_44),
.A2(n_51),
.B1(n_150),
.B2(n_181),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_44),
.A2(n_51),
.B1(n_221),
.B2(n_222),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_44),
.A2(n_51),
.B1(n_222),
.B2(n_229),
.Y(n_228)
);

AND2x2_ASAP7_75t_L g44 ( 
.A(n_45),
.B(n_48),
.Y(n_44)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_46),
.Y(n_47)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_48),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_48),
.A2(n_114),
.B1(n_149),
.B2(n_151),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_48),
.A2(n_151),
.B1(n_180),
.B2(n_260),
.Y(n_259)
);

CKINVDCx14_ASAP7_75t_R g101 ( 
.A(n_52),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g52 ( 
.A1(n_53),
.A2(n_54),
.B1(n_63),
.B2(n_65),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_53),
.A2(n_54),
.B1(n_65),
.B2(n_85),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_53),
.A2(n_54),
.B1(n_63),
.B2(n_119),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_53),
.A2(n_54),
.B1(n_85),
.B2(n_133),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_53),
.A2(n_54),
.B1(n_119),
.B2(n_155),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_53),
.A2(n_54),
.B1(n_195),
.B2(n_198),
.Y(n_194)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_53),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_54),
.B(n_59),
.Y(n_53)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_54),
.Y(n_174)
);

OA22x2_ASAP7_75t_L g54 ( 
.A1(n_55),
.A2(n_56),
.B1(n_57),
.B2(n_58),
.Y(n_54)
);

INVx5_ASAP7_75t_L g58 ( 
.A(n_55),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_55),
.A2(n_58),
.B1(n_75),
.B2(n_76),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_55),
.B(n_187),
.Y(n_186)
);

OAI32xp33_ASAP7_75t_L g210 ( 
.A1(n_55),
.A2(n_57),
.A3(n_60),
.B1(n_197),
.B2(n_211),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_56),
.A2(n_57),
.B1(n_60),
.B2(n_61),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_56),
.B(n_58),
.Y(n_211)
);

INVx11_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_61),
.B(n_187),
.Y(n_197)
);

BUFx16f_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g67 ( 
.A1(n_68),
.A2(n_82),
.B1(n_94),
.B2(n_95),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_68),
.Y(n_94)
);

OAI21xp33_ASAP7_75t_L g103 ( 
.A1(n_68),
.A2(n_69),
.B(n_80),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_69),
.B(n_80),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_70),
.A2(n_73),
.B1(n_78),
.B2(n_79),
.Y(n_69)
);

INVxp67_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_71),
.A2(n_77),
.B1(n_116),
.B2(n_117),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_73),
.A2(n_78),
.B1(n_79),
.B2(n_91),
.Y(n_90)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_73),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_73),
.A2(n_79),
.B1(n_167),
.B2(n_170),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_73),
.A2(n_79),
.B1(n_280),
.B2(n_281),
.Y(n_279)
);

OAI21xp5_ASAP7_75t_SL g313 ( 
.A1(n_73),
.A2(n_79),
.B(n_314),
.Y(n_313)
);

AND2x2_ASAP7_75t_L g73 ( 
.A(n_74),
.B(n_77),
.Y(n_73)
);

INVx8_ASAP7_75t_L g76 ( 
.A(n_75),
.Y(n_76)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_77),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_77),
.A2(n_92),
.B1(n_116),
.B2(n_131),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_77),
.A2(n_116),
.B1(n_117),
.B2(n_153),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_77),
.A2(n_116),
.B1(n_171),
.B2(n_201),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_L g256 ( 
.A1(n_77),
.A2(n_168),
.B(n_257),
.Y(n_256)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_82),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_83),
.A2(n_84),
.B1(n_86),
.B2(n_87),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_83),
.A2(n_84),
.B1(n_126),
.B2(n_127),
.Y(n_125)
);

CKINVDCx14_ASAP7_75t_R g83 ( 
.A(n_84),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_84),
.B(n_88),
.C(n_90),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_84),
.B(n_124),
.C(n_127),
.Y(n_310)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_88),
.A2(n_89),
.B1(n_90),
.B2(n_93),
.Y(n_87)
);

CKINVDCx16_ASAP7_75t_R g93 ( 
.A(n_88),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_88),
.A2(n_93),
.B1(n_129),
.B2(n_130),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_88),
.B(n_130),
.C(n_132),
.Y(n_320)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

CKINVDCx14_ASAP7_75t_R g91 ( 
.A(n_92),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_102),
.C(n_104),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_97),
.A2(n_98),
.B1(n_102),
.B2(n_103),
.Y(n_158)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

XOR2xp5_ASAP7_75t_L g157 ( 
.A(n_104),
.B(n_158),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_105),
.B(n_115),
.C(n_118),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_105),
.A2(n_106),
.B1(n_138),
.B2(n_139),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_106),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_107),
.B(n_111),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g291 ( 
.A1(n_107),
.A2(n_108),
.B1(n_111),
.B2(n_112),
.Y(n_291)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVxp67_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

XOR2xp5_ASAP7_75t_L g139 ( 
.A(n_115),
.B(n_118),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_L g306 ( 
.A1(n_121),
.A2(n_307),
.B(n_308),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_122),
.B(n_123),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_122),
.B(n_123),
.Y(n_308)
);

XNOR2xp5_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_125),
.Y(n_123)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

XNOR2xp5_ASAP7_75t_L g127 ( 
.A(n_128),
.B(n_132),
.Y(n_127)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

CKINVDCx16_ASAP7_75t_R g314 ( 
.A(n_131),
.Y(n_314)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_133),
.Y(n_316)
);

OAI21xp5_ASAP7_75t_L g134 ( 
.A1(n_135),
.A2(n_159),
.B(n_305),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_136),
.B(n_157),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_136),
.B(n_157),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_140),
.C(n_141),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_L g303 ( 
.A(n_137),
.B(n_140),
.Y(n_303)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_L g302 ( 
.A(n_141),
.B(n_303),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_152),
.C(n_154),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_142),
.A2(n_143),
.B1(n_293),
.B2(n_294),
.Y(n_292)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_148),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_144),
.B(n_148),
.Y(n_276)
);

CKINVDCx16_ASAP7_75t_R g146 ( 
.A(n_147),
.Y(n_146)
);

CKINVDCx16_ASAP7_75t_R g149 ( 
.A(n_150),
.Y(n_149)
);

XOR2xp5_ASAP7_75t_L g294 ( 
.A(n_152),
.B(n_154),
.Y(n_294)
);

INVxp67_ASAP7_75t_L g281 ( 
.A(n_153),
.Y(n_281)
);

INVxp67_ASAP7_75t_L g285 ( 
.A(n_155),
.Y(n_285)
);

AOI21xp5_ASAP7_75t_L g159 ( 
.A1(n_160),
.A2(n_300),
.B(n_304),
.Y(n_159)
);

OAI221xp5_ASAP7_75t_L g160 ( 
.A1(n_161),
.A2(n_287),
.B1(n_298),
.B2(n_299),
.C(n_331),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_162),
.B(n_271),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_L g162 ( 
.A1(n_163),
.A2(n_214),
.B(n_270),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_164),
.B(n_191),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g270 ( 
.A(n_164),
.B(n_191),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_165),
.B(n_178),
.C(n_182),
.Y(n_164)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_165),
.B(n_267),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_SL g165 ( 
.A(n_166),
.B(n_172),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_166),
.B(n_173),
.C(n_175),
.Y(n_212)
);

INVxp67_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

INVxp67_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_L g172 ( 
.A(n_173),
.B(n_175),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g282 ( 
.A1(n_174),
.A2(n_283),
.B1(n_284),
.B2(n_285),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g315 ( 
.A1(n_174),
.A2(n_284),
.B1(n_316),
.B2(n_317),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_SL g325 ( 
.A1(n_174),
.A2(n_284),
.B1(n_317),
.B2(n_326),
.Y(n_325)
);

OAI22xp5_ASAP7_75t_L g267 ( 
.A1(n_178),
.A2(n_182),
.B1(n_183),
.B2(n_268),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_178),
.Y(n_268)
);

INVxp67_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_189),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_184),
.A2(n_185),
.B1(n_189),
.B2(n_262),
.Y(n_261)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

CKINVDCx16_ASAP7_75t_R g258 ( 
.A(n_186),
.Y(n_258)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_189),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_192),
.A2(n_193),
.B1(n_205),
.B2(n_213),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_192),
.B(n_206),
.C(n_212),
.Y(n_272)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g193 ( 
.A(n_194),
.B(n_199),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_194),
.B(n_200),
.C(n_204),
.Y(n_275)
);

CKINVDCx16_ASAP7_75t_R g196 ( 
.A(n_197),
.Y(n_196)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_198),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_200),
.A2(n_202),
.B1(n_203),
.B2(n_204),
.Y(n_199)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_200),
.Y(n_203)
);

INVxp67_ASAP7_75t_L g280 ( 
.A(n_201),
.Y(n_280)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_202),
.Y(n_204)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_205),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_SL g205 ( 
.A(n_206),
.B(n_212),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_207),
.A2(n_208),
.B1(n_209),
.B2(n_210),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g286 ( 
.A(n_207),
.B(n_210),
.Y(n_286)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

AOI21xp5_ASAP7_75t_L g214 ( 
.A1(n_215),
.A2(n_264),
.B(n_269),
.Y(n_214)
);

OAI21xp5_ASAP7_75t_SL g215 ( 
.A1(n_216),
.A2(n_252),
.B(n_263),
.Y(n_215)
);

AOI21xp5_ASAP7_75t_L g216 ( 
.A1(n_217),
.A2(n_232),
.B(n_251),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_225),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_SL g251 ( 
.A(n_218),
.B(n_225),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_219),
.B(n_223),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_219),
.A2(n_220),
.B1(n_223),
.B2(n_239),
.Y(n_238)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_223),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_230),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_227),
.B(n_228),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_227),
.B(n_228),
.C(n_230),
.Y(n_253)
);

INVxp67_ASAP7_75t_L g260 ( 
.A(n_229),
.Y(n_260)
);

INVxp67_ASAP7_75t_L g237 ( 
.A(n_231),
.Y(n_237)
);

OAI21xp5_ASAP7_75t_SL g232 ( 
.A1(n_233),
.A2(n_240),
.B(n_250),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_234),
.B(n_238),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_SL g250 ( 
.A(n_234),
.B(n_238),
.Y(n_250)
);

INVxp67_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

AOI21xp5_ASAP7_75t_L g240 ( 
.A1(n_241),
.A2(n_246),
.B(n_249),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_SL g241 ( 
.A(n_242),
.B(n_244),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_247),
.B(n_248),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_SL g249 ( 
.A(n_247),
.B(n_248),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_253),
.B(n_254),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_SL g263 ( 
.A(n_253),
.B(n_254),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_255),
.B(n_261),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_256),
.B(n_259),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_256),
.B(n_259),
.C(n_261),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_265),
.B(n_266),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_SL g269 ( 
.A(n_265),
.B(n_266),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_272),
.B(n_273),
.Y(n_271)
);

OR2x2_ASAP7_75t_L g298 ( 
.A(n_272),
.B(n_273),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_274),
.B(n_277),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_275),
.B(n_276),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_275),
.B(n_276),
.C(n_277),
.Y(n_288)
);

XOR2xp5_ASAP7_75t_L g277 ( 
.A(n_278),
.B(n_286),
.Y(n_277)
);

XOR2xp5_ASAP7_75t_L g278 ( 
.A(n_279),
.B(n_282),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_279),
.B(n_282),
.C(n_286),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_288),
.B(n_289),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_288),
.B(n_289),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_L g289 ( 
.A(n_290),
.B(n_297),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_291),
.A2(n_292),
.B1(n_295),
.B2(n_296),
.Y(n_290)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_291),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_291),
.B(n_296),
.C(n_297),
.Y(n_301)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_292),
.Y(n_296)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_301),
.B(n_302),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_301),
.B(n_302),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_SL g309 ( 
.A(n_310),
.B(n_311),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_310),
.B(n_311),
.Y(n_321)
);

XNOR2xp5_ASAP7_75t_L g311 ( 
.A(n_312),
.B(n_320),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_L g312 ( 
.A1(n_313),
.A2(n_315),
.B1(n_318),
.B2(n_319),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_313),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_315),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_315),
.B(n_318),
.C(n_320),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_323),
.B(n_329),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_324),
.B(n_327),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g324 ( 
.A(n_325),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_325),
.B(n_328),
.Y(n_329)
);

CKINVDCx14_ASAP7_75t_R g327 ( 
.A(n_328),
.Y(n_327)
);


endmodule