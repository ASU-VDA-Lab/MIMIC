module fake_netlist_6_375_n_1438 (n_52, n_1, n_91, n_326, n_256, n_209, n_63, n_223, n_278, n_341, n_148, n_226, n_161, n_22, n_208, n_68, n_316, n_28, n_304, n_212, n_50, n_7, n_144, n_125, n_168, n_297, n_342, n_77, n_106, n_160, n_131, n_188, n_310, n_186, n_245, n_0, n_350, n_78, n_84, n_142, n_143, n_180, n_62, n_349, n_233, n_255, n_284, n_140, n_337, n_214, n_67, n_15, n_246, n_38, n_289, n_59, n_181, n_182, n_238, n_202, n_320, n_108, n_327, n_280, n_287, n_353, n_65, n_230, n_141, n_200, n_176, n_114, n_86, n_198, n_104, n_222, n_179, n_248, n_300, n_71, n_74, n_229, n_305, n_72, n_173, n_250, n_111, n_314, n_35, n_183, n_79, n_338, n_56, n_119, n_235, n_147, n_191, n_340, n_39, n_344, n_73, n_101, n_167, n_174, n_127, n_153, n_156, n_145, n_42, n_133, n_96, n_8, n_189, n_213, n_294, n_302, n_129, n_197, n_11, n_137, n_17, n_343, n_20, n_155, n_109, n_122, n_45, n_34, n_218, n_70, n_234, n_37, n_82, n_27, n_236, n_112, n_172, n_270, n_239, n_126, n_97, n_58, n_290, n_220, n_118, n_224, n_48, n_25, n_93, n_80, n_196, n_352, n_9, n_107, n_6, n_14, n_89, n_103, n_272, n_185, n_348, n_69, n_293, n_31, n_334, n_53, n_44, n_232, n_16, n_163, n_46, n_330, n_298, n_18, n_281, n_258, n_154, n_98, n_260, n_265, n_313, n_279, n_252, n_228, n_166, n_184, n_216, n_83, n_323, n_152, n_92, n_321, n_331, n_105, n_227, n_132, n_102, n_204, n_261, n_312, n_32, n_66, n_130, n_164, n_292, n_100, n_121, n_307, n_23, n_2, n_291, n_219, n_150, n_264, n_263, n_325, n_329, n_33, n_61, n_237, n_244, n_76, n_243, n_124, n_94, n_282, n_116, n_211, n_117, n_175, n_322, n_345, n_231, n_354, n_40, n_240, n_139, n_319, n_41, n_134, n_273, n_95, n_311, n_10, n_253, n_123, n_136, n_249, n_201, n_159, n_157, n_162, n_115, n_128, n_241, n_30, n_275, n_43, n_276, n_221, n_146, n_318, n_303, n_306, n_21, n_193, n_269, n_346, n_88, n_3, n_277, n_113, n_4, n_199, n_138, n_266, n_296, n_268, n_271, n_158, n_217, n_49, n_210, n_299, n_206, n_5, n_333, n_215, n_178, n_247, n_225, n_308, n_309, n_355, n_317, n_149, n_90, n_347, n_24, n_54, n_328, n_87, n_195, n_285, n_85, n_99, n_257, n_13, n_203, n_286, n_254, n_207, n_242, n_19, n_47, n_29, n_75, n_324, n_335, n_205, n_120, n_251, n_301, n_274, n_110, n_151, n_81, n_36, n_26, n_55, n_267, n_339, n_315, n_64, n_288, n_135, n_165, n_351, n_259, n_177, n_295, n_190, n_262, n_187, n_60, n_170, n_332, n_336, n_12, n_194, n_171, n_192, n_57, n_169, n_51, n_283, n_1438);

input n_52;
input n_1;
input n_91;
input n_326;
input n_256;
input n_209;
input n_63;
input n_223;
input n_278;
input n_341;
input n_148;
input n_226;
input n_161;
input n_22;
input n_208;
input n_68;
input n_316;
input n_28;
input n_304;
input n_212;
input n_50;
input n_7;
input n_144;
input n_125;
input n_168;
input n_297;
input n_342;
input n_77;
input n_106;
input n_160;
input n_131;
input n_188;
input n_310;
input n_186;
input n_245;
input n_0;
input n_350;
input n_78;
input n_84;
input n_142;
input n_143;
input n_180;
input n_62;
input n_349;
input n_233;
input n_255;
input n_284;
input n_140;
input n_337;
input n_214;
input n_67;
input n_15;
input n_246;
input n_38;
input n_289;
input n_59;
input n_181;
input n_182;
input n_238;
input n_202;
input n_320;
input n_108;
input n_327;
input n_280;
input n_287;
input n_353;
input n_65;
input n_230;
input n_141;
input n_200;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_222;
input n_179;
input n_248;
input n_300;
input n_71;
input n_74;
input n_229;
input n_305;
input n_72;
input n_173;
input n_250;
input n_111;
input n_314;
input n_35;
input n_183;
input n_79;
input n_338;
input n_56;
input n_119;
input n_235;
input n_147;
input n_191;
input n_340;
input n_39;
input n_344;
input n_73;
input n_101;
input n_167;
input n_174;
input n_127;
input n_153;
input n_156;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_189;
input n_213;
input n_294;
input n_302;
input n_129;
input n_197;
input n_11;
input n_137;
input n_17;
input n_343;
input n_20;
input n_155;
input n_109;
input n_122;
input n_45;
input n_34;
input n_218;
input n_70;
input n_234;
input n_37;
input n_82;
input n_27;
input n_236;
input n_112;
input n_172;
input n_270;
input n_239;
input n_126;
input n_97;
input n_58;
input n_290;
input n_220;
input n_118;
input n_224;
input n_48;
input n_25;
input n_93;
input n_80;
input n_196;
input n_352;
input n_9;
input n_107;
input n_6;
input n_14;
input n_89;
input n_103;
input n_272;
input n_185;
input n_348;
input n_69;
input n_293;
input n_31;
input n_334;
input n_53;
input n_44;
input n_232;
input n_16;
input n_163;
input n_46;
input n_330;
input n_298;
input n_18;
input n_281;
input n_258;
input n_154;
input n_98;
input n_260;
input n_265;
input n_313;
input n_279;
input n_252;
input n_228;
input n_166;
input n_184;
input n_216;
input n_83;
input n_323;
input n_152;
input n_92;
input n_321;
input n_331;
input n_105;
input n_227;
input n_132;
input n_102;
input n_204;
input n_261;
input n_312;
input n_32;
input n_66;
input n_130;
input n_164;
input n_292;
input n_100;
input n_121;
input n_307;
input n_23;
input n_2;
input n_291;
input n_219;
input n_150;
input n_264;
input n_263;
input n_325;
input n_329;
input n_33;
input n_61;
input n_237;
input n_244;
input n_76;
input n_243;
input n_124;
input n_94;
input n_282;
input n_116;
input n_211;
input n_117;
input n_175;
input n_322;
input n_345;
input n_231;
input n_354;
input n_40;
input n_240;
input n_139;
input n_319;
input n_41;
input n_134;
input n_273;
input n_95;
input n_311;
input n_10;
input n_253;
input n_123;
input n_136;
input n_249;
input n_201;
input n_159;
input n_157;
input n_162;
input n_115;
input n_128;
input n_241;
input n_30;
input n_275;
input n_43;
input n_276;
input n_221;
input n_146;
input n_318;
input n_303;
input n_306;
input n_21;
input n_193;
input n_269;
input n_346;
input n_88;
input n_3;
input n_277;
input n_113;
input n_4;
input n_199;
input n_138;
input n_266;
input n_296;
input n_268;
input n_271;
input n_158;
input n_217;
input n_49;
input n_210;
input n_299;
input n_206;
input n_5;
input n_333;
input n_215;
input n_178;
input n_247;
input n_225;
input n_308;
input n_309;
input n_355;
input n_317;
input n_149;
input n_90;
input n_347;
input n_24;
input n_54;
input n_328;
input n_87;
input n_195;
input n_285;
input n_85;
input n_99;
input n_257;
input n_13;
input n_203;
input n_286;
input n_254;
input n_207;
input n_242;
input n_19;
input n_47;
input n_29;
input n_75;
input n_324;
input n_335;
input n_205;
input n_120;
input n_251;
input n_301;
input n_274;
input n_110;
input n_151;
input n_81;
input n_36;
input n_26;
input n_55;
input n_267;
input n_339;
input n_315;
input n_64;
input n_288;
input n_135;
input n_165;
input n_351;
input n_259;
input n_177;
input n_295;
input n_190;
input n_262;
input n_187;
input n_60;
input n_170;
input n_332;
input n_336;
input n_12;
input n_194;
input n_171;
input n_192;
input n_57;
input n_169;
input n_51;
input n_283;

output n_1438;

wire n_992;
wire n_801;
wire n_1234;
wire n_1199;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_1212;
wire n_726;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_783;
wire n_798;
wire n_509;
wire n_1342;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_805;
wire n_1151;
wire n_396;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1009;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1032;
wire n_1247;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_424;
wire n_1415;
wire n_1370;
wire n_369;
wire n_415;
wire n_830;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_447;
wire n_1172;
wire n_852;
wire n_1393;
wire n_1078;
wire n_544;
wire n_1140;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_616;
wire n_658;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1163;
wire n_1180;
wire n_943;
wire n_491;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_405;
wire n_538;
wire n_1106;
wire n_886;
wire n_953;
wire n_1094;
wire n_1345;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1280;
wire n_713;
wire n_1400;
wire n_976;
wire n_734;
wire n_1088;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_659;
wire n_407;
wire n_913;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_686;
wire n_757;
wire n_594;
wire n_577;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_606;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_916;
wire n_483;
wire n_608;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_1162;
wire n_860;
wire n_788;
wire n_939;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_982;
wire n_549;
wire n_1075;
wire n_408;
wire n_932;
wire n_979;
wire n_905;
wire n_993;
wire n_689;
wire n_1330;
wire n_1413;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_692;
wire n_733;
wire n_1233;
wire n_1289;
wire n_487;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1111;
wire n_715;
wire n_1251;
wire n_1265;
wire n_530;
wire n_618;
wire n_1297;
wire n_1312;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_1335;
wire n_1069;
wire n_612;
wire n_1165;
wire n_702;
wire n_1175;
wire n_1386;
wire n_429;
wire n_1012;
wire n_780;
wire n_675;
wire n_903;
wire n_835;
wire n_1214;
wire n_928;
wire n_690;
wire n_850;
wire n_816;
wire n_1157;
wire n_1188;
wire n_877;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1124;
wire n_515;
wire n_598;
wire n_696;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_697;
wire n_687;
wire n_890;
wire n_637;
wire n_701;
wire n_950;
wire n_388;
wire n_484;
wire n_891;
wire n_1412;
wire n_949;
wire n_678;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_590;
wire n_362;
wire n_1052;
wire n_462;
wire n_1033;
wire n_1296;
wire n_694;
wire n_1294;
wire n_1420;
wire n_595;
wire n_627;
wire n_524;
wire n_1044;
wire n_1391;
wire n_449;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1072;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_840;
wire n_874;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_898;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_963;
wire n_639;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_605;
wire n_826;
wire n_872;
wire n_1139;
wire n_718;
wire n_1018;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_996;
wire n_532;
wire n_1308;
wire n_1376;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_622;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1340;
wire n_631;
wire n_720;
wire n_842;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1246;
wire n_899;
wire n_738;
wire n_1304;
wire n_1035;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1181;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_648;
wire n_657;
wire n_1049;
wire n_803;
wire n_926;
wire n_927;
wire n_919;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_777;
wire n_1299;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_1195;
wire n_552;
wire n_1358;
wire n_1388;
wire n_912;
wire n_745;
wire n_1284;
wire n_1142;
wire n_716;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1395;
wire n_731;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_683;
wire n_811;
wire n_1207;
wire n_527;
wire n_1368;
wire n_1418;
wire n_958;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1382;
wire n_1372;
wire n_505;
wire n_1339;
wire n_537;
wire n_1427;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1220;
wire n_556;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_1159;
wire n_1092;
wire n_441;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1223;
wire n_511;
wire n_1286;
wire n_1053;
wire n_416;
wire n_520;
wire n_418;
wire n_1093;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_518;
wire n_1185;
wire n_453;
wire n_914;
wire n_759;
wire n_426;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1224;
wire n_1135;
wire n_1179;
wire n_1169;
wire n_401;
wire n_463;
wire n_1243;
wire n_848;
wire n_1096;
wire n_1091;
wire n_1425;
wire n_1281;
wire n_1267;
wire n_983;
wire n_427;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1419;
wire n_1437;
wire n_385;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_664;
wire n_1429;
wire n_435;
wire n_793;
wire n_587;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1079;
wire n_828;
wire n_607;
wire n_419;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_368;
wire n_575;
wire n_994;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_557;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1275;
wire n_485;
wire n_443;
wire n_892;
wire n_768;
wire n_421;
wire n_1095;
wire n_597;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1024;
wire n_517;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1015;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1126;
wire n_710;
wire n_1108;
wire n_1182;
wire n_1298;
wire n_785;
wire n_746;
wire n_609;
wire n_1356;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_380;
wire n_1190;
wire n_397;
wire n_1262;
wire n_1213;
wire n_1350;
wire n_1272;
wire n_782;
wire n_490;
wire n_809;
wire n_1043;
wire n_986;
wire n_1081;
wire n_402;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1361;
wire n_662;
wire n_374;
wire n_1152;
wire n_450;
wire n_921;
wire n_1346;
wire n_711;
wire n_579;
wire n_1352;
wire n_937;
wire n_370;
wire n_650;
wire n_1046;
wire n_1145;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_1406;
wire n_456;
wire n_1332;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_934;
wire n_482;
wire n_1407;
wire n_420;
wire n_1341;
wire n_394;
wire n_942;
wire n_543;
wire n_1271;
wire n_1355;
wire n_1225;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_1343;
wire n_548;
wire n_833;
wire n_523;
wire n_1319;
wire n_707;
wire n_799;
wire n_1155;
wire n_787;
wire n_1416;
wire n_1146;
wire n_1086;
wire n_1066;
wire n_1282;
wire n_550;
wire n_652;
wire n_560;
wire n_1241;
wire n_1321;
wire n_569;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_1292;
wire n_1373;
wire n_1029;
wire n_790;
wire n_1210;
wire n_1248;
wire n_902;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_786;
wire n_1236;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1325;
wire n_1002;
wire n_545;
wire n_489;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1360;
wire n_1200;
wire n_479;
wire n_1353;
wire n_869;
wire n_1154;
wire n_1113;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_897;
wire n_846;
wire n_841;
wire n_1001;
wire n_508;
wire n_1050;
wire n_1411;
wire n_1177;
wire n_1150;
wire n_398;
wire n_1191;
wire n_566;
wire n_1023;
wire n_1076;
wire n_1118;
wire n_1007;
wire n_1378;
wire n_855;
wire n_591;
wire n_1377;
wire n_853;
wire n_440;
wire n_695;
wire n_875;
wire n_367;
wire n_680;
wire n_661;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_1074;
wire n_698;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_1379;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1130;
wire n_573;
wire n_769;
wire n_676;
wire n_1120;
wire n_832;
wire n_555;
wire n_389;
wire n_814;
wire n_669;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_863;
wire n_601;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_763;
wire n_1147;
wire n_360;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_1173;
wire n_525;
wire n_1116;
wire n_611;
wire n_1219;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_930;
wire n_888;
wire n_1112;
wire n_910;
wire n_911;
wire n_653;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_414;
wire n_563;
wire n_1011;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_779;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1109;
wire n_712;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_1161;
wire n_1085;
wire n_1239;
wire n_771;
wire n_470;
wire n_475;
wire n_924;
wire n_492;
wire n_1149;
wire n_1184;
wire n_719;
wire n_455;
wire n_363;
wire n_1090;
wire n_592;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_503;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_878;
wire n_620;
wire n_519;
wire n_469;
wire n_1218;
wire n_500;
wire n_981;
wire n_714;
wire n_1349;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1198;
wire n_436;
wire n_409;
wire n_1244;
wire n_756;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_583;
wire n_1039;
wire n_1034;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_467;
wire n_359;
wire n_973;
wire n_1055;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_404;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_588;
wire n_1260;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_534;
wire n_1006;
wire n_373;
wire n_730;
wire n_1311;
wire n_670;
wire n_1089;
wire n_1365;
wire n_1417;
wire n_1242;
wire n_681;
wire n_1226;
wire n_1274;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_784;
wire n_434;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_900;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_1013;
wire n_1259;
wire n_649;
wire n_1240;

CKINVDCx14_ASAP7_75t_R g356 ( 
.A(n_79),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_246),
.Y(n_357)
);

INVx2_ASAP7_75t_SL g358 ( 
.A(n_296),
.Y(n_358)
);

BUFx10_ASAP7_75t_L g359 ( 
.A(n_107),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_201),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_83),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_343),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_81),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_281),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_179),
.Y(n_365)
);

BUFx3_ASAP7_75t_L g366 ( 
.A(n_213),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_73),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_312),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_6),
.Y(n_369)
);

HB1xp67_ASAP7_75t_L g370 ( 
.A(n_310),
.Y(n_370)
);

INVx2_ASAP7_75t_SL g371 ( 
.A(n_77),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_20),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_60),
.Y(n_373)
);

INVx2_ASAP7_75t_L g374 ( 
.A(n_348),
.Y(n_374)
);

CKINVDCx16_ASAP7_75t_R g375 ( 
.A(n_48),
.Y(n_375)
);

INVx1_ASAP7_75t_SL g376 ( 
.A(n_17),
.Y(n_376)
);

BUFx6f_ASAP7_75t_L g377 ( 
.A(n_134),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_282),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_198),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_132),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_114),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_340),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_279),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_350),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_53),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_196),
.Y(n_386)
);

BUFx6f_ASAP7_75t_L g387 ( 
.A(n_122),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_184),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_335),
.Y(n_389)
);

CKINVDCx16_ASAP7_75t_R g390 ( 
.A(n_101),
.Y(n_390)
);

INVx2_ASAP7_75t_L g391 ( 
.A(n_244),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_193),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_178),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_219),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_344),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_129),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_324),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_338),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_316),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_283),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_259),
.Y(n_401)
);

BUFx10_ASAP7_75t_L g402 ( 
.A(n_288),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_19),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_154),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_263),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_17),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_141),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_88),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_212),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_157),
.Y(n_410)
);

CKINVDCx14_ASAP7_75t_R g411 ( 
.A(n_5),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_26),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_115),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_131),
.Y(n_414)
);

INVx1_ASAP7_75t_SL g415 ( 
.A(n_10),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_266),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_108),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_251),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_286),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_225),
.Y(n_420)
);

CKINVDCx20_ASAP7_75t_R g421 ( 
.A(n_208),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_90),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_243),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_238),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_71),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_209),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_105),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_200),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_34),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_7),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_321),
.Y(n_431)
);

CKINVDCx5p33_ASAP7_75t_R g432 ( 
.A(n_44),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_218),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_317),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_153),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_124),
.Y(n_436)
);

INVx2_ASAP7_75t_SL g437 ( 
.A(n_216),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_126),
.Y(n_438)
);

BUFx10_ASAP7_75t_L g439 ( 
.A(n_125),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_138),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_99),
.Y(n_441)
);

CKINVDCx5p33_ASAP7_75t_R g442 ( 
.A(n_82),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_62),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_151),
.Y(n_444)
);

INVx2_ASAP7_75t_L g445 ( 
.A(n_267),
.Y(n_445)
);

HB1xp67_ASAP7_75t_L g446 ( 
.A(n_355),
.Y(n_446)
);

CKINVDCx16_ASAP7_75t_R g447 ( 
.A(n_248),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_242),
.Y(n_448)
);

INVx1_ASAP7_75t_SL g449 ( 
.A(n_110),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_117),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_56),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_289),
.Y(n_452)
);

CKINVDCx20_ASAP7_75t_R g453 ( 
.A(n_42),
.Y(n_453)
);

INVx2_ASAP7_75t_L g454 ( 
.A(n_334),
.Y(n_454)
);

CKINVDCx5p33_ASAP7_75t_R g455 ( 
.A(n_258),
.Y(n_455)
);

CKINVDCx5p33_ASAP7_75t_R g456 ( 
.A(n_195),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_164),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_128),
.Y(n_458)
);

CKINVDCx5p33_ASAP7_75t_R g459 ( 
.A(n_65),
.Y(n_459)
);

CKINVDCx5p33_ASAP7_75t_R g460 ( 
.A(n_185),
.Y(n_460)
);

BUFx5_ASAP7_75t_L g461 ( 
.A(n_330),
.Y(n_461)
);

CKINVDCx5p33_ASAP7_75t_R g462 ( 
.A(n_158),
.Y(n_462)
);

CKINVDCx5p33_ASAP7_75t_R g463 ( 
.A(n_301),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_223),
.Y(n_464)
);

CKINVDCx20_ASAP7_75t_R g465 ( 
.A(n_85),
.Y(n_465)
);

BUFx6f_ASAP7_75t_L g466 ( 
.A(n_277),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_50),
.Y(n_467)
);

CKINVDCx5p33_ASAP7_75t_R g468 ( 
.A(n_323),
.Y(n_468)
);

INVxp67_ASAP7_75t_L g469 ( 
.A(n_34),
.Y(n_469)
);

CKINVDCx5p33_ASAP7_75t_R g470 ( 
.A(n_294),
.Y(n_470)
);

CKINVDCx20_ASAP7_75t_R g471 ( 
.A(n_197),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_347),
.Y(n_472)
);

CKINVDCx5p33_ASAP7_75t_R g473 ( 
.A(n_127),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_285),
.Y(n_474)
);

INVx2_ASAP7_75t_L g475 ( 
.A(n_74),
.Y(n_475)
);

CKINVDCx5p33_ASAP7_75t_R g476 ( 
.A(n_44),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_25),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_176),
.Y(n_478)
);

CKINVDCx5p33_ASAP7_75t_R g479 ( 
.A(n_303),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_311),
.Y(n_480)
);

CKINVDCx5p33_ASAP7_75t_R g481 ( 
.A(n_166),
.Y(n_481)
);

CKINVDCx5p33_ASAP7_75t_R g482 ( 
.A(n_337),
.Y(n_482)
);

CKINVDCx5p33_ASAP7_75t_R g483 ( 
.A(n_104),
.Y(n_483)
);

CKINVDCx5p33_ASAP7_75t_R g484 ( 
.A(n_149),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_271),
.Y(n_485)
);

CKINVDCx5p33_ASAP7_75t_R g486 ( 
.A(n_284),
.Y(n_486)
);

BUFx6f_ASAP7_75t_L g487 ( 
.A(n_237),
.Y(n_487)
);

CKINVDCx20_ASAP7_75t_R g488 ( 
.A(n_181),
.Y(n_488)
);

CKINVDCx5p33_ASAP7_75t_R g489 ( 
.A(n_121),
.Y(n_489)
);

CKINVDCx5p33_ASAP7_75t_R g490 ( 
.A(n_260),
.Y(n_490)
);

CKINVDCx5p33_ASAP7_75t_R g491 ( 
.A(n_57),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_80),
.Y(n_492)
);

CKINVDCx5p33_ASAP7_75t_R g493 ( 
.A(n_264),
.Y(n_493)
);

CKINVDCx5p33_ASAP7_75t_R g494 ( 
.A(n_119),
.Y(n_494)
);

CKINVDCx5p33_ASAP7_75t_R g495 ( 
.A(n_328),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_23),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_146),
.Y(n_497)
);

CKINVDCx5p33_ASAP7_75t_R g498 ( 
.A(n_172),
.Y(n_498)
);

INVx2_ASAP7_75t_L g499 ( 
.A(n_57),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_304),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_342),
.Y(n_501)
);

CKINVDCx5p33_ASAP7_75t_R g502 ( 
.A(n_8),
.Y(n_502)
);

BUFx3_ASAP7_75t_L g503 ( 
.A(n_106),
.Y(n_503)
);

CKINVDCx5p33_ASAP7_75t_R g504 ( 
.A(n_174),
.Y(n_504)
);

CKINVDCx5p33_ASAP7_75t_R g505 ( 
.A(n_269),
.Y(n_505)
);

CKINVDCx5p33_ASAP7_75t_R g506 ( 
.A(n_91),
.Y(n_506)
);

CKINVDCx5p33_ASAP7_75t_R g507 ( 
.A(n_5),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_160),
.Y(n_508)
);

CKINVDCx5p33_ASAP7_75t_R g509 ( 
.A(n_92),
.Y(n_509)
);

CKINVDCx5p33_ASAP7_75t_R g510 ( 
.A(n_306),
.Y(n_510)
);

CKINVDCx5p33_ASAP7_75t_R g511 ( 
.A(n_341),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_118),
.Y(n_512)
);

CKINVDCx5p33_ASAP7_75t_R g513 ( 
.A(n_332),
.Y(n_513)
);

INVx2_ASAP7_75t_L g514 ( 
.A(n_69),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_322),
.Y(n_515)
);

CKINVDCx5p33_ASAP7_75t_R g516 ( 
.A(n_346),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_291),
.Y(n_517)
);

CKINVDCx5p33_ASAP7_75t_R g518 ( 
.A(n_254),
.Y(n_518)
);

CKINVDCx5p33_ASAP7_75t_R g519 ( 
.A(n_235),
.Y(n_519)
);

CKINVDCx16_ASAP7_75t_R g520 ( 
.A(n_325),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_50),
.Y(n_521)
);

CKINVDCx20_ASAP7_75t_R g522 ( 
.A(n_190),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_308),
.Y(n_523)
);

CKINVDCx5p33_ASAP7_75t_R g524 ( 
.A(n_299),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_327),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_287),
.Y(n_526)
);

CKINVDCx5p33_ASAP7_75t_R g527 ( 
.A(n_349),
.Y(n_527)
);

CKINVDCx5p33_ASAP7_75t_R g528 ( 
.A(n_318),
.Y(n_528)
);

CKINVDCx5p33_ASAP7_75t_R g529 ( 
.A(n_24),
.Y(n_529)
);

CKINVDCx5p33_ASAP7_75t_R g530 ( 
.A(n_234),
.Y(n_530)
);

INVx2_ASAP7_75t_SL g531 ( 
.A(n_49),
.Y(n_531)
);

CKINVDCx5p33_ASAP7_75t_R g532 ( 
.A(n_102),
.Y(n_532)
);

CKINVDCx5p33_ASAP7_75t_R g533 ( 
.A(n_314),
.Y(n_533)
);

INVx2_ASAP7_75t_L g534 ( 
.A(n_309),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_55),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_293),
.Y(n_536)
);

CKINVDCx5p33_ASAP7_75t_R g537 ( 
.A(n_275),
.Y(n_537)
);

CKINVDCx5p33_ASAP7_75t_R g538 ( 
.A(n_253),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_48),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_353),
.Y(n_540)
);

CKINVDCx5p33_ASAP7_75t_R g541 ( 
.A(n_97),
.Y(n_541)
);

CKINVDCx5p33_ASAP7_75t_R g542 ( 
.A(n_162),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_30),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_140),
.Y(n_544)
);

CKINVDCx5p33_ASAP7_75t_R g545 ( 
.A(n_4),
.Y(n_545)
);

INVx1_ASAP7_75t_SL g546 ( 
.A(n_100),
.Y(n_546)
);

CKINVDCx5p33_ASAP7_75t_R g547 ( 
.A(n_298),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_130),
.Y(n_548)
);

CKINVDCx5p33_ASAP7_75t_R g549 ( 
.A(n_177),
.Y(n_549)
);

CKINVDCx20_ASAP7_75t_R g550 ( 
.A(n_211),
.Y(n_550)
);

INVx2_ASAP7_75t_SL g551 ( 
.A(n_76),
.Y(n_551)
);

CKINVDCx5p33_ASAP7_75t_R g552 ( 
.A(n_14),
.Y(n_552)
);

CKINVDCx5p33_ASAP7_75t_R g553 ( 
.A(n_300),
.Y(n_553)
);

CKINVDCx5p33_ASAP7_75t_R g554 ( 
.A(n_194),
.Y(n_554)
);

CKINVDCx5p33_ASAP7_75t_R g555 ( 
.A(n_150),
.Y(n_555)
);

CKINVDCx5p33_ASAP7_75t_R g556 ( 
.A(n_220),
.Y(n_556)
);

NOR2xp33_ASAP7_75t_L g557 ( 
.A(n_370),
.B(n_0),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_403),
.Y(n_558)
);

CKINVDCx20_ASAP7_75t_R g559 ( 
.A(n_453),
.Y(n_559)
);

CKINVDCx5p33_ASAP7_75t_R g560 ( 
.A(n_357),
.Y(n_560)
);

CKINVDCx16_ASAP7_75t_R g561 ( 
.A(n_375),
.Y(n_561)
);

HB1xp67_ASAP7_75t_L g562 ( 
.A(n_369),
.Y(n_562)
);

CKINVDCx5p33_ASAP7_75t_R g563 ( 
.A(n_360),
.Y(n_563)
);

CKINVDCx5p33_ASAP7_75t_R g564 ( 
.A(n_361),
.Y(n_564)
);

INVx2_ASAP7_75t_L g565 ( 
.A(n_461),
.Y(n_565)
);

CKINVDCx5p33_ASAP7_75t_R g566 ( 
.A(n_362),
.Y(n_566)
);

HB1xp67_ASAP7_75t_L g567 ( 
.A(n_372),
.Y(n_567)
);

CKINVDCx5p33_ASAP7_75t_R g568 ( 
.A(n_364),
.Y(n_568)
);

CKINVDCx5p33_ASAP7_75t_R g569 ( 
.A(n_365),
.Y(n_569)
);

NOR2xp33_ASAP7_75t_L g570 ( 
.A(n_446),
.B(n_0),
.Y(n_570)
);

INVxp67_ASAP7_75t_L g571 ( 
.A(n_412),
.Y(n_571)
);

BUFx2_ASAP7_75t_L g572 ( 
.A(n_411),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_451),
.Y(n_573)
);

CKINVDCx5p33_ASAP7_75t_R g574 ( 
.A(n_367),
.Y(n_574)
);

NOR2xp33_ASAP7_75t_L g575 ( 
.A(n_411),
.B(n_1),
.Y(n_575)
);

CKINVDCx5p33_ASAP7_75t_R g576 ( 
.A(n_368),
.Y(n_576)
);

CKINVDCx5p33_ASAP7_75t_R g577 ( 
.A(n_378),
.Y(n_577)
);

INVxp33_ASAP7_75t_SL g578 ( 
.A(n_373),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_467),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_477),
.Y(n_580)
);

CKINVDCx5p33_ASAP7_75t_R g581 ( 
.A(n_379),
.Y(n_581)
);

CKINVDCx5p33_ASAP7_75t_R g582 ( 
.A(n_380),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_496),
.Y(n_583)
);

CKINVDCx5p33_ASAP7_75t_R g584 ( 
.A(n_381),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_521),
.Y(n_585)
);

CKINVDCx5p33_ASAP7_75t_R g586 ( 
.A(n_382),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_535),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_539),
.Y(n_588)
);

CKINVDCx20_ASAP7_75t_R g589 ( 
.A(n_465),
.Y(n_589)
);

CKINVDCx5p33_ASAP7_75t_R g590 ( 
.A(n_383),
.Y(n_590)
);

BUFx3_ASAP7_75t_L g591 ( 
.A(n_366),
.Y(n_591)
);

CKINVDCx20_ASAP7_75t_R g592 ( 
.A(n_465),
.Y(n_592)
);

CKINVDCx5p33_ASAP7_75t_R g593 ( 
.A(n_384),
.Y(n_593)
);

INVxp67_ASAP7_75t_SL g594 ( 
.A(n_366),
.Y(n_594)
);

CKINVDCx5p33_ASAP7_75t_R g595 ( 
.A(n_386),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_543),
.Y(n_596)
);

INVxp67_ASAP7_75t_L g597 ( 
.A(n_531),
.Y(n_597)
);

NOR2xp67_ASAP7_75t_L g598 ( 
.A(n_469),
.B(n_1),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_503),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_503),
.Y(n_600)
);

CKINVDCx5p33_ASAP7_75t_R g601 ( 
.A(n_389),
.Y(n_601)
);

CKINVDCx20_ASAP7_75t_R g602 ( 
.A(n_550),
.Y(n_602)
);

INVxp67_ASAP7_75t_L g603 ( 
.A(n_376),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_363),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_388),
.Y(n_605)
);

CKINVDCx20_ASAP7_75t_R g606 ( 
.A(n_550),
.Y(n_606)
);

CKINVDCx5p33_ASAP7_75t_R g607 ( 
.A(n_392),
.Y(n_607)
);

CKINVDCx5p33_ASAP7_75t_R g608 ( 
.A(n_393),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_398),
.Y(n_609)
);

CKINVDCx16_ASAP7_75t_R g610 ( 
.A(n_390),
.Y(n_610)
);

NOR2xp67_ASAP7_75t_L g611 ( 
.A(n_499),
.B(n_2),
.Y(n_611)
);

CKINVDCx5p33_ASAP7_75t_R g612 ( 
.A(n_394),
.Y(n_612)
);

HB1xp67_ASAP7_75t_L g613 ( 
.A(n_385),
.Y(n_613)
);

CKINVDCx5p33_ASAP7_75t_R g614 ( 
.A(n_395),
.Y(n_614)
);

CKINVDCx20_ASAP7_75t_R g615 ( 
.A(n_406),
.Y(n_615)
);

INVxp67_ASAP7_75t_SL g616 ( 
.A(n_399),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_404),
.Y(n_617)
);

INVxp33_ASAP7_75t_L g618 ( 
.A(n_499),
.Y(n_618)
);

CKINVDCx20_ASAP7_75t_R g619 ( 
.A(n_429),
.Y(n_619)
);

NOR2xp67_ASAP7_75t_L g620 ( 
.A(n_374),
.B(n_2),
.Y(n_620)
);

NOR2xp33_ASAP7_75t_L g621 ( 
.A(n_358),
.B(n_3),
.Y(n_621)
);

CKINVDCx5p33_ASAP7_75t_R g622 ( 
.A(n_396),
.Y(n_622)
);

INVxp67_ASAP7_75t_L g623 ( 
.A(n_415),
.Y(n_623)
);

CKINVDCx20_ASAP7_75t_R g624 ( 
.A(n_430),
.Y(n_624)
);

BUFx2_ASAP7_75t_L g625 ( 
.A(n_432),
.Y(n_625)
);

CKINVDCx5p33_ASAP7_75t_R g626 ( 
.A(n_397),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_405),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_407),
.Y(n_628)
);

INVx2_ASAP7_75t_L g629 ( 
.A(n_461),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_408),
.Y(n_630)
);

INVx2_ASAP7_75t_L g631 ( 
.A(n_461),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_409),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_417),
.Y(n_633)
);

CKINVDCx20_ASAP7_75t_R g634 ( 
.A(n_421),
.Y(n_634)
);

INVxp67_ASAP7_75t_SL g635 ( 
.A(n_418),
.Y(n_635)
);

CKINVDCx5p33_ASAP7_75t_R g636 ( 
.A(n_400),
.Y(n_636)
);

CKINVDCx5p33_ASAP7_75t_R g637 ( 
.A(n_401),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_422),
.Y(n_638)
);

CKINVDCx16_ASAP7_75t_R g639 ( 
.A(n_447),
.Y(n_639)
);

CKINVDCx20_ASAP7_75t_R g640 ( 
.A(n_471),
.Y(n_640)
);

CKINVDCx5p33_ASAP7_75t_R g641 ( 
.A(n_410),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_423),
.Y(n_642)
);

CKINVDCx5p33_ASAP7_75t_R g643 ( 
.A(n_413),
.Y(n_643)
);

BUFx3_ASAP7_75t_L g644 ( 
.A(n_359),
.Y(n_644)
);

CKINVDCx20_ASAP7_75t_R g645 ( 
.A(n_443),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_425),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_427),
.Y(n_647)
);

CKINVDCx5p33_ASAP7_75t_R g648 ( 
.A(n_414),
.Y(n_648)
);

NOR2xp33_ASAP7_75t_L g649 ( 
.A(n_371),
.B(n_3),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_434),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_436),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_440),
.Y(n_652)
);

CKINVDCx20_ASAP7_75t_R g653 ( 
.A(n_476),
.Y(n_653)
);

CKINVDCx20_ASAP7_75t_R g654 ( 
.A(n_491),
.Y(n_654)
);

INVxp67_ASAP7_75t_L g655 ( 
.A(n_502),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_441),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_L g657 ( 
.A(n_437),
.B(n_4),
.Y(n_657)
);

CKINVDCx5p33_ASAP7_75t_R g658 ( 
.A(n_416),
.Y(n_658)
);

CKINVDCx16_ASAP7_75t_R g659 ( 
.A(n_520),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_448),
.Y(n_660)
);

BUFx2_ASAP7_75t_L g661 ( 
.A(n_615),
.Y(n_661)
);

AND2x2_ASAP7_75t_L g662 ( 
.A(n_572),
.B(n_356),
.Y(n_662)
);

AND2x2_ASAP7_75t_L g663 ( 
.A(n_655),
.B(n_356),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_604),
.Y(n_664)
);

CKINVDCx5p33_ASAP7_75t_R g665 ( 
.A(n_560),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_L g666 ( 
.A(n_563),
.B(n_551),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_L g667 ( 
.A(n_564),
.B(n_374),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_L g668 ( 
.A(n_566),
.B(n_391),
.Y(n_668)
);

INVx2_ASAP7_75t_L g669 ( 
.A(n_565),
.Y(n_669)
);

CKINVDCx20_ASAP7_75t_R g670 ( 
.A(n_634),
.Y(n_670)
);

CKINVDCx5p33_ASAP7_75t_R g671 ( 
.A(n_568),
.Y(n_671)
);

INVx3_ASAP7_75t_L g672 ( 
.A(n_591),
.Y(n_672)
);

CKINVDCx5p33_ASAP7_75t_R g673 ( 
.A(n_569),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_L g674 ( 
.A(n_574),
.B(n_391),
.Y(n_674)
);

HB1xp67_ASAP7_75t_L g675 ( 
.A(n_603),
.Y(n_675)
);

BUFx8_ASAP7_75t_L g676 ( 
.A(n_625),
.Y(n_676)
);

BUFx6f_ASAP7_75t_L g677 ( 
.A(n_558),
.Y(n_677)
);

AND2x2_ASAP7_75t_L g678 ( 
.A(n_562),
.B(n_359),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_L g679 ( 
.A(n_576),
.B(n_577),
.Y(n_679)
);

BUFx6f_ASAP7_75t_L g680 ( 
.A(n_573),
.Y(n_680)
);

AND2x2_ASAP7_75t_L g681 ( 
.A(n_567),
.B(n_402),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_605),
.Y(n_682)
);

AND2x2_ASAP7_75t_L g683 ( 
.A(n_613),
.B(n_402),
.Y(n_683)
);

HB1xp67_ASAP7_75t_L g684 ( 
.A(n_623),
.Y(n_684)
);

INVx1_ASAP7_75t_SL g685 ( 
.A(n_589),
.Y(n_685)
);

INVxp67_ASAP7_75t_L g686 ( 
.A(n_644),
.Y(n_686)
);

AND2x2_ASAP7_75t_L g687 ( 
.A(n_594),
.B(n_439),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_609),
.Y(n_688)
);

AND2x4_ASAP7_75t_L g689 ( 
.A(n_644),
.B(n_445),
.Y(n_689)
);

NAND2xp33_ASAP7_75t_SL g690 ( 
.A(n_657),
.B(n_507),
.Y(n_690)
);

CKINVDCx20_ASAP7_75t_R g691 ( 
.A(n_640),
.Y(n_691)
);

INVxp67_ASAP7_75t_L g692 ( 
.A(n_591),
.Y(n_692)
);

INVx2_ASAP7_75t_L g693 ( 
.A(n_565),
.Y(n_693)
);

HB1xp67_ASAP7_75t_L g694 ( 
.A(n_597),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_617),
.Y(n_695)
);

CKINVDCx20_ASAP7_75t_R g696 ( 
.A(n_589),
.Y(n_696)
);

NOR2xp33_ASAP7_75t_R g697 ( 
.A(n_581),
.B(n_488),
.Y(n_697)
);

CKINVDCx20_ASAP7_75t_R g698 ( 
.A(n_592),
.Y(n_698)
);

CKINVDCx5p33_ASAP7_75t_R g699 ( 
.A(n_582),
.Y(n_699)
);

BUFx6f_ASAP7_75t_L g700 ( 
.A(n_579),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_627),
.Y(n_701)
);

CKINVDCx5p33_ASAP7_75t_R g702 ( 
.A(n_584),
.Y(n_702)
);

NOR2xp33_ASAP7_75t_R g703 ( 
.A(n_586),
.B(n_522),
.Y(n_703)
);

INVx2_ASAP7_75t_L g704 ( 
.A(n_629),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_628),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_630),
.Y(n_706)
);

CKINVDCx5p33_ASAP7_75t_R g707 ( 
.A(n_590),
.Y(n_707)
);

AND3x1_ASAP7_75t_L g708 ( 
.A(n_557),
.B(n_454),
.C(n_445),
.Y(n_708)
);

CKINVDCx5p33_ASAP7_75t_R g709 ( 
.A(n_593),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_632),
.Y(n_710)
);

AND2x4_ASAP7_75t_L g711 ( 
.A(n_616),
.B(n_454),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_633),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_638),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_642),
.Y(n_714)
);

BUFx6f_ASAP7_75t_L g715 ( 
.A(n_580),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_646),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_647),
.Y(n_717)
);

AND2x2_ASAP7_75t_L g718 ( 
.A(n_618),
.B(n_439),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_650),
.Y(n_719)
);

XNOR2xp5_ASAP7_75t_L g720 ( 
.A(n_592),
.B(n_529),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_651),
.Y(n_721)
);

INVx2_ASAP7_75t_L g722 ( 
.A(n_629),
.Y(n_722)
);

CKINVDCx5p33_ASAP7_75t_R g723 ( 
.A(n_595),
.Y(n_723)
);

CKINVDCx5p33_ASAP7_75t_R g724 ( 
.A(n_601),
.Y(n_724)
);

CKINVDCx5p33_ASAP7_75t_R g725 ( 
.A(n_607),
.Y(n_725)
);

INVx2_ASAP7_75t_L g726 ( 
.A(n_631),
.Y(n_726)
);

CKINVDCx20_ASAP7_75t_R g727 ( 
.A(n_602),
.Y(n_727)
);

INVx3_ASAP7_75t_L g728 ( 
.A(n_583),
.Y(n_728)
);

CKINVDCx20_ASAP7_75t_R g729 ( 
.A(n_602),
.Y(n_729)
);

CKINVDCx5p33_ASAP7_75t_R g730 ( 
.A(n_608),
.Y(n_730)
);

INVxp67_ASAP7_75t_L g731 ( 
.A(n_570),
.Y(n_731)
);

NAND2xp33_ASAP7_75t_R g732 ( 
.A(n_578),
.B(n_545),
.Y(n_732)
);

CKINVDCx5p33_ASAP7_75t_R g733 ( 
.A(n_612),
.Y(n_733)
);

BUFx6f_ASAP7_75t_L g734 ( 
.A(n_585),
.Y(n_734)
);

INVx2_ASAP7_75t_L g735 ( 
.A(n_631),
.Y(n_735)
);

CKINVDCx5p33_ASAP7_75t_R g736 ( 
.A(n_614),
.Y(n_736)
);

CKINVDCx5p33_ASAP7_75t_R g737 ( 
.A(n_622),
.Y(n_737)
);

INVx2_ASAP7_75t_L g738 ( 
.A(n_652),
.Y(n_738)
);

CKINVDCx5p33_ASAP7_75t_R g739 ( 
.A(n_626),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_656),
.Y(n_740)
);

HB1xp67_ASAP7_75t_L g741 ( 
.A(n_598),
.Y(n_741)
);

BUFx10_ASAP7_75t_L g742 ( 
.A(n_636),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_660),
.Y(n_743)
);

INVx2_ASAP7_75t_L g744 ( 
.A(n_587),
.Y(n_744)
);

INVx2_ASAP7_75t_L g745 ( 
.A(n_588),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_596),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_746),
.Y(n_747)
);

INVx2_ASAP7_75t_L g748 ( 
.A(n_669),
.Y(n_748)
);

INVx4_ASAP7_75t_L g749 ( 
.A(n_672),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_L g750 ( 
.A(n_669),
.B(n_635),
.Y(n_750)
);

BUFx3_ASAP7_75t_L g751 ( 
.A(n_672),
.Y(n_751)
);

INVx2_ASAP7_75t_SL g752 ( 
.A(n_718),
.Y(n_752)
);

OR2x6_ASAP7_75t_L g753 ( 
.A(n_675),
.B(n_571),
.Y(n_753)
);

AND2x2_ASAP7_75t_L g754 ( 
.A(n_675),
.B(n_610),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_664),
.Y(n_755)
);

INVx4_ASAP7_75t_SL g756 ( 
.A(n_711),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_682),
.Y(n_757)
);

INVx2_ASAP7_75t_L g758 ( 
.A(n_693),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_688),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_695),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_701),
.Y(n_761)
);

INVx2_ASAP7_75t_L g762 ( 
.A(n_693),
.Y(n_762)
);

OR2x6_ASAP7_75t_L g763 ( 
.A(n_684),
.B(n_575),
.Y(n_763)
);

AND2x4_ASAP7_75t_L g764 ( 
.A(n_692),
.B(n_599),
.Y(n_764)
);

INVx2_ASAP7_75t_SL g765 ( 
.A(n_684),
.Y(n_765)
);

HB1xp67_ASAP7_75t_L g766 ( 
.A(n_694),
.Y(n_766)
);

INVx2_ASAP7_75t_L g767 ( 
.A(n_704),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_SL g768 ( 
.A(n_678),
.B(n_659),
.Y(n_768)
);

INVx2_ASAP7_75t_SL g769 ( 
.A(n_681),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_L g770 ( 
.A(n_704),
.B(n_722),
.Y(n_770)
);

AND3x1_ASAP7_75t_L g771 ( 
.A(n_683),
.B(n_649),
.C(n_621),
.Y(n_771)
);

INVxp67_ASAP7_75t_L g772 ( 
.A(n_694),
.Y(n_772)
);

NOR2xp33_ASAP7_75t_L g773 ( 
.A(n_731),
.B(n_637),
.Y(n_773)
);

AND2x2_ASAP7_75t_L g774 ( 
.A(n_662),
.B(n_639),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_705),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_SL g776 ( 
.A(n_697),
.B(n_641),
.Y(n_776)
);

AND2x2_ASAP7_75t_SL g777 ( 
.A(n_708),
.B(n_561),
.Y(n_777)
);

BUFx6f_ASAP7_75t_L g778 ( 
.A(n_677),
.Y(n_778)
);

AND2x2_ASAP7_75t_SL g779 ( 
.A(n_661),
.B(n_475),
.Y(n_779)
);

INVx4_ASAP7_75t_L g780 ( 
.A(n_677),
.Y(n_780)
);

AOI22xp33_ASAP7_75t_L g781 ( 
.A1(n_711),
.A2(n_620),
.B1(n_618),
.B2(n_611),
.Y(n_781)
);

NOR2xp33_ASAP7_75t_L g782 ( 
.A(n_667),
.B(n_643),
.Y(n_782)
);

INVx8_ASAP7_75t_L g783 ( 
.A(n_665),
.Y(n_783)
);

INVx2_ASAP7_75t_L g784 ( 
.A(n_722),
.Y(n_784)
);

AND2x2_ASAP7_75t_L g785 ( 
.A(n_741),
.B(n_648),
.Y(n_785)
);

OR2x6_ASAP7_75t_L g786 ( 
.A(n_679),
.B(n_600),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_L g787 ( 
.A(n_726),
.B(n_735),
.Y(n_787)
);

CKINVDCx5p33_ASAP7_75t_R g788 ( 
.A(n_671),
.Y(n_788)
);

INVx2_ASAP7_75t_L g789 ( 
.A(n_726),
.Y(n_789)
);

CKINVDCx5p33_ASAP7_75t_R g790 ( 
.A(n_673),
.Y(n_790)
);

INVx2_ASAP7_75t_L g791 ( 
.A(n_735),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_L g792 ( 
.A(n_706),
.B(n_475),
.Y(n_792)
);

INVx3_ASAP7_75t_L g793 ( 
.A(n_677),
.Y(n_793)
);

INVx2_ASAP7_75t_L g794 ( 
.A(n_677),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_710),
.Y(n_795)
);

INVx2_ASAP7_75t_L g796 ( 
.A(n_680),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_712),
.Y(n_797)
);

BUFx6f_ASAP7_75t_L g798 ( 
.A(n_680),
.Y(n_798)
);

NOR2xp33_ASAP7_75t_L g799 ( 
.A(n_668),
.B(n_658),
.Y(n_799)
);

NOR3xp33_ASAP7_75t_SL g800 ( 
.A(n_732),
.B(n_552),
.C(n_420),
.Y(n_800)
);

NAND2xp33_ASAP7_75t_L g801 ( 
.A(n_674),
.B(n_377),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_713),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_SL g803 ( 
.A(n_697),
.B(n_615),
.Y(n_803)
);

NOR2xp33_ASAP7_75t_L g804 ( 
.A(n_666),
.B(n_619),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_714),
.Y(n_805)
);

BUFx2_ASAP7_75t_L g806 ( 
.A(n_703),
.Y(n_806)
);

NOR2xp33_ASAP7_75t_L g807 ( 
.A(n_663),
.B(n_619),
.Y(n_807)
);

NAND2xp33_ASAP7_75t_L g808 ( 
.A(n_741),
.B(n_377),
.Y(n_808)
);

INVx3_ASAP7_75t_L g809 ( 
.A(n_680),
.Y(n_809)
);

INVx2_ASAP7_75t_SL g810 ( 
.A(n_687),
.Y(n_810)
);

INVx2_ASAP7_75t_L g811 ( 
.A(n_680),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_L g812 ( 
.A(n_716),
.B(n_514),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_SL g813 ( 
.A(n_703),
.B(n_624),
.Y(n_813)
);

INVxp67_ASAP7_75t_L g814 ( 
.A(n_732),
.Y(n_814)
);

INVx2_ASAP7_75t_L g815 ( 
.A(n_700),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_L g816 ( 
.A(n_717),
.B(n_514),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_719),
.Y(n_817)
);

INVx5_ASAP7_75t_L g818 ( 
.A(n_700),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_721),
.Y(n_819)
);

BUFx6f_ASAP7_75t_SL g820 ( 
.A(n_742),
.Y(n_820)
);

INVx3_ASAP7_75t_L g821 ( 
.A(n_700),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_740),
.Y(n_822)
);

INVx2_ASAP7_75t_L g823 ( 
.A(n_700),
.Y(n_823)
);

BUFx10_ASAP7_75t_L g824 ( 
.A(n_699),
.Y(n_824)
);

NAND3xp33_ASAP7_75t_L g825 ( 
.A(n_743),
.B(n_534),
.C(n_452),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_715),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_SL g827 ( 
.A(n_686),
.B(n_624),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_SL g828 ( 
.A(n_702),
.B(n_654),
.Y(n_828)
);

INVx2_ASAP7_75t_L g829 ( 
.A(n_715),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_SL g830 ( 
.A(n_707),
.B(n_654),
.Y(n_830)
);

AND2x4_ASAP7_75t_L g831 ( 
.A(n_689),
.B(n_450),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_715),
.Y(n_832)
);

AOI22xp33_ASAP7_75t_L g833 ( 
.A1(n_690),
.A2(n_534),
.B1(n_458),
.B2(n_464),
.Y(n_833)
);

INVx1_ASAP7_75t_SL g834 ( 
.A(n_685),
.Y(n_834)
);

BUFx2_ASAP7_75t_L g835 ( 
.A(n_720),
.Y(n_835)
);

INVx3_ASAP7_75t_L g836 ( 
.A(n_715),
.Y(n_836)
);

BUFx10_ASAP7_75t_L g837 ( 
.A(n_709),
.Y(n_837)
);

INVx4_ASAP7_75t_L g838 ( 
.A(n_734),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_L g839 ( 
.A(n_738),
.B(n_461),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_L g840 ( 
.A(n_781),
.B(n_689),
.Y(n_840)
);

INVx3_ASAP7_75t_L g841 ( 
.A(n_749),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_L g842 ( 
.A(n_781),
.B(n_738),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_SL g843 ( 
.A(n_769),
.B(n_742),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_L g844 ( 
.A(n_750),
.B(n_728),
.Y(n_844)
);

NOR2xp33_ASAP7_75t_L g845 ( 
.A(n_773),
.B(n_782),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_747),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_L g847 ( 
.A(n_750),
.B(n_728),
.Y(n_847)
);

AOI22xp33_ASAP7_75t_L g848 ( 
.A1(n_833),
.A2(n_472),
.B1(n_474),
.B2(n_457),
.Y(n_848)
);

INVx2_ASAP7_75t_L g849 ( 
.A(n_748),
.Y(n_849)
);

OR2x2_ASAP7_75t_SL g850 ( 
.A(n_766),
.B(n_606),
.Y(n_850)
);

AO22x1_ASAP7_75t_L g851 ( 
.A1(n_785),
.A2(n_723),
.B1(n_725),
.B2(n_724),
.Y(n_851)
);

INVx2_ASAP7_75t_SL g852 ( 
.A(n_765),
.Y(n_852)
);

NAND2xp5_ASAP7_75t_L g853 ( 
.A(n_799),
.B(n_730),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_L g854 ( 
.A(n_749),
.B(n_733),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_755),
.Y(n_855)
);

AND2x6_ASAP7_75t_SL g856 ( 
.A(n_753),
.B(n_478),
.Y(n_856)
);

INVx1_ASAP7_75t_L g857 ( 
.A(n_757),
.Y(n_857)
);

AND2x2_ASAP7_75t_L g858 ( 
.A(n_772),
.B(n_736),
.Y(n_858)
);

AOI22xp33_ASAP7_75t_L g859 ( 
.A1(n_833),
.A2(n_831),
.B1(n_762),
.B2(n_767),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_SL g860 ( 
.A(n_752),
.B(n_737),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_L g861 ( 
.A(n_756),
.B(n_739),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_L g862 ( 
.A(n_756),
.B(n_734),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_L g863 ( 
.A(n_756),
.B(n_734),
.Y(n_863)
);

AND2x2_ASAP7_75t_L g864 ( 
.A(n_772),
.B(n_645),
.Y(n_864)
);

BUFx3_ASAP7_75t_L g865 ( 
.A(n_751),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_SL g866 ( 
.A(n_810),
.B(n_645),
.Y(n_866)
);

BUFx6f_ASAP7_75t_L g867 ( 
.A(n_778),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_L g868 ( 
.A(n_770),
.B(n_744),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_L g869 ( 
.A(n_759),
.B(n_734),
.Y(n_869)
);

NAND2xp5_ASAP7_75t_L g870 ( 
.A(n_760),
.B(n_480),
.Y(n_870)
);

NOR2xp33_ASAP7_75t_L g871 ( 
.A(n_814),
.B(n_653),
.Y(n_871)
);

OR2x2_ASAP7_75t_L g872 ( 
.A(n_766),
.B(n_744),
.Y(n_872)
);

AOI22xp5_ASAP7_75t_L g873 ( 
.A1(n_771),
.A2(n_653),
.B1(n_546),
.B2(n_449),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_L g874 ( 
.A(n_761),
.B(n_485),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_SL g875 ( 
.A(n_814),
.B(n_676),
.Y(n_875)
);

NAND3xp33_ASAP7_75t_SL g876 ( 
.A(n_804),
.B(n_606),
.C(n_559),
.Y(n_876)
);

NOR2xp33_ASAP7_75t_L g877 ( 
.A(n_786),
.B(n_768),
.Y(n_877)
);

INVx2_ASAP7_75t_SL g878 ( 
.A(n_764),
.Y(n_878)
);

AOI22xp5_ASAP7_75t_L g879 ( 
.A1(n_771),
.A2(n_424),
.B1(n_426),
.B2(n_419),
.Y(n_879)
);

AND2x4_ASAP7_75t_L g880 ( 
.A(n_775),
.B(n_745),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_SL g881 ( 
.A(n_774),
.B(n_676),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_L g882 ( 
.A(n_795),
.B(n_492),
.Y(n_882)
);

NAND2xp5_ASAP7_75t_L g883 ( 
.A(n_797),
.B(n_497),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_SL g884 ( 
.A(n_806),
.B(n_428),
.Y(n_884)
);

NOR2xp33_ASAP7_75t_L g885 ( 
.A(n_786),
.B(n_559),
.Y(n_885)
);

INVx2_ASAP7_75t_L g886 ( 
.A(n_758),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_802),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_L g888 ( 
.A(n_770),
.B(n_745),
.Y(n_888)
);

NOR2xp33_ASAP7_75t_L g889 ( 
.A(n_786),
.B(n_670),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_805),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_L g891 ( 
.A(n_787),
.B(n_461),
.Y(n_891)
);

INVx1_ASAP7_75t_L g892 ( 
.A(n_817),
.Y(n_892)
);

INVxp67_ASAP7_75t_L g893 ( 
.A(n_754),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_SL g894 ( 
.A(n_777),
.B(n_431),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_L g895 ( 
.A(n_787),
.B(n_461),
.Y(n_895)
);

OAI21xp5_ASAP7_75t_L g896 ( 
.A1(n_831),
.A2(n_501),
.B(n_500),
.Y(n_896)
);

INVx1_ASAP7_75t_L g897 ( 
.A(n_819),
.Y(n_897)
);

INVx1_ASAP7_75t_L g898 ( 
.A(n_822),
.Y(n_898)
);

INVx2_ASAP7_75t_L g899 ( 
.A(n_784),
.Y(n_899)
);

NOR2xp33_ASAP7_75t_L g900 ( 
.A(n_776),
.B(n_763),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_L g901 ( 
.A(n_793),
.B(n_508),
.Y(n_901)
);

INVx1_ASAP7_75t_L g902 ( 
.A(n_764),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_SL g903 ( 
.A(n_800),
.B(n_433),
.Y(n_903)
);

INVx1_ASAP7_75t_L g904 ( 
.A(n_792),
.Y(n_904)
);

INVx3_ASAP7_75t_L g905 ( 
.A(n_778),
.Y(n_905)
);

INVx2_ASAP7_75t_L g906 ( 
.A(n_789),
.Y(n_906)
);

NOR2xp33_ASAP7_75t_L g907 ( 
.A(n_763),
.B(n_691),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_SL g908 ( 
.A(n_800),
.B(n_435),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_SL g909 ( 
.A(n_779),
.B(n_438),
.Y(n_909)
);

BUFx3_ASAP7_75t_L g910 ( 
.A(n_783),
.Y(n_910)
);

AND2x4_ASAP7_75t_L g911 ( 
.A(n_794),
.B(n_512),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_L g912 ( 
.A(n_793),
.B(n_515),
.Y(n_912)
);

NOR2xp33_ASAP7_75t_L g913 ( 
.A(n_763),
.B(n_696),
.Y(n_913)
);

NOR3xp33_ASAP7_75t_SL g914 ( 
.A(n_827),
.B(n_444),
.C(n_442),
.Y(n_914)
);

AOI22xp5_ASAP7_75t_L g915 ( 
.A1(n_807),
.A2(n_456),
.B1(n_459),
.B2(n_455),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_SL g916 ( 
.A(n_778),
.B(n_460),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_792),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_L g918 ( 
.A(n_791),
.B(n_517),
.Y(n_918)
);

INVx8_ASAP7_75t_L g919 ( 
.A(n_783),
.Y(n_919)
);

INVx1_ASAP7_75t_L g920 ( 
.A(n_812),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_812),
.Y(n_921)
);

INVx2_ASAP7_75t_L g922 ( 
.A(n_809),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_816),
.Y(n_923)
);

BUFx12f_ASAP7_75t_L g924 ( 
.A(n_824),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_L g925 ( 
.A(n_816),
.B(n_523),
.Y(n_925)
);

AOI21xp5_ASAP7_75t_L g926 ( 
.A1(n_826),
.A2(n_832),
.B(n_811),
.Y(n_926)
);

HB1xp67_ASAP7_75t_L g927 ( 
.A(n_834),
.Y(n_927)
);

NOR2xp67_ASAP7_75t_L g928 ( 
.A(n_788),
.B(n_462),
.Y(n_928)
);

INVx2_ASAP7_75t_L g929 ( 
.A(n_809),
.Y(n_929)
);

INVx2_ASAP7_75t_L g930 ( 
.A(n_821),
.Y(n_930)
);

AND2x4_ASAP7_75t_L g931 ( 
.A(n_796),
.B(n_525),
.Y(n_931)
);

NAND2xp5_ASAP7_75t_L g932 ( 
.A(n_821),
.B(n_526),
.Y(n_932)
);

INVx2_ASAP7_75t_L g933 ( 
.A(n_836),
.Y(n_933)
);

INVx4_ASAP7_75t_L g934 ( 
.A(n_919),
.Y(n_934)
);

INVx1_ASAP7_75t_L g935 ( 
.A(n_846),
.Y(n_935)
);

BUFx6f_ASAP7_75t_L g936 ( 
.A(n_867),
.Y(n_936)
);

INVx1_ASAP7_75t_L g937 ( 
.A(n_855),
.Y(n_937)
);

AND2x4_ASAP7_75t_L g938 ( 
.A(n_865),
.B(n_815),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_L g939 ( 
.A(n_845),
.B(n_836),
.Y(n_939)
);

NAND3xp33_ASAP7_75t_SL g940 ( 
.A(n_873),
.B(n_834),
.C(n_727),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_SL g941 ( 
.A(n_853),
.B(n_824),
.Y(n_941)
);

INVx2_ASAP7_75t_L g942 ( 
.A(n_880),
.Y(n_942)
);

NOR3xp33_ASAP7_75t_SL g943 ( 
.A(n_876),
.B(n_830),
.C(n_828),
.Y(n_943)
);

HB1xp67_ASAP7_75t_L g944 ( 
.A(n_927),
.Y(n_944)
);

NOR2xp33_ASAP7_75t_R g945 ( 
.A(n_919),
.B(n_790),
.Y(n_945)
);

HB1xp67_ASAP7_75t_L g946 ( 
.A(n_893),
.Y(n_946)
);

INVx1_ASAP7_75t_L g947 ( 
.A(n_857),
.Y(n_947)
);

CKINVDCx6p67_ASAP7_75t_R g948 ( 
.A(n_910),
.Y(n_948)
);

BUFx3_ASAP7_75t_L g949 ( 
.A(n_924),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_L g950 ( 
.A(n_904),
.B(n_823),
.Y(n_950)
);

BUFx2_ASAP7_75t_L g951 ( 
.A(n_864),
.Y(n_951)
);

BUFx6f_ASAP7_75t_L g952 ( 
.A(n_867),
.Y(n_952)
);

O2A1O1Ixp5_ASAP7_75t_L g953 ( 
.A1(n_917),
.A2(n_921),
.B(n_923),
.C(n_920),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_L g954 ( 
.A(n_844),
.B(n_829),
.Y(n_954)
);

AND2x6_ASAP7_75t_SL g955 ( 
.A(n_913),
.B(n_753),
.Y(n_955)
);

INVx2_ASAP7_75t_L g956 ( 
.A(n_880),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_SL g957 ( 
.A(n_858),
.B(n_837),
.Y(n_957)
);

NAND2xp5_ASAP7_75t_SL g958 ( 
.A(n_854),
.B(n_837),
.Y(n_958)
);

BUFx2_ASAP7_75t_L g959 ( 
.A(n_850),
.Y(n_959)
);

A2O1A1Ixp33_ASAP7_75t_L g960 ( 
.A1(n_896),
.A2(n_825),
.B(n_803),
.C(n_813),
.Y(n_960)
);

BUFx3_ASAP7_75t_L g961 ( 
.A(n_919),
.Y(n_961)
);

BUFx3_ASAP7_75t_L g962 ( 
.A(n_852),
.Y(n_962)
);

NOR3xp33_ASAP7_75t_SL g963 ( 
.A(n_871),
.B(n_825),
.C(n_468),
.Y(n_963)
);

NAND2xp5_ASAP7_75t_L g964 ( 
.A(n_844),
.B(n_839),
.Y(n_964)
);

BUFx2_ASAP7_75t_L g965 ( 
.A(n_872),
.Y(n_965)
);

INVx1_ASAP7_75t_L g966 ( 
.A(n_887),
.Y(n_966)
);

NAND2xp5_ASAP7_75t_L g967 ( 
.A(n_847),
.B(n_839),
.Y(n_967)
);

BUFx3_ASAP7_75t_L g968 ( 
.A(n_902),
.Y(n_968)
);

AOI22xp5_ASAP7_75t_L g969 ( 
.A1(n_900),
.A2(n_780),
.B1(n_838),
.B2(n_801),
.Y(n_969)
);

NOR2xp33_ASAP7_75t_L g970 ( 
.A(n_866),
.B(n_698),
.Y(n_970)
);

NOR2xp33_ASAP7_75t_R g971 ( 
.A(n_861),
.B(n_729),
.Y(n_971)
);

INVx2_ASAP7_75t_L g972 ( 
.A(n_849),
.Y(n_972)
);

INVx5_ASAP7_75t_L g973 ( 
.A(n_841),
.Y(n_973)
);

NOR2xp33_ASAP7_75t_L g974 ( 
.A(n_877),
.B(n_860),
.Y(n_974)
);

NAND2xp5_ASAP7_75t_L g975 ( 
.A(n_847),
.B(n_780),
.Y(n_975)
);

AOI22xp5_ASAP7_75t_L g976 ( 
.A1(n_842),
.A2(n_838),
.B1(n_798),
.B2(n_808),
.Y(n_976)
);

NAND2xp5_ASAP7_75t_L g977 ( 
.A(n_868),
.B(n_798),
.Y(n_977)
);

BUFx2_ASAP7_75t_L g978 ( 
.A(n_878),
.Y(n_978)
);

OR2x2_ASAP7_75t_SL g979 ( 
.A(n_840),
.B(n_835),
.Y(n_979)
);

INVx2_ASAP7_75t_L g980 ( 
.A(n_886),
.Y(n_980)
);

BUFx12f_ASAP7_75t_L g981 ( 
.A(n_856),
.Y(n_981)
);

INVx2_ASAP7_75t_L g982 ( 
.A(n_899),
.Y(n_982)
);

INVx1_ASAP7_75t_L g983 ( 
.A(n_890),
.Y(n_983)
);

OAI22xp5_ASAP7_75t_L g984 ( 
.A1(n_848),
.A2(n_753),
.B1(n_540),
.B2(n_544),
.Y(n_984)
);

NAND3xp33_ASAP7_75t_SL g985 ( 
.A(n_879),
.B(n_470),
.C(n_463),
.Y(n_985)
);

BUFx12f_ASAP7_75t_L g986 ( 
.A(n_911),
.Y(n_986)
);

BUFx4f_ASAP7_75t_L g987 ( 
.A(n_892),
.Y(n_987)
);

NOR3xp33_ASAP7_75t_SL g988 ( 
.A(n_885),
.B(n_479),
.C(n_473),
.Y(n_988)
);

NAND2xp5_ASAP7_75t_SL g989 ( 
.A(n_840),
.B(n_783),
.Y(n_989)
);

BUFx6f_ASAP7_75t_L g990 ( 
.A(n_867),
.Y(n_990)
);

BUFx2_ASAP7_75t_L g991 ( 
.A(n_842),
.Y(n_991)
);

AND2x2_ASAP7_75t_L g992 ( 
.A(n_928),
.B(n_798),
.Y(n_992)
);

NAND2xp5_ASAP7_75t_L g993 ( 
.A(n_868),
.B(n_818),
.Y(n_993)
);

NAND2xp5_ASAP7_75t_L g994 ( 
.A(n_888),
.B(n_818),
.Y(n_994)
);

OR2x2_ASAP7_75t_L g995 ( 
.A(n_851),
.B(n_536),
.Y(n_995)
);

AOI21xp5_ASAP7_75t_L g996 ( 
.A1(n_841),
.A2(n_818),
.B(n_548),
.Y(n_996)
);

AND2x4_ASAP7_75t_L g997 ( 
.A(n_897),
.B(n_818),
.Y(n_997)
);

AND2x2_ASAP7_75t_L g998 ( 
.A(n_898),
.B(n_820),
.Y(n_998)
);

AOI22xp33_ASAP7_75t_SL g999 ( 
.A1(n_889),
.A2(n_820),
.B1(n_387),
.B2(n_466),
.Y(n_999)
);

A2O1A1Ixp33_ASAP7_75t_L g1000 ( 
.A1(n_896),
.A2(n_482),
.B(n_483),
.C(n_481),
.Y(n_1000)
);

BUFx2_ASAP7_75t_L g1001 ( 
.A(n_911),
.Y(n_1001)
);

BUFx3_ASAP7_75t_L g1002 ( 
.A(n_907),
.Y(n_1002)
);

INVx1_ASAP7_75t_L g1003 ( 
.A(n_906),
.Y(n_1003)
);

INVx3_ASAP7_75t_L g1004 ( 
.A(n_905),
.Y(n_1004)
);

AND2x4_ASAP7_75t_L g1005 ( 
.A(n_931),
.B(n_64),
.Y(n_1005)
);

NAND2xp33_ASAP7_75t_L g1006 ( 
.A(n_945),
.B(n_914),
.Y(n_1006)
);

NAND2xp5_ASAP7_75t_L g1007 ( 
.A(n_991),
.B(n_888),
.Y(n_1007)
);

INVx1_ASAP7_75t_L g1008 ( 
.A(n_935),
.Y(n_1008)
);

NAND2xp5_ASAP7_75t_L g1009 ( 
.A(n_964),
.B(n_925),
.Y(n_1009)
);

NAND2xp5_ASAP7_75t_L g1010 ( 
.A(n_939),
.B(n_925),
.Y(n_1010)
);

NOR3xp33_ASAP7_75t_L g1011 ( 
.A(n_940),
.B(n_875),
.C(n_894),
.Y(n_1011)
);

BUFx12f_ASAP7_75t_L g1012 ( 
.A(n_986),
.Y(n_1012)
);

OR2x2_ASAP7_75t_L g1013 ( 
.A(n_965),
.B(n_884),
.Y(n_1013)
);

AND2x2_ASAP7_75t_L g1014 ( 
.A(n_951),
.B(n_843),
.Y(n_1014)
);

NAND2xp5_ASAP7_75t_L g1015 ( 
.A(n_964),
.B(n_891),
.Y(n_1015)
);

OAI21xp5_ASAP7_75t_L g1016 ( 
.A1(n_953),
.A2(n_895),
.B(n_891),
.Y(n_1016)
);

OAI21x1_ASAP7_75t_L g1017 ( 
.A1(n_996),
.A2(n_954),
.B(n_950),
.Y(n_1017)
);

INVx6_ASAP7_75t_L g1018 ( 
.A(n_934),
.Y(n_1018)
);

NAND2xp5_ASAP7_75t_L g1019 ( 
.A(n_939),
.B(n_870),
.Y(n_1019)
);

OAI22xp5_ASAP7_75t_L g1020 ( 
.A1(n_960),
.A2(n_859),
.B1(n_909),
.B2(n_895),
.Y(n_1020)
);

AO21x1_ASAP7_75t_L g1021 ( 
.A1(n_967),
.A2(n_932),
.B(n_908),
.Y(n_1021)
);

NAND2xp5_ASAP7_75t_L g1022 ( 
.A(n_967),
.B(n_874),
.Y(n_1022)
);

OAI21x1_ASAP7_75t_L g1023 ( 
.A1(n_996),
.A2(n_926),
.B(n_905),
.Y(n_1023)
);

OAI21xp5_ASAP7_75t_L g1024 ( 
.A1(n_954),
.A2(n_932),
.B(n_883),
.Y(n_1024)
);

AOI21x1_ASAP7_75t_L g1025 ( 
.A1(n_975),
.A2(n_912),
.B(n_901),
.Y(n_1025)
);

OAI21x1_ASAP7_75t_L g1026 ( 
.A1(n_950),
.A2(n_929),
.B(n_922),
.Y(n_1026)
);

NAND3x1_ASAP7_75t_L g1027 ( 
.A(n_970),
.B(n_974),
.C(n_998),
.Y(n_1027)
);

BUFx6f_ASAP7_75t_L g1028 ( 
.A(n_936),
.Y(n_1028)
);

NAND2xp5_ASAP7_75t_L g1029 ( 
.A(n_977),
.B(n_882),
.Y(n_1029)
);

CKINVDCx5p33_ASAP7_75t_R g1030 ( 
.A(n_971),
.Y(n_1030)
);

AND2x2_ASAP7_75t_L g1031 ( 
.A(n_944),
.B(n_946),
.Y(n_1031)
);

NAND2xp33_ASAP7_75t_SL g1032 ( 
.A(n_943),
.B(n_881),
.Y(n_1032)
);

A2O1A1Ixp33_ASAP7_75t_L g1033 ( 
.A1(n_987),
.A2(n_915),
.B(n_869),
.C(n_903),
.Y(n_1033)
);

NAND2xp5_ASAP7_75t_L g1034 ( 
.A(n_977),
.B(n_931),
.Y(n_1034)
);

NAND2xp5_ASAP7_75t_SL g1035 ( 
.A(n_987),
.B(n_862),
.Y(n_1035)
);

NAND2x1_ASAP7_75t_L g1036 ( 
.A(n_936),
.B(n_952),
.Y(n_1036)
);

OAI21xp5_ASAP7_75t_L g1037 ( 
.A1(n_975),
.A2(n_918),
.B(n_863),
.Y(n_1037)
);

INVx1_ASAP7_75t_L g1038 ( 
.A(n_937),
.Y(n_1038)
);

INVx1_ASAP7_75t_L g1039 ( 
.A(n_947),
.Y(n_1039)
);

OAI21x1_ASAP7_75t_L g1040 ( 
.A1(n_993),
.A2(n_933),
.B(n_930),
.Y(n_1040)
);

AND2x2_ASAP7_75t_L g1041 ( 
.A(n_1001),
.B(n_918),
.Y(n_1041)
);

NAND2xp5_ASAP7_75t_L g1042 ( 
.A(n_966),
.B(n_916),
.Y(n_1042)
);

OAI21x1_ASAP7_75t_L g1043 ( 
.A1(n_993),
.A2(n_67),
.B(n_66),
.Y(n_1043)
);

OAI21x1_ASAP7_75t_L g1044 ( 
.A1(n_994),
.A2(n_70),
.B(n_68),
.Y(n_1044)
);

AOI21x1_ASAP7_75t_L g1045 ( 
.A1(n_994),
.A2(n_387),
.B(n_377),
.Y(n_1045)
);

OAI22xp5_ASAP7_75t_L g1046 ( 
.A1(n_973),
.A2(n_387),
.B1(n_466),
.B2(n_377),
.Y(n_1046)
);

OAI21xp5_ASAP7_75t_L g1047 ( 
.A1(n_1000),
.A2(n_963),
.B(n_976),
.Y(n_1047)
);

OAI21xp5_ASAP7_75t_L g1048 ( 
.A1(n_985),
.A2(n_486),
.B(n_484),
.Y(n_1048)
);

OAI21x1_ASAP7_75t_L g1049 ( 
.A1(n_1004),
.A2(n_75),
.B(n_72),
.Y(n_1049)
);

INVx2_ASAP7_75t_SL g1050 ( 
.A(n_962),
.Y(n_1050)
);

AOI21xp5_ASAP7_75t_L g1051 ( 
.A1(n_973),
.A2(n_466),
.B(n_387),
.Y(n_1051)
);

INVx3_ASAP7_75t_L g1052 ( 
.A(n_1004),
.Y(n_1052)
);

INVx2_ASAP7_75t_L g1053 ( 
.A(n_972),
.Y(n_1053)
);

OAI21x1_ASAP7_75t_L g1054 ( 
.A1(n_1003),
.A2(n_84),
.B(n_78),
.Y(n_1054)
);

AO31x2_ASAP7_75t_L g1055 ( 
.A1(n_984),
.A2(n_487),
.A3(n_466),
.B(n_8),
.Y(n_1055)
);

INVx2_ASAP7_75t_L g1056 ( 
.A(n_980),
.Y(n_1056)
);

INVx5_ASAP7_75t_L g1057 ( 
.A(n_936),
.Y(n_1057)
);

OAI21x1_ASAP7_75t_L g1058 ( 
.A1(n_982),
.A2(n_87),
.B(n_86),
.Y(n_1058)
);

NAND2xp5_ASAP7_75t_L g1059 ( 
.A(n_983),
.B(n_489),
.Y(n_1059)
);

HB1xp67_ASAP7_75t_L g1060 ( 
.A(n_978),
.Y(n_1060)
);

AND2x2_ASAP7_75t_L g1061 ( 
.A(n_942),
.B(n_490),
.Y(n_1061)
);

INVx1_ASAP7_75t_L g1062 ( 
.A(n_956),
.Y(n_1062)
);

AND2x4_ASAP7_75t_L g1063 ( 
.A(n_938),
.B(n_89),
.Y(n_1063)
);

A2O1A1Ixp33_ASAP7_75t_L g1064 ( 
.A1(n_1005),
.A2(n_556),
.B(n_493),
.C(n_495),
.Y(n_1064)
);

NAND2xp5_ASAP7_75t_L g1065 ( 
.A(n_973),
.B(n_494),
.Y(n_1065)
);

NAND2xp5_ASAP7_75t_L g1066 ( 
.A(n_1007),
.B(n_941),
.Y(n_1066)
);

INVx2_ASAP7_75t_L g1067 ( 
.A(n_1008),
.Y(n_1067)
);

NAND2x1p5_ASAP7_75t_L g1068 ( 
.A(n_1057),
.B(n_973),
.Y(n_1068)
);

OAI21x1_ASAP7_75t_L g1069 ( 
.A1(n_1040),
.A2(n_989),
.B(n_992),
.Y(n_1069)
);

OAI21xp5_ASAP7_75t_L g1070 ( 
.A1(n_1020),
.A2(n_1009),
.B(n_1022),
.Y(n_1070)
);

INVx1_ASAP7_75t_L g1071 ( 
.A(n_1038),
.Y(n_1071)
);

AO31x2_ASAP7_75t_L g1072 ( 
.A1(n_1021),
.A2(n_984),
.A3(n_959),
.B(n_979),
.Y(n_1072)
);

OA21x2_ASAP7_75t_L g1073 ( 
.A1(n_1016),
.A2(n_969),
.B(n_995),
.Y(n_1073)
);

OAI222xp33_ASAP7_75t_L g1074 ( 
.A1(n_1020),
.A2(n_999),
.B1(n_957),
.B2(n_1005),
.C1(n_958),
.C2(n_1002),
.Y(n_1074)
);

HB1xp67_ASAP7_75t_L g1075 ( 
.A(n_1060),
.Y(n_1075)
);

INVxp67_ASAP7_75t_L g1076 ( 
.A(n_1031),
.Y(n_1076)
);

BUFx3_ASAP7_75t_L g1077 ( 
.A(n_1057),
.Y(n_1077)
);

AND2x4_ASAP7_75t_L g1078 ( 
.A(n_1063),
.B(n_934),
.Y(n_1078)
);

CKINVDCx5p33_ASAP7_75t_R g1079 ( 
.A(n_1030),
.Y(n_1079)
);

OAI21xp5_ASAP7_75t_L g1080 ( 
.A1(n_1009),
.A2(n_988),
.B(n_997),
.Y(n_1080)
);

BUFx2_ASAP7_75t_L g1081 ( 
.A(n_1014),
.Y(n_1081)
);

AOI21xp5_ASAP7_75t_L g1082 ( 
.A1(n_1015),
.A2(n_997),
.B(n_990),
.Y(n_1082)
);

O2A1O1Ixp33_ASAP7_75t_L g1083 ( 
.A1(n_1011),
.A2(n_968),
.B(n_938),
.C(n_961),
.Y(n_1083)
);

OAI22xp5_ASAP7_75t_L g1084 ( 
.A1(n_1015),
.A2(n_952),
.B1(n_990),
.B2(n_948),
.Y(n_1084)
);

AND2x2_ASAP7_75t_L g1085 ( 
.A(n_1041),
.B(n_949),
.Y(n_1085)
);

OAI21x1_ASAP7_75t_L g1086 ( 
.A1(n_1026),
.A2(n_990),
.B(n_952),
.Y(n_1086)
);

NOR2xp33_ASAP7_75t_L g1087 ( 
.A(n_1042),
.B(n_955),
.Y(n_1087)
);

INVx2_ASAP7_75t_L g1088 ( 
.A(n_1039),
.Y(n_1088)
);

INVx2_ASAP7_75t_SL g1089 ( 
.A(n_1050),
.Y(n_1089)
);

INVx3_ASAP7_75t_L g1090 ( 
.A(n_1018),
.Y(n_1090)
);

INVx1_ASAP7_75t_L g1091 ( 
.A(n_1053),
.Y(n_1091)
);

AND2x4_ASAP7_75t_L g1092 ( 
.A(n_1063),
.B(n_93),
.Y(n_1092)
);

OAI21x1_ASAP7_75t_L g1093 ( 
.A1(n_1023),
.A2(n_487),
.B(n_95),
.Y(n_1093)
);

OAI21x1_ASAP7_75t_L g1094 ( 
.A1(n_1017),
.A2(n_487),
.B(n_96),
.Y(n_1094)
);

OAI21x1_ASAP7_75t_L g1095 ( 
.A1(n_1058),
.A2(n_487),
.B(n_98),
.Y(n_1095)
);

AOI21xp5_ASAP7_75t_L g1096 ( 
.A1(n_1016),
.A2(n_504),
.B(n_498),
.Y(n_1096)
);

OA21x2_ASAP7_75t_L g1097 ( 
.A1(n_1024),
.A2(n_506),
.B(n_505),
.Y(n_1097)
);

OAI21x1_ASAP7_75t_L g1098 ( 
.A1(n_1025),
.A2(n_103),
.B(n_94),
.Y(n_1098)
);

INVx2_ASAP7_75t_L g1099 ( 
.A(n_1052),
.Y(n_1099)
);

NAND2xp5_ASAP7_75t_L g1100 ( 
.A(n_1010),
.B(n_509),
.Y(n_1100)
);

A2O1A1Ixp33_ASAP7_75t_L g1101 ( 
.A1(n_1047),
.A2(n_510),
.B(n_511),
.C(n_513),
.Y(n_1101)
);

NAND2x1p5_ASAP7_75t_L g1102 ( 
.A(n_1057),
.B(n_109),
.Y(n_1102)
);

AND2x4_ASAP7_75t_L g1103 ( 
.A(n_1056),
.B(n_1062),
.Y(n_1103)
);

OAI21x1_ASAP7_75t_SL g1104 ( 
.A1(n_1047),
.A2(n_112),
.B(n_111),
.Y(n_1104)
);

INVx5_ASAP7_75t_SL g1105 ( 
.A(n_1028),
.Y(n_1105)
);

HB1xp67_ASAP7_75t_L g1106 ( 
.A(n_1028),
.Y(n_1106)
);

INVx1_ASAP7_75t_L g1107 ( 
.A(n_1052),
.Y(n_1107)
);

OAI21x1_ASAP7_75t_L g1108 ( 
.A1(n_1049),
.A2(n_116),
.B(n_113),
.Y(n_1108)
);

AOI22xp33_ASAP7_75t_L g1109 ( 
.A1(n_1032),
.A2(n_537),
.B1(n_555),
.B2(n_554),
.Y(n_1109)
);

OA21x2_ASAP7_75t_L g1110 ( 
.A1(n_1024),
.A2(n_518),
.B(n_516),
.Y(n_1110)
);

NOR2xp33_ASAP7_75t_L g1111 ( 
.A(n_1013),
.B(n_981),
.Y(n_1111)
);

NAND2x1p5_ASAP7_75t_L g1112 ( 
.A(n_1028),
.B(n_120),
.Y(n_1112)
);

AOI22xp33_ASAP7_75t_L g1113 ( 
.A1(n_1019),
.A2(n_553),
.B1(n_549),
.B2(n_547),
.Y(n_1113)
);

INVx2_ASAP7_75t_L g1114 ( 
.A(n_1029),
.Y(n_1114)
);

OAI21x1_ASAP7_75t_L g1115 ( 
.A1(n_1037),
.A2(n_133),
.B(n_123),
.Y(n_1115)
);

AOI22xp33_ASAP7_75t_L g1116 ( 
.A1(n_1048),
.A2(n_542),
.B1(n_541),
.B2(n_538),
.Y(n_1116)
);

OA21x2_ASAP7_75t_L g1117 ( 
.A1(n_1037),
.A2(n_524),
.B(n_519),
.Y(n_1117)
);

OAI21x1_ASAP7_75t_L g1118 ( 
.A1(n_1054),
.A2(n_136),
.B(n_135),
.Y(n_1118)
);

BUFx3_ASAP7_75t_L g1119 ( 
.A(n_1018),
.Y(n_1119)
);

CKINVDCx5p33_ASAP7_75t_R g1120 ( 
.A(n_1079),
.Y(n_1120)
);

AOI22xp5_ASAP7_75t_L g1121 ( 
.A1(n_1087),
.A2(n_1027),
.B1(n_1006),
.B2(n_1061),
.Y(n_1121)
);

CKINVDCx6p67_ASAP7_75t_R g1122 ( 
.A(n_1119),
.Y(n_1122)
);

AOI21xp33_ASAP7_75t_L g1123 ( 
.A1(n_1070),
.A2(n_1101),
.B(n_1073),
.Y(n_1123)
);

INVx3_ASAP7_75t_L g1124 ( 
.A(n_1068),
.Y(n_1124)
);

BUFx6f_ASAP7_75t_L g1125 ( 
.A(n_1077),
.Y(n_1125)
);

OR2x6_ASAP7_75t_L g1126 ( 
.A(n_1083),
.B(n_1034),
.Y(n_1126)
);

BUFx8_ASAP7_75t_SL g1127 ( 
.A(n_1079),
.Y(n_1127)
);

INVx2_ASAP7_75t_SL g1128 ( 
.A(n_1119),
.Y(n_1128)
);

HB1xp67_ASAP7_75t_L g1129 ( 
.A(n_1075),
.Y(n_1129)
);

AOI22xp33_ASAP7_75t_SL g1130 ( 
.A1(n_1087),
.A2(n_1048),
.B1(n_1046),
.B2(n_1059),
.Y(n_1130)
);

AND2x2_ASAP7_75t_L g1131 ( 
.A(n_1081),
.B(n_1059),
.Y(n_1131)
);

AND2x4_ASAP7_75t_L g1132 ( 
.A(n_1078),
.B(n_1092),
.Y(n_1132)
);

NAND2xp5_ASAP7_75t_L g1133 ( 
.A(n_1114),
.B(n_1033),
.Y(n_1133)
);

NAND2xp5_ASAP7_75t_L g1134 ( 
.A(n_1114),
.B(n_1055),
.Y(n_1134)
);

CKINVDCx5p33_ASAP7_75t_R g1135 ( 
.A(n_1075),
.Y(n_1135)
);

NAND3xp33_ASAP7_75t_SL g1136 ( 
.A(n_1116),
.B(n_1064),
.C(n_1065),
.Y(n_1136)
);

INVx1_ASAP7_75t_L g1137 ( 
.A(n_1067),
.Y(n_1137)
);

AOI22xp33_ASAP7_75t_L g1138 ( 
.A1(n_1116),
.A2(n_1035),
.B1(n_1012),
.B2(n_1046),
.Y(n_1138)
);

INVx2_ASAP7_75t_L g1139 ( 
.A(n_1067),
.Y(n_1139)
);

NOR2x1p5_ASAP7_75t_L g1140 ( 
.A(n_1092),
.B(n_1090),
.Y(n_1140)
);

OAI22xp33_ASAP7_75t_L g1141 ( 
.A1(n_1066),
.A2(n_1036),
.B1(n_527),
.B2(n_533),
.Y(n_1141)
);

AOI22xp33_ASAP7_75t_L g1142 ( 
.A1(n_1109),
.A2(n_528),
.B1(n_530),
.B2(n_532),
.Y(n_1142)
);

NAND2x1_ASAP7_75t_L g1143 ( 
.A(n_1088),
.B(n_1051),
.Y(n_1143)
);

INVx2_ASAP7_75t_L g1144 ( 
.A(n_1088),
.Y(n_1144)
);

AOI22xp33_ASAP7_75t_L g1145 ( 
.A1(n_1109),
.A2(n_1044),
.B1(n_1043),
.B2(n_1055),
.Y(n_1145)
);

NOR2x1_ASAP7_75t_R g1146 ( 
.A(n_1077),
.B(n_1055),
.Y(n_1146)
);

INVx1_ASAP7_75t_L g1147 ( 
.A(n_1071),
.Y(n_1147)
);

BUFx2_ASAP7_75t_L g1148 ( 
.A(n_1085),
.Y(n_1148)
);

AOI22xp33_ASAP7_75t_L g1149 ( 
.A1(n_1080),
.A2(n_1045),
.B1(n_7),
.B2(n_9),
.Y(n_1149)
);

CKINVDCx5p33_ASAP7_75t_R g1150 ( 
.A(n_1089),
.Y(n_1150)
);

OAI22xp5_ASAP7_75t_SL g1151 ( 
.A1(n_1111),
.A2(n_6),
.B1(n_9),
.B2(n_10),
.Y(n_1151)
);

INVx2_ASAP7_75t_SL g1152 ( 
.A(n_1090),
.Y(n_1152)
);

OAI21xp5_ASAP7_75t_L g1153 ( 
.A1(n_1101),
.A2(n_139),
.B(n_137),
.Y(n_1153)
);

AOI22xp33_ASAP7_75t_L g1154 ( 
.A1(n_1113),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_1154)
);

AOI22xp33_ASAP7_75t_L g1155 ( 
.A1(n_1113),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_1155)
);

AND2x2_ASAP7_75t_L g1156 ( 
.A(n_1076),
.B(n_14),
.Y(n_1156)
);

OR2x2_ASAP7_75t_L g1157 ( 
.A(n_1091),
.B(n_15),
.Y(n_1157)
);

INVxp67_ASAP7_75t_SL g1158 ( 
.A(n_1068),
.Y(n_1158)
);

INVx1_ASAP7_75t_L g1159 ( 
.A(n_1103),
.Y(n_1159)
);

AND2x2_ASAP7_75t_L g1160 ( 
.A(n_1092),
.B(n_15),
.Y(n_1160)
);

NAND2xp5_ASAP7_75t_L g1161 ( 
.A(n_1082),
.B(n_16),
.Y(n_1161)
);

INVx1_ASAP7_75t_L g1162 ( 
.A(n_1103),
.Y(n_1162)
);

INVx1_ASAP7_75t_L g1163 ( 
.A(n_1103),
.Y(n_1163)
);

INVx3_ASAP7_75t_L g1164 ( 
.A(n_1078),
.Y(n_1164)
);

BUFx6f_ASAP7_75t_L g1165 ( 
.A(n_1078),
.Y(n_1165)
);

NAND2x1p5_ASAP7_75t_L g1166 ( 
.A(n_1099),
.B(n_1107),
.Y(n_1166)
);

INVx3_ASAP7_75t_L g1167 ( 
.A(n_1105),
.Y(n_1167)
);

BUFx3_ASAP7_75t_L g1168 ( 
.A(n_1106),
.Y(n_1168)
);

INVx1_ASAP7_75t_L g1169 ( 
.A(n_1099),
.Y(n_1169)
);

INVx1_ASAP7_75t_L g1170 ( 
.A(n_1106),
.Y(n_1170)
);

AOI22xp33_ASAP7_75t_SL g1171 ( 
.A1(n_1104),
.A2(n_16),
.B1(n_18),
.B2(n_19),
.Y(n_1171)
);

BUFx3_ASAP7_75t_L g1172 ( 
.A(n_1111),
.Y(n_1172)
);

OR2x6_ASAP7_75t_SL g1173 ( 
.A(n_1084),
.B(n_18),
.Y(n_1173)
);

INVx1_ASAP7_75t_L g1174 ( 
.A(n_1072),
.Y(n_1174)
);

AOI22xp33_ASAP7_75t_SL g1175 ( 
.A1(n_1073),
.A2(n_20),
.B1(n_21),
.B2(n_22),
.Y(n_1175)
);

AOI211x1_ASAP7_75t_L g1176 ( 
.A1(n_1074),
.A2(n_21),
.B(n_22),
.C(n_23),
.Y(n_1176)
);

OAI22xp5_ASAP7_75t_L g1177 ( 
.A1(n_1100),
.A2(n_24),
.B1(n_25),
.B2(n_26),
.Y(n_1177)
);

AOI21xp5_ASAP7_75t_L g1178 ( 
.A1(n_1073),
.A2(n_354),
.B(n_143),
.Y(n_1178)
);

CKINVDCx20_ASAP7_75t_R g1179 ( 
.A(n_1105),
.Y(n_1179)
);

AND2x2_ASAP7_75t_L g1180 ( 
.A(n_1131),
.B(n_1072),
.Y(n_1180)
);

AND2x2_ASAP7_75t_L g1181 ( 
.A(n_1160),
.B(n_1072),
.Y(n_1181)
);

AOI22xp33_ASAP7_75t_SL g1182 ( 
.A1(n_1153),
.A2(n_1151),
.B1(n_1177),
.B2(n_1161),
.Y(n_1182)
);

AOI222xp33_ASAP7_75t_L g1183 ( 
.A1(n_1177),
.A2(n_27),
.B1(n_28),
.B2(n_29),
.C1(n_30),
.C2(n_31),
.Y(n_1183)
);

INVx1_ASAP7_75t_L g1184 ( 
.A(n_1147),
.Y(n_1184)
);

AOI22xp33_ASAP7_75t_L g1185 ( 
.A1(n_1130),
.A2(n_1096),
.B1(n_1097),
.B2(n_1110),
.Y(n_1185)
);

AOI22xp33_ASAP7_75t_L g1186 ( 
.A1(n_1153),
.A2(n_1110),
.B1(n_1097),
.B2(n_1117),
.Y(n_1186)
);

AOI22xp33_ASAP7_75t_L g1187 ( 
.A1(n_1154),
.A2(n_1110),
.B1(n_1097),
.B2(n_1117),
.Y(n_1187)
);

OAI22xp33_ASAP7_75t_L g1188 ( 
.A1(n_1121),
.A2(n_1102),
.B1(n_1112),
.B2(n_1117),
.Y(n_1188)
);

AOI22xp33_ASAP7_75t_SL g1189 ( 
.A1(n_1161),
.A2(n_1112),
.B1(n_1115),
.B2(n_1102),
.Y(n_1189)
);

INVx1_ASAP7_75t_L g1190 ( 
.A(n_1137),
.Y(n_1190)
);

INVx2_ASAP7_75t_L g1191 ( 
.A(n_1139),
.Y(n_1191)
);

BUFx2_ASAP7_75t_L g1192 ( 
.A(n_1135),
.Y(n_1192)
);

INVx1_ASAP7_75t_L g1193 ( 
.A(n_1144),
.Y(n_1193)
);

AOI22xp33_ASAP7_75t_L g1194 ( 
.A1(n_1155),
.A2(n_1069),
.B1(n_1098),
.B2(n_1118),
.Y(n_1194)
);

INVx1_ASAP7_75t_L g1195 ( 
.A(n_1134),
.Y(n_1195)
);

BUFx2_ASAP7_75t_L g1196 ( 
.A(n_1148),
.Y(n_1196)
);

NAND2xp5_ASAP7_75t_L g1197 ( 
.A(n_1133),
.B(n_1072),
.Y(n_1197)
);

OAI221xp5_ASAP7_75t_L g1198 ( 
.A1(n_1171),
.A2(n_27),
.B1(n_28),
.B2(n_29),
.C(n_31),
.Y(n_1198)
);

AOI221xp5_ASAP7_75t_L g1199 ( 
.A1(n_1176),
.A2(n_32),
.B1(n_33),
.B2(n_35),
.C(n_36),
.Y(n_1199)
);

AOI21xp5_ASAP7_75t_L g1200 ( 
.A1(n_1123),
.A2(n_1093),
.B(n_1094),
.Y(n_1200)
);

BUFx3_ASAP7_75t_L g1201 ( 
.A(n_1179),
.Y(n_1201)
);

INVx2_ASAP7_75t_L g1202 ( 
.A(n_1169),
.Y(n_1202)
);

AOI22xp33_ASAP7_75t_L g1203 ( 
.A1(n_1136),
.A2(n_1108),
.B1(n_1105),
.B2(n_1095),
.Y(n_1203)
);

AOI21xp5_ASAP7_75t_L g1204 ( 
.A1(n_1123),
.A2(n_1086),
.B(n_144),
.Y(n_1204)
);

BUFx6f_ASAP7_75t_L g1205 ( 
.A(n_1125),
.Y(n_1205)
);

INVx1_ASAP7_75t_L g1206 ( 
.A(n_1134),
.Y(n_1206)
);

AOI22xp33_ASAP7_75t_L g1207 ( 
.A1(n_1126),
.A2(n_32),
.B1(n_33),
.B2(n_35),
.Y(n_1207)
);

AOI221xp5_ASAP7_75t_L g1208 ( 
.A1(n_1175),
.A2(n_36),
.B1(n_37),
.B2(n_38),
.C(n_39),
.Y(n_1208)
);

AOI21xp5_ASAP7_75t_L g1209 ( 
.A1(n_1133),
.A2(n_221),
.B(n_351),
.Y(n_1209)
);

INVx1_ASAP7_75t_L g1210 ( 
.A(n_1170),
.Y(n_1210)
);

AOI22xp33_ASAP7_75t_SL g1211 ( 
.A1(n_1172),
.A2(n_37),
.B1(n_38),
.B2(n_39),
.Y(n_1211)
);

AOI22xp33_ASAP7_75t_SL g1212 ( 
.A1(n_1132),
.A2(n_40),
.B1(n_41),
.B2(n_42),
.Y(n_1212)
);

NAND2xp5_ASAP7_75t_L g1213 ( 
.A(n_1174),
.B(n_40),
.Y(n_1213)
);

OAI221xp5_ASAP7_75t_L g1214 ( 
.A1(n_1149),
.A2(n_1138),
.B1(n_1142),
.B2(n_1126),
.C(n_1145),
.Y(n_1214)
);

BUFx3_ASAP7_75t_L g1215 ( 
.A(n_1122),
.Y(n_1215)
);

AND2x2_ASAP7_75t_L g1216 ( 
.A(n_1159),
.B(n_142),
.Y(n_1216)
);

OR2x2_ASAP7_75t_L g1217 ( 
.A(n_1129),
.B(n_41),
.Y(n_1217)
);

AOI22xp33_ASAP7_75t_L g1218 ( 
.A1(n_1126),
.A2(n_43),
.B1(n_45),
.B2(n_46),
.Y(n_1218)
);

AOI22xp33_ASAP7_75t_L g1219 ( 
.A1(n_1140),
.A2(n_43),
.B1(n_45),
.B2(n_46),
.Y(n_1219)
);

INVx1_ASAP7_75t_L g1220 ( 
.A(n_1162),
.Y(n_1220)
);

OAI22xp5_ASAP7_75t_L g1221 ( 
.A1(n_1173),
.A2(n_47),
.B1(n_49),
.B2(n_51),
.Y(n_1221)
);

AND2x4_ASAP7_75t_L g1222 ( 
.A(n_1132),
.B(n_145),
.Y(n_1222)
);

CKINVDCx20_ASAP7_75t_R g1223 ( 
.A(n_1127),
.Y(n_1223)
);

OAI22xp33_ASAP7_75t_L g1224 ( 
.A1(n_1150),
.A2(n_47),
.B1(n_51),
.B2(n_52),
.Y(n_1224)
);

NAND2xp5_ASAP7_75t_SL g1225 ( 
.A(n_1165),
.B(n_147),
.Y(n_1225)
);

OR2x6_ASAP7_75t_SL g1226 ( 
.A(n_1120),
.B(n_52),
.Y(n_1226)
);

OAI211xp5_ASAP7_75t_L g1227 ( 
.A1(n_1156),
.A2(n_53),
.B(n_54),
.C(n_55),
.Y(n_1227)
);

A2O1A1Ixp33_ASAP7_75t_L g1228 ( 
.A1(n_1178),
.A2(n_54),
.B(n_56),
.C(n_58),
.Y(n_1228)
);

OAI22xp5_ASAP7_75t_L g1229 ( 
.A1(n_1157),
.A2(n_58),
.B1(n_59),
.B2(n_60),
.Y(n_1229)
);

INVx2_ASAP7_75t_L g1230 ( 
.A(n_1163),
.Y(n_1230)
);

OAI22xp5_ASAP7_75t_L g1231 ( 
.A1(n_1167),
.A2(n_59),
.B1(n_61),
.B2(n_62),
.Y(n_1231)
);

INVx2_ASAP7_75t_L g1232 ( 
.A(n_1166),
.Y(n_1232)
);

AO31x2_ASAP7_75t_L g1233 ( 
.A1(n_1146),
.A2(n_239),
.A3(n_345),
.B(n_148),
.Y(n_1233)
);

INVx3_ASAP7_75t_L g1234 ( 
.A(n_1165),
.Y(n_1234)
);

INVx2_ASAP7_75t_L g1235 ( 
.A(n_1166),
.Y(n_1235)
);

AOI22xp33_ASAP7_75t_L g1236 ( 
.A1(n_1182),
.A2(n_1164),
.B1(n_1141),
.B2(n_1165),
.Y(n_1236)
);

NOR2xp33_ASAP7_75t_L g1237 ( 
.A(n_1192),
.B(n_1152),
.Y(n_1237)
);

INVx2_ASAP7_75t_L g1238 ( 
.A(n_1184),
.Y(n_1238)
);

AND2x2_ASAP7_75t_L g1239 ( 
.A(n_1180),
.B(n_1164),
.Y(n_1239)
);

INVx4_ASAP7_75t_R g1240 ( 
.A(n_1215),
.Y(n_1240)
);

INVx1_ASAP7_75t_L g1241 ( 
.A(n_1195),
.Y(n_1241)
);

HB1xp67_ASAP7_75t_L g1242 ( 
.A(n_1196),
.Y(n_1242)
);

INVx3_ASAP7_75t_L g1243 ( 
.A(n_1232),
.Y(n_1243)
);

INVx4_ASAP7_75t_L g1244 ( 
.A(n_1205),
.Y(n_1244)
);

AND2x4_ASAP7_75t_L g1245 ( 
.A(n_1190),
.B(n_1168),
.Y(n_1245)
);

BUFx3_ASAP7_75t_L g1246 ( 
.A(n_1205),
.Y(n_1246)
);

AO31x2_ASAP7_75t_L g1247 ( 
.A1(n_1200),
.A2(n_1143),
.A3(n_1158),
.B(n_63),
.Y(n_1247)
);

INVx1_ASAP7_75t_L g1248 ( 
.A(n_1206),
.Y(n_1248)
);

INVx1_ASAP7_75t_L g1249 ( 
.A(n_1202),
.Y(n_1249)
);

INVx1_ASAP7_75t_L g1250 ( 
.A(n_1197),
.Y(n_1250)
);

INVx2_ASAP7_75t_L g1251 ( 
.A(n_1210),
.Y(n_1251)
);

BUFx3_ASAP7_75t_L g1252 ( 
.A(n_1205),
.Y(n_1252)
);

AND2x2_ASAP7_75t_L g1253 ( 
.A(n_1181),
.B(n_1197),
.Y(n_1253)
);

AND2x2_ASAP7_75t_L g1254 ( 
.A(n_1220),
.B(n_1124),
.Y(n_1254)
);

AOI22xp33_ASAP7_75t_L g1255 ( 
.A1(n_1198),
.A2(n_1124),
.B1(n_1167),
.B2(n_1128),
.Y(n_1255)
);

OR2x2_ASAP7_75t_L g1256 ( 
.A(n_1213),
.B(n_1125),
.Y(n_1256)
);

AOI22xp33_ASAP7_75t_L g1257 ( 
.A1(n_1198),
.A2(n_1125),
.B1(n_63),
.B2(n_61),
.Y(n_1257)
);

INVx2_ASAP7_75t_L g1258 ( 
.A(n_1193),
.Y(n_1258)
);

OR2x2_ASAP7_75t_L g1259 ( 
.A(n_1213),
.B(n_152),
.Y(n_1259)
);

AND2x4_ASAP7_75t_L g1260 ( 
.A(n_1235),
.B(n_155),
.Y(n_1260)
);

AND2x4_ASAP7_75t_L g1261 ( 
.A(n_1230),
.B(n_156),
.Y(n_1261)
);

BUFx2_ASAP7_75t_L g1262 ( 
.A(n_1233),
.Y(n_1262)
);

NOR2x1_ASAP7_75t_L g1263 ( 
.A(n_1188),
.B(n_159),
.Y(n_1263)
);

OAI22xp5_ASAP7_75t_L g1264 ( 
.A1(n_1219),
.A2(n_161),
.B1(n_163),
.B2(n_165),
.Y(n_1264)
);

INVx1_ASAP7_75t_L g1265 ( 
.A(n_1191),
.Y(n_1265)
);

NAND2xp5_ASAP7_75t_L g1266 ( 
.A(n_1217),
.B(n_167),
.Y(n_1266)
);

OR2x2_ASAP7_75t_L g1267 ( 
.A(n_1186),
.B(n_168),
.Y(n_1267)
);

AND2x2_ASAP7_75t_L g1268 ( 
.A(n_1185),
.B(n_169),
.Y(n_1268)
);

AND2x2_ASAP7_75t_L g1269 ( 
.A(n_1233),
.B(n_170),
.Y(n_1269)
);

BUFx6f_ASAP7_75t_SL g1270 ( 
.A(n_1222),
.Y(n_1270)
);

HB1xp67_ASAP7_75t_L g1271 ( 
.A(n_1234),
.Y(n_1271)
);

OR2x2_ASAP7_75t_L g1272 ( 
.A(n_1187),
.B(n_171),
.Y(n_1272)
);

INVx2_ASAP7_75t_L g1273 ( 
.A(n_1233),
.Y(n_1273)
);

AND2x2_ASAP7_75t_L g1274 ( 
.A(n_1234),
.B(n_173),
.Y(n_1274)
);

BUFx3_ASAP7_75t_L g1275 ( 
.A(n_1201),
.Y(n_1275)
);

AND2x2_ASAP7_75t_L g1276 ( 
.A(n_1189),
.B(n_175),
.Y(n_1276)
);

AND2x4_ASAP7_75t_L g1277 ( 
.A(n_1204),
.B(n_180),
.Y(n_1277)
);

AO21x2_ASAP7_75t_L g1278 ( 
.A1(n_1228),
.A2(n_182),
.B(n_183),
.Y(n_1278)
);

INVx2_ASAP7_75t_L g1279 ( 
.A(n_1216),
.Y(n_1279)
);

AOI211xp5_ASAP7_75t_L g1280 ( 
.A1(n_1276),
.A2(n_1221),
.B(n_1224),
.C(n_1231),
.Y(n_1280)
);

NOR4xp25_ASAP7_75t_SL g1281 ( 
.A(n_1262),
.B(n_1214),
.C(n_1208),
.D(n_1199),
.Y(n_1281)
);

AOI33xp33_ASAP7_75t_L g1282 ( 
.A1(n_1257),
.A2(n_1211),
.A3(n_1212),
.B1(n_1207),
.B2(n_1218),
.B3(n_1226),
.Y(n_1282)
);

INVx2_ASAP7_75t_L g1283 ( 
.A(n_1238),
.Y(n_1283)
);

AND2x4_ASAP7_75t_L g1284 ( 
.A(n_1238),
.B(n_1222),
.Y(n_1284)
);

INVx1_ASAP7_75t_L g1285 ( 
.A(n_1251),
.Y(n_1285)
);

AOI33xp33_ASAP7_75t_L g1286 ( 
.A1(n_1255),
.A2(n_1221),
.A3(n_1183),
.B1(n_1203),
.B2(n_1227),
.B3(n_1231),
.Y(n_1286)
);

OAI22xp5_ASAP7_75t_SL g1287 ( 
.A1(n_1263),
.A2(n_1223),
.B1(n_1214),
.B2(n_1229),
.Y(n_1287)
);

OAI33xp33_ASAP7_75t_L g1288 ( 
.A1(n_1250),
.A2(n_1229),
.A3(n_1183),
.B1(n_1225),
.B2(n_1209),
.B3(n_1194),
.Y(n_1288)
);

INVx2_ASAP7_75t_L g1289 ( 
.A(n_1258),
.Y(n_1289)
);

AOI221xp5_ASAP7_75t_L g1290 ( 
.A1(n_1242),
.A2(n_352),
.B1(n_187),
.B2(n_188),
.C(n_189),
.Y(n_1290)
);

INVx1_ASAP7_75t_L g1291 ( 
.A(n_1251),
.Y(n_1291)
);

INVx2_ASAP7_75t_L g1292 ( 
.A(n_1258),
.Y(n_1292)
);

AO22x1_ASAP7_75t_L g1293 ( 
.A1(n_1263),
.A2(n_186),
.B1(n_191),
.B2(n_192),
.Y(n_1293)
);

INVx1_ASAP7_75t_L g1294 ( 
.A(n_1249),
.Y(n_1294)
);

AOI22xp33_ASAP7_75t_L g1295 ( 
.A1(n_1278),
.A2(n_1268),
.B1(n_1276),
.B2(n_1277),
.Y(n_1295)
);

OAI31xp33_ASAP7_75t_L g1296 ( 
.A1(n_1264),
.A2(n_199),
.A3(n_202),
.B(n_203),
.Y(n_1296)
);

NAND3xp33_ASAP7_75t_L g1297 ( 
.A(n_1259),
.B(n_204),
.C(n_205),
.Y(n_1297)
);

OAI22xp5_ASAP7_75t_L g1298 ( 
.A1(n_1236),
.A2(n_1270),
.B1(n_1256),
.B2(n_1272),
.Y(n_1298)
);

INVx2_ASAP7_75t_L g1299 ( 
.A(n_1249),
.Y(n_1299)
);

INVx1_ASAP7_75t_L g1300 ( 
.A(n_1241),
.Y(n_1300)
);

INVx2_ASAP7_75t_SL g1301 ( 
.A(n_1245),
.Y(n_1301)
);

BUFx2_ASAP7_75t_L g1302 ( 
.A(n_1245),
.Y(n_1302)
);

HB1xp67_ASAP7_75t_L g1303 ( 
.A(n_1245),
.Y(n_1303)
);

INVx1_ASAP7_75t_L g1304 ( 
.A(n_1241),
.Y(n_1304)
);

AND2x2_ASAP7_75t_L g1305 ( 
.A(n_1253),
.B(n_206),
.Y(n_1305)
);

AO21x2_ASAP7_75t_L g1306 ( 
.A1(n_1273),
.A2(n_207),
.B(n_210),
.Y(n_1306)
);

AOI221xp5_ASAP7_75t_L g1307 ( 
.A1(n_1266),
.A2(n_214),
.B1(n_215),
.B2(n_217),
.C(n_222),
.Y(n_1307)
);

NAND2x1p5_ASAP7_75t_L g1308 ( 
.A(n_1284),
.B(n_1262),
.Y(n_1308)
);

INVx1_ASAP7_75t_L g1309 ( 
.A(n_1299),
.Y(n_1309)
);

AND2x2_ASAP7_75t_L g1310 ( 
.A(n_1302),
.B(n_1253),
.Y(n_1310)
);

INVx1_ASAP7_75t_L g1311 ( 
.A(n_1299),
.Y(n_1311)
);

INVx1_ASAP7_75t_L g1312 ( 
.A(n_1285),
.Y(n_1312)
);

INVx1_ASAP7_75t_SL g1313 ( 
.A(n_1302),
.Y(n_1313)
);

NOR2xp33_ASAP7_75t_L g1314 ( 
.A(n_1301),
.B(n_1275),
.Y(n_1314)
);

AND2x2_ASAP7_75t_L g1315 ( 
.A(n_1303),
.B(n_1239),
.Y(n_1315)
);

OR2x2_ASAP7_75t_L g1316 ( 
.A(n_1301),
.B(n_1250),
.Y(n_1316)
);

INVx1_ASAP7_75t_L g1317 ( 
.A(n_1291),
.Y(n_1317)
);

NAND2xp5_ASAP7_75t_L g1318 ( 
.A(n_1289),
.B(n_1248),
.Y(n_1318)
);

AND2x2_ASAP7_75t_L g1319 ( 
.A(n_1289),
.B(n_1239),
.Y(n_1319)
);

INVx4_ASAP7_75t_L g1320 ( 
.A(n_1305),
.Y(n_1320)
);

AND2x2_ASAP7_75t_L g1321 ( 
.A(n_1292),
.B(n_1275),
.Y(n_1321)
);

AND2x4_ASAP7_75t_L g1322 ( 
.A(n_1284),
.B(n_1245),
.Y(n_1322)
);

AOI32xp33_ASAP7_75t_L g1323 ( 
.A1(n_1280),
.A2(n_1295),
.A3(n_1298),
.B1(n_1269),
.B2(n_1305),
.Y(n_1323)
);

NAND2xp5_ASAP7_75t_SL g1324 ( 
.A(n_1287),
.B(n_1256),
.Y(n_1324)
);

NOR3xp33_ASAP7_75t_L g1325 ( 
.A(n_1293),
.B(n_1269),
.C(n_1268),
.Y(n_1325)
);

NAND2x1_ASAP7_75t_L g1326 ( 
.A(n_1292),
.B(n_1240),
.Y(n_1326)
);

INVx2_ASAP7_75t_SL g1327 ( 
.A(n_1321),
.Y(n_1327)
);

INVx1_ASAP7_75t_SL g1328 ( 
.A(n_1313),
.Y(n_1328)
);

INVx1_ASAP7_75t_L g1329 ( 
.A(n_1312),
.Y(n_1329)
);

INVx1_ASAP7_75t_L g1330 ( 
.A(n_1317),
.Y(n_1330)
);

INVxp67_ASAP7_75t_L g1331 ( 
.A(n_1324),
.Y(n_1331)
);

AND2x4_ASAP7_75t_L g1332 ( 
.A(n_1322),
.B(n_1284),
.Y(n_1332)
);

NAND2xp5_ASAP7_75t_L g1333 ( 
.A(n_1309),
.B(n_1300),
.Y(n_1333)
);

OAI21xp33_ASAP7_75t_L g1334 ( 
.A1(n_1323),
.A2(n_1286),
.B(n_1282),
.Y(n_1334)
);

AND2x4_ASAP7_75t_L g1335 ( 
.A(n_1322),
.B(n_1294),
.Y(n_1335)
);

INVx2_ASAP7_75t_L g1336 ( 
.A(n_1316),
.Y(n_1336)
);

AND2x2_ASAP7_75t_L g1337 ( 
.A(n_1310),
.B(n_1283),
.Y(n_1337)
);

NAND2xp5_ASAP7_75t_L g1338 ( 
.A(n_1331),
.B(n_1311),
.Y(n_1338)
);

INVx2_ASAP7_75t_L g1339 ( 
.A(n_1335),
.Y(n_1339)
);

INVx1_ASAP7_75t_L g1340 ( 
.A(n_1329),
.Y(n_1340)
);

INVx4_ASAP7_75t_L g1341 ( 
.A(n_1332),
.Y(n_1341)
);

AND2x2_ASAP7_75t_L g1342 ( 
.A(n_1332),
.B(n_1315),
.Y(n_1342)
);

INVx1_ASAP7_75t_L g1343 ( 
.A(n_1330),
.Y(n_1343)
);

OR2x6_ASAP7_75t_L g1344 ( 
.A(n_1331),
.B(n_1293),
.Y(n_1344)
);

AND2x2_ASAP7_75t_L g1345 ( 
.A(n_1335),
.B(n_1319),
.Y(n_1345)
);

INVx2_ASAP7_75t_L g1346 ( 
.A(n_1327),
.Y(n_1346)
);

AND2x4_ASAP7_75t_L g1347 ( 
.A(n_1328),
.B(n_1320),
.Y(n_1347)
);

NAND2xp5_ASAP7_75t_L g1348 ( 
.A(n_1328),
.B(n_1318),
.Y(n_1348)
);

INVx1_ASAP7_75t_L g1349 ( 
.A(n_1333),
.Y(n_1349)
);

INVx2_ASAP7_75t_L g1350 ( 
.A(n_1336),
.Y(n_1350)
);

INVx2_ASAP7_75t_L g1351 ( 
.A(n_1333),
.Y(n_1351)
);

INVxp67_ASAP7_75t_SL g1352 ( 
.A(n_1347),
.Y(n_1352)
);

INVx1_ASAP7_75t_L g1353 ( 
.A(n_1340),
.Y(n_1353)
);

OR2x2_ASAP7_75t_L g1354 ( 
.A(n_1350),
.B(n_1337),
.Y(n_1354)
);

INVx1_ASAP7_75t_L g1355 ( 
.A(n_1343),
.Y(n_1355)
);

INVx1_ASAP7_75t_L g1356 ( 
.A(n_1338),
.Y(n_1356)
);

INVx2_ASAP7_75t_L g1357 ( 
.A(n_1341),
.Y(n_1357)
);

INVx1_ASAP7_75t_L g1358 ( 
.A(n_1338),
.Y(n_1358)
);

NAND2xp5_ASAP7_75t_L g1359 ( 
.A(n_1349),
.B(n_1351),
.Y(n_1359)
);

INVx1_ASAP7_75t_L g1360 ( 
.A(n_1351),
.Y(n_1360)
);

OAI22xp33_ASAP7_75t_L g1361 ( 
.A1(n_1352),
.A2(n_1344),
.B1(n_1341),
.B2(n_1339),
.Y(n_1361)
);

NOR2xp33_ASAP7_75t_L g1362 ( 
.A(n_1357),
.B(n_1334),
.Y(n_1362)
);

AOI32xp33_ASAP7_75t_L g1363 ( 
.A1(n_1356),
.A2(n_1325),
.A3(n_1347),
.B1(n_1346),
.B2(n_1344),
.Y(n_1363)
);

OAI31xp33_ASAP7_75t_L g1364 ( 
.A1(n_1358),
.A2(n_1325),
.A3(n_1344),
.B(n_1297),
.Y(n_1364)
);

A2O1A1Ixp33_ASAP7_75t_L g1365 ( 
.A1(n_1353),
.A2(n_1282),
.B(n_1286),
.C(n_1326),
.Y(n_1365)
);

NOR2xp33_ASAP7_75t_SL g1366 ( 
.A(n_1355),
.B(n_1288),
.Y(n_1366)
);

AO21x1_ASAP7_75t_L g1367 ( 
.A1(n_1360),
.A2(n_1348),
.B(n_1237),
.Y(n_1367)
);

AND2x2_ASAP7_75t_L g1368 ( 
.A(n_1362),
.B(n_1342),
.Y(n_1368)
);

AND2x2_ASAP7_75t_SL g1369 ( 
.A(n_1366),
.B(n_1364),
.Y(n_1369)
);

INVx1_ASAP7_75t_SL g1370 ( 
.A(n_1363),
.Y(n_1370)
);

OAI211xp5_ASAP7_75t_SL g1371 ( 
.A1(n_1361),
.A2(n_1359),
.B(n_1354),
.C(n_1290),
.Y(n_1371)
);

A2O1A1Ixp33_ASAP7_75t_L g1372 ( 
.A1(n_1365),
.A2(n_1359),
.B(n_1348),
.C(n_1314),
.Y(n_1372)
);

AOI22xp33_ASAP7_75t_SL g1373 ( 
.A1(n_1367),
.A2(n_1270),
.B1(n_1320),
.B2(n_1278),
.Y(n_1373)
);

NAND2xp5_ASAP7_75t_L g1374 ( 
.A(n_1362),
.B(n_1345),
.Y(n_1374)
);

INVx1_ASAP7_75t_L g1375 ( 
.A(n_1368),
.Y(n_1375)
);

INVx1_ASAP7_75t_L g1376 ( 
.A(n_1374),
.Y(n_1376)
);

NAND2xp5_ASAP7_75t_L g1377 ( 
.A(n_1369),
.B(n_1313),
.Y(n_1377)
);

NOR2xp33_ASAP7_75t_L g1378 ( 
.A(n_1370),
.B(n_1318),
.Y(n_1378)
);

OAI211xp5_ASAP7_75t_L g1379 ( 
.A1(n_1372),
.A2(n_1281),
.B(n_1296),
.C(n_1307),
.Y(n_1379)
);

NAND2xp5_ASAP7_75t_L g1380 ( 
.A(n_1373),
.B(n_1304),
.Y(n_1380)
);

NAND2xp5_ASAP7_75t_L g1381 ( 
.A(n_1371),
.B(n_1308),
.Y(n_1381)
);

NAND3xp33_ASAP7_75t_SL g1382 ( 
.A(n_1370),
.B(n_1259),
.C(n_1267),
.Y(n_1382)
);

AOI211xp5_ASAP7_75t_L g1383 ( 
.A1(n_1370),
.A2(n_1272),
.B(n_1267),
.C(n_1277),
.Y(n_1383)
);

OAI221xp5_ASAP7_75t_L g1384 ( 
.A1(n_1379),
.A2(n_1308),
.B1(n_1240),
.B2(n_1271),
.C(n_1265),
.Y(n_1384)
);

INVx1_ASAP7_75t_L g1385 ( 
.A(n_1375),
.Y(n_1385)
);

OAI211xp5_ASAP7_75t_L g1386 ( 
.A1(n_1381),
.A2(n_1274),
.B(n_1244),
.C(n_1273),
.Y(n_1386)
);

NOR3xp33_ASAP7_75t_L g1387 ( 
.A(n_1376),
.B(n_1277),
.C(n_1274),
.Y(n_1387)
);

AOI211xp5_ASAP7_75t_L g1388 ( 
.A1(n_1377),
.A2(n_1277),
.B(n_1261),
.C(n_1260),
.Y(n_1388)
);

INVx1_ASAP7_75t_L g1389 ( 
.A(n_1378),
.Y(n_1389)
);

NAND2xp5_ASAP7_75t_L g1390 ( 
.A(n_1383),
.B(n_1283),
.Y(n_1390)
);

OAI21xp5_ASAP7_75t_SL g1391 ( 
.A1(n_1382),
.A2(n_1261),
.B(n_1260),
.Y(n_1391)
);

AOI21xp5_ASAP7_75t_L g1392 ( 
.A1(n_1389),
.A2(n_1380),
.B(n_1278),
.Y(n_1392)
);

NAND2xp5_ASAP7_75t_L g1393 ( 
.A(n_1385),
.B(n_1387),
.Y(n_1393)
);

BUFx2_ASAP7_75t_R g1394 ( 
.A(n_1390),
.Y(n_1394)
);

OAI21xp5_ASAP7_75t_L g1395 ( 
.A1(n_1384),
.A2(n_1261),
.B(n_1260),
.Y(n_1395)
);

BUFx2_ASAP7_75t_L g1396 ( 
.A(n_1391),
.Y(n_1396)
);

AOI22xp5_ASAP7_75t_L g1397 ( 
.A1(n_1386),
.A2(n_1270),
.B1(n_1246),
.B2(n_1244),
.Y(n_1397)
);

AOI22xp5_ASAP7_75t_L g1398 ( 
.A1(n_1388),
.A2(n_1246),
.B1(n_1244),
.B2(n_1306),
.Y(n_1398)
);

XOR2x2_ASAP7_75t_L g1399 ( 
.A(n_1389),
.B(n_1261),
.Y(n_1399)
);

AND3x4_ASAP7_75t_L g1400 ( 
.A(n_1394),
.B(n_1252),
.C(n_1260),
.Y(n_1400)
);

OR2x2_ASAP7_75t_L g1401 ( 
.A(n_1393),
.B(n_1247),
.Y(n_1401)
);

NAND2xp5_ASAP7_75t_L g1402 ( 
.A(n_1396),
.B(n_1248),
.Y(n_1402)
);

INVx1_ASAP7_75t_L g1403 ( 
.A(n_1399),
.Y(n_1403)
);

AND2x2_ASAP7_75t_L g1404 ( 
.A(n_1397),
.B(n_1252),
.Y(n_1404)
);

NAND4xp25_ASAP7_75t_L g1405 ( 
.A(n_1392),
.B(n_1252),
.C(n_1244),
.D(n_1279),
.Y(n_1405)
);

AOI221xp5_ASAP7_75t_L g1406 ( 
.A1(n_1398),
.A2(n_1306),
.B1(n_1265),
.B2(n_1243),
.C(n_1254),
.Y(n_1406)
);

NOR3xp33_ASAP7_75t_SL g1407 ( 
.A(n_1395),
.B(n_1306),
.C(n_226),
.Y(n_1407)
);

INVx2_ASAP7_75t_L g1408 ( 
.A(n_1400),
.Y(n_1408)
);

NAND2xp5_ASAP7_75t_SL g1409 ( 
.A(n_1407),
.B(n_1243),
.Y(n_1409)
);

NAND3xp33_ASAP7_75t_SL g1410 ( 
.A(n_1403),
.B(n_1401),
.C(n_1402),
.Y(n_1410)
);

INVx1_ASAP7_75t_L g1411 ( 
.A(n_1404),
.Y(n_1411)
);

AO22x2_ASAP7_75t_L g1412 ( 
.A1(n_1405),
.A2(n_1243),
.B1(n_1279),
.B2(n_1254),
.Y(n_1412)
);

NAND5xp2_ASAP7_75t_L g1413 ( 
.A(n_1406),
.B(n_1247),
.C(n_227),
.D(n_228),
.E(n_229),
.Y(n_1413)
);

A2O1A1Ixp33_ASAP7_75t_L g1414 ( 
.A1(n_1407),
.A2(n_1247),
.B(n_230),
.C(n_231),
.Y(n_1414)
);

OAI221xp5_ASAP7_75t_L g1415 ( 
.A1(n_1407),
.A2(n_1247),
.B1(n_232),
.B2(n_233),
.C(n_236),
.Y(n_1415)
);

OAI221xp5_ASAP7_75t_L g1416 ( 
.A1(n_1414),
.A2(n_1247),
.B1(n_240),
.B2(n_241),
.C(n_245),
.Y(n_1416)
);

OAI222xp33_ASAP7_75t_L g1417 ( 
.A1(n_1411),
.A2(n_224),
.B1(n_247),
.B2(n_249),
.C1(n_250),
.C2(n_252),
.Y(n_1417)
);

AOI21xp5_ASAP7_75t_L g1418 ( 
.A1(n_1410),
.A2(n_255),
.B(n_256),
.Y(n_1418)
);

NAND2xp5_ASAP7_75t_L g1419 ( 
.A(n_1408),
.B(n_257),
.Y(n_1419)
);

OAI22xp5_ASAP7_75t_L g1420 ( 
.A1(n_1415),
.A2(n_261),
.B1(n_262),
.B2(n_265),
.Y(n_1420)
);

INVx1_ASAP7_75t_L g1421 ( 
.A(n_1409),
.Y(n_1421)
);

AND2x4_ASAP7_75t_L g1422 ( 
.A(n_1412),
.B(n_268),
.Y(n_1422)
);

INVx1_ASAP7_75t_L g1423 ( 
.A(n_1419),
.Y(n_1423)
);

AOI22xp5_ASAP7_75t_SL g1424 ( 
.A1(n_1421),
.A2(n_1418),
.B1(n_1420),
.B2(n_1422),
.Y(n_1424)
);

INVx1_ASAP7_75t_L g1425 ( 
.A(n_1416),
.Y(n_1425)
);

A2O1A1Ixp33_ASAP7_75t_L g1426 ( 
.A1(n_1417),
.A2(n_1413),
.B(n_272),
.C(n_273),
.Y(n_1426)
);

INVx1_ASAP7_75t_L g1427 ( 
.A(n_1424),
.Y(n_1427)
);

AOI22xp33_ASAP7_75t_L g1428 ( 
.A1(n_1425),
.A2(n_270),
.B1(n_274),
.B2(n_276),
.Y(n_1428)
);

INVx1_ASAP7_75t_L g1429 ( 
.A(n_1427),
.Y(n_1429)
);

INVx2_ASAP7_75t_L g1430 ( 
.A(n_1428),
.Y(n_1430)
);

AOI21xp5_ASAP7_75t_L g1431 ( 
.A1(n_1429),
.A2(n_1423),
.B(n_1430),
.Y(n_1431)
);

AOI21xp5_ASAP7_75t_L g1432 ( 
.A1(n_1429),
.A2(n_1426),
.B(n_280),
.Y(n_1432)
);

INVx1_ASAP7_75t_L g1433 ( 
.A(n_1431),
.Y(n_1433)
);

OAI22xp5_ASAP7_75t_L g1434 ( 
.A1(n_1432),
.A2(n_278),
.B1(n_290),
.B2(n_292),
.Y(n_1434)
);

AOI222xp33_ASAP7_75t_L g1435 ( 
.A1(n_1431),
.A2(n_295),
.B1(n_297),
.B2(n_302),
.C1(n_305),
.C2(n_307),
.Y(n_1435)
);

AOI322xp5_ASAP7_75t_L g1436 ( 
.A1(n_1433),
.A2(n_313),
.A3(n_315),
.B1(n_319),
.B2(n_320),
.C1(n_326),
.C2(n_329),
.Y(n_1436)
);

AOI22xp5_ASAP7_75t_L g1437 ( 
.A1(n_1436),
.A2(n_1434),
.B1(n_1435),
.B2(n_336),
.Y(n_1437)
);

AOI211xp5_ASAP7_75t_L g1438 ( 
.A1(n_1437),
.A2(n_331),
.B(n_333),
.C(n_339),
.Y(n_1438)
);


endmodule