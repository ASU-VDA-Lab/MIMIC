module fake_jpeg_23446_n_112 (n_3, n_2, n_1, n_0, n_4, n_8, n_6, n_5, n_7, n_112);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_6;
input n_5;
input n_7;

output n_112;

wire n_10;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_9;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

INVx1_ASAP7_75t_L g9 ( 
.A(n_4),
.Y(n_9)
);

INVx1_ASAP7_75t_L g10 ( 
.A(n_4),
.Y(n_10)
);

BUFx12_ASAP7_75t_L g11 ( 
.A(n_4),
.Y(n_11)
);

BUFx12f_ASAP7_75t_L g12 ( 
.A(n_8),
.Y(n_12)
);

BUFx12f_ASAP7_75t_L g13 ( 
.A(n_3),
.Y(n_13)
);

BUFx16f_ASAP7_75t_L g14 ( 
.A(n_8),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_5),
.Y(n_15)
);

INVx4_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_9),
.B(n_0),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_SL g31 ( 
.A(n_20),
.B(n_19),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_14),
.B(n_0),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_21),
.B(n_26),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_22),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_23),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_24),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

AOI22xp33_ASAP7_75t_SL g28 ( 
.A1(n_25),
.A2(n_27),
.B1(n_16),
.B2(n_13),
.Y(n_28)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_28),
.B(n_11),
.Y(n_37)
);

AND2x2_ASAP7_75t_L g30 ( 
.A(n_22),
.B(n_13),
.Y(n_30)
);

AND2x2_ASAP7_75t_L g50 ( 
.A(n_30),
.B(n_33),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_SL g41 ( 
.A(n_31),
.B(n_35),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_23),
.B(n_18),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_SL g35 ( 
.A(n_26),
.B(n_15),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_L g64 ( 
.A1(n_37),
.A2(n_39),
.B1(n_32),
.B2(n_29),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g38 ( 
.A(n_31),
.B(n_19),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_38),
.B(n_46),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g39 ( 
.A1(n_33),
.A2(n_16),
.B1(n_13),
.B2(n_27),
.Y(n_39)
);

MAJx2_ASAP7_75t_L g40 ( 
.A(n_35),
.B(n_13),
.C(n_24),
.Y(n_40)
);

XNOR2xp5_ASAP7_75t_L g59 ( 
.A(n_40),
.B(n_43),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g42 ( 
.A1(n_33),
.A2(n_9),
.B1(n_15),
.B2(n_10),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_L g62 ( 
.A1(n_42),
.A2(n_10),
.B1(n_32),
.B2(n_34),
.Y(n_62)
);

AND2x6_ASAP7_75t_L g43 ( 
.A(n_30),
.B(n_0),
.Y(n_43)
);

INVx11_ASAP7_75t_L g44 ( 
.A(n_29),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_44),
.B(n_45),
.Y(n_54)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_29),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_29),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_47),
.B(n_34),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_36),
.B(n_11),
.Y(n_48)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_48),
.Y(n_55)
);

AOI32xp33_ASAP7_75t_L g49 ( 
.A1(n_30),
.A2(n_36),
.A3(n_34),
.B1(n_32),
.B2(n_28),
.Y(n_49)
);

AOI21xp5_ASAP7_75t_SL g52 ( 
.A1(n_49),
.A2(n_30),
.B(n_29),
.Y(n_52)
);

INVxp67_ASAP7_75t_L g51 ( 
.A(n_39),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_51),
.B(n_62),
.Y(n_68)
);

OAI21xp5_ASAP7_75t_SL g75 ( 
.A1(n_52),
.A2(n_57),
.B(n_43),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g56 ( 
.A(n_41),
.B(n_31),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_SL g76 ( 
.A(n_56),
.B(n_60),
.Y(n_76)
);

AND2x2_ASAP7_75t_L g57 ( 
.A(n_50),
.B(n_30),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_50),
.B(n_18),
.Y(n_58)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_58),
.Y(n_66)
);

NOR2x1_ASAP7_75t_L g60 ( 
.A(n_41),
.B(n_29),
.Y(n_60)
);

CKINVDCx16_ASAP7_75t_R g65 ( 
.A(n_61),
.Y(n_65)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_47),
.Y(n_63)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_63),
.Y(n_71)
);

INVxp67_ASAP7_75t_L g72 ( 
.A(n_64),
.Y(n_72)
);

AOI21xp33_ASAP7_75t_SL g67 ( 
.A1(n_60),
.A2(n_40),
.B(n_50),
.Y(n_67)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_67),
.B(n_69),
.C(n_75),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g69 ( 
.A(n_58),
.B(n_46),
.C(n_49),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_54),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_70),
.B(n_73),
.Y(n_80)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_62),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_53),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_74),
.B(n_25),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_63),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_77),
.Y(n_84)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_68),
.Y(n_78)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_78),
.Y(n_90)
);

AOI322xp5_ASAP7_75t_SL g79 ( 
.A1(n_76),
.A2(n_59),
.A3(n_57),
.B1(n_55),
.B2(n_52),
.C1(n_42),
.C2(n_51),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_79),
.B(n_74),
.C(n_66),
.Y(n_91)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_71),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_81),
.A2(n_72),
.B1(n_73),
.B2(n_65),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_L g82 ( 
.A1(n_69),
.A2(n_57),
.B(n_59),
.Y(n_82)
);

XOR2xp5_ASAP7_75t_L g88 ( 
.A(n_82),
.B(n_86),
.Y(n_88)
);

XOR2xp5_ASAP7_75t_L g87 ( 
.A(n_85),
.B(n_75),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_L g86 ( 
.A1(n_66),
.A2(n_18),
.B(n_17),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_87),
.B(n_88),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_89),
.B(n_80),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_91),
.B(n_85),
.C(n_86),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_83),
.B(n_70),
.C(n_72),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_92),
.B(n_83),
.C(n_82),
.Y(n_95)
);

BUFx2_ASAP7_75t_L g93 ( 
.A(n_84),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_93),
.B(n_44),
.Y(n_94)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_94),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_95),
.B(n_96),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_97),
.A2(n_90),
.B1(n_93),
.B2(n_45),
.Y(n_102)
);

OR2x2_ASAP7_75t_L g101 ( 
.A(n_98),
.B(n_88),
.Y(n_101)
);

A2O1A1O1Ixp25_ASAP7_75t_L g105 ( 
.A1(n_101),
.A2(n_14),
.B(n_17),
.C(n_3),
.D(n_5),
.Y(n_105)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_102),
.Y(n_103)
);

AND2x2_ASAP7_75t_L g104 ( 
.A(n_100),
.B(n_95),
.Y(n_104)
);

AOI322xp5_ASAP7_75t_L g107 ( 
.A1(n_104),
.A2(n_99),
.A3(n_2),
.B1(n_3),
.B2(n_6),
.C1(n_7),
.C2(n_1),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_105),
.B(n_2),
.C(n_6),
.Y(n_109)
);

XNOR2x1_ASAP7_75t_L g106 ( 
.A(n_100),
.B(n_14),
.Y(n_106)
);

AO21x2_ASAP7_75t_L g108 ( 
.A1(n_106),
.A2(n_2),
.B(n_6),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_107),
.B(n_108),
.C(n_109),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_110),
.B(n_103),
.Y(n_111)
);

XOR2xp5_ASAP7_75t_L g112 ( 
.A(n_111),
.B(n_7),
.Y(n_112)
);


endmodule