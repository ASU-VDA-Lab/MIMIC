module fake_ariane_2417_n_1806 (n_83, n_8, n_56, n_60, n_64, n_119, n_124, n_90, n_38, n_47, n_110, n_153, n_18, n_86, n_75, n_89, n_67, n_149, n_34, n_158, n_69, n_95, n_92, n_143, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_152, n_120, n_106, n_12, n_53, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_156, n_49, n_20, n_100, n_17, n_50, n_132, n_62, n_147, n_51, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_11, n_129, n_126, n_137, n_122, n_148, n_52, n_157, n_135, n_73, n_77, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_125, n_22, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_151, n_136, n_28, n_80, n_146, n_97, n_154, n_142, n_14, n_88, n_141, n_68, n_116, n_104, n_145, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_1806);

input n_83;
input n_8;
input n_56;
input n_60;
input n_64;
input n_119;
input n_124;
input n_90;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_149;
input n_34;
input n_158;
input n_69;
input n_95;
input n_92;
input n_143;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_152;
input n_120;
input n_106;
input n_12;
input n_53;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_156;
input n_49;
input n_20;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_147;
input n_51;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_52;
input n_157;
input n_135;
input n_73;
input n_77;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_125;
input n_22;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_151;
input n_136;
input n_28;
input n_80;
input n_146;
input n_97;
input n_154;
input n_142;
input n_14;
input n_88;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_1806;

wire n_913;
wire n_1681;
wire n_1507;
wire n_1486;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_1250;
wire n_1169;
wire n_789;
wire n_850;
wire n_610;
wire n_245;
wire n_1713;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_187;
wire n_1463;
wire n_1238;
wire n_1515;
wire n_817;
wire n_924;
wire n_781;
wire n_1566;
wire n_189;
wire n_717;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_1706;
wire n_524;
wire n_1214;
wire n_634;
wire n_1246;
wire n_1138;
wire n_214;
wire n_764;
wire n_1503;
wire n_462;
wire n_1196;
wire n_1181;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1745;
wire n_1366;
wire n_232;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1457;
wire n_377;
wire n_1682;
wire n_520;
wire n_870;
wire n_1453;
wire n_279;
wire n_945;
wire n_958;
wire n_813;
wire n_419;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1184;
wire n_202;
wire n_1535;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_1277;
wire n_1746;
wire n_829;
wire n_1761;
wire n_1062;
wire n_339;
wire n_738;
wire n_1690;
wire n_672;
wire n_740;
wire n_1283;
wire n_167;
wire n_1736;
wire n_1018;
wire n_259;
wire n_953;
wire n_1364;
wire n_1224;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_1688;
wire n_989;
wire n_645;
wire n_242;
wire n_331;
wire n_559;
wire n_495;
wire n_267;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_200;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_1522;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_1404;
wire n_868;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_1676;
wire n_1085;
wire n_277;
wire n_1636;
wire n_432;
wire n_293;
wire n_823;
wire n_620;
wire n_1074;
wire n_859;
wire n_1765;
wire n_587;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_352;
wire n_206;
wire n_899;
wire n_1703;
wire n_611;
wire n_1295;
wire n_365;
wire n_238;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_334;
wire n_192;
wire n_661;
wire n_1751;
wire n_300;
wire n_533;
wire n_438;
wire n_1560;
wire n_1654;
wire n_1548;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_376;
wire n_512;
wire n_1597;
wire n_1771;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1354;
wire n_1790;
wire n_1213;
wire n_237;
wire n_780;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_209;
wire n_490;
wire n_1461;
wire n_1391;
wire n_225;
wire n_1599;
wire n_1006;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_1594;
wire n_680;
wire n_287;
wire n_1716;
wire n_302;
wire n_380;
wire n_1585;
wire n_1432;
wire n_249;
wire n_1108;
wire n_355;
wire n_212;
wire n_444;
wire n_851;
wire n_1590;
wire n_1351;
wire n_1274;
wire n_257;
wire n_652;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_182;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_407;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_460;
wire n_1555;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_966;
wire n_992;
wire n_955;
wire n_1182;
wire n_794;
wire n_1692;
wire n_1562;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_288;
wire n_179;
wire n_1292;
wire n_1178;
wire n_1435;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_306;
wire n_203;
wire n_436;
wire n_324;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_967;
wire n_1083;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1787;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_1717;
wire n_824;
wire n_428;
wire n_159;
wire n_892;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_990;
wire n_1623;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_1780;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1680;
wire n_964;
wire n_1627;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_1731;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_934;
wire n_1447;
wire n_1220;
wire n_356;
wire n_698;
wire n_1674;
wire n_307;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_1633;
wire n_404;
wire n_172;
wire n_1058;
wire n_347;
wire n_1042;
wire n_183;
wire n_1234;
wire n_479;
wire n_1578;
wire n_1455;
wire n_299;
wire n_836;
wire n_1279;
wire n_564;
wire n_205;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_1689;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_1728;
wire n_370;
wire n_706;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_348;
wire n_552;
wire n_670;
wire n_379;
wire n_162;
wire n_264;
wire n_441;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_1618;
wire n_1743;
wire n_905;
wire n_207;
wire n_720;
wire n_926;
wire n_194;
wire n_1802;
wire n_1163;
wire n_186;
wire n_1795;
wire n_1384;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1648;
wire n_1413;
wire n_855;
wire n_808;
wire n_1365;
wire n_553;
wire n_1439;
wire n_814;
wire n_578;
wire n_1665;
wire n_1287;
wire n_405;
wire n_1611;
wire n_320;
wire n_1414;
wire n_1134;
wire n_1484;
wire n_647;
wire n_1423;
wire n_481;
wire n_600;
wire n_1053;
wire n_1609;
wire n_529;
wire n_502;
wire n_218;
wire n_1467;
wire n_247;
wire n_1798;
wire n_1304;
wire n_1608;
wire n_1744;
wire n_1105;
wire n_547;
wire n_439;
wire n_604;
wire n_677;
wire n_478;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_1278;
wire n_707;
wire n_983;
wire n_727;
wire n_699;
wire n_590;
wire n_301;
wire n_1726;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_325;
wire n_1740;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_729;
wire n_887;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_163;
wire n_1693;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_233;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_321;
wire n_221;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1763;
wire n_1666;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_281;
wire n_262;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_1667;
wire n_845;
wire n_888;
wire n_1649;
wire n_1677;
wire n_1297;
wire n_178;
wire n_551;
wire n_417;
wire n_1708;
wire n_343;
wire n_1222;
wire n_582;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_534;
wire n_1791;
wire n_1460;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_451;
wire n_745;
wire n_1741;
wire n_1572;
wire n_1793;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_769;
wire n_1797;
wire n_1753;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_982;
wire n_1800;
wire n_915;
wire n_215;
wire n_1075;
wire n_454;
wire n_298;
wire n_1331;
wire n_1529;
wire n_1227;
wire n_655;
wire n_1734;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_1700;
wire n_659;
wire n_1332;
wire n_509;
wire n_666;
wire n_1747;
wire n_430;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1766;
wire n_1338;
wire n_1342;
wire n_456;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_521;
wire n_873;
wire n_1301;
wire n_1748;
wire n_1243;
wire n_1400;
wire n_342;
wire n_1466;
wire n_1513;
wire n_1527;
wire n_358;
wire n_1783;
wire n_608;
wire n_1538;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1668;
wire n_1605;
wire n_1078;
wire n_266;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_687;
wire n_797;
wire n_1786;
wire n_480;
wire n_1327;
wire n_1475;
wire n_211;
wire n_642;
wire n_1804;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_1757;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_393;
wire n_1632;
wire n_1769;
wire n_474;
wire n_805;
wire n_295;
wire n_1658;
wire n_190;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_180;
wire n_730;
wire n_386;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1137;
wire n_1258;
wire n_197;
wire n_640;
wire n_463;
wire n_1476;
wire n_1524;
wire n_1733;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_1784;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_283;
wire n_806;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_643;
wire n_1492;
wire n_226;
wire n_1441;
wire n_682;
wire n_1616;
wire n_819;
wire n_586;
wire n_1324;
wire n_1429;
wire n_1778;
wire n_1776;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1759;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_198;
wire n_1208;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1577;
wire n_1448;
wire n_1009;
wire n_230;
wire n_1133;
wire n_883;
wire n_473;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_594;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_169;
wire n_1201;
wire n_1288;
wire n_173;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_426;
wire n_433;
wire n_398;
wire n_210;
wire n_1090;
wire n_1367;
wire n_253;
wire n_166;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_224;
wire n_894;
wire n_1380;
wire n_1624;
wire n_1801;
wire n_420;
wire n_1291;
wire n_562;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1023;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_467;
wire n_1511;
wire n_1422;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_1641;
wire n_168;
wire n_538;
wire n_1517;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_1307;
wire n_1128;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1773;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_810;
wire n_1290;
wire n_181;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_628;
wire n_1300;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_414;
wire n_571;
wire n_1521;
wire n_1694;
wire n_284;
wire n_593;
wire n_1695;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_1774;
wire n_409;
wire n_171;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_526;
wire n_1767;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1444;
wire n_1803;
wire n_820;
wire n_1749;
wire n_872;
wire n_1653;
wire n_254;
wire n_1157;
wire n_1584;
wire n_234;
wire n_848;
wire n_1664;
wire n_280;
wire n_629;
wire n_1739;
wire n_161;
wire n_532;
wire n_1789;
wire n_763;
wire n_540;
wire n_216;
wire n_692;
wire n_984;
wire n_1687;
wire n_223;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_1756;
wire n_1606;
wire n_395;
wire n_621;
wire n_1587;
wire n_213;
wire n_1772;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_493;
wire n_1311;
wire n_1589;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_697;
wire n_622;
wire n_1626;
wire n_1335;
wire n_1715;
wire n_296;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_1785;
wire n_792;
wire n_1262;
wire n_580;
wire n_1579;
wire n_494;
wire n_434;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1183;
wire n_1326;
wire n_1805;
wire n_981;
wire n_1110;
wire n_1758;
wire n_243;
wire n_1407;
wire n_185;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_164;
wire n_184;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_1054;
wire n_508;
wire n_1679;
wire n_353;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_191;
wire n_1011;
wire n_978;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_1721;
wire n_653;
wire n_1445;
wire n_1317;
wire n_783;
wire n_556;
wire n_1127;
wire n_170;
wire n_1536;
wire n_1471;
wire n_160;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_176;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_541;
wire n_499;
wire n_1775;
wire n_788;
wire n_908;
wire n_1036;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_1663;
wire n_1625;
wire n_318;
wire n_1458;
wire n_244;
wire n_679;
wire n_1630;
wire n_220;
wire n_663;
wire n_1720;
wire n_443;
wire n_1412;
wire n_1738;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_1735;
wire n_1788;
wire n_391;
wire n_940;
wire n_1537;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_765;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_1530;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_857;
wire n_898;
wire n_363;
wire n_1067;
wire n_968;
wire n_1235;
wire n_1323;
wire n_1462;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_1755;
wire n_1285;
wire n_193;
wire n_733;
wire n_761;
wire n_731;
wire n_336;
wire n_315;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_1106;
wire n_648;
wire n_784;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_1348;
wire n_753;
wire n_1770;
wire n_701;
wire n_1003;
wire n_1125;
wire n_1710;
wire n_309;
wire n_1344;
wire n_1390;
wire n_401;
wire n_485;
wire n_1792;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_291;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1510;
wire n_1099;
wire n_839;
wire n_1754;
wire n_759;
wire n_567;
wire n_369;
wire n_240;
wire n_1727;
wire n_1575;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_188;
wire n_323;
wire n_550;
wire n_1315;
wire n_1660;
wire n_997;
wire n_635;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_248;
wire n_1152;
wire n_921;
wire n_1615;
wire n_1236;
wire n_228;
wire n_1265;
wire n_1576;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1684;
wire n_1673;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_1696;
wire n_498;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1497;
wire n_459;
wire n_1136;
wire n_1782;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_383;
wire n_838;
wire n_1558;
wire n_1316;
wire n_175;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_1781;
wire n_709;
wire n_809;
wire n_1686;
wire n_235;
wire n_881;
wire n_1019;
wire n_1477;
wire n_1777;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_199;
wire n_217;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_708;
wire n_308;
wire n_1223;
wire n_201;
wire n_1768;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1041;
wire n_993;
wire n_948;
wire n_922;
wire n_1004;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_1764;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_196;
wire n_1337;
wire n_774;
wire n_933;
wire n_1779;
wire n_596;
wire n_954;
wire n_1168;
wire n_219;
wire n_1310;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_252;
wire n_664;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_1732;
wire n_415;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1724;
wire n_1670;
wire n_1707;
wire n_1799;
wire n_1126;
wire n_195;
wire n_938;
wire n_1328;
wire n_895;
wire n_304;
wire n_1639;
wire n_583;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_946;
wire n_757;
wire n_375;
wire n_1655;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_472;
wire n_937;
wire n_1474;
wire n_265;
wire n_1583;
wire n_1604;
wire n_208;
wire n_1631;
wire n_1702;
wire n_174;
wire n_275;
wire n_1794;
wire n_1375;
wire n_204;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_496;
wire n_866;
wire n_246;
wire n_925;
wire n_1752;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_1129;
wire n_1252;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_165;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_329;
wire n_718;
wire n_1434;
wire n_340;
wire n_1569;
wire n_548;
wire n_289;
wire n_523;
wire n_1662;
wire n_457;
wire n_1299;
wire n_177;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1228;
wire n_1244;
wire n_1796;
wire n_411;
wire n_484;
wire n_849;
wire n_357;
wire n_412;
wire n_1251;
wire n_447;
wire n_1421;
wire n_1762;
wire n_1233;
wire n_1574;
wire n_1672;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_1487;
wire n_675;

INVx1_ASAP7_75t_L g159 ( 
.A(n_31),
.Y(n_159)
);

CKINVDCx5p33_ASAP7_75t_R g160 ( 
.A(n_58),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_54),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_148),
.Y(n_162)
);

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_144),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_43),
.Y(n_164)
);

CKINVDCx5p33_ASAP7_75t_R g165 ( 
.A(n_44),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_137),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_81),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_95),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_8),
.Y(n_169)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_131),
.Y(n_170)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_149),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_105),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_46),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_27),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_122),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_59),
.Y(n_176)
);

BUFx2_ASAP7_75t_L g177 ( 
.A(n_66),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_113),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_109),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_25),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_130),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_39),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_15),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_21),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_129),
.Y(n_185)
);

INVxp67_ASAP7_75t_L g186 ( 
.A(n_53),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_90),
.Y(n_187)
);

INVx1_ASAP7_75t_SL g188 ( 
.A(n_154),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_44),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_133),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_17),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_7),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_135),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_151),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_33),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_30),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_146),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_20),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_134),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_32),
.Y(n_200)
);

BUFx3_ASAP7_75t_L g201 ( 
.A(n_126),
.Y(n_201)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_41),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_124),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_52),
.Y(n_204)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_40),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_114),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_156),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_50),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_6),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_140),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_121),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_76),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_89),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_43),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_73),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_12),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_6),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_24),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_158),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_125),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_30),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_23),
.Y(n_222)
);

BUFx8_ASAP7_75t_SL g223 ( 
.A(n_99),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_48),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_10),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_82),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_26),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_51),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_55),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_93),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_108),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_112),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_110),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_7),
.Y(n_234)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_145),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_37),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_92),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_107),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_69),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_100),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_116),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_94),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_36),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_96),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_77),
.Y(n_245)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_50),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_102),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_152),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_71),
.Y(n_249)
);

BUFx3_ASAP7_75t_L g250 ( 
.A(n_74),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_8),
.Y(n_251)
);

CKINVDCx16_ASAP7_75t_R g252 ( 
.A(n_67),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_101),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_91),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_142),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_36),
.Y(n_256)
);

INVx2_ASAP7_75t_SL g257 ( 
.A(n_20),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_10),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_48),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_56),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_40),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_13),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_49),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_12),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_3),
.Y(n_265)
);

BUFx6f_ASAP7_75t_L g266 ( 
.A(n_34),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_45),
.Y(n_267)
);

BUFx2_ASAP7_75t_L g268 ( 
.A(n_31),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_34),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_85),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_0),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_72),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_87),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_78),
.Y(n_274)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_79),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_0),
.Y(n_276)
);

INVx1_ASAP7_75t_SL g277 ( 
.A(n_16),
.Y(n_277)
);

HB1xp67_ASAP7_75t_L g278 ( 
.A(n_86),
.Y(n_278)
);

BUFx2_ASAP7_75t_SL g279 ( 
.A(n_26),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_153),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_119),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_115),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_4),
.Y(n_283)
);

BUFx3_ASAP7_75t_L g284 ( 
.A(n_60),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_68),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_23),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_117),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_35),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_47),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_11),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_46),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_138),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_118),
.Y(n_293)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_2),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_29),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_141),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_139),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_147),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_47),
.Y(n_299)
);

INVx2_ASAP7_75t_L g300 ( 
.A(n_14),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_157),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_37),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_1),
.Y(n_303)
);

INVx2_ASAP7_75t_SL g304 ( 
.A(n_83),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_27),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_22),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_25),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_155),
.Y(n_308)
);

INVx2_ASAP7_75t_L g309 ( 
.A(n_62),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_61),
.Y(n_310)
);

BUFx3_ASAP7_75t_L g311 ( 
.A(n_128),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_19),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_132),
.Y(n_313)
);

INVxp33_ASAP7_75t_SL g314 ( 
.A(n_268),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_223),
.Y(n_315)
);

BUFx6f_ASAP7_75t_L g316 ( 
.A(n_266),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_161),
.Y(n_317)
);

INVx2_ASAP7_75t_L g318 ( 
.A(n_266),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_161),
.Y(n_319)
);

INVxp67_ASAP7_75t_L g320 ( 
.A(n_268),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_194),
.Y(n_321)
);

HB1xp67_ASAP7_75t_L g322 ( 
.A(n_165),
.Y(n_322)
);

INVxp67_ASAP7_75t_L g323 ( 
.A(n_279),
.Y(n_323)
);

BUFx2_ASAP7_75t_L g324 ( 
.A(n_205),
.Y(n_324)
);

INVxp67_ASAP7_75t_SL g325 ( 
.A(n_205),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_167),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_194),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_204),
.Y(n_328)
);

INVxp67_ASAP7_75t_L g329 ( 
.A(n_279),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_204),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_213),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_213),
.Y(n_332)
);

INVxp33_ASAP7_75t_SL g333 ( 
.A(n_169),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_215),
.Y(n_334)
);

CKINVDCx16_ASAP7_75t_R g335 ( 
.A(n_252),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g336 ( 
.A(n_179),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_181),
.Y(n_337)
);

INVxp33_ASAP7_75t_SL g338 ( 
.A(n_182),
.Y(n_338)
);

CKINVDCx20_ASAP7_75t_R g339 ( 
.A(n_187),
.Y(n_339)
);

INVxp67_ASAP7_75t_L g340 ( 
.A(n_159),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_215),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_219),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_210),
.Y(n_343)
);

CKINVDCx20_ASAP7_75t_R g344 ( 
.A(n_253),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_219),
.Y(n_345)
);

INVx2_ASAP7_75t_L g346 ( 
.A(n_266),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_229),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_229),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_230),
.Y(n_349)
);

HB1xp67_ASAP7_75t_L g350 ( 
.A(n_183),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_282),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_230),
.Y(n_352)
);

INVx2_ASAP7_75t_L g353 ( 
.A(n_266),
.Y(n_353)
);

CKINVDCx20_ASAP7_75t_R g354 ( 
.A(n_313),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_237),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_237),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_239),
.Y(n_357)
);

INVx2_ASAP7_75t_L g358 ( 
.A(n_266),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_239),
.Y(n_359)
);

INVx2_ASAP7_75t_L g360 ( 
.A(n_266),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_244),
.Y(n_361)
);

CKINVDCx20_ASAP7_75t_R g362 ( 
.A(n_198),
.Y(n_362)
);

INVxp67_ASAP7_75t_L g363 ( 
.A(n_159),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_244),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_248),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_248),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_270),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_270),
.Y(n_368)
);

CKINVDCx20_ASAP7_75t_R g369 ( 
.A(n_217),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_293),
.Y(n_370)
);

INVxp67_ASAP7_75t_SL g371 ( 
.A(n_246),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_293),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_184),
.Y(n_373)
);

CKINVDCx20_ASAP7_75t_R g374 ( 
.A(n_262),
.Y(n_374)
);

INVxp33_ASAP7_75t_SL g375 ( 
.A(n_191),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_296),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_296),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_298),
.Y(n_378)
);

INVxp67_ASAP7_75t_SL g379 ( 
.A(n_246),
.Y(n_379)
);

CKINVDCx20_ASAP7_75t_R g380 ( 
.A(n_312),
.Y(n_380)
);

INVxp33_ASAP7_75t_SL g381 ( 
.A(n_192),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_298),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_301),
.Y(n_383)
);

INVx2_ASAP7_75t_L g384 ( 
.A(n_201),
.Y(n_384)
);

INVxp67_ASAP7_75t_L g385 ( 
.A(n_164),
.Y(n_385)
);

INVxp33_ASAP7_75t_SL g386 ( 
.A(n_195),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_301),
.Y(n_387)
);

CKINVDCx16_ASAP7_75t_R g388 ( 
.A(n_252),
.Y(n_388)
);

XNOR2x2_ASAP7_75t_L g389 ( 
.A(n_314),
.B(n_277),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_317),
.Y(n_390)
);

BUFx6f_ASAP7_75t_L g391 ( 
.A(n_316),
.Y(n_391)
);

INVx3_ASAP7_75t_L g392 ( 
.A(n_316),
.Y(n_392)
);

INVx2_ASAP7_75t_L g393 ( 
.A(n_316),
.Y(n_393)
);

INVx3_ASAP7_75t_L g394 ( 
.A(n_316),
.Y(n_394)
);

AND2x2_ASAP7_75t_L g395 ( 
.A(n_324),
.B(n_177),
.Y(n_395)
);

BUFx6f_ASAP7_75t_L g396 ( 
.A(n_316),
.Y(n_396)
);

BUFx6f_ASAP7_75t_L g397 ( 
.A(n_318),
.Y(n_397)
);

INVx3_ASAP7_75t_L g398 ( 
.A(n_318),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_317),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_384),
.B(n_177),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_326),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_319),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_319),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_321),
.Y(n_404)
);

INVx3_ASAP7_75t_L g405 ( 
.A(n_346),
.Y(n_405)
);

INVx2_ASAP7_75t_L g406 ( 
.A(n_346),
.Y(n_406)
);

OAI22xp5_ASAP7_75t_L g407 ( 
.A1(n_320),
.A2(n_257),
.B1(n_174),
.B2(n_180),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_384),
.B(n_278),
.Y(n_408)
);

AND2x4_ASAP7_75t_L g409 ( 
.A(n_321),
.B(n_327),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_327),
.Y(n_410)
);

INVx2_ASAP7_75t_L g411 ( 
.A(n_353),
.Y(n_411)
);

NAND2x1p5_ASAP7_75t_L g412 ( 
.A(n_328),
.B(n_201),
.Y(n_412)
);

HB1xp67_ASAP7_75t_L g413 ( 
.A(n_373),
.Y(n_413)
);

BUFx6f_ASAP7_75t_L g414 ( 
.A(n_353),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_328),
.Y(n_415)
);

BUFx6f_ASAP7_75t_L g416 ( 
.A(n_358),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_330),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_330),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_331),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_331),
.Y(n_420)
);

AND2x6_ASAP7_75t_L g421 ( 
.A(n_332),
.B(n_275),
.Y(n_421)
);

INVx3_ASAP7_75t_L g422 ( 
.A(n_358),
.Y(n_422)
);

NOR2x1_ASAP7_75t_L g423 ( 
.A(n_332),
.B(n_201),
.Y(n_423)
);

INVxp67_ASAP7_75t_L g424 ( 
.A(n_322),
.Y(n_424)
);

BUFx6f_ASAP7_75t_L g425 ( 
.A(n_360),
.Y(n_425)
);

INVx2_ASAP7_75t_L g426 ( 
.A(n_360),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_334),
.Y(n_427)
);

HB1xp67_ASAP7_75t_L g428 ( 
.A(n_350),
.Y(n_428)
);

NAND2xp33_ASAP7_75t_R g429 ( 
.A(n_333),
.B(n_196),
.Y(n_429)
);

INVx2_ASAP7_75t_L g430 ( 
.A(n_334),
.Y(n_430)
);

BUFx6f_ASAP7_75t_L g431 ( 
.A(n_341),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_341),
.Y(n_432)
);

OAI21x1_ASAP7_75t_L g433 ( 
.A1(n_342),
.A2(n_309),
.B(n_275),
.Y(n_433)
);

AND2x4_ASAP7_75t_L g434 ( 
.A(n_342),
.B(n_246),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_337),
.Y(n_435)
);

INVx2_ASAP7_75t_L g436 ( 
.A(n_345),
.Y(n_436)
);

CKINVDCx5p33_ASAP7_75t_R g437 ( 
.A(n_343),
.Y(n_437)
);

INVx3_ASAP7_75t_L g438 ( 
.A(n_345),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_347),
.Y(n_439)
);

OAI21x1_ASAP7_75t_L g440 ( 
.A1(n_347),
.A2(n_309),
.B(n_275),
.Y(n_440)
);

OAI22xp5_ASAP7_75t_L g441 ( 
.A1(n_388),
.A2(n_257),
.B1(n_174),
.B2(n_164),
.Y(n_441)
);

NOR2xp33_ASAP7_75t_L g442 ( 
.A(n_338),
.B(n_375),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_348),
.B(n_304),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_348),
.Y(n_444)
);

INVx2_ASAP7_75t_L g445 ( 
.A(n_349),
.Y(n_445)
);

CKINVDCx20_ASAP7_75t_R g446 ( 
.A(n_362),
.Y(n_446)
);

NOR2xp67_ASAP7_75t_L g447 ( 
.A(n_349),
.B(n_304),
.Y(n_447)
);

INVx3_ASAP7_75t_L g448 ( 
.A(n_352),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_352),
.Y(n_449)
);

NOR2xp33_ASAP7_75t_L g450 ( 
.A(n_381),
.B(n_186),
.Y(n_450)
);

BUFx6f_ASAP7_75t_L g451 ( 
.A(n_355),
.Y(n_451)
);

BUFx6f_ASAP7_75t_L g452 ( 
.A(n_355),
.Y(n_452)
);

BUFx6f_ASAP7_75t_L g453 ( 
.A(n_356),
.Y(n_453)
);

INVx4_ASAP7_75t_L g454 ( 
.A(n_356),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_357),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_357),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_L g457 ( 
.A(n_359),
.B(n_188),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_359),
.Y(n_458)
);

AND2x2_ASAP7_75t_L g459 ( 
.A(n_324),
.B(n_294),
.Y(n_459)
);

BUFx3_ASAP7_75t_L g460 ( 
.A(n_409),
.Y(n_460)
);

AOI22xp33_ASAP7_75t_L g461 ( 
.A1(n_441),
.A2(n_376),
.B1(n_387),
.B2(n_364),
.Y(n_461)
);

CKINVDCx20_ASAP7_75t_R g462 ( 
.A(n_446),
.Y(n_462)
);

AND2x2_ASAP7_75t_L g463 ( 
.A(n_409),
.B(n_325),
.Y(n_463)
);

INVx2_ASAP7_75t_L g464 ( 
.A(n_406),
.Y(n_464)
);

NOR2xp33_ASAP7_75t_L g465 ( 
.A(n_450),
.B(n_335),
.Y(n_465)
);

INVxp67_ASAP7_75t_L g466 ( 
.A(n_429),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_L g467 ( 
.A(n_409),
.B(n_388),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_431),
.Y(n_468)
);

AOI22xp33_ASAP7_75t_L g469 ( 
.A1(n_441),
.A2(n_387),
.B1(n_361),
.B2(n_364),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_431),
.Y(n_470)
);

INVx6_ASAP7_75t_L g471 ( 
.A(n_454),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_431),
.Y(n_472)
);

INVx2_ASAP7_75t_L g473 ( 
.A(n_406),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_431),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_431),
.Y(n_475)
);

BUFx6f_ASAP7_75t_L g476 ( 
.A(n_431),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_431),
.Y(n_477)
);

OAI22xp33_ASAP7_75t_SL g478 ( 
.A1(n_407),
.A2(n_385),
.B1(n_340),
.B2(n_363),
.Y(n_478)
);

HB1xp67_ASAP7_75t_L g479 ( 
.A(n_401),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_451),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_SL g481 ( 
.A(n_442),
.B(n_386),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_451),
.Y(n_482)
);

INVx2_ASAP7_75t_L g483 ( 
.A(n_411),
.Y(n_483)
);

BUFx2_ASAP7_75t_L g484 ( 
.A(n_435),
.Y(n_484)
);

NOR2xp33_ASAP7_75t_L g485 ( 
.A(n_454),
.B(n_323),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_451),
.Y(n_486)
);

OR2x6_ASAP7_75t_L g487 ( 
.A(n_412),
.B(n_361),
.Y(n_487)
);

HB1xp67_ASAP7_75t_L g488 ( 
.A(n_437),
.Y(n_488)
);

INVx3_ASAP7_75t_L g489 ( 
.A(n_451),
.Y(n_489)
);

NOR2xp33_ASAP7_75t_L g490 ( 
.A(n_454),
.B(n_329),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_451),
.Y(n_491)
);

INVx2_ASAP7_75t_L g492 ( 
.A(n_411),
.Y(n_492)
);

AOI22xp5_ASAP7_75t_L g493 ( 
.A1(n_424),
.A2(n_227),
.B1(n_200),
.B2(n_208),
.Y(n_493)
);

AND2x2_ASAP7_75t_L g494 ( 
.A(n_434),
.B(n_371),
.Y(n_494)
);

INVx2_ASAP7_75t_SL g495 ( 
.A(n_412),
.Y(n_495)
);

INVx2_ASAP7_75t_SL g496 ( 
.A(n_412),
.Y(n_496)
);

INVx2_ASAP7_75t_L g497 ( 
.A(n_411),
.Y(n_497)
);

CKINVDCx5p33_ASAP7_75t_R g498 ( 
.A(n_413),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_L g499 ( 
.A(n_457),
.B(n_379),
.Y(n_499)
);

AO21x2_ASAP7_75t_L g500 ( 
.A1(n_433),
.A2(n_366),
.B(n_365),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_451),
.Y(n_501)
);

BUFx4f_ASAP7_75t_L g502 ( 
.A(n_451),
.Y(n_502)
);

INVx4_ASAP7_75t_L g503 ( 
.A(n_438),
.Y(n_503)
);

INVx2_ASAP7_75t_L g504 ( 
.A(n_426),
.Y(n_504)
);

INVx2_ASAP7_75t_L g505 ( 
.A(n_426),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_452),
.Y(n_506)
);

OR2x6_ASAP7_75t_L g507 ( 
.A(n_412),
.B(n_365),
.Y(n_507)
);

INVx2_ASAP7_75t_SL g508 ( 
.A(n_428),
.Y(n_508)
);

INVx2_ASAP7_75t_L g509 ( 
.A(n_426),
.Y(n_509)
);

INVx2_ASAP7_75t_L g510 ( 
.A(n_452),
.Y(n_510)
);

INVx2_ASAP7_75t_L g511 ( 
.A(n_452),
.Y(n_511)
);

INVx2_ASAP7_75t_L g512 ( 
.A(n_452),
.Y(n_512)
);

BUFx6f_ASAP7_75t_L g513 ( 
.A(n_452),
.Y(n_513)
);

INVx2_ASAP7_75t_SL g514 ( 
.A(n_395),
.Y(n_514)
);

AO22x2_ASAP7_75t_L g515 ( 
.A1(n_407),
.A2(n_383),
.B1(n_382),
.B2(n_368),
.Y(n_515)
);

INVx2_ASAP7_75t_L g516 ( 
.A(n_452),
.Y(n_516)
);

INVx3_ASAP7_75t_L g517 ( 
.A(n_452),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_453),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_SL g519 ( 
.A(n_424),
.B(n_315),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_453),
.Y(n_520)
);

NAND2xp33_ASAP7_75t_R g521 ( 
.A(n_395),
.B(n_351),
.Y(n_521)
);

AO21x2_ASAP7_75t_L g522 ( 
.A1(n_433),
.A2(n_368),
.B(n_367),
.Y(n_522)
);

INVx3_ASAP7_75t_L g523 ( 
.A(n_453),
.Y(n_523)
);

BUFx10_ASAP7_75t_L g524 ( 
.A(n_434),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_453),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_453),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_L g527 ( 
.A(n_454),
.B(n_367),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_453),
.Y(n_528)
);

INVx2_ASAP7_75t_SL g529 ( 
.A(n_459),
.Y(n_529)
);

INVx3_ASAP7_75t_L g530 ( 
.A(n_453),
.Y(n_530)
);

INVx4_ASAP7_75t_L g531 ( 
.A(n_438),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_438),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_438),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_448),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_SL g535 ( 
.A(n_448),
.B(n_370),
.Y(n_535)
);

NAND2xp33_ASAP7_75t_R g536 ( 
.A(n_459),
.B(n_336),
.Y(n_536)
);

INVx2_ASAP7_75t_L g537 ( 
.A(n_398),
.Y(n_537)
);

INVx4_ASAP7_75t_L g538 ( 
.A(n_448),
.Y(n_538)
);

INVx2_ASAP7_75t_L g539 ( 
.A(n_398),
.Y(n_539)
);

INVx2_ASAP7_75t_L g540 ( 
.A(n_398),
.Y(n_540)
);

NOR3xp33_ASAP7_75t_L g541 ( 
.A(n_448),
.B(n_180),
.C(n_173),
.Y(n_541)
);

INVx2_ASAP7_75t_L g542 ( 
.A(n_398),
.Y(n_542)
);

BUFx2_ASAP7_75t_L g543 ( 
.A(n_389),
.Y(n_543)
);

BUFx3_ASAP7_75t_L g544 ( 
.A(n_390),
.Y(n_544)
);

INVx2_ASAP7_75t_L g545 ( 
.A(n_405),
.Y(n_545)
);

AO22x2_ASAP7_75t_L g546 ( 
.A1(n_389),
.A2(n_383),
.B1(n_382),
.B2(n_378),
.Y(n_546)
);

INVx3_ASAP7_75t_L g547 ( 
.A(n_430),
.Y(n_547)
);

INVx1_ASAP7_75t_SL g548 ( 
.A(n_400),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_433),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_L g550 ( 
.A(n_390),
.B(n_370),
.Y(n_550)
);

INVx2_ASAP7_75t_SL g551 ( 
.A(n_400),
.Y(n_551)
);

INVx4_ASAP7_75t_L g552 ( 
.A(n_434),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_SL g553 ( 
.A(n_443),
.B(n_372),
.Y(n_553)
);

BUFx2_ASAP7_75t_L g554 ( 
.A(n_389),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_440),
.Y(n_555)
);

INVx2_ASAP7_75t_SL g556 ( 
.A(n_408),
.Y(n_556)
);

INVx2_ASAP7_75t_L g557 ( 
.A(n_405),
.Y(n_557)
);

INVx3_ASAP7_75t_L g558 ( 
.A(n_430),
.Y(n_558)
);

NOR2xp33_ASAP7_75t_L g559 ( 
.A(n_408),
.B(n_372),
.Y(n_559)
);

INVx2_ASAP7_75t_SL g560 ( 
.A(n_423),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_SL g561 ( 
.A(n_443),
.B(n_376),
.Y(n_561)
);

BUFx3_ASAP7_75t_L g562 ( 
.A(n_399),
.Y(n_562)
);

INVxp33_ASAP7_75t_SL g563 ( 
.A(n_423),
.Y(n_563)
);

AOI22xp5_ASAP7_75t_L g564 ( 
.A1(n_434),
.A2(n_251),
.B1(n_259),
.B2(n_261),
.Y(n_564)
);

CKINVDCx5p33_ASAP7_75t_R g565 ( 
.A(n_421),
.Y(n_565)
);

BUFx10_ASAP7_75t_L g566 ( 
.A(n_399),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_440),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_SL g568 ( 
.A(n_402),
.B(n_403),
.Y(n_568)
);

BUFx3_ASAP7_75t_L g569 ( 
.A(n_402),
.Y(n_569)
);

INVx2_ASAP7_75t_L g570 ( 
.A(n_405),
.Y(n_570)
);

AND2x2_ASAP7_75t_L g571 ( 
.A(n_403),
.B(n_377),
.Y(n_571)
);

INVx2_ASAP7_75t_L g572 ( 
.A(n_405),
.Y(n_572)
);

INVx2_ASAP7_75t_L g573 ( 
.A(n_422),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_440),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_430),
.Y(n_575)
);

BUFx6f_ASAP7_75t_L g576 ( 
.A(n_397),
.Y(n_576)
);

INVx2_ASAP7_75t_L g577 ( 
.A(n_422),
.Y(n_577)
);

INVx2_ASAP7_75t_L g578 ( 
.A(n_422),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_SL g579 ( 
.A(n_404),
.B(n_410),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_436),
.Y(n_580)
);

INVx4_ASAP7_75t_L g581 ( 
.A(n_421),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_436),
.Y(n_582)
);

NOR2xp33_ASAP7_75t_L g583 ( 
.A(n_404),
.B(n_377),
.Y(n_583)
);

INVx2_ASAP7_75t_L g584 ( 
.A(n_422),
.Y(n_584)
);

INVx2_ASAP7_75t_L g585 ( 
.A(n_397),
.Y(n_585)
);

INVx2_ASAP7_75t_SL g586 ( 
.A(n_410),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_L g587 ( 
.A(n_415),
.B(n_417),
.Y(n_587)
);

CKINVDCx5p33_ASAP7_75t_R g588 ( 
.A(n_421),
.Y(n_588)
);

INVx8_ASAP7_75t_L g589 ( 
.A(n_421),
.Y(n_589)
);

INVx2_ASAP7_75t_L g590 ( 
.A(n_397),
.Y(n_590)
);

INVx2_ASAP7_75t_L g591 ( 
.A(n_397),
.Y(n_591)
);

NOR2xp33_ASAP7_75t_L g592 ( 
.A(n_415),
.B(n_378),
.Y(n_592)
);

OAI22xp33_ASAP7_75t_SL g593 ( 
.A1(n_417),
.A2(n_256),
.B1(n_258),
.B2(n_236),
.Y(n_593)
);

INVxp67_ASAP7_75t_L g594 ( 
.A(n_447),
.Y(n_594)
);

INVx2_ASAP7_75t_L g595 ( 
.A(n_397),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_436),
.Y(n_596)
);

OR2x6_ASAP7_75t_L g597 ( 
.A(n_447),
.B(n_202),
.Y(n_597)
);

BUFx6f_ASAP7_75t_L g598 ( 
.A(n_397),
.Y(n_598)
);

INVx2_ASAP7_75t_L g599 ( 
.A(n_414),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_445),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_SL g601 ( 
.A(n_418),
.B(n_209),
.Y(n_601)
);

AOI22xp5_ASAP7_75t_L g602 ( 
.A1(n_421),
.A2(n_243),
.B1(n_263),
.B2(n_269),
.Y(n_602)
);

INVxp67_ASAP7_75t_L g603 ( 
.A(n_418),
.Y(n_603)
);

NAND2xp33_ASAP7_75t_L g604 ( 
.A(n_419),
.B(n_309),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_445),
.Y(n_605)
);

AND2x4_ASAP7_75t_L g606 ( 
.A(n_419),
.B(n_173),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_SL g607 ( 
.A(n_566),
.B(n_420),
.Y(n_607)
);

INVx4_ASAP7_75t_L g608 ( 
.A(n_589),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_L g609 ( 
.A(n_556),
.B(n_420),
.Y(n_609)
);

INVx2_ASAP7_75t_L g610 ( 
.A(n_464),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_L g611 ( 
.A(n_556),
.B(n_427),
.Y(n_611)
);

NOR2xp33_ASAP7_75t_L g612 ( 
.A(n_563),
.B(n_427),
.Y(n_612)
);

AND2x4_ASAP7_75t_L g613 ( 
.A(n_460),
.B(n_432),
.Y(n_613)
);

A2O1A1Ixp33_ASAP7_75t_L g614 ( 
.A1(n_559),
.A2(n_458),
.B(n_456),
.C(n_455),
.Y(n_614)
);

BUFx6f_ASAP7_75t_L g615 ( 
.A(n_460),
.Y(n_615)
);

INVx2_ASAP7_75t_SL g616 ( 
.A(n_508),
.Y(n_616)
);

INVx2_ASAP7_75t_SL g617 ( 
.A(n_508),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_SL g618 ( 
.A(n_566),
.B(n_432),
.Y(n_618)
);

BUFx6f_ASAP7_75t_SL g619 ( 
.A(n_514),
.Y(n_619)
);

AOI22xp33_ASAP7_75t_L g620 ( 
.A1(n_546),
.A2(n_421),
.B1(n_445),
.B2(n_455),
.Y(n_620)
);

NOR2xp33_ASAP7_75t_L g621 ( 
.A(n_563),
.B(n_439),
.Y(n_621)
);

NOR2xp33_ASAP7_75t_L g622 ( 
.A(n_548),
.B(n_439),
.Y(n_622)
);

NOR2xp33_ASAP7_75t_L g623 ( 
.A(n_551),
.B(n_444),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_SL g624 ( 
.A(n_566),
.B(n_444),
.Y(n_624)
);

OR2x2_ASAP7_75t_L g625 ( 
.A(n_484),
.B(n_339),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_544),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_SL g627 ( 
.A(n_503),
.B(n_449),
.Y(n_627)
);

INVx2_ASAP7_75t_SL g628 ( 
.A(n_514),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_SL g629 ( 
.A(n_503),
.B(n_449),
.Y(n_629)
);

O2A1O1Ixp33_ASAP7_75t_L g630 ( 
.A1(n_553),
.A2(n_458),
.B(n_456),
.C(n_294),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_SL g631 ( 
.A(n_503),
.B(n_170),
.Y(n_631)
);

INVx2_ASAP7_75t_SL g632 ( 
.A(n_498),
.Y(n_632)
);

NOR2xp33_ASAP7_75t_L g633 ( 
.A(n_551),
.B(n_216),
.Y(n_633)
);

NOR2xp33_ASAP7_75t_L g634 ( 
.A(n_467),
.B(n_218),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_544),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_562),
.Y(n_636)
);

OAI22xp5_ASAP7_75t_SL g637 ( 
.A1(n_462),
.A2(n_380),
.B1(n_374),
.B2(n_369),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_SL g638 ( 
.A(n_531),
.B(n_170),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_SL g639 ( 
.A(n_531),
.B(n_171),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_562),
.Y(n_640)
);

NAND3xp33_ASAP7_75t_L g641 ( 
.A(n_465),
.B(n_225),
.C(n_221),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_SL g642 ( 
.A(n_531),
.B(n_171),
.Y(n_642)
);

O2A1O1Ixp5_ASAP7_75t_L g643 ( 
.A1(n_568),
.A2(n_394),
.B(n_392),
.C(n_294),
.Y(n_643)
);

NOR3xp33_ASAP7_75t_L g644 ( 
.A(n_481),
.B(n_214),
.C(n_189),
.Y(n_644)
);

AOI22xp33_ASAP7_75t_L g645 ( 
.A1(n_546),
.A2(n_421),
.B1(n_300),
.B2(n_202),
.Y(n_645)
);

INVx3_ASAP7_75t_L g646 ( 
.A(n_538),
.Y(n_646)
);

NOR2xp33_ASAP7_75t_L g647 ( 
.A(n_466),
.B(n_228),
.Y(n_647)
);

NOR2xp33_ASAP7_75t_L g648 ( 
.A(n_552),
.B(n_276),
.Y(n_648)
);

AND2x2_ASAP7_75t_L g649 ( 
.A(n_484),
.B(n_344),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_569),
.Y(n_650)
);

AOI22xp5_ASAP7_75t_L g651 ( 
.A1(n_586),
.A2(n_507),
.B1(n_487),
.B2(n_463),
.Y(n_651)
);

BUFx3_ASAP7_75t_L g652 ( 
.A(n_479),
.Y(n_652)
);

NOR2xp33_ASAP7_75t_L g653 ( 
.A(n_552),
.B(n_283),
.Y(n_653)
);

NAND3xp33_ASAP7_75t_L g654 ( 
.A(n_485),
.B(n_289),
.C(n_288),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_L g655 ( 
.A(n_499),
.B(n_421),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_569),
.Y(n_656)
);

NOR2xp67_ASAP7_75t_L g657 ( 
.A(n_488),
.B(n_392),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_532),
.Y(n_658)
);

INVx2_ASAP7_75t_L g659 ( 
.A(n_473),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_532),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_SL g661 ( 
.A(n_538),
.B(n_235),
.Y(n_661)
);

AND2x4_ASAP7_75t_L g662 ( 
.A(n_529),
.B(n_354),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_L g663 ( 
.A(n_586),
.B(n_300),
.Y(n_663)
);

CKINVDCx5p33_ASAP7_75t_R g664 ( 
.A(n_498),
.Y(n_664)
);

INVx2_ASAP7_75t_SL g665 ( 
.A(n_571),
.Y(n_665)
);

AND2x4_ASAP7_75t_L g666 ( 
.A(n_529),
.B(n_189),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_L g667 ( 
.A(n_490),
.B(n_214),
.Y(n_667)
);

BUFx3_ASAP7_75t_L g668 ( 
.A(n_606),
.Y(n_668)
);

NOR2xp33_ASAP7_75t_L g669 ( 
.A(n_552),
.B(n_290),
.Y(n_669)
);

INVx2_ASAP7_75t_L g670 ( 
.A(n_473),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_L g671 ( 
.A(n_603),
.B(n_222),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_L g672 ( 
.A(n_463),
.B(n_222),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_533),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_L g674 ( 
.A(n_571),
.B(n_224),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_L g675 ( 
.A(n_583),
.B(n_224),
.Y(n_675)
);

AND2x2_ASAP7_75t_L g676 ( 
.A(n_494),
.B(n_234),
.Y(n_676)
);

NOR2xp33_ASAP7_75t_L g677 ( 
.A(n_560),
.B(n_538),
.Y(n_677)
);

NOR2xp33_ASAP7_75t_L g678 ( 
.A(n_560),
.B(n_291),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_L g679 ( 
.A(n_592),
.B(n_234),
.Y(n_679)
);

BUFx6f_ASAP7_75t_L g680 ( 
.A(n_589),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_SL g681 ( 
.A(n_581),
.B(n_235),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_SL g682 ( 
.A(n_581),
.B(n_391),
.Y(n_682)
);

NOR3xp33_ASAP7_75t_L g683 ( 
.A(n_519),
.B(n_264),
.C(n_302),
.Y(n_683)
);

BUFx6f_ASAP7_75t_L g684 ( 
.A(n_589),
.Y(n_684)
);

INVx2_ASAP7_75t_L g685 ( 
.A(n_483),
.Y(n_685)
);

AND2x2_ASAP7_75t_L g686 ( 
.A(n_494),
.B(n_264),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_533),
.Y(n_687)
);

AND2x2_ASAP7_75t_L g688 ( 
.A(n_493),
.B(n_265),
.Y(n_688)
);

INVx2_ASAP7_75t_L g689 ( 
.A(n_483),
.Y(n_689)
);

INVx2_ASAP7_75t_SL g690 ( 
.A(n_597),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_SL g691 ( 
.A(n_581),
.B(n_391),
.Y(n_691)
);

INVx2_ASAP7_75t_SL g692 ( 
.A(n_597),
.Y(n_692)
);

NOR2xp67_ASAP7_75t_L g693 ( 
.A(n_594),
.B(n_602),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_534),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_L g695 ( 
.A(n_561),
.B(n_265),
.Y(n_695)
);

AOI22xp5_ASAP7_75t_L g696 ( 
.A1(n_487),
.A2(n_185),
.B1(n_190),
.B2(n_310),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_SL g697 ( 
.A(n_495),
.B(n_391),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_L g698 ( 
.A(n_606),
.B(n_267),
.Y(n_698)
);

INVx3_ASAP7_75t_L g699 ( 
.A(n_524),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_SL g700 ( 
.A(n_495),
.B(n_496),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_L g701 ( 
.A(n_606),
.B(n_267),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_534),
.Y(n_702)
);

BUFx6f_ASAP7_75t_SL g703 ( 
.A(n_597),
.Y(n_703)
);

OR2x2_ASAP7_75t_L g704 ( 
.A(n_543),
.B(n_271),
.Y(n_704)
);

BUFx3_ASAP7_75t_L g705 ( 
.A(n_597),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_L g706 ( 
.A(n_527),
.B(n_271),
.Y(n_706)
);

NOR2xp33_ASAP7_75t_L g707 ( 
.A(n_601),
.B(n_471),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_587),
.Y(n_708)
);

INVx2_ASAP7_75t_L g709 ( 
.A(n_492),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_L g710 ( 
.A(n_550),
.B(n_286),
.Y(n_710)
);

INVx2_ASAP7_75t_L g711 ( 
.A(n_492),
.Y(n_711)
);

BUFx6f_ASAP7_75t_L g712 ( 
.A(n_589),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_L g713 ( 
.A(n_461),
.B(n_286),
.Y(n_713)
);

INVx2_ASAP7_75t_SL g714 ( 
.A(n_515),
.Y(n_714)
);

AOI21xp5_ASAP7_75t_L g715 ( 
.A1(n_502),
.A2(n_393),
.B(n_394),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_L g716 ( 
.A(n_469),
.B(n_496),
.Y(n_716)
);

NOR2xp33_ASAP7_75t_L g717 ( 
.A(n_471),
.B(n_299),
.Y(n_717)
);

NAND2x1_ASAP7_75t_L g718 ( 
.A(n_471),
.B(n_392),
.Y(n_718)
);

AOI22xp5_ASAP7_75t_L g719 ( 
.A1(n_487),
.A2(n_175),
.B1(n_166),
.B2(n_308),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_575),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_SL g721 ( 
.A(n_476),
.B(n_513),
.Y(n_721)
);

NOR2xp33_ASAP7_75t_SL g722 ( 
.A(n_543),
.B(n_303),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_575),
.Y(n_723)
);

AND2x6_ASAP7_75t_SL g724 ( 
.A(n_593),
.B(n_295),
.Y(n_724)
);

NOR2xp33_ASAP7_75t_L g725 ( 
.A(n_478),
.B(n_306),
.Y(n_725)
);

NAND3xp33_ASAP7_75t_L g726 ( 
.A(n_602),
.B(n_307),
.C(n_302),
.Y(n_726)
);

BUFx3_ASAP7_75t_L g727 ( 
.A(n_537),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_L g728 ( 
.A(n_547),
.B(n_295),
.Y(n_728)
);

INVx3_ASAP7_75t_L g729 ( 
.A(n_524),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_580),
.Y(n_730)
);

OAI22xp5_ASAP7_75t_L g731 ( 
.A1(n_487),
.A2(n_305),
.B1(n_284),
.B2(n_250),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_SL g732 ( 
.A(n_524),
.B(n_160),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_L g733 ( 
.A(n_547),
.B(n_305),
.Y(n_733)
);

OAI22xp5_ASAP7_75t_SL g734 ( 
.A1(n_554),
.A2(n_250),
.B1(n_311),
.B2(n_284),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_580),
.Y(n_735)
);

INVx2_ASAP7_75t_L g736 ( 
.A(n_497),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_L g737 ( 
.A(n_547),
.B(n_162),
.Y(n_737)
);

NOR2xp67_ASAP7_75t_L g738 ( 
.A(n_564),
.B(n_392),
.Y(n_738)
);

AO221x1_ASAP7_75t_L g739 ( 
.A1(n_546),
.A2(n_416),
.B1(n_414),
.B2(n_425),
.C(n_394),
.Y(n_739)
);

INVx2_ASAP7_75t_L g740 ( 
.A(n_497),
.Y(n_740)
);

NOR2xp33_ASAP7_75t_L g741 ( 
.A(n_579),
.B(n_1),
.Y(n_741)
);

INVx2_ASAP7_75t_SL g742 ( 
.A(n_515),
.Y(n_742)
);

INVx4_ASAP7_75t_L g743 ( 
.A(n_507),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_L g744 ( 
.A(n_558),
.B(n_163),
.Y(n_744)
);

NAND2xp33_ASAP7_75t_L g745 ( 
.A(n_476),
.B(n_513),
.Y(n_745)
);

AOI22xp33_ASAP7_75t_L g746 ( 
.A1(n_546),
.A2(n_311),
.B1(n_284),
.B2(n_250),
.Y(n_746)
);

INVxp67_ASAP7_75t_L g747 ( 
.A(n_521),
.Y(n_747)
);

AO22x2_ASAP7_75t_L g748 ( 
.A1(n_554),
.A2(n_311),
.B1(n_3),
.B2(n_4),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_582),
.Y(n_749)
);

NOR2xp33_ASAP7_75t_L g750 ( 
.A(n_507),
.B(n_2),
.Y(n_750)
);

OAI21xp33_ASAP7_75t_L g751 ( 
.A1(n_515),
.A2(n_245),
.B(n_172),
.Y(n_751)
);

BUFx2_ASAP7_75t_L g752 ( 
.A(n_515),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_L g753 ( 
.A(n_558),
.B(n_168),
.Y(n_753)
);

INVx1_ASAP7_75t_SL g754 ( 
.A(n_536),
.Y(n_754)
);

INVx2_ASAP7_75t_L g755 ( 
.A(n_504),
.Y(n_755)
);

NOR2xp67_ASAP7_75t_L g756 ( 
.A(n_537),
.B(n_394),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_SL g757 ( 
.A(n_476),
.B(n_391),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_L g758 ( 
.A(n_558),
.B(n_176),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_L g759 ( 
.A(n_535),
.B(n_178),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_582),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_L g761 ( 
.A(n_596),
.B(n_193),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_L g762 ( 
.A(n_596),
.B(n_197),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_L g763 ( 
.A(n_600),
.B(n_199),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_L g764 ( 
.A(n_600),
.B(n_203),
.Y(n_764)
);

BUFx6f_ASAP7_75t_L g765 ( 
.A(n_476),
.Y(n_765)
);

INVx2_ASAP7_75t_L g766 ( 
.A(n_504),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_SL g767 ( 
.A(n_565),
.B(n_206),
.Y(n_767)
);

NOR2x1p5_ASAP7_75t_L g768 ( 
.A(n_565),
.B(n_207),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_SL g769 ( 
.A(n_588),
.B(n_211),
.Y(n_769)
);

AOI21xp5_ASAP7_75t_L g770 ( 
.A1(n_502),
.A2(n_470),
.B(n_468),
.Y(n_770)
);

AND2x6_ASAP7_75t_SL g771 ( 
.A(n_507),
.B(n_605),
.Y(n_771)
);

NOR2xp33_ASAP7_75t_L g772 ( 
.A(n_489),
.B(n_5),
.Y(n_772)
);

NOR2x1p5_ASAP7_75t_L g773 ( 
.A(n_588),
.B(n_212),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_658),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_L g775 ( 
.A(n_622),
.B(n_541),
.Y(n_775)
);

BUFx8_ASAP7_75t_L g776 ( 
.A(n_619),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_660),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_673),
.Y(n_778)
);

AND2x4_ASAP7_75t_L g779 ( 
.A(n_705),
.B(n_605),
.Y(n_779)
);

NOR2x2_ASAP7_75t_L g780 ( 
.A(n_664),
.B(n_539),
.Y(n_780)
);

INVx2_ASAP7_75t_L g781 ( 
.A(n_727),
.Y(n_781)
);

INVx1_ASAP7_75t_L g782 ( 
.A(n_687),
.Y(n_782)
);

AOI22xp5_ASAP7_75t_SL g783 ( 
.A1(n_649),
.A2(n_287),
.B1(n_297),
.B2(n_292),
.Y(n_783)
);

INVx2_ASAP7_75t_L g784 ( 
.A(n_610),
.Y(n_784)
);

INVx1_ASAP7_75t_L g785 ( 
.A(n_694),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_L g786 ( 
.A(n_622),
.B(n_539),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_702),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_613),
.Y(n_788)
);

BUFx3_ASAP7_75t_L g789 ( 
.A(n_615),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_L g790 ( 
.A(n_623),
.B(n_540),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_613),
.Y(n_791)
);

A2O1A1Ixp33_ASAP7_75t_L g792 ( 
.A1(n_750),
.A2(n_604),
.B(n_567),
.C(n_574),
.Y(n_792)
);

AND2x4_ASAP7_75t_L g793 ( 
.A(n_668),
.B(n_489),
.Y(n_793)
);

A2O1A1Ixp33_ASAP7_75t_L g794 ( 
.A1(n_750),
.A2(n_623),
.B(n_741),
.C(n_621),
.Y(n_794)
);

AND2x2_ASAP7_75t_SL g795 ( 
.A(n_746),
.B(n_604),
.Y(n_795)
);

AOI22xp33_ASAP7_75t_L g796 ( 
.A1(n_645),
.A2(n_746),
.B1(n_620),
.B2(n_752),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_720),
.Y(n_797)
);

BUFx2_ASAP7_75t_L g798 ( 
.A(n_662),
.Y(n_798)
);

BUFx6f_ASAP7_75t_L g799 ( 
.A(n_680),
.Y(n_799)
);

AND2x6_ASAP7_75t_SL g800 ( 
.A(n_725),
.B(n_468),
.Y(n_800)
);

NOR2xp67_ASAP7_75t_L g801 ( 
.A(n_747),
.B(n_540),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_L g802 ( 
.A(n_612),
.B(n_542),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_723),
.Y(n_803)
);

AOI22xp33_ASAP7_75t_L g804 ( 
.A1(n_645),
.A2(n_505),
.B1(n_509),
.B2(n_557),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_730),
.Y(n_805)
);

AOI22xp5_ASAP7_75t_L g806 ( 
.A1(n_612),
.A2(n_489),
.B1(n_517),
.B2(n_523),
.Y(n_806)
);

AND2x4_ASAP7_75t_L g807 ( 
.A(n_743),
.B(n_517),
.Y(n_807)
);

NOR2xp33_ASAP7_75t_R g808 ( 
.A(n_632),
.B(n_517),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_SL g809 ( 
.A(n_646),
.B(n_476),
.Y(n_809)
);

OR2x2_ASAP7_75t_L g810 ( 
.A(n_625),
.B(n_542),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_SL g811 ( 
.A(n_646),
.B(n_651),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_L g812 ( 
.A(n_621),
.B(n_545),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_SL g813 ( 
.A(n_677),
.B(n_513),
.Y(n_813)
);

CKINVDCx5p33_ASAP7_75t_R g814 ( 
.A(n_637),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_735),
.Y(n_815)
);

OR2x2_ASAP7_75t_L g816 ( 
.A(n_662),
.B(n_545),
.Y(n_816)
);

AOI22xp5_ASAP7_75t_L g817 ( 
.A1(n_722),
.A2(n_523),
.B1(n_530),
.B2(n_470),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_749),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_L g819 ( 
.A(n_708),
.B(n_557),
.Y(n_819)
);

OR2x6_ASAP7_75t_L g820 ( 
.A(n_714),
.B(n_570),
.Y(n_820)
);

INVx1_ASAP7_75t_L g821 ( 
.A(n_760),
.Y(n_821)
);

NOR2xp33_ASAP7_75t_L g822 ( 
.A(n_616),
.B(n_523),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_665),
.Y(n_823)
);

AOI22xp33_ASAP7_75t_L g824 ( 
.A1(n_620),
.A2(n_505),
.B1(n_509),
.B2(n_573),
.Y(n_824)
);

AOI21xp5_ASAP7_75t_L g825 ( 
.A1(n_721),
.A2(n_502),
.B(n_549),
.Y(n_825)
);

BUFx3_ASAP7_75t_L g826 ( 
.A(n_615),
.Y(n_826)
);

AOI22xp33_ASAP7_75t_L g827 ( 
.A1(n_748),
.A2(n_572),
.B1(n_573),
.B2(n_577),
.Y(n_827)
);

INVx5_ASAP7_75t_L g828 ( 
.A(n_680),
.Y(n_828)
);

HB1xp67_ASAP7_75t_L g829 ( 
.A(n_742),
.Y(n_829)
);

AOI22xp5_ASAP7_75t_L g830 ( 
.A1(n_634),
.A2(n_530),
.B1(n_472),
.B2(n_526),
.Y(n_830)
);

INVx3_ASAP7_75t_L g831 ( 
.A(n_680),
.Y(n_831)
);

AND2x4_ASAP7_75t_L g832 ( 
.A(n_743),
.B(n_530),
.Y(n_832)
);

NOR2xp67_ASAP7_75t_L g833 ( 
.A(n_617),
.B(n_577),
.Y(n_833)
);

BUFx3_ASAP7_75t_L g834 ( 
.A(n_615),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_L g835 ( 
.A(n_609),
.B(n_578),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_SL g836 ( 
.A(n_615),
.B(n_699),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_728),
.Y(n_837)
);

A2O1A1Ixp33_ASAP7_75t_L g838 ( 
.A1(n_741),
.A2(n_555),
.B(n_549),
.C(n_567),
.Y(n_838)
);

CKINVDCx20_ASAP7_75t_R g839 ( 
.A(n_652),
.Y(n_839)
);

BUFx2_ASAP7_75t_L g840 ( 
.A(n_771),
.Y(n_840)
);

OAI22xp5_ASAP7_75t_L g841 ( 
.A1(n_611),
.A2(n_555),
.B1(n_574),
.B2(n_472),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_L g842 ( 
.A(n_633),
.B(n_584),
.Y(n_842)
);

OR2x2_ASAP7_75t_L g843 ( 
.A(n_704),
.B(n_584),
.Y(n_843)
);

OAI22xp5_ASAP7_75t_SL g844 ( 
.A1(n_725),
.A2(n_238),
.B1(n_226),
.B2(n_231),
.Y(n_844)
);

BUFx3_ASAP7_75t_L g845 ( 
.A(n_754),
.Y(n_845)
);

INVx2_ASAP7_75t_L g846 ( 
.A(n_659),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_733),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_L g848 ( 
.A(n_634),
.B(n_474),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_L g849 ( 
.A(n_678),
.B(n_474),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_L g850 ( 
.A(n_678),
.B(n_475),
.Y(n_850)
);

INVxp67_ASAP7_75t_SL g851 ( 
.A(n_680),
.Y(n_851)
);

INVx5_ASAP7_75t_L g852 ( 
.A(n_684),
.Y(n_852)
);

INVx1_ASAP7_75t_L g853 ( 
.A(n_626),
.Y(n_853)
);

NOR2xp33_ASAP7_75t_L g854 ( 
.A(n_628),
.B(n_647),
.Y(n_854)
);

AND2x6_ASAP7_75t_SL g855 ( 
.A(n_647),
.B(n_475),
.Y(n_855)
);

INVx2_ASAP7_75t_L g856 ( 
.A(n_670),
.Y(n_856)
);

BUFx3_ASAP7_75t_L g857 ( 
.A(n_666),
.Y(n_857)
);

AND2x4_ASAP7_75t_L g858 ( 
.A(n_690),
.B(n_510),
.Y(n_858)
);

AND2x4_ASAP7_75t_L g859 ( 
.A(n_692),
.B(n_510),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_L g860 ( 
.A(n_648),
.B(n_653),
.Y(n_860)
);

OAI22xp33_ASAP7_75t_L g861 ( 
.A1(n_713),
.A2(n_512),
.B1(n_511),
.B2(n_516),
.Y(n_861)
);

INVx2_ASAP7_75t_L g862 ( 
.A(n_685),
.Y(n_862)
);

AOI22xp33_ASAP7_75t_L g863 ( 
.A1(n_748),
.A2(n_516),
.B1(n_511),
.B2(n_512),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_L g864 ( 
.A(n_648),
.B(n_477),
.Y(n_864)
);

INVx2_ASAP7_75t_L g865 ( 
.A(n_689),
.Y(n_865)
);

INVx5_ASAP7_75t_L g866 ( 
.A(n_684),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_635),
.Y(n_867)
);

AND2x4_ASAP7_75t_L g868 ( 
.A(n_699),
.B(n_477),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_636),
.Y(n_869)
);

OAI22xp5_ASAP7_75t_L g870 ( 
.A1(n_607),
.A2(n_525),
.B1(n_482),
.B2(n_486),
.Y(n_870)
);

AND2x2_ASAP7_75t_L g871 ( 
.A(n_688),
.B(n_500),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_SL g872 ( 
.A(n_729),
.B(n_513),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_SL g873 ( 
.A(n_729),
.B(n_480),
.Y(n_873)
);

O2A1O1Ixp33_ASAP7_75t_L g874 ( 
.A1(n_607),
.A2(n_520),
.B(n_480),
.C(n_482),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_L g875 ( 
.A(n_653),
.B(n_486),
.Y(n_875)
);

INVx1_ASAP7_75t_L g876 ( 
.A(n_640),
.Y(n_876)
);

BUFx6f_ASAP7_75t_L g877 ( 
.A(n_684),
.Y(n_877)
);

AOI22xp33_ASAP7_75t_L g878 ( 
.A1(n_748),
.A2(n_522),
.B1(n_500),
.B2(n_501),
.Y(n_878)
);

CKINVDCx5p33_ASAP7_75t_R g879 ( 
.A(n_619),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_650),
.Y(n_880)
);

INVx3_ASAP7_75t_L g881 ( 
.A(n_712),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_L g882 ( 
.A(n_669),
.B(n_491),
.Y(n_882)
);

AOI22xp5_ASAP7_75t_SL g883 ( 
.A1(n_731),
.A2(n_285),
.B1(n_232),
.B2(n_233),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_656),
.Y(n_884)
);

AND2x2_ASAP7_75t_L g885 ( 
.A(n_676),
.B(n_500),
.Y(n_885)
);

CKINVDCx16_ASAP7_75t_R g886 ( 
.A(n_703),
.Y(n_886)
);

AND2x2_ASAP7_75t_SL g887 ( 
.A(n_716),
.B(n_491),
.Y(n_887)
);

NOR2xp33_ASAP7_75t_L g888 ( 
.A(n_641),
.B(n_654),
.Y(n_888)
);

INVx2_ASAP7_75t_L g889 ( 
.A(n_709),
.Y(n_889)
);

INVx4_ASAP7_75t_L g890 ( 
.A(n_712),
.Y(n_890)
);

BUFx2_ASAP7_75t_L g891 ( 
.A(n_666),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_L g892 ( 
.A(n_669),
.B(n_501),
.Y(n_892)
);

OAI21xp33_ASAP7_75t_L g893 ( 
.A1(n_667),
.A2(n_525),
.B(n_506),
.Y(n_893)
);

INVx2_ASAP7_75t_SL g894 ( 
.A(n_686),
.Y(n_894)
);

INVx2_ASAP7_75t_L g895 ( 
.A(n_711),
.Y(n_895)
);

A2O1A1Ixp33_ASAP7_75t_SL g896 ( 
.A1(n_772),
.A2(n_528),
.B(n_506),
.C(n_518),
.Y(n_896)
);

NOR2xp33_ASAP7_75t_L g897 ( 
.A(n_618),
.B(n_518),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_L g898 ( 
.A(n_717),
.B(n_520),
.Y(n_898)
);

BUFx6f_ASAP7_75t_L g899 ( 
.A(n_712),
.Y(n_899)
);

NAND3xp33_ASAP7_75t_SL g900 ( 
.A(n_644),
.B(n_274),
.C(n_240),
.Y(n_900)
);

INVx1_ASAP7_75t_L g901 ( 
.A(n_736),
.Y(n_901)
);

INVx1_ASAP7_75t_L g902 ( 
.A(n_740),
.Y(n_902)
);

INVx2_ASAP7_75t_L g903 ( 
.A(n_755),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_L g904 ( 
.A(n_717),
.B(n_526),
.Y(n_904)
);

INVx2_ASAP7_75t_L g905 ( 
.A(n_766),
.Y(n_905)
);

AND2x4_ASAP7_75t_L g906 ( 
.A(n_657),
.B(n_528),
.Y(n_906)
);

INVx2_ASAP7_75t_L g907 ( 
.A(n_718),
.Y(n_907)
);

AO22x1_ASAP7_75t_L g908 ( 
.A1(n_683),
.A2(n_281),
.B1(n_241),
.B2(n_242),
.Y(n_908)
);

CKINVDCx5p33_ASAP7_75t_R g909 ( 
.A(n_703),
.Y(n_909)
);

INVx4_ASAP7_75t_L g910 ( 
.A(n_608),
.Y(n_910)
);

BUFx2_ASAP7_75t_L g911 ( 
.A(n_698),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_L g912 ( 
.A(n_675),
.B(n_585),
.Y(n_912)
);

OAI21xp33_ASAP7_75t_L g913 ( 
.A1(n_679),
.A2(n_220),
.B(n_247),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_SL g914 ( 
.A(n_618),
.B(n_624),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_L g915 ( 
.A(n_672),
.B(n_701),
.Y(n_915)
);

BUFx3_ASAP7_75t_L g916 ( 
.A(n_695),
.Y(n_916)
);

NAND2x1p5_ASAP7_75t_L g917 ( 
.A(n_608),
.B(n_576),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_L g918 ( 
.A(n_674),
.B(n_585),
.Y(n_918)
);

AND2x4_ASAP7_75t_L g919 ( 
.A(n_768),
.B(n_590),
.Y(n_919)
);

O2A1O1Ixp5_ASAP7_75t_L g920 ( 
.A1(n_614),
.A2(n_599),
.B(n_595),
.C(n_591),
.Y(n_920)
);

OAI22xp5_ASAP7_75t_L g921 ( 
.A1(n_624),
.A2(n_598),
.B1(n_576),
.B2(n_595),
.Y(n_921)
);

INVx1_ASAP7_75t_L g922 ( 
.A(n_663),
.Y(n_922)
);

AOI21xp5_ASAP7_75t_L g923 ( 
.A1(n_721),
.A2(n_627),
.B(n_629),
.Y(n_923)
);

INVxp67_ASAP7_75t_L g924 ( 
.A(n_707),
.Y(n_924)
);

INVx1_ASAP7_75t_L g925 ( 
.A(n_630),
.Y(n_925)
);

INVx2_ASAP7_75t_L g926 ( 
.A(n_765),
.Y(n_926)
);

INVx2_ASAP7_75t_L g927 ( 
.A(n_765),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_SL g928 ( 
.A(n_765),
.B(n_598),
.Y(n_928)
);

INVx2_ASAP7_75t_L g929 ( 
.A(n_765),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_L g930 ( 
.A(n_693),
.B(n_599),
.Y(n_930)
);

BUFx3_ASAP7_75t_L g931 ( 
.A(n_707),
.Y(n_931)
);

INVx5_ASAP7_75t_L g932 ( 
.A(n_724),
.Y(n_932)
);

NOR2xp33_ASAP7_75t_SL g933 ( 
.A(n_734),
.B(n_751),
.Y(n_933)
);

AND2x2_ASAP7_75t_L g934 ( 
.A(n_671),
.B(n_522),
.Y(n_934)
);

INVx4_ASAP7_75t_L g935 ( 
.A(n_739),
.Y(n_935)
);

NAND2xp5_ASAP7_75t_L g936 ( 
.A(n_710),
.B(n_591),
.Y(n_936)
);

NOR2xp33_ASAP7_75t_L g937 ( 
.A(n_627),
.B(n_590),
.Y(n_937)
);

NOR2xp33_ASAP7_75t_L g938 ( 
.A(n_629),
.B(n_598),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_L g939 ( 
.A(n_706),
.B(n_522),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_L g940 ( 
.A(n_696),
.B(n_719),
.Y(n_940)
);

BUFx3_ASAP7_75t_L g941 ( 
.A(n_772),
.Y(n_941)
);

BUFx2_ASAP7_75t_L g942 ( 
.A(n_726),
.Y(n_942)
);

INVx1_ASAP7_75t_L g943 ( 
.A(n_756),
.Y(n_943)
);

BUFx6f_ASAP7_75t_L g944 ( 
.A(n_682),
.Y(n_944)
);

INVx1_ASAP7_75t_L g945 ( 
.A(n_761),
.Y(n_945)
);

INVx2_ASAP7_75t_L g946 ( 
.A(n_643),
.Y(n_946)
);

INVx2_ASAP7_75t_L g947 ( 
.A(n_697),
.Y(n_947)
);

INVxp67_ASAP7_75t_L g948 ( 
.A(n_738),
.Y(n_948)
);

NOR2xp33_ASAP7_75t_L g949 ( 
.A(n_732),
.B(n_598),
.Y(n_949)
);

AOI22xp33_ASAP7_75t_L g950 ( 
.A1(n_681),
.A2(n_773),
.B1(n_655),
.B2(n_700),
.Y(n_950)
);

BUFx6f_ASAP7_75t_L g951 ( 
.A(n_682),
.Y(n_951)
);

NAND2x1p5_ASAP7_75t_L g952 ( 
.A(n_700),
.B(n_576),
.Y(n_952)
);

INVx1_ASAP7_75t_L g953 ( 
.A(n_762),
.Y(n_953)
);

AND2x2_ASAP7_75t_L g954 ( 
.A(n_763),
.B(n_425),
.Y(n_954)
);

NAND2xp5_ASAP7_75t_L g955 ( 
.A(n_775),
.B(n_764),
.Y(n_955)
);

INVx1_ASAP7_75t_SL g956 ( 
.A(n_839),
.Y(n_956)
);

BUFx6f_ASAP7_75t_L g957 ( 
.A(n_789),
.Y(n_957)
);

NAND2xp5_ASAP7_75t_SL g958 ( 
.A(n_860),
.B(n_737),
.Y(n_958)
);

INVx1_ASAP7_75t_L g959 ( 
.A(n_774),
.Y(n_959)
);

OAI22xp5_ASAP7_75t_L g960 ( 
.A1(n_794),
.A2(n_642),
.B1(n_631),
.B2(n_638),
.Y(n_960)
);

AOI21xp5_ASAP7_75t_L g961 ( 
.A1(n_838),
.A2(n_745),
.B(n_770),
.Y(n_961)
);

AOI21xp5_ASAP7_75t_L g962 ( 
.A1(n_838),
.A2(n_631),
.B(n_638),
.Y(n_962)
);

INVx1_ASAP7_75t_L g963 ( 
.A(n_777),
.Y(n_963)
);

BUFx2_ASAP7_75t_L g964 ( 
.A(n_798),
.Y(n_964)
);

NOR3xp33_ASAP7_75t_SL g965 ( 
.A(n_879),
.B(n_759),
.C(n_758),
.Y(n_965)
);

NAND2xp5_ASAP7_75t_L g966 ( 
.A(n_794),
.B(n_639),
.Y(n_966)
);

NAND2xp5_ASAP7_75t_L g967 ( 
.A(n_915),
.B(n_639),
.Y(n_967)
);

NAND2xp5_ASAP7_75t_SL g968 ( 
.A(n_854),
.B(n_744),
.Y(n_968)
);

O2A1O1Ixp5_ASAP7_75t_L g969 ( 
.A1(n_813),
.A2(n_661),
.B(n_642),
.C(n_757),
.Y(n_969)
);

AO21x1_ASAP7_75t_L g970 ( 
.A1(n_811),
.A2(n_875),
.B(n_864),
.Y(n_970)
);

AND2x2_ASAP7_75t_L g971 ( 
.A(n_891),
.B(n_753),
.Y(n_971)
);

NOR2xp33_ASAP7_75t_L g972 ( 
.A(n_854),
.B(n_767),
.Y(n_972)
);

AND2x4_ASAP7_75t_SL g973 ( 
.A(n_779),
.B(n_576),
.Y(n_973)
);

A2O1A1Ixp33_ASAP7_75t_L g974 ( 
.A1(n_924),
.A2(n_661),
.B(n_681),
.C(n_697),
.Y(n_974)
);

OAI22xp5_ASAP7_75t_L g975 ( 
.A1(n_796),
.A2(n_757),
.B1(n_769),
.B2(n_691),
.Y(n_975)
);

A2O1A1Ixp33_ASAP7_75t_L g976 ( 
.A1(n_924),
.A2(n_691),
.B(n_715),
.C(n_576),
.Y(n_976)
);

CKINVDCx5p33_ASAP7_75t_R g977 ( 
.A(n_776),
.Y(n_977)
);

OR2x2_ASAP7_75t_L g978 ( 
.A(n_894),
.B(n_425),
.Y(n_978)
);

O2A1O1Ixp33_ASAP7_75t_L g979 ( 
.A1(n_940),
.A2(n_393),
.B(n_9),
.C(n_11),
.Y(n_979)
);

OR2x2_ASAP7_75t_L g980 ( 
.A(n_857),
.B(n_425),
.Y(n_980)
);

BUFx12f_ASAP7_75t_L g981 ( 
.A(n_776),
.Y(n_981)
);

NOR2xp33_ASAP7_75t_L g982 ( 
.A(n_945),
.B(n_249),
.Y(n_982)
);

INVxp67_ASAP7_75t_L g983 ( 
.A(n_810),
.Y(n_983)
);

AOI21xp5_ASAP7_75t_L g984 ( 
.A1(n_882),
.A2(n_892),
.B(n_841),
.Y(n_984)
);

BUFx12f_ASAP7_75t_L g985 ( 
.A(n_909),
.Y(n_985)
);

OR2x2_ASAP7_75t_L g986 ( 
.A(n_911),
.B(n_425),
.Y(n_986)
);

NOR2xp33_ASAP7_75t_R g987 ( 
.A(n_814),
.B(n_254),
.Y(n_987)
);

OAI22xp5_ASAP7_75t_SL g988 ( 
.A1(n_844),
.A2(n_255),
.B1(n_260),
.B2(n_272),
.Y(n_988)
);

INVx5_ASAP7_75t_L g989 ( 
.A(n_820),
.Y(n_989)
);

BUFx6f_ASAP7_75t_L g990 ( 
.A(n_789),
.Y(n_990)
);

NAND2xp5_ASAP7_75t_L g991 ( 
.A(n_788),
.B(n_5),
.Y(n_991)
);

INVx1_ASAP7_75t_SL g992 ( 
.A(n_845),
.Y(n_992)
);

A2O1A1Ixp33_ASAP7_75t_L g993 ( 
.A1(n_888),
.A2(n_393),
.B(n_416),
.C(n_414),
.Y(n_993)
);

NAND2xp5_ASAP7_75t_L g994 ( 
.A(n_791),
.B(n_9),
.Y(n_994)
);

OAI22xp5_ASAP7_75t_L g995 ( 
.A1(n_796),
.A2(n_280),
.B1(n_273),
.B2(n_414),
.Y(n_995)
);

INVx4_ASAP7_75t_L g996 ( 
.A(n_828),
.Y(n_996)
);

AOI21xp5_ASAP7_75t_L g997 ( 
.A1(n_898),
.A2(n_904),
.B(n_848),
.Y(n_997)
);

CKINVDCx11_ASAP7_75t_R g998 ( 
.A(n_886),
.Y(n_998)
);

NOR2xp33_ASAP7_75t_L g999 ( 
.A(n_953),
.B(n_13),
.Y(n_999)
);

BUFx2_ASAP7_75t_L g1000 ( 
.A(n_808),
.Y(n_1000)
);

INVx2_ASAP7_75t_L g1001 ( 
.A(n_784),
.Y(n_1001)
);

INVx4_ASAP7_75t_L g1002 ( 
.A(n_828),
.Y(n_1002)
);

AND2x2_ASAP7_75t_L g1003 ( 
.A(n_783),
.B(n_425),
.Y(n_1003)
);

HB1xp67_ASAP7_75t_L g1004 ( 
.A(n_843),
.Y(n_1004)
);

O2A1O1Ixp33_ASAP7_75t_L g1005 ( 
.A1(n_888),
.A2(n_16),
.B(n_17),
.C(n_18),
.Y(n_1005)
);

NAND2xp5_ASAP7_75t_L g1006 ( 
.A(n_916),
.B(n_18),
.Y(n_1006)
);

HB1xp67_ASAP7_75t_L g1007 ( 
.A(n_816),
.Y(n_1007)
);

NAND2xp5_ASAP7_75t_L g1008 ( 
.A(n_829),
.B(n_931),
.Y(n_1008)
);

INVx1_ASAP7_75t_L g1009 ( 
.A(n_778),
.Y(n_1009)
);

AOI21xp5_ASAP7_75t_L g1010 ( 
.A1(n_790),
.A2(n_396),
.B(n_391),
.Y(n_1010)
);

INVx1_ASAP7_75t_L g1011 ( 
.A(n_782),
.Y(n_1011)
);

A2O1A1Ixp33_ASAP7_75t_L g1012 ( 
.A1(n_897),
.A2(n_425),
.B(n_416),
.C(n_414),
.Y(n_1012)
);

INVx1_ASAP7_75t_L g1013 ( 
.A(n_785),
.Y(n_1013)
);

O2A1O1Ixp5_ASAP7_75t_SL g1014 ( 
.A1(n_948),
.A2(n_416),
.B(n_414),
.C(n_396),
.Y(n_1014)
);

NOR3xp33_ASAP7_75t_SL g1015 ( 
.A(n_900),
.B(n_19),
.C(n_21),
.Y(n_1015)
);

NOR2xp33_ASAP7_75t_L g1016 ( 
.A(n_931),
.B(n_22),
.Y(n_1016)
);

OAI21x1_ASAP7_75t_L g1017 ( 
.A1(n_825),
.A2(n_416),
.B(n_414),
.Y(n_1017)
);

NOR2xp33_ASAP7_75t_R g1018 ( 
.A(n_855),
.B(n_75),
.Y(n_1018)
);

OAI21x1_ASAP7_75t_L g1019 ( 
.A1(n_920),
.A2(n_416),
.B(n_396),
.Y(n_1019)
);

OAI22xp5_ASAP7_75t_L g1020 ( 
.A1(n_795),
.A2(n_416),
.B1(n_28),
.B2(n_29),
.Y(n_1020)
);

BUFx6f_ASAP7_75t_L g1021 ( 
.A(n_826),
.Y(n_1021)
);

INVxp67_ASAP7_75t_L g1022 ( 
.A(n_823),
.Y(n_1022)
);

AOI22xp33_ASAP7_75t_L g1023 ( 
.A1(n_795),
.A2(n_396),
.B1(n_391),
.B2(n_32),
.Y(n_1023)
);

AOI21xp5_ASAP7_75t_L g1024 ( 
.A1(n_849),
.A2(n_391),
.B(n_396),
.Y(n_1024)
);

NOR2xp33_ASAP7_75t_R g1025 ( 
.A(n_900),
.B(n_80),
.Y(n_1025)
);

NOR2x1p5_ASAP7_75t_L g1026 ( 
.A(n_935),
.B(n_396),
.Y(n_1026)
);

NAND2xp5_ASAP7_75t_SL g1027 ( 
.A(n_808),
.B(n_396),
.Y(n_1027)
);

INVx1_ASAP7_75t_L g1028 ( 
.A(n_787),
.Y(n_1028)
);

HB1xp67_ASAP7_75t_L g1029 ( 
.A(n_779),
.Y(n_1029)
);

AOI21xp5_ASAP7_75t_L g1030 ( 
.A1(n_850),
.A2(n_70),
.B(n_143),
.Y(n_1030)
);

INVx1_ASAP7_75t_L g1031 ( 
.A(n_797),
.Y(n_1031)
);

NAND3xp33_ASAP7_75t_L g1032 ( 
.A(n_883),
.B(n_24),
.C(n_28),
.Y(n_1032)
);

AND2x2_ASAP7_75t_L g1033 ( 
.A(n_932),
.B(n_33),
.Y(n_1033)
);

NAND2xp5_ASAP7_75t_SL g1034 ( 
.A(n_802),
.B(n_35),
.Y(n_1034)
);

AND2x2_ASAP7_75t_L g1035 ( 
.A(n_932),
.B(n_38),
.Y(n_1035)
);

O2A1O1Ixp5_ASAP7_75t_SL g1036 ( 
.A1(n_948),
.A2(n_38),
.B(n_39),
.C(n_41),
.Y(n_1036)
);

NAND2xp5_ASAP7_75t_L g1037 ( 
.A(n_829),
.B(n_42),
.Y(n_1037)
);

AOI21xp5_ASAP7_75t_L g1038 ( 
.A1(n_939),
.A2(n_97),
.B(n_136),
.Y(n_1038)
);

NAND2xp5_ASAP7_75t_L g1039 ( 
.A(n_812),
.B(n_42),
.Y(n_1039)
);

INVx1_ASAP7_75t_L g1040 ( 
.A(n_803),
.Y(n_1040)
);

HB1xp67_ASAP7_75t_L g1041 ( 
.A(n_781),
.Y(n_1041)
);

AOI22xp5_ASAP7_75t_L g1042 ( 
.A1(n_933),
.A2(n_45),
.B1(n_49),
.B2(n_51),
.Y(n_1042)
);

NOR2xp33_ASAP7_75t_L g1043 ( 
.A(n_942),
.B(n_57),
.Y(n_1043)
);

BUFx4f_ASAP7_75t_L g1044 ( 
.A(n_807),
.Y(n_1044)
);

NAND2xp5_ASAP7_75t_L g1045 ( 
.A(n_871),
.B(n_63),
.Y(n_1045)
);

NAND2xp5_ASAP7_75t_L g1046 ( 
.A(n_885),
.B(n_64),
.Y(n_1046)
);

AOI21xp5_ASAP7_75t_L g1047 ( 
.A1(n_813),
.A2(n_65),
.B(n_84),
.Y(n_1047)
);

NOR2xp33_ASAP7_75t_L g1048 ( 
.A(n_800),
.B(n_88),
.Y(n_1048)
);

INVx1_ASAP7_75t_L g1049 ( 
.A(n_805),
.Y(n_1049)
);

NAND2xp5_ASAP7_75t_L g1050 ( 
.A(n_837),
.B(n_98),
.Y(n_1050)
);

INVx4_ASAP7_75t_L g1051 ( 
.A(n_828),
.Y(n_1051)
);

NAND2xp5_ASAP7_75t_L g1052 ( 
.A(n_847),
.B(n_103),
.Y(n_1052)
);

BUFx6f_ASAP7_75t_L g1053 ( 
.A(n_826),
.Y(n_1053)
);

NOR2xp33_ASAP7_75t_L g1054 ( 
.A(n_922),
.B(n_853),
.Y(n_1054)
);

INVx1_ASAP7_75t_L g1055 ( 
.A(n_815),
.Y(n_1055)
);

INVx1_ASAP7_75t_L g1056 ( 
.A(n_818),
.Y(n_1056)
);

NOR3xp33_ASAP7_75t_SL g1057 ( 
.A(n_913),
.B(n_104),
.C(n_106),
.Y(n_1057)
);

NAND2xp5_ASAP7_75t_SL g1058 ( 
.A(n_807),
.B(n_111),
.Y(n_1058)
);

NAND2xp5_ASAP7_75t_L g1059 ( 
.A(n_786),
.B(n_120),
.Y(n_1059)
);

NAND2xp5_ASAP7_75t_L g1060 ( 
.A(n_821),
.B(n_123),
.Y(n_1060)
);

AND2x2_ASAP7_75t_L g1061 ( 
.A(n_932),
.B(n_127),
.Y(n_1061)
);

INVx1_ASAP7_75t_L g1062 ( 
.A(n_901),
.Y(n_1062)
);

O2A1O1Ixp33_ASAP7_75t_L g1063 ( 
.A1(n_914),
.A2(n_150),
.B(n_811),
.C(n_842),
.Y(n_1063)
);

INVx1_ASAP7_75t_L g1064 ( 
.A(n_902),
.Y(n_1064)
);

OAI22xp5_ASAP7_75t_L g1065 ( 
.A1(n_863),
.A2(n_941),
.B1(n_827),
.B2(n_792),
.Y(n_1065)
);

NOR2xp33_ASAP7_75t_R g1066 ( 
.A(n_828),
.B(n_852),
.Y(n_1066)
);

NAND2xp5_ASAP7_75t_L g1067 ( 
.A(n_887),
.B(n_941),
.Y(n_1067)
);

O2A1O1Ixp33_ASAP7_75t_SL g1068 ( 
.A1(n_914),
.A2(n_872),
.B(n_896),
.C(n_809),
.Y(n_1068)
);

INVx1_ASAP7_75t_L g1069 ( 
.A(n_867),
.Y(n_1069)
);

OAI21x1_ASAP7_75t_L g1070 ( 
.A1(n_920),
.A2(n_923),
.B(n_921),
.Y(n_1070)
);

BUFx8_ASAP7_75t_L g1071 ( 
.A(n_840),
.Y(n_1071)
);

OA22x2_ASAP7_75t_L g1072 ( 
.A1(n_869),
.A2(n_880),
.B1(n_876),
.B2(n_884),
.Y(n_1072)
);

NAND2xp5_ASAP7_75t_SL g1073 ( 
.A(n_832),
.B(n_793),
.Y(n_1073)
);

A2O1A1Ixp33_ASAP7_75t_L g1074 ( 
.A1(n_949),
.A2(n_893),
.B(n_938),
.C(n_934),
.Y(n_1074)
);

AOI21xp5_ASAP7_75t_L g1075 ( 
.A1(n_928),
.A2(n_835),
.B(n_912),
.Y(n_1075)
);

NOR2xp33_ASAP7_75t_L g1076 ( 
.A(n_935),
.B(n_793),
.Y(n_1076)
);

NAND2xp5_ASAP7_75t_SL g1077 ( 
.A(n_832),
.B(n_910),
.Y(n_1077)
);

INVx2_ASAP7_75t_L g1078 ( 
.A(n_846),
.Y(n_1078)
);

INVx2_ASAP7_75t_L g1079 ( 
.A(n_856),
.Y(n_1079)
);

CKINVDCx6p67_ASAP7_75t_R g1080 ( 
.A(n_932),
.Y(n_1080)
);

INVx4_ASAP7_75t_L g1081 ( 
.A(n_852),
.Y(n_1081)
);

CKINVDCx20_ASAP7_75t_R g1082 ( 
.A(n_834),
.Y(n_1082)
);

NAND2x1p5_ASAP7_75t_L g1083 ( 
.A(n_834),
.B(n_852),
.Y(n_1083)
);

AOI21xp5_ASAP7_75t_L g1084 ( 
.A1(n_896),
.A2(n_918),
.B(n_872),
.Y(n_1084)
);

NAND2xp5_ASAP7_75t_SL g1085 ( 
.A(n_910),
.B(n_852),
.Y(n_1085)
);

AND2x4_ASAP7_75t_L g1086 ( 
.A(n_820),
.B(n_866),
.Y(n_1086)
);

HB1xp67_ASAP7_75t_L g1087 ( 
.A(n_820),
.Y(n_1087)
);

INVx2_ASAP7_75t_L g1088 ( 
.A(n_862),
.Y(n_1088)
);

AND2x4_ASAP7_75t_L g1089 ( 
.A(n_866),
.B(n_833),
.Y(n_1089)
);

AOI21xp5_ASAP7_75t_L g1090 ( 
.A1(n_936),
.A2(n_819),
.B(n_836),
.Y(n_1090)
);

AOI22xp33_ASAP7_75t_L g1091 ( 
.A1(n_863),
.A2(n_827),
.B1(n_887),
.B2(n_895),
.Y(n_1091)
);

INVx4_ASAP7_75t_L g1092 ( 
.A(n_866),
.Y(n_1092)
);

INVx1_ASAP7_75t_L g1093 ( 
.A(n_865),
.Y(n_1093)
);

O2A1O1Ixp33_ASAP7_75t_SL g1094 ( 
.A1(n_873),
.A2(n_836),
.B(n_938),
.C(n_870),
.Y(n_1094)
);

NOR2xp33_ASAP7_75t_R g1095 ( 
.A(n_866),
.B(n_799),
.Y(n_1095)
);

NOR2xp33_ASAP7_75t_R g1096 ( 
.A(n_799),
.B(n_899),
.Y(n_1096)
);

OAI22xp5_ASAP7_75t_L g1097 ( 
.A1(n_806),
.A2(n_878),
.B1(n_830),
.B2(n_925),
.Y(n_1097)
);

NOR2xp33_ASAP7_75t_L g1098 ( 
.A(n_822),
.B(n_930),
.Y(n_1098)
);

O2A1O1Ixp33_ASAP7_75t_L g1099 ( 
.A1(n_822),
.A2(n_873),
.B(n_874),
.C(n_937),
.Y(n_1099)
);

A2O1A1Ixp33_ASAP7_75t_L g1100 ( 
.A1(n_949),
.A2(n_937),
.B(n_950),
.C(n_947),
.Y(n_1100)
);

BUFx6f_ASAP7_75t_L g1101 ( 
.A(n_799),
.Y(n_1101)
);

NAND2xp5_ASAP7_75t_L g1102 ( 
.A(n_955),
.B(n_908),
.Y(n_1102)
);

NOR4xp25_ASAP7_75t_L g1103 ( 
.A(n_1020),
.B(n_878),
.C(n_861),
.D(n_950),
.Y(n_1103)
);

OA22x2_ASAP7_75t_L g1104 ( 
.A1(n_956),
.A2(n_919),
.B1(n_943),
.B2(n_859),
.Y(n_1104)
);

OAI21xp5_ASAP7_75t_SL g1105 ( 
.A1(n_1020),
.A2(n_817),
.B(n_868),
.Y(n_1105)
);

OAI21x1_ASAP7_75t_L g1106 ( 
.A1(n_1019),
.A2(n_952),
.B(n_946),
.Y(n_1106)
);

INVx1_ASAP7_75t_L g1107 ( 
.A(n_963),
.Y(n_1107)
);

NAND2xp5_ASAP7_75t_SL g1108 ( 
.A(n_972),
.B(n_868),
.Y(n_1108)
);

BUFx2_ASAP7_75t_L g1109 ( 
.A(n_956),
.Y(n_1109)
);

BUFx6f_ASAP7_75t_L g1110 ( 
.A(n_1044),
.Y(n_1110)
);

BUFx3_ASAP7_75t_L g1111 ( 
.A(n_985),
.Y(n_1111)
);

OAI21x1_ASAP7_75t_L g1112 ( 
.A1(n_1017),
.A2(n_952),
.B(n_954),
.Y(n_1112)
);

NAND2xp5_ASAP7_75t_L g1113 ( 
.A(n_1098),
.B(n_927),
.Y(n_1113)
);

BUFx10_ASAP7_75t_L g1114 ( 
.A(n_977),
.Y(n_1114)
);

AOI21xp5_ASAP7_75t_L g1115 ( 
.A1(n_961),
.A2(n_958),
.B(n_966),
.Y(n_1115)
);

AOI21xp5_ASAP7_75t_L g1116 ( 
.A1(n_966),
.A2(n_851),
.B(n_926),
.Y(n_1116)
);

INVx2_ASAP7_75t_SL g1117 ( 
.A(n_1082),
.Y(n_1117)
);

OAI21x1_ASAP7_75t_L g1118 ( 
.A1(n_1070),
.A2(n_917),
.B(n_929),
.Y(n_1118)
);

A2O1A1Ixp33_ASAP7_75t_L g1119 ( 
.A1(n_999),
.A2(n_801),
.B(n_919),
.C(n_906),
.Y(n_1119)
);

OAI21x1_ASAP7_75t_SL g1120 ( 
.A1(n_1067),
.A2(n_907),
.B(n_890),
.Y(n_1120)
);

NAND2xp5_ASAP7_75t_SL g1121 ( 
.A(n_1044),
.B(n_951),
.Y(n_1121)
);

NOR2xp33_ASAP7_75t_L g1122 ( 
.A(n_1008),
.B(n_1016),
.Y(n_1122)
);

NAND2xp5_ASAP7_75t_L g1123 ( 
.A(n_1004),
.B(n_859),
.Y(n_1123)
);

NOR2xp33_ASAP7_75t_R g1124 ( 
.A(n_998),
.B(n_877),
.Y(n_1124)
);

AOI21xp5_ASAP7_75t_L g1125 ( 
.A1(n_1075),
.A2(n_917),
.B(n_906),
.Y(n_1125)
);

OR2x2_ASAP7_75t_L g1126 ( 
.A(n_983),
.B(n_905),
.Y(n_1126)
);

OAI21x1_ASAP7_75t_L g1127 ( 
.A1(n_1010),
.A2(n_824),
.B(n_881),
.Y(n_1127)
);

OAI21x1_ASAP7_75t_L g1128 ( 
.A1(n_1024),
.A2(n_824),
.B(n_881),
.Y(n_1128)
);

INVx2_ASAP7_75t_L g1129 ( 
.A(n_1001),
.Y(n_1129)
);

AOI21xp5_ASAP7_75t_L g1130 ( 
.A1(n_1094),
.A2(n_951),
.B(n_944),
.Y(n_1130)
);

INVxp67_ASAP7_75t_SL g1131 ( 
.A(n_1029),
.Y(n_1131)
);

NAND2xp5_ASAP7_75t_L g1132 ( 
.A(n_1007),
.B(n_858),
.Y(n_1132)
);

BUFx5_ASAP7_75t_L g1133 ( 
.A(n_1086),
.Y(n_1133)
);

NAND2xp5_ASAP7_75t_L g1134 ( 
.A(n_992),
.B(n_858),
.Y(n_1134)
);

AOI22xp5_ASAP7_75t_L g1135 ( 
.A1(n_1065),
.A2(n_1042),
.B1(n_1023),
.B2(n_1043),
.Y(n_1135)
);

NAND2xp5_ASAP7_75t_L g1136 ( 
.A(n_992),
.B(n_889),
.Y(n_1136)
);

AND2x2_ASAP7_75t_L g1137 ( 
.A(n_964),
.B(n_903),
.Y(n_1137)
);

AOI21xp33_ASAP7_75t_L g1138 ( 
.A1(n_1097),
.A2(n_951),
.B(n_944),
.Y(n_1138)
);

AOI21xp5_ASAP7_75t_L g1139 ( 
.A1(n_1059),
.A2(n_951),
.B(n_944),
.Y(n_1139)
);

BUFx6f_ASAP7_75t_L g1140 ( 
.A(n_957),
.Y(n_1140)
);

NAND2xp5_ASAP7_75t_L g1141 ( 
.A(n_1054),
.B(n_944),
.Y(n_1141)
);

OAI22xp5_ASAP7_75t_L g1142 ( 
.A1(n_1065),
.A2(n_804),
.B1(n_799),
.B2(n_877),
.Y(n_1142)
);

AND2x2_ASAP7_75t_L g1143 ( 
.A(n_987),
.B(n_804),
.Y(n_1143)
);

INVx5_ASAP7_75t_L g1144 ( 
.A(n_989),
.Y(n_1144)
);

INVx1_ASAP7_75t_L g1145 ( 
.A(n_1009),
.Y(n_1145)
);

NAND2xp5_ASAP7_75t_L g1146 ( 
.A(n_971),
.B(n_831),
.Y(n_1146)
);

INVx6_ASAP7_75t_L g1147 ( 
.A(n_1071),
.Y(n_1147)
);

AOI21x1_ASAP7_75t_L g1148 ( 
.A1(n_1084),
.A2(n_780),
.B(n_831),
.Y(n_1148)
);

NOR4xp25_ASAP7_75t_L g1149 ( 
.A(n_1005),
.B(n_890),
.C(n_899),
.D(n_877),
.Y(n_1149)
);

AOI211x1_ASAP7_75t_L g1150 ( 
.A1(n_1032),
.A2(n_877),
.B(n_899),
.C(n_991),
.Y(n_1150)
);

OAI21x1_ASAP7_75t_L g1151 ( 
.A1(n_1014),
.A2(n_962),
.B(n_1090),
.Y(n_1151)
);

INVx3_ASAP7_75t_L g1152 ( 
.A(n_1086),
.Y(n_1152)
);

INVx4_ASAP7_75t_L g1153 ( 
.A(n_996),
.Y(n_1153)
);

OAI21x1_ASAP7_75t_L g1154 ( 
.A1(n_1063),
.A2(n_899),
.B(n_969),
.Y(n_1154)
);

A2O1A1Ixp33_ASAP7_75t_L g1155 ( 
.A1(n_982),
.A2(n_1039),
.B(n_1057),
.C(n_979),
.Y(n_1155)
);

NOR2xp33_ASAP7_75t_L g1156 ( 
.A(n_1076),
.B(n_988),
.Y(n_1156)
);

BUFx6f_ASAP7_75t_L g1157 ( 
.A(n_957),
.Y(n_1157)
);

NOR2x1_ASAP7_75t_SL g1158 ( 
.A(n_989),
.B(n_996),
.Y(n_1158)
);

AOI21xp33_ASAP7_75t_L g1159 ( 
.A1(n_1097),
.A2(n_995),
.B(n_1045),
.Y(n_1159)
);

OAI21x1_ASAP7_75t_L g1160 ( 
.A1(n_1047),
.A2(n_960),
.B(n_1038),
.Y(n_1160)
);

OAI21x1_ASAP7_75t_L g1161 ( 
.A1(n_960),
.A2(n_1099),
.B(n_1030),
.Y(n_1161)
);

NAND2xp5_ASAP7_75t_L g1162 ( 
.A(n_967),
.B(n_1091),
.Y(n_1162)
);

OAI21x1_ASAP7_75t_L g1163 ( 
.A1(n_1046),
.A2(n_970),
.B(n_1045),
.Y(n_1163)
);

OAI21x1_ASAP7_75t_SL g1164 ( 
.A1(n_967),
.A2(n_1037),
.B(n_1060),
.Y(n_1164)
);

OAI21x1_ASAP7_75t_L g1165 ( 
.A1(n_1046),
.A2(n_1072),
.B(n_1050),
.Y(n_1165)
);

OAI21x1_ASAP7_75t_L g1166 ( 
.A1(n_1072),
.A2(n_1050),
.B(n_1052),
.Y(n_1166)
);

INVxp67_ASAP7_75t_SL g1167 ( 
.A(n_973),
.Y(n_1167)
);

NAND2xp5_ASAP7_75t_L g1168 ( 
.A(n_1100),
.B(n_1011),
.Y(n_1168)
);

OR2x6_ASAP7_75t_L g1169 ( 
.A(n_1073),
.B(n_1089),
.Y(n_1169)
);

OA21x2_ASAP7_75t_L g1170 ( 
.A1(n_1074),
.A2(n_993),
.B(n_1012),
.Y(n_1170)
);

NOR2xp33_ASAP7_75t_SL g1171 ( 
.A(n_989),
.B(n_1048),
.Y(n_1171)
);

INVx1_ASAP7_75t_L g1172 ( 
.A(n_1013),
.Y(n_1172)
);

OAI21xp33_ASAP7_75t_SL g1173 ( 
.A1(n_1026),
.A2(n_968),
.B(n_1034),
.Y(n_1173)
);

INVx1_ASAP7_75t_L g1174 ( 
.A(n_1028),
.Y(n_1174)
);

INVx1_ASAP7_75t_L g1175 ( 
.A(n_1031),
.Y(n_1175)
);

OAI22xp5_ASAP7_75t_L g1176 ( 
.A1(n_1040),
.A2(n_1049),
.B1(n_1056),
.B2(n_1055),
.Y(n_1176)
);

NAND2xp5_ASAP7_75t_L g1177 ( 
.A(n_989),
.B(n_975),
.Y(n_1177)
);

OAI21x1_ASAP7_75t_SL g1178 ( 
.A1(n_1052),
.A2(n_994),
.B(n_975),
.Y(n_1178)
);

AND2x2_ASAP7_75t_L g1179 ( 
.A(n_1033),
.B(n_1035),
.Y(n_1179)
);

NAND2xp5_ASAP7_75t_L g1180 ( 
.A(n_1093),
.B(n_1069),
.Y(n_1180)
);

INVx1_ASAP7_75t_L g1181 ( 
.A(n_1062),
.Y(n_1181)
);

AOI21x1_ASAP7_75t_L g1182 ( 
.A1(n_1027),
.A2(n_1003),
.B(n_1087),
.Y(n_1182)
);

BUFx2_ASAP7_75t_L g1183 ( 
.A(n_1096),
.Y(n_1183)
);

OAI21x1_ASAP7_75t_L g1184 ( 
.A1(n_1083),
.A2(n_1036),
.B(n_1058),
.Y(n_1184)
);

NOR2xp33_ASAP7_75t_R g1185 ( 
.A(n_981),
.B(n_1080),
.Y(n_1185)
);

OAI22xp5_ASAP7_75t_L g1186 ( 
.A1(n_1015),
.A2(n_1006),
.B1(n_974),
.B2(n_995),
.Y(n_1186)
);

OAI21x1_ASAP7_75t_L g1187 ( 
.A1(n_1083),
.A2(n_1085),
.B(n_1064),
.Y(n_1187)
);

INVx2_ASAP7_75t_SL g1188 ( 
.A(n_1071),
.Y(n_1188)
);

AND2x2_ASAP7_75t_L g1189 ( 
.A(n_1041),
.B(n_1022),
.Y(n_1189)
);

AOI21xp5_ASAP7_75t_L g1190 ( 
.A1(n_1068),
.A2(n_976),
.B(n_1077),
.Y(n_1190)
);

NOR2xp67_ASAP7_75t_L g1191 ( 
.A(n_1002),
.B(n_1051),
.Y(n_1191)
);

NOR2xp33_ASAP7_75t_L g1192 ( 
.A(n_1000),
.B(n_957),
.Y(n_1192)
);

AOI21xp5_ASAP7_75t_L g1193 ( 
.A1(n_1101),
.A2(n_1081),
.B(n_1051),
.Y(n_1193)
);

BUFx3_ASAP7_75t_L g1194 ( 
.A(n_990),
.Y(n_1194)
);

AO31x2_ASAP7_75t_L g1195 ( 
.A1(n_1078),
.A2(n_1079),
.A3(n_1088),
.B(n_1002),
.Y(n_1195)
);

OAI21xp5_ASAP7_75t_L g1196 ( 
.A1(n_965),
.A2(n_978),
.B(n_986),
.Y(n_1196)
);

NAND2xp5_ASAP7_75t_L g1197 ( 
.A(n_990),
.B(n_1021),
.Y(n_1197)
);

HB1xp67_ASAP7_75t_L g1198 ( 
.A(n_1021),
.Y(n_1198)
);

NAND3xp33_ASAP7_75t_SL g1199 ( 
.A(n_1025),
.B(n_1018),
.C(n_1061),
.Y(n_1199)
);

AND2x2_ASAP7_75t_L g1200 ( 
.A(n_1053),
.B(n_980),
.Y(n_1200)
);

O2A1O1Ixp5_ASAP7_75t_L g1201 ( 
.A1(n_1081),
.A2(n_1092),
.B(n_1089),
.C(n_1101),
.Y(n_1201)
);

OAI22x1_ASAP7_75t_L g1202 ( 
.A1(n_1092),
.A2(n_1066),
.B1(n_1095),
.B2(n_1053),
.Y(n_1202)
);

NOR2xp67_ASAP7_75t_L g1203 ( 
.A(n_1053),
.B(n_1101),
.Y(n_1203)
);

INVx1_ASAP7_75t_L g1204 ( 
.A(n_959),
.Y(n_1204)
);

AND2x2_ASAP7_75t_L g1205 ( 
.A(n_1004),
.B(n_543),
.Y(n_1205)
);

NAND2xp5_ASAP7_75t_L g1206 ( 
.A(n_955),
.B(n_794),
.Y(n_1206)
);

AOI22xp5_ASAP7_75t_L g1207 ( 
.A1(n_1020),
.A2(n_794),
.B1(n_748),
.B2(n_933),
.Y(n_1207)
);

NAND3xp33_ASAP7_75t_SL g1208 ( 
.A(n_1042),
.B(n_664),
.C(n_435),
.Y(n_1208)
);

OA21x2_ASAP7_75t_L g1209 ( 
.A1(n_1070),
.A2(n_1019),
.B(n_1084),
.Y(n_1209)
);

CKINVDCx8_ASAP7_75t_R g1210 ( 
.A(n_977),
.Y(n_1210)
);

NOR2xp33_ASAP7_75t_L g1211 ( 
.A(n_956),
.B(n_664),
.Y(n_1211)
);

A2O1A1Ixp33_ASAP7_75t_L g1212 ( 
.A1(n_972),
.A2(n_860),
.B(n_794),
.C(n_888),
.Y(n_1212)
);

CKINVDCx8_ASAP7_75t_R g1213 ( 
.A(n_977),
.Y(n_1213)
);

AO31x2_ASAP7_75t_L g1214 ( 
.A1(n_970),
.A2(n_1074),
.A3(n_1097),
.B(n_997),
.Y(n_1214)
);

AOI21xp33_ASAP7_75t_L g1215 ( 
.A1(n_1020),
.A2(n_860),
.B(n_794),
.Y(n_1215)
);

NAND2xp33_ASAP7_75t_R g1216 ( 
.A(n_987),
.B(n_401),
.Y(n_1216)
);

NAND2xp5_ASAP7_75t_L g1217 ( 
.A(n_955),
.B(n_548),
.Y(n_1217)
);

AOI21xp5_ASAP7_75t_L g1218 ( 
.A1(n_984),
.A2(n_860),
.B(n_997),
.Y(n_1218)
);

OAI21x1_ASAP7_75t_L g1219 ( 
.A1(n_1019),
.A2(n_1017),
.B(n_1070),
.Y(n_1219)
);

BUFx2_ASAP7_75t_L g1220 ( 
.A(n_956),
.Y(n_1220)
);

AND2x4_ASAP7_75t_L g1221 ( 
.A(n_1073),
.B(n_1086),
.Y(n_1221)
);

INVx1_ASAP7_75t_L g1222 ( 
.A(n_959),
.Y(n_1222)
);

INVx1_ASAP7_75t_L g1223 ( 
.A(n_959),
.Y(n_1223)
);

AOI21xp5_ASAP7_75t_L g1224 ( 
.A1(n_984),
.A2(n_860),
.B(n_997),
.Y(n_1224)
);

AO31x2_ASAP7_75t_L g1225 ( 
.A1(n_970),
.A2(n_1074),
.A3(n_1097),
.B(n_997),
.Y(n_1225)
);

BUFx2_ASAP7_75t_L g1226 ( 
.A(n_956),
.Y(n_1226)
);

NOR2x1_ASAP7_75t_L g1227 ( 
.A(n_1008),
.B(n_839),
.Y(n_1227)
);

AOI21xp5_ASAP7_75t_L g1228 ( 
.A1(n_984),
.A2(n_860),
.B(n_997),
.Y(n_1228)
);

AOI21x1_ASAP7_75t_L g1229 ( 
.A1(n_984),
.A2(n_1084),
.B(n_961),
.Y(n_1229)
);

AOI21xp5_ASAP7_75t_L g1230 ( 
.A1(n_984),
.A2(n_860),
.B(n_997),
.Y(n_1230)
);

AOI21xp5_ASAP7_75t_L g1231 ( 
.A1(n_984),
.A2(n_860),
.B(n_997),
.Y(n_1231)
);

INVx1_ASAP7_75t_L g1232 ( 
.A(n_959),
.Y(n_1232)
);

AOI22xp5_ASAP7_75t_L g1233 ( 
.A1(n_1020),
.A2(n_794),
.B1(n_748),
.B2(n_933),
.Y(n_1233)
);

INVx1_ASAP7_75t_SL g1234 ( 
.A(n_992),
.Y(n_1234)
);

NOR2xp33_ASAP7_75t_L g1235 ( 
.A(n_956),
.B(n_664),
.Y(n_1235)
);

AOI21xp5_ASAP7_75t_L g1236 ( 
.A1(n_984),
.A2(n_860),
.B(n_997),
.Y(n_1236)
);

AND2x2_ASAP7_75t_L g1237 ( 
.A(n_1004),
.B(n_543),
.Y(n_1237)
);

INVx2_ASAP7_75t_SL g1238 ( 
.A(n_956),
.Y(n_1238)
);

NAND2xp5_ASAP7_75t_L g1239 ( 
.A(n_955),
.B(n_794),
.Y(n_1239)
);

AOI211x1_ASAP7_75t_L g1240 ( 
.A1(n_1032),
.A2(n_1020),
.B(n_940),
.C(n_955),
.Y(n_1240)
);

AO31x2_ASAP7_75t_L g1241 ( 
.A1(n_970),
.A2(n_1074),
.A3(n_1097),
.B(n_997),
.Y(n_1241)
);

NOR2xp33_ASAP7_75t_L g1242 ( 
.A(n_956),
.B(n_664),
.Y(n_1242)
);

BUFx3_ASAP7_75t_L g1243 ( 
.A(n_985),
.Y(n_1243)
);

O2A1O1Ixp5_ASAP7_75t_L g1244 ( 
.A1(n_1020),
.A2(n_860),
.B(n_794),
.C(n_970),
.Y(n_1244)
);

AOI21xp5_ASAP7_75t_L g1245 ( 
.A1(n_984),
.A2(n_860),
.B(n_997),
.Y(n_1245)
);

INVx1_ASAP7_75t_L g1246 ( 
.A(n_1180),
.Y(n_1246)
);

OAI21xp5_ASAP7_75t_L g1247 ( 
.A1(n_1212),
.A2(n_1244),
.B(n_1215),
.Y(n_1247)
);

O2A1O1Ixp5_ASAP7_75t_L g1248 ( 
.A1(n_1215),
.A2(n_1159),
.B(n_1155),
.C(n_1186),
.Y(n_1248)
);

INVx1_ASAP7_75t_L g1249 ( 
.A(n_1180),
.Y(n_1249)
);

AO21x2_ASAP7_75t_L g1250 ( 
.A1(n_1159),
.A2(n_1178),
.B(n_1163),
.Y(n_1250)
);

BUFx3_ASAP7_75t_L g1251 ( 
.A(n_1183),
.Y(n_1251)
);

INVx1_ASAP7_75t_L g1252 ( 
.A(n_1176),
.Y(n_1252)
);

OA21x2_ASAP7_75t_L g1253 ( 
.A1(n_1151),
.A2(n_1161),
.B(n_1219),
.Y(n_1253)
);

NOR2xp33_ASAP7_75t_L g1254 ( 
.A(n_1122),
.B(n_1108),
.Y(n_1254)
);

INVx3_ASAP7_75t_L g1255 ( 
.A(n_1148),
.Y(n_1255)
);

BUFx3_ASAP7_75t_L g1256 ( 
.A(n_1194),
.Y(n_1256)
);

NOR2xp33_ASAP7_75t_L g1257 ( 
.A(n_1207),
.B(n_1233),
.Y(n_1257)
);

NOR2xp33_ASAP7_75t_L g1258 ( 
.A(n_1207),
.B(n_1233),
.Y(n_1258)
);

NAND2xp5_ASAP7_75t_L g1259 ( 
.A(n_1217),
.B(n_1206),
.Y(n_1259)
);

AO21x2_ASAP7_75t_L g1260 ( 
.A1(n_1164),
.A2(n_1166),
.B(n_1182),
.Y(n_1260)
);

AO32x2_ASAP7_75t_L g1261 ( 
.A1(n_1186),
.A2(n_1176),
.A3(n_1142),
.B1(n_1238),
.B2(n_1103),
.Y(n_1261)
);

AND2x2_ASAP7_75t_L g1262 ( 
.A(n_1206),
.B(n_1239),
.Y(n_1262)
);

AND2x4_ASAP7_75t_L g1263 ( 
.A(n_1152),
.B(n_1221),
.Y(n_1263)
);

OR2x6_ASAP7_75t_L g1264 ( 
.A(n_1177),
.B(n_1150),
.Y(n_1264)
);

AOI22xp33_ASAP7_75t_SL g1265 ( 
.A1(n_1143),
.A2(n_1171),
.B1(n_1156),
.B2(n_1104),
.Y(n_1265)
);

INVx1_ASAP7_75t_L g1266 ( 
.A(n_1107),
.Y(n_1266)
);

O2A1O1Ixp33_ASAP7_75t_SL g1267 ( 
.A1(n_1239),
.A2(n_1102),
.B(n_1135),
.C(n_1105),
.Y(n_1267)
);

AOI22xp33_ASAP7_75t_L g1268 ( 
.A1(n_1135),
.A2(n_1199),
.B1(n_1205),
.B2(n_1237),
.Y(n_1268)
);

OAI21x1_ASAP7_75t_L g1269 ( 
.A1(n_1229),
.A2(n_1160),
.B(n_1236),
.Y(n_1269)
);

INVx2_ASAP7_75t_L g1270 ( 
.A(n_1214),
.Y(n_1270)
);

OAI21x1_ASAP7_75t_L g1271 ( 
.A1(n_1218),
.A2(n_1245),
.B(n_1231),
.Y(n_1271)
);

OAI21x1_ASAP7_75t_L g1272 ( 
.A1(n_1224),
.A2(n_1228),
.B(n_1230),
.Y(n_1272)
);

INVx1_ASAP7_75t_L g1273 ( 
.A(n_1145),
.Y(n_1273)
);

INVx1_ASAP7_75t_L g1274 ( 
.A(n_1172),
.Y(n_1274)
);

OA21x2_ASAP7_75t_L g1275 ( 
.A1(n_1165),
.A2(n_1106),
.B(n_1177),
.Y(n_1275)
);

OAI21xp5_ASAP7_75t_L g1276 ( 
.A1(n_1173),
.A2(n_1115),
.B(n_1130),
.Y(n_1276)
);

OAI21x1_ASAP7_75t_L g1277 ( 
.A1(n_1112),
.A2(n_1118),
.B(n_1154),
.Y(n_1277)
);

INVx2_ASAP7_75t_L g1278 ( 
.A(n_1214),
.Y(n_1278)
);

HB1xp67_ASAP7_75t_L g1279 ( 
.A(n_1141),
.Y(n_1279)
);

OAI21x1_ASAP7_75t_L g1280 ( 
.A1(n_1190),
.A2(n_1127),
.B(n_1128),
.Y(n_1280)
);

AOI221xp5_ASAP7_75t_L g1281 ( 
.A1(n_1103),
.A2(n_1240),
.B1(n_1208),
.B2(n_1149),
.C(n_1222),
.Y(n_1281)
);

AND2x2_ASAP7_75t_L g1282 ( 
.A(n_1174),
.B(n_1175),
.Y(n_1282)
);

AOI22xp33_ASAP7_75t_L g1283 ( 
.A1(n_1162),
.A2(n_1179),
.B1(n_1171),
.B2(n_1129),
.Y(n_1283)
);

INVx1_ASAP7_75t_L g1284 ( 
.A(n_1204),
.Y(n_1284)
);

OAI21x1_ASAP7_75t_L g1285 ( 
.A1(n_1209),
.A2(n_1139),
.B(n_1125),
.Y(n_1285)
);

INVx1_ASAP7_75t_L g1286 ( 
.A(n_1223),
.Y(n_1286)
);

OAI21x1_ASAP7_75t_L g1287 ( 
.A1(n_1209),
.A2(n_1116),
.B(n_1184),
.Y(n_1287)
);

NAND2xp5_ASAP7_75t_L g1288 ( 
.A(n_1234),
.B(n_1137),
.Y(n_1288)
);

AO31x2_ASAP7_75t_L g1289 ( 
.A1(n_1142),
.A2(n_1162),
.A3(n_1168),
.B(n_1113),
.Y(n_1289)
);

OAI21xp33_ASAP7_75t_SL g1290 ( 
.A1(n_1168),
.A2(n_1113),
.B(n_1138),
.Y(n_1290)
);

OAI21xp5_ASAP7_75t_L g1291 ( 
.A1(n_1105),
.A2(n_1119),
.B(n_1149),
.Y(n_1291)
);

INVxp67_ASAP7_75t_L g1292 ( 
.A(n_1211),
.Y(n_1292)
);

OAI211xp5_ASAP7_75t_L g1293 ( 
.A1(n_1235),
.A2(n_1242),
.B(n_1109),
.C(n_1220),
.Y(n_1293)
);

INVx2_ASAP7_75t_L g1294 ( 
.A(n_1225),
.Y(n_1294)
);

OAI21xp5_ASAP7_75t_L g1295 ( 
.A1(n_1138),
.A2(n_1196),
.B(n_1193),
.Y(n_1295)
);

INVx1_ASAP7_75t_L g1296 ( 
.A(n_1232),
.Y(n_1296)
);

OAI21x1_ASAP7_75t_L g1297 ( 
.A1(n_1170),
.A2(n_1120),
.B(n_1187),
.Y(n_1297)
);

AOI21xp5_ASAP7_75t_SL g1298 ( 
.A1(n_1202),
.A2(n_1167),
.B(n_1158),
.Y(n_1298)
);

AOI22xp33_ASAP7_75t_SL g1299 ( 
.A1(n_1234),
.A2(n_1131),
.B1(n_1134),
.B2(n_1189),
.Y(n_1299)
);

INVx2_ASAP7_75t_L g1300 ( 
.A(n_1225),
.Y(n_1300)
);

HB1xp67_ASAP7_75t_L g1301 ( 
.A(n_1200),
.Y(n_1301)
);

INVx1_ASAP7_75t_L g1302 ( 
.A(n_1181),
.Y(n_1302)
);

O2A1O1Ixp33_ASAP7_75t_L g1303 ( 
.A1(n_1196),
.A2(n_1226),
.B(n_1146),
.C(n_1117),
.Y(n_1303)
);

OAI21x1_ASAP7_75t_L g1304 ( 
.A1(n_1170),
.A2(n_1201),
.B(n_1197),
.Y(n_1304)
);

NAND2xp5_ASAP7_75t_L g1305 ( 
.A(n_1123),
.B(n_1132),
.Y(n_1305)
);

BUFx6f_ASAP7_75t_L g1306 ( 
.A(n_1110),
.Y(n_1306)
);

INVx2_ASAP7_75t_L g1307 ( 
.A(n_1225),
.Y(n_1307)
);

OAI21x1_ASAP7_75t_L g1308 ( 
.A1(n_1197),
.A2(n_1121),
.B(n_1152),
.Y(n_1308)
);

A2O1A1Ixp33_ASAP7_75t_L g1309 ( 
.A1(n_1227),
.A2(n_1241),
.B(n_1192),
.C(n_1221),
.Y(n_1309)
);

OAI22xp5_ASAP7_75t_L g1310 ( 
.A1(n_1169),
.A2(n_1110),
.B1(n_1153),
.B2(n_1136),
.Y(n_1310)
);

OAI22xp5_ASAP7_75t_L g1311 ( 
.A1(n_1169),
.A2(n_1110),
.B1(n_1153),
.B2(n_1210),
.Y(n_1311)
);

BUFx8_ASAP7_75t_L g1312 ( 
.A(n_1188),
.Y(n_1312)
);

INVx2_ASAP7_75t_L g1313 ( 
.A(n_1241),
.Y(n_1313)
);

INVx1_ASAP7_75t_L g1314 ( 
.A(n_1126),
.Y(n_1314)
);

INVx1_ASAP7_75t_L g1315 ( 
.A(n_1198),
.Y(n_1315)
);

INVx6_ASAP7_75t_L g1316 ( 
.A(n_1144),
.Y(n_1316)
);

INVx3_ASAP7_75t_L g1317 ( 
.A(n_1241),
.Y(n_1317)
);

O2A1O1Ixp33_ASAP7_75t_SL g1318 ( 
.A1(n_1191),
.A2(n_1144),
.B(n_1124),
.C(n_1133),
.Y(n_1318)
);

OAI21xp5_ASAP7_75t_L g1319 ( 
.A1(n_1203),
.A2(n_1169),
.B(n_1216),
.Y(n_1319)
);

CKINVDCx11_ASAP7_75t_R g1320 ( 
.A(n_1213),
.Y(n_1320)
);

NAND2xp5_ASAP7_75t_L g1321 ( 
.A(n_1133),
.B(n_1140),
.Y(n_1321)
);

INVx2_ASAP7_75t_SL g1322 ( 
.A(n_1157),
.Y(n_1322)
);

INVx1_ASAP7_75t_L g1323 ( 
.A(n_1157),
.Y(n_1323)
);

INVx1_ASAP7_75t_L g1324 ( 
.A(n_1157),
.Y(n_1324)
);

INVx1_ASAP7_75t_L g1325 ( 
.A(n_1133),
.Y(n_1325)
);

NAND2xp33_ASAP7_75t_L g1326 ( 
.A(n_1133),
.B(n_1185),
.Y(n_1326)
);

OAI21x1_ASAP7_75t_L g1327 ( 
.A1(n_1133),
.A2(n_1147),
.B(n_1114),
.Y(n_1327)
);

OAI21x1_ASAP7_75t_L g1328 ( 
.A1(n_1147),
.A2(n_1114),
.B(n_1111),
.Y(n_1328)
);

INVx2_ASAP7_75t_L g1329 ( 
.A(n_1243),
.Y(n_1329)
);

INVx1_ASAP7_75t_L g1330 ( 
.A(n_1180),
.Y(n_1330)
);

OAI21x1_ASAP7_75t_L g1331 ( 
.A1(n_1229),
.A2(n_1151),
.B(n_1219),
.Y(n_1331)
);

OAI21x1_ASAP7_75t_L g1332 ( 
.A1(n_1229),
.A2(n_1151),
.B(n_1219),
.Y(n_1332)
);

HB1xp67_ASAP7_75t_L g1333 ( 
.A(n_1141),
.Y(n_1333)
);

OAI21x1_ASAP7_75t_SL g1334 ( 
.A1(n_1207),
.A2(n_1233),
.B(n_1164),
.Y(n_1334)
);

CKINVDCx5p33_ASAP7_75t_R g1335 ( 
.A(n_1216),
.Y(n_1335)
);

NAND2xp5_ASAP7_75t_L g1336 ( 
.A(n_1217),
.B(n_1122),
.Y(n_1336)
);

INVx2_ASAP7_75t_L g1337 ( 
.A(n_1195),
.Y(n_1337)
);

OAI21x1_ASAP7_75t_L g1338 ( 
.A1(n_1229),
.A2(n_1151),
.B(n_1219),
.Y(n_1338)
);

OAI21xp5_ASAP7_75t_L g1339 ( 
.A1(n_1212),
.A2(n_860),
.B(n_794),
.Y(n_1339)
);

OAI21x1_ASAP7_75t_L g1340 ( 
.A1(n_1229),
.A2(n_1151),
.B(n_1219),
.Y(n_1340)
);

NAND2xp5_ASAP7_75t_L g1341 ( 
.A(n_1217),
.B(n_1122),
.Y(n_1341)
);

OAI21x1_ASAP7_75t_L g1342 ( 
.A1(n_1229),
.A2(n_1151),
.B(n_1219),
.Y(n_1342)
);

OAI21x1_ASAP7_75t_L g1343 ( 
.A1(n_1229),
.A2(n_1151),
.B(n_1219),
.Y(n_1343)
);

INVx6_ASAP7_75t_L g1344 ( 
.A(n_1110),
.Y(n_1344)
);

AOI21x1_ASAP7_75t_L g1345 ( 
.A1(n_1229),
.A2(n_1224),
.B(n_1218),
.Y(n_1345)
);

OAI21x1_ASAP7_75t_L g1346 ( 
.A1(n_1229),
.A2(n_1151),
.B(n_1219),
.Y(n_1346)
);

INVx2_ASAP7_75t_L g1347 ( 
.A(n_1195),
.Y(n_1347)
);

OAI21x1_ASAP7_75t_L g1348 ( 
.A1(n_1229),
.A2(n_1151),
.B(n_1219),
.Y(n_1348)
);

INVx1_ASAP7_75t_L g1349 ( 
.A(n_1180),
.Y(n_1349)
);

INVx1_ASAP7_75t_L g1350 ( 
.A(n_1180),
.Y(n_1350)
);

OA21x2_ASAP7_75t_L g1351 ( 
.A1(n_1151),
.A2(n_1161),
.B(n_1163),
.Y(n_1351)
);

AOI22xp33_ASAP7_75t_L g1352 ( 
.A1(n_1207),
.A2(n_543),
.B1(n_554),
.B2(n_1233),
.Y(n_1352)
);

INVx1_ASAP7_75t_L g1353 ( 
.A(n_1180),
.Y(n_1353)
);

INVx3_ASAP7_75t_L g1354 ( 
.A(n_1148),
.Y(n_1354)
);

INVx4_ASAP7_75t_L g1355 ( 
.A(n_1144),
.Y(n_1355)
);

OR2x6_ASAP7_75t_L g1356 ( 
.A(n_1177),
.B(n_1150),
.Y(n_1356)
);

AOI22xp33_ASAP7_75t_L g1357 ( 
.A1(n_1207),
.A2(n_543),
.B1(n_554),
.B2(n_1233),
.Y(n_1357)
);

INVx2_ASAP7_75t_SL g1358 ( 
.A(n_1144),
.Y(n_1358)
);

NAND2x1p5_ASAP7_75t_L g1359 ( 
.A(n_1144),
.B(n_989),
.Y(n_1359)
);

OAI22xp33_ASAP7_75t_L g1360 ( 
.A1(n_1207),
.A2(n_1233),
.B1(n_1135),
.B2(n_933),
.Y(n_1360)
);

O2A1O1Ixp5_ASAP7_75t_L g1361 ( 
.A1(n_1215),
.A2(n_1159),
.B(n_1244),
.C(n_860),
.Y(n_1361)
);

AO31x2_ASAP7_75t_L g1362 ( 
.A1(n_1177),
.A2(n_970),
.A3(n_1097),
.B(n_1074),
.Y(n_1362)
);

AOI22xp33_ASAP7_75t_SL g1363 ( 
.A1(n_1143),
.A2(n_554),
.B1(n_543),
.B2(n_933),
.Y(n_1363)
);

BUFx4_ASAP7_75t_SL g1364 ( 
.A(n_1111),
.Y(n_1364)
);

INVx2_ASAP7_75t_L g1365 ( 
.A(n_1195),
.Y(n_1365)
);

HB1xp67_ASAP7_75t_L g1366 ( 
.A(n_1141),
.Y(n_1366)
);

OAI21x1_ASAP7_75t_L g1367 ( 
.A1(n_1229),
.A2(n_1151),
.B(n_1219),
.Y(n_1367)
);

AND2x2_ASAP7_75t_L g1368 ( 
.A(n_1122),
.B(n_1179),
.Y(n_1368)
);

NAND2xp5_ASAP7_75t_SL g1369 ( 
.A(n_1207),
.B(n_1233),
.Y(n_1369)
);

OAI21x1_ASAP7_75t_L g1370 ( 
.A1(n_1229),
.A2(n_1151),
.B(n_1219),
.Y(n_1370)
);

BUFx2_ASAP7_75t_L g1371 ( 
.A(n_1109),
.Y(n_1371)
);

OA21x2_ASAP7_75t_L g1372 ( 
.A1(n_1151),
.A2(n_1161),
.B(n_1163),
.Y(n_1372)
);

NOR2xp33_ASAP7_75t_L g1373 ( 
.A(n_1212),
.B(n_1122),
.Y(n_1373)
);

INVx1_ASAP7_75t_L g1374 ( 
.A(n_1180),
.Y(n_1374)
);

INVx1_ASAP7_75t_L g1375 ( 
.A(n_1180),
.Y(n_1375)
);

NAND2xp5_ASAP7_75t_L g1376 ( 
.A(n_1217),
.B(n_1122),
.Y(n_1376)
);

OAI21x1_ASAP7_75t_L g1377 ( 
.A1(n_1229),
.A2(n_1151),
.B(n_1219),
.Y(n_1377)
);

AOI221xp5_ASAP7_75t_SL g1378 ( 
.A1(n_1212),
.A2(n_1005),
.B1(n_1186),
.B2(n_1020),
.C(n_794),
.Y(n_1378)
);

OAI21x1_ASAP7_75t_L g1379 ( 
.A1(n_1229),
.A2(n_1151),
.B(n_1219),
.Y(n_1379)
);

NAND3x1_ASAP7_75t_L g1380 ( 
.A(n_1207),
.B(n_1233),
.C(n_1135),
.Y(n_1380)
);

NAND2x1_ASAP7_75t_L g1381 ( 
.A(n_1164),
.B(n_1120),
.Y(n_1381)
);

INVx2_ASAP7_75t_L g1382 ( 
.A(n_1195),
.Y(n_1382)
);

AND2x2_ASAP7_75t_L g1383 ( 
.A(n_1207),
.B(n_1233),
.Y(n_1383)
);

NAND2xp5_ASAP7_75t_L g1384 ( 
.A(n_1373),
.B(n_1336),
.Y(n_1384)
);

AND2x2_ASAP7_75t_L g1385 ( 
.A(n_1368),
.B(n_1301),
.Y(n_1385)
);

BUFx6f_ASAP7_75t_L g1386 ( 
.A(n_1256),
.Y(n_1386)
);

OAI22xp5_ASAP7_75t_L g1387 ( 
.A1(n_1373),
.A2(n_1380),
.B1(n_1258),
.B2(n_1257),
.Y(n_1387)
);

HB1xp67_ASAP7_75t_L g1388 ( 
.A(n_1315),
.Y(n_1388)
);

CKINVDCx20_ASAP7_75t_R g1389 ( 
.A(n_1320),
.Y(n_1389)
);

AND2x2_ASAP7_75t_L g1390 ( 
.A(n_1262),
.B(n_1371),
.Y(n_1390)
);

AOI221x1_ASAP7_75t_SL g1391 ( 
.A1(n_1360),
.A2(n_1341),
.B1(n_1376),
.B2(n_1257),
.C(n_1258),
.Y(n_1391)
);

OR2x2_ASAP7_75t_L g1392 ( 
.A(n_1288),
.B(n_1262),
.Y(n_1392)
);

AND2x2_ASAP7_75t_L g1393 ( 
.A(n_1282),
.B(n_1254),
.Y(n_1393)
);

INVx3_ASAP7_75t_L g1394 ( 
.A(n_1327),
.Y(n_1394)
);

A2O1A1Ixp33_ASAP7_75t_L g1395 ( 
.A1(n_1291),
.A2(n_1248),
.B(n_1369),
.C(n_1339),
.Y(n_1395)
);

AOI221xp5_ASAP7_75t_L g1396 ( 
.A1(n_1267),
.A2(n_1369),
.B1(n_1383),
.B2(n_1357),
.C(n_1352),
.Y(n_1396)
);

OA21x2_ASAP7_75t_L g1397 ( 
.A1(n_1331),
.A2(n_1332),
.B(n_1346),
.Y(n_1397)
);

AOI21x1_ASAP7_75t_SL g1398 ( 
.A1(n_1321),
.A2(n_1378),
.B(n_1259),
.Y(n_1398)
);

AND2x2_ASAP7_75t_L g1399 ( 
.A(n_1254),
.B(n_1383),
.Y(n_1399)
);

OAI22xp5_ASAP7_75t_L g1400 ( 
.A1(n_1380),
.A2(n_1292),
.B1(n_1363),
.B2(n_1293),
.Y(n_1400)
);

AND2x2_ASAP7_75t_L g1401 ( 
.A(n_1251),
.B(n_1268),
.Y(n_1401)
);

CKINVDCx16_ASAP7_75t_R g1402 ( 
.A(n_1256),
.Y(n_1402)
);

OR2x2_ASAP7_75t_L g1403 ( 
.A(n_1279),
.B(n_1333),
.Y(n_1403)
);

OA21x2_ASAP7_75t_L g1404 ( 
.A1(n_1331),
.A2(n_1367),
.B(n_1343),
.Y(n_1404)
);

OAI22xp5_ASAP7_75t_SL g1405 ( 
.A1(n_1335),
.A2(n_1265),
.B1(n_1329),
.B2(n_1247),
.Y(n_1405)
);

OA21x2_ASAP7_75t_L g1406 ( 
.A1(n_1332),
.A2(n_1340),
.B(n_1343),
.Y(n_1406)
);

OR2x2_ASAP7_75t_L g1407 ( 
.A(n_1366),
.B(n_1266),
.Y(n_1407)
);

CKINVDCx12_ASAP7_75t_R g1408 ( 
.A(n_1364),
.Y(n_1408)
);

OAI22xp5_ASAP7_75t_L g1409 ( 
.A1(n_1281),
.A2(n_1252),
.B1(n_1283),
.B2(n_1299),
.Y(n_1409)
);

AND2x2_ASAP7_75t_L g1410 ( 
.A(n_1273),
.B(n_1274),
.Y(n_1410)
);

AOI21x1_ASAP7_75t_SL g1411 ( 
.A1(n_1361),
.A2(n_1261),
.B(n_1351),
.Y(n_1411)
);

AND2x2_ASAP7_75t_L g1412 ( 
.A(n_1284),
.B(n_1286),
.Y(n_1412)
);

O2A1O1Ixp33_ASAP7_75t_L g1413 ( 
.A1(n_1267),
.A2(n_1334),
.B(n_1303),
.C(n_1290),
.Y(n_1413)
);

INVx1_ASAP7_75t_L g1414 ( 
.A(n_1296),
.Y(n_1414)
);

NAND2xp5_ASAP7_75t_L g1415 ( 
.A(n_1246),
.B(n_1249),
.Y(n_1415)
);

O2A1O1Ixp33_ASAP7_75t_L g1416 ( 
.A1(n_1276),
.A2(n_1295),
.B(n_1311),
.C(n_1309),
.Y(n_1416)
);

O2A1O1Ixp33_ASAP7_75t_L g1417 ( 
.A1(n_1309),
.A2(n_1326),
.B(n_1310),
.C(n_1329),
.Y(n_1417)
);

OAI22xp5_ASAP7_75t_L g1418 ( 
.A1(n_1264),
.A2(n_1356),
.B1(n_1335),
.B2(n_1330),
.Y(n_1418)
);

AOI21xp5_ASAP7_75t_L g1419 ( 
.A1(n_1271),
.A2(n_1272),
.B(n_1269),
.Y(n_1419)
);

HB1xp67_ASAP7_75t_L g1420 ( 
.A(n_1264),
.Y(n_1420)
);

HB1xp67_ASAP7_75t_L g1421 ( 
.A(n_1264),
.Y(n_1421)
);

CKINVDCx5p33_ASAP7_75t_R g1422 ( 
.A(n_1320),
.Y(n_1422)
);

OAI22xp5_ASAP7_75t_L g1423 ( 
.A1(n_1356),
.A2(n_1353),
.B1(n_1375),
.B2(n_1350),
.Y(n_1423)
);

OA21x2_ASAP7_75t_L g1424 ( 
.A1(n_1338),
.A2(n_1379),
.B(n_1377),
.Y(n_1424)
);

AND2x2_ASAP7_75t_L g1425 ( 
.A(n_1302),
.B(n_1263),
.Y(n_1425)
);

AOI21xp5_ASAP7_75t_L g1426 ( 
.A1(n_1269),
.A2(n_1285),
.B(n_1381),
.Y(n_1426)
);

NAND2xp5_ASAP7_75t_L g1427 ( 
.A(n_1349),
.B(n_1374),
.Y(n_1427)
);

INVx1_ASAP7_75t_L g1428 ( 
.A(n_1314),
.Y(n_1428)
);

INVx1_ASAP7_75t_SL g1429 ( 
.A(n_1305),
.Y(n_1429)
);

AOI21x1_ASAP7_75t_SL g1430 ( 
.A1(n_1261),
.A2(n_1372),
.B(n_1345),
.Y(n_1430)
);

A2O1A1Ixp33_ASAP7_75t_L g1431 ( 
.A1(n_1319),
.A2(n_1326),
.B(n_1317),
.C(n_1327),
.Y(n_1431)
);

NOR2xp67_ASAP7_75t_L g1432 ( 
.A(n_1355),
.B(n_1358),
.Y(n_1432)
);

NAND2xp5_ASAP7_75t_L g1433 ( 
.A(n_1323),
.B(n_1324),
.Y(n_1433)
);

BUFx2_ASAP7_75t_L g1434 ( 
.A(n_1356),
.Y(n_1434)
);

AOI21x1_ASAP7_75t_SL g1435 ( 
.A1(n_1312),
.A2(n_1253),
.B(n_1250),
.Y(n_1435)
);

OAI22xp5_ASAP7_75t_L g1436 ( 
.A1(n_1344),
.A2(n_1325),
.B1(n_1354),
.B2(n_1255),
.Y(n_1436)
);

AOI21x1_ASAP7_75t_SL g1437 ( 
.A1(n_1312),
.A2(n_1253),
.B(n_1250),
.Y(n_1437)
);

CKINVDCx5p33_ASAP7_75t_R g1438 ( 
.A(n_1312),
.Y(n_1438)
);

O2A1O1Ixp5_ASAP7_75t_L g1439 ( 
.A1(n_1317),
.A2(n_1255),
.B(n_1354),
.C(n_1300),
.Y(n_1439)
);

INVx1_ASAP7_75t_L g1440 ( 
.A(n_1289),
.Y(n_1440)
);

NAND2xp5_ASAP7_75t_L g1441 ( 
.A(n_1322),
.B(n_1289),
.Y(n_1441)
);

AND2x2_ASAP7_75t_L g1442 ( 
.A(n_1322),
.B(n_1308),
.Y(n_1442)
);

OAI22xp5_ASAP7_75t_L g1443 ( 
.A1(n_1306),
.A2(n_1316),
.B1(n_1298),
.B2(n_1359),
.Y(n_1443)
);

AND2x4_ASAP7_75t_L g1444 ( 
.A(n_1328),
.B(n_1358),
.Y(n_1444)
);

NAND2xp5_ASAP7_75t_L g1445 ( 
.A(n_1362),
.B(n_1306),
.Y(n_1445)
);

NAND2xp5_ASAP7_75t_L g1446 ( 
.A(n_1362),
.B(n_1306),
.Y(n_1446)
);

AOI21xp5_ASAP7_75t_SL g1447 ( 
.A1(n_1355),
.A2(n_1359),
.B(n_1313),
.Y(n_1447)
);

CKINVDCx5p33_ASAP7_75t_R g1448 ( 
.A(n_1316),
.Y(n_1448)
);

O2A1O1Ixp5_ASAP7_75t_L g1449 ( 
.A1(n_1270),
.A2(n_1307),
.B(n_1300),
.C(n_1294),
.Y(n_1449)
);

INVx3_ASAP7_75t_L g1450 ( 
.A(n_1308),
.Y(n_1450)
);

AOI21x1_ASAP7_75t_SL g1451 ( 
.A1(n_1338),
.A2(n_1346),
.B(n_1379),
.Y(n_1451)
);

AND2x2_ASAP7_75t_L g1452 ( 
.A(n_1328),
.B(n_1304),
.Y(n_1452)
);

AOI21x1_ASAP7_75t_SL g1453 ( 
.A1(n_1340),
.A2(n_1342),
.B(n_1370),
.Y(n_1453)
);

OAI22xp5_ASAP7_75t_L g1454 ( 
.A1(n_1316),
.A2(n_1307),
.B1(n_1278),
.B2(n_1275),
.Y(n_1454)
);

O2A1O1Ixp33_ASAP7_75t_L g1455 ( 
.A1(n_1318),
.A2(n_1278),
.B(n_1260),
.C(n_1275),
.Y(n_1455)
);

OR2x2_ASAP7_75t_L g1456 ( 
.A(n_1304),
.B(n_1275),
.Y(n_1456)
);

OA21x2_ASAP7_75t_L g1457 ( 
.A1(n_1342),
.A2(n_1370),
.B(n_1367),
.Y(n_1457)
);

OAI22xp5_ASAP7_75t_SL g1458 ( 
.A1(n_1318),
.A2(n_1337),
.B1(n_1365),
.B2(n_1347),
.Y(n_1458)
);

O2A1O1Ixp5_ASAP7_75t_L g1459 ( 
.A1(n_1382),
.A2(n_1297),
.B(n_1280),
.C(n_1277),
.Y(n_1459)
);

AND2x4_ASAP7_75t_L g1460 ( 
.A(n_1297),
.B(n_1277),
.Y(n_1460)
);

O2A1O1Ixp33_ASAP7_75t_L g1461 ( 
.A1(n_1280),
.A2(n_1212),
.B(n_794),
.C(n_1373),
.Y(n_1461)
);

NAND2xp5_ASAP7_75t_L g1462 ( 
.A(n_1348),
.B(n_1287),
.Y(n_1462)
);

AND2x2_ASAP7_75t_L g1463 ( 
.A(n_1348),
.B(n_1368),
.Y(n_1463)
);

O2A1O1Ixp33_ASAP7_75t_L g1464 ( 
.A1(n_1373),
.A2(n_1212),
.B(n_794),
.C(n_1215),
.Y(n_1464)
);

AOI21xp5_ASAP7_75t_L g1465 ( 
.A1(n_1339),
.A2(n_1224),
.B(n_1218),
.Y(n_1465)
);

AND2x2_ASAP7_75t_L g1466 ( 
.A(n_1368),
.B(n_1301),
.Y(n_1466)
);

AOI221x1_ASAP7_75t_SL g1467 ( 
.A1(n_1373),
.A2(n_164),
.B1(n_174),
.B2(n_173),
.C(n_159),
.Y(n_1467)
);

AND2x4_ASAP7_75t_L g1468 ( 
.A(n_1301),
.B(n_1251),
.Y(n_1468)
);

AOI21x1_ASAP7_75t_SL g1469 ( 
.A1(n_1336),
.A2(n_860),
.B(n_1039),
.Y(n_1469)
);

OAI31xp33_ASAP7_75t_L g1470 ( 
.A1(n_1360),
.A2(n_748),
.A3(n_1258),
.B(n_1257),
.Y(n_1470)
);

NAND2xp5_ASAP7_75t_L g1471 ( 
.A(n_1373),
.B(n_1336),
.Y(n_1471)
);

OA21x2_ASAP7_75t_L g1472 ( 
.A1(n_1331),
.A2(n_1338),
.B(n_1332),
.Y(n_1472)
);

INVx5_ASAP7_75t_L g1473 ( 
.A(n_1316),
.Y(n_1473)
);

OR2x2_ASAP7_75t_L g1474 ( 
.A(n_1301),
.B(n_1288),
.Y(n_1474)
);

NAND2xp5_ASAP7_75t_L g1475 ( 
.A(n_1373),
.B(n_1336),
.Y(n_1475)
);

BUFx2_ASAP7_75t_L g1476 ( 
.A(n_1371),
.Y(n_1476)
);

A2O1A1Ixp33_ASAP7_75t_L g1477 ( 
.A1(n_1257),
.A2(n_1258),
.B(n_1207),
.C(n_1233),
.Y(n_1477)
);

INVx2_ASAP7_75t_SL g1478 ( 
.A(n_1452),
.Y(n_1478)
);

INVxp67_ASAP7_75t_L g1479 ( 
.A(n_1441),
.Y(n_1479)
);

HB1xp67_ASAP7_75t_L g1480 ( 
.A(n_1388),
.Y(n_1480)
);

HB1xp67_ASAP7_75t_L g1481 ( 
.A(n_1456),
.Y(n_1481)
);

AND2x2_ASAP7_75t_L g1482 ( 
.A(n_1463),
.B(n_1390),
.Y(n_1482)
);

AOI22xp5_ASAP7_75t_L g1483 ( 
.A1(n_1387),
.A2(n_1477),
.B1(n_1396),
.B2(n_1400),
.Y(n_1483)
);

BUFx6f_ASAP7_75t_L g1484 ( 
.A(n_1460),
.Y(n_1484)
);

BUFx2_ASAP7_75t_L g1485 ( 
.A(n_1460),
.Y(n_1485)
);

INVx1_ASAP7_75t_L g1486 ( 
.A(n_1414),
.Y(n_1486)
);

INVx3_ASAP7_75t_L g1487 ( 
.A(n_1397),
.Y(n_1487)
);

INVx2_ASAP7_75t_L g1488 ( 
.A(n_1449),
.Y(n_1488)
);

INVx1_ASAP7_75t_L g1489 ( 
.A(n_1410),
.Y(n_1489)
);

INVx1_ASAP7_75t_L g1490 ( 
.A(n_1412),
.Y(n_1490)
);

AND2x2_ASAP7_75t_L g1491 ( 
.A(n_1393),
.B(n_1450),
.Y(n_1491)
);

INVx2_ASAP7_75t_L g1492 ( 
.A(n_1449),
.Y(n_1492)
);

INVx1_ASAP7_75t_L g1493 ( 
.A(n_1415),
.Y(n_1493)
);

INVx1_ASAP7_75t_L g1494 ( 
.A(n_1427),
.Y(n_1494)
);

INVx1_ASAP7_75t_L g1495 ( 
.A(n_1440),
.Y(n_1495)
);

INVx3_ASAP7_75t_L g1496 ( 
.A(n_1397),
.Y(n_1496)
);

INVx1_ASAP7_75t_L g1497 ( 
.A(n_1428),
.Y(n_1497)
);

INVx1_ASAP7_75t_L g1498 ( 
.A(n_1445),
.Y(n_1498)
);

INVx1_ASAP7_75t_L g1499 ( 
.A(n_1446),
.Y(n_1499)
);

NAND2xp5_ASAP7_75t_L g1500 ( 
.A(n_1384),
.B(n_1471),
.Y(n_1500)
);

INVx1_ASAP7_75t_L g1501 ( 
.A(n_1442),
.Y(n_1501)
);

OAI21x1_ASAP7_75t_L g1502 ( 
.A1(n_1451),
.A2(n_1453),
.B(n_1430),
.Y(n_1502)
);

OR2x2_ASAP7_75t_L g1503 ( 
.A(n_1392),
.B(n_1474),
.Y(n_1503)
);

HB1xp67_ASAP7_75t_SL g1504 ( 
.A(n_1391),
.Y(n_1504)
);

AND2x2_ASAP7_75t_L g1505 ( 
.A(n_1385),
.B(n_1466),
.Y(n_1505)
);

INVx1_ASAP7_75t_L g1506 ( 
.A(n_1407),
.Y(n_1506)
);

OR2x2_ASAP7_75t_L g1507 ( 
.A(n_1403),
.B(n_1476),
.Y(n_1507)
);

OAI21xp5_ASAP7_75t_L g1508 ( 
.A1(n_1395),
.A2(n_1464),
.B(n_1461),
.Y(n_1508)
);

INVx1_ASAP7_75t_L g1509 ( 
.A(n_1420),
.Y(n_1509)
);

OR2x2_ASAP7_75t_L g1510 ( 
.A(n_1421),
.B(n_1434),
.Y(n_1510)
);

INVx1_ASAP7_75t_L g1511 ( 
.A(n_1439),
.Y(n_1511)
);

AO21x2_ASAP7_75t_L g1512 ( 
.A1(n_1419),
.A2(n_1465),
.B(n_1455),
.Y(n_1512)
);

NAND2xp5_ASAP7_75t_L g1513 ( 
.A(n_1475),
.B(n_1399),
.Y(n_1513)
);

AND2x2_ASAP7_75t_L g1514 ( 
.A(n_1404),
.B(n_1424),
.Y(n_1514)
);

AND2x2_ASAP7_75t_L g1515 ( 
.A(n_1404),
.B(n_1424),
.Y(n_1515)
);

INVx2_ASAP7_75t_SL g1516 ( 
.A(n_1444),
.Y(n_1516)
);

HB1xp67_ASAP7_75t_L g1517 ( 
.A(n_1462),
.Y(n_1517)
);

OR2x2_ASAP7_75t_L g1518 ( 
.A(n_1423),
.B(n_1418),
.Y(n_1518)
);

AO21x2_ASAP7_75t_L g1519 ( 
.A1(n_1455),
.A2(n_1454),
.B(n_1426),
.Y(n_1519)
);

OR2x2_ASAP7_75t_L g1520 ( 
.A(n_1468),
.B(n_1425),
.Y(n_1520)
);

INVx1_ASAP7_75t_L g1521 ( 
.A(n_1436),
.Y(n_1521)
);

NAND2xp5_ASAP7_75t_L g1522 ( 
.A(n_1429),
.B(n_1464),
.Y(n_1522)
);

NOR2xp33_ASAP7_75t_L g1523 ( 
.A(n_1413),
.B(n_1402),
.Y(n_1523)
);

AND2x4_ASAP7_75t_L g1524 ( 
.A(n_1394),
.B(n_1431),
.Y(n_1524)
);

AOI222xp33_ASAP7_75t_L g1525 ( 
.A1(n_1405),
.A2(n_1409),
.B1(n_1470),
.B2(n_1467),
.C1(n_1401),
.C2(n_1389),
.Y(n_1525)
);

AND2x2_ASAP7_75t_L g1526 ( 
.A(n_1406),
.B(n_1472),
.Y(n_1526)
);

AO21x2_ASAP7_75t_L g1527 ( 
.A1(n_1426),
.A2(n_1416),
.B(n_1461),
.Y(n_1527)
);

OR2x2_ASAP7_75t_L g1528 ( 
.A(n_1394),
.B(n_1433),
.Y(n_1528)
);

AND2x2_ASAP7_75t_L g1529 ( 
.A(n_1457),
.B(n_1472),
.Y(n_1529)
);

INVx2_ASAP7_75t_SL g1530 ( 
.A(n_1386),
.Y(n_1530)
);

BUFx2_ASAP7_75t_L g1531 ( 
.A(n_1457),
.Y(n_1531)
);

AO21x2_ASAP7_75t_L g1532 ( 
.A1(n_1416),
.A2(n_1413),
.B(n_1447),
.Y(n_1532)
);

AND2x2_ASAP7_75t_L g1533 ( 
.A(n_1482),
.B(n_1459),
.Y(n_1533)
);

NAND2xp5_ASAP7_75t_SL g1534 ( 
.A(n_1508),
.B(n_1386),
.Y(n_1534)
);

INVx1_ASAP7_75t_L g1535 ( 
.A(n_1495),
.Y(n_1535)
);

OA21x2_ASAP7_75t_L g1536 ( 
.A1(n_1502),
.A2(n_1531),
.B(n_1515),
.Y(n_1536)
);

HB1xp67_ASAP7_75t_L g1537 ( 
.A(n_1481),
.Y(n_1537)
);

AND2x4_ASAP7_75t_L g1538 ( 
.A(n_1484),
.B(n_1473),
.Y(n_1538)
);

AOI22xp33_ASAP7_75t_L g1539 ( 
.A1(n_1525),
.A2(n_1483),
.B1(n_1508),
.B2(n_1522),
.Y(n_1539)
);

INVx2_ASAP7_75t_L g1540 ( 
.A(n_1487),
.Y(n_1540)
);

BUFx3_ASAP7_75t_L g1541 ( 
.A(n_1484),
.Y(n_1541)
);

AND2x2_ASAP7_75t_L g1542 ( 
.A(n_1514),
.B(n_1430),
.Y(n_1542)
);

BUFx2_ASAP7_75t_SL g1543 ( 
.A(n_1524),
.Y(n_1543)
);

HB1xp67_ASAP7_75t_L g1544 ( 
.A(n_1517),
.Y(n_1544)
);

OR2x2_ASAP7_75t_L g1545 ( 
.A(n_1507),
.B(n_1386),
.Y(n_1545)
);

AND2x2_ASAP7_75t_L g1546 ( 
.A(n_1515),
.B(n_1411),
.Y(n_1546)
);

AND2x2_ASAP7_75t_L g1547 ( 
.A(n_1526),
.B(n_1411),
.Y(n_1547)
);

INVx2_ASAP7_75t_L g1548 ( 
.A(n_1496),
.Y(n_1548)
);

HB1xp67_ASAP7_75t_L g1549 ( 
.A(n_1480),
.Y(n_1549)
);

HB1xp67_ASAP7_75t_L g1550 ( 
.A(n_1480),
.Y(n_1550)
);

NAND2xp5_ASAP7_75t_L g1551 ( 
.A(n_1479),
.B(n_1417),
.Y(n_1551)
);

AOI21xp33_ASAP7_75t_L g1552 ( 
.A1(n_1525),
.A2(n_1417),
.B(n_1443),
.Y(n_1552)
);

AND2x4_ASAP7_75t_L g1553 ( 
.A(n_1484),
.B(n_1485),
.Y(n_1553)
);

AND2x2_ASAP7_75t_L g1554 ( 
.A(n_1529),
.B(n_1491),
.Y(n_1554)
);

OAI321xp33_ASAP7_75t_L g1555 ( 
.A1(n_1483),
.A2(n_1469),
.A3(n_1458),
.B1(n_1398),
.B2(n_1437),
.C(n_1435),
.Y(n_1555)
);

AO21x2_ASAP7_75t_L g1556 ( 
.A1(n_1546),
.A2(n_1492),
.B(n_1488),
.Y(n_1556)
);

INVx3_ASAP7_75t_L g1557 ( 
.A(n_1536),
.Y(n_1557)
);

BUFx3_ASAP7_75t_L g1558 ( 
.A(n_1538),
.Y(n_1558)
);

INVx1_ASAP7_75t_L g1559 ( 
.A(n_1535),
.Y(n_1559)
);

AND2x2_ASAP7_75t_L g1560 ( 
.A(n_1554),
.B(n_1491),
.Y(n_1560)
);

BUFx3_ASAP7_75t_L g1561 ( 
.A(n_1538),
.Y(n_1561)
);

INVx2_ASAP7_75t_SL g1562 ( 
.A(n_1541),
.Y(n_1562)
);

AOI222xp33_ASAP7_75t_L g1563 ( 
.A1(n_1539),
.A2(n_1522),
.B1(n_1500),
.B2(n_1523),
.C1(n_1504),
.C2(n_1513),
.Y(n_1563)
);

OAI221xp5_ASAP7_75t_L g1564 ( 
.A1(n_1539),
.A2(n_1523),
.B1(n_1504),
.B2(n_1518),
.C(n_1500),
.Y(n_1564)
);

AO21x2_ASAP7_75t_L g1565 ( 
.A1(n_1546),
.A2(n_1511),
.B(n_1492),
.Y(n_1565)
);

INVxp67_ASAP7_75t_L g1566 ( 
.A(n_1549),
.Y(n_1566)
);

INVx1_ASAP7_75t_L g1567 ( 
.A(n_1535),
.Y(n_1567)
);

OAI221xp5_ASAP7_75t_L g1568 ( 
.A1(n_1552),
.A2(n_1518),
.B1(n_1511),
.B2(n_1513),
.C(n_1521),
.Y(n_1568)
);

AO21x2_ASAP7_75t_L g1569 ( 
.A1(n_1546),
.A2(n_1492),
.B(n_1488),
.Y(n_1569)
);

INVx2_ASAP7_75t_SL g1570 ( 
.A(n_1541),
.Y(n_1570)
);

AOI33xp33_ASAP7_75t_L g1571 ( 
.A1(n_1546),
.A2(n_1521),
.A3(n_1486),
.B1(n_1506),
.B2(n_1490),
.B3(n_1489),
.Y(n_1571)
);

OAI221xp5_ASAP7_75t_L g1572 ( 
.A1(n_1552),
.A2(n_1518),
.B1(n_1506),
.B2(n_1509),
.C(n_1499),
.Y(n_1572)
);

AND2x2_ASAP7_75t_L g1573 ( 
.A(n_1554),
.B(n_1491),
.Y(n_1573)
);

AOI33xp33_ASAP7_75t_L g1574 ( 
.A1(n_1547),
.A2(n_1489),
.A3(n_1490),
.B1(n_1497),
.B2(n_1529),
.B3(n_1501),
.Y(n_1574)
);

OR2x2_ASAP7_75t_L g1575 ( 
.A(n_1537),
.B(n_1507),
.Y(n_1575)
);

NOR2xp67_ASAP7_75t_SL g1576 ( 
.A(n_1543),
.B(n_1473),
.Y(n_1576)
);

OAI22xp5_ASAP7_75t_L g1577 ( 
.A1(n_1551),
.A2(n_1505),
.B1(n_1520),
.B2(n_1503),
.Y(n_1577)
);

OAI221xp5_ASAP7_75t_L g1578 ( 
.A1(n_1551),
.A2(n_1509),
.B1(n_1498),
.B2(n_1499),
.C(n_1510),
.Y(n_1578)
);

INVxp67_ASAP7_75t_L g1579 ( 
.A(n_1549),
.Y(n_1579)
);

NOR2xp33_ASAP7_75t_R g1580 ( 
.A(n_1545),
.B(n_1408),
.Y(n_1580)
);

BUFx2_ASAP7_75t_L g1581 ( 
.A(n_1550),
.Y(n_1581)
);

AOI22xp33_ASAP7_75t_L g1582 ( 
.A1(n_1547),
.A2(n_1532),
.B1(n_1527),
.B2(n_1488),
.Y(n_1582)
);

AO21x2_ASAP7_75t_L g1583 ( 
.A1(n_1547),
.A2(n_1519),
.B(n_1512),
.Y(n_1583)
);

BUFx2_ASAP7_75t_L g1584 ( 
.A(n_1550),
.Y(n_1584)
);

OAI221xp5_ASAP7_75t_L g1585 ( 
.A1(n_1534),
.A2(n_1498),
.B1(n_1510),
.B2(n_1497),
.C(n_1516),
.Y(n_1585)
);

INVx1_ASAP7_75t_L g1586 ( 
.A(n_1535),
.Y(n_1586)
);

AOI221xp5_ASAP7_75t_L g1587 ( 
.A1(n_1547),
.A2(n_1532),
.B1(n_1527),
.B2(n_1494),
.C(n_1493),
.Y(n_1587)
);

OR2x2_ASAP7_75t_L g1588 ( 
.A(n_1537),
.B(n_1503),
.Y(n_1588)
);

OAI21xp5_ASAP7_75t_L g1589 ( 
.A1(n_1555),
.A2(n_1524),
.B(n_1528),
.Y(n_1589)
);

AND2x2_ASAP7_75t_L g1590 ( 
.A(n_1533),
.B(n_1478),
.Y(n_1590)
);

INVx1_ASAP7_75t_SL g1591 ( 
.A(n_1580),
.Y(n_1591)
);

INVx1_ASAP7_75t_L g1592 ( 
.A(n_1559),
.Y(n_1592)
);

NAND2xp5_ASAP7_75t_L g1593 ( 
.A(n_1571),
.B(n_1544),
.Y(n_1593)
);

INVxp67_ASAP7_75t_SL g1594 ( 
.A(n_1557),
.Y(n_1594)
);

INVxp67_ASAP7_75t_L g1595 ( 
.A(n_1572),
.Y(n_1595)
);

INVxp67_ASAP7_75t_L g1596 ( 
.A(n_1572),
.Y(n_1596)
);

INVx2_ASAP7_75t_L g1597 ( 
.A(n_1583),
.Y(n_1597)
);

NAND3xp33_ASAP7_75t_L g1598 ( 
.A(n_1587),
.B(n_1536),
.C(n_1542),
.Y(n_1598)
);

INVx2_ASAP7_75t_SL g1599 ( 
.A(n_1558),
.Y(n_1599)
);

HB1xp67_ASAP7_75t_L g1600 ( 
.A(n_1581),
.Y(n_1600)
);

INVx1_ASAP7_75t_L g1601 ( 
.A(n_1559),
.Y(n_1601)
);

INVx1_ASAP7_75t_L g1602 ( 
.A(n_1567),
.Y(n_1602)
);

OR2x2_ASAP7_75t_L g1603 ( 
.A(n_1588),
.B(n_1544),
.Y(n_1603)
);

INVx2_ASAP7_75t_SL g1604 ( 
.A(n_1557),
.Y(n_1604)
);

INVx2_ASAP7_75t_L g1605 ( 
.A(n_1583),
.Y(n_1605)
);

INVx1_ASAP7_75t_L g1606 ( 
.A(n_1567),
.Y(n_1606)
);

NOR2x1p5_ASAP7_75t_L g1607 ( 
.A(n_1558),
.B(n_1561),
.Y(n_1607)
);

INVx1_ASAP7_75t_L g1608 ( 
.A(n_1586),
.Y(n_1608)
);

INVx2_ASAP7_75t_L g1609 ( 
.A(n_1583),
.Y(n_1609)
);

INVx1_ASAP7_75t_L g1610 ( 
.A(n_1586),
.Y(n_1610)
);

INVx2_ASAP7_75t_L g1611 ( 
.A(n_1583),
.Y(n_1611)
);

INVx2_ASAP7_75t_L g1612 ( 
.A(n_1583),
.Y(n_1612)
);

INVx3_ASAP7_75t_L g1613 ( 
.A(n_1557),
.Y(n_1613)
);

INVx3_ASAP7_75t_L g1614 ( 
.A(n_1557),
.Y(n_1614)
);

AO21x2_ASAP7_75t_L g1615 ( 
.A1(n_1565),
.A2(n_1519),
.B(n_1542),
.Y(n_1615)
);

INVx1_ASAP7_75t_SL g1616 ( 
.A(n_1580),
.Y(n_1616)
);

AND2x4_ASAP7_75t_L g1617 ( 
.A(n_1558),
.B(n_1561),
.Y(n_1617)
);

INVx2_ASAP7_75t_L g1618 ( 
.A(n_1556),
.Y(n_1618)
);

AND2x4_ASAP7_75t_L g1619 ( 
.A(n_1561),
.B(n_1553),
.Y(n_1619)
);

OA21x2_ASAP7_75t_L g1620 ( 
.A1(n_1587),
.A2(n_1540),
.B(n_1548),
.Y(n_1620)
);

NOR2x1_ASAP7_75t_L g1621 ( 
.A(n_1589),
.B(n_1534),
.Y(n_1621)
);

INVx2_ASAP7_75t_L g1622 ( 
.A(n_1556),
.Y(n_1622)
);

INVx2_ASAP7_75t_L g1623 ( 
.A(n_1556),
.Y(n_1623)
);

INVx3_ASAP7_75t_L g1624 ( 
.A(n_1556),
.Y(n_1624)
);

INVx1_ASAP7_75t_L g1625 ( 
.A(n_1588),
.Y(n_1625)
);

INVx2_ASAP7_75t_L g1626 ( 
.A(n_1556),
.Y(n_1626)
);

INVx4_ASAP7_75t_L g1627 ( 
.A(n_1565),
.Y(n_1627)
);

AND2x2_ASAP7_75t_L g1628 ( 
.A(n_1607),
.B(n_1590),
.Y(n_1628)
);

INVx2_ASAP7_75t_L g1629 ( 
.A(n_1627),
.Y(n_1629)
);

NAND2xp5_ASAP7_75t_L g1630 ( 
.A(n_1595),
.B(n_1571),
.Y(n_1630)
);

INVx1_ASAP7_75t_L g1631 ( 
.A(n_1592),
.Y(n_1631)
);

AND2x4_ASAP7_75t_L g1632 ( 
.A(n_1607),
.B(n_1589),
.Y(n_1632)
);

NAND3xp33_ASAP7_75t_SL g1633 ( 
.A(n_1595),
.B(n_1596),
.C(n_1598),
.Y(n_1633)
);

INVx1_ASAP7_75t_L g1634 ( 
.A(n_1592),
.Y(n_1634)
);

AND2x2_ASAP7_75t_L g1635 ( 
.A(n_1607),
.B(n_1590),
.Y(n_1635)
);

INVxp67_ASAP7_75t_SL g1636 ( 
.A(n_1621),
.Y(n_1636)
);

INVx1_ASAP7_75t_L g1637 ( 
.A(n_1592),
.Y(n_1637)
);

INVx2_ASAP7_75t_SL g1638 ( 
.A(n_1617),
.Y(n_1638)
);

AND2x2_ASAP7_75t_L g1639 ( 
.A(n_1617),
.B(n_1590),
.Y(n_1639)
);

INVx1_ASAP7_75t_L g1640 ( 
.A(n_1601),
.Y(n_1640)
);

NAND2xp5_ASAP7_75t_L g1641 ( 
.A(n_1596),
.B(n_1574),
.Y(n_1641)
);

NAND2xp5_ASAP7_75t_L g1642 ( 
.A(n_1621),
.B(n_1574),
.Y(n_1642)
);

INVx3_ASAP7_75t_L g1643 ( 
.A(n_1627),
.Y(n_1643)
);

NOR2xp33_ASAP7_75t_L g1644 ( 
.A(n_1591),
.B(n_1422),
.Y(n_1644)
);

A2O1A1Ixp33_ASAP7_75t_L g1645 ( 
.A1(n_1598),
.A2(n_1564),
.B(n_1568),
.C(n_1582),
.Y(n_1645)
);

OR2x2_ASAP7_75t_L g1646 ( 
.A(n_1593),
.B(n_1603),
.Y(n_1646)
);

INVx1_ASAP7_75t_SL g1647 ( 
.A(n_1591),
.Y(n_1647)
);

INVxp67_ASAP7_75t_L g1648 ( 
.A(n_1616),
.Y(n_1648)
);

AND2x2_ASAP7_75t_L g1649 ( 
.A(n_1617),
.B(n_1560),
.Y(n_1649)
);

OR2x2_ASAP7_75t_L g1650 ( 
.A(n_1593),
.B(n_1575),
.Y(n_1650)
);

OR2x2_ASAP7_75t_L g1651 ( 
.A(n_1603),
.B(n_1625),
.Y(n_1651)
);

NAND2xp5_ASAP7_75t_SL g1652 ( 
.A(n_1616),
.B(n_1577),
.Y(n_1652)
);

NAND2xp5_ASAP7_75t_SL g1653 ( 
.A(n_1617),
.B(n_1577),
.Y(n_1653)
);

AOI31xp33_ASAP7_75t_L g1654 ( 
.A1(n_1599),
.A2(n_1563),
.A3(n_1564),
.B(n_1568),
.Y(n_1654)
);

AND2x2_ASAP7_75t_L g1655 ( 
.A(n_1617),
.B(n_1560),
.Y(n_1655)
);

HB1xp67_ASAP7_75t_L g1656 ( 
.A(n_1600),
.Y(n_1656)
);

INVx1_ASAP7_75t_L g1657 ( 
.A(n_1601),
.Y(n_1657)
);

OR2x2_ASAP7_75t_L g1658 ( 
.A(n_1603),
.B(n_1625),
.Y(n_1658)
);

INVx1_ASAP7_75t_L g1659 ( 
.A(n_1601),
.Y(n_1659)
);

AOI22xp33_ASAP7_75t_L g1660 ( 
.A1(n_1615),
.A2(n_1563),
.B1(n_1582),
.B2(n_1565),
.Y(n_1660)
);

INVx1_ASAP7_75t_L g1661 ( 
.A(n_1602),
.Y(n_1661)
);

OR2x2_ASAP7_75t_L g1662 ( 
.A(n_1625),
.B(n_1575),
.Y(n_1662)
);

NAND2xp33_ASAP7_75t_SL g1663 ( 
.A(n_1599),
.B(n_1576),
.Y(n_1663)
);

INVx1_ASAP7_75t_L g1664 ( 
.A(n_1602),
.Y(n_1664)
);

INVx2_ASAP7_75t_L g1665 ( 
.A(n_1627),
.Y(n_1665)
);

NAND2x1_ASAP7_75t_L g1666 ( 
.A(n_1627),
.B(n_1581),
.Y(n_1666)
);

INVx1_ASAP7_75t_L g1667 ( 
.A(n_1602),
.Y(n_1667)
);

NOR2xp33_ASAP7_75t_SL g1668 ( 
.A(n_1617),
.B(n_1438),
.Y(n_1668)
);

INVx1_ASAP7_75t_L g1669 ( 
.A(n_1606),
.Y(n_1669)
);

AND2x2_ASAP7_75t_L g1670 ( 
.A(n_1599),
.B(n_1560),
.Y(n_1670)
);

NAND2xp5_ASAP7_75t_L g1671 ( 
.A(n_1647),
.B(n_1600),
.Y(n_1671)
);

AOI21xp33_ASAP7_75t_L g1672 ( 
.A1(n_1654),
.A2(n_1615),
.B(n_1627),
.Y(n_1672)
);

AND2x2_ASAP7_75t_L g1673 ( 
.A(n_1632),
.B(n_1619),
.Y(n_1673)
);

OR2x2_ASAP7_75t_L g1674 ( 
.A(n_1646),
.B(n_1575),
.Y(n_1674)
);

INVx1_ASAP7_75t_L g1675 ( 
.A(n_1664),
.Y(n_1675)
);

AOI22xp5_ASAP7_75t_L g1676 ( 
.A1(n_1633),
.A2(n_1615),
.B1(n_1620),
.B2(n_1627),
.Y(n_1676)
);

OR2x2_ASAP7_75t_L g1677 ( 
.A(n_1646),
.B(n_1615),
.Y(n_1677)
);

NAND2xp5_ASAP7_75t_L g1678 ( 
.A(n_1648),
.B(n_1565),
.Y(n_1678)
);

INVx2_ASAP7_75t_L g1679 ( 
.A(n_1643),
.Y(n_1679)
);

AND2x2_ASAP7_75t_L g1680 ( 
.A(n_1632),
.B(n_1619),
.Y(n_1680)
);

INVx1_ASAP7_75t_L g1681 ( 
.A(n_1664),
.Y(n_1681)
);

OR2x2_ASAP7_75t_L g1682 ( 
.A(n_1641),
.B(n_1588),
.Y(n_1682)
);

NAND2xp33_ASAP7_75t_L g1683 ( 
.A(n_1630),
.B(n_1604),
.Y(n_1683)
);

OR2x2_ASAP7_75t_L g1684 ( 
.A(n_1650),
.B(n_1569),
.Y(n_1684)
);

OR2x2_ASAP7_75t_L g1685 ( 
.A(n_1650),
.B(n_1569),
.Y(n_1685)
);

AO22x1_ASAP7_75t_L g1686 ( 
.A1(n_1636),
.A2(n_1594),
.B1(n_1624),
.B2(n_1623),
.Y(n_1686)
);

NOR2xp33_ASAP7_75t_L g1687 ( 
.A(n_1644),
.B(n_1615),
.Y(n_1687)
);

AOI32xp33_ASAP7_75t_L g1688 ( 
.A1(n_1642),
.A2(n_1624),
.A3(n_1594),
.B1(n_1626),
.B2(n_1623),
.Y(n_1688)
);

INVx1_ASAP7_75t_SL g1689 ( 
.A(n_1652),
.Y(n_1689)
);

INVx1_ASAP7_75t_L g1690 ( 
.A(n_1667),
.Y(n_1690)
);

AND2x2_ASAP7_75t_L g1691 ( 
.A(n_1632),
.B(n_1619),
.Y(n_1691)
);

INVx1_ASAP7_75t_L g1692 ( 
.A(n_1667),
.Y(n_1692)
);

NOR2x1p5_ASAP7_75t_SL g1693 ( 
.A(n_1629),
.B(n_1618),
.Y(n_1693)
);

AND2x2_ASAP7_75t_L g1694 ( 
.A(n_1628),
.B(n_1619),
.Y(n_1694)
);

NAND2xp33_ASAP7_75t_L g1695 ( 
.A(n_1645),
.B(n_1604),
.Y(n_1695)
);

AND2x2_ASAP7_75t_L g1696 ( 
.A(n_1628),
.B(n_1619),
.Y(n_1696)
);

INVxp67_ASAP7_75t_L g1697 ( 
.A(n_1656),
.Y(n_1697)
);

INVx2_ASAP7_75t_L g1698 ( 
.A(n_1643),
.Y(n_1698)
);

OR2x2_ASAP7_75t_L g1699 ( 
.A(n_1651),
.B(n_1569),
.Y(n_1699)
);

INVx1_ASAP7_75t_L g1700 ( 
.A(n_1631),
.Y(n_1700)
);

AND2x2_ASAP7_75t_L g1701 ( 
.A(n_1635),
.B(n_1619),
.Y(n_1701)
);

INVx1_ASAP7_75t_L g1702 ( 
.A(n_1634),
.Y(n_1702)
);

NAND2xp5_ASAP7_75t_L g1703 ( 
.A(n_1651),
.B(n_1533),
.Y(n_1703)
);

INVx1_ASAP7_75t_L g1704 ( 
.A(n_1637),
.Y(n_1704)
);

INVx1_ASAP7_75t_L g1705 ( 
.A(n_1640),
.Y(n_1705)
);

AND2x2_ASAP7_75t_L g1706 ( 
.A(n_1635),
.B(n_1573),
.Y(n_1706)
);

NAND2x1p5_ASAP7_75t_L g1707 ( 
.A(n_1689),
.B(n_1576),
.Y(n_1707)
);

OAI21xp5_ASAP7_75t_L g1708 ( 
.A1(n_1695),
.A2(n_1676),
.B(n_1672),
.Y(n_1708)
);

INVx1_ASAP7_75t_SL g1709 ( 
.A(n_1671),
.Y(n_1709)
);

AND2x2_ASAP7_75t_L g1710 ( 
.A(n_1673),
.B(n_1649),
.Y(n_1710)
);

INVx1_ASAP7_75t_SL g1711 ( 
.A(n_1683),
.Y(n_1711)
);

OR2x6_ASAP7_75t_L g1712 ( 
.A(n_1686),
.B(n_1638),
.Y(n_1712)
);

OR2x2_ASAP7_75t_L g1713 ( 
.A(n_1682),
.B(n_1658),
.Y(n_1713)
);

OR2x2_ASAP7_75t_L g1714 ( 
.A(n_1674),
.B(n_1658),
.Y(n_1714)
);

INVxp67_ASAP7_75t_L g1715 ( 
.A(n_1695),
.Y(n_1715)
);

NOR2xp33_ASAP7_75t_L g1716 ( 
.A(n_1697),
.B(n_1668),
.Y(n_1716)
);

INVx1_ASAP7_75t_L g1717 ( 
.A(n_1675),
.Y(n_1717)
);

NAND2xp5_ASAP7_75t_L g1718 ( 
.A(n_1700),
.B(n_1660),
.Y(n_1718)
);

AND2x2_ASAP7_75t_L g1719 ( 
.A(n_1673),
.B(n_1649),
.Y(n_1719)
);

INVx2_ASAP7_75t_L g1720 ( 
.A(n_1677),
.Y(n_1720)
);

NAND2xp33_ASAP7_75t_SL g1721 ( 
.A(n_1680),
.B(n_1666),
.Y(n_1721)
);

INVx1_ASAP7_75t_L g1722 ( 
.A(n_1681),
.Y(n_1722)
);

AND2x2_ASAP7_75t_L g1723 ( 
.A(n_1680),
.B(n_1655),
.Y(n_1723)
);

OR2x2_ASAP7_75t_L g1724 ( 
.A(n_1703),
.B(n_1662),
.Y(n_1724)
);

OAI22xp5_ASAP7_75t_L g1725 ( 
.A1(n_1687),
.A2(n_1653),
.B1(n_1638),
.B2(n_1655),
.Y(n_1725)
);

INVx1_ASAP7_75t_L g1726 ( 
.A(n_1690),
.Y(n_1726)
);

NOR2xp33_ASAP7_75t_L g1727 ( 
.A(n_1683),
.B(n_1663),
.Y(n_1727)
);

INVx1_ASAP7_75t_L g1728 ( 
.A(n_1692),
.Y(n_1728)
);

INVx1_ASAP7_75t_L g1729 ( 
.A(n_1702),
.Y(n_1729)
);

INVx1_ASAP7_75t_L g1730 ( 
.A(n_1704),
.Y(n_1730)
);

INVx1_ASAP7_75t_SL g1731 ( 
.A(n_1691),
.Y(n_1731)
);

INVxp67_ASAP7_75t_SL g1732 ( 
.A(n_1715),
.Y(n_1732)
);

OAI322xp33_ASAP7_75t_L g1733 ( 
.A1(n_1715),
.A2(n_1677),
.A3(n_1687),
.B1(n_1678),
.B2(n_1685),
.C1(n_1684),
.C2(n_1699),
.Y(n_1733)
);

OAI21xp5_ASAP7_75t_L g1734 ( 
.A1(n_1708),
.A2(n_1666),
.B(n_1620),
.Y(n_1734)
);

OAI21xp5_ASAP7_75t_SL g1735 ( 
.A1(n_1711),
.A2(n_1688),
.B(n_1691),
.Y(n_1735)
);

NAND2xp5_ASAP7_75t_L g1736 ( 
.A(n_1731),
.B(n_1706),
.Y(n_1736)
);

OAI322xp33_ASAP7_75t_L g1737 ( 
.A1(n_1718),
.A2(n_1629),
.A3(n_1665),
.B1(n_1643),
.B2(n_1618),
.C1(n_1623),
.C2(n_1622),
.Y(n_1737)
);

OAI21xp33_ASAP7_75t_SL g1738 ( 
.A1(n_1712),
.A2(n_1696),
.B(n_1694),
.Y(n_1738)
);

NAND3xp33_ASAP7_75t_L g1739 ( 
.A(n_1727),
.B(n_1698),
.C(n_1679),
.Y(n_1739)
);

NAND2xp5_ASAP7_75t_L g1740 ( 
.A(n_1709),
.B(n_1706),
.Y(n_1740)
);

OAI221xp5_ASAP7_75t_SL g1741 ( 
.A1(n_1712),
.A2(n_1665),
.B1(n_1624),
.B2(n_1679),
.C(n_1698),
.Y(n_1741)
);

OAI221xp5_ASAP7_75t_SL g1742 ( 
.A1(n_1712),
.A2(n_1624),
.B1(n_1604),
.B2(n_1626),
.C(n_1623),
.Y(n_1742)
);

INVx1_ASAP7_75t_L g1743 ( 
.A(n_1713),
.Y(n_1743)
);

INVx1_ASAP7_75t_L g1744 ( 
.A(n_1714),
.Y(n_1744)
);

AOI21xp5_ASAP7_75t_L g1745 ( 
.A1(n_1727),
.A2(n_1663),
.B(n_1605),
.Y(n_1745)
);

OAI32xp33_ASAP7_75t_L g1746 ( 
.A1(n_1707),
.A2(n_1725),
.A3(n_1721),
.B1(n_1716),
.B2(n_1724),
.Y(n_1746)
);

INVxp67_ASAP7_75t_SL g1747 ( 
.A(n_1716),
.Y(n_1747)
);

INVx2_ASAP7_75t_L g1748 ( 
.A(n_1719),
.Y(n_1748)
);

NAND3xp33_ASAP7_75t_L g1749 ( 
.A(n_1729),
.B(n_1730),
.C(n_1722),
.Y(n_1749)
);

AO22x1_ASAP7_75t_L g1750 ( 
.A1(n_1719),
.A2(n_1624),
.B1(n_1705),
.B2(n_1696),
.Y(n_1750)
);

OAI222xp33_ASAP7_75t_L g1751 ( 
.A1(n_1742),
.A2(n_1707),
.B1(n_1624),
.B2(n_1720),
.C1(n_1618),
.C2(n_1622),
.Y(n_1751)
);

NOR2x1_ASAP7_75t_L g1752 ( 
.A(n_1739),
.B(n_1717),
.Y(n_1752)
);

INVx2_ASAP7_75t_L g1753 ( 
.A(n_1748),
.Y(n_1753)
);

NOR2x1_ASAP7_75t_L g1754 ( 
.A(n_1749),
.B(n_1726),
.Y(n_1754)
);

AOI22xp5_ASAP7_75t_L g1755 ( 
.A1(n_1735),
.A2(n_1734),
.B1(n_1747),
.B2(n_1738),
.Y(n_1755)
);

NOR2xp33_ASAP7_75t_L g1756 ( 
.A(n_1732),
.B(n_1710),
.Y(n_1756)
);

OR2x6_ASAP7_75t_L g1757 ( 
.A(n_1743),
.B(n_1728),
.Y(n_1757)
);

INVx2_ASAP7_75t_L g1758 ( 
.A(n_1744),
.Y(n_1758)
);

OR2x2_ASAP7_75t_L g1759 ( 
.A(n_1740),
.B(n_1662),
.Y(n_1759)
);

INVx1_ASAP7_75t_L g1760 ( 
.A(n_1736),
.Y(n_1760)
);

NOR2x1_ASAP7_75t_L g1761 ( 
.A(n_1737),
.B(n_1723),
.Y(n_1761)
);

OR2x2_ASAP7_75t_L g1762 ( 
.A(n_1757),
.B(n_1759),
.Y(n_1762)
);

AOI221xp5_ASAP7_75t_L g1763 ( 
.A1(n_1751),
.A2(n_1733),
.B1(n_1746),
.B2(n_1742),
.C(n_1741),
.Y(n_1763)
);

OAI21xp33_ASAP7_75t_L g1764 ( 
.A1(n_1756),
.A2(n_1741),
.B(n_1745),
.Y(n_1764)
);

OAI211xp5_ASAP7_75t_L g1765 ( 
.A1(n_1755),
.A2(n_1721),
.B(n_1701),
.C(n_1694),
.Y(n_1765)
);

AOI211xp5_ASAP7_75t_L g1766 ( 
.A1(n_1760),
.A2(n_1750),
.B(n_1720),
.C(n_1555),
.Y(n_1766)
);

AOI222xp33_ASAP7_75t_L g1767 ( 
.A1(n_1761),
.A2(n_1693),
.B1(n_1609),
.B2(n_1605),
.C1(n_1612),
.C2(n_1611),
.Y(n_1767)
);

AOI222xp33_ASAP7_75t_L g1768 ( 
.A1(n_1754),
.A2(n_1612),
.B1(n_1611),
.B2(n_1597),
.C1(n_1609),
.C2(n_1605),
.Y(n_1768)
);

NOR3xp33_ASAP7_75t_L g1769 ( 
.A(n_1758),
.B(n_1605),
.C(n_1597),
.Y(n_1769)
);

O2A1O1Ixp33_ASAP7_75t_L g1770 ( 
.A1(n_1752),
.A2(n_1604),
.B(n_1618),
.C(n_1622),
.Y(n_1770)
);

OAI221xp5_ASAP7_75t_L g1771 ( 
.A1(n_1757),
.A2(n_1620),
.B1(n_1622),
.B2(n_1626),
.C(n_1611),
.Y(n_1771)
);

AND2x2_ASAP7_75t_L g1772 ( 
.A(n_1753),
.B(n_1701),
.Y(n_1772)
);

OAI21xp33_ASAP7_75t_L g1773 ( 
.A1(n_1765),
.A2(n_1669),
.B(n_1661),
.Y(n_1773)
);

AOI22xp5_ASAP7_75t_L g1774 ( 
.A1(n_1767),
.A2(n_1620),
.B1(n_1609),
.B2(n_1612),
.Y(n_1774)
);

OAI221xp5_ASAP7_75t_L g1775 ( 
.A1(n_1763),
.A2(n_1626),
.B1(n_1620),
.B2(n_1612),
.C(n_1597),
.Y(n_1775)
);

OAI211xp5_ASAP7_75t_L g1776 ( 
.A1(n_1764),
.A2(n_1766),
.B(n_1762),
.C(n_1770),
.Y(n_1776)
);

OAI22xp33_ASAP7_75t_L g1777 ( 
.A1(n_1771),
.A2(n_1620),
.B1(n_1597),
.B2(n_1611),
.Y(n_1777)
);

O2A1O1Ixp33_ASAP7_75t_L g1778 ( 
.A1(n_1772),
.A2(n_1609),
.B(n_1614),
.C(n_1613),
.Y(n_1778)
);

NAND3xp33_ASAP7_75t_L g1779 ( 
.A(n_1776),
.B(n_1769),
.C(n_1768),
.Y(n_1779)
);

NAND2xp5_ASAP7_75t_L g1780 ( 
.A(n_1773),
.B(n_1670),
.Y(n_1780)
);

INVx1_ASAP7_75t_L g1781 ( 
.A(n_1775),
.Y(n_1781)
);

OR2x2_ASAP7_75t_L g1782 ( 
.A(n_1777),
.B(n_1670),
.Y(n_1782)
);

NAND2xp5_ASAP7_75t_SL g1783 ( 
.A(n_1778),
.B(n_1657),
.Y(n_1783)
);

AND2x4_ASAP7_75t_L g1784 ( 
.A(n_1774),
.B(n_1639),
.Y(n_1784)
);

OAI21xp5_ASAP7_75t_SL g1785 ( 
.A1(n_1779),
.A2(n_1614),
.B(n_1613),
.Y(n_1785)
);

NOR2xp33_ASAP7_75t_L g1786 ( 
.A(n_1780),
.B(n_1659),
.Y(n_1786)
);

OAI21xp5_ASAP7_75t_SL g1787 ( 
.A1(n_1784),
.A2(n_1614),
.B(n_1613),
.Y(n_1787)
);

NAND4xp75_ASAP7_75t_L g1788 ( 
.A(n_1781),
.B(n_1639),
.C(n_1562),
.D(n_1570),
.Y(n_1788)
);

AOI22xp33_ASAP7_75t_L g1789 ( 
.A1(n_1782),
.A2(n_1569),
.B1(n_1614),
.B2(n_1613),
.Y(n_1789)
);

AND2x4_ASAP7_75t_L g1790 ( 
.A(n_1786),
.B(n_1783),
.Y(n_1790)
);

OAI22xp5_ASAP7_75t_SL g1791 ( 
.A1(n_1789),
.A2(n_1613),
.B1(n_1614),
.B2(n_1585),
.Y(n_1791)
);

NOR3xp33_ASAP7_75t_L g1792 ( 
.A(n_1785),
.B(n_1555),
.C(n_1613),
.Y(n_1792)
);

NOR3xp33_ASAP7_75t_L g1793 ( 
.A(n_1790),
.B(n_1788),
.C(n_1787),
.Y(n_1793)
);

OAI221xp5_ASAP7_75t_L g1794 ( 
.A1(n_1793),
.A2(n_1791),
.B1(n_1792),
.B2(n_1614),
.C(n_1585),
.Y(n_1794)
);

OR5x1_ASAP7_75t_L g1795 ( 
.A(n_1794),
.B(n_1579),
.C(n_1566),
.D(n_1584),
.E(n_1608),
.Y(n_1795)
);

INVx1_ASAP7_75t_L g1796 ( 
.A(n_1794),
.Y(n_1796)
);

INVx2_ASAP7_75t_L g1797 ( 
.A(n_1795),
.Y(n_1797)
);

NOR2xp67_ASAP7_75t_L g1798 ( 
.A(n_1796),
.B(n_1566),
.Y(n_1798)
);

NAND2xp5_ASAP7_75t_SL g1799 ( 
.A(n_1798),
.B(n_1606),
.Y(n_1799)
);

OR2x6_ASAP7_75t_L g1800 ( 
.A(n_1797),
.B(n_1530),
.Y(n_1800)
);

INVx2_ASAP7_75t_SL g1801 ( 
.A(n_1800),
.Y(n_1801)
);

AOI21xp5_ASAP7_75t_L g1802 ( 
.A1(n_1801),
.A2(n_1799),
.B(n_1606),
.Y(n_1802)
);

NAND2xp5_ASAP7_75t_L g1803 ( 
.A(n_1802),
.B(n_1608),
.Y(n_1803)
);

AOI322xp5_ASAP7_75t_L g1804 ( 
.A1(n_1803),
.A2(n_1610),
.A3(n_1608),
.B1(n_1570),
.B2(n_1562),
.C1(n_1579),
.C2(n_1584),
.Y(n_1804)
);

AOI22xp5_ASAP7_75t_L g1805 ( 
.A1(n_1804),
.A2(n_1610),
.B1(n_1569),
.B2(n_1448),
.Y(n_1805)
);

AOI211xp5_ASAP7_75t_L g1806 ( 
.A1(n_1805),
.A2(n_1578),
.B(n_1610),
.C(n_1432),
.Y(n_1806)
);


endmodule