module real_aes_6975_n_103 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_103);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_103;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_357;
wire n_287;
wire n_635;
wire n_503;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_693;
wire n_496;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_178;
wire n_409;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_725;
wire n_455;
wire n_310;
wire n_504;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_733;
wire n_402;
wire n_602;
wire n_552;
wire n_617;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_713;
wire n_598;
wire n_735;
wire n_728;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_397;
wire n_193;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_420;
wire n_336;
wire n_349;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_741;
wire n_283;
wire n_314;
wire n_249;
wire n_623;
wire n_721;
wire n_446;
wire n_221;
wire n_681;
wire n_156;
wire n_456;
wire n_359;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_241;
wire n_175;
wire n_687;
wire n_729;
wire n_646;
wire n_710;
wire n_650;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
AOI222xp33_ASAP7_75t_SL g125 ( .A1(n_0), .A2(n_126), .B1(n_132), .B2(n_721), .C1(n_722), .C2(n_725), .Y(n_125) );
NAND3xp33_ASAP7_75t_SL g109 ( .A(n_1), .B(n_86), .C(n_110), .Y(n_109) );
INVx1_ASAP7_75t_L g123 ( .A(n_1), .Y(n_123) );
INVx1_ASAP7_75t_L g462 ( .A(n_2), .Y(n_462) );
INVx1_ASAP7_75t_L g265 ( .A(n_3), .Y(n_265) );
AOI22xp33_ASAP7_75t_L g537 ( .A1(n_4), .A2(n_38), .B1(n_215), .B2(n_501), .Y(n_537) );
AOI21xp33_ASAP7_75t_L g226 ( .A1(n_5), .A2(n_148), .B(n_227), .Y(n_226) );
NAND2xp5_ASAP7_75t_L g487 ( .A(n_6), .B(n_170), .Y(n_487) );
AND2x6_ASAP7_75t_L g153 ( .A(n_7), .B(n_154), .Y(n_153) );
AOI21xp5_ASAP7_75t_L g146 ( .A1(n_8), .A2(n_147), .B(n_155), .Y(n_146) );
NOR2xp33_ASAP7_75t_L g107 ( .A(n_9), .B(n_39), .Y(n_107) );
NAND2xp5_ASAP7_75t_L g212 ( .A(n_10), .B(n_213), .Y(n_212) );
INVx1_ASAP7_75t_L g232 ( .A(n_11), .Y(n_232) );
INVx1_ASAP7_75t_L g145 ( .A(n_12), .Y(n_145) );
INVx1_ASAP7_75t_L g456 ( .A(n_13), .Y(n_456) );
INVx1_ASAP7_75t_L g165 ( .A(n_14), .Y(n_165) );
NAND2xp5_ASAP7_75t_L g518 ( .A(n_15), .B(n_239), .Y(n_518) );
NAND2xp5_ASAP7_75t_L g489 ( .A(n_16), .B(n_171), .Y(n_489) );
AO32x2_ASAP7_75t_L g535 ( .A1(n_17), .A2(n_170), .A3(n_186), .B1(n_475), .B2(n_536), .Y(n_535) );
NAND2xp5_ASAP7_75t_SL g521 ( .A(n_18), .B(n_215), .Y(n_521) );
NAND2xp5_ASAP7_75t_L g198 ( .A(n_19), .B(n_182), .Y(n_198) );
NAND2xp5_ASAP7_75t_L g465 ( .A(n_20), .B(n_171), .Y(n_465) );
AOI22xp33_ASAP7_75t_L g538 ( .A1(n_21), .A2(n_49), .B1(n_215), .B2(n_501), .Y(n_538) );
NAND2xp5_ASAP7_75t_SL g175 ( .A(n_22), .B(n_148), .Y(n_175) );
AOI22xp33_ASAP7_75t_SL g502 ( .A1(n_23), .A2(n_77), .B1(n_215), .B2(n_239), .Y(n_502) );
NAND2xp5_ASAP7_75t_SL g511 ( .A(n_24), .B(n_215), .Y(n_511) );
NAND2xp5_ASAP7_75t_L g255 ( .A(n_25), .B(n_225), .Y(n_255) );
A2O1A1Ixp33_ASAP7_75t_L g161 ( .A1(n_26), .A2(n_162), .B(n_164), .C(n_166), .Y(n_161) );
AOI22xp33_ASAP7_75t_L g103 ( .A1(n_27), .A2(n_104), .B1(n_113), .B2(n_741), .Y(n_103) );
BUFx6f_ASAP7_75t_L g152 ( .A(n_28), .Y(n_152) );
NAND2xp5_ASAP7_75t_L g476 ( .A(n_29), .B(n_141), .Y(n_476) );
NAND2xp5_ASAP7_75t_L g266 ( .A(n_30), .B(n_197), .Y(n_266) );
OAI22xp5_ASAP7_75t_L g127 ( .A1(n_31), .A2(n_101), .B1(n_128), .B2(n_129), .Y(n_127) );
INVx1_ASAP7_75t_L g129 ( .A(n_31), .Y(n_129) );
INVx1_ASAP7_75t_L g244 ( .A(n_32), .Y(n_244) );
NAND2xp5_ASAP7_75t_L g513 ( .A(n_33), .B(n_141), .Y(n_513) );
INVx2_ASAP7_75t_L g151 ( .A(n_34), .Y(n_151) );
NAND2xp5_ASAP7_75t_SL g470 ( .A(n_35), .B(n_215), .Y(n_470) );
NAND2xp5_ASAP7_75t_L g523 ( .A(n_36), .B(n_141), .Y(n_523) );
A2O1A1Ixp33_ASAP7_75t_L g176 ( .A1(n_37), .A2(n_153), .B(n_158), .C(n_177), .Y(n_176) );
INVx1_ASAP7_75t_L g242 ( .A(n_40), .Y(n_242) );
NAND2xp5_ASAP7_75t_SL g196 ( .A(n_41), .B(n_197), .Y(n_196) );
NAND2xp5_ASAP7_75t_SL g482 ( .A(n_42), .B(n_215), .Y(n_482) );
AOI22xp33_ASAP7_75t_L g500 ( .A1(n_43), .A2(n_87), .B1(n_167), .B2(n_501), .Y(n_500) );
NAND2xp5_ASAP7_75t_SL g485 ( .A(n_44), .B(n_215), .Y(n_485) );
NAND2xp5_ASAP7_75t_L g457 ( .A(n_45), .B(n_215), .Y(n_457) );
CKINVDCx16_ASAP7_75t_R g245 ( .A(n_46), .Y(n_245) );
NAND2xp5_ASAP7_75t_L g486 ( .A(n_47), .B(n_461), .Y(n_486) );
NAND2xp5_ASAP7_75t_L g216 ( .A(n_48), .B(n_148), .Y(n_216) );
AOI22xp33_ASAP7_75t_SL g493 ( .A1(n_50), .A2(n_60), .B1(n_215), .B2(n_239), .Y(n_493) );
OAI22xp5_ASAP7_75t_SL g733 ( .A1(n_51), .A2(n_734), .B1(n_737), .B2(n_738), .Y(n_733) );
CKINVDCx20_ASAP7_75t_R g737 ( .A(n_51), .Y(n_737) );
AOI22xp5_ASAP7_75t_L g238 ( .A1(n_52), .A2(n_158), .B1(n_239), .B2(n_241), .Y(n_238) );
CKINVDCx20_ASAP7_75t_R g188 ( .A(n_53), .Y(n_188) );
NAND2xp5_ASAP7_75t_SL g474 ( .A(n_54), .B(n_215), .Y(n_474) );
CKINVDCx16_ASAP7_75t_R g262 ( .A(n_55), .Y(n_262) );
NAND2xp5_ASAP7_75t_SL g517 ( .A(n_56), .B(n_215), .Y(n_517) );
A2O1A1Ixp33_ASAP7_75t_L g229 ( .A1(n_57), .A2(n_230), .B(n_231), .C(n_233), .Y(n_229) );
CKINVDCx20_ASAP7_75t_R g201 ( .A(n_58), .Y(n_201) );
INVx1_ASAP7_75t_L g228 ( .A(n_59), .Y(n_228) );
INVx1_ASAP7_75t_L g154 ( .A(n_61), .Y(n_154) );
OAI22xp5_ASAP7_75t_SL g126 ( .A1(n_62), .A2(n_127), .B1(n_130), .B2(n_131), .Y(n_126) );
CKINVDCx20_ASAP7_75t_R g131 ( .A(n_62), .Y(n_131) );
NAND2xp5_ASAP7_75t_L g463 ( .A(n_63), .B(n_215), .Y(n_463) );
INVx1_ASAP7_75t_L g144 ( .A(n_64), .Y(n_144) );
OAI22xp5_ASAP7_75t_SL g734 ( .A1(n_65), .A2(n_76), .B1(n_735), .B2(n_736), .Y(n_734) );
CKINVDCx20_ASAP7_75t_R g735 ( .A(n_65), .Y(n_735) );
CKINVDCx20_ASAP7_75t_R g117 ( .A(n_66), .Y(n_117) );
AO32x2_ASAP7_75t_L g498 ( .A1(n_67), .A2(n_170), .A3(n_207), .B1(n_475), .B2(n_499), .Y(n_498) );
INVx1_ASAP7_75t_L g473 ( .A(n_68), .Y(n_473) );
INVx1_ASAP7_75t_L g508 ( .A(n_69), .Y(n_508) );
A2O1A1Ixp33_ASAP7_75t_SL g252 ( .A1(n_70), .A2(n_182), .B(n_233), .C(n_253), .Y(n_252) );
INVxp67_ASAP7_75t_L g254 ( .A(n_71), .Y(n_254) );
NAND2xp5_ASAP7_75t_SL g509 ( .A(n_72), .B(n_239), .Y(n_509) );
INVx1_ASAP7_75t_L g112 ( .A(n_73), .Y(n_112) );
CKINVDCx20_ASAP7_75t_R g247 ( .A(n_74), .Y(n_247) );
INVx1_ASAP7_75t_L g192 ( .A(n_75), .Y(n_192) );
CKINVDCx20_ASAP7_75t_R g736 ( .A(n_76), .Y(n_736) );
A2O1A1Ixp33_ASAP7_75t_L g194 ( .A1(n_78), .A2(n_153), .B(n_158), .C(n_195), .Y(n_194) );
NAND2xp5_ASAP7_75t_L g522 ( .A(n_79), .B(n_501), .Y(n_522) );
NAND2xp5_ASAP7_75t_SL g512 ( .A(n_80), .B(n_239), .Y(n_512) );
NAND2xp5_ASAP7_75t_SL g178 ( .A(n_81), .B(n_179), .Y(n_178) );
INVx2_ASAP7_75t_L g142 ( .A(n_82), .Y(n_142) );
NAND2xp5_ASAP7_75t_L g181 ( .A(n_83), .B(n_182), .Y(n_181) );
NAND2xp5_ASAP7_75t_L g483 ( .A(n_84), .B(n_239), .Y(n_483) );
A2O1A1Ixp33_ASAP7_75t_L g263 ( .A1(n_85), .A2(n_153), .B(n_158), .C(n_264), .Y(n_263) );
OR2x2_ASAP7_75t_L g120 ( .A(n_86), .B(n_121), .Y(n_120) );
OR2x2_ASAP7_75t_L g133 ( .A(n_86), .B(n_122), .Y(n_133) );
INVx2_ASAP7_75t_L g445 ( .A(n_86), .Y(n_445) );
AOI22xp33_ASAP7_75t_L g492 ( .A1(n_88), .A2(n_102), .B1(n_239), .B2(n_240), .Y(n_492) );
NAND2xp5_ASAP7_75t_L g234 ( .A(n_89), .B(n_141), .Y(n_234) );
CKINVDCx20_ASAP7_75t_R g269 ( .A(n_90), .Y(n_269) );
A2O1A1Ixp33_ASAP7_75t_L g209 ( .A1(n_91), .A2(n_153), .B(n_158), .C(n_210), .Y(n_209) );
CKINVDCx20_ASAP7_75t_R g218 ( .A(n_92), .Y(n_218) );
INVx1_ASAP7_75t_L g251 ( .A(n_93), .Y(n_251) );
CKINVDCx16_ASAP7_75t_R g156 ( .A(n_94), .Y(n_156) );
CKINVDCx20_ASAP7_75t_R g124 ( .A(n_95), .Y(n_124) );
NAND2xp5_ASAP7_75t_SL g211 ( .A(n_96), .B(n_179), .Y(n_211) );
NAND2xp5_ASAP7_75t_L g471 ( .A(n_97), .B(n_239), .Y(n_471) );
NAND2xp5_ASAP7_75t_L g169 ( .A(n_98), .B(n_170), .Y(n_169) );
NAND2xp5_ASAP7_75t_L g111 ( .A(n_99), .B(n_112), .Y(n_111) );
AOI21xp5_ASAP7_75t_L g249 ( .A1(n_100), .A2(n_148), .B(n_250), .Y(n_249) );
CKINVDCx20_ASAP7_75t_R g128 ( .A(n_101), .Y(n_128) );
INVx1_ASAP7_75t_L g104 ( .A(n_105), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_106), .Y(n_105) );
CKINVDCx12_ASAP7_75t_R g743 ( .A(n_106), .Y(n_743) );
AND2x2_ASAP7_75t_L g106 ( .A(n_107), .B(n_108), .Y(n_106) );
AND2x2_ASAP7_75t_L g122 ( .A(n_107), .B(n_123), .Y(n_122) );
INVx1_ASAP7_75t_L g108 ( .A(n_109), .Y(n_108) );
INVx1_ASAP7_75t_SL g110 ( .A(n_111), .Y(n_110) );
AOI22x1_ASAP7_75t_L g113 ( .A1(n_114), .A2(n_125), .B1(n_728), .B2(n_730), .Y(n_113) );
NOR2xp33_ASAP7_75t_L g114 ( .A(n_115), .B(n_118), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_116), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
INVx2_ASAP7_75t_L g729 ( .A(n_117), .Y(n_729) );
AOI21xp5_ASAP7_75t_L g730 ( .A1(n_118), .A2(n_731), .B(n_739), .Y(n_730) );
NOR2xp33_ASAP7_75t_SL g118 ( .A(n_119), .B(n_124), .Y(n_118) );
HB1xp67_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
INVx1_ASAP7_75t_SL g740 ( .A(n_120), .Y(n_740) );
NOR2x2_ASAP7_75t_L g727 ( .A(n_121), .B(n_445), .Y(n_727) );
INVx2_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
OR2x2_ASAP7_75t_L g444 ( .A(n_122), .B(n_445), .Y(n_444) );
INVx1_ASAP7_75t_L g721 ( .A(n_126), .Y(n_721) );
INVx1_ASAP7_75t_L g130 ( .A(n_127), .Y(n_130) );
OAI22xp5_ASAP7_75t_L g132 ( .A1(n_133), .A2(n_134), .B1(n_442), .B2(n_446), .Y(n_132) );
OAI22xp5_ASAP7_75t_SL g722 ( .A1(n_133), .A2(n_444), .B1(n_723), .B2(n_724), .Y(n_722) );
INVx2_ASAP7_75t_SL g723 ( .A(n_134), .Y(n_723) );
OAI22xp5_ASAP7_75t_SL g731 ( .A1(n_134), .A2(n_723), .B1(n_732), .B2(n_733), .Y(n_731) );
OR4x2_ASAP7_75t_L g134 ( .A(n_135), .B(n_338), .C(n_397), .D(n_424), .Y(n_134) );
NAND3xp33_ASAP7_75t_SL g135 ( .A(n_136), .B(n_280), .C(n_305), .Y(n_135) );
O2A1O1Ixp33_ASAP7_75t_L g136 ( .A1(n_137), .A2(n_203), .B(n_223), .C(n_256), .Y(n_136) );
AOI211xp5_ASAP7_75t_SL g428 ( .A1(n_137), .A2(n_429), .B(n_431), .C(n_434), .Y(n_428) );
AND2x2_ASAP7_75t_L g137 ( .A(n_138), .B(n_172), .Y(n_137) );
INVx1_ASAP7_75t_L g303 ( .A(n_138), .Y(n_303) );
INVx1_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
OR2x2_ASAP7_75t_L g278 ( .A(n_139), .B(n_279), .Y(n_278) );
INVx2_ASAP7_75t_L g310 ( .A(n_139), .Y(n_310) );
AND2x2_ASAP7_75t_L g365 ( .A(n_139), .B(n_334), .Y(n_365) );
NAND2xp5_ASAP7_75t_L g388 ( .A(n_139), .B(n_221), .Y(n_388) );
NAND2xp5_ASAP7_75t_L g423 ( .A(n_139), .B(n_222), .Y(n_423) );
INVx2_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
INVx1_ASAP7_75t_L g284 ( .A(n_140), .Y(n_284) );
AND2x2_ASAP7_75t_L g327 ( .A(n_140), .B(n_190), .Y(n_327) );
AND2x2_ASAP7_75t_L g345 ( .A(n_140), .B(n_222), .Y(n_345) );
OA21x2_ASAP7_75t_L g140 ( .A1(n_141), .A2(n_146), .B(n_169), .Y(n_140) );
INVx1_ASAP7_75t_L g202 ( .A(n_141), .Y(n_202) );
INVx2_ASAP7_75t_L g207 ( .A(n_141), .Y(n_207) );
OA21x2_ASAP7_75t_L g505 ( .A1(n_141), .A2(n_506), .B(n_513), .Y(n_505) );
OA21x2_ASAP7_75t_L g514 ( .A1(n_141), .A2(n_515), .B(n_523), .Y(n_514) );
AND2x2_ASAP7_75t_SL g141 ( .A(n_142), .B(n_143), .Y(n_141) );
AND2x2_ASAP7_75t_L g171 ( .A(n_142), .B(n_143), .Y(n_171) );
NAND2xp5_ASAP7_75t_L g143 ( .A(n_144), .B(n_145), .Y(n_143) );
BUFx2_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
AND2x4_ASAP7_75t_L g148 ( .A(n_149), .B(n_153), .Y(n_148) );
NAND2x1p5_ASAP7_75t_L g193 ( .A(n_149), .B(n_153), .Y(n_193) );
AND2x2_ASAP7_75t_L g149 ( .A(n_150), .B(n_152), .Y(n_149) );
INVx1_ASAP7_75t_L g461 ( .A(n_150), .Y(n_461) );
INVx1_ASAP7_75t_L g150 ( .A(n_151), .Y(n_150) );
INVx2_ASAP7_75t_L g159 ( .A(n_151), .Y(n_159) );
INVx1_ASAP7_75t_L g240 ( .A(n_151), .Y(n_240) );
INVx1_ASAP7_75t_L g160 ( .A(n_152), .Y(n_160) );
BUFx6f_ASAP7_75t_L g163 ( .A(n_152), .Y(n_163) );
INVx3_ASAP7_75t_L g180 ( .A(n_152), .Y(n_180) );
INVx1_ASAP7_75t_L g182 ( .A(n_152), .Y(n_182) );
BUFx6f_ASAP7_75t_L g197 ( .A(n_152), .Y(n_197) );
INVx4_ASAP7_75t_SL g168 ( .A(n_153), .Y(n_168) );
OAI21xp5_ASAP7_75t_L g454 ( .A1(n_153), .A2(n_455), .B(n_459), .Y(n_454) );
BUFx3_ASAP7_75t_L g475 ( .A(n_153), .Y(n_475) );
OAI21xp5_ASAP7_75t_L g480 ( .A1(n_153), .A2(n_481), .B(n_484), .Y(n_480) );
OAI21xp5_ASAP7_75t_L g506 ( .A1(n_153), .A2(n_507), .B(n_510), .Y(n_506) );
OAI21xp5_ASAP7_75t_L g515 ( .A1(n_153), .A2(n_516), .B(n_520), .Y(n_515) );
O2A1O1Ixp33_ASAP7_75t_L g155 ( .A1(n_156), .A2(n_157), .B(n_161), .C(n_168), .Y(n_155) );
O2A1O1Ixp33_ASAP7_75t_L g227 ( .A1(n_157), .A2(n_168), .B(n_228), .C(n_229), .Y(n_227) );
O2A1O1Ixp33_ASAP7_75t_L g250 ( .A1(n_157), .A2(n_168), .B(n_251), .C(n_252), .Y(n_250) );
INVx5_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
AND2x6_ASAP7_75t_L g158 ( .A(n_159), .B(n_160), .Y(n_158) );
BUFx3_ASAP7_75t_L g167 ( .A(n_159), .Y(n_167) );
BUFx6f_ASAP7_75t_L g215 ( .A(n_159), .Y(n_215) );
INVx1_ASAP7_75t_L g501 ( .A(n_159), .Y(n_501) );
NOR2xp33_ASAP7_75t_L g164 ( .A(n_162), .B(n_165), .Y(n_164) );
INVx1_ASAP7_75t_L g458 ( .A(n_162), .Y(n_458) );
AOI21xp5_ASAP7_75t_L g510 ( .A1(n_162), .A2(n_511), .B(n_512), .Y(n_510) );
INVx4_ASAP7_75t_L g162 ( .A(n_163), .Y(n_162) );
OAI22xp5_ASAP7_75t_SL g241 ( .A1(n_163), .A2(n_242), .B1(n_243), .B2(n_244), .Y(n_241) );
INVx2_ASAP7_75t_L g243 ( .A(n_163), .Y(n_243) );
INVx1_ASAP7_75t_L g166 ( .A(n_167), .Y(n_166) );
INVx2_ASAP7_75t_L g184 ( .A(n_167), .Y(n_184) );
OAI22xp33_ASAP7_75t_L g237 ( .A1(n_168), .A2(n_193), .B1(n_238), .B2(n_245), .Y(n_237) );
INVx4_ASAP7_75t_L g189 ( .A(n_170), .Y(n_189) );
OA21x2_ASAP7_75t_L g248 ( .A1(n_170), .A2(n_249), .B(n_255), .Y(n_248) );
OA21x2_ASAP7_75t_L g479 ( .A1(n_170), .A2(n_480), .B(n_487), .Y(n_479) );
BUFx6f_ASAP7_75t_L g170 ( .A(n_171), .Y(n_170) );
INVx1_ASAP7_75t_L g186 ( .A(n_171), .Y(n_186) );
INVx4_ASAP7_75t_L g277 ( .A(n_172), .Y(n_277) );
OAI21xp5_ASAP7_75t_L g332 ( .A1(n_172), .A2(n_333), .B(n_335), .Y(n_332) );
AND2x2_ASAP7_75t_L g413 ( .A(n_172), .B(n_414), .Y(n_413) );
AND2x2_ASAP7_75t_L g172 ( .A(n_173), .B(n_190), .Y(n_172) );
INVx1_ASAP7_75t_L g220 ( .A(n_173), .Y(n_220) );
AND2x2_ASAP7_75t_L g282 ( .A(n_173), .B(n_222), .Y(n_282) );
OR2x2_ASAP7_75t_L g311 ( .A(n_173), .B(n_312), .Y(n_311) );
INVx2_ASAP7_75t_L g325 ( .A(n_173), .Y(n_325) );
INVx3_ASAP7_75t_L g334 ( .A(n_173), .Y(n_334) );
AND2x2_ASAP7_75t_L g344 ( .A(n_173), .B(n_345), .Y(n_344) );
AND2x2_ASAP7_75t_L g377 ( .A(n_173), .B(n_283), .Y(n_377) );
AND2x2_ASAP7_75t_L g401 ( .A(n_173), .B(n_357), .Y(n_401) );
OR2x6_ASAP7_75t_L g173 ( .A(n_174), .B(n_187), .Y(n_173) );
AOI21xp5_ASAP7_75t_SL g174 ( .A1(n_175), .A2(n_176), .B(n_185), .Y(n_174) );
AOI21xp5_ASAP7_75t_L g177 ( .A1(n_178), .A2(n_181), .B(n_183), .Y(n_177) );
O2A1O1Ixp33_ASAP7_75t_L g264 ( .A1(n_179), .A2(n_265), .B(n_266), .C(n_267), .Y(n_264) );
INVx2_ASAP7_75t_L g464 ( .A(n_179), .Y(n_464) );
AOI21xp5_ASAP7_75t_L g469 ( .A1(n_179), .A2(n_470), .B(n_471), .Y(n_469) );
AOI21xp5_ASAP7_75t_L g481 ( .A1(n_179), .A2(n_482), .B(n_483), .Y(n_481) );
O2A1O1Ixp5_ASAP7_75t_SL g507 ( .A1(n_179), .A2(n_233), .B(n_508), .C(n_509), .Y(n_507) );
INVx5_ASAP7_75t_L g179 ( .A(n_180), .Y(n_179) );
NOR2xp33_ASAP7_75t_L g231 ( .A(n_180), .B(n_232), .Y(n_231) );
NOR2xp33_ASAP7_75t_L g253 ( .A(n_180), .B(n_254), .Y(n_253) );
OAI22xp5_ASAP7_75t_SL g499 ( .A1(n_180), .A2(n_197), .B1(n_500), .B2(n_502), .Y(n_499) );
INVx1_ASAP7_75t_L g519 ( .A(n_182), .Y(n_519) );
AOI21xp5_ASAP7_75t_L g195 ( .A1(n_183), .A2(n_196), .B(n_198), .Y(n_195) );
INVx2_ASAP7_75t_L g183 ( .A(n_184), .Y(n_183) );
INVx1_ASAP7_75t_L g199 ( .A(n_185), .Y(n_199) );
OA21x2_ASAP7_75t_L g453 ( .A1(n_185), .A2(n_454), .B(n_465), .Y(n_453) );
OA21x2_ASAP7_75t_L g467 ( .A1(n_185), .A2(n_468), .B(n_476), .Y(n_467) );
INVx2_ASAP7_75t_L g185 ( .A(n_186), .Y(n_185) );
AO21x2_ASAP7_75t_L g236 ( .A1(n_186), .A2(n_237), .B(n_246), .Y(n_236) );
NOR2xp33_ASAP7_75t_L g246 ( .A(n_186), .B(n_247), .Y(n_246) );
AO21x2_ASAP7_75t_L g260 ( .A1(n_186), .A2(n_261), .B(n_268), .Y(n_260) );
NOR2xp33_ASAP7_75t_SL g187 ( .A(n_188), .B(n_189), .Y(n_187) );
INVx3_ASAP7_75t_L g225 ( .A(n_189), .Y(n_225) );
NAND3xp33_ASAP7_75t_L g490 ( .A(n_189), .B(n_475), .C(n_491), .Y(n_490) );
AO21x1_ASAP7_75t_L g569 ( .A1(n_189), .A2(n_491), .B(n_570), .Y(n_569) );
INVx2_ASAP7_75t_L g222 ( .A(n_190), .Y(n_222) );
AND2x2_ASAP7_75t_L g437 ( .A(n_190), .B(n_279), .Y(n_437) );
AO21x2_ASAP7_75t_L g190 ( .A1(n_191), .A2(n_199), .B(n_200), .Y(n_190) );
OAI21xp5_ASAP7_75t_L g191 ( .A1(n_192), .A2(n_193), .B(n_194), .Y(n_191) );
OAI21xp5_ASAP7_75t_L g261 ( .A1(n_193), .A2(n_262), .B(n_263), .Y(n_261) );
INVx4_ASAP7_75t_L g213 ( .A(n_197), .Y(n_213) );
INVx2_ASAP7_75t_L g230 ( .A(n_197), .Y(n_230) );
OAI22xp5_ASAP7_75t_L g491 ( .A1(n_197), .A2(n_464), .B1(n_492), .B2(n_493), .Y(n_491) );
OAI22xp5_ASAP7_75t_L g536 ( .A1(n_197), .A2(n_464), .B1(n_537), .B2(n_538), .Y(n_536) );
NOR2xp33_ASAP7_75t_L g200 ( .A(n_201), .B(n_202), .Y(n_200) );
NOR2xp33_ASAP7_75t_L g217 ( .A(n_202), .B(n_218), .Y(n_217) );
NOR2xp33_ASAP7_75t_L g268 ( .A(n_202), .B(n_269), .Y(n_268) );
AND2x2_ASAP7_75t_L g203 ( .A(n_204), .B(n_219), .Y(n_203) );
INVx1_ASAP7_75t_L g204 ( .A(n_205), .Y(n_204) );
NOR2xp33_ASAP7_75t_L g333 ( .A(n_205), .B(n_334), .Y(n_333) );
AND2x2_ASAP7_75t_L g357 ( .A(n_205), .B(n_345), .Y(n_357) );
NAND2xp5_ASAP7_75t_L g419 ( .A(n_205), .B(n_334), .Y(n_419) );
INVx1_ASAP7_75t_L g205 ( .A(n_206), .Y(n_205) );
INVx2_ASAP7_75t_L g279 ( .A(n_206), .Y(n_279) );
AND2x2_ASAP7_75t_L g283 ( .A(n_206), .B(n_284), .Y(n_283) );
AND2x2_ASAP7_75t_L g324 ( .A(n_206), .B(n_325), .Y(n_324) );
AO21x2_ASAP7_75t_L g206 ( .A1(n_207), .A2(n_208), .B(n_217), .Y(n_206) );
NAND2xp5_ASAP7_75t_L g208 ( .A(n_209), .B(n_216), .Y(n_208) );
AOI21xp5_ASAP7_75t_L g210 ( .A1(n_211), .A2(n_212), .B(n_214), .Y(n_210) );
HB1xp67_ASAP7_75t_L g214 ( .A(n_215), .Y(n_214) );
INVx3_ASAP7_75t_L g233 ( .A(n_215), .Y(n_233) );
NAND2xp5_ASAP7_75t_L g342 ( .A(n_219), .B(n_320), .Y(n_342) );
INVx1_ASAP7_75t_L g381 ( .A(n_219), .Y(n_381) );
NAND2xp5_ASAP7_75t_L g425 ( .A(n_219), .B(n_308), .Y(n_425) );
AND2x2_ASAP7_75t_L g219 ( .A(n_220), .B(n_221), .Y(n_219) );
AND2x2_ASAP7_75t_L g288 ( .A(n_220), .B(n_283), .Y(n_288) );
INVx2_ASAP7_75t_L g221 ( .A(n_222), .Y(n_221) );
NAND2xp5_ASAP7_75t_L g312 ( .A(n_222), .B(n_279), .Y(n_312) );
INVx1_ASAP7_75t_L g391 ( .A(n_222), .Y(n_391) );
AOI322xp5_ASAP7_75t_L g415 ( .A1(n_223), .A2(n_330), .A3(n_390), .B1(n_416), .B2(n_418), .C1(n_420), .C2(n_422), .Y(n_415) );
AND2x2_ASAP7_75t_SL g223 ( .A(n_224), .B(n_235), .Y(n_223) );
AND2x2_ASAP7_75t_L g270 ( .A(n_224), .B(n_248), .Y(n_270) );
INVx1_ASAP7_75t_SL g273 ( .A(n_224), .Y(n_273) );
AND2x2_ASAP7_75t_L g275 ( .A(n_224), .B(n_236), .Y(n_275) );
NAND2xp5_ASAP7_75t_L g298 ( .A(n_224), .B(n_292), .Y(n_298) );
INVx2_ASAP7_75t_L g317 ( .A(n_224), .Y(n_317) );
AND2x2_ASAP7_75t_L g330 ( .A(n_224), .B(n_331), .Y(n_330) );
OR2x2_ASAP7_75t_L g368 ( .A(n_224), .B(n_292), .Y(n_368) );
BUFx2_ASAP7_75t_L g385 ( .A(n_224), .Y(n_385) );
AND2x2_ASAP7_75t_L g399 ( .A(n_224), .B(n_259), .Y(n_399) );
OA21x2_ASAP7_75t_L g224 ( .A1(n_225), .A2(n_226), .B(n_234), .Y(n_224) );
O2A1O1Ixp5_ASAP7_75t_L g472 ( .A1(n_230), .A2(n_460), .B(n_473), .C(n_474), .Y(n_472) );
AOI21xp5_ASAP7_75t_L g520 ( .A1(n_230), .A2(n_521), .B(n_522), .Y(n_520) );
NAND2xp5_ASAP7_75t_L g314 ( .A(n_235), .B(n_287), .Y(n_314) );
AND2x2_ASAP7_75t_L g441 ( .A(n_235), .B(n_317), .Y(n_441) );
AND2x2_ASAP7_75t_L g235 ( .A(n_236), .B(n_248), .Y(n_235) );
OR2x2_ASAP7_75t_L g286 ( .A(n_236), .B(n_287), .Y(n_286) );
INVx3_ASAP7_75t_L g292 ( .A(n_236), .Y(n_292) );
AND2x2_ASAP7_75t_L g337 ( .A(n_236), .B(n_260), .Y(n_337) );
NOR2xp33_ASAP7_75t_L g384 ( .A(n_236), .B(n_385), .Y(n_384) );
HB1xp67_ASAP7_75t_L g421 ( .A(n_236), .Y(n_421) );
INVx2_ASAP7_75t_L g267 ( .A(n_239), .Y(n_267) );
INVx3_ASAP7_75t_L g239 ( .A(n_240), .Y(n_239) );
AND2x2_ASAP7_75t_L g272 ( .A(n_248), .B(n_273), .Y(n_272) );
INVx1_ASAP7_75t_L g294 ( .A(n_248), .Y(n_294) );
BUFx2_ASAP7_75t_L g300 ( .A(n_248), .Y(n_300) );
AND2x2_ASAP7_75t_L g319 ( .A(n_248), .B(n_292), .Y(n_319) );
INVx3_ASAP7_75t_L g331 ( .A(n_248), .Y(n_331) );
OR2x2_ASAP7_75t_L g341 ( .A(n_248), .B(n_292), .Y(n_341) );
AOI31xp33_ASAP7_75t_SL g256 ( .A1(n_257), .A2(n_271), .A3(n_274), .B(n_276), .Y(n_256) );
NAND2xp5_ASAP7_75t_L g257 ( .A(n_258), .B(n_270), .Y(n_257) );
NAND2xp5_ASAP7_75t_L g304 ( .A(n_258), .B(n_293), .Y(n_304) );
OR2x2_ASAP7_75t_L g328 ( .A(n_258), .B(n_298), .Y(n_328) );
INVx1_ASAP7_75t_SL g258 ( .A(n_259), .Y(n_258) );
NAND2xp5_ASAP7_75t_L g271 ( .A(n_259), .B(n_272), .Y(n_271) );
OR2x2_ASAP7_75t_L g349 ( .A(n_259), .B(n_341), .Y(n_349) );
NOR2xp33_ASAP7_75t_L g359 ( .A(n_259), .B(n_331), .Y(n_359) );
AND2x2_ASAP7_75t_L g366 ( .A(n_259), .B(n_367), .Y(n_366) );
NAND2x1_ASAP7_75t_L g394 ( .A(n_259), .B(n_330), .Y(n_394) );
NOR2xp33_ASAP7_75t_L g395 ( .A(n_259), .B(n_385), .Y(n_395) );
AND2x2_ASAP7_75t_L g407 ( .A(n_259), .B(n_292), .Y(n_407) );
INVx3_ASAP7_75t_L g259 ( .A(n_260), .Y(n_259) );
INVx3_ASAP7_75t_L g287 ( .A(n_260), .Y(n_287) );
O2A1O1Ixp33_ASAP7_75t_L g455 ( .A1(n_267), .A2(n_456), .B(n_457), .C(n_458), .Y(n_455) );
INVx1_ASAP7_75t_L g353 ( .A(n_270), .Y(n_353) );
NAND2xp5_ASAP7_75t_L g406 ( .A(n_270), .B(n_407), .Y(n_406) );
NAND2xp5_ASAP7_75t_L g382 ( .A(n_272), .B(n_348), .Y(n_382) );
AND2x4_ASAP7_75t_L g293 ( .A(n_273), .B(n_294), .Y(n_293) );
CKINVDCx16_ASAP7_75t_R g274 ( .A(n_275), .Y(n_274) );
OR2x2_ASAP7_75t_L g276 ( .A(n_277), .B(n_278), .Y(n_276) );
INVx2_ASAP7_75t_L g372 ( .A(n_278), .Y(n_372) );
NOR2xp33_ASAP7_75t_L g389 ( .A(n_278), .B(n_390), .Y(n_389) );
AND2x2_ASAP7_75t_L g320 ( .A(n_279), .B(n_310), .Y(n_320) );
AND2x2_ASAP7_75t_L g414 ( .A(n_279), .B(n_284), .Y(n_414) );
INVx1_ASAP7_75t_L g439 ( .A(n_279), .Y(n_439) );
AOI221xp5_ASAP7_75t_L g280 ( .A1(n_281), .A2(n_285), .B1(n_288), .B2(n_289), .C(n_295), .Y(n_280) );
CKINVDCx14_ASAP7_75t_R g301 ( .A(n_281), .Y(n_301) );
AND2x2_ASAP7_75t_L g281 ( .A(n_282), .B(n_283), .Y(n_281) );
NAND2xp5_ASAP7_75t_L g302 ( .A(n_282), .B(n_303), .Y(n_302) );
NAND2xp5_ASAP7_75t_L g355 ( .A(n_285), .B(n_336), .Y(n_355) );
INVx3_ASAP7_75t_SL g285 ( .A(n_286), .Y(n_285) );
OR2x2_ASAP7_75t_L g404 ( .A(n_286), .B(n_300), .Y(n_404) );
AND2x2_ASAP7_75t_L g318 ( .A(n_287), .B(n_319), .Y(n_318) );
INVx1_ASAP7_75t_L g348 ( .A(n_287), .Y(n_348) );
NAND2xp5_ASAP7_75t_L g376 ( .A(n_287), .B(n_331), .Y(n_376) );
NOR3xp33_ASAP7_75t_L g418 ( .A(n_287), .B(n_388), .C(n_419), .Y(n_418) );
AOI211xp5_ASAP7_75t_SL g351 ( .A1(n_288), .A2(n_352), .B(n_354), .C(n_362), .Y(n_351) );
INVx1_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
OAI22xp33_ASAP7_75t_L g340 ( .A1(n_290), .A2(n_341), .B1(n_342), .B2(n_343), .Y(n_340) );
NAND2xp5_ASAP7_75t_L g290 ( .A(n_291), .B(n_293), .Y(n_290) );
NAND2xp5_ASAP7_75t_L g329 ( .A(n_291), .B(n_330), .Y(n_329) );
NAND2xp5_ASAP7_75t_L g374 ( .A(n_291), .B(n_375), .Y(n_374) );
BUFx2_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
AND2x2_ASAP7_75t_L g433 ( .A(n_293), .B(n_407), .Y(n_433) );
OAI22xp5_ASAP7_75t_L g295 ( .A1(n_296), .A2(n_301), .B1(n_302), .B2(n_304), .Y(n_295) );
NOR2xp33_ASAP7_75t_SL g296 ( .A(n_297), .B(n_299), .Y(n_296) );
INVx1_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
NAND2xp5_ASAP7_75t_L g379 ( .A(n_299), .B(n_348), .Y(n_379) );
INVx1_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
OAI22xp5_ASAP7_75t_L g431 ( .A1(n_302), .A2(n_394), .B1(n_425), .B2(n_432), .Y(n_431) );
AOI221xp5_ASAP7_75t_L g305 ( .A1(n_306), .A2(n_313), .B1(n_315), .B2(n_320), .C(n_321), .Y(n_305) );
INVx1_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
OR2x2_ASAP7_75t_L g307 ( .A(n_308), .B(n_311), .Y(n_307) );
HB1xp67_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
INVxp67_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
OAI221xp5_ASAP7_75t_L g321 ( .A1(n_311), .A2(n_322), .B1(n_328), .B2(n_329), .C(n_332), .Y(n_321) );
INVx1_ASAP7_75t_L g364 ( .A(n_312), .Y(n_364) );
INVx1_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
INVx1_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
NAND2xp5_ASAP7_75t_L g316 ( .A(n_317), .B(n_318), .Y(n_316) );
INVx1_ASAP7_75t_SL g336 ( .A(n_317), .Y(n_336) );
OR2x2_ASAP7_75t_L g409 ( .A(n_317), .B(n_341), .Y(n_409) );
AND2x2_ASAP7_75t_L g411 ( .A(n_317), .B(n_319), .Y(n_411) );
INVx1_ASAP7_75t_L g350 ( .A(n_320), .Y(n_350) );
OR2x2_ASAP7_75t_L g322 ( .A(n_323), .B(n_326), .Y(n_322) );
AOI21xp33_ASAP7_75t_SL g380 ( .A1(n_323), .A2(n_381), .B(n_382), .Y(n_380) );
OR2x2_ASAP7_75t_L g387 ( .A(n_323), .B(n_388), .Y(n_387) );
INVx1_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
AND2x2_ASAP7_75t_L g361 ( .A(n_324), .B(n_345), .Y(n_361) );
INVx1_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
NAND2xp33_ASAP7_75t_SL g378 ( .A(n_329), .B(n_379), .Y(n_378) );
NAND2xp5_ASAP7_75t_L g347 ( .A(n_330), .B(n_348), .Y(n_347) );
NAND2xp5_ASAP7_75t_L g430 ( .A(n_331), .B(n_367), .Y(n_430) );
O2A1O1Ixp33_ASAP7_75t_L g346 ( .A1(n_334), .A2(n_347), .B(n_349), .C(n_350), .Y(n_346) );
NAND2x1_ASAP7_75t_SL g371 ( .A(n_334), .B(n_372), .Y(n_371) );
AOI22xp5_ASAP7_75t_L g383 ( .A1(n_335), .A2(n_384), .B1(n_386), .B2(n_389), .Y(n_383) );
AND2x2_ASAP7_75t_L g335 ( .A(n_336), .B(n_337), .Y(n_335) );
NAND2xp5_ASAP7_75t_L g426 ( .A(n_337), .B(n_427), .Y(n_426) );
NAND5xp2_ASAP7_75t_L g338 ( .A(n_339), .B(n_351), .C(n_369), .D(n_383), .E(n_392), .Y(n_338) );
NOR2xp33_ASAP7_75t_L g339 ( .A(n_340), .B(n_346), .Y(n_339) );
INVx1_ASAP7_75t_L g396 ( .A(n_342), .Y(n_396) );
INVx1_ASAP7_75t_SL g343 ( .A(n_344), .Y(n_343) );
AOI221xp5_ASAP7_75t_L g402 ( .A1(n_344), .A2(n_363), .B1(n_403), .B2(n_405), .C(n_408), .Y(n_402) );
NAND2xp5_ASAP7_75t_L g438 ( .A(n_345), .B(n_439), .Y(n_438) );
NOR2xp33_ASAP7_75t_L g352 ( .A(n_348), .B(n_353), .Y(n_352) );
NAND2xp5_ASAP7_75t_L g417 ( .A(n_348), .B(n_414), .Y(n_417) );
OAI22xp5_ASAP7_75t_L g354 ( .A1(n_355), .A2(n_356), .B1(n_358), .B2(n_360), .Y(n_354) );
INVx1_ASAP7_75t_SL g356 ( .A(n_357), .Y(n_356) );
INVx1_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
INVx1_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
AND2x2_ASAP7_75t_L g362 ( .A(n_363), .B(n_366), .Y(n_362) );
AND2x2_ASAP7_75t_L g363 ( .A(n_364), .B(n_365), .Y(n_363) );
AND2x2_ASAP7_75t_L g436 ( .A(n_365), .B(n_437), .Y(n_436) );
INVx1_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
AOI221xp5_ASAP7_75t_L g369 ( .A1(n_370), .A2(n_373), .B1(n_377), .B2(n_378), .C(n_380), .Y(n_369) );
INVx1_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
INVx1_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
AND2x2_ASAP7_75t_L g420 ( .A(n_375), .B(n_421), .Y(n_420) );
INVx1_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
INVx1_ASAP7_75t_SL g427 ( .A(n_385), .Y(n_427) );
INVx1_ASAP7_75t_SL g386 ( .A(n_387), .Y(n_386) );
INVx1_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
OAI21xp5_ASAP7_75t_SL g392 ( .A1(n_393), .A2(n_395), .B(n_396), .Y(n_392) );
INVx1_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
OAI211xp5_ASAP7_75t_SL g397 ( .A1(n_398), .A2(n_400), .B(n_402), .C(n_415), .Y(n_397) );
INVx1_ASAP7_75t_SL g398 ( .A(n_399), .Y(n_398) );
A2O1A1Ixp33_ASAP7_75t_L g424 ( .A1(n_400), .A2(n_425), .B(n_426), .C(n_428), .Y(n_424) );
INVx1_ASAP7_75t_SL g400 ( .A(n_401), .Y(n_400) );
INVx1_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
NAND2xp5_ASAP7_75t_SL g405 ( .A(n_404), .B(n_406), .Y(n_405) );
AOI21xp33_ASAP7_75t_L g408 ( .A1(n_409), .A2(n_410), .B(n_412), .Y(n_408) );
INVx1_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
INVx1_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
INVx1_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
INVx1_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
INVx1_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
INVx2_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
AOI21xp33_ASAP7_75t_L g434 ( .A1(n_435), .A2(n_438), .B(n_440), .Y(n_434) );
INVx1_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
INVx2_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
INVx2_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
INVx1_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
INVx1_ASAP7_75t_L g724 ( .A(n_446), .Y(n_724) );
INVx1_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
INVx2_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
OR5x1_ASAP7_75t_L g448 ( .A(n_449), .B(n_612), .C(n_670), .D(n_706), .E(n_713), .Y(n_448) );
NAND3xp33_ASAP7_75t_SL g449 ( .A(n_450), .B(n_558), .C(n_582), .Y(n_449) );
AOI221xp5_ASAP7_75t_L g450 ( .A1(n_451), .A2(n_494), .B1(n_524), .B2(n_529), .C(n_539), .Y(n_450) );
OAI21xp5_ASAP7_75t_SL g692 ( .A1(n_451), .A2(n_693), .B(n_695), .Y(n_692) );
AND2x2_ASAP7_75t_L g451 ( .A(n_452), .B(n_477), .Y(n_451) );
NAND2x1p5_ASAP7_75t_L g682 ( .A(n_452), .B(n_683), .Y(n_682) );
AND2x2_ASAP7_75t_L g452 ( .A(n_453), .B(n_466), .Y(n_452) );
INVx2_ASAP7_75t_L g528 ( .A(n_453), .Y(n_528) );
AND2x2_ASAP7_75t_L g541 ( .A(n_453), .B(n_479), .Y(n_541) );
AND2x2_ASAP7_75t_L g595 ( .A(n_453), .B(n_478), .Y(n_595) );
NAND2xp5_ASAP7_75t_L g610 ( .A(n_453), .B(n_467), .Y(n_610) );
O2A1O1Ixp33_ASAP7_75t_L g459 ( .A1(n_460), .A2(n_462), .B(n_463), .C(n_464), .Y(n_459) );
INVx2_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
AOI21xp5_ASAP7_75t_L g484 ( .A1(n_464), .A2(n_485), .B(n_486), .Y(n_484) );
AND2x2_ASAP7_75t_L g628 ( .A(n_466), .B(n_569), .Y(n_628) );
AND2x2_ASAP7_75t_L g661 ( .A(n_466), .B(n_479), .Y(n_661) );
INVx2_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
OR2x2_ASAP7_75t_L g568 ( .A(n_467), .B(n_569), .Y(n_568) );
AND2x2_ASAP7_75t_L g581 ( .A(n_467), .B(n_479), .Y(n_581) );
AND2x2_ASAP7_75t_L g588 ( .A(n_467), .B(n_569), .Y(n_588) );
HB1xp67_ASAP7_75t_L g597 ( .A(n_467), .Y(n_597) );
AND2x2_ASAP7_75t_L g604 ( .A(n_467), .B(n_478), .Y(n_604) );
INVx1_ASAP7_75t_L g635 ( .A(n_467), .Y(n_635) );
OAI21xp5_ASAP7_75t_L g468 ( .A1(n_469), .A2(n_472), .B(n_475), .Y(n_468) );
INVx1_ASAP7_75t_L g611 ( .A(n_477), .Y(n_611) );
AND2x2_ASAP7_75t_L g477 ( .A(n_478), .B(n_488), .Y(n_477) );
INVx2_ASAP7_75t_L g567 ( .A(n_478), .Y(n_567) );
AND2x2_ASAP7_75t_L g589 ( .A(n_478), .B(n_528), .Y(n_589) );
NAND2xp5_ASAP7_75t_L g640 ( .A(n_478), .B(n_635), .Y(n_640) );
INVx3_ASAP7_75t_L g478 ( .A(n_479), .Y(n_478) );
NAND2xp5_ASAP7_75t_L g527 ( .A(n_479), .B(n_528), .Y(n_527) );
AND2x2_ASAP7_75t_L g712 ( .A(n_479), .B(n_676), .Y(n_712) );
INVx2_ASAP7_75t_L g526 ( .A(n_488), .Y(n_526) );
INVx3_ASAP7_75t_L g627 ( .A(n_488), .Y(n_627) );
OR2x2_ASAP7_75t_L g657 ( .A(n_488), .B(n_658), .Y(n_657) );
NOR2x1_ASAP7_75t_L g683 ( .A(n_488), .B(n_567), .Y(n_683) );
AND2x4_ASAP7_75t_L g488 ( .A(n_489), .B(n_490), .Y(n_488) );
INVx1_ASAP7_75t_L g570 ( .A(n_489), .Y(n_570) );
AOI33xp33_ASAP7_75t_L g703 ( .A1(n_494), .A2(n_541), .A3(n_555), .B1(n_627), .B2(n_704), .B3(n_705), .Y(n_703) );
INVx1_ASAP7_75t_L g494 ( .A(n_495), .Y(n_494) );
OR2x2_ASAP7_75t_L g495 ( .A(n_496), .B(n_503), .Y(n_495) );
OR2x2_ASAP7_75t_L g556 ( .A(n_496), .B(n_557), .Y(n_556) );
NOR2xp33_ASAP7_75t_L g615 ( .A(n_496), .B(n_553), .Y(n_615) );
OR2x2_ASAP7_75t_L g668 ( .A(n_496), .B(n_669), .Y(n_668) );
INVx2_ASAP7_75t_L g496 ( .A(n_497), .Y(n_496) );
AND2x2_ASAP7_75t_L g594 ( .A(n_497), .B(n_595), .Y(n_594) );
OR2x2_ASAP7_75t_L g619 ( .A(n_497), .B(n_503), .Y(n_619) );
AND2x2_ASAP7_75t_L g686 ( .A(n_497), .B(n_531), .Y(n_686) );
AOI21xp5_ASAP7_75t_L g711 ( .A1(n_497), .A2(n_586), .B(n_712), .Y(n_711) );
BUFx6f_ASAP7_75t_L g497 ( .A(n_498), .Y(n_497) );
INVx1_ASAP7_75t_L g533 ( .A(n_498), .Y(n_533) );
INVx1_ASAP7_75t_L g546 ( .A(n_498), .Y(n_546) );
AND2x2_ASAP7_75t_L g565 ( .A(n_498), .B(n_535), .Y(n_565) );
AND2x2_ASAP7_75t_L g614 ( .A(n_498), .B(n_534), .Y(n_614) );
INVx2_ASAP7_75t_SL g656 ( .A(n_503), .Y(n_656) );
OR2x2_ASAP7_75t_L g503 ( .A(n_504), .B(n_514), .Y(n_503) );
INVx2_ASAP7_75t_L g576 ( .A(n_504), .Y(n_576) );
INVx1_ASAP7_75t_L g707 ( .A(n_504), .Y(n_707) );
AND2x2_ASAP7_75t_L g720 ( .A(n_504), .B(n_601), .Y(n_720) );
INVx2_ASAP7_75t_L g504 ( .A(n_505), .Y(n_504) );
INVx2_ASAP7_75t_L g547 ( .A(n_505), .Y(n_547) );
OR2x2_ASAP7_75t_L g553 ( .A(n_505), .B(n_554), .Y(n_553) );
HB1xp67_ASAP7_75t_L g564 ( .A(n_505), .Y(n_564) );
HB1xp67_ASAP7_75t_L g531 ( .A(n_514), .Y(n_531) );
AND2x2_ASAP7_75t_L g548 ( .A(n_514), .B(n_534), .Y(n_548) );
INVx1_ASAP7_75t_L g554 ( .A(n_514), .Y(n_554) );
INVx1_ASAP7_75t_L g561 ( .A(n_514), .Y(n_561) );
AND2x2_ASAP7_75t_L g586 ( .A(n_514), .B(n_535), .Y(n_586) );
INVx2_ASAP7_75t_L g602 ( .A(n_514), .Y(n_602) );
AND2x2_ASAP7_75t_L g695 ( .A(n_514), .B(n_696), .Y(n_695) );
NAND2xp5_ASAP7_75t_L g716 ( .A(n_514), .B(n_576), .Y(n_716) );
AOI21xp5_ASAP7_75t_L g516 ( .A1(n_517), .A2(n_518), .B(n_519), .Y(n_516) );
INVx1_ASAP7_75t_SL g524 ( .A(n_525), .Y(n_524) );
OR2x2_ASAP7_75t_L g525 ( .A(n_526), .B(n_527), .Y(n_525) );
INVx2_ASAP7_75t_L g550 ( .A(n_526), .Y(n_550) );
INVx1_ASAP7_75t_L g579 ( .A(n_526), .Y(n_579) );
NOR2xp33_ASAP7_75t_L g676 ( .A(n_526), .B(n_610), .Y(n_676) );
INVx1_ASAP7_75t_SL g636 ( .A(n_527), .Y(n_636) );
INVx2_ASAP7_75t_L g557 ( .A(n_528), .Y(n_557) );
AND2x2_ASAP7_75t_L g626 ( .A(n_528), .B(n_627), .Y(n_626) );
AND2x2_ASAP7_75t_L g642 ( .A(n_528), .B(n_643), .Y(n_642) );
AND2x2_ASAP7_75t_L g529 ( .A(n_530), .B(n_532), .Y(n_529) );
INVx1_ASAP7_75t_L g704 ( .A(n_530), .Y(n_704) );
INVx1_ASAP7_75t_L g530 ( .A(n_531), .Y(n_530) );
AND2x2_ASAP7_75t_L g559 ( .A(n_532), .B(n_560), .Y(n_559) );
AND2x2_ASAP7_75t_L g662 ( .A(n_532), .B(n_652), .Y(n_662) );
AOI21xp5_ASAP7_75t_L g714 ( .A1(n_532), .A2(n_673), .B(n_715), .Y(n_714) );
AND2x2_ASAP7_75t_L g532 ( .A(n_533), .B(n_534), .Y(n_532) );
AND2x2_ASAP7_75t_L g575 ( .A(n_533), .B(n_576), .Y(n_575) );
BUFx2_ASAP7_75t_L g600 ( .A(n_533), .Y(n_600) );
INVx1_ASAP7_75t_L g624 ( .A(n_533), .Y(n_624) );
OR2x2_ASAP7_75t_L g688 ( .A(n_534), .B(n_547), .Y(n_688) );
NOR2xp67_ASAP7_75t_L g696 ( .A(n_534), .B(n_697), .Y(n_696) );
INVx2_ASAP7_75t_L g534 ( .A(n_535), .Y(n_534) );
AND2x2_ASAP7_75t_L g601 ( .A(n_535), .B(n_602), .Y(n_601) );
BUFx2_ASAP7_75t_L g608 ( .A(n_535), .Y(n_608) );
OAI22xp5_ASAP7_75t_L g539 ( .A1(n_540), .A2(n_542), .B1(n_549), .B2(n_551), .Y(n_539) );
OR2x2_ASAP7_75t_L g618 ( .A(n_540), .B(n_568), .Y(n_618) );
INVx1_ASAP7_75t_SL g540 ( .A(n_541), .Y(n_540) );
AOI222xp33_ASAP7_75t_L g659 ( .A1(n_541), .A2(n_660), .B1(n_662), .B2(n_663), .C1(n_664), .C2(n_667), .Y(n_659) );
INVx1_ASAP7_75t_L g542 ( .A(n_543), .Y(n_542) );
AND2x2_ASAP7_75t_L g543 ( .A(n_544), .B(n_548), .Y(n_543) );
INVx1_ASAP7_75t_SL g544 ( .A(n_545), .Y(n_544) );
OR2x2_ASAP7_75t_L g606 ( .A(n_545), .B(n_607), .Y(n_606) );
NAND2xp5_ASAP7_75t_L g545 ( .A(n_546), .B(n_547), .Y(n_545) );
AND2x2_ASAP7_75t_SL g560 ( .A(n_547), .B(n_561), .Y(n_560) );
HB1xp67_ASAP7_75t_L g631 ( .A(n_547), .Y(n_631) );
AND2x2_ASAP7_75t_L g679 ( .A(n_547), .B(n_548), .Y(n_679) );
INVx1_ASAP7_75t_L g697 ( .A(n_547), .Y(n_697) );
INVx1_ASAP7_75t_L g549 ( .A(n_550), .Y(n_549) );
AND2x2_ASAP7_75t_L g663 ( .A(n_550), .B(n_589), .Y(n_663) );
AND2x2_ASAP7_75t_L g705 ( .A(n_550), .B(n_581), .Y(n_705) );
NAND2xp5_ASAP7_75t_L g551 ( .A(n_552), .B(n_555), .Y(n_551) );
NAND2xp5_ASAP7_75t_L g687 ( .A(n_552), .B(n_600), .Y(n_687) );
INVx2_ASAP7_75t_L g552 ( .A(n_553), .Y(n_552) );
NAND2xp5_ASAP7_75t_SL g584 ( .A(n_553), .B(n_585), .Y(n_584) );
INVx1_ASAP7_75t_L g555 ( .A(n_556), .Y(n_555) );
AND2x2_ASAP7_75t_L g580 ( .A(n_557), .B(n_581), .Y(n_580) );
INVx3_ASAP7_75t_L g648 ( .A(n_557), .Y(n_648) );
O2A1O1Ixp33_ASAP7_75t_L g558 ( .A1(n_559), .A2(n_562), .B(n_566), .C(n_571), .Y(n_558) );
INVxp67_ASAP7_75t_L g572 ( .A(n_559), .Y(n_572) );
NAND2xp5_ASAP7_75t_L g623 ( .A(n_560), .B(n_624), .Y(n_623) );
NAND2xp5_ASAP7_75t_L g702 ( .A(n_560), .B(n_607), .Y(n_702) );
BUFx3_ASAP7_75t_L g666 ( .A(n_561), .Y(n_666) );
INVx1_ASAP7_75t_L g573 ( .A(n_562), .Y(n_573) );
AND2x2_ASAP7_75t_L g562 ( .A(n_563), .B(n_565), .Y(n_562) );
INVx1_ASAP7_75t_L g563 ( .A(n_564), .Y(n_563) );
AND2x2_ASAP7_75t_L g592 ( .A(n_564), .B(n_586), .Y(n_592) );
INVx1_ASAP7_75t_SL g632 ( .A(n_565), .Y(n_632) );
NOR2xp33_ASAP7_75t_L g566 ( .A(n_567), .B(n_568), .Y(n_566) );
INVx1_ASAP7_75t_L g622 ( .A(n_567), .Y(n_622) );
AND2x2_ASAP7_75t_L g645 ( .A(n_567), .B(n_628), .Y(n_645) );
INVx1_ASAP7_75t_SL g616 ( .A(n_568), .Y(n_616) );
INVx1_ASAP7_75t_L g643 ( .A(n_569), .Y(n_643) );
AOI31xp33_ASAP7_75t_L g571 ( .A1(n_572), .A2(n_573), .A3(n_574), .B(n_577), .Y(n_571) );
INVx1_ASAP7_75t_L g574 ( .A(n_575), .Y(n_574) );
AND2x2_ASAP7_75t_L g664 ( .A(n_575), .B(n_665), .Y(n_664) );
INVx1_ASAP7_75t_L g638 ( .A(n_576), .Y(n_638) );
BUFx2_ASAP7_75t_L g652 ( .A(n_576), .Y(n_652) );
AND2x2_ASAP7_75t_L g680 ( .A(n_576), .B(n_601), .Y(n_680) );
NAND2xp5_ASAP7_75t_L g577 ( .A(n_578), .B(n_580), .Y(n_577) );
INVx1_ASAP7_75t_L g578 ( .A(n_579), .Y(n_578) );
INVx1_ASAP7_75t_SL g653 ( .A(n_580), .Y(n_653) );
NAND2xp5_ASAP7_75t_L g694 ( .A(n_581), .B(n_648), .Y(n_694) );
AND2x2_ASAP7_75t_L g701 ( .A(n_581), .B(n_627), .Y(n_701) );
AOI211xp5_ASAP7_75t_L g582 ( .A1(n_583), .A2(n_587), .B(n_590), .C(n_605), .Y(n_582) );
INVxp67_ASAP7_75t_L g583 ( .A(n_584), .Y(n_583) );
INVx2_ASAP7_75t_L g585 ( .A(n_586), .Y(n_585) );
AOI221xp5_ASAP7_75t_L g613 ( .A1(n_587), .A2(n_614), .B1(n_615), .B2(n_616), .C(n_617), .Y(n_613) );
AND2x2_ASAP7_75t_L g587 ( .A(n_588), .B(n_589), .Y(n_587) );
AND2x2_ASAP7_75t_L g621 ( .A(n_588), .B(n_622), .Y(n_621) );
INVx2_ASAP7_75t_L g658 ( .A(n_589), .Y(n_658) );
OAI32xp33_ASAP7_75t_L g590 ( .A1(n_591), .A2(n_593), .A3(n_596), .B1(n_598), .B2(n_603), .Y(n_590) );
INVx1_ASAP7_75t_L g591 ( .A(n_592), .Y(n_591) );
O2A1O1Ixp33_ASAP7_75t_L g644 ( .A1(n_592), .A2(n_645), .B(n_646), .C(n_649), .Y(n_644) );
INVx1_ASAP7_75t_L g593 ( .A(n_594), .Y(n_593) );
INVx1_ASAP7_75t_L g596 ( .A(n_597), .Y(n_596) );
INVx1_ASAP7_75t_L g598 ( .A(n_599), .Y(n_598) );
AND2x2_ASAP7_75t_L g599 ( .A(n_600), .B(n_601), .Y(n_599) );
OAI21xp5_ASAP7_75t_SL g708 ( .A1(n_600), .A2(n_709), .B(n_710), .Y(n_708) );
INVx1_ASAP7_75t_L g669 ( .A(n_601), .Y(n_669) );
INVxp67_ASAP7_75t_L g603 ( .A(n_604), .Y(n_603) );
NOR2xp33_ASAP7_75t_L g605 ( .A(n_606), .B(n_609), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g637 ( .A(n_607), .B(n_638), .Y(n_637) );
AND2x2_ASAP7_75t_L g655 ( .A(n_607), .B(n_656), .Y(n_655) );
INVx2_ASAP7_75t_L g607 ( .A(n_608), .Y(n_607) );
INVx1_ASAP7_75t_L g672 ( .A(n_609), .Y(n_672) );
OR2x2_ASAP7_75t_L g609 ( .A(n_610), .B(n_611), .Y(n_609) );
NAND4xp25_ASAP7_75t_SL g612 ( .A(n_613), .B(n_625), .C(n_644), .D(n_659), .Y(n_612) );
AND2x2_ASAP7_75t_L g651 ( .A(n_614), .B(n_652), .Y(n_651) );
AND2x4_ASAP7_75t_L g673 ( .A(n_614), .B(n_666), .Y(n_673) );
NAND2xp5_ASAP7_75t_L g647 ( .A(n_616), .B(n_648), .Y(n_647) );
OAI22xp5_ASAP7_75t_L g617 ( .A1(n_618), .A2(n_619), .B1(n_620), .B2(n_623), .Y(n_617) );
OAI22xp5_ASAP7_75t_L g699 ( .A1(n_618), .A2(n_669), .B1(n_700), .B2(n_702), .Y(n_699) );
O2A1O1Ixp33_ASAP7_75t_L g706 ( .A1(n_618), .A2(n_707), .B(n_708), .C(n_711), .Y(n_706) );
INVx2_ASAP7_75t_L g677 ( .A(n_619), .Y(n_677) );
INVx1_ASAP7_75t_L g620 ( .A(n_621), .Y(n_620) );
AOI222xp33_ASAP7_75t_L g671 ( .A1(n_621), .A2(n_655), .B1(n_672), .B2(n_673), .C1(n_674), .C2(n_677), .Y(n_671) );
O2A1O1Ixp33_ASAP7_75t_L g625 ( .A1(n_626), .A2(n_628), .B(n_629), .C(n_633), .Y(n_625) );
INVx1_ASAP7_75t_L g691 ( .A(n_626), .Y(n_691) );
INVx1_ASAP7_75t_L g629 ( .A(n_630), .Y(n_629) );
OAI22xp33_ASAP7_75t_L g633 ( .A1(n_630), .A2(n_634), .B1(n_637), .B2(n_639), .Y(n_633) );
OR2x2_ASAP7_75t_L g630 ( .A(n_631), .B(n_632), .Y(n_630) );
NAND2xp5_ASAP7_75t_L g634 ( .A(n_635), .B(n_636), .Y(n_634) );
OR2x2_ASAP7_75t_L g639 ( .A(n_640), .B(n_641), .Y(n_639) );
INVx1_ASAP7_75t_L g641 ( .A(n_642), .Y(n_641) );
AND2x2_ASAP7_75t_L g660 ( .A(n_642), .B(n_661), .Y(n_660) );
INVx1_ASAP7_75t_L g718 ( .A(n_645), .Y(n_718) );
INVx1_ASAP7_75t_L g646 ( .A(n_647), .Y(n_646) );
OAI22xp33_ASAP7_75t_L g649 ( .A1(n_650), .A2(n_653), .B1(n_654), .B2(n_657), .Y(n_649) );
INVx1_ASAP7_75t_L g650 ( .A(n_651), .Y(n_650) );
NAND2xp5_ASAP7_75t_L g685 ( .A(n_652), .B(n_686), .Y(n_685) );
INVx1_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
INVx1_ASAP7_75t_L g709 ( .A(n_657), .Y(n_709) );
INVx1_ASAP7_75t_L g690 ( .A(n_661), .Y(n_690) );
CKINVDCx16_ASAP7_75t_R g717 ( .A(n_663), .Y(n_717) );
INVxp67_ASAP7_75t_L g665 ( .A(n_666), .Y(n_665) );
INVx1_ASAP7_75t_L g667 ( .A(n_668), .Y(n_667) );
NAND5xp2_ASAP7_75t_L g670 ( .A(n_671), .B(n_678), .C(n_692), .D(n_698), .E(n_703), .Y(n_670) );
INVx1_ASAP7_75t_SL g674 ( .A(n_675), .Y(n_674) );
INVx1_ASAP7_75t_L g675 ( .A(n_676), .Y(n_675) );
O2A1O1Ixp33_ASAP7_75t_L g678 ( .A1(n_679), .A2(n_680), .B(n_681), .C(n_684), .Y(n_678) );
INVx1_ASAP7_75t_L g681 ( .A(n_682), .Y(n_681) );
AOI31xp33_ASAP7_75t_L g684 ( .A1(n_685), .A2(n_687), .A3(n_688), .B(n_689), .Y(n_684) );
INVx1_ASAP7_75t_L g710 ( .A(n_686), .Y(n_710) );
OR2x2_ASAP7_75t_L g689 ( .A(n_690), .B(n_691), .Y(n_689) );
INVx1_ASAP7_75t_L g693 ( .A(n_694), .Y(n_693) );
INVx1_ASAP7_75t_L g698 ( .A(n_699), .Y(n_698) );
OAI222xp33_ASAP7_75t_L g713 ( .A1(n_700), .A2(n_702), .B1(n_714), .B2(n_717), .C1(n_718), .C2(n_719), .Y(n_713) );
INVx1_ASAP7_75t_L g700 ( .A(n_701), .Y(n_700) );
INVx1_ASAP7_75t_L g715 ( .A(n_716), .Y(n_715) );
INVx2_ASAP7_75t_SL g719 ( .A(n_720), .Y(n_719) );
INVx1_ASAP7_75t_L g725 ( .A(n_726), .Y(n_725) );
INVx2_ASAP7_75t_L g726 ( .A(n_727), .Y(n_726) );
INVx2_ASAP7_75t_SL g728 ( .A(n_729), .Y(n_728) );
CKINVDCx20_ASAP7_75t_R g732 ( .A(n_733), .Y(n_732) );
CKINVDCx14_ASAP7_75t_R g738 ( .A(n_734), .Y(n_738) );
INVx1_ASAP7_75t_SL g739 ( .A(n_740), .Y(n_739) );
INVx1_ASAP7_75t_L g741 ( .A(n_742), .Y(n_741) );
INVx1_ASAP7_75t_L g742 ( .A(n_743), .Y(n_742) );
endmodule