module fake_aes_11441_n_632 (n_44, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_6, n_4, n_40, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_632);
input n_44;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_6;
input n_4;
input n_40;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_632;
wire n_117;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_612;
wire n_154;
wire n_328;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_162;
wire n_387;
wire n_163;
wire n_476;
wire n_105;
wire n_227;
wire n_384;
wire n_434;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_586;
wire n_244;
wire n_540;
wire n_563;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_367;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_108;
wire n_91;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_293;
wire n_533;
wire n_506;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_307;
wire n_191;
wire n_610;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_482;
wire n_394;
wire n_415;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_77;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_172;
wire n_329;
wire n_251;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_621;
wire n_370;
wire n_589;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_90;
wire n_357;
wire n_260;
wire n_78;
wire n_539;
wire n_201;
wire n_197;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_208;
wire n_200;
wire n_573;
wire n_126;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_295;
wire n_143;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_552;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_438;
wire n_134;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_618;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_84;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_132;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx4_ASAP7_75t_R g77 ( .A(n_17), .Y(n_77) );
HB1xp67_ASAP7_75t_L g78 ( .A(n_14), .Y(n_78) );
INVx1_ASAP7_75t_SL g79 ( .A(n_53), .Y(n_79) );
INVx1_ASAP7_75t_L g80 ( .A(n_9), .Y(n_80) );
INVx1_ASAP7_75t_L g81 ( .A(n_20), .Y(n_81) );
INVxp33_ASAP7_75t_SL g82 ( .A(n_47), .Y(n_82) );
INVx1_ASAP7_75t_L g83 ( .A(n_10), .Y(n_83) );
INVx1_ASAP7_75t_L g84 ( .A(n_56), .Y(n_84) );
INVx1_ASAP7_75t_L g85 ( .A(n_43), .Y(n_85) );
INVx1_ASAP7_75t_L g86 ( .A(n_72), .Y(n_86) );
BUFx3_ASAP7_75t_L g87 ( .A(n_0), .Y(n_87) );
CKINVDCx5p33_ASAP7_75t_R g88 ( .A(n_38), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_18), .Y(n_89) );
INVx1_ASAP7_75t_L g90 ( .A(n_24), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_3), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_12), .Y(n_92) );
CKINVDCx5p33_ASAP7_75t_R g93 ( .A(n_11), .Y(n_93) );
CKINVDCx5p33_ASAP7_75t_R g94 ( .A(n_69), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_36), .Y(n_95) );
CKINVDCx5p33_ASAP7_75t_R g96 ( .A(n_34), .Y(n_96) );
CKINVDCx20_ASAP7_75t_R g97 ( .A(n_18), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_12), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_67), .Y(n_99) );
CKINVDCx5p33_ASAP7_75t_R g100 ( .A(n_32), .Y(n_100) );
NAND2xp5_ASAP7_75t_L g101 ( .A(n_14), .B(n_51), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_65), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_29), .Y(n_103) );
CKINVDCx5p33_ASAP7_75t_R g104 ( .A(n_71), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_11), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_27), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_45), .Y(n_107) );
BUFx6f_ASAP7_75t_L g108 ( .A(n_10), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_57), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_4), .Y(n_110) );
CKINVDCx5p33_ASAP7_75t_R g111 ( .A(n_37), .Y(n_111) );
INVxp33_ASAP7_75t_SL g112 ( .A(n_76), .Y(n_112) );
INVxp67_ASAP7_75t_L g113 ( .A(n_8), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_70), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_7), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_25), .Y(n_116) );
CKINVDCx16_ASAP7_75t_R g117 ( .A(n_4), .Y(n_117) );
CKINVDCx20_ASAP7_75t_R g118 ( .A(n_1), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_22), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_0), .Y(n_120) );
INVx2_ASAP7_75t_L g121 ( .A(n_90), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_90), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_87), .Y(n_123) );
BUFx6f_ASAP7_75t_L g124 ( .A(n_108), .Y(n_124) );
INVx1_ASAP7_75t_L g125 ( .A(n_87), .Y(n_125) );
INVx3_ASAP7_75t_L g126 ( .A(n_108), .Y(n_126) );
INVx2_ASAP7_75t_L g127 ( .A(n_81), .Y(n_127) );
INVx1_ASAP7_75t_L g128 ( .A(n_84), .Y(n_128) );
INVx1_ASAP7_75t_L g129 ( .A(n_85), .Y(n_129) );
HB1xp67_ASAP7_75t_L g130 ( .A(n_78), .Y(n_130) );
BUFx6f_ASAP7_75t_L g131 ( .A(n_108), .Y(n_131) );
INVx1_ASAP7_75t_L g132 ( .A(n_86), .Y(n_132) );
INVx2_ASAP7_75t_L g133 ( .A(n_95), .Y(n_133) );
HB1xp67_ASAP7_75t_L g134 ( .A(n_93), .Y(n_134) );
BUFx6f_ASAP7_75t_L g135 ( .A(n_108), .Y(n_135) );
AND2x4_ASAP7_75t_L g136 ( .A(n_89), .B(n_1), .Y(n_136) );
AND2x4_ASAP7_75t_L g137 ( .A(n_89), .B(n_2), .Y(n_137) );
INVx4_ASAP7_75t_L g138 ( .A(n_88), .Y(n_138) );
BUFx8_ASAP7_75t_L g139 ( .A(n_99), .Y(n_139) );
INVx1_ASAP7_75t_L g140 ( .A(n_102), .Y(n_140) );
INVx4_ASAP7_75t_L g141 ( .A(n_88), .Y(n_141) );
INVx1_ASAP7_75t_L g142 ( .A(n_103), .Y(n_142) );
INVx2_ASAP7_75t_L g143 ( .A(n_106), .Y(n_143) );
BUFx8_ASAP7_75t_L g144 ( .A(n_107), .Y(n_144) );
HB1xp67_ASAP7_75t_L g145 ( .A(n_93), .Y(n_145) );
INVx1_ASAP7_75t_L g146 ( .A(n_109), .Y(n_146) );
AND2x2_ASAP7_75t_L g147 ( .A(n_117), .B(n_2), .Y(n_147) );
AND2x2_ASAP7_75t_L g148 ( .A(n_91), .B(n_3), .Y(n_148) );
OAI21x1_ASAP7_75t_L g149 ( .A1(n_114), .A2(n_119), .B(n_116), .Y(n_149) );
AND3x2_ASAP7_75t_L g150 ( .A(n_113), .B(n_91), .C(n_98), .Y(n_150) );
INVx1_ASAP7_75t_L g151 ( .A(n_108), .Y(n_151) );
AND2x4_ASAP7_75t_L g152 ( .A(n_120), .B(n_5), .Y(n_152) );
INVx4_ASAP7_75t_L g153 ( .A(n_94), .Y(n_153) );
INVx1_ASAP7_75t_L g154 ( .A(n_80), .Y(n_154) );
INVx1_ASAP7_75t_L g155 ( .A(n_83), .Y(n_155) );
BUFx2_ASAP7_75t_L g156 ( .A(n_94), .Y(n_156) );
INVx1_ASAP7_75t_L g157 ( .A(n_92), .Y(n_157) );
BUFx6f_ASAP7_75t_L g158 ( .A(n_105), .Y(n_158) );
AND2x2_ASAP7_75t_L g159 ( .A(n_156), .B(n_111), .Y(n_159) );
NAND2xp5_ASAP7_75t_L g160 ( .A(n_138), .B(n_96), .Y(n_160) );
INVx2_ASAP7_75t_L g161 ( .A(n_124), .Y(n_161) );
NAND2xp5_ASAP7_75t_L g162 ( .A(n_138), .B(n_96), .Y(n_162) );
INVx1_ASAP7_75t_L g163 ( .A(n_121), .Y(n_163) );
INVx1_ASAP7_75t_L g164 ( .A(n_121), .Y(n_164) );
AND2x4_ASAP7_75t_L g165 ( .A(n_136), .B(n_115), .Y(n_165) );
BUFx6f_ASAP7_75t_L g166 ( .A(n_124), .Y(n_166) );
AND2x4_ASAP7_75t_L g167 ( .A(n_136), .B(n_110), .Y(n_167) );
NAND2xp5_ASAP7_75t_L g168 ( .A(n_138), .B(n_111), .Y(n_168) );
CKINVDCx5p33_ASAP7_75t_R g169 ( .A(n_156), .Y(n_169) );
INVx1_ASAP7_75t_L g170 ( .A(n_121), .Y(n_170) );
INVx4_ASAP7_75t_L g171 ( .A(n_136), .Y(n_171) );
AND2x4_ASAP7_75t_L g172 ( .A(n_136), .B(n_104), .Y(n_172) );
INVx1_ASAP7_75t_L g173 ( .A(n_158), .Y(n_173) );
INVx1_ASAP7_75t_L g174 ( .A(n_158), .Y(n_174) );
AND2x2_ASAP7_75t_L g175 ( .A(n_130), .B(n_138), .Y(n_175) );
INVx2_ASAP7_75t_L g176 ( .A(n_124), .Y(n_176) );
AND2x6_ASAP7_75t_L g177 ( .A(n_137), .B(n_101), .Y(n_177) );
BUFx6f_ASAP7_75t_L g178 ( .A(n_124), .Y(n_178) );
AND2x4_ASAP7_75t_L g179 ( .A(n_137), .B(n_104), .Y(n_179) );
INVx2_ASAP7_75t_L g180 ( .A(n_124), .Y(n_180) );
NOR2xp33_ASAP7_75t_L g181 ( .A(n_141), .B(n_112), .Y(n_181) );
INVx2_ASAP7_75t_L g182 ( .A(n_124), .Y(n_182) );
INVx3_ASAP7_75t_L g183 ( .A(n_137), .Y(n_183) );
AND2x6_ASAP7_75t_L g184 ( .A(n_137), .B(n_79), .Y(n_184) );
NAND2xp5_ASAP7_75t_SL g185 ( .A(n_141), .B(n_100), .Y(n_185) );
INVx1_ASAP7_75t_L g186 ( .A(n_158), .Y(n_186) );
INVx2_ASAP7_75t_SL g187 ( .A(n_141), .Y(n_187) );
INVx1_ASAP7_75t_L g188 ( .A(n_158), .Y(n_188) );
INVx1_ASAP7_75t_L g189 ( .A(n_158), .Y(n_189) );
NAND2xp5_ASAP7_75t_L g190 ( .A(n_141), .B(n_100), .Y(n_190) );
INVx2_ASAP7_75t_L g191 ( .A(n_131), .Y(n_191) );
NAND2xp5_ASAP7_75t_L g192 ( .A(n_153), .B(n_112), .Y(n_192) );
INVx3_ASAP7_75t_L g193 ( .A(n_152), .Y(n_193) );
INVx1_ASAP7_75t_L g194 ( .A(n_158), .Y(n_194) );
INVx1_ASAP7_75t_L g195 ( .A(n_126), .Y(n_195) );
INVx1_ASAP7_75t_L g196 ( .A(n_126), .Y(n_196) );
INVx2_ASAP7_75t_SL g197 ( .A(n_153), .Y(n_197) );
NOR2xp33_ASAP7_75t_L g198 ( .A(n_153), .B(n_82), .Y(n_198) );
INVx1_ASAP7_75t_SL g199 ( .A(n_134), .Y(n_199) );
INVx2_ASAP7_75t_L g200 ( .A(n_131), .Y(n_200) );
AND2x2_ASAP7_75t_L g201 ( .A(n_130), .B(n_118), .Y(n_201) );
OAI22xp5_ASAP7_75t_L g202 ( .A1(n_134), .A2(n_118), .B1(n_97), .B2(n_82), .Y(n_202) );
AO22x2_ASAP7_75t_L g203 ( .A1(n_152), .A2(n_77), .B1(n_97), .B2(n_7), .Y(n_203) );
INVx1_ASAP7_75t_L g204 ( .A(n_126), .Y(n_204) );
INVx1_ASAP7_75t_L g205 ( .A(n_163), .Y(n_205) );
INVx3_ASAP7_75t_L g206 ( .A(n_171), .Y(n_206) );
INVx1_ASAP7_75t_L g207 ( .A(n_163), .Y(n_207) );
BUFx6f_ASAP7_75t_L g208 ( .A(n_164), .Y(n_208) );
INVx2_ASAP7_75t_SL g209 ( .A(n_159), .Y(n_209) );
INVx3_ASAP7_75t_L g210 ( .A(n_171), .Y(n_210) );
BUFx4f_ASAP7_75t_L g211 ( .A(n_184), .Y(n_211) );
INVx1_ASAP7_75t_L g212 ( .A(n_164), .Y(n_212) );
AO22x1_ASAP7_75t_L g213 ( .A1(n_184), .A2(n_144), .B1(n_139), .B2(n_152), .Y(n_213) );
INVx2_ASAP7_75t_L g214 ( .A(n_170), .Y(n_214) );
INVx2_ASAP7_75t_SL g215 ( .A(n_159), .Y(n_215) );
OR2x6_ASAP7_75t_L g216 ( .A(n_203), .B(n_147), .Y(n_216) );
BUFx3_ASAP7_75t_L g217 ( .A(n_184), .Y(n_217) );
INVx1_ASAP7_75t_L g218 ( .A(n_170), .Y(n_218) );
AND2x4_ASAP7_75t_SL g219 ( .A(n_175), .B(n_201), .Y(n_219) );
NAND2xp5_ASAP7_75t_L g220 ( .A(n_175), .B(n_153), .Y(n_220) );
CKINVDCx5p33_ASAP7_75t_R g221 ( .A(n_169), .Y(n_221) );
AOI21xp5_ASAP7_75t_L g222 ( .A1(n_183), .A2(n_149), .B(n_122), .Y(n_222) );
HB1xp67_ASAP7_75t_L g223 ( .A(n_199), .Y(n_223) );
BUFx6f_ASAP7_75t_L g224 ( .A(n_171), .Y(n_224) );
NAND2xp5_ASAP7_75t_SL g225 ( .A(n_172), .B(n_139), .Y(n_225) );
INVx1_ASAP7_75t_L g226 ( .A(n_165), .Y(n_226) );
NAND3xp33_ASAP7_75t_L g227 ( .A(n_169), .B(n_145), .C(n_144), .Y(n_227) );
INVx1_ASAP7_75t_L g228 ( .A(n_165), .Y(n_228) );
NAND2xp5_ASAP7_75t_SL g229 ( .A(n_172), .B(n_139), .Y(n_229) );
NAND2xp5_ASAP7_75t_L g230 ( .A(n_181), .B(n_145), .Y(n_230) );
INVxp67_ASAP7_75t_SL g231 ( .A(n_183), .Y(n_231) );
NAND2xp5_ASAP7_75t_SL g232 ( .A(n_172), .B(n_139), .Y(n_232) );
INVx1_ASAP7_75t_L g233 ( .A(n_165), .Y(n_233) );
INVx5_ASAP7_75t_L g234 ( .A(n_184), .Y(n_234) );
NOR2xp33_ASAP7_75t_L g235 ( .A(n_192), .B(n_150), .Y(n_235) );
AND2x2_ASAP7_75t_L g236 ( .A(n_172), .B(n_147), .Y(n_236) );
AND2x4_ASAP7_75t_L g237 ( .A(n_179), .B(n_152), .Y(n_237) );
INVx1_ASAP7_75t_L g238 ( .A(n_165), .Y(n_238) );
INVxp67_ASAP7_75t_SL g239 ( .A(n_183), .Y(n_239) );
INVx2_ASAP7_75t_L g240 ( .A(n_173), .Y(n_240) );
INVx1_ASAP7_75t_L g241 ( .A(n_193), .Y(n_241) );
AND2x6_ASAP7_75t_L g242 ( .A(n_193), .B(n_148), .Y(n_242) );
INVx3_ASAP7_75t_L g243 ( .A(n_171), .Y(n_243) );
INVx2_ASAP7_75t_L g244 ( .A(n_173), .Y(n_244) );
NAND2xp5_ASAP7_75t_L g245 ( .A(n_198), .B(n_144), .Y(n_245) );
AND2x4_ASAP7_75t_L g246 ( .A(n_179), .B(n_148), .Y(n_246) );
BUFx3_ASAP7_75t_L g247 ( .A(n_184), .Y(n_247) );
NAND2xp5_ASAP7_75t_L g248 ( .A(n_179), .B(n_144), .Y(n_248) );
INVx1_ASAP7_75t_L g249 ( .A(n_193), .Y(n_249) );
BUFx3_ASAP7_75t_L g250 ( .A(n_184), .Y(n_250) );
BUFx2_ASAP7_75t_L g251 ( .A(n_203), .Y(n_251) );
NAND2xp5_ASAP7_75t_SL g252 ( .A(n_179), .B(n_128), .Y(n_252) );
OR2x6_ASAP7_75t_L g253 ( .A(n_203), .B(n_154), .Y(n_253) );
NOR2xp33_ASAP7_75t_R g254 ( .A(n_184), .B(n_150), .Y(n_254) );
INVx1_ASAP7_75t_L g255 ( .A(n_167), .Y(n_255) );
INVx1_ASAP7_75t_L g256 ( .A(n_167), .Y(n_256) );
INVx2_ASAP7_75t_SL g257 ( .A(n_167), .Y(n_257) );
HB1xp67_ASAP7_75t_L g258 ( .A(n_201), .Y(n_258) );
NAND2xp5_ASAP7_75t_SL g259 ( .A(n_167), .B(n_128), .Y(n_259) );
HB1xp67_ASAP7_75t_L g260 ( .A(n_223), .Y(n_260) );
OAI22xp5_ASAP7_75t_L g261 ( .A1(n_216), .A2(n_203), .B1(n_202), .B2(n_160), .Y(n_261) );
NAND2xp5_ASAP7_75t_L g262 ( .A(n_246), .B(n_177), .Y(n_262) );
NOR2xp33_ASAP7_75t_L g263 ( .A(n_209), .B(n_185), .Y(n_263) );
BUFx3_ASAP7_75t_L g264 ( .A(n_224), .Y(n_264) );
INVx1_ASAP7_75t_L g265 ( .A(n_218), .Y(n_265) );
BUFx4f_ASAP7_75t_L g266 ( .A(n_242), .Y(n_266) );
OAI22xp5_ASAP7_75t_L g267 ( .A1(n_216), .A2(n_162), .B1(n_168), .B2(n_190), .Y(n_267) );
NAND2xp33_ASAP7_75t_SL g268 ( .A(n_251), .B(n_187), .Y(n_268) );
BUFx12f_ASAP7_75t_L g269 ( .A(n_221), .Y(n_269) );
AND3x1_ASAP7_75t_SL g270 ( .A(n_221), .B(n_154), .C(n_155), .Y(n_270) );
INVx1_ASAP7_75t_L g271 ( .A(n_255), .Y(n_271) );
NAND2xp5_ASAP7_75t_L g272 ( .A(n_246), .B(n_177), .Y(n_272) );
INVx1_ASAP7_75t_L g273 ( .A(n_218), .Y(n_273) );
BUFx12f_ASAP7_75t_L g274 ( .A(n_253), .Y(n_274) );
AOI222xp33_ASAP7_75t_L g275 ( .A1(n_258), .A2(n_155), .B1(n_157), .B2(n_146), .C1(n_142), .C2(n_129), .Y(n_275) );
INVx1_ASAP7_75t_L g276 ( .A(n_255), .Y(n_276) );
INVx1_ASAP7_75t_SL g277 ( .A(n_219), .Y(n_277) );
CKINVDCx5p33_ASAP7_75t_R g278 ( .A(n_216), .Y(n_278) );
INVx1_ASAP7_75t_L g279 ( .A(n_226), .Y(n_279) );
NAND3xp33_ASAP7_75t_L g280 ( .A(n_235), .B(n_197), .C(n_187), .Y(n_280) );
BUFx6f_ASAP7_75t_L g281 ( .A(n_224), .Y(n_281) );
INVx2_ASAP7_75t_L g282 ( .A(n_208), .Y(n_282) );
AOI22xp5_ASAP7_75t_L g283 ( .A1(n_216), .A2(n_177), .B1(n_197), .B2(n_142), .Y(n_283) );
INVx2_ASAP7_75t_L g284 ( .A(n_208), .Y(n_284) );
NAND2xp5_ASAP7_75t_L g285 ( .A(n_246), .B(n_177), .Y(n_285) );
AOI22xp33_ASAP7_75t_L g286 ( .A1(n_253), .A2(n_177), .B1(n_146), .B2(n_140), .Y(n_286) );
INVx3_ASAP7_75t_L g287 ( .A(n_224), .Y(n_287) );
BUFx3_ASAP7_75t_L g288 ( .A(n_224), .Y(n_288) );
BUFx6f_ASAP7_75t_L g289 ( .A(n_224), .Y(n_289) );
INVx3_ASAP7_75t_L g290 ( .A(n_206), .Y(n_290) );
INVx1_ASAP7_75t_L g291 ( .A(n_228), .Y(n_291) );
OR2x2_ASAP7_75t_L g292 ( .A(n_253), .B(n_129), .Y(n_292) );
INVx2_ASAP7_75t_L g293 ( .A(n_208), .Y(n_293) );
HB1xp67_ASAP7_75t_L g294 ( .A(n_253), .Y(n_294) );
BUFx6f_ASAP7_75t_L g295 ( .A(n_208), .Y(n_295) );
INVx2_ASAP7_75t_L g296 ( .A(n_208), .Y(n_296) );
AOI22xp5_ASAP7_75t_L g297 ( .A1(n_236), .A2(n_177), .B1(n_140), .B2(n_132), .Y(n_297) );
INVx1_ASAP7_75t_L g298 ( .A(n_233), .Y(n_298) );
BUFx2_ASAP7_75t_L g299 ( .A(n_242), .Y(n_299) );
AOI22xp5_ASAP7_75t_L g300 ( .A1(n_236), .A2(n_177), .B1(n_132), .B2(n_122), .Y(n_300) );
BUFx12f_ASAP7_75t_L g301 ( .A(n_251), .Y(n_301) );
INVx2_ASAP7_75t_SL g302 ( .A(n_257), .Y(n_302) );
HB1xp67_ASAP7_75t_L g303 ( .A(n_209), .Y(n_303) );
INVx1_ASAP7_75t_L g304 ( .A(n_238), .Y(n_304) );
INVx5_ASAP7_75t_L g305 ( .A(n_242), .Y(n_305) );
INVx2_ASAP7_75t_L g306 ( .A(n_214), .Y(n_306) );
INVx1_ASAP7_75t_L g307 ( .A(n_256), .Y(n_307) );
CKINVDCx8_ASAP7_75t_R g308 ( .A(n_242), .Y(n_308) );
OAI22xp33_ASAP7_75t_SL g309 ( .A1(n_261), .A2(n_232), .B1(n_225), .B2(n_229), .Y(n_309) );
INVx1_ASAP7_75t_SL g310 ( .A(n_260), .Y(n_310) );
INVx3_ASAP7_75t_L g311 ( .A(n_281), .Y(n_311) );
AND2x2_ASAP7_75t_L g312 ( .A(n_275), .B(n_219), .Y(n_312) );
AOI21xp5_ASAP7_75t_L g313 ( .A1(n_265), .A2(n_222), .B(n_248), .Y(n_313) );
AOI22xp33_ASAP7_75t_L g314 ( .A1(n_274), .A2(n_237), .B1(n_215), .B2(n_242), .Y(n_314) );
OAI21x1_ASAP7_75t_L g315 ( .A1(n_267), .A2(n_149), .B(n_214), .Y(n_315) );
CKINVDCx8_ASAP7_75t_R g316 ( .A(n_305), .Y(n_316) );
BUFx2_ASAP7_75t_L g317 ( .A(n_269), .Y(n_317) );
AOI22xp33_ASAP7_75t_L g318 ( .A1(n_274), .A2(n_237), .B1(n_215), .B2(n_242), .Y(n_318) );
OAI22xp33_ASAP7_75t_L g319 ( .A1(n_278), .A2(n_230), .B1(n_257), .B2(n_227), .Y(n_319) );
HB1xp67_ASAP7_75t_L g320 ( .A(n_277), .Y(n_320) );
INVx4_ASAP7_75t_L g321 ( .A(n_305), .Y(n_321) );
INVx1_ASAP7_75t_L g322 ( .A(n_303), .Y(n_322) );
OAI22xp5_ASAP7_75t_L g323 ( .A1(n_292), .A2(n_237), .B1(n_211), .B2(n_205), .Y(n_323) );
INVx4_ASAP7_75t_L g324 ( .A(n_305), .Y(n_324) );
AND2x4_ASAP7_75t_L g325 ( .A(n_305), .B(n_252), .Y(n_325) );
INVx2_ASAP7_75t_L g326 ( .A(n_306), .Y(n_326) );
INVx1_ASAP7_75t_L g327 ( .A(n_279), .Y(n_327) );
NAND2xp5_ASAP7_75t_L g328 ( .A(n_297), .B(n_220), .Y(n_328) );
OAI21x1_ASAP7_75t_L g329 ( .A1(n_282), .A2(n_149), .B(n_212), .Y(n_329) );
CKINVDCx6p67_ASAP7_75t_R g330 ( .A(n_305), .Y(n_330) );
AOI22xp33_ASAP7_75t_SL g331 ( .A1(n_278), .A2(n_211), .B1(n_254), .B2(n_250), .Y(n_331) );
NAND2xp5_ASAP7_75t_L g332 ( .A(n_300), .B(n_259), .Y(n_332) );
AOI22xp5_ASAP7_75t_L g333 ( .A1(n_292), .A2(n_245), .B1(n_213), .B2(n_239), .Y(n_333) );
OAI22xp5_ASAP7_75t_L g334 ( .A1(n_286), .A2(n_211), .B1(n_207), .B2(n_247), .Y(n_334) );
AND2x4_ASAP7_75t_L g335 ( .A(n_299), .B(n_206), .Y(n_335) );
AOI22xp5_ASAP7_75t_L g336 ( .A1(n_294), .A2(n_270), .B1(n_272), .B2(n_285), .Y(n_336) );
OAI22xp33_ASAP7_75t_SL g337 ( .A1(n_308), .A2(n_250), .B1(n_217), .B2(n_247), .Y(n_337) );
AOI22xp33_ASAP7_75t_SL g338 ( .A1(n_301), .A2(n_217), .B1(n_234), .B2(n_213), .Y(n_338) );
AND2x2_ASAP7_75t_L g339 ( .A(n_299), .B(n_157), .Y(n_339) );
NAND2xp5_ASAP7_75t_L g340 ( .A(n_291), .B(n_231), .Y(n_340) );
OAI22xp33_ASAP7_75t_L g341 ( .A1(n_308), .A2(n_234), .B1(n_206), .B2(n_243), .Y(n_341) );
OAI221xp5_ASAP7_75t_L g342 ( .A1(n_312), .A2(n_263), .B1(n_283), .B2(n_262), .C(n_268), .Y(n_342) );
INVx2_ASAP7_75t_L g343 ( .A(n_326), .Y(n_343) );
AOI22xp33_ASAP7_75t_L g344 ( .A1(n_309), .A2(n_301), .B1(n_268), .B2(n_266), .Y(n_344) );
OAI22x1_ASAP7_75t_L g345 ( .A1(n_310), .A2(n_273), .B1(n_265), .B2(n_234), .Y(n_345) );
OR2x2_ASAP7_75t_L g346 ( .A(n_326), .B(n_306), .Y(n_346) );
OAI211xp5_ASAP7_75t_L g347 ( .A1(n_314), .A2(n_318), .B(n_336), .C(n_320), .Y(n_347) );
AOI22xp33_ASAP7_75t_L g348 ( .A1(n_319), .A2(n_266), .B1(n_273), .B2(n_276), .Y(n_348) );
AOI221xp5_ASAP7_75t_L g349 ( .A1(n_322), .A2(n_307), .B1(n_304), .B2(n_298), .C(n_271), .Y(n_349) );
AOI22xp33_ASAP7_75t_SL g350 ( .A1(n_323), .A2(n_266), .B1(n_234), .B2(n_302), .Y(n_350) );
INVx2_ASAP7_75t_L g351 ( .A(n_329), .Y(n_351) );
BUFx6f_ASAP7_75t_L g352 ( .A(n_316), .Y(n_352) );
OAI22xp33_ASAP7_75t_L g353 ( .A1(n_333), .A2(n_234), .B1(n_302), .B2(n_264), .Y(n_353) );
NAND3xp33_ASAP7_75t_L g354 ( .A(n_313), .B(n_289), .C(n_281), .Y(n_354) );
HB1xp67_ASAP7_75t_L g355 ( .A(n_317), .Y(n_355) );
OAI22xp5_ASAP7_75t_L g356 ( .A1(n_328), .A2(n_295), .B1(n_127), .B2(n_133), .Y(n_356) );
AO31x2_ASAP7_75t_L g357 ( .A1(n_334), .A2(n_127), .A3(n_133), .B(n_143), .Y(n_357) );
AOI22xp33_ASAP7_75t_L g358 ( .A1(n_332), .A2(n_290), .B1(n_249), .B2(n_241), .Y(n_358) );
NAND2xp5_ASAP7_75t_L g359 ( .A(n_327), .B(n_287), .Y(n_359) );
AOI22xp33_ASAP7_75t_L g360 ( .A1(n_339), .A2(n_290), .B1(n_249), .B2(n_241), .Y(n_360) );
AND2x2_ASAP7_75t_L g361 ( .A(n_314), .B(n_290), .Y(n_361) );
AOI221xp5_ASAP7_75t_L g362 ( .A1(n_318), .A2(n_143), .B1(n_125), .B2(n_123), .C(n_280), .Y(n_362) );
A2O1A1Ixp33_ASAP7_75t_L g363 ( .A1(n_340), .A2(n_287), .B(n_288), .C(n_264), .Y(n_363) );
AOI221xp5_ASAP7_75t_SL g364 ( .A1(n_337), .A2(n_123), .B1(n_125), .B2(n_289), .C(n_281), .Y(n_364) );
AO21x1_ASAP7_75t_L g365 ( .A1(n_315), .A2(n_151), .B(n_194), .Y(n_365) );
INVx2_ASAP7_75t_L g366 ( .A(n_329), .Y(n_366) );
BUFx2_ASAP7_75t_L g367 ( .A(n_330), .Y(n_367) );
AND2x2_ASAP7_75t_L g368 ( .A(n_335), .B(n_281), .Y(n_368) );
AO21x2_ASAP7_75t_L g369 ( .A1(n_354), .A2(n_315), .B(n_341), .Y(n_369) );
OAI22xp33_ASAP7_75t_L g370 ( .A1(n_342), .A2(n_330), .B1(n_316), .B2(n_321), .Y(n_370) );
INVx1_ASAP7_75t_L g371 ( .A(n_343), .Y(n_371) );
OAI22xp5_ASAP7_75t_L g372 ( .A1(n_344), .A2(n_338), .B1(n_331), .B2(n_321), .Y(n_372) );
INVx4_ASAP7_75t_L g373 ( .A(n_352), .Y(n_373) );
NAND3xp33_ASAP7_75t_L g374 ( .A(n_364), .B(n_135), .C(n_131), .Y(n_374) );
INVx1_ASAP7_75t_L g375 ( .A(n_343), .Y(n_375) );
AOI211xp5_ASAP7_75t_L g376 ( .A1(n_347), .A2(n_325), .B(n_335), .C(n_151), .Y(n_376) );
OAI221xp5_ASAP7_75t_L g377 ( .A1(n_348), .A2(n_287), .B1(n_288), .B2(n_324), .C(n_321), .Y(n_377) );
HB1xp67_ASAP7_75t_L g378 ( .A(n_355), .Y(n_378) );
INVx2_ASAP7_75t_L g379 ( .A(n_346), .Y(n_379) );
INVx1_ASAP7_75t_L g380 ( .A(n_346), .Y(n_380) );
OAI31xp33_ASAP7_75t_L g381 ( .A1(n_353), .A2(n_325), .A3(n_335), .B(n_243), .Y(n_381) );
INVx2_ASAP7_75t_L g382 ( .A(n_351), .Y(n_382) );
AND2x4_ASAP7_75t_L g383 ( .A(n_361), .B(n_311), .Y(n_383) );
INVx1_ASAP7_75t_L g384 ( .A(n_359), .Y(n_384) );
OAI22xp5_ASAP7_75t_L g385 ( .A1(n_356), .A2(n_324), .B1(n_325), .B2(n_311), .Y(n_385) );
AOI222xp33_ASAP7_75t_L g386 ( .A1(n_349), .A2(n_131), .B1(n_135), .B2(n_289), .C1(n_284), .C2(n_282), .Y(n_386) );
INVx2_ASAP7_75t_L g387 ( .A(n_351), .Y(n_387) );
AOI21xp5_ASAP7_75t_SL g388 ( .A1(n_356), .A2(n_295), .B(n_289), .Y(n_388) );
OAI221xp5_ASAP7_75t_L g389 ( .A1(n_358), .A2(n_289), .B1(n_293), .B2(n_296), .C(n_284), .Y(n_389) );
AND2x2_ASAP7_75t_L g390 ( .A(n_368), .B(n_293), .Y(n_390) );
OAI211xp5_ASAP7_75t_L g391 ( .A1(n_367), .A2(n_131), .B(n_135), .C(n_189), .Y(n_391) );
NAND3xp33_ASAP7_75t_L g392 ( .A(n_364), .B(n_131), .C(n_135), .Y(n_392) );
AND2x2_ASAP7_75t_L g393 ( .A(n_368), .B(n_296), .Y(n_393) );
INVxp67_ASAP7_75t_R g394 ( .A(n_345), .Y(n_394) );
INVx2_ASAP7_75t_L g395 ( .A(n_366), .Y(n_395) );
OAI31xp33_ASAP7_75t_L g396 ( .A1(n_361), .A2(n_243), .A3(n_210), .B(n_186), .Y(n_396) );
AOI22xp33_ASAP7_75t_SL g397 ( .A1(n_367), .A2(n_295), .B1(n_210), .B2(n_135), .Y(n_397) );
OAI332xp33_ASAP7_75t_L g398 ( .A1(n_366), .A2(n_194), .A3(n_189), .B1(n_188), .B2(n_186), .B3(n_174), .C1(n_15), .C2(n_5), .Y(n_398) );
AND2x2_ASAP7_75t_L g399 ( .A(n_383), .B(n_357), .Y(n_399) );
AND2x4_ASAP7_75t_L g400 ( .A(n_383), .B(n_354), .Y(n_400) );
INVx2_ASAP7_75t_L g401 ( .A(n_382), .Y(n_401) );
INVx1_ASAP7_75t_L g402 ( .A(n_371), .Y(n_402) );
INVx3_ASAP7_75t_L g403 ( .A(n_373), .Y(n_403) );
HB1xp67_ASAP7_75t_L g404 ( .A(n_382), .Y(n_404) );
AND2x2_ASAP7_75t_L g405 ( .A(n_383), .B(n_357), .Y(n_405) );
INVx1_ASAP7_75t_SL g406 ( .A(n_378), .Y(n_406) );
OR2x2_ASAP7_75t_L g407 ( .A(n_380), .B(n_357), .Y(n_407) );
OAI221xp5_ASAP7_75t_L g408 ( .A1(n_376), .A2(n_360), .B1(n_362), .B2(n_350), .C(n_363), .Y(n_408) );
INVx1_ASAP7_75t_L g409 ( .A(n_371), .Y(n_409) );
INVx1_ASAP7_75t_SL g410 ( .A(n_373), .Y(n_410) );
NAND3xp33_ASAP7_75t_L g411 ( .A(n_376), .B(n_135), .C(n_352), .Y(n_411) );
INVx1_ASAP7_75t_L g412 ( .A(n_375), .Y(n_412) );
INVx1_ASAP7_75t_L g413 ( .A(n_375), .Y(n_413) );
OR2x2_ASAP7_75t_L g414 ( .A(n_380), .B(n_357), .Y(n_414) );
INVx1_ASAP7_75t_L g415 ( .A(n_387), .Y(n_415) );
NAND2xp5_ASAP7_75t_L g416 ( .A(n_379), .B(n_357), .Y(n_416) );
INVx1_ASAP7_75t_L g417 ( .A(n_387), .Y(n_417) );
INVx2_ASAP7_75t_L g418 ( .A(n_395), .Y(n_418) );
INVx2_ASAP7_75t_L g419 ( .A(n_395), .Y(n_419) );
OAI31xp33_ASAP7_75t_L g420 ( .A1(n_370), .A2(n_374), .A3(n_392), .B(n_372), .Y(n_420) );
AND2x2_ASAP7_75t_L g421 ( .A(n_383), .B(n_379), .Y(n_421) );
INVx3_ASAP7_75t_L g422 ( .A(n_373), .Y(n_422) );
HB1xp67_ASAP7_75t_L g423 ( .A(n_374), .Y(n_423) );
INVx2_ASAP7_75t_L g424 ( .A(n_369), .Y(n_424) );
INVx1_ASAP7_75t_L g425 ( .A(n_384), .Y(n_425) );
AND2x2_ASAP7_75t_L g426 ( .A(n_394), .B(n_365), .Y(n_426) );
INVx1_ASAP7_75t_L g427 ( .A(n_384), .Y(n_427) );
INVx4_ASAP7_75t_L g428 ( .A(n_390), .Y(n_428) );
AND2x2_ASAP7_75t_L g429 ( .A(n_390), .B(n_345), .Y(n_429) );
OAI22xp5_ASAP7_75t_L g430 ( .A1(n_392), .A2(n_352), .B1(n_295), .B2(n_365), .Y(n_430) );
NAND2xp5_ASAP7_75t_L g431 ( .A(n_393), .B(n_352), .Y(n_431) );
NAND2xp5_ASAP7_75t_SL g432 ( .A(n_386), .B(n_352), .Y(n_432) );
AND2x2_ASAP7_75t_L g433 ( .A(n_393), .B(n_6), .Y(n_433) );
INVx2_ASAP7_75t_L g434 ( .A(n_369), .Y(n_434) );
AND2x2_ASAP7_75t_L g435 ( .A(n_394), .B(n_6), .Y(n_435) );
BUFx3_ASAP7_75t_L g436 ( .A(n_377), .Y(n_436) );
NAND2xp5_ASAP7_75t_L g437 ( .A(n_385), .B(n_295), .Y(n_437) );
INVx3_ASAP7_75t_L g438 ( .A(n_369), .Y(n_438) );
AOI221xp5_ASAP7_75t_L g439 ( .A1(n_398), .A2(n_188), .B1(n_174), .B2(n_204), .C(n_196), .Y(n_439) );
INVx2_ASAP7_75t_SL g440 ( .A(n_388), .Y(n_440) );
AND2x2_ASAP7_75t_L g441 ( .A(n_388), .B(n_8), .Y(n_441) );
AOI33xp33_ASAP7_75t_L g442 ( .A1(n_397), .A2(n_196), .A3(n_195), .B1(n_204), .B2(n_16), .B3(n_17), .Y(n_442) );
INVx1_ASAP7_75t_SL g443 ( .A(n_406), .Y(n_443) );
AND2x2_ASAP7_75t_L g444 ( .A(n_428), .B(n_9), .Y(n_444) );
INVx1_ASAP7_75t_L g445 ( .A(n_425), .Y(n_445) );
AND2x2_ASAP7_75t_L g446 ( .A(n_421), .B(n_13), .Y(n_446) );
OAI33xp33_ASAP7_75t_L g447 ( .A1(n_427), .A2(n_13), .A3(n_15), .B1(n_16), .B2(n_200), .B3(n_191), .Y(n_447) );
AOI22xp33_ASAP7_75t_L g448 ( .A1(n_439), .A2(n_381), .B1(n_396), .B2(n_389), .Y(n_448) );
HB1xp67_ASAP7_75t_L g449 ( .A(n_410), .Y(n_449) );
NAND2xp5_ASAP7_75t_L g450 ( .A(n_427), .B(n_391), .Y(n_450) );
INVx1_ASAP7_75t_SL g451 ( .A(n_410), .Y(n_451) );
HB1xp67_ASAP7_75t_L g452 ( .A(n_404), .Y(n_452) );
AO21x2_ASAP7_75t_L g453 ( .A1(n_441), .A2(n_430), .B(n_424), .Y(n_453) );
AND2x2_ASAP7_75t_L g454 ( .A(n_421), .B(n_19), .Y(n_454) );
NAND2xp5_ASAP7_75t_L g455 ( .A(n_433), .B(n_21), .Y(n_455) );
INVx1_ASAP7_75t_L g456 ( .A(n_402), .Y(n_456) );
INVx1_ASAP7_75t_L g457 ( .A(n_402), .Y(n_457) );
NAND2xp5_ASAP7_75t_SL g458 ( .A(n_420), .B(n_166), .Y(n_458) );
NOR3xp33_ASAP7_75t_SL g459 ( .A(n_411), .B(n_195), .C(n_26), .Y(n_459) );
NOR2xp67_ASAP7_75t_L g460 ( .A(n_411), .B(n_23), .Y(n_460) );
INVx1_ASAP7_75t_L g461 ( .A(n_409), .Y(n_461) );
BUFx2_ASAP7_75t_L g462 ( .A(n_428), .Y(n_462) );
AND2x4_ASAP7_75t_L g463 ( .A(n_399), .B(n_28), .Y(n_463) );
INVx1_ASAP7_75t_L g464 ( .A(n_412), .Y(n_464) );
INVx2_ASAP7_75t_SL g465 ( .A(n_403), .Y(n_465) );
INVx1_ASAP7_75t_L g466 ( .A(n_412), .Y(n_466) );
INVxp67_ASAP7_75t_SL g467 ( .A(n_404), .Y(n_467) );
OR2x2_ASAP7_75t_L g468 ( .A(n_428), .B(n_30), .Y(n_468) );
INVx1_ASAP7_75t_L g469 ( .A(n_413), .Y(n_469) );
NAND2xp5_ASAP7_75t_L g470 ( .A(n_433), .B(n_31), .Y(n_470) );
AND2x2_ASAP7_75t_L g471 ( .A(n_399), .B(n_33), .Y(n_471) );
OR2x2_ASAP7_75t_L g472 ( .A(n_428), .B(n_35), .Y(n_472) );
AND2x2_ASAP7_75t_L g473 ( .A(n_399), .B(n_39), .Y(n_473) );
INVxp67_ASAP7_75t_L g474 ( .A(n_441), .Y(n_474) );
AOI22xp5_ASAP7_75t_L g475 ( .A1(n_439), .A2(n_210), .B1(n_244), .B2(n_240), .Y(n_475) );
INVx2_ASAP7_75t_SL g476 ( .A(n_403), .Y(n_476) );
AND2x2_ASAP7_75t_L g477 ( .A(n_405), .B(n_40), .Y(n_477) );
HB1xp67_ASAP7_75t_L g478 ( .A(n_403), .Y(n_478) );
NAND3xp33_ASAP7_75t_L g479 ( .A(n_441), .B(n_166), .C(n_178), .Y(n_479) );
AOI22xp33_ASAP7_75t_L g480 ( .A1(n_436), .A2(n_166), .B1(n_178), .B2(n_200), .Y(n_480) );
OR2x2_ASAP7_75t_L g481 ( .A(n_431), .B(n_41), .Y(n_481) );
NOR2xp33_ASAP7_75t_L g482 ( .A(n_435), .B(n_42), .Y(n_482) );
OR2x2_ASAP7_75t_L g483 ( .A(n_431), .B(n_44), .Y(n_483) );
NAND2xp5_ASAP7_75t_SL g484 ( .A(n_420), .B(n_166), .Y(n_484) );
OR2x2_ASAP7_75t_L g485 ( .A(n_407), .B(n_46), .Y(n_485) );
O2A1O1Ixp5_ASAP7_75t_L g486 ( .A1(n_432), .A2(n_191), .B(n_182), .C(n_180), .Y(n_486) );
INVx1_ASAP7_75t_SL g487 ( .A(n_403), .Y(n_487) );
NAND2xp5_ASAP7_75t_L g488 ( .A(n_435), .B(n_48), .Y(n_488) );
INVx3_ASAP7_75t_L g489 ( .A(n_422), .Y(n_489) );
NAND3xp33_ASAP7_75t_SL g490 ( .A(n_442), .B(n_182), .C(n_180), .Y(n_490) );
INVx2_ASAP7_75t_SL g491 ( .A(n_422), .Y(n_491) );
NAND2xp5_ASAP7_75t_L g492 ( .A(n_443), .B(n_414), .Y(n_492) );
OAI21xp5_ASAP7_75t_L g493 ( .A1(n_460), .A2(n_423), .B(n_430), .Y(n_493) );
INVxp67_ASAP7_75t_L g494 ( .A(n_449), .Y(n_494) );
NOR2xp33_ASAP7_75t_L g495 ( .A(n_474), .B(n_422), .Y(n_495) );
NAND4xp25_ASAP7_75t_L g496 ( .A(n_482), .B(n_436), .C(n_426), .D(n_408), .Y(n_496) );
AOI322xp5_ASAP7_75t_L g497 ( .A1(n_444), .A2(n_426), .A3(n_405), .B1(n_429), .B2(n_423), .C1(n_436), .C2(n_440), .Y(n_497) );
AND2x2_ASAP7_75t_L g498 ( .A(n_462), .B(n_451), .Y(n_498) );
NAND2xp5_ASAP7_75t_L g499 ( .A(n_445), .B(n_414), .Y(n_499) );
INVx2_ASAP7_75t_SL g500 ( .A(n_465), .Y(n_500) );
OAI31xp33_ASAP7_75t_L g501 ( .A1(n_482), .A2(n_408), .A3(n_426), .B(n_440), .Y(n_501) );
INVx1_ASAP7_75t_L g502 ( .A(n_456), .Y(n_502) );
NAND2xp5_ASAP7_75t_L g503 ( .A(n_446), .B(n_416), .Y(n_503) );
NAND2xp5_ASAP7_75t_L g504 ( .A(n_446), .B(n_416), .Y(n_504) );
INVx1_ASAP7_75t_L g505 ( .A(n_457), .Y(n_505) );
INVx1_ASAP7_75t_L g506 ( .A(n_461), .Y(n_506) );
AOI22xp5_ASAP7_75t_SL g507 ( .A1(n_463), .A2(n_422), .B1(n_440), .B2(n_400), .Y(n_507) );
INVx1_ASAP7_75t_SL g508 ( .A(n_487), .Y(n_508) );
NAND2xp5_ASAP7_75t_L g509 ( .A(n_464), .B(n_415), .Y(n_509) );
AND3x2_ASAP7_75t_L g510 ( .A(n_478), .B(n_400), .C(n_415), .Y(n_510) );
NOR2xp33_ASAP7_75t_L g511 ( .A(n_488), .B(n_400), .Y(n_511) );
NAND2xp5_ASAP7_75t_L g512 ( .A(n_466), .B(n_417), .Y(n_512) );
A2O1A1Ixp33_ASAP7_75t_L g513 ( .A1(n_459), .A2(n_400), .B(n_417), .C(n_437), .Y(n_513) );
CKINVDCx20_ASAP7_75t_R g514 ( .A(n_477), .Y(n_514) );
OR2x2_ASAP7_75t_L g515 ( .A(n_452), .B(n_419), .Y(n_515) );
INVx1_ASAP7_75t_SL g516 ( .A(n_489), .Y(n_516) );
NAND2xp5_ASAP7_75t_L g517 ( .A(n_469), .B(n_419), .Y(n_517) );
INVx1_ASAP7_75t_L g518 ( .A(n_467), .Y(n_518) );
INVx3_ASAP7_75t_SL g519 ( .A(n_468), .Y(n_519) );
OR2x2_ASAP7_75t_L g520 ( .A(n_465), .B(n_418), .Y(n_520) );
OR2x2_ASAP7_75t_L g521 ( .A(n_476), .B(n_401), .Y(n_521) );
AND2x2_ASAP7_75t_L g522 ( .A(n_471), .B(n_438), .Y(n_522) );
NAND2xp5_ASAP7_75t_L g523 ( .A(n_473), .B(n_434), .Y(n_523) );
NAND4xp25_ASAP7_75t_L g524 ( .A(n_448), .B(n_438), .C(n_434), .D(n_424), .Y(n_524) );
INVx1_ASAP7_75t_SL g525 ( .A(n_489), .Y(n_525) );
INVxp67_ASAP7_75t_L g526 ( .A(n_476), .Y(n_526) );
INVx1_ASAP7_75t_SL g527 ( .A(n_489), .Y(n_527) );
OAI21xp33_ASAP7_75t_L g528 ( .A1(n_458), .A2(n_438), .B(n_434), .Y(n_528) );
NAND3xp33_ASAP7_75t_L g529 ( .A(n_479), .B(n_438), .C(n_424), .Y(n_529) );
AND2x2_ASAP7_75t_L g530 ( .A(n_477), .B(n_49), .Y(n_530) );
INVx2_ASAP7_75t_L g531 ( .A(n_491), .Y(n_531) );
AND2x6_ASAP7_75t_L g532 ( .A(n_463), .B(n_50), .Y(n_532) );
INVx1_ASAP7_75t_L g533 ( .A(n_450), .Y(n_533) );
INVx2_ASAP7_75t_L g534 ( .A(n_491), .Y(n_534) );
AND2x2_ASAP7_75t_L g535 ( .A(n_463), .B(n_52), .Y(n_535) );
INVx1_ASAP7_75t_L g536 ( .A(n_485), .Y(n_536) );
AND2x2_ASAP7_75t_L g537 ( .A(n_522), .B(n_453), .Y(n_537) );
OAI21xp5_ASAP7_75t_L g538 ( .A1(n_501), .A2(n_458), .B(n_484), .Y(n_538) );
INVx1_ASAP7_75t_L g539 ( .A(n_502), .Y(n_539) );
INVxp67_ASAP7_75t_SL g540 ( .A(n_494), .Y(n_540) );
INVx1_ASAP7_75t_SL g541 ( .A(n_498), .Y(n_541) );
NAND2xp5_ASAP7_75t_L g542 ( .A(n_533), .B(n_453), .Y(n_542) );
INVx1_ASAP7_75t_L g543 ( .A(n_505), .Y(n_543) );
INVx2_ASAP7_75t_SL g544 ( .A(n_508), .Y(n_544) );
INVx1_ASAP7_75t_L g545 ( .A(n_506), .Y(n_545) );
HB1xp67_ASAP7_75t_L g546 ( .A(n_508), .Y(n_546) );
INVx1_ASAP7_75t_SL g547 ( .A(n_514), .Y(n_547) );
INVx1_ASAP7_75t_SL g548 ( .A(n_519), .Y(n_548) );
NAND2xp5_ASAP7_75t_SL g549 ( .A(n_507), .B(n_472), .Y(n_549) );
INVx1_ASAP7_75t_SL g550 ( .A(n_492), .Y(n_550) );
NAND2x1p5_ASAP7_75t_L g551 ( .A(n_535), .B(n_454), .Y(n_551) );
NAND2xp5_ASAP7_75t_L g552 ( .A(n_518), .B(n_499), .Y(n_552) );
INVx1_ASAP7_75t_L g553 ( .A(n_509), .Y(n_553) );
NAND2xp5_ASAP7_75t_L g554 ( .A(n_499), .B(n_483), .Y(n_554) );
INVx1_ASAP7_75t_L g555 ( .A(n_512), .Y(n_555) );
AOI21xp33_ASAP7_75t_L g556 ( .A1(n_495), .A2(n_470), .B(n_455), .Y(n_556) );
INVx3_ASAP7_75t_L g557 ( .A(n_510), .Y(n_557) );
AOI211xp5_ASAP7_75t_L g558 ( .A1(n_496), .A2(n_447), .B(n_481), .C(n_475), .Y(n_558) );
INVx1_ASAP7_75t_L g559 ( .A(n_517), .Y(n_559) );
AND2x4_ASAP7_75t_L g560 ( .A(n_500), .B(n_480), .Y(n_560) );
INVx1_ASAP7_75t_L g561 ( .A(n_515), .Y(n_561) );
INVxp67_ASAP7_75t_L g562 ( .A(n_531), .Y(n_562) );
INVx1_ASAP7_75t_L g563 ( .A(n_520), .Y(n_563) );
INVx2_ASAP7_75t_SL g564 ( .A(n_521), .Y(n_564) );
NOR2x1_ASAP7_75t_L g565 ( .A(n_493), .B(n_490), .Y(n_565) );
AOI221xp5_ASAP7_75t_L g566 ( .A1(n_496), .A2(n_448), .B1(n_486), .B2(n_161), .C(n_176), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g567 ( .A(n_503), .B(n_54), .Y(n_567) );
OR2x2_ASAP7_75t_L g568 ( .A(n_504), .B(n_176), .Y(n_568) );
INVx2_ASAP7_75t_SL g569 ( .A(n_534), .Y(n_569) );
NAND2xp5_ASAP7_75t_SL g570 ( .A(n_493), .B(n_178), .Y(n_570) );
INVx1_ASAP7_75t_L g571 ( .A(n_526), .Y(n_571) );
NAND2xp5_ASAP7_75t_L g572 ( .A(n_497), .B(n_55), .Y(n_572) );
NAND3xp33_ASAP7_75t_L g573 ( .A(n_524), .B(n_178), .C(n_166), .Y(n_573) );
AOI21xp5_ASAP7_75t_L g574 ( .A1(n_528), .A2(n_513), .B(n_524), .Y(n_574) );
OAI21xp5_ASAP7_75t_L g575 ( .A1(n_532), .A2(n_58), .B(n_59), .Y(n_575) );
HB1xp67_ASAP7_75t_L g576 ( .A(n_516), .Y(n_576) );
AND4x1_ASAP7_75t_SL g577 ( .A(n_532), .B(n_60), .C(n_61), .D(n_62), .Y(n_577) );
INVx2_ASAP7_75t_SL g578 ( .A(n_532), .Y(n_578) );
AND2x2_ASAP7_75t_L g579 ( .A(n_511), .B(n_63), .Y(n_579) );
INVx1_ASAP7_75t_L g580 ( .A(n_536), .Y(n_580) );
NAND3xp33_ASAP7_75t_L g581 ( .A(n_529), .B(n_64), .C(n_66), .Y(n_581) );
NAND2xp33_ASAP7_75t_SL g582 ( .A(n_530), .B(n_68), .Y(n_582) );
INVx1_ASAP7_75t_L g583 ( .A(n_523), .Y(n_583) );
OAI211xp5_ASAP7_75t_SL g584 ( .A1(n_516), .A2(n_73), .B(n_74), .C(n_75), .Y(n_584) );
AOI22xp5_ASAP7_75t_L g585 ( .A1(n_532), .A2(n_496), .B1(n_474), .B2(n_514), .Y(n_585) );
INVxp67_ASAP7_75t_SL g586 ( .A(n_525), .Y(n_586) );
AOI221xp5_ASAP7_75t_L g587 ( .A1(n_527), .A2(n_533), .B1(n_496), .B2(n_524), .C(n_406), .Y(n_587) );
OA22x2_ASAP7_75t_L g588 ( .A1(n_510), .A2(n_519), .B1(n_462), .B2(n_443), .Y(n_588) );
OAI22xp5_ASAP7_75t_SL g589 ( .A1(n_514), .A2(n_519), .B1(n_462), .B2(n_474), .Y(n_589) );
CKINVDCx5p33_ASAP7_75t_R g590 ( .A(n_514), .Y(n_590) );
INVx1_ASAP7_75t_L g591 ( .A(n_502), .Y(n_591) );
AOI21xp33_ASAP7_75t_SL g592 ( .A1(n_519), .A2(n_501), .B(n_411), .Y(n_592) );
INVx1_ASAP7_75t_L g593 ( .A(n_502), .Y(n_593) );
BUFx6f_ASAP7_75t_L g594 ( .A(n_568), .Y(n_594) );
OAI21xp5_ASAP7_75t_L g595 ( .A1(n_565), .A2(n_538), .B(n_592), .Y(n_595) );
INVx1_ASAP7_75t_L g596 ( .A(n_552), .Y(n_596) );
OAI221xp5_ASAP7_75t_SL g597 ( .A1(n_585), .A2(n_587), .B1(n_548), .B2(n_574), .C(n_547), .Y(n_597) );
NOR3xp33_ASAP7_75t_L g598 ( .A(n_572), .B(n_577), .C(n_549), .Y(n_598) );
OAI321xp33_ASAP7_75t_L g599 ( .A1(n_549), .A2(n_589), .A3(n_578), .B1(n_542), .B2(n_575), .C(n_551), .Y(n_599) );
AND2x2_ASAP7_75t_L g600 ( .A(n_537), .B(n_546), .Y(n_600) );
NOR4xp25_ASAP7_75t_L g601 ( .A(n_540), .B(n_580), .C(n_570), .D(n_571), .Y(n_601) );
OAI221xp5_ASAP7_75t_L g602 ( .A1(n_588), .A2(n_558), .B1(n_557), .B2(n_582), .C(n_551), .Y(n_602) );
NAND4xp25_ASAP7_75t_L g603 ( .A(n_556), .B(n_573), .C(n_582), .D(n_570), .Y(n_603) );
AND2x2_ASAP7_75t_L g604 ( .A(n_537), .B(n_546), .Y(n_604) );
INVx1_ASAP7_75t_L g605 ( .A(n_559), .Y(n_605) );
HB1xp67_ASAP7_75t_L g606 ( .A(n_544), .Y(n_606) );
NAND4xp75_ASAP7_75t_L g607 ( .A(n_579), .B(n_567), .C(n_544), .D(n_566), .Y(n_607) );
AOI21xp5_ASAP7_75t_L g608 ( .A1(n_588), .A2(n_557), .B(n_590), .Y(n_608) );
AND2x2_ASAP7_75t_L g609 ( .A(n_608), .B(n_541), .Y(n_609) );
AOI221xp5_ASAP7_75t_L g610 ( .A1(n_595), .A2(n_555), .B1(n_553), .B2(n_550), .C(n_583), .Y(n_610) );
O2A1O1Ixp33_ASAP7_75t_L g611 ( .A1(n_597), .A2(n_584), .B(n_557), .C(n_576), .Y(n_611) );
NOR2x1_ASAP7_75t_SL g612 ( .A(n_594), .B(n_569), .Y(n_612) );
INVx2_ASAP7_75t_SL g613 ( .A(n_606), .Y(n_613) );
XOR2xp5_ASAP7_75t_L g614 ( .A(n_607), .B(n_554), .Y(n_614) );
AOI221xp5_ASAP7_75t_L g615 ( .A1(n_599), .A2(n_563), .B1(n_593), .B2(n_539), .C(n_545), .Y(n_615) );
NOR2x1_ASAP7_75t_L g616 ( .A(n_602), .B(n_581), .Y(n_616) );
INVx2_ASAP7_75t_SL g617 ( .A(n_594), .Y(n_617) );
AOI22xp33_ASAP7_75t_SL g618 ( .A1(n_609), .A2(n_600), .B1(n_604), .B2(n_594), .Y(n_618) );
NAND4xp25_ASAP7_75t_L g619 ( .A(n_616), .B(n_598), .C(n_603), .D(n_604), .Y(n_619) );
OAI222xp33_ASAP7_75t_L g620 ( .A1(n_614), .A2(n_600), .B1(n_596), .B2(n_605), .C1(n_564), .C2(n_562), .Y(n_620) );
OR5x1_ASAP7_75t_L g621 ( .A(n_615), .B(n_601), .C(n_607), .D(n_594), .E(n_586), .Y(n_621) );
OAI22xp33_ASAP7_75t_SL g622 ( .A1(n_613), .A2(n_586), .B1(n_564), .B2(n_576), .Y(n_622) );
NAND3xp33_ASAP7_75t_L g623 ( .A(n_619), .B(n_611), .C(n_610), .Y(n_623) );
OAI22xp5_ASAP7_75t_L g624 ( .A1(n_618), .A2(n_617), .B1(n_612), .B2(n_561), .Y(n_624) );
AOI22xp5_ASAP7_75t_L g625 ( .A1(n_622), .A2(n_560), .B1(n_591), .B2(n_543), .Y(n_625) );
INVx1_ASAP7_75t_L g626 ( .A(n_625), .Y(n_626) );
INVx1_ASAP7_75t_L g627 ( .A(n_623), .Y(n_627) );
INVxp67_ASAP7_75t_SL g628 ( .A(n_627), .Y(n_628) );
INVx2_ASAP7_75t_L g629 ( .A(n_626), .Y(n_629) );
OAI21xp5_ASAP7_75t_L g630 ( .A1(n_628), .A2(n_624), .B(n_620), .Y(n_630) );
XNOR2xp5_ASAP7_75t_L g631 ( .A(n_630), .B(n_629), .Y(n_631) );
OAI21xp5_ASAP7_75t_L g632 ( .A1(n_631), .A2(n_621), .B(n_568), .Y(n_632) );
endmodule