module fake_jpeg_1066_n_189 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_189);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_189;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_186;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx3_ASAP7_75t_L g42 ( 
.A(n_11),
.Y(n_42)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_25),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_34),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_1),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_19),
.Y(n_46)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_41),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_20),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_36),
.Y(n_49)
);

INVx1_ASAP7_75t_SL g50 ( 
.A(n_11),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_29),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_5),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_0),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_28),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_37),
.Y(n_55)
);

BUFx12_ASAP7_75t_L g56 ( 
.A(n_23),
.Y(n_56)
);

CKINVDCx16_ASAP7_75t_R g57 ( 
.A(n_9),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_15),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_26),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_16),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_24),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_33),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_47),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_63),
.Y(n_74)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_42),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_64),
.Y(n_79)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_44),
.Y(n_65)
);

INVx3_ASAP7_75t_SL g80 ( 
.A(n_65),
.Y(n_80)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_43),
.Y(n_66)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_66),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_53),
.B(n_0),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_67),
.B(n_57),
.Y(n_83)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_42),
.Y(n_68)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_68),
.Y(n_76)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_45),
.Y(n_69)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_69),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_47),
.Y(n_70)
);

NAND2xp33_ASAP7_75t_SL g78 ( 
.A(n_70),
.B(n_52),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_64),
.B(n_45),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_71),
.B(n_75),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_68),
.A2(n_52),
.B1(n_47),
.B2(n_50),
.Y(n_72)
);

AOI21xp5_ASAP7_75t_L g93 ( 
.A1(n_72),
.A2(n_59),
.B(n_55),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_63),
.B(n_58),
.Y(n_75)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_70),
.B(n_50),
.Y(n_77)
);

OR2x2_ASAP7_75t_L g102 ( 
.A(n_77),
.B(n_54),
.Y(n_102)
);

AND2x2_ASAP7_75t_L g98 ( 
.A(n_78),
.B(n_83),
.Y(n_98)
);

BUFx16f_ASAP7_75t_L g82 ( 
.A(n_65),
.Y(n_82)
);

BUFx3_ASAP7_75t_L g90 ( 
.A(n_82),
.Y(n_90)
);

AO22x2_ASAP7_75t_SL g84 ( 
.A1(n_66),
.A2(n_62),
.B1(n_48),
.B2(n_51),
.Y(n_84)
);

O2A1O1Ixp33_ASAP7_75t_L g91 ( 
.A1(n_84),
.A2(n_61),
.B(n_62),
.C(n_51),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_82),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_85),
.B(n_100),
.Y(n_109)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_76),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_86),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_L g87 ( 
.A1(n_73),
.A2(n_60),
.B1(n_43),
.B2(n_61),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_87),
.A2(n_93),
.B1(n_49),
.B2(n_46),
.Y(n_107)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_81),
.Y(n_88)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_88),
.Y(n_112)
);

XNOR2xp5_ASAP7_75t_SL g89 ( 
.A(n_77),
.B(n_48),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_89),
.B(n_92),
.C(n_56),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_L g115 ( 
.A1(n_91),
.A2(n_84),
.B(n_56),
.Y(n_115)
);

XNOR2xp5_ASAP7_75t_L g92 ( 
.A(n_80),
.B(n_54),
.Y(n_92)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_76),
.Y(n_95)
);

AND2x2_ASAP7_75t_L g113 ( 
.A(n_95),
.B(n_96),
.Y(n_113)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_79),
.Y(n_96)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_80),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_97),
.B(n_72),
.Y(n_106)
);

BUFx3_ASAP7_75t_L g99 ( 
.A(n_79),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_99),
.B(n_101),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_74),
.Y(n_100)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_74),
.Y(n_101)
);

AND2x2_ASAP7_75t_L g122 ( 
.A(n_102),
.B(n_4),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_91),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_103),
.B(n_106),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_98),
.A2(n_94),
.B1(n_96),
.B2(n_99),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_SL g125 ( 
.A1(n_105),
.A2(n_5),
.B(n_6),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_107),
.B(n_108),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_102),
.B(n_84),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_90),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_110),
.B(n_114),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_SL g111 ( 
.A(n_98),
.B(n_1),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_111),
.B(n_116),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_90),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_115),
.B(n_118),
.Y(n_144)
);

A2O1A1Ixp33_ASAP7_75t_L g118 ( 
.A1(n_87),
.A2(n_2),
.B(n_3),
.C(n_4),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_102),
.B(n_2),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_119),
.B(n_120),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_102),
.B(n_3),
.Y(n_120)
);

XNOR2xp5_ASAP7_75t_L g121 ( 
.A(n_89),
.B(n_56),
.Y(n_121)
);

XNOR2xp5_ASAP7_75t_L g129 ( 
.A(n_121),
.B(n_6),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_122),
.B(n_7),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_104),
.A2(n_22),
.B1(n_39),
.B2(n_38),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_SL g150 ( 
.A1(n_123),
.A2(n_125),
.B(n_128),
.Y(n_150)
);

HB1xp67_ASAP7_75t_L g124 ( 
.A(n_117),
.Y(n_124)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_124),
.Y(n_146)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_109),
.Y(n_127)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_127),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_113),
.A2(n_21),
.B1(n_35),
.B2(n_32),
.Y(n_128)
);

XOR2xp5_ASAP7_75t_L g147 ( 
.A(n_129),
.B(n_10),
.Y(n_147)
);

BUFx24_ASAP7_75t_SL g130 ( 
.A(n_122),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_130),
.B(n_134),
.Y(n_155)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_112),
.Y(n_133)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_133),
.Y(n_152)
);

XNOR2xp5_ASAP7_75t_L g135 ( 
.A(n_121),
.B(n_18),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_135),
.B(n_12),
.C(n_13),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_116),
.B(n_7),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_136),
.B(n_137),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_113),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_107),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_140),
.A2(n_12),
.B1(n_13),
.B2(n_14),
.Y(n_148)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_117),
.Y(n_141)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_141),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_105),
.B(n_8),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_142),
.B(n_14),
.Y(n_159)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_118),
.Y(n_143)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_143),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_147),
.B(n_162),
.C(n_149),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_148),
.B(n_151),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_SL g164 ( 
.A(n_149),
.B(n_160),
.Y(n_164)
);

O2A1O1Ixp33_ASAP7_75t_L g151 ( 
.A1(n_126),
.A2(n_27),
.B(n_31),
.C(n_30),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_139),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_153),
.B(n_159),
.Y(n_169)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_144),
.Y(n_158)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_158),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_131),
.B(n_15),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_125),
.B(n_16),
.Y(n_161)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_161),
.Y(n_171)
);

XOR2xp5_ASAP7_75t_L g162 ( 
.A(n_129),
.B(n_40),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_163),
.B(n_165),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_156),
.B(n_135),
.C(n_138),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_145),
.A2(n_132),
.B1(n_140),
.B2(n_123),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g173 ( 
.A1(n_166),
.A2(n_157),
.B1(n_146),
.B2(n_148),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_152),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_167),
.B(n_155),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_L g172 ( 
.A1(n_168),
.A2(n_151),
.B(n_150),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_172),
.B(n_177),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_173),
.A2(n_175),
.B1(n_171),
.B2(n_169),
.Y(n_179)
);

FAx1_ASAP7_75t_SL g174 ( 
.A(n_165),
.B(n_150),
.CI(n_147),
.CON(n_174),
.SN(n_174)
);

NOR2xp33_ASAP7_75t_SL g181 ( 
.A(n_174),
.B(n_164),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_170),
.A2(n_146),
.B1(n_154),
.B2(n_162),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_L g178 ( 
.A(n_176),
.B(n_163),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g182 ( 
.A(n_178),
.B(n_181),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_179),
.B(n_175),
.Y(n_183)
);

XOR2xp5_ASAP7_75t_L g184 ( 
.A(n_183),
.B(n_180),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_184),
.B(n_182),
.Y(n_185)
);

AOI21xp5_ASAP7_75t_L g186 ( 
.A1(n_185),
.A2(n_178),
.B(n_172),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g187 ( 
.A(n_186),
.B(n_174),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_187),
.B(n_128),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_L g189 ( 
.A(n_188),
.B(n_17),
.Y(n_189)
);


endmodule