module real_jpeg_2140_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_166;
wire n_176;
wire n_221;
wire n_215;
wire n_104;
wire n_194;
wire n_153;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_227;
wire n_126;
wire n_214;
wire n_13;
wire n_120;
wire n_113;
wire n_155;
wire n_199;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_136;
wire n_44;
wire n_28;
wire n_208;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_203;
wire n_192;
wire n_100;
wire n_198;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_195;
wire n_110;
wire n_205;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_103;
wire n_225;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_185;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_167;
wire n_213;
wire n_179;
wire n_202;
wire n_216;
wire n_133;
wire n_138;
wire n_25;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;
wire n_16;

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_0),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_1),
.A2(n_64),
.B1(n_65),
.B2(n_68),
.Y(n_63)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_1),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_1),
.A2(n_25),
.B1(n_26),
.B2(n_68),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g30 ( 
.A1(n_2),
.A2(n_31),
.B1(n_33),
.B2(n_34),
.Y(n_30)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_2),
.Y(n_33)
);

MAJIxp5_ASAP7_75t_L g59 ( 
.A(n_2),
.B(n_31),
.C(n_46),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_2),
.A2(n_25),
.B1(n_26),
.B2(n_33),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_2),
.A2(n_33),
.B1(n_48),
.B2(n_50),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_2),
.A2(n_33),
.B1(n_64),
.B2(n_65),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_2),
.B(n_44),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_2),
.B(n_24),
.C(n_26),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_2),
.B(n_65),
.C(n_82),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_2),
.B(n_22),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_2),
.B(n_62),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_2),
.B(n_164),
.Y(n_217)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_3),
.Y(n_62)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

OAI22xp33_ASAP7_75t_SL g38 ( 
.A1(n_5),
.A2(n_31),
.B1(n_34),
.B2(n_39),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_5),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_SL g54 ( 
.A1(n_5),
.A2(n_39),
.B1(n_48),
.B2(n_50),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_5),
.A2(n_25),
.B1(n_26),
.B2(n_39),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_5),
.A2(n_39),
.B1(n_64),
.B2(n_65),
.Y(n_195)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_6),
.Y(n_48)
);

BUFx16f_ASAP7_75t_L g83 ( 
.A(n_7),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_8),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_SL g47 ( 
.A1(n_9),
.A2(n_48),
.B1(n_49),
.B2(n_50),
.Y(n_47)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_9),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_L g70 ( 
.A1(n_9),
.A2(n_49),
.B1(n_64),
.B2(n_65),
.Y(n_70)
);

OAI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_9),
.A2(n_25),
.B1(n_26),
.B2(n_49),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_L g101 ( 
.A1(n_9),
.A2(n_31),
.B1(n_34),
.B2(n_49),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_10),
.Y(n_46)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

XOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_127),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_126),
.Y(n_13)
);

INVxp67_ASAP7_75t_L g14 ( 
.A(n_15),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_104),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_16),
.B(n_104),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_72),
.C(n_87),
.Y(n_16)
);

XNOR2xp5_ASAP7_75t_L g145 ( 
.A(n_17),
.B(n_146),
.Y(n_145)
);

XOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_56),
.Y(n_17)
);

AOI22xp5_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_20),
.B1(n_42),
.B2(n_55),
.Y(n_18)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_19),
.B(n_55),
.C(n_56),
.Y(n_105)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_35),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_30),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_22),
.B(n_38),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_L g113 ( 
.A1(n_22),
.A2(n_30),
.B(n_114),
.Y(n_113)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_23),
.B(n_41),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_23),
.B(n_101),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_25),
.B1(n_26),
.B2(n_29),
.Y(n_23)
);

INVx3_ASAP7_75t_SL g29 ( 
.A(n_24),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_L g41 ( 
.A1(n_24),
.A2(n_29),
.B1(n_31),
.B2(n_34),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_25),
.A2(n_26),
.B1(n_81),
.B2(n_82),
.Y(n_80)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_26),
.B(n_189),
.Y(n_188)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_SL g180 ( 
.A(n_30),
.B(n_114),
.Y(n_180)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_31),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_SL g44 ( 
.A1(n_31),
.A2(n_34),
.B1(n_45),
.B2(n_46),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_31),
.B(n_159),
.Y(n_158)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVxp67_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_36),
.B(n_139),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_37),
.B(n_40),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_SL g100 ( 
.A(n_40),
.B(n_101),
.Y(n_100)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_40),
.Y(n_114)
);

CKINVDCx14_ASAP7_75t_R g55 ( 
.A(n_42),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_43),
.B(n_51),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_44),
.B(n_47),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_44),
.B(n_53),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_44),
.B(n_54),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_L g53 ( 
.A1(n_45),
.A2(n_46),
.B1(n_48),
.B2(n_50),
.Y(n_53)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_47),
.B(n_52),
.Y(n_112)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_48),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_48),
.B(n_59),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_52),
.B(n_54),
.Y(n_51)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_52),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_57),
.B(n_60),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_57),
.A2(n_58),
.B1(n_60),
.B2(n_136),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_58),
.Y(n_57)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_60),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_L g60 ( 
.A1(n_61),
.A2(n_63),
.B(n_69),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_61),
.B(n_65),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_61),
.B(n_70),
.Y(n_75)
);

AOI21xp5_ASAP7_75t_L g160 ( 
.A1(n_61),
.A2(n_71),
.B(n_125),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_SL g209 ( 
.A(n_61),
.B(n_195),
.Y(n_209)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_62),
.B(n_124),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_SL g73 ( 
.A1(n_63),
.A2(n_71),
.B(n_74),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_64),
.A2(n_65),
.B1(n_81),
.B2(n_82),
.Y(n_84)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_65),
.B(n_213),
.Y(n_212)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

BUFx12f_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_69),
.B(n_123),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_69),
.B(n_208),
.Y(n_207)
);

OR2x2_ASAP7_75t_L g69 ( 
.A(n_70),
.B(n_71),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_71),
.B(n_125),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_71),
.B(n_195),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_L g146 ( 
.A(n_72),
.B(n_87),
.Y(n_146)
);

XOR2xp5_ASAP7_75t_L g72 ( 
.A(n_73),
.B(n_76),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_73),
.B(n_76),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_74),
.B(n_143),
.Y(n_142)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g216 ( 
.A(n_75),
.B(n_194),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_77),
.B(n_85),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_77),
.B(n_178),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_78),
.B(n_79),
.Y(n_77)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_78),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_78),
.B(n_164),
.Y(n_163)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_79),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_79),
.B(n_86),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_79),
.B(n_166),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_80),
.B(n_84),
.Y(n_79)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

BUFx3_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_84),
.B(n_86),
.Y(n_85)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_84),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_85),
.B(n_165),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_88),
.B(n_94),
.C(n_99),
.Y(n_87)
);

XOR2xp5_ASAP7_75t_L g132 ( 
.A(n_88),
.B(n_133),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_91),
.Y(n_88)
);

INVxp33_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_90),
.B(n_112),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_SL g91 ( 
.A(n_92),
.B(n_93),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_94),
.A2(n_95),
.B1(n_99),
.B2(n_134),
.Y(n_133)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

AOI21x1_ASAP7_75t_SL g95 ( 
.A1(n_96),
.A2(n_97),
.B(n_98),
.Y(n_95)
);

OAI21xp5_ASAP7_75t_L g119 ( 
.A1(n_96),
.A2(n_120),
.B(n_121),
.Y(n_119)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_96),
.Y(n_164)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_99),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_SL g99 ( 
.A(n_100),
.B(n_102),
.Y(n_99)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_103),
.B(n_180),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g104 ( 
.A(n_105),
.B(n_106),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_107),
.A2(n_108),
.B1(n_117),
.B2(n_118),
.Y(n_106)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

XOR2xp5_ASAP7_75t_L g108 ( 
.A(n_109),
.B(n_110),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_111),
.A2(n_113),
.B1(n_115),
.B2(n_116),
.Y(n_110)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_111),
.Y(n_115)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_113),
.Y(n_116)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

XOR2xp5_ASAP7_75t_L g118 ( 
.A(n_119),
.B(n_122),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_121),
.B(n_178),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_123),
.B(n_193),
.Y(n_192)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_128),
.B(n_147),
.Y(n_127)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_145),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_130),
.B(n_145),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_135),
.C(n_137),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_131),
.A2(n_132),
.B1(n_168),
.B2(n_169),
.Y(n_167)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

XOR2xp5_ASAP7_75t_L g169 ( 
.A(n_135),
.B(n_137),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_140),
.C(n_141),
.Y(n_137)
);

XOR2xp5_ASAP7_75t_L g153 ( 
.A(n_138),
.B(n_154),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_140),
.A2(n_141),
.B1(n_142),
.B2(n_155),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_140),
.Y(n_155)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

INVxp67_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_SL g214 ( 
.A(n_144),
.B(n_209),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_148),
.B(n_149),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_L g149 ( 
.A1(n_150),
.A2(n_170),
.B(n_227),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_167),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_151),
.B(n_167),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_156),
.C(n_161),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_152),
.A2(n_153),
.B1(n_173),
.B2(n_175),
.Y(n_172)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_156),
.A2(n_161),
.B1(n_162),
.B2(n_174),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_156),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_160),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_157),
.A2(n_158),
.B1(n_160),
.B2(n_182),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_158),
.Y(n_157)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_160),
.Y(n_182)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_165),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_164),
.B(n_166),
.Y(n_178)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

AOI21x1_ASAP7_75t_SL g170 ( 
.A1(n_171),
.A2(n_183),
.B(n_226),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_172),
.B(n_176),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_172),
.B(n_176),
.Y(n_226)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_173),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_177),
.B(n_179),
.C(n_181),
.Y(n_176)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_177),
.B(n_179),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_181),
.B(n_224),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_L g183 ( 
.A1(n_184),
.A2(n_221),
.B(n_225),
.Y(n_183)
);

AOI21xp5_ASAP7_75t_L g184 ( 
.A1(n_185),
.A2(n_203),
.B(n_220),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_191),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_186),
.B(n_191),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_187),
.B(n_190),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_L g205 ( 
.A1(n_187),
.A2(n_188),
.B1(n_190),
.B2(n_206),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_188),
.Y(n_187)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_190),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_192),
.A2(n_196),
.B1(n_197),
.B2(n_202),
.Y(n_191)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_192),
.Y(n_202)
);

INVxp67_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_198),
.A2(n_199),
.B1(n_200),
.B2(n_201),
.Y(n_197)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_198),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_199),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_199),
.B(n_200),
.C(n_202),
.Y(n_222)
);

OAI21xp5_ASAP7_75t_SL g203 ( 
.A1(n_204),
.A2(n_210),
.B(n_219),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_SL g204 ( 
.A(n_205),
.B(n_207),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_205),
.B(n_207),
.Y(n_219)
);

INVxp67_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

AOI21xp5_ASAP7_75t_L g210 ( 
.A1(n_211),
.A2(n_215),
.B(n_218),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_212),
.B(n_214),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_216),
.B(n_217),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_216),
.B(n_217),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_223),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_222),
.B(n_223),
.Y(n_225)
);


endmodule