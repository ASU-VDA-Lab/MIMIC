module fake_ariane_1696_n_1079 (n_83, n_8, n_56, n_60, n_170, n_160, n_64, n_119, n_124, n_167, n_90, n_38, n_47, n_110, n_153, n_18, n_86, n_75, n_89, n_67, n_176, n_149, n_34, n_158, n_172, n_69, n_95, n_175, n_92, n_143, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_152, n_120, n_169, n_106, n_12, n_53, n_173, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_156, n_49, n_20, n_174, n_100, n_17, n_50, n_132, n_62, n_147, n_51, n_166, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_159, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_178, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_148, n_164, n_52, n_157, n_177, n_135, n_73, n_77, n_171, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_151, n_136, n_28, n_80, n_146, n_97, n_154, n_142, n_161, n_14, n_163, n_88, n_141, n_68, n_116, n_104, n_145, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_1079);

input n_83;
input n_8;
input n_56;
input n_60;
input n_170;
input n_160;
input n_64;
input n_119;
input n_124;
input n_167;
input n_90;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_176;
input n_149;
input n_34;
input n_158;
input n_172;
input n_69;
input n_95;
input n_175;
input n_92;
input n_143;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_152;
input n_120;
input n_169;
input n_106;
input n_12;
input n_53;
input n_173;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_156;
input n_49;
input n_20;
input n_174;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_147;
input n_51;
input n_166;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_159;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_178;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_164;
input n_52;
input n_157;
input n_177;
input n_135;
input n_73;
input n_77;
input n_171;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_151;
input n_136;
input n_28;
input n_80;
input n_146;
input n_97;
input n_154;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_1079;

wire n_295;
wire n_356;
wire n_556;
wire n_190;
wire n_698;
wire n_1072;
wire n_695;
wire n_913;
wire n_180;
wire n_730;
wire n_386;
wire n_307;
wire n_516;
wire n_589;
wire n_332;
wire n_1008;
wire n_581;
wire n_294;
wire n_1020;
wire n_646;
wire n_197;
wire n_640;
wire n_463;
wire n_1024;
wire n_830;
wire n_691;
wire n_404;
wire n_943;
wire n_678;
wire n_1058;
wire n_651;
wire n_987;
wire n_936;
wire n_423;
wire n_347;
wire n_1042;
wire n_961;
wire n_183;
wire n_469;
wire n_1046;
wire n_479;
wire n_726;
wire n_603;
wire n_878;
wire n_373;
wire n_299;
wire n_836;
wire n_541;
wire n_499;
wire n_789;
wire n_788;
wire n_908;
wire n_850;
wire n_771;
wire n_1036;
wire n_564;
wire n_610;
wire n_205;
wire n_752;
wire n_341;
wire n_1029;
wire n_985;
wire n_421;
wire n_245;
wire n_549;
wire n_760;
wire n_522;
wire n_319;
wire n_591;
wire n_690;
wire n_906;
wire n_416;
wire n_969;
wire n_283;
wire n_919;
wire n_525;
wire n_187;
wire n_806;
wire n_367;
wire n_970;
wire n_713;
wire n_649;
wire n_598;
wire n_374;
wire n_345;
wire n_318;
wire n_817;
wire n_244;
wire n_643;
wire n_679;
wire n_226;
wire n_924;
wire n_927;
wire n_781;
wire n_261;
wire n_220;
wire n_682;
wire n_663;
wire n_370;
wire n_706;
wire n_189;
wire n_717;
wire n_819;
wire n_286;
wire n_443;
wire n_586;
wire n_952;
wire n_864;
wire n_686;
wire n_605;
wire n_776;
wire n_424;
wire n_528;
wire n_584;
wire n_387;
wire n_406;
wire n_826;
wire n_524;
wire n_634;
wire n_391;
wire n_349;
wire n_756;
wire n_466;
wire n_940;
wire n_1016;
wire n_346;
wire n_214;
wire n_764;
wire n_979;
wire n_348;
wire n_552;
wire n_1077;
wire n_462;
wire n_607;
wire n_670;
wire n_897;
wire n_949;
wire n_956;
wire n_410;
wire n_445;
wire n_515;
wire n_379;
wire n_807;
wire n_765;
wire n_264;
wire n_891;
wire n_737;
wire n_885;
wire n_198;
wire n_232;
wire n_441;
wire n_568;
wire n_1032;
wire n_385;
wire n_637;
wire n_917;
wire n_327;
wire n_766;
wire n_372;
wire n_377;
wire n_396;
wire n_802;
wire n_631;
wire n_399;
wire n_554;
wire n_960;
wire n_520;
wire n_980;
wire n_870;
wire n_714;
wire n_279;
wire n_945;
wire n_702;
wire n_958;
wire n_905;
wire n_207;
wire n_790;
wire n_898;
wire n_857;
wire n_363;
wire n_720;
wire n_968;
wire n_1067;
wire n_354;
wire n_813;
wire n_926;
wire n_725;
wire n_419;
wire n_1009;
wire n_230;
wire n_270;
wire n_194;
wire n_1064;
wire n_633;
wire n_900;
wire n_883;
wire n_338;
wire n_995;
wire n_285;
wire n_473;
wire n_186;
wire n_801;
wire n_202;
wire n_193;
wire n_733;
wire n_818;
wire n_761;
wire n_500;
wire n_665;
wire n_336;
wire n_754;
wire n_731;
wire n_779;
wire n_871;
wire n_315;
wire n_903;
wire n_1073;
wire n_594;
wire n_311;
wire n_239;
wire n_402;
wire n_1052;
wire n_1068;
wire n_272;
wire n_829;
wire n_1062;
wire n_668;
wire n_339;
wire n_738;
wire n_758;
wire n_833;
wire n_672;
wire n_487;
wire n_740;
wire n_879;
wire n_422;
wire n_648;
wire n_784;
wire n_269;
wire n_597;
wire n_816;
wire n_1018;
wire n_855;
wire n_1047;
wire n_259;
wire n_835;
wire n_808;
wire n_953;
wire n_446;
wire n_553;
wire n_1076;
wire n_753;
wire n_1050;
wire n_566;
wire n_814;
wire n_578;
wire n_701;
wire n_1003;
wire n_625;
wire n_405;
wire n_557;
wire n_989;
wire n_242;
wire n_645;
wire n_858;
wire n_320;
wire n_331;
wire n_309;
wire n_559;
wire n_401;
wire n_485;
wire n_267;
wire n_495;
wire n_504;
wire n_647;
wire n_483;
wire n_335;
wire n_435;
wire n_1035;
wire n_350;
wire n_291;
wire n_822;
wire n_381;
wire n_344;
wire n_795;
wire n_426;
wire n_433;
wire n_481;
wire n_600;
wire n_721;
wire n_1053;
wire n_840;
wire n_398;
wire n_210;
wire n_200;
wire n_529;
wire n_502;
wire n_253;
wire n_561;
wire n_770;
wire n_218;
wire n_821;
wire n_928;
wire n_839;
wire n_271;
wire n_465;
wire n_486;
wire n_507;
wire n_901;
wire n_759;
wire n_247;
wire n_569;
wire n_567;
wire n_825;
wire n_732;
wire n_971;
wire n_240;
wire n_369;
wire n_224;
wire n_787;
wire n_894;
wire n_547;
wire n_420;
wire n_562;
wire n_518;
wire n_439;
wire n_604;
wire n_614;
wire n_677;
wire n_222;
wire n_478;
wire n_703;
wire n_748;
wire n_786;
wire n_510;
wire n_1061;
wire n_1045;
wire n_868;
wire n_256;
wire n_831;
wire n_326;
wire n_681;
wire n_778;
wire n_227;
wire n_874;
wire n_188;
wire n_323;
wire n_550;
wire n_1023;
wire n_988;
wire n_635;
wire n_707;
wire n_997;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_694;
wire n_884;
wire n_983;
wire n_282;
wire n_328;
wire n_368;
wire n_1034;
wire n_590;
wire n_699;
wire n_727;
wire n_277;
wire n_248;
wire n_301;
wire n_467;
wire n_432;
wire n_545;
wire n_1015;
wire n_536;
wire n_644;
wire n_293;
wire n_823;
wire n_921;
wire n_620;
wire n_228;
wire n_325;
wire n_276;
wire n_688;
wire n_1074;
wire n_859;
wire n_636;
wire n_427;
wire n_587;
wire n_497;
wire n_693;
wire n_863;
wire n_303;
wire n_671;
wire n_442;
wire n_777;
wire n_929;
wire n_206;
wire n_352;
wire n_538;
wire n_899;
wire n_920;
wire n_576;
wire n_843;
wire n_511;
wire n_611;
wire n_455;
wire n_365;
wire n_429;
wire n_654;
wire n_238;
wire n_588;
wire n_1013;
wire n_986;
wire n_638;
wire n_334;
wire n_192;
wire n_729;
wire n_887;
wire n_661;
wire n_488;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_300;
wire n_533;
wire n_904;
wire n_505;
wire n_869;
wire n_846;
wire n_390;
wire n_498;
wire n_501;
wire n_438;
wire n_1059;
wire n_314;
wire n_684;
wire n_440;
wire n_627;
wire n_1039;
wire n_273;
wire n_305;
wire n_539;
wire n_312;
wire n_233;
wire n_728;
wire n_388;
wire n_333;
wire n_449;
wire n_612;
wire n_413;
wire n_392;
wire n_376;
wire n_957;
wire n_977;
wire n_512;
wire n_715;
wire n_889;
wire n_1066;
wire n_935;
wire n_579;
wire n_844;
wire n_1012;
wire n_459;
wire n_685;
wire n_221;
wire n_321;
wire n_911;
wire n_458;
wire n_361;
wire n_383;
wire n_623;
wire n_838;
wire n_237;
wire n_780;
wire n_861;
wire n_950;
wire n_1017;
wire n_711;
wire n_877;
wire n_1021;
wire n_1065;
wire n_453;
wire n_734;
wire n_491;
wire n_810;
wire n_181;
wire n_723;
wire n_617;
wire n_616;
wire n_658;
wire n_630;
wire n_705;
wire n_570;
wire n_1055;
wire n_260;
wire n_362;
wire n_543;
wire n_942;
wire n_310;
wire n_709;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_281;
wire n_628;
wire n_809;
wire n_461;
wire n_490;
wire n_262;
wire n_209;
wire n_743;
wire n_225;
wire n_907;
wire n_235;
wire n_1006;
wire n_881;
wire n_660;
wire n_464;
wire n_735;
wire n_575;
wire n_546;
wire n_1019;
wire n_297;
wire n_962;
wire n_662;
wire n_641;
wire n_1005;
wire n_503;
wire n_941;
wire n_700;
wire n_910;
wire n_290;
wire n_527;
wire n_747;
wire n_741;
wire n_772;
wire n_847;
wire n_939;
wire n_371;
wire n_845;
wire n_888;
wire n_199;
wire n_918;
wire n_639;
wire n_217;
wire n_452;
wire n_673;
wire n_676;
wire n_551;
wire n_308;
wire n_708;
wire n_417;
wire n_201;
wire n_1038;
wire n_572;
wire n_343;
wire n_865;
wire n_1041;
wire n_414;
wire n_571;
wire n_680;
wire n_287;
wire n_302;
wire n_993;
wire n_380;
wire n_948;
wire n_582;
wire n_284;
wire n_922;
wire n_1004;
wire n_448;
wire n_593;
wire n_755;
wire n_710;
wire n_860;
wire n_249;
wire n_534;
wire n_212;
wire n_444;
wire n_355;
wire n_609;
wire n_278;
wire n_851;
wire n_1043;
wire n_255;
wire n_560;
wire n_450;
wire n_890;
wire n_257;
wire n_842;
wire n_652;
wire n_451;
wire n_613;
wire n_745;
wire n_475;
wire n_1022;
wire n_1033;
wire n_896;
wire n_409;
wire n_947;
wire n_930;
wire n_519;
wire n_902;
wire n_384;
wire n_1031;
wire n_468;
wire n_1056;
wire n_853;
wire n_526;
wire n_716;
wire n_742;
wire n_182;
wire n_696;
wire n_1040;
wire n_674;
wire n_482;
wire n_316;
wire n_196;
wire n_798;
wire n_769;
wire n_820;
wire n_577;
wire n_407;
wire n_774;
wire n_933;
wire n_872;
wire n_916;
wire n_254;
wire n_596;
wire n_954;
wire n_912;
wire n_476;
wire n_460;
wire n_219;
wire n_832;
wire n_535;
wire n_231;
wire n_366;
wire n_744;
wire n_762;
wire n_656;
wire n_555;
wire n_234;
wire n_492;
wire n_574;
wire n_848;
wire n_804;
wire n_280;
wire n_982;
wire n_915;
wire n_215;
wire n_252;
wire n_629;
wire n_664;
wire n_1075;
wire n_454;
wire n_966;
wire n_992;
wire n_298;
wire n_955;
wire n_532;
wire n_415;
wire n_794;
wire n_763;
wire n_655;
wire n_544;
wire n_540;
wire n_216;
wire n_692;
wire n_599;
wire n_768;
wire n_514;
wire n_418;
wire n_984;
wire n_537;
wire n_1063;
wire n_223;
wire n_403;
wire n_750;
wire n_834;
wire n_991;
wire n_389;
wire n_1007;
wire n_800;
wire n_657;
wire n_513;
wire n_837;
wire n_288;
wire n_179;
wire n_812;
wire n_395;
wire n_621;
wire n_195;
wire n_606;
wire n_951;
wire n_1026;
wire n_213;
wire n_938;
wire n_862;
wire n_304;
wire n_895;
wire n_659;
wire n_583;
wire n_509;
wire n_1014;
wire n_724;
wire n_306;
wire n_666;
wire n_1000;
wire n_313;
wire n_430;
wire n_626;
wire n_493;
wire n_722;
wire n_203;
wire n_378;
wire n_436;
wire n_946;
wire n_757;
wire n_375;
wire n_324;
wire n_1030;
wire n_585;
wire n_875;
wire n_669;
wire n_785;
wire n_827;
wire n_931;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_622;
wire n_697;
wire n_967;
wire n_998;
wire n_999;
wire n_472;
wire n_937;
wire n_296;
wire n_265;
wire n_746;
wire n_208;
wire n_456;
wire n_292;
wire n_880;
wire n_793;
wire n_852;
wire n_275;
wire n_704;
wire n_1060;
wire n_1044;
wire n_204;
wire n_751;
wire n_615;
wire n_1027;
wire n_1070;
wire n_996;
wire n_521;
wire n_963;
wire n_873;
wire n_496;
wire n_739;
wire n_1028;
wire n_342;
wire n_866;
wire n_246;
wire n_517;
wire n_925;
wire n_530;
wire n_792;
wire n_1001;
wire n_824;
wire n_428;
wire n_1002;
wire n_358;
wire n_580;
wire n_892;
wire n_608;
wire n_959;
wire n_494;
wire n_1051;
wire n_719;
wire n_263;
wire n_434;
wire n_360;
wire n_975;
wire n_563;
wire n_229;
wire n_394;
wire n_923;
wire n_250;
wire n_932;
wire n_773;
wire n_1037;
wire n_981;
wire n_1010;
wire n_882;
wire n_990;
wire n_317;
wire n_867;
wire n_243;
wire n_803;
wire n_329;
wire n_718;
wire n_185;
wire n_340;
wire n_944;
wire n_749;
wire n_994;
wire n_289;
wire n_548;
wire n_542;
wire n_815;
wire n_973;
wire n_523;
wire n_1078;
wire n_268;
wire n_972;
wire n_266;
wire n_470;
wire n_457;
wire n_632;
wire n_184;
wire n_477;
wire n_364;
wire n_258;
wire n_650;
wire n_782;
wire n_856;
wire n_425;
wire n_431;
wire n_811;
wire n_1054;
wire n_508;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1071;
wire n_411;
wire n_484;
wire n_712;
wire n_976;
wire n_909;
wire n_849;
wire n_353;
wire n_736;
wire n_767;
wire n_1025;
wire n_241;
wire n_357;
wire n_412;
wire n_687;
wire n_447;
wire n_964;
wire n_1057;
wire n_191;
wire n_382;
wire n_797;
wire n_489;
wire n_480;
wire n_978;
wire n_642;
wire n_211;
wire n_1011;
wire n_408;
wire n_828;
wire n_595;
wire n_322;
wire n_251;
wire n_974;
wire n_506;
wire n_893;
wire n_602;
wire n_799;
wire n_558;
wire n_592;
wire n_397;
wire n_841;
wire n_854;
wire n_471;
wire n_351;
wire n_886;
wire n_965;
wire n_393;
wire n_1069;
wire n_474;
wire n_653;
wire n_359;
wire n_573;
wire n_796;
wire n_805;
wire n_531;
wire n_934;
wire n_783;
wire n_675;

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_84),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_156),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_169),
.Y(n_181)
);

BUFx3_ASAP7_75t_L g182 ( 
.A(n_2),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_109),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_173),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_168),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_172),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_47),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_56),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_146),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_128),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_167),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_49),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_107),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_159),
.Y(n_194)
);

INVxp67_ASAP7_75t_L g195 ( 
.A(n_22),
.Y(n_195)
);

BUFx8_ASAP7_75t_SL g196 ( 
.A(n_162),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_143),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_118),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_127),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_35),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_12),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_102),
.Y(n_202)
);

BUFx10_ASAP7_75t_L g203 ( 
.A(n_9),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_142),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_88),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_25),
.Y(n_206)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_153),
.Y(n_207)
);

BUFx10_ASAP7_75t_L g208 ( 
.A(n_51),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_161),
.Y(n_209)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_64),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_39),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_11),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_23),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_89),
.Y(n_214)
);

INVx1_ASAP7_75t_SL g215 ( 
.A(n_2),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_65),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_123),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_59),
.Y(n_218)
);

BUFx10_ASAP7_75t_L g219 ( 
.A(n_166),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_119),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_157),
.Y(n_221)
);

BUFx3_ASAP7_75t_L g222 ( 
.A(n_163),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_58),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_48),
.Y(n_224)
);

BUFx3_ASAP7_75t_L g225 ( 
.A(n_24),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_141),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_46),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_165),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_151),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_170),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_0),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_72),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_164),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_20),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_43),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_100),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_66),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_113),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_104),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_68),
.Y(n_240)
);

INVx1_ASAP7_75t_SL g241 ( 
.A(n_93),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_38),
.Y(n_242)
);

BUFx10_ASAP7_75t_L g243 ( 
.A(n_174),
.Y(n_243)
);

INVx1_ASAP7_75t_SL g244 ( 
.A(n_101),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_24),
.Y(n_245)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_27),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_14),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_27),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_114),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_160),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_171),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_246),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_182),
.Y(n_253)
);

HB1xp67_ASAP7_75t_L g254 ( 
.A(n_182),
.Y(n_254)
);

BUFx2_ASAP7_75t_L g255 ( 
.A(n_225),
.Y(n_255)
);

BUFx2_ASAP7_75t_L g256 ( 
.A(n_225),
.Y(n_256)
);

CKINVDCx16_ASAP7_75t_R g257 ( 
.A(n_203),
.Y(n_257)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_222),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_246),
.Y(n_259)
);

INVxp33_ASAP7_75t_L g260 ( 
.A(n_201),
.Y(n_260)
);

INVxp67_ASAP7_75t_SL g261 ( 
.A(n_195),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_207),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_196),
.Y(n_263)
);

BUFx2_ASAP7_75t_SL g264 ( 
.A(n_237),
.Y(n_264)
);

INVxp33_ASAP7_75t_SL g265 ( 
.A(n_206),
.Y(n_265)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_222),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_207),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_196),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_210),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_210),
.Y(n_270)
);

HB1xp67_ASAP7_75t_L g271 ( 
.A(n_212),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_237),
.Y(n_272)
);

BUFx2_ASAP7_75t_L g273 ( 
.A(n_213),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_208),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_208),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_180),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_208),
.Y(n_277)
);

INVxp67_ASAP7_75t_L g278 ( 
.A(n_203),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_219),
.Y(n_279)
);

INVxp67_ASAP7_75t_SL g280 ( 
.A(n_183),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_219),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_219),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_234),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_243),
.Y(n_284)
);

INVxp67_ASAP7_75t_L g285 ( 
.A(n_203),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_243),
.Y(n_286)
);

INVx1_ASAP7_75t_SL g287 ( 
.A(n_245),
.Y(n_287)
);

INVxp67_ASAP7_75t_L g288 ( 
.A(n_231),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_243),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_185),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_187),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_188),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_197),
.Y(n_293)
);

INVxp67_ASAP7_75t_SL g294 ( 
.A(n_200),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_205),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_189),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_216),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_217),
.Y(n_298)
);

INVxp67_ASAP7_75t_SL g299 ( 
.A(n_221),
.Y(n_299)
);

CKINVDCx14_ASAP7_75t_R g300 ( 
.A(n_232),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_262),
.Y(n_301)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_262),
.Y(n_302)
);

INVxp67_ASAP7_75t_L g303 ( 
.A(n_273),
.Y(n_303)
);

INVx2_ASAP7_75t_L g304 ( 
.A(n_267),
.Y(n_304)
);

OAI21x1_ASAP7_75t_L g305 ( 
.A1(n_276),
.A2(n_224),
.B(n_223),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_267),
.Y(n_306)
);

AND2x2_ASAP7_75t_L g307 ( 
.A(n_255),
.B(n_215),
.Y(n_307)
);

BUFx3_ASAP7_75t_L g308 ( 
.A(n_258),
.Y(n_308)
);

INVxp33_ASAP7_75t_SL g309 ( 
.A(n_263),
.Y(n_309)
);

AND2x2_ASAP7_75t_L g310 ( 
.A(n_255),
.B(n_256),
.Y(n_310)
);

INVx2_ASAP7_75t_L g311 ( 
.A(n_269),
.Y(n_311)
);

AND2x4_ASAP7_75t_L g312 ( 
.A(n_280),
.B(n_230),
.Y(n_312)
);

AND2x2_ASAP7_75t_L g313 ( 
.A(n_256),
.B(n_247),
.Y(n_313)
);

HB1xp67_ASAP7_75t_L g314 ( 
.A(n_263),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_L g315 ( 
.A1(n_265),
.A2(n_234),
.B1(n_249),
.B2(n_248),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_269),
.Y(n_316)
);

BUFx12f_ASAP7_75t_L g317 ( 
.A(n_268),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_270),
.Y(n_318)
);

BUFx6f_ASAP7_75t_L g319 ( 
.A(n_270),
.Y(n_319)
);

AND2x6_ASAP7_75t_L g320 ( 
.A(n_276),
.B(n_233),
.Y(n_320)
);

AND2x6_ASAP7_75t_L g321 ( 
.A(n_295),
.B(n_235),
.Y(n_321)
);

OA21x2_ASAP7_75t_L g322 ( 
.A1(n_295),
.A2(n_251),
.B(n_236),
.Y(n_322)
);

INVxp33_ASAP7_75t_SL g323 ( 
.A(n_268),
.Y(n_323)
);

INVx4_ASAP7_75t_L g324 ( 
.A(n_258),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_296),
.Y(n_325)
);

INVx2_ASAP7_75t_L g326 ( 
.A(n_252),
.Y(n_326)
);

INVx2_ASAP7_75t_L g327 ( 
.A(n_266),
.Y(n_327)
);

BUFx2_ASAP7_75t_L g328 ( 
.A(n_273),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_274),
.B(n_241),
.Y(n_329)
);

AND2x4_ASAP7_75t_L g330 ( 
.A(n_294),
.B(n_244),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_297),
.Y(n_331)
);

AND2x2_ASAP7_75t_L g332 ( 
.A(n_260),
.B(n_179),
.Y(n_332)
);

BUFx6f_ASAP7_75t_L g333 ( 
.A(n_266),
.Y(n_333)
);

INVx2_ASAP7_75t_L g334 ( 
.A(n_252),
.Y(n_334)
);

INVx3_ASAP7_75t_L g335 ( 
.A(n_297),
.Y(n_335)
);

OA21x2_ASAP7_75t_L g336 ( 
.A1(n_298),
.A2(n_184),
.B(n_181),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_298),
.Y(n_337)
);

BUFx12f_ASAP7_75t_L g338 ( 
.A(n_296),
.Y(n_338)
);

INVx2_ASAP7_75t_L g339 ( 
.A(n_259),
.Y(n_339)
);

BUFx6f_ASAP7_75t_L g340 ( 
.A(n_259),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_300),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_290),
.Y(n_342)
);

AND2x4_ASAP7_75t_L g343 ( 
.A(n_299),
.B(n_291),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_292),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_293),
.Y(n_345)
);

INVx5_ASAP7_75t_L g346 ( 
.A(n_257),
.Y(n_346)
);

INVxp67_ASAP7_75t_L g347 ( 
.A(n_271),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_SL g348 ( 
.A(n_275),
.B(n_186),
.Y(n_348)
);

BUFx2_ASAP7_75t_L g349 ( 
.A(n_272),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_253),
.Y(n_350)
);

INVx2_ASAP7_75t_L g351 ( 
.A(n_254),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_277),
.Y(n_352)
);

INVx2_ASAP7_75t_L g353 ( 
.A(n_279),
.Y(n_353)
);

OAI22x1_ASAP7_75t_SL g354 ( 
.A1(n_283),
.A2(n_250),
.B1(n_242),
.B2(n_240),
.Y(n_354)
);

AND2x2_ASAP7_75t_L g355 ( 
.A(n_281),
.B(n_190),
.Y(n_355)
);

INVx2_ASAP7_75t_L g356 ( 
.A(n_319),
.Y(n_356)
);

INVx2_ASAP7_75t_L g357 ( 
.A(n_319),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_335),
.Y(n_358)
);

INVx2_ASAP7_75t_SL g359 ( 
.A(n_346),
.Y(n_359)
);

INVxp33_ASAP7_75t_L g360 ( 
.A(n_328),
.Y(n_360)
);

INVx2_ASAP7_75t_L g361 ( 
.A(n_319),
.Y(n_361)
);

INVx8_ASAP7_75t_L g362 ( 
.A(n_320),
.Y(n_362)
);

INVx2_ASAP7_75t_L g363 ( 
.A(n_319),
.Y(n_363)
);

INVx2_ASAP7_75t_L g364 ( 
.A(n_319),
.Y(n_364)
);

INVx2_ASAP7_75t_L g365 ( 
.A(n_340),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_SL g366 ( 
.A(n_332),
.B(n_346),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_335),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_335),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_335),
.Y(n_369)
);

INVx1_ASAP7_75t_SL g370 ( 
.A(n_328),
.Y(n_370)
);

INVx3_ASAP7_75t_L g371 ( 
.A(n_333),
.Y(n_371)
);

INVx2_ASAP7_75t_SL g372 ( 
.A(n_346),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_331),
.Y(n_373)
);

NOR2xp33_ASAP7_75t_L g374 ( 
.A(n_352),
.B(n_265),
.Y(n_374)
);

INVx2_ASAP7_75t_SL g375 ( 
.A(n_346),
.Y(n_375)
);

BUFx3_ASAP7_75t_L g376 ( 
.A(n_308),
.Y(n_376)
);

INVx2_ASAP7_75t_L g377 ( 
.A(n_340),
.Y(n_377)
);

INVx2_ASAP7_75t_L g378 ( 
.A(n_340),
.Y(n_378)
);

INVx2_ASAP7_75t_L g379 ( 
.A(n_340),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_331),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_SL g381 ( 
.A(n_332),
.B(n_278),
.Y(n_381)
);

INVx2_ASAP7_75t_L g382 ( 
.A(n_340),
.Y(n_382)
);

INVx2_ASAP7_75t_L g383 ( 
.A(n_333),
.Y(n_383)
);

INVx2_ASAP7_75t_L g384 ( 
.A(n_333),
.Y(n_384)
);

INVx2_ASAP7_75t_L g385 ( 
.A(n_333),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_337),
.Y(n_386)
);

INVx2_ASAP7_75t_L g387 ( 
.A(n_333),
.Y(n_387)
);

INVx3_ASAP7_75t_L g388 ( 
.A(n_324),
.Y(n_388)
);

INVx2_ASAP7_75t_L g389 ( 
.A(n_326),
.Y(n_389)
);

BUFx6f_ASAP7_75t_SL g390 ( 
.A(n_330),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_337),
.Y(n_391)
);

INVx3_ASAP7_75t_L g392 ( 
.A(n_324),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_302),
.Y(n_393)
);

BUFx6f_ASAP7_75t_SL g394 ( 
.A(n_330),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_302),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_330),
.B(n_282),
.Y(n_396)
);

BUFx10_ASAP7_75t_L g397 ( 
.A(n_341),
.Y(n_397)
);

INVx2_ASAP7_75t_SL g398 ( 
.A(n_346),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_304),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_330),
.B(n_284),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_343),
.B(n_286),
.Y(n_401)
);

HB1xp67_ASAP7_75t_L g402 ( 
.A(n_349),
.Y(n_402)
);

INVxp67_ASAP7_75t_L g403 ( 
.A(n_349),
.Y(n_403)
);

NOR2x1p5_ASAP7_75t_L g404 ( 
.A(n_317),
.B(n_313),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_SL g405 ( 
.A(n_346),
.B(n_285),
.Y(n_405)
);

INVx2_ASAP7_75t_L g406 ( 
.A(n_326),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_304),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_311),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_311),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_301),
.Y(n_410)
);

AND3x2_ASAP7_75t_L g411 ( 
.A(n_314),
.B(n_261),
.C(n_289),
.Y(n_411)
);

NOR2xp33_ASAP7_75t_L g412 ( 
.A(n_352),
.B(n_288),
.Y(n_412)
);

AND2x2_ASAP7_75t_L g413 ( 
.A(n_343),
.B(n_264),
.Y(n_413)
);

INVx2_ASAP7_75t_L g414 ( 
.A(n_326),
.Y(n_414)
);

INVx11_ASAP7_75t_L g415 ( 
.A(n_317),
.Y(n_415)
);

INVx2_ASAP7_75t_L g416 ( 
.A(n_334),
.Y(n_416)
);

INVxp33_ASAP7_75t_L g417 ( 
.A(n_307),
.Y(n_417)
);

INVx2_ASAP7_75t_L g418 ( 
.A(n_334),
.Y(n_418)
);

BUFx6f_ASAP7_75t_SL g419 ( 
.A(n_343),
.Y(n_419)
);

OAI22xp33_ASAP7_75t_L g420 ( 
.A1(n_315),
.A2(n_272),
.B1(n_287),
.B2(n_264),
.Y(n_420)
);

AND2x2_ASAP7_75t_L g421 ( 
.A(n_343),
.B(n_191),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_SL g422 ( 
.A(n_329),
.B(n_192),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_301),
.Y(n_423)
);

INVx2_ASAP7_75t_SL g424 ( 
.A(n_310),
.Y(n_424)
);

INVx2_ASAP7_75t_L g425 ( 
.A(n_339),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_312),
.B(n_193),
.Y(n_426)
);

AND3x2_ASAP7_75t_L g427 ( 
.A(n_303),
.B(n_0),
.C(n_1),
.Y(n_427)
);

INVx2_ASAP7_75t_SL g428 ( 
.A(n_310),
.Y(n_428)
);

INVx2_ASAP7_75t_L g429 ( 
.A(n_339),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_358),
.Y(n_430)
);

NOR2xp33_ASAP7_75t_SL g431 ( 
.A(n_362),
.B(n_338),
.Y(n_431)
);

CKINVDCx20_ASAP7_75t_R g432 ( 
.A(n_397),
.Y(n_432)
);

AOI21xp5_ASAP7_75t_L g433 ( 
.A1(n_358),
.A2(n_368),
.B(n_367),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_367),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_368),
.Y(n_435)
);

XNOR2xp5_ASAP7_75t_L g436 ( 
.A(n_404),
.B(n_325),
.Y(n_436)
);

INVx2_ASAP7_75t_L g437 ( 
.A(n_376),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_415),
.Y(n_438)
);

NOR2xp33_ASAP7_75t_L g439 ( 
.A(n_417),
.B(n_309),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_369),
.Y(n_440)
);

CKINVDCx20_ASAP7_75t_R g441 ( 
.A(n_397),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_369),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_373),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_373),
.Y(n_444)
);

INVxp33_ASAP7_75t_L g445 ( 
.A(n_360),
.Y(n_445)
);

INVx2_ASAP7_75t_SL g446 ( 
.A(n_413),
.Y(n_446)
);

AND2x2_ASAP7_75t_L g447 ( 
.A(n_370),
.B(n_307),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_380),
.Y(n_448)
);

NOR2xp33_ASAP7_75t_L g449 ( 
.A(n_374),
.B(n_355),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_380),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_386),
.Y(n_451)
);

OR2x2_ASAP7_75t_L g452 ( 
.A(n_370),
.B(n_402),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_386),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_391),
.Y(n_454)
);

INVx2_ASAP7_75t_L g455 ( 
.A(n_376),
.Y(n_455)
);

AND2x4_ASAP7_75t_L g456 ( 
.A(n_413),
.B(n_353),
.Y(n_456)
);

CKINVDCx16_ASAP7_75t_R g457 ( 
.A(n_397),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_391),
.Y(n_458)
);

CKINVDCx16_ASAP7_75t_R g459 ( 
.A(n_419),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_410),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_410),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_423),
.Y(n_462)
);

CKINVDCx20_ASAP7_75t_R g463 ( 
.A(n_403),
.Y(n_463)
);

AOI21xp5_ASAP7_75t_L g464 ( 
.A1(n_423),
.A2(n_336),
.B(n_305),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_393),
.Y(n_465)
);

XOR2xp5_ASAP7_75t_L g466 ( 
.A(n_420),
.B(n_323),
.Y(n_466)
);

AND2x2_ASAP7_75t_L g467 ( 
.A(n_424),
.B(n_313),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_393),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_395),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_395),
.Y(n_470)
);

NOR2xp33_ASAP7_75t_L g471 ( 
.A(n_419),
.B(n_355),
.Y(n_471)
);

NAND2xp33_ASAP7_75t_R g472 ( 
.A(n_411),
.B(n_336),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_399),
.Y(n_473)
);

XOR2xp5_ASAP7_75t_L g474 ( 
.A(n_381),
.B(n_315),
.Y(n_474)
);

BUFx8_ASAP7_75t_L g475 ( 
.A(n_390),
.Y(n_475)
);

NOR2xp33_ASAP7_75t_L g476 ( 
.A(n_419),
.B(n_348),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_399),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_407),
.Y(n_478)
);

INVx2_ASAP7_75t_L g479 ( 
.A(n_389),
.Y(n_479)
);

NOR2xp33_ASAP7_75t_L g480 ( 
.A(n_396),
.B(n_353),
.Y(n_480)
);

XOR2xp5_ASAP7_75t_L g481 ( 
.A(n_424),
.B(n_354),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_407),
.Y(n_482)
);

CKINVDCx20_ASAP7_75t_R g483 ( 
.A(n_428),
.Y(n_483)
);

XOR2xp5_ASAP7_75t_L g484 ( 
.A(n_428),
.B(n_354),
.Y(n_484)
);

NOR2xp33_ASAP7_75t_L g485 ( 
.A(n_400),
.B(n_412),
.Y(n_485)
);

BUFx6f_ASAP7_75t_L g486 ( 
.A(n_362),
.Y(n_486)
);

AND2x2_ASAP7_75t_L g487 ( 
.A(n_421),
.B(n_347),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_408),
.Y(n_488)
);

CKINVDCx5p33_ASAP7_75t_R g489 ( 
.A(n_415),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_408),
.Y(n_490)
);

BUFx6f_ASAP7_75t_SL g491 ( 
.A(n_404),
.Y(n_491)
);

INVxp33_ASAP7_75t_L g492 ( 
.A(n_421),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_409),
.Y(n_493)
);

AND2x4_ASAP7_75t_L g494 ( 
.A(n_401),
.B(n_312),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_409),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_416),
.Y(n_496)
);

INVx2_ASAP7_75t_L g497 ( 
.A(n_389),
.Y(n_497)
);

CKINVDCx5p33_ASAP7_75t_R g498 ( 
.A(n_390),
.Y(n_498)
);

CKINVDCx5p33_ASAP7_75t_R g499 ( 
.A(n_390),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_416),
.Y(n_500)
);

XOR2xp5_ASAP7_75t_L g501 ( 
.A(n_405),
.B(n_338),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_418),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_418),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_425),
.Y(n_504)
);

XNOR2xp5_ASAP7_75t_L g505 ( 
.A(n_422),
.B(n_351),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_L g506 ( 
.A(n_406),
.B(n_312),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_425),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_429),
.Y(n_508)
);

BUFx2_ASAP7_75t_L g509 ( 
.A(n_426),
.Y(n_509)
);

OR2x2_ASAP7_75t_L g510 ( 
.A(n_429),
.B(n_351),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_406),
.Y(n_511)
);

INVx2_ASAP7_75t_L g512 ( 
.A(n_414),
.Y(n_512)
);

NAND2x1p5_ASAP7_75t_L g513 ( 
.A(n_486),
.B(n_359),
.Y(n_513)
);

NOR2xp33_ASAP7_75t_L g514 ( 
.A(n_492),
.B(n_394),
.Y(n_514)
);

AND2x4_ASAP7_75t_L g515 ( 
.A(n_446),
.B(n_312),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_443),
.Y(n_516)
);

AND2x4_ASAP7_75t_L g517 ( 
.A(n_456),
.B(n_494),
.Y(n_517)
);

AND2x2_ASAP7_75t_L g518 ( 
.A(n_447),
.B(n_351),
.Y(n_518)
);

INVx2_ASAP7_75t_SL g519 ( 
.A(n_452),
.Y(n_519)
);

OAI22xp33_ASAP7_75t_L g520 ( 
.A1(n_449),
.A2(n_344),
.B1(n_345),
.B2(n_342),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_L g521 ( 
.A(n_485),
.B(n_388),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_444),
.Y(n_522)
);

NAND2x1_ASAP7_75t_L g523 ( 
.A(n_486),
.B(n_371),
.Y(n_523)
);

NOR2x2_ASAP7_75t_L g524 ( 
.A(n_463),
.B(n_427),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_SL g525 ( 
.A(n_486),
.B(n_359),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_448),
.Y(n_526)
);

HB1xp67_ASAP7_75t_L g527 ( 
.A(n_456),
.Y(n_527)
);

INVx2_ASAP7_75t_L g528 ( 
.A(n_479),
.Y(n_528)
);

INVx2_ASAP7_75t_L g529 ( 
.A(n_497),
.Y(n_529)
);

INVx3_ASAP7_75t_L g530 ( 
.A(n_437),
.Y(n_530)
);

AOI22xp33_ASAP7_75t_L g531 ( 
.A1(n_474),
.A2(n_321),
.B1(n_320),
.B2(n_394),
.Y(n_531)
);

AND2x2_ASAP7_75t_L g532 ( 
.A(n_487),
.B(n_342),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_L g533 ( 
.A(n_485),
.B(n_388),
.Y(n_533)
);

AOI22xp5_ASAP7_75t_L g534 ( 
.A1(n_449),
.A2(n_394),
.B1(n_366),
.B2(n_375),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_SL g535 ( 
.A(n_450),
.B(n_372),
.Y(n_535)
);

NOR2xp67_ASAP7_75t_L g536 ( 
.A(n_438),
.B(n_324),
.Y(n_536)
);

INVx2_ASAP7_75t_SL g537 ( 
.A(n_475),
.Y(n_537)
);

INVx2_ASAP7_75t_L g538 ( 
.A(n_512),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_451),
.Y(n_539)
);

HB1xp67_ASAP7_75t_L g540 ( 
.A(n_483),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_L g541 ( 
.A(n_494),
.B(n_388),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_SL g542 ( 
.A(n_453),
.B(n_372),
.Y(n_542)
);

OAI22xp5_ASAP7_75t_L g543 ( 
.A1(n_454),
.A2(n_392),
.B1(n_362),
.B2(n_375),
.Y(n_543)
);

HB1xp67_ASAP7_75t_L g544 ( 
.A(n_467),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_458),
.Y(n_545)
);

AOI21xp5_ASAP7_75t_L g546 ( 
.A1(n_433),
.A2(n_392),
.B(n_362),
.Y(n_546)
);

NOR2xp33_ASAP7_75t_L g547 ( 
.A(n_509),
.B(n_392),
.Y(n_547)
);

INVx2_ASAP7_75t_L g548 ( 
.A(n_511),
.Y(n_548)
);

AOI22xp33_ASAP7_75t_L g549 ( 
.A1(n_506),
.A2(n_321),
.B1(n_320),
.B2(n_414),
.Y(n_549)
);

INVx2_ASAP7_75t_SL g550 ( 
.A(n_475),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_L g551 ( 
.A(n_480),
.B(n_398),
.Y(n_551)
);

AOI22xp33_ASAP7_75t_L g552 ( 
.A1(n_506),
.A2(n_321),
.B1(n_320),
.B2(n_336),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_L g553 ( 
.A(n_480),
.B(n_398),
.Y(n_553)
);

A2O1A1Ixp33_ASAP7_75t_L g554 ( 
.A1(n_460),
.A2(n_305),
.B(n_345),
.C(n_344),
.Y(n_554)
);

AOI22xp33_ASAP7_75t_SL g555 ( 
.A1(n_459),
.A2(n_362),
.B1(n_321),
.B2(n_320),
.Y(n_555)
);

INVx2_ASAP7_75t_L g556 ( 
.A(n_496),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_L g557 ( 
.A(n_510),
.B(n_308),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_461),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_L g559 ( 
.A(n_462),
.B(n_308),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_430),
.Y(n_560)
);

AND2x4_ASAP7_75t_L g561 ( 
.A(n_471),
.B(n_498),
.Y(n_561)
);

INVx2_ASAP7_75t_L g562 ( 
.A(n_500),
.Y(n_562)
);

INVxp67_ASAP7_75t_SL g563 ( 
.A(n_445),
.Y(n_563)
);

BUFx6f_ASAP7_75t_L g564 ( 
.A(n_455),
.Y(n_564)
);

NOR2xp33_ASAP7_75t_L g565 ( 
.A(n_471),
.B(n_371),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_434),
.Y(n_566)
);

AOI22xp33_ASAP7_75t_L g567 ( 
.A1(n_465),
.A2(n_321),
.B1(n_320),
.B2(n_336),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_L g568 ( 
.A(n_468),
.B(n_324),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_L g569 ( 
.A(n_469),
.B(n_320),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_435),
.Y(n_570)
);

AND2x2_ASAP7_75t_L g571 ( 
.A(n_439),
.B(n_350),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_L g572 ( 
.A(n_470),
.B(n_321),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_SL g573 ( 
.A(n_440),
.B(n_356),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_442),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_516),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_L g576 ( 
.A(n_521),
.B(n_473),
.Y(n_576)
);

NOR2xp33_ASAP7_75t_L g577 ( 
.A(n_519),
.B(n_466),
.Y(n_577)
);

BUFx3_ASAP7_75t_L g578 ( 
.A(n_537),
.Y(n_578)
);

BUFx8_ASAP7_75t_L g579 ( 
.A(n_550),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_522),
.Y(n_580)
);

NOR3xp33_ASAP7_75t_SL g581 ( 
.A(n_520),
.B(n_457),
.C(n_489),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_526),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_L g583 ( 
.A(n_533),
.B(n_477),
.Y(n_583)
);

INVx4_ASAP7_75t_L g584 ( 
.A(n_517),
.Y(n_584)
);

BUFx3_ASAP7_75t_L g585 ( 
.A(n_540),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_L g586 ( 
.A(n_520),
.B(n_478),
.Y(n_586)
);

BUFx2_ASAP7_75t_L g587 ( 
.A(n_540),
.Y(n_587)
);

NOR3xp33_ASAP7_75t_SL g588 ( 
.A(n_539),
.B(n_436),
.C(n_472),
.Y(n_588)
);

OR2x6_ASAP7_75t_L g589 ( 
.A(n_517),
.B(n_476),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_SL g590 ( 
.A(n_547),
.B(n_431),
.Y(n_590)
);

NAND3xp33_ASAP7_75t_SL g591 ( 
.A(n_571),
.B(n_441),
.C(n_432),
.Y(n_591)
);

CKINVDCx20_ASAP7_75t_R g592 ( 
.A(n_544),
.Y(n_592)
);

AO21x2_ASAP7_75t_L g593 ( 
.A1(n_554),
.A2(n_464),
.B(n_482),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_545),
.Y(n_594)
);

AND2x4_ASAP7_75t_L g595 ( 
.A(n_527),
.B(n_499),
.Y(n_595)
);

INVx4_ASAP7_75t_L g596 ( 
.A(n_564),
.Y(n_596)
);

INVxp67_ASAP7_75t_SL g597 ( 
.A(n_527),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_558),
.Y(n_598)
);

HB1xp67_ASAP7_75t_L g599 ( 
.A(n_544),
.Y(n_599)
);

BUFx3_ASAP7_75t_L g600 ( 
.A(n_561),
.Y(n_600)
);

HB1xp67_ASAP7_75t_L g601 ( 
.A(n_518),
.Y(n_601)
);

NOR3xp33_ASAP7_75t_SL g602 ( 
.A(n_560),
.B(n_505),
.C(n_476),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_566),
.Y(n_603)
);

INVx2_ASAP7_75t_L g604 ( 
.A(n_548),
.Y(n_604)
);

INVx3_ASAP7_75t_SL g605 ( 
.A(n_524),
.Y(n_605)
);

INVx2_ASAP7_75t_SL g606 ( 
.A(n_561),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_L g607 ( 
.A(n_532),
.B(n_488),
.Y(n_607)
);

BUFx3_ASAP7_75t_L g608 ( 
.A(n_564),
.Y(n_608)
);

BUFx6f_ASAP7_75t_L g609 ( 
.A(n_564),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_L g610 ( 
.A(n_547),
.B(n_490),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_570),
.Y(n_611)
);

OR2x6_ASAP7_75t_L g612 ( 
.A(n_515),
.B(n_514),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_574),
.Y(n_613)
);

INVx2_ASAP7_75t_L g614 ( 
.A(n_556),
.Y(n_614)
);

NOR3xp33_ASAP7_75t_SL g615 ( 
.A(n_563),
.B(n_433),
.C(n_350),
.Y(n_615)
);

CKINVDCx5p33_ASAP7_75t_R g616 ( 
.A(n_564),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_L g617 ( 
.A(n_565),
.B(n_493),
.Y(n_617)
);

AND2x4_ASAP7_75t_L g618 ( 
.A(n_515),
.B(n_495),
.Y(n_618)
);

AND2x4_ASAP7_75t_L g619 ( 
.A(n_514),
.B(n_502),
.Y(n_619)
);

NOR3xp33_ASAP7_75t_SL g620 ( 
.A(n_565),
.B(n_316),
.C(n_306),
.Y(n_620)
);

AND2x4_ASAP7_75t_L g621 ( 
.A(n_530),
.B(n_503),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_L g622 ( 
.A(n_541),
.B(n_504),
.Y(n_622)
);

INVx2_ASAP7_75t_L g623 ( 
.A(n_562),
.Y(n_623)
);

BUFx6f_ASAP7_75t_L g624 ( 
.A(n_523),
.Y(n_624)
);

INVx3_ASAP7_75t_L g625 ( 
.A(n_513),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_528),
.Y(n_626)
);

INVx2_ASAP7_75t_SL g627 ( 
.A(n_530),
.Y(n_627)
);

AO22x1_ASAP7_75t_L g628 ( 
.A1(n_529),
.A2(n_491),
.B1(n_431),
.B2(n_484),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_538),
.Y(n_629)
);

AND2x4_ASAP7_75t_L g630 ( 
.A(n_536),
.B(n_507),
.Y(n_630)
);

HB1xp67_ASAP7_75t_L g631 ( 
.A(n_557),
.Y(n_631)
);

A2O1A1Ixp33_ASAP7_75t_L g632 ( 
.A1(n_586),
.A2(n_534),
.B(n_553),
.C(n_551),
.Y(n_632)
);

OAI21xp5_ASAP7_75t_L g633 ( 
.A1(n_617),
.A2(n_464),
.B(n_554),
.Y(n_633)
);

OAI21x1_ASAP7_75t_L g634 ( 
.A1(n_576),
.A2(n_546),
.B(n_573),
.Y(n_634)
);

OAI21xp5_ASAP7_75t_L g635 ( 
.A1(n_617),
.A2(n_572),
.B(n_569),
.Y(n_635)
);

AOI21x1_ASAP7_75t_L g636 ( 
.A1(n_590),
.A2(n_573),
.B(n_542),
.Y(n_636)
);

OAI21x1_ASAP7_75t_L g637 ( 
.A1(n_576),
.A2(n_525),
.B(n_535),
.Y(n_637)
);

A2O1A1Ixp33_ASAP7_75t_L g638 ( 
.A1(n_586),
.A2(n_531),
.B(n_567),
.C(n_552),
.Y(n_638)
);

INVx3_ASAP7_75t_SL g639 ( 
.A(n_605),
.Y(n_639)
);

O2A1O1Ixp5_ASAP7_75t_L g640 ( 
.A1(n_610),
.A2(n_525),
.B(n_543),
.C(n_542),
.Y(n_640)
);

AOI21xp5_ASAP7_75t_L g641 ( 
.A1(n_583),
.A2(n_535),
.B(n_559),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_575),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_580),
.Y(n_643)
);

OAI21xp5_ASAP7_75t_L g644 ( 
.A1(n_583),
.A2(n_552),
.B(n_567),
.Y(n_644)
);

OAI21x1_ASAP7_75t_L g645 ( 
.A1(n_622),
.A2(n_513),
.B(n_508),
.Y(n_645)
);

OAI22x1_ASAP7_75t_L g646 ( 
.A1(n_619),
.A2(n_481),
.B1(n_501),
.B2(n_491),
.Y(n_646)
);

NOR2xp33_ASAP7_75t_L g647 ( 
.A(n_592),
.B(n_306),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_L g648 ( 
.A(n_601),
.B(n_327),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_L g649 ( 
.A(n_610),
.B(n_531),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_L g650 ( 
.A(n_607),
.B(n_568),
.Y(n_650)
);

OAI21x1_ASAP7_75t_L g651 ( 
.A1(n_622),
.A2(n_384),
.B(n_383),
.Y(n_651)
);

OAI21x1_ASAP7_75t_L g652 ( 
.A1(n_625),
.A2(n_384),
.B(n_383),
.Y(n_652)
);

AOI21xp5_ASAP7_75t_L g653 ( 
.A1(n_593),
.A2(n_549),
.B(n_555),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_582),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_L g655 ( 
.A(n_607),
.B(n_327),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_L g656 ( 
.A(n_597),
.B(n_316),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_594),
.Y(n_657)
);

AOI21xp5_ASAP7_75t_L g658 ( 
.A1(n_593),
.A2(n_549),
.B(n_371),
.Y(n_658)
);

AOI21xp5_ASAP7_75t_L g659 ( 
.A1(n_630),
.A2(n_387),
.B(n_385),
.Y(n_659)
);

INVxp67_ASAP7_75t_SL g660 ( 
.A(n_597),
.Y(n_660)
);

BUFx4f_ASAP7_75t_L g661 ( 
.A(n_595),
.Y(n_661)
);

OAI22xp5_ASAP7_75t_L g662 ( 
.A1(n_581),
.A2(n_318),
.B1(n_364),
.B2(n_382),
.Y(n_662)
);

OAI21xp5_ASAP7_75t_L g663 ( 
.A1(n_620),
.A2(n_357),
.B(n_356),
.Y(n_663)
);

OAI21x1_ASAP7_75t_L g664 ( 
.A1(n_625),
.A2(n_387),
.B(n_385),
.Y(n_664)
);

INVx2_ASAP7_75t_SL g665 ( 
.A(n_579),
.Y(n_665)
);

NOR2xp33_ASAP7_75t_L g666 ( 
.A(n_591),
.B(n_318),
.Y(n_666)
);

OAI21x1_ASAP7_75t_L g667 ( 
.A1(n_598),
.A2(n_361),
.B(n_357),
.Y(n_667)
);

INVx2_ASAP7_75t_L g668 ( 
.A(n_604),
.Y(n_668)
);

AND2x2_ASAP7_75t_L g669 ( 
.A(n_599),
.B(n_322),
.Y(n_669)
);

BUFx8_ASAP7_75t_L g670 ( 
.A(n_587),
.Y(n_670)
);

A2O1A1Ixp33_ASAP7_75t_L g671 ( 
.A1(n_615),
.A2(n_382),
.B(n_379),
.C(n_378),
.Y(n_671)
);

NOR2xp33_ASAP7_75t_L g672 ( 
.A(n_591),
.B(n_194),
.Y(n_672)
);

INVxp67_ASAP7_75t_SL g673 ( 
.A(n_618),
.Y(n_673)
);

OAI22x1_ASAP7_75t_L g674 ( 
.A1(n_619),
.A2(n_322),
.B1(n_378),
.B2(n_377),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_L g675 ( 
.A(n_577),
.B(n_321),
.Y(n_675)
);

HB1xp67_ASAP7_75t_L g676 ( 
.A(n_618),
.Y(n_676)
);

AND2x2_ASAP7_75t_L g677 ( 
.A(n_595),
.B(n_322),
.Y(n_677)
);

AND2x4_ASAP7_75t_L g678 ( 
.A(n_584),
.B(n_361),
.Y(n_678)
);

INVx2_ASAP7_75t_L g679 ( 
.A(n_614),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_SL g680 ( 
.A(n_581),
.B(n_363),
.Y(n_680)
);

OAI21xp5_ASAP7_75t_L g681 ( 
.A1(n_603),
.A2(n_364),
.B(n_363),
.Y(n_681)
);

OAI21x1_ASAP7_75t_L g682 ( 
.A1(n_611),
.A2(n_377),
.B(n_365),
.Y(n_682)
);

INVxp67_ASAP7_75t_L g683 ( 
.A(n_585),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_631),
.B(n_379),
.Y(n_684)
);

OAI21x1_ASAP7_75t_L g685 ( 
.A1(n_613),
.A2(n_365),
.B(n_322),
.Y(n_685)
);

AOI21xp33_ASAP7_75t_L g686 ( 
.A1(n_612),
.A2(n_199),
.B(n_198),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_623),
.Y(n_687)
);

OAI21xp5_ASAP7_75t_L g688 ( 
.A1(n_630),
.A2(n_621),
.B(n_626),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_L g689 ( 
.A(n_647),
.B(n_676),
.Y(n_689)
);

AO22x2_ASAP7_75t_L g690 ( 
.A1(n_660),
.A2(n_629),
.B1(n_621),
.B2(n_606),
.Y(n_690)
);

AOI22xp33_ASAP7_75t_L g691 ( 
.A1(n_644),
.A2(n_612),
.B1(n_589),
.B2(n_584),
.Y(n_691)
);

INVx2_ASAP7_75t_L g692 ( 
.A(n_668),
.Y(n_692)
);

OAI22x1_ASAP7_75t_L g693 ( 
.A1(n_666),
.A2(n_627),
.B1(n_616),
.B2(n_602),
.Y(n_693)
);

OR2x2_ASAP7_75t_L g694 ( 
.A(n_642),
.B(n_600),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_L g695 ( 
.A(n_673),
.B(n_588),
.Y(n_695)
);

OAI21x1_ASAP7_75t_L g696 ( 
.A1(n_651),
.A2(n_596),
.B(n_609),
.Y(n_696)
);

AOI31xp67_ASAP7_75t_L g697 ( 
.A1(n_680),
.A2(n_649),
.A3(n_650),
.B(n_655),
.Y(n_697)
);

BUFx5_ASAP7_75t_L g698 ( 
.A(n_643),
.Y(n_698)
);

INVx2_ASAP7_75t_L g699 ( 
.A(n_679),
.Y(n_699)
);

OAI21xp5_ASAP7_75t_L g700 ( 
.A1(n_632),
.A2(n_640),
.B(n_641),
.Y(n_700)
);

OAI21xp5_ASAP7_75t_L g701 ( 
.A1(n_637),
.A2(n_612),
.B(n_596),
.Y(n_701)
);

BUFx6f_ASAP7_75t_L g702 ( 
.A(n_661),
.Y(n_702)
);

AOI21xp5_ASAP7_75t_L g703 ( 
.A1(n_638),
.A2(n_609),
.B(n_589),
.Y(n_703)
);

O2A1O1Ixp33_ASAP7_75t_SL g704 ( 
.A1(n_650),
.A2(n_628),
.B(n_3),
.C(n_4),
.Y(n_704)
);

NOR2xp67_ASAP7_75t_SL g705 ( 
.A(n_665),
.B(n_578),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_654),
.Y(n_706)
);

INVx2_ASAP7_75t_L g707 ( 
.A(n_687),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_657),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_669),
.Y(n_709)
);

OAI21x1_ASAP7_75t_L g710 ( 
.A1(n_634),
.A2(n_609),
.B(n_608),
.Y(n_710)
);

NOR2xp33_ASAP7_75t_L g711 ( 
.A(n_683),
.B(n_579),
.Y(n_711)
);

A2O1A1Ixp33_ASAP7_75t_L g712 ( 
.A1(n_644),
.A2(n_624),
.B(n_226),
.C(n_239),
.Y(n_712)
);

BUFx2_ASAP7_75t_L g713 ( 
.A(n_670),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_L g714 ( 
.A(n_649),
.B(n_589),
.Y(n_714)
);

AND2x4_ASAP7_75t_L g715 ( 
.A(n_688),
.B(n_624),
.Y(n_715)
);

AND2x2_ASAP7_75t_L g716 ( 
.A(n_661),
.B(n_1),
.Y(n_716)
);

A2O1A1Ixp33_ASAP7_75t_L g717 ( 
.A1(n_672),
.A2(n_653),
.B(n_686),
.C(n_675),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_656),
.Y(n_718)
);

AO21x2_ASAP7_75t_L g719 ( 
.A1(n_633),
.A2(n_658),
.B(n_681),
.Y(n_719)
);

INVxp67_ASAP7_75t_L g720 ( 
.A(n_670),
.Y(n_720)
);

AO31x2_ASAP7_75t_L g721 ( 
.A1(n_674),
.A2(n_624),
.A3(n_116),
.B(n_117),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_L g722 ( 
.A(n_648),
.B(n_3),
.Y(n_722)
);

AOI21xp5_ASAP7_75t_L g723 ( 
.A1(n_633),
.A2(n_204),
.B(n_202),
.Y(n_723)
);

AOI21xp5_ASAP7_75t_L g724 ( 
.A1(n_635),
.A2(n_211),
.B(n_209),
.Y(n_724)
);

NOR2xp33_ASAP7_75t_L g725 ( 
.A(n_639),
.B(n_4),
.Y(n_725)
);

BUFx10_ASAP7_75t_L g726 ( 
.A(n_678),
.Y(n_726)
);

AOI221xp5_ASAP7_75t_L g727 ( 
.A1(n_686),
.A2(n_238),
.B1(n_229),
.B2(n_228),
.C(n_227),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_L g728 ( 
.A(n_677),
.B(n_5),
.Y(n_728)
);

AO31x2_ASAP7_75t_L g729 ( 
.A1(n_671),
.A2(n_108),
.A3(n_178),
.B(n_177),
.Y(n_729)
);

NOR2xp33_ASAP7_75t_L g730 ( 
.A(n_678),
.B(n_5),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_684),
.Y(n_731)
);

BUFx2_ASAP7_75t_L g732 ( 
.A(n_688),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_685),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_636),
.Y(n_734)
);

AOI22xp5_ASAP7_75t_L g735 ( 
.A1(n_646),
.A2(n_220),
.B1(n_218),
.B2(n_214),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_667),
.Y(n_736)
);

BUFx3_ASAP7_75t_L g737 ( 
.A(n_645),
.Y(n_737)
);

OR2x2_ASAP7_75t_L g738 ( 
.A(n_681),
.B(n_6),
.Y(n_738)
);

INVx3_ASAP7_75t_L g739 ( 
.A(n_682),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_L g740 ( 
.A(n_662),
.B(n_6),
.Y(n_740)
);

OAI22xp33_ASAP7_75t_L g741 ( 
.A1(n_662),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_741)
);

INVx1_ASAP7_75t_SL g742 ( 
.A(n_659),
.Y(n_742)
);

OAI21x1_ASAP7_75t_L g743 ( 
.A1(n_652),
.A2(n_32),
.B(n_31),
.Y(n_743)
);

OAI21x1_ASAP7_75t_SL g744 ( 
.A1(n_663),
.A2(n_7),
.B(n_8),
.Y(n_744)
);

OAI21x1_ASAP7_75t_L g745 ( 
.A1(n_664),
.A2(n_34),
.B(n_33),
.Y(n_745)
);

AOI21xp33_ASAP7_75t_L g746 ( 
.A1(n_663),
.A2(n_10),
.B(n_11),
.Y(n_746)
);

CKINVDCx5p33_ASAP7_75t_R g747 ( 
.A(n_635),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_642),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_642),
.Y(n_749)
);

OAI21x1_ASAP7_75t_L g750 ( 
.A1(n_651),
.A2(n_37),
.B(n_36),
.Y(n_750)
);

AO31x2_ASAP7_75t_L g751 ( 
.A1(n_674),
.A2(n_115),
.A3(n_176),
.B(n_175),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_L g752 ( 
.A(n_647),
.B(n_10),
.Y(n_752)
);

OAI21x1_ASAP7_75t_L g753 ( 
.A1(n_651),
.A2(n_41),
.B(n_40),
.Y(n_753)
);

BUFx2_ASAP7_75t_L g754 ( 
.A(n_670),
.Y(n_754)
);

AOI21xp5_ASAP7_75t_L g755 ( 
.A1(n_632),
.A2(n_12),
.B(n_13),
.Y(n_755)
);

INVxp67_ASAP7_75t_SL g756 ( 
.A(n_660),
.Y(n_756)
);

BUFx12f_ASAP7_75t_L g757 ( 
.A(n_713),
.Y(n_757)
);

OAI22xp33_ASAP7_75t_L g758 ( 
.A1(n_752),
.A2(n_13),
.B1(n_14),
.B2(n_15),
.Y(n_758)
);

INVx8_ASAP7_75t_L g759 ( 
.A(n_702),
.Y(n_759)
);

OAI22xp5_ASAP7_75t_L g760 ( 
.A1(n_747),
.A2(n_15),
.B1(n_16),
.B2(n_17),
.Y(n_760)
);

AOI22xp5_ASAP7_75t_L g761 ( 
.A1(n_741),
.A2(n_740),
.B1(n_689),
.B2(n_691),
.Y(n_761)
);

INVx6_ASAP7_75t_L g762 ( 
.A(n_702),
.Y(n_762)
);

AND2x4_ASAP7_75t_L g763 ( 
.A(n_756),
.B(n_42),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_L g764 ( 
.A(n_718),
.B(n_16),
.Y(n_764)
);

BUFx4_ASAP7_75t_SL g765 ( 
.A(n_754),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_L g766 ( 
.A(n_731),
.B(n_706),
.Y(n_766)
);

INVx1_ASAP7_75t_SL g767 ( 
.A(n_732),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_708),
.Y(n_768)
);

AOI22xp33_ASAP7_75t_L g769 ( 
.A1(n_690),
.A2(n_17),
.B1(n_18),
.B2(n_19),
.Y(n_769)
);

AOI22xp33_ASAP7_75t_L g770 ( 
.A1(n_690),
.A2(n_18),
.B1(n_19),
.B2(n_20),
.Y(n_770)
);

AOI22xp33_ASAP7_75t_L g771 ( 
.A1(n_695),
.A2(n_21),
.B1(n_22),
.B2(n_23),
.Y(n_771)
);

INVx6_ASAP7_75t_L g772 ( 
.A(n_702),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_748),
.Y(n_773)
);

CKINVDCx6p67_ASAP7_75t_R g774 ( 
.A(n_693),
.Y(n_774)
);

CKINVDCx20_ASAP7_75t_R g775 ( 
.A(n_720),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_749),
.Y(n_776)
);

AOI22xp33_ASAP7_75t_SL g777 ( 
.A1(n_744),
.A2(n_21),
.B1(n_25),
.B2(n_26),
.Y(n_777)
);

CKINVDCx11_ASAP7_75t_R g778 ( 
.A(n_726),
.Y(n_778)
);

INVx2_ASAP7_75t_L g779 ( 
.A(n_707),
.Y(n_779)
);

AOI22xp5_ASAP7_75t_L g780 ( 
.A1(n_714),
.A2(n_26),
.B1(n_28),
.B2(n_29),
.Y(n_780)
);

CKINVDCx5p33_ASAP7_75t_R g781 ( 
.A(n_711),
.Y(n_781)
);

BUFx12f_ASAP7_75t_L g782 ( 
.A(n_694),
.Y(n_782)
);

INVx2_ASAP7_75t_L g783 ( 
.A(n_692),
.Y(n_783)
);

INVx2_ASAP7_75t_L g784 ( 
.A(n_699),
.Y(n_784)
);

INVx2_ASAP7_75t_L g785 ( 
.A(n_734),
.Y(n_785)
);

OAI22xp5_ASAP7_75t_L g786 ( 
.A1(n_755),
.A2(n_28),
.B1(n_29),
.B2(n_30),
.Y(n_786)
);

INVx8_ASAP7_75t_L g787 ( 
.A(n_715),
.Y(n_787)
);

BUFx2_ASAP7_75t_SL g788 ( 
.A(n_716),
.Y(n_788)
);

AOI22xp33_ASAP7_75t_SL g789 ( 
.A1(n_700),
.A2(n_30),
.B1(n_44),
.B2(n_45),
.Y(n_789)
);

AOI22xp33_ASAP7_75t_L g790 ( 
.A1(n_709),
.A2(n_50),
.B1(n_52),
.B2(n_53),
.Y(n_790)
);

BUFx12f_ASAP7_75t_L g791 ( 
.A(n_726),
.Y(n_791)
);

AOI22xp33_ASAP7_75t_L g792 ( 
.A1(n_715),
.A2(n_54),
.B1(n_55),
.B2(n_57),
.Y(n_792)
);

BUFx6f_ASAP7_75t_SL g793 ( 
.A(n_705),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_698),
.Y(n_794)
);

BUFx2_ASAP7_75t_L g795 ( 
.A(n_698),
.Y(n_795)
);

INVx2_ASAP7_75t_L g796 ( 
.A(n_698),
.Y(n_796)
);

AOI22xp33_ASAP7_75t_L g797 ( 
.A1(n_703),
.A2(n_60),
.B1(n_61),
.B2(n_62),
.Y(n_797)
);

BUFx2_ASAP7_75t_SL g798 ( 
.A(n_698),
.Y(n_798)
);

AOI22xp5_ASAP7_75t_L g799 ( 
.A1(n_704),
.A2(n_63),
.B1(n_67),
.B2(n_69),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_697),
.Y(n_800)
);

CKINVDCx20_ASAP7_75t_R g801 ( 
.A(n_735),
.Y(n_801)
);

INVx1_ASAP7_75t_SL g802 ( 
.A(n_742),
.Y(n_802)
);

CKINVDCx6p67_ASAP7_75t_R g803 ( 
.A(n_728),
.Y(n_803)
);

AOI22xp33_ASAP7_75t_L g804 ( 
.A1(n_746),
.A2(n_70),
.B1(n_71),
.B2(n_73),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_738),
.Y(n_805)
);

BUFx2_ASAP7_75t_L g806 ( 
.A(n_701),
.Y(n_806)
);

AOI22xp33_ASAP7_75t_L g807 ( 
.A1(n_723),
.A2(n_74),
.B1(n_75),
.B2(n_76),
.Y(n_807)
);

CKINVDCx6p67_ASAP7_75t_R g808 ( 
.A(n_722),
.Y(n_808)
);

CKINVDCx11_ASAP7_75t_R g809 ( 
.A(n_737),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_733),
.Y(n_810)
);

AOI22xp33_ASAP7_75t_SL g811 ( 
.A1(n_730),
.A2(n_77),
.B1(n_78),
.B2(n_79),
.Y(n_811)
);

BUFx2_ASAP7_75t_L g812 ( 
.A(n_710),
.Y(n_812)
);

OAI21xp5_ASAP7_75t_SL g813 ( 
.A1(n_725),
.A2(n_80),
.B(n_81),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_736),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_L g815 ( 
.A(n_717),
.B(n_719),
.Y(n_815)
);

BUFx2_ASAP7_75t_SL g816 ( 
.A(n_739),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_721),
.Y(n_817)
);

INVx2_ASAP7_75t_L g818 ( 
.A(n_721),
.Y(n_818)
);

INVx2_ASAP7_75t_L g819 ( 
.A(n_810),
.Y(n_819)
);

AOI221xp5_ASAP7_75t_L g820 ( 
.A1(n_758),
.A2(n_727),
.B1(n_712),
.B2(n_724),
.C(n_739),
.Y(n_820)
);

OAI21x1_ASAP7_75t_L g821 ( 
.A1(n_815),
.A2(n_696),
.B(n_753),
.Y(n_821)
);

INVx2_ASAP7_75t_L g822 ( 
.A(n_785),
.Y(n_822)
);

INVx3_ASAP7_75t_L g823 ( 
.A(n_796),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_768),
.Y(n_824)
);

HB1xp67_ASAP7_75t_L g825 ( 
.A(n_767),
.Y(n_825)
);

AOI22xp33_ASAP7_75t_SL g826 ( 
.A1(n_801),
.A2(n_721),
.B1(n_751),
.B2(n_729),
.Y(n_826)
);

OAI21x1_ASAP7_75t_L g827 ( 
.A1(n_800),
.A2(n_818),
.B(n_817),
.Y(n_827)
);

OAI22xp33_ASAP7_75t_L g828 ( 
.A1(n_813),
.A2(n_729),
.B1(n_751),
.B2(n_745),
.Y(n_828)
);

OA21x2_ASAP7_75t_L g829 ( 
.A1(n_812),
.A2(n_814),
.B(n_794),
.Y(n_829)
);

OR2x2_ASAP7_75t_L g830 ( 
.A(n_767),
.B(n_802),
.Y(n_830)
);

INVx2_ASAP7_75t_L g831 ( 
.A(n_779),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_773),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_776),
.Y(n_833)
);

HB1xp67_ASAP7_75t_L g834 ( 
.A(n_805),
.Y(n_834)
);

NOR2xp33_ASAP7_75t_L g835 ( 
.A(n_781),
.B(n_82),
.Y(n_835)
);

BUFx6f_ASAP7_75t_L g836 ( 
.A(n_809),
.Y(n_836)
);

AO21x2_ASAP7_75t_L g837 ( 
.A1(n_799),
.A2(n_750),
.B(n_743),
.Y(n_837)
);

HB1xp67_ASAP7_75t_L g838 ( 
.A(n_802),
.Y(n_838)
);

INVx2_ASAP7_75t_L g839 ( 
.A(n_783),
.Y(n_839)
);

INVx2_ASAP7_75t_L g840 ( 
.A(n_784),
.Y(n_840)
);

AND2x2_ASAP7_75t_L g841 ( 
.A(n_795),
.B(n_751),
.Y(n_841)
);

OR2x6_ASAP7_75t_L g842 ( 
.A(n_806),
.B(n_729),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_766),
.Y(n_843)
);

NOR2xp33_ASAP7_75t_R g844 ( 
.A(n_775),
.B(n_83),
.Y(n_844)
);

OAI21x1_ASAP7_75t_L g845 ( 
.A1(n_797),
.A2(n_85),
.B(n_86),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_798),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_816),
.Y(n_847)
);

INVx2_ASAP7_75t_L g848 ( 
.A(n_787),
.Y(n_848)
);

OAI21x1_ASAP7_75t_L g849 ( 
.A1(n_799),
.A2(n_790),
.B(n_792),
.Y(n_849)
);

INVx3_ASAP7_75t_L g850 ( 
.A(n_763),
.Y(n_850)
);

BUFx2_ASAP7_75t_L g851 ( 
.A(n_763),
.Y(n_851)
);

HB1xp67_ASAP7_75t_L g852 ( 
.A(n_764),
.Y(n_852)
);

INVx1_ASAP7_75t_L g853 ( 
.A(n_787),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_L g854 ( 
.A(n_808),
.B(n_87),
.Y(n_854)
);

NAND2x1p5_ASAP7_75t_L g855 ( 
.A(n_761),
.B(n_780),
.Y(n_855)
);

BUFx2_ASAP7_75t_L g856 ( 
.A(n_791),
.Y(n_856)
);

BUFx2_ASAP7_75t_L g857 ( 
.A(n_774),
.Y(n_857)
);

INVx2_ASAP7_75t_L g858 ( 
.A(n_787),
.Y(n_858)
);

OAI21x1_ASAP7_75t_L g859 ( 
.A1(n_807),
.A2(n_770),
.B(n_769),
.Y(n_859)
);

INVx1_ASAP7_75t_L g860 ( 
.A(n_761),
.Y(n_860)
);

INVx1_ASAP7_75t_L g861 ( 
.A(n_780),
.Y(n_861)
);

INVx1_ASAP7_75t_L g862 ( 
.A(n_788),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_786),
.Y(n_863)
);

INVx2_ASAP7_75t_L g864 ( 
.A(n_782),
.Y(n_864)
);

OAI22xp33_ASAP7_75t_L g865 ( 
.A1(n_813),
.A2(n_90),
.B1(n_91),
.B2(n_92),
.Y(n_865)
);

AND2x2_ASAP7_75t_L g866 ( 
.A(n_803),
.B(n_94),
.Y(n_866)
);

INVx2_ASAP7_75t_L g867 ( 
.A(n_762),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_819),
.Y(n_868)
);

INVx2_ASAP7_75t_SL g869 ( 
.A(n_830),
.Y(n_869)
);

AO21x2_ASAP7_75t_L g870 ( 
.A1(n_828),
.A2(n_827),
.B(n_821),
.Y(n_870)
);

OR2x2_ASAP7_75t_L g871 ( 
.A(n_830),
.B(n_760),
.Y(n_871)
);

OR2x2_ASAP7_75t_L g872 ( 
.A(n_838),
.B(n_771),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_L g873 ( 
.A(n_825),
.B(n_834),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_L g874 ( 
.A(n_843),
.B(n_778),
.Y(n_874)
);

HB1xp67_ASAP7_75t_L g875 ( 
.A(n_824),
.Y(n_875)
);

INVx2_ASAP7_75t_SL g876 ( 
.A(n_851),
.Y(n_876)
);

HB1xp67_ASAP7_75t_L g877 ( 
.A(n_824),
.Y(n_877)
);

CKINVDCx6p67_ASAP7_75t_R g878 ( 
.A(n_836),
.Y(n_878)
);

AOI222xp33_ASAP7_75t_L g879 ( 
.A1(n_861),
.A2(n_793),
.B1(n_804),
.B2(n_757),
.C1(n_777),
.C2(n_772),
.Y(n_879)
);

AND2x2_ASAP7_75t_L g880 ( 
.A(n_841),
.B(n_789),
.Y(n_880)
);

AND2x2_ASAP7_75t_L g881 ( 
.A(n_841),
.B(n_762),
.Y(n_881)
);

AOI22xp33_ASAP7_75t_L g882 ( 
.A1(n_855),
.A2(n_793),
.B1(n_811),
.B2(n_772),
.Y(n_882)
);

AND2x2_ASAP7_75t_L g883 ( 
.A(n_851),
.B(n_823),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_819),
.Y(n_884)
);

INVx2_ASAP7_75t_L g885 ( 
.A(n_819),
.Y(n_885)
);

HB1xp67_ASAP7_75t_L g886 ( 
.A(n_832),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_832),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_833),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_L g889 ( 
.A(n_843),
.B(n_759),
.Y(n_889)
);

OA21x2_ASAP7_75t_L g890 ( 
.A1(n_827),
.A2(n_759),
.B(n_96),
.Y(n_890)
);

INVx1_ASAP7_75t_L g891 ( 
.A(n_833),
.Y(n_891)
);

OA21x2_ASAP7_75t_L g892 ( 
.A1(n_821),
.A2(n_759),
.B(n_97),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_822),
.Y(n_893)
);

AND2x2_ASAP7_75t_L g894 ( 
.A(n_823),
.B(n_829),
.Y(n_894)
);

INVx1_ASAP7_75t_L g895 ( 
.A(n_822),
.Y(n_895)
);

OR2x2_ASAP7_75t_L g896 ( 
.A(n_860),
.B(n_765),
.Y(n_896)
);

BUFx3_ASAP7_75t_L g897 ( 
.A(n_836),
.Y(n_897)
);

INVx1_ASAP7_75t_L g898 ( 
.A(n_829),
.Y(n_898)
);

INVx2_ASAP7_75t_L g899 ( 
.A(n_829),
.Y(n_899)
);

BUFx3_ASAP7_75t_L g900 ( 
.A(n_897),
.Y(n_900)
);

INVxp67_ASAP7_75t_SL g901 ( 
.A(n_899),
.Y(n_901)
);

AND2x2_ASAP7_75t_L g902 ( 
.A(n_894),
.B(n_883),
.Y(n_902)
);

INVx2_ASAP7_75t_L g903 ( 
.A(n_899),
.Y(n_903)
);

INVx1_ASAP7_75t_SL g904 ( 
.A(n_883),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_L g905 ( 
.A(n_875),
.B(n_829),
.Y(n_905)
);

HB1xp67_ASAP7_75t_L g906 ( 
.A(n_869),
.Y(n_906)
);

INVxp67_ASAP7_75t_SL g907 ( 
.A(n_899),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_868),
.Y(n_908)
);

INVx2_ASAP7_75t_L g909 ( 
.A(n_898),
.Y(n_909)
);

OAI222xp33_ASAP7_75t_L g910 ( 
.A1(n_880),
.A2(n_855),
.B1(n_861),
.B2(n_860),
.C1(n_826),
.C2(n_842),
.Y(n_910)
);

INVx2_ASAP7_75t_SL g911 ( 
.A(n_894),
.Y(n_911)
);

INVx3_ASAP7_75t_L g912 ( 
.A(n_870),
.Y(n_912)
);

AND2x2_ASAP7_75t_L g913 ( 
.A(n_876),
.B(n_862),
.Y(n_913)
);

AND2x2_ASAP7_75t_L g914 ( 
.A(n_876),
.B(n_823),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_L g915 ( 
.A(n_877),
.B(n_852),
.Y(n_915)
);

BUFx3_ASAP7_75t_L g916 ( 
.A(n_897),
.Y(n_916)
);

AND2x2_ASAP7_75t_L g917 ( 
.A(n_869),
.B(n_823),
.Y(n_917)
);

BUFx2_ASAP7_75t_L g918 ( 
.A(n_897),
.Y(n_918)
);

NAND2xp5_ASAP7_75t_L g919 ( 
.A(n_886),
.B(n_847),
.Y(n_919)
);

INVx2_ASAP7_75t_SL g920 ( 
.A(n_898),
.Y(n_920)
);

INVx2_ASAP7_75t_L g921 ( 
.A(n_885),
.Y(n_921)
);

HB1xp67_ASAP7_75t_L g922 ( 
.A(n_873),
.Y(n_922)
);

HB1xp67_ASAP7_75t_L g923 ( 
.A(n_922),
.Y(n_923)
);

INVx2_ASAP7_75t_L g924 ( 
.A(n_920),
.Y(n_924)
);

INVx2_ASAP7_75t_L g925 ( 
.A(n_920),
.Y(n_925)
);

INVx1_ASAP7_75t_L g926 ( 
.A(n_915),
.Y(n_926)
);

HB1xp67_ASAP7_75t_L g927 ( 
.A(n_906),
.Y(n_927)
);

AOI22xp5_ASAP7_75t_L g928 ( 
.A1(n_912),
.A2(n_855),
.B1(n_880),
.B2(n_879),
.Y(n_928)
);

INVx1_ASAP7_75t_L g929 ( 
.A(n_915),
.Y(n_929)
);

AND2x2_ASAP7_75t_L g930 ( 
.A(n_918),
.B(n_874),
.Y(n_930)
);

AND2x2_ASAP7_75t_L g931 ( 
.A(n_918),
.B(n_878),
.Y(n_931)
);

HB1xp67_ASAP7_75t_L g932 ( 
.A(n_919),
.Y(n_932)
);

INVx1_ASAP7_75t_L g933 ( 
.A(n_919),
.Y(n_933)
);

BUFx2_ASAP7_75t_L g934 ( 
.A(n_900),
.Y(n_934)
);

OR2x2_ASAP7_75t_L g935 ( 
.A(n_904),
.B(n_887),
.Y(n_935)
);

INVx1_ASAP7_75t_L g936 ( 
.A(n_908),
.Y(n_936)
);

AND2x2_ASAP7_75t_L g937 ( 
.A(n_904),
.B(n_878),
.Y(n_937)
);

INVx4_ASAP7_75t_L g938 ( 
.A(n_900),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_L g939 ( 
.A(n_913),
.B(n_887),
.Y(n_939)
);

NOR2xp33_ASAP7_75t_SL g940 ( 
.A(n_910),
.B(n_836),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_L g941 ( 
.A(n_933),
.B(n_908),
.Y(n_941)
);

OR2x2_ASAP7_75t_L g942 ( 
.A(n_926),
.B(n_871),
.Y(n_942)
);

INVxp67_ASAP7_75t_L g943 ( 
.A(n_934),
.Y(n_943)
);

NAND2xp5_ASAP7_75t_L g944 ( 
.A(n_929),
.B(n_932),
.Y(n_944)
);

AND2x4_ASAP7_75t_L g945 ( 
.A(n_930),
.B(n_836),
.Y(n_945)
);

INVx1_ASAP7_75t_L g946 ( 
.A(n_923),
.Y(n_946)
);

INVx2_ASAP7_75t_L g947 ( 
.A(n_935),
.Y(n_947)
);

INVx1_ASAP7_75t_L g948 ( 
.A(n_936),
.Y(n_948)
);

INVx2_ASAP7_75t_SL g949 ( 
.A(n_930),
.Y(n_949)
);

AND2x2_ASAP7_75t_L g950 ( 
.A(n_931),
.B(n_900),
.Y(n_950)
);

AND2x2_ASAP7_75t_L g951 ( 
.A(n_931),
.B(n_916),
.Y(n_951)
);

INVxp67_ASAP7_75t_L g952 ( 
.A(n_946),
.Y(n_952)
);

INVx2_ASAP7_75t_L g953 ( 
.A(n_945),
.Y(n_953)
);

INVxp67_ASAP7_75t_L g954 ( 
.A(n_945),
.Y(n_954)
);

HB1xp67_ASAP7_75t_L g955 ( 
.A(n_943),
.Y(n_955)
);

INVx1_ASAP7_75t_L g956 ( 
.A(n_948),
.Y(n_956)
);

OR2x2_ASAP7_75t_L g957 ( 
.A(n_942),
.B(n_944),
.Y(n_957)
);

NAND2xp5_ASAP7_75t_SL g958 ( 
.A(n_949),
.B(n_940),
.Y(n_958)
);

INVx1_ASAP7_75t_SL g959 ( 
.A(n_950),
.Y(n_959)
);

NAND2xp5_ASAP7_75t_L g960 ( 
.A(n_959),
.B(n_943),
.Y(n_960)
);

AO221x2_ASAP7_75t_L g961 ( 
.A1(n_953),
.A2(n_944),
.B1(n_910),
.B2(n_924),
.C(n_925),
.Y(n_961)
);

OAI221xp5_ASAP7_75t_L g962 ( 
.A1(n_958),
.A2(n_928),
.B1(n_912),
.B2(n_901),
.C(n_907),
.Y(n_962)
);

NAND2xp5_ASAP7_75t_L g963 ( 
.A(n_955),
.B(n_947),
.Y(n_963)
);

NAND2xp33_ASAP7_75t_SL g964 ( 
.A(n_957),
.B(n_836),
.Y(n_964)
);

AND2x4_ASAP7_75t_SL g965 ( 
.A(n_956),
.B(n_951),
.Y(n_965)
);

OAI221xp5_ASAP7_75t_L g966 ( 
.A1(n_954),
.A2(n_912),
.B1(n_907),
.B2(n_901),
.C(n_905),
.Y(n_966)
);

OR2x2_ASAP7_75t_L g967 ( 
.A(n_963),
.B(n_952),
.Y(n_967)
);

NAND2xp5_ASAP7_75t_L g968 ( 
.A(n_965),
.B(n_952),
.Y(n_968)
);

INVx1_ASAP7_75t_L g969 ( 
.A(n_960),
.Y(n_969)
);

INVx1_ASAP7_75t_SL g970 ( 
.A(n_964),
.Y(n_970)
);

AOI21xp5_ASAP7_75t_L g971 ( 
.A1(n_961),
.A2(n_934),
.B(n_912),
.Y(n_971)
);

NAND2xp5_ASAP7_75t_SL g972 ( 
.A(n_962),
.B(n_938),
.Y(n_972)
);

OR2x2_ASAP7_75t_L g973 ( 
.A(n_966),
.B(n_941),
.Y(n_973)
);

NAND2xp5_ASAP7_75t_L g974 ( 
.A(n_965),
.B(n_927),
.Y(n_974)
);

NAND2xp5_ASAP7_75t_L g975 ( 
.A(n_965),
.B(n_941),
.Y(n_975)
);

NAND2xp5_ASAP7_75t_L g976 ( 
.A(n_965),
.B(n_924),
.Y(n_976)
);

INVx1_ASAP7_75t_L g977 ( 
.A(n_963),
.Y(n_977)
);

NOR2xp33_ASAP7_75t_L g978 ( 
.A(n_970),
.B(n_938),
.Y(n_978)
);

OAI221xp5_ASAP7_75t_L g979 ( 
.A1(n_971),
.A2(n_857),
.B1(n_905),
.B2(n_854),
.C(n_920),
.Y(n_979)
);

INVx1_ASAP7_75t_L g980 ( 
.A(n_969),
.Y(n_980)
);

NAND3x2_ASAP7_75t_L g981 ( 
.A(n_967),
.B(n_857),
.C(n_856),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_L g982 ( 
.A(n_977),
.B(n_925),
.Y(n_982)
);

NOR2xp33_ASAP7_75t_L g983 ( 
.A(n_974),
.B(n_938),
.Y(n_983)
);

INVx1_ASAP7_75t_L g984 ( 
.A(n_975),
.Y(n_984)
);

OAI322xp33_ASAP7_75t_L g985 ( 
.A1(n_973),
.A2(n_871),
.A3(n_872),
.B1(n_865),
.B2(n_863),
.C1(n_896),
.C2(n_911),
.Y(n_985)
);

AOI21xp5_ASAP7_75t_L g986 ( 
.A1(n_985),
.A2(n_968),
.B(n_972),
.Y(n_986)
);

INVx1_ASAP7_75t_L g987 ( 
.A(n_982),
.Y(n_987)
);

INVx1_ASAP7_75t_L g988 ( 
.A(n_984),
.Y(n_988)
);

INVx2_ASAP7_75t_L g989 ( 
.A(n_980),
.Y(n_989)
);

AOI21xp33_ASAP7_75t_L g990 ( 
.A1(n_978),
.A2(n_976),
.B(n_835),
.Y(n_990)
);

AND2x2_ASAP7_75t_L g991 ( 
.A(n_983),
.B(n_937),
.Y(n_991)
);

OAI221xp5_ASAP7_75t_L g992 ( 
.A1(n_979),
.A2(n_862),
.B1(n_892),
.B2(n_882),
.C(n_872),
.Y(n_992)
);

OAI22xp33_ASAP7_75t_SL g993 ( 
.A1(n_988),
.A2(n_981),
.B1(n_864),
.B2(n_896),
.Y(n_993)
);

OAI321xp33_ASAP7_75t_L g994 ( 
.A1(n_986),
.A2(n_866),
.A3(n_842),
.B1(n_856),
.B2(n_864),
.C(n_820),
.Y(n_994)
);

AOI21xp5_ASAP7_75t_L g995 ( 
.A1(n_990),
.A2(n_937),
.B(n_939),
.Y(n_995)
);

AOI21xp5_ASAP7_75t_L g996 ( 
.A1(n_990),
.A2(n_911),
.B(n_935),
.Y(n_996)
);

OR2x2_ASAP7_75t_L g997 ( 
.A(n_989),
.B(n_911),
.Y(n_997)
);

AOI211xp5_ASAP7_75t_SL g998 ( 
.A1(n_987),
.A2(n_866),
.B(n_847),
.C(n_863),
.Y(n_998)
);

INVxp67_ASAP7_75t_L g999 ( 
.A(n_997),
.Y(n_999)
);

INVx1_ASAP7_75t_L g1000 ( 
.A(n_993),
.Y(n_1000)
);

BUFx2_ASAP7_75t_L g1001 ( 
.A(n_998),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_L g1002 ( 
.A(n_995),
.B(n_991),
.Y(n_1002)
);

INVx2_ASAP7_75t_L g1003 ( 
.A(n_994),
.Y(n_1003)
);

HB1xp67_ASAP7_75t_L g1004 ( 
.A(n_996),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_L g1005 ( 
.A(n_1001),
.B(n_992),
.Y(n_1005)
);

NOR2xp33_ASAP7_75t_L g1006 ( 
.A(n_1002),
.B(n_916),
.Y(n_1006)
);

NAND2xp5_ASAP7_75t_L g1007 ( 
.A(n_999),
.B(n_909),
.Y(n_1007)
);

NAND2xp5_ASAP7_75t_L g1008 ( 
.A(n_1004),
.B(n_909),
.Y(n_1008)
);

INVx1_ASAP7_75t_L g1009 ( 
.A(n_1000),
.Y(n_1009)
);

NOR3xp33_ASAP7_75t_L g1010 ( 
.A(n_1003),
.B(n_844),
.C(n_903),
.Y(n_1010)
);

OAI211xp5_ASAP7_75t_L g1011 ( 
.A1(n_1006),
.A2(n_916),
.B(n_913),
.C(n_902),
.Y(n_1011)
);

NAND4xp75_ASAP7_75t_L g1012 ( 
.A(n_1009),
.B(n_892),
.C(n_890),
.D(n_902),
.Y(n_1012)
);

NOR4xp25_ASAP7_75t_L g1013 ( 
.A(n_1005),
.B(n_909),
.C(n_902),
.D(n_903),
.Y(n_1013)
);

AOI322xp5_ASAP7_75t_L g1014 ( 
.A1(n_1010),
.A2(n_903),
.A3(n_850),
.B1(n_881),
.B2(n_917),
.C1(n_892),
.C2(n_859),
.Y(n_1014)
);

OAI211xp5_ASAP7_75t_L g1015 ( 
.A1(n_1008),
.A2(n_914),
.B(n_846),
.C(n_892),
.Y(n_1015)
);

NOR3xp33_ASAP7_75t_L g1016 ( 
.A(n_1007),
.B(n_845),
.C(n_859),
.Y(n_1016)
);

AOI21xp33_ASAP7_75t_SL g1017 ( 
.A1(n_1009),
.A2(n_890),
.B(n_870),
.Y(n_1017)
);

NAND2xp5_ASAP7_75t_L g1018 ( 
.A(n_1013),
.B(n_870),
.Y(n_1018)
);

NAND3xp33_ASAP7_75t_L g1019 ( 
.A(n_1016),
.B(n_890),
.C(n_888),
.Y(n_1019)
);

AOI211xp5_ASAP7_75t_L g1020 ( 
.A1(n_1015),
.A2(n_846),
.B(n_891),
.C(n_888),
.Y(n_1020)
);

INVx1_ASAP7_75t_SL g1021 ( 
.A(n_1012),
.Y(n_1021)
);

NOR2xp33_ASAP7_75t_L g1022 ( 
.A(n_1011),
.B(n_890),
.Y(n_1022)
);

NAND4xp75_ASAP7_75t_L g1023 ( 
.A(n_1014),
.B(n_917),
.C(n_881),
.D(n_889),
.Y(n_1023)
);

NOR3xp33_ASAP7_75t_L g1024 ( 
.A(n_1017),
.B(n_845),
.C(n_849),
.Y(n_1024)
);

OAI21xp33_ASAP7_75t_SL g1025 ( 
.A1(n_1013),
.A2(n_914),
.B(n_917),
.Y(n_1025)
);

INVx2_ASAP7_75t_L g1026 ( 
.A(n_1012),
.Y(n_1026)
);

NAND2xp5_ASAP7_75t_SL g1027 ( 
.A(n_1026),
.B(n_914),
.Y(n_1027)
);

BUFx2_ASAP7_75t_L g1028 ( 
.A(n_1021),
.Y(n_1028)
);

OAI211xp5_ASAP7_75t_L g1029 ( 
.A1(n_1020),
.A2(n_891),
.B(n_850),
.C(n_921),
.Y(n_1029)
);

OR2x2_ASAP7_75t_L g1030 ( 
.A(n_1018),
.B(n_921),
.Y(n_1030)
);

NOR2x1_ASAP7_75t_L g1031 ( 
.A(n_1023),
.B(n_1022),
.Y(n_1031)
);

NAND2xp5_ASAP7_75t_L g1032 ( 
.A(n_1024),
.B(n_921),
.Y(n_1032)
);

INVx1_ASAP7_75t_L g1033 ( 
.A(n_1019),
.Y(n_1033)
);

OAI22xp33_ASAP7_75t_L g1034 ( 
.A1(n_1025),
.A2(n_850),
.B1(n_842),
.B2(n_867),
.Y(n_1034)
);

OAI22xp5_ASAP7_75t_SL g1035 ( 
.A1(n_1021),
.A2(n_850),
.B1(n_842),
.B2(n_867),
.Y(n_1035)
);

OAI221xp5_ASAP7_75t_L g1036 ( 
.A1(n_1021),
.A2(n_842),
.B1(n_868),
.B2(n_884),
.C(n_885),
.Y(n_1036)
);

NOR2x1_ASAP7_75t_L g1037 ( 
.A(n_1026),
.B(n_837),
.Y(n_1037)
);

NAND4xp25_ASAP7_75t_L g1038 ( 
.A(n_1028),
.B(n_1031),
.C(n_1033),
.D(n_1027),
.Y(n_1038)
);

NOR4xp25_ASAP7_75t_L g1039 ( 
.A(n_1030),
.B(n_884),
.C(n_853),
.D(n_885),
.Y(n_1039)
);

NAND4xp75_ASAP7_75t_L g1040 ( 
.A(n_1037),
.B(n_853),
.C(n_858),
.D(n_848),
.Y(n_1040)
);

NOR4xp75_ASAP7_75t_L g1041 ( 
.A(n_1036),
.B(n_95),
.C(n_98),
.D(n_99),
.Y(n_1041)
);

OAI21xp5_ASAP7_75t_L g1042 ( 
.A1(n_1034),
.A2(n_1029),
.B(n_1032),
.Y(n_1042)
);

AND2x4_ASAP7_75t_L g1043 ( 
.A(n_1035),
.B(n_848),
.Y(n_1043)
);

INVx2_ASAP7_75t_L g1044 ( 
.A(n_1028),
.Y(n_1044)
);

INVx1_ASAP7_75t_L g1045 ( 
.A(n_1028),
.Y(n_1045)
);

NOR3xp33_ASAP7_75t_SL g1046 ( 
.A(n_1033),
.B(n_103),
.C(n_105),
.Y(n_1046)
);

AND3x1_ASAP7_75t_L g1047 ( 
.A(n_1031),
.B(n_858),
.C(n_110),
.Y(n_1047)
);

NAND4xp75_ASAP7_75t_L g1048 ( 
.A(n_1031),
.B(n_106),
.C(n_111),
.D(n_112),
.Y(n_1048)
);

AND3x1_ASAP7_75t_L g1049 ( 
.A(n_1031),
.B(n_120),
.C(n_121),
.Y(n_1049)
);

AND2x2_ASAP7_75t_L g1050 ( 
.A(n_1028),
.B(n_837),
.Y(n_1050)
);

NAND4xp75_ASAP7_75t_L g1051 ( 
.A(n_1045),
.B(n_122),
.C(n_124),
.D(n_125),
.Y(n_1051)
);

NOR2xp67_ASAP7_75t_R g1052 ( 
.A(n_1044),
.B(n_126),
.Y(n_1052)
);

OAI22xp5_ASAP7_75t_SL g1053 ( 
.A1(n_1047),
.A2(n_1049),
.B1(n_1038),
.B2(n_1042),
.Y(n_1053)
);

INVx2_ASAP7_75t_L g1054 ( 
.A(n_1048),
.Y(n_1054)
);

INVx2_ASAP7_75t_L g1055 ( 
.A(n_1040),
.Y(n_1055)
);

NOR2xp67_ASAP7_75t_L g1056 ( 
.A(n_1050),
.B(n_129),
.Y(n_1056)
);

INVx2_ASAP7_75t_L g1057 ( 
.A(n_1043),
.Y(n_1057)
);

INVx1_ASAP7_75t_L g1058 ( 
.A(n_1046),
.Y(n_1058)
);

AOI222xp33_ASAP7_75t_L g1059 ( 
.A1(n_1041),
.A2(n_849),
.B1(n_893),
.B2(n_895),
.C1(n_831),
.C2(n_839),
.Y(n_1059)
);

OAI22x1_ASAP7_75t_L g1060 ( 
.A1(n_1058),
.A2(n_1039),
.B1(n_895),
.B2(n_893),
.Y(n_1060)
);

INVx1_ASAP7_75t_L g1061 ( 
.A(n_1053),
.Y(n_1061)
);

INVx1_ASAP7_75t_L g1062 ( 
.A(n_1052),
.Y(n_1062)
);

AO22x1_ASAP7_75t_L g1063 ( 
.A1(n_1054),
.A2(n_130),
.B1(n_131),
.B2(n_132),
.Y(n_1063)
);

OAI22xp5_ASAP7_75t_L g1064 ( 
.A1(n_1055),
.A2(n_831),
.B1(n_839),
.B2(n_840),
.Y(n_1064)
);

AOI22xp5_ASAP7_75t_L g1065 ( 
.A1(n_1056),
.A2(n_837),
.B1(n_840),
.B2(n_839),
.Y(n_1065)
);

OAI22xp5_ASAP7_75t_L g1066 ( 
.A1(n_1057),
.A2(n_840),
.B1(n_134),
.B2(n_135),
.Y(n_1066)
);

HB1xp67_ASAP7_75t_L g1067 ( 
.A(n_1051),
.Y(n_1067)
);

AOI22x1_ASAP7_75t_L g1068 ( 
.A1(n_1061),
.A2(n_1059),
.B1(n_136),
.B2(n_137),
.Y(n_1068)
);

NOR2xp67_ASAP7_75t_L g1069 ( 
.A(n_1062),
.B(n_133),
.Y(n_1069)
);

OAI22xp5_ASAP7_75t_L g1070 ( 
.A1(n_1067),
.A2(n_138),
.B1(n_139),
.B2(n_140),
.Y(n_1070)
);

INVx2_ASAP7_75t_L g1071 ( 
.A(n_1060),
.Y(n_1071)
);

AOI22xp5_ASAP7_75t_SL g1072 ( 
.A1(n_1071),
.A2(n_1063),
.B1(n_1066),
.B2(n_1064),
.Y(n_1072)
);

INVx1_ASAP7_75t_SL g1073 ( 
.A(n_1072),
.Y(n_1073)
);

AND2x2_ASAP7_75t_L g1074 ( 
.A(n_1073),
.B(n_1069),
.Y(n_1074)
);

AOI22xp5_ASAP7_75t_SL g1075 ( 
.A1(n_1074),
.A2(n_1070),
.B1(n_1068),
.B2(n_1065),
.Y(n_1075)
);

NAND2xp5_ASAP7_75t_L g1076 ( 
.A(n_1075),
.B(n_144),
.Y(n_1076)
);

AOI22xp33_ASAP7_75t_L g1077 ( 
.A1(n_1076),
.A2(n_145),
.B1(n_147),
.B2(n_148),
.Y(n_1077)
);

OAI22xp5_ASAP7_75t_L g1078 ( 
.A1(n_1077),
.A2(n_149),
.B1(n_150),
.B2(n_152),
.Y(n_1078)
);

AOI211xp5_ASAP7_75t_L g1079 ( 
.A1(n_1078),
.A2(n_154),
.B(n_155),
.C(n_158),
.Y(n_1079)
);


endmodule