module fake_jpeg_31480_n_467 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_467);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_467;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_145;
wire n_20;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

INVx4_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

BUFx10_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_11),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

INVx8_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_7),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

BUFx12_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

CKINVDCx16_ASAP7_75t_R g33 ( 
.A(n_14),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_3),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_13),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_0),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_5),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_15),
.Y(n_38)
);

BUFx4f_ASAP7_75t_L g39 ( 
.A(n_8),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_6),
.Y(n_40)
);

BUFx8_ASAP7_75t_L g41 ( 
.A(n_5),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_9),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_4),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_0),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_15),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_5),
.Y(n_46)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_13),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_14),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_27),
.Y(n_49)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_49),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_35),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_50),
.B(n_51),
.Y(n_111)
);

OR2x2_ASAP7_75t_L g51 ( 
.A(n_38),
.B(n_29),
.Y(n_51)
);

INVx11_ASAP7_75t_L g52 ( 
.A(n_26),
.Y(n_52)
);

INVx5_ASAP7_75t_L g106 ( 
.A(n_52),
.Y(n_106)
);

INVx6_ASAP7_75t_SL g53 ( 
.A(n_48),
.Y(n_53)
);

CKINVDCx16_ASAP7_75t_R g107 ( 
.A(n_53),
.Y(n_107)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_27),
.Y(n_54)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_54),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_35),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_55),
.B(n_60),
.Y(n_129)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_41),
.Y(n_56)
);

INVx8_ASAP7_75t_L g136 ( 
.A(n_56),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_16),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_57),
.Y(n_98)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_16),
.Y(n_58)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_58),
.Y(n_97)
);

INVx2_ASAP7_75t_SL g59 ( 
.A(n_39),
.Y(n_59)
);

INVx2_ASAP7_75t_SL g121 ( 
.A(n_59),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_19),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_16),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_61),
.Y(n_123)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_22),
.Y(n_62)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_62),
.Y(n_100)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_41),
.Y(n_63)
);

INVx5_ASAP7_75t_L g115 ( 
.A(n_63),
.Y(n_115)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_26),
.Y(n_64)
);

INVx5_ASAP7_75t_L g131 ( 
.A(n_64),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_16),
.Y(n_65)
);

INVx6_ASAP7_75t_L g110 ( 
.A(n_65),
.Y(n_110)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_26),
.Y(n_66)
);

BUFx3_ASAP7_75t_L g139 ( 
.A(n_66),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_19),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_67),
.B(n_72),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_28),
.Y(n_68)
);

INVx6_ASAP7_75t_L g128 ( 
.A(n_68),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_28),
.Y(n_69)
);

INVx6_ASAP7_75t_L g145 ( 
.A(n_69),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_28),
.Y(n_70)
);

INVx4_ASAP7_75t_L g105 ( 
.A(n_70),
.Y(n_105)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_45),
.Y(n_71)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_71),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_19),
.Y(n_72)
);

CKINVDCx9p33_ASAP7_75t_R g73 ( 
.A(n_39),
.Y(n_73)
);

INVx4_ASAP7_75t_L g140 ( 
.A(n_73),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_22),
.B(n_1),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_74),
.B(n_83),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_28),
.Y(n_75)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_75),
.Y(n_104)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_47),
.Y(n_76)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_76),
.Y(n_99)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_47),
.Y(n_77)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_77),
.Y(n_101)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_45),
.Y(n_78)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_78),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_38),
.B(n_15),
.Y(n_79)
);

AND2x2_ASAP7_75t_L g137 ( 
.A(n_79),
.B(n_80),
.Y(n_137)
);

INVx1_ASAP7_75t_SL g80 ( 
.A(n_18),
.Y(n_80)
);

BUFx12_ASAP7_75t_L g81 ( 
.A(n_39),
.Y(n_81)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_81),
.Y(n_120)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_18),
.Y(n_82)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_82),
.Y(n_118)
);

INVx1_ASAP7_75t_SL g83 ( 
.A(n_18),
.Y(n_83)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_17),
.Y(n_84)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_84),
.Y(n_127)
);

BUFx3_ASAP7_75t_L g85 ( 
.A(n_30),
.Y(n_85)
);

INVx3_ASAP7_75t_L g143 ( 
.A(n_85),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_35),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_86),
.B(n_89),
.Y(n_124)
);

INVx8_ASAP7_75t_L g87 ( 
.A(n_41),
.Y(n_87)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_87),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_48),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_88),
.A2(n_43),
.B1(n_42),
.B2(n_37),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_33),
.B(n_14),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_SL g90 ( 
.A(n_33),
.B(n_12),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_90),
.B(n_93),
.Y(n_141)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_30),
.Y(n_91)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_91),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_30),
.Y(n_92)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_92),
.Y(n_146)
);

INVx5_ASAP7_75t_L g93 ( 
.A(n_47),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_19),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_94),
.B(n_95),
.Y(n_149)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_17),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_53),
.A2(n_36),
.B1(n_30),
.B2(n_32),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g171 ( 
.A1(n_96),
.A2(n_125),
.B1(n_126),
.B2(n_133),
.Y(n_171)
);

AOI22xp33_ASAP7_75t_L g103 ( 
.A1(n_62),
.A2(n_48),
.B1(n_40),
.B2(n_29),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_103),
.A2(n_112),
.B1(n_122),
.B2(n_132),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_49),
.A2(n_48),
.B1(n_40),
.B2(n_24),
.Y(n_112)
);

OAI22xp33_ASAP7_75t_L g113 ( 
.A1(n_57),
.A2(n_34),
.B1(n_32),
.B2(n_39),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_113),
.A2(n_116),
.B1(n_147),
.B2(n_59),
.Y(n_197)
);

OAI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_74),
.A2(n_34),
.B1(n_32),
.B2(n_39),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_54),
.A2(n_24),
.B1(n_46),
.B2(n_23),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_56),
.A2(n_87),
.B1(n_63),
.B2(n_85),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_73),
.A2(n_36),
.B1(n_34),
.B2(n_32),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_L g132 ( 
.A1(n_61),
.A2(n_34),
.B1(n_46),
.B2(n_23),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_64),
.A2(n_36),
.B1(n_44),
.B2(n_21),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_66),
.A2(n_36),
.B1(n_44),
.B2(n_21),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_SL g194 ( 
.A1(n_134),
.A2(n_59),
.B1(n_58),
.B2(n_93),
.Y(n_194)
);

AND2x2_ASAP7_75t_SL g135 ( 
.A(n_82),
.B(n_2),
.Y(n_135)
);

AND2x2_ASAP7_75t_L g198 ( 
.A(n_135),
.B(n_148),
.Y(n_198)
);

AOI22xp33_ASAP7_75t_L g138 ( 
.A1(n_65),
.A2(n_43),
.B1(n_42),
.B2(n_37),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_L g186 ( 
.A1(n_138),
.A2(n_69),
.B1(n_92),
.B2(n_68),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_51),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_SL g178 ( 
.A(n_144),
.B(n_25),
.Y(n_178)
);

AND2x4_ASAP7_75t_L g148 ( 
.A(n_88),
.B(n_41),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_109),
.B(n_95),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_150),
.B(n_154),
.Y(n_204)
);

BUFx6f_ASAP7_75t_L g152 ( 
.A(n_98),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g214 ( 
.A(n_152),
.Y(n_214)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_102),
.Y(n_153)
);

CKINVDCx16_ASAP7_75t_R g205 ( 
.A(n_153),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_135),
.B(n_84),
.Y(n_154)
);

CKINVDCx16_ASAP7_75t_R g155 ( 
.A(n_142),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_155),
.B(n_162),
.Y(n_224)
);

BUFx12f_ASAP7_75t_L g156 ( 
.A(n_115),
.Y(n_156)
);

INVx3_ASAP7_75t_L g227 ( 
.A(n_156),
.Y(n_227)
);

INVx6_ASAP7_75t_L g157 ( 
.A(n_98),
.Y(n_157)
);

INVx5_ASAP7_75t_L g241 ( 
.A(n_157),
.Y(n_241)
);

BUFx3_ASAP7_75t_L g158 ( 
.A(n_139),
.Y(n_158)
);

CKINVDCx14_ASAP7_75t_R g206 ( 
.A(n_158),
.Y(n_206)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_108),
.Y(n_159)
);

CKINVDCx16_ASAP7_75t_R g233 ( 
.A(n_159),
.Y(n_233)
);

INVx5_ASAP7_75t_L g160 ( 
.A(n_115),
.Y(n_160)
);

INVx1_ASAP7_75t_SL g232 ( 
.A(n_160),
.Y(n_232)
);

AOI21xp5_ASAP7_75t_L g161 ( 
.A1(n_148),
.A2(n_83),
.B(n_80),
.Y(n_161)
);

AOI21xp5_ASAP7_75t_L g228 ( 
.A1(n_161),
.A2(n_163),
.B(n_131),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_107),
.Y(n_162)
);

O2A1O1Ixp33_ASAP7_75t_L g163 ( 
.A1(n_148),
.A2(n_60),
.B(n_72),
.C(n_67),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_149),
.B(n_124),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_164),
.B(n_168),
.Y(n_218)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_114),
.Y(n_165)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_165),
.Y(n_212)
);

HB1xp67_ASAP7_75t_L g166 ( 
.A(n_99),
.Y(n_166)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_166),
.Y(n_202)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_130),
.Y(n_167)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_167),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_111),
.B(n_71),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_129),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_169),
.B(n_177),
.Y(n_231)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_100),
.Y(n_170)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_170),
.Y(n_215)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_127),
.Y(n_172)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_172),
.Y(n_229)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_117),
.Y(n_173)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_173),
.Y(n_235)
);

INVx6_ASAP7_75t_L g174 ( 
.A(n_123),
.Y(n_174)
);

INVx2_ASAP7_75t_SL g238 ( 
.A(n_174),
.Y(n_238)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_118),
.Y(n_175)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_175),
.Y(n_239)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_146),
.Y(n_176)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_176),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_141),
.B(n_78),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_178),
.Y(n_201)
);

BUFx6f_ASAP7_75t_L g179 ( 
.A(n_123),
.Y(n_179)
);

INVxp67_ASAP7_75t_L g210 ( 
.A(n_179),
.Y(n_210)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_99),
.Y(n_180)
);

INVxp67_ASAP7_75t_L g222 ( 
.A(n_180),
.Y(n_222)
);

OR2x2_ASAP7_75t_L g181 ( 
.A(n_137),
.B(n_31),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_181),
.Y(n_217)
);

XNOR2x1_ASAP7_75t_L g182 ( 
.A(n_135),
.B(n_41),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_182),
.B(n_199),
.C(n_121),
.Y(n_216)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_104),
.Y(n_183)
);

NAND2xp33_ASAP7_75t_SL g209 ( 
.A(n_183),
.B(n_188),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_148),
.B(n_91),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_184),
.B(n_187),
.Y(n_236)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_101),
.Y(n_185)
);

AND2x2_ASAP7_75t_L g207 ( 
.A(n_185),
.B(n_193),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_186),
.A2(n_126),
.B1(n_134),
.B2(n_133),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_137),
.B(n_121),
.Y(n_187)
);

INVx4_ASAP7_75t_SL g188 ( 
.A(n_140),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_101),
.Y(n_189)
);

INVxp67_ASAP7_75t_L g225 ( 
.A(n_189),
.Y(n_225)
);

CKINVDCx14_ASAP7_75t_R g190 ( 
.A(n_119),
.Y(n_190)
);

INVxp67_ASAP7_75t_L g234 ( 
.A(n_190),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_139),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_191),
.Y(n_203)
);

INVx4_ASAP7_75t_L g192 ( 
.A(n_97),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_192),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_120),
.B(n_31),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g208 ( 
.A1(n_194),
.A2(n_125),
.B1(n_96),
.B2(n_140),
.Y(n_208)
);

INVx2_ASAP7_75t_SL g195 ( 
.A(n_97),
.Y(n_195)
);

AND2x2_ASAP7_75t_L g220 ( 
.A(n_195),
.B(n_196),
.Y(n_220)
);

INVx3_ASAP7_75t_L g196 ( 
.A(n_120),
.Y(n_196)
);

AND2x2_ASAP7_75t_L g223 ( 
.A(n_197),
.B(n_105),
.Y(n_223)
);

AND2x2_ASAP7_75t_SL g199 ( 
.A(n_131),
.B(n_76),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_200),
.A2(n_211),
.B1(n_219),
.B2(n_221),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_208),
.A2(n_162),
.B1(n_143),
.B2(n_136),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_L g211 ( 
.A1(n_197),
.A2(n_145),
.B1(n_110),
.B2(n_128),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_151),
.A2(n_113),
.B1(n_110),
.B2(n_145),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_213),
.A2(n_236),
.B1(n_200),
.B2(n_234),
.Y(n_275)
);

AND2x2_ASAP7_75t_L g255 ( 
.A(n_216),
.B(n_226),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_184),
.A2(n_171),
.B1(n_150),
.B2(n_154),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_163),
.A2(n_70),
.B1(n_75),
.B2(n_128),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_223),
.A2(n_199),
.B1(n_161),
.B2(n_151),
.Y(n_245)
);

AND2x2_ASAP7_75t_L g226 ( 
.A(n_198),
.B(n_77),
.Y(n_226)
);

OAI21xp5_ASAP7_75t_SL g267 ( 
.A1(n_228),
.A2(n_185),
.B(n_195),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_198),
.B(n_105),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_240),
.B(n_182),
.Y(n_249)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_229),
.Y(n_243)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_243),
.Y(n_284)
);

INVx1_ASAP7_75t_SL g299 ( 
.A(n_245),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_224),
.B(n_201),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_SL g302 ( 
.A(n_246),
.B(n_247),
.Y(n_302)
);

CKINVDCx14_ASAP7_75t_R g247 ( 
.A(n_207),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_L g248 ( 
.A1(n_213),
.A2(n_187),
.B1(n_198),
.B2(n_181),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_248),
.A2(n_251),
.B1(n_275),
.B2(n_217),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_249),
.B(n_265),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_220),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_250),
.B(n_252),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_L g251 ( 
.A1(n_223),
.A2(n_172),
.B1(n_199),
.B2(n_157),
.Y(n_251)
);

INVxp67_ASAP7_75t_L g252 ( 
.A(n_220),
.Y(n_252)
);

INVx4_ASAP7_75t_L g253 ( 
.A(n_227),
.Y(n_253)
);

BUFx2_ASAP7_75t_L g286 ( 
.A(n_253),
.Y(n_286)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_229),
.Y(n_254)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_254),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_L g293 ( 
.A1(n_256),
.A2(n_272),
.B1(n_232),
.B2(n_206),
.Y(n_293)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_212),
.Y(n_257)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_257),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_220),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_258),
.B(n_261),
.Y(n_312)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_242),
.Y(n_259)
);

CKINVDCx16_ASAP7_75t_R g287 ( 
.A(n_259),
.Y(n_287)
);

INVx5_ASAP7_75t_L g260 ( 
.A(n_241),
.Y(n_260)
);

HB1xp67_ASAP7_75t_L g288 ( 
.A(n_260),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_201),
.B(n_196),
.Y(n_261)
);

AND2x2_ASAP7_75t_L g262 ( 
.A(n_226),
.B(n_170),
.Y(n_262)
);

INVxp67_ASAP7_75t_L g304 ( 
.A(n_262),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_205),
.B(n_192),
.Y(n_263)
);

CKINVDCx16_ASAP7_75t_R g313 ( 
.A(n_263),
.Y(n_313)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_237),
.Y(n_264)
);

BUFx4f_ASAP7_75t_L g307 ( 
.A(n_264),
.Y(n_307)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_212),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_235),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_266),
.B(n_270),
.Y(n_303)
);

OAI21xp5_ASAP7_75t_SL g305 ( 
.A1(n_267),
.A2(n_268),
.B(n_277),
.Y(n_305)
);

AOI32xp33_ASAP7_75t_L g268 ( 
.A1(n_217),
.A2(n_143),
.A3(n_174),
.B1(n_160),
.B2(n_156),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_204),
.B(n_236),
.C(n_216),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_L g290 ( 
.A(n_269),
.B(n_271),
.Y(n_290)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_235),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_204),
.B(n_175),
.Y(n_271)
);

AOI22xp33_ASAP7_75t_L g272 ( 
.A1(n_223),
.A2(n_152),
.B1(n_179),
.B2(n_188),
.Y(n_272)
);

INVx1_ASAP7_75t_SL g273 ( 
.A(n_207),
.Y(n_273)
);

OR2x2_ASAP7_75t_L g292 ( 
.A(n_273),
.B(n_209),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_219),
.A2(n_167),
.B1(n_183),
.B2(n_106),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_SL g298 ( 
.A1(n_274),
.A2(n_278),
.B1(n_238),
.B2(n_232),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_240),
.B(n_20),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_276),
.B(n_279),
.Y(n_297)
);

AND2x2_ASAP7_75t_L g277 ( 
.A(n_226),
.B(n_158),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_228),
.A2(n_106),
.B1(n_136),
.B2(n_52),
.Y(n_278)
);

AND2x2_ASAP7_75t_L g279 ( 
.A(n_221),
.B(n_20),
.Y(n_279)
);

INVxp67_ASAP7_75t_L g280 ( 
.A(n_207),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g300 ( 
.A(n_280),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_203),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_281),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_L g324 ( 
.A1(n_283),
.A2(n_279),
.B1(n_256),
.B2(n_278),
.Y(n_324)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_275),
.A2(n_234),
.B1(n_231),
.B2(n_233),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_SL g319 ( 
.A1(n_289),
.A2(n_315),
.B1(n_274),
.B2(n_280),
.Y(n_319)
);

OR2x2_ASAP7_75t_L g317 ( 
.A(n_292),
.B(n_301),
.Y(n_317)
);

AOI22xp5_ASAP7_75t_L g320 ( 
.A1(n_293),
.A2(n_298),
.B1(n_311),
.B2(n_252),
.Y(n_320)
);

OAI21xp5_ASAP7_75t_L g294 ( 
.A1(n_273),
.A2(n_242),
.B(n_225),
.Y(n_294)
);

AND2x2_ASAP7_75t_L g333 ( 
.A(n_294),
.B(n_296),
.Y(n_333)
);

XOR2xp5_ASAP7_75t_L g295 ( 
.A(n_269),
.B(n_218),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_295),
.B(n_310),
.C(n_255),
.Y(n_322)
);

OAI21xp5_ASAP7_75t_L g296 ( 
.A1(n_249),
.A2(n_225),
.B(n_222),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g301 ( 
.A(n_264),
.Y(n_301)
);

OAI21xp5_ASAP7_75t_L g308 ( 
.A1(n_245),
.A2(n_222),
.B(n_230),
.Y(n_308)
);

XNOR2xp5_ASAP7_75t_SL g336 ( 
.A(n_308),
.B(n_314),
.Y(n_336)
);

XOR2xp5_ASAP7_75t_L g310 ( 
.A(n_255),
.B(n_215),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_L g311 ( 
.A1(n_244),
.A2(n_238),
.B1(n_210),
.B2(n_241),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_L g314 ( 
.A(n_255),
.B(n_239),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_L g315 ( 
.A1(n_244),
.A2(n_238),
.B1(n_210),
.B2(n_239),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_257),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_SL g339 ( 
.A(n_316),
.B(n_215),
.Y(n_339)
);

CKINVDCx14_ASAP7_75t_R g318 ( 
.A(n_302),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_318),
.B(n_338),
.Y(n_349)
);

AOI22xp5_ASAP7_75t_L g347 ( 
.A1(n_319),
.A2(n_324),
.B1(n_334),
.B2(n_345),
.Y(n_347)
);

OAI22xp5_ASAP7_75t_L g372 ( 
.A1(n_320),
.A2(n_343),
.B1(n_286),
.B2(n_25),
.Y(n_372)
);

AOI21xp33_ASAP7_75t_L g321 ( 
.A1(n_313),
.A2(n_276),
.B(n_267),
.Y(n_321)
);

OAI21xp33_ASAP7_75t_L g373 ( 
.A1(n_321),
.A2(n_326),
.B(n_156),
.Y(n_373)
);

XOR2xp5_ASAP7_75t_L g354 ( 
.A(n_322),
.B(n_297),
.Y(n_354)
);

XOR2xp5_ASAP7_75t_L g323 ( 
.A(n_290),
.B(n_271),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g350 ( 
.A(n_323),
.B(n_327),
.C(n_331),
.Y(n_350)
);

OAI22xp5_ASAP7_75t_L g325 ( 
.A1(n_289),
.A2(n_279),
.B1(n_254),
.B2(n_243),
.Y(n_325)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_325),
.Y(n_368)
);

NOR2xp33_ASAP7_75t_SL g326 ( 
.A(n_291),
.B(n_295),
.Y(n_326)
);

XOR2xp5_ASAP7_75t_L g327 ( 
.A(n_290),
.B(n_277),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_303),
.Y(n_328)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_328),
.Y(n_352)
);

INVx2_ASAP7_75t_L g329 ( 
.A(n_307),
.Y(n_329)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_329),
.Y(n_364)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_303),
.Y(n_330)
);

CKINVDCx16_ASAP7_75t_R g362 ( 
.A(n_330),
.Y(n_362)
);

XOR2xp5_ASAP7_75t_L g331 ( 
.A(n_310),
.B(n_277),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g332 ( 
.A(n_307),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g358 ( 
.A(n_332),
.Y(n_358)
);

OAI22xp5_ASAP7_75t_SL g334 ( 
.A1(n_299),
.A2(n_270),
.B1(n_266),
.B2(n_265),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_314),
.B(n_262),
.C(n_202),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g356 ( 
.A(n_335),
.B(n_342),
.C(n_346),
.Y(n_356)
);

NOR2xp33_ASAP7_75t_L g337 ( 
.A(n_312),
.B(n_253),
.Y(n_337)
);

CKINVDCx20_ASAP7_75t_R g360 ( 
.A(n_337),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_282),
.B(n_262),
.Y(n_338)
);

CKINVDCx20_ASAP7_75t_R g361 ( 
.A(n_339),
.Y(n_361)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_306),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_340),
.B(n_344),
.Y(n_351)
);

CKINVDCx16_ASAP7_75t_R g341 ( 
.A(n_306),
.Y(n_341)
);

CKINVDCx20_ASAP7_75t_R g365 ( 
.A(n_341),
.Y(n_365)
);

XOR2xp5_ASAP7_75t_L g342 ( 
.A(n_282),
.B(n_202),
.Y(n_342)
);

OAI22xp5_ASAP7_75t_L g343 ( 
.A1(n_315),
.A2(n_283),
.B1(n_299),
.B2(n_308),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_284),
.Y(n_344)
);

OAI22xp5_ASAP7_75t_SL g345 ( 
.A1(n_305),
.A2(n_260),
.B1(n_214),
.B2(n_237),
.Y(n_345)
);

XOR2xp5_ASAP7_75t_L g346 ( 
.A(n_296),
.B(n_227),
.Y(n_346)
);

INVx3_ASAP7_75t_L g348 ( 
.A(n_329),
.Y(n_348)
);

BUFx2_ASAP7_75t_L g384 ( 
.A(n_348),
.Y(n_384)
);

OAI21xp5_ASAP7_75t_SL g353 ( 
.A1(n_317),
.A2(n_305),
.B(n_292),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_SL g374 ( 
.A(n_353),
.B(n_366),
.Y(n_374)
);

XOR2xp5_ASAP7_75t_L g388 ( 
.A(n_354),
.B(n_370),
.Y(n_388)
);

XNOR2xp5_ASAP7_75t_L g355 ( 
.A(n_323),
.B(n_297),
.Y(n_355)
);

XNOR2xp5_ASAP7_75t_L g392 ( 
.A(n_355),
.B(n_81),
.Y(n_392)
);

MAJIxp5_ASAP7_75t_L g357 ( 
.A(n_322),
.B(n_304),
.C(n_300),
.Y(n_357)
);

MAJIxp5_ASAP7_75t_L g379 ( 
.A(n_357),
.B(n_367),
.C(n_346),
.Y(n_379)
);

OAI22xp5_ASAP7_75t_SL g359 ( 
.A1(n_328),
.A2(n_304),
.B1(n_300),
.B2(n_294),
.Y(n_359)
);

AOI22xp5_ASAP7_75t_L g378 ( 
.A1(n_359),
.A2(n_363),
.B1(n_372),
.B2(n_333),
.Y(n_378)
);

OAI22xp5_ASAP7_75t_SL g363 ( 
.A1(n_330),
.A2(n_298),
.B1(n_309),
.B2(n_285),
.Y(n_363)
);

OAI21xp5_ASAP7_75t_SL g366 ( 
.A1(n_317),
.A2(n_288),
.B(n_285),
.Y(n_366)
);

MAJIxp5_ASAP7_75t_L g367 ( 
.A(n_327),
.B(n_284),
.C(n_287),
.Y(n_367)
);

FAx1_ASAP7_75t_SL g369 ( 
.A(n_336),
.B(n_333),
.CI(n_338),
.CON(n_369),
.SN(n_369)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_369),
.Y(n_387)
);

XOR2xp5_ASAP7_75t_L g370 ( 
.A(n_336),
.B(n_307),
.Y(n_370)
);

AOI22xp5_ASAP7_75t_L g371 ( 
.A1(n_319),
.A2(n_301),
.B1(n_286),
.B2(n_214),
.Y(n_371)
);

OAI22xp5_ASAP7_75t_SL g382 ( 
.A1(n_371),
.A2(n_332),
.B1(n_335),
.B2(n_334),
.Y(n_382)
);

NOR2xp67_ASAP7_75t_SL g381 ( 
.A(n_373),
.B(n_331),
.Y(n_381)
);

CKINVDCx20_ASAP7_75t_R g375 ( 
.A(n_351),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_375),
.B(n_383),
.Y(n_402)
);

OAI21xp5_ASAP7_75t_L g376 ( 
.A1(n_349),
.A2(n_333),
.B(n_320),
.Y(n_376)
);

OAI21xp5_ASAP7_75t_L g404 ( 
.A1(n_376),
.A2(n_347),
.B(n_371),
.Y(n_404)
);

OAI22xp33_ASAP7_75t_SL g377 ( 
.A1(n_352),
.A2(n_340),
.B1(n_344),
.B2(n_345),
.Y(n_377)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_377),
.Y(n_398)
);

NOR2xp33_ASAP7_75t_L g406 ( 
.A(n_378),
.B(n_394),
.Y(n_406)
);

XOR2xp5_ASAP7_75t_L g399 ( 
.A(n_379),
.B(n_392),
.Y(n_399)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_351),
.Y(n_380)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_380),
.Y(n_401)
);

BUFx12_ASAP7_75t_L g413 ( 
.A(n_381),
.Y(n_413)
);

AND2x2_ASAP7_75t_L g410 ( 
.A(n_382),
.B(n_359),
.Y(n_410)
);

OAI22xp5_ASAP7_75t_SL g383 ( 
.A1(n_347),
.A2(n_342),
.B1(n_58),
.B2(n_36),
.Y(n_383)
);

CKINVDCx20_ASAP7_75t_R g385 ( 
.A(n_349),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_385),
.B(n_393),
.Y(n_409)
);

OAI22xp5_ASAP7_75t_L g386 ( 
.A1(n_361),
.A2(n_12),
.B1(n_31),
.B2(n_4),
.Y(n_386)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_386),
.Y(n_405)
);

XNOR2xp5_ASAP7_75t_SL g389 ( 
.A(n_370),
.B(n_81),
.Y(n_389)
);

XNOR2xp5_ASAP7_75t_SL g403 ( 
.A(n_389),
.B(n_356),
.Y(n_403)
);

OAI22xp5_ASAP7_75t_L g390 ( 
.A1(n_368),
.A2(n_31),
.B1(n_3),
.B2(n_6),
.Y(n_390)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_390),
.Y(n_411)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_352),
.Y(n_391)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_391),
.Y(n_414)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_366),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_363),
.Y(n_394)
);

XOR2xp5_ASAP7_75t_L g395 ( 
.A(n_350),
.B(n_31),
.Y(n_395)
);

XOR2xp5_ASAP7_75t_L g407 ( 
.A(n_395),
.B(n_396),
.Y(n_407)
);

XOR2xp5_ASAP7_75t_L g396 ( 
.A(n_350),
.B(n_19),
.Y(n_396)
);

OAI21xp33_ASAP7_75t_L g397 ( 
.A1(n_374),
.A2(n_353),
.B(n_369),
.Y(n_397)
);

XOR2xp5_ASAP7_75t_L g417 ( 
.A(n_397),
.B(n_403),
.Y(n_417)
);

MAJIxp5_ASAP7_75t_L g400 ( 
.A(n_379),
.B(n_356),
.C(n_354),
.Y(n_400)
);

MAJIxp5_ASAP7_75t_L g415 ( 
.A(n_400),
.B(n_388),
.C(n_396),
.Y(n_415)
);

XOR2xp5_ASAP7_75t_L g428 ( 
.A(n_404),
.B(n_383),
.Y(n_428)
);

NOR2xp33_ASAP7_75t_L g408 ( 
.A(n_378),
.B(n_365),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_408),
.B(n_410),
.Y(n_416)
);

XOR2xp5_ASAP7_75t_L g412 ( 
.A(n_388),
.B(n_355),
.Y(n_412)
);

XOR2xp5_ASAP7_75t_L g425 ( 
.A(n_412),
.B(n_389),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_L g436 ( 
.A(n_415),
.B(n_418),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g418 ( 
.A(n_414),
.B(n_360),
.Y(n_418)
);

XNOR2xp5_ASAP7_75t_L g419 ( 
.A(n_400),
.B(n_399),
.Y(n_419)
);

XOR2xp5_ASAP7_75t_L g433 ( 
.A(n_419),
.B(n_420),
.Y(n_433)
);

XNOR2xp5_ASAP7_75t_L g420 ( 
.A(n_399),
.B(n_367),
.Y(n_420)
);

NOR2xp33_ASAP7_75t_L g421 ( 
.A(n_402),
.B(n_393),
.Y(n_421)
);

CKINVDCx20_ASAP7_75t_R g439 ( 
.A(n_421),
.Y(n_439)
);

NOR2xp33_ASAP7_75t_L g422 ( 
.A(n_406),
.B(n_382),
.Y(n_422)
);

NOR2xp33_ASAP7_75t_SL g440 ( 
.A(n_422),
.B(n_423),
.Y(n_440)
);

NOR2xp33_ASAP7_75t_L g423 ( 
.A(n_409),
.B(n_362),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_SL g424 ( 
.A(n_410),
.B(n_376),
.Y(n_424)
);

AOI21xp5_ASAP7_75t_L g431 ( 
.A1(n_424),
.A2(n_425),
.B(n_426),
.Y(n_431)
);

XOR2xp5_ASAP7_75t_L g426 ( 
.A(n_412),
.B(n_357),
.Y(n_426)
);

OAI22xp5_ASAP7_75t_L g427 ( 
.A1(n_405),
.A2(n_380),
.B1(n_391),
.B2(n_358),
.Y(n_427)
);

HB1xp67_ASAP7_75t_L g435 ( 
.A(n_427),
.Y(n_435)
);

AOI21xp5_ASAP7_75t_L g432 ( 
.A1(n_428),
.A2(n_410),
.B(n_387),
.Y(n_432)
);

OAI22xp5_ASAP7_75t_L g429 ( 
.A1(n_416),
.A2(n_398),
.B1(n_404),
.B2(n_411),
.Y(n_429)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_429),
.Y(n_445)
);

AND2x2_ASAP7_75t_L g430 ( 
.A(n_428),
.B(n_401),
.Y(n_430)
);

OR2x2_ASAP7_75t_L g441 ( 
.A(n_430),
.B(n_369),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_SL g444 ( 
.A(n_432),
.B(n_440),
.Y(n_444)
);

OAI22xp5_ASAP7_75t_SL g434 ( 
.A1(n_415),
.A2(n_397),
.B1(n_413),
.B2(n_364),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_434),
.B(n_438),
.Y(n_449)
);

AOI21xp5_ASAP7_75t_L g437 ( 
.A1(n_417),
.A2(n_413),
.B(n_395),
.Y(n_437)
);

OAI21xp5_ASAP7_75t_SL g446 ( 
.A1(n_437),
.A2(n_431),
.B(n_436),
.Y(n_446)
);

OAI21xp5_ASAP7_75t_L g438 ( 
.A1(n_417),
.A2(n_413),
.B(n_403),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_441),
.B(n_443),
.Y(n_452)
);

MAJIxp5_ASAP7_75t_L g442 ( 
.A(n_433),
.B(n_426),
.C(n_407),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_SL g455 ( 
.A(n_442),
.B(n_448),
.Y(n_455)
);

NOR2xp33_ASAP7_75t_L g443 ( 
.A(n_439),
.B(n_384),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_444),
.B(n_447),
.Y(n_456)
);

XNOR2xp5_ASAP7_75t_L g454 ( 
.A(n_446),
.B(n_443),
.Y(n_454)
);

NOR2xp33_ASAP7_75t_SL g447 ( 
.A(n_430),
.B(n_425),
.Y(n_447)
);

MAJIxp5_ASAP7_75t_L g448 ( 
.A(n_435),
.B(n_407),
.C(n_392),
.Y(n_448)
);

BUFx6f_ASAP7_75t_L g450 ( 
.A(n_435),
.Y(n_450)
);

NOR2xp33_ASAP7_75t_SL g451 ( 
.A(n_450),
.B(n_364),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_451),
.B(n_453),
.Y(n_459)
);

OAI21xp5_ASAP7_75t_L g453 ( 
.A1(n_449),
.A2(n_348),
.B(n_384),
.Y(n_453)
);

AND2x2_ASAP7_75t_L g461 ( 
.A(n_454),
.B(n_19),
.Y(n_461)
);

NOR2xp33_ASAP7_75t_L g457 ( 
.A(n_450),
.B(n_2),
.Y(n_457)
);

OAI21xp5_ASAP7_75t_L g458 ( 
.A1(n_457),
.A2(n_441),
.B(n_445),
.Y(n_458)
);

A2O1A1O1Ixp25_ASAP7_75t_L g463 ( 
.A1(n_458),
.A2(n_452),
.B(n_459),
.C(n_455),
.D(n_10),
.Y(n_463)
);

NOR2xp67_ASAP7_75t_SL g460 ( 
.A(n_456),
.B(n_6),
.Y(n_460)
);

OAI21xp5_ASAP7_75t_SL g462 ( 
.A1(n_460),
.A2(n_461),
.B(n_457),
.Y(n_462)
);

OAI321xp33_ASAP7_75t_L g464 ( 
.A1(n_462),
.A2(n_463),
.A3(n_6),
.B1(n_7),
.B2(n_9),
.C(n_10),
.Y(n_464)
);

AO22x1_ASAP7_75t_L g465 ( 
.A1(n_464),
.A2(n_7),
.B1(n_9),
.B2(n_10),
.Y(n_465)
);

AOI221xp5_ASAP7_75t_L g466 ( 
.A1(n_465),
.A2(n_7),
.B1(n_9),
.B2(n_10),
.C(n_11),
.Y(n_466)
);

XOR2xp5_ASAP7_75t_L g467 ( 
.A(n_466),
.B(n_11),
.Y(n_467)
);


endmodule