module fake_jpeg_31263_n_492 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_492);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_492;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_490;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_8),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_4),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_0),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

BUFx16f_ASAP7_75t_L g21 ( 
.A(n_15),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_6),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

BUFx10_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_6),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_4),
.Y(n_33)
);

CKINVDCx16_ASAP7_75t_R g34 ( 
.A(n_2),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_12),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_4),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_3),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_5),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_13),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_13),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_7),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_14),
.Y(n_42)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_6),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_2),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_5),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_7),
.B(n_15),
.Y(n_46)
);

INVx2_ASAP7_75t_SL g47 ( 
.A(n_12),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_8),
.Y(n_48)
);

INVxp67_ASAP7_75t_L g49 ( 
.A(n_4),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_11),
.Y(n_50)
);

INVx11_ASAP7_75t_L g51 ( 
.A(n_21),
.Y(n_51)
);

INVx5_ASAP7_75t_L g106 ( 
.A(n_51),
.Y(n_106)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_26),
.Y(n_52)
);

INVx5_ASAP7_75t_L g119 ( 
.A(n_52),
.Y(n_119)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_25),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_53),
.Y(n_107)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_43),
.Y(n_54)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_54),
.Y(n_104)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_25),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_55),
.Y(n_128)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_25),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g148 ( 
.A(n_56),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_46),
.B(n_8),
.Y(n_57)
);

AND2x2_ASAP7_75t_L g115 ( 
.A(n_57),
.B(n_74),
.Y(n_115)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_26),
.Y(n_58)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_58),
.Y(n_100)
);

BUFx24_ASAP7_75t_L g59 ( 
.A(n_21),
.Y(n_59)
);

INVx5_ASAP7_75t_L g123 ( 
.A(n_59),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_25),
.Y(n_60)
);

INVx6_ASAP7_75t_L g146 ( 
.A(n_60),
.Y(n_146)
);

INVx13_ASAP7_75t_L g61 ( 
.A(n_21),
.Y(n_61)
);

INVx5_ASAP7_75t_L g135 ( 
.A(n_61),
.Y(n_135)
);

INVx13_ASAP7_75t_L g62 ( 
.A(n_21),
.Y(n_62)
);

INVx5_ASAP7_75t_L g145 ( 
.A(n_62),
.Y(n_145)
);

INVx11_ASAP7_75t_L g63 ( 
.A(n_21),
.Y(n_63)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_63),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_30),
.Y(n_64)
);

INVx8_ASAP7_75t_L g101 ( 
.A(n_64),
.Y(n_101)
);

BUFx12f_ASAP7_75t_L g65 ( 
.A(n_30),
.Y(n_65)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_65),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_46),
.B(n_8),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_66),
.B(n_17),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_30),
.Y(n_67)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_67),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_SL g68 ( 
.A(n_46),
.B(n_9),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_68),
.B(n_88),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_30),
.Y(n_69)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_69),
.Y(n_121)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_26),
.Y(n_70)
);

INVx3_ASAP7_75t_L g130 ( 
.A(n_70),
.Y(n_130)
);

BUFx5_ASAP7_75t_L g71 ( 
.A(n_35),
.Y(n_71)
);

INVx4_ASAP7_75t_L g105 ( 
.A(n_71),
.Y(n_105)
);

INVx11_ASAP7_75t_L g72 ( 
.A(n_24),
.Y(n_72)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_72),
.Y(n_103)
);

INVx5_ASAP7_75t_L g73 ( 
.A(n_35),
.Y(n_73)
);

INVx4_ASAP7_75t_L g127 ( 
.A(n_73),
.Y(n_127)
);

AND2x2_ASAP7_75t_L g74 ( 
.A(n_43),
.B(n_9),
.Y(n_74)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_43),
.Y(n_75)
);

INVx3_ASAP7_75t_L g131 ( 
.A(n_75),
.Y(n_131)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_35),
.Y(n_76)
);

INVx3_ASAP7_75t_L g134 ( 
.A(n_76),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_35),
.Y(n_77)
);

INVx3_ASAP7_75t_L g137 ( 
.A(n_77),
.Y(n_137)
);

BUFx2_ASAP7_75t_L g78 ( 
.A(n_24),
.Y(n_78)
);

INVx3_ASAP7_75t_L g138 ( 
.A(n_78),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_24),
.Y(n_79)
);

INVx3_ASAP7_75t_L g139 ( 
.A(n_79),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_24),
.Y(n_80)
);

INVx3_ASAP7_75t_L g140 ( 
.A(n_80),
.Y(n_140)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_44),
.Y(n_81)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_81),
.Y(n_116)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_44),
.Y(n_82)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_82),
.Y(n_132)
);

INVx5_ASAP7_75t_L g83 ( 
.A(n_44),
.Y(n_83)
);

INVx4_ASAP7_75t_L g141 ( 
.A(n_83),
.Y(n_141)
);

BUFx3_ASAP7_75t_L g84 ( 
.A(n_44),
.Y(n_84)
);

INVx4_ASAP7_75t_L g150 ( 
.A(n_84),
.Y(n_150)
);

INVx8_ASAP7_75t_L g85 ( 
.A(n_27),
.Y(n_85)
);

INVx4_ASAP7_75t_L g155 ( 
.A(n_85),
.Y(n_155)
);

INVx11_ASAP7_75t_L g86 ( 
.A(n_34),
.Y(n_86)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_86),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_47),
.Y(n_87)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_87),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_49),
.B(n_9),
.Y(n_88)
);

BUFx12_ASAP7_75t_L g89 ( 
.A(n_34),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_89),
.B(n_95),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_47),
.Y(n_90)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_90),
.Y(n_110)
);

BUFx5_ASAP7_75t_L g91 ( 
.A(n_47),
.Y(n_91)
);

OR2x2_ASAP7_75t_L g112 ( 
.A(n_91),
.B(n_19),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_47),
.Y(n_92)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_92),
.Y(n_124)
);

BUFx3_ASAP7_75t_L g93 ( 
.A(n_20),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_93),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_27),
.Y(n_94)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_94),
.Y(n_153)
);

INVx13_ASAP7_75t_L g95 ( 
.A(n_27),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_27),
.Y(n_96)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_96),
.Y(n_154)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_23),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_97),
.B(n_98),
.Y(n_143)
);

INVx5_ASAP7_75t_L g98 ( 
.A(n_27),
.Y(n_98)
);

INVx11_ASAP7_75t_L g99 ( 
.A(n_27),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_99),
.B(n_19),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_L g108 ( 
.A1(n_53),
.A2(n_22),
.B1(n_48),
.B2(n_42),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g177 ( 
.A1(n_108),
.A2(n_111),
.B1(n_114),
.B2(n_117),
.Y(n_177)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_78),
.A2(n_45),
.B1(n_29),
.B2(n_18),
.Y(n_111)
);

CKINVDCx16_ASAP7_75t_R g176 ( 
.A(n_112),
.Y(n_176)
);

AOI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_76),
.A2(n_45),
.B1(n_29),
.B2(n_18),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_84),
.A2(n_45),
.B1(n_29),
.B2(n_18),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_52),
.A2(n_17),
.B1(n_50),
.B2(n_22),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_122),
.A2(n_126),
.B1(n_92),
.B2(n_90),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_125),
.B(n_129),
.Y(n_159)
);

AOI22xp33_ASAP7_75t_L g126 ( 
.A1(n_55),
.A2(n_20),
.B1(n_48),
.B2(n_42),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_97),
.B(n_41),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_74),
.B(n_41),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_133),
.B(n_144),
.Y(n_192)
);

NAND2x1_ASAP7_75t_L g136 ( 
.A(n_89),
.B(n_59),
.Y(n_136)
);

AO22x1_ASAP7_75t_L g168 ( 
.A1(n_136),
.A2(n_86),
.B1(n_59),
.B2(n_95),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_75),
.B(n_40),
.Y(n_144)
);

INVxp67_ASAP7_75t_L g161 ( 
.A(n_151),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_93),
.B(n_40),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_152),
.B(n_37),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_109),
.B(n_89),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_156),
.B(n_157),
.Y(n_212)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_116),
.Y(n_158)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_158),
.Y(n_229)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_132),
.Y(n_160)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_160),
.Y(n_243)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_104),
.Y(n_162)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_162),
.Y(n_223)
);

INVx3_ASAP7_75t_L g163 ( 
.A(n_123),
.Y(n_163)
);

INVx4_ASAP7_75t_L g208 ( 
.A(n_163),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_115),
.B(n_37),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_SL g215 ( 
.A(n_164),
.B(n_167),
.Y(n_215)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_147),
.Y(n_165)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_165),
.Y(n_234)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_131),
.Y(n_166)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_166),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_115),
.B(n_112),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_L g216 ( 
.A(n_168),
.B(n_136),
.Y(n_216)
);

INVx3_ASAP7_75t_L g169 ( 
.A(n_123),
.Y(n_169)
);

INVx4_ASAP7_75t_L g217 ( 
.A(n_169),
.Y(n_217)
);

INVx3_ASAP7_75t_L g170 ( 
.A(n_102),
.Y(n_170)
);

INVx3_ASAP7_75t_L g231 ( 
.A(n_170),
.Y(n_231)
);

INVx3_ASAP7_75t_L g171 ( 
.A(n_106),
.Y(n_171)
);

INVx3_ASAP7_75t_L g244 ( 
.A(n_171),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_143),
.A2(n_56),
.B1(n_60),
.B2(n_64),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_L g211 ( 
.A1(n_172),
.A2(n_117),
.B1(n_122),
.B2(n_168),
.Y(n_211)
);

AOI22xp33_ASAP7_75t_SL g173 ( 
.A1(n_120),
.A2(n_70),
.B1(n_73),
.B2(n_58),
.Y(n_173)
);

AOI22xp33_ASAP7_75t_SL g236 ( 
.A1(n_173),
.A2(n_190),
.B1(n_199),
.B2(n_203),
.Y(n_236)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_110),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_174),
.B(n_182),
.Y(n_218)
);

INVx3_ASAP7_75t_L g175 ( 
.A(n_106),
.Y(n_175)
);

INVx6_ASAP7_75t_L g241 ( 
.A(n_175),
.Y(n_241)
);

A2O1A1Ixp33_ASAP7_75t_L g178 ( 
.A1(n_142),
.A2(n_39),
.B(n_33),
.C(n_31),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_178),
.B(n_32),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_179),
.A2(n_201),
.B1(n_177),
.B2(n_101),
.Y(n_222)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_103),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_180),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_114),
.A2(n_77),
.B1(n_67),
.B2(n_69),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_181),
.A2(n_196),
.B1(n_99),
.B2(n_105),
.Y(n_251)
);

INVxp67_ASAP7_75t_L g182 ( 
.A(n_130),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_124),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_183),
.B(n_186),
.Y(n_221)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_134),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_184),
.Y(n_210)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_139),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_185),
.Y(n_219)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_153),
.Y(n_186)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_140),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_187),
.Y(n_230)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_121),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_188),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_SL g189 ( 
.A(n_135),
.B(n_23),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_189),
.B(n_191),
.Y(n_227)
);

BUFx6f_ASAP7_75t_L g190 ( 
.A(n_146),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_154),
.Y(n_191)
);

AOI22xp33_ASAP7_75t_L g193 ( 
.A1(n_146),
.A2(n_72),
.B1(n_79),
.B2(n_80),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_193),
.A2(n_172),
.B1(n_101),
.B2(n_128),
.Y(n_220)
);

INVx3_ASAP7_75t_L g194 ( 
.A(n_135),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_194),
.B(n_195),
.Y(n_242)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_100),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_111),
.A2(n_17),
.B1(n_83),
.B2(n_19),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_149),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_197),
.B(n_198),
.Y(n_249)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_108),
.Y(n_198)
);

INVx3_ASAP7_75t_L g199 ( 
.A(n_145),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_113),
.B(n_33),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_200),
.B(n_202),
.Y(n_214)
);

OAI22xp33_ASAP7_75t_SL g201 ( 
.A1(n_107),
.A2(n_87),
.B1(n_96),
.B2(n_94),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_145),
.B(n_31),
.Y(n_202)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_137),
.Y(n_203)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_138),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_204),
.B(n_205),
.Y(n_224)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_126),
.Y(n_205)
);

INVx2_ASAP7_75t_SL g206 ( 
.A(n_118),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_206),
.B(n_207),
.Y(n_246)
);

HB1xp67_ASAP7_75t_L g207 ( 
.A(n_150),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_211),
.A2(n_216),
.B1(n_220),
.B2(n_232),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_161),
.B(n_176),
.C(n_192),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g269 ( 
.A(n_213),
.B(n_226),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_222),
.A2(n_225),
.B1(n_228),
.B2(n_190),
.Y(n_258)
);

AOI22xp33_ASAP7_75t_L g225 ( 
.A1(n_185),
.A2(n_128),
.B1(n_148),
.B2(n_107),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_159),
.B(n_61),
.Y(n_226)
);

AOI22xp33_ASAP7_75t_L g228 ( 
.A1(n_187),
.A2(n_148),
.B1(n_203),
.B2(n_188),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_161),
.A2(n_65),
.B1(n_150),
.B2(n_141),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_SL g279 ( 
.A(n_235),
.B(n_248),
.Y(n_279)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_200),
.B(n_62),
.Y(n_237)
);

XOR2xp5_ASAP7_75t_L g275 ( 
.A(n_237),
.B(n_239),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_178),
.B(n_33),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_238),
.B(n_32),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_202),
.B(n_48),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_L g240 ( 
.A1(n_158),
.A2(n_127),
.B1(n_141),
.B2(n_155),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_240),
.A2(n_247),
.B1(n_182),
.B2(n_163),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_SL g245 ( 
.A(n_194),
.B(n_199),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_SL g277 ( 
.A(n_245),
.B(n_36),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_L g247 ( 
.A1(n_160),
.A2(n_127),
.B1(n_155),
.B2(n_119),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_166),
.B(n_28),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_L g267 ( 
.A1(n_251),
.A2(n_169),
.B1(n_85),
.B2(n_98),
.Y(n_267)
);

AOI22xp33_ASAP7_75t_SL g252 ( 
.A1(n_236),
.A2(n_119),
.B1(n_105),
.B2(n_175),
.Y(n_252)
);

OAI21xp5_ASAP7_75t_SL g309 ( 
.A1(n_252),
.A2(n_267),
.B(n_282),
.Y(n_309)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_246),
.Y(n_253)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_253),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_SL g300 ( 
.A(n_254),
.B(n_278),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_214),
.B(n_239),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_255),
.B(n_257),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_214),
.B(n_170),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_258),
.A2(n_261),
.B1(n_267),
.B2(n_271),
.Y(n_293)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_259),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_227),
.B(n_212),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_260),
.B(n_265),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_222),
.A2(n_184),
.B1(n_65),
.B2(n_204),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_211),
.A2(n_216),
.B1(n_220),
.B2(n_235),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_262),
.A2(n_263),
.B1(n_272),
.B2(n_270),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_238),
.A2(n_180),
.B1(n_171),
.B2(n_206),
.Y(n_263)
);

INVxp67_ASAP7_75t_L g264 ( 
.A(n_245),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_264),
.B(n_274),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_215),
.B(n_206),
.Y(n_265)
);

BUFx3_ASAP7_75t_L g266 ( 
.A(n_241),
.Y(n_266)
);

INVx4_ASAP7_75t_L g295 ( 
.A(n_266),
.Y(n_295)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_246),
.Y(n_268)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_268),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_237),
.B(n_38),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_270),
.B(n_280),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_251),
.A2(n_63),
.B1(n_51),
.B2(n_32),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_226),
.A2(n_50),
.B1(n_42),
.B2(n_39),
.Y(n_272)
);

AOI22x1_ASAP7_75t_SL g273 ( 
.A1(n_249),
.A2(n_50),
.B1(n_39),
.B2(n_38),
.Y(n_273)
);

OAI31xp33_ASAP7_75t_SL g326 ( 
.A1(n_273),
.A2(n_278),
.A3(n_1),
.B(n_3),
.Y(n_326)
);

INVxp67_ASAP7_75t_L g274 ( 
.A(n_218),
.Y(n_274)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_224),
.Y(n_276)
);

INVx1_ASAP7_75t_SL g306 ( 
.A(n_276),
.Y(n_306)
);

OAI21xp33_ASAP7_75t_L g316 ( 
.A1(n_277),
.A2(n_217),
.B(n_250),
.Y(n_316)
);

O2A1O1Ixp33_ASAP7_75t_L g278 ( 
.A1(n_224),
.A2(n_38),
.B(n_36),
.C(n_31),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_215),
.B(n_36),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_232),
.A2(n_28),
.B1(n_22),
.B2(n_20),
.Y(n_281)
);

AOI21xp5_ASAP7_75t_L g297 ( 
.A1(n_281),
.A2(n_282),
.B(n_0),
.Y(n_297)
);

AOI21xp5_ASAP7_75t_L g282 ( 
.A1(n_242),
.A2(n_28),
.B(n_10),
.Y(n_282)
);

INVx4_ASAP7_75t_L g283 ( 
.A(n_208),
.Y(n_283)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_283),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_221),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_284),
.B(n_291),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_213),
.A2(n_248),
.B1(n_223),
.B2(n_219),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_285),
.A2(n_286),
.B1(n_247),
.B2(n_240),
.Y(n_303)
);

OAI22xp33_ASAP7_75t_SL g286 ( 
.A1(n_223),
.A2(n_7),
.B1(n_15),
.B2(n_13),
.Y(n_286)
);

AND2x2_ASAP7_75t_SL g287 ( 
.A(n_234),
.B(n_0),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_L g311 ( 
.A(n_287),
.B(n_243),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_234),
.B(n_6),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_288),
.B(n_289),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_209),
.B(n_0),
.Y(n_289)
);

BUFx3_ASAP7_75t_L g290 ( 
.A(n_241),
.Y(n_290)
);

INVx2_ASAP7_75t_L g318 ( 
.A(n_290),
.Y(n_318)
);

INVx2_ASAP7_75t_L g291 ( 
.A(n_250),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_L g328 ( 
.A1(n_292),
.A2(n_296),
.B1(n_298),
.B2(n_313),
.Y(n_328)
);

OAI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_262),
.A2(n_233),
.B1(n_219),
.B2(n_230),
.Y(n_296)
);

OAI21xp5_ASAP7_75t_SL g344 ( 
.A1(n_297),
.A2(n_317),
.B(n_286),
.Y(n_344)
);

OAI22xp5_ASAP7_75t_L g298 ( 
.A1(n_256),
.A2(n_230),
.B1(n_233),
.B2(n_210),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_300),
.B(n_327),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_SL g301 ( 
.A(n_280),
.B(n_210),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_SL g333 ( 
.A(n_301),
.B(n_260),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_303),
.B(n_259),
.Y(n_330)
);

XNOR2x1_ASAP7_75t_L g305 ( 
.A(n_269),
.B(n_209),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_L g338 ( 
.A(n_305),
.B(n_311),
.Y(n_338)
);

AOI22xp5_ASAP7_75t_SL g307 ( 
.A1(n_261),
.A2(n_217),
.B1(n_208),
.B2(n_244),
.Y(n_307)
);

INVxp67_ASAP7_75t_L g348 ( 
.A(n_307),
.Y(n_348)
);

AOI21x1_ASAP7_75t_L g331 ( 
.A1(n_309),
.A2(n_252),
.B(n_273),
.Y(n_331)
);

OAI22xp5_ASAP7_75t_SL g313 ( 
.A1(n_256),
.A2(n_243),
.B1(n_229),
.B2(n_231),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_L g314 ( 
.A1(n_253),
.A2(n_231),
.B1(n_229),
.B2(n_244),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_L g335 ( 
.A1(n_314),
.A2(n_271),
.B1(n_283),
.B2(n_290),
.Y(n_335)
);

NAND3xp33_ASAP7_75t_L g329 ( 
.A(n_316),
.B(n_277),
.C(n_265),
.Y(n_329)
);

AOI21xp5_ASAP7_75t_L g317 ( 
.A1(n_268),
.A2(n_10),
.B(n_15),
.Y(n_317)
);

AOI22xp5_ASAP7_75t_L g320 ( 
.A1(n_258),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_320)
);

OAI22xp5_ASAP7_75t_SL g334 ( 
.A1(n_320),
.A2(n_323),
.B1(n_263),
.B2(n_288),
.Y(n_334)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_289),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g332 ( 
.A(n_321),
.Y(n_332)
);

XNOR2xp5_ASAP7_75t_SL g322 ( 
.A(n_269),
.B(n_3),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g358 ( 
.A(n_322),
.B(n_275),
.C(n_290),
.Y(n_358)
);

AOI22xp5_ASAP7_75t_L g323 ( 
.A1(n_276),
.A2(n_1),
.B1(n_3),
.B2(n_5),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g325 ( 
.A(n_266),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g341 ( 
.A(n_325),
.Y(n_341)
);

OA22x2_ASAP7_75t_L g351 ( 
.A1(n_326),
.A2(n_278),
.B1(n_287),
.B2(n_291),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_257),
.B(n_1),
.Y(n_327)
);

INVxp67_ASAP7_75t_L g370 ( 
.A(n_329),
.Y(n_370)
);

OAI22xp5_ASAP7_75t_L g368 ( 
.A1(n_330),
.A2(n_335),
.B1(n_304),
.B2(n_303),
.Y(n_368)
);

OAI21xp5_ASAP7_75t_L g366 ( 
.A1(n_331),
.A2(n_342),
.B(n_317),
.Y(n_366)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_333),
.Y(n_382)
);

AOI22xp5_ASAP7_75t_L g361 ( 
.A1(n_334),
.A2(n_343),
.B1(n_350),
.B2(n_292),
.Y(n_361)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_319),
.Y(n_336)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_336),
.Y(n_387)
);

NOR2xp33_ASAP7_75t_L g337 ( 
.A(n_308),
.B(n_284),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_SL g369 ( 
.A(n_337),
.B(n_340),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_SL g340 ( 
.A(n_310),
.B(n_285),
.Y(n_340)
);

OAI21xp5_ASAP7_75t_L g342 ( 
.A1(n_297),
.A2(n_254),
.B(n_279),
.Y(n_342)
);

OAI22xp5_ASAP7_75t_SL g343 ( 
.A1(n_293),
.A2(n_279),
.B1(n_255),
.B2(n_273),
.Y(n_343)
);

AOI21xp5_ASAP7_75t_L g373 ( 
.A1(n_344),
.A2(n_326),
.B(n_309),
.Y(n_373)
);

AOI22xp5_ASAP7_75t_L g345 ( 
.A1(n_298),
.A2(n_275),
.B1(n_287),
.B2(n_283),
.Y(n_345)
);

OAI22xp5_ASAP7_75t_SL g386 ( 
.A1(n_345),
.A2(n_327),
.B1(n_324),
.B2(n_323),
.Y(n_386)
);

CKINVDCx20_ASAP7_75t_R g346 ( 
.A(n_319),
.Y(n_346)
);

CKINVDCx20_ASAP7_75t_R g365 ( 
.A(n_346),
.Y(n_365)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_294),
.Y(n_347)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_347),
.Y(n_372)
);

INVxp67_ASAP7_75t_L g349 ( 
.A(n_314),
.Y(n_349)
);

INVxp67_ASAP7_75t_L g384 ( 
.A(n_349),
.Y(n_384)
);

OAI22xp5_ASAP7_75t_SL g350 ( 
.A1(n_293),
.A2(n_281),
.B1(n_272),
.B2(n_287),
.Y(n_350)
);

AND2x2_ASAP7_75t_L g376 ( 
.A(n_351),
.B(n_307),
.Y(n_376)
);

CKINVDCx16_ASAP7_75t_R g352 ( 
.A(n_315),
.Y(n_352)
);

NOR2xp33_ASAP7_75t_L g367 ( 
.A(n_352),
.B(n_356),
.Y(n_367)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_294),
.Y(n_353)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_353),
.Y(n_374)
);

INVx2_ASAP7_75t_L g354 ( 
.A(n_318),
.Y(n_354)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_354),
.Y(n_377)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_312),
.Y(n_355)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_355),
.Y(n_378)
);

NOR2xp33_ASAP7_75t_L g356 ( 
.A(n_308),
.B(n_315),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_312),
.Y(n_357)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_357),
.Y(n_388)
);

MAJx2_ASAP7_75t_L g363 ( 
.A(n_358),
.B(n_310),
.C(n_306),
.Y(n_363)
);

BUFx12f_ASAP7_75t_L g359 ( 
.A(n_295),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_L g380 ( 
.A(n_359),
.B(n_295),
.Y(n_380)
);

XNOR2xp5_ASAP7_75t_L g360 ( 
.A(n_338),
.B(n_305),
.Y(n_360)
);

XNOR2xp5_ASAP7_75t_L g392 ( 
.A(n_360),
.B(n_362),
.Y(n_392)
);

OAI22xp5_ASAP7_75t_SL g404 ( 
.A1(n_361),
.A2(n_371),
.B1(n_381),
.B2(n_328),
.Y(n_404)
);

XNOR2xp5_ASAP7_75t_L g362 ( 
.A(n_338),
.B(n_322),
.Y(n_362)
);

XOR2xp5_ASAP7_75t_L g400 ( 
.A(n_363),
.B(n_366),
.Y(n_400)
);

MAJIxp5_ASAP7_75t_L g364 ( 
.A(n_358),
.B(n_299),
.C(n_311),
.Y(n_364)
);

MAJIxp5_ASAP7_75t_L g402 ( 
.A(n_364),
.B(n_375),
.C(n_339),
.Y(n_402)
);

AOI22xp5_ASAP7_75t_L g391 ( 
.A1(n_368),
.A2(n_386),
.B1(n_334),
.B2(n_348),
.Y(n_391)
);

AOI22xp5_ASAP7_75t_L g371 ( 
.A1(n_349),
.A2(n_296),
.B1(n_304),
.B2(n_313),
.Y(n_371)
);

CKINVDCx14_ASAP7_75t_R g393 ( 
.A(n_373),
.Y(n_393)
);

MAJIxp5_ASAP7_75t_L g375 ( 
.A(n_345),
.B(n_299),
.C(n_306),
.Y(n_375)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_376),
.Y(n_394)
);

AOI21xp5_ASAP7_75t_L g379 ( 
.A1(n_348),
.A2(n_300),
.B(n_301),
.Y(n_379)
);

NOR2xp33_ASAP7_75t_L g401 ( 
.A(n_379),
.B(n_351),
.Y(n_401)
);

CKINVDCx20_ASAP7_75t_R g403 ( 
.A(n_380),
.Y(n_403)
);

AOI22xp5_ASAP7_75t_L g381 ( 
.A1(n_350),
.A2(n_321),
.B1(n_325),
.B2(n_320),
.Y(n_381)
);

NOR2xp33_ASAP7_75t_L g383 ( 
.A(n_333),
.B(n_324),
.Y(n_383)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_383),
.Y(n_406)
);

CKINVDCx20_ASAP7_75t_R g385 ( 
.A(n_341),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_SL g389 ( 
.A(n_385),
.B(n_332),
.Y(n_389)
);

CKINVDCx16_ASAP7_75t_R g428 ( 
.A(n_389),
.Y(n_428)
);

OAI22xp5_ASAP7_75t_L g390 ( 
.A1(n_382),
.A2(n_332),
.B1(n_328),
.B2(n_335),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_390),
.B(n_410),
.Y(n_421)
);

OAI22xp5_ASAP7_75t_SL g427 ( 
.A1(n_391),
.A2(n_396),
.B1(n_409),
.B2(n_377),
.Y(n_427)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_372),
.Y(n_395)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_395),
.Y(n_414)
);

AOI22xp5_ASAP7_75t_L g396 ( 
.A1(n_384),
.A2(n_343),
.B1(n_336),
.B2(n_346),
.Y(n_396)
);

XNOR2xp5_ASAP7_75t_L g397 ( 
.A(n_364),
.B(n_342),
.Y(n_397)
);

MAJIxp5_ASAP7_75t_L g415 ( 
.A(n_397),
.B(n_398),
.C(n_402),
.Y(n_415)
);

XNOR2xp5_ASAP7_75t_L g398 ( 
.A(n_363),
.B(n_339),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_372),
.Y(n_399)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_399),
.Y(n_419)
);

OAI21xp33_ASAP7_75t_L g420 ( 
.A1(n_401),
.A2(n_376),
.B(n_378),
.Y(n_420)
);

AOI22xp5_ASAP7_75t_L g423 ( 
.A1(n_404),
.A2(n_408),
.B1(n_388),
.B2(n_374),
.Y(n_423)
);

XOR2xp5_ASAP7_75t_L g405 ( 
.A(n_360),
.B(n_331),
.Y(n_405)
);

MAJIxp5_ASAP7_75t_L g416 ( 
.A(n_405),
.B(n_375),
.C(n_366),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_365),
.B(n_353),
.Y(n_407)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_407),
.Y(n_424)
);

OAI22xp5_ASAP7_75t_SL g408 ( 
.A1(n_361),
.A2(n_357),
.B1(n_355),
.B2(n_347),
.Y(n_408)
);

AOI22xp5_ASAP7_75t_L g409 ( 
.A1(n_384),
.A2(n_341),
.B1(n_344),
.B2(n_351),
.Y(n_409)
);

OAI22xp5_ASAP7_75t_L g410 ( 
.A1(n_369),
.A2(n_370),
.B1(n_381),
.B2(n_367),
.Y(n_410)
);

HB1xp67_ASAP7_75t_L g411 ( 
.A(n_387),
.Y(n_411)
);

NOR2xp33_ASAP7_75t_L g426 ( 
.A(n_411),
.B(n_412),
.Y(n_426)
);

OAI22xp5_ASAP7_75t_L g412 ( 
.A1(n_370),
.A2(n_351),
.B1(n_354),
.B2(n_318),
.Y(n_412)
);

OAI22xp5_ASAP7_75t_L g413 ( 
.A1(n_409),
.A2(n_376),
.B1(n_373),
.B2(n_371),
.Y(n_413)
);

AOI22xp5_ASAP7_75t_L g438 ( 
.A1(n_413),
.A2(n_427),
.B1(n_404),
.B2(n_394),
.Y(n_438)
);

XOR2xp5_ASAP7_75t_L g432 ( 
.A(n_416),
.B(n_420),
.Y(n_432)
);

NOR2xp33_ASAP7_75t_SL g417 ( 
.A(n_406),
.B(n_379),
.Y(n_417)
);

OAI22xp5_ASAP7_75t_L g433 ( 
.A1(n_417),
.A2(n_418),
.B1(n_393),
.B2(n_403),
.Y(n_433)
);

AOI21xp33_ASAP7_75t_L g418 ( 
.A1(n_407),
.A2(n_388),
.B(n_378),
.Y(n_418)
);

MAJIxp5_ASAP7_75t_L g422 ( 
.A(n_402),
.B(n_386),
.C(n_362),
.Y(n_422)
);

MAJIxp5_ASAP7_75t_L g440 ( 
.A(n_422),
.B(n_425),
.C(n_398),
.Y(n_440)
);

OAI22xp5_ASAP7_75t_SL g436 ( 
.A1(n_423),
.A2(n_391),
.B1(n_429),
.B2(n_426),
.Y(n_436)
);

MAJIxp5_ASAP7_75t_L g425 ( 
.A(n_397),
.B(n_374),
.C(n_377),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_SL g429 ( 
.A(n_396),
.B(n_302),
.Y(n_429)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_429),
.Y(n_434)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_395),
.Y(n_430)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_430),
.Y(n_435)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_399),
.Y(n_431)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_431),
.Y(n_437)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_433),
.Y(n_456)
);

XOR2xp5_ASAP7_75t_L g453 ( 
.A(n_436),
.B(n_419),
.Y(n_453)
);

OAI22xp5_ASAP7_75t_SL g449 ( 
.A1(n_438),
.A2(n_427),
.B1(n_425),
.B2(n_416),
.Y(n_449)
);

OR2x2_ASAP7_75t_L g439 ( 
.A(n_424),
.B(n_394),
.Y(n_439)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_439),
.Y(n_461)
);

XNOR2xp5_ASAP7_75t_L g460 ( 
.A(n_440),
.B(n_441),
.Y(n_460)
);

XNOR2xp5_ASAP7_75t_L g441 ( 
.A(n_422),
.B(n_400),
.Y(n_441)
);

OAI22xp5_ASAP7_75t_SL g442 ( 
.A1(n_421),
.A2(n_408),
.B1(n_400),
.B2(n_405),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_SL g452 ( 
.A(n_442),
.B(n_443),
.Y(n_452)
);

OAI22xp5_ASAP7_75t_SL g443 ( 
.A1(n_421),
.A2(n_359),
.B1(n_302),
.B2(n_392),
.Y(n_443)
);

AOI21xp5_ASAP7_75t_L g444 ( 
.A1(n_417),
.A2(n_392),
.B(n_266),
.Y(n_444)
);

NAND3xp33_ASAP7_75t_SL g450 ( 
.A(n_444),
.B(n_445),
.C(n_446),
.Y(n_450)
);

OAI21xp5_ASAP7_75t_SL g445 ( 
.A1(n_413),
.A2(n_424),
.B(n_426),
.Y(n_445)
);

OAI21xp5_ASAP7_75t_L g446 ( 
.A1(n_423),
.A2(n_359),
.B(n_10),
.Y(n_446)
);

MAJIxp5_ASAP7_75t_L g447 ( 
.A(n_415),
.B(n_359),
.C(n_10),
.Y(n_447)
);

MAJIxp5_ASAP7_75t_L g451 ( 
.A(n_447),
.B(n_414),
.C(n_419),
.Y(n_451)
);

AOI22xp33_ASAP7_75t_SL g448 ( 
.A1(n_435),
.A2(n_431),
.B1(n_430),
.B2(n_414),
.Y(n_448)
);

CKINVDCx20_ASAP7_75t_R g471 ( 
.A(n_448),
.Y(n_471)
);

AOI22xp5_ASAP7_75t_L g472 ( 
.A1(n_449),
.A2(n_446),
.B1(n_11),
.B2(n_16),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_SL g462 ( 
.A(n_451),
.B(n_457),
.Y(n_462)
);

XOR2xp5_ASAP7_75t_L g463 ( 
.A(n_453),
.B(n_445),
.Y(n_463)
);

OAI22xp5_ASAP7_75t_SL g454 ( 
.A1(n_438),
.A2(n_428),
.B1(n_415),
.B2(n_12),
.Y(n_454)
);

AOI22xp5_ASAP7_75t_L g468 ( 
.A1(n_454),
.A2(n_437),
.B1(n_435),
.B2(n_434),
.Y(n_468)
);

MAJIxp5_ASAP7_75t_L g455 ( 
.A(n_440),
.B(n_428),
.C(n_11),
.Y(n_455)
);

MAJIxp5_ASAP7_75t_L g466 ( 
.A(n_455),
.B(n_458),
.C(n_437),
.Y(n_466)
);

NOR2xp33_ASAP7_75t_L g457 ( 
.A(n_447),
.B(n_5),
.Y(n_457)
);

MAJIxp5_ASAP7_75t_L g458 ( 
.A(n_441),
.B(n_11),
.C(n_16),
.Y(n_458)
);

NOR2xp33_ASAP7_75t_L g459 ( 
.A(n_443),
.B(n_436),
.Y(n_459)
);

NOR2xp33_ASAP7_75t_L g470 ( 
.A(n_459),
.B(n_442),
.Y(n_470)
);

XNOR2xp5_ASAP7_75t_L g476 ( 
.A(n_463),
.B(n_468),
.Y(n_476)
);

NOR2xp33_ASAP7_75t_SL g464 ( 
.A(n_455),
.B(n_432),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_SL g479 ( 
.A(n_464),
.B(n_465),
.Y(n_479)
);

NOR2xp33_ASAP7_75t_SL g465 ( 
.A(n_456),
.B(n_432),
.Y(n_465)
);

NOR2xp33_ASAP7_75t_L g473 ( 
.A(n_466),
.B(n_467),
.Y(n_473)
);

NOR2xp33_ASAP7_75t_SL g467 ( 
.A(n_460),
.B(n_444),
.Y(n_467)
);

OAI21xp5_ASAP7_75t_L g469 ( 
.A1(n_461),
.A2(n_439),
.B(n_434),
.Y(n_469)
);

OR2x2_ASAP7_75t_L g477 ( 
.A(n_469),
.B(n_470),
.Y(n_477)
);

MAJIxp5_ASAP7_75t_L g478 ( 
.A(n_472),
.B(n_453),
.C(n_451),
.Y(n_478)
);

OAI21xp5_ASAP7_75t_L g474 ( 
.A1(n_471),
.A2(n_461),
.B(n_452),
.Y(n_474)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_474),
.Y(n_480)
);

NOR2xp33_ASAP7_75t_SL g475 ( 
.A(n_462),
.B(n_460),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_SL g481 ( 
.A(n_475),
.B(n_454),
.Y(n_481)
);

NOR2xp33_ASAP7_75t_L g482 ( 
.A(n_478),
.B(n_463),
.Y(n_482)
);

AOI21x1_ASAP7_75t_L g485 ( 
.A1(n_481),
.A2(n_473),
.B(n_469),
.Y(n_485)
);

NOR2xp33_ASAP7_75t_L g484 ( 
.A(n_482),
.B(n_483),
.Y(n_484)
);

INVxp67_ASAP7_75t_L g483 ( 
.A(n_479),
.Y(n_483)
);

OAI21xp5_ASAP7_75t_SL g488 ( 
.A1(n_485),
.A2(n_484),
.B(n_458),
.Y(n_488)
);

OAI21xp33_ASAP7_75t_L g486 ( 
.A1(n_480),
.A2(n_477),
.B(n_476),
.Y(n_486)
);

NOR3xp33_ASAP7_75t_L g487 ( 
.A(n_486),
.B(n_478),
.C(n_477),
.Y(n_487)
);

AOI22xp5_ASAP7_75t_SL g489 ( 
.A1(n_487),
.A2(n_488),
.B1(n_449),
.B2(n_450),
.Y(n_489)
);

BUFx24_ASAP7_75t_SL g490 ( 
.A(n_489),
.Y(n_490)
);

OAI21xp5_ASAP7_75t_L g491 ( 
.A1(n_490),
.A2(n_466),
.B(n_472),
.Y(n_491)
);

AOI21xp5_ASAP7_75t_L g492 ( 
.A1(n_491),
.A2(n_16),
.B(n_484),
.Y(n_492)
);


endmodule