module fake_netlist_6_3271_n_1037 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_235, n_256, n_298, n_18, n_21, n_193, n_147, n_269, n_258, n_281, n_154, n_191, n_88, n_3, n_209, n_98, n_277, n_260, n_265, n_283, n_113, n_39, n_63, n_223, n_278, n_270, n_73, n_279, n_4, n_148, n_199, n_138, n_22, n_161, n_208, n_68, n_226, n_228, n_252, n_266, n_296, n_166, n_28, n_184, n_212, n_268, n_271, n_50, n_158, n_49, n_7, n_210, n_216, n_83, n_206, n_217, n_299, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_215, n_297, n_178, n_247, n_225, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_227, n_132, n_188, n_102, n_186, n_204, n_245, n_0, n_87, n_195, n_285, n_261, n_189, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_213, n_164, n_257, n_100, n_292, n_129, n_13, n_121, n_294, n_197, n_11, n_137, n_17, n_23, n_203, n_254, n_142, n_286, n_20, n_143, n_207, n_2, n_242, n_180, n_19, n_47, n_62, n_29, n_155, n_219, n_291, n_75, n_109, n_150, n_233, n_263, n_122, n_264, n_45, n_255, n_284, n_205, n_34, n_140, n_218, n_70, n_120, n_234, n_251, n_301, n_214, n_274, n_37, n_15, n_67, n_33, n_82, n_27, n_236, n_246, n_38, n_110, n_151, n_289, n_61, n_112, n_172, n_237, n_81, n_59, n_244, n_181, n_76, n_36, n_182, n_26, n_124, n_238, n_239, n_55, n_126, n_202, n_94, n_97, n_108, n_267, n_282, n_58, n_116, n_280, n_211, n_287, n_64, n_220, n_288, n_290, n_117, n_118, n_175, n_224, n_48, n_231, n_65, n_230, n_25, n_40, n_93, n_80, n_141, n_240, n_135, n_196, n_200, n_165, n_139, n_41, n_134, n_259, n_177, n_176, n_273, n_114, n_86, n_198, n_104, n_222, n_95, n_179, n_243, n_9, n_248, n_300, n_107, n_10, n_295, n_71, n_74, n_229, n_253, n_6, n_190, n_14, n_123, n_262, n_136, n_72, n_187, n_89, n_249, n_173, n_201, n_250, n_103, n_111, n_60, n_159, n_272, n_157, n_162, n_170, n_185, n_35, n_183, n_232, n_115, n_12, n_69, n_128, n_241, n_30, n_79, n_275, n_43, n_194, n_171, n_293, n_31, n_192, n_57, n_169, n_53, n_276, n_51, n_44, n_56, n_221, n_1037);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_235;
input n_256;
input n_298;
input n_18;
input n_21;
input n_193;
input n_147;
input n_269;
input n_258;
input n_281;
input n_154;
input n_191;
input n_88;
input n_3;
input n_209;
input n_98;
input n_277;
input n_260;
input n_265;
input n_283;
input n_113;
input n_39;
input n_63;
input n_223;
input n_278;
input n_270;
input n_73;
input n_279;
input n_4;
input n_148;
input n_199;
input n_138;
input n_22;
input n_161;
input n_208;
input n_68;
input n_226;
input n_228;
input n_252;
input n_266;
input n_296;
input n_166;
input n_28;
input n_184;
input n_212;
input n_268;
input n_271;
input n_50;
input n_158;
input n_49;
input n_7;
input n_210;
input n_216;
input n_83;
input n_206;
input n_217;
input n_299;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_215;
input n_297;
input n_178;
input n_247;
input n_225;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_227;
input n_132;
input n_188;
input n_102;
input n_186;
input n_204;
input n_245;
input n_0;
input n_87;
input n_195;
input n_285;
input n_261;
input n_189;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_213;
input n_164;
input n_257;
input n_100;
input n_292;
input n_129;
input n_13;
input n_121;
input n_294;
input n_197;
input n_11;
input n_137;
input n_17;
input n_23;
input n_203;
input n_254;
input n_142;
input n_286;
input n_20;
input n_143;
input n_207;
input n_2;
input n_242;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_219;
input n_291;
input n_75;
input n_109;
input n_150;
input n_233;
input n_263;
input n_122;
input n_264;
input n_45;
input n_255;
input n_284;
input n_205;
input n_34;
input n_140;
input n_218;
input n_70;
input n_120;
input n_234;
input n_251;
input n_301;
input n_214;
input n_274;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_236;
input n_246;
input n_38;
input n_110;
input n_151;
input n_289;
input n_61;
input n_112;
input n_172;
input n_237;
input n_81;
input n_59;
input n_244;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_238;
input n_239;
input n_55;
input n_126;
input n_202;
input n_94;
input n_97;
input n_108;
input n_267;
input n_282;
input n_58;
input n_116;
input n_280;
input n_211;
input n_287;
input n_64;
input n_220;
input n_288;
input n_290;
input n_117;
input n_118;
input n_175;
input n_224;
input n_48;
input n_231;
input n_65;
input n_230;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_240;
input n_135;
input n_196;
input n_200;
input n_165;
input n_139;
input n_41;
input n_134;
input n_259;
input n_177;
input n_176;
input n_273;
input n_114;
input n_86;
input n_198;
input n_104;
input n_222;
input n_95;
input n_179;
input n_243;
input n_9;
input n_248;
input n_300;
input n_107;
input n_10;
input n_295;
input n_71;
input n_74;
input n_229;
input n_253;
input n_6;
input n_190;
input n_14;
input n_123;
input n_262;
input n_136;
input n_72;
input n_187;
input n_89;
input n_249;
input n_173;
input n_201;
input n_250;
input n_103;
input n_111;
input n_60;
input n_159;
input n_272;
input n_157;
input n_162;
input n_170;
input n_185;
input n_35;
input n_183;
input n_232;
input n_115;
input n_12;
input n_69;
input n_128;
input n_241;
input n_30;
input n_79;
input n_275;
input n_43;
input n_194;
input n_171;
input n_293;
input n_31;
input n_192;
input n_57;
input n_169;
input n_53;
input n_276;
input n_51;
input n_44;
input n_56;
input n_221;

output n_1037;

wire n_992;
wire n_591;
wire n_435;
wire n_793;
wire n_326;
wire n_801;
wire n_853;
wire n_440;
wire n_587;
wire n_695;
wire n_507;
wire n_968;
wire n_909;
wire n_580;
wire n_762;
wire n_1030;
wire n_881;
wire n_875;
wire n_465;
wire n_680;
wire n_367;
wire n_760;
wire n_741;
wire n_1008;
wire n_1027;
wire n_590;
wire n_625;
wire n_661;
wire n_362;
wire n_341;
wire n_828;
wire n_462;
wire n_671;
wire n_607;
wire n_726;
wire n_1033;
wire n_316;
wire n_419;
wire n_304;
wire n_700;
wire n_694;
wire n_933;
wire n_740;
wire n_578;
wire n_703;
wire n_1003;
wire n_365;
wire n_978;
wire n_384;
wire n_595;
wire n_627;
wire n_524;
wire n_342;
wire n_820;
wire n_951;
wire n_783;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_751;
wire n_449;
wire n_749;
wire n_798;
wire n_310;
wire n_509;
wire n_368;
wire n_575;
wire n_994;
wire n_677;
wire n_969;
wire n_988;
wire n_805;
wire n_396;
wire n_495;
wire n_815;
wire n_350;
wire n_585;
wire n_732;
wire n_974;
wire n_568;
wire n_392;
wire n_840;
wire n_442;
wire n_874;
wire n_480;
wire n_724;
wire n_382;
wire n_673;
wire n_1020;
wire n_1009;
wire n_628;
wire n_883;
wire n_557;
wire n_823;
wire n_349;
wire n_643;
wire n_617;
wire n_698;
wire n_898;
wire n_1032;
wire n_845;
wire n_807;
wire n_1036;
wire n_739;
wire n_400;
wire n_337;
wire n_955;
wire n_865;
wire n_893;
wire n_925;
wire n_485;
wire n_1026;
wire n_443;
wire n_892;
wire n_768;
wire n_471;
wire n_935;
wire n_421;
wire n_781;
wire n_424;
wire n_789;
wire n_615;
wire n_573;
wire n_769;
wire n_320;
wire n_639;
wire n_676;
wire n_327;
wire n_794;
wire n_963;
wire n_727;
wire n_894;
wire n_369;
wire n_597;
wire n_685;
wire n_832;
wire n_353;
wire n_610;
wire n_555;
wire n_389;
wire n_814;
wire n_415;
wire n_830;
wire n_605;
wire n_461;
wire n_873;
wire n_383;
wire n_826;
wire n_1024;
wire n_669;
wire n_447;
wire n_872;
wire n_517;
wire n_718;
wire n_1018;
wire n_747;
wire n_852;
wire n_667;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_621;
wire n_305;
wire n_721;
wire n_996;
wire n_750;
wire n_532;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_468;
wire n_544;
wire n_901;
wire n_504;
wire n_923;
wire n_314;
wire n_378;
wire n_413;
wire n_377;
wire n_791;
wire n_510;
wire n_837;
wire n_836;
wire n_1015;
wire n_863;
wire n_375;
wire n_601;
wire n_338;
wire n_522;
wire n_948;
wire n_466;
wire n_704;
wire n_918;
wire n_748;
wire n_506;
wire n_763;
wire n_360;
wire n_945;
wire n_977;
wire n_603;
wire n_1005;
wire n_991;
wire n_957;
wire n_536;
wire n_895;
wire n_866;
wire n_622;
wire n_340;
wire n_710;
wire n_387;
wire n_452;
wire n_658;
wire n_616;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_581;
wire n_761;
wire n_428;
wire n_785;
wire n_746;
wire n_609;
wire n_765;
wire n_432;
wire n_987;
wire n_641;
wire n_822;
wire n_693;
wire n_631;
wire n_516;
wire n_720;
wire n_525;
wire n_758;
wire n_842;
wire n_611;
wire n_943;
wire n_491;
wire n_843;
wire n_656;
wire n_772;
wire n_989;
wire n_797;
wire n_666;
wire n_1016;
wire n_371;
wire n_795;
wire n_770;
wire n_940;
wire n_567;
wire n_899;
wire n_738;
wire n_405;
wire n_538;
wire n_1035;
wire n_838;
wire n_302;
wire n_499;
wire n_380;
wire n_705;
wire n_647;
wire n_343;
wire n_844;
wire n_448;
wire n_886;
wire n_953;
wire n_1004;
wire n_1017;
wire n_494;
wire n_539;
wire n_493;
wire n_397;
wire n_1022;
wire n_614;
wire n_529;
wire n_445;
wire n_425;
wire n_684;
wire n_930;
wire n_888;
wire n_454;
wire n_638;
wire n_910;
wire n_486;
wire n_911;
wire n_381;
wire n_947;
wire n_653;
wire n_887;
wire n_752;
wire n_908;
wire n_944;
wire n_713;
wire n_648;
wire n_657;
wire n_576;
wire n_1028;
wire n_472;
wire n_414;
wire n_563;
wire n_782;
wire n_976;
wire n_490;
wire n_803;
wire n_809;
wire n_1011;
wire n_926;
wire n_927;
wire n_839;
wire n_986;
wire n_734;
wire n_708;
wire n_919;
wire n_402;
wire n_352;
wire n_917;
wire n_668;
wire n_478;
wire n_626;
wire n_990;
wire n_574;
wire n_779;
wire n_800;
wire n_929;
wire n_460;
wire n_907;
wire n_854;
wire n_417;
wire n_446;
wire n_498;
wire n_662;
wire n_374;
wire n_659;
wire n_709;
wire n_870;
wire n_366;
wire n_904;
wire n_777;
wire n_407;
wire n_913;
wire n_450;
wire n_808;
wire n_867;
wire n_526;
wire n_921;
wire n_712;
wire n_348;
wire n_711;
wire n_579;
wire n_376;
wire n_937;
wire n_390;
wire n_473;
wire n_334;
wire n_559;
wire n_370;
wire n_458;
wire n_650;
wire n_998;
wire n_717;
wire n_330;
wire n_771;
wire n_470;
wire n_475;
wire n_924;
wire n_492;
wire n_972;
wire n_551;
wire n_699;
wire n_456;
wire n_564;
wire n_313;
wire n_624;
wire n_451;
wire n_824;
wire n_962;
wire n_1000;
wire n_686;
wire n_796;
wire n_757;
wire n_565;
wire n_594;
wire n_719;
wire n_356;
wire n_577;
wire n_936;
wire n_552;
wire n_619;
wire n_885;
wire n_455;
wire n_896;
wire n_521;
wire n_363;
wire n_572;
wire n_912;
wire n_395;
wire n_813;
wire n_592;
wire n_745;
wire n_654;
wire n_323;
wire n_829;
wire n_606;
wire n_393;
wire n_818;
wire n_984;
wire n_411;
wire n_503;
wire n_716;
wire n_623;
wire n_884;
wire n_599;
wire n_513;
wire n_776;
wire n_321;
wire n_645;
wire n_331;
wire n_916;
wire n_868;
wire n_570;
wire n_731;
wire n_859;
wire n_406;
wire n_483;
wire n_735;
wire n_482;
wire n_934;
wire n_755;
wire n_931;
wire n_1021;
wire n_527;
wire n_608;
wire n_683;
wire n_474;
wire n_620;
wire n_420;
wire n_878;
wire n_630;
wire n_312;
wire n_394;
wire n_519;
wire n_541;
wire n_512;
wire n_958;
wire n_307;
wire n_469;
wire n_433;
wire n_500;
wire n_942;
wire n_792;
wire n_880;
wire n_476;
wire n_981;
wire n_714;
wire n_543;
wire n_889;
wire n_357;
wire n_985;
wire n_589;
wire n_860;
wire n_481;
wire n_788;
wire n_819;
wire n_939;
wire n_997;
wire n_821;
wire n_325;
wire n_938;
wire n_767;
wire n_804;
wire n_329;
wire n_600;
wire n_464;
wire n_831;
wire n_802;
wire n_982;
wire n_964;
wire n_561;
wire n_477;
wire n_549;
wire n_980;
wire n_533;
wire n_954;
wire n_408;
wire n_932;
wire n_806;
wire n_864;
wire n_879;
wire n_959;
wire n_584;
wire n_399;
wire n_979;
wire n_548;
wire n_905;
wire n_436;
wire n_833;
wire n_523;
wire n_707;
wire n_322;
wire n_993;
wire n_345;
wire n_409;
wire n_354;
wire n_689;
wire n_799;
wire n_505;
wire n_756;
wire n_319;
wire n_547;
wire n_537;
wire n_558;
wire n_810;
wire n_635;
wire n_787;
wire n_311;
wire n_403;
wire n_723;
wire n_634;
wire n_583;
wire n_596;
wire n_966;
wire n_546;
wire n_562;
wire n_386;
wire n_764;
wire n_556;
wire n_1034;
wire n_692;
wire n_733;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_487;
wire n_550;
wire n_553;
wire n_652;
wire n_849;
wire n_970;
wire n_560;
wire n_1014;
wire n_753;
wire n_642;
wire n_995;
wire n_569;
wire n_441;
wire n_811;
wire n_882;
wire n_444;
wire n_586;
wire n_423;
wire n_737;
wire n_318;
wire n_303;
wire n_511;
wire n_715;
wire n_467;
wire n_306;
wire n_359;
wire n_973;
wire n_346;
wire n_416;
wire n_530;
wire n_520;
wire n_1029;
wire n_418;
wire n_618;
wire n_790;
wire n_582;
wire n_861;
wire n_674;
wire n_857;
wire n_871;
wire n_967;
wire n_775;
wire n_922;
wire n_571;
wire n_404;
wire n_651;
wire n_439;
wire n_518;
wire n_679;
wire n_612;
wire n_453;
wire n_633;
wire n_665;
wire n_902;
wire n_333;
wire n_588;
wire n_308;
wire n_309;
wire n_914;
wire n_759;
wire n_1010;
wire n_355;
wire n_426;
wire n_317;
wire n_915;
wire n_632;
wire n_702;
wire n_431;
wire n_347;
wire n_812;
wire n_459;
wire n_502;
wire n_328;
wire n_672;
wire n_534;
wire n_488;
wire n_429;
wire n_1006;
wire n_373;
wire n_1012;
wire n_497;
wire n_780;
wire n_773;
wire n_675;
wire n_920;
wire n_903;
wire n_730;
wire n_655;
wire n_706;
wire n_786;
wire n_670;
wire n_834;
wire n_835;
wire n_928;
wire n_690;
wire n_850;
wire n_401;
wire n_324;
wire n_743;
wire n_766;
wire n_816;
wire n_335;
wire n_430;
wire n_1002;
wire n_463;
wire n_545;
wire n_489;
wire n_877;
wire n_604;
wire n_848;
wire n_1019;
wire n_825;
wire n_636;
wire n_728;
wire n_681;
wire n_729;
wire n_876;
wire n_774;
wire n_412;
wire n_640;
wire n_660;
wire n_965;
wire n_438;
wire n_339;
wire n_784;
wire n_315;
wire n_515;
wire n_434;
wire n_983;
wire n_427;
wire n_479;
wire n_598;
wire n_496;
wire n_422;
wire n_696;
wire n_906;
wire n_688;
wire n_722;
wire n_961;
wire n_862;
wire n_869;
wire n_351;
wire n_437;
wire n_540;
wire n_593;
wire n_514;
wire n_646;
wire n_528;
wire n_391;
wire n_457;
wire n_687;
wire n_697;
wire n_364;
wire n_890;
wire n_637;
wire n_385;
wire n_701;
wire n_817;
wire n_950;
wire n_629;
wire n_388;
wire n_858;
wire n_484;
wire n_613;
wire n_736;
wire n_897;
wire n_900;
wire n_846;
wire n_501;
wire n_841;
wire n_956;
wire n_960;
wire n_531;
wire n_827;
wire n_1001;
wire n_361;
wire n_508;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1025;
wire n_332;
wire n_891;
wire n_336;
wire n_410;
wire n_398;
wire n_566;
wire n_554;
wire n_602;
wire n_1023;
wire n_1013;
wire n_664;
wire n_949;
wire n_678;
wire n_1007;
wire n_649;
wire n_855;

INVxp67_ASAP7_75t_L g302 ( 
.A(n_19),
.Y(n_302)
);

CKINVDCx16_ASAP7_75t_R g303 ( 
.A(n_74),
.Y(n_303)
);

INVxp67_ASAP7_75t_L g304 ( 
.A(n_178),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_211),
.Y(n_305)
);

BUFx3_ASAP7_75t_L g306 ( 
.A(n_301),
.Y(n_306)
);

INVx2_ASAP7_75t_L g307 ( 
.A(n_13),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_158),
.Y(n_308)
);

INVxp33_ASAP7_75t_L g309 ( 
.A(n_10),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_147),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_275),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_218),
.Y(n_312)
);

INVx2_ASAP7_75t_L g313 ( 
.A(n_234),
.Y(n_313)
);

INVxp67_ASAP7_75t_L g314 ( 
.A(n_133),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_204),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_107),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_220),
.Y(n_317)
);

INVx2_ASAP7_75t_L g318 ( 
.A(n_138),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_70),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_66),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_299),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_127),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_108),
.Y(n_323)
);

INVxp67_ASAP7_75t_L g324 ( 
.A(n_254),
.Y(n_324)
);

INVx2_ASAP7_75t_L g325 ( 
.A(n_189),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_157),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_267),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_82),
.Y(n_328)
);

BUFx3_ASAP7_75t_L g329 ( 
.A(n_185),
.Y(n_329)
);

INVxp67_ASAP7_75t_L g330 ( 
.A(n_10),
.Y(n_330)
);

BUFx6f_ASAP7_75t_L g331 ( 
.A(n_271),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_2),
.Y(n_332)
);

INVx2_ASAP7_75t_L g333 ( 
.A(n_288),
.Y(n_333)
);

INVx2_ASAP7_75t_L g334 ( 
.A(n_60),
.Y(n_334)
);

INVx2_ASAP7_75t_L g335 ( 
.A(n_153),
.Y(n_335)
);

INVxp33_ASAP7_75t_SL g336 ( 
.A(n_202),
.Y(n_336)
);

INVx2_ASAP7_75t_L g337 ( 
.A(n_36),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_247),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_194),
.Y(n_339)
);

CKINVDCx14_ASAP7_75t_R g340 ( 
.A(n_273),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_110),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_175),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_237),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_276),
.Y(n_344)
);

HB1xp67_ASAP7_75t_L g345 ( 
.A(n_135),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_236),
.Y(n_346)
);

INVxp67_ASAP7_75t_SL g347 ( 
.A(n_228),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_73),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_22),
.Y(n_349)
);

INVxp33_ASAP7_75t_L g350 ( 
.A(n_69),
.Y(n_350)
);

INVx2_ASAP7_75t_L g351 ( 
.A(n_243),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_129),
.Y(n_352)
);

INVxp33_ASAP7_75t_SL g353 ( 
.A(n_199),
.Y(n_353)
);

INVx2_ASAP7_75t_L g354 ( 
.A(n_143),
.Y(n_354)
);

INVxp33_ASAP7_75t_SL g355 ( 
.A(n_90),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_131),
.Y(n_356)
);

CKINVDCx20_ASAP7_75t_R g357 ( 
.A(n_38),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_286),
.Y(n_358)
);

CKINVDCx14_ASAP7_75t_R g359 ( 
.A(n_251),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_113),
.Y(n_360)
);

CKINVDCx14_ASAP7_75t_R g361 ( 
.A(n_119),
.Y(n_361)
);

BUFx6f_ASAP7_75t_L g362 ( 
.A(n_246),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_39),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_48),
.Y(n_364)
);

INVxp67_ASAP7_75t_L g365 ( 
.A(n_156),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_31),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_28),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_277),
.Y(n_368)
);

BUFx2_ASAP7_75t_L g369 ( 
.A(n_222),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_284),
.Y(n_370)
);

BUFx2_ASAP7_75t_L g371 ( 
.A(n_103),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_64),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_268),
.Y(n_373)
);

INVxp67_ASAP7_75t_SL g374 ( 
.A(n_109),
.Y(n_374)
);

INVx3_ASAP7_75t_L g375 ( 
.A(n_184),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_1),
.Y(n_376)
);

INVxp67_ASAP7_75t_SL g377 ( 
.A(n_77),
.Y(n_377)
);

CKINVDCx20_ASAP7_75t_R g378 ( 
.A(n_215),
.Y(n_378)
);

INVxp67_ASAP7_75t_SL g379 ( 
.A(n_249),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_176),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_231),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_50),
.Y(n_382)
);

INVxp33_ASAP7_75t_SL g383 ( 
.A(n_45),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_160),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_97),
.Y(n_385)
);

CKINVDCx20_ASAP7_75t_R g386 ( 
.A(n_76),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_161),
.Y(n_387)
);

INVx2_ASAP7_75t_L g388 ( 
.A(n_270),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_244),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_126),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_14),
.Y(n_391)
);

INVxp67_ASAP7_75t_L g392 ( 
.A(n_219),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_100),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_272),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_144),
.Y(n_395)
);

INVxp67_ASAP7_75t_SL g396 ( 
.A(n_188),
.Y(n_396)
);

BUFx3_ASAP7_75t_L g397 ( 
.A(n_150),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_35),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_289),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_279),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_125),
.Y(n_401)
);

INVx1_ASAP7_75t_SL g402 ( 
.A(n_163),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_212),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_101),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_34),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_173),
.Y(n_406)
);

INVxp67_ASAP7_75t_L g407 ( 
.A(n_6),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_151),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_68),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_134),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_72),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_6),
.Y(n_412)
);

INVxp67_ASAP7_75t_SL g413 ( 
.A(n_136),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_5),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_269),
.Y(n_415)
);

INVxp33_ASAP7_75t_L g416 ( 
.A(n_182),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_79),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_298),
.Y(n_418)
);

CKINVDCx20_ASAP7_75t_R g419 ( 
.A(n_198),
.Y(n_419)
);

INVxp33_ASAP7_75t_SL g420 ( 
.A(n_83),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_122),
.Y(n_421)
);

CKINVDCx20_ASAP7_75t_R g422 ( 
.A(n_104),
.Y(n_422)
);

INVxp67_ASAP7_75t_SL g423 ( 
.A(n_89),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_214),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_281),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_259),
.Y(n_426)
);

INVx2_ASAP7_75t_L g427 ( 
.A(n_87),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_37),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_179),
.Y(n_429)
);

CKINVDCx20_ASAP7_75t_R g430 ( 
.A(n_25),
.Y(n_430)
);

CKINVDCx20_ASAP7_75t_R g431 ( 
.A(n_300),
.Y(n_431)
);

BUFx2_ASAP7_75t_L g432 ( 
.A(n_105),
.Y(n_432)
);

INVxp67_ASAP7_75t_L g433 ( 
.A(n_291),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_137),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_278),
.Y(n_435)
);

CKINVDCx20_ASAP7_75t_R g436 ( 
.A(n_32),
.Y(n_436)
);

INVx2_ASAP7_75t_L g437 ( 
.A(n_258),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_106),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_167),
.Y(n_439)
);

INVx2_ASAP7_75t_L g440 ( 
.A(n_210),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_250),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_142),
.Y(n_442)
);

INVxp67_ASAP7_75t_SL g443 ( 
.A(n_123),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_55),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_12),
.Y(n_445)
);

INVxp33_ASAP7_75t_L g446 ( 
.A(n_116),
.Y(n_446)
);

INVxp67_ASAP7_75t_SL g447 ( 
.A(n_95),
.Y(n_447)
);

OR2x2_ASAP7_75t_L g448 ( 
.A(n_213),
.B(n_260),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_155),
.Y(n_449)
);

CKINVDCx16_ASAP7_75t_R g450 ( 
.A(n_67),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_232),
.Y(n_451)
);

CKINVDCx20_ASAP7_75t_R g452 ( 
.A(n_280),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_196),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_230),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_208),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_49),
.Y(n_456)
);

CKINVDCx14_ASAP7_75t_R g457 ( 
.A(n_297),
.Y(n_457)
);

INVxp33_ASAP7_75t_L g458 ( 
.A(n_27),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_248),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_145),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_92),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_111),
.Y(n_462)
);

INVxp67_ASAP7_75t_SL g463 ( 
.A(n_148),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_86),
.Y(n_464)
);

CKINVDCx20_ASAP7_75t_R g465 ( 
.A(n_63),
.Y(n_465)
);

BUFx5_ASAP7_75t_L g466 ( 
.A(n_140),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_43),
.Y(n_467)
);

INVxp33_ASAP7_75t_L g468 ( 
.A(n_139),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_168),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_174),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_290),
.Y(n_471)
);

CKINVDCx14_ASAP7_75t_R g472 ( 
.A(n_217),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_229),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_132),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_264),
.Y(n_475)
);

CKINVDCx20_ASAP7_75t_R g476 ( 
.A(n_65),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_245),
.Y(n_477)
);

BUFx3_ASAP7_75t_L g478 ( 
.A(n_233),
.Y(n_478)
);

CKINVDCx16_ASAP7_75t_R g479 ( 
.A(n_12),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_61),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_4),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_221),
.Y(n_482)
);

INVx2_ASAP7_75t_L g483 ( 
.A(n_225),
.Y(n_483)
);

INVxp33_ASAP7_75t_SL g484 ( 
.A(n_2),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_192),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_154),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_88),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_203),
.Y(n_488)
);

INVxp67_ASAP7_75t_L g489 ( 
.A(n_285),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_52),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_146),
.Y(n_491)
);

BUFx2_ASAP7_75t_SL g492 ( 
.A(n_209),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_293),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_307),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_332),
.Y(n_495)
);

INVx2_ASAP7_75t_L g496 ( 
.A(n_466),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_376),
.Y(n_497)
);

INVx2_ASAP7_75t_L g498 ( 
.A(n_466),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_412),
.Y(n_499)
);

INVx2_ASAP7_75t_L g500 ( 
.A(n_466),
.Y(n_500)
);

INVx3_ASAP7_75t_L g501 ( 
.A(n_414),
.Y(n_501)
);

AND2x4_ASAP7_75t_L g502 ( 
.A(n_306),
.B(n_0),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_445),
.Y(n_503)
);

OAI22xp5_ASAP7_75t_SL g504 ( 
.A1(n_479),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_504)
);

INVx2_ASAP7_75t_L g505 ( 
.A(n_466),
.Y(n_505)
);

INVx2_ASAP7_75t_L g506 ( 
.A(n_466),
.Y(n_506)
);

INVx2_ASAP7_75t_L g507 ( 
.A(n_481),
.Y(n_507)
);

INVx2_ASAP7_75t_L g508 ( 
.A(n_329),
.Y(n_508)
);

NOR2x1_ASAP7_75t_L g509 ( 
.A(n_375),
.B(n_23),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_305),
.Y(n_510)
);

OA21x2_ASAP7_75t_L g511 ( 
.A1(n_308),
.A2(n_3),
.B(n_4),
.Y(n_511)
);

AND2x2_ASAP7_75t_L g512 ( 
.A(n_369),
.B(n_5),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_310),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_L g514 ( 
.A(n_375),
.B(n_7),
.Y(n_514)
);

INVx3_ASAP7_75t_L g515 ( 
.A(n_391),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_311),
.Y(n_516)
);

OR2x2_ASAP7_75t_L g517 ( 
.A(n_302),
.B(n_7),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_L g518 ( 
.A(n_371),
.B(n_8),
.Y(n_518)
);

INVx2_ASAP7_75t_L g519 ( 
.A(n_397),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_312),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_315),
.Y(n_521)
);

INVxp67_ASAP7_75t_L g522 ( 
.A(n_302),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_SL g523 ( 
.A(n_303),
.B(n_8),
.Y(n_523)
);

INVx2_ASAP7_75t_L g524 ( 
.A(n_478),
.Y(n_524)
);

HB1xp67_ASAP7_75t_L g525 ( 
.A(n_330),
.Y(n_525)
);

INVx3_ASAP7_75t_L g526 ( 
.A(n_331),
.Y(n_526)
);

BUFx6f_ASAP7_75t_L g527 ( 
.A(n_331),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_L g528 ( 
.A(n_432),
.B(n_9),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_316),
.Y(n_529)
);

NAND2xp33_ASAP7_75t_SL g530 ( 
.A(n_309),
.B(n_9),
.Y(n_530)
);

INVx2_ASAP7_75t_L g531 ( 
.A(n_331),
.Y(n_531)
);

INVx2_ASAP7_75t_L g532 ( 
.A(n_362),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_317),
.Y(n_533)
);

NOR2xp33_ASAP7_75t_L g534 ( 
.A(n_350),
.B(n_11),
.Y(n_534)
);

NAND2xp33_ASAP7_75t_L g535 ( 
.A(n_345),
.B(n_11),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_319),
.Y(n_536)
);

AND2x2_ASAP7_75t_L g537 ( 
.A(n_340),
.B(n_13),
.Y(n_537)
);

AND2x4_ASAP7_75t_L g538 ( 
.A(n_313),
.B(n_14),
.Y(n_538)
);

BUFx2_ASAP7_75t_L g539 ( 
.A(n_330),
.Y(n_539)
);

INVx2_ASAP7_75t_L g540 ( 
.A(n_362),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_SL g541 ( 
.A(n_450),
.B(n_15),
.Y(n_541)
);

AND2x4_ASAP7_75t_L g542 ( 
.A(n_318),
.B(n_15),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_L g543 ( 
.A(n_325),
.B(n_16),
.Y(n_543)
);

BUFx6f_ASAP7_75t_L g544 ( 
.A(n_362),
.Y(n_544)
);

BUFx6f_ASAP7_75t_L g545 ( 
.A(n_333),
.Y(n_545)
);

HB1xp67_ASAP7_75t_L g546 ( 
.A(n_407),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_320),
.Y(n_547)
);

INVx2_ASAP7_75t_L g548 ( 
.A(n_321),
.Y(n_548)
);

BUFx6f_ASAP7_75t_L g549 ( 
.A(n_334),
.Y(n_549)
);

INVxp67_ASAP7_75t_L g550 ( 
.A(n_407),
.Y(n_550)
);

NOR2xp33_ASAP7_75t_L g551 ( 
.A(n_416),
.B(n_446),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_322),
.Y(n_552)
);

HB1xp67_ASAP7_75t_L g553 ( 
.A(n_484),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_326),
.Y(n_554)
);

BUFx2_ASAP7_75t_L g555 ( 
.A(n_357),
.Y(n_555)
);

AND2x4_ASAP7_75t_L g556 ( 
.A(n_335),
.B(n_16),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_328),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_339),
.Y(n_558)
);

INVx2_ASAP7_75t_L g559 ( 
.A(n_341),
.Y(n_559)
);

INVx3_ASAP7_75t_L g560 ( 
.A(n_342),
.Y(n_560)
);

INVx3_ASAP7_75t_L g561 ( 
.A(n_343),
.Y(n_561)
);

INVx2_ASAP7_75t_L g562 ( 
.A(n_344),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_346),
.Y(n_563)
);

INVx2_ASAP7_75t_L g564 ( 
.A(n_348),
.Y(n_564)
);

INVx2_ASAP7_75t_L g565 ( 
.A(n_349),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_356),
.Y(n_566)
);

INVx2_ASAP7_75t_L g567 ( 
.A(n_358),
.Y(n_567)
);

BUFx3_ASAP7_75t_L g568 ( 
.A(n_323),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_360),
.Y(n_569)
);

NOR2xp33_ASAP7_75t_L g570 ( 
.A(n_458),
.B(n_17),
.Y(n_570)
);

INVx1_ASAP7_75t_SL g571 ( 
.A(n_378),
.Y(n_571)
);

INVx2_ASAP7_75t_SL g572 ( 
.A(n_327),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_363),
.Y(n_573)
);

AND2x4_ASAP7_75t_L g574 ( 
.A(n_337),
.B(n_17),
.Y(n_574)
);

BUFx6f_ASAP7_75t_L g575 ( 
.A(n_351),
.Y(n_575)
);

INVx2_ASAP7_75t_L g576 ( 
.A(n_364),
.Y(n_576)
);

INVx3_ASAP7_75t_L g577 ( 
.A(n_366),
.Y(n_577)
);

NAND2xp33_ASAP7_75t_L g578 ( 
.A(n_468),
.B(n_18),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_368),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_L g580 ( 
.A(n_354),
.B(n_18),
.Y(n_580)
);

INVx2_ASAP7_75t_L g581 ( 
.A(n_372),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_373),
.Y(n_582)
);

NOR2xp33_ASAP7_75t_L g583 ( 
.A(n_304),
.B(n_19),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_381),
.Y(n_584)
);

INVx3_ASAP7_75t_L g585 ( 
.A(n_382),
.Y(n_585)
);

INVx2_ASAP7_75t_L g586 ( 
.A(n_385),
.Y(n_586)
);

NOR2xp33_ASAP7_75t_SL g587 ( 
.A(n_402),
.B(n_20),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_SL g588 ( 
.A(n_402),
.B(n_20),
.Y(n_588)
);

AND2x4_ASAP7_75t_L g589 ( 
.A(n_388),
.B(n_21),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_L g590 ( 
.A(n_427),
.B(n_21),
.Y(n_590)
);

AND2x6_ASAP7_75t_L g591 ( 
.A(n_437),
.B(n_24),
.Y(n_591)
);

HB1xp67_ASAP7_75t_L g592 ( 
.A(n_387),
.Y(n_592)
);

AND2x2_ASAP7_75t_L g593 ( 
.A(n_359),
.B(n_26),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_389),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_L g595 ( 
.A(n_440),
.B(n_29),
.Y(n_595)
);

INVx2_ASAP7_75t_L g596 ( 
.A(n_390),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_SL g597 ( 
.A(n_336),
.B(n_30),
.Y(n_597)
);

INVx2_ASAP7_75t_L g598 ( 
.A(n_393),
.Y(n_598)
);

AND2x4_ASAP7_75t_L g599 ( 
.A(n_483),
.B(n_33),
.Y(n_599)
);

INVx2_ASAP7_75t_L g600 ( 
.A(n_394),
.Y(n_600)
);

NOR2x1p5_ASAP7_75t_L g601 ( 
.A(n_518),
.B(n_528),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_526),
.Y(n_602)
);

AND2x2_ASAP7_75t_L g603 ( 
.A(n_551),
.B(n_361),
.Y(n_603)
);

BUFx3_ASAP7_75t_L g604 ( 
.A(n_568),
.Y(n_604)
);

INVx5_ASAP7_75t_L g605 ( 
.A(n_527),
.Y(n_605)
);

INVx2_ASAP7_75t_SL g606 ( 
.A(n_515),
.Y(n_606)
);

BUFx8_ASAP7_75t_SL g607 ( 
.A(n_555),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_L g608 ( 
.A(n_572),
.B(n_457),
.Y(n_608)
);

OR2x6_ASAP7_75t_L g609 ( 
.A(n_553),
.B(n_492),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_527),
.Y(n_610)
);

INVx3_ASAP7_75t_L g611 ( 
.A(n_545),
.Y(n_611)
);

AND2x6_ASAP7_75t_L g612 ( 
.A(n_599),
.B(n_395),
.Y(n_612)
);

CKINVDCx5p33_ASAP7_75t_R g613 ( 
.A(n_571),
.Y(n_613)
);

INVx2_ASAP7_75t_L g614 ( 
.A(n_527),
.Y(n_614)
);

INVx3_ASAP7_75t_L g615 ( 
.A(n_545),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_526),
.Y(n_616)
);

INVx2_ASAP7_75t_L g617 ( 
.A(n_544),
.Y(n_617)
);

INVx2_ASAP7_75t_L g618 ( 
.A(n_544),
.Y(n_618)
);

CKINVDCx5p33_ASAP7_75t_R g619 ( 
.A(n_515),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_544),
.Y(n_620)
);

INVx2_ASAP7_75t_L g621 ( 
.A(n_531),
.Y(n_621)
);

INVx4_ASAP7_75t_L g622 ( 
.A(n_593),
.Y(n_622)
);

NOR2xp33_ASAP7_75t_L g623 ( 
.A(n_512),
.B(n_534),
.Y(n_623)
);

INVx5_ASAP7_75t_L g624 ( 
.A(n_591),
.Y(n_624)
);

INVxp67_ASAP7_75t_L g625 ( 
.A(n_525),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_532),
.Y(n_626)
);

BUFx4f_ASAP7_75t_L g627 ( 
.A(n_591),
.Y(n_627)
);

OAI22xp5_ASAP7_75t_SL g628 ( 
.A1(n_504),
.A2(n_430),
.B1(n_386),
.B2(n_419),
.Y(n_628)
);

OR2x2_ASAP7_75t_L g629 ( 
.A(n_508),
.B(n_399),
.Y(n_629)
);

BUFx3_ASAP7_75t_L g630 ( 
.A(n_519),
.Y(n_630)
);

OAI22xp33_ASAP7_75t_SL g631 ( 
.A1(n_523),
.A2(n_353),
.B1(n_355),
.B2(n_383),
.Y(n_631)
);

HB1xp67_ASAP7_75t_L g632 ( 
.A(n_524),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_L g633 ( 
.A(n_599),
.B(n_472),
.Y(n_633)
);

BUFx3_ASAP7_75t_L g634 ( 
.A(n_545),
.Y(n_634)
);

INVx2_ASAP7_75t_L g635 ( 
.A(n_540),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_495),
.Y(n_636)
);

NOR2xp33_ASAP7_75t_L g637 ( 
.A(n_570),
.B(n_420),
.Y(n_637)
);

BUFx6f_ASAP7_75t_L g638 ( 
.A(n_549),
.Y(n_638)
);

BUFx3_ASAP7_75t_L g639 ( 
.A(n_549),
.Y(n_639)
);

HB1xp67_ASAP7_75t_L g640 ( 
.A(n_546),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_SL g641 ( 
.A(n_537),
.B(n_304),
.Y(n_641)
);

INVx3_ASAP7_75t_L g642 ( 
.A(n_549),
.Y(n_642)
);

CKINVDCx5p33_ASAP7_75t_R g643 ( 
.A(n_592),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_548),
.Y(n_644)
);

AOI22xp5_ASAP7_75t_L g645 ( 
.A1(n_541),
.A2(n_452),
.B1(n_476),
.B2(n_436),
.Y(n_645)
);

INVx2_ASAP7_75t_L g646 ( 
.A(n_575),
.Y(n_646)
);

INVx3_ASAP7_75t_L g647 ( 
.A(n_575),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_559),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_495),
.Y(n_649)
);

INVx1_ASAP7_75t_SL g650 ( 
.A(n_539),
.Y(n_650)
);

NAND3xp33_ASAP7_75t_L g651 ( 
.A(n_578),
.B(n_365),
.C(n_324),
.Y(n_651)
);

INVx4_ASAP7_75t_L g652 ( 
.A(n_575),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_L g653 ( 
.A(n_510),
.B(n_400),
.Y(n_653)
);

INVx2_ASAP7_75t_SL g654 ( 
.A(n_503),
.Y(n_654)
);

AND2x4_ASAP7_75t_L g655 ( 
.A(n_502),
.B(n_314),
.Y(n_655)
);

INVx4_ASAP7_75t_L g656 ( 
.A(n_591),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_562),
.Y(n_657)
);

AOI22xp33_ASAP7_75t_L g658 ( 
.A1(n_538),
.A2(n_556),
.B1(n_574),
.B2(n_542),
.Y(n_658)
);

HB1xp67_ASAP7_75t_L g659 ( 
.A(n_522),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_L g660 ( 
.A(n_513),
.B(n_516),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_564),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_SL g662 ( 
.A(n_502),
.B(n_324),
.Y(n_662)
);

NAND3x1_ASAP7_75t_L g663 ( 
.A(n_583),
.B(n_403),
.C(n_401),
.Y(n_663)
);

INVx2_ASAP7_75t_SL g664 ( 
.A(n_507),
.Y(n_664)
);

BUFx6f_ASAP7_75t_L g665 ( 
.A(n_538),
.Y(n_665)
);

INVx2_ASAP7_75t_L g666 ( 
.A(n_565),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_567),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_L g668 ( 
.A(n_520),
.B(n_404),
.Y(n_668)
);

AND2x4_ASAP7_75t_L g669 ( 
.A(n_542),
.B(n_556),
.Y(n_669)
);

AND2x6_ASAP7_75t_L g670 ( 
.A(n_509),
.B(n_405),
.Y(n_670)
);

AND2x4_ASAP7_75t_L g671 ( 
.A(n_574),
.B(n_347),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_L g672 ( 
.A(n_521),
.B(n_409),
.Y(n_672)
);

AND2x2_ASAP7_75t_L g673 ( 
.A(n_550),
.B(n_365),
.Y(n_673)
);

INVx3_ASAP7_75t_L g674 ( 
.A(n_501),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_576),
.Y(n_675)
);

INVx2_ASAP7_75t_SL g676 ( 
.A(n_497),
.Y(n_676)
);

INVx3_ASAP7_75t_L g677 ( 
.A(n_501),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_L g678 ( 
.A(n_529),
.B(n_533),
.Y(n_678)
);

INVx4_ASAP7_75t_L g679 ( 
.A(n_591),
.Y(n_679)
);

AND2x4_ASAP7_75t_L g680 ( 
.A(n_589),
.B(n_374),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_L g681 ( 
.A(n_536),
.B(n_410),
.Y(n_681)
);

AO22x2_ASAP7_75t_L g682 ( 
.A1(n_517),
.A2(n_448),
.B1(n_433),
.B2(n_392),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_581),
.Y(n_683)
);

INVx2_ASAP7_75t_SL g684 ( 
.A(n_497),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_586),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_L g686 ( 
.A(n_547),
.B(n_552),
.Y(n_686)
);

INVx2_ASAP7_75t_L g687 ( 
.A(n_596),
.Y(n_687)
);

NAND3xp33_ASAP7_75t_L g688 ( 
.A(n_514),
.B(n_433),
.C(n_392),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_598),
.Y(n_689)
);

NOR2xp33_ASAP7_75t_L g690 ( 
.A(n_543),
.B(n_489),
.Y(n_690)
);

INVx1_ASAP7_75t_SL g691 ( 
.A(n_554),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_L g692 ( 
.A(n_623),
.B(n_597),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_632),
.Y(n_693)
);

OR2x6_ASAP7_75t_L g694 ( 
.A(n_609),
.B(n_625),
.Y(n_694)
);

BUFx3_ASAP7_75t_L g695 ( 
.A(n_634),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_630),
.Y(n_696)
);

CKINVDCx5p33_ASAP7_75t_R g697 ( 
.A(n_613),
.Y(n_697)
);

BUFx6f_ASAP7_75t_L g698 ( 
.A(n_638),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_611),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_615),
.Y(n_700)
);

BUFx2_ASAP7_75t_L g701 ( 
.A(n_643),
.Y(n_701)
);

AND2x2_ASAP7_75t_SL g702 ( 
.A(n_645),
.B(n_535),
.Y(n_702)
);

INVxp67_ASAP7_75t_L g703 ( 
.A(n_659),
.Y(n_703)
);

INVx2_ASAP7_75t_SL g704 ( 
.A(n_650),
.Y(n_704)
);

INVxp67_ASAP7_75t_SL g705 ( 
.A(n_638),
.Y(n_705)
);

CKINVDCx11_ASAP7_75t_R g706 ( 
.A(n_609),
.Y(n_706)
);

AOI22xp5_ASAP7_75t_L g707 ( 
.A1(n_637),
.A2(n_530),
.B1(n_422),
.B2(n_431),
.Y(n_707)
);

AOI22xp5_ASAP7_75t_L g708 ( 
.A1(n_601),
.A2(n_465),
.B1(n_587),
.B2(n_588),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_642),
.Y(n_709)
);

AO22x1_ASAP7_75t_L g710 ( 
.A1(n_690),
.A2(n_589),
.B1(n_580),
.B2(n_590),
.Y(n_710)
);

BUFx6f_ASAP7_75t_L g711 ( 
.A(n_639),
.Y(n_711)
);

INVx2_ASAP7_75t_SL g712 ( 
.A(n_640),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_647),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_L g714 ( 
.A(n_603),
.B(n_557),
.Y(n_714)
);

AND2x2_ASAP7_75t_L g715 ( 
.A(n_691),
.B(n_600),
.Y(n_715)
);

OR2x4_ASAP7_75t_L g716 ( 
.A(n_629),
.B(n_499),
.Y(n_716)
);

OR2x2_ASAP7_75t_SL g717 ( 
.A(n_651),
.B(n_511),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_SL g718 ( 
.A(n_665),
.B(n_338),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_646),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_L g720 ( 
.A(n_622),
.B(n_558),
.Y(n_720)
);

INVx3_ASAP7_75t_L g721 ( 
.A(n_652),
.Y(n_721)
);

AOI22xp33_ASAP7_75t_L g722 ( 
.A1(n_671),
.A2(n_511),
.B1(n_569),
.B2(n_563),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_610),
.Y(n_723)
);

INVx2_ASAP7_75t_SL g724 ( 
.A(n_673),
.Y(n_724)
);

BUFx6f_ASAP7_75t_L g725 ( 
.A(n_665),
.Y(n_725)
);

INVx2_ASAP7_75t_L g726 ( 
.A(n_614),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_610),
.Y(n_727)
);

INVx2_ASAP7_75t_L g728 ( 
.A(n_617),
.Y(n_728)
);

INVx4_ASAP7_75t_L g729 ( 
.A(n_619),
.Y(n_729)
);

INVx5_ASAP7_75t_L g730 ( 
.A(n_670),
.Y(n_730)
);

INVx2_ASAP7_75t_L g731 ( 
.A(n_618),
.Y(n_731)
);

AOI22xp5_ASAP7_75t_L g732 ( 
.A1(n_631),
.A2(n_489),
.B1(n_595),
.B2(n_352),
.Y(n_732)
);

BUFx6f_ASAP7_75t_SL g733 ( 
.A(n_604),
.Y(n_733)
);

INVx1_ASAP7_75t_SL g734 ( 
.A(n_607),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_664),
.Y(n_735)
);

AND2x4_ASAP7_75t_L g736 ( 
.A(n_669),
.B(n_499),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_L g737 ( 
.A(n_622),
.B(n_566),
.Y(n_737)
);

INVx6_ASAP7_75t_L g738 ( 
.A(n_652),
.Y(n_738)
);

AND2x4_ASAP7_75t_L g739 ( 
.A(n_669),
.B(n_494),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_L g740 ( 
.A(n_612),
.B(n_573),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_620),
.Y(n_741)
);

AOI22xp33_ASAP7_75t_L g742 ( 
.A1(n_671),
.A2(n_594),
.B1(n_573),
.B2(n_584),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_666),
.Y(n_743)
);

INVx2_ASAP7_75t_L g744 ( 
.A(n_621),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_687),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_636),
.Y(n_746)
);

AND2x4_ASAP7_75t_L g747 ( 
.A(n_606),
.B(n_494),
.Y(n_747)
);

NOR2xp33_ASAP7_75t_L g748 ( 
.A(n_608),
.B(n_579),
.Y(n_748)
);

AND2x4_ASAP7_75t_L g749 ( 
.A(n_680),
.B(n_579),
.Y(n_749)
);

INVx2_ASAP7_75t_L g750 ( 
.A(n_635),
.Y(n_750)
);

BUFx6f_ASAP7_75t_L g751 ( 
.A(n_605),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_L g752 ( 
.A(n_612),
.B(n_582),
.Y(n_752)
);

INVx2_ASAP7_75t_L g753 ( 
.A(n_626),
.Y(n_753)
);

AND2x2_ASAP7_75t_L g754 ( 
.A(n_658),
.B(n_582),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_L g755 ( 
.A(n_612),
.B(n_584),
.Y(n_755)
);

OR2x2_ASAP7_75t_L g756 ( 
.A(n_662),
.B(n_560),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_636),
.Y(n_757)
);

BUFx2_ASAP7_75t_L g758 ( 
.A(n_682),
.Y(n_758)
);

BUFx6f_ASAP7_75t_L g759 ( 
.A(n_605),
.Y(n_759)
);

INVx2_ASAP7_75t_L g760 ( 
.A(n_644),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_649),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_SL g762 ( 
.A(n_680),
.B(n_367),
.Y(n_762)
);

AND2x2_ASAP7_75t_L g763 ( 
.A(n_674),
.B(n_594),
.Y(n_763)
);

INVx2_ASAP7_75t_L g764 ( 
.A(n_648),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_649),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_654),
.Y(n_766)
);

AND2x6_ASAP7_75t_SL g767 ( 
.A(n_628),
.B(n_411),
.Y(n_767)
);

INVx2_ASAP7_75t_L g768 ( 
.A(n_657),
.Y(n_768)
);

OAI22xp5_ASAP7_75t_L g769 ( 
.A1(n_641),
.A2(n_463),
.B1(n_377),
.B2(n_379),
.Y(n_769)
);

HB1xp67_ASAP7_75t_L g770 ( 
.A(n_677),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_L g771 ( 
.A(n_633),
.B(n_560),
.Y(n_771)
);

CKINVDCx8_ASAP7_75t_R g772 ( 
.A(n_670),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_602),
.Y(n_773)
);

BUFx2_ASAP7_75t_L g774 ( 
.A(n_704),
.Y(n_774)
);

AND2x4_ASAP7_75t_L g775 ( 
.A(n_736),
.B(n_655),
.Y(n_775)
);

OAI22xp33_ASAP7_75t_SL g776 ( 
.A1(n_692),
.A2(n_655),
.B1(n_454),
.B2(n_444),
.Y(n_776)
);

INVx2_ASAP7_75t_L g777 ( 
.A(n_744),
.Y(n_777)
);

AND2x4_ASAP7_75t_L g778 ( 
.A(n_736),
.B(n_676),
.Y(n_778)
);

NOR2xp33_ASAP7_75t_R g779 ( 
.A(n_697),
.B(n_370),
.Y(n_779)
);

INVx3_ASAP7_75t_L g780 ( 
.A(n_725),
.Y(n_780)
);

INVx3_ASAP7_75t_SL g781 ( 
.A(n_734),
.Y(n_781)
);

AOI21x1_ASAP7_75t_L g782 ( 
.A1(n_771),
.A2(n_668),
.B(n_653),
.Y(n_782)
);

AND2x2_ASAP7_75t_L g783 ( 
.A(n_715),
.B(n_684),
.Y(n_783)
);

INVx1_ASAP7_75t_SL g784 ( 
.A(n_701),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_L g785 ( 
.A(n_748),
.B(n_670),
.Y(n_785)
);

OR2x2_ASAP7_75t_L g786 ( 
.A(n_724),
.B(n_712),
.Y(n_786)
);

BUFx12f_ASAP7_75t_L g787 ( 
.A(n_706),
.Y(n_787)
);

AOI21xp5_ASAP7_75t_L g788 ( 
.A1(n_720),
.A2(n_627),
.B(n_656),
.Y(n_788)
);

INVx1_ASAP7_75t_L g789 ( 
.A(n_746),
.Y(n_789)
);

BUFx2_ASAP7_75t_L g790 ( 
.A(n_758),
.Y(n_790)
);

BUFx3_ASAP7_75t_L g791 ( 
.A(n_725),
.Y(n_791)
);

NOR2xp33_ASAP7_75t_L g792 ( 
.A(n_703),
.B(n_688),
.Y(n_792)
);

AOI221xp5_ASAP7_75t_L g793 ( 
.A1(n_708),
.A2(n_682),
.B1(n_672),
.B2(n_681),
.C(n_585),
.Y(n_793)
);

O2A1O1Ixp33_ASAP7_75t_L g794 ( 
.A1(n_769),
.A2(n_686),
.B(n_660),
.C(n_678),
.Y(n_794)
);

AND2x4_ASAP7_75t_L g795 ( 
.A(n_739),
.B(n_661),
.Y(n_795)
);

HB1xp67_ASAP7_75t_L g796 ( 
.A(n_701),
.Y(n_796)
);

INVx2_ASAP7_75t_L g797 ( 
.A(n_750),
.Y(n_797)
);

BUFx6f_ASAP7_75t_L g798 ( 
.A(n_698),
.Y(n_798)
);

AOI22xp5_ASAP7_75t_L g799 ( 
.A1(n_702),
.A2(n_663),
.B1(n_656),
.B2(n_679),
.Y(n_799)
);

NOR2xp33_ASAP7_75t_L g800 ( 
.A(n_729),
.B(n_679),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_757),
.Y(n_801)
);

BUFx6f_ASAP7_75t_L g802 ( 
.A(n_698),
.Y(n_802)
);

BUFx2_ASAP7_75t_L g803 ( 
.A(n_758),
.Y(n_803)
);

INVxp67_ASAP7_75t_SL g804 ( 
.A(n_721),
.Y(n_804)
);

HB1xp67_ASAP7_75t_L g805 ( 
.A(n_693),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_761),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_765),
.Y(n_807)
);

AOI21xp5_ASAP7_75t_L g808 ( 
.A1(n_737),
.A2(n_624),
.B(n_413),
.Y(n_808)
);

AOI22xp5_ASAP7_75t_L g809 ( 
.A1(n_749),
.A2(n_447),
.B1(n_443),
.B2(n_396),
.Y(n_809)
);

INVx5_ASAP7_75t_L g810 ( 
.A(n_751),
.Y(n_810)
);

OR2x6_ASAP7_75t_L g811 ( 
.A(n_694),
.B(n_689),
.Y(n_811)
);

INVx2_ASAP7_75t_L g812 ( 
.A(n_760),
.Y(n_812)
);

BUFx6f_ASAP7_75t_L g813 ( 
.A(n_711),
.Y(n_813)
);

OAI22xp5_ASAP7_75t_L g814 ( 
.A1(n_722),
.A2(n_423),
.B1(n_417),
.B2(n_418),
.Y(n_814)
);

INVx3_ASAP7_75t_L g815 ( 
.A(n_695),
.Y(n_815)
);

INVx3_ASAP7_75t_L g816 ( 
.A(n_711),
.Y(n_816)
);

AND2x4_ASAP7_75t_SL g817 ( 
.A(n_754),
.B(n_749),
.Y(n_817)
);

INVx2_ASAP7_75t_L g818 ( 
.A(n_764),
.Y(n_818)
);

INVx8_ASAP7_75t_L g819 ( 
.A(n_733),
.Y(n_819)
);

AOI22xp33_ASAP7_75t_L g820 ( 
.A1(n_739),
.A2(n_469),
.B1(n_421),
.B2(n_424),
.Y(n_820)
);

AOI22xp5_ASAP7_75t_L g821 ( 
.A1(n_710),
.A2(n_380),
.B1(n_384),
.B2(n_398),
.Y(n_821)
);

AOI22xp33_ASAP7_75t_L g822 ( 
.A1(n_714),
.A2(n_473),
.B1(n_425),
.B2(n_426),
.Y(n_822)
);

AOI22xp33_ASAP7_75t_L g823 ( 
.A1(n_740),
.A2(n_475),
.B1(n_428),
.B2(n_429),
.Y(n_823)
);

INVx3_ASAP7_75t_L g824 ( 
.A(n_747),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_L g825 ( 
.A(n_710),
.B(n_624),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_L g826 ( 
.A(n_752),
.B(n_624),
.Y(n_826)
);

NOR2xp33_ASAP7_75t_L g827 ( 
.A(n_707),
.B(n_762),
.Y(n_827)
);

INVx2_ASAP7_75t_SL g828 ( 
.A(n_716),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_L g829 ( 
.A(n_755),
.B(n_667),
.Y(n_829)
);

CKINVDCx20_ASAP7_75t_R g830 ( 
.A(n_772),
.Y(n_830)
);

INVx2_ASAP7_75t_L g831 ( 
.A(n_768),
.Y(n_831)
);

CKINVDCx8_ASAP7_75t_R g832 ( 
.A(n_767),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_743),
.Y(n_833)
);

OAI21x1_ASAP7_75t_SL g834 ( 
.A1(n_732),
.A2(n_435),
.B(n_434),
.Y(n_834)
);

AND2x2_ASAP7_75t_L g835 ( 
.A(n_747),
.B(n_675),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_745),
.Y(n_836)
);

INVx2_ASAP7_75t_L g837 ( 
.A(n_753),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_763),
.Y(n_838)
);

INVx1_ASAP7_75t_SL g839 ( 
.A(n_770),
.Y(n_839)
);

AOI21xp5_ASAP7_75t_L g840 ( 
.A1(n_718),
.A2(n_685),
.B(n_683),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_L g841 ( 
.A(n_838),
.B(n_742),
.Y(n_841)
);

BUFx12f_ASAP7_75t_L g842 ( 
.A(n_787),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_789),
.Y(n_843)
);

OAI22xp5_ASAP7_75t_L g844 ( 
.A1(n_827),
.A2(n_717),
.B1(n_756),
.B2(n_694),
.Y(n_844)
);

OAI22xp5_ASAP7_75t_L g845 ( 
.A1(n_799),
.A2(n_730),
.B1(n_766),
.B2(n_723),
.Y(n_845)
);

BUFx2_ASAP7_75t_L g846 ( 
.A(n_774),
.Y(n_846)
);

AND2x4_ASAP7_75t_L g847 ( 
.A(n_775),
.B(n_696),
.Y(n_847)
);

INVx1_ASAP7_75t_L g848 ( 
.A(n_801),
.Y(n_848)
);

OAI22xp5_ASAP7_75t_L g849 ( 
.A1(n_817),
.A2(n_730),
.B1(n_738),
.B2(n_727),
.Y(n_849)
);

INVx2_ASAP7_75t_L g850 ( 
.A(n_806),
.Y(n_850)
);

BUFx2_ASAP7_75t_L g851 ( 
.A(n_774),
.Y(n_851)
);

HB1xp67_ASAP7_75t_L g852 ( 
.A(n_796),
.Y(n_852)
);

OAI21x1_ASAP7_75t_L g853 ( 
.A1(n_788),
.A2(n_728),
.B(n_726),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_807),
.Y(n_854)
);

AOI22xp5_ASAP7_75t_L g855 ( 
.A1(n_814),
.A2(n_773),
.B1(n_488),
.B2(n_487),
.Y(n_855)
);

AND2x2_ASAP7_75t_L g856 ( 
.A(n_783),
.B(n_735),
.Y(n_856)
);

AND2x4_ASAP7_75t_SL g857 ( 
.A(n_813),
.B(n_731),
.Y(n_857)
);

BUFx3_ASAP7_75t_L g858 ( 
.A(n_813),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_833),
.Y(n_859)
);

INVx2_ASAP7_75t_L g860 ( 
.A(n_777),
.Y(n_860)
);

AND2x2_ASAP7_75t_L g861 ( 
.A(n_784),
.B(n_730),
.Y(n_861)
);

INVx2_ASAP7_75t_L g862 ( 
.A(n_797),
.Y(n_862)
);

OAI22xp5_ASAP7_75t_L g863 ( 
.A1(n_820),
.A2(n_485),
.B1(n_438),
.B2(n_451),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_L g864 ( 
.A(n_785),
.B(n_719),
.Y(n_864)
);

INVxp67_ASAP7_75t_L g865 ( 
.A(n_786),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_SL g866 ( 
.A(n_824),
.B(n_741),
.Y(n_866)
);

OAI221xp5_ASAP7_75t_L g867 ( 
.A1(n_793),
.A2(n_822),
.B1(n_809),
.B2(n_792),
.C(n_821),
.Y(n_867)
);

AND2x4_ASAP7_75t_L g868 ( 
.A(n_775),
.B(n_705),
.Y(n_868)
);

INVx2_ASAP7_75t_SL g869 ( 
.A(n_828),
.Y(n_869)
);

INVx2_ASAP7_75t_SL g870 ( 
.A(n_798),
.Y(n_870)
);

OAI22xp33_ASAP7_75t_L g871 ( 
.A1(n_829),
.A2(n_482),
.B1(n_439),
.B2(n_467),
.Y(n_871)
);

OR2x2_ASAP7_75t_L g872 ( 
.A(n_790),
.B(n_699),
.Y(n_872)
);

OAI22xp5_ASAP7_75t_L g873 ( 
.A1(n_804),
.A2(n_738),
.B1(n_441),
.B2(n_486),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_L g874 ( 
.A(n_794),
.B(n_442),
.Y(n_874)
);

AOI22xp33_ASAP7_75t_L g875 ( 
.A1(n_823),
.A2(n_490),
.B1(n_449),
.B2(n_460),
.Y(n_875)
);

OAI31xp33_ASAP7_75t_SL g876 ( 
.A1(n_836),
.A2(n_491),
.A3(n_455),
.B(n_456),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_835),
.Y(n_877)
);

CKINVDCx5p33_ASAP7_75t_R g878 ( 
.A(n_779),
.Y(n_878)
);

INVx2_ASAP7_75t_L g879 ( 
.A(n_812),
.Y(n_879)
);

AOI221xp5_ASAP7_75t_L g880 ( 
.A1(n_790),
.A2(n_561),
.B1(n_577),
.B2(n_585),
.C(n_470),
.Y(n_880)
);

AND2x2_ASAP7_75t_L g881 ( 
.A(n_839),
.B(n_700),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_818),
.Y(n_882)
);

OR2x2_ASAP7_75t_L g883 ( 
.A(n_803),
.B(n_709),
.Y(n_883)
);

AOI22xp33_ASAP7_75t_L g884 ( 
.A1(n_834),
.A2(n_493),
.B1(n_453),
.B2(n_471),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_831),
.Y(n_885)
);

AOI22xp5_ASAP7_75t_L g886 ( 
.A1(n_778),
.A2(n_462),
.B1(n_477),
.B2(n_474),
.Y(n_886)
);

HB1xp67_ASAP7_75t_L g887 ( 
.A(n_803),
.Y(n_887)
);

BUFx6f_ASAP7_75t_L g888 ( 
.A(n_798),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_837),
.Y(n_889)
);

HB1xp67_ASAP7_75t_L g890 ( 
.A(n_887),
.Y(n_890)
);

OAI211xp5_ASAP7_75t_L g891 ( 
.A1(n_876),
.A2(n_832),
.B(n_805),
.C(n_815),
.Y(n_891)
);

AOI22xp33_ASAP7_75t_L g892 ( 
.A1(n_867),
.A2(n_778),
.B1(n_834),
.B2(n_795),
.Y(n_892)
);

AOI21xp5_ASAP7_75t_L g893 ( 
.A1(n_874),
.A2(n_826),
.B(n_800),
.Y(n_893)
);

AOI22xp5_ASAP7_75t_L g894 ( 
.A1(n_844),
.A2(n_795),
.B1(n_776),
.B2(n_825),
.Y(n_894)
);

OAI22xp5_ASAP7_75t_SL g895 ( 
.A1(n_878),
.A2(n_830),
.B1(n_781),
.B2(n_811),
.Y(n_895)
);

AOI22xp33_ASAP7_75t_SL g896 ( 
.A1(n_844),
.A2(n_819),
.B1(n_791),
.B2(n_780),
.Y(n_896)
);

AND2x2_ASAP7_75t_L g897 ( 
.A(n_877),
.B(n_816),
.Y(n_897)
);

OAI221xp5_ASAP7_75t_SL g898 ( 
.A1(n_876),
.A2(n_811),
.B1(n_840),
.B2(n_819),
.C(n_808),
.Y(n_898)
);

AND2x2_ASAP7_75t_L g899 ( 
.A(n_856),
.B(n_802),
.Y(n_899)
);

AOI22xp33_ASAP7_75t_L g900 ( 
.A1(n_850),
.A2(n_480),
.B1(n_464),
.B2(n_461),
.Y(n_900)
);

AOI221xp5_ASAP7_75t_L g901 ( 
.A1(n_863),
.A2(n_802),
.B1(n_561),
.B2(n_577),
.C(n_459),
.Y(n_901)
);

AOI22xp33_ASAP7_75t_L g902 ( 
.A1(n_843),
.A2(n_713),
.B1(n_408),
.B2(n_415),
.Y(n_902)
);

AND2x2_ASAP7_75t_L g903 ( 
.A(n_881),
.B(n_782),
.Y(n_903)
);

INVxp67_ASAP7_75t_L g904 ( 
.A(n_852),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_848),
.Y(n_905)
);

AOI221xp5_ASAP7_75t_L g906 ( 
.A1(n_863),
.A2(n_865),
.B1(n_854),
.B2(n_886),
.C(n_871),
.Y(n_906)
);

AOI22xp33_ASAP7_75t_L g907 ( 
.A1(n_841),
.A2(n_406),
.B1(n_506),
.B2(n_505),
.Y(n_907)
);

OAI22xp5_ASAP7_75t_L g908 ( 
.A1(n_864),
.A2(n_859),
.B1(n_849),
.B2(n_846),
.Y(n_908)
);

AOI22xp33_ASAP7_75t_SL g909 ( 
.A1(n_851),
.A2(n_810),
.B1(n_500),
.B2(n_498),
.Y(n_909)
);

OAI22xp5_ASAP7_75t_L g910 ( 
.A1(n_882),
.A2(n_810),
.B1(n_496),
.B2(n_616),
.Y(n_910)
);

AOI22xp33_ASAP7_75t_L g911 ( 
.A1(n_879),
.A2(n_810),
.B1(n_759),
.B2(n_751),
.Y(n_911)
);

AOI22xp33_ASAP7_75t_L g912 ( 
.A1(n_885),
.A2(n_759),
.B1(n_605),
.B2(n_42),
.Y(n_912)
);

OAI21xp33_ASAP7_75t_L g913 ( 
.A1(n_886),
.A2(n_40),
.B(n_41),
.Y(n_913)
);

AOI22xp33_ASAP7_75t_L g914 ( 
.A1(n_889),
.A2(n_860),
.B1(n_862),
.B2(n_855),
.Y(n_914)
);

AOI22xp33_ASAP7_75t_L g915 ( 
.A1(n_855),
.A2(n_44),
.B1(n_46),
.B2(n_47),
.Y(n_915)
);

AOI21xp33_ASAP7_75t_L g916 ( 
.A1(n_872),
.A2(n_51),
.B(n_53),
.Y(n_916)
);

AOI22xp33_ASAP7_75t_L g917 ( 
.A1(n_875),
.A2(n_54),
.B1(n_56),
.B2(n_57),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_L g918 ( 
.A(n_868),
.B(n_58),
.Y(n_918)
);

INVx2_ASAP7_75t_L g919 ( 
.A(n_853),
.Y(n_919)
);

NOR2xp33_ASAP7_75t_L g920 ( 
.A(n_883),
.B(n_59),
.Y(n_920)
);

AND2x2_ASAP7_75t_L g921 ( 
.A(n_861),
.B(n_62),
.Y(n_921)
);

OAI22xp5_ASAP7_75t_L g922 ( 
.A1(n_845),
.A2(n_71),
.B1(n_75),
.B2(n_78),
.Y(n_922)
);

NAND2x1_ASAP7_75t_L g923 ( 
.A(n_888),
.B(n_80),
.Y(n_923)
);

OAI221xp5_ASAP7_75t_L g924 ( 
.A1(n_869),
.A2(n_884),
.B1(n_880),
.B2(n_866),
.C(n_858),
.Y(n_924)
);

OAI21xp33_ASAP7_75t_L g925 ( 
.A1(n_847),
.A2(n_81),
.B(n_84),
.Y(n_925)
);

AOI21xp33_ASAP7_75t_L g926 ( 
.A1(n_847),
.A2(n_85),
.B(n_91),
.Y(n_926)
);

AND2x2_ASAP7_75t_L g927 ( 
.A(n_868),
.B(n_93),
.Y(n_927)
);

AOI22xp33_ASAP7_75t_SL g928 ( 
.A1(n_891),
.A2(n_888),
.B1(n_845),
.B2(n_842),
.Y(n_928)
);

AOI221xp5_ASAP7_75t_L g929 ( 
.A1(n_906),
.A2(n_873),
.B1(n_870),
.B2(n_888),
.C(n_857),
.Y(n_929)
);

AOI22xp5_ASAP7_75t_L g930 ( 
.A1(n_920),
.A2(n_94),
.B1(n_96),
.B2(n_98),
.Y(n_930)
);

INVx2_ASAP7_75t_L g931 ( 
.A(n_905),
.Y(n_931)
);

AND2x2_ASAP7_75t_L g932 ( 
.A(n_899),
.B(n_99),
.Y(n_932)
);

OAI221xp5_ASAP7_75t_SL g933 ( 
.A1(n_913),
.A2(n_102),
.B1(n_112),
.B2(n_114),
.C(n_115),
.Y(n_933)
);

NAND3xp33_ASAP7_75t_L g934 ( 
.A(n_894),
.B(n_117),
.C(n_118),
.Y(n_934)
);

OAI21xp5_ASAP7_75t_L g935 ( 
.A1(n_903),
.A2(n_120),
.B(n_121),
.Y(n_935)
);

A2O1A1Ixp33_ASAP7_75t_L g936 ( 
.A1(n_892),
.A2(n_124),
.B(n_128),
.C(n_130),
.Y(n_936)
);

OAI21xp5_ASAP7_75t_SL g937 ( 
.A1(n_915),
.A2(n_141),
.B(n_149),
.Y(n_937)
);

INVxp67_ASAP7_75t_L g938 ( 
.A(n_890),
.Y(n_938)
);

AOI22xp33_ASAP7_75t_SL g939 ( 
.A1(n_922),
.A2(n_152),
.B1(n_159),
.B2(n_162),
.Y(n_939)
);

OAI211xp5_ASAP7_75t_L g940 ( 
.A1(n_896),
.A2(n_904),
.B(n_925),
.C(n_890),
.Y(n_940)
);

AND2x4_ASAP7_75t_SL g941 ( 
.A(n_927),
.B(n_164),
.Y(n_941)
);

INVx2_ASAP7_75t_L g942 ( 
.A(n_897),
.Y(n_942)
);

AOI21x1_ASAP7_75t_L g943 ( 
.A1(n_893),
.A2(n_296),
.B(n_166),
.Y(n_943)
);

NAND3xp33_ASAP7_75t_L g944 ( 
.A(n_898),
.B(n_165),
.C(n_169),
.Y(n_944)
);

INVx2_ASAP7_75t_L g945 ( 
.A(n_919),
.Y(n_945)
);

NAND2xp5_ASAP7_75t_L g946 ( 
.A(n_908),
.B(n_170),
.Y(n_946)
);

HB1xp67_ASAP7_75t_L g947 ( 
.A(n_904),
.Y(n_947)
);

OAI33xp33_ASAP7_75t_L g948 ( 
.A1(n_910),
.A2(n_171),
.A3(n_172),
.B1(n_177),
.B2(n_180),
.B3(n_181),
.Y(n_948)
);

AOI22xp33_ASAP7_75t_L g949 ( 
.A1(n_924),
.A2(n_183),
.B1(n_186),
.B2(n_187),
.Y(n_949)
);

OR2x2_ASAP7_75t_L g950 ( 
.A(n_921),
.B(n_190),
.Y(n_950)
);

INVx2_ASAP7_75t_L g951 ( 
.A(n_918),
.Y(n_951)
);

INVx1_ASAP7_75t_L g952 ( 
.A(n_914),
.Y(n_952)
);

HB1xp67_ASAP7_75t_L g953 ( 
.A(n_895),
.Y(n_953)
);

AND2x2_ASAP7_75t_L g954 ( 
.A(n_896),
.B(n_191),
.Y(n_954)
);

AND2x2_ASAP7_75t_L g955 ( 
.A(n_909),
.B(n_193),
.Y(n_955)
);

OAI21x1_ASAP7_75t_L g956 ( 
.A1(n_923),
.A2(n_195),
.B(n_197),
.Y(n_956)
);

HB1xp67_ASAP7_75t_L g957 ( 
.A(n_911),
.Y(n_957)
);

OR2x2_ASAP7_75t_L g958 ( 
.A(n_947),
.B(n_938),
.Y(n_958)
);

OAI31xp33_ASAP7_75t_L g959 ( 
.A1(n_933),
.A2(n_916),
.A3(n_926),
.B(n_917),
.Y(n_959)
);

NAND4xp25_ASAP7_75t_L g960 ( 
.A(n_938),
.B(n_901),
.C(n_902),
.D(n_909),
.Y(n_960)
);

AO31x2_ASAP7_75t_L g961 ( 
.A1(n_945),
.A2(n_907),
.A3(n_900),
.B(n_912),
.Y(n_961)
);

AO21x2_ASAP7_75t_L g962 ( 
.A1(n_944),
.A2(n_200),
.B(n_201),
.Y(n_962)
);

OAI21xp5_ASAP7_75t_L g963 ( 
.A1(n_934),
.A2(n_205),
.B(n_206),
.Y(n_963)
);

NAND2xp5_ASAP7_75t_SL g964 ( 
.A(n_951),
.B(n_207),
.Y(n_964)
);

AND2x4_ASAP7_75t_L g965 ( 
.A(n_942),
.B(n_216),
.Y(n_965)
);

INVx2_ASAP7_75t_L g966 ( 
.A(n_931),
.Y(n_966)
);

AND2x2_ASAP7_75t_L g967 ( 
.A(n_932),
.B(n_223),
.Y(n_967)
);

INVx1_ASAP7_75t_L g968 ( 
.A(n_952),
.Y(n_968)
);

AOI22xp5_ASAP7_75t_L g969 ( 
.A1(n_940),
.A2(n_224),
.B1(n_226),
.B2(n_227),
.Y(n_969)
);

OR2x2_ASAP7_75t_L g970 ( 
.A(n_947),
.B(n_950),
.Y(n_970)
);

INVx2_ASAP7_75t_L g971 ( 
.A(n_956),
.Y(n_971)
);

INVx3_ASAP7_75t_L g972 ( 
.A(n_941),
.Y(n_972)
);

OAI221xp5_ASAP7_75t_L g973 ( 
.A1(n_937),
.A2(n_235),
.B1(n_238),
.B2(n_239),
.C(n_240),
.Y(n_973)
);

OR2x2_ASAP7_75t_L g974 ( 
.A(n_957),
.B(n_241),
.Y(n_974)
);

OR2x2_ASAP7_75t_L g975 ( 
.A(n_957),
.B(n_242),
.Y(n_975)
);

OAI31xp33_ASAP7_75t_SL g976 ( 
.A1(n_954),
.A2(n_252),
.A3(n_253),
.B(n_255),
.Y(n_976)
);

INVx3_ASAP7_75t_L g977 ( 
.A(n_943),
.Y(n_977)
);

INVx2_ASAP7_75t_L g978 ( 
.A(n_946),
.Y(n_978)
);

AND2x2_ASAP7_75t_L g979 ( 
.A(n_970),
.B(n_928),
.Y(n_979)
);

OR2x2_ASAP7_75t_L g980 ( 
.A(n_958),
.B(n_953),
.Y(n_980)
);

AND2x2_ASAP7_75t_L g981 ( 
.A(n_968),
.B(n_955),
.Y(n_981)
);

BUFx2_ASAP7_75t_L g982 ( 
.A(n_966),
.Y(n_982)
);

BUFx3_ASAP7_75t_L g983 ( 
.A(n_972),
.Y(n_983)
);

OR2x2_ASAP7_75t_L g984 ( 
.A(n_968),
.B(n_935),
.Y(n_984)
);

NAND2xp5_ASAP7_75t_L g985 ( 
.A(n_978),
.B(n_928),
.Y(n_985)
);

AND2x2_ASAP7_75t_L g986 ( 
.A(n_974),
.B(n_939),
.Y(n_986)
);

INVx2_ASAP7_75t_L g987 ( 
.A(n_971),
.Y(n_987)
);

INVx1_ASAP7_75t_L g988 ( 
.A(n_975),
.Y(n_988)
);

INVx1_ASAP7_75t_L g989 ( 
.A(n_977),
.Y(n_989)
);

AND2x2_ASAP7_75t_L g990 ( 
.A(n_965),
.B(n_939),
.Y(n_990)
);

AND2x2_ASAP7_75t_L g991 ( 
.A(n_965),
.B(n_949),
.Y(n_991)
);

AND2x2_ASAP7_75t_L g992 ( 
.A(n_976),
.B(n_936),
.Y(n_992)
);

NAND2xp5_ASAP7_75t_L g993 ( 
.A(n_967),
.B(n_929),
.Y(n_993)
);

AND2x2_ASAP7_75t_L g994 ( 
.A(n_969),
.B(n_930),
.Y(n_994)
);

INVx1_ASAP7_75t_L g995 ( 
.A(n_977),
.Y(n_995)
);

NAND2xp5_ASAP7_75t_L g996 ( 
.A(n_972),
.B(n_256),
.Y(n_996)
);

INVx1_ASAP7_75t_L g997 ( 
.A(n_989),
.Y(n_997)
);

OR2x2_ASAP7_75t_L g998 ( 
.A(n_988),
.B(n_962),
.Y(n_998)
);

AND2x2_ASAP7_75t_L g999 ( 
.A(n_979),
.B(n_969),
.Y(n_999)
);

NAND2xp5_ASAP7_75t_L g1000 ( 
.A(n_982),
.B(n_959),
.Y(n_1000)
);

INVx1_ASAP7_75t_L g1001 ( 
.A(n_995),
.Y(n_1001)
);

BUFx2_ASAP7_75t_SL g1002 ( 
.A(n_983),
.Y(n_1002)
);

NAND2xp5_ASAP7_75t_L g1003 ( 
.A(n_981),
.B(n_964),
.Y(n_1003)
);

NAND2xp5_ASAP7_75t_L g1004 ( 
.A(n_981),
.B(n_962),
.Y(n_1004)
);

NOR2xp33_ASAP7_75t_L g1005 ( 
.A(n_980),
.B(n_960),
.Y(n_1005)
);

AND2x2_ASAP7_75t_L g1006 ( 
.A(n_990),
.B(n_963),
.Y(n_1006)
);

AND2x4_ASAP7_75t_L g1007 ( 
.A(n_983),
.B(n_961),
.Y(n_1007)
);

INVx1_ASAP7_75t_SL g1008 ( 
.A(n_985),
.Y(n_1008)
);

INVx1_ASAP7_75t_L g1009 ( 
.A(n_997),
.Y(n_1009)
);

INVx1_ASAP7_75t_L g1010 ( 
.A(n_1001),
.Y(n_1010)
);

XNOR2x2_ASAP7_75t_L g1011 ( 
.A(n_1008),
.B(n_986),
.Y(n_1011)
);

INVx1_ASAP7_75t_L g1012 ( 
.A(n_998),
.Y(n_1012)
);

OR2x2_ASAP7_75t_L g1013 ( 
.A(n_1004),
.B(n_987),
.Y(n_1013)
);

INVx1_ASAP7_75t_L g1014 ( 
.A(n_1007),
.Y(n_1014)
);

AND2x2_ASAP7_75t_L g1015 ( 
.A(n_1008),
.B(n_986),
.Y(n_1015)
);

OAI21xp5_ASAP7_75t_SL g1016 ( 
.A1(n_1015),
.A2(n_1006),
.B(n_999),
.Y(n_1016)
);

XNOR2xp5_ASAP7_75t_L g1017 ( 
.A(n_1011),
.B(n_1000),
.Y(n_1017)
);

INVx1_ASAP7_75t_L g1018 ( 
.A(n_1009),
.Y(n_1018)
);

OR2x2_ASAP7_75t_L g1019 ( 
.A(n_1012),
.B(n_1003),
.Y(n_1019)
);

AOI211xp5_ASAP7_75t_L g1020 ( 
.A1(n_1011),
.A2(n_1005),
.B(n_994),
.C(n_992),
.Y(n_1020)
);

AND2x2_ASAP7_75t_L g1021 ( 
.A(n_1016),
.B(n_1014),
.Y(n_1021)
);

AOI21xp5_ASAP7_75t_L g1022 ( 
.A1(n_1020),
.A2(n_994),
.B(n_992),
.Y(n_1022)
);

INVx2_ASAP7_75t_L g1023 ( 
.A(n_1018),
.Y(n_1023)
);

CKINVDCx20_ASAP7_75t_R g1024 ( 
.A(n_1017),
.Y(n_1024)
);

OAI221xp5_ASAP7_75t_SL g1025 ( 
.A1(n_1022),
.A2(n_993),
.B1(n_973),
.B2(n_1019),
.C(n_984),
.Y(n_1025)
);

AOI322xp5_ASAP7_75t_L g1026 ( 
.A1(n_1024),
.A2(n_991),
.A3(n_1010),
.B1(n_1007),
.B2(n_996),
.C1(n_933),
.C2(n_987),
.Y(n_1026)
);

AND2x2_ASAP7_75t_L g1027 ( 
.A(n_1021),
.B(n_1002),
.Y(n_1027)
);

NOR2x1_ASAP7_75t_L g1028 ( 
.A(n_1023),
.B(n_1013),
.Y(n_1028)
);

OAI211xp5_ASAP7_75t_L g1029 ( 
.A1(n_1024),
.A2(n_991),
.B(n_948),
.C(n_262),
.Y(n_1029)
);

NAND3xp33_ASAP7_75t_L g1030 ( 
.A(n_1026),
.B(n_948),
.C(n_261),
.Y(n_1030)
);

AOI221x1_ASAP7_75t_L g1031 ( 
.A1(n_1027),
.A2(n_961),
.B1(n_263),
.B2(n_265),
.C(n_266),
.Y(n_1031)
);

XNOR2xp5_ASAP7_75t_L g1032 ( 
.A(n_1030),
.B(n_1029),
.Y(n_1032)
);

OAI221xp5_ASAP7_75t_L g1033 ( 
.A1(n_1032),
.A2(n_1025),
.B1(n_1028),
.B2(n_1031),
.C(n_283),
.Y(n_1033)
);

AND3x4_ASAP7_75t_L g1034 ( 
.A(n_1033),
.B(n_257),
.C(n_274),
.Y(n_1034)
);

INVx1_ASAP7_75t_L g1035 ( 
.A(n_1034),
.Y(n_1035)
);

AOI22xp33_ASAP7_75t_L g1036 ( 
.A1(n_1035),
.A2(n_282),
.B1(n_287),
.B2(n_292),
.Y(n_1036)
);

AOI21xp5_ASAP7_75t_L g1037 ( 
.A1(n_1036),
.A2(n_294),
.B(n_295),
.Y(n_1037)
);


endmodule