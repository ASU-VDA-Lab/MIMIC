module fake_jpeg_2199_n_653 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_653);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_653;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_182;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_620;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_417;
wire n_362;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_635;
wire n_517;
wire n_629;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_643;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_647;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_641;
wire n_48;
wire n_465;
wire n_638;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_623;
wire n_579;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_637;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_624;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_646;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_393;
wire n_349;
wire n_234;
wire n_530;
wire n_634;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_639;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_645;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_622;
wire n_463;
wire n_92;
wire n_332;
wire n_640;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_626;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_511;
wire n_486;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_642;
wire n_101;
wire n_226;
wire n_509;
wire n_644;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_649;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_615;
wire n_598;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_648;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_631;
wire n_433;
wire n_636;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_650;
wire n_218;
wire n_63;
wire n_652;
wire n_599;
wire n_239;
wire n_243;
wire n_481;
wire n_628;
wire n_619;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_260;
wire n_199;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_625;
wire n_147;
wire n_449;
wire n_627;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_613;
wire n_630;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_633;
wire n_112;
wire n_632;
wire n_616;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_651;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_621;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

CKINVDCx14_ASAP7_75t_R g21 ( 
.A(n_11),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

INVx8_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_11),
.Y(n_25)
);

INVx8_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

INVx13_ASAP7_75t_L g27 ( 
.A(n_18),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_19),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_4),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_6),
.Y(n_31)
);

BUFx12_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_10),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_18),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_10),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_10),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_1),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_9),
.Y(n_38)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_17),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_7),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_0),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_11),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_9),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_12),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_16),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_1),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_9),
.Y(n_47)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_18),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_2),
.Y(n_49)
);

BUFx5_ASAP7_75t_L g50 ( 
.A(n_8),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_7),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_11),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_16),
.Y(n_53)
);

INVxp33_ASAP7_75t_L g54 ( 
.A(n_19),
.Y(n_54)
);

INVx8_ASAP7_75t_L g55 ( 
.A(n_16),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_14),
.Y(n_56)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_14),
.Y(n_57)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_38),
.Y(n_58)
);

BUFx2_ASAP7_75t_L g155 ( 
.A(n_58),
.Y(n_155)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_37),
.Y(n_59)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_59),
.Y(n_131)
);

CKINVDCx9p33_ASAP7_75t_R g60 ( 
.A(n_21),
.Y(n_60)
);

INVx8_ASAP7_75t_L g172 ( 
.A(n_60),
.Y(n_172)
);

INVx11_ASAP7_75t_L g61 ( 
.A(n_38),
.Y(n_61)
);

INVx4_ASAP7_75t_L g133 ( 
.A(n_61),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_22),
.B(n_9),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_62),
.B(n_90),
.Y(n_145)
);

AND2x4_ASAP7_75t_SL g63 ( 
.A(n_37),
.B(n_41),
.Y(n_63)
);

NAND2xp33_ASAP7_75t_SL g222 ( 
.A(n_63),
.B(n_83),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_35),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_64),
.B(n_80),
.Y(n_148)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_33),
.Y(n_65)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_65),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_35),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_66),
.Y(n_134)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_33),
.Y(n_67)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_67),
.Y(n_165)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_22),
.Y(n_68)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_68),
.Y(n_138)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_36),
.Y(n_69)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_69),
.Y(n_171)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_39),
.Y(n_70)
);

INVx3_ASAP7_75t_L g132 ( 
.A(n_70),
.Y(n_132)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_36),
.Y(n_71)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_71),
.Y(n_176)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_48),
.Y(n_72)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_72),
.Y(n_177)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_35),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g142 ( 
.A(n_73),
.Y(n_142)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_48),
.Y(n_74)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_74),
.Y(n_179)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_39),
.Y(n_75)
);

INVx3_ASAP7_75t_L g136 ( 
.A(n_75),
.Y(n_136)
);

INVx8_ASAP7_75t_L g76 ( 
.A(n_38),
.Y(n_76)
);

BUFx2_ASAP7_75t_L g180 ( 
.A(n_76),
.Y(n_180)
);

BUFx5_ASAP7_75t_L g77 ( 
.A(n_50),
.Y(n_77)
);

INVx4_ASAP7_75t_L g144 ( 
.A(n_77),
.Y(n_144)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_28),
.Y(n_78)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_78),
.Y(n_169)
);

BUFx5_ASAP7_75t_L g79 ( 
.A(n_50),
.Y(n_79)
);

INVx4_ASAP7_75t_L g168 ( 
.A(n_79),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_35),
.Y(n_80)
);

BUFx3_ASAP7_75t_L g81 ( 
.A(n_24),
.Y(n_81)
);

BUFx3_ASAP7_75t_L g140 ( 
.A(n_81),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_34),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_82),
.B(n_96),
.Y(n_149)
);

OR2x2_ASAP7_75t_L g83 ( 
.A(n_54),
.B(n_10),
.Y(n_83)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_48),
.Y(n_84)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_84),
.Y(n_185)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_28),
.Y(n_85)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_85),
.Y(n_189)
);

BUFx12f_ASAP7_75t_L g86 ( 
.A(n_32),
.Y(n_86)
);

INVx5_ASAP7_75t_L g152 ( 
.A(n_86),
.Y(n_152)
);

INVx8_ASAP7_75t_L g87 ( 
.A(n_38),
.Y(n_87)
);

INVx5_ASAP7_75t_L g159 ( 
.A(n_87),
.Y(n_159)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_39),
.Y(n_88)
);

INVx3_ASAP7_75t_L g206 ( 
.A(n_88),
.Y(n_206)
);

INVx8_ASAP7_75t_L g89 ( 
.A(n_38),
.Y(n_89)
);

INVx5_ASAP7_75t_L g161 ( 
.A(n_89),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_31),
.B(n_8),
.Y(n_90)
);

INVx13_ASAP7_75t_L g91 ( 
.A(n_27),
.Y(n_91)
);

INVx13_ASAP7_75t_L g224 ( 
.A(n_91),
.Y(n_224)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_31),
.Y(n_92)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_92),
.Y(n_209)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_34),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g143 ( 
.A(n_93),
.Y(n_143)
);

BUFx12f_ASAP7_75t_L g94 ( 
.A(n_32),
.Y(n_94)
);

INVx5_ASAP7_75t_L g182 ( 
.A(n_94),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_54),
.B(n_19),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_95),
.B(n_125),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_34),
.Y(n_96)
);

INVx4_ASAP7_75t_L g97 ( 
.A(n_41),
.Y(n_97)
);

INVx4_ASAP7_75t_L g170 ( 
.A(n_97),
.Y(n_170)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_41),
.Y(n_98)
);

INVx4_ASAP7_75t_L g178 ( 
.A(n_98),
.Y(n_178)
);

INVx8_ASAP7_75t_L g99 ( 
.A(n_52),
.Y(n_99)
);

INVx5_ASAP7_75t_L g188 ( 
.A(n_99),
.Y(n_188)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_52),
.Y(n_100)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_100),
.Y(n_191)
);

BUFx12f_ASAP7_75t_L g101 ( 
.A(n_32),
.Y(n_101)
);

INVx5_ASAP7_75t_L g205 ( 
.A(n_101),
.Y(n_205)
);

BUFx3_ASAP7_75t_L g102 ( 
.A(n_24),
.Y(n_102)
);

BUFx3_ASAP7_75t_L g160 ( 
.A(n_102),
.Y(n_160)
);

INVx6_ASAP7_75t_L g103 ( 
.A(n_45),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g147 ( 
.A(n_103),
.Y(n_147)
);

INVx8_ASAP7_75t_L g104 ( 
.A(n_52),
.Y(n_104)
);

BUFx3_ASAP7_75t_L g181 ( 
.A(n_104),
.Y(n_181)
);

BUFx12f_ASAP7_75t_L g105 ( 
.A(n_32),
.Y(n_105)
);

INVx8_ASAP7_75t_L g194 ( 
.A(n_105),
.Y(n_194)
);

INVx13_ASAP7_75t_L g106 ( 
.A(n_27),
.Y(n_106)
);

BUFx3_ASAP7_75t_L g213 ( 
.A(n_106),
.Y(n_213)
);

INVx11_ASAP7_75t_L g107 ( 
.A(n_52),
.Y(n_107)
);

INVx4_ASAP7_75t_L g183 ( 
.A(n_107),
.Y(n_183)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_45),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g154 ( 
.A(n_108),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_SL g109 ( 
.A(n_25),
.B(n_8),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_109),
.B(n_130),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_45),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g164 ( 
.A(n_110),
.Y(n_164)
);

BUFx3_ASAP7_75t_L g111 ( 
.A(n_24),
.Y(n_111)
);

INVx4_ASAP7_75t_L g195 ( 
.A(n_111),
.Y(n_195)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_20),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g197 ( 
.A(n_112),
.Y(n_197)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_20),
.Y(n_113)
);

INVx6_ASAP7_75t_L g166 ( 
.A(n_113),
.Y(n_166)
);

INVx8_ASAP7_75t_L g114 ( 
.A(n_52),
.Y(n_114)
);

INVx4_ASAP7_75t_L g198 ( 
.A(n_114),
.Y(n_198)
);

INVx8_ASAP7_75t_L g115 ( 
.A(n_57),
.Y(n_115)
);

INVx4_ASAP7_75t_L g203 ( 
.A(n_115),
.Y(n_203)
);

INVx8_ASAP7_75t_L g116 ( 
.A(n_57),
.Y(n_116)
);

INVx4_ASAP7_75t_L g214 ( 
.A(n_116),
.Y(n_214)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_40),
.Y(n_117)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_117),
.Y(n_219)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_20),
.Y(n_118)
);

INVx6_ASAP7_75t_L g200 ( 
.A(n_118),
.Y(n_200)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_57),
.Y(n_119)
);

INVx4_ASAP7_75t_L g217 ( 
.A(n_119),
.Y(n_217)
);

INVx6_ASAP7_75t_L g120 ( 
.A(n_23),
.Y(n_120)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_120),
.Y(n_196)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_57),
.Y(n_121)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_121),
.Y(n_199)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_57),
.Y(n_122)
);

INVx6_ASAP7_75t_L g218 ( 
.A(n_122),
.Y(n_218)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_23),
.Y(n_123)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_123),
.Y(n_221)
);

INVx11_ASAP7_75t_L g124 ( 
.A(n_27),
.Y(n_124)
);

INVx6_ASAP7_75t_L g220 ( 
.A(n_124),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_40),
.B(n_12),
.Y(n_125)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_49),
.Y(n_126)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_126),
.Y(n_223)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_32),
.Y(n_127)
);

INVx6_ASAP7_75t_L g228 ( 
.A(n_127),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_46),
.B(n_12),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_128),
.B(n_15),
.Y(n_162)
);

BUFx5_ASAP7_75t_L g129 ( 
.A(n_50),
.Y(n_129)
);

AOI21xp33_ASAP7_75t_L g229 ( 
.A1(n_129),
.A2(n_4),
.B(n_5),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_21),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_83),
.B(n_53),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_SL g255 ( 
.A(n_135),
.B(n_139),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_103),
.A2(n_44),
.B1(n_25),
.B2(n_29),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g253 ( 
.A1(n_137),
.A2(n_150),
.B1(n_156),
.B2(n_175),
.Y(n_253)
);

AND2x2_ASAP7_75t_L g139 ( 
.A(n_119),
.B(n_56),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_84),
.B(n_56),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_SL g247 ( 
.A(n_141),
.B(n_158),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_60),
.A2(n_44),
.B1(n_42),
.B2(n_51),
.Y(n_146)
);

OAI22xp33_ASAP7_75t_SL g282 ( 
.A1(n_146),
.A2(n_127),
.B1(n_87),
.B2(n_89),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_63),
.A2(n_49),
.B1(n_53),
.B2(n_51),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_63),
.A2(n_42),
.B1(n_47),
.B2(n_29),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_86),
.B(n_47),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g233 ( 
.A(n_162),
.B(n_167),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_86),
.B(n_43),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_163),
.B(n_173),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_70),
.B(n_46),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_94),
.B(n_43),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_88),
.B(n_30),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_174),
.B(n_208),
.Y(n_236)
);

AOI22xp33_ASAP7_75t_SL g175 ( 
.A1(n_123),
.A2(n_55),
.B1(n_26),
.B2(n_23),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_94),
.B(n_30),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_184),
.B(n_187),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_98),
.B(n_55),
.C(n_26),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g308 ( 
.A(n_186),
.B(n_175),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_101),
.B(n_55),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_101),
.B(n_26),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_190),
.B(n_193),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_93),
.A2(n_12),
.B1(n_18),
.B2(n_2),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_192),
.A2(n_204),
.B1(n_115),
.B2(n_15),
.Y(n_298)
);

AND2x2_ASAP7_75t_L g193 ( 
.A(n_97),
.B(n_7),
.Y(n_193)
);

OA22x2_ASAP7_75t_L g201 ( 
.A1(n_120),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_201)
);

AOI22x1_ASAP7_75t_L g313 ( 
.A1(n_201),
.A2(n_216),
.B1(n_215),
.B2(n_210),
.Y(n_313)
);

AND2x2_ASAP7_75t_L g202 ( 
.A(n_75),
.B(n_6),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_202),
.B(n_207),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_L g204 ( 
.A1(n_108),
.A2(n_6),
.B1(n_17),
.B2(n_2),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_105),
.B(n_19),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_112),
.B(n_13),
.Y(n_208)
);

AOI22xp33_ASAP7_75t_SL g210 ( 
.A1(n_61),
.A2(n_13),
.B1(n_16),
.B2(n_3),
.Y(n_210)
);

AOI22xp33_ASAP7_75t_SL g234 ( 
.A1(n_210),
.A2(n_215),
.B1(n_225),
.B2(n_111),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_105),
.B(n_17),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_211),
.B(n_212),
.Y(n_266)
);

AND2x2_ASAP7_75t_L g212 ( 
.A(n_58),
.B(n_5),
.Y(n_212)
);

AOI22xp33_ASAP7_75t_SL g215 ( 
.A1(n_107),
.A2(n_5),
.B1(n_15),
.B2(n_3),
.Y(n_215)
);

OAI22xp33_ASAP7_75t_SL g216 ( 
.A1(n_113),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_216)
);

AOI22xp33_ASAP7_75t_SL g225 ( 
.A1(n_81),
.A2(n_13),
.B1(n_3),
.B2(n_4),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_73),
.Y(n_226)
);

INVx1_ASAP7_75t_SL g249 ( 
.A(n_226),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_118),
.B(n_4),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_SL g251 ( 
.A(n_227),
.B(n_66),
.Y(n_251)
);

OR2x4_ASAP7_75t_L g309 ( 
.A(n_229),
.B(n_225),
.Y(n_309)
);

CKINVDCx16_ASAP7_75t_R g230 ( 
.A(n_155),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_SL g347 ( 
.A(n_230),
.B(n_232),
.Y(n_347)
);

INVx3_ASAP7_75t_L g231 ( 
.A(n_213),
.Y(n_231)
);

BUFx2_ASAP7_75t_L g358 ( 
.A(n_231),
.Y(n_358)
);

A2O1A1Ixp33_ASAP7_75t_L g232 ( 
.A1(n_222),
.A2(n_91),
.B(n_106),
.C(n_124),
.Y(n_232)
);

INVxp67_ASAP7_75t_L g329 ( 
.A(n_234),
.Y(n_329)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_148),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_SL g359 ( 
.A(n_235),
.B(n_252),
.Y(n_359)
);

INVx13_ASAP7_75t_L g237 ( 
.A(n_224),
.Y(n_237)
);

INVx1_ASAP7_75t_SL g339 ( 
.A(n_237),
.Y(n_339)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_223),
.Y(n_238)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_238),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_145),
.B(n_0),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_241),
.B(n_279),
.Y(n_321)
);

INVx3_ASAP7_75t_SL g242 ( 
.A(n_172),
.Y(n_242)
);

INVx2_ASAP7_75t_L g327 ( 
.A(n_242),
.Y(n_327)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_196),
.Y(n_243)
);

INVx2_ASAP7_75t_L g342 ( 
.A(n_243),
.Y(n_342)
);

INVx3_ASAP7_75t_L g244 ( 
.A(n_213),
.Y(n_244)
);

INVx3_ASAP7_75t_L g351 ( 
.A(n_244),
.Y(n_351)
);

INVxp67_ASAP7_75t_L g246 ( 
.A(n_139),
.Y(n_246)
);

BUFx3_ASAP7_75t_L g330 ( 
.A(n_246),
.Y(n_330)
);

BUFx2_ASAP7_75t_L g248 ( 
.A(n_155),
.Y(n_248)
);

BUFx3_ASAP7_75t_L g344 ( 
.A(n_248),
.Y(n_344)
);

BUFx6f_ASAP7_75t_L g250 ( 
.A(n_143),
.Y(n_250)
);

BUFx6f_ASAP7_75t_L g371 ( 
.A(n_250),
.Y(n_371)
);

NAND3xp33_ASAP7_75t_L g362 ( 
.A(n_251),
.B(n_287),
.C(n_291),
.Y(n_362)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_149),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_157),
.B(n_153),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_SL g317 ( 
.A(n_254),
.B(n_267),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_180),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_SL g360 ( 
.A(n_256),
.B(n_261),
.Y(n_360)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_221),
.Y(n_257)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_257),
.Y(n_325)
);

BUFx6f_ASAP7_75t_L g258 ( 
.A(n_143),
.Y(n_258)
);

INVx5_ASAP7_75t_L g353 ( 
.A(n_258),
.Y(n_353)
);

AOI22xp33_ASAP7_75t_SL g259 ( 
.A1(n_172),
.A2(n_144),
.B1(n_168),
.B2(n_212),
.Y(n_259)
);

AOI22xp33_ASAP7_75t_SL g338 ( 
.A1(n_259),
.A2(n_260),
.B1(n_181),
.B2(n_161),
.Y(n_338)
);

O2A1O1Ixp33_ASAP7_75t_SL g260 ( 
.A1(n_201),
.A2(n_129),
.B(n_79),
.C(n_77),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_180),
.Y(n_261)
);

BUFx12f_ASAP7_75t_L g262 ( 
.A(n_194),
.Y(n_262)
);

INVx5_ASAP7_75t_L g366 ( 
.A(n_262),
.Y(n_366)
);

INVx13_ASAP7_75t_L g263 ( 
.A(n_224),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g345 ( 
.A(n_263),
.Y(n_345)
);

INVxp67_ASAP7_75t_L g264 ( 
.A(n_136),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_264),
.B(n_281),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_SL g267 ( 
.A(n_138),
.B(n_102),
.Y(n_267)
);

INVx6_ASAP7_75t_L g268 ( 
.A(n_154),
.Y(n_268)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_268),
.Y(n_336)
);

INVx5_ASAP7_75t_L g269 ( 
.A(n_194),
.Y(n_269)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_269),
.Y(n_367)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_185),
.Y(n_270)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_270),
.Y(n_369)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_178),
.Y(n_271)
);

AND2x2_ASAP7_75t_L g322 ( 
.A(n_271),
.B(n_273),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_169),
.B(n_189),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_SL g365 ( 
.A(n_272),
.B(n_275),
.Y(n_365)
);

INVx2_ASAP7_75t_SL g273 ( 
.A(n_170),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_209),
.Y(n_274)
);

AND2x2_ASAP7_75t_L g323 ( 
.A(n_274),
.B(n_276),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_219),
.B(n_99),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_217),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_218),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_SL g368 ( 
.A(n_277),
.B(n_278),
.Y(n_368)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_151),
.B(n_104),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_193),
.B(n_110),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_202),
.B(n_122),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_280),
.B(n_288),
.Y(n_332)
);

BUFx3_ASAP7_75t_L g281 ( 
.A(n_152),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_SL g373 ( 
.A1(n_282),
.A2(n_164),
.B1(n_242),
.B2(n_260),
.Y(n_373)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_217),
.Y(n_283)
);

AND2x2_ASAP7_75t_L g349 ( 
.A(n_283),
.B(n_285),
.Y(n_349)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_165),
.B(n_76),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_284),
.B(n_289),
.Y(n_328)
);

INVx3_ASAP7_75t_L g285 ( 
.A(n_198),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_178),
.Y(n_286)
);

OR2x2_ASAP7_75t_L g331 ( 
.A(n_286),
.B(n_290),
.Y(n_331)
);

BUFx4f_ASAP7_75t_SL g287 ( 
.A(n_132),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_131),
.B(n_13),
.Y(n_288)
);

CKINVDCx16_ASAP7_75t_R g289 ( 
.A(n_133),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_170),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_218),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g292 ( 
.A(n_159),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_292),
.B(n_293),
.Y(n_333)
);

INVxp33_ASAP7_75t_L g293 ( 
.A(n_216),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_171),
.B(n_14),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_294),
.B(n_297),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_176),
.B(n_116),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_295),
.B(n_296),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_177),
.B(n_114),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_201),
.B(n_15),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_L g363 ( 
.A1(n_298),
.A2(n_313),
.B1(n_297),
.B2(n_308),
.Y(n_363)
);

INVxp67_ASAP7_75t_L g299 ( 
.A(n_206),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g352 ( 
.A(n_299),
.B(n_302),
.Y(n_352)
);

MAJx2_ASAP7_75t_L g300 ( 
.A(n_179),
.B(n_17),
.C(n_199),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_300),
.B(n_160),
.C(n_140),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_191),
.B(n_147),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_301),
.B(n_310),
.Y(n_337)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_147),
.Y(n_302)
);

BUFx3_ASAP7_75t_L g303 ( 
.A(n_182),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g355 ( 
.A(n_303),
.B(n_304),
.Y(n_355)
);

INVx2_ASAP7_75t_L g304 ( 
.A(n_195),
.Y(n_304)
);

INVx5_ASAP7_75t_L g305 ( 
.A(n_140),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g348 ( 
.A(n_305),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_195),
.B(n_160),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g370 ( 
.A(n_306),
.B(n_307),
.Y(n_370)
);

BUFx3_ASAP7_75t_L g307 ( 
.A(n_205),
.Y(n_307)
);

XNOR2x1_ASAP7_75t_L g375 ( 
.A(n_308),
.B(n_309),
.Y(n_375)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_198),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_203),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_311),
.B(n_312),
.Y(n_346)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_203),
.Y(n_312)
);

INVx3_ASAP7_75t_L g314 ( 
.A(n_214),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g374 ( 
.A(n_314),
.B(n_164),
.Y(n_374)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_214),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_315),
.B(n_228),
.Y(n_356)
);

AOI21xp5_ASAP7_75t_L g318 ( 
.A1(n_232),
.A2(n_168),
.B(n_144),
.Y(n_318)
);

OAI21xp5_ASAP7_75t_SL g390 ( 
.A1(n_318),
.A2(n_343),
.B(n_329),
.Y(n_390)
);

XNOR2xp5_ASAP7_75t_L g378 ( 
.A(n_320),
.B(n_280),
.Y(n_378)
);

XNOR2xp5_ASAP7_75t_L g324 ( 
.A(n_233),
.B(n_300),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g380 ( 
.A(n_324),
.B(n_326),
.C(n_265),
.Y(n_380)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_246),
.B(n_181),
.C(n_133),
.Y(n_326)
);

OAI21x1_ASAP7_75t_R g396 ( 
.A1(n_338),
.A2(n_292),
.B(n_242),
.Y(n_396)
);

NOR3xp33_ASAP7_75t_SL g340 ( 
.A(n_247),
.B(n_188),
.C(n_220),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_L g383 ( 
.A(n_340),
.B(n_354),
.Y(n_383)
);

AOI22xp33_ASAP7_75t_SL g341 ( 
.A1(n_253),
.A2(n_183),
.B1(n_197),
.B2(n_154),
.Y(n_341)
);

INVxp67_ASAP7_75t_L g382 ( 
.A(n_341),
.Y(n_382)
);

FAx1_ASAP7_75t_SL g343 ( 
.A(n_309),
.B(n_183),
.CI(n_220),
.CON(n_343),
.SN(n_343)
);

NOR2xp33_ASAP7_75t_SL g397 ( 
.A(n_343),
.B(n_252),
.Y(n_397)
);

OAI22xp5_ASAP7_75t_SL g350 ( 
.A1(n_293),
.A2(n_166),
.B1(n_200),
.B2(n_142),
.Y(n_350)
);

AOI22xp5_ASAP7_75t_L g405 ( 
.A1(n_350),
.A2(n_250),
.B1(n_258),
.B2(n_256),
.Y(n_405)
);

AOI32xp33_ASAP7_75t_L g354 ( 
.A1(n_245),
.A2(n_228),
.A3(n_166),
.B1(n_200),
.B2(n_142),
.Y(n_354)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_356),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_288),
.B(n_197),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_357),
.B(n_361),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_294),
.B(n_134),
.Y(n_361)
);

OAI22xp5_ASAP7_75t_L g422 ( 
.A1(n_363),
.A2(n_373),
.B1(n_287),
.B2(n_305),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_236),
.B(n_134),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_364),
.B(n_376),
.Y(n_395)
);

BUFx24_ASAP7_75t_SL g372 ( 
.A(n_235),
.Y(n_372)
);

NOR2xp33_ASAP7_75t_L g387 ( 
.A(n_372),
.B(n_255),
.Y(n_387)
);

CKINVDCx16_ASAP7_75t_R g411 ( 
.A(n_374),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_241),
.B(n_266),
.Y(n_376)
);

OR2x2_ASAP7_75t_L g377 ( 
.A(n_347),
.B(n_240),
.Y(n_377)
);

CKINVDCx14_ASAP7_75t_R g464 ( 
.A(n_377),
.Y(n_464)
);

XOR2xp5_ASAP7_75t_L g438 ( 
.A(n_378),
.B(n_370),
.Y(n_438)
);

OAI22xp5_ASAP7_75t_SL g379 ( 
.A1(n_363),
.A2(n_298),
.B1(n_313),
.B2(n_260),
.Y(n_379)
);

AOI22xp5_ASAP7_75t_L g457 ( 
.A1(n_379),
.A2(n_388),
.B1(n_406),
.B2(n_418),
.Y(n_457)
);

XNOR2xp5_ASAP7_75t_L g442 ( 
.A(n_380),
.B(n_378),
.Y(n_442)
);

AOI21xp5_ASAP7_75t_SL g381 ( 
.A1(n_375),
.A2(n_239),
.B(n_255),
.Y(n_381)
);

OAI21xp5_ASAP7_75t_SL g429 ( 
.A1(n_381),
.A2(n_390),
.B(n_399),
.Y(n_429)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_346),
.Y(n_385)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_385),
.Y(n_425)
);

AOI22xp33_ASAP7_75t_L g386 ( 
.A1(n_333),
.A2(n_291),
.B1(n_277),
.B2(n_238),
.Y(n_386)
);

OAI22xp5_ASAP7_75t_L g459 ( 
.A1(n_386),
.A2(n_410),
.B1(n_327),
.B2(n_325),
.Y(n_459)
);

NOR2xp33_ASAP7_75t_L g431 ( 
.A(n_387),
.B(n_392),
.Y(n_431)
);

OAI22xp5_ASAP7_75t_SL g388 ( 
.A1(n_373),
.A2(n_313),
.B1(n_279),
.B2(n_301),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_346),
.Y(n_389)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_389),
.Y(n_436)
);

CKINVDCx20_ASAP7_75t_R g392 ( 
.A(n_323),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_323),
.Y(n_393)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_393),
.Y(n_449)
);

INVx4_ASAP7_75t_L g394 ( 
.A(n_353),
.Y(n_394)
);

HB1xp67_ASAP7_75t_L g447 ( 
.A(n_394),
.Y(n_447)
);

AOI22xp5_ASAP7_75t_SL g452 ( 
.A1(n_396),
.A2(n_419),
.B1(n_422),
.B2(n_330),
.Y(n_452)
);

INVxp67_ASAP7_75t_L g458 ( 
.A(n_397),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_335),
.B(n_274),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_398),
.B(n_401),
.Y(n_437)
);

AOI21xp5_ASAP7_75t_SL g399 ( 
.A1(n_375),
.A2(n_263),
.B(n_237),
.Y(n_399)
);

OAI21xp5_ASAP7_75t_SL g400 ( 
.A1(n_318),
.A2(n_249),
.B(n_286),
.Y(n_400)
);

OAI21xp5_ASAP7_75t_SL g440 ( 
.A1(n_400),
.A2(n_414),
.B(n_392),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_335),
.B(n_243),
.Y(n_401)
);

MAJIxp5_ASAP7_75t_L g402 ( 
.A(n_324),
.B(n_270),
.C(n_257),
.Y(n_402)
);

MAJIxp5_ASAP7_75t_L g439 ( 
.A(n_402),
.B(n_349),
.C(n_331),
.Y(n_439)
);

NOR2xp33_ASAP7_75t_SL g403 ( 
.A(n_376),
.B(n_261),
.Y(n_403)
);

NOR2xp33_ASAP7_75t_L g433 ( 
.A(n_403),
.B(n_409),
.Y(n_433)
);

INVx3_ASAP7_75t_L g404 ( 
.A(n_353),
.Y(n_404)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_404),
.Y(n_460)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_405),
.Y(n_462)
);

OAI22xp5_ASAP7_75t_SL g406 ( 
.A1(n_329),
.A2(n_337),
.B1(n_332),
.B2(n_361),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_357),
.B(n_249),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g441 ( 
.A(n_407),
.B(n_412),
.Y(n_441)
);

AOI22xp33_ASAP7_75t_SL g408 ( 
.A1(n_350),
.A2(n_314),
.B1(n_285),
.B2(n_310),
.Y(n_408)
);

OAI21xp33_ASAP7_75t_SL g426 ( 
.A1(n_408),
.A2(n_421),
.B(n_423),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_SL g409 ( 
.A(n_365),
.B(n_290),
.Y(n_409)
);

AOI22xp5_ASAP7_75t_L g410 ( 
.A1(n_337),
.A2(n_302),
.B1(n_312),
.B2(n_311),
.Y(n_410)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_323),
.Y(n_412)
);

CKINVDCx20_ASAP7_75t_R g413 ( 
.A(n_360),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_413),
.B(n_415),
.Y(n_453)
);

OAI21x1_ASAP7_75t_L g414 ( 
.A1(n_343),
.A2(n_315),
.B(n_276),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_319),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_319),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_416),
.B(n_417),
.Y(n_463)
);

INVx2_ASAP7_75t_L g417 ( 
.A(n_336),
.Y(n_417)
);

OAI22xp5_ASAP7_75t_SL g418 ( 
.A1(n_332),
.A2(n_268),
.B1(n_283),
.B2(n_271),
.Y(n_418)
);

OAI22xp5_ASAP7_75t_SL g419 ( 
.A1(n_364),
.A2(n_321),
.B1(n_354),
.B2(n_334),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_321),
.B(n_320),
.Y(n_420)
);

XNOR2xp5_ASAP7_75t_SL g430 ( 
.A(n_420),
.B(n_326),
.Y(n_430)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_369),
.Y(n_421)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_369),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_356),
.Y(n_424)
);

CKINVDCx20_ASAP7_75t_R g432 ( 
.A(n_424),
.Y(n_432)
);

OAI21xp5_ASAP7_75t_L g427 ( 
.A1(n_399),
.A2(n_368),
.B(n_362),
.Y(n_427)
);

OAI21xp5_ASAP7_75t_SL g477 ( 
.A1(n_427),
.A2(n_440),
.B(n_444),
.Y(n_477)
);

OAI32xp33_ASAP7_75t_L g428 ( 
.A1(n_398),
.A2(n_317),
.A3(n_368),
.B1(n_328),
.B2(n_365),
.Y(n_428)
);

INVxp67_ASAP7_75t_L g478 ( 
.A(n_428),
.Y(n_478)
);

XOR2xp5_ASAP7_75t_L g488 ( 
.A(n_430),
.B(n_446),
.Y(n_488)
);

CKINVDCx20_ASAP7_75t_R g434 ( 
.A(n_410),
.Y(n_434)
);

NOR2xp33_ASAP7_75t_SL g492 ( 
.A(n_434),
.B(n_445),
.Y(n_492)
);

CKINVDCx16_ASAP7_75t_R g435 ( 
.A(n_418),
.Y(n_435)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_435),
.Y(n_468)
);

MAJIxp5_ASAP7_75t_L g475 ( 
.A(n_438),
.B(n_439),
.C(n_442),
.Y(n_475)
);

XOR2xp5_ASAP7_75t_L g443 ( 
.A(n_420),
.B(n_317),
.Y(n_443)
);

MAJIxp5_ASAP7_75t_L g486 ( 
.A(n_443),
.B(n_455),
.C(n_456),
.Y(n_486)
);

OAI21xp5_ASAP7_75t_SL g444 ( 
.A1(n_390),
.A2(n_345),
.B(n_355),
.Y(n_444)
);

CKINVDCx20_ASAP7_75t_R g445 ( 
.A(n_403),
.Y(n_445)
);

XNOR2xp5_ASAP7_75t_SL g446 ( 
.A(n_380),
.B(n_359),
.Y(n_446)
);

OAI22xp5_ASAP7_75t_SL g448 ( 
.A1(n_383),
.A2(n_340),
.B1(n_331),
.B2(n_330),
.Y(n_448)
);

AOI22xp5_ASAP7_75t_L g474 ( 
.A1(n_448),
.A2(n_397),
.B1(n_419),
.B2(n_388),
.Y(n_474)
);

OAI21xp5_ASAP7_75t_SL g450 ( 
.A1(n_414),
.A2(n_345),
.B(n_316),
.Y(n_450)
);

OAI21xp5_ASAP7_75t_L g472 ( 
.A1(n_450),
.A2(n_454),
.B(n_377),
.Y(n_472)
);

CKINVDCx20_ASAP7_75t_R g451 ( 
.A(n_407),
.Y(n_451)
);

AND2x2_ASAP7_75t_L g502 ( 
.A(n_451),
.B(n_452),
.Y(n_502)
);

AOI22xp5_ASAP7_75t_SL g454 ( 
.A1(n_422),
.A2(n_348),
.B1(n_367),
.B2(n_352),
.Y(n_454)
);

XOR2xp5_ASAP7_75t_L g455 ( 
.A(n_402),
.B(n_349),
.Y(n_455)
);

XOR2xp5_ASAP7_75t_L g456 ( 
.A(n_395),
.B(n_349),
.Y(n_456)
);

INVxp33_ASAP7_75t_L g491 ( 
.A(n_459),
.Y(n_491)
);

AOI21xp5_ASAP7_75t_L g461 ( 
.A1(n_400),
.A2(n_339),
.B(n_348),
.Y(n_461)
);

AOI21xp5_ASAP7_75t_L g503 ( 
.A1(n_461),
.A2(n_322),
.B(n_244),
.Y(n_503)
);

XNOR2xp5_ASAP7_75t_L g465 ( 
.A(n_395),
.B(n_325),
.Y(n_465)
);

MAJIxp5_ASAP7_75t_L g493 ( 
.A(n_465),
.B(n_446),
.C(n_430),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_L g466 ( 
.A(n_453),
.B(n_391),
.Y(n_466)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_466),
.Y(n_519)
);

XNOR2x2_ASAP7_75t_L g467 ( 
.A(n_441),
.B(n_377),
.Y(n_467)
);

XNOR2xp5_ASAP7_75t_L g516 ( 
.A(n_467),
.B(n_493),
.Y(n_516)
);

CKINVDCx20_ASAP7_75t_R g469 ( 
.A(n_463),
.Y(n_469)
);

INVxp67_ASAP7_75t_SL g512 ( 
.A(n_469),
.Y(n_512)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_463),
.Y(n_470)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_470),
.Y(n_507)
);

OAI22xp5_ASAP7_75t_SL g471 ( 
.A1(n_457),
.A2(n_379),
.B1(n_424),
.B2(n_384),
.Y(n_471)
);

AOI22xp5_ASAP7_75t_L g520 ( 
.A1(n_471),
.A2(n_456),
.B1(n_459),
.B2(n_433),
.Y(n_520)
);

INVx1_ASAP7_75t_SL g531 ( 
.A(n_472),
.Y(n_531)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_453),
.Y(n_473)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_473),
.Y(n_525)
);

OAI22xp5_ASAP7_75t_L g508 ( 
.A1(n_474),
.A2(n_481),
.B1(n_485),
.B2(n_487),
.Y(n_508)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_425),
.Y(n_476)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_476),
.Y(n_523)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_425),
.Y(n_479)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_479),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_SL g480 ( 
.A(n_458),
.B(n_413),
.Y(n_480)
);

NAND3xp33_ASAP7_75t_L g510 ( 
.A(n_480),
.B(n_484),
.C(n_431),
.Y(n_510)
);

AOI22xp5_ASAP7_75t_L g481 ( 
.A1(n_457),
.A2(n_406),
.B1(n_389),
.B2(n_385),
.Y(n_481)
);

CKINVDCx16_ASAP7_75t_R g482 ( 
.A(n_447),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_SL g505 ( 
.A(n_482),
.B(n_460),
.Y(n_505)
);

BUFx6f_ASAP7_75t_L g483 ( 
.A(n_460),
.Y(n_483)
);

INVx3_ASAP7_75t_L g537 ( 
.A(n_483),
.Y(n_537)
);

NOR2xp33_ASAP7_75t_L g484 ( 
.A(n_443),
.B(n_411),
.Y(n_484)
);

AOI22xp5_ASAP7_75t_L g485 ( 
.A1(n_435),
.A2(n_384),
.B1(n_382),
.B2(n_396),
.Y(n_485)
);

OAI22xp5_ASAP7_75t_L g487 ( 
.A1(n_431),
.A2(n_382),
.B1(n_396),
.B2(n_401),
.Y(n_487)
);

AOI22xp5_ASAP7_75t_L g489 ( 
.A1(n_434),
.A2(n_391),
.B1(n_393),
.B2(n_412),
.Y(n_489)
);

OAI22xp5_ASAP7_75t_L g509 ( 
.A1(n_489),
.A2(n_494),
.B1(n_496),
.B2(n_498),
.Y(n_509)
);

MAJIxp5_ASAP7_75t_R g490 ( 
.A(n_429),
.B(n_381),
.C(n_415),
.Y(n_490)
);

NOR2xp33_ASAP7_75t_L g513 ( 
.A(n_490),
.B(n_429),
.Y(n_513)
);

AOI22xp5_ASAP7_75t_L g494 ( 
.A1(n_432),
.A2(n_436),
.B1(n_451),
.B2(n_462),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_436),
.Y(n_495)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_495),
.Y(n_532)
);

AOI22xp5_ASAP7_75t_L g496 ( 
.A1(n_432),
.A2(n_416),
.B1(n_405),
.B2(n_423),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_L g497 ( 
.A(n_437),
.B(n_421),
.Y(n_497)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_497),
.Y(n_533)
);

AOI22xp5_ASAP7_75t_L g498 ( 
.A1(n_462),
.A2(n_417),
.B1(n_404),
.B2(n_394),
.Y(n_498)
);

AOI22xp5_ASAP7_75t_SL g499 ( 
.A1(n_464),
.A2(n_367),
.B1(n_366),
.B2(n_339),
.Y(n_499)
);

AND2x2_ASAP7_75t_L g529 ( 
.A(n_499),
.B(n_366),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_437),
.B(n_336),
.Y(n_500)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_500),
.Y(n_539)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_449),
.Y(n_501)
);

INVxp67_ASAP7_75t_L g535 ( 
.A(n_501),
.Y(n_535)
);

AOI21xp5_ASAP7_75t_L g538 ( 
.A1(n_503),
.A2(n_231),
.B(n_358),
.Y(n_538)
);

OAI22xp5_ASAP7_75t_SL g504 ( 
.A1(n_481),
.A2(n_452),
.B1(n_454),
.B2(n_464),
.Y(n_504)
);

AOI22xp5_ASAP7_75t_L g549 ( 
.A1(n_504),
.A2(n_517),
.B1(n_468),
.B2(n_472),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_L g568 ( 
.A(n_505),
.B(n_515),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_L g506 ( 
.A(n_497),
.B(n_441),
.Y(n_506)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_506),
.Y(n_550)
);

OAI22xp5_ASAP7_75t_L g547 ( 
.A1(n_510),
.A2(n_520),
.B1(n_522),
.B2(n_527),
.Y(n_547)
);

MAJIxp5_ASAP7_75t_L g511 ( 
.A(n_475),
.B(n_442),
.C(n_455),
.Y(n_511)
);

MAJIxp5_ASAP7_75t_L g551 ( 
.A(n_511),
.B(n_526),
.C(n_493),
.Y(n_551)
);

OAI21xp5_ASAP7_75t_SL g545 ( 
.A1(n_513),
.A2(n_524),
.B(n_538),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_L g514 ( 
.A(n_466),
.B(n_465),
.Y(n_514)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_514),
.Y(n_562)
);

CKINVDCx16_ASAP7_75t_R g515 ( 
.A(n_502),
.Y(n_515)
);

OAI22xp5_ASAP7_75t_SL g517 ( 
.A1(n_478),
.A2(n_445),
.B1(n_461),
.B2(n_449),
.Y(n_517)
);

NOR2xp33_ASAP7_75t_L g518 ( 
.A(n_478),
.B(n_433),
.Y(n_518)
);

CKINVDCx16_ASAP7_75t_R g554 ( 
.A(n_518),
.Y(n_554)
);

XNOR2xp5_ASAP7_75t_L g521 ( 
.A(n_488),
.B(n_438),
.Y(n_521)
);

XOR2xp5_ASAP7_75t_L g558 ( 
.A(n_521),
.B(n_514),
.Y(n_558)
);

AOI22xp5_ASAP7_75t_L g522 ( 
.A1(n_471),
.A2(n_426),
.B1(n_448),
.B2(n_427),
.Y(n_522)
);

OAI21xp5_ASAP7_75t_L g524 ( 
.A1(n_477),
.A2(n_444),
.B(n_440),
.Y(n_524)
);

MAJIxp5_ASAP7_75t_L g526 ( 
.A(n_475),
.B(n_439),
.C(n_450),
.Y(n_526)
);

OAI22xp5_ASAP7_75t_L g527 ( 
.A1(n_474),
.A2(n_428),
.B1(n_371),
.B2(n_327),
.Y(n_527)
);

FAx1_ASAP7_75t_SL g528 ( 
.A(n_467),
.B(n_322),
.CI(n_287),
.CON(n_528),
.SN(n_528)
);

NAND2xp5_ASAP7_75t_SL g543 ( 
.A(n_528),
.B(n_534),
.Y(n_543)
);

AND2x2_ASAP7_75t_L g566 ( 
.A(n_529),
.B(n_483),
.Y(n_566)
);

NOR2xp33_ASAP7_75t_L g534 ( 
.A(n_490),
.B(n_351),
.Y(n_534)
);

HB1xp67_ASAP7_75t_L g536 ( 
.A(n_489),
.Y(n_536)
);

HB1xp67_ASAP7_75t_L g560 ( 
.A(n_536),
.Y(n_560)
);

INVx11_ASAP7_75t_L g540 ( 
.A(n_528),
.Y(n_540)
);

INVx2_ASAP7_75t_L g580 ( 
.A(n_540),
.Y(n_580)
);

XNOR2xp5_ASAP7_75t_L g541 ( 
.A(n_511),
.B(n_526),
.Y(n_541)
);

XOR2xp5_ASAP7_75t_L g588 ( 
.A(n_541),
.B(n_542),
.Y(n_588)
);

XNOR2xp5_ASAP7_75t_SL g542 ( 
.A(n_521),
.B(n_488),
.Y(n_542)
);

XNOR2xp5_ASAP7_75t_L g544 ( 
.A(n_516),
.B(n_486),
.Y(n_544)
);

NOR2xp33_ASAP7_75t_L g581 ( 
.A(n_544),
.B(n_557),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_SL g546 ( 
.A(n_517),
.B(n_486),
.Y(n_546)
);

NAND3xp33_ASAP7_75t_L g591 ( 
.A(n_546),
.B(n_548),
.C(n_358),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_SL g548 ( 
.A(n_520),
.B(n_492),
.Y(n_548)
);

OAI22xp5_ASAP7_75t_L g572 ( 
.A1(n_549),
.A2(n_538),
.B1(n_519),
.B2(n_529),
.Y(n_572)
);

MAJIxp5_ASAP7_75t_L g578 ( 
.A(n_551),
.B(n_558),
.C(n_559),
.Y(n_578)
);

AOI22xp5_ASAP7_75t_L g552 ( 
.A1(n_508),
.A2(n_473),
.B1(n_502),
.B2(n_468),
.Y(n_552)
);

OAI22xp5_ASAP7_75t_SL g570 ( 
.A1(n_552),
.A2(n_553),
.B1(n_556),
.B2(n_564),
.Y(n_570)
);

AOI22xp5_ASAP7_75t_L g553 ( 
.A1(n_509),
.A2(n_502),
.B1(n_491),
.B2(n_492),
.Y(n_553)
);

OAI22xp5_ASAP7_75t_L g555 ( 
.A1(n_522),
.A2(n_494),
.B1(n_496),
.B2(n_469),
.Y(n_555)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_555),
.Y(n_587)
);

AOI22xp5_ASAP7_75t_L g556 ( 
.A1(n_504),
.A2(n_470),
.B1(n_500),
.B2(n_485),
.Y(n_556)
);

XNOR2xp5_ASAP7_75t_L g557 ( 
.A(n_516),
.B(n_477),
.Y(n_557)
);

MAJIxp5_ASAP7_75t_L g559 ( 
.A(n_531),
.B(n_479),
.C(n_476),
.Y(n_559)
);

MAJIxp5_ASAP7_75t_L g561 ( 
.A(n_531),
.B(n_495),
.C(n_501),
.Y(n_561)
);

MAJIxp5_ASAP7_75t_L g582 ( 
.A(n_561),
.B(n_563),
.C(n_532),
.Y(n_582)
);

XOR2xp5_ASAP7_75t_L g563 ( 
.A(n_524),
.B(n_499),
.Y(n_563)
);

AOI22xp5_ASAP7_75t_L g564 ( 
.A1(n_512),
.A2(n_533),
.B1(n_539),
.B2(n_525),
.Y(n_564)
);

OAI22xp5_ASAP7_75t_SL g565 ( 
.A1(n_533),
.A2(n_503),
.B1(n_498),
.B2(n_483),
.Y(n_565)
);

AOI22xp5_ASAP7_75t_SL g579 ( 
.A1(n_565),
.A2(n_532),
.B1(n_530),
.B2(n_523),
.Y(n_579)
);

AND2x2_ASAP7_75t_L g571 ( 
.A(n_566),
.B(n_537),
.Y(n_571)
);

BUFx2_ASAP7_75t_L g567 ( 
.A(n_537),
.Y(n_567)
);

INVx1_ASAP7_75t_SL g573 ( 
.A(n_567),
.Y(n_573)
);

OAI21xp5_ASAP7_75t_L g569 ( 
.A1(n_549),
.A2(n_507),
.B(n_539),
.Y(n_569)
);

AOI21xp5_ASAP7_75t_L g600 ( 
.A1(n_569),
.A2(n_590),
.B(n_545),
.Y(n_600)
);

INVxp67_ASAP7_75t_L g598 ( 
.A(n_571),
.Y(n_598)
);

XOR2xp5_ASAP7_75t_L g596 ( 
.A(n_572),
.B(n_563),
.Y(n_596)
);

AOI221xp5_ASAP7_75t_L g574 ( 
.A1(n_554),
.A2(n_562),
.B1(n_568),
.B2(n_550),
.C(n_559),
.Y(n_574)
);

AOI21xp33_ASAP7_75t_L g609 ( 
.A1(n_574),
.A2(n_585),
.B(n_586),
.Y(n_609)
);

OAI22xp5_ASAP7_75t_SL g575 ( 
.A1(n_553),
.A2(n_519),
.B1(n_506),
.B2(n_529),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_L g602 ( 
.A(n_575),
.B(n_583),
.Y(n_602)
);

NOR2xp33_ASAP7_75t_L g576 ( 
.A(n_560),
.B(n_535),
.Y(n_576)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_576),
.Y(n_592)
);

OAI22xp5_ASAP7_75t_L g577 ( 
.A1(n_556),
.A2(n_528),
.B1(n_535),
.B2(n_530),
.Y(n_577)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_577),
.Y(n_597)
);

XNOR2xp5_ASAP7_75t_L g593 ( 
.A(n_579),
.B(n_582),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_L g583 ( 
.A(n_564),
.B(n_523),
.Y(n_583)
);

OAI22xp5_ASAP7_75t_SL g584 ( 
.A1(n_552),
.A2(n_543),
.B1(n_547),
.B2(n_566),
.Y(n_584)
);

NOR2xp33_ASAP7_75t_L g595 ( 
.A(n_584),
.B(n_591),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_L g585 ( 
.A(n_561),
.B(n_322),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_L g586 ( 
.A(n_565),
.B(n_566),
.Y(n_586)
);

MAJIxp5_ASAP7_75t_L g589 ( 
.A(n_541),
.B(n_351),
.C(n_358),
.Y(n_589)
);

MAJIxp5_ASAP7_75t_L g594 ( 
.A(n_589),
.B(n_558),
.C(n_588),
.Y(n_594)
);

OAI21xp5_ASAP7_75t_SL g590 ( 
.A1(n_545),
.A2(n_269),
.B(n_304),
.Y(n_590)
);

XNOR2xp5_ASAP7_75t_L g611 ( 
.A(n_594),
.B(n_607),
.Y(n_611)
);

XOR2xp5_ASAP7_75t_L g622 ( 
.A(n_596),
.B(n_590),
.Y(n_622)
);

NOR2xp33_ASAP7_75t_SL g599 ( 
.A(n_578),
.B(n_581),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_L g612 ( 
.A(n_599),
.B(n_601),
.Y(n_612)
);

OR2x2_ASAP7_75t_L g616 ( 
.A(n_600),
.B(n_579),
.Y(n_616)
);

MAJIxp5_ASAP7_75t_L g601 ( 
.A(n_578),
.B(n_551),
.C(n_544),
.Y(n_601)
);

MAJIxp5_ASAP7_75t_L g603 ( 
.A(n_582),
.B(n_557),
.C(n_542),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_L g620 ( 
.A(n_603),
.B(n_604),
.Y(n_620)
);

XNOR2xp5_ASAP7_75t_L g604 ( 
.A(n_589),
.B(n_567),
.Y(n_604)
);

MAJIxp5_ASAP7_75t_L g605 ( 
.A(n_588),
.B(n_540),
.C(n_342),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_L g624 ( 
.A(n_605),
.B(n_606),
.Y(n_624)
);

MAJIxp5_ASAP7_75t_L g606 ( 
.A(n_585),
.B(n_342),
.C(n_371),
.Y(n_606)
);

XNOR2xp5_ASAP7_75t_L g607 ( 
.A(n_569),
.B(n_584),
.Y(n_607)
);

MAJIxp5_ASAP7_75t_L g608 ( 
.A(n_587),
.B(n_248),
.C(n_281),
.Y(n_608)
);

MAJIxp5_ASAP7_75t_L g625 ( 
.A(n_608),
.B(n_344),
.C(n_273),
.Y(n_625)
);

XOR2xp5_ASAP7_75t_L g610 ( 
.A(n_570),
.B(n_299),
.Y(n_610)
);

XNOR2xp5_ASAP7_75t_L g615 ( 
.A(n_610),
.B(n_577),
.Y(n_615)
);

AOI22xp5_ASAP7_75t_SL g613 ( 
.A1(n_595),
.A2(n_587),
.B1(n_570),
.B2(n_580),
.Y(n_613)
);

XNOR2xp5_ASAP7_75t_L g633 ( 
.A(n_613),
.B(n_625),
.Y(n_633)
);

OAI21x1_ASAP7_75t_L g614 ( 
.A1(n_592),
.A2(n_576),
.B(n_580),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_L g632 ( 
.A(n_614),
.B(n_616),
.Y(n_632)
);

XOR2xp5_ASAP7_75t_L g630 ( 
.A(n_615),
.B(n_622),
.Y(n_630)
);

AOI22xp5_ASAP7_75t_L g617 ( 
.A1(n_597),
.A2(n_575),
.B1(n_586),
.B2(n_583),
.Y(n_617)
);

OAI22xp5_ASAP7_75t_L g627 ( 
.A1(n_617),
.A2(n_618),
.B1(n_596),
.B2(n_605),
.Y(n_627)
);

AOI22xp5_ASAP7_75t_L g618 ( 
.A1(n_602),
.A2(n_572),
.B1(n_573),
.B2(n_571),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_598),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_L g635 ( 
.A(n_619),
.B(n_621),
.Y(n_635)
);

XNOR2xp5_ASAP7_75t_L g621 ( 
.A(n_593),
.B(n_571),
.Y(n_621)
);

OAI22xp5_ASAP7_75t_SL g623 ( 
.A1(n_598),
.A2(n_573),
.B1(n_344),
.B2(n_303),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_SL g631 ( 
.A(n_623),
.B(n_610),
.Y(n_631)
);

MAJIxp5_ASAP7_75t_L g626 ( 
.A(n_611),
.B(n_601),
.C(n_593),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_L g641 ( 
.A(n_626),
.B(n_627),
.Y(n_641)
);

NOR2xp33_ASAP7_75t_L g628 ( 
.A(n_612),
.B(n_608),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_SL g640 ( 
.A(n_628),
.B(n_629),
.Y(n_640)
);

NOR2xp33_ASAP7_75t_L g629 ( 
.A(n_611),
.B(n_594),
.Y(n_629)
);

NOR2xp33_ASAP7_75t_L g642 ( 
.A(n_631),
.B(n_615),
.Y(n_642)
);

MAJIxp5_ASAP7_75t_L g634 ( 
.A(n_620),
.B(n_603),
.C(n_606),
.Y(n_634)
);

XNOR2xp5_ASAP7_75t_L g639 ( 
.A(n_634),
.B(n_636),
.Y(n_639)
);

OAI21xp5_ASAP7_75t_SL g636 ( 
.A1(n_613),
.A2(n_609),
.B(n_273),
.Y(n_636)
);

MAJIxp5_ASAP7_75t_L g637 ( 
.A(n_626),
.B(n_621),
.C(n_624),
.Y(n_637)
);

NOR2xp33_ASAP7_75t_L g647 ( 
.A(n_637),
.B(n_638),
.Y(n_647)
);

MAJx2_ASAP7_75t_L g638 ( 
.A(n_632),
.B(n_616),
.C(n_622),
.Y(n_638)
);

AO21x1_ASAP7_75t_L g644 ( 
.A1(n_642),
.A2(n_643),
.B(n_633),
.Y(n_644)
);

BUFx24_ASAP7_75t_SL g643 ( 
.A(n_635),
.Y(n_643)
);

OAI21xp33_ASAP7_75t_L g648 ( 
.A1(n_644),
.A2(n_645),
.B(n_630),
.Y(n_648)
);

AND2x2_ASAP7_75t_L g645 ( 
.A(n_641),
.B(n_634),
.Y(n_645)
);

OAI22xp5_ASAP7_75t_SL g646 ( 
.A1(n_640),
.A2(n_633),
.B1(n_630),
.B2(n_625),
.Y(n_646)
);

INVxp33_ASAP7_75t_L g649 ( 
.A(n_646),
.Y(n_649)
);

NAND4xp25_ASAP7_75t_SL g650 ( 
.A(n_648),
.B(n_647),
.C(n_639),
.D(n_262),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_L g651 ( 
.A(n_650),
.B(n_647),
.Y(n_651)
);

OAI22xp5_ASAP7_75t_L g652 ( 
.A1(n_651),
.A2(n_649),
.B1(n_262),
.B2(n_307),
.Y(n_652)
);

MAJIxp5_ASAP7_75t_L g653 ( 
.A(n_652),
.B(n_264),
.C(n_262),
.Y(n_653)
);


endmodule