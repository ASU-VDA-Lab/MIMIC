module fake_jpeg_1117_n_556 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_556);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_556;

wire n_529;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_417;
wire n_362;
wire n_470;
wire n_172;
wire n_547;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_384;
wire n_296;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_541;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g19 ( 
.A(n_16),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

BUFx24_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_15),
.Y(n_25)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_18),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_1),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

BUFx4f_ASAP7_75t_L g31 ( 
.A(n_15),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_8),
.Y(n_32)
);

INVxp67_ASAP7_75t_L g33 ( 
.A(n_6),
.Y(n_33)
);

CKINVDCx14_ASAP7_75t_R g34 ( 
.A(n_15),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_10),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_10),
.Y(n_36)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_2),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_9),
.Y(n_38)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_3),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_8),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_7),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_13),
.Y(n_42)
);

CKINVDCx14_ASAP7_75t_R g43 ( 
.A(n_13),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_3),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_16),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_16),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_8),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_4),
.Y(n_48)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_14),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_8),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_12),
.Y(n_51)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_4),
.Y(n_52)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_20),
.Y(n_53)
);

INVx5_ASAP7_75t_L g168 ( 
.A(n_53),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_21),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_54),
.Y(n_106)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_19),
.Y(n_55)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_55),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_21),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_56),
.Y(n_116)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_52),
.Y(n_57)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_57),
.Y(n_109)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_52),
.Y(n_58)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_58),
.Y(n_123)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_26),
.Y(n_59)
);

BUFx2_ASAP7_75t_L g127 ( 
.A(n_59),
.Y(n_127)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_31),
.Y(n_60)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_60),
.Y(n_125)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_31),
.Y(n_61)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_61),
.Y(n_136)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_31),
.Y(n_62)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_62),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_28),
.B(n_45),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_63),
.B(n_68),
.Y(n_121)
);

INVx5_ASAP7_75t_L g64 ( 
.A(n_22),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g132 ( 
.A(n_64),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_34),
.Y(n_65)
);

CKINVDCx5p33_ASAP7_75t_R g107 ( 
.A(n_65),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_21),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_66),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_24),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_67),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_28),
.B(n_18),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_24),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_69),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_24),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g152 ( 
.A(n_70),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_25),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_71),
.B(n_74),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_45),
.B(n_18),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_SL g117 ( 
.A(n_72),
.B(n_84),
.Y(n_117)
);

BUFx5_ASAP7_75t_L g73 ( 
.A(n_23),
.Y(n_73)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_73),
.Y(n_108)
);

AND2x2_ASAP7_75t_L g74 ( 
.A(n_31),
.B(n_17),
.Y(n_74)
);

INVx6_ASAP7_75t_L g75 ( 
.A(n_42),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g163 ( 
.A(n_75),
.Y(n_163)
);

INVx6_ASAP7_75t_L g76 ( 
.A(n_42),
.Y(n_76)
);

INVx8_ASAP7_75t_L g126 ( 
.A(n_76),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_42),
.Y(n_77)
);

INVx6_ASAP7_75t_L g165 ( 
.A(n_77),
.Y(n_165)
);

AOI22xp33_ASAP7_75t_L g78 ( 
.A1(n_43),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_78)
);

OAI21xp5_ASAP7_75t_SL g141 ( 
.A1(n_78),
.A2(n_41),
.B(n_48),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_25),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_79),
.B(n_81),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_50),
.Y(n_80)
);

BUFx3_ASAP7_75t_L g149 ( 
.A(n_80),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_25),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_33),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_82),
.B(n_88),
.Y(n_146)
);

INVx5_ASAP7_75t_L g83 ( 
.A(n_22),
.Y(n_83)
);

BUFx3_ASAP7_75t_L g156 ( 
.A(n_83),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_19),
.B(n_46),
.Y(n_84)
);

BUFx3_ASAP7_75t_L g85 ( 
.A(n_36),
.Y(n_85)
);

INVx5_ASAP7_75t_L g110 ( 
.A(n_85),
.Y(n_110)
);

BUFx12f_ASAP7_75t_L g86 ( 
.A(n_37),
.Y(n_86)
);

BUFx4f_ASAP7_75t_SL g133 ( 
.A(n_86),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_50),
.Y(n_87)
);

INVx5_ASAP7_75t_L g112 ( 
.A(n_87),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_39),
.Y(n_88)
);

INVx13_ASAP7_75t_L g89 ( 
.A(n_23),
.Y(n_89)
);

BUFx24_ASAP7_75t_L g115 ( 
.A(n_89),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_39),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_90),
.B(n_40),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_50),
.Y(n_91)
);

INVx5_ASAP7_75t_L g118 ( 
.A(n_91),
.Y(n_118)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_26),
.Y(n_92)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_92),
.Y(n_139)
);

INVx2_ASAP7_75t_SL g93 ( 
.A(n_23),
.Y(n_93)
);

INVx4_ASAP7_75t_L g122 ( 
.A(n_93),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_39),
.Y(n_94)
);

INVx5_ASAP7_75t_L g142 ( 
.A(n_94),
.Y(n_142)
);

BUFx3_ASAP7_75t_L g95 ( 
.A(n_36),
.Y(n_95)
);

INVx5_ASAP7_75t_L g143 ( 
.A(n_95),
.Y(n_143)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_37),
.Y(n_96)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_96),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_20),
.Y(n_97)
);

INVx4_ASAP7_75t_L g134 ( 
.A(n_97),
.Y(n_134)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_46),
.Y(n_98)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_98),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_20),
.Y(n_99)
);

INVx4_ASAP7_75t_L g153 ( 
.A(n_99),
.Y(n_153)
);

INVx1_ASAP7_75t_SL g100 ( 
.A(n_20),
.Y(n_100)
);

AND2x2_ASAP7_75t_L g160 ( 
.A(n_100),
.B(n_40),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_27),
.Y(n_101)
);

INVx4_ASAP7_75t_L g158 ( 
.A(n_101),
.Y(n_158)
);

INVx6_ASAP7_75t_L g102 ( 
.A(n_27),
.Y(n_102)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_102),
.Y(n_148)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_27),
.Y(n_103)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_103),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_27),
.Y(n_104)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_104),
.Y(n_161)
);

INVx8_ASAP7_75t_SL g105 ( 
.A(n_23),
.Y(n_105)
);

BUFx2_ASAP7_75t_SL g155 ( 
.A(n_105),
.Y(n_155)
);

NAND2x1p5_ASAP7_75t_L g111 ( 
.A(n_74),
.B(n_49),
.Y(n_111)
);

AND2x2_ASAP7_75t_L g201 ( 
.A(n_111),
.B(n_160),
.Y(n_201)
);

BUFx4f_ASAP7_75t_L g113 ( 
.A(n_93),
.Y(n_113)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_113),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_94),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_SL g204 ( 
.A(n_114),
.B(n_128),
.Y(n_204)
);

AOI21xp33_ASAP7_75t_L g128 ( 
.A1(n_57),
.A2(n_51),
.B(n_30),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_102),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_SL g216 ( 
.A(n_129),
.B(n_138),
.Y(n_216)
);

INVx11_ASAP7_75t_L g130 ( 
.A(n_86),
.Y(n_130)
);

INVx4_ASAP7_75t_L g173 ( 
.A(n_130),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_58),
.B(n_30),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_100),
.A2(n_49),
.B1(n_40),
.B2(n_35),
.Y(n_140)
);

OA22x2_ASAP7_75t_L g186 ( 
.A1(n_140),
.A2(n_167),
.B1(n_64),
.B2(n_73),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_141),
.A2(n_77),
.B1(n_70),
.B2(n_69),
.Y(n_226)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_92),
.Y(n_151)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_151),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_75),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_154),
.B(n_166),
.Y(n_169)
);

A2O1A1Ixp33_ASAP7_75t_L g157 ( 
.A1(n_96),
.A2(n_41),
.B(n_48),
.C(n_38),
.Y(n_157)
);

HAxp5_ASAP7_75t_SL g210 ( 
.A(n_157),
.B(n_101),
.CON(n_210),
.SN(n_210)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_159),
.Y(n_193)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_61),
.Y(n_162)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_162),
.Y(n_219)
);

CKINVDCx12_ASAP7_75t_R g164 ( 
.A(n_89),
.Y(n_164)
);

BUFx8_ASAP7_75t_L g195 ( 
.A(n_164),
.Y(n_195)
);

OR2x2_ASAP7_75t_L g166 ( 
.A(n_78),
.B(n_51),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_SL g167 ( 
.A1(n_59),
.A2(n_40),
.B1(n_44),
.B2(n_35),
.Y(n_167)
);

BUFx3_ASAP7_75t_L g170 ( 
.A(n_110),
.Y(n_170)
);

BUFx3_ASAP7_75t_L g262 ( 
.A(n_170),
.Y(n_262)
);

INVx11_ASAP7_75t_L g171 ( 
.A(n_115),
.Y(n_171)
);

INVx1_ASAP7_75t_SL g235 ( 
.A(n_171),
.Y(n_235)
);

INVx8_ASAP7_75t_L g172 ( 
.A(n_106),
.Y(n_172)
);

INVx3_ASAP7_75t_L g250 ( 
.A(n_172),
.Y(n_250)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_136),
.Y(n_175)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_175),
.Y(n_231)
);

OR2x2_ASAP7_75t_L g177 ( 
.A(n_121),
.B(n_103),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g259 ( 
.A(n_177),
.B(n_178),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_107),
.Y(n_178)
);

BUFx10_ASAP7_75t_L g179 ( 
.A(n_115),
.Y(n_179)
);

INVx1_ASAP7_75t_SL g249 ( 
.A(n_179),
.Y(n_249)
);

BUFx3_ASAP7_75t_L g180 ( 
.A(n_143),
.Y(n_180)
);

INVx1_ASAP7_75t_SL g254 ( 
.A(n_180),
.Y(n_254)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_125),
.Y(n_181)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_181),
.Y(n_240)
);

OR2x4_ASAP7_75t_L g182 ( 
.A(n_111),
.B(n_43),
.Y(n_182)
);

NAND2xp33_ASAP7_75t_SL g266 ( 
.A(n_182),
.B(n_210),
.Y(n_266)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_137),
.Y(n_183)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_183),
.Y(n_248)
);

INVx3_ASAP7_75t_L g184 ( 
.A(n_168),
.Y(n_184)
);

INVx3_ASAP7_75t_L g251 ( 
.A(n_184),
.Y(n_251)
);

AOI22xp33_ASAP7_75t_SL g185 ( 
.A1(n_113),
.A2(n_44),
.B1(n_47),
.B2(n_83),
.Y(n_185)
);

AOI22xp33_ASAP7_75t_SL g246 ( 
.A1(n_185),
.A2(n_186),
.B1(n_206),
.B2(n_214),
.Y(n_246)
);

INVx8_ASAP7_75t_L g187 ( 
.A(n_106),
.Y(n_187)
);

INVx3_ASAP7_75t_L g280 ( 
.A(n_187),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_146),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_188),
.B(n_191),
.Y(n_233)
);

BUFx6f_ASAP7_75t_L g189 ( 
.A(n_116),
.Y(n_189)
);

INVx6_ASAP7_75t_L g232 ( 
.A(n_189),
.Y(n_232)
);

INVx11_ASAP7_75t_L g190 ( 
.A(n_115),
.Y(n_190)
);

INVx1_ASAP7_75t_SL g269 ( 
.A(n_190),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_117),
.B(n_86),
.Y(n_191)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_148),
.Y(n_192)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_192),
.Y(n_253)
);

INVx11_ASAP7_75t_L g194 ( 
.A(n_155),
.Y(n_194)
);

INVx2_ASAP7_75t_SL g263 ( 
.A(n_194),
.Y(n_263)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_124),
.Y(n_196)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_196),
.Y(n_238)
);

INVx11_ASAP7_75t_L g197 ( 
.A(n_130),
.Y(n_197)
);

CKINVDCx16_ASAP7_75t_R g261 ( 
.A(n_197),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_147),
.B(n_47),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_198),
.B(n_203),
.Y(n_244)
);

AOI22xp33_ASAP7_75t_L g199 ( 
.A1(n_157),
.A2(n_29),
.B1(n_32),
.B2(n_38),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_L g241 ( 
.A1(n_199),
.A2(n_112),
.B1(n_118),
.B2(n_165),
.Y(n_241)
);

BUFx5_ASAP7_75t_L g200 ( 
.A(n_150),
.Y(n_200)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_200),
.Y(n_271)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_120),
.Y(n_202)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_202),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_119),
.B(n_32),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_109),
.B(n_29),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_205),
.B(n_208),
.Y(n_247)
);

AOI22xp33_ASAP7_75t_SL g206 ( 
.A1(n_160),
.A2(n_85),
.B1(n_95),
.B2(n_122),
.Y(n_206)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_123),
.Y(n_207)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_207),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_122),
.B(n_53),
.Y(n_208)
);

AND2x2_ASAP7_75t_SL g209 ( 
.A(n_139),
.B(n_104),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_209),
.B(n_140),
.C(n_167),
.Y(n_237)
);

BUFx12_ASAP7_75t_L g211 ( 
.A(n_133),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_211),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_144),
.B(n_17),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_212),
.B(n_222),
.Y(n_258)
);

BUFx3_ASAP7_75t_L g213 ( 
.A(n_168),
.Y(n_213)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_213),
.Y(n_256)
);

INVx11_ASAP7_75t_L g214 ( 
.A(n_108),
.Y(n_214)
);

BUFx2_ASAP7_75t_L g215 ( 
.A(n_132),
.Y(n_215)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_215),
.Y(n_273)
);

INVx3_ASAP7_75t_L g217 ( 
.A(n_132),
.Y(n_217)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_217),
.Y(n_274)
);

INVx4_ASAP7_75t_L g218 ( 
.A(n_134),
.Y(n_218)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_218),
.Y(n_277)
);

INVx6_ASAP7_75t_L g220 ( 
.A(n_116),
.Y(n_220)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_220),
.Y(n_282)
);

BUFx6f_ASAP7_75t_L g221 ( 
.A(n_131),
.Y(n_221)
);

AOI22xp33_ASAP7_75t_SL g279 ( 
.A1(n_221),
.A2(n_225),
.B1(n_227),
.B2(n_0),
.Y(n_279)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_127),
.Y(n_222)
);

AND2x2_ASAP7_75t_L g223 ( 
.A(n_127),
.B(n_99),
.Y(n_223)
);

AND2x2_ASAP7_75t_L g236 ( 
.A(n_223),
.B(n_226),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_156),
.B(n_97),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_224),
.B(n_229),
.Y(n_260)
);

AOI22xp33_ASAP7_75t_SL g225 ( 
.A1(n_108),
.A2(n_91),
.B1(n_87),
.B2(n_80),
.Y(n_225)
);

AOI22xp33_ASAP7_75t_SL g227 ( 
.A1(n_156),
.A2(n_67),
.B1(n_66),
.B2(n_56),
.Y(n_227)
);

INVx4_ASAP7_75t_L g228 ( 
.A(n_134),
.Y(n_228)
);

AND2x2_ASAP7_75t_L g243 ( 
.A(n_228),
.B(n_230),
.Y(n_243)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_161),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_166),
.A2(n_54),
.B1(n_76),
.B2(n_17),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_204),
.B(n_163),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_234),
.B(n_252),
.Y(n_287)
);

AND2x2_ASAP7_75t_L g298 ( 
.A(n_237),
.B(n_241),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_201),
.A2(n_163),
.B1(n_126),
.B2(n_145),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_L g303 ( 
.A1(n_242),
.A2(n_268),
.B1(n_171),
.B2(n_190),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_216),
.B(n_165),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_201),
.A2(n_142),
.B1(n_153),
.B2(n_158),
.Y(n_255)
);

OR2x2_ASAP7_75t_L g293 ( 
.A(n_255),
.B(n_265),
.Y(n_293)
);

XOR2xp5_ASAP7_75t_L g257 ( 
.A(n_201),
.B(n_133),
.Y(n_257)
);

XOR2xp5_ASAP7_75t_L g295 ( 
.A(n_257),
.B(n_264),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_177),
.B(n_158),
.C(n_153),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_182),
.A2(n_169),
.B1(n_193),
.B2(n_210),
.Y(n_265)
);

AO22x2_ASAP7_75t_L g267 ( 
.A1(n_186),
.A2(n_126),
.B1(n_149),
.B2(n_145),
.Y(n_267)
);

INVx2_ASAP7_75t_L g314 ( 
.A(n_267),
.Y(n_314)
);

OAI22xp5_ASAP7_75t_L g268 ( 
.A1(n_226),
.A2(n_152),
.B1(n_135),
.B2(n_131),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_209),
.B(n_149),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_270),
.B(n_272),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_209),
.B(n_152),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_176),
.B(n_135),
.Y(n_276)
);

INVxp67_ASAP7_75t_L g296 ( 
.A(n_276),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_207),
.B(n_0),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_278),
.B(n_1),
.Y(n_324)
);

INVxp67_ASAP7_75t_L g306 ( 
.A(n_279),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_230),
.B(n_0),
.Y(n_281)
);

XOR2xp5_ASAP7_75t_L g320 ( 
.A(n_281),
.B(n_179),
.Y(n_320)
);

A2O1A1Ixp33_ASAP7_75t_L g283 ( 
.A1(n_195),
.A2(n_1),
.B(n_3),
.C(n_4),
.Y(n_283)
);

A2O1A1Ixp33_ASAP7_75t_L g308 ( 
.A1(n_283),
.A2(n_179),
.B(n_174),
.C(n_211),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_233),
.B(n_183),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_SL g348 ( 
.A(n_284),
.B(n_285),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_247),
.B(n_181),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_245),
.Y(n_286)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_286),
.Y(n_338)
);

OAI21xp33_ASAP7_75t_L g288 ( 
.A1(n_266),
.A2(n_195),
.B(n_179),
.Y(n_288)
);

INVxp33_ASAP7_75t_L g350 ( 
.A(n_288),
.Y(n_350)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_231),
.Y(n_289)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_289),
.Y(n_345)
);

OAI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_234),
.A2(n_186),
.B1(n_220),
.B2(n_223),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g340 ( 
.A1(n_290),
.A2(n_294),
.B1(n_305),
.B2(n_307),
.Y(n_340)
);

INVx13_ASAP7_75t_L g291 ( 
.A(n_275),
.Y(n_291)
);

BUFx12f_ASAP7_75t_L g356 ( 
.A(n_291),
.Y(n_356)
);

OAI21xp5_ASAP7_75t_L g292 ( 
.A1(n_266),
.A2(n_195),
.B(n_186),
.Y(n_292)
);

OAI21xp5_ASAP7_75t_SL g337 ( 
.A1(n_292),
.A2(n_269),
.B(n_263),
.Y(n_337)
);

OAI22xp5_ASAP7_75t_SL g294 ( 
.A1(n_265),
.A2(n_223),
.B1(n_189),
.B2(n_221),
.Y(n_294)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_231),
.Y(n_297)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_297),
.Y(n_346)
);

INVx13_ASAP7_75t_L g299 ( 
.A(n_249),
.Y(n_299)
);

INVxp67_ASAP7_75t_L g333 ( 
.A(n_299),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_SL g301 ( 
.A(n_259),
.B(n_184),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_SL g363 ( 
.A(n_301),
.B(n_313),
.Y(n_363)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_240),
.Y(n_302)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_302),
.Y(n_347)
);

AOI22xp33_ASAP7_75t_L g332 ( 
.A1(n_303),
.A2(n_309),
.B1(n_269),
.B2(n_263),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g304 ( 
.A(n_260),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g353 ( 
.A(n_304),
.B(n_310),
.Y(n_353)
);

OAI22xp5_ASAP7_75t_SL g305 ( 
.A1(n_236),
.A2(n_246),
.B1(n_252),
.B2(n_243),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_SL g307 ( 
.A1(n_236),
.A2(n_192),
.B1(n_187),
.B2(n_172),
.Y(n_307)
);

OAI21xp5_ASAP7_75t_L g351 ( 
.A1(n_308),
.A2(n_271),
.B(n_262),
.Y(n_351)
);

OAI22xp33_ASAP7_75t_SL g309 ( 
.A1(n_255),
.A2(n_228),
.B1(n_218),
.B2(n_213),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_278),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_SL g311 ( 
.A(n_264),
.B(n_175),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_311),
.B(n_315),
.Y(n_358)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_240),
.Y(n_312)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_312),
.Y(n_361)
);

NOR2xp33_ASAP7_75t_SL g313 ( 
.A(n_244),
.B(n_219),
.Y(n_313)
);

OAI32xp33_ASAP7_75t_L g315 ( 
.A1(n_243),
.A2(n_174),
.A3(n_214),
.B1(n_197),
.B2(n_200),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_SL g316 ( 
.A1(n_236),
.A2(n_243),
.B1(n_272),
.B2(n_242),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_L g342 ( 
.A1(n_316),
.A2(n_328),
.B1(n_329),
.B2(n_261),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_258),
.B(n_217),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_317),
.B(n_324),
.Y(n_367)
);

OAI22xp5_ASAP7_75t_L g318 ( 
.A1(n_237),
.A2(n_180),
.B1(n_170),
.B2(n_215),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_L g372 ( 
.A1(n_318),
.A2(n_330),
.B1(n_14),
.B2(n_306),
.Y(n_372)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_248),
.Y(n_319)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_319),
.Y(n_362)
);

XNOR2xp5_ASAP7_75t_L g349 ( 
.A(n_320),
.B(n_325),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_283),
.Y(n_321)
);

OR2x2_ASAP7_75t_L g370 ( 
.A(n_321),
.B(n_12),
.Y(n_370)
);

INVx13_ASAP7_75t_L g322 ( 
.A(n_249),
.Y(n_322)
);

INVxp67_ASAP7_75t_L g357 ( 
.A(n_322),
.Y(n_357)
);

INVx13_ASAP7_75t_L g323 ( 
.A(n_235),
.Y(n_323)
);

AOI22xp33_ASAP7_75t_SL g341 ( 
.A1(n_323),
.A2(n_327),
.B1(n_254),
.B2(n_262),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_270),
.B(n_173),
.Y(n_325)
);

INVx2_ASAP7_75t_L g326 ( 
.A(n_251),
.Y(n_326)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_326),
.Y(n_365)
);

INVx13_ASAP7_75t_L g327 ( 
.A(n_235),
.Y(n_327)
);

OAI22xp5_ASAP7_75t_SL g328 ( 
.A1(n_267),
.A2(n_173),
.B1(n_211),
.B2(n_194),
.Y(n_328)
);

OAI22xp5_ASAP7_75t_SL g329 ( 
.A1(n_267),
.A2(n_257),
.B1(n_281),
.B2(n_238),
.Y(n_329)
);

OAI22xp5_ASAP7_75t_L g330 ( 
.A1(n_267),
.A2(n_3),
.B1(n_5),
.B2(n_6),
.Y(n_330)
);

INVxp67_ASAP7_75t_L g331 ( 
.A(n_248),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g335 ( 
.A(n_331),
.Y(n_335)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_332),
.Y(n_375)
);

AOI22xp33_ASAP7_75t_L g334 ( 
.A1(n_314),
.A2(n_250),
.B1(n_280),
.B2(n_251),
.Y(n_334)
);

OAI22xp5_ASAP7_75t_L g389 ( 
.A1(n_334),
.A2(n_371),
.B1(n_303),
.B2(n_340),
.Y(n_389)
);

OAI22xp5_ASAP7_75t_SL g336 ( 
.A1(n_314),
.A2(n_282),
.B1(n_280),
.B2(n_250),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_336),
.B(n_344),
.Y(n_374)
);

OAI21xp5_ASAP7_75t_L g376 ( 
.A1(n_337),
.A2(n_339),
.B(n_354),
.Y(n_376)
);

AOI21xp5_ASAP7_75t_L g339 ( 
.A1(n_292),
.A2(n_263),
.B(n_254),
.Y(n_339)
);

BUFx2_ASAP7_75t_L g405 ( 
.A(n_341),
.Y(n_405)
);

AND2x2_ASAP7_75t_L g390 ( 
.A(n_342),
.B(n_372),
.Y(n_390)
);

AOI22xp5_ASAP7_75t_L g343 ( 
.A1(n_298),
.A2(n_274),
.B1(n_256),
.B2(n_273),
.Y(n_343)
);

OAI22xp5_ASAP7_75t_SL g392 ( 
.A1(n_343),
.A2(n_352),
.B1(n_364),
.B2(n_366),
.Y(n_392)
);

OAI22xp5_ASAP7_75t_SL g344 ( 
.A1(n_298),
.A2(n_232),
.B1(n_277),
.B2(n_253),
.Y(n_344)
);

OR2x2_ASAP7_75t_L g378 ( 
.A(n_351),
.B(n_339),
.Y(n_378)
);

AOI22xp5_ASAP7_75t_L g352 ( 
.A1(n_298),
.A2(n_253),
.B1(n_239),
.B2(n_271),
.Y(n_352)
);

OAI21xp5_ASAP7_75t_SL g354 ( 
.A1(n_293),
.A2(n_232),
.B(n_6),
.Y(n_354)
);

OAI22xp5_ASAP7_75t_SL g355 ( 
.A1(n_287),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_355),
.B(n_369),
.Y(n_385)
);

MAJIxp5_ASAP7_75t_L g359 ( 
.A(n_295),
.B(n_5),
.C(n_9),
.Y(n_359)
);

MAJIxp5_ASAP7_75t_L g380 ( 
.A(n_359),
.B(n_360),
.C(n_308),
.Y(n_380)
);

MAJIxp5_ASAP7_75t_L g360 ( 
.A(n_295),
.B(n_5),
.C(n_9),
.Y(n_360)
);

AOI22xp5_ASAP7_75t_L g364 ( 
.A1(n_329),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_364)
);

AOI22xp5_ASAP7_75t_L g366 ( 
.A1(n_290),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_366)
);

XNOR2xp5_ASAP7_75t_L g368 ( 
.A(n_311),
.B(n_11),
.Y(n_368)
);

XNOR2xp5_ASAP7_75t_SL g377 ( 
.A(n_368),
.B(n_320),
.Y(n_377)
);

OAI22xp5_ASAP7_75t_SL g369 ( 
.A1(n_287),
.A2(n_12),
.B1(n_14),
.B2(n_293),
.Y(n_369)
);

OAI21xp5_ASAP7_75t_L g397 ( 
.A1(n_370),
.A2(n_373),
.B(n_333),
.Y(n_397)
);

AOI22xp5_ASAP7_75t_L g371 ( 
.A1(n_305),
.A2(n_316),
.B1(n_293),
.B2(n_294),
.Y(n_371)
);

OR2x2_ASAP7_75t_L g373 ( 
.A(n_301),
.B(n_14),
.Y(n_373)
);

OAI21xp33_ASAP7_75t_L g384 ( 
.A1(n_373),
.A2(n_308),
.B(n_321),
.Y(n_384)
);

XNOR2xp5_ASAP7_75t_L g441 ( 
.A(n_377),
.B(n_382),
.Y(n_441)
);

OAI21xp5_ASAP7_75t_L g432 ( 
.A1(n_378),
.A2(n_350),
.B(n_370),
.Y(n_432)
);

INVx11_ASAP7_75t_L g379 ( 
.A(n_356),
.Y(n_379)
);

INVx4_ASAP7_75t_L g429 ( 
.A(n_379),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_SL g423 ( 
.A(n_380),
.B(n_400),
.Y(n_423)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_338),
.Y(n_381)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_381),
.Y(n_422)
);

MAJIxp5_ASAP7_75t_L g382 ( 
.A(n_349),
.B(n_310),
.C(n_318),
.Y(n_382)
);

BUFx6f_ASAP7_75t_L g383 ( 
.A(n_356),
.Y(n_383)
);

BUFx6f_ASAP7_75t_L g421 ( 
.A(n_383),
.Y(n_421)
);

CKINVDCx14_ASAP7_75t_R g410 ( 
.A(n_384),
.Y(n_410)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_338),
.Y(n_386)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_386),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_353),
.B(n_324),
.Y(n_387)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_387),
.Y(n_438)
);

CKINVDCx16_ASAP7_75t_R g388 ( 
.A(n_363),
.Y(n_388)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_388),
.Y(n_439)
);

OAI22xp5_ASAP7_75t_L g427 ( 
.A1(n_389),
.A2(n_406),
.B1(n_366),
.B2(n_346),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_367),
.B(n_300),
.Y(n_391)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_391),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_367),
.B(n_300),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_393),
.B(n_402),
.Y(n_424)
);

NOR2xp33_ASAP7_75t_L g394 ( 
.A(n_348),
.B(n_313),
.Y(n_394)
);

NOR2xp33_ASAP7_75t_SL g430 ( 
.A(n_394),
.B(n_395),
.Y(n_430)
);

NOR2xp33_ASAP7_75t_L g395 ( 
.A(n_348),
.B(n_304),
.Y(n_395)
);

NOR2xp33_ASAP7_75t_SL g396 ( 
.A(n_369),
.B(n_285),
.Y(n_396)
);

NAND3xp33_ASAP7_75t_L g425 ( 
.A(n_396),
.B(n_398),
.C(n_399),
.Y(n_425)
);

INVx1_ASAP7_75t_SL g431 ( 
.A(n_397),
.Y(n_431)
);

NOR2xp33_ASAP7_75t_L g398 ( 
.A(n_335),
.B(n_296),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_SL g399 ( 
.A(n_335),
.B(n_317),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_SL g400 ( 
.A(n_352),
.B(n_284),
.Y(n_400)
);

MAJIxp5_ASAP7_75t_SL g401 ( 
.A(n_371),
.B(n_328),
.C(n_330),
.Y(n_401)
);

OAI21xp5_ASAP7_75t_SL g419 ( 
.A1(n_401),
.A2(n_354),
.B(n_337),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_344),
.B(n_325),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_364),
.B(n_286),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g436 ( 
.A(n_403),
.B(n_404),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_358),
.B(n_315),
.Y(n_404)
);

OAI22xp5_ASAP7_75t_L g406 ( 
.A1(n_342),
.A2(n_307),
.B1(n_326),
.B2(n_297),
.Y(n_406)
);

CKINVDCx20_ASAP7_75t_R g407 ( 
.A(n_333),
.Y(n_407)
);

CKINVDCx20_ASAP7_75t_R g416 ( 
.A(n_407),
.Y(n_416)
);

INVx2_ASAP7_75t_L g408 ( 
.A(n_345),
.Y(n_408)
);

INVxp67_ASAP7_75t_L g412 ( 
.A(n_408),
.Y(n_412)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_345),
.Y(n_409)
);

NOR2xp33_ASAP7_75t_L g411 ( 
.A(n_409),
.B(n_365),
.Y(n_411)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_411),
.Y(n_447)
);

XOR2xp5_ASAP7_75t_L g413 ( 
.A(n_382),
.B(n_349),
.Y(n_413)
);

XOR2xp5_ASAP7_75t_L g451 ( 
.A(n_413),
.B(n_420),
.Y(n_451)
);

AO22x1_ASAP7_75t_L g414 ( 
.A1(n_389),
.A2(n_358),
.B1(n_336),
.B2(n_351),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g455 ( 
.A(n_414),
.B(n_432),
.Y(n_455)
);

OAI22xp5_ASAP7_75t_SL g415 ( 
.A1(n_404),
.A2(n_340),
.B1(n_370),
.B2(n_343),
.Y(n_415)
);

AOI22xp5_ASAP7_75t_L g448 ( 
.A1(n_415),
.A2(n_435),
.B1(n_402),
.B2(n_406),
.Y(n_448)
);

NOR2xp33_ASAP7_75t_L g417 ( 
.A(n_388),
.B(n_356),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_SL g456 ( 
.A(n_417),
.B(n_418),
.Y(n_456)
);

CKINVDCx20_ASAP7_75t_R g418 ( 
.A(n_383),
.Y(n_418)
);

NOR2xp33_ASAP7_75t_L g445 ( 
.A(n_419),
.B(n_433),
.Y(n_445)
);

XOR2xp5_ASAP7_75t_L g420 ( 
.A(n_377),
.B(n_368),
.Y(n_420)
);

BUFx6f_ASAP7_75t_L g426 ( 
.A(n_383),
.Y(n_426)
);

CKINVDCx20_ASAP7_75t_R g449 ( 
.A(n_426),
.Y(n_449)
);

OAI22xp5_ASAP7_75t_L g444 ( 
.A1(n_427),
.A2(n_375),
.B1(n_390),
.B2(n_403),
.Y(n_444)
);

NOR2xp33_ASAP7_75t_L g433 ( 
.A(n_387),
.B(n_396),
.Y(n_433)
);

NOR2xp33_ASAP7_75t_L g434 ( 
.A(n_391),
.B(n_356),
.Y(n_434)
);

CKINVDCx20_ASAP7_75t_R g462 ( 
.A(n_434),
.Y(n_462)
);

OAI22xp5_ASAP7_75t_SL g435 ( 
.A1(n_390),
.A2(n_346),
.B1(n_362),
.B2(n_361),
.Y(n_435)
);

BUFx3_ASAP7_75t_L g437 ( 
.A(n_405),
.Y(n_437)
);

AOI22xp33_ASAP7_75t_SL g453 ( 
.A1(n_437),
.A2(n_405),
.B1(n_379),
.B2(n_375),
.Y(n_453)
);

MAJIxp5_ASAP7_75t_L g442 ( 
.A(n_413),
.B(n_380),
.C(n_393),
.Y(n_442)
);

MAJIxp5_ASAP7_75t_L g475 ( 
.A(n_442),
.B(n_446),
.C(n_463),
.Y(n_475)
);

OAI22xp5_ASAP7_75t_SL g443 ( 
.A1(n_436),
.A2(n_378),
.B1(n_390),
.B2(n_376),
.Y(n_443)
);

AOI22xp5_ASAP7_75t_L g477 ( 
.A1(n_443),
.A2(n_444),
.B1(n_431),
.B2(n_416),
.Y(n_477)
);

MAJIxp5_ASAP7_75t_L g446 ( 
.A(n_441),
.B(n_407),
.C(n_359),
.Y(n_446)
);

OAI22xp5_ASAP7_75t_SL g486 ( 
.A1(n_448),
.A2(n_457),
.B1(n_465),
.B2(n_428),
.Y(n_486)
);

XNOR2xp5_ASAP7_75t_SL g450 ( 
.A(n_441),
.B(n_360),
.Y(n_450)
);

XOR2xp5_ASAP7_75t_L g470 ( 
.A(n_450),
.B(n_452),
.Y(n_470)
);

XOR2xp5_ASAP7_75t_L g452 ( 
.A(n_420),
.B(n_378),
.Y(n_452)
);

OAI21xp5_ASAP7_75t_SL g479 ( 
.A1(n_453),
.A2(n_419),
.B(n_426),
.Y(n_479)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_422),
.Y(n_454)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_454),
.Y(n_469)
);

AOI22xp5_ASAP7_75t_L g457 ( 
.A1(n_414),
.A2(n_415),
.B1(n_436),
.B2(n_376),
.Y(n_457)
);

XNOR2xp5_ASAP7_75t_SL g458 ( 
.A(n_423),
.B(n_397),
.Y(n_458)
);

XOR2xp5_ASAP7_75t_L g473 ( 
.A(n_458),
.B(n_459),
.Y(n_473)
);

XOR2xp5_ASAP7_75t_L g459 ( 
.A(n_440),
.B(n_409),
.Y(n_459)
);

OAI22xp5_ASAP7_75t_L g460 ( 
.A1(n_425),
.A2(n_385),
.B1(n_374),
.B2(n_405),
.Y(n_460)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_460),
.Y(n_482)
);

OAI22xp5_ASAP7_75t_L g461 ( 
.A1(n_430),
.A2(n_385),
.B1(n_374),
.B2(n_386),
.Y(n_461)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_461),
.Y(n_485)
);

MAJIxp5_ASAP7_75t_L g463 ( 
.A(n_440),
.B(n_401),
.C(n_381),
.Y(n_463)
);

OAI22xp5_ASAP7_75t_L g464 ( 
.A1(n_439),
.A2(n_408),
.B1(n_392),
.B2(n_361),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_464),
.B(n_466),
.Y(n_471)
);

AOI22xp5_ASAP7_75t_L g465 ( 
.A1(n_414),
.A2(n_392),
.B1(n_362),
.B2(n_347),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_422),
.Y(n_466)
);

XNOR2xp5_ASAP7_75t_L g467 ( 
.A(n_424),
.B(n_291),
.Y(n_467)
);

XNOR2xp5_ASAP7_75t_L g490 ( 
.A(n_467),
.B(n_357),
.Y(n_490)
);

XOR2xp5_ASAP7_75t_L g468 ( 
.A(n_424),
.B(n_291),
.Y(n_468)
);

XOR2xp5_ASAP7_75t_L g476 ( 
.A(n_468),
.B(n_435),
.Y(n_476)
);

CKINVDCx20_ASAP7_75t_R g472 ( 
.A(n_456),
.Y(n_472)
);

NOR2xp33_ASAP7_75t_SL g501 ( 
.A(n_472),
.B(n_474),
.Y(n_501)
);

CKINVDCx20_ASAP7_75t_R g474 ( 
.A(n_462),
.Y(n_474)
);

XNOR2xp5_ASAP7_75t_SL g493 ( 
.A(n_476),
.B(n_465),
.Y(n_493)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_477),
.Y(n_500)
);

AOI22xp5_ASAP7_75t_L g478 ( 
.A1(n_448),
.A2(n_431),
.B1(n_416),
.B2(n_410),
.Y(n_478)
);

AOI22xp5_ASAP7_75t_L g496 ( 
.A1(n_478),
.A2(n_483),
.B1(n_443),
.B2(n_468),
.Y(n_496)
);

NOR2xp33_ASAP7_75t_L g499 ( 
.A(n_479),
.B(n_489),
.Y(n_499)
);

MAJIxp5_ASAP7_75t_L g480 ( 
.A(n_442),
.B(n_412),
.C(n_438),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_SL g492 ( 
.A(n_480),
.B(n_481),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_SL g481 ( 
.A(n_447),
.B(n_439),
.Y(n_481)
);

AOI22xp5_ASAP7_75t_L g483 ( 
.A1(n_457),
.A2(n_438),
.B1(n_432),
.B2(n_412),
.Y(n_483)
);

MAJIxp5_ASAP7_75t_L g484 ( 
.A(n_451),
.B(n_428),
.C(n_347),
.Y(n_484)
);

MAJIxp5_ASAP7_75t_L g497 ( 
.A(n_484),
.B(n_487),
.C(n_488),
.Y(n_497)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_486),
.Y(n_505)
);

MAJIxp5_ASAP7_75t_L g487 ( 
.A(n_451),
.B(n_365),
.C(n_357),
.Y(n_487)
);

MAJIxp5_ASAP7_75t_L g488 ( 
.A(n_446),
.B(n_450),
.C(n_452),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_SL g489 ( 
.A(n_447),
.B(n_289),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_L g498 ( 
.A(n_490),
.B(n_467),
.Y(n_498)
);

AOI21xp5_ASAP7_75t_L g491 ( 
.A1(n_455),
.A2(n_429),
.B(n_437),
.Y(n_491)
);

OAI21xp5_ASAP7_75t_L g494 ( 
.A1(n_491),
.A2(n_455),
.B(n_463),
.Y(n_494)
);

XNOR2xp5_ASAP7_75t_L g511 ( 
.A(n_493),
.B(n_495),
.Y(n_511)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_494),
.Y(n_510)
);

XNOR2xp5_ASAP7_75t_L g495 ( 
.A(n_484),
.B(n_458),
.Y(n_495)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_496),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_L g514 ( 
.A(n_498),
.B(n_502),
.Y(n_514)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_469),
.Y(n_502)
);

CKINVDCx20_ASAP7_75t_R g503 ( 
.A(n_471),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_L g519 ( 
.A(n_503),
.B(n_507),
.Y(n_519)
);

AOI22xp5_ASAP7_75t_L g504 ( 
.A1(n_485),
.A2(n_445),
.B1(n_459),
.B2(n_454),
.Y(n_504)
);

OAI22xp5_ASAP7_75t_L g522 ( 
.A1(n_504),
.A2(n_506),
.B1(n_491),
.B2(n_476),
.Y(n_522)
);

AOI22xp5_ASAP7_75t_L g506 ( 
.A1(n_482),
.A2(n_466),
.B1(n_449),
.B2(n_421),
.Y(n_506)
);

NOR2xp33_ASAP7_75t_L g507 ( 
.A(n_480),
.B(n_429),
.Y(n_507)
);

NOR2xp33_ASAP7_75t_L g508 ( 
.A(n_475),
.B(n_421),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_L g521 ( 
.A(n_508),
.B(n_509),
.Y(n_521)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_478),
.Y(n_509)
);

MAJIxp5_ASAP7_75t_L g512 ( 
.A(n_497),
.B(n_475),
.C(n_487),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_512),
.B(n_513),
.Y(n_525)
);

MAJIxp5_ASAP7_75t_L g513 ( 
.A(n_497),
.B(n_488),
.C(n_486),
.Y(n_513)
);

XNOR2xp5_ASAP7_75t_L g516 ( 
.A(n_495),
.B(n_473),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_L g535 ( 
.A(n_516),
.B(n_518),
.Y(n_535)
);

AOI22xp5_ASAP7_75t_L g517 ( 
.A1(n_505),
.A2(n_471),
.B1(n_477),
.B2(n_483),
.Y(n_517)
);

INVxp67_ASAP7_75t_L g532 ( 
.A(n_517),
.Y(n_532)
);

CKINVDCx16_ASAP7_75t_R g518 ( 
.A(n_492),
.Y(n_518)
);

NOR2xp33_ASAP7_75t_L g520 ( 
.A(n_501),
.B(n_504),
.Y(n_520)
);

CKINVDCx14_ASAP7_75t_R g534 ( 
.A(n_520),
.Y(n_534)
);

XOR2xp5_ASAP7_75t_L g528 ( 
.A(n_522),
.B(n_523),
.Y(n_528)
);

AOI22xp5_ASAP7_75t_L g523 ( 
.A1(n_505),
.A2(n_473),
.B1(n_479),
.B2(n_490),
.Y(n_523)
);

MAJIxp5_ASAP7_75t_L g524 ( 
.A(n_500),
.B(n_470),
.C(n_302),
.Y(n_524)
);

MAJIxp5_ASAP7_75t_L g530 ( 
.A(n_524),
.B(n_498),
.C(n_493),
.Y(n_530)
);

NOR2xp33_ASAP7_75t_L g526 ( 
.A(n_515),
.B(n_506),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_L g541 ( 
.A(n_526),
.B(n_529),
.Y(n_541)
);

OAI21xp5_ASAP7_75t_SL g527 ( 
.A1(n_510),
.A2(n_499),
.B(n_494),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_SL g536 ( 
.A(n_527),
.B(n_530),
.Y(n_536)
);

NOR2xp33_ASAP7_75t_L g529 ( 
.A(n_513),
.B(n_500),
.Y(n_529)
);

BUFx24_ASAP7_75t_SL g531 ( 
.A(n_521),
.Y(n_531)
);

NOR2xp33_ASAP7_75t_SL g537 ( 
.A(n_531),
.B(n_512),
.Y(n_537)
);

OAI21xp5_ASAP7_75t_L g533 ( 
.A1(n_519),
.A2(n_496),
.B(n_470),
.Y(n_533)
);

CKINVDCx20_ASAP7_75t_R g542 ( 
.A(n_533),
.Y(n_542)
);

NAND3xp33_ASAP7_75t_L g546 ( 
.A(n_537),
.B(n_516),
.C(n_312),
.Y(n_546)
);

MAJIxp5_ASAP7_75t_L g538 ( 
.A(n_525),
.B(n_524),
.C(n_517),
.Y(n_538)
);

AOI21xp5_ASAP7_75t_L g543 ( 
.A1(n_538),
.A2(n_539),
.B(n_540),
.Y(n_543)
);

NOR2xp33_ASAP7_75t_L g539 ( 
.A(n_532),
.B(n_514),
.Y(n_539)
);

NOR2xp33_ASAP7_75t_L g540 ( 
.A(n_532),
.B(n_511),
.Y(n_540)
);

OAI22xp5_ASAP7_75t_L g544 ( 
.A1(n_542),
.A2(n_534),
.B1(n_535),
.B2(n_528),
.Y(n_544)
);

XOR2xp5_ASAP7_75t_L g548 ( 
.A(n_544),
.B(n_538),
.Y(n_548)
);

AO22x1_ASAP7_75t_L g545 ( 
.A1(n_541),
.A2(n_528),
.B1(n_523),
.B2(n_511),
.Y(n_545)
);

OAI21xp5_ASAP7_75t_L g547 ( 
.A1(n_545),
.A2(n_546),
.B(n_536),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_L g550 ( 
.A(n_547),
.B(n_548),
.Y(n_550)
);

OAI21xp5_ASAP7_75t_L g549 ( 
.A1(n_543),
.A2(n_319),
.B(n_355),
.Y(n_549)
);

NOR2xp33_ASAP7_75t_L g551 ( 
.A(n_549),
.B(n_299),
.Y(n_551)
);

AOI21xp5_ASAP7_75t_SL g552 ( 
.A1(n_551),
.A2(n_299),
.B(n_322),
.Y(n_552)
);

MAJIxp5_ASAP7_75t_L g553 ( 
.A(n_552),
.B(n_322),
.C(n_323),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_SL g554 ( 
.A(n_553),
.B(n_550),
.Y(n_554)
);

NOR2xp33_ASAP7_75t_L g555 ( 
.A(n_554),
.B(n_323),
.Y(n_555)
);

OAI21x1_ASAP7_75t_L g556 ( 
.A1(n_555),
.A2(n_327),
.B(n_501),
.Y(n_556)
);


endmodule