module fake_jpeg_8130_n_70 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_26, n_9, n_5, n_11, n_17, n_25, n_2, n_12, n_8, n_15, n_7, n_70);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_70;

wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_69;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_40;
wire n_59;
wire n_35;
wire n_48;
wire n_68;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_65;
wire n_63;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_44;
wire n_38;
wire n_28;
wire n_36;
wire n_62;
wire n_31;
wire n_56;
wire n_67;
wire n_37;
wire n_29;
wire n_43;
wire n_50;
wire n_32;
wire n_66;

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_18),
.B(n_25),
.Y(n_28)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_27),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_21),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_22),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_24),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_16),
.Y(n_33)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_19),
.Y(n_34)
);

AOI22xp33_ASAP7_75t_SL g35 ( 
.A1(n_31),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_35)
);

AOI21xp5_ASAP7_75t_L g44 ( 
.A1(n_35),
.A2(n_4),
.B(n_5),
.Y(n_44)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_33),
.Y(n_36)
);

INVx5_ASAP7_75t_L g45 ( 
.A(n_36),
.Y(n_45)
);

BUFx2_ASAP7_75t_L g37 ( 
.A(n_30),
.Y(n_37)
);

INVx1_ASAP7_75t_SL g49 ( 
.A(n_37),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_L g38 ( 
.A1(n_31),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_L g51 ( 
.A1(n_38),
.A2(n_42),
.B1(n_6),
.B2(n_7),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_29),
.B(n_3),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_SL g52 ( 
.A(n_39),
.B(n_6),
.Y(n_52)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_30),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_40),
.B(n_9),
.Y(n_55)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_29),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_41),
.B(n_34),
.Y(n_43)
);

OAI22xp33_ASAP7_75t_L g42 ( 
.A1(n_34),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_43),
.B(n_46),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_44),
.A2(n_53),
.B1(n_55),
.B2(n_26),
.Y(n_61)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_39),
.Y(n_46)
);

BUFx10_ASAP7_75t_L g47 ( 
.A(n_37),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_47),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_41),
.B(n_32),
.Y(n_48)
);

A2O1A1O1Ixp25_ASAP7_75t_L g56 ( 
.A1(n_48),
.A2(n_52),
.B(n_28),
.C(n_10),
.D(n_12),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_36),
.A2(n_33),
.B1(n_7),
.B2(n_8),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_50),
.A2(n_51),
.B1(n_11),
.B2(n_15),
.Y(n_59)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_36),
.Y(n_53)
);

OA22x2_ASAP7_75t_L g54 ( 
.A1(n_37),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g58 ( 
.A1(n_54),
.A2(n_40),
.B1(n_13),
.B2(n_14),
.Y(n_58)
);

XOR2xp5_ASAP7_75t_L g64 ( 
.A(n_56),
.B(n_58),
.Y(n_64)
);

MAJIxp5_ASAP7_75t_L g63 ( 
.A(n_59),
.B(n_60),
.C(n_61),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_51),
.A2(n_17),
.B1(n_20),
.B2(n_23),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g65 ( 
.A1(n_64),
.A2(n_58),
.B1(n_45),
.B2(n_54),
.Y(n_65)
);

MAJIxp5_ASAP7_75t_L g66 ( 
.A(n_65),
.B(n_63),
.C(n_44),
.Y(n_66)
);

XNOR2xp5_ASAP7_75t_L g67 ( 
.A(n_66),
.B(n_56),
.Y(n_67)
);

OR2x2_ASAP7_75t_L g68 ( 
.A(n_67),
.B(n_57),
.Y(n_68)
);

AOI322xp5_ASAP7_75t_L g69 ( 
.A1(n_68),
.A2(n_61),
.A3(n_62),
.B1(n_54),
.B2(n_49),
.C1(n_47),
.C2(n_45),
.Y(n_69)
);

OAI221xp5_ASAP7_75t_L g70 ( 
.A1(n_69),
.A2(n_47),
.B1(n_49),
.B2(n_54),
.C(n_65),
.Y(n_70)
);


endmodule