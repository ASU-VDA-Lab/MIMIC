module fake_jpeg_11388_n_374 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_374);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_374;

wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx5_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_16),
.Y(n_19)
);

BUFx12_ASAP7_75t_L g20 ( 
.A(n_16),
.Y(n_20)
);

INVx6_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_14),
.Y(n_22)
);

BUFx10_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_15),
.Y(n_25)
);

INVx8_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_16),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_3),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_4),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_15),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_14),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_1),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_14),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_6),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_5),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_7),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_10),
.Y(n_41)
);

CKINVDCx16_ASAP7_75t_R g42 ( 
.A(n_15),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_4),
.B(n_5),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_9),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_3),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_8),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_6),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_2),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_4),
.Y(n_49)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_6),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_3),
.Y(n_51)
);

INVx11_ASAP7_75t_L g52 ( 
.A(n_4),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_10),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_13),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_51),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_55),
.Y(n_113)
);

INVx4_ASAP7_75t_SL g56 ( 
.A(n_23),
.Y(n_56)
);

CKINVDCx6p67_ASAP7_75t_R g143 ( 
.A(n_56),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g57 ( 
.A1(n_29),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_57),
.A2(n_101),
.B1(n_39),
.B2(n_48),
.Y(n_148)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_30),
.Y(n_58)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_58),
.Y(n_118)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_22),
.Y(n_59)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_59),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_20),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_60),
.B(n_61),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_20),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_20),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_62),
.B(n_65),
.Y(n_122)
);

BUFx5_ASAP7_75t_L g63 ( 
.A(n_17),
.Y(n_63)
);

INVx4_ASAP7_75t_L g112 ( 
.A(n_63),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_43),
.B(n_13),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_64),
.B(n_103),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_20),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_25),
.B(n_7),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_66),
.B(n_88),
.Y(n_137)
);

INVx8_ASAP7_75t_L g67 ( 
.A(n_17),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_67),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_51),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g142 ( 
.A(n_68),
.Y(n_142)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_29),
.Y(n_69)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_69),
.Y(n_117)
);

CKINVDCx16_ASAP7_75t_R g70 ( 
.A(n_23),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_70),
.B(n_71),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_23),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_51),
.Y(n_72)
);

INVx6_ASAP7_75t_L g120 ( 
.A(n_72),
.Y(n_120)
);

INVx8_ASAP7_75t_L g73 ( 
.A(n_23),
.Y(n_73)
);

INVx3_ASAP7_75t_SL g116 ( 
.A(n_73),
.Y(n_116)
);

INVx8_ASAP7_75t_L g74 ( 
.A(n_23),
.Y(n_74)
);

INVx3_ASAP7_75t_L g133 ( 
.A(n_74),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_19),
.Y(n_75)
);

INVx8_ASAP7_75t_L g152 ( 
.A(n_75),
.Y(n_152)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_30),
.Y(n_76)
);

INVx3_ASAP7_75t_L g145 ( 
.A(n_76),
.Y(n_145)
);

INVx6_ASAP7_75t_L g77 ( 
.A(n_19),
.Y(n_77)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_77),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_19),
.Y(n_78)
);

INVx4_ASAP7_75t_L g149 ( 
.A(n_78),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_28),
.Y(n_79)
);

INVx4_ASAP7_75t_L g159 ( 
.A(n_79),
.Y(n_159)
);

BUFx4f_ASAP7_75t_L g80 ( 
.A(n_52),
.Y(n_80)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_80),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_28),
.Y(n_81)
);

INVx4_ASAP7_75t_L g173 ( 
.A(n_81),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_43),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_82),
.B(n_84),
.Y(n_130)
);

BUFx12f_ASAP7_75t_L g83 ( 
.A(n_33),
.Y(n_83)
);

CKINVDCx9p33_ASAP7_75t_R g115 ( 
.A(n_83),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_SL g84 ( 
.A(n_25),
.B(n_7),
.Y(n_84)
);

NAND2x1_ASAP7_75t_SL g85 ( 
.A(n_35),
.B(n_40),
.Y(n_85)
);

CKINVDCx16_ASAP7_75t_R g111 ( 
.A(n_85),
.Y(n_111)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_50),
.Y(n_86)
);

HB1xp67_ASAP7_75t_L g119 ( 
.A(n_86),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_28),
.Y(n_87)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_87),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_37),
.B(n_12),
.Y(n_88)
);

INVx5_ASAP7_75t_L g89 ( 
.A(n_30),
.Y(n_89)
);

HB1xp67_ASAP7_75t_L g153 ( 
.A(n_89),
.Y(n_153)
);

NAND2x1_ASAP7_75t_L g90 ( 
.A(n_35),
.B(n_0),
.Y(n_90)
);

A2O1A1Ixp33_ASAP7_75t_L g129 ( 
.A1(n_90),
.A2(n_18),
.B(n_24),
.C(n_36),
.Y(n_129)
);

BUFx2_ASAP7_75t_L g91 ( 
.A(n_50),
.Y(n_91)
);

INVxp67_ASAP7_75t_L g135 ( 
.A(n_91),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_33),
.Y(n_92)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_92),
.Y(n_170)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_22),
.Y(n_93)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_93),
.Y(n_139)
);

BUFx12_ASAP7_75t_L g94 ( 
.A(n_52),
.Y(n_94)
);

CKINVDCx12_ASAP7_75t_R g154 ( 
.A(n_94),
.Y(n_154)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_33),
.Y(n_95)
);

HB1xp67_ASAP7_75t_L g162 ( 
.A(n_95),
.Y(n_162)
);

INVx1_ASAP7_75t_SL g96 ( 
.A(n_49),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g141 ( 
.A(n_96),
.B(n_98),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_49),
.Y(n_97)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_97),
.Y(n_171)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_40),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_37),
.B(n_11),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_99),
.B(n_110),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_49),
.Y(n_100)
);

CKINVDCx9p33_ASAP7_75t_R g169 ( 
.A(n_100),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_21),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_101)
);

BUFx3_ASAP7_75t_L g102 ( 
.A(n_34),
.Y(n_102)
);

AND2x2_ASAP7_75t_L g164 ( 
.A(n_102),
.B(n_108),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_41),
.B(n_53),
.Y(n_103)
);

CKINVDCx16_ASAP7_75t_R g104 ( 
.A(n_42),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_104),
.B(n_106),
.Y(n_144)
);

AOI21xp33_ASAP7_75t_L g105 ( 
.A1(n_41),
.A2(n_8),
.B(n_10),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_SL g124 ( 
.A(n_105),
.B(n_1),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_SL g106 ( 
.A(n_53),
.B(n_8),
.Y(n_106)
);

AND2x2_ASAP7_75t_L g107 ( 
.A(n_34),
.B(n_11),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_107),
.B(n_32),
.Y(n_157)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_34),
.Y(n_108)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_18),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_109),
.B(n_36),
.Y(n_147)
);

HB1xp67_ASAP7_75t_L g110 ( 
.A(n_27),
.Y(n_110)
);

O2A1O1Ixp33_ASAP7_75t_SL g114 ( 
.A1(n_90),
.A2(n_42),
.B(n_48),
.C(n_47),
.Y(n_114)
);

A2O1A1Ixp33_ASAP7_75t_L g202 ( 
.A1(n_114),
.A2(n_102),
.B(n_74),
.C(n_92),
.Y(n_202)
);

AOI21xp33_ASAP7_75t_L g174 ( 
.A1(n_124),
.A2(n_45),
.B(n_6),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_107),
.B(n_44),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_125),
.B(n_126),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_85),
.B(n_44),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_94),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_128),
.B(n_136),
.Y(n_182)
);

OAI21xp33_ASAP7_75t_L g224 ( 
.A1(n_129),
.A2(n_143),
.B(n_154),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_57),
.B(n_46),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_131),
.B(n_156),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_SL g136 ( 
.A(n_56),
.B(n_54),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_91),
.A2(n_26),
.B1(n_21),
.B2(n_46),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_SL g177 ( 
.A1(n_146),
.A2(n_155),
.B1(n_115),
.B2(n_169),
.Y(n_177)
);

AND2x2_ASAP7_75t_L g196 ( 
.A(n_147),
.B(n_166),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_148),
.A2(n_150),
.B1(n_165),
.B2(n_73),
.Y(n_195)
);

OAI22xp33_ASAP7_75t_SL g150 ( 
.A1(n_101),
.A2(n_27),
.B1(n_24),
.B2(n_21),
.Y(n_150)
);

CKINVDCx11_ASAP7_75t_R g151 ( 
.A(n_67),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_151),
.B(n_163),
.Y(n_185)
);

AOI22xp33_ASAP7_75t_SL g155 ( 
.A1(n_86),
.A2(n_26),
.B1(n_54),
.B2(n_38),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_95),
.B(n_32),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_SL g178 ( 
.A(n_157),
.B(n_63),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_77),
.B(n_38),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_158),
.B(n_125),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_94),
.Y(n_163)
);

OAI22xp33_ASAP7_75t_SL g165 ( 
.A1(n_75),
.A2(n_26),
.B1(n_31),
.B2(n_39),
.Y(n_165)
);

AND2x2_ASAP7_75t_SL g166 ( 
.A(n_58),
.B(n_76),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_96),
.B(n_31),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_167),
.B(n_135),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_89),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_168),
.B(n_83),
.Y(n_192)
);

AOI22xp33_ASAP7_75t_L g172 ( 
.A1(n_55),
.A2(n_45),
.B1(n_47),
.B2(n_3),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_172),
.A2(n_68),
.B1(n_72),
.B2(n_81),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_SL g230 ( 
.A(n_174),
.B(n_179),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_162),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_175),
.B(n_178),
.Y(n_233)
);

CKINVDCx16_ASAP7_75t_R g176 ( 
.A(n_115),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_176),
.B(n_194),
.Y(n_248)
);

INVxp67_ASAP7_75t_L g249 ( 
.A(n_177),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_SL g179 ( 
.A(n_130),
.B(n_83),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_180),
.A2(n_184),
.B1(n_213),
.B2(n_221),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_123),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_181),
.B(n_188),
.Y(n_241)
);

BUFx6f_ASAP7_75t_L g183 ( 
.A(n_113),
.Y(n_183)
);

INVx3_ASAP7_75t_L g260 ( 
.A(n_183),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_L g184 ( 
.A1(n_131),
.A2(n_87),
.B1(n_79),
.B2(n_78),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_SL g186 ( 
.A(n_144),
.B(n_140),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_SL g236 ( 
.A(n_186),
.B(n_201),
.Y(n_236)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_158),
.Y(n_187)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_187),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_156),
.Y(n_188)
);

BUFx6f_ASAP7_75t_L g190 ( 
.A(n_113),
.Y(n_190)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_190),
.Y(n_252)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_170),
.Y(n_191)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_191),
.Y(n_250)
);

CKINVDCx16_ASAP7_75t_R g258 ( 
.A(n_192),
.Y(n_258)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_170),
.Y(n_193)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_193),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_160),
.B(n_137),
.Y(n_194)
);

OR2x2_ASAP7_75t_L g231 ( 
.A(n_195),
.B(n_212),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_198),
.B(n_206),
.Y(n_234)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_171),
.Y(n_199)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_199),
.Y(n_254)
);

BUFx8_ASAP7_75t_L g200 ( 
.A(n_169),
.Y(n_200)
);

CKINVDCx16_ASAP7_75t_R g245 ( 
.A(n_200),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_132),
.B(n_108),
.Y(n_201)
);

AO22x1_ASAP7_75t_L g243 ( 
.A1(n_202),
.A2(n_223),
.B1(n_196),
.B2(n_178),
.Y(n_243)
);

INVx8_ASAP7_75t_L g203 ( 
.A(n_127),
.Y(n_203)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_203),
.Y(n_256)
);

BUFx6f_ASAP7_75t_L g204 ( 
.A(n_142),
.Y(n_204)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_204),
.Y(n_255)
);

AOI22xp33_ASAP7_75t_L g205 ( 
.A1(n_111),
.A2(n_97),
.B1(n_100),
.B2(n_80),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_L g232 ( 
.A1(n_205),
.A2(n_116),
.B1(n_142),
.B2(n_133),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_129),
.B(n_80),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_126),
.B(n_139),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_207),
.B(n_208),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_117),
.B(n_166),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_121),
.B(n_122),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_209),
.B(n_211),
.Y(n_244)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_138),
.Y(n_210)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_210),
.Y(n_261)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_138),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_L g213 ( 
.A1(n_114),
.A2(n_117),
.B1(n_120),
.B2(n_134),
.Y(n_213)
);

INVx3_ASAP7_75t_L g214 ( 
.A(n_127),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_214),
.B(n_215),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_143),
.B(n_141),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_166),
.A2(n_164),
.B1(n_141),
.B2(n_112),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_SL g238 ( 
.A1(n_216),
.A2(n_224),
.B(n_208),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_141),
.B(n_134),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_217),
.B(n_220),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_143),
.B(n_119),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_218),
.B(n_219),
.Y(n_264)
);

INVxp67_ASAP7_75t_L g219 ( 
.A(n_164),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_143),
.B(n_153),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_161),
.A2(n_120),
.B1(n_173),
.B2(n_149),
.Y(n_221)
);

BUFx2_ASAP7_75t_L g222 ( 
.A(n_152),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_222),
.A2(n_223),
.B1(n_225),
.B2(n_219),
.Y(n_237)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_164),
.Y(n_223)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_161),
.Y(n_225)
);

OAI32xp33_ASAP7_75t_L g226 ( 
.A1(n_197),
.A2(n_112),
.A3(n_173),
.B1(n_159),
.B2(n_149),
.Y(n_226)
);

AOI32xp33_ASAP7_75t_L g277 ( 
.A1(n_226),
.A2(n_200),
.A3(n_190),
.B1(n_183),
.B2(n_204),
.Y(n_277)
);

OA22x2_ASAP7_75t_L g227 ( 
.A1(n_195),
.A2(n_159),
.B1(n_152),
.B2(n_133),
.Y(n_227)
);

A2O1A1Ixp33_ASAP7_75t_SL g278 ( 
.A1(n_227),
.A2(n_235),
.B(n_243),
.C(n_200),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_188),
.B(n_118),
.C(n_145),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_228),
.B(n_229),
.C(n_246),
.Y(n_274)
);

OAI21xp5_ASAP7_75t_L g229 ( 
.A1(n_206),
.A2(n_135),
.B(n_118),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g291 ( 
.A1(n_232),
.A2(n_240),
.B1(n_251),
.B2(n_259),
.Y(n_291)
);

OA22x2_ASAP7_75t_L g235 ( 
.A1(n_202),
.A2(n_116),
.B1(n_145),
.B2(n_187),
.Y(n_235)
);

CKINVDCx16_ASAP7_75t_R g281 ( 
.A(n_237),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_SL g265 ( 
.A(n_238),
.B(n_175),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_197),
.A2(n_198),
.B1(n_216),
.B2(n_207),
.Y(n_240)
);

OAI21xp5_ASAP7_75t_L g246 ( 
.A1(n_196),
.A2(n_189),
.B(n_182),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_189),
.A2(n_196),
.B1(n_217),
.B2(n_186),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_199),
.A2(n_193),
.B1(n_191),
.B2(n_214),
.Y(n_259)
);

A2O1A1Ixp33_ASAP7_75t_L g262 ( 
.A1(n_185),
.A2(n_181),
.B(n_179),
.C(n_212),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_262),
.B(n_200),
.Y(n_268)
);

OAI21xp5_ASAP7_75t_SL g305 ( 
.A1(n_265),
.A2(n_288),
.B(n_290),
.Y(n_305)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_254),
.Y(n_266)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_266),
.Y(n_297)
);

INVx3_ASAP7_75t_L g267 ( 
.A(n_256),
.Y(n_267)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_267),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_SL g299 ( 
.A(n_268),
.B(n_269),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_SL g269 ( 
.A(n_241),
.B(n_210),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_248),
.B(n_222),
.Y(n_270)
);

INVxp67_ASAP7_75t_L g298 ( 
.A(n_270),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_234),
.B(n_225),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_271),
.B(n_276),
.C(n_283),
.Y(n_303)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_254),
.Y(n_272)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_272),
.Y(n_314)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_250),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_273),
.B(n_275),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_SL g275 ( 
.A(n_236),
.B(n_203),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_257),
.B(n_221),
.C(n_222),
.Y(n_276)
);

AO21x1_ASAP7_75t_L g302 ( 
.A1(n_277),
.A2(n_278),
.B(n_281),
.Y(n_302)
);

AOI22xp33_ASAP7_75t_L g279 ( 
.A1(n_231),
.A2(n_183),
.B1(n_190),
.B2(n_204),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_L g295 ( 
.A1(n_279),
.A2(n_292),
.B1(n_242),
.B2(n_237),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_259),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_280),
.B(n_284),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_L g282 ( 
.A1(n_231),
.A2(n_234),
.B1(n_239),
.B2(n_242),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g315 ( 
.A1(n_282),
.A2(n_287),
.B1(n_272),
.B2(n_266),
.Y(n_315)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_251),
.B(n_240),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_SL g284 ( 
.A(n_244),
.B(n_236),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_258),
.B(n_233),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_285),
.B(n_286),
.Y(n_308)
);

HB1xp67_ASAP7_75t_L g286 ( 
.A(n_256),
.Y(n_286)
);

BUFx6f_ASAP7_75t_L g287 ( 
.A(n_252),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_246),
.B(n_230),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_L g289 ( 
.A(n_257),
.B(n_263),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_289),
.B(n_250),
.C(n_227),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_SL g290 ( 
.A(n_239),
.B(n_263),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_229),
.A2(n_231),
.B1(n_235),
.B2(n_243),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_SL g293 ( 
.A(n_230),
.B(n_243),
.C(n_264),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_293),
.B(n_235),
.C(n_247),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_228),
.B(n_238),
.Y(n_294)
);

XOR2xp5_ASAP7_75t_L g311 ( 
.A(n_294),
.B(n_232),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_L g329 ( 
.A1(n_295),
.A2(n_301),
.B1(n_311),
.B2(n_313),
.Y(n_329)
);

OAI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_292),
.A2(n_249),
.B1(n_235),
.B2(n_227),
.Y(n_301)
);

AOI21xp5_ASAP7_75t_L g325 ( 
.A1(n_302),
.A2(n_306),
.B(n_307),
.Y(n_325)
);

MAJx2_ASAP7_75t_L g319 ( 
.A(n_304),
.B(n_313),
.C(n_274),
.Y(n_319)
);

OAI21xp5_ASAP7_75t_SL g306 ( 
.A1(n_294),
.A2(n_249),
.B(n_262),
.Y(n_306)
);

AOI21xp5_ASAP7_75t_L g307 ( 
.A1(n_293),
.A2(n_226),
.B(n_227),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_289),
.B(n_261),
.C(n_253),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_310),
.B(n_311),
.C(n_274),
.Y(n_318)
);

OAI21xp5_ASAP7_75t_L g312 ( 
.A1(n_268),
.A2(n_261),
.B(n_253),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_312),
.B(n_291),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_315),
.B(n_273),
.Y(n_327)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_297),
.Y(n_316)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_316),
.Y(n_340)
);

CKINVDCx20_ASAP7_75t_R g317 ( 
.A(n_296),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_317),
.B(n_323),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_318),
.B(n_319),
.C(n_321),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_SL g338 ( 
.A(n_320),
.B(n_324),
.Y(n_338)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_303),
.B(n_283),
.C(n_271),
.Y(n_321)
);

OAI21xp33_ASAP7_75t_L g322 ( 
.A1(n_299),
.A2(n_278),
.B(n_276),
.Y(n_322)
);

NAND3xp33_ASAP7_75t_L g335 ( 
.A(n_322),
.B(n_326),
.C(n_330),
.Y(n_335)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_297),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_SL g324 ( 
.A(n_296),
.B(n_305),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_SL g326 ( 
.A(n_305),
.B(n_291),
.Y(n_326)
);

OAI22xp5_ASAP7_75t_L g342 ( 
.A1(n_327),
.A2(n_329),
.B1(n_331),
.B2(n_313),
.Y(n_342)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_303),
.B(n_278),
.C(n_267),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_328),
.B(n_303),
.C(n_311),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_308),
.B(n_287),
.Y(n_330)
);

AOI221xp5_ASAP7_75t_L g331 ( 
.A1(n_312),
.A2(n_278),
.B1(n_255),
.B2(n_245),
.C(n_260),
.Y(n_331)
);

AOI21xp5_ASAP7_75t_L g333 ( 
.A1(n_325),
.A2(n_302),
.B(n_306),
.Y(n_333)
);

AOI21xp5_ASAP7_75t_SL g349 ( 
.A1(n_333),
.A2(n_341),
.B(n_343),
.Y(n_349)
);

MAJIxp5_ASAP7_75t_L g346 ( 
.A(n_334),
.B(n_321),
.C(n_318),
.Y(n_346)
);

CKINVDCx20_ASAP7_75t_R g336 ( 
.A(n_327),
.Y(n_336)
);

AND2x2_ASAP7_75t_L g345 ( 
.A(n_336),
.B(n_315),
.Y(n_345)
);

OAI22xp5_ASAP7_75t_SL g339 ( 
.A1(n_329),
.A2(n_302),
.B1(n_307),
.B2(n_304),
.Y(n_339)
);

AOI22xp5_ASAP7_75t_L g352 ( 
.A1(n_339),
.A2(n_342),
.B1(n_308),
.B2(n_323),
.Y(n_352)
);

AOI21xp5_ASAP7_75t_L g341 ( 
.A1(n_325),
.A2(n_320),
.B(n_328),
.Y(n_341)
);

AOI22xp5_ASAP7_75t_SL g343 ( 
.A1(n_326),
.A2(n_301),
.B1(n_295),
.B2(n_298),
.Y(n_343)
);

OAI21xp5_ASAP7_75t_SL g344 ( 
.A1(n_341),
.A2(n_317),
.B(n_299),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_SL g356 ( 
.A(n_344),
.B(n_345),
.Y(n_356)
);

MAJIxp5_ASAP7_75t_L g353 ( 
.A(n_346),
.B(n_350),
.C(n_338),
.Y(n_353)
);

XNOR2xp5_ASAP7_75t_L g347 ( 
.A(n_332),
.B(n_319),
.Y(n_347)
);

XOR2xp5_ASAP7_75t_L g354 ( 
.A(n_347),
.B(n_348),
.Y(n_354)
);

XNOR2xp5_ASAP7_75t_L g348 ( 
.A(n_332),
.B(n_334),
.Y(n_348)
);

MAJIxp5_ASAP7_75t_L g350 ( 
.A(n_339),
.B(n_319),
.C(n_310),
.Y(n_350)
);

OAI21xp5_ASAP7_75t_L g351 ( 
.A1(n_335),
.A2(n_324),
.B(n_309),
.Y(n_351)
);

XOR2xp5_ASAP7_75t_L g359 ( 
.A(n_351),
.B(n_352),
.Y(n_359)
);

MAJIxp5_ASAP7_75t_L g363 ( 
.A(n_353),
.B(n_314),
.C(n_300),
.Y(n_363)
);

AOI21xp5_ASAP7_75t_L g355 ( 
.A1(n_345),
.A2(n_333),
.B(n_343),
.Y(n_355)
);

OAI21xp5_ASAP7_75t_SL g361 ( 
.A1(n_355),
.A2(n_349),
.B(n_337),
.Y(n_361)
);

OAI31xp33_ASAP7_75t_L g357 ( 
.A1(n_349),
.A2(n_336),
.A3(n_337),
.B(n_340),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_357),
.B(n_358),
.Y(n_360)
);

INVx6_ASAP7_75t_L g358 ( 
.A(n_348),
.Y(n_358)
);

OAI21xp5_ASAP7_75t_L g367 ( 
.A1(n_361),
.A2(n_356),
.B(n_355),
.Y(n_367)
);

AOI322xp5_ASAP7_75t_L g362 ( 
.A1(n_356),
.A2(n_309),
.A3(n_350),
.B1(n_340),
.B2(n_316),
.C1(n_314),
.C2(n_346),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_SL g366 ( 
.A(n_362),
.B(n_363),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_SL g364 ( 
.A(n_359),
.B(n_300),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_L g365 ( 
.A(n_364),
.B(n_359),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_365),
.B(n_367),
.Y(n_368)
);

INVxp67_ASAP7_75t_L g369 ( 
.A(n_366),
.Y(n_369)
);

OAI22xp33_ASAP7_75t_L g371 ( 
.A1(n_369),
.A2(n_360),
.B1(n_358),
.B2(n_357),
.Y(n_371)
);

MAJIxp5_ASAP7_75t_L g370 ( 
.A(n_366),
.B(n_353),
.C(n_354),
.Y(n_370)
);

AOI211xp5_ASAP7_75t_L g372 ( 
.A1(n_370),
.A2(n_354),
.B(n_255),
.C(n_260),
.Y(n_372)
);

MAJIxp5_ASAP7_75t_L g373 ( 
.A(n_371),
.B(n_372),
.C(n_368),
.Y(n_373)
);

XNOR2xp5_ASAP7_75t_L g374 ( 
.A(n_373),
.B(n_252),
.Y(n_374)
);


endmodule