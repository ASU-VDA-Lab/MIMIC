module fake_jpeg_27337_n_196 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_196);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_196;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_140;
wire n_96;

BUFx5_ASAP7_75t_L g14 ( 
.A(n_1),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_13),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_2),
.Y(n_16)
);

BUFx5_ASAP7_75t_L g17 ( 
.A(n_13),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_9),
.Y(n_20)
);

INVx13_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

INVx5_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_0),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_1),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_SL g32 ( 
.A(n_16),
.B(n_0),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_SL g51 ( 
.A(n_32),
.B(n_42),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g33 ( 
.A1(n_26),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_33),
.B(n_39),
.Y(n_53)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_19),
.Y(n_34)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_34),
.Y(n_68)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_19),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_35),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_27),
.Y(n_36)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_36),
.Y(n_46)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_19),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_37),
.Y(n_69)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_21),
.Y(n_38)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_38),
.Y(n_59)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_16),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_19),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g76 ( 
.A(n_40),
.Y(n_76)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_25),
.Y(n_41)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_41),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_20),
.B(n_12),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_25),
.B(n_4),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_43),
.B(n_25),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_SL g44 ( 
.A(n_20),
.B(n_31),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_44),
.B(n_31),
.Y(n_66)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_25),
.Y(n_45)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_45),
.Y(n_65)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_36),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_47),
.B(n_57),
.Y(n_77)
);

INVx5_ASAP7_75t_L g48 ( 
.A(n_40),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_48),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g49 ( 
.A(n_43),
.B(n_27),
.C(n_15),
.Y(n_49)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_49),
.B(n_15),
.C(n_14),
.Y(n_99)
);

BUFx16f_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

INVx13_ASAP7_75t_L g85 ( 
.A(n_50),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_L g52 ( 
.A1(n_34),
.A2(n_45),
.B1(n_37),
.B2(n_35),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_52),
.A2(n_15),
.B1(n_14),
.B2(n_6),
.Y(n_97)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_55),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_39),
.A2(n_27),
.B1(n_26),
.B2(n_21),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_56),
.A2(n_70),
.B1(n_24),
.B2(n_23),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_44),
.B(n_30),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_58),
.B(n_66),
.Y(n_100)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_40),
.Y(n_60)
);

BUFx2_ASAP7_75t_L g94 ( 
.A(n_60),
.Y(n_94)
);

BUFx2_ASAP7_75t_L g61 ( 
.A(n_41),
.Y(n_61)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_61),
.Y(n_83)
);

INVx5_ASAP7_75t_L g62 ( 
.A(n_41),
.Y(n_62)
);

INVx5_ASAP7_75t_SL g98 ( 
.A(n_62),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_32),
.B(n_30),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_64),
.B(n_67),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_41),
.B(n_29),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_34),
.A2(n_26),
.B1(n_21),
.B2(n_29),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_44),
.B(n_17),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_71),
.B(n_72),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_42),
.Y(n_72)
);

INVx1_ASAP7_75t_SL g73 ( 
.A(n_43),
.Y(n_73)
);

INVx13_ASAP7_75t_L g91 ( 
.A(n_73),
.Y(n_91)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_40),
.Y(n_74)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_74),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_44),
.B(n_17),
.Y(n_75)
);

INVxp67_ASAP7_75t_L g80 ( 
.A(n_75),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_73),
.B(n_28),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_78),
.B(n_63),
.Y(n_107)
);

OAI21xp5_ASAP7_75t_L g79 ( 
.A1(n_53),
.A2(n_28),
.B(n_24),
.Y(n_79)
);

OAI21xp5_ASAP7_75t_L g113 ( 
.A1(n_79),
.A2(n_95),
.B(n_56),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_81),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_46),
.A2(n_68),
.B1(n_65),
.B2(n_52),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_86),
.A2(n_102),
.B1(n_60),
.B2(n_62),
.Y(n_117)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_61),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_88),
.B(n_101),
.Y(n_125)
);

BUFx5_ASAP7_75t_L g89 ( 
.A(n_76),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_89),
.B(n_76),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_46),
.A2(n_23),
.B1(n_22),
.B2(n_18),
.Y(n_92)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_92),
.Y(n_119)
);

A2O1A1Ixp33_ASAP7_75t_L g95 ( 
.A1(n_51),
.A2(n_18),
.B(n_22),
.C(n_17),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_54),
.A2(n_15),
.B1(n_14),
.B2(n_6),
.Y(n_96)
);

A2O1A1Ixp33_ASAP7_75t_SL g124 ( 
.A1(n_96),
.A2(n_4),
.B(n_7),
.C(n_8),
.Y(n_124)
);

AND2x2_ASAP7_75t_L g103 ( 
.A(n_97),
.B(n_99),
.Y(n_103)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_63),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_70),
.A2(n_4),
.B1(n_5),
.B2(n_7),
.Y(n_102)
);

CKINVDCx16_ASAP7_75t_R g135 ( 
.A(n_104),
.Y(n_135)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_82),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_105),
.B(n_109),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_77),
.B(n_59),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_106),
.B(n_108),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_SL g126 ( 
.A(n_107),
.B(n_112),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_87),
.B(n_59),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_90),
.B(n_12),
.Y(n_109)
);

AND2x2_ASAP7_75t_L g111 ( 
.A(n_99),
.B(n_69),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_L g141 ( 
.A1(n_111),
.A2(n_113),
.B(n_119),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_94),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_80),
.B(n_74),
.Y(n_114)
);

CKINVDCx16_ASAP7_75t_R g137 ( 
.A(n_114),
.Y(n_137)
);

INVx6_ASAP7_75t_L g115 ( 
.A(n_82),
.Y(n_115)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_115),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_80),
.B(n_55),
.Y(n_116)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_116),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_117),
.A2(n_118),
.B1(n_93),
.B2(n_85),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_86),
.A2(n_54),
.B1(n_69),
.B2(n_7),
.Y(n_118)
);

MAJx2_ASAP7_75t_L g120 ( 
.A(n_91),
.B(n_50),
.C(n_5),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_120),
.B(n_84),
.C(n_98),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_79),
.B(n_10),
.Y(n_121)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_121),
.Y(n_142)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_94),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_122),
.B(n_123),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_94),
.Y(n_123)
);

AOI21xp5_ASAP7_75t_L g131 ( 
.A1(n_124),
.A2(n_102),
.B(n_97),
.Y(n_131)
);

BUFx5_ASAP7_75t_L g127 ( 
.A(n_105),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_127),
.B(n_89),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_L g152 ( 
.A1(n_131),
.A2(n_141),
.B(n_119),
.Y(n_152)
);

AOI22xp33_ASAP7_75t_L g132 ( 
.A1(n_113),
.A2(n_91),
.B1(n_101),
.B2(n_78),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_132),
.A2(n_134),
.B1(n_143),
.B2(n_144),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_110),
.A2(n_100),
.B1(n_98),
.B2(n_84),
.Y(n_134)
);

XNOR2xp5_ASAP7_75t_SL g138 ( 
.A(n_107),
.B(n_95),
.Y(n_138)
);

XOR2xp5_ASAP7_75t_L g154 ( 
.A(n_138),
.B(n_139),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_111),
.B(n_83),
.C(n_88),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_140),
.B(n_111),
.C(n_120),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_110),
.A2(n_98),
.B1(n_83),
.B2(n_93),
.Y(n_143)
);

INVxp67_ASAP7_75t_L g164 ( 
.A(n_145),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_L g162 ( 
.A(n_146),
.B(n_155),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_SL g147 ( 
.A(n_129),
.B(n_117),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_147),
.B(n_148),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_128),
.B(n_125),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_130),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_149),
.B(n_150),
.Y(n_160)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_130),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_SL g159 ( 
.A(n_152),
.B(n_158),
.Y(n_159)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_126),
.Y(n_153)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_153),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_140),
.B(n_103),
.C(n_120),
.Y(n_155)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_127),
.Y(n_156)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_156),
.Y(n_167)
);

AOI21xp5_ASAP7_75t_L g157 ( 
.A1(n_141),
.A2(n_103),
.B(n_124),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_157),
.A2(n_131),
.B1(n_144),
.B2(n_129),
.Y(n_163)
);

A2O1A1O1Ixp25_ASAP7_75t_L g158 ( 
.A1(n_138),
.A2(n_139),
.B(n_103),
.C(n_126),
.D(n_134),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_163),
.B(n_151),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_SL g166 ( 
.A(n_154),
.B(n_155),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_166),
.B(n_154),
.C(n_146),
.Y(n_172)
);

AOI322xp5_ASAP7_75t_L g168 ( 
.A1(n_152),
.A2(n_143),
.A3(n_137),
.B1(n_135),
.B2(n_118),
.C1(n_142),
.C2(n_136),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_168),
.B(n_149),
.Y(n_174)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_147),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_169),
.B(n_170),
.Y(n_176)
);

HB1xp67_ASAP7_75t_L g170 ( 
.A(n_156),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_SL g181 ( 
.A1(n_171),
.A2(n_142),
.B(n_160),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_172),
.B(n_174),
.C(n_177),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_L g173 ( 
.A1(n_161),
.A2(n_165),
.B1(n_153),
.B2(n_157),
.Y(n_173)
);

INVxp67_ASAP7_75t_L g184 ( 
.A(n_173),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_164),
.B(n_136),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_175),
.B(n_178),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_166),
.B(n_150),
.C(n_158),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_164),
.B(n_137),
.Y(n_178)
);

BUFx24_ASAP7_75t_SL g179 ( 
.A(n_176),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_179),
.B(n_183),
.Y(n_187)
);

AOI21xp5_ASAP7_75t_L g189 ( 
.A1(n_181),
.A2(n_167),
.B(n_124),
.Y(n_189)
);

AOI21xp5_ASAP7_75t_SL g183 ( 
.A1(n_177),
.A2(n_159),
.B(n_135),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_182),
.B(n_184),
.Y(n_185)
);

AOI21xp5_ASAP7_75t_L g192 ( 
.A1(n_185),
.A2(n_186),
.B(n_133),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g186 ( 
.A(n_180),
.B(n_172),
.Y(n_186)
);

NOR2x1_ASAP7_75t_L g188 ( 
.A(n_181),
.B(n_159),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_188),
.A2(n_189),
.B1(n_124),
.B2(n_162),
.Y(n_190)
);

INVxp67_ASAP7_75t_L g193 ( 
.A(n_190),
.Y(n_193)
);

AOI322xp5_ASAP7_75t_L g191 ( 
.A1(n_188),
.A2(n_162),
.A3(n_123),
.B1(n_112),
.B2(n_124),
.C1(n_125),
.C2(n_133),
.Y(n_191)
);

AOI21xp5_ASAP7_75t_SL g194 ( 
.A1(n_191),
.A2(n_192),
.B(n_187),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_L g195 ( 
.A1(n_194),
.A2(n_186),
.B(n_122),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g196 ( 
.A(n_195),
.B(n_193),
.Y(n_196)
);


endmodule