module fake_jpeg_12463_n_159 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_159);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_159;

wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_93;
wire n_91;
wire n_54;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx11_ASAP7_75t_L g48 ( 
.A(n_36),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_9),
.Y(n_49)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_42),
.Y(n_50)
);

BUFx12_ASAP7_75t_L g51 ( 
.A(n_14),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_0),
.B(n_34),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_38),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_29),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_45),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_44),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_47),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_40),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_41),
.B(n_33),
.Y(n_59)
);

BUFx10_ASAP7_75t_L g60 ( 
.A(n_2),
.Y(n_60)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_11),
.Y(n_61)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_11),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_3),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_12),
.B(n_7),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_27),
.Y(n_65)
);

BUFx5_ASAP7_75t_L g66 ( 
.A(n_31),
.Y(n_66)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_8),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_32),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_21),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_L g70 ( 
.A1(n_62),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_70)
);

OA22x2_ASAP7_75t_L g83 ( 
.A1(n_70),
.A2(n_67),
.B1(n_60),
.B2(n_49),
.Y(n_83)
);

INVx5_ASAP7_75t_L g71 ( 
.A(n_48),
.Y(n_71)
);

INVx5_ASAP7_75t_L g85 ( 
.A(n_71),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_52),
.B(n_19),
.Y(n_72)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_72),
.B(n_59),
.C(n_60),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_56),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_73),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_48),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_74),
.B(n_75),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_63),
.B(n_1),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_51),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_76),
.B(n_79),
.Y(n_87)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_66),
.Y(n_77)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_77),
.Y(n_84)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_66),
.Y(n_78)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_78),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_64),
.B(n_3),
.Y(n_79)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_73),
.Y(n_80)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_80),
.Y(n_107)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_73),
.Y(n_81)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_81),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_72),
.A2(n_67),
.B1(n_62),
.B2(n_61),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_82),
.A2(n_49),
.B1(n_60),
.B2(n_50),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_83),
.B(n_93),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_76),
.B(n_57),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_SL g106 ( 
.A(n_88),
.B(n_92),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_91),
.B(n_94),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_74),
.B(n_55),
.Y(n_92)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_71),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_77),
.B(n_58),
.Y(n_94)
);

OR2x2_ASAP7_75t_L g96 ( 
.A(n_84),
.B(n_78),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_96),
.B(n_100),
.Y(n_128)
);

HB1xp67_ASAP7_75t_L g97 ( 
.A(n_84),
.Y(n_97)
);

CKINVDCx16_ASAP7_75t_R g121 ( 
.A(n_97),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_86),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_98),
.B(n_101),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_87),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_SL g102 ( 
.A1(n_83),
.A2(n_69),
.B(n_68),
.Y(n_102)
);

AOI21xp5_ASAP7_75t_L g117 ( 
.A1(n_102),
.A2(n_114),
.B(n_5),
.Y(n_117)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_89),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_103),
.B(n_107),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_89),
.A2(n_50),
.B1(n_56),
.B2(n_53),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_104),
.A2(n_109),
.B1(n_9),
.B2(n_10),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_80),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_105),
.B(n_24),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_83),
.B(n_54),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_SL g119 ( 
.A(n_108),
.B(n_110),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_90),
.A2(n_65),
.B1(n_51),
.B2(n_6),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_85),
.B(n_4),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_90),
.B(n_51),
.C(n_22),
.Y(n_112)
);

XOR2x2_ASAP7_75t_L g132 ( 
.A(n_112),
.B(n_13),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_85),
.B(n_4),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_SL g120 ( 
.A(n_113),
.B(n_5),
.Y(n_120)
);

AOI21xp5_ASAP7_75t_L g114 ( 
.A1(n_84),
.A2(n_20),
.B(n_43),
.Y(n_114)
);

OAI32xp33_ASAP7_75t_L g115 ( 
.A1(n_99),
.A2(n_18),
.A3(n_39),
.B1(n_37),
.B2(n_35),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_115),
.B(n_120),
.Y(n_135)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_95),
.Y(n_116)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_116),
.Y(n_146)
);

AOI21xp5_ASAP7_75t_L g138 ( 
.A1(n_117),
.A2(n_126),
.B(n_106),
.Y(n_138)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_95),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_118),
.B(n_124),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_102),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_122),
.A2(n_133),
.B1(n_26),
.B2(n_28),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_111),
.B(n_46),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_125),
.B(n_127),
.Y(n_145)
);

NAND2x1_ASAP7_75t_SL g126 ( 
.A(n_96),
.B(n_10),
.Y(n_126)
);

XNOR2xp5_ASAP7_75t_L g136 ( 
.A(n_129),
.B(n_130),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_114),
.B(n_30),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_100),
.B(n_12),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_131),
.B(n_132),
.C(n_134),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_109),
.A2(n_13),
.B1(n_15),
.B2(n_16),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_107),
.B(n_17),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_121),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_137),
.B(n_143),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_L g151 ( 
.A1(n_138),
.A2(n_126),
.B(n_119),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_124),
.B(n_112),
.C(n_103),
.Y(n_141)
);

XOR2xp5_ASAP7_75t_L g148 ( 
.A(n_141),
.B(n_142),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_123),
.B(n_23),
.C(n_25),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_132),
.B(n_117),
.C(n_130),
.Y(n_143)
);

OR2x2_ASAP7_75t_L g150 ( 
.A(n_144),
.B(n_122),
.Y(n_150)
);

BUFx24_ASAP7_75t_SL g149 ( 
.A(n_136),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_149),
.B(n_150),
.Y(n_154)
);

AO221x1_ASAP7_75t_L g153 ( 
.A1(n_151),
.A2(n_135),
.B1(n_139),
.B2(n_146),
.C(n_115),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_147),
.A2(n_145),
.B1(n_128),
.B2(n_140),
.Y(n_152)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_152),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_155),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_156),
.Y(n_157)
);

AOI322xp5_ASAP7_75t_L g158 ( 
.A1(n_157),
.A2(n_135),
.A3(n_153),
.B1(n_152),
.B2(n_154),
.C1(n_137),
.C2(n_134),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_L g159 ( 
.A(n_158),
.B(n_148),
.Y(n_159)
);


endmodule