module fake_netlist_6_3203_n_112 (n_16, n_1, n_9, n_8, n_18, n_10, n_6, n_15, n_3, n_14, n_0, n_4, n_13, n_11, n_17, n_12, n_7, n_2, n_5, n_19, n_112);

input n_16;
input n_1;
input n_9;
input n_8;
input n_18;
input n_10;
input n_6;
input n_15;
input n_3;
input n_14;
input n_0;
input n_4;
input n_13;
input n_11;
input n_17;
input n_12;
input n_7;
input n_2;
input n_5;
input n_19;

output n_112;

wire n_52;
wire n_91;
wire n_46;
wire n_21;
wire n_88;
wire n_98;
wire n_39;
wire n_63;
wire n_73;
wire n_22;
wire n_68;
wire n_28;
wire n_50;
wire n_49;
wire n_83;
wire n_101;
wire n_77;
wire n_106;
wire n_92;
wire n_42;
wire n_96;
wire n_90;
wire n_24;
wire n_105;
wire n_54;
wire n_102;
wire n_87;
wire n_32;
wire n_66;
wire n_85;
wire n_99;
wire n_78;
wire n_84;
wire n_100;
wire n_23;
wire n_20;
wire n_47;
wire n_62;
wire n_29;
wire n_75;
wire n_109;
wire n_45;
wire n_34;
wire n_70;
wire n_67;
wire n_37;
wire n_33;
wire n_82;
wire n_27;
wire n_38;
wire n_110;
wire n_61;
wire n_81;
wire n_59;
wire n_76;
wire n_36;
wire n_26;
wire n_55;
wire n_94;
wire n_97;
wire n_108;
wire n_58;
wire n_64;
wire n_48;
wire n_65;
wire n_25;
wire n_40;
wire n_93;
wire n_80;
wire n_41;
wire n_86;
wire n_104;
wire n_95;
wire n_107;
wire n_71;
wire n_74;
wire n_72;
wire n_89;
wire n_103;
wire n_111;
wire n_60;
wire n_35;
wire n_69;
wire n_30;
wire n_79;
wire n_43;
wire n_31;
wire n_57;
wire n_53;
wire n_51;
wire n_44;
wire n_56;

INVxp33_ASAP7_75t_SL g20 ( 
.A(n_12),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_10),
.Y(n_21)
);

CKINVDCx5p33_ASAP7_75t_R g22 ( 
.A(n_8),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_17),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_15),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

CKINVDCx5p33_ASAP7_75t_R g26 ( 
.A(n_9),
.Y(n_26)
);

INVxp67_ASAP7_75t_SL g27 ( 
.A(n_18),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

CKINVDCx16_ASAP7_75t_R g29 ( 
.A(n_3),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_4),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

CKINVDCx16_ASAP7_75t_R g33 ( 
.A(n_3),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_11),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_14),
.Y(n_35)
);

CKINVDCx5p33_ASAP7_75t_R g36 ( 
.A(n_29),
.Y(n_36)
);

CKINVDCx5p33_ASAP7_75t_R g37 ( 
.A(n_33),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_21),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_25),
.Y(n_39)
);

CKINVDCx5p33_ASAP7_75t_R g40 ( 
.A(n_21),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_30),
.Y(n_41)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_23),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_28),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_32),
.Y(n_44)
);

NOR2x1p5_ASAP7_75t_L g45 ( 
.A(n_23),
.B(n_0),
.Y(n_45)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_24),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g47 ( 
.A(n_20),
.B(n_1),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_22),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_43),
.B(n_26),
.Y(n_49)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_46),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g51 ( 
.A1(n_36),
.A2(n_31),
.B1(n_27),
.B2(n_35),
.Y(n_51)
);

BUFx8_ASAP7_75t_L g52 ( 
.A(n_39),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_41),
.Y(n_53)
);

INVx2_ASAP7_75t_SL g54 ( 
.A(n_36),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_44),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_44),
.Y(n_56)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_46),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_50),
.Y(n_58)
);

AND2x2_ASAP7_75t_L g59 ( 
.A(n_55),
.B(n_43),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_49),
.B(n_46),
.Y(n_60)
);

OR2x6_ASAP7_75t_L g61 ( 
.A(n_54),
.B(n_45),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_53),
.Y(n_62)
);

AOI21xp5_ASAP7_75t_L g63 ( 
.A1(n_49),
.A2(n_57),
.B(n_50),
.Y(n_63)
);

AOI21xp5_ASAP7_75t_L g64 ( 
.A1(n_60),
.A2(n_57),
.B(n_47),
.Y(n_64)
);

OAI21x1_ASAP7_75t_L g65 ( 
.A1(n_63),
.A2(n_42),
.B(n_34),
.Y(n_65)
);

OA21x2_ASAP7_75t_L g66 ( 
.A1(n_62),
.A2(n_56),
.B(n_51),
.Y(n_66)
);

OAI21x1_ASAP7_75t_L g67 ( 
.A1(n_59),
.A2(n_42),
.B(n_24),
.Y(n_67)
);

OAI21x1_ASAP7_75t_L g68 ( 
.A1(n_59),
.A2(n_42),
.B(n_24),
.Y(n_68)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_58),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_69),
.B(n_58),
.Y(n_70)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_69),
.Y(n_71)
);

INVx5_ASAP7_75t_SL g72 ( 
.A(n_66),
.Y(n_72)
);

NAND2xp33_ASAP7_75t_R g73 ( 
.A(n_66),
.B(n_40),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_67),
.Y(n_74)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_71),
.B(n_61),
.Y(n_75)
);

OA21x2_ASAP7_75t_L g76 ( 
.A1(n_70),
.A2(n_65),
.B(n_68),
.Y(n_76)
);

BUFx3_ASAP7_75t_L g77 ( 
.A(n_74),
.Y(n_77)
);

OAI21x1_ASAP7_75t_L g78 ( 
.A1(n_72),
.A2(n_64),
.B(n_24),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_72),
.Y(n_79)
);

OR2x2_ASAP7_75t_L g80 ( 
.A(n_75),
.B(n_40),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_75),
.Y(n_81)
);

NOR2xp67_ASAP7_75t_L g82 ( 
.A(n_79),
.B(n_64),
.Y(n_82)
);

AND2x2_ASAP7_75t_L g83 ( 
.A(n_79),
.B(n_61),
.Y(n_83)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_82),
.Y(n_84)
);

INVx1_ASAP7_75t_SL g85 ( 
.A(n_80),
.Y(n_85)
);

NOR2xp67_ASAP7_75t_L g86 ( 
.A(n_81),
.B(n_77),
.Y(n_86)
);

HB1xp67_ASAP7_75t_L g87 ( 
.A(n_83),
.Y(n_87)
);

INVx1_ASAP7_75t_SL g88 ( 
.A(n_83),
.Y(n_88)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_81),
.Y(n_89)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_89),
.Y(n_90)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_87),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_88),
.B(n_38),
.Y(n_92)
);

AND2x2_ASAP7_75t_L g93 ( 
.A(n_84),
.B(n_78),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_91),
.B(n_85),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_92),
.B(n_48),
.Y(n_95)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_90),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_93),
.B(n_37),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_93),
.B(n_37),
.Y(n_98)
);

NAND4xp25_ASAP7_75t_SL g99 ( 
.A(n_94),
.B(n_84),
.C(n_73),
.D(n_1),
.Y(n_99)
);

AOI221xp5_ASAP7_75t_L g100 ( 
.A1(n_97),
.A2(n_4),
.B1(n_61),
.B2(n_77),
.C(n_52),
.Y(n_100)
);

OAI21xp33_ASAP7_75t_L g101 ( 
.A1(n_98),
.A2(n_86),
.B(n_78),
.Y(n_101)
);

A2O1A1Ixp33_ASAP7_75t_L g102 ( 
.A1(n_95),
.A2(n_78),
.B(n_77),
.C(n_52),
.Y(n_102)
);

NOR2x1p5_ASAP7_75t_L g103 ( 
.A(n_99),
.B(n_96),
.Y(n_103)
);

AOI21xp33_ASAP7_75t_L g104 ( 
.A1(n_101),
.A2(n_76),
.B(n_7),
.Y(n_104)
);

OR2x2_ASAP7_75t_L g105 ( 
.A(n_102),
.B(n_76),
.Y(n_105)
);

HB1xp67_ASAP7_75t_L g106 ( 
.A(n_105),
.Y(n_106)
);

CKINVDCx5p33_ASAP7_75t_R g107 ( 
.A(n_103),
.Y(n_107)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_106),
.Y(n_108)
);

AOI21xp5_ASAP7_75t_L g109 ( 
.A1(n_108),
.A2(n_107),
.B(n_100),
.Y(n_109)
);

AND3x1_ASAP7_75t_L g110 ( 
.A(n_109),
.B(n_104),
.C(n_13),
.Y(n_110)
);

AOI222xp33_ASAP7_75t_L g111 ( 
.A1(n_110),
.A2(n_5),
.B1(n_16),
.B2(n_19),
.C1(n_74),
.C2(n_76),
.Y(n_111)
);

AOI21xp5_ASAP7_75t_L g112 ( 
.A1(n_111),
.A2(n_76),
.B(n_74),
.Y(n_112)
);


endmodule