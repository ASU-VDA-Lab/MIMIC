module fake_jpeg_9294_n_108 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_108);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_108;

wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_49;
wire n_76;
wire n_88;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_81;
wire n_106;
wire n_44;
wire n_75;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_93;
wire n_91;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_62;
wire n_43;
wire n_100;
wire n_82;
wire n_96;

INVx5_ASAP7_75t_L g43 ( 
.A(n_40),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_29),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_15),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_42),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_34),
.Y(n_47)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_5),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_23),
.Y(n_49)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_19),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_2),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_4),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_16),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_20),
.B(n_24),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_33),
.Y(n_56)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_37),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_27),
.Y(n_58)
);

BUFx10_ASAP7_75t_L g59 ( 
.A(n_39),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_8),
.Y(n_60)
);

BUFx5_ASAP7_75t_L g61 ( 
.A(n_6),
.Y(n_61)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_41),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_26),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_7),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_50),
.Y(n_65)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_65),
.Y(n_77)
);

BUFx5_ASAP7_75t_L g66 ( 
.A(n_61),
.Y(n_66)
);

BUFx2_ASAP7_75t_L g82 ( 
.A(n_66),
.Y(n_82)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_59),
.Y(n_67)
);

INVx2_ASAP7_75t_SL g76 ( 
.A(n_67),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_44),
.Y(n_68)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_68),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_45),
.B(n_0),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_69),
.B(n_70),
.Y(n_86)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_43),
.Y(n_70)
);

INVx8_ASAP7_75t_L g71 ( 
.A(n_57),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_71),
.A2(n_75),
.B1(n_58),
.B2(n_53),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_51),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_72),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_52),
.Y(n_73)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_73),
.Y(n_84)
);

BUFx3_ASAP7_75t_L g74 ( 
.A(n_63),
.Y(n_74)
);

INVx1_ASAP7_75t_SL g85 ( 
.A(n_74),
.Y(n_85)
);

INVx6_ASAP7_75t_L g75 ( 
.A(n_48),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_75),
.A2(n_62),
.B1(n_64),
.B2(n_54),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_79),
.A2(n_46),
.B1(n_3),
.B2(n_9),
.Y(n_90)
);

BUFx2_ASAP7_75t_L g91 ( 
.A(n_80),
.Y(n_91)
);

AOI21xp33_ASAP7_75t_L g83 ( 
.A1(n_69),
.A2(n_55),
.B(n_56),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_83),
.A2(n_60),
.B1(n_49),
.B2(n_47),
.Y(n_88)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_66),
.Y(n_87)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_87),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_88),
.B(n_89),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_81),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_90),
.A2(n_93),
.B1(n_78),
.B2(n_84),
.Y(n_94)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_77),
.Y(n_93)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_94),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_96),
.B(n_95),
.C(n_86),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_97),
.B(n_91),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_98),
.B(n_85),
.C(n_92),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_99),
.A2(n_82),
.B1(n_76),
.B2(n_11),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_100),
.B(n_1),
.C(n_10),
.Y(n_101)
);

AOI21xp5_ASAP7_75t_L g102 ( 
.A1(n_101),
.A2(n_12),
.B(n_13),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_102),
.B(n_14),
.Y(n_103)
);

A2O1A1O1Ixp25_ASAP7_75t_L g104 ( 
.A1(n_103),
.A2(n_17),
.B(n_18),
.C(n_21),
.D(n_22),
.Y(n_104)
);

XOR2xp5_ASAP7_75t_L g105 ( 
.A(n_104),
.B(n_25),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_105),
.B(n_28),
.C(n_30),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_106),
.B(n_31),
.C(n_32),
.Y(n_107)
);

AOI21xp5_ASAP7_75t_L g108 ( 
.A1(n_107),
.A2(n_35),
.B(n_36),
.Y(n_108)
);


endmodule