module fake_jpeg_2812_n_118 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_118);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_118;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_1),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_2),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_6),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_5),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_9),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

BUFx10_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

BUFx16f_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_0),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_4),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

BUFx2_ASAP7_75t_L g26 ( 
.A(n_20),
.Y(n_26)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_26),
.Y(n_44)
);

INVx5_ASAP7_75t_L g27 ( 
.A(n_24),
.Y(n_27)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_27),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_20),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_28),
.Y(n_37)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_19),
.Y(n_29)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_29),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_20),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_30),
.Y(n_43)
);

INVx1_ASAP7_75t_SL g31 ( 
.A(n_24),
.Y(n_31)
);

BUFx16f_ASAP7_75t_L g46 ( 
.A(n_31),
.Y(n_46)
);

INVx11_ASAP7_75t_L g32 ( 
.A(n_24),
.Y(n_32)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_32),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_24),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_SL g39 ( 
.A(n_33),
.B(n_22),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_16),
.B(n_4),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_SL g35 ( 
.A(n_34),
.B(n_23),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_35),
.B(n_41),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g36 ( 
.A1(n_31),
.A2(n_13),
.B1(n_21),
.B2(n_12),
.Y(n_36)
);

CKINVDCx16_ASAP7_75t_R g57 ( 
.A(n_36),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g38 ( 
.A1(n_29),
.A2(n_19),
.B1(n_17),
.B2(n_14),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_38),
.B(n_42),
.Y(n_49)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_39),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_SL g41 ( 
.A1(n_31),
.A2(n_13),
.B1(n_21),
.B2(n_12),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_34),
.B(n_25),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_46),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_50),
.B(n_54),
.Y(n_62)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_45),
.Y(n_51)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_51),
.Y(n_70)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_45),
.Y(n_53)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_53),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_46),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_46),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_55),
.B(n_28),
.Y(n_66)
);

MAJIxp5_ASAP7_75t_L g56 ( 
.A(n_38),
.B(n_26),
.C(n_44),
.Y(n_56)
);

XOR2xp5_ASAP7_75t_L g72 ( 
.A(n_56),
.B(n_32),
.Y(n_72)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_44),
.Y(n_58)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_58),
.Y(n_63)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_47),
.Y(n_59)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_59),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_42),
.B(n_25),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_60),
.B(n_35),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_61),
.B(n_65),
.Y(n_76)
);

OAI21xp5_ASAP7_75t_L g64 ( 
.A1(n_48),
.A2(n_26),
.B(n_40),
.Y(n_64)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_64),
.B(n_54),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_52),
.B(n_15),
.Y(n_65)
);

CKINVDCx16_ASAP7_75t_R g78 ( 
.A(n_66),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_52),
.B(n_15),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_67),
.B(n_60),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_57),
.A2(n_32),
.B1(n_40),
.B2(n_28),
.Y(n_68)
);

INVxp67_ASAP7_75t_L g79 ( 
.A(n_68),
.Y(n_79)
);

XNOR2xp5_ASAP7_75t_L g84 ( 
.A(n_72),
.B(n_59),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_49),
.A2(n_33),
.B1(n_27),
.B2(n_14),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_73),
.A2(n_49),
.B1(n_47),
.B2(n_33),
.Y(n_74)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_74),
.Y(n_89)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_69),
.Y(n_75)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_75),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_77),
.B(n_80),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_72),
.A2(n_56),
.B1(n_53),
.B2(n_51),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_SL g93 ( 
.A(n_81),
.B(n_83),
.Y(n_93)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_71),
.Y(n_82)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_82),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_61),
.B(n_58),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_84),
.B(n_64),
.C(n_67),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_77),
.Y(n_85)
);

OAI21xp5_ASAP7_75t_L g94 ( 
.A1(n_85),
.A2(n_86),
.B(n_80),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_77),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_87),
.B(n_78),
.C(n_84),
.Y(n_95)
);

AOI322xp5_ASAP7_75t_L g90 ( 
.A1(n_76),
.A2(n_65),
.A3(n_18),
.B1(n_73),
.B2(n_17),
.C1(n_62),
.C2(n_70),
.Y(n_90)
);

AOI322xp5_ASAP7_75t_L g100 ( 
.A1(n_90),
.A2(n_89),
.A3(n_91),
.B1(n_86),
.B2(n_18),
.C1(n_93),
.C2(n_88),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_94),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_95),
.B(n_96),
.C(n_97),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_87),
.B(n_55),
.C(n_63),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_92),
.B(n_63),
.C(n_69),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_L g98 ( 
.A1(n_85),
.A2(n_79),
.B(n_74),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_98),
.A2(n_88),
.B1(n_37),
.B2(n_43),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_89),
.A2(n_79),
.B1(n_22),
.B2(n_43),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_99),
.A2(n_100),
.B1(n_37),
.B2(n_91),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_SL g106 ( 
.A1(n_103),
.A2(n_104),
.B(n_37),
.Y(n_106)
);

XOR2xp5_ASAP7_75t_L g105 ( 
.A(n_94),
.B(n_28),
.Y(n_105)
);

XOR2xp5_ASAP7_75t_L g109 ( 
.A(n_105),
.B(n_0),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_106),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_112)
);

AOI21x1_ASAP7_75t_L g107 ( 
.A1(n_101),
.A2(n_30),
.B(n_18),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_107),
.B(n_108),
.C(n_109),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_102),
.B(n_30),
.C(n_18),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_108),
.B(n_102),
.C(n_105),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_SL g113 ( 
.A(n_111),
.B(n_112),
.Y(n_113)
);

AOI21xp5_ASAP7_75t_SL g114 ( 
.A1(n_110),
.A2(n_6),
.B(n_7),
.Y(n_114)
);

AOI21xp5_ASAP7_75t_L g115 ( 
.A1(n_114),
.A2(n_8),
.B(n_10),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_SL g116 ( 
.A1(n_115),
.A2(n_113),
.B(n_2),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_116),
.B(n_1),
.Y(n_117)
);

XOR2xp5_ASAP7_75t_L g118 ( 
.A(n_117),
.B(n_3),
.Y(n_118)
);


endmodule