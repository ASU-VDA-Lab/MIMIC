module real_aes_15895_n_4 (n_0, n_3, n_2, n_1, n_4);
input n_0;
input n_3;
input n_2;
input n_1;
output n_4;
wire n_5;
wire n_7;
wire n_8;
wire n_6;
wire n_9;
wire n_10;
wire n_11;
INVx1_ASAP7_75t_L g9 ( .A(n_0), .Y(n_9) );
HB1xp67_ASAP7_75t_L g5 ( .A(n_1), .Y(n_5) );
HB1xp67_ASAP7_75t_L g10 ( .A(n_2), .Y(n_10) );
NAND2xp5_ASAP7_75t_L g11 ( .A(n_3), .B(n_8), .Y(n_11) );
AOI22xp33_ASAP7_75t_L g4 ( .A1(n_5), .A2(n_6), .B1(n_10), .B2(n_11), .Y(n_4) );
NOR2xp33_ASAP7_75t_L g6 ( .A(n_7), .B(n_10), .Y(n_6) );
CKINVDCx16_ASAP7_75t_R g7 ( .A(n_8), .Y(n_7) );
HB1xp67_ASAP7_75t_L g8 ( .A(n_9), .Y(n_8) );
endmodule