module fake_jpeg_6667_n_317 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_317);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_317;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_137;
wire n_74;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g15 ( 
.A(n_9),
.Y(n_15)
);

BUFx3_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_7),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

INVx3_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_3),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_31),
.B(n_33),
.Y(n_46)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_22),
.Y(n_32)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_32),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_19),
.B(n_14),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_17),
.B(n_0),
.Y(n_34)
);

AND2x2_ASAP7_75t_L g51 ( 
.A(n_34),
.B(n_24),
.Y(n_51)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_22),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_35),
.B(n_36),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_19),
.B(n_14),
.Y(n_36)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_22),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_37),
.B(n_38),
.Y(n_63)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_25),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_16),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_39),
.B(n_26),
.Y(n_42)
);

INVx5_ASAP7_75t_L g40 ( 
.A(n_30),
.Y(n_40)
);

INVx5_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_19),
.B(n_14),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_41),
.B(n_13),
.Y(n_58)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_42),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g43 ( 
.A1(n_31),
.A2(n_24),
.B1(n_17),
.B2(n_30),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_43),
.A2(n_41),
.B1(n_15),
.B2(n_37),
.Y(n_73)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_40),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_44),
.B(n_47),
.Y(n_80)
);

OAI21xp33_ASAP7_75t_L g45 ( 
.A1(n_34),
.A2(n_30),
.B(n_25),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_45),
.A2(n_29),
.B1(n_28),
.B2(n_27),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_34),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_33),
.Y(n_48)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_48),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_33),
.B(n_21),
.Y(n_49)
);

MAJIxp5_ASAP7_75t_L g69 ( 
.A(n_49),
.B(n_41),
.C(n_36),
.Y(n_69)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_40),
.Y(n_50)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_50),
.Y(n_75)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_51),
.Y(n_84)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_40),
.Y(n_52)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_52),
.Y(n_86)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_32),
.Y(n_54)
);

INVxp67_ASAP7_75t_L g79 ( 
.A(n_54),
.Y(n_79)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_36),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_55),
.A2(n_65),
.B1(n_35),
.B2(n_38),
.Y(n_66)
);

BUFx12f_ASAP7_75t_L g56 ( 
.A(n_32),
.Y(n_56)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_56),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_58),
.A2(n_37),
.B1(n_39),
.B2(n_12),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_L g59 ( 
.A1(n_31),
.A2(n_21),
.B1(n_18),
.B2(n_20),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_L g72 ( 
.A1(n_59),
.A2(n_15),
.B1(n_31),
.B2(n_38),
.Y(n_72)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_39),
.Y(n_60)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_60),
.Y(n_68)
);

INVx4_ASAP7_75t_SL g61 ( 
.A(n_32),
.Y(n_61)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_61),
.Y(n_87)
);

BUFx5_ASAP7_75t_L g64 ( 
.A(n_32),
.Y(n_64)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_64),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_35),
.A2(n_25),
.B1(n_18),
.B2(n_20),
.Y(n_65)
);

AOI21xp5_ASAP7_75t_L g95 ( 
.A1(n_66),
.A2(n_77),
.B(n_83),
.Y(n_95)
);

AND2x2_ASAP7_75t_L g107 ( 
.A(n_69),
.B(n_49),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_48),
.A2(n_38),
.B1(n_37),
.B2(n_35),
.Y(n_70)
);

INVxp67_ASAP7_75t_L g92 ( 
.A(n_70),
.Y(n_92)
);

CKINVDCx16_ASAP7_75t_R g94 ( 
.A(n_72),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_L g104 ( 
.A1(n_73),
.A2(n_82),
.B1(n_88),
.B2(n_50),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_76),
.B(n_11),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_47),
.A2(n_28),
.B1(n_27),
.B2(n_23),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_78),
.A2(n_81),
.B1(n_85),
.B2(n_53),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_43),
.A2(n_28),
.B1(n_27),
.B2(n_23),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_L g82 ( 
.A1(n_55),
.A2(n_23),
.B1(n_26),
.B2(n_16),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_44),
.A2(n_32),
.B1(n_13),
.B2(n_12),
.Y(n_83)
);

OA22x2_ASAP7_75t_L g85 ( 
.A1(n_61),
.A2(n_32),
.B1(n_29),
.B2(n_26),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_L g88 ( 
.A1(n_52),
.A2(n_29),
.B1(n_1),
.B2(n_2),
.Y(n_88)
);

CKINVDCx14_ASAP7_75t_R g90 ( 
.A(n_80),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_90),
.B(n_93),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_91),
.A2(n_109),
.B1(n_104),
.B2(n_94),
.Y(n_118)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_80),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_78),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_96),
.B(n_97),
.Y(n_137)
);

HB1xp67_ASAP7_75t_L g97 ( 
.A(n_85),
.Y(n_97)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_73),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_98),
.B(n_99),
.Y(n_122)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_72),
.Y(n_99)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_82),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_100),
.B(n_102),
.Y(n_134)
);

O2A1O1Ixp33_ASAP7_75t_SL g101 ( 
.A1(n_85),
.A2(n_61),
.B(n_53),
.C(n_64),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_101),
.A2(n_62),
.B1(n_68),
.B2(n_75),
.Y(n_141)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_70),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_85),
.Y(n_103)
);

INVxp67_ASAP7_75t_SL g130 ( 
.A(n_103),
.Y(n_130)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_104),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_71),
.B(n_51),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_105),
.B(n_108),
.Y(n_123)
);

INVx1_ASAP7_75t_SL g106 ( 
.A(n_85),
.Y(n_106)
);

AND2x2_ASAP7_75t_L g128 ( 
.A(n_106),
.B(n_87),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_107),
.A2(n_111),
.B1(n_110),
.B2(n_90),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_71),
.B(n_51),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_88),
.Y(n_109)
);

AO21x1_ASAP7_75t_L g139 ( 
.A1(n_109),
.A2(n_112),
.B(n_63),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_84),
.B(n_46),
.Y(n_110)
);

XNOR2xp5_ASAP7_75t_L g121 ( 
.A(n_110),
.B(n_105),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_84),
.B(n_46),
.Y(n_111)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_111),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_67),
.B(n_57),
.Y(n_113)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_113),
.Y(n_131)
);

CKINVDCx16_ASAP7_75t_R g114 ( 
.A(n_83),
.Y(n_114)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_114),
.Y(n_135)
);

OAI21xp33_ASAP7_75t_L g115 ( 
.A1(n_111),
.A2(n_77),
.B(n_57),
.Y(n_115)
);

XNOR2xp5_ASAP7_75t_L g163 ( 
.A(n_115),
.B(n_121),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_SL g146 ( 
.A(n_116),
.B(n_126),
.Y(n_146)
);

BUFx5_ASAP7_75t_L g117 ( 
.A(n_92),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_117),
.B(n_127),
.Y(n_158)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_118),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_98),
.A2(n_81),
.B1(n_66),
.B2(n_60),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_119),
.A2(n_124),
.B1(n_129),
.B2(n_141),
.Y(n_167)
);

AO22x1_ASAP7_75t_L g124 ( 
.A1(n_97),
.A2(n_62),
.B1(n_87),
.B2(n_68),
.Y(n_124)
);

NAND2xp33_ASAP7_75t_R g126 ( 
.A(n_93),
.B(n_63),
.Y(n_126)
);

BUFx12_ASAP7_75t_L g127 ( 
.A(n_101),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_128),
.B(n_138),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_95),
.A2(n_67),
.B1(n_86),
.B2(n_62),
.Y(n_129)
);

AND2x2_ASAP7_75t_L g133 ( 
.A(n_108),
.B(n_69),
.Y(n_133)
);

AND2x2_ASAP7_75t_L g145 ( 
.A(n_133),
.B(n_136),
.Y(n_145)
);

AND2x2_ASAP7_75t_L g136 ( 
.A(n_106),
.B(n_107),
.Y(n_136)
);

INVxp67_ASAP7_75t_L g138 ( 
.A(n_95),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_139),
.B(n_103),
.Y(n_166)
);

AOI21xp5_ASAP7_75t_L g140 ( 
.A1(n_95),
.A2(n_75),
.B(n_86),
.Y(n_140)
);

XOR2xp5_ASAP7_75t_L g151 ( 
.A(n_140),
.B(n_91),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_125),
.B(n_107),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_142),
.B(n_147),
.Y(n_178)
);

OR2x2_ASAP7_75t_L g143 ( 
.A(n_124),
.B(n_96),
.Y(n_143)
);

AND2x2_ASAP7_75t_L g186 ( 
.A(n_143),
.B(n_151),
.Y(n_186)
);

BUFx24_ASAP7_75t_SL g144 ( 
.A(n_121),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_144),
.B(n_159),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_125),
.B(n_107),
.Y(n_147)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_137),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_149),
.B(n_156),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_116),
.B(n_113),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_150),
.B(n_152),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_133),
.B(n_136),
.Y(n_152)
);

AND2x2_ASAP7_75t_L g153 ( 
.A(n_136),
.B(n_106),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_L g179 ( 
.A1(n_153),
.A2(n_164),
.B(n_122),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_133),
.B(n_102),
.Y(n_154)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_154),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_123),
.B(n_131),
.Y(n_155)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_155),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_SL g156 ( 
.A(n_131),
.B(n_94),
.Y(n_156)
);

AND2x6_ASAP7_75t_L g157 ( 
.A(n_138),
.B(n_101),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_L g188 ( 
.A(n_157),
.B(n_58),
.Y(n_188)
);

CKINVDCx16_ASAP7_75t_R g159 ( 
.A(n_132),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_123),
.B(n_91),
.C(n_114),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_160),
.B(n_134),
.C(n_141),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_140),
.B(n_101),
.Y(n_161)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_161),
.Y(n_187)
);

AND2x2_ASAP7_75t_L g164 ( 
.A(n_127),
.B(n_103),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_124),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_165),
.Y(n_170)
);

AO21x1_ASAP7_75t_L g177 ( 
.A1(n_166),
.A2(n_158),
.B(n_162),
.Y(n_177)
);

AOI322xp5_ASAP7_75t_L g168 ( 
.A1(n_157),
.A2(n_129),
.A3(n_118),
.B1(n_120),
.B2(n_134),
.C1(n_128),
.C2(n_127),
.Y(n_168)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_168),
.B(n_173),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_148),
.A2(n_119),
.B1(n_120),
.B2(n_130),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_171),
.A2(n_179),
.B1(n_184),
.B2(n_153),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_148),
.A2(n_128),
.B1(n_127),
.B2(n_135),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_174),
.A2(n_176),
.B1(n_180),
.B2(n_68),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_167),
.A2(n_135),
.B1(n_99),
.B2(n_100),
.Y(n_176)
);

O2A1O1Ixp33_ASAP7_75t_L g196 ( 
.A1(n_177),
.A2(n_161),
.B(n_153),
.C(n_143),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_167),
.A2(n_117),
.B1(n_139),
.B2(n_103),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_155),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_181),
.Y(n_199)
);

CKINVDCx16_ASAP7_75t_R g182 ( 
.A(n_151),
.Y(n_182)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_182),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_SL g183 ( 
.A(n_152),
.B(n_139),
.Y(n_183)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_183),
.Y(n_209)
);

XNOR2x1_ASAP7_75t_SL g184 ( 
.A(n_145),
.B(n_112),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_154),
.B(n_54),
.C(n_56),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_185),
.B(n_190),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_L g200 ( 
.A1(n_188),
.A2(n_160),
.B1(n_163),
.B2(n_146),
.Y(n_200)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_150),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_142),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_191),
.B(n_193),
.Y(n_210)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_147),
.Y(n_193)
);

XOR2xp5_ASAP7_75t_L g194 ( 
.A(n_163),
.B(n_56),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_194),
.B(n_185),
.Y(n_211)
);

CKINVDCx14_ASAP7_75t_R g195 ( 
.A(n_176),
.Y(n_195)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_195),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_196),
.A2(n_204),
.B1(n_212),
.B2(n_215),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_197),
.A2(n_202),
.B1(n_187),
.B2(n_193),
.Y(n_226)
);

INVxp67_ASAP7_75t_L g198 ( 
.A(n_174),
.Y(n_198)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_198),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_200),
.B(n_173),
.Y(n_223)
);

AO22x1_ASAP7_75t_L g202 ( 
.A1(n_186),
.A2(n_164),
.B1(n_146),
.B2(n_145),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_170),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_SL g221 ( 
.A(n_203),
.B(n_213),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_L g204 ( 
.A1(n_180),
.A2(n_149),
.B1(n_164),
.B2(n_145),
.Y(n_204)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_178),
.Y(n_206)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_206),
.Y(n_233)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_178),
.Y(n_207)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_207),
.Y(n_234)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_189),
.Y(n_208)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_208),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_211),
.B(n_194),
.C(n_169),
.Y(n_224)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_172),
.Y(n_213)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_191),
.Y(n_214)
);

INVxp67_ASAP7_75t_L g237 ( 
.A(n_214),
.Y(n_237)
);

INVx1_ASAP7_75t_SL g215 ( 
.A(n_184),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_189),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_216),
.A2(n_218),
.B1(n_219),
.B2(n_175),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_187),
.A2(n_74),
.B1(n_89),
.B2(n_79),
.Y(n_218)
);

INVx5_ASAP7_75t_L g219 ( 
.A(n_188),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_223),
.B(n_226),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_224),
.B(n_225),
.C(n_209),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_201),
.B(n_169),
.C(n_183),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_219),
.B(n_186),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_227),
.B(n_228),
.Y(n_246)
);

XNOR2x1_ASAP7_75t_L g228 ( 
.A(n_202),
.B(n_186),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_211),
.B(n_179),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_229),
.B(n_230),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_197),
.B(n_171),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_198),
.A2(n_175),
.B1(n_177),
.B2(n_192),
.Y(n_232)
);

CKINVDCx16_ASAP7_75t_R g253 ( 
.A(n_232),
.Y(n_253)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_235),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_217),
.B(n_56),
.Y(n_236)
);

XOR2xp5_ASAP7_75t_L g248 ( 
.A(n_236),
.B(n_238),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_217),
.B(n_54),
.Y(n_238)
);

XOR2xp5_ASAP7_75t_L g239 ( 
.A(n_202),
.B(n_54),
.Y(n_239)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_239),
.B(n_218),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_L g241 ( 
.A1(n_231),
.A2(n_199),
.B1(n_214),
.B2(n_205),
.Y(n_241)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_241),
.Y(n_261)
);

OAI21xp5_ASAP7_75t_SL g242 ( 
.A1(n_220),
.A2(n_210),
.B(n_205),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_242),
.A2(n_243),
.B1(n_215),
.B2(n_236),
.Y(n_266)
);

OAI21xp5_ASAP7_75t_SL g243 ( 
.A1(n_228),
.A2(n_237),
.B(n_210),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_237),
.B(n_216),
.Y(n_244)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_244),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_249),
.B(n_254),
.C(n_258),
.Y(n_260)
);

INVx13_ASAP7_75t_L g250 ( 
.A(n_233),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_250),
.B(n_251),
.Y(n_263)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_221),
.Y(n_251)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_222),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_255),
.B(n_257),
.Y(n_271)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_239),
.Y(n_256)
);

AOI22xp33_ASAP7_75t_SL g262 ( 
.A1(n_256),
.A2(n_227),
.B1(n_196),
.B2(n_223),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_234),
.B(n_208),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_224),
.B(n_207),
.C(n_206),
.Y(n_258)
);

AOI21xp5_ASAP7_75t_L g259 ( 
.A1(n_240),
.A2(n_212),
.B(n_225),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_L g267 ( 
.A1(n_259),
.A2(n_238),
.B1(n_89),
.B2(n_13),
.Y(n_267)
);

OAI21xp33_ASAP7_75t_SL g284 ( 
.A1(n_262),
.A2(n_275),
.B(n_246),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_258),
.B(n_245),
.C(n_254),
.Y(n_264)
);

OAI21xp5_ASAP7_75t_L g280 ( 
.A1(n_264),
.A2(n_269),
.B(n_272),
.Y(n_280)
);

INVxp67_ASAP7_75t_SL g265 ( 
.A(n_243),
.Y(n_265)
);

OAI21x1_ASAP7_75t_L g276 ( 
.A1(n_265),
.A2(n_249),
.B(n_259),
.Y(n_276)
);

XOR2xp5_ASAP7_75t_L g285 ( 
.A(n_266),
.B(n_267),
.Y(n_285)
);

A2O1A1Ixp33_ASAP7_75t_L g268 ( 
.A1(n_253),
.A2(n_12),
.B(n_11),
.C(n_2),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_SL g283 ( 
.A(n_268),
.B(n_256),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_245),
.B(n_74),
.C(n_29),
.Y(n_269)
);

HB1xp67_ASAP7_75t_L g270 ( 
.A(n_242),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_270),
.B(n_250),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_244),
.B(n_74),
.C(n_29),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_252),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_SL g279 ( 
.A(n_274),
.B(n_11),
.Y(n_279)
);

AOI22xp33_ASAP7_75t_L g275 ( 
.A1(n_252),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_275)
);

AOI21xp5_ASAP7_75t_L g290 ( 
.A1(n_276),
.A2(n_277),
.B(n_284),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_273),
.B(n_247),
.Y(n_278)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_278),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_279),
.B(n_282),
.Y(n_289)
);

INVx3_ASAP7_75t_L g281 ( 
.A(n_272),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_SL g293 ( 
.A(n_281),
.B(n_269),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_273),
.B(n_247),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_SL g294 ( 
.A(n_283),
.B(n_287),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_261),
.B(n_246),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_286),
.B(n_288),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_274),
.B(n_248),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_263),
.B(n_248),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_280),
.B(n_264),
.C(n_260),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_291),
.B(n_293),
.C(n_4),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_285),
.B(n_271),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_295),
.B(n_296),
.C(n_297),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_285),
.B(n_268),
.Y(n_296)
);

XOR2xp5_ASAP7_75t_L g297 ( 
.A(n_284),
.B(n_266),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_281),
.B(n_260),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_L g305 ( 
.A(n_298),
.B(n_289),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_299),
.B(n_0),
.Y(n_300)
);

AOI21xp5_ASAP7_75t_L g312 ( 
.A1(n_300),
.A2(n_301),
.B(n_304),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_290),
.B(n_1),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_SL g302 ( 
.A1(n_294),
.A2(n_291),
.B1(n_292),
.B2(n_290),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_L g311 ( 
.A1(n_302),
.A2(n_6),
.B1(n_8),
.B2(n_9),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_SL g303 ( 
.A1(n_297),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_303),
.B(n_305),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_291),
.B(n_4),
.C(n_5),
.Y(n_306)
);

XOR2xp5_ASAP7_75t_L g309 ( 
.A(n_306),
.B(n_5),
.Y(n_309)
);

AOI21x1_ASAP7_75t_SL g308 ( 
.A1(n_304),
.A2(n_307),
.B(n_306),
.Y(n_308)
);

AOI21xp5_ASAP7_75t_SL g314 ( 
.A1(n_308),
.A2(n_6),
.B(n_8),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_309),
.B(n_311),
.C(n_6),
.Y(n_313)
);

OAI321xp33_ASAP7_75t_L g315 ( 
.A1(n_313),
.A2(n_314),
.A3(n_312),
.B1(n_10),
.B2(n_6),
.C(n_310),
.Y(n_315)
);

BUFx24_ASAP7_75t_SL g316 ( 
.A(n_315),
.Y(n_316)
);

XOR2xp5_ASAP7_75t_L g317 ( 
.A(n_316),
.B(n_310),
.Y(n_317)
);


endmodule