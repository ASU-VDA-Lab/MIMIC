module real_aes_1588_n_8 (n_4, n_0, n_3, n_5, n_2, n_7, n_6, n_1, n_8);
input n_4;
input n_0;
input n_3;
input n_5;
input n_2;
input n_7;
input n_6;
input n_1;
output n_8;
wire n_17;
wire n_22;
wire n_13;
wire n_24;
wire n_12;
wire n_19;
wire n_25;
wire n_14;
wire n_11;
wire n_16;
wire n_15;
wire n_23;
wire n_9;
wire n_20;
wire n_18;
wire n_26;
wire n_21;
wire n_10;
INVxp33_ASAP7_75t_L g17 ( .A(n_0), .Y(n_17) );
INVxp67_ASAP7_75t_L g16 ( .A(n_1), .Y(n_16) );
NAND3xp33_ASAP7_75t_SL g21 ( .A(n_2), .B(n_22), .C(n_23), .Y(n_21) );
INVx3_ASAP7_75t_L g25 ( .A(n_3), .Y(n_25) );
INVx1_ASAP7_75t_L g22 ( .A(n_4), .Y(n_22) );
INVx1_ASAP7_75t_L g10 ( .A(n_5), .Y(n_10) );
NOR2xp33_ASAP7_75t_L g26 ( .A(n_5), .B(n_11), .Y(n_26) );
AOI32xp33_ASAP7_75t_L g8 ( .A1(n_6), .A2(n_9), .A3(n_15), .B1(n_18), .B2(n_19), .Y(n_8) );
INVx1_ASAP7_75t_L g18 ( .A(n_6), .Y(n_18) );
INVx1_ASAP7_75t_L g14 ( .A(n_7), .Y(n_14) );
NOR2xp33_ASAP7_75t_L g9 ( .A(n_10), .B(n_11), .Y(n_9) );
OAI21xp33_ASAP7_75t_SL g19 ( .A1(n_11), .A2(n_15), .B(n_20), .Y(n_19) );
AOI21xp5_ASAP7_75t_SL g20 ( .A1(n_11), .A2(n_21), .B(n_26), .Y(n_20) );
CKINVDCx16_ASAP7_75t_R g11 ( .A(n_12), .Y(n_11) );
INVx1_ASAP7_75t_L g12 ( .A(n_13), .Y(n_12) );
HB1xp67_ASAP7_75t_L g13 ( .A(n_14), .Y(n_13) );
NOR2xp33_ASAP7_75t_L g15 ( .A(n_16), .B(n_17), .Y(n_15) );
INVx2_ASAP7_75t_L g23 ( .A(n_24), .Y(n_23) );
HB1xp67_ASAP7_75t_L g24 ( .A(n_25), .Y(n_24) );
endmodule