module fake_jpeg_25915_n_200 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_200);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_200;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g15 ( 
.A(n_14),
.Y(n_15)
);

BUFx5_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_8),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_8),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

INVx8_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_9),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_10),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_7),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

AOI22xp5_ASAP7_75t_L g32 ( 
.A1(n_26),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_SL g47 ( 
.A1(n_32),
.A2(n_19),
.B1(n_29),
.B2(n_28),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_26),
.B(n_0),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_33),
.B(n_35),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_30),
.Y(n_34)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_34),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_SL g35 ( 
.A(n_18),
.B(n_1),
.Y(n_35)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_30),
.Y(n_36)
);

HB1xp67_ASAP7_75t_L g49 ( 
.A(n_36),
.Y(n_49)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_30),
.Y(n_37)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_37),
.Y(n_57)
);

BUFx12_ASAP7_75t_L g38 ( 
.A(n_30),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_38),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_30),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_39),
.Y(n_52)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_21),
.Y(n_40)
);

OR2x2_ASAP7_75t_L g43 ( 
.A(n_40),
.B(n_41),
.Y(n_43)
);

CKINVDCx16_ASAP7_75t_R g41 ( 
.A(n_16),
.Y(n_41)
);

INVx5_ASAP7_75t_L g44 ( 
.A(n_34),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_44),
.B(n_39),
.Y(n_62)
);

INVx2_ASAP7_75t_SL g45 ( 
.A(n_34),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_45),
.B(n_54),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g46 ( 
.A1(n_33),
.A2(n_25),
.B1(n_22),
.B2(n_24),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_46),
.A2(n_47),
.B1(n_16),
.B2(n_23),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_36),
.A2(n_25),
.B1(n_29),
.B2(n_28),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_50),
.A2(n_51),
.B1(n_40),
.B2(n_17),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_37),
.A2(n_25),
.B1(n_27),
.B2(n_19),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_32),
.A2(n_27),
.B1(n_18),
.B2(n_24),
.Y(n_53)
);

OAI21xp5_ASAP7_75t_SL g73 ( 
.A1(n_53),
.A2(n_55),
.B(n_31),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_35),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_41),
.A2(n_17),
.B1(n_22),
.B2(n_20),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_58),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_90)
);

CKINVDCx16_ASAP7_75t_R g59 ( 
.A(n_49),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_59),
.B(n_60),
.Y(n_86)
);

OAI21xp33_ASAP7_75t_L g60 ( 
.A1(n_48),
.A2(n_31),
.B(n_20),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_49),
.Y(n_61)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_61),
.Y(n_94)
);

INVxp67_ASAP7_75t_L g80 ( 
.A(n_62),
.Y(n_80)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_57),
.Y(n_64)
);

BUFx24_ASAP7_75t_L g85 ( 
.A(n_64),
.Y(n_85)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_55),
.Y(n_65)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_65),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_48),
.B(n_54),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_66),
.B(n_75),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_47),
.B(n_15),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_SL g100 ( 
.A(n_67),
.B(n_68),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_46),
.B(n_15),
.Y(n_68)
);

INVxp67_ASAP7_75t_L g69 ( 
.A(n_56),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_69),
.B(n_72),
.Y(n_82)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_43),
.Y(n_70)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_70),
.Y(n_91)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_43),
.Y(n_71)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_71),
.Y(n_98)
);

CKINVDCx16_ASAP7_75t_R g72 ( 
.A(n_43),
.Y(n_72)
);

OAI21xp5_ASAP7_75t_L g97 ( 
.A1(n_73),
.A2(n_2),
.B(n_4),
.Y(n_97)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_52),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_74),
.B(n_79),
.Y(n_93)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_53),
.Y(n_75)
);

OA22x2_ASAP7_75t_L g76 ( 
.A1(n_42),
.A2(n_38),
.B1(n_39),
.B2(n_21),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_76),
.A2(n_45),
.B1(n_42),
.B2(n_44),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_57),
.B(n_38),
.C(n_21),
.Y(n_77)
);

XOR2xp5_ASAP7_75t_L g87 ( 
.A(n_77),
.B(n_45),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_78),
.A2(n_44),
.B1(n_23),
.B2(n_4),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_56),
.B(n_21),
.Y(n_79)
);

AOI21xp5_ASAP7_75t_L g81 ( 
.A1(n_65),
.A2(n_38),
.B(n_3),
.Y(n_81)
);

OAI21xp5_ASAP7_75t_SL g121 ( 
.A1(n_81),
.A2(n_90),
.B(n_76),
.Y(n_121)
);

AND2x2_ASAP7_75t_L g118 ( 
.A(n_83),
.B(n_87),
.Y(n_118)
);

AO21x2_ASAP7_75t_L g84 ( 
.A1(n_76),
.A2(n_42),
.B(n_45),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_84),
.A2(n_89),
.B1(n_92),
.B2(n_72),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_75),
.A2(n_52),
.B1(n_56),
.B2(n_5),
.Y(n_92)
);

INVxp67_ASAP7_75t_L g95 ( 
.A(n_63),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_95),
.B(n_76),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_L g106 ( 
.A1(n_97),
.A2(n_73),
.B(n_68),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_67),
.B(n_13),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_SL g115 ( 
.A(n_99),
.B(n_11),
.Y(n_115)
);

XOR2xp5_ASAP7_75t_L g101 ( 
.A(n_66),
.B(n_6),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_101),
.B(n_71),
.C(n_70),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_63),
.B(n_52),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_102),
.B(n_95),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_103),
.A2(n_84),
.B1(n_96),
.B2(n_80),
.Y(n_132)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_102),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_104),
.B(n_107),
.Y(n_124)
);

BUFx5_ASAP7_75t_L g105 ( 
.A(n_85),
.Y(n_105)
);

BUFx2_ASAP7_75t_L g130 ( 
.A(n_105),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_L g133 ( 
.A1(n_106),
.A2(n_121),
.B(n_97),
.Y(n_133)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_93),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_108),
.B(n_114),
.Y(n_131)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_85),
.Y(n_109)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_109),
.Y(n_127)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_88),
.Y(n_110)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_110),
.Y(n_129)
);

INVxp67_ASAP7_75t_L g111 ( 
.A(n_82),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_SL g141 ( 
.A1(n_111),
.A2(n_116),
.B(n_120),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_SL g135 ( 
.A(n_112),
.B(n_84),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_100),
.B(n_59),
.Y(n_113)
);

CKINVDCx16_ASAP7_75t_R g123 ( 
.A(n_113),
.Y(n_123)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_83),
.Y(n_114)
);

BUFx24_ASAP7_75t_SL g140 ( 
.A(n_115),
.Y(n_140)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_92),
.Y(n_116)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_84),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_117),
.B(n_119),
.Y(n_136)
);

AOI21xp5_ASAP7_75t_L g120 ( 
.A1(n_96),
.A2(n_61),
.B(n_78),
.Y(n_120)
);

BUFx4f_ASAP7_75t_SL g122 ( 
.A(n_85),
.Y(n_122)
);

CKINVDCx16_ASAP7_75t_R g126 ( 
.A(n_122),
.Y(n_126)
);

AOI21x1_ASAP7_75t_L g125 ( 
.A1(n_120),
.A2(n_84),
.B(n_81),
.Y(n_125)
);

INVxp67_ASAP7_75t_L g148 ( 
.A(n_125),
.Y(n_148)
);

CKINVDCx16_ASAP7_75t_R g128 ( 
.A(n_119),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_128),
.B(n_134),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_132),
.A2(n_137),
.B1(n_114),
.B2(n_116),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_SL g152 ( 
.A(n_133),
.B(n_138),
.Y(n_152)
);

CKINVDCx16_ASAP7_75t_R g134 ( 
.A(n_122),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_135),
.B(n_103),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_117),
.A2(n_89),
.B1(n_88),
.B2(n_87),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_L g138 ( 
.A1(n_118),
.A2(n_86),
.B(n_98),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_118),
.B(n_101),
.C(n_77),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_139),
.B(n_108),
.C(n_106),
.Y(n_144)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_130),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_142),
.B(n_143),
.Y(n_167)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_130),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_144),
.B(n_146),
.C(n_153),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_145),
.A2(n_94),
.B1(n_127),
.B2(n_64),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_139),
.B(n_118),
.C(n_104),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g147 ( 
.A(n_126),
.Y(n_147)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_147),
.Y(n_157)
);

MAJx2_ASAP7_75t_L g149 ( 
.A(n_131),
.B(n_133),
.C(n_141),
.Y(n_149)
);

MAJx2_ASAP7_75t_L g164 ( 
.A(n_149),
.B(n_129),
.C(n_91),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_124),
.Y(n_150)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_150),
.Y(n_165)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_124),
.Y(n_151)
);

AOI21xp5_ASAP7_75t_L g161 ( 
.A1(n_151),
.A2(n_136),
.B(n_141),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_131),
.B(n_107),
.C(n_121),
.Y(n_153)
);

FAx1_ASAP7_75t_SL g158 ( 
.A(n_155),
.B(n_132),
.CI(n_137),
.CON(n_158),
.SN(n_158)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_123),
.B(n_105),
.Y(n_156)
);

AOI322xp5_ASAP7_75t_L g163 ( 
.A1(n_156),
.A2(n_140),
.A3(n_122),
.B1(n_111),
.B2(n_80),
.C1(n_135),
.C2(n_127),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_158),
.B(n_161),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_148),
.A2(n_136),
.B1(n_153),
.B2(n_125),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_159),
.A2(n_166),
.B1(n_76),
.B2(n_74),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_146),
.B(n_138),
.C(n_129),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_162),
.B(n_109),
.C(n_52),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_163),
.B(n_168),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_L g171 ( 
.A(n_164),
.B(n_152),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_145),
.A2(n_148),
.B1(n_149),
.B2(n_154),
.Y(n_166)
);

AOI21xp5_ASAP7_75t_L g170 ( 
.A1(n_166),
.A2(n_152),
.B(n_147),
.Y(n_170)
);

XOR2xp5_ASAP7_75t_L g179 ( 
.A(n_170),
.B(n_171),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_165),
.B(n_94),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_173),
.B(n_176),
.Y(n_181)
);

XOR2xp5_ASAP7_75t_L g174 ( 
.A(n_160),
.B(n_144),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_174),
.B(n_175),
.C(n_159),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g177 ( 
.A(n_160),
.B(n_74),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_177),
.B(n_161),
.C(n_157),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_178),
.B(n_180),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_169),
.B(n_162),
.C(n_164),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_172),
.B(n_167),
.Y(n_182)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_182),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_175),
.B(n_168),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_183),
.A2(n_184),
.B1(n_181),
.B2(n_179),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_185),
.B(n_186),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_183),
.A2(n_171),
.B1(n_158),
.B2(n_177),
.Y(n_186)
);

NOR3xp33_ASAP7_75t_SL g189 ( 
.A(n_180),
.B(n_158),
.C(n_174),
.Y(n_189)
);

OR2x2_ASAP7_75t_L g193 ( 
.A(n_189),
.B(n_52),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_188),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_190),
.B(n_191),
.Y(n_195)
);

OAI21x1_ASAP7_75t_L g191 ( 
.A1(n_189),
.A2(n_12),
.B(n_7),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_193),
.B(n_186),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_194),
.B(n_187),
.C(n_192),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_196),
.B(n_197),
.C(n_6),
.Y(n_198)
);

HB1xp67_ASAP7_75t_L g197 ( 
.A(n_195),
.Y(n_197)
);

A2O1A1Ixp33_ASAP7_75t_L g199 ( 
.A1(n_198),
.A2(n_6),
.B(n_8),
.C(n_9),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_199),
.B(n_9),
.Y(n_200)
);


endmodule