module fake_jpeg_9675_n_176 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_176);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_176;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_175;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_12),
.Y(n_13)
);

BUFx12f_ASAP7_75t_L g14 ( 
.A(n_5),
.Y(n_14)
);

INVx6_ASAP7_75t_SL g15 ( 
.A(n_11),
.Y(n_15)
);

INVx3_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_8),
.B(n_0),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

INVx4_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_6),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_9),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

BUFx10_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_28),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_14),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_29),
.B(n_31),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

BUFx2_ASAP7_75t_L g39 ( 
.A(n_30),
.Y(n_39)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_20),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_14),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_SL g44 ( 
.A(n_32),
.B(n_33),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_17),
.B(n_0),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_23),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_34),
.B(n_27),
.Y(n_38)
);

INVx4_ASAP7_75t_SL g35 ( 
.A(n_27),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_SL g37 ( 
.A1(n_35),
.A2(n_20),
.B1(n_16),
.B2(n_24),
.Y(n_37)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_23),
.Y(n_36)
);

AND2x2_ASAP7_75t_L g40 ( 
.A(n_36),
.B(n_24),
.Y(n_40)
);

OAI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_37),
.A2(n_35),
.B1(n_31),
.B2(n_34),
.Y(n_48)
);

OAI21xp33_ASAP7_75t_L g65 ( 
.A1(n_38),
.A2(n_40),
.B(n_36),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_28),
.Y(n_41)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_41),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g42 ( 
.A1(n_35),
.A2(n_16),
.B1(n_18),
.B2(n_15),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_L g66 ( 
.A1(n_42),
.A2(n_46),
.B1(n_13),
.B2(n_26),
.Y(n_66)
);

BUFx12_ASAP7_75t_L g45 ( 
.A(n_28),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_45),
.B(n_34),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g46 ( 
.A1(n_35),
.A2(n_22),
.B1(n_21),
.B2(n_18),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_48),
.A2(n_49),
.B1(n_67),
.B2(n_63),
.Y(n_88)
);

OA22x2_ASAP7_75t_L g49 ( 
.A1(n_40),
.A2(n_29),
.B1(n_32),
.B2(n_30),
.Y(n_49)
);

INVxp67_ASAP7_75t_L g75 ( 
.A(n_50),
.Y(n_75)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_47),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_51),
.B(n_52),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g52 ( 
.A(n_47),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_38),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_53),
.B(n_65),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_40),
.A2(n_15),
.B1(n_31),
.B2(n_22),
.Y(n_54)
);

AOI21xp5_ASAP7_75t_L g81 ( 
.A1(n_54),
.A2(n_57),
.B(n_59),
.Y(n_81)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_41),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_55),
.B(n_68),
.Y(n_72)
);

INVx4_ASAP7_75t_SL g56 ( 
.A(n_43),
.Y(n_56)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_56),
.Y(n_74)
);

OR2x2_ASAP7_75t_SL g57 ( 
.A(n_40),
.B(n_19),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_44),
.B(n_30),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_58),
.B(n_64),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_37),
.A2(n_31),
.B1(n_21),
.B2(n_19),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_44),
.B(n_33),
.Y(n_60)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_60),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_45),
.B(n_17),
.Y(n_61)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_61),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_45),
.B(n_1),
.Y(n_62)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_62),
.Y(n_91)
);

OAI22xp33_ASAP7_75t_L g63 ( 
.A1(n_46),
.A2(n_36),
.B1(n_30),
.B2(n_28),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_63),
.A2(n_25),
.B1(n_13),
.B2(n_26),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_43),
.B(n_27),
.Y(n_64)
);

AOI21xp5_ASAP7_75t_L g82 ( 
.A1(n_66),
.A2(n_67),
.B(n_45),
.Y(n_82)
);

OR2x2_ASAP7_75t_SL g67 ( 
.A(n_39),
.B(n_25),
.Y(n_67)
);

CKINVDCx16_ASAP7_75t_R g68 ( 
.A(n_39),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_39),
.B(n_13),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_69),
.B(n_70),
.Y(n_79)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_41),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_53),
.B(n_43),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_76),
.B(n_78),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_77),
.B(n_87),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_58),
.B(n_52),
.Y(n_78)
);

XNOR2xp5_ASAP7_75t_L g101 ( 
.A(n_82),
.B(n_25),
.Y(n_101)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_55),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_83),
.B(n_70),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_51),
.A2(n_25),
.B1(n_45),
.B2(n_10),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_84),
.A2(n_88),
.B1(n_89),
.B2(n_56),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_49),
.B(n_1),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_49),
.A2(n_25),
.B1(n_10),
.B2(n_4),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_56),
.Y(n_92)
);

CKINVDCx10_ASAP7_75t_R g104 ( 
.A(n_92),
.Y(n_104)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_64),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_93),
.B(n_2),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_SL g94 ( 
.A(n_80),
.B(n_57),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_94),
.B(n_97),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_78),
.B(n_90),
.C(n_73),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_95),
.B(n_105),
.C(n_98),
.Y(n_115)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_72),
.Y(n_96)
);

INVxp67_ASAP7_75t_SL g125 ( 
.A(n_96),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_76),
.Y(n_97)
);

NOR2x1_ASAP7_75t_L g99 ( 
.A(n_87),
.B(n_49),
.Y(n_99)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_99),
.Y(n_114)
);

XNOR2xp5_ASAP7_75t_L g123 ( 
.A(n_101),
.B(n_81),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_SL g124 ( 
.A1(n_102),
.A2(n_108),
.B(n_111),
.Y(n_124)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_103),
.Y(n_117)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_73),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_105),
.B(n_109),
.Y(n_118)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_106),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_75),
.B(n_2),
.Y(n_107)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_107),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_88),
.A2(n_71),
.B1(n_3),
.B2(n_4),
.Y(n_108)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_85),
.Y(n_109)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_79),
.Y(n_110)
);

INVxp33_ASAP7_75t_L g121 ( 
.A(n_110),
.Y(n_121)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_84),
.Y(n_111)
);

INVx13_ASAP7_75t_L g112 ( 
.A(n_83),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_112),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_89),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_SL g127 ( 
.A1(n_113),
.A2(n_77),
.B(n_75),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_115),
.B(n_120),
.C(n_122),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_95),
.B(n_93),
.C(n_82),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_98),
.B(n_81),
.C(n_86),
.Y(n_122)
);

XOR2xp5_ASAP7_75t_L g140 ( 
.A(n_123),
.B(n_92),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_127),
.B(n_108),
.Y(n_130)
);

AOI21xp5_ASAP7_75t_L g129 ( 
.A1(n_99),
.A2(n_74),
.B(n_91),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_129),
.B(n_111),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_L g144 ( 
.A(n_130),
.B(n_132),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_118),
.B(n_97),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_131),
.B(n_133),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_SL g133 ( 
.A(n_119),
.B(n_109),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_125),
.B(n_104),
.Y(n_135)
);

CKINVDCx16_ASAP7_75t_R g147 ( 
.A(n_135),
.Y(n_147)
);

OAI322xp33_ASAP7_75t_L g136 ( 
.A1(n_118),
.A2(n_101),
.A3(n_113),
.B1(n_110),
.B2(n_102),
.C1(n_100),
.C2(n_96),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_L g149 ( 
.A(n_136),
.B(n_138),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_114),
.B(n_104),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_137),
.B(n_139),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_117),
.B(n_126),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_124),
.A2(n_74),
.B1(n_112),
.B2(n_71),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_140),
.B(n_141),
.C(n_122),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_SL g141 ( 
.A(n_128),
.B(n_2),
.Y(n_141)
);

INVx1_ASAP7_75t_SL g142 ( 
.A(n_137),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_142),
.B(n_150),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_SL g146 ( 
.A(n_140),
.B(n_123),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_SL g155 ( 
.A(n_146),
.B(n_3),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_148),
.B(n_4),
.C(n_5),
.Y(n_156)
);

BUFx12_ASAP7_75t_L g150 ( 
.A(n_134),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_143),
.A2(n_124),
.B1(n_139),
.B2(n_127),
.Y(n_151)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_151),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_145),
.A2(n_129),
.B1(n_120),
.B2(n_121),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_152),
.B(n_154),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_146),
.B(n_134),
.C(n_115),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_153),
.B(n_156),
.C(n_157),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_SL g154 ( 
.A1(n_147),
.A2(n_121),
.B(n_116),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_L g164 ( 
.A(n_155),
.B(n_6),
.Y(n_164)
);

XOR2xp5_ASAP7_75t_L g157 ( 
.A(n_149),
.B(n_5),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_L g162 ( 
.A1(n_158),
.A2(n_142),
.B(n_150),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_162),
.B(n_155),
.C(n_153),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_SL g163 ( 
.A(n_157),
.B(n_144),
.Y(n_163)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_163),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_164),
.B(n_7),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_165),
.B(n_166),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_159),
.B(n_150),
.C(n_8),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_168),
.B(n_164),
.Y(n_171)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_167),
.Y(n_169)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_169),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_171),
.B(n_159),
.Y(n_172)
);

AOI322xp5_ASAP7_75t_L g174 ( 
.A1(n_172),
.A2(n_170),
.A3(n_169),
.B1(n_160),
.B2(n_161),
.C1(n_173),
.C2(n_7),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_174),
.Y(n_175)
);

XOR2xp5_ASAP7_75t_L g176 ( 
.A(n_175),
.B(n_9),
.Y(n_176)
);


endmodule