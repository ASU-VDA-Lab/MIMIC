module real_jpeg_5107_n_14 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_2, n_13, n_6, n_7, n_3, n_10, n_9, n_14);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_2;
input n_13;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_14;

wire n_384;
wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_50;
wire n_409;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_366;
wire n_328;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_417;
wire n_128;
wire n_202;
wire n_216;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_393;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_387;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_402;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_420;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_404;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_273;
wire n_253;
wire n_16;
wire n_54;
wire n_168;
wire n_38;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_343;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_299;
wire n_243;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_32;
wire n_228;
wire n_389;
wire n_15;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_364;

INVx8_ASAP7_75t_L g70 ( 
.A(n_0),
.Y(n_70)
);

OAI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_1),
.A2(n_86),
.B1(n_89),
.B2(n_90),
.Y(n_85)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_1),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_1),
.A2(n_127),
.B1(n_128),
.B2(n_129),
.Y(n_126)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_1),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_1),
.A2(n_129),
.B1(n_163),
.B2(n_166),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_1),
.A2(n_129),
.B1(n_204),
.B2(n_206),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g46 ( 
.A1(n_2),
.A2(n_47),
.B1(n_49),
.B2(n_50),
.Y(n_46)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_2),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_2),
.A2(n_49),
.B1(n_156),
.B2(n_159),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_2),
.A2(n_49),
.B1(n_191),
.B2(n_193),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g220 ( 
.A1(n_2),
.A2(n_49),
.B1(n_221),
.B2(n_222),
.Y(n_220)
);

O2A1O1Ixp33_ASAP7_75t_L g258 ( 
.A1(n_2),
.A2(n_259),
.B(n_262),
.C(n_265),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_2),
.B(n_186),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_2),
.B(n_55),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_2),
.B(n_299),
.C(n_302),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_2),
.B(n_119),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_2),
.B(n_296),
.C(n_324),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_2),
.B(n_28),
.Y(n_342)
);

AOI22xp5_ASAP7_75t_L g21 ( 
.A1(n_3),
.A2(n_22),
.B1(n_24),
.B2(n_25),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_3),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_3),
.A2(n_24),
.B1(n_153),
.B2(n_155),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_3),
.A2(n_24),
.B1(n_34),
.B2(n_197),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_L g268 ( 
.A1(n_3),
.A2(n_24),
.B1(n_269),
.B2(n_270),
.Y(n_268)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_4),
.Y(n_59)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_4),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g180 ( 
.A(n_4),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g423 ( 
.A(n_5),
.Y(n_423)
);

OAI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_6),
.A2(n_79),
.B1(n_81),
.B2(n_82),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_6),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_6),
.A2(n_81),
.B1(n_121),
.B2(n_122),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_6),
.A2(n_81),
.B1(n_128),
.B2(n_134),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_6),
.A2(n_81),
.B1(n_178),
.B2(n_181),
.Y(n_177)
);

INVx6_ASAP7_75t_L g99 ( 
.A(n_7),
.Y(n_99)
);

INVx8_ASAP7_75t_L g175 ( 
.A(n_8),
.Y(n_175)
);

BUFx6f_ASAP7_75t_L g186 ( 
.A(n_8),
.Y(n_186)
);

BUFx6f_ASAP7_75t_L g212 ( 
.A(n_8),
.Y(n_212)
);

BUFx5_ASAP7_75t_L g287 ( 
.A(n_8),
.Y(n_287)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_9),
.Y(n_37)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_9),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g261 ( 
.A(n_9),
.Y(n_261)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

INVx3_ASAP7_75t_L g419 ( 
.A(n_11),
.Y(n_419)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

INVx6_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_12),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_12),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_12),
.Y(n_48)
);

BUFx5_ASAP7_75t_L g50 ( 
.A(n_12),
.Y(n_50)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_12),
.Y(n_138)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_13),
.Y(n_57)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_13),
.Y(n_64)
);

AOI21xp5_ASAP7_75t_L g14 ( 
.A1(n_15),
.A2(n_418),
.B(n_420),
.Y(n_14)
);

XNOR2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_141),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_SL g16 ( 
.A(n_17),
.B(n_139),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_SL g17 ( 
.A(n_18),
.B(n_132),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_18),
.B(n_132),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_125),
.C(n_130),
.Y(n_18)
);

XOR2xp5_ASAP7_75t_L g414 ( 
.A(n_19),
.B(n_415),
.Y(n_414)
);

MAJIxp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_52),
.C(n_84),
.Y(n_19)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_20),
.A2(n_188),
.B1(n_189),
.B2(n_199),
.Y(n_187)
);

CKINVDCx16_ASAP7_75t_R g199 ( 
.A(n_20),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_20),
.B(n_148),
.C(n_189),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_20),
.B(n_240),
.C(n_257),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g366 ( 
.A1(n_20),
.A2(n_199),
.B1(n_240),
.B2(n_343),
.Y(n_366)
);

AOI22xp5_ASAP7_75t_L g389 ( 
.A1(n_20),
.A2(n_199),
.B1(n_390),
.B2(n_391),
.Y(n_389)
);

OA22x2_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_27),
.B1(n_46),
.B2(n_51),
.Y(n_20)
);

OA22x2_ASAP7_75t_L g228 ( 
.A1(n_21),
.A2(n_27),
.B1(n_46),
.B2(n_51),
.Y(n_228)
);

INVx4_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

INVx8_ASAP7_75t_L g127 ( 
.A(n_23),
.Y(n_127)
);

INVx8_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_27),
.A2(n_46),
.B1(n_51),
.B2(n_126),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_27),
.A2(n_51),
.B1(n_126),
.B2(n_133),
.Y(n_132)
);

AOI21xp5_ASAP7_75t_L g235 ( 
.A1(n_27),
.A2(n_46),
.B(n_51),
.Y(n_235)
);

OR2x2_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_38),
.Y(n_27)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_28),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g28 ( 
.A1(n_29),
.A2(n_32),
.B1(n_34),
.B2(n_36),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_30),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_30),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g322 ( 
.A(n_30),
.Y(n_322)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g88 ( 
.A(n_31),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_31),
.Y(n_92)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_31),
.Y(n_108)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_31),
.Y(n_195)
);

AOI22xp33_ASAP7_75t_L g38 ( 
.A1(n_32),
.A2(n_39),
.B1(n_41),
.B2(n_43),
.Y(n_38)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx3_ASAP7_75t_SL g263 ( 
.A(n_33),
.Y(n_263)
);

INVx5_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx5_ASAP7_75t_L g265 ( 
.A(n_39),
.Y(n_265)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

OAI21xp33_ASAP7_75t_L g262 ( 
.A1(n_49),
.A2(n_263),
.B(n_264),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_SL g391 ( 
.A1(n_52),
.A2(n_84),
.B1(n_392),
.B2(n_393),
.Y(n_391)
);

CKINVDCx14_ASAP7_75t_R g393 ( 
.A(n_52),
.Y(n_393)
);

MAJIxp5_ASAP7_75t_L g394 ( 
.A(n_52),
.B(n_228),
.C(n_395),
.Y(n_394)
);

OAI22xp5_ASAP7_75t_SL g401 ( 
.A1(n_52),
.A2(n_393),
.B1(n_395),
.B2(n_402),
.Y(n_401)
);

AND2x2_ASAP7_75t_SL g52 ( 
.A(n_53),
.B(n_78),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_53),
.B(n_158),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_54),
.B(n_65),
.Y(n_53)
);

OA22x2_ASAP7_75t_L g150 ( 
.A1(n_54),
.A2(n_65),
.B1(n_151),
.B2(n_157),
.Y(n_150)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

NOR2x1_ASAP7_75t_L g66 ( 
.A(n_55),
.B(n_67),
.Y(n_66)
);

AOI21xp5_ASAP7_75t_L g202 ( 
.A1(n_55),
.A2(n_203),
.B(n_207),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_55),
.B(n_152),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_55),
.A2(n_66),
.B1(n_78),
.B2(n_203),
.Y(n_239)
);

AO22x1_ASAP7_75t_SL g55 ( 
.A1(n_56),
.A2(n_58),
.B1(n_60),
.B2(n_63),
.Y(n_55)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx5_ASAP7_75t_L g72 ( 
.A(n_57),
.Y(n_72)
);

INVx4_ASAP7_75t_L g301 ( 
.A(n_57),
.Y(n_301)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_58),
.Y(n_223)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

BUFx5_ASAP7_75t_L g171 ( 
.A(n_59),
.Y(n_171)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx4_ASAP7_75t_L g167 ( 
.A(n_61),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g165 ( 
.A(n_62),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g182 ( 
.A(n_62),
.Y(n_182)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx1_ASAP7_75t_SL g65 ( 
.A(n_66),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_66),
.B(n_158),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g67 ( 
.A1(n_68),
.A2(n_71),
.B1(n_73),
.B2(n_74),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx3_ASAP7_75t_L g159 ( 
.A(n_69),
.Y(n_159)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx11_ASAP7_75t_L g77 ( 
.A(n_70),
.Y(n_77)
);

BUFx5_ASAP7_75t_L g115 ( 
.A(n_70),
.Y(n_115)
);

INVx3_ASAP7_75t_L g156 ( 
.A(n_70),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g297 ( 
.A(n_70),
.Y(n_297)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_71),
.Y(n_73)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_75),
.Y(n_205)
);

INVx5_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx5_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_77),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_77),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_77),
.Y(n_111)
);

INVx3_ASAP7_75t_L g206 ( 
.A(n_79),
.Y(n_206)
);

INVx6_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVx11_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_84),
.Y(n_392)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_85),
.A2(n_93),
.B1(n_119),
.B2(n_120),
.Y(n_84)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_85),
.Y(n_396)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

BUFx3_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_88),
.Y(n_124)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_88),
.Y(n_192)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_92),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g198 ( 
.A(n_92),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g397 ( 
.A(n_93),
.B(n_227),
.Y(n_397)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_94),
.B(n_109),
.Y(n_131)
);

OA22x2_ASAP7_75t_L g189 ( 
.A1(n_94),
.A2(n_109),
.B1(n_190),
.B2(n_196),
.Y(n_189)
);

OA22x2_ASAP7_75t_L g240 ( 
.A1(n_94),
.A2(n_109),
.B1(n_190),
.B2(n_196),
.Y(n_240)
);

NAND2x1_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_109),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_96),
.A2(n_100),
.B1(n_104),
.B2(n_106),
.Y(n_95)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_99),
.Y(n_105)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_99),
.Y(n_113)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx5_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx4_ASAP7_75t_L g264 ( 
.A(n_103),
.Y(n_264)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx4_ASAP7_75t_L g327 ( 
.A(n_105),
.Y(n_327)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_109),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_L g395 ( 
.A1(n_109),
.A2(n_396),
.B(n_397),
.Y(n_395)
);

AOI22x1_ASAP7_75t_L g109 ( 
.A1(n_110),
.A2(n_112),
.B1(n_114),
.B2(n_116),
.Y(n_109)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_111),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx4_ASAP7_75t_L g118 ( 
.A(n_113),
.Y(n_118)
);

INVx5_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_120),
.B(n_131),
.Y(n_130)
);

HB1xp67_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

XOR2xp5_ASAP7_75t_L g415 ( 
.A(n_125),
.B(n_130),
.Y(n_415)
);

INVx8_ASAP7_75t_L g128 ( 
.A(n_127),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_131),
.B(n_227),
.Y(n_226)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx3_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

INVx4_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

INVxp67_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_SL g141 ( 
.A1(n_142),
.A2(n_413),
.B(n_417),
.Y(n_141)
);

AOI21xp5_ASAP7_75t_L g142 ( 
.A1(n_143),
.A2(n_384),
.B(n_410),
.Y(n_142)
);

OAI211xp5_ASAP7_75t_L g143 ( 
.A1(n_144),
.A2(n_273),
.B(n_378),
.C(n_383),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_245),
.Y(n_144)
);

A2O1A1Ixp33_ASAP7_75t_L g378 ( 
.A1(n_145),
.A2(n_245),
.B(n_379),
.C(n_382),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_146),
.B(n_229),
.Y(n_145)
);

OR2x2_ASAP7_75t_L g383 ( 
.A(n_146),
.B(n_229),
.Y(n_383)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_200),
.C(n_214),
.Y(n_146)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_147),
.B(n_200),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g147 ( 
.A(n_148),
.B(n_187),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_149),
.B(n_160),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g254 ( 
.A1(n_149),
.A2(n_150),
.B1(n_160),
.B2(n_255),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_L g309 ( 
.A1(n_149),
.A2(n_150),
.B1(n_310),
.B2(n_311),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_SL g334 ( 
.A1(n_149),
.A2(n_150),
.B1(n_335),
.B2(n_336),
.Y(n_334)
);

INVx3_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_150),
.B(n_267),
.C(n_310),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g348 ( 
.A(n_150),
.B(n_335),
.C(n_337),
.Y(n_348)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

INVx3_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

INVx4_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

INVxp67_ASAP7_75t_L g255 ( 
.A(n_160),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_161),
.A2(n_168),
.B1(n_176),
.B2(n_183),
.Y(n_160)
);

INVxp67_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

AOI21xp5_ASAP7_75t_L g217 ( 
.A1(n_162),
.A2(n_184),
.B(n_218),
.Y(n_217)
);

INVx4_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

INVx2_ASAP7_75t_L g303 ( 
.A(n_165),
.Y(n_303)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_166),
.Y(n_221)
);

INVx4_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_168),
.B(n_211),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_168),
.B(n_219),
.Y(n_218)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_169),
.A2(n_220),
.B1(n_268),
.B2(n_271),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_169),
.A2(n_220),
.B1(n_268),
.B2(n_285),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_172),
.Y(n_169)
);

INVx3_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

INVx3_ASAP7_75t_L g270 ( 
.A(n_171),
.Y(n_270)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

INVx4_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

BUFx6f_ASAP7_75t_L g272 ( 
.A(n_175),
.Y(n_272)
);

INVxp67_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_177),
.B(n_210),
.Y(n_209)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

INVx3_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

BUFx6f_ASAP7_75t_L g269 ( 
.A(n_180),
.Y(n_269)
);

BUFx6f_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_184),
.Y(n_183)
);

BUFx3_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

BUFx6f_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g330 ( 
.A1(n_188),
.A2(n_189),
.B1(n_224),
.B2(n_294),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g345 ( 
.A(n_188),
.B(n_294),
.C(n_317),
.Y(n_345)
);

OAI22xp5_ASAP7_75t_SL g352 ( 
.A1(n_188),
.A2(n_189),
.B1(n_353),
.B2(n_354),
.Y(n_352)
);

CKINVDCx16_ASAP7_75t_R g188 ( 
.A(n_189),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g370 ( 
.A(n_189),
.B(n_228),
.C(n_353),
.Y(n_370)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_190),
.Y(n_227)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

INVx5_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

INVx6_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

INVx5_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_201),
.A2(n_202),
.B1(n_209),
.B2(n_213),
.Y(n_200)
);

INVxp67_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_202),
.B(n_209),
.Y(n_236)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

INVxp67_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

AND2x2_ASAP7_75t_SL g224 ( 
.A(n_208),
.B(n_225),
.Y(n_224)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_209),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_209),
.A2(n_213),
.B1(n_234),
.B2(n_235),
.Y(n_233)
);

OAI21xp5_ASAP7_75t_L g404 ( 
.A1(n_209),
.A2(n_235),
.B(n_236),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_210),
.B(n_220),
.Y(n_328)
);

INVx3_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_214),
.B(n_247),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_215),
.B(n_226),
.C(n_228),
.Y(n_214)
);

INVxp67_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_216),
.B(n_251),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_217),
.B(n_224),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_L g368 ( 
.A1(n_217),
.A2(n_224),
.B1(n_294),
.B2(n_369),
.Y(n_368)
);

INVxp67_ASAP7_75t_L g369 ( 
.A(n_217),
.Y(n_369)
);

INVxp67_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_224),
.A2(n_294),
.B1(n_295),
.B2(n_304),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_224),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_226),
.A2(n_228),
.B1(n_252),
.B2(n_253),
.Y(n_251)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_226),
.Y(n_253)
);

INVx2_ASAP7_75t_SL g252 ( 
.A(n_228),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g350 ( 
.A1(n_228),
.A2(n_252),
.B1(n_351),
.B2(n_352),
.Y(n_350)
);

OAI22xp5_ASAP7_75t_SL g387 ( 
.A1(n_228),
.A2(n_252),
.B1(n_388),
.B2(n_389),
.Y(n_387)
);

AOI22xp5_ASAP7_75t_L g399 ( 
.A1(n_228),
.A2(n_252),
.B1(n_400),
.B2(n_401),
.Y(n_399)
);

MAJIxp5_ASAP7_75t_L g416 ( 
.A(n_228),
.B(n_389),
.C(n_394),
.Y(n_416)
);

AOI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_230),
.A2(n_231),
.B1(n_243),
.B2(n_244),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_232),
.A2(n_237),
.B1(n_238),
.B2(n_242),
.Y(n_231)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_232),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g232 ( 
.A(n_233),
.B(n_236),
.Y(n_232)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g409 ( 
.A(n_237),
.B(n_242),
.C(n_244),
.Y(n_409)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

OAI21xp5_ASAP7_75t_L g238 ( 
.A1(n_239),
.A2(n_240),
.B(n_241),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_239),
.B(n_240),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g338 ( 
.A1(n_240),
.A2(n_339),
.B1(n_340),
.B2(n_343),
.Y(n_338)
);

CKINVDCx16_ASAP7_75t_R g343 ( 
.A(n_240),
.Y(n_343)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_241),
.Y(n_403)
);

OAI22xp5_ASAP7_75t_SL g407 ( 
.A1(n_241),
.A2(n_399),
.B1(n_403),
.B2(n_408),
.Y(n_407)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_243),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_SL g245 ( 
.A(n_246),
.B(n_248),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g382 ( 
.A(n_246),
.B(n_248),
.Y(n_382)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_249),
.B(n_254),
.C(n_256),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_L g376 ( 
.A1(n_249),
.A2(n_250),
.B1(n_254),
.B2(n_377),
.Y(n_376)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_254),
.Y(n_377)
);

XNOR2xp5_ASAP7_75t_L g375 ( 
.A(n_256),
.B(n_376),
.Y(n_375)
);

XOR2xp5_ASAP7_75t_L g365 ( 
.A(n_257),
.B(n_366),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_258),
.B(n_266),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_SL g359 ( 
.A1(n_258),
.A2(n_266),
.B1(n_267),
.B2(n_360),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_258),
.Y(n_360)
);

INVx6_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

INVx4_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_266),
.A2(n_267),
.B1(n_308),
.B2(n_309),
.Y(n_307)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_267),
.B(n_289),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_267),
.B(n_289),
.Y(n_290)
);

INVx1_ASAP7_75t_SL g282 ( 
.A(n_270),
.Y(n_282)
);

INVx8_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_SL g273 ( 
.A(n_274),
.B(n_362),
.Y(n_273)
);

OAI21xp5_ASAP7_75t_SL g274 ( 
.A1(n_275),
.A2(n_347),
.B(n_361),
.Y(n_274)
);

AOI21xp5_ASAP7_75t_L g275 ( 
.A1(n_276),
.A2(n_332),
.B(n_346),
.Y(n_275)
);

OAI21xp5_ASAP7_75t_SL g276 ( 
.A1(n_277),
.A2(n_314),
.B(n_331),
.Y(n_276)
);

AOI21xp5_ASAP7_75t_L g277 ( 
.A1(n_278),
.A2(n_306),
.B(n_313),
.Y(n_277)
);

OAI21xp5_ASAP7_75t_L g278 ( 
.A1(n_279),
.A2(n_291),
.B(n_305),
.Y(n_278)
);

AOI21xp5_ASAP7_75t_SL g279 ( 
.A1(n_280),
.A2(n_288),
.B(n_290),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_281),
.B(n_284),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_282),
.B(n_283),
.Y(n_281)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_284),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_L g340 ( 
.A1(n_284),
.A2(n_292),
.B1(n_341),
.B2(n_342),
.Y(n_340)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_292),
.B(n_293),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_292),
.B(n_293),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g357 ( 
.A(n_292),
.B(n_341),
.C(n_343),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_294),
.B(n_304),
.Y(n_312)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_295),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_296),
.B(n_298),
.Y(n_295)
);

INVx5_ASAP7_75t_L g296 ( 
.A(n_297),
.Y(n_296)
);

INVx3_ASAP7_75t_L g299 ( 
.A(n_300),
.Y(n_299)
);

INVx4_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

BUFx3_ASAP7_75t_L g302 ( 
.A(n_303),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_SL g306 ( 
.A(n_307),
.B(n_312),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_307),
.B(n_312),
.Y(n_313)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_309),
.Y(n_308)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_310),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_315),
.B(n_316),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_315),
.B(n_316),
.Y(n_331)
);

XOR2xp5_ASAP7_75t_L g316 ( 
.A(n_317),
.B(n_330),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_L g317 ( 
.A1(n_318),
.A2(n_319),
.B1(n_328),
.B2(n_329),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_318),
.B(n_329),
.Y(n_335)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_319),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_320),
.B(n_323),
.Y(n_319)
);

INVx2_ASAP7_75t_L g320 ( 
.A(n_321),
.Y(n_320)
);

INVx2_ASAP7_75t_L g321 ( 
.A(n_322),
.Y(n_321)
);

INVx2_ASAP7_75t_L g324 ( 
.A(n_325),
.Y(n_324)
);

INVx3_ASAP7_75t_L g325 ( 
.A(n_326),
.Y(n_325)
);

INVx6_ASAP7_75t_L g326 ( 
.A(n_327),
.Y(n_326)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_328),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_SL g332 ( 
.A(n_333),
.B(n_345),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g346 ( 
.A(n_333),
.B(n_345),
.Y(n_346)
);

AOI22xp5_ASAP7_75t_L g333 ( 
.A1(n_334),
.A2(n_337),
.B1(n_338),
.B2(n_344),
.Y(n_333)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_334),
.Y(n_344)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_335),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_338),
.Y(n_337)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_340),
.Y(n_339)
);

CKINVDCx14_ASAP7_75t_R g341 ( 
.A(n_342),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_L g347 ( 
.A(n_348),
.B(n_349),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_348),
.B(n_349),
.Y(n_361)
);

XNOR2xp5_ASAP7_75t_L g349 ( 
.A(n_350),
.B(n_355),
.Y(n_349)
);

MAJIxp5_ASAP7_75t_L g371 ( 
.A(n_350),
.B(n_357),
.C(n_358),
.Y(n_371)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_352),
.Y(n_351)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_353),
.Y(n_354)
);

OAI22xp5_ASAP7_75t_SL g355 ( 
.A1(n_356),
.A2(n_357),
.B1(n_358),
.B2(n_359),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_357),
.Y(n_356)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_359),
.Y(n_358)
);

NOR2x1_ASAP7_75t_L g362 ( 
.A(n_363),
.B(n_372),
.Y(n_362)
);

NOR2xp33_ASAP7_75t_SL g363 ( 
.A(n_364),
.B(n_371),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_364),
.B(n_371),
.Y(n_380)
);

XNOR2xp5_ASAP7_75t_L g364 ( 
.A(n_365),
.B(n_367),
.Y(n_364)
);

INVxp67_ASAP7_75t_L g374 ( 
.A(n_365),
.Y(n_374)
);

XOR2xp5_ASAP7_75t_L g367 ( 
.A(n_368),
.B(n_370),
.Y(n_367)
);

MAJIxp5_ASAP7_75t_L g373 ( 
.A(n_368),
.B(n_370),
.C(n_374),
.Y(n_373)
);

OAI21xp5_ASAP7_75t_L g379 ( 
.A1(n_372),
.A2(n_380),
.B(n_381),
.Y(n_379)
);

AND2x2_ASAP7_75t_L g372 ( 
.A(n_373),
.B(n_375),
.Y(n_372)
);

OR2x2_ASAP7_75t_L g381 ( 
.A(n_373),
.B(n_375),
.Y(n_381)
);

NOR2xp33_ASAP7_75t_L g384 ( 
.A(n_385),
.B(n_405),
.Y(n_384)
);

OAI21xp5_ASAP7_75t_L g410 ( 
.A1(n_385),
.A2(n_411),
.B(n_412),
.Y(n_410)
);

NOR2xp33_ASAP7_75t_SL g385 ( 
.A(n_386),
.B(n_398),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_386),
.B(n_398),
.Y(n_412)
);

XNOR2xp5_ASAP7_75t_L g386 ( 
.A(n_387),
.B(n_394),
.Y(n_386)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_389),
.Y(n_388)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_391),
.Y(n_390)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_395),
.Y(n_402)
);

MAJIxp5_ASAP7_75t_L g398 ( 
.A(n_399),
.B(n_403),
.C(n_404),
.Y(n_398)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_399),
.Y(n_408)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_401),
.Y(n_400)
);

XNOR2xp5_ASAP7_75t_L g406 ( 
.A(n_404),
.B(n_407),
.Y(n_406)
);

NOR2xp33_ASAP7_75t_SL g405 ( 
.A(n_406),
.B(n_409),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_406),
.B(n_409),
.Y(n_411)
);

NOR2xp33_ASAP7_75t_L g413 ( 
.A(n_414),
.B(n_416),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g417 ( 
.A(n_414),
.B(n_416),
.Y(n_417)
);

INVx6_ASAP7_75t_L g418 ( 
.A(n_419),
.Y(n_418)
);

INVx13_ASAP7_75t_L g422 ( 
.A(n_419),
.Y(n_422)
);

NOR2xp33_ASAP7_75t_L g420 ( 
.A(n_421),
.B(n_423),
.Y(n_420)
);

BUFx4f_ASAP7_75t_SL g421 ( 
.A(n_422),
.Y(n_421)
);


endmodule