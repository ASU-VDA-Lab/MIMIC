module fake_netlist_5_1235_n_4853 (n_137, n_294, n_431, n_318, n_380, n_419, n_444, n_469, n_82, n_194, n_316, n_389, n_418, n_248, n_124, n_86, n_136, n_146, n_315, n_268, n_523, n_451, n_532, n_408, n_61, n_376, n_503, n_127, n_75, n_235, n_226, n_74, n_515, n_57, n_353, n_351, n_367, n_452, n_397, n_493, n_111, n_525, n_483, n_155, n_43, n_116, n_22, n_467, n_423, n_284, n_46, n_245, n_21, n_501, n_139, n_38, n_105, n_280, n_4, n_378, n_17, n_382, n_254, n_33, n_23, n_302, n_265, n_526, n_293, n_372, n_443, n_244, n_47, n_173, n_198, n_447, n_247, n_314, n_368, n_433, n_8, n_321, n_292, n_100, n_455, n_417, n_212, n_385, n_498, n_516, n_507, n_119, n_497, n_275, n_252, n_26, n_295, n_133, n_330, n_508, n_506, n_2, n_6, n_509, n_39, n_147, n_373, n_67, n_307, n_439, n_87, n_150, n_530, n_106, n_209, n_259, n_448, n_375, n_301, n_68, n_93, n_186, n_537, n_134, n_191, n_51, n_63, n_492, n_171, n_153, n_524, n_399, n_341, n_204, n_394, n_250, n_543, n_260, n_298, n_320, n_518, n_505, n_286, n_122, n_282, n_331, n_10, n_24, n_406, n_519, n_470, n_325, n_449, n_132, n_90, n_101, n_281, n_240, n_381, n_189, n_220, n_291, n_231, n_257, n_390, n_31, n_456, n_13, n_371, n_481, n_535, n_152, n_540, n_317, n_9, n_323, n_195, n_42, n_356, n_227, n_45, n_271, n_94, n_335, n_123, n_370, n_167, n_234, n_343, n_308, n_379, n_428, n_267, n_514, n_457, n_297, n_156, n_5, n_225, n_377, n_484, n_219, n_442, n_157, n_131, n_192, n_223, n_392, n_158, n_138, n_264, n_109, n_472, n_454, n_387, n_374, n_163, n_276, n_339, n_95, n_183, n_185, n_243, n_398, n_396, n_347, n_169, n_59, n_522, n_255, n_215, n_350, n_196, n_459, n_211, n_218, n_400, n_181, n_436, n_3, n_290, n_221, n_178, n_386, n_287, n_344, n_473, n_422, n_475, n_72, n_104, n_41, n_415, n_56, n_141, n_485, n_496, n_355, n_486, n_15, n_336, n_145, n_48, n_521, n_50, n_337, n_430, n_313, n_88, n_479, n_528, n_510, n_216, n_168, n_395, n_164, n_432, n_311, n_208, n_142, n_214, n_328, n_140, n_299, n_303, n_369, n_296, n_241, n_357, n_184, n_446, n_445, n_65, n_78, n_144, n_114, n_96, n_165, n_468, n_499, n_213, n_129, n_342, n_482, n_517, n_98, n_361, n_464, n_363, n_402, n_413, n_197, n_107, n_69, n_236, n_388, n_1, n_249, n_304, n_329, n_203, n_274, n_384, n_460, n_80, n_35, n_73, n_277, n_92, n_19, n_338, n_149, n_477, n_461, n_333, n_309, n_30, n_512, n_14, n_84, n_462, n_130, n_322, n_258, n_29, n_79, n_151, n_25, n_306, n_458, n_288, n_188, n_190, n_201, n_263, n_471, n_44, n_224, n_40, n_34, n_228, n_283, n_383, n_474, n_112, n_542, n_85, n_463, n_488, n_502, n_239, n_466, n_420, n_489, n_55, n_49, n_310, n_54, n_504, n_511, n_12, n_465, n_76, n_358, n_362, n_170, n_332, n_27, n_77, n_102, n_161, n_273, n_349, n_270, n_230, n_81, n_118, n_279, n_70, n_253, n_261, n_174, n_289, n_172, n_206, n_217, n_440, n_478, n_441, n_450, n_312, n_476, n_429, n_534, n_345, n_210, n_494, n_365, n_91, n_176, n_182, n_143, n_83, n_354, n_480, n_237, n_425, n_513, n_407, n_527, n_180, n_340, n_207, n_37, n_346, n_393, n_229, n_108, n_487, n_495, n_437, n_66, n_177, n_60, n_403, n_453, n_421, n_16, n_0, n_58, n_405, n_18, n_359, n_490, n_117, n_326, n_233, n_404, n_205, n_366, n_113, n_246, n_179, n_125, n_410, n_269, n_529, n_128, n_285, n_412, n_120, n_232, n_327, n_135, n_126, n_202, n_266, n_272, n_491, n_427, n_193, n_251, n_352, n_53, n_160, n_426, n_520, n_409, n_500, n_154, n_62, n_148, n_71, n_300, n_435, n_159, n_334, n_541, n_391, n_434, n_539, n_175, n_538, n_262, n_238, n_99, n_411, n_414, n_319, n_364, n_20, n_536, n_531, n_121, n_242, n_360, n_36, n_200, n_162, n_64, n_222, n_28, n_89, n_438, n_115, n_324, n_416, n_199, n_187, n_32, n_401, n_103, n_348, n_97, n_166, n_11, n_424, n_7, n_256, n_305, n_533, n_52, n_278, n_110, n_4853);

input n_137;
input n_294;
input n_431;
input n_318;
input n_380;
input n_419;
input n_444;
input n_469;
input n_82;
input n_194;
input n_316;
input n_389;
input n_418;
input n_248;
input n_124;
input n_86;
input n_136;
input n_146;
input n_315;
input n_268;
input n_523;
input n_451;
input n_532;
input n_408;
input n_61;
input n_376;
input n_503;
input n_127;
input n_75;
input n_235;
input n_226;
input n_74;
input n_515;
input n_57;
input n_353;
input n_351;
input n_367;
input n_452;
input n_397;
input n_493;
input n_111;
input n_525;
input n_483;
input n_155;
input n_43;
input n_116;
input n_22;
input n_467;
input n_423;
input n_284;
input n_46;
input n_245;
input n_21;
input n_501;
input n_139;
input n_38;
input n_105;
input n_280;
input n_4;
input n_378;
input n_17;
input n_382;
input n_254;
input n_33;
input n_23;
input n_302;
input n_265;
input n_526;
input n_293;
input n_372;
input n_443;
input n_244;
input n_47;
input n_173;
input n_198;
input n_447;
input n_247;
input n_314;
input n_368;
input n_433;
input n_8;
input n_321;
input n_292;
input n_100;
input n_455;
input n_417;
input n_212;
input n_385;
input n_498;
input n_516;
input n_507;
input n_119;
input n_497;
input n_275;
input n_252;
input n_26;
input n_295;
input n_133;
input n_330;
input n_508;
input n_506;
input n_2;
input n_6;
input n_509;
input n_39;
input n_147;
input n_373;
input n_67;
input n_307;
input n_439;
input n_87;
input n_150;
input n_530;
input n_106;
input n_209;
input n_259;
input n_448;
input n_375;
input n_301;
input n_68;
input n_93;
input n_186;
input n_537;
input n_134;
input n_191;
input n_51;
input n_63;
input n_492;
input n_171;
input n_153;
input n_524;
input n_399;
input n_341;
input n_204;
input n_394;
input n_250;
input n_543;
input n_260;
input n_298;
input n_320;
input n_518;
input n_505;
input n_286;
input n_122;
input n_282;
input n_331;
input n_10;
input n_24;
input n_406;
input n_519;
input n_470;
input n_325;
input n_449;
input n_132;
input n_90;
input n_101;
input n_281;
input n_240;
input n_381;
input n_189;
input n_220;
input n_291;
input n_231;
input n_257;
input n_390;
input n_31;
input n_456;
input n_13;
input n_371;
input n_481;
input n_535;
input n_152;
input n_540;
input n_317;
input n_9;
input n_323;
input n_195;
input n_42;
input n_356;
input n_227;
input n_45;
input n_271;
input n_94;
input n_335;
input n_123;
input n_370;
input n_167;
input n_234;
input n_343;
input n_308;
input n_379;
input n_428;
input n_267;
input n_514;
input n_457;
input n_297;
input n_156;
input n_5;
input n_225;
input n_377;
input n_484;
input n_219;
input n_442;
input n_157;
input n_131;
input n_192;
input n_223;
input n_392;
input n_158;
input n_138;
input n_264;
input n_109;
input n_472;
input n_454;
input n_387;
input n_374;
input n_163;
input n_276;
input n_339;
input n_95;
input n_183;
input n_185;
input n_243;
input n_398;
input n_396;
input n_347;
input n_169;
input n_59;
input n_522;
input n_255;
input n_215;
input n_350;
input n_196;
input n_459;
input n_211;
input n_218;
input n_400;
input n_181;
input n_436;
input n_3;
input n_290;
input n_221;
input n_178;
input n_386;
input n_287;
input n_344;
input n_473;
input n_422;
input n_475;
input n_72;
input n_104;
input n_41;
input n_415;
input n_56;
input n_141;
input n_485;
input n_496;
input n_355;
input n_486;
input n_15;
input n_336;
input n_145;
input n_48;
input n_521;
input n_50;
input n_337;
input n_430;
input n_313;
input n_88;
input n_479;
input n_528;
input n_510;
input n_216;
input n_168;
input n_395;
input n_164;
input n_432;
input n_311;
input n_208;
input n_142;
input n_214;
input n_328;
input n_140;
input n_299;
input n_303;
input n_369;
input n_296;
input n_241;
input n_357;
input n_184;
input n_446;
input n_445;
input n_65;
input n_78;
input n_144;
input n_114;
input n_96;
input n_165;
input n_468;
input n_499;
input n_213;
input n_129;
input n_342;
input n_482;
input n_517;
input n_98;
input n_361;
input n_464;
input n_363;
input n_402;
input n_413;
input n_197;
input n_107;
input n_69;
input n_236;
input n_388;
input n_1;
input n_249;
input n_304;
input n_329;
input n_203;
input n_274;
input n_384;
input n_460;
input n_80;
input n_35;
input n_73;
input n_277;
input n_92;
input n_19;
input n_338;
input n_149;
input n_477;
input n_461;
input n_333;
input n_309;
input n_30;
input n_512;
input n_14;
input n_84;
input n_462;
input n_130;
input n_322;
input n_258;
input n_29;
input n_79;
input n_151;
input n_25;
input n_306;
input n_458;
input n_288;
input n_188;
input n_190;
input n_201;
input n_263;
input n_471;
input n_44;
input n_224;
input n_40;
input n_34;
input n_228;
input n_283;
input n_383;
input n_474;
input n_112;
input n_542;
input n_85;
input n_463;
input n_488;
input n_502;
input n_239;
input n_466;
input n_420;
input n_489;
input n_55;
input n_49;
input n_310;
input n_54;
input n_504;
input n_511;
input n_12;
input n_465;
input n_76;
input n_358;
input n_362;
input n_170;
input n_332;
input n_27;
input n_77;
input n_102;
input n_161;
input n_273;
input n_349;
input n_270;
input n_230;
input n_81;
input n_118;
input n_279;
input n_70;
input n_253;
input n_261;
input n_174;
input n_289;
input n_172;
input n_206;
input n_217;
input n_440;
input n_478;
input n_441;
input n_450;
input n_312;
input n_476;
input n_429;
input n_534;
input n_345;
input n_210;
input n_494;
input n_365;
input n_91;
input n_176;
input n_182;
input n_143;
input n_83;
input n_354;
input n_480;
input n_237;
input n_425;
input n_513;
input n_407;
input n_527;
input n_180;
input n_340;
input n_207;
input n_37;
input n_346;
input n_393;
input n_229;
input n_108;
input n_487;
input n_495;
input n_437;
input n_66;
input n_177;
input n_60;
input n_403;
input n_453;
input n_421;
input n_16;
input n_0;
input n_58;
input n_405;
input n_18;
input n_359;
input n_490;
input n_117;
input n_326;
input n_233;
input n_404;
input n_205;
input n_366;
input n_113;
input n_246;
input n_179;
input n_125;
input n_410;
input n_269;
input n_529;
input n_128;
input n_285;
input n_412;
input n_120;
input n_232;
input n_327;
input n_135;
input n_126;
input n_202;
input n_266;
input n_272;
input n_491;
input n_427;
input n_193;
input n_251;
input n_352;
input n_53;
input n_160;
input n_426;
input n_520;
input n_409;
input n_500;
input n_154;
input n_62;
input n_148;
input n_71;
input n_300;
input n_435;
input n_159;
input n_334;
input n_541;
input n_391;
input n_434;
input n_539;
input n_175;
input n_538;
input n_262;
input n_238;
input n_99;
input n_411;
input n_414;
input n_319;
input n_364;
input n_20;
input n_536;
input n_531;
input n_121;
input n_242;
input n_360;
input n_36;
input n_200;
input n_162;
input n_64;
input n_222;
input n_28;
input n_89;
input n_438;
input n_115;
input n_324;
input n_416;
input n_199;
input n_187;
input n_32;
input n_401;
input n_103;
input n_348;
input n_97;
input n_166;
input n_11;
input n_424;
input n_7;
input n_256;
input n_305;
input n_533;
input n_52;
input n_278;
input n_110;

output n_4853;

wire n_924;
wire n_1263;
wire n_3304;
wire n_977;
wire n_1378;
wire n_2417;
wire n_2756;
wire n_611;
wire n_2253;
wire n_3912;
wire n_1126;
wire n_1423;
wire n_1729;
wire n_4706;
wire n_2739;
wire n_1166;
wire n_2380;
wire n_1751;
wire n_2771;
wire n_3241;
wire n_785;
wire n_1508;
wire n_4129;
wire n_4604;
wire n_549;
wire n_2617;
wire n_2200;
wire n_3261;
wire n_3006;
wire n_4798;
wire n_1161;
wire n_3795;
wire n_3863;
wire n_3027;
wire n_1859;
wire n_4419;
wire n_2746;
wire n_1677;
wire n_4477;
wire n_1150;
wire n_2327;
wire n_3179;
wire n_3127;
wire n_3256;
wire n_1780;
wire n_3732;
wire n_1488;
wire n_4250;
wire n_667;
wire n_2899;
wire n_2955;
wire n_790;
wire n_3619;
wire n_1055;
wire n_3541;
wire n_3622;
wire n_4112;
wire n_2386;
wire n_3596;
wire n_1501;
wire n_4699;
wire n_4337;
wire n_2395;
wire n_3906;
wire n_4138;
wire n_880;
wire n_4127;
wire n_3086;
wire n_3297;
wire n_544;
wire n_1007;
wire n_2369;
wire n_2927;
wire n_552;
wire n_1528;
wire n_4217;
wire n_4395;
wire n_2683;
wire n_1370;
wire n_1292;
wire n_2347;
wire n_2520;
wire n_2821;
wire n_1198;
wire n_1360;
wire n_2388;
wire n_1099;
wire n_4292;
wire n_2568;
wire n_3641;
wire n_4577;
wire n_956;
wire n_564;
wire n_4240;
wire n_4508;
wire n_1738;
wire n_2021;
wire n_3728;
wire n_2134;
wire n_3064;
wire n_2391;
wire n_4236;
wire n_3088;
wire n_4202;
wire n_1021;
wire n_1960;
wire n_2843;
wire n_2185;
wire n_3270;
wire n_4639;
wire n_551;
wire n_2143;
wire n_3713;
wire n_2853;
wire n_3615;
wire n_2059;
wire n_1323;
wire n_3663;
wire n_1466;
wire n_688;
wire n_1695;
wire n_2487;
wire n_3766;
wire n_1353;
wire n_800;
wire n_3595;
wire n_3246;
wire n_3202;
wire n_1347;
wire n_2495;
wire n_2880;
wire n_1535;
wire n_3813;
wire n_1789;
wire n_1666;
wire n_3350;
wire n_2389;
wire n_4165;
wire n_671;
wire n_4238;
wire n_819;
wire n_1451;
wire n_1022;
wire n_4038;
wire n_2302;
wire n_915;
wire n_4109;
wire n_1545;
wire n_2374;
wire n_864;
wire n_859;
wire n_951;
wire n_3341;
wire n_1947;
wire n_1264;
wire n_3587;
wire n_2114;
wire n_4128;
wire n_3445;
wire n_4412;
wire n_2001;
wire n_1494;
wire n_3407;
wire n_3571;
wire n_3599;
wire n_3785;
wire n_4145;
wire n_625;
wire n_854;
wire n_1462;
wire n_2069;
wire n_1799;
wire n_2396;
wire n_3621;
wire n_4211;
wire n_1580;
wire n_4734;
wire n_674;
wire n_1939;
wire n_2486;
wire n_3434;
wire n_1806;
wire n_933;
wire n_2244;
wire n_3815;
wire n_2257;
wire n_4635;
wire n_1152;
wire n_3501;
wire n_3448;
wire n_1869;
wire n_1607;
wire n_1563;
wire n_606;
wire n_3039;
wire n_3019;
wire n_2011;
wire n_2096;
wire n_4013;
wire n_4227;
wire n_4033;
wire n_4289;
wire n_877;
wire n_2105;
wire n_2538;
wire n_3776;
wire n_2024;
wire n_2530;
wire n_4242;
wire n_4517;
wire n_1696;
wire n_2483;
wire n_4780;
wire n_3163;
wire n_4425;
wire n_755;
wire n_1118;
wire n_1686;
wire n_947;
wire n_1285;
wire n_3710;
wire n_4243;
wire n_3851;
wire n_2543;
wire n_4155;
wire n_4615;
wire n_1359;
wire n_1728;
wire n_2076;
wire n_2031;
wire n_556;
wire n_1107;
wire n_3036;
wire n_2482;
wire n_3695;
wire n_3891;
wire n_2677;
wire n_1230;
wire n_4144;
wire n_668;
wire n_2165;
wire n_1896;
wire n_2147;
wire n_929;
wire n_3010;
wire n_3180;
wire n_3379;
wire n_3832;
wire n_4374;
wire n_3532;
wire n_2770;
wire n_1124;
wire n_3987;
wire n_4061;
wire n_4131;
wire n_2127;
wire n_1818;
wire n_902;
wire n_1576;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1705;
wire n_2584;
wire n_4561;
wire n_1257;
wire n_2639;
wire n_1182;
wire n_3188;
wire n_3325;
wire n_3107;
wire n_3531;
wire n_3403;
wire n_4021;
wire n_579;
wire n_1698;
wire n_3880;
wire n_1261;
wire n_2329;
wire n_938;
wire n_1098;
wire n_2963;
wire n_3624;
wire n_3834;
wire n_2142;
wire n_3186;
wire n_3461;
wire n_3082;
wire n_4548;
wire n_1154;
wire n_2189;
wire n_3796;
wire n_3332;
wire n_1242;
wire n_3283;
wire n_1135;
wire n_3048;
wire n_3258;
wire n_4501;
wire n_3937;
wire n_3696;
wire n_2323;
wire n_2203;
wire n_2597;
wire n_4525;
wire n_4622;
wire n_1016;
wire n_1243;
wire n_4315;
wire n_546;
wire n_2959;
wire n_3340;
wire n_2047;
wire n_1280;
wire n_3277;
wire n_3782;
wire n_1845;
wire n_2052;
wire n_2193;
wire n_2978;
wire n_2058;
wire n_2458;
wire n_4208;
wire n_4499;
wire n_2478;
wire n_3650;
wire n_3786;
wire n_4816;
wire n_2761;
wire n_731;
wire n_1483;
wire n_2888;
wire n_3638;
wire n_1314;
wire n_1512;
wire n_3157;
wire n_709;
wire n_1490;
wire n_1236;
wire n_1633;
wire n_4177;
wire n_2537;
wire n_2983;
wire n_3763;
wire n_569;
wire n_2669;
wire n_2144;
wire n_1778;
wire n_3214;
wire n_2306;
wire n_920;
wire n_2515;
wire n_3022;
wire n_3810;
wire n_1289;
wire n_1517;
wire n_2091;
wire n_2652;
wire n_2635;
wire n_2466;
wire n_4311;
wire n_4264;
wire n_3631;
wire n_2715;
wire n_3806;
wire n_4691;
wire n_3087;
wire n_4197;
wire n_2085;
wire n_4829;
wire n_3489;
wire n_1669;
wire n_2566;
wire n_976;
wire n_1949;
wire n_1449;
wire n_1946;
wire n_2936;
wire n_4678;
wire n_1566;
wire n_2032;
wire n_2587;
wire n_4483;
wire n_2149;
wire n_1078;
wire n_2782;
wire n_1670;
wire n_2672;
wire n_775;
wire n_3060;
wire n_4276;
wire n_2651;
wire n_3947;
wire n_4358;
wire n_3490;
wire n_3656;
wire n_600;
wire n_1484;
wire n_2071;
wire n_2643;
wire n_1374;
wire n_1328;
wire n_2561;
wire n_4715;
wire n_4793;
wire n_2141;
wire n_1948;
wire n_3013;
wire n_3183;
wire n_1984;
wire n_3437;
wire n_3868;
wire n_4369;
wire n_4543;
wire n_2099;
wire n_2408;
wire n_4168;
wire n_3446;
wire n_3353;
wire n_1877;
wire n_4203;
wire n_3687;
wire n_1831;
wire n_1598;
wire n_3049;
wire n_4394;
wire n_1723;
wire n_955;
wire n_1850;
wire n_3028;
wire n_1146;
wire n_4350;
wire n_882;
wire n_2384;
wire n_4485;
wire n_4626;
wire n_1036;
wire n_1749;
wire n_1097;
wire n_3156;
wire n_550;
wire n_696;
wire n_3101;
wire n_3669;
wire n_897;
wire n_798;
wire n_3376;
wire n_646;
wire n_1428;
wire n_2663;
wire n_1394;
wire n_4468;
wire n_2659;
wire n_3653;
wire n_1414;
wire n_1216;
wire n_580;
wire n_2693;
wire n_3798;
wire n_3702;
wire n_1040;
wire n_4065;
wire n_3836;
wire n_2202;
wire n_2648;
wire n_3963;
wire n_1872;
wire n_3389;
wire n_1852;
wire n_2159;
wire n_578;
wire n_2976;
wire n_3876;
wire n_926;
wire n_2180;
wire n_2249;
wire n_2353;
wire n_4135;
wire n_1218;
wire n_1931;
wire n_2439;
wire n_4811;
wire n_2632;
wire n_2276;
wire n_3089;
wire n_4187;
wire n_777;
wire n_1070;
wire n_1547;
wire n_4166;
wire n_2089;
wire n_3420;
wire n_1030;
wire n_2470;
wire n_1755;
wire n_3222;
wire n_1071;
wire n_1165;
wire n_1267;
wire n_1561;
wire n_1801;
wire n_3985;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_4760;
wire n_4652;
wire n_1513;
wire n_2908;
wire n_2970;
wire n_3361;
wire n_1600;
wire n_4624;
wire n_4758;
wire n_3744;
wire n_663;
wire n_845;
wire n_2235;
wire n_4263;
wire n_1862;
wire n_673;
wire n_837;
wire n_3980;
wire n_1239;
wire n_2915;
wire n_2300;
wire n_2791;
wire n_1796;
wire n_2551;
wire n_3291;
wire n_4255;
wire n_4716;
wire n_680;
wire n_1587;
wire n_1473;
wire n_2682;
wire n_553;
wire n_901;
wire n_3755;
wire n_4484;
wire n_2432;
wire n_3668;
wire n_813;
wire n_4258;
wire n_1521;
wire n_4498;
wire n_1284;
wire n_1590;
wire n_3440;
wire n_3405;
wire n_2174;
wire n_2714;
wire n_1748;
wire n_4745;
wire n_3563;
wire n_2934;
wire n_1672;
wire n_4237;
wire n_4569;
wire n_2506;
wire n_675;
wire n_2699;
wire n_4064;
wire n_888;
wire n_1880;
wire n_2769;
wire n_3542;
wire n_2337;
wire n_3436;
wire n_1167;
wire n_1626;
wire n_3550;
wire n_637;
wire n_2615;
wire n_3940;
wire n_1384;
wire n_1556;
wire n_3907;
wire n_1863;
wire n_1064;
wire n_858;
wire n_2079;
wire n_3841;
wire n_2238;
wire n_923;
wire n_2118;
wire n_691;
wire n_1151;
wire n_2985;
wire n_2944;
wire n_881;
wire n_4770;
wire n_1405;
wire n_2407;
wire n_1706;
wire n_3418;
wire n_4629;
wire n_2932;
wire n_2980;
wire n_2753;
wire n_1582;
wire n_3637;
wire n_1069;
wire n_3306;
wire n_1784;
wire n_2859;
wire n_2842;
wire n_1075;
wire n_3262;
wire n_3136;
wire n_4523;
wire n_3395;
wire n_2868;
wire n_1836;
wire n_1450;
wire n_4080;
wire n_4006;
wire n_3141;
wire n_4226;
wire n_4741;
wire n_1322;
wire n_2101;
wire n_1471;
wire n_1986;
wire n_2863;
wire n_4752;
wire n_2072;
wire n_3164;
wire n_2738;
wire n_1750;
wire n_3570;
wire n_3690;
wire n_1459;
wire n_889;
wire n_2358;
wire n_973;
wire n_3986;
wire n_4376;
wire n_4753;
wire n_3716;
wire n_4025;
wire n_2968;
wire n_1700;
wire n_2833;
wire n_4712;
wire n_3191;
wire n_571;
wire n_1585;
wire n_2712;
wire n_2684;
wire n_3837;
wire n_3593;
wire n_3193;
wire n_3885;
wire n_3936;
wire n_1971;
wire n_1599;
wire n_4552;
wire n_3252;
wire n_4421;
wire n_2275;
wire n_2855;
wire n_4503;
wire n_3507;
wire n_3273;
wire n_3821;
wire n_2713;
wire n_3544;
wire n_2644;
wire n_2700;
wire n_4310;
wire n_1211;
wire n_1197;
wire n_4836;
wire n_3367;
wire n_4464;
wire n_4020;
wire n_2951;
wire n_1523;
wire n_2730;
wire n_1950;
wire n_3008;
wire n_3709;
wire n_907;
wire n_3096;
wire n_2251;
wire n_1447;
wire n_1377;
wire n_3915;
wire n_4469;
wire n_2370;
wire n_3496;
wire n_4414;
wire n_3954;
wire n_4114;
wire n_989;
wire n_2544;
wire n_1039;
wire n_4532;
wire n_2214;
wire n_3339;
wire n_3427;
wire n_2055;
wire n_3735;
wire n_3025;
wire n_3349;
wire n_1403;
wire n_4067;
wire n_4674;
wire n_2248;
wire n_4042;
wire n_4176;
wire n_2356;
wire n_736;
wire n_892;
wire n_4385;
wire n_3320;
wire n_4556;
wire n_3007;
wire n_2688;
wire n_1000;
wire n_1202;
wire n_2750;
wire n_3899;
wire n_2620;
wire n_1278;
wire n_2622;
wire n_2062;
wire n_2668;
wire n_4159;
wire n_3714;
wire n_1002;
wire n_1581;
wire n_1463;
wire n_2100;
wire n_3071;
wire n_3739;
wire n_4089;
wire n_3651;
wire n_3310;
wire n_593;
wire n_3487;
wire n_4333;
wire n_2258;
wire n_4069;
wire n_748;
wire n_586;
wire n_1058;
wire n_1667;
wire n_3359;
wire n_838;
wire n_2784;
wire n_3718;
wire n_3983;
wire n_2919;
wire n_3092;
wire n_1053;
wire n_3470;
wire n_1224;
wire n_2865;
wire n_4327;
wire n_4405;
wire n_2557;
wire n_1926;
wire n_2706;
wire n_1248;
wire n_1331;
wire n_4195;
wire n_953;
wire n_1014;
wire n_4218;
wire n_1241;
wire n_3676;
wire n_2150;
wire n_3146;
wire n_4375;
wire n_4504;
wire n_2241;
wire n_4717;
wire n_4788;
wire n_2757;
wire n_3789;
wire n_2152;
wire n_3598;
wire n_963;
wire n_1052;
wire n_4850;
wire n_954;
wire n_627;
wire n_3781;
wire n_4813;
wire n_1385;
wire n_793;
wire n_2590;
wire n_4815;
wire n_2776;
wire n_4408;
wire n_2140;
wire n_2385;
wire n_3580;
wire n_4246;
wire n_1819;
wire n_4531;
wire n_2330;
wire n_2139;
wire n_2942;
wire n_4353;
wire n_4609;
wire n_2987;
wire n_1527;
wire n_2042;
wire n_4567;
wire n_3106;
wire n_1882;
wire n_4164;
wire n_884;
wire n_3328;
wire n_944;
wire n_4130;
wire n_1754;
wire n_4234;
wire n_3889;
wire n_3611;
wire n_1623;
wire n_2862;
wire n_4256;
wire n_2175;
wire n_2921;
wire n_2720;
wire n_2324;
wire n_1854;
wire n_2606;
wire n_2674;
wire n_3187;
wire n_1565;
wire n_4088;
wire n_4224;
wire n_3508;
wire n_2828;
wire n_3682;
wire n_4357;
wire n_3371;
wire n_1809;
wire n_1856;
wire n_4471;
wire n_4161;
wire n_4462;
wire n_4472;
wire n_647;
wire n_3433;
wire n_4024;
wire n_3392;
wire n_1072;
wire n_2267;
wire n_2218;
wire n_857;
wire n_2305;
wire n_832;
wire n_3430;
wire n_3975;
wire n_4444;
wire n_2636;
wire n_2450;
wire n_3208;
wire n_1319;
wire n_561;
wire n_2379;
wire n_3331;
wire n_3447;
wire n_2616;
wire n_2911;
wire n_3992;
wire n_3305;
wire n_2154;
wire n_1951;
wire n_1825;
wire n_4148;
wire n_4151;
wire n_1906;
wire n_1883;
wire n_4103;
wire n_2759;
wire n_1712;
wire n_4415;
wire n_1387;
wire n_4466;
wire n_3528;
wire n_3649;
wire n_2262;
wire n_4702;
wire n_4302;
wire n_2462;
wire n_2514;
wire n_4373;
wire n_1532;
wire n_4806;
wire n_4252;
wire n_2322;
wire n_4457;
wire n_2271;
wire n_2625;
wire n_3257;
wire n_3625;
wire n_4786;
wire n_1027;
wire n_971;
wire n_1156;
wire n_794;
wire n_4630;
wire n_4643;
wire n_4331;
wire n_4160;
wire n_2945;
wire n_2798;
wire n_2331;
wire n_2293;
wire n_686;
wire n_3989;
wire n_4475;
wire n_2837;
wire n_847;
wire n_3804;
wire n_4051;
wire n_4344;
wire n_4846;
wire n_1393;
wire n_2319;
wire n_4844;
wire n_596;
wire n_1775;
wire n_2979;
wire n_3296;
wire n_2028;
wire n_1368;
wire n_3481;
wire n_2762;
wire n_558;
wire n_3655;
wire n_4688;
wire n_4765;
wire n_2808;
wire n_702;
wire n_1276;
wire n_3009;
wire n_2548;
wire n_822;
wire n_1412;
wire n_2679;
wire n_2676;
wire n_1709;
wire n_3981;
wire n_4683;
wire n_2108;
wire n_3640;
wire n_728;
wire n_4491;
wire n_4388;
wire n_2930;
wire n_1162;
wire n_1538;
wire n_4206;
wire n_1838;
wire n_1199;
wire n_1847;
wire n_1779;
wire n_2767;
wire n_2777;
wire n_2603;
wire n_3514;
wire n_3116;
wire n_1884;
wire n_2434;
wire n_4132;
wire n_2660;
wire n_3602;
wire n_1038;
wire n_2967;
wire n_1369;
wire n_3909;
wire n_4738;
wire n_2611;
wire n_4261;
wire n_1841;
wire n_1660;
wire n_887;
wire n_1905;
wire n_2553;
wire n_3706;
wire n_3207;
wire n_2581;
wire n_3944;
wire n_2195;
wire n_2529;
wire n_3224;
wire n_2698;
wire n_3752;
wire n_4090;
wire n_4647;
wire n_809;
wire n_3923;
wire n_870;
wire n_931;
wire n_599;
wire n_1891;
wire n_1711;
wire n_1662;
wire n_1481;
wire n_2626;
wire n_3441;
wire n_3042;
wire n_4696;
wire n_4837;
wire n_1942;
wire n_1978;
wire n_1544;
wire n_4001;
wire n_2510;
wire n_3047;
wire n_3526;
wire n_4219;
wire n_868;
wire n_2454;
wire n_4371;
wire n_639;
wire n_2804;
wire n_914;
wire n_3659;
wire n_2120;
wire n_2546;
wire n_1629;
wire n_1293;
wire n_2801;
wire n_3120;
wire n_4473;
wire n_965;
wire n_1876;
wire n_1743;
wire n_4007;
wire n_4620;
wire n_3790;
wire n_4011;
wire n_4268;
wire n_3491;
wire n_935;
wire n_1175;
wire n_2763;
wire n_817;
wire n_4613;
wire n_1479;
wire n_1810;
wire n_4480;
wire n_4649;
wire n_2350;
wire n_2813;
wire n_2825;
wire n_2009;
wire n_1888;
wire n_759;
wire n_3643;
wire n_3895;
wire n_4194;
wire n_2222;
wire n_4438;
wire n_4824;
wire n_1892;
wire n_4120;
wire n_3510;
wire n_4427;
wire n_3745;
wire n_806;
wire n_2990;
wire n_1997;
wire n_2667;
wire n_1766;
wire n_3218;
wire n_3748;
wire n_1477;
wire n_3142;
wire n_4278;
wire n_1635;
wire n_1963;
wire n_4795;
wire n_2226;
wire n_1571;
wire n_2891;
wire n_3119;
wire n_4623;
wire n_4142;
wire n_1189;
wire n_2690;
wire n_4028;
wire n_4082;
wire n_4410;
wire n_3370;
wire n_1860;
wire n_2215;
wire n_3479;
wire n_4085;
wire n_1259;
wire n_4073;
wire n_1690;
wire n_4260;
wire n_4553;
wire n_3819;
wire n_706;
wire n_746;
wire n_1649;
wire n_3150;
wire n_4163;
wire n_747;
wire n_4439;
wire n_2064;
wire n_784;
wire n_3978;
wire n_4325;
wire n_4832;
wire n_2449;
wire n_3867;
wire n_1733;
wire n_4809;
wire n_4372;
wire n_1244;
wire n_3500;
wire n_2413;
wire n_1194;
wire n_1925;
wire n_3660;
wire n_2297;
wire n_4186;
wire n_1815;
wire n_3279;
wire n_2621;
wire n_615;
wire n_851;
wire n_4731;
wire n_1759;
wire n_843;
wire n_1788;
wire n_2491;
wire n_2177;
wire n_3747;
wire n_913;
wire n_1537;
wire n_705;
wire n_3833;
wire n_865;
wire n_2227;
wire n_3775;
wire n_4133;
wire n_678;
wire n_2671;
wire n_697;
wire n_4262;
wire n_4184;
wire n_4618;
wire n_1222;
wire n_1679;
wire n_2190;
wire n_3346;
wire n_4742;
wire n_4841;
wire n_776;
wire n_2022;
wire n_1798;
wire n_3814;
wire n_1790;
wire n_2518;
wire n_4585;
wire n_2876;
wire n_4720;
wire n_1415;
wire n_2629;
wire n_4099;
wire n_4481;
wire n_2592;
wire n_3416;
wire n_4379;
wire n_3484;
wire n_3620;
wire n_1260;
wire n_1746;
wire n_1647;
wire n_2181;
wire n_2479;
wire n_2838;
wire n_4842;
wire n_4340;
wire n_1829;
wire n_1464;
wire n_3133;
wire n_3513;
wire n_4295;
wire n_4685;
wire n_649;
wire n_547;
wire n_2563;
wire n_1444;
wire n_4030;
wire n_1191;
wire n_4645;
wire n_2387;
wire n_2992;
wire n_4334;
wire n_1674;
wire n_3725;
wire n_1833;
wire n_4490;
wire n_3138;
wire n_1830;
wire n_2517;
wire n_4397;
wire n_2073;
wire n_1710;
wire n_1128;
wire n_4511;
wire n_2928;
wire n_3128;
wire n_4694;
wire n_1734;
wire n_4533;
wire n_3038;
wire n_4820;
wire n_744;
wire n_629;
wire n_590;
wire n_3770;
wire n_4014;
wire n_2631;
wire n_1308;
wire n_3068;
wire n_2178;
wire n_2871;
wire n_1767;
wire n_3144;
wire n_4244;
wire n_4757;
wire n_4603;
wire n_2943;
wire n_2913;
wire n_4254;
wire n_2336;
wire n_3143;
wire n_3168;
wire n_1680;
wire n_4697;
wire n_1233;
wire n_4179;
wire n_3469;
wire n_2607;
wire n_3994;
wire n_4190;
wire n_1615;
wire n_4175;
wire n_4810;
wire n_1529;
wire n_2005;
wire n_1916;
wire n_3317;
wire n_677;
wire n_4648;
wire n_1333;
wire n_2469;
wire n_1121;
wire n_2723;
wire n_3355;
wire n_604;
wire n_2007;
wire n_3220;
wire n_4641;
wire n_4391;
wire n_949;
wire n_2539;
wire n_3917;
wire n_3942;
wire n_3263;
wire n_2582;
wire n_1443;
wire n_1008;
wire n_3855;
wire n_946;
wire n_1539;
wire n_2736;
wire n_4157;
wire n_4283;
wire n_4681;
wire n_1001;
wire n_1503;
wire n_2054;
wire n_3765;
wire n_4638;
wire n_1468;
wire n_1559;
wire n_3823;
wire n_1765;
wire n_3455;
wire n_1866;
wire n_4173;
wire n_689;
wire n_3158;
wire n_738;
wire n_1624;
wire n_3000;
wire n_640;
wire n_3452;
wire n_1510;
wire n_624;
wire n_1380;
wire n_1744;
wire n_3816;
wire n_2623;
wire n_1617;
wire n_1010;
wire n_1994;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_3108;
wire n_3113;
wire n_3111;
wire n_2718;
wire n_1195;
wire n_1839;
wire n_1837;
wire n_2577;
wire n_610;
wire n_3760;
wire n_4108;
wire n_4486;
wire n_4557;
wire n_4707;
wire n_4078;
wire n_4451;
wire n_1760;
wire n_2875;
wire n_936;
wire n_568;
wire n_1500;
wire n_2960;
wire n_1090;
wire n_2796;
wire n_4527;
wire n_757;
wire n_3844;
wire n_3280;
wire n_2342;
wire n_633;
wire n_2856;
wire n_4054;
wire n_3471;
wire n_1832;
wire n_4627;
wire n_1851;
wire n_758;
wire n_999;
wire n_3205;
wire n_4156;
wire n_4848;
wire n_2046;
wire n_4146;
wire n_2848;
wire n_2741;
wire n_4360;
wire n_2937;
wire n_3666;
wire n_3003;
wire n_3610;
wire n_1933;
wire n_3828;
wire n_2290;
wire n_1656;
wire n_3564;
wire n_3288;
wire n_1158;
wire n_3095;
wire n_4404;
wire n_2045;
wire n_3369;
wire n_3783;
wire n_3988;
wire n_1509;
wire n_1874;
wire n_2040;
wire n_563;
wire n_4787;
wire n_2060;
wire n_3199;
wire n_2613;
wire n_2805;
wire n_1987;
wire n_3667;
wire n_1145;
wire n_878;
wire n_4541;
wire n_3843;
wire n_3457;
wire n_1678;
wire n_1049;
wire n_1153;
wire n_3856;
wire n_2145;
wire n_741;
wire n_1639;
wire n_1306;
wire n_3703;
wire n_4324;
wire n_1068;
wire n_3030;
wire n_3558;
wire n_4821;
wire n_1871;
wire n_2580;
wire n_3630;
wire n_2545;
wire n_2787;
wire n_3685;
wire n_4249;
wire n_2914;
wire n_1964;
wire n_2869;
wire n_4002;
wire n_1163;
wire n_906;
wire n_3271;
wire n_4771;
wire n_2039;
wire n_1207;
wire n_919;
wire n_908;
wire n_4086;
wire n_2412;
wire n_4356;
wire n_2406;
wire n_4814;
wire n_3623;
wire n_2846;
wire n_724;
wire n_3753;
wire n_1781;
wire n_2084;
wire n_2925;
wire n_3648;
wire n_2035;
wire n_658;
wire n_2061;
wire n_3773;
wire n_4718;
wire n_3555;
wire n_3579;
wire n_3918;
wire n_3075;
wire n_3173;
wire n_4432;
wire n_2378;
wire n_2509;
wire n_1740;
wire n_3236;
wire n_2398;
wire n_1362;
wire n_4317;
wire n_3969;
wire n_2857;
wire n_4528;
wire n_3932;
wire n_1586;
wire n_4291;
wire n_959;
wire n_2459;
wire n_3031;
wire n_4692;
wire n_4154;
wire n_4619;
wire n_4673;
wire n_3396;
wire n_3701;
wire n_940;
wire n_4386;
wire n_1445;
wire n_3516;
wire n_4023;
wire n_4149;
wire n_4822;
wire n_1492;
wire n_2155;
wire n_2516;
wire n_3797;
wire n_1923;
wire n_4420;
wire n_1773;
wire n_592;
wire n_3243;
wire n_1169;
wire n_1596;
wire n_1692;
wire n_2666;
wire n_2982;
wire n_3385;
wire n_1017;
wire n_2481;
wire n_2947;
wire n_3545;
wire n_2171;
wire n_4708;
wire n_978;
wire n_2768;
wire n_4299;
wire n_2116;
wire n_2314;
wire n_1434;
wire n_4801;
wire n_1054;
wire n_2507;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_4019;
wire n_4826;
wire n_2420;
wire n_2900;
wire n_1095;
wire n_3343;
wire n_3515;
wire n_1828;
wire n_1614;
wire n_2886;
wire n_2093;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_2339;
wire n_2038;
wire n_2320;
wire n_2473;
wire n_3287;
wire n_4637;
wire n_2137;
wire n_3378;
wire n_603;
wire n_4640;
wire n_1431;
wire n_2583;
wire n_1593;
wire n_1033;
wire n_3767;
wire n_4279;
wire n_4769;
wire n_4785;
wire n_4396;
wire n_3426;
wire n_3454;
wire n_2299;
wire n_2540;
wire n_2873;
wire n_3820;
wire n_636;
wire n_4589;
wire n_4632;
wire n_4367;
wire n_3741;
wire n_660;
wire n_3410;
wire n_4578;
wire n_2087;
wire n_1640;
wire n_4294;
wire n_2162;
wire n_1732;
wire n_1009;
wire n_2847;
wire n_1148;
wire n_2051;
wire n_3221;
wire n_742;
wire n_750;
wire n_2029;
wire n_995;
wire n_4125;
wire n_2168;
wire n_2790;
wire n_1609;
wire n_4232;
wire n_3629;
wire n_3021;
wire n_1989;
wire n_3818;
wire n_2359;
wire n_2941;
wire n_3674;
wire n_1887;
wire n_4413;
wire n_3502;
wire n_2523;
wire n_1383;
wire n_3098;
wire n_1073;
wire n_2457;
wire n_2346;
wire n_4387;
wire n_662;
wire n_2312;
wire n_3990;
wire n_4493;
wire n_4790;
wire n_962;
wire n_3475;
wire n_1215;
wire n_3015;
wire n_4453;
wire n_4170;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1920;
wire n_1065;
wire n_1592;
wire n_2536;
wire n_1336;
wire n_2882;
wire n_3719;
wire n_1721;
wire n_1959;
wire n_1758;
wire n_2338;
wire n_3681;
wire n_2952;
wire n_2737;
wire n_1574;
wire n_3672;
wire n_4847;
wire n_2399;
wire n_3058;
wire n_4147;
wire n_4308;
wire n_2812;
wire n_2048;
wire n_3197;
wire n_3109;
wire n_3607;
wire n_2355;
wire n_2133;
wire n_4365;
wire n_1921;
wire n_2721;
wire n_1309;
wire n_1878;
wire n_1426;
wire n_3830;
wire n_1043;
wire n_2585;
wire n_3505;
wire n_3002;
wire n_1800;
wire n_1548;
wire n_2725;
wire n_614;
wire n_1421;
wire n_4510;
wire n_4610;
wire n_2571;
wire n_1286;
wire n_3730;
wire n_3883;
wire n_4489;
wire n_1177;
wire n_3276;
wire n_1355;
wire n_974;
wire n_2565;
wire n_4152;
wire n_727;
wire n_3897;
wire n_1159;
wire n_3845;
wire n_957;
wire n_3787;
wire n_773;
wire n_2124;
wire n_743;
wire n_3001;
wire n_2081;
wire n_3945;
wire n_4392;
wire n_4660;
wire n_3149;
wire n_4570;
wire n_4542;
wire n_613;
wire n_1119;
wire n_2261;
wire n_1240;
wire n_2156;
wire n_1820;
wire n_2729;
wire n_3268;
wire n_3597;
wire n_4296;
wire n_2418;
wire n_3827;
wire n_829;
wire n_2519;
wire n_3354;
wire n_4281;
wire n_2724;
wire n_4661;
wire n_4447;
wire n_1612;
wire n_2179;
wire n_4200;
wire n_1416;
wire n_2077;
wire n_2897;
wire n_3614;
wire n_4198;
wire n_2909;
wire n_1724;
wire n_2111;
wire n_2521;
wire n_3301;
wire n_4285;
wire n_4651;
wire n_3466;
wire n_4534;
wire n_4500;
wire n_3458;
wire n_1237;
wire n_700;
wire n_573;
wire n_1420;
wire n_3185;
wire n_1132;
wire n_3330;
wire n_4818;
wire n_4514;
wire n_1366;
wire n_4606;
wire n_4800;
wire n_1300;
wire n_3960;
wire n_4774;
wire n_2595;
wire n_1127;
wire n_3248;
wire n_2477;
wire n_761;
wire n_2277;
wire n_3523;
wire n_1785;
wire n_1568;
wire n_2829;
wire n_4597;
wire n_3905;
wire n_4329;
wire n_1006;
wire n_3411;
wire n_3887;
wire n_4087;
wire n_2110;
wire n_3811;
wire n_4093;
wire n_1270;
wire n_1664;
wire n_3200;
wire n_4271;
wire n_1486;
wire n_582;
wire n_3586;
wire n_4672;
wire n_1332;
wire n_3519;
wire n_4433;
wire n_2231;
wire n_1390;
wire n_4682;
wire n_2017;
wire n_2474;
wire n_2879;
wire n_2604;
wire n_4174;
wire n_2090;
wire n_3374;
wire n_3153;
wire n_3045;
wire n_2367;
wire n_1870;
wire n_1591;
wire n_2033;
wire n_4071;
wire n_4330;
wire n_4341;
wire n_4257;
wire n_4766;
wire n_3453;
wire n_1682;
wire n_1980;
wire n_2628;
wire n_2390;
wire n_1249;
wire n_3399;
wire n_4312;
wire n_2896;
wire n_652;
wire n_1111;
wire n_3213;
wire n_1365;
wire n_4074;
wire n_4600;
wire n_1927;
wire n_3065;
wire n_4361;
wire n_2132;
wire n_1349;
wire n_1093;
wire n_4460;
wire n_2400;
wire n_4633;
wire n_1031;
wire n_3645;
wire n_4614;
wire n_609;
wire n_1041;
wire n_1265;
wire n_3223;
wire n_1909;
wire n_3838;
wire n_3929;
wire n_3077;
wire n_4277;
wire n_2681;
wire n_1562;
wire n_3103;
wire n_834;
wire n_3474;
wire n_765;
wire n_4140;
wire n_3675;
wire n_2255;
wire n_2424;
wire n_4732;
wire n_2272;
wire n_893;
wire n_3984;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_1965;
wire n_3387;
wire n_630;
wire n_1902;
wire n_2151;
wire n_1941;
wire n_2106;
wire n_2775;
wire n_2716;
wire n_3938;
wire n_4665;
wire n_1913;
wire n_2878;
wire n_4693;
wire n_1823;
wire n_4434;
wire n_4662;
wire n_3679;
wire n_3779;
wire n_874;
wire n_2464;
wire n_3422;
wire n_3888;
wire n_1101;
wire n_2831;
wire n_1106;
wire n_4326;
wire n_1456;
wire n_3557;
wire n_2230;
wire n_3498;
wire n_4189;
wire n_2015;
wire n_2365;
wire n_1875;
wire n_1982;
wire n_4744;
wire n_4110;
wire n_1304;
wire n_2803;
wire n_1324;
wire n_2851;
wire n_3707;
wire n_987;
wire n_4207;
wire n_3189;
wire n_1846;
wire n_3037;
wire n_4305;
wire n_4545;
wire n_2066;
wire n_1885;
wire n_1455;
wire n_3429;
wire n_767;
wire n_993;
wire n_1903;
wire n_2490;
wire n_1407;
wire n_3849;
wire n_3946;
wire n_2452;
wire n_1551;
wire n_3154;
wire n_545;
wire n_3229;
wire n_860;
wire n_4213;
wire n_4463;
wire n_2849;
wire n_1805;
wire n_3925;
wire n_2176;
wire n_2204;
wire n_2905;
wire n_1816;
wire n_3692;
wire n_4687;
wire n_948;
wire n_3965;
wire n_3566;
wire n_1217;
wire n_2220;
wire n_4059;
wire n_2455;
wire n_4349;
wire n_4595;
wire n_628;
wire n_1849;
wire n_3788;
wire n_4670;
wire n_4084;
wire n_4703;
wire n_2410;
wire n_729;
wire n_1131;
wire n_1084;
wire n_1961;
wire n_4313;
wire n_970;
wire n_4037;
wire n_1935;
wire n_911;
wire n_2922;
wire n_1430;
wire n_3275;
wire n_3499;
wire n_2645;
wire n_4802;
wire n_2467;
wire n_3366;
wire n_2727;
wire n_1094;
wire n_1534;
wire n_560;
wire n_1354;
wire n_2288;
wire n_3421;
wire n_4139;
wire n_1351;
wire n_2696;
wire n_2240;
wire n_4063;
wire n_4428;
wire n_1205;
wire n_1044;
wire n_2436;
wire n_1209;
wire n_3029;
wire n_3242;
wire n_1552;
wire n_2508;
wire n_3592;
wire n_3618;
wire n_4031;
wire n_4650;
wire n_602;
wire n_3525;
wire n_574;
wire n_2593;
wire n_3486;
wire n_1435;
wire n_879;
wire n_3394;
wire n_3793;
wire n_3683;
wire n_2416;
wire n_2405;
wire n_3642;
wire n_623;
wire n_3995;
wire n_4669;
wire n_3286;
wire n_2088;
wire n_2953;
wire n_3808;
wire n_824;
wire n_4036;
wire n_1645;
wire n_3881;
wire n_4339;
wire n_4041;
wire n_2461;
wire n_1327;
wire n_2858;
wire n_2243;
wire n_4583;
wire n_4060;
wire n_996;
wire n_1684;
wire n_2658;
wire n_921;
wire n_3590;
wire n_1717;
wire n_4763;
wire n_572;
wire n_2895;
wire n_815;
wire n_1795;
wire n_2128;
wire n_4210;
wire n_2578;
wire n_4594;
wire n_3097;
wire n_3483;
wire n_1821;
wire n_3894;
wire n_4666;
wire n_2929;
wire n_3424;
wire n_3478;
wire n_1381;
wire n_2555;
wire n_4015;
wire n_2662;
wire n_2740;
wire n_3824;
wire n_3751;
wire n_1611;
wire n_1037;
wire n_2368;
wire n_3890;
wire n_3388;
wire n_2656;
wire n_1080;
wire n_2301;
wire n_1274;
wire n_3583;
wire n_4494;
wire n_2890;
wire n_3560;
wire n_3059;
wire n_3524;
wire n_4076;
wire n_2554;
wire n_4714;
wire n_3465;
wire n_1316;
wire n_1708;
wire n_2419;
wire n_3215;
wire n_4796;
wire n_1438;
wire n_3698;
wire n_3927;
wire n_1082;
wire n_1840;
wire n_589;
wire n_3961;
wire n_716;
wire n_1630;
wire n_2122;
wire n_2512;
wire n_3589;
wire n_4540;
wire n_4102;
wire n_4776;
wire n_562;
wire n_1436;
wire n_3549;
wire n_1691;
wire n_952;
wire n_2786;
wire n_2534;
wire n_2092;
wire n_3171;
wire n_1229;
wire n_4799;
wire n_701;
wire n_1437;
wire n_1023;
wire n_2075;
wire n_645;
wire n_3658;
wire n_3449;
wire n_803;
wire n_1092;
wire n_2694;
wire n_1776;
wire n_3559;
wire n_4807;
wire n_2198;
wire n_2610;
wire n_2661;
wire n_2572;
wire n_2989;
wire n_2281;
wire n_2131;
wire n_2789;
wire n_3026;
wire n_4775;
wire n_3993;
wire n_2216;
wire n_3020;
wire n_3677;
wire n_1757;
wire n_890;
wire n_1897;
wire n_764;
wire n_1919;
wire n_1056;
wire n_1424;
wire n_960;
wire n_3588;
wire n_3462;
wire n_2933;
wire n_4230;
wire n_2308;
wire n_3468;
wire n_4590;
wire n_1893;
wire n_2910;
wire n_3419;
wire n_4381;
wire n_4266;
wire n_3886;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_4455;
wire n_2053;
wire n_2163;
wire n_4830;
wire n_634;
wire n_2328;
wire n_1958;
wire n_4664;
wire n_2254;
wire n_1252;
wire n_3860;
wire n_1382;
wire n_1029;
wire n_925;
wire n_3546;
wire n_1206;
wire n_4248;
wire n_2647;
wire n_3784;
wire n_3160;
wire n_2969;
wire n_2191;
wire n_1311;
wire n_2864;
wire n_3941;
wire n_4754;
wire n_3195;
wire n_1519;
wire n_3190;
wire n_950;
wire n_2428;
wire n_1553;
wire n_3678;
wire n_4443;
wire n_3847;
wire n_2664;
wire n_4507;
wire n_4554;
wire n_1811;
wire n_2443;
wire n_2624;
wire n_3012;
wire n_3456;
wire n_4575;
wire n_4845;
wire n_1346;
wire n_3053;
wire n_1299;
wire n_3244;
wire n_2158;
wire n_1808;
wire n_3893;
wire n_3290;
wire n_4663;
wire n_1060;
wire n_1141;
wire n_2266;
wire n_3130;
wire n_2824;
wire n_2465;
wire n_3033;
wire n_2650;
wire n_3298;
wire n_3569;
wire n_912;
wire n_968;
wire n_3548;
wire n_4452;
wire n_4348;
wire n_619;
wire n_2440;
wire n_1386;
wire n_1699;
wire n_3334;
wire n_967;
wire n_2923;
wire n_4162;
wire n_1442;
wire n_3665;
wire n_4355;
wire n_3494;
wire n_2541;
wire n_4383;
wire n_2731;
wire n_1139;
wire n_3264;
wire n_2333;
wire n_3953;
wire n_2916;
wire n_3166;
wire n_885;
wire n_1432;
wire n_3875;
wire n_3976;
wire n_4122;
wire n_1357;
wire n_2125;
wire n_3771;
wire n_3979;
wire n_4297;
wire n_683;
wire n_3110;
wire n_1632;
wire n_4582;
wire n_2998;
wire n_1057;
wire n_4684;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_4003;
wire n_3800;
wire n_721;
wire n_2402;
wire n_1157;
wire n_3073;
wire n_2403;
wire n_4301;
wire n_4572;
wire n_841;
wire n_1050;
wire n_4586;
wire n_802;
wire n_1954;
wire n_4048;
wire n_4608;
wire n_4840;
wire n_4026;
wire n_2265;
wire n_3162;
wire n_1608;
wire n_983;
wire n_1844;
wire n_4104;
wire n_4512;
wire n_2760;
wire n_2792;
wire n_3554;
wire n_3377;
wire n_2870;
wire n_3777;
wire n_4377;
wire n_1305;
wire n_3749;
wire n_3178;
wire n_873;
wire n_1826;
wire n_3962;
wire n_3991;
wire n_4784;
wire n_1112;
wire n_3134;
wire n_2999;
wire n_2304;
wire n_762;
wire n_1283;
wire n_1644;
wire n_4172;
wire n_2637;
wire n_2334;
wire n_4791;
wire n_4384;
wire n_4536;
wire n_690;
wire n_4046;
wire n_1974;
wire n_2463;
wire n_4521;
wire n_583;
wire n_4488;
wire n_2086;
wire n_3537;
wire n_4423;
wire n_4773;
wire n_2289;
wire n_3080;
wire n_3051;
wire n_4096;
wire n_4199;
wire n_1343;
wire n_2701;
wire n_2783;
wire n_4497;
wire n_2263;
wire n_3362;
wire n_2881;
wire n_1203;
wire n_1631;
wire n_3750;
wire n_3282;
wire n_2472;
wire n_821;
wire n_4611;
wire n_1763;
wire n_4755;
wire n_2341;
wire n_3105;
wire n_3231;
wire n_1966;
wire n_3632;
wire n_1768;
wire n_2294;
wire n_1179;
wire n_4588;
wire n_621;
wire n_753;
wire n_2475;
wire n_2733;
wire n_1048;
wire n_1719;
wire n_2993;
wire n_4598;
wire n_3864;
wire n_1288;
wire n_4286;
wire n_4478;
wire n_2785;
wire n_4658;
wire n_2556;
wire n_2269;
wire n_2732;
wire n_2309;
wire n_2415;
wire n_2948;
wire n_3274;
wire n_3041;
wire n_3299;
wire n_4519;
wire n_2646;
wire n_1560;
wire n_3715;
wire n_1605;
wire n_4362;
wire n_2236;
wire n_4470;
wire n_1228;
wire n_2816;
wire n_4306;
wire n_2123;
wire n_3209;
wire n_972;
wire n_3504;
wire n_692;
wire n_2685;
wire n_2037;
wire n_3920;
wire n_3040;
wire n_1953;
wire n_1938;
wire n_820;
wire n_1200;
wire n_2499;
wire n_4422;
wire n_1911;
wire n_3616;
wire n_2460;
wire n_4058;
wire n_3568;
wire n_3664;
wire n_2589;
wire n_3203;
wire n_1363;
wire n_1301;
wire n_1668;
wire n_3737;
wire n_3913;
wire n_1185;
wire n_991;
wire n_2903;
wire n_3417;
wire n_3482;
wire n_3866;
wire n_828;
wire n_1967;
wire n_779;
wire n_576;
wire n_1143;
wire n_1579;
wire n_2233;
wire n_3717;
wire n_4106;
wire n_4034;
wire n_1329;
wire n_2743;
wire n_2675;
wire n_3255;
wire n_1312;
wire n_1439;
wire n_804;
wire n_4555;
wire n_3052;
wire n_1688;
wire n_2827;
wire n_945;
wire n_2997;
wire n_3743;
wire n_3327;
wire n_1504;
wire n_4400;
wire n_943;
wire n_3326;
wire n_4689;
wire n_3956;
wire n_3572;
wire n_992;
wire n_3067;
wire n_4215;
wire n_1932;
wire n_4280;
wire n_3375;
wire n_2755;
wire n_4721;
wire n_4047;
wire n_842;
wire n_3734;
wire n_650;
wire n_984;
wire n_694;
wire n_3237;
wire n_2082;
wire n_4778;
wire n_1992;
wire n_2429;
wire n_1643;
wire n_1983;
wire n_883;
wire n_4402;
wire n_3167;
wire n_4239;
wire n_4029;
wire n_3400;
wire n_1594;
wire n_4550;
wire n_1214;
wire n_1400;
wire n_1342;
wire n_3423;
wire n_900;
wire n_2362;
wire n_856;
wire n_2609;
wire n_3870;
wire n_1793;
wire n_3382;
wire n_1976;
wire n_2223;
wire n_3044;
wire n_3574;
wire n_4352;
wire n_4441;
wire n_4496;
wire n_918;
wire n_4761;
wire n_3529;
wire n_3854;
wire n_942;
wire n_2169;
wire n_1804;
wire n_1977;
wire n_1557;
wire n_2468;
wire n_2153;
wire n_1147;
wire n_4201;
wire n_1610;
wire n_4347;
wire n_1077;
wire n_1422;
wire n_3196;
wire n_4095;
wire n_3078;
wire n_4593;
wire n_2533;
wire n_2364;
wire n_4338;
wire n_3492;
wire n_618;
wire n_3094;
wire n_896;
wire n_2310;
wire n_2780;
wire n_4727;
wire n_3952;
wire n_4568;
wire n_2287;
wire n_2860;
wire n_3316;
wire n_2291;
wire n_3099;
wire n_4043;
wire n_3704;
wire n_2596;
wire n_894;
wire n_1636;
wire n_2056;
wire n_3253;
wire n_1730;
wire n_3601;
wire n_3603;
wire n_4027;
wire n_831;
wire n_2280;
wire n_4123;
wire n_2192;
wire n_4599;
wire n_964;
wire n_3633;
wire n_3363;
wire n_4479;
wire n_1373;
wire n_4812;
wire n_1350;
wire n_1511;
wire n_1865;
wire n_2973;
wire n_1470;
wire n_2094;
wire n_2670;
wire n_1096;
wire n_1575;
wire n_1735;
wire n_1697;
wire n_2318;
wire n_833;
wire n_2393;
wire n_3689;
wire n_2020;
wire n_4628;
wire n_3831;
wire n_1646;
wire n_2502;
wire n_3801;
wire n_2504;
wire n_1307;
wire n_4495;
wire n_4762;
wire n_1881;
wire n_4416;
wire n_2974;
wire n_988;
wire n_2749;
wire n_2043;
wire n_2901;
wire n_1940;
wire n_814;
wire n_2751;
wire n_2707;
wire n_2793;
wire n_3372;
wire n_3451;
wire n_4539;
wire n_2971;
wire n_4657;
wire n_3442;
wire n_1549;
wire n_1934;
wire n_2311;
wire n_1201;
wire n_1114;
wire n_3950;
wire n_4000;
wire n_655;
wire n_4458;
wire n_3240;
wire n_2025;
wire n_1616;
wire n_4121;
wire n_3998;
wire n_1446;
wire n_2285;
wire n_4406;
wire n_3147;
wire n_2758;
wire n_4141;
wire n_1458;
wire n_669;
wire n_2471;
wire n_1176;
wire n_1472;
wire n_2298;
wire n_4476;
wire n_1807;
wire n_4756;
wire n_3869;
wire n_4307;
wire n_1149;
wire n_2618;
wire n_4359;
wire n_1671;
wire n_635;
wire n_2559;
wire n_763;
wire n_3230;
wire n_1020;
wire n_1062;
wire n_3342;
wire n_4748;
wire n_2303;
wire n_1824;
wire n_1917;
wire n_2295;
wire n_1219;
wire n_3386;
wire n_3931;
wire n_3708;
wire n_1204;
wire n_4010;
wire n_4107;
wire n_2840;
wire n_4667;
wire n_3729;
wire n_2810;
wire n_2325;
wire n_2747;
wire n_2446;
wire n_3488;
wire n_4690;
wire n_1814;
wire n_1035;
wire n_2822;
wire n_4437;
wire n_4710;
wire n_3861;
wire n_4736;
wire n_3780;
wire n_555;
wire n_783;
wire n_1928;
wire n_1848;
wire n_4607;
wire n_2126;
wire n_4547;
wire n_4117;
wire n_2893;
wire n_4573;
wire n_3636;
wire n_1188;
wire n_2588;
wire n_2962;
wire n_4004;
wire n_4118;
wire n_1722;
wire n_3957;
wire n_661;
wire n_4803;
wire n_2441;
wire n_3848;
wire n_1802;
wire n_3083;
wire n_4284;
wire n_4668;
wire n_2600;
wire n_4487;
wire n_3919;
wire n_4079;
wire n_3898;
wire n_849;
wire n_2795;
wire n_4091;
wire n_584;
wire n_681;
wire n_1638;
wire n_1786;
wire n_2981;
wire n_2282;
wire n_2002;
wire n_3608;
wire n_2800;
wire n_3712;
wire n_4817;
wire n_2371;
wire n_2935;
wire n_4513;
wire n_3233;
wire n_3829;
wire n_3380;
wire n_3177;
wire n_4053;
wire n_830;
wire n_4274;
wire n_2098;
wire n_1296;
wire n_2627;
wire n_3409;
wire n_3460;
wire n_2352;
wire n_4759;
wire n_3538;
wire n_1413;
wire n_801;
wire n_4040;
wire n_2207;
wire n_4467;
wire n_2080;
wire n_2377;
wire n_2619;
wire n_3085;
wire n_2340;
wire n_2444;
wire n_2068;
wire n_3552;
wire n_4849;
wire n_875;
wire n_1110;
wire n_4474;
wire n_1655;
wire n_2641;
wire n_3198;
wire n_749;
wire n_1895;
wire n_3123;
wire n_3684;
wire n_4735;
wire n_3137;
wire n_2574;
wire n_1134;
wire n_1358;
wire n_717;
wire n_4728;
wire n_4316;
wire n_939;
wire n_3697;
wire n_2361;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_3393;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_4247;
wire n_2638;
wire n_866;
wire n_969;
wire n_1401;
wire n_4018;
wire n_4044;
wire n_3900;
wire n_4617;
wire n_4062;
wire n_4524;
wire n_4113;
wire n_3520;
wire n_3971;
wire n_4843;
wire n_2492;
wire n_1019;
wire n_1998;
wire n_1105;
wire n_4686;
wire n_4518;
wire n_3759;
wire n_1338;
wire n_577;
wire n_4409;
wire n_4411;
wire n_4005;
wire n_2016;
wire n_1522;
wire n_4321;
wire n_4342;
wire n_3872;
wire n_2949;
wire n_1687;
wire n_1637;
wire n_2034;
wire n_1419;
wire n_2711;
wire n_4631;
wire n_4336;
wire n_3933;
wire n_1653;
wire n_693;
wire n_2270;
wire n_1506;
wire n_3206;
wire n_4777;
wire n_4792;
wire n_2653;
wire n_3578;
wire n_3966;
wire n_990;
wire n_836;
wire n_2867;
wire n_3812;
wire n_2496;
wire n_1886;
wire n_1389;
wire n_1894;
wire n_975;
wire n_1908;
wire n_1256;
wire n_1702;
wire n_2259;
wire n_2794;
wire n_567;
wire n_1465;
wire n_3145;
wire n_4183;
wire n_3124;
wire n_778;
wire n_1122;
wire n_4068;
wire n_4253;
wire n_4290;
wire n_4233;
wire n_3192;
wire n_2608;
wire n_3877;
wire n_3764;
wire n_2657;
wire n_770;
wire n_4709;
wire n_2995;
wire n_1375;
wire n_2494;
wire n_3547;
wire n_2649;
wire n_3977;
wire n_1102;
wire n_3727;
wire n_2852;
wire n_3774;
wire n_4052;
wire n_2392;
wire n_3459;
wire n_3093;
wire n_1843;
wire n_711;
wire n_1499;
wire n_3061;
wire n_4398;
wire n_3155;
wire n_1187;
wire n_3517;
wire n_2633;
wire n_1441;
wire n_3100;
wire n_2522;
wire n_2435;
wire n_1597;
wire n_1929;
wire n_1392;
wire n_2807;
wire n_1164;
wire n_1659;
wire n_2097;
wire n_2542;
wire n_2313;
wire n_1834;
wire n_1174;
wire n_2431;
wire n_3356;
wire n_3324;
wire n_3914;
wire n_2835;
wire n_3758;
wire n_4304;
wire n_3911;
wire n_4625;
wire n_2558;
wire n_1371;
wire n_617;
wire n_1303;
wire n_2206;
wire n_2063;
wire n_3803;
wire n_3182;
wire n_4431;
wire n_1572;
wire n_1968;
wire n_4192;
wire n_3742;
wire n_3269;
wire n_2564;
wire n_2252;
wire n_876;
wire n_1516;
wire n_3736;
wire n_4656;
wire n_4805;
wire n_1190;
wire n_3506;
wire n_3896;
wire n_1736;
wire n_3605;
wire n_1685;
wire n_3958;
wire n_4819;
wire n_2409;
wire n_601;
wire n_917;
wire n_3450;
wire n_1714;
wire n_966;
wire n_4729;
wire n_1116;
wire n_2000;
wire n_1661;
wire n_3402;
wire n_1212;
wire n_2074;
wire n_1541;
wire n_2576;
wire n_3565;
wire n_4679;
wire n_4115;
wire n_726;
wire n_3174;
wire n_982;
wire n_4701;
wire n_2575;
wire n_2988;
wire n_3390;
wire n_1573;
wire n_1453;
wire n_1731;
wire n_2217;
wire n_3746;
wire n_818;
wire n_2373;
wire n_1970;
wire n_861;
wire n_1713;
wire n_1183;
wire n_3398;
wire n_2307;
wire n_2766;
wire n_3817;
wire n_1658;
wire n_899;
wire n_1253;
wire n_2722;
wire n_1737;
wire n_2745;
wire n_2201;
wire n_2117;
wire n_3408;
wire n_4167;
wire n_1904;
wire n_2640;
wire n_1993;
wire n_4823;
wire n_774;
wire n_3835;
wire n_1628;
wire n_2493;
wire n_2205;
wire n_3432;
wire n_1335;
wire n_1514;
wire n_1777;
wire n_1957;
wire n_1059;
wire n_1345;
wire n_3967;
wire n_1133;
wire n_1912;
wire n_1771;
wire n_3401;
wire n_1899;
wire n_3226;
wire n_557;
wire n_1410;
wire n_4537;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_3090;
wire n_2067;
wire n_707;
wire n_1168;
wire n_2437;
wire n_2219;
wire n_2885;
wire n_3762;
wire n_3902;
wire n_4730;
wire n_3533;
wire n_2877;
wire n_3318;
wire n_4070;
wire n_2148;
wire n_4282;
wire n_937;
wire n_2445;
wire n_1427;
wire n_2779;
wire n_3485;
wire n_4180;
wire n_1584;
wire n_665;
wire n_1726;
wire n_3035;
wire n_1835;
wire n_3839;
wire n_1440;
wire n_3654;
wire n_2164;
wire n_1988;
wire n_3333;
wire n_2115;
wire n_1853;
wire n_1356;
wire n_2845;
wire n_1787;
wire n_4137;
wire n_2634;
wire n_4529;
wire n_910;
wire n_2232;
wire n_3034;
wire n_2212;
wire n_4143;
wire n_4323;
wire n_4659;
wire n_2602;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1302;
wire n_1774;
wire n_4713;
wire n_1725;
wire n_1313;
wire n_1136;
wire n_3972;
wire n_1491;
wire n_754;
wire n_4579;
wire n_4616;
wire n_2811;
wire n_1496;
wire n_3348;
wire n_3014;
wire n_2547;
wire n_1125;
wire n_3639;
wire n_708;
wire n_1812;
wire n_735;
wire n_2501;
wire n_3079;
wire n_4105;
wire n_1915;
wire n_1109;
wire n_2532;
wire n_895;
wire n_1310;
wire n_2605;
wire n_3358;
wire n_2121;
wire n_1803;
wire n_4747;
wire n_3791;
wire n_4204;
wire n_3308;
wire n_2665;
wire n_1991;
wire n_2224;
wire n_1543;
wire n_1979;
wire n_791;
wire n_732;
wire n_1533;
wire n_3368;
wire n_1399;
wire n_2924;
wire n_4772;
wire n_3467;
wire n_808;
wire n_2484;
wire n_4111;
wire n_797;
wire n_3530;
wire n_1025;
wire n_1930;
wire n_1955;
wire n_4587;
wire n_3731;
wire n_2765;
wire n_3329;
wire n_4322;
wire n_4743;
wire n_2994;
wire n_1067;
wire n_3805;
wire n_3825;
wire n_2946;
wire n_1720;
wire n_2830;
wire n_4538;
wire n_2401;
wire n_3135;
wire n_4354;
wire n_3657;
wire n_2003;
wire n_1457;
wire n_766;
wire n_3928;
wire n_4653;
wire n_2692;
wire n_3573;
wire n_3148;
wire n_2354;
wire n_2246;
wire n_2008;
wire n_1117;
wire n_4654;
wire n_799;
wire n_2264;
wire n_4677;
wire n_2754;
wire n_687;
wire n_3534;
wire n_715;
wire n_3901;
wire n_1742;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_2489;
wire n_4275;
wire n_1266;
wire n_3970;
wire n_3757;
wire n_3438;
wire n_4098;
wire n_872;
wire n_2012;
wire n_594;
wire n_3792;
wire n_4733;
wire n_4272;
wire n_1291;
wire n_3974;
wire n_3381;
wire n_3871;
wire n_4094;
wire n_3503;
wire n_1297;
wire n_1753;
wire n_2283;
wire n_2866;
wire n_3278;
wire n_1782;
wire n_2245;
wire n_3561;
wire n_1155;
wire n_1418;
wire n_4789;
wire n_1972;
wire n_1689;
wire n_1524;
wire n_1485;
wire n_2806;
wire n_4269;
wire n_1011;
wire n_1184;
wire n_2184;
wire n_4695;
wire n_985;
wire n_2917;
wire n_2425;
wire n_1855;
wire n_869;
wire n_810;
wire n_2965;
wire n_3536;
wire n_3661;
wire n_3635;
wire n_4150;
wire n_3217;
wire n_3425;
wire n_827;
wire n_3404;
wire n_1703;
wire n_3312;
wire n_4055;
wire n_1352;
wire n_2926;
wire n_626;
wire n_2197;
wire n_2199;
wire n_3540;
wire n_1650;
wire n_3670;
wire n_1144;
wire n_3973;
wire n_1137;
wire n_1570;
wire n_2814;
wire n_3046;
wire n_3882;
wire n_3934;
wire n_1170;
wire n_2213;
wire n_2023;
wire n_3826;
wire n_3249;
wire n_3211;
wire n_3285;
wire n_2351;
wire n_2211;
wire n_2095;
wire n_3121;
wire n_3922;
wire n_3846;
wire n_676;
wire n_2103;
wire n_653;
wire n_4442;
wire n_3968;
wire n_4698;
wire n_4634;
wire n_2160;
wire n_642;
wire n_3337;
wire n_2228;
wire n_2527;
wire n_4704;
wire n_1602;
wire n_2498;
wire n_855;
wire n_1178;
wire n_1461;
wire n_2697;
wire n_4551;
wire n_850;
wire n_684;
wire n_3074;
wire n_3204;
wire n_4779;
wire n_2421;
wire n_2286;
wire n_2902;
wire n_664;
wire n_1999;
wire n_2372;
wire n_2065;
wire n_2136;
wire n_3673;
wire n_2480;
wire n_4017;
wire n_3768;
wire n_1372;
wire n_2861;
wire n_605;
wire n_2630;
wire n_1273;
wire n_3943;
wire n_1822;
wire n_3397;
wire n_3740;
wire n_620;
wire n_643;
wire n_2430;
wire n_2363;
wire n_4072;
wire n_916;
wire n_1081;
wire n_4418;
wire n_2549;
wire n_2705;
wire n_3005;
wire n_2332;
wire n_1235;
wire n_4380;
wire n_703;
wire n_698;
wire n_1115;
wire n_980;
wire n_2433;
wire n_3293;
wire n_3129;
wire n_4126;
wire n_1282;
wire n_1318;
wire n_1783;
wire n_780;
wire n_4781;
wire n_2977;
wire n_3606;
wire n_2601;
wire n_3043;
wire n_4022;
wire n_998;
wire n_3802;
wire n_2375;
wire n_4506;
wire n_2550;
wire n_1454;
wire n_3723;
wire n_1227;
wire n_1531;
wire n_840;
wire n_4424;
wire n_1334;
wire n_4852;
wire n_1907;
wire n_3600;
wire n_823;
wire n_2686;
wire n_2528;
wire n_4134;
wire n_725;
wire n_2344;
wire n_3892;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_4700;
wire n_2836;
wire n_4035;
wire n_2316;
wire n_672;
wire n_1985;
wire n_3055;
wire n_1898;
wire n_2107;
wire n_3294;
wire n_3219;
wire n_3711;
wire n_4426;
wire n_3315;
wire n_581;
wire n_2906;
wire n_554;
wire n_1625;
wire n_2130;
wire n_3415;
wire n_2284;
wire n_2187;
wire n_898;
wire n_2817;
wire n_3172;
wire n_3139;
wire n_2773;
wire n_3292;
wire n_3239;
wire n_2598;
wire n_4436;
wire n_3878;
wire n_1762;
wire n_1013;
wire n_4450;
wire n_3365;
wire n_3476;
wire n_3686;
wire n_1452;
wire n_718;
wire n_4601;
wire n_2687;
wire n_3023;
wire n_3553;
wire n_1120;
wire n_719;
wire n_4746;
wire n_1791;
wire n_1890;
wire n_1747;
wire n_714;
wire n_2850;
wire n_4220;
wire n_4251;
wire n_1817;
wire n_1944;
wire n_909;
wire n_1683;
wire n_1530;
wire n_1497;
wire n_4075;
wire n_4193;
wire n_3982;
wire n_2654;
wire n_997;
wire n_3431;
wire n_4621;
wire n_3104;
wire n_932;
wire n_3169;
wire n_3151;
wire n_612;
wire n_3822;
wire n_3131;
wire n_2078;
wire n_1409;
wire n_3850;
wire n_4737;
wire n_788;
wire n_1326;
wire n_3070;
wire n_3284;
wire n_4066;
wire n_3647;
wire n_4459;
wire n_3176;
wire n_2884;
wire n_1268;
wire n_2996;
wire n_559;
wire n_825;
wire n_4515;
wire n_4351;
wire n_2819;
wire n_3126;
wire n_4559;
wire n_4403;
wire n_1981;
wire n_2186;
wire n_1320;
wire n_4368;
wire n_1663;
wire n_737;
wire n_1718;
wire n_4050;
wire n_3700;
wire n_4509;
wire n_4740;
wire n_3609;
wire n_4136;
wire n_986;
wire n_2315;
wire n_3228;
wire n_1317;
wire n_1518;
wire n_1715;
wire n_2102;
wire n_3581;
wire n_2562;
wire n_1281;
wire n_1952;
wire n_4077;
wire n_4223;
wire n_4642;
wire n_4393;
wire n_1192;
wire n_2221;
wire n_1024;
wire n_3576;
wire n_1063;
wire n_3720;
wire n_1889;
wire n_1792;
wire n_1564;
wire n_4535;
wire n_1868;
wire n_1613;
wire n_733;
wire n_1489;
wire n_1922;
wire n_2966;
wire n_4049;
wire n_1376;
wire n_941;
wire n_2560;
wire n_981;
wire n_2326;
wire n_3862;
wire n_1569;
wire n_4522;
wire n_2188;
wire n_4794;
wire n_3495;
wire n_3879;
wire n_867;
wire n_2348;
wire n_2422;
wire n_3959;
wire n_2239;
wire n_587;
wire n_2950;
wire n_792;
wire n_756;
wire n_1429;
wire n_4724;
wire n_4644;
wire n_4456;
wire n_1238;
wire n_2448;
wire n_3140;
wire n_4346;
wire n_3852;
wire n_548;
wire n_3170;
wire n_3724;
wire n_812;
wire n_2104;
wire n_4520;
wire n_2748;
wire n_3311;
wire n_2057;
wire n_3272;
wire n_4008;
wire n_3011;
wire n_1772;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_2898;
wire n_782;
wire n_2717;
wire n_4196;
wire n_2818;
wire n_1100;
wire n_3646;
wire n_2129;
wire n_3345;
wire n_1395;
wire n_1861;
wire n_4546;
wire n_862;
wire n_3584;
wire n_1425;
wire n_4592;
wire n_760;
wire n_3858;
wire n_4675;
wire n_1901;
wire n_3069;
wire n_4502;
wire n_3756;
wire n_4370;
wire n_1900;
wire n_1620;
wire n_3032;
wire n_3628;
wire n_3691;
wire n_2889;
wire n_4851;
wire n_4235;
wire n_1330;
wire n_1867;
wire n_1945;
wire n_2772;
wire n_3018;
wire n_1675;
wire n_3072;
wire n_1924;
wire n_2573;
wire n_3084;
wire n_3081;
wire n_3313;
wire n_1727;
wire n_2710;
wire n_1554;
wire n_4382;
wire n_4435;
wire n_2939;
wire n_1745;
wire n_3924;
wire n_2735;
wire n_769;
wire n_2497;
wire n_2006;
wire n_3412;
wire n_3999;
wire n_4571;
wire n_2844;
wire n_1995;
wire n_2411;
wire n_3807;
wire n_2138;
wire n_1046;
wire n_934;
wire n_1618;
wire n_2260;
wire n_826;
wire n_2343;
wire n_1813;
wire n_2447;
wire n_3761;
wire n_4764;
wire n_886;
wire n_4833;
wire n_3439;
wire n_2014;
wire n_3056;
wire n_1221;
wire n_2345;
wire n_2986;
wire n_654;
wire n_1172;
wire n_2535;
wire n_4205;
wire n_1341;
wire n_2774;
wire n_570;
wire n_2726;
wire n_3295;
wire n_1641;
wire n_1361;
wire n_3184;
wire n_4723;
wire n_2382;
wire n_4719;
wire n_1707;
wire n_4828;
wire n_853;
wire n_4178;
wire n_4655;
wire n_3062;
wire n_3161;
wire n_4581;
wire n_2317;
wire n_751;
wire n_3289;
wire n_4558;
wire n_4827;
wire n_2799;
wire n_4454;
wire n_2172;
wire n_1973;
wire n_4229;
wire n_786;
wire n_1083;
wire n_1142;
wire n_4739;
wire n_2376;
wire n_2488;
wire n_4722;
wire n_1129;
wire n_2579;
wire n_3477;
wire n_3017;
wire n_3626;
wire n_2476;
wire n_704;
wire n_4768;
wire n_787;
wire n_4399;
wire n_1770;
wire n_2781;
wire n_4100;
wire n_4228;
wire n_2456;
wire n_4401;
wire n_3904;
wire n_961;
wire n_2250;
wire n_2678;
wire n_1756;
wire n_771;
wire n_2778;
wire n_4782;
wire n_1716;
wire n_2788;
wire n_4838;
wire n_2872;
wire n_1225;
wire n_2984;
wire n_1520;
wire n_2451;
wire n_2887;
wire n_3364;
wire n_1287;
wire n_4363;
wire n_1262;
wire n_2691;
wire n_930;
wire n_4092;
wire n_3908;
wire n_1873;
wire n_1411;
wire n_3926;
wire n_3201;
wire n_3054;
wire n_4335;
wire n_1962;
wire n_622;
wire n_3996;
wire n_4221;
wire n_1577;
wire n_2423;
wire n_3671;
wire n_1087;
wire n_3472;
wire n_2526;
wire n_2854;
wire n_994;
wire n_1701;
wire n_3344;
wire n_2194;
wire n_4181;
wire n_848;
wire n_1550;
wire n_4465;
wire n_2874;
wire n_2764;
wire n_2703;
wire n_1498;
wire n_2167;
wire n_4605;
wire n_3302;
wire n_3235;
wire n_1223;
wire n_1272;
wire n_2680;
wire n_4225;
wire n_3391;
wire n_682;
wire n_1567;
wire n_4259;
wire n_2567;
wire n_3949;
wire n_3543;
wire n_1247;
wire n_2709;
wire n_3102;
wire n_922;
wire n_3122;
wire n_816;
wire n_4808;
wire n_1648;
wire n_591;
wire n_3842;
wire n_1536;
wire n_3050;
wire n_3265;
wire n_1857;
wire n_4056;
wire n_4482;
wire n_4153;
wire n_1344;
wire n_2041;
wire n_631;
wire n_3627;
wire n_4564;
wire n_1246;
wire n_3840;
wire n_4300;
wire n_1478;
wire n_1339;
wire n_1797;
wire n_2957;
wire n_1769;
wire n_3551;
wire n_839;
wire n_3903;
wire n_4783;
wire n_4834;
wire n_1210;
wire n_3518;
wire n_2964;
wire n_3769;
wire n_1364;
wire n_2956;
wire n_2357;
wire n_3733;
wire n_2183;
wire n_2673;
wire n_2742;
wire n_3314;
wire n_4158;
wire n_4530;
wire n_2360;
wire n_3254;
wire n_4267;
wire n_2292;
wire n_1250;
wire n_2173;
wire n_3859;
wire n_3722;
wire n_3865;
wire n_4171;
wire n_1842;
wire n_871;
wire n_2442;
wire n_3309;
wire n_3738;
wire n_4045;
wire n_685;
wire n_598;
wire n_608;
wire n_928;
wire n_1367;
wire n_4562;
wire n_1943;
wire n_3634;
wire n_1460;
wire n_772;
wire n_2018;
wire n_3464;
wire n_3260;
wire n_4526;
wire n_1555;
wire n_3117;
wire n_2834;
wire n_3245;
wire n_4417;
wire n_3357;
wire n_2531;
wire n_1589;
wire n_4116;
wire n_3428;
wire n_2961;
wire n_1086;
wire n_2570;
wire n_2702;
wire n_796;
wire n_1858;
wire n_3351;
wire n_1619;
wire n_3527;
wire n_2815;
wire n_2119;
wire n_1502;
wire n_2552;
wire n_2157;
wire n_3754;
wire n_4612;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_2744;
wire n_1348;
wire n_2030;
wire n_2453;
wire n_2883;
wire n_1752;
wire n_1525;
wire n_2397;
wire n_740;
wire n_3115;
wire n_903;
wire n_4287;
wire n_4749;
wire n_3509;
wire n_3352;
wire n_4390;
wire n_2208;
wire n_3076;
wire n_1404;
wire n_4182;
wire n_3063;
wire n_3617;
wire n_2912;
wire n_1794;
wire n_3535;
wire n_2182;
wire n_1315;
wire n_2234;
wire n_4825;
wire n_1061;
wire n_3251;
wire n_4440;
wire n_4549;
wire n_4804;
wire n_1910;
wire n_1298;
wire n_3955;
wire n_2931;
wire n_1652;
wire n_4516;
wire n_2209;
wire n_3794;
wire n_2050;
wire n_2809;
wire n_4270;
wire n_4505;
wire n_1193;
wire n_2797;
wire n_1676;
wire n_1255;
wire n_1113;
wire n_3118;
wire n_4565;
wire n_4039;
wire n_3227;
wire n_3300;
wire n_4303;
wire n_2321;
wire n_3511;
wire n_1226;
wire n_4574;
wire n_722;
wire n_1277;
wire n_3680;
wire n_2591;
wire n_3443;
wire n_2146;
wire n_844;
wire n_3384;
wire n_852;
wire n_4839;
wire n_3497;
wire n_4602;
wire n_1487;
wire n_4449;
wire n_1864;
wire n_3644;
wire n_1028;
wire n_1601;
wire n_4016;
wire n_3336;
wire n_3935;
wire n_781;
wire n_2940;
wire n_3435;
wire n_3521;
wire n_3575;
wire n_1546;
wire n_595;
wire n_3562;
wire n_3948;
wire n_2612;
wire n_4750;
wire n_1337;
wire n_1495;
wire n_4445;
wire n_632;
wire n_699;
wire n_4566;
wire n_4231;
wire n_979;
wire n_1515;
wire n_2841;
wire n_3165;
wire n_1627;
wire n_2918;
wire n_3232;
wire n_3322;
wire n_4576;
wire n_3652;
wire n_1245;
wire n_846;
wire n_2427;
wire n_2438;
wire n_2505;
wire n_1673;
wire n_2832;
wire n_1321;
wire n_1975;
wire n_4097;
wire n_2296;
wire n_2070;
wire n_3250;
wire n_1937;
wire n_585;
wire n_2112;
wire n_4083;
wire n_1739;
wire n_3181;
wire n_2958;
wire n_616;
wire n_2278;
wire n_2594;
wire n_3114;
wire n_3125;
wire n_2394;
wire n_3234;
wire n_1914;
wire n_3612;
wire n_4461;
wire n_2954;
wire n_2135;
wire n_2335;
wire n_2904;
wire n_3493;
wire n_4835;
wire n_4430;
wire n_745;
wire n_2381;
wire n_4767;
wire n_3303;
wire n_1654;
wire n_4328;
wire n_3004;
wire n_3323;
wire n_3916;
wire n_2569;
wire n_3112;
wire n_2349;
wire n_1103;
wire n_3921;
wire n_4081;
wire n_3132;
wire n_3556;
wire n_648;
wire n_1379;
wire n_2734;
wire n_3874;
wire n_4101;
wire n_4407;
wire n_2196;
wire n_3591;
wire n_4676;
wire n_4273;
wire n_3951;
wire n_3024;
wire n_4544;
wire n_2170;
wire n_1076;
wire n_2823;
wire n_1091;
wire n_1408;
wire n_3512;
wire n_1761;
wire n_641;
wire n_3238;
wire n_3210;
wire n_4389;
wire n_3930;
wire n_730;
wire n_4448;
wire n_3175;
wire n_3522;
wire n_2036;
wire n_1325;
wire n_3267;
wire n_1595;
wire n_2161;
wire n_4429;
wire n_575;
wire n_795;
wire n_2404;
wire n_4345;
wire n_2083;
wire n_695;
wire n_4591;
wire n_3281;
wire n_656;
wire n_3307;
wire n_1606;
wire n_2503;
wire n_1220;
wire n_1694;
wire n_1540;
wire n_3964;
wire n_3266;
wire n_2485;
wire n_4318;
wire n_3772;
wire n_1956;
wire n_1936;
wire n_4646;
wire n_1642;
wire n_2279;
wire n_3373;
wire n_2655;
wire n_2027;
wire n_3884;
wire n_4446;
wire n_4185;
wire n_2642;
wire n_1130;
wire n_720;
wire n_2500;
wire n_4797;
wire n_2366;
wire n_4563;
wire n_4725;
wire n_1918;
wire n_1526;
wire n_863;
wire n_3726;
wire n_2210;
wire n_4169;
wire n_805;
wire n_3247;
wire n_3997;
wire n_1604;
wire n_1275;
wire n_2525;
wire n_2513;
wire n_3091;
wire n_4831;
wire n_2695;
wire n_1764;
wire n_3480;
wire n_2892;
wire n_4032;
wire n_3057;
wire n_3194;
wire n_3582;
wire n_3066;
wire n_712;
wire n_2414;
wire n_2907;
wire n_1583;
wire n_2426;
wire n_2826;
wire n_3577;
wire n_3539;
wire n_1042;
wire n_1402;
wire n_2820;
wire n_3662;
wire n_2049;
wire n_2273;
wire n_2719;
wire n_4319;
wire n_4343;
wire n_1493;
wire n_4212;
wire n_657;
wire n_4320;
wire n_644;
wire n_1741;
wire n_2229;
wire n_4124;
wire n_1160;
wire n_1397;
wire n_4057;
wire n_4332;
wire n_1258;
wire n_4314;
wire n_4596;
wire n_1074;
wire n_3347;
wire n_2004;
wire n_3216;
wire n_4492;
wire n_1621;
wire n_2708;
wire n_3809;
wire n_2113;
wire n_566;
wire n_565;
wire n_2586;
wire n_3694;
wire n_1448;
wire n_4288;
wire n_4245;
wire n_4364;
wire n_2225;
wire n_3613;
wire n_3567;
wire n_1507;
wire n_4378;
wire n_4726;
wire n_1398;
wire n_2383;
wire n_1996;
wire n_597;
wire n_1879;
wire n_3406;
wire n_3604;
wire n_3444;
wire n_3853;
wire n_4751;
wire n_1181;
wire n_1505;
wire n_4222;
wire n_4216;
wire n_1634;
wire n_3939;
wire n_1196;
wire n_4012;
wire n_2019;
wire n_651;
wire n_4636;
wire n_1340;
wire n_2274;
wire n_2972;
wire n_811;
wire n_1558;
wire n_3225;
wire n_4584;
wire n_4241;
wire n_807;
wire n_3321;
wire n_2166;
wire n_3910;
wire n_4711;
wire n_2938;
wire n_3212;
wire n_835;
wire n_666;
wire n_3319;
wire n_3594;
wire n_1433;
wire n_4309;
wire n_1704;
wire n_2256;
wire n_3152;
wire n_3721;
wire n_3335;
wire n_1254;
wire n_3799;
wire n_4119;
wire n_4298;
wire n_1026;
wire n_3413;
wire n_2026;
wire n_1969;
wire n_1234;
wire n_4680;
wire n_2109;
wire n_2044;
wire n_927;
wire n_1089;
wire n_2689;
wire n_1138;
wire n_1990;
wire n_2920;
wire n_2013;
wire n_3259;
wire n_4265;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_2614;
wire n_4191;
wire n_2511;
wire n_4293;
wire n_1681;
wire n_2991;
wire n_2010;
wire n_3688;
wire n_3383;
wire n_1018;
wire n_2242;
wire n_2752;
wire n_2247;
wire n_2894;
wire n_3016;
wire n_1693;
wire n_3585;
wire n_2975;
wire n_3473;
wire n_4188;
wire n_4560;
wire n_2599;
wire n_713;
wire n_2704;
wire n_904;
wire n_2839;
wire n_3338;
wire n_1588;
wire n_4214;
wire n_1622;
wire n_2237;
wire n_3414;
wire n_3463;
wire n_3699;
wire n_1180;
wire n_1827;
wire n_4671;
wire n_3360;
wire n_4209;
wire n_2524;
wire n_3873;
wire n_1271;
wire n_3705;
wire n_2802;
wire n_1542;
wire n_1251;
wire n_3693;
wire n_4366;
wire n_4009;
wire n_3159;
wire n_4705;
wire n_2728;
wire n_3857;
wire n_2268;
wire n_3778;
wire n_4580;

CKINVDCx5p33_ASAP7_75t_R g544 ( 
.A(n_428),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_494),
.Y(n_545)
);

INVx1_ASAP7_75t_SL g546 ( 
.A(n_27),
.Y(n_546)
);

INVx1_ASAP7_75t_SL g547 ( 
.A(n_541),
.Y(n_547)
);

CKINVDCx20_ASAP7_75t_R g548 ( 
.A(n_394),
.Y(n_548)
);

CKINVDCx5p33_ASAP7_75t_R g549 ( 
.A(n_465),
.Y(n_549)
);

CKINVDCx5p33_ASAP7_75t_R g550 ( 
.A(n_456),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_27),
.Y(n_551)
);

CKINVDCx5p33_ASAP7_75t_R g552 ( 
.A(n_281),
.Y(n_552)
);

CKINVDCx5p33_ASAP7_75t_R g553 ( 
.A(n_534),
.Y(n_553)
);

CKINVDCx5p33_ASAP7_75t_R g554 ( 
.A(n_188),
.Y(n_554)
);

CKINVDCx5p33_ASAP7_75t_R g555 ( 
.A(n_220),
.Y(n_555)
);

CKINVDCx5p33_ASAP7_75t_R g556 ( 
.A(n_156),
.Y(n_556)
);

CKINVDCx5p33_ASAP7_75t_R g557 ( 
.A(n_19),
.Y(n_557)
);

CKINVDCx5p33_ASAP7_75t_R g558 ( 
.A(n_182),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_480),
.Y(n_559)
);

CKINVDCx5p33_ASAP7_75t_R g560 ( 
.A(n_171),
.Y(n_560)
);

CKINVDCx5p33_ASAP7_75t_R g561 ( 
.A(n_491),
.Y(n_561)
);

INVx1_ASAP7_75t_SL g562 ( 
.A(n_125),
.Y(n_562)
);

INVx1_ASAP7_75t_SL g563 ( 
.A(n_238),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_148),
.Y(n_564)
);

CKINVDCx5p33_ASAP7_75t_R g565 ( 
.A(n_207),
.Y(n_565)
);

CKINVDCx5p33_ASAP7_75t_R g566 ( 
.A(n_460),
.Y(n_566)
);

CKINVDCx5p33_ASAP7_75t_R g567 ( 
.A(n_131),
.Y(n_567)
);

CKINVDCx5p33_ASAP7_75t_R g568 ( 
.A(n_341),
.Y(n_568)
);

CKINVDCx5p33_ASAP7_75t_R g569 ( 
.A(n_451),
.Y(n_569)
);

CKINVDCx5p33_ASAP7_75t_R g570 ( 
.A(n_365),
.Y(n_570)
);

INVx1_ASAP7_75t_SL g571 ( 
.A(n_426),
.Y(n_571)
);

CKINVDCx5p33_ASAP7_75t_R g572 ( 
.A(n_128),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_161),
.Y(n_573)
);

CKINVDCx5p33_ASAP7_75t_R g574 ( 
.A(n_157),
.Y(n_574)
);

CKINVDCx5p33_ASAP7_75t_R g575 ( 
.A(n_11),
.Y(n_575)
);

INVx1_ASAP7_75t_SL g576 ( 
.A(n_174),
.Y(n_576)
);

BUFx10_ASAP7_75t_L g577 ( 
.A(n_218),
.Y(n_577)
);

CKINVDCx5p33_ASAP7_75t_R g578 ( 
.A(n_404),
.Y(n_578)
);

CKINVDCx5p33_ASAP7_75t_R g579 ( 
.A(n_405),
.Y(n_579)
);

CKINVDCx5p33_ASAP7_75t_R g580 ( 
.A(n_44),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_248),
.Y(n_581)
);

INVx1_ASAP7_75t_SL g582 ( 
.A(n_163),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_253),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_264),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_129),
.Y(n_585)
);

BUFx10_ASAP7_75t_L g586 ( 
.A(n_48),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_268),
.Y(n_587)
);

CKINVDCx16_ASAP7_75t_R g588 ( 
.A(n_431),
.Y(n_588)
);

CKINVDCx5p33_ASAP7_75t_R g589 ( 
.A(n_293),
.Y(n_589)
);

CKINVDCx5p33_ASAP7_75t_R g590 ( 
.A(n_268),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_510),
.Y(n_591)
);

CKINVDCx5p33_ASAP7_75t_R g592 ( 
.A(n_533),
.Y(n_592)
);

CKINVDCx5p33_ASAP7_75t_R g593 ( 
.A(n_386),
.Y(n_593)
);

CKINVDCx5p33_ASAP7_75t_R g594 ( 
.A(n_159),
.Y(n_594)
);

CKINVDCx5p33_ASAP7_75t_R g595 ( 
.A(n_43),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_528),
.Y(n_596)
);

BUFx3_ASAP7_75t_L g597 ( 
.A(n_40),
.Y(n_597)
);

CKINVDCx5p33_ASAP7_75t_R g598 ( 
.A(n_419),
.Y(n_598)
);

HB1xp67_ASAP7_75t_L g599 ( 
.A(n_542),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_532),
.Y(n_600)
);

CKINVDCx20_ASAP7_75t_R g601 ( 
.A(n_127),
.Y(n_601)
);

CKINVDCx5p33_ASAP7_75t_R g602 ( 
.A(n_366),
.Y(n_602)
);

BUFx10_ASAP7_75t_L g603 ( 
.A(n_501),
.Y(n_603)
);

CKINVDCx5p33_ASAP7_75t_R g604 ( 
.A(n_370),
.Y(n_604)
);

INVx2_ASAP7_75t_L g605 ( 
.A(n_539),
.Y(n_605)
);

CKINVDCx5p33_ASAP7_75t_R g606 ( 
.A(n_83),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_209),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_254),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_515),
.Y(n_609)
);

CKINVDCx5p33_ASAP7_75t_R g610 ( 
.A(n_279),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_416),
.Y(n_611)
);

CKINVDCx5p33_ASAP7_75t_R g612 ( 
.A(n_105),
.Y(n_612)
);

CKINVDCx5p33_ASAP7_75t_R g613 ( 
.A(n_202),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_207),
.Y(n_614)
);

CKINVDCx20_ASAP7_75t_R g615 ( 
.A(n_201),
.Y(n_615)
);

CKINVDCx5p33_ASAP7_75t_R g616 ( 
.A(n_369),
.Y(n_616)
);

BUFx10_ASAP7_75t_L g617 ( 
.A(n_162),
.Y(n_617)
);

CKINVDCx5p33_ASAP7_75t_R g618 ( 
.A(n_306),
.Y(n_618)
);

INVx1_ASAP7_75t_SL g619 ( 
.A(n_427),
.Y(n_619)
);

CKINVDCx5p33_ASAP7_75t_R g620 ( 
.A(n_7),
.Y(n_620)
);

INVxp67_ASAP7_75t_L g621 ( 
.A(n_232),
.Y(n_621)
);

CKINVDCx5p33_ASAP7_75t_R g622 ( 
.A(n_99),
.Y(n_622)
);

INVx2_ASAP7_75t_L g623 ( 
.A(n_134),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_520),
.Y(n_624)
);

CKINVDCx5p33_ASAP7_75t_R g625 ( 
.A(n_121),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_35),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_192),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_203),
.Y(n_628)
);

CKINVDCx5p33_ASAP7_75t_R g629 ( 
.A(n_163),
.Y(n_629)
);

INVx1_ASAP7_75t_SL g630 ( 
.A(n_519),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_198),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_339),
.Y(n_632)
);

CKINVDCx20_ASAP7_75t_R g633 ( 
.A(n_508),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_512),
.Y(n_634)
);

INVx2_ASAP7_75t_L g635 ( 
.A(n_31),
.Y(n_635)
);

CKINVDCx5p33_ASAP7_75t_R g636 ( 
.A(n_483),
.Y(n_636)
);

CKINVDCx5p33_ASAP7_75t_R g637 ( 
.A(n_83),
.Y(n_637)
);

BUFx10_ASAP7_75t_L g638 ( 
.A(n_52),
.Y(n_638)
);

CKINVDCx5p33_ASAP7_75t_R g639 ( 
.A(n_44),
.Y(n_639)
);

CKINVDCx5p33_ASAP7_75t_R g640 ( 
.A(n_202),
.Y(n_640)
);

CKINVDCx5p33_ASAP7_75t_R g641 ( 
.A(n_161),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_523),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_505),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_462),
.Y(n_644)
);

INVx2_ASAP7_75t_SL g645 ( 
.A(n_197),
.Y(n_645)
);

INVx2_ASAP7_75t_L g646 ( 
.A(n_39),
.Y(n_646)
);

CKINVDCx5p33_ASAP7_75t_R g647 ( 
.A(n_478),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_120),
.Y(n_648)
);

CKINVDCx5p33_ASAP7_75t_R g649 ( 
.A(n_204),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_525),
.Y(n_650)
);

CKINVDCx5p33_ASAP7_75t_R g651 ( 
.A(n_538),
.Y(n_651)
);

CKINVDCx5p33_ASAP7_75t_R g652 ( 
.A(n_364),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_315),
.Y(n_653)
);

CKINVDCx5p33_ASAP7_75t_R g654 ( 
.A(n_401),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_67),
.Y(n_655)
);

CKINVDCx5p33_ASAP7_75t_R g656 ( 
.A(n_232),
.Y(n_656)
);

CKINVDCx5p33_ASAP7_75t_R g657 ( 
.A(n_412),
.Y(n_657)
);

CKINVDCx5p33_ASAP7_75t_R g658 ( 
.A(n_352),
.Y(n_658)
);

CKINVDCx5p33_ASAP7_75t_R g659 ( 
.A(n_271),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_226),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_516),
.Y(n_661)
);

CKINVDCx5p33_ASAP7_75t_R g662 ( 
.A(n_360),
.Y(n_662)
);

CKINVDCx5p33_ASAP7_75t_R g663 ( 
.A(n_77),
.Y(n_663)
);

CKINVDCx5p33_ASAP7_75t_R g664 ( 
.A(n_10),
.Y(n_664)
);

CKINVDCx5p33_ASAP7_75t_R g665 ( 
.A(n_7),
.Y(n_665)
);

BUFx10_ASAP7_75t_L g666 ( 
.A(n_103),
.Y(n_666)
);

CKINVDCx5p33_ASAP7_75t_R g667 ( 
.A(n_484),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_182),
.Y(n_668)
);

INVx2_ASAP7_75t_SL g669 ( 
.A(n_361),
.Y(n_669)
);

CKINVDCx5p33_ASAP7_75t_R g670 ( 
.A(n_351),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_299),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_130),
.Y(n_672)
);

BUFx6f_ASAP7_75t_L g673 ( 
.A(n_165),
.Y(n_673)
);

BUFx10_ASAP7_75t_L g674 ( 
.A(n_180),
.Y(n_674)
);

CKINVDCx5p33_ASAP7_75t_R g675 ( 
.A(n_241),
.Y(n_675)
);

CKINVDCx5p33_ASAP7_75t_R g676 ( 
.A(n_108),
.Y(n_676)
);

BUFx3_ASAP7_75t_L g677 ( 
.A(n_23),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_487),
.Y(n_678)
);

BUFx6f_ASAP7_75t_L g679 ( 
.A(n_387),
.Y(n_679)
);

CKINVDCx16_ASAP7_75t_R g680 ( 
.A(n_113),
.Y(n_680)
);

CKINVDCx5p33_ASAP7_75t_R g681 ( 
.A(n_255),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_128),
.Y(n_682)
);

CKINVDCx5p33_ASAP7_75t_R g683 ( 
.A(n_212),
.Y(n_683)
);

INVx2_ASAP7_75t_L g684 ( 
.A(n_434),
.Y(n_684)
);

CKINVDCx5p33_ASAP7_75t_R g685 ( 
.A(n_194),
.Y(n_685)
);

CKINVDCx5p33_ASAP7_75t_R g686 ( 
.A(n_527),
.Y(n_686)
);

CKINVDCx20_ASAP7_75t_R g687 ( 
.A(n_286),
.Y(n_687)
);

CKINVDCx5p33_ASAP7_75t_R g688 ( 
.A(n_62),
.Y(n_688)
);

HB1xp67_ASAP7_75t_L g689 ( 
.A(n_279),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_454),
.Y(n_690)
);

CKINVDCx5p33_ASAP7_75t_R g691 ( 
.A(n_249),
.Y(n_691)
);

INVx1_ASAP7_75t_SL g692 ( 
.A(n_444),
.Y(n_692)
);

CKINVDCx5p33_ASAP7_75t_R g693 ( 
.A(n_518),
.Y(n_693)
);

INVx2_ASAP7_75t_L g694 ( 
.A(n_406),
.Y(n_694)
);

CKINVDCx5p33_ASAP7_75t_R g695 ( 
.A(n_93),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_183),
.Y(n_696)
);

CKINVDCx5p33_ASAP7_75t_R g697 ( 
.A(n_275),
.Y(n_697)
);

INVx2_ASAP7_75t_SL g698 ( 
.A(n_191),
.Y(n_698)
);

CKINVDCx20_ASAP7_75t_R g699 ( 
.A(n_55),
.Y(n_699)
);

CKINVDCx5p33_ASAP7_75t_R g700 ( 
.A(n_496),
.Y(n_700)
);

CKINVDCx5p33_ASAP7_75t_R g701 ( 
.A(n_537),
.Y(n_701)
);

INVx2_ASAP7_75t_L g702 ( 
.A(n_152),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_0),
.Y(n_703)
);

CKINVDCx5p33_ASAP7_75t_R g704 ( 
.A(n_258),
.Y(n_704)
);

CKINVDCx5p33_ASAP7_75t_R g705 ( 
.A(n_213),
.Y(n_705)
);

CKINVDCx20_ASAP7_75t_R g706 ( 
.A(n_345),
.Y(n_706)
);

INVx1_ASAP7_75t_SL g707 ( 
.A(n_334),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_540),
.Y(n_708)
);

CKINVDCx5p33_ASAP7_75t_R g709 ( 
.A(n_105),
.Y(n_709)
);

CKINVDCx20_ASAP7_75t_R g710 ( 
.A(n_73),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_259),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_77),
.Y(n_712)
);

CKINVDCx5p33_ASAP7_75t_R g713 ( 
.A(n_325),
.Y(n_713)
);

CKINVDCx5p33_ASAP7_75t_R g714 ( 
.A(n_321),
.Y(n_714)
);

CKINVDCx5p33_ASAP7_75t_R g715 ( 
.A(n_471),
.Y(n_715)
);

CKINVDCx5p33_ASAP7_75t_R g716 ( 
.A(n_291),
.Y(n_716)
);

BUFx10_ASAP7_75t_L g717 ( 
.A(n_457),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_52),
.Y(n_718)
);

CKINVDCx5p33_ASAP7_75t_R g719 ( 
.A(n_300),
.Y(n_719)
);

CKINVDCx5p33_ASAP7_75t_R g720 ( 
.A(n_5),
.Y(n_720)
);

CKINVDCx20_ASAP7_75t_R g721 ( 
.A(n_198),
.Y(n_721)
);

CKINVDCx20_ASAP7_75t_R g722 ( 
.A(n_173),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_507),
.Y(n_723)
);

BUFx6f_ASAP7_75t_L g724 ( 
.A(n_119),
.Y(n_724)
);

INVx2_ASAP7_75t_SL g725 ( 
.A(n_96),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_312),
.Y(n_726)
);

CKINVDCx5p33_ASAP7_75t_R g727 ( 
.A(n_490),
.Y(n_727)
);

INVx2_ASAP7_75t_SL g728 ( 
.A(n_322),
.Y(n_728)
);

CKINVDCx5p33_ASAP7_75t_R g729 ( 
.A(n_203),
.Y(n_729)
);

CKINVDCx5p33_ASAP7_75t_R g730 ( 
.A(n_391),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_476),
.Y(n_731)
);

BUFx10_ASAP7_75t_L g732 ( 
.A(n_216),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_340),
.Y(n_733)
);

CKINVDCx5p33_ASAP7_75t_R g734 ( 
.A(n_53),
.Y(n_734)
);

INVx2_ASAP7_75t_SL g735 ( 
.A(n_46),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_121),
.Y(n_736)
);

CKINVDCx20_ASAP7_75t_R g737 ( 
.A(n_19),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_137),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_439),
.Y(n_739)
);

CKINVDCx5p33_ASAP7_75t_R g740 ( 
.A(n_499),
.Y(n_740)
);

CKINVDCx5p33_ASAP7_75t_R g741 ( 
.A(n_376),
.Y(n_741)
);

CKINVDCx5p33_ASAP7_75t_R g742 ( 
.A(n_233),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_36),
.Y(n_743)
);

CKINVDCx14_ASAP7_75t_R g744 ( 
.A(n_38),
.Y(n_744)
);

CKINVDCx5p33_ASAP7_75t_R g745 ( 
.A(n_294),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_53),
.Y(n_746)
);

CKINVDCx5p33_ASAP7_75t_R g747 ( 
.A(n_240),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_86),
.Y(n_748)
);

INVxp67_ASAP7_75t_L g749 ( 
.A(n_17),
.Y(n_749)
);

CKINVDCx5p33_ASAP7_75t_R g750 ( 
.A(n_402),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_514),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_127),
.Y(n_752)
);

CKINVDCx5p33_ASAP7_75t_R g753 ( 
.A(n_133),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_464),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_81),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_31),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_178),
.Y(n_757)
);

CKINVDCx5p33_ASAP7_75t_R g758 ( 
.A(n_82),
.Y(n_758)
);

INVx2_ASAP7_75t_L g759 ( 
.A(n_503),
.Y(n_759)
);

INVx2_ASAP7_75t_SL g760 ( 
.A(n_168),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_373),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_216),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_208),
.Y(n_763)
);

BUFx3_ASAP7_75t_L g764 ( 
.A(n_440),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_61),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_327),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_122),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_475),
.Y(n_768)
);

CKINVDCx20_ASAP7_75t_R g769 ( 
.A(n_14),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_72),
.Y(n_770)
);

CKINVDCx5p33_ASAP7_75t_R g771 ( 
.A(n_60),
.Y(n_771)
);

CKINVDCx5p33_ASAP7_75t_R g772 ( 
.A(n_132),
.Y(n_772)
);

INVx1_ASAP7_75t_SL g773 ( 
.A(n_536),
.Y(n_773)
);

INVx1_ASAP7_75t_SL g774 ( 
.A(n_129),
.Y(n_774)
);

CKINVDCx5p33_ASAP7_75t_R g775 ( 
.A(n_495),
.Y(n_775)
);

INVx1_ASAP7_75t_SL g776 ( 
.A(n_194),
.Y(n_776)
);

CKINVDCx5p33_ASAP7_75t_R g777 ( 
.A(n_11),
.Y(n_777)
);

BUFx3_ASAP7_75t_L g778 ( 
.A(n_130),
.Y(n_778)
);

CKINVDCx20_ASAP7_75t_R g779 ( 
.A(n_463),
.Y(n_779)
);

CKINVDCx5p33_ASAP7_75t_R g780 ( 
.A(n_332),
.Y(n_780)
);

CKINVDCx5p33_ASAP7_75t_R g781 ( 
.A(n_342),
.Y(n_781)
);

CKINVDCx5p33_ASAP7_75t_R g782 ( 
.A(n_115),
.Y(n_782)
);

CKINVDCx5p33_ASAP7_75t_R g783 ( 
.A(n_253),
.Y(n_783)
);

INVx2_ASAP7_75t_SL g784 ( 
.A(n_385),
.Y(n_784)
);

CKINVDCx5p33_ASAP7_75t_R g785 ( 
.A(n_326),
.Y(n_785)
);

BUFx5_ASAP7_75t_L g786 ( 
.A(n_113),
.Y(n_786)
);

CKINVDCx5p33_ASAP7_75t_R g787 ( 
.A(n_392),
.Y(n_787)
);

CKINVDCx5p33_ASAP7_75t_R g788 ( 
.A(n_99),
.Y(n_788)
);

CKINVDCx5p33_ASAP7_75t_R g789 ( 
.A(n_145),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_230),
.Y(n_790)
);

BUFx6f_ASAP7_75t_L g791 ( 
.A(n_181),
.Y(n_791)
);

BUFx3_ASAP7_75t_L g792 ( 
.A(n_448),
.Y(n_792)
);

CKINVDCx5p33_ASAP7_75t_R g793 ( 
.A(n_269),
.Y(n_793)
);

INVx2_ASAP7_75t_L g794 ( 
.A(n_126),
.Y(n_794)
);

CKINVDCx16_ASAP7_75t_R g795 ( 
.A(n_187),
.Y(n_795)
);

BUFx5_ASAP7_75t_L g796 ( 
.A(n_335),
.Y(n_796)
);

CKINVDCx16_ASAP7_75t_R g797 ( 
.A(n_158),
.Y(n_797)
);

CKINVDCx5p33_ASAP7_75t_R g798 ( 
.A(n_436),
.Y(n_798)
);

CKINVDCx5p33_ASAP7_75t_R g799 ( 
.A(n_382),
.Y(n_799)
);

BUFx2_ASAP7_75t_L g800 ( 
.A(n_18),
.Y(n_800)
);

CKINVDCx5p33_ASAP7_75t_R g801 ( 
.A(n_98),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_139),
.Y(n_802)
);

CKINVDCx5p33_ASAP7_75t_R g803 ( 
.A(n_186),
.Y(n_803)
);

CKINVDCx5p33_ASAP7_75t_R g804 ( 
.A(n_29),
.Y(n_804)
);

CKINVDCx5p33_ASAP7_75t_R g805 ( 
.A(n_529),
.Y(n_805)
);

BUFx10_ASAP7_75t_L g806 ( 
.A(n_153),
.Y(n_806)
);

CKINVDCx5p33_ASAP7_75t_R g807 ( 
.A(n_260),
.Y(n_807)
);

CKINVDCx5p33_ASAP7_75t_R g808 ( 
.A(n_543),
.Y(n_808)
);

BUFx2_ASAP7_75t_L g809 ( 
.A(n_60),
.Y(n_809)
);

CKINVDCx5p33_ASAP7_75t_R g810 ( 
.A(n_297),
.Y(n_810)
);

INVx2_ASAP7_75t_SL g811 ( 
.A(n_437),
.Y(n_811)
);

BUFx6f_ASAP7_75t_L g812 ( 
.A(n_337),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_530),
.Y(n_813)
);

INVx2_ASAP7_75t_SL g814 ( 
.A(n_102),
.Y(n_814)
);

CKINVDCx5p33_ASAP7_75t_R g815 ( 
.A(n_144),
.Y(n_815)
);

CKINVDCx5p33_ASAP7_75t_R g816 ( 
.A(n_191),
.Y(n_816)
);

CKINVDCx5p33_ASAP7_75t_R g817 ( 
.A(n_274),
.Y(n_817)
);

CKINVDCx5p33_ASAP7_75t_R g818 ( 
.A(n_153),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_301),
.Y(n_819)
);

BUFx3_ASAP7_75t_L g820 ( 
.A(n_155),
.Y(n_820)
);

BUFx6f_ASAP7_75t_L g821 ( 
.A(n_485),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_282),
.Y(n_822)
);

CKINVDCx16_ASAP7_75t_R g823 ( 
.A(n_222),
.Y(n_823)
);

CKINVDCx5p33_ASAP7_75t_R g824 ( 
.A(n_139),
.Y(n_824)
);

CKINVDCx5p33_ASAP7_75t_R g825 ( 
.A(n_249),
.Y(n_825)
);

CKINVDCx5p33_ASAP7_75t_R g826 ( 
.A(n_3),
.Y(n_826)
);

CKINVDCx5p33_ASAP7_75t_R g827 ( 
.A(n_50),
.Y(n_827)
);

CKINVDCx5p33_ASAP7_75t_R g828 ( 
.A(n_137),
.Y(n_828)
);

INVx1_ASAP7_75t_SL g829 ( 
.A(n_40),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_281),
.Y(n_830)
);

CKINVDCx5p33_ASAP7_75t_R g831 ( 
.A(n_347),
.Y(n_831)
);

CKINVDCx5p33_ASAP7_75t_R g832 ( 
.A(n_290),
.Y(n_832)
);

CKINVDCx5p33_ASAP7_75t_R g833 ( 
.A(n_488),
.Y(n_833)
);

CKINVDCx5p33_ASAP7_75t_R g834 ( 
.A(n_173),
.Y(n_834)
);

BUFx10_ASAP7_75t_L g835 ( 
.A(n_493),
.Y(n_835)
);

CKINVDCx5p33_ASAP7_75t_R g836 ( 
.A(n_378),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_468),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_84),
.Y(n_838)
);

CKINVDCx5p33_ASAP7_75t_R g839 ( 
.A(n_438),
.Y(n_839)
);

CKINVDCx5p33_ASAP7_75t_R g840 ( 
.A(n_218),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_254),
.Y(n_841)
);

BUFx3_ASAP7_75t_L g842 ( 
.A(n_259),
.Y(n_842)
);

INVx2_ASAP7_75t_L g843 ( 
.A(n_87),
.Y(n_843)
);

CKINVDCx5p33_ASAP7_75t_R g844 ( 
.A(n_368),
.Y(n_844)
);

CKINVDCx5p33_ASAP7_75t_R g845 ( 
.A(n_243),
.Y(n_845)
);

CKINVDCx5p33_ASAP7_75t_R g846 ( 
.A(n_16),
.Y(n_846)
);

CKINVDCx5p33_ASAP7_75t_R g847 ( 
.A(n_276),
.Y(n_847)
);

CKINVDCx5p33_ASAP7_75t_R g848 ( 
.A(n_13),
.Y(n_848)
);

CKINVDCx5p33_ASAP7_75t_R g849 ( 
.A(n_297),
.Y(n_849)
);

CKINVDCx20_ASAP7_75t_R g850 ( 
.A(n_9),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_69),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_175),
.Y(n_852)
);

CKINVDCx5p33_ASAP7_75t_R g853 ( 
.A(n_291),
.Y(n_853)
);

INVx2_ASAP7_75t_L g854 ( 
.A(n_242),
.Y(n_854)
);

INVx2_ASAP7_75t_L g855 ( 
.A(n_152),
.Y(n_855)
);

CKINVDCx5p33_ASAP7_75t_R g856 ( 
.A(n_317),
.Y(n_856)
);

INVx1_ASAP7_75t_L g857 ( 
.A(n_455),
.Y(n_857)
);

CKINVDCx5p33_ASAP7_75t_R g858 ( 
.A(n_396),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_521),
.Y(n_859)
);

CKINVDCx5p33_ASAP7_75t_R g860 ( 
.A(n_269),
.Y(n_860)
);

CKINVDCx20_ASAP7_75t_R g861 ( 
.A(n_176),
.Y(n_861)
);

CKINVDCx5p33_ASAP7_75t_R g862 ( 
.A(n_450),
.Y(n_862)
);

CKINVDCx5p33_ASAP7_75t_R g863 ( 
.A(n_239),
.Y(n_863)
);

INVx2_ASAP7_75t_SL g864 ( 
.A(n_400),
.Y(n_864)
);

CKINVDCx14_ASAP7_75t_R g865 ( 
.A(n_146),
.Y(n_865)
);

BUFx2_ASAP7_75t_L g866 ( 
.A(n_230),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_28),
.Y(n_867)
);

CKINVDCx5p33_ASAP7_75t_R g868 ( 
.A(n_513),
.Y(n_868)
);

CKINVDCx5p33_ASAP7_75t_R g869 ( 
.A(n_415),
.Y(n_869)
);

BUFx8_ASAP7_75t_SL g870 ( 
.A(n_193),
.Y(n_870)
);

CKINVDCx5p33_ASAP7_75t_R g871 ( 
.A(n_466),
.Y(n_871)
);

INVx1_ASAP7_75t_SL g872 ( 
.A(n_302),
.Y(n_872)
);

CKINVDCx5p33_ASAP7_75t_R g873 ( 
.A(n_251),
.Y(n_873)
);

CKINVDCx5p33_ASAP7_75t_R g874 ( 
.A(n_90),
.Y(n_874)
);

INVx3_ASAP7_75t_L g875 ( 
.A(n_486),
.Y(n_875)
);

CKINVDCx5p33_ASAP7_75t_R g876 ( 
.A(n_328),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_41),
.Y(n_877)
);

CKINVDCx5p33_ASAP7_75t_R g878 ( 
.A(n_42),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_175),
.Y(n_879)
);

CKINVDCx20_ASAP7_75t_R g880 ( 
.A(n_48),
.Y(n_880)
);

INVx1_ASAP7_75t_L g881 ( 
.A(n_111),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_123),
.Y(n_882)
);

CKINVDCx5p33_ASAP7_75t_R g883 ( 
.A(n_263),
.Y(n_883)
);

CKINVDCx5p33_ASAP7_75t_R g884 ( 
.A(n_3),
.Y(n_884)
);

CKINVDCx5p33_ASAP7_75t_R g885 ( 
.A(n_290),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_295),
.Y(n_886)
);

CKINVDCx5p33_ASAP7_75t_R g887 ( 
.A(n_37),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_126),
.Y(n_888)
);

CKINVDCx5p33_ASAP7_75t_R g889 ( 
.A(n_204),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_489),
.Y(n_890)
);

CKINVDCx5p33_ASAP7_75t_R g891 ( 
.A(n_220),
.Y(n_891)
);

CKINVDCx5p33_ASAP7_75t_R g892 ( 
.A(n_535),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_423),
.Y(n_893)
);

INVx2_ASAP7_75t_L g894 ( 
.A(n_85),
.Y(n_894)
);

CKINVDCx5p33_ASAP7_75t_R g895 ( 
.A(n_266),
.Y(n_895)
);

CKINVDCx5p33_ASAP7_75t_R g896 ( 
.A(n_531),
.Y(n_896)
);

INVx1_ASAP7_75t_L g897 ( 
.A(n_13),
.Y(n_897)
);

CKINVDCx5p33_ASAP7_75t_R g898 ( 
.A(n_155),
.Y(n_898)
);

CKINVDCx5p33_ASAP7_75t_R g899 ( 
.A(n_319),
.Y(n_899)
);

INVx1_ASAP7_75t_L g900 ( 
.A(n_449),
.Y(n_900)
);

CKINVDCx5p33_ASAP7_75t_R g901 ( 
.A(n_33),
.Y(n_901)
);

CKINVDCx5p33_ASAP7_75t_R g902 ( 
.A(n_417),
.Y(n_902)
);

CKINVDCx5p33_ASAP7_75t_R g903 ( 
.A(n_239),
.Y(n_903)
);

BUFx3_ASAP7_75t_L g904 ( 
.A(n_223),
.Y(n_904)
);

INVx2_ASAP7_75t_L g905 ( 
.A(n_277),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_458),
.Y(n_906)
);

INVx1_ASAP7_75t_SL g907 ( 
.A(n_403),
.Y(n_907)
);

CKINVDCx5p33_ASAP7_75t_R g908 ( 
.A(n_122),
.Y(n_908)
);

CKINVDCx5p33_ASAP7_75t_R g909 ( 
.A(n_131),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_107),
.Y(n_910)
);

BUFx10_ASAP7_75t_L g911 ( 
.A(n_272),
.Y(n_911)
);

BUFx2_ASAP7_75t_L g912 ( 
.A(n_98),
.Y(n_912)
);

BUFx2_ASAP7_75t_L g913 ( 
.A(n_9),
.Y(n_913)
);

INVx1_ASAP7_75t_L g914 ( 
.A(n_304),
.Y(n_914)
);

BUFx6f_ASAP7_75t_L g915 ( 
.A(n_349),
.Y(n_915)
);

CKINVDCx5p33_ASAP7_75t_R g916 ( 
.A(n_82),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_270),
.Y(n_917)
);

INVx1_ASAP7_75t_L g918 ( 
.A(n_270),
.Y(n_918)
);

CKINVDCx5p33_ASAP7_75t_R g919 ( 
.A(n_68),
.Y(n_919)
);

INVx1_ASAP7_75t_L g920 ( 
.A(n_223),
.Y(n_920)
);

CKINVDCx5p33_ASAP7_75t_R g921 ( 
.A(n_88),
.Y(n_921)
);

INVx1_ASAP7_75t_L g922 ( 
.A(n_226),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_421),
.Y(n_923)
);

CKINVDCx5p33_ASAP7_75t_R g924 ( 
.A(n_524),
.Y(n_924)
);

INVx1_ASAP7_75t_L g925 ( 
.A(n_511),
.Y(n_925)
);

CKINVDCx5p33_ASAP7_75t_R g926 ( 
.A(n_395),
.Y(n_926)
);

CKINVDCx5p33_ASAP7_75t_R g927 ( 
.A(n_522),
.Y(n_927)
);

CKINVDCx5p33_ASAP7_75t_R g928 ( 
.A(n_414),
.Y(n_928)
);

INVx1_ASAP7_75t_L g929 ( 
.A(n_266),
.Y(n_929)
);

CKINVDCx5p33_ASAP7_75t_R g930 ( 
.A(n_358),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_265),
.Y(n_931)
);

CKINVDCx5p33_ASAP7_75t_R g932 ( 
.A(n_526),
.Y(n_932)
);

CKINVDCx5p33_ASAP7_75t_R g933 ( 
.A(n_388),
.Y(n_933)
);

CKINVDCx5p33_ASAP7_75t_R g934 ( 
.A(n_70),
.Y(n_934)
);

CKINVDCx5p33_ASAP7_75t_R g935 ( 
.A(n_318),
.Y(n_935)
);

INVx2_ASAP7_75t_L g936 ( 
.A(n_356),
.Y(n_936)
);

CKINVDCx5p33_ASAP7_75t_R g937 ( 
.A(n_236),
.Y(n_937)
);

CKINVDCx5p33_ASAP7_75t_R g938 ( 
.A(n_408),
.Y(n_938)
);

CKINVDCx5p33_ASAP7_75t_R g939 ( 
.A(n_158),
.Y(n_939)
);

CKINVDCx5p33_ASAP7_75t_R g940 ( 
.A(n_243),
.Y(n_940)
);

CKINVDCx5p33_ASAP7_75t_R g941 ( 
.A(n_459),
.Y(n_941)
);

INVx2_ASAP7_75t_SL g942 ( 
.A(n_308),
.Y(n_942)
);

CKINVDCx5p33_ASAP7_75t_R g943 ( 
.A(n_294),
.Y(n_943)
);

INVx1_ASAP7_75t_L g944 ( 
.A(n_445),
.Y(n_944)
);

BUFx8_ASAP7_75t_SL g945 ( 
.A(n_110),
.Y(n_945)
);

INVx1_ASAP7_75t_SL g946 ( 
.A(n_422),
.Y(n_946)
);

CKINVDCx5p33_ASAP7_75t_R g947 ( 
.A(n_284),
.Y(n_947)
);

CKINVDCx5p33_ASAP7_75t_R g948 ( 
.A(n_114),
.Y(n_948)
);

CKINVDCx20_ASAP7_75t_R g949 ( 
.A(n_85),
.Y(n_949)
);

CKINVDCx5p33_ASAP7_75t_R g950 ( 
.A(n_5),
.Y(n_950)
);

BUFx5_ASAP7_75t_L g951 ( 
.A(n_300),
.Y(n_951)
);

INVx1_ASAP7_75t_L g952 ( 
.A(n_94),
.Y(n_952)
);

INVx1_ASAP7_75t_L g953 ( 
.A(n_39),
.Y(n_953)
);

INVx1_ASAP7_75t_L g954 ( 
.A(n_145),
.Y(n_954)
);

CKINVDCx14_ASAP7_75t_R g955 ( 
.A(n_221),
.Y(n_955)
);

INVx1_ASAP7_75t_L g956 ( 
.A(n_179),
.Y(n_956)
);

INVx1_ASAP7_75t_SL g957 ( 
.A(n_504),
.Y(n_957)
);

INVx1_ASAP7_75t_L g958 ( 
.A(n_435),
.Y(n_958)
);

CKINVDCx5p33_ASAP7_75t_R g959 ( 
.A(n_92),
.Y(n_959)
);

INVxp33_ASAP7_75t_L g960 ( 
.A(n_689),
.Y(n_960)
);

INVx1_ASAP7_75t_L g961 ( 
.A(n_786),
.Y(n_961)
);

INVx1_ASAP7_75t_L g962 ( 
.A(n_786),
.Y(n_962)
);

INVx1_ASAP7_75t_L g963 ( 
.A(n_786),
.Y(n_963)
);

INVxp33_ASAP7_75t_SL g964 ( 
.A(n_552),
.Y(n_964)
);

CKINVDCx16_ASAP7_75t_R g965 ( 
.A(n_680),
.Y(n_965)
);

INVx1_ASAP7_75t_L g966 ( 
.A(n_786),
.Y(n_966)
);

INVx1_ASAP7_75t_L g967 ( 
.A(n_786),
.Y(n_967)
);

INVx1_ASAP7_75t_L g968 ( 
.A(n_786),
.Y(n_968)
);

INVx1_ASAP7_75t_L g969 ( 
.A(n_786),
.Y(n_969)
);

CKINVDCx5p33_ASAP7_75t_R g970 ( 
.A(n_870),
.Y(n_970)
);

INVxp67_ASAP7_75t_SL g971 ( 
.A(n_599),
.Y(n_971)
);

CKINVDCx5p33_ASAP7_75t_R g972 ( 
.A(n_945),
.Y(n_972)
);

INVx1_ASAP7_75t_L g973 ( 
.A(n_951),
.Y(n_973)
);

INVx1_ASAP7_75t_L g974 ( 
.A(n_951),
.Y(n_974)
);

NAND2xp5_ASAP7_75t_L g975 ( 
.A(n_744),
.B(n_0),
.Y(n_975)
);

INVx1_ASAP7_75t_L g976 ( 
.A(n_951),
.Y(n_976)
);

INVx1_ASAP7_75t_L g977 ( 
.A(n_951),
.Y(n_977)
);

CKINVDCx5p33_ASAP7_75t_R g978 ( 
.A(n_865),
.Y(n_978)
);

BUFx2_ASAP7_75t_L g979 ( 
.A(n_800),
.Y(n_979)
);

INVx1_ASAP7_75t_L g980 ( 
.A(n_951),
.Y(n_980)
);

INVx1_ASAP7_75t_L g981 ( 
.A(n_951),
.Y(n_981)
);

INVx1_ASAP7_75t_L g982 ( 
.A(n_951),
.Y(n_982)
);

INVx1_ASAP7_75t_L g983 ( 
.A(n_951),
.Y(n_983)
);

INVx1_ASAP7_75t_L g984 ( 
.A(n_597),
.Y(n_984)
);

CKINVDCx20_ASAP7_75t_R g985 ( 
.A(n_601),
.Y(n_985)
);

INVx1_ASAP7_75t_L g986 ( 
.A(n_597),
.Y(n_986)
);

CKINVDCx5p33_ASAP7_75t_R g987 ( 
.A(n_955),
.Y(n_987)
);

INVx1_ASAP7_75t_L g988 ( 
.A(n_677),
.Y(n_988)
);

INVx1_ASAP7_75t_L g989 ( 
.A(n_677),
.Y(n_989)
);

INVxp67_ASAP7_75t_L g990 ( 
.A(n_809),
.Y(n_990)
);

INVx1_ASAP7_75t_L g991 ( 
.A(n_778),
.Y(n_991)
);

INVxp33_ASAP7_75t_SL g992 ( 
.A(n_552),
.Y(n_992)
);

INVxp67_ASAP7_75t_L g993 ( 
.A(n_866),
.Y(n_993)
);

HB1xp67_ASAP7_75t_L g994 ( 
.A(n_795),
.Y(n_994)
);

INVx1_ASAP7_75t_L g995 ( 
.A(n_778),
.Y(n_995)
);

INVx1_ASAP7_75t_L g996 ( 
.A(n_820),
.Y(n_996)
);

BUFx3_ASAP7_75t_L g997 ( 
.A(n_764),
.Y(n_997)
);

INVx1_ASAP7_75t_L g998 ( 
.A(n_673),
.Y(n_998)
);

INVxp67_ASAP7_75t_L g999 ( 
.A(n_912),
.Y(n_999)
);

INVx2_ASAP7_75t_L g1000 ( 
.A(n_673),
.Y(n_1000)
);

INVx2_ASAP7_75t_L g1001 ( 
.A(n_673),
.Y(n_1001)
);

INVx1_ASAP7_75t_L g1002 ( 
.A(n_820),
.Y(n_1002)
);

CKINVDCx5p33_ASAP7_75t_R g1003 ( 
.A(n_797),
.Y(n_1003)
);

BUFx3_ASAP7_75t_L g1004 ( 
.A(n_764),
.Y(n_1004)
);

BUFx3_ASAP7_75t_L g1005 ( 
.A(n_792),
.Y(n_1005)
);

INVx1_ASAP7_75t_L g1006 ( 
.A(n_842),
.Y(n_1006)
);

INVx1_ASAP7_75t_L g1007 ( 
.A(n_842),
.Y(n_1007)
);

INVx1_ASAP7_75t_L g1008 ( 
.A(n_904),
.Y(n_1008)
);

INVx1_ASAP7_75t_L g1009 ( 
.A(n_904),
.Y(n_1009)
);

HB1xp67_ASAP7_75t_L g1010 ( 
.A(n_823),
.Y(n_1010)
);

INVx1_ASAP7_75t_L g1011 ( 
.A(n_673),
.Y(n_1011)
);

INVx1_ASAP7_75t_L g1012 ( 
.A(n_673),
.Y(n_1012)
);

INVx1_ASAP7_75t_L g1013 ( 
.A(n_724),
.Y(n_1013)
);

INVx1_ASAP7_75t_L g1014 ( 
.A(n_724),
.Y(n_1014)
);

INVx2_ASAP7_75t_L g1015 ( 
.A(n_724),
.Y(n_1015)
);

INVxp67_ASAP7_75t_SL g1016 ( 
.A(n_792),
.Y(n_1016)
);

CKINVDCx20_ASAP7_75t_R g1017 ( 
.A(n_615),
.Y(n_1017)
);

INVx1_ASAP7_75t_L g1018 ( 
.A(n_724),
.Y(n_1018)
);

INVx1_ASAP7_75t_L g1019 ( 
.A(n_724),
.Y(n_1019)
);

INVx1_ASAP7_75t_L g1020 ( 
.A(n_791),
.Y(n_1020)
);

INVx1_ASAP7_75t_L g1021 ( 
.A(n_791),
.Y(n_1021)
);

CKINVDCx5p33_ASAP7_75t_R g1022 ( 
.A(n_625),
.Y(n_1022)
);

INVxp67_ASAP7_75t_L g1023 ( 
.A(n_913),
.Y(n_1023)
);

INVx3_ASAP7_75t_L g1024 ( 
.A(n_791),
.Y(n_1024)
);

INVx1_ASAP7_75t_L g1025 ( 
.A(n_791),
.Y(n_1025)
);

INVx1_ASAP7_75t_L g1026 ( 
.A(n_791),
.Y(n_1026)
);

INVx1_ASAP7_75t_L g1027 ( 
.A(n_551),
.Y(n_1027)
);

CKINVDCx5p33_ASAP7_75t_R g1028 ( 
.A(n_629),
.Y(n_1028)
);

INVx1_ASAP7_75t_L g1029 ( 
.A(n_564),
.Y(n_1029)
);

INVx2_ASAP7_75t_SL g1030 ( 
.A(n_577),
.Y(n_1030)
);

INVx2_ASAP7_75t_L g1031 ( 
.A(n_796),
.Y(n_1031)
);

INVx1_ASAP7_75t_L g1032 ( 
.A(n_573),
.Y(n_1032)
);

INVx1_ASAP7_75t_L g1033 ( 
.A(n_581),
.Y(n_1033)
);

INVx1_ASAP7_75t_L g1034 ( 
.A(n_583),
.Y(n_1034)
);

INVx1_ASAP7_75t_L g1035 ( 
.A(n_584),
.Y(n_1035)
);

INVx1_ASAP7_75t_L g1036 ( 
.A(n_585),
.Y(n_1036)
);

INVx2_ASAP7_75t_SL g1037 ( 
.A(n_577),
.Y(n_1037)
);

INVx1_ASAP7_75t_L g1038 ( 
.A(n_587),
.Y(n_1038)
);

CKINVDCx16_ASAP7_75t_R g1039 ( 
.A(n_588),
.Y(n_1039)
);

INVx1_ASAP7_75t_L g1040 ( 
.A(n_607),
.Y(n_1040)
);

CKINVDCx20_ASAP7_75t_R g1041 ( 
.A(n_687),
.Y(n_1041)
);

CKINVDCx14_ASAP7_75t_R g1042 ( 
.A(n_603),
.Y(n_1042)
);

INVx1_ASAP7_75t_L g1043 ( 
.A(n_608),
.Y(n_1043)
);

INVx1_ASAP7_75t_L g1044 ( 
.A(n_614),
.Y(n_1044)
);

CKINVDCx5p33_ASAP7_75t_R g1045 ( 
.A(n_637),
.Y(n_1045)
);

CKINVDCx20_ASAP7_75t_R g1046 ( 
.A(n_699),
.Y(n_1046)
);

INVx1_ASAP7_75t_L g1047 ( 
.A(n_626),
.Y(n_1047)
);

CKINVDCx5p33_ASAP7_75t_R g1048 ( 
.A(n_639),
.Y(n_1048)
);

INVx1_ASAP7_75t_L g1049 ( 
.A(n_623),
.Y(n_1049)
);

BUFx2_ASAP7_75t_L g1050 ( 
.A(n_554),
.Y(n_1050)
);

INVxp67_ASAP7_75t_SL g1051 ( 
.A(n_875),
.Y(n_1051)
);

INVxp33_ASAP7_75t_SL g1052 ( 
.A(n_554),
.Y(n_1052)
);

INVx1_ASAP7_75t_L g1053 ( 
.A(n_623),
.Y(n_1053)
);

INVx1_ASAP7_75t_L g1054 ( 
.A(n_635),
.Y(n_1054)
);

CKINVDCx20_ASAP7_75t_R g1055 ( 
.A(n_710),
.Y(n_1055)
);

NOR2xp67_ASAP7_75t_L g1056 ( 
.A(n_875),
.B(n_1),
.Y(n_1056)
);

INVxp67_ASAP7_75t_SL g1057 ( 
.A(n_875),
.Y(n_1057)
);

INVx1_ASAP7_75t_L g1058 ( 
.A(n_627),
.Y(n_1058)
);

CKINVDCx5p33_ASAP7_75t_R g1059 ( 
.A(n_640),
.Y(n_1059)
);

INVx1_ASAP7_75t_L g1060 ( 
.A(n_628),
.Y(n_1060)
);

INVx1_ASAP7_75t_L g1061 ( 
.A(n_631),
.Y(n_1061)
);

INVx2_ASAP7_75t_SL g1062 ( 
.A(n_577),
.Y(n_1062)
);

INVxp33_ASAP7_75t_SL g1063 ( 
.A(n_555),
.Y(n_1063)
);

CKINVDCx16_ASAP7_75t_R g1064 ( 
.A(n_586),
.Y(n_1064)
);

INVx1_ASAP7_75t_L g1065 ( 
.A(n_648),
.Y(n_1065)
);

INVxp67_ASAP7_75t_SL g1066 ( 
.A(n_545),
.Y(n_1066)
);

INVx1_ASAP7_75t_L g1067 ( 
.A(n_655),
.Y(n_1067)
);

INVx1_ASAP7_75t_L g1068 ( 
.A(n_660),
.Y(n_1068)
);

CKINVDCx5p33_ASAP7_75t_R g1069 ( 
.A(n_641),
.Y(n_1069)
);

INVx1_ASAP7_75t_L g1070 ( 
.A(n_668),
.Y(n_1070)
);

HB1xp67_ASAP7_75t_L g1071 ( 
.A(n_555),
.Y(n_1071)
);

INVx1_ASAP7_75t_L g1072 ( 
.A(n_671),
.Y(n_1072)
);

INVx1_ASAP7_75t_L g1073 ( 
.A(n_672),
.Y(n_1073)
);

CKINVDCx20_ASAP7_75t_R g1074 ( 
.A(n_721),
.Y(n_1074)
);

CKINVDCx5p33_ASAP7_75t_R g1075 ( 
.A(n_649),
.Y(n_1075)
);

INVx1_ASAP7_75t_L g1076 ( 
.A(n_682),
.Y(n_1076)
);

INVx2_ASAP7_75t_L g1077 ( 
.A(n_796),
.Y(n_1077)
);

CKINVDCx5p33_ASAP7_75t_R g1078 ( 
.A(n_656),
.Y(n_1078)
);

INVxp67_ASAP7_75t_SL g1079 ( 
.A(n_559),
.Y(n_1079)
);

INVx1_ASAP7_75t_L g1080 ( 
.A(n_696),
.Y(n_1080)
);

INVx1_ASAP7_75t_L g1081 ( 
.A(n_703),
.Y(n_1081)
);

HB1xp67_ASAP7_75t_L g1082 ( 
.A(n_556),
.Y(n_1082)
);

HB1xp67_ASAP7_75t_L g1083 ( 
.A(n_556),
.Y(n_1083)
);

INVx1_ASAP7_75t_L g1084 ( 
.A(n_711),
.Y(n_1084)
);

INVx1_ASAP7_75t_L g1085 ( 
.A(n_712),
.Y(n_1085)
);

BUFx3_ASAP7_75t_L g1086 ( 
.A(n_603),
.Y(n_1086)
);

INVxp33_ASAP7_75t_L g1087 ( 
.A(n_635),
.Y(n_1087)
);

INVxp33_ASAP7_75t_SL g1088 ( 
.A(n_557),
.Y(n_1088)
);

CKINVDCx20_ASAP7_75t_R g1089 ( 
.A(n_722),
.Y(n_1089)
);

INVx1_ASAP7_75t_L g1090 ( 
.A(n_718),
.Y(n_1090)
);

INVx1_ASAP7_75t_L g1091 ( 
.A(n_736),
.Y(n_1091)
);

INVx1_ASAP7_75t_L g1092 ( 
.A(n_738),
.Y(n_1092)
);

INVx1_ASAP7_75t_L g1093 ( 
.A(n_743),
.Y(n_1093)
);

CKINVDCx20_ASAP7_75t_R g1094 ( 
.A(n_737),
.Y(n_1094)
);

INVxp33_ASAP7_75t_SL g1095 ( 
.A(n_557),
.Y(n_1095)
);

INVx1_ASAP7_75t_L g1096 ( 
.A(n_746),
.Y(n_1096)
);

INVx1_ASAP7_75t_L g1097 ( 
.A(n_748),
.Y(n_1097)
);

INVx1_ASAP7_75t_L g1098 ( 
.A(n_752),
.Y(n_1098)
);

OR2x2_ASAP7_75t_L g1099 ( 
.A(n_755),
.B(n_1),
.Y(n_1099)
);

INVx1_ASAP7_75t_L g1100 ( 
.A(n_756),
.Y(n_1100)
);

CKINVDCx5p33_ASAP7_75t_R g1101 ( 
.A(n_659),
.Y(n_1101)
);

INVx1_ASAP7_75t_L g1102 ( 
.A(n_757),
.Y(n_1102)
);

BUFx3_ASAP7_75t_L g1103 ( 
.A(n_603),
.Y(n_1103)
);

INVx2_ASAP7_75t_L g1104 ( 
.A(n_796),
.Y(n_1104)
);

INVx1_ASAP7_75t_L g1105 ( 
.A(n_762),
.Y(n_1105)
);

INVx1_ASAP7_75t_L g1106 ( 
.A(n_763),
.Y(n_1106)
);

INVx1_ASAP7_75t_L g1107 ( 
.A(n_765),
.Y(n_1107)
);

INVx1_ASAP7_75t_L g1108 ( 
.A(n_767),
.Y(n_1108)
);

INVx1_ASAP7_75t_L g1109 ( 
.A(n_770),
.Y(n_1109)
);

INVx2_ASAP7_75t_SL g1110 ( 
.A(n_586),
.Y(n_1110)
);

INVx1_ASAP7_75t_L g1111 ( 
.A(n_790),
.Y(n_1111)
);

INVx1_ASAP7_75t_L g1112 ( 
.A(n_802),
.Y(n_1112)
);

INVx1_ASAP7_75t_L g1113 ( 
.A(n_822),
.Y(n_1113)
);

CKINVDCx5p33_ASAP7_75t_R g1114 ( 
.A(n_663),
.Y(n_1114)
);

CKINVDCx16_ASAP7_75t_R g1115 ( 
.A(n_586),
.Y(n_1115)
);

INVx1_ASAP7_75t_L g1116 ( 
.A(n_830),
.Y(n_1116)
);

INVx1_ASAP7_75t_L g1117 ( 
.A(n_838),
.Y(n_1117)
);

INVx1_ASAP7_75t_L g1118 ( 
.A(n_841),
.Y(n_1118)
);

CKINVDCx5p33_ASAP7_75t_R g1119 ( 
.A(n_664),
.Y(n_1119)
);

CKINVDCx5p33_ASAP7_75t_R g1120 ( 
.A(n_665),
.Y(n_1120)
);

INVx1_ASAP7_75t_L g1121 ( 
.A(n_851),
.Y(n_1121)
);

INVx1_ASAP7_75t_L g1122 ( 
.A(n_852),
.Y(n_1122)
);

INVx1_ASAP7_75t_L g1123 ( 
.A(n_867),
.Y(n_1123)
);

INVx2_ASAP7_75t_L g1124 ( 
.A(n_796),
.Y(n_1124)
);

INVx1_ASAP7_75t_L g1125 ( 
.A(n_877),
.Y(n_1125)
);

INVx2_ASAP7_75t_L g1126 ( 
.A(n_796),
.Y(n_1126)
);

HB1xp67_ASAP7_75t_L g1127 ( 
.A(n_558),
.Y(n_1127)
);

CKINVDCx5p33_ASAP7_75t_R g1128 ( 
.A(n_675),
.Y(n_1128)
);

INVx1_ASAP7_75t_L g1129 ( 
.A(n_879),
.Y(n_1129)
);

INVxp67_ASAP7_75t_SL g1130 ( 
.A(n_591),
.Y(n_1130)
);

INVx1_ASAP7_75t_L g1131 ( 
.A(n_881),
.Y(n_1131)
);

INVx1_ASAP7_75t_L g1132 ( 
.A(n_882),
.Y(n_1132)
);

CKINVDCx16_ASAP7_75t_R g1133 ( 
.A(n_617),
.Y(n_1133)
);

INVx1_ASAP7_75t_L g1134 ( 
.A(n_886),
.Y(n_1134)
);

INVx1_ASAP7_75t_L g1135 ( 
.A(n_888),
.Y(n_1135)
);

INVxp33_ASAP7_75t_SL g1136 ( 
.A(n_558),
.Y(n_1136)
);

INVx2_ASAP7_75t_L g1137 ( 
.A(n_796),
.Y(n_1137)
);

INVx1_ASAP7_75t_L g1138 ( 
.A(n_897),
.Y(n_1138)
);

INVx1_ASAP7_75t_L g1139 ( 
.A(n_910),
.Y(n_1139)
);

INVx1_ASAP7_75t_L g1140 ( 
.A(n_917),
.Y(n_1140)
);

CKINVDCx5p33_ASAP7_75t_R g1141 ( 
.A(n_676),
.Y(n_1141)
);

INVxp67_ASAP7_75t_SL g1142 ( 
.A(n_596),
.Y(n_1142)
);

INVxp67_ASAP7_75t_SL g1143 ( 
.A(n_600),
.Y(n_1143)
);

CKINVDCx5p33_ASAP7_75t_R g1144 ( 
.A(n_681),
.Y(n_1144)
);

CKINVDCx20_ASAP7_75t_R g1145 ( 
.A(n_769),
.Y(n_1145)
);

INVxp33_ASAP7_75t_SL g1146 ( 
.A(n_560),
.Y(n_1146)
);

INVx1_ASAP7_75t_L g1147 ( 
.A(n_918),
.Y(n_1147)
);

CKINVDCx5p33_ASAP7_75t_R g1148 ( 
.A(n_683),
.Y(n_1148)
);

CKINVDCx5p33_ASAP7_75t_R g1149 ( 
.A(n_685),
.Y(n_1149)
);

CKINVDCx5p33_ASAP7_75t_R g1150 ( 
.A(n_688),
.Y(n_1150)
);

CKINVDCx5p33_ASAP7_75t_R g1151 ( 
.A(n_691),
.Y(n_1151)
);

INVx1_ASAP7_75t_L g1152 ( 
.A(n_920),
.Y(n_1152)
);

INVx1_ASAP7_75t_L g1153 ( 
.A(n_922),
.Y(n_1153)
);

INVx1_ASAP7_75t_L g1154 ( 
.A(n_929),
.Y(n_1154)
);

INVx2_ASAP7_75t_L g1155 ( 
.A(n_796),
.Y(n_1155)
);

INVxp67_ASAP7_75t_SL g1156 ( 
.A(n_609),
.Y(n_1156)
);

INVx1_ASAP7_75t_L g1157 ( 
.A(n_931),
.Y(n_1157)
);

INVx1_ASAP7_75t_L g1158 ( 
.A(n_952),
.Y(n_1158)
);

CKINVDCx5p33_ASAP7_75t_R g1159 ( 
.A(n_695),
.Y(n_1159)
);

CKINVDCx16_ASAP7_75t_R g1160 ( 
.A(n_617),
.Y(n_1160)
);

INVx1_ASAP7_75t_L g1161 ( 
.A(n_953),
.Y(n_1161)
);

INVx1_ASAP7_75t_L g1162 ( 
.A(n_954),
.Y(n_1162)
);

INVx1_ASAP7_75t_L g1163 ( 
.A(n_956),
.Y(n_1163)
);

CKINVDCx5p33_ASAP7_75t_R g1164 ( 
.A(n_697),
.Y(n_1164)
);

INVx1_ASAP7_75t_L g1165 ( 
.A(n_611),
.Y(n_1165)
);

INVx1_ASAP7_75t_L g1166 ( 
.A(n_624),
.Y(n_1166)
);

INVx1_ASAP7_75t_L g1167 ( 
.A(n_632),
.Y(n_1167)
);

INVx1_ASAP7_75t_L g1168 ( 
.A(n_634),
.Y(n_1168)
);

INVx1_ASAP7_75t_L g1169 ( 
.A(n_642),
.Y(n_1169)
);

CKINVDCx5p33_ASAP7_75t_R g1170 ( 
.A(n_704),
.Y(n_1170)
);

INVxp33_ASAP7_75t_SL g1171 ( 
.A(n_560),
.Y(n_1171)
);

CKINVDCx20_ASAP7_75t_R g1172 ( 
.A(n_850),
.Y(n_1172)
);

CKINVDCx16_ASAP7_75t_R g1173 ( 
.A(n_617),
.Y(n_1173)
);

INVx2_ASAP7_75t_L g1174 ( 
.A(n_646),
.Y(n_1174)
);

INVxp67_ASAP7_75t_SL g1175 ( 
.A(n_643),
.Y(n_1175)
);

INVxp33_ASAP7_75t_L g1176 ( 
.A(n_646),
.Y(n_1176)
);

INVx1_ASAP7_75t_L g1177 ( 
.A(n_644),
.Y(n_1177)
);

INVx1_ASAP7_75t_L g1178 ( 
.A(n_650),
.Y(n_1178)
);

INVx1_ASAP7_75t_L g1179 ( 
.A(n_653),
.Y(n_1179)
);

INVx1_ASAP7_75t_L g1180 ( 
.A(n_661),
.Y(n_1180)
);

BUFx3_ASAP7_75t_L g1181 ( 
.A(n_717),
.Y(n_1181)
);

INVx1_ASAP7_75t_L g1182 ( 
.A(n_678),
.Y(n_1182)
);

INVx1_ASAP7_75t_L g1183 ( 
.A(n_690),
.Y(n_1183)
);

INVx1_ASAP7_75t_L g1184 ( 
.A(n_708),
.Y(n_1184)
);

INVx1_ASAP7_75t_L g1185 ( 
.A(n_723),
.Y(n_1185)
);

INVx1_ASAP7_75t_SL g1186 ( 
.A(n_861),
.Y(n_1186)
);

INVx1_ASAP7_75t_L g1187 ( 
.A(n_726),
.Y(n_1187)
);

BUFx3_ASAP7_75t_L g1188 ( 
.A(n_717),
.Y(n_1188)
);

INVx1_ASAP7_75t_L g1189 ( 
.A(n_731),
.Y(n_1189)
);

CKINVDCx20_ASAP7_75t_R g1190 ( 
.A(n_880),
.Y(n_1190)
);

INVxp33_ASAP7_75t_SL g1191 ( 
.A(n_565),
.Y(n_1191)
);

INVx1_ASAP7_75t_L g1192 ( 
.A(n_733),
.Y(n_1192)
);

INVx1_ASAP7_75t_L g1193 ( 
.A(n_739),
.Y(n_1193)
);

INVx1_ASAP7_75t_L g1194 ( 
.A(n_702),
.Y(n_1194)
);

CKINVDCx5p33_ASAP7_75t_R g1195 ( 
.A(n_705),
.Y(n_1195)
);

INVxp33_ASAP7_75t_SL g1196 ( 
.A(n_565),
.Y(n_1196)
);

INVx1_ASAP7_75t_L g1197 ( 
.A(n_751),
.Y(n_1197)
);

INVx1_ASAP7_75t_L g1198 ( 
.A(n_754),
.Y(n_1198)
);

CKINVDCx5p33_ASAP7_75t_R g1199 ( 
.A(n_709),
.Y(n_1199)
);

INVxp33_ASAP7_75t_SL g1200 ( 
.A(n_567),
.Y(n_1200)
);

INVx1_ASAP7_75t_L g1201 ( 
.A(n_761),
.Y(n_1201)
);

INVxp67_ASAP7_75t_L g1202 ( 
.A(n_638),
.Y(n_1202)
);

INVx1_ASAP7_75t_L g1203 ( 
.A(n_766),
.Y(n_1203)
);

INVxp67_ASAP7_75t_L g1204 ( 
.A(n_638),
.Y(n_1204)
);

INVx1_ASAP7_75t_L g1205 ( 
.A(n_768),
.Y(n_1205)
);

INVx1_ASAP7_75t_L g1206 ( 
.A(n_813),
.Y(n_1206)
);

INVx1_ASAP7_75t_L g1207 ( 
.A(n_819),
.Y(n_1207)
);

INVx2_ASAP7_75t_L g1208 ( 
.A(n_702),
.Y(n_1208)
);

INVxp33_ASAP7_75t_SL g1209 ( 
.A(n_567),
.Y(n_1209)
);

INVxp67_ASAP7_75t_SL g1210 ( 
.A(n_837),
.Y(n_1210)
);

INVx1_ASAP7_75t_L g1211 ( 
.A(n_857),
.Y(n_1211)
);

INVxp67_ASAP7_75t_L g1212 ( 
.A(n_638),
.Y(n_1212)
);

INVx1_ASAP7_75t_L g1213 ( 
.A(n_859),
.Y(n_1213)
);

INVx1_ASAP7_75t_L g1214 ( 
.A(n_890),
.Y(n_1214)
);

INVx1_ASAP7_75t_L g1215 ( 
.A(n_893),
.Y(n_1215)
);

INVx1_ASAP7_75t_L g1216 ( 
.A(n_900),
.Y(n_1216)
);

INVx1_ASAP7_75t_L g1217 ( 
.A(n_906),
.Y(n_1217)
);

INVx2_ASAP7_75t_SL g1218 ( 
.A(n_666),
.Y(n_1218)
);

INVxp67_ASAP7_75t_SL g1219 ( 
.A(n_914),
.Y(n_1219)
);

INVxp67_ASAP7_75t_L g1220 ( 
.A(n_666),
.Y(n_1220)
);

INVx1_ASAP7_75t_L g1221 ( 
.A(n_923),
.Y(n_1221)
);

INVx1_ASAP7_75t_L g1222 ( 
.A(n_925),
.Y(n_1222)
);

INVx2_ASAP7_75t_L g1223 ( 
.A(n_794),
.Y(n_1223)
);

INVx2_ASAP7_75t_SL g1224 ( 
.A(n_666),
.Y(n_1224)
);

CKINVDCx16_ASAP7_75t_R g1225 ( 
.A(n_674),
.Y(n_1225)
);

INVx1_ASAP7_75t_L g1226 ( 
.A(n_944),
.Y(n_1226)
);

INVx1_ASAP7_75t_L g1227 ( 
.A(n_958),
.Y(n_1227)
);

INVx1_ASAP7_75t_L g1228 ( 
.A(n_605),
.Y(n_1228)
);

BUFx3_ASAP7_75t_L g1229 ( 
.A(n_717),
.Y(n_1229)
);

INVx1_ASAP7_75t_L g1230 ( 
.A(n_605),
.Y(n_1230)
);

INVx2_ASAP7_75t_L g1231 ( 
.A(n_794),
.Y(n_1231)
);

INVx2_ASAP7_75t_L g1232 ( 
.A(n_843),
.Y(n_1232)
);

CKINVDCx16_ASAP7_75t_R g1233 ( 
.A(n_674),
.Y(n_1233)
);

INVx1_ASAP7_75t_L g1234 ( 
.A(n_684),
.Y(n_1234)
);

BUFx6f_ASAP7_75t_L g1235 ( 
.A(n_679),
.Y(n_1235)
);

INVx2_ASAP7_75t_L g1236 ( 
.A(n_843),
.Y(n_1236)
);

INVx1_ASAP7_75t_L g1237 ( 
.A(n_684),
.Y(n_1237)
);

CKINVDCx20_ASAP7_75t_R g1238 ( 
.A(n_949),
.Y(n_1238)
);

CKINVDCx16_ASAP7_75t_R g1239 ( 
.A(n_674),
.Y(n_1239)
);

INVx1_ASAP7_75t_L g1240 ( 
.A(n_694),
.Y(n_1240)
);

INVxp67_ASAP7_75t_SL g1241 ( 
.A(n_694),
.Y(n_1241)
);

INVx1_ASAP7_75t_L g1242 ( 
.A(n_759),
.Y(n_1242)
);

CKINVDCx20_ASAP7_75t_R g1243 ( 
.A(n_572),
.Y(n_1243)
);

INVx1_ASAP7_75t_L g1244 ( 
.A(n_759),
.Y(n_1244)
);

CKINVDCx14_ASAP7_75t_R g1245 ( 
.A(n_835),
.Y(n_1245)
);

INVx1_ASAP7_75t_L g1246 ( 
.A(n_936),
.Y(n_1246)
);

INVx2_ASAP7_75t_L g1247 ( 
.A(n_854),
.Y(n_1247)
);

CKINVDCx14_ASAP7_75t_R g1248 ( 
.A(n_835),
.Y(n_1248)
);

BUFx6f_ASAP7_75t_L g1249 ( 
.A(n_679),
.Y(n_1249)
);

INVx2_ASAP7_75t_L g1250 ( 
.A(n_854),
.Y(n_1250)
);

INVxp67_ASAP7_75t_L g1251 ( 
.A(n_732),
.Y(n_1251)
);

INVx1_ASAP7_75t_L g1252 ( 
.A(n_936),
.Y(n_1252)
);

INVx1_ASAP7_75t_L g1253 ( 
.A(n_855),
.Y(n_1253)
);

CKINVDCx5p33_ASAP7_75t_R g1254 ( 
.A(n_716),
.Y(n_1254)
);

INVx1_ASAP7_75t_L g1255 ( 
.A(n_855),
.Y(n_1255)
);

CKINVDCx5p33_ASAP7_75t_R g1256 ( 
.A(n_719),
.Y(n_1256)
);

INVx1_ASAP7_75t_L g1257 ( 
.A(n_894),
.Y(n_1257)
);

INVx1_ASAP7_75t_L g1258 ( 
.A(n_894),
.Y(n_1258)
);

HB1xp67_ASAP7_75t_L g1259 ( 
.A(n_572),
.Y(n_1259)
);

CKINVDCx5p33_ASAP7_75t_R g1260 ( 
.A(n_720),
.Y(n_1260)
);

INVx1_ASAP7_75t_L g1261 ( 
.A(n_905),
.Y(n_1261)
);

BUFx3_ASAP7_75t_L g1262 ( 
.A(n_835),
.Y(n_1262)
);

CKINVDCx5p33_ASAP7_75t_R g1263 ( 
.A(n_729),
.Y(n_1263)
);

INVx1_ASAP7_75t_L g1264 ( 
.A(n_905),
.Y(n_1264)
);

INVx1_ASAP7_75t_L g1265 ( 
.A(n_669),
.Y(n_1265)
);

INVx1_ASAP7_75t_L g1266 ( 
.A(n_669),
.Y(n_1266)
);

INVx1_ASAP7_75t_L g1267 ( 
.A(n_728),
.Y(n_1267)
);

INVxp33_ASAP7_75t_L g1268 ( 
.A(n_679),
.Y(n_1268)
);

INVx1_ASAP7_75t_L g1269 ( 
.A(n_728),
.Y(n_1269)
);

INVx1_ASAP7_75t_L g1270 ( 
.A(n_784),
.Y(n_1270)
);

INVx1_ASAP7_75t_L g1271 ( 
.A(n_784),
.Y(n_1271)
);

INVx1_ASAP7_75t_L g1272 ( 
.A(n_811),
.Y(n_1272)
);

INVx1_ASAP7_75t_L g1273 ( 
.A(n_811),
.Y(n_1273)
);

INVx1_ASAP7_75t_L g1274 ( 
.A(n_864),
.Y(n_1274)
);

INVx1_ASAP7_75t_L g1275 ( 
.A(n_864),
.Y(n_1275)
);

INVx1_ASAP7_75t_L g1276 ( 
.A(n_942),
.Y(n_1276)
);

INVx1_ASAP7_75t_L g1277 ( 
.A(n_942),
.Y(n_1277)
);

INVx1_ASAP7_75t_L g1278 ( 
.A(n_732),
.Y(n_1278)
);

INVx1_ASAP7_75t_L g1279 ( 
.A(n_732),
.Y(n_1279)
);

CKINVDCx5p33_ASAP7_75t_R g1280 ( 
.A(n_734),
.Y(n_1280)
);

INVx1_ASAP7_75t_L g1281 ( 
.A(n_806),
.Y(n_1281)
);

INVxp33_ASAP7_75t_SL g1282 ( 
.A(n_574),
.Y(n_1282)
);

INVx2_ASAP7_75t_L g1283 ( 
.A(n_679),
.Y(n_1283)
);

INVx1_ASAP7_75t_L g1284 ( 
.A(n_806),
.Y(n_1284)
);

INVx1_ASAP7_75t_L g1285 ( 
.A(n_806),
.Y(n_1285)
);

INVx1_ASAP7_75t_L g1286 ( 
.A(n_911),
.Y(n_1286)
);

INVx1_ASAP7_75t_L g1287 ( 
.A(n_911),
.Y(n_1287)
);

INVx1_ASAP7_75t_L g1288 ( 
.A(n_911),
.Y(n_1288)
);

INVxp33_ASAP7_75t_L g1289 ( 
.A(n_679),
.Y(n_1289)
);

BUFx6f_ASAP7_75t_L g1290 ( 
.A(n_812),
.Y(n_1290)
);

INVx2_ASAP7_75t_L g1291 ( 
.A(n_812),
.Y(n_1291)
);

INVx2_ASAP7_75t_L g1292 ( 
.A(n_812),
.Y(n_1292)
);

CKINVDCx14_ASAP7_75t_R g1293 ( 
.A(n_544),
.Y(n_1293)
);

NOR2xp33_ASAP7_75t_L g1294 ( 
.A(n_547),
.B(n_2),
.Y(n_1294)
);

CKINVDCx20_ASAP7_75t_R g1295 ( 
.A(n_574),
.Y(n_1295)
);

INVx1_ASAP7_75t_L g1296 ( 
.A(n_645),
.Y(n_1296)
);

INVx1_ASAP7_75t_L g1297 ( 
.A(n_645),
.Y(n_1297)
);

INVx1_ASAP7_75t_L g1298 ( 
.A(n_698),
.Y(n_1298)
);

INVx1_ASAP7_75t_L g1299 ( 
.A(n_698),
.Y(n_1299)
);

INVx1_ASAP7_75t_L g1300 ( 
.A(n_725),
.Y(n_1300)
);

INVx1_ASAP7_75t_L g1301 ( 
.A(n_725),
.Y(n_1301)
);

INVx1_ASAP7_75t_L g1302 ( 
.A(n_735),
.Y(n_1302)
);

INVx1_ASAP7_75t_L g1303 ( 
.A(n_735),
.Y(n_1303)
);

INVx1_ASAP7_75t_L g1304 ( 
.A(n_760),
.Y(n_1304)
);

INVx2_ASAP7_75t_L g1305 ( 
.A(n_812),
.Y(n_1305)
);

INVx1_ASAP7_75t_SL g1306 ( 
.A(n_546),
.Y(n_1306)
);

INVx1_ASAP7_75t_L g1307 ( 
.A(n_760),
.Y(n_1307)
);

INVx1_ASAP7_75t_L g1308 ( 
.A(n_814),
.Y(n_1308)
);

INVxp67_ASAP7_75t_SL g1309 ( 
.A(n_621),
.Y(n_1309)
);

CKINVDCx20_ASAP7_75t_R g1310 ( 
.A(n_575),
.Y(n_1310)
);

INVx1_ASAP7_75t_L g1311 ( 
.A(n_814),
.Y(n_1311)
);

INVx2_ASAP7_75t_L g1312 ( 
.A(n_812),
.Y(n_1312)
);

CKINVDCx5p33_ASAP7_75t_R g1313 ( 
.A(n_742),
.Y(n_1313)
);

BUFx3_ASAP7_75t_L g1314 ( 
.A(n_544),
.Y(n_1314)
);

INVx1_ASAP7_75t_L g1315 ( 
.A(n_745),
.Y(n_1315)
);

INVx1_ASAP7_75t_L g1316 ( 
.A(n_747),
.Y(n_1316)
);

CKINVDCx5p33_ASAP7_75t_R g1317 ( 
.A(n_753),
.Y(n_1317)
);

INVx1_ASAP7_75t_L g1318 ( 
.A(n_758),
.Y(n_1318)
);

INVx1_ASAP7_75t_L g1319 ( 
.A(n_771),
.Y(n_1319)
);

INVxp67_ASAP7_75t_SL g1320 ( 
.A(n_749),
.Y(n_1320)
);

CKINVDCx5p33_ASAP7_75t_R g1321 ( 
.A(n_772),
.Y(n_1321)
);

HB1xp67_ASAP7_75t_L g1322 ( 
.A(n_575),
.Y(n_1322)
);

CKINVDCx14_ASAP7_75t_R g1323 ( 
.A(n_549),
.Y(n_1323)
);

CKINVDCx16_ASAP7_75t_R g1324 ( 
.A(n_548),
.Y(n_1324)
);

INVx1_ASAP7_75t_L g1325 ( 
.A(n_777),
.Y(n_1325)
);

INVx2_ASAP7_75t_L g1326 ( 
.A(n_821),
.Y(n_1326)
);

INVxp67_ASAP7_75t_L g1327 ( 
.A(n_580),
.Y(n_1327)
);

INVx1_ASAP7_75t_L g1328 ( 
.A(n_782),
.Y(n_1328)
);

CKINVDCx20_ASAP7_75t_R g1329 ( 
.A(n_580),
.Y(n_1329)
);

BUFx2_ASAP7_75t_L g1330 ( 
.A(n_589),
.Y(n_1330)
);

INVx1_ASAP7_75t_L g1331 ( 
.A(n_783),
.Y(n_1331)
);

INVx1_ASAP7_75t_L g1332 ( 
.A(n_788),
.Y(n_1332)
);

INVx2_ASAP7_75t_L g1333 ( 
.A(n_821),
.Y(n_1333)
);

INVx1_ASAP7_75t_L g1334 ( 
.A(n_789),
.Y(n_1334)
);

INVx1_ASAP7_75t_L g1335 ( 
.A(n_821),
.Y(n_1335)
);

CKINVDCx20_ASAP7_75t_R g1336 ( 
.A(n_589),
.Y(n_1336)
);

INVxp67_ASAP7_75t_L g1337 ( 
.A(n_590),
.Y(n_1337)
);

CKINVDCx16_ASAP7_75t_R g1338 ( 
.A(n_633),
.Y(n_1338)
);

BUFx12f_ASAP7_75t_L g1339 ( 
.A(n_970),
.Y(n_1339)
);

INVx4_ASAP7_75t_L g1340 ( 
.A(n_1022),
.Y(n_1340)
);

AND2x2_ASAP7_75t_L g1341 ( 
.A(n_1314),
.B(n_571),
.Y(n_1341)
);

AND2x2_ASAP7_75t_L g1342 ( 
.A(n_1314),
.B(n_619),
.Y(n_1342)
);

BUFx2_ASAP7_75t_L g1343 ( 
.A(n_1003),
.Y(n_1343)
);

AND2x2_ASAP7_75t_L g1344 ( 
.A(n_1042),
.B(n_630),
.Y(n_1344)
);

BUFx8_ASAP7_75t_SL g1345 ( 
.A(n_970),
.Y(n_1345)
);

BUFx6f_ASAP7_75t_L g1346 ( 
.A(n_1235),
.Y(n_1346)
);

AND2x2_ASAP7_75t_L g1347 ( 
.A(n_1042),
.B(n_692),
.Y(n_1347)
);

AND2x4_ASAP7_75t_L g1348 ( 
.A(n_1086),
.B(n_707),
.Y(n_1348)
);

NOR2xp33_ASAP7_75t_L g1349 ( 
.A(n_1051),
.B(n_773),
.Y(n_1349)
);

BUFx2_ASAP7_75t_L g1350 ( 
.A(n_1003),
.Y(n_1350)
);

AND2x2_ASAP7_75t_L g1351 ( 
.A(n_1245),
.B(n_1248),
.Y(n_1351)
);

INVx3_ASAP7_75t_L g1352 ( 
.A(n_1024),
.Y(n_1352)
);

BUFx6f_ASAP7_75t_L g1353 ( 
.A(n_1235),
.Y(n_1353)
);

AND2x6_ASAP7_75t_L g1354 ( 
.A(n_961),
.B(n_821),
.Y(n_1354)
);

NAND2xp5_ASAP7_75t_L g1355 ( 
.A(n_1016),
.B(n_636),
.Y(n_1355)
);

INVx1_ASAP7_75t_L g1356 ( 
.A(n_1011),
.Y(n_1356)
);

NAND2xp5_ASAP7_75t_L g1357 ( 
.A(n_1057),
.B(n_647),
.Y(n_1357)
);

BUFx3_ASAP7_75t_L g1358 ( 
.A(n_997),
.Y(n_1358)
);

NAND2xp5_ASAP7_75t_L g1359 ( 
.A(n_1315),
.B(n_651),
.Y(n_1359)
);

BUFx8_ASAP7_75t_L g1360 ( 
.A(n_1030),
.Y(n_1360)
);

HB1xp67_ASAP7_75t_L g1361 ( 
.A(n_1306),
.Y(n_1361)
);

INVx2_ASAP7_75t_L g1362 ( 
.A(n_1000),
.Y(n_1362)
);

NAND2xp5_ASAP7_75t_L g1363 ( 
.A(n_1316),
.B(n_652),
.Y(n_1363)
);

AND2x4_ASAP7_75t_L g1364 ( 
.A(n_1086),
.B(n_1103),
.Y(n_1364)
);

AND2x4_ASAP7_75t_L g1365 ( 
.A(n_1103),
.B(n_872),
.Y(n_1365)
);

AND2x4_ASAP7_75t_L g1366 ( 
.A(n_1181),
.B(n_907),
.Y(n_1366)
);

BUFx2_ASAP7_75t_L g1367 ( 
.A(n_1243),
.Y(n_1367)
);

BUFx6f_ASAP7_75t_L g1368 ( 
.A(n_1235),
.Y(n_1368)
);

NAND2xp5_ASAP7_75t_L g1369 ( 
.A(n_1318),
.B(n_654),
.Y(n_1369)
);

AND2x2_ASAP7_75t_L g1370 ( 
.A(n_1245),
.B(n_946),
.Y(n_1370)
);

INVx2_ASAP7_75t_L g1371 ( 
.A(n_1000),
.Y(n_1371)
);

AND2x2_ASAP7_75t_L g1372 ( 
.A(n_1248),
.B(n_957),
.Y(n_1372)
);

INVx2_ASAP7_75t_L g1373 ( 
.A(n_1001),
.Y(n_1373)
);

BUFx6f_ASAP7_75t_L g1374 ( 
.A(n_1235),
.Y(n_1374)
);

INVx1_ASAP7_75t_L g1375 ( 
.A(n_1012),
.Y(n_1375)
);

BUFx6f_ASAP7_75t_L g1376 ( 
.A(n_1249),
.Y(n_1376)
);

BUFx6f_ASAP7_75t_L g1377 ( 
.A(n_1249),
.Y(n_1377)
);

INVx2_ASAP7_75t_L g1378 ( 
.A(n_1001),
.Y(n_1378)
);

INVx2_ASAP7_75t_L g1379 ( 
.A(n_1015),
.Y(n_1379)
);

NAND2xp5_ASAP7_75t_L g1380 ( 
.A(n_1319),
.B(n_1325),
.Y(n_1380)
);

AND2x4_ASAP7_75t_L g1381 ( 
.A(n_1181),
.B(n_549),
.Y(n_1381)
);

NAND2xp5_ASAP7_75t_L g1382 ( 
.A(n_1328),
.B(n_657),
.Y(n_1382)
);

NAND2xp5_ASAP7_75t_L g1383 ( 
.A(n_1331),
.B(n_658),
.Y(n_1383)
);

AND2x4_ASAP7_75t_L g1384 ( 
.A(n_1188),
.B(n_1229),
.Y(n_1384)
);

BUFx6f_ASAP7_75t_L g1385 ( 
.A(n_1249),
.Y(n_1385)
);

HB1xp67_ASAP7_75t_L g1386 ( 
.A(n_994),
.Y(n_1386)
);

AND2x2_ASAP7_75t_L g1387 ( 
.A(n_1327),
.B(n_550),
.Y(n_1387)
);

INVx1_ASAP7_75t_L g1388 ( 
.A(n_1013),
.Y(n_1388)
);

NAND2xp5_ASAP7_75t_L g1389 ( 
.A(n_1332),
.B(n_1334),
.Y(n_1389)
);

NAND2xp5_ASAP7_75t_L g1390 ( 
.A(n_1293),
.B(n_662),
.Y(n_1390)
);

NOR2xp33_ASAP7_75t_L g1391 ( 
.A(n_975),
.B(n_550),
.Y(n_1391)
);

AND2x4_ASAP7_75t_L g1392 ( 
.A(n_1188),
.B(n_553),
.Y(n_1392)
);

NAND2xp5_ASAP7_75t_L g1393 ( 
.A(n_1293),
.B(n_667),
.Y(n_1393)
);

BUFx6f_ASAP7_75t_L g1394 ( 
.A(n_1249),
.Y(n_1394)
);

NAND2xp5_ASAP7_75t_L g1395 ( 
.A(n_1323),
.B(n_670),
.Y(n_1395)
);

BUFx3_ASAP7_75t_L g1396 ( 
.A(n_997),
.Y(n_1396)
);

INVx4_ASAP7_75t_L g1397 ( 
.A(n_1022),
.Y(n_1397)
);

AND2x2_ASAP7_75t_L g1398 ( 
.A(n_1337),
.B(n_553),
.Y(n_1398)
);

AND2x6_ASAP7_75t_L g1399 ( 
.A(n_961),
.B(n_821),
.Y(n_1399)
);

BUFx3_ASAP7_75t_L g1400 ( 
.A(n_1004),
.Y(n_1400)
);

BUFx6f_ASAP7_75t_L g1401 ( 
.A(n_1290),
.Y(n_1401)
);

NAND2xp5_ASAP7_75t_SL g1402 ( 
.A(n_1056),
.B(n_793),
.Y(n_1402)
);

BUFx3_ASAP7_75t_L g1403 ( 
.A(n_1004),
.Y(n_1403)
);

INVx1_ASAP7_75t_L g1404 ( 
.A(n_1014),
.Y(n_1404)
);

NAND2xp5_ASAP7_75t_L g1405 ( 
.A(n_1323),
.B(n_686),
.Y(n_1405)
);

BUFx3_ASAP7_75t_L g1406 ( 
.A(n_1005),
.Y(n_1406)
);

BUFx6f_ASAP7_75t_L g1407 ( 
.A(n_1290),
.Y(n_1407)
);

BUFx3_ASAP7_75t_L g1408 ( 
.A(n_1005),
.Y(n_1408)
);

BUFx6f_ASAP7_75t_L g1409 ( 
.A(n_1290),
.Y(n_1409)
);

AND2x2_ASAP7_75t_L g1410 ( 
.A(n_971),
.B(n_561),
.Y(n_1410)
);

NAND2xp5_ASAP7_75t_L g1411 ( 
.A(n_1066),
.B(n_693),
.Y(n_1411)
);

INVx5_ASAP7_75t_L g1412 ( 
.A(n_1024),
.Y(n_1412)
);

BUFx3_ASAP7_75t_L g1413 ( 
.A(n_1024),
.Y(n_1413)
);

INVx2_ASAP7_75t_L g1414 ( 
.A(n_1015),
.Y(n_1414)
);

NOR2xp33_ASAP7_75t_L g1415 ( 
.A(n_1241),
.B(n_561),
.Y(n_1415)
);

AND2x4_ASAP7_75t_L g1416 ( 
.A(n_1229),
.B(n_1262),
.Y(n_1416)
);

NOR2xp33_ASAP7_75t_L g1417 ( 
.A(n_1294),
.B(n_566),
.Y(n_1417)
);

BUFx6f_ASAP7_75t_L g1418 ( 
.A(n_1283),
.Y(n_1418)
);

INVx2_ASAP7_75t_L g1419 ( 
.A(n_998),
.Y(n_1419)
);

BUFx6f_ASAP7_75t_L g1420 ( 
.A(n_1283),
.Y(n_1420)
);

AND2x4_ASAP7_75t_L g1421 ( 
.A(n_1262),
.B(n_1278),
.Y(n_1421)
);

AND2x2_ASAP7_75t_L g1422 ( 
.A(n_1087),
.B(n_566),
.Y(n_1422)
);

NOR2xp33_ASAP7_75t_L g1423 ( 
.A(n_1079),
.B(n_568),
.Y(n_1423)
);

BUFx6f_ASAP7_75t_L g1424 ( 
.A(n_1291),
.Y(n_1424)
);

INVx5_ASAP7_75t_L g1425 ( 
.A(n_1291),
.Y(n_1425)
);

NOR2xp33_ASAP7_75t_L g1426 ( 
.A(n_1130),
.B(n_568),
.Y(n_1426)
);

AND2x2_ASAP7_75t_L g1427 ( 
.A(n_1087),
.B(n_569),
.Y(n_1427)
);

BUFx3_ASAP7_75t_L g1428 ( 
.A(n_984),
.Y(n_1428)
);

NAND2xp5_ASAP7_75t_L g1429 ( 
.A(n_1142),
.B(n_700),
.Y(n_1429)
);

BUFx6f_ASAP7_75t_L g1430 ( 
.A(n_1292),
.Y(n_1430)
);

HB1xp67_ASAP7_75t_L g1431 ( 
.A(n_1010),
.Y(n_1431)
);

BUFx6f_ASAP7_75t_L g1432 ( 
.A(n_1292),
.Y(n_1432)
);

AND2x4_ASAP7_75t_L g1433 ( 
.A(n_1279),
.B(n_569),
.Y(n_1433)
);

INVx3_ASAP7_75t_L g1434 ( 
.A(n_1174),
.Y(n_1434)
);

NOR2xp33_ASAP7_75t_L g1435 ( 
.A(n_1143),
.B(n_570),
.Y(n_1435)
);

NOR2xp33_ASAP7_75t_L g1436 ( 
.A(n_1156),
.B(n_1175),
.Y(n_1436)
);

AND2x4_ASAP7_75t_L g1437 ( 
.A(n_1281),
.B(n_570),
.Y(n_1437)
);

NAND2xp5_ASAP7_75t_L g1438 ( 
.A(n_1210),
.B(n_701),
.Y(n_1438)
);

INVx2_ASAP7_75t_L g1439 ( 
.A(n_998),
.Y(n_1439)
);

BUFx12f_ASAP7_75t_L g1440 ( 
.A(n_972),
.Y(n_1440)
);

INVx2_ASAP7_75t_L g1441 ( 
.A(n_1305),
.Y(n_1441)
);

INVx5_ASAP7_75t_L g1442 ( 
.A(n_1305),
.Y(n_1442)
);

BUFx6f_ASAP7_75t_L g1443 ( 
.A(n_1312),
.Y(n_1443)
);

BUFx12f_ASAP7_75t_L g1444 ( 
.A(n_972),
.Y(n_1444)
);

CKINVDCx5p33_ASAP7_75t_R g1445 ( 
.A(n_1028),
.Y(n_1445)
);

INVx1_ASAP7_75t_L g1446 ( 
.A(n_1018),
.Y(n_1446)
);

INVx3_ASAP7_75t_L g1447 ( 
.A(n_1174),
.Y(n_1447)
);

NAND2xp5_ASAP7_75t_L g1448 ( 
.A(n_1219),
.B(n_713),
.Y(n_1448)
);

NAND2xp5_ASAP7_75t_L g1449 ( 
.A(n_1309),
.B(n_714),
.Y(n_1449)
);

INVx5_ASAP7_75t_L g1450 ( 
.A(n_1312),
.Y(n_1450)
);

INVx5_ASAP7_75t_L g1451 ( 
.A(n_1326),
.Y(n_1451)
);

BUFx6f_ASAP7_75t_L g1452 ( 
.A(n_1326),
.Y(n_1452)
);

NOR2xp33_ASAP7_75t_L g1453 ( 
.A(n_964),
.B(n_578),
.Y(n_1453)
);

INVx1_ASAP7_75t_L g1454 ( 
.A(n_1019),
.Y(n_1454)
);

AND2x2_ASAP7_75t_L g1455 ( 
.A(n_1176),
.B(n_578),
.Y(n_1455)
);

INVx1_ASAP7_75t_L g1456 ( 
.A(n_1020),
.Y(n_1456)
);

CKINVDCx5p33_ASAP7_75t_R g1457 ( 
.A(n_1028),
.Y(n_1457)
);

NOR2xp33_ASAP7_75t_L g1458 ( 
.A(n_964),
.B(n_579),
.Y(n_1458)
);

BUFx3_ASAP7_75t_L g1459 ( 
.A(n_986),
.Y(n_1459)
);

BUFx6f_ASAP7_75t_L g1460 ( 
.A(n_1333),
.Y(n_1460)
);

AND2x4_ASAP7_75t_L g1461 ( 
.A(n_1284),
.B(n_579),
.Y(n_1461)
);

AND2x2_ASAP7_75t_L g1462 ( 
.A(n_1176),
.B(n_592),
.Y(n_1462)
);

NOR2xp33_ASAP7_75t_L g1463 ( 
.A(n_992),
.B(n_592),
.Y(n_1463)
);

BUFx6f_ASAP7_75t_L g1464 ( 
.A(n_1333),
.Y(n_1464)
);

INVxp67_ASAP7_75t_L g1465 ( 
.A(n_1071),
.Y(n_1465)
);

HB1xp67_ASAP7_75t_L g1466 ( 
.A(n_1082),
.Y(n_1466)
);

INVx1_ASAP7_75t_L g1467 ( 
.A(n_1021),
.Y(n_1467)
);

AND2x4_ASAP7_75t_L g1468 ( 
.A(n_1285),
.B(n_593),
.Y(n_1468)
);

AND2x4_ASAP7_75t_L g1469 ( 
.A(n_1286),
.B(n_593),
.Y(n_1469)
);

BUFx6f_ASAP7_75t_L g1470 ( 
.A(n_1025),
.Y(n_1470)
);

INVx1_ASAP7_75t_L g1471 ( 
.A(n_1026),
.Y(n_1471)
);

NAND2xp5_ASAP7_75t_L g1472 ( 
.A(n_1320),
.B(n_715),
.Y(n_1472)
);

AND2x2_ASAP7_75t_L g1473 ( 
.A(n_978),
.B(n_987),
.Y(n_1473)
);

NAND2xp5_ASAP7_75t_L g1474 ( 
.A(n_1268),
.B(n_727),
.Y(n_1474)
);

CKINVDCx5p33_ASAP7_75t_R g1475 ( 
.A(n_1045),
.Y(n_1475)
);

NAND2xp5_ASAP7_75t_SL g1476 ( 
.A(n_978),
.B(n_801),
.Y(n_1476)
);

BUFx6f_ASAP7_75t_L g1477 ( 
.A(n_1208),
.Y(n_1477)
);

BUFx6f_ASAP7_75t_L g1478 ( 
.A(n_1208),
.Y(n_1478)
);

INVx5_ASAP7_75t_L g1479 ( 
.A(n_1223),
.Y(n_1479)
);

INVx5_ASAP7_75t_L g1480 ( 
.A(n_1223),
.Y(n_1480)
);

AND2x4_ASAP7_75t_L g1481 ( 
.A(n_1287),
.B(n_598),
.Y(n_1481)
);

INVx2_ASAP7_75t_SL g1482 ( 
.A(n_1045),
.Y(n_1482)
);

HB1xp67_ASAP7_75t_L g1483 ( 
.A(n_1083),
.Y(n_1483)
);

NOR2xp33_ASAP7_75t_L g1484 ( 
.A(n_992),
.B(n_598),
.Y(n_1484)
);

INVx2_ASAP7_75t_L g1485 ( 
.A(n_962),
.Y(n_1485)
);

AND2x4_ASAP7_75t_L g1486 ( 
.A(n_1288),
.B(n_602),
.Y(n_1486)
);

INVxp67_ASAP7_75t_L g1487 ( 
.A(n_1127),
.Y(n_1487)
);

INVx4_ASAP7_75t_L g1488 ( 
.A(n_1048),
.Y(n_1488)
);

INVx1_ASAP7_75t_L g1489 ( 
.A(n_1165),
.Y(n_1489)
);

INVx2_ASAP7_75t_SL g1490 ( 
.A(n_1048),
.Y(n_1490)
);

BUFx6f_ASAP7_75t_L g1491 ( 
.A(n_1231),
.Y(n_1491)
);

BUFx6f_ASAP7_75t_L g1492 ( 
.A(n_1231),
.Y(n_1492)
);

HB1xp67_ASAP7_75t_L g1493 ( 
.A(n_1259),
.Y(n_1493)
);

INVx1_ASAP7_75t_L g1494 ( 
.A(n_1166),
.Y(n_1494)
);

AND2x2_ASAP7_75t_L g1495 ( 
.A(n_987),
.B(n_602),
.Y(n_1495)
);

NAND2xp5_ASAP7_75t_L g1496 ( 
.A(n_1268),
.B(n_730),
.Y(n_1496)
);

AND2x2_ASAP7_75t_L g1497 ( 
.A(n_1322),
.B(n_604),
.Y(n_1497)
);

INVx2_ASAP7_75t_SL g1498 ( 
.A(n_1059),
.Y(n_1498)
);

BUFx3_ASAP7_75t_L g1499 ( 
.A(n_988),
.Y(n_1499)
);

NAND2xp5_ASAP7_75t_L g1500 ( 
.A(n_1289),
.B(n_740),
.Y(n_1500)
);

AND2x2_ASAP7_75t_L g1501 ( 
.A(n_1059),
.B(n_604),
.Y(n_1501)
);

BUFx6f_ASAP7_75t_L g1502 ( 
.A(n_1232),
.Y(n_1502)
);

INVx2_ASAP7_75t_L g1503 ( 
.A(n_963),
.Y(n_1503)
);

BUFx12f_ASAP7_75t_L g1504 ( 
.A(n_1069),
.Y(n_1504)
);

AND2x2_ASAP7_75t_L g1505 ( 
.A(n_1069),
.B(n_616),
.Y(n_1505)
);

INVxp67_ASAP7_75t_L g1506 ( 
.A(n_1050),
.Y(n_1506)
);

INVx2_ASAP7_75t_L g1507 ( 
.A(n_966),
.Y(n_1507)
);

INVx5_ASAP7_75t_L g1508 ( 
.A(n_1232),
.Y(n_1508)
);

INVx1_ASAP7_75t_L g1509 ( 
.A(n_1167),
.Y(n_1509)
);

BUFx2_ASAP7_75t_L g1510 ( 
.A(n_1243),
.Y(n_1510)
);

CKINVDCx5p33_ASAP7_75t_R g1511 ( 
.A(n_1075),
.Y(n_1511)
);

BUFx12f_ASAP7_75t_L g1512 ( 
.A(n_1075),
.Y(n_1512)
);

NOR2xp33_ASAP7_75t_L g1513 ( 
.A(n_1052),
.B(n_1063),
.Y(n_1513)
);

BUFx6f_ASAP7_75t_L g1514 ( 
.A(n_1236),
.Y(n_1514)
);

HB1xp67_ASAP7_75t_L g1515 ( 
.A(n_1050),
.Y(n_1515)
);

NAND2xp5_ASAP7_75t_L g1516 ( 
.A(n_1289),
.B(n_741),
.Y(n_1516)
);

NAND2xp5_ASAP7_75t_L g1517 ( 
.A(n_1168),
.B(n_1169),
.Y(n_1517)
);

NOR2xp33_ASAP7_75t_L g1518 ( 
.A(n_1052),
.B(n_616),
.Y(n_1518)
);

INVx1_ASAP7_75t_L g1519 ( 
.A(n_1177),
.Y(n_1519)
);

NAND2xp5_ASAP7_75t_L g1520 ( 
.A(n_1178),
.B(n_750),
.Y(n_1520)
);

HB1xp67_ASAP7_75t_L g1521 ( 
.A(n_1330),
.Y(n_1521)
);

AND2x2_ASAP7_75t_L g1522 ( 
.A(n_1078),
.B(n_618),
.Y(n_1522)
);

BUFx6f_ASAP7_75t_L g1523 ( 
.A(n_1236),
.Y(n_1523)
);

INVx5_ASAP7_75t_L g1524 ( 
.A(n_1247),
.Y(n_1524)
);

BUFx12f_ASAP7_75t_L g1525 ( 
.A(n_1078),
.Y(n_1525)
);

INVx2_ASAP7_75t_L g1526 ( 
.A(n_967),
.Y(n_1526)
);

INVx1_ASAP7_75t_L g1527 ( 
.A(n_1179),
.Y(n_1527)
);

NOR2xp33_ASAP7_75t_L g1528 ( 
.A(n_1063),
.B(n_618),
.Y(n_1528)
);

BUFx3_ASAP7_75t_L g1529 ( 
.A(n_989),
.Y(n_1529)
);

NOR2xp33_ASAP7_75t_SL g1530 ( 
.A(n_1039),
.B(n_706),
.Y(n_1530)
);

NAND2xp5_ASAP7_75t_L g1531 ( 
.A(n_1180),
.B(n_775),
.Y(n_1531)
);

AND2x4_ASAP7_75t_L g1532 ( 
.A(n_1030),
.B(n_876),
.Y(n_1532)
);

AND2x4_ASAP7_75t_L g1533 ( 
.A(n_1037),
.B(n_876),
.Y(n_1533)
);

INVx1_ASAP7_75t_L g1534 ( 
.A(n_1182),
.Y(n_1534)
);

NOR2xp33_ASAP7_75t_SL g1535 ( 
.A(n_965),
.B(n_1064),
.Y(n_1535)
);

NAND2xp5_ASAP7_75t_L g1536 ( 
.A(n_1183),
.B(n_780),
.Y(n_1536)
);

BUFx3_ASAP7_75t_L g1537 ( 
.A(n_991),
.Y(n_1537)
);

INVx5_ASAP7_75t_L g1538 ( 
.A(n_1247),
.Y(n_1538)
);

AND2x4_ASAP7_75t_L g1539 ( 
.A(n_1037),
.B(n_892),
.Y(n_1539)
);

AND2x2_ASAP7_75t_L g1540 ( 
.A(n_1101),
.B(n_892),
.Y(n_1540)
);

BUFx6f_ASAP7_75t_L g1541 ( 
.A(n_1250),
.Y(n_1541)
);

BUFx6f_ASAP7_75t_L g1542 ( 
.A(n_1250),
.Y(n_1542)
);

BUFx6f_ASAP7_75t_L g1543 ( 
.A(n_1335),
.Y(n_1543)
);

INVx1_ASAP7_75t_L g1544 ( 
.A(n_1184),
.Y(n_1544)
);

AND2x4_ASAP7_75t_L g1545 ( 
.A(n_1062),
.B(n_1110),
.Y(n_1545)
);

BUFx6f_ASAP7_75t_L g1546 ( 
.A(n_1335),
.Y(n_1546)
);

INVx2_ASAP7_75t_SL g1547 ( 
.A(n_1101),
.Y(n_1547)
);

INVx5_ASAP7_75t_L g1548 ( 
.A(n_1031),
.Y(n_1548)
);

INVx1_ASAP7_75t_L g1549 ( 
.A(n_1185),
.Y(n_1549)
);

INVx1_ASAP7_75t_L g1550 ( 
.A(n_1187),
.Y(n_1550)
);

NAND2xp5_ASAP7_75t_L g1551 ( 
.A(n_1189),
.B(n_781),
.Y(n_1551)
);

BUFx6f_ASAP7_75t_L g1552 ( 
.A(n_968),
.Y(n_1552)
);

NAND2xp5_ASAP7_75t_SL g1553 ( 
.A(n_1062),
.B(n_1110),
.Y(n_1553)
);

BUFx2_ASAP7_75t_L g1554 ( 
.A(n_1295),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_1192),
.Y(n_1555)
);

NOR2xp33_ASAP7_75t_L g1556 ( 
.A(n_1088),
.B(n_896),
.Y(n_1556)
);

BUFx6f_ASAP7_75t_L g1557 ( 
.A(n_969),
.Y(n_1557)
);

INVx3_ASAP7_75t_L g1558 ( 
.A(n_1027),
.Y(n_1558)
);

BUFx12f_ASAP7_75t_L g1559 ( 
.A(n_1114),
.Y(n_1559)
);

AND2x6_ASAP7_75t_L g1560 ( 
.A(n_973),
.B(n_915),
.Y(n_1560)
);

BUFx12f_ASAP7_75t_L g1561 ( 
.A(n_1114),
.Y(n_1561)
);

NAND2xp5_ASAP7_75t_L g1562 ( 
.A(n_1193),
.B(n_785),
.Y(n_1562)
);

NOR2xp33_ASAP7_75t_SL g1563 ( 
.A(n_1115),
.B(n_779),
.Y(n_1563)
);

BUFx6f_ASAP7_75t_L g1564 ( 
.A(n_974),
.Y(n_1564)
);

BUFx2_ASAP7_75t_L g1565 ( 
.A(n_1295),
.Y(n_1565)
);

BUFx3_ASAP7_75t_L g1566 ( 
.A(n_995),
.Y(n_1566)
);

INVx2_ASAP7_75t_L g1567 ( 
.A(n_976),
.Y(n_1567)
);

INVx1_ASAP7_75t_L g1568 ( 
.A(n_1197),
.Y(n_1568)
);

BUFx8_ASAP7_75t_SL g1569 ( 
.A(n_985),
.Y(n_1569)
);

INVx1_ASAP7_75t_L g1570 ( 
.A(n_1198),
.Y(n_1570)
);

INVx2_ASAP7_75t_SL g1571 ( 
.A(n_1119),
.Y(n_1571)
);

NOR2xp33_ASAP7_75t_L g1572 ( 
.A(n_1088),
.B(n_1095),
.Y(n_1572)
);

INVx3_ASAP7_75t_L g1573 ( 
.A(n_1029),
.Y(n_1573)
);

NOR2xp33_ASAP7_75t_L g1574 ( 
.A(n_1095),
.B(n_896),
.Y(n_1574)
);

NAND2xp5_ASAP7_75t_L g1575 ( 
.A(n_1201),
.B(n_787),
.Y(n_1575)
);

INVx2_ASAP7_75t_L g1576 ( 
.A(n_977),
.Y(n_1576)
);

NOR2xp33_ASAP7_75t_L g1577 ( 
.A(n_1136),
.B(n_899),
.Y(n_1577)
);

AND2x2_ASAP7_75t_L g1578 ( 
.A(n_1119),
.B(n_899),
.Y(n_1578)
);

BUFx6f_ASAP7_75t_L g1579 ( 
.A(n_980),
.Y(n_1579)
);

BUFx12f_ASAP7_75t_L g1580 ( 
.A(n_1120),
.Y(n_1580)
);

INVx1_ASAP7_75t_L g1581 ( 
.A(n_1203),
.Y(n_1581)
);

BUFx12f_ASAP7_75t_L g1582 ( 
.A(n_1120),
.Y(n_1582)
);

BUFx12f_ASAP7_75t_L g1583 ( 
.A(n_1128),
.Y(n_1583)
);

INVx1_ASAP7_75t_L g1584 ( 
.A(n_1205),
.Y(n_1584)
);

BUFx6f_ASAP7_75t_L g1585 ( 
.A(n_981),
.Y(n_1585)
);

INVx1_ASAP7_75t_L g1586 ( 
.A(n_1206),
.Y(n_1586)
);

BUFx6f_ASAP7_75t_L g1587 ( 
.A(n_982),
.Y(n_1587)
);

AND2x4_ASAP7_75t_L g1588 ( 
.A(n_1218),
.B(n_902),
.Y(n_1588)
);

AND2x2_ASAP7_75t_L g1589 ( 
.A(n_1128),
.B(n_902),
.Y(n_1589)
);

INVx4_ASAP7_75t_L g1590 ( 
.A(n_1141),
.Y(n_1590)
);

NAND2xp5_ASAP7_75t_L g1591 ( 
.A(n_1207),
.B(n_798),
.Y(n_1591)
);

BUFx6f_ASAP7_75t_L g1592 ( 
.A(n_983),
.Y(n_1592)
);

AND2x4_ASAP7_75t_L g1593 ( 
.A(n_1218),
.B(n_924),
.Y(n_1593)
);

AND2x2_ASAP7_75t_L g1594 ( 
.A(n_1141),
.B(n_924),
.Y(n_1594)
);

INVx1_ASAP7_75t_L g1595 ( 
.A(n_1211),
.Y(n_1595)
);

INVx2_ASAP7_75t_L g1596 ( 
.A(n_1228),
.Y(n_1596)
);

INVx4_ASAP7_75t_L g1597 ( 
.A(n_1144),
.Y(n_1597)
);

NAND2xp5_ASAP7_75t_L g1598 ( 
.A(n_1213),
.B(n_799),
.Y(n_1598)
);

BUFx6f_ASAP7_75t_L g1599 ( 
.A(n_1049),
.Y(n_1599)
);

BUFx6f_ASAP7_75t_L g1600 ( 
.A(n_1049),
.Y(n_1600)
);

NOR2xp33_ASAP7_75t_L g1601 ( 
.A(n_1136),
.B(n_926),
.Y(n_1601)
);

AND2x2_ASAP7_75t_L g1602 ( 
.A(n_1144),
.B(n_926),
.Y(n_1602)
);

INVx2_ASAP7_75t_L g1603 ( 
.A(n_1230),
.Y(n_1603)
);

HB1xp67_ASAP7_75t_L g1604 ( 
.A(n_1330),
.Y(n_1604)
);

AND2x4_ASAP7_75t_L g1605 ( 
.A(n_1224),
.B(n_927),
.Y(n_1605)
);

INVxp67_ASAP7_75t_L g1606 ( 
.A(n_979),
.Y(n_1606)
);

BUFx6f_ASAP7_75t_L g1607 ( 
.A(n_1053),
.Y(n_1607)
);

BUFx8_ASAP7_75t_SL g1608 ( 
.A(n_985),
.Y(n_1608)
);

INVx1_ASAP7_75t_L g1609 ( 
.A(n_1214),
.Y(n_1609)
);

HB1xp67_ASAP7_75t_L g1610 ( 
.A(n_1148),
.Y(n_1610)
);

BUFx6f_ASAP7_75t_L g1611 ( 
.A(n_1053),
.Y(n_1611)
);

BUFx8_ASAP7_75t_SL g1612 ( 
.A(n_1017),
.Y(n_1612)
);

NAND2xp5_ASAP7_75t_L g1613 ( 
.A(n_1215),
.B(n_805),
.Y(n_1613)
);

NAND2xp5_ASAP7_75t_L g1614 ( 
.A(n_1216),
.B(n_808),
.Y(n_1614)
);

INVx2_ASAP7_75t_SL g1615 ( 
.A(n_1148),
.Y(n_1615)
);

NAND2xp5_ASAP7_75t_L g1616 ( 
.A(n_1217),
.B(n_1221),
.Y(n_1616)
);

AND2x4_ASAP7_75t_L g1617 ( 
.A(n_1224),
.B(n_927),
.Y(n_1617)
);

INVx3_ASAP7_75t_L g1618 ( 
.A(n_1032),
.Y(n_1618)
);

AND2x4_ASAP7_75t_L g1619 ( 
.A(n_990),
.B(n_928),
.Y(n_1619)
);

AND2x6_ASAP7_75t_L g1620 ( 
.A(n_1077),
.B(n_915),
.Y(n_1620)
);

CKINVDCx5p33_ASAP7_75t_R g1621 ( 
.A(n_1149),
.Y(n_1621)
);

BUFx8_ASAP7_75t_L g1622 ( 
.A(n_979),
.Y(n_1622)
);

BUFx6f_ASAP7_75t_L g1623 ( 
.A(n_1054),
.Y(n_1623)
);

NAND2xp5_ASAP7_75t_L g1624 ( 
.A(n_1222),
.B(n_831),
.Y(n_1624)
);

AND2x4_ASAP7_75t_L g1625 ( 
.A(n_993),
.B(n_928),
.Y(n_1625)
);

CKINVDCx6p67_ASAP7_75t_R g1626 ( 
.A(n_1133),
.Y(n_1626)
);

BUFx8_ASAP7_75t_SL g1627 ( 
.A(n_1017),
.Y(n_1627)
);

BUFx12f_ASAP7_75t_L g1628 ( 
.A(n_1149),
.Y(n_1628)
);

NAND2xp5_ASAP7_75t_L g1629 ( 
.A(n_1226),
.B(n_833),
.Y(n_1629)
);

NAND2xp5_ASAP7_75t_SL g1630 ( 
.A(n_1150),
.B(n_803),
.Y(n_1630)
);

NOR2xp33_ASAP7_75t_L g1631 ( 
.A(n_1146),
.B(n_930),
.Y(n_1631)
);

BUFx6f_ASAP7_75t_L g1632 ( 
.A(n_1054),
.Y(n_1632)
);

AND2x2_ASAP7_75t_L g1633 ( 
.A(n_1150),
.B(n_930),
.Y(n_1633)
);

INVx4_ASAP7_75t_L g1634 ( 
.A(n_1151),
.Y(n_1634)
);

BUFx3_ASAP7_75t_L g1635 ( 
.A(n_996),
.Y(n_1635)
);

NOR2xp33_ASAP7_75t_SL g1636 ( 
.A(n_1160),
.B(n_932),
.Y(n_1636)
);

BUFx2_ASAP7_75t_L g1637 ( 
.A(n_1310),
.Y(n_1637)
);

AND2x2_ASAP7_75t_L g1638 ( 
.A(n_1151),
.B(n_932),
.Y(n_1638)
);

NAND2xp5_ASAP7_75t_L g1639 ( 
.A(n_1227),
.B(n_836),
.Y(n_1639)
);

NOR2xp33_ASAP7_75t_L g1640 ( 
.A(n_1146),
.B(n_933),
.Y(n_1640)
);

BUFx2_ASAP7_75t_L g1641 ( 
.A(n_1310),
.Y(n_1641)
);

NOR2xp33_ASAP7_75t_L g1642 ( 
.A(n_1171),
.B(n_933),
.Y(n_1642)
);

INVx2_ASAP7_75t_SL g1643 ( 
.A(n_1159),
.Y(n_1643)
);

BUFx8_ASAP7_75t_SL g1644 ( 
.A(n_1041),
.Y(n_1644)
);

NOR2xp33_ASAP7_75t_L g1645 ( 
.A(n_1171),
.B(n_935),
.Y(n_1645)
);

INVx2_ASAP7_75t_L g1646 ( 
.A(n_1234),
.Y(n_1646)
);

CKINVDCx5p33_ASAP7_75t_R g1647 ( 
.A(n_1159),
.Y(n_1647)
);

NAND2xp33_ASAP7_75t_L g1648 ( 
.A(n_1099),
.B(n_915),
.Y(n_1648)
);

BUFx3_ASAP7_75t_L g1649 ( 
.A(n_1002),
.Y(n_1649)
);

HB1xp67_ASAP7_75t_L g1650 ( 
.A(n_1164),
.Y(n_1650)
);

INVx4_ASAP7_75t_L g1651 ( 
.A(n_1164),
.Y(n_1651)
);

INVx1_ASAP7_75t_L g1652 ( 
.A(n_1033),
.Y(n_1652)
);

AND2x4_ASAP7_75t_L g1653 ( 
.A(n_999),
.B(n_935),
.Y(n_1653)
);

AND2x6_ASAP7_75t_L g1654 ( 
.A(n_1104),
.B(n_915),
.Y(n_1654)
);

AND2x4_ASAP7_75t_L g1655 ( 
.A(n_1023),
.B(n_938),
.Y(n_1655)
);

NAND2xp5_ASAP7_75t_L g1656 ( 
.A(n_1006),
.B(n_839),
.Y(n_1656)
);

NOR2xp33_ASAP7_75t_L g1657 ( 
.A(n_1191),
.B(n_938),
.Y(n_1657)
);

AND2x4_ASAP7_75t_L g1658 ( 
.A(n_1007),
.B(n_941),
.Y(n_1658)
);

INVx1_ASAP7_75t_L g1659 ( 
.A(n_1413),
.Y(n_1659)
);

INVx6_ASAP7_75t_L g1660 ( 
.A(n_1364),
.Y(n_1660)
);

INVx1_ASAP7_75t_L g1661 ( 
.A(n_1413),
.Y(n_1661)
);

NAND2x1_ASAP7_75t_L g1662 ( 
.A(n_1620),
.B(n_915),
.Y(n_1662)
);

BUFx6f_ASAP7_75t_L g1663 ( 
.A(n_1346),
.Y(n_1663)
);

INVx1_ASAP7_75t_L g1664 ( 
.A(n_1652),
.Y(n_1664)
);

INVx1_ASAP7_75t_L g1665 ( 
.A(n_1489),
.Y(n_1665)
);

AND2x2_ASAP7_75t_L g1666 ( 
.A(n_1361),
.B(n_1170),
.Y(n_1666)
);

INVx1_ASAP7_75t_L g1667 ( 
.A(n_1494),
.Y(n_1667)
);

INVx1_ASAP7_75t_L g1668 ( 
.A(n_1509),
.Y(n_1668)
);

CKINVDCx8_ASAP7_75t_R g1669 ( 
.A(n_1367),
.Y(n_1669)
);

NAND2xp5_ASAP7_75t_L g1670 ( 
.A(n_1391),
.B(n_1170),
.Y(n_1670)
);

BUFx2_ASAP7_75t_L g1671 ( 
.A(n_1361),
.Y(n_1671)
);

BUFx6f_ASAP7_75t_L g1672 ( 
.A(n_1346),
.Y(n_1672)
);

AND2x2_ASAP7_75t_L g1673 ( 
.A(n_1422),
.B(n_1195),
.Y(n_1673)
);

INVx1_ASAP7_75t_L g1674 ( 
.A(n_1519),
.Y(n_1674)
);

BUFx2_ASAP7_75t_L g1675 ( 
.A(n_1622),
.Y(n_1675)
);

HB1xp67_ASAP7_75t_L g1676 ( 
.A(n_1427),
.Y(n_1676)
);

INVx2_ASAP7_75t_L g1677 ( 
.A(n_1362),
.Y(n_1677)
);

INVx1_ASAP7_75t_L g1678 ( 
.A(n_1527),
.Y(n_1678)
);

INVx2_ASAP7_75t_L g1679 ( 
.A(n_1362),
.Y(n_1679)
);

BUFx6f_ASAP7_75t_L g1680 ( 
.A(n_1346),
.Y(n_1680)
);

INVx3_ASAP7_75t_L g1681 ( 
.A(n_1346),
.Y(n_1681)
);

BUFx6f_ASAP7_75t_L g1682 ( 
.A(n_1353),
.Y(n_1682)
);

BUFx6f_ASAP7_75t_L g1683 ( 
.A(n_1353),
.Y(n_1683)
);

AND3x2_ASAP7_75t_L g1684 ( 
.A(n_1636),
.B(n_1204),
.C(n_1202),
.Y(n_1684)
);

INVx2_ASAP7_75t_L g1685 ( 
.A(n_1371),
.Y(n_1685)
);

BUFx8_ASAP7_75t_L g1686 ( 
.A(n_1510),
.Y(n_1686)
);

BUFx2_ASAP7_75t_L g1687 ( 
.A(n_1622),
.Y(n_1687)
);

INVx3_ASAP7_75t_L g1688 ( 
.A(n_1353),
.Y(n_1688)
);

INVx3_ASAP7_75t_L g1689 ( 
.A(n_1353),
.Y(n_1689)
);

OA21x2_ASAP7_75t_L g1690 ( 
.A1(n_1485),
.A2(n_1240),
.B(n_1237),
.Y(n_1690)
);

BUFx6f_ASAP7_75t_L g1691 ( 
.A(n_1368),
.Y(n_1691)
);

NAND2xp5_ASAP7_75t_L g1692 ( 
.A(n_1391),
.B(n_1195),
.Y(n_1692)
);

INVx2_ASAP7_75t_L g1693 ( 
.A(n_1371),
.Y(n_1693)
);

AND2x4_ASAP7_75t_L g1694 ( 
.A(n_1358),
.B(n_1265),
.Y(n_1694)
);

INVx1_ASAP7_75t_L g1695 ( 
.A(n_1534),
.Y(n_1695)
);

INVx2_ASAP7_75t_L g1696 ( 
.A(n_1373),
.Y(n_1696)
);

INVx2_ASAP7_75t_L g1697 ( 
.A(n_1373),
.Y(n_1697)
);

BUFx6f_ASAP7_75t_L g1698 ( 
.A(n_1368),
.Y(n_1698)
);

BUFx6f_ASAP7_75t_L g1699 ( 
.A(n_1368),
.Y(n_1699)
);

AND2x6_ASAP7_75t_L g1700 ( 
.A(n_1351),
.B(n_1124),
.Y(n_1700)
);

INVx1_ASAP7_75t_L g1701 ( 
.A(n_1544),
.Y(n_1701)
);

INVx1_ASAP7_75t_L g1702 ( 
.A(n_1549),
.Y(n_1702)
);

BUFx6f_ASAP7_75t_L g1703 ( 
.A(n_1368),
.Y(n_1703)
);

INVx1_ASAP7_75t_L g1704 ( 
.A(n_1550),
.Y(n_1704)
);

INVx2_ASAP7_75t_L g1705 ( 
.A(n_1378),
.Y(n_1705)
);

BUFx8_ASAP7_75t_L g1706 ( 
.A(n_1554),
.Y(n_1706)
);

NAND2xp5_ASAP7_75t_L g1707 ( 
.A(n_1349),
.B(n_1199),
.Y(n_1707)
);

INVx1_ASAP7_75t_L g1708 ( 
.A(n_1555),
.Y(n_1708)
);

BUFx6f_ASAP7_75t_L g1709 ( 
.A(n_1374),
.Y(n_1709)
);

AOI22xp5_ASAP7_75t_L g1710 ( 
.A1(n_1417),
.A2(n_1254),
.B1(n_1256),
.B2(n_1199),
.Y(n_1710)
);

INVx1_ASAP7_75t_L g1711 ( 
.A(n_1568),
.Y(n_1711)
);

INVx2_ASAP7_75t_L g1712 ( 
.A(n_1378),
.Y(n_1712)
);

INVx3_ASAP7_75t_L g1713 ( 
.A(n_1374),
.Y(n_1713)
);

INVxp67_ASAP7_75t_L g1714 ( 
.A(n_1453),
.Y(n_1714)
);

INVx1_ASAP7_75t_L g1715 ( 
.A(n_1570),
.Y(n_1715)
);

INVx1_ASAP7_75t_L g1716 ( 
.A(n_1581),
.Y(n_1716)
);

INVx2_ASAP7_75t_L g1717 ( 
.A(n_1379),
.Y(n_1717)
);

INVx3_ASAP7_75t_L g1718 ( 
.A(n_1374),
.Y(n_1718)
);

AND2x2_ASAP7_75t_L g1719 ( 
.A(n_1455),
.B(n_1266),
.Y(n_1719)
);

AND2x4_ASAP7_75t_L g1720 ( 
.A(n_1358),
.B(n_1267),
.Y(n_1720)
);

BUFx6f_ASAP7_75t_L g1721 ( 
.A(n_1374),
.Y(n_1721)
);

INVx3_ASAP7_75t_L g1722 ( 
.A(n_1376),
.Y(n_1722)
);

NAND2xp5_ASAP7_75t_L g1723 ( 
.A(n_1349),
.B(n_1357),
.Y(n_1723)
);

INVx1_ASAP7_75t_L g1724 ( 
.A(n_1584),
.Y(n_1724)
);

NAND2xp5_ASAP7_75t_L g1725 ( 
.A(n_1355),
.B(n_1254),
.Y(n_1725)
);

INVx2_ASAP7_75t_L g1726 ( 
.A(n_1379),
.Y(n_1726)
);

INVx1_ASAP7_75t_L g1727 ( 
.A(n_1586),
.Y(n_1727)
);

INVx1_ASAP7_75t_L g1728 ( 
.A(n_1595),
.Y(n_1728)
);

INVx3_ASAP7_75t_L g1729 ( 
.A(n_1376),
.Y(n_1729)
);

AND2x4_ASAP7_75t_L g1730 ( 
.A(n_1396),
.B(n_1269),
.Y(n_1730)
);

AND2x2_ASAP7_75t_L g1731 ( 
.A(n_1462),
.B(n_1256),
.Y(n_1731)
);

INVx1_ASAP7_75t_L g1732 ( 
.A(n_1609),
.Y(n_1732)
);

INVx1_ASAP7_75t_L g1733 ( 
.A(n_1485),
.Y(n_1733)
);

AND2x2_ASAP7_75t_L g1734 ( 
.A(n_1545),
.B(n_1260),
.Y(n_1734)
);

AND2x4_ASAP7_75t_L g1735 ( 
.A(n_1396),
.B(n_1270),
.Y(n_1735)
);

AND2x4_ASAP7_75t_L g1736 ( 
.A(n_1400),
.B(n_1271),
.Y(n_1736)
);

INVx2_ASAP7_75t_L g1737 ( 
.A(n_1414),
.Y(n_1737)
);

INVx1_ASAP7_75t_L g1738 ( 
.A(n_1503),
.Y(n_1738)
);

INVx1_ASAP7_75t_L g1739 ( 
.A(n_1503),
.Y(n_1739)
);

INVx1_ASAP7_75t_L g1740 ( 
.A(n_1507),
.Y(n_1740)
);

NAND2xp5_ASAP7_75t_L g1741 ( 
.A(n_1341),
.B(n_1260),
.Y(n_1741)
);

BUFx6f_ASAP7_75t_L g1742 ( 
.A(n_1376),
.Y(n_1742)
);

INVx3_ASAP7_75t_L g1743 ( 
.A(n_1376),
.Y(n_1743)
);

INVx2_ASAP7_75t_L g1744 ( 
.A(n_1414),
.Y(n_1744)
);

INVx2_ASAP7_75t_L g1745 ( 
.A(n_1441),
.Y(n_1745)
);

NAND2xp5_ASAP7_75t_SL g1746 ( 
.A(n_1545),
.B(n_1263),
.Y(n_1746)
);

OA21x2_ASAP7_75t_L g1747 ( 
.A1(n_1507),
.A2(n_1244),
.B(n_1242),
.Y(n_1747)
);

AND2x2_ASAP7_75t_L g1748 ( 
.A(n_1344),
.B(n_1263),
.Y(n_1748)
);

AND2x4_ASAP7_75t_L g1749 ( 
.A(n_1400),
.B(n_1272),
.Y(n_1749)
);

BUFx6f_ASAP7_75t_L g1750 ( 
.A(n_1377),
.Y(n_1750)
);

INVx2_ASAP7_75t_L g1751 ( 
.A(n_1441),
.Y(n_1751)
);

INVx1_ASAP7_75t_L g1752 ( 
.A(n_1526),
.Y(n_1752)
);

INVxp67_ASAP7_75t_L g1753 ( 
.A(n_1453),
.Y(n_1753)
);

INVx1_ASAP7_75t_L g1754 ( 
.A(n_1526),
.Y(n_1754)
);

INVx1_ASAP7_75t_L g1755 ( 
.A(n_1567),
.Y(n_1755)
);

INVx1_ASAP7_75t_L g1756 ( 
.A(n_1567),
.Y(n_1756)
);

INVx4_ASAP7_75t_L g1757 ( 
.A(n_1548),
.Y(n_1757)
);

INVx1_ASAP7_75t_L g1758 ( 
.A(n_1576),
.Y(n_1758)
);

NOR2xp33_ASAP7_75t_L g1759 ( 
.A(n_1380),
.B(n_1191),
.Y(n_1759)
);

NOR2xp33_ASAP7_75t_SL g1760 ( 
.A(n_1340),
.B(n_1324),
.Y(n_1760)
);

INVx1_ASAP7_75t_L g1761 ( 
.A(n_1576),
.Y(n_1761)
);

INVx1_ASAP7_75t_L g1762 ( 
.A(n_1552),
.Y(n_1762)
);

INVx1_ASAP7_75t_L g1763 ( 
.A(n_1552),
.Y(n_1763)
);

INVx1_ASAP7_75t_L g1764 ( 
.A(n_1552),
.Y(n_1764)
);

INVxp67_ASAP7_75t_L g1765 ( 
.A(n_1458),
.Y(n_1765)
);

INVx3_ASAP7_75t_L g1766 ( 
.A(n_1377),
.Y(n_1766)
);

NAND2xp5_ASAP7_75t_L g1767 ( 
.A(n_1342),
.B(n_1280),
.Y(n_1767)
);

INVx4_ASAP7_75t_L g1768 ( 
.A(n_1548),
.Y(n_1768)
);

INVx1_ASAP7_75t_L g1769 ( 
.A(n_1552),
.Y(n_1769)
);

NAND2xp5_ASAP7_75t_SL g1770 ( 
.A(n_1348),
.B(n_1280),
.Y(n_1770)
);

CKINVDCx8_ASAP7_75t_R g1771 ( 
.A(n_1565),
.Y(n_1771)
);

BUFx6f_ASAP7_75t_L g1772 ( 
.A(n_1377),
.Y(n_1772)
);

AND2x2_ASAP7_75t_L g1773 ( 
.A(n_1347),
.B(n_1313),
.Y(n_1773)
);

OAI22xp5_ASAP7_75t_SL g1774 ( 
.A1(n_1513),
.A2(n_1336),
.B1(n_1329),
.B2(n_1046),
.Y(n_1774)
);

AND2x2_ASAP7_75t_L g1775 ( 
.A(n_1370),
.B(n_1313),
.Y(n_1775)
);

NAND2xp5_ASAP7_75t_L g1776 ( 
.A(n_1474),
.B(n_1317),
.Y(n_1776)
);

BUFx8_ASAP7_75t_L g1777 ( 
.A(n_1637),
.Y(n_1777)
);

HB1xp67_ASAP7_75t_L g1778 ( 
.A(n_1515),
.Y(n_1778)
);

INVx1_ASAP7_75t_L g1779 ( 
.A(n_1557),
.Y(n_1779)
);

BUFx6f_ASAP7_75t_L g1780 ( 
.A(n_1377),
.Y(n_1780)
);

NOR2x1_ASAP7_75t_L g1781 ( 
.A(n_1340),
.B(n_1273),
.Y(n_1781)
);

INVx2_ASAP7_75t_L g1782 ( 
.A(n_1419),
.Y(n_1782)
);

NAND2xp5_ASAP7_75t_SL g1783 ( 
.A(n_1348),
.B(n_1317),
.Y(n_1783)
);

BUFx6f_ASAP7_75t_L g1784 ( 
.A(n_1385),
.Y(n_1784)
);

INVx1_ASAP7_75t_L g1785 ( 
.A(n_1557),
.Y(n_1785)
);

NAND2xp5_ASAP7_75t_L g1786 ( 
.A(n_1496),
.B(n_1321),
.Y(n_1786)
);

BUFx6f_ASAP7_75t_L g1787 ( 
.A(n_1385),
.Y(n_1787)
);

AND2x2_ASAP7_75t_L g1788 ( 
.A(n_1436),
.B(n_1274),
.Y(n_1788)
);

INVx2_ASAP7_75t_L g1789 ( 
.A(n_1419),
.Y(n_1789)
);

NAND2xp5_ASAP7_75t_L g1790 ( 
.A(n_1500),
.B(n_1321),
.Y(n_1790)
);

NAND2xp5_ASAP7_75t_SL g1791 ( 
.A(n_1365),
.B(n_844),
.Y(n_1791)
);

INVx1_ASAP7_75t_L g1792 ( 
.A(n_1557),
.Y(n_1792)
);

INVx2_ASAP7_75t_L g1793 ( 
.A(n_1439),
.Y(n_1793)
);

BUFx6f_ASAP7_75t_L g1794 ( 
.A(n_1385),
.Y(n_1794)
);

XOR2xp5_ASAP7_75t_L g1795 ( 
.A(n_1445),
.B(n_1338),
.Y(n_1795)
);

INVx2_ASAP7_75t_L g1796 ( 
.A(n_1439),
.Y(n_1796)
);

INVx2_ASAP7_75t_L g1797 ( 
.A(n_1477),
.Y(n_1797)
);

BUFx6f_ASAP7_75t_L g1798 ( 
.A(n_1385),
.Y(n_1798)
);

INVx1_ASAP7_75t_L g1799 ( 
.A(n_1557),
.Y(n_1799)
);

NOR2xp33_ASAP7_75t_L g1800 ( 
.A(n_1389),
.B(n_1196),
.Y(n_1800)
);

INVx1_ASAP7_75t_L g1801 ( 
.A(n_1564),
.Y(n_1801)
);

INVx1_ASAP7_75t_L g1802 ( 
.A(n_1564),
.Y(n_1802)
);

NAND2xp5_ASAP7_75t_L g1803 ( 
.A(n_1516),
.B(n_1246),
.Y(n_1803)
);

AND2x2_ASAP7_75t_L g1804 ( 
.A(n_1372),
.B(n_960),
.Y(n_1804)
);

INVx1_ASAP7_75t_L g1805 ( 
.A(n_1564),
.Y(n_1805)
);

INVx2_ASAP7_75t_L g1806 ( 
.A(n_1477),
.Y(n_1806)
);

NAND2xp5_ASAP7_75t_L g1807 ( 
.A(n_1411),
.B(n_1252),
.Y(n_1807)
);

INVx1_ASAP7_75t_L g1808 ( 
.A(n_1564),
.Y(n_1808)
);

AND2x2_ASAP7_75t_L g1809 ( 
.A(n_1410),
.B(n_960),
.Y(n_1809)
);

BUFx2_ASAP7_75t_L g1810 ( 
.A(n_1386),
.Y(n_1810)
);

INVx1_ASAP7_75t_L g1811 ( 
.A(n_1579),
.Y(n_1811)
);

NAND2xp33_ASAP7_75t_L g1812 ( 
.A(n_1354),
.B(n_1099),
.Y(n_1812)
);

CKINVDCx20_ASAP7_75t_R g1813 ( 
.A(n_1569),
.Y(n_1813)
);

INVx1_ASAP7_75t_L g1814 ( 
.A(n_1579),
.Y(n_1814)
);

AND2x4_ASAP7_75t_L g1815 ( 
.A(n_1403),
.B(n_1275),
.Y(n_1815)
);

INVx1_ASAP7_75t_L g1816 ( 
.A(n_1579),
.Y(n_1816)
);

INVx2_ASAP7_75t_L g1817 ( 
.A(n_1477),
.Y(n_1817)
);

INVx1_ASAP7_75t_L g1818 ( 
.A(n_1579),
.Y(n_1818)
);

BUFx6f_ASAP7_75t_L g1819 ( 
.A(n_1394),
.Y(n_1819)
);

AND2x2_ASAP7_75t_L g1820 ( 
.A(n_1415),
.B(n_1173),
.Y(n_1820)
);

HB1xp67_ASAP7_75t_L g1821 ( 
.A(n_1515),
.Y(n_1821)
);

INVx1_ASAP7_75t_L g1822 ( 
.A(n_1585),
.Y(n_1822)
);

NAND2xp5_ASAP7_75t_SL g1823 ( 
.A(n_1365),
.B(n_856),
.Y(n_1823)
);

BUFx6f_ASAP7_75t_L g1824 ( 
.A(n_1394),
.Y(n_1824)
);

BUFx3_ASAP7_75t_L g1825 ( 
.A(n_1403),
.Y(n_1825)
);

OA21x2_ASAP7_75t_L g1826 ( 
.A1(n_1356),
.A2(n_1126),
.B(n_1124),
.Y(n_1826)
);

HB1xp67_ASAP7_75t_L g1827 ( 
.A(n_1521),
.Y(n_1827)
);

INVx3_ASAP7_75t_L g1828 ( 
.A(n_1394),
.Y(n_1828)
);

BUFx2_ASAP7_75t_L g1829 ( 
.A(n_1386),
.Y(n_1829)
);

AND2x4_ASAP7_75t_L g1830 ( 
.A(n_1406),
.B(n_1276),
.Y(n_1830)
);

INVx1_ASAP7_75t_L g1831 ( 
.A(n_1585),
.Y(n_1831)
);

NOR2xp33_ASAP7_75t_L g1832 ( 
.A(n_1359),
.B(n_1196),
.Y(n_1832)
);

INVx3_ASAP7_75t_L g1833 ( 
.A(n_1394),
.Y(n_1833)
);

INVx1_ASAP7_75t_L g1834 ( 
.A(n_1585),
.Y(n_1834)
);

INVx3_ASAP7_75t_L g1835 ( 
.A(n_1401),
.Y(n_1835)
);

BUFx6f_ASAP7_75t_L g1836 ( 
.A(n_1401),
.Y(n_1836)
);

NAND2xp5_ASAP7_75t_L g1837 ( 
.A(n_1429),
.B(n_1277),
.Y(n_1837)
);

INVx3_ASAP7_75t_L g1838 ( 
.A(n_1401),
.Y(n_1838)
);

INVxp67_ASAP7_75t_L g1839 ( 
.A(n_1458),
.Y(n_1839)
);

NAND2xp5_ASAP7_75t_L g1840 ( 
.A(n_1438),
.B(n_858),
.Y(n_1840)
);

INVx3_ASAP7_75t_L g1841 ( 
.A(n_1401),
.Y(n_1841)
);

AOI22xp5_ASAP7_75t_L g1842 ( 
.A1(n_1417),
.A2(n_1200),
.B1(n_1282),
.B2(n_1209),
.Y(n_1842)
);

AND2x4_ASAP7_75t_L g1843 ( 
.A(n_1406),
.B(n_1034),
.Y(n_1843)
);

INVx1_ASAP7_75t_L g1844 ( 
.A(n_1585),
.Y(n_1844)
);

AND2x6_ASAP7_75t_L g1845 ( 
.A(n_1387),
.B(n_1126),
.Y(n_1845)
);

INVx2_ASAP7_75t_L g1846 ( 
.A(n_1477),
.Y(n_1846)
);

BUFx8_ASAP7_75t_L g1847 ( 
.A(n_1641),
.Y(n_1847)
);

INVx1_ASAP7_75t_L g1848 ( 
.A(n_1587),
.Y(n_1848)
);

NOR2xp33_ASAP7_75t_L g1849 ( 
.A(n_1363),
.B(n_1369),
.Y(n_1849)
);

OA21x2_ASAP7_75t_L g1850 ( 
.A1(n_1375),
.A2(n_1155),
.B(n_1137),
.Y(n_1850)
);

AND2x2_ASAP7_75t_L g1851 ( 
.A(n_1415),
.B(n_1225),
.Y(n_1851)
);

INVx1_ASAP7_75t_L g1852 ( 
.A(n_1587),
.Y(n_1852)
);

CKINVDCx5p33_ASAP7_75t_R g1853 ( 
.A(n_1569),
.Y(n_1853)
);

INVx1_ASAP7_75t_L g1854 ( 
.A(n_1587),
.Y(n_1854)
);

INVx1_ASAP7_75t_L g1855 ( 
.A(n_1587),
.Y(n_1855)
);

NOR2xp33_ASAP7_75t_L g1856 ( 
.A(n_1382),
.B(n_1200),
.Y(n_1856)
);

NAND2xp5_ASAP7_75t_L g1857 ( 
.A(n_1448),
.B(n_862),
.Y(n_1857)
);

OAI22xp5_ASAP7_75t_L g1858 ( 
.A1(n_1506),
.A2(n_1282),
.B1(n_1209),
.B2(n_807),
.Y(n_1858)
);

BUFx6f_ASAP7_75t_L g1859 ( 
.A(n_1407),
.Y(n_1859)
);

BUFx6f_ASAP7_75t_L g1860 ( 
.A(n_1407),
.Y(n_1860)
);

INVx1_ASAP7_75t_L g1861 ( 
.A(n_1592),
.Y(n_1861)
);

INVx2_ASAP7_75t_L g1862 ( 
.A(n_1478),
.Y(n_1862)
);

BUFx6f_ASAP7_75t_L g1863 ( 
.A(n_1407),
.Y(n_1863)
);

AND2x2_ASAP7_75t_L g1864 ( 
.A(n_1532),
.B(n_1233),
.Y(n_1864)
);

NAND2xp5_ASAP7_75t_L g1865 ( 
.A(n_1383),
.B(n_868),
.Y(n_1865)
);

OA21x2_ASAP7_75t_L g1866 ( 
.A1(n_1388),
.A2(n_1446),
.B(n_1404),
.Y(n_1866)
);

INVx1_ASAP7_75t_L g1867 ( 
.A(n_1592),
.Y(n_1867)
);

AND2x2_ASAP7_75t_L g1868 ( 
.A(n_1436),
.B(n_1008),
.Y(n_1868)
);

INVx1_ASAP7_75t_L g1869 ( 
.A(n_1592),
.Y(n_1869)
);

BUFx6f_ASAP7_75t_L g1870 ( 
.A(n_1407),
.Y(n_1870)
);

INVxp67_ASAP7_75t_L g1871 ( 
.A(n_1463),
.Y(n_1871)
);

INVx1_ASAP7_75t_L g1872 ( 
.A(n_1592),
.Y(n_1872)
);

INVx1_ASAP7_75t_L g1873 ( 
.A(n_1428),
.Y(n_1873)
);

INVx1_ASAP7_75t_L g1874 ( 
.A(n_1428),
.Y(n_1874)
);

AND2x2_ASAP7_75t_L g1875 ( 
.A(n_1596),
.B(n_1009),
.Y(n_1875)
);

INVx3_ASAP7_75t_L g1876 ( 
.A(n_1409),
.Y(n_1876)
);

INVx2_ASAP7_75t_L g1877 ( 
.A(n_1478),
.Y(n_1877)
);

INVx2_ASAP7_75t_L g1878 ( 
.A(n_1478),
.Y(n_1878)
);

NAND2xp5_ASAP7_75t_L g1879 ( 
.A(n_1520),
.B(n_869),
.Y(n_1879)
);

AND2x4_ASAP7_75t_L g1880 ( 
.A(n_1408),
.B(n_1035),
.Y(n_1880)
);

INVx1_ASAP7_75t_L g1881 ( 
.A(n_1459),
.Y(n_1881)
);

INVx2_ASAP7_75t_L g1882 ( 
.A(n_1478),
.Y(n_1882)
);

INVx1_ASAP7_75t_L g1883 ( 
.A(n_1459),
.Y(n_1883)
);

NAND2xp5_ASAP7_75t_L g1884 ( 
.A(n_1531),
.B(n_871),
.Y(n_1884)
);

AND2x2_ASAP7_75t_L g1885 ( 
.A(n_1532),
.B(n_1239),
.Y(n_1885)
);

INVx1_ASAP7_75t_L g1886 ( 
.A(n_1499),
.Y(n_1886)
);

INVx2_ASAP7_75t_L g1887 ( 
.A(n_1491),
.Y(n_1887)
);

NAND2xp5_ASAP7_75t_L g1888 ( 
.A(n_1536),
.B(n_941),
.Y(n_1888)
);

INVx1_ASAP7_75t_L g1889 ( 
.A(n_1499),
.Y(n_1889)
);

HB1xp67_ASAP7_75t_L g1890 ( 
.A(n_1521),
.Y(n_1890)
);

NAND2xp5_ASAP7_75t_L g1891 ( 
.A(n_1551),
.B(n_1137),
.Y(n_1891)
);

NAND2xp33_ASAP7_75t_SL g1892 ( 
.A(n_1553),
.B(n_590),
.Y(n_1892)
);

INVx1_ASAP7_75t_L g1893 ( 
.A(n_1529),
.Y(n_1893)
);

NAND2xp5_ASAP7_75t_L g1894 ( 
.A(n_1562),
.B(n_1155),
.Y(n_1894)
);

INVx2_ASAP7_75t_L g1895 ( 
.A(n_1491),
.Y(n_1895)
);

INVx2_ASAP7_75t_L g1896 ( 
.A(n_1491),
.Y(n_1896)
);

AND2x4_ASAP7_75t_L g1897 ( 
.A(n_1408),
.B(n_1036),
.Y(n_1897)
);

BUFx6f_ASAP7_75t_L g1898 ( 
.A(n_1409),
.Y(n_1898)
);

INVx2_ASAP7_75t_L g1899 ( 
.A(n_1491),
.Y(n_1899)
);

INVx2_ASAP7_75t_L g1900 ( 
.A(n_1492),
.Y(n_1900)
);

AOI22xp5_ASAP7_75t_L g1901 ( 
.A1(n_1630),
.A2(n_1336),
.B1(n_1329),
.B2(n_1212),
.Y(n_1901)
);

OA21x2_ASAP7_75t_L g1902 ( 
.A1(n_1454),
.A2(n_1194),
.B(n_1253),
.Y(n_1902)
);

INVx2_ASAP7_75t_L g1903 ( 
.A(n_1492),
.Y(n_1903)
);

INVx1_ASAP7_75t_L g1904 ( 
.A(n_1529),
.Y(n_1904)
);

AND2x6_ASAP7_75t_L g1905 ( 
.A(n_1398),
.B(n_1038),
.Y(n_1905)
);

HB1xp67_ASAP7_75t_L g1906 ( 
.A(n_1604),
.Y(n_1906)
);

AND2x2_ASAP7_75t_L g1907 ( 
.A(n_1533),
.B(n_1220),
.Y(n_1907)
);

INVx1_ASAP7_75t_L g1908 ( 
.A(n_1537),
.Y(n_1908)
);

INVx3_ASAP7_75t_L g1909 ( 
.A(n_1409),
.Y(n_1909)
);

BUFx3_ASAP7_75t_L g1910 ( 
.A(n_1537),
.Y(n_1910)
);

AND2x2_ASAP7_75t_L g1911 ( 
.A(n_1533),
.B(n_1251),
.Y(n_1911)
);

AND2x2_ASAP7_75t_L g1912 ( 
.A(n_1539),
.B(n_1186),
.Y(n_1912)
);

INVx1_ASAP7_75t_L g1913 ( 
.A(n_1566),
.Y(n_1913)
);

OAI21x1_ASAP7_75t_L g1914 ( 
.A1(n_1656),
.A2(n_1194),
.B(n_1255),
.Y(n_1914)
);

INVx1_ASAP7_75t_L g1915 ( 
.A(n_1566),
.Y(n_1915)
);

NAND2xp5_ASAP7_75t_L g1916 ( 
.A(n_1575),
.B(n_1257),
.Y(n_1916)
);

INVx1_ASAP7_75t_L g1917 ( 
.A(n_1635),
.Y(n_1917)
);

INVx1_ASAP7_75t_L g1918 ( 
.A(n_1635),
.Y(n_1918)
);

INVx1_ASAP7_75t_L g1919 ( 
.A(n_1649),
.Y(n_1919)
);

INVx1_ASAP7_75t_L g1920 ( 
.A(n_1649),
.Y(n_1920)
);

INVx1_ASAP7_75t_L g1921 ( 
.A(n_1352),
.Y(n_1921)
);

NAND2xp5_ASAP7_75t_SL g1922 ( 
.A(n_1366),
.B(n_804),
.Y(n_1922)
);

INVx1_ASAP7_75t_L g1923 ( 
.A(n_1352),
.Y(n_1923)
);

HB1xp67_ASAP7_75t_L g1924 ( 
.A(n_1604),
.Y(n_1924)
);

BUFx6f_ASAP7_75t_L g1925 ( 
.A(n_1409),
.Y(n_1925)
);

INVx6_ASAP7_75t_L g1926 ( 
.A(n_1364),
.Y(n_1926)
);

AND2x2_ASAP7_75t_L g1927 ( 
.A(n_1596),
.B(n_1258),
.Y(n_1927)
);

HB1xp67_ASAP7_75t_L g1928 ( 
.A(n_1431),
.Y(n_1928)
);

NOR2xp33_ASAP7_75t_SL g1929 ( 
.A(n_1397),
.B(n_562),
.Y(n_1929)
);

NAND2xp5_ASAP7_75t_L g1930 ( 
.A(n_1591),
.B(n_1261),
.Y(n_1930)
);

NAND2xp5_ASAP7_75t_L g1931 ( 
.A(n_1598),
.B(n_1264),
.Y(n_1931)
);

NAND2xp5_ASAP7_75t_SL g1932 ( 
.A(n_1366),
.B(n_810),
.Y(n_1932)
);

INVx1_ASAP7_75t_L g1933 ( 
.A(n_1456),
.Y(n_1933)
);

NAND2xp5_ASAP7_75t_L g1934 ( 
.A(n_1613),
.B(n_1040),
.Y(n_1934)
);

BUFx6f_ASAP7_75t_L g1935 ( 
.A(n_1418),
.Y(n_1935)
);

INVx2_ASAP7_75t_L g1936 ( 
.A(n_1492),
.Y(n_1936)
);

BUFx6f_ASAP7_75t_L g1937 ( 
.A(n_1418),
.Y(n_1937)
);

INVx2_ASAP7_75t_L g1938 ( 
.A(n_1492),
.Y(n_1938)
);

NAND2xp5_ASAP7_75t_L g1939 ( 
.A(n_1614),
.B(n_1043),
.Y(n_1939)
);

AND2x4_ASAP7_75t_L g1940 ( 
.A(n_1558),
.B(n_1044),
.Y(n_1940)
);

BUFx6f_ASAP7_75t_L g1941 ( 
.A(n_1418),
.Y(n_1941)
);

BUFx2_ASAP7_75t_L g1942 ( 
.A(n_1431),
.Y(n_1942)
);

NAND2xp5_ASAP7_75t_L g1943 ( 
.A(n_1624),
.B(n_1047),
.Y(n_1943)
);

INVx2_ASAP7_75t_L g1944 ( 
.A(n_1502),
.Y(n_1944)
);

INVx1_ASAP7_75t_L g1945 ( 
.A(n_1467),
.Y(n_1945)
);

NAND2xp5_ASAP7_75t_L g1946 ( 
.A(n_1629),
.B(n_1058),
.Y(n_1946)
);

INVx1_ASAP7_75t_L g1947 ( 
.A(n_1471),
.Y(n_1947)
);

INVx2_ASAP7_75t_L g1948 ( 
.A(n_1502),
.Y(n_1948)
);

AND2x2_ASAP7_75t_L g1949 ( 
.A(n_1539),
.B(n_1296),
.Y(n_1949)
);

AND3x2_ASAP7_75t_L g1950 ( 
.A(n_1343),
.B(n_1298),
.C(n_1297),
.Y(n_1950)
);

INVx1_ASAP7_75t_L g1951 ( 
.A(n_1558),
.Y(n_1951)
);

INVx1_ASAP7_75t_L g1952 ( 
.A(n_1573),
.Y(n_1952)
);

INVx2_ASAP7_75t_L g1953 ( 
.A(n_1502),
.Y(n_1953)
);

BUFx3_ASAP7_75t_L g1954 ( 
.A(n_1384),
.Y(n_1954)
);

HB1xp67_ASAP7_75t_L g1955 ( 
.A(n_1466),
.Y(n_1955)
);

INVxp67_ASAP7_75t_L g1956 ( 
.A(n_1463),
.Y(n_1956)
);

NAND2xp5_ASAP7_75t_L g1957 ( 
.A(n_1639),
.B(n_1060),
.Y(n_1957)
);

AND2x2_ASAP7_75t_L g1958 ( 
.A(n_1588),
.B(n_1299),
.Y(n_1958)
);

CKINVDCx6p67_ASAP7_75t_R g1959 ( 
.A(n_1626),
.Y(n_1959)
);

INVx2_ASAP7_75t_L g1960 ( 
.A(n_1502),
.Y(n_1960)
);

INVx2_ASAP7_75t_L g1961 ( 
.A(n_1514),
.Y(n_1961)
);

AND2x2_ASAP7_75t_L g1962 ( 
.A(n_1588),
.B(n_1300),
.Y(n_1962)
);

AND2x4_ASAP7_75t_L g1963 ( 
.A(n_1573),
.B(n_1061),
.Y(n_1963)
);

INVx1_ASAP7_75t_L g1964 ( 
.A(n_1618),
.Y(n_1964)
);

BUFx6f_ASAP7_75t_L g1965 ( 
.A(n_1418),
.Y(n_1965)
);

INVx1_ASAP7_75t_L g1966 ( 
.A(n_1618),
.Y(n_1966)
);

NAND2xp5_ASAP7_75t_L g1967 ( 
.A(n_1449),
.B(n_1065),
.Y(n_1967)
);

INVx1_ASAP7_75t_L g1968 ( 
.A(n_1470),
.Y(n_1968)
);

INVx3_ASAP7_75t_L g1969 ( 
.A(n_1420),
.Y(n_1969)
);

INVx1_ASAP7_75t_L g1970 ( 
.A(n_1470),
.Y(n_1970)
);

INVxp67_ASAP7_75t_L g1971 ( 
.A(n_1484),
.Y(n_1971)
);

INVx1_ASAP7_75t_L g1972 ( 
.A(n_1470),
.Y(n_1972)
);

INVx2_ASAP7_75t_L g1973 ( 
.A(n_1514),
.Y(n_1973)
);

BUFx6f_ASAP7_75t_L g1974 ( 
.A(n_1420),
.Y(n_1974)
);

BUFx6f_ASAP7_75t_L g1975 ( 
.A(n_1420),
.Y(n_1975)
);

AND2x4_ASAP7_75t_L g1976 ( 
.A(n_1384),
.B(n_1067),
.Y(n_1976)
);

XNOR2xp5_ASAP7_75t_L g1977 ( 
.A(n_1457),
.B(n_1041),
.Y(n_1977)
);

BUFx6f_ASAP7_75t_L g1978 ( 
.A(n_1420),
.Y(n_1978)
);

BUFx12f_ASAP7_75t_L g1979 ( 
.A(n_1360),
.Y(n_1979)
);

INVx2_ASAP7_75t_L g1980 ( 
.A(n_1514),
.Y(n_1980)
);

INVx1_ASAP7_75t_L g1981 ( 
.A(n_1470),
.Y(n_1981)
);

BUFx6f_ASAP7_75t_L g1982 ( 
.A(n_1424),
.Y(n_1982)
);

INVx1_ASAP7_75t_L g1983 ( 
.A(n_1514),
.Y(n_1983)
);

INVx2_ASAP7_75t_L g1984 ( 
.A(n_1523),
.Y(n_1984)
);

INVx3_ASAP7_75t_L g1985 ( 
.A(n_1424),
.Y(n_1985)
);

AND2x2_ASAP7_75t_L g1986 ( 
.A(n_1603),
.B(n_1301),
.Y(n_1986)
);

BUFx6f_ASAP7_75t_L g1987 ( 
.A(n_1424),
.Y(n_1987)
);

AND2x4_ASAP7_75t_L g1988 ( 
.A(n_1416),
.B(n_1068),
.Y(n_1988)
);

AND2x2_ASAP7_75t_L g1989 ( 
.A(n_1593),
.B(n_1302),
.Y(n_1989)
);

BUFx2_ASAP7_75t_L g1990 ( 
.A(n_1350),
.Y(n_1990)
);

NAND2xp5_ASAP7_75t_L g1991 ( 
.A(n_1472),
.B(n_1070),
.Y(n_1991)
);

INVx3_ASAP7_75t_L g1992 ( 
.A(n_1424),
.Y(n_1992)
);

CKINVDCx5p33_ASAP7_75t_R g1993 ( 
.A(n_1608),
.Y(n_1993)
);

OA21x2_ASAP7_75t_L g1994 ( 
.A1(n_1517),
.A2(n_1073),
.B(n_1072),
.Y(n_1994)
);

INVx3_ASAP7_75t_L g1995 ( 
.A(n_1430),
.Y(n_1995)
);

BUFx12f_ASAP7_75t_L g1996 ( 
.A(n_1360),
.Y(n_1996)
);

INVx2_ASAP7_75t_L g1997 ( 
.A(n_1523),
.Y(n_1997)
);

INVx3_ASAP7_75t_L g1998 ( 
.A(n_1430),
.Y(n_1998)
);

INVx1_ASAP7_75t_L g1999 ( 
.A(n_1523),
.Y(n_1999)
);

INVx1_ASAP7_75t_L g2000 ( 
.A(n_1523),
.Y(n_2000)
);

INVx1_ASAP7_75t_L g2001 ( 
.A(n_1541),
.Y(n_2001)
);

BUFx6f_ASAP7_75t_L g2002 ( 
.A(n_1430),
.Y(n_2002)
);

NAND2xp5_ASAP7_75t_L g2003 ( 
.A(n_1423),
.B(n_1076),
.Y(n_2003)
);

NAND2xp5_ASAP7_75t_SL g2004 ( 
.A(n_1593),
.B(n_1605),
.Y(n_2004)
);

INVx1_ASAP7_75t_L g2005 ( 
.A(n_1541),
.Y(n_2005)
);

INVx1_ASAP7_75t_L g2006 ( 
.A(n_1541),
.Y(n_2006)
);

NAND2xp5_ASAP7_75t_L g2007 ( 
.A(n_1423),
.B(n_1080),
.Y(n_2007)
);

BUFx6f_ASAP7_75t_L g2008 ( 
.A(n_1430),
.Y(n_2008)
);

INVx2_ASAP7_75t_L g2009 ( 
.A(n_1541),
.Y(n_2009)
);

INVx1_ASAP7_75t_L g2010 ( 
.A(n_1542),
.Y(n_2010)
);

INVx2_ASAP7_75t_L g2011 ( 
.A(n_1542),
.Y(n_2011)
);

NAND2xp5_ASAP7_75t_L g2012 ( 
.A(n_1426),
.B(n_1081),
.Y(n_2012)
);

INVx1_ASAP7_75t_L g2013 ( 
.A(n_1542),
.Y(n_2013)
);

INVx8_ASAP7_75t_L g2014 ( 
.A(n_1905),
.Y(n_2014)
);

OR2x2_ASAP7_75t_L g2015 ( 
.A(n_1671),
.B(n_1466),
.Y(n_2015)
);

INVx1_ASAP7_75t_L g2016 ( 
.A(n_1690),
.Y(n_2016)
);

INVx2_ASAP7_75t_L g2017 ( 
.A(n_1826),
.Y(n_2017)
);

BUFx10_ASAP7_75t_L g2018 ( 
.A(n_1759),
.Y(n_2018)
);

INVx1_ASAP7_75t_L g2019 ( 
.A(n_1690),
.Y(n_2019)
);

INVx2_ASAP7_75t_L g2020 ( 
.A(n_1826),
.Y(n_2020)
);

INVx1_ASAP7_75t_L g2021 ( 
.A(n_1690),
.Y(n_2021)
);

INVx1_ASAP7_75t_L g2022 ( 
.A(n_1747),
.Y(n_2022)
);

NOR2xp33_ASAP7_75t_L g2023 ( 
.A(n_1714),
.B(n_1484),
.Y(n_2023)
);

INVx1_ASAP7_75t_L g2024 ( 
.A(n_1747),
.Y(n_2024)
);

INVx8_ASAP7_75t_L g2025 ( 
.A(n_1905),
.Y(n_2025)
);

INVx3_ASAP7_75t_L g2026 ( 
.A(n_1747),
.Y(n_2026)
);

BUFx6f_ASAP7_75t_L g2027 ( 
.A(n_1826),
.Y(n_2027)
);

NAND3xp33_ASAP7_75t_L g2028 ( 
.A(n_1849),
.B(n_1648),
.C(n_1435),
.Y(n_2028)
);

INVx2_ASAP7_75t_L g2029 ( 
.A(n_1850),
.Y(n_2029)
);

INVx2_ASAP7_75t_L g2030 ( 
.A(n_1850),
.Y(n_2030)
);

NAND2xp5_ASAP7_75t_SL g2031 ( 
.A(n_1670),
.B(n_1651),
.Y(n_2031)
);

INVx2_ASAP7_75t_L g2032 ( 
.A(n_1850),
.Y(n_2032)
);

CKINVDCx5p33_ASAP7_75t_R g2033 ( 
.A(n_1853),
.Y(n_2033)
);

INVx1_ASAP7_75t_L g2034 ( 
.A(n_1902),
.Y(n_2034)
);

BUFx3_ASAP7_75t_L g2035 ( 
.A(n_1954),
.Y(n_2035)
);

INVx2_ASAP7_75t_L g2036 ( 
.A(n_1677),
.Y(n_2036)
);

NOR2x1p5_ASAP7_75t_L g2037 ( 
.A(n_1979),
.B(n_1996),
.Y(n_2037)
);

INVx1_ASAP7_75t_L g2038 ( 
.A(n_1902),
.Y(n_2038)
);

INVx1_ASAP7_75t_L g2039 ( 
.A(n_1902),
.Y(n_2039)
);

NAND2xp5_ASAP7_75t_SL g2040 ( 
.A(n_1692),
.B(n_1651),
.Y(n_2040)
);

NAND2xp5_ASAP7_75t_SL g2041 ( 
.A(n_1707),
.B(n_1397),
.Y(n_2041)
);

INVx2_ASAP7_75t_SL g2042 ( 
.A(n_1843),
.Y(n_2042)
);

INVx1_ASAP7_75t_L g2043 ( 
.A(n_1866),
.Y(n_2043)
);

INVx8_ASAP7_75t_L g2044 ( 
.A(n_1905),
.Y(n_2044)
);

INVx1_ASAP7_75t_L g2045 ( 
.A(n_1866),
.Y(n_2045)
);

NAND2xp5_ASAP7_75t_SL g2046 ( 
.A(n_1832),
.B(n_1488),
.Y(n_2046)
);

INVx2_ASAP7_75t_L g2047 ( 
.A(n_1677),
.Y(n_2047)
);

INVx2_ASAP7_75t_L g2048 ( 
.A(n_1679),
.Y(n_2048)
);

INVx1_ASAP7_75t_L g2049 ( 
.A(n_1866),
.Y(n_2049)
);

INVx2_ASAP7_75t_L g2050 ( 
.A(n_1679),
.Y(n_2050)
);

BUFx3_ASAP7_75t_L g2051 ( 
.A(n_1954),
.Y(n_2051)
);

OAI22xp5_ASAP7_75t_L g2052 ( 
.A1(n_1753),
.A2(n_1506),
.B1(n_1606),
.B2(n_1487),
.Y(n_2052)
);

INVx2_ASAP7_75t_L g2053 ( 
.A(n_1685),
.Y(n_2053)
);

NOR2xp33_ASAP7_75t_L g2054 ( 
.A(n_1765),
.B(n_1518),
.Y(n_2054)
);

AND2x2_ASAP7_75t_L g2055 ( 
.A(n_1719),
.B(n_1605),
.Y(n_2055)
);

INVx1_ASAP7_75t_L g2056 ( 
.A(n_1782),
.Y(n_2056)
);

NAND2xp5_ASAP7_75t_L g2057 ( 
.A(n_1849),
.B(n_1648),
.Y(n_2057)
);

INVx2_ASAP7_75t_L g2058 ( 
.A(n_1685),
.Y(n_2058)
);

NAND2xp5_ASAP7_75t_L g2059 ( 
.A(n_1723),
.B(n_1617),
.Y(n_2059)
);

INVxp67_ASAP7_75t_L g2060 ( 
.A(n_1666),
.Y(n_2060)
);

INVxp33_ASAP7_75t_L g2061 ( 
.A(n_1928),
.Y(n_2061)
);

INVx1_ASAP7_75t_L g2062 ( 
.A(n_1782),
.Y(n_2062)
);

INVx1_ASAP7_75t_L g2063 ( 
.A(n_1789),
.Y(n_2063)
);

INVx2_ASAP7_75t_L g2064 ( 
.A(n_1693),
.Y(n_2064)
);

HB1xp67_ASAP7_75t_L g2065 ( 
.A(n_1928),
.Y(n_2065)
);

INVx2_ASAP7_75t_L g2066 ( 
.A(n_1693),
.Y(n_2066)
);

INVx1_ASAP7_75t_L g2067 ( 
.A(n_1789),
.Y(n_2067)
);

OR2x2_ASAP7_75t_L g2068 ( 
.A(n_1778),
.B(n_1483),
.Y(n_2068)
);

INVx1_ASAP7_75t_L g2069 ( 
.A(n_1793),
.Y(n_2069)
);

INVx1_ASAP7_75t_SL g2070 ( 
.A(n_1804),
.Y(n_2070)
);

INVx1_ASAP7_75t_L g2071 ( 
.A(n_1793),
.Y(n_2071)
);

NAND2xp5_ASAP7_75t_SL g2072 ( 
.A(n_1832),
.B(n_1856),
.Y(n_2072)
);

AND3x2_ASAP7_75t_L g2073 ( 
.A(n_1929),
.B(n_1563),
.C(n_1535),
.Y(n_2073)
);

INVx1_ASAP7_75t_L g2074 ( 
.A(n_1796),
.Y(n_2074)
);

INVx2_ASAP7_75t_L g2075 ( 
.A(n_1696),
.Y(n_2075)
);

INVx2_ASAP7_75t_SL g2076 ( 
.A(n_1843),
.Y(n_2076)
);

INVx1_ASAP7_75t_L g2077 ( 
.A(n_1796),
.Y(n_2077)
);

OAI22xp33_ASAP7_75t_L g2078 ( 
.A1(n_1839),
.A2(n_1530),
.B1(n_1487),
.B2(n_1465),
.Y(n_2078)
);

BUFx6f_ASAP7_75t_L g2079 ( 
.A(n_1700),
.Y(n_2079)
);

BUFx6f_ASAP7_75t_SL g2080 ( 
.A(n_1976),
.Y(n_2080)
);

INVx3_ASAP7_75t_L g2081 ( 
.A(n_1696),
.Y(n_2081)
);

INVx2_ASAP7_75t_L g2082 ( 
.A(n_1697),
.Y(n_2082)
);

NAND2xp5_ASAP7_75t_SL g2083 ( 
.A(n_1856),
.B(n_1488),
.Y(n_2083)
);

INVx3_ASAP7_75t_L g2084 ( 
.A(n_1697),
.Y(n_2084)
);

INVx1_ASAP7_75t_L g2085 ( 
.A(n_1705),
.Y(n_2085)
);

BUFx6f_ASAP7_75t_L g2086 ( 
.A(n_1700),
.Y(n_2086)
);

NOR2xp33_ASAP7_75t_L g2087 ( 
.A(n_1871),
.B(n_1518),
.Y(n_2087)
);

INVx2_ASAP7_75t_L g2088 ( 
.A(n_1705),
.Y(n_2088)
);

AO21x2_ASAP7_75t_L g2089 ( 
.A1(n_1812),
.A2(n_1630),
.B(n_1402),
.Y(n_2089)
);

AND2x2_ASAP7_75t_L g2090 ( 
.A(n_1719),
.B(n_1617),
.Y(n_2090)
);

INVx3_ASAP7_75t_L g2091 ( 
.A(n_1712),
.Y(n_2091)
);

INVx2_ASAP7_75t_L g2092 ( 
.A(n_1712),
.Y(n_2092)
);

NOR2xp33_ASAP7_75t_SL g2093 ( 
.A(n_1759),
.B(n_1800),
.Y(n_2093)
);

AND2x2_ASAP7_75t_L g2094 ( 
.A(n_1809),
.B(n_1497),
.Y(n_2094)
);

NAND2xp5_ASAP7_75t_SL g2095 ( 
.A(n_1800),
.B(n_1590),
.Y(n_2095)
);

INVx2_ASAP7_75t_L g2096 ( 
.A(n_1717),
.Y(n_2096)
);

AO21x2_ASAP7_75t_L g2097 ( 
.A1(n_1812),
.A2(n_1402),
.B(n_1476),
.Y(n_2097)
);

HB1xp67_ASAP7_75t_L g2098 ( 
.A(n_1912),
.Y(n_2098)
);

INVx2_ASAP7_75t_L g2099 ( 
.A(n_1717),
.Y(n_2099)
);

INVx2_ASAP7_75t_SL g2100 ( 
.A(n_1843),
.Y(n_2100)
);

AND2x2_ASAP7_75t_L g2101 ( 
.A(n_1676),
.B(n_1416),
.Y(n_2101)
);

INVx2_ASAP7_75t_L g2102 ( 
.A(n_1726),
.Y(n_2102)
);

INVx2_ASAP7_75t_L g2103 ( 
.A(n_1726),
.Y(n_2103)
);

INVx1_ASAP7_75t_L g2104 ( 
.A(n_1737),
.Y(n_2104)
);

INVx1_ASAP7_75t_L g2105 ( 
.A(n_1737),
.Y(n_2105)
);

INVx2_ASAP7_75t_L g2106 ( 
.A(n_1744),
.Y(n_2106)
);

INVx1_ASAP7_75t_L g2107 ( 
.A(n_1744),
.Y(n_2107)
);

NAND2xp5_ASAP7_75t_SL g2108 ( 
.A(n_1956),
.B(n_1971),
.Y(n_2108)
);

AND2x2_ASAP7_75t_L g2109 ( 
.A(n_1676),
.B(n_1658),
.Y(n_2109)
);

INVx1_ASAP7_75t_L g2110 ( 
.A(n_1745),
.Y(n_2110)
);

INVx2_ASAP7_75t_L g2111 ( 
.A(n_1745),
.Y(n_2111)
);

NOR2x1p5_ASAP7_75t_L g2112 ( 
.A(n_1979),
.B(n_1504),
.Y(n_2112)
);

NAND2xp5_ASAP7_75t_SL g2113 ( 
.A(n_1741),
.B(n_1590),
.Y(n_2113)
);

INVx2_ASAP7_75t_L g2114 ( 
.A(n_1751),
.Y(n_2114)
);

AO21x2_ASAP7_75t_L g2115 ( 
.A1(n_1914),
.A2(n_1476),
.B(n_1393),
.Y(n_2115)
);

INVx11_ASAP7_75t_L g2116 ( 
.A(n_1686),
.Y(n_2116)
);

INVx2_ASAP7_75t_L g2117 ( 
.A(n_1751),
.Y(n_2117)
);

NAND2xp5_ASAP7_75t_L g2118 ( 
.A(n_1891),
.B(n_1426),
.Y(n_2118)
);

INVx2_ASAP7_75t_L g2119 ( 
.A(n_1733),
.Y(n_2119)
);

INVx1_ASAP7_75t_L g2120 ( 
.A(n_1738),
.Y(n_2120)
);

NAND2xp5_ASAP7_75t_L g2121 ( 
.A(n_1894),
.B(n_1435),
.Y(n_2121)
);

AND2x2_ASAP7_75t_SL g2122 ( 
.A(n_1725),
.B(n_1528),
.Y(n_2122)
);

INVx1_ASAP7_75t_L g2123 ( 
.A(n_1739),
.Y(n_2123)
);

INVx2_ASAP7_75t_L g2124 ( 
.A(n_1740),
.Y(n_2124)
);

INVx2_ASAP7_75t_L g2125 ( 
.A(n_1752),
.Y(n_2125)
);

INVx3_ASAP7_75t_L g2126 ( 
.A(n_1797),
.Y(n_2126)
);

INVx4_ASAP7_75t_L g2127 ( 
.A(n_1935),
.Y(n_2127)
);

INVx1_ASAP7_75t_L g2128 ( 
.A(n_1754),
.Y(n_2128)
);

INVx1_ASAP7_75t_L g2129 ( 
.A(n_1755),
.Y(n_2129)
);

CKINVDCx16_ASAP7_75t_R g2130 ( 
.A(n_1774),
.Y(n_2130)
);

OR2x2_ASAP7_75t_L g2131 ( 
.A(n_1778),
.B(n_1483),
.Y(n_2131)
);

NAND2xp5_ASAP7_75t_SL g2132 ( 
.A(n_1767),
.B(n_1597),
.Y(n_2132)
);

INVx1_ASAP7_75t_L g2133 ( 
.A(n_1756),
.Y(n_2133)
);

NAND2xp5_ASAP7_75t_L g2134 ( 
.A(n_1967),
.B(n_1991),
.Y(n_2134)
);

INVx1_ASAP7_75t_L g2135 ( 
.A(n_1758),
.Y(n_2135)
);

INVx2_ASAP7_75t_SL g2136 ( 
.A(n_1880),
.Y(n_2136)
);

NAND2xp5_ASAP7_75t_SL g2137 ( 
.A(n_2004),
.B(n_1597),
.Y(n_2137)
);

INVx2_ASAP7_75t_L g2138 ( 
.A(n_1761),
.Y(n_2138)
);

INVx2_ASAP7_75t_L g2139 ( 
.A(n_1927),
.Y(n_2139)
);

INVx1_ASAP7_75t_L g2140 ( 
.A(n_1921),
.Y(n_2140)
);

NAND2xp5_ASAP7_75t_SL g2141 ( 
.A(n_2004),
.B(n_1634),
.Y(n_2141)
);

INVx2_ASAP7_75t_L g2142 ( 
.A(n_1927),
.Y(n_2142)
);

INVx2_ASAP7_75t_L g2143 ( 
.A(n_1923),
.Y(n_2143)
);

INVx2_ASAP7_75t_L g2144 ( 
.A(n_1797),
.Y(n_2144)
);

NAND2xp5_ASAP7_75t_SL g2145 ( 
.A(n_1673),
.B(n_1634),
.Y(n_2145)
);

NAND2xp5_ASAP7_75t_SL g2146 ( 
.A(n_1731),
.B(n_1482),
.Y(n_2146)
);

INVx1_ASAP7_75t_L g2147 ( 
.A(n_1951),
.Y(n_2147)
);

INVx3_ASAP7_75t_L g2148 ( 
.A(n_1806),
.Y(n_2148)
);

AND2x2_ASAP7_75t_L g2149 ( 
.A(n_1868),
.B(n_1788),
.Y(n_2149)
);

INVx2_ASAP7_75t_L g2150 ( 
.A(n_1806),
.Y(n_2150)
);

NAND2xp5_ASAP7_75t_L g2151 ( 
.A(n_1807),
.B(n_1528),
.Y(n_2151)
);

INVx2_ASAP7_75t_L g2152 ( 
.A(n_1817),
.Y(n_2152)
);

INVx2_ASAP7_75t_L g2153 ( 
.A(n_1817),
.Y(n_2153)
);

NAND2xp5_ASAP7_75t_SL g2154 ( 
.A(n_1748),
.B(n_1490),
.Y(n_2154)
);

NAND2xp5_ASAP7_75t_L g2155 ( 
.A(n_1803),
.B(n_1556),
.Y(n_2155)
);

INVx1_ASAP7_75t_L g2156 ( 
.A(n_1952),
.Y(n_2156)
);

INVx2_ASAP7_75t_L g2157 ( 
.A(n_1846),
.Y(n_2157)
);

BUFx2_ASAP7_75t_L g2158 ( 
.A(n_1810),
.Y(n_2158)
);

INVx2_ASAP7_75t_L g2159 ( 
.A(n_1846),
.Y(n_2159)
);

OR2x2_ASAP7_75t_L g2160 ( 
.A(n_1821),
.B(n_1493),
.Y(n_2160)
);

INVx1_ASAP7_75t_L g2161 ( 
.A(n_1964),
.Y(n_2161)
);

INVx2_ASAP7_75t_L g2162 ( 
.A(n_1862),
.Y(n_2162)
);

NAND2xp5_ASAP7_75t_SL g2163 ( 
.A(n_1773),
.B(n_1498),
.Y(n_2163)
);

AO21x2_ASAP7_75t_L g2164 ( 
.A1(n_1914),
.A2(n_1395),
.B(n_1390),
.Y(n_2164)
);

INVx2_ASAP7_75t_L g2165 ( 
.A(n_1862),
.Y(n_2165)
);

INVx1_ASAP7_75t_L g2166 ( 
.A(n_1966),
.Y(n_2166)
);

NAND2xp5_ASAP7_75t_L g2167 ( 
.A(n_1934),
.B(n_1556),
.Y(n_2167)
);

INVx2_ASAP7_75t_L g2168 ( 
.A(n_1877),
.Y(n_2168)
);

CKINVDCx6p67_ASAP7_75t_R g2169 ( 
.A(n_1996),
.Y(n_2169)
);

INVx4_ASAP7_75t_L g2170 ( 
.A(n_1935),
.Y(n_2170)
);

NAND2xp5_ASAP7_75t_L g2171 ( 
.A(n_1939),
.B(n_1943),
.Y(n_2171)
);

INVx2_ASAP7_75t_L g2172 ( 
.A(n_1877),
.Y(n_2172)
);

NAND2xp5_ASAP7_75t_L g2173 ( 
.A(n_1946),
.B(n_1957),
.Y(n_2173)
);

INVx2_ASAP7_75t_L g2174 ( 
.A(n_1878),
.Y(n_2174)
);

INVx2_ASAP7_75t_L g2175 ( 
.A(n_1878),
.Y(n_2175)
);

AND2x4_ASAP7_75t_L g2176 ( 
.A(n_1825),
.B(n_1421),
.Y(n_2176)
);

INVx2_ASAP7_75t_L g2177 ( 
.A(n_1882),
.Y(n_2177)
);

INVx2_ASAP7_75t_L g2178 ( 
.A(n_1882),
.Y(n_2178)
);

INVx2_ASAP7_75t_L g2179 ( 
.A(n_1887),
.Y(n_2179)
);

AND3x2_ASAP7_75t_L g2180 ( 
.A(n_1675),
.B(n_1650),
.C(n_1610),
.Y(n_2180)
);

INVx3_ASAP7_75t_L g2181 ( 
.A(n_1887),
.Y(n_2181)
);

AND2x2_ASAP7_75t_L g2182 ( 
.A(n_1868),
.B(n_1658),
.Y(n_2182)
);

INVx1_ASAP7_75t_L g2183 ( 
.A(n_1895),
.Y(n_2183)
);

NAND2xp5_ASAP7_75t_L g2184 ( 
.A(n_1837),
.B(n_1574),
.Y(n_2184)
);

INVx1_ASAP7_75t_L g2185 ( 
.A(n_1895),
.Y(n_2185)
);

INVx2_ASAP7_75t_SL g2186 ( 
.A(n_1880),
.Y(n_2186)
);

INVx1_ASAP7_75t_L g2187 ( 
.A(n_1896),
.Y(n_2187)
);

BUFx6f_ASAP7_75t_L g2188 ( 
.A(n_1700),
.Y(n_2188)
);

INVx2_ASAP7_75t_SL g2189 ( 
.A(n_1880),
.Y(n_2189)
);

INVx4_ASAP7_75t_L g2190 ( 
.A(n_1935),
.Y(n_2190)
);

INVx1_ASAP7_75t_L g2191 ( 
.A(n_1896),
.Y(n_2191)
);

INVx2_ASAP7_75t_L g2192 ( 
.A(n_1899),
.Y(n_2192)
);

INVx1_ASAP7_75t_L g2193 ( 
.A(n_1899),
.Y(n_2193)
);

INVx1_ASAP7_75t_L g2194 ( 
.A(n_1900),
.Y(n_2194)
);

INVx1_ASAP7_75t_L g2195 ( 
.A(n_1900),
.Y(n_2195)
);

INVx2_ASAP7_75t_L g2196 ( 
.A(n_1903),
.Y(n_2196)
);

INVxp33_ASAP7_75t_L g2197 ( 
.A(n_1955),
.Y(n_2197)
);

AOI22xp33_ASAP7_75t_L g2198 ( 
.A1(n_1845),
.A2(n_1437),
.B1(n_1461),
.B2(n_1433),
.Y(n_2198)
);

INVx1_ASAP7_75t_L g2199 ( 
.A(n_1903),
.Y(n_2199)
);

INVx1_ASAP7_75t_L g2200 ( 
.A(n_1936),
.Y(n_2200)
);

INVx2_ASAP7_75t_L g2201 ( 
.A(n_1936),
.Y(n_2201)
);

BUFx2_ASAP7_75t_L g2202 ( 
.A(n_1829),
.Y(n_2202)
);

INVx2_ASAP7_75t_L g2203 ( 
.A(n_1938),
.Y(n_2203)
);

AND2x2_ASAP7_75t_L g2204 ( 
.A(n_1788),
.B(n_1949),
.Y(n_2204)
);

INVx2_ASAP7_75t_SL g2205 ( 
.A(n_1897),
.Y(n_2205)
);

INVx4_ASAP7_75t_L g2206 ( 
.A(n_1935),
.Y(n_2206)
);

INVx3_ASAP7_75t_L g2207 ( 
.A(n_1938),
.Y(n_2207)
);

OAI22xp5_ASAP7_75t_L g2208 ( 
.A1(n_2003),
.A2(n_1606),
.B1(n_1465),
.B2(n_1572),
.Y(n_2208)
);

INVx3_ASAP7_75t_L g2209 ( 
.A(n_1944),
.Y(n_2209)
);

NAND2xp33_ASAP7_75t_L g2210 ( 
.A(n_1700),
.B(n_1405),
.Y(n_2210)
);

INVx2_ASAP7_75t_L g2211 ( 
.A(n_1944),
.Y(n_2211)
);

INVx2_ASAP7_75t_L g2212 ( 
.A(n_1948),
.Y(n_2212)
);

NOR2xp33_ASAP7_75t_L g2213 ( 
.A(n_1776),
.B(n_1574),
.Y(n_2213)
);

BUFx3_ASAP7_75t_L g2214 ( 
.A(n_1660),
.Y(n_2214)
);

NAND2xp5_ASAP7_75t_L g2215 ( 
.A(n_1905),
.B(n_1840),
.Y(n_2215)
);

INVx2_ASAP7_75t_L g2216 ( 
.A(n_1948),
.Y(n_2216)
);

NOR2xp33_ASAP7_75t_L g2217 ( 
.A(n_1786),
.B(n_1577),
.Y(n_2217)
);

NAND2xp5_ASAP7_75t_SL g2218 ( 
.A(n_1775),
.B(n_1547),
.Y(n_2218)
);

INVx3_ASAP7_75t_L g2219 ( 
.A(n_1953),
.Y(n_2219)
);

NAND3xp33_ASAP7_75t_L g2220 ( 
.A(n_2007),
.B(n_1657),
.C(n_1645),
.Y(n_2220)
);

BUFx10_ASAP7_75t_L g2221 ( 
.A(n_1684),
.Y(n_2221)
);

INVx2_ASAP7_75t_L g2222 ( 
.A(n_1953),
.Y(n_2222)
);

INVx1_ASAP7_75t_L g2223 ( 
.A(n_1960),
.Y(n_2223)
);

INVx2_ASAP7_75t_L g2224 ( 
.A(n_1960),
.Y(n_2224)
);

INVx1_ASAP7_75t_L g2225 ( 
.A(n_1961),
.Y(n_2225)
);

NAND2xp5_ASAP7_75t_L g2226 ( 
.A(n_1905),
.B(n_1577),
.Y(n_2226)
);

INVx1_ASAP7_75t_L g2227 ( 
.A(n_1961),
.Y(n_2227)
);

INVx2_ASAP7_75t_L g2228 ( 
.A(n_1973),
.Y(n_2228)
);

INVx2_ASAP7_75t_L g2229 ( 
.A(n_1973),
.Y(n_2229)
);

INVx1_ASAP7_75t_L g2230 ( 
.A(n_1980),
.Y(n_2230)
);

AND2x2_ASAP7_75t_L g2231 ( 
.A(n_1958),
.B(n_1421),
.Y(n_2231)
);

OR2x2_ASAP7_75t_L g2232 ( 
.A(n_1821),
.B(n_1493),
.Y(n_2232)
);

OR2x2_ASAP7_75t_L g2233 ( 
.A(n_1827),
.B(n_1650),
.Y(n_2233)
);

INVx2_ASAP7_75t_L g2234 ( 
.A(n_1980),
.Y(n_2234)
);

AND2x2_ASAP7_75t_L g2235 ( 
.A(n_1962),
.B(n_1653),
.Y(n_2235)
);

INVx1_ASAP7_75t_L g2236 ( 
.A(n_1984),
.Y(n_2236)
);

NOR2xp33_ASAP7_75t_L g2237 ( 
.A(n_1790),
.B(n_1601),
.Y(n_2237)
);

INVx1_ASAP7_75t_SL g2238 ( 
.A(n_1942),
.Y(n_2238)
);

NAND2xp5_ASAP7_75t_SL g2239 ( 
.A(n_1820),
.B(n_1571),
.Y(n_2239)
);

INVx2_ASAP7_75t_L g2240 ( 
.A(n_1984),
.Y(n_2240)
);

INVx2_ASAP7_75t_L g2241 ( 
.A(n_1997),
.Y(n_2241)
);

INVx1_ASAP7_75t_L g2242 ( 
.A(n_1997),
.Y(n_2242)
);

NAND2xp5_ASAP7_75t_SL g2243 ( 
.A(n_1851),
.B(n_1615),
.Y(n_2243)
);

INVx2_ASAP7_75t_L g2244 ( 
.A(n_2009),
.Y(n_2244)
);

INVx4_ASAP7_75t_L g2245 ( 
.A(n_1937),
.Y(n_2245)
);

NAND2xp5_ASAP7_75t_SL g2246 ( 
.A(n_1842),
.B(n_1643),
.Y(n_2246)
);

INVx2_ASAP7_75t_L g2247 ( 
.A(n_2009),
.Y(n_2247)
);

BUFx2_ASAP7_75t_L g2248 ( 
.A(n_1827),
.Y(n_2248)
);

BUFx10_ASAP7_75t_L g2249 ( 
.A(n_1684),
.Y(n_2249)
);

INVx4_ASAP7_75t_L g2250 ( 
.A(n_1937),
.Y(n_2250)
);

AND2x2_ASAP7_75t_L g2251 ( 
.A(n_1989),
.B(n_1655),
.Y(n_2251)
);

NAND2xp5_ASAP7_75t_SL g2252 ( 
.A(n_1710),
.B(n_1475),
.Y(n_2252)
);

INVx2_ASAP7_75t_L g2253 ( 
.A(n_2011),
.Y(n_2253)
);

INVx3_ASAP7_75t_L g2254 ( 
.A(n_2011),
.Y(n_2254)
);

INVx2_ASAP7_75t_L g2255 ( 
.A(n_1875),
.Y(n_2255)
);

NAND2xp33_ASAP7_75t_L g2256 ( 
.A(n_1700),
.B(n_1511),
.Y(n_2256)
);

NAND2xp5_ASAP7_75t_L g2257 ( 
.A(n_2012),
.B(n_1601),
.Y(n_2257)
);

INVx2_ASAP7_75t_SL g2258 ( 
.A(n_1897),
.Y(n_2258)
);

INVx1_ASAP7_75t_SL g2259 ( 
.A(n_1955),
.Y(n_2259)
);

INVx3_ASAP7_75t_L g2260 ( 
.A(n_1969),
.Y(n_2260)
);

INVx1_ASAP7_75t_L g2261 ( 
.A(n_1933),
.Y(n_2261)
);

NAND2xp5_ASAP7_75t_L g2262 ( 
.A(n_1845),
.B(n_1631),
.Y(n_2262)
);

BUFx3_ASAP7_75t_L g2263 ( 
.A(n_1660),
.Y(n_2263)
);

INVx2_ASAP7_75t_L g2264 ( 
.A(n_1875),
.Y(n_2264)
);

INVx2_ASAP7_75t_L g2265 ( 
.A(n_1986),
.Y(n_2265)
);

NAND2xp5_ASAP7_75t_L g2266 ( 
.A(n_1845),
.B(n_1631),
.Y(n_2266)
);

INVx2_ASAP7_75t_L g2267 ( 
.A(n_1986),
.Y(n_2267)
);

INVx1_ASAP7_75t_L g2268 ( 
.A(n_1945),
.Y(n_2268)
);

NAND2xp5_ASAP7_75t_SL g2269 ( 
.A(n_1907),
.B(n_1647),
.Y(n_2269)
);

NAND2xp5_ASAP7_75t_L g2270 ( 
.A(n_1845),
.B(n_1640),
.Y(n_2270)
);

INVx3_ASAP7_75t_L g2271 ( 
.A(n_1969),
.Y(n_2271)
);

INVx2_ASAP7_75t_L g2272 ( 
.A(n_1947),
.Y(n_2272)
);

INVx2_ASAP7_75t_L g2273 ( 
.A(n_1994),
.Y(n_2273)
);

INVx2_ASAP7_75t_L g2274 ( 
.A(n_1994),
.Y(n_2274)
);

INVx2_ASAP7_75t_L g2275 ( 
.A(n_1994),
.Y(n_2275)
);

INVx1_ASAP7_75t_L g2276 ( 
.A(n_1664),
.Y(n_2276)
);

NAND2xp5_ASAP7_75t_L g2277 ( 
.A(n_1845),
.B(n_1640),
.Y(n_2277)
);

NAND2xp33_ASAP7_75t_L g2278 ( 
.A(n_1865),
.B(n_1621),
.Y(n_2278)
);

BUFx6f_ASAP7_75t_L g2279 ( 
.A(n_1663),
.Y(n_2279)
);

NAND2xp5_ASAP7_75t_SL g2280 ( 
.A(n_1911),
.B(n_1513),
.Y(n_2280)
);

INVx1_ASAP7_75t_L g2281 ( 
.A(n_1665),
.Y(n_2281)
);

INVx3_ASAP7_75t_L g2282 ( 
.A(n_1969),
.Y(n_2282)
);

NAND2xp5_ASAP7_75t_L g2283 ( 
.A(n_1916),
.B(n_1642),
.Y(n_2283)
);

INVx1_ASAP7_75t_L g2284 ( 
.A(n_1667),
.Y(n_2284)
);

INVx2_ASAP7_75t_L g2285 ( 
.A(n_1985),
.Y(n_2285)
);

NAND2xp5_ASAP7_75t_L g2286 ( 
.A(n_1930),
.B(n_1642),
.Y(n_2286)
);

INVx3_ASAP7_75t_L g2287 ( 
.A(n_1985),
.Y(n_2287)
);

INVx1_ASAP7_75t_L g2288 ( 
.A(n_1668),
.Y(n_2288)
);

AND3x2_ASAP7_75t_L g2289 ( 
.A(n_1687),
.B(n_1760),
.C(n_1610),
.Y(n_2289)
);

INVx2_ASAP7_75t_L g2290 ( 
.A(n_1985),
.Y(n_2290)
);

INVx1_ASAP7_75t_L g2291 ( 
.A(n_1674),
.Y(n_2291)
);

INVx3_ASAP7_75t_L g2292 ( 
.A(n_1992),
.Y(n_2292)
);

NAND2xp5_ASAP7_75t_SL g2293 ( 
.A(n_1734),
.B(n_1572),
.Y(n_2293)
);

XOR2xp5_ASAP7_75t_L g2294 ( 
.A(n_1977),
.B(n_1046),
.Y(n_2294)
);

AND2x2_ASAP7_75t_L g2295 ( 
.A(n_1976),
.B(n_1653),
.Y(n_2295)
);

INVx2_ASAP7_75t_L g2296 ( 
.A(n_1992),
.Y(n_2296)
);

INVx2_ASAP7_75t_L g2297 ( 
.A(n_1992),
.Y(n_2297)
);

AOI22xp33_ASAP7_75t_L g2298 ( 
.A1(n_1892),
.A2(n_1931),
.B1(n_1695),
.B2(n_1701),
.Y(n_2298)
);

INVx8_ASAP7_75t_L g2299 ( 
.A(n_1976),
.Y(n_2299)
);

INVx3_ASAP7_75t_L g2300 ( 
.A(n_1995),
.Y(n_2300)
);

INVx2_ASAP7_75t_L g2301 ( 
.A(n_1995),
.Y(n_2301)
);

INVx2_ASAP7_75t_SL g2302 ( 
.A(n_1897),
.Y(n_2302)
);

INVx2_ASAP7_75t_L g2303 ( 
.A(n_1995),
.Y(n_2303)
);

INVx2_ASAP7_75t_L g2304 ( 
.A(n_1998),
.Y(n_2304)
);

AND2x2_ASAP7_75t_L g2305 ( 
.A(n_1988),
.B(n_1655),
.Y(n_2305)
);

INVx2_ASAP7_75t_SL g2306 ( 
.A(n_1694),
.Y(n_2306)
);

INVx2_ASAP7_75t_L g2307 ( 
.A(n_1998),
.Y(n_2307)
);

INVx2_ASAP7_75t_L g2308 ( 
.A(n_1998),
.Y(n_2308)
);

NAND2xp5_ASAP7_75t_L g2309 ( 
.A(n_1857),
.B(n_1645),
.Y(n_2309)
);

INVx2_ASAP7_75t_L g2310 ( 
.A(n_1681),
.Y(n_2310)
);

BUFx10_ASAP7_75t_L g2311 ( 
.A(n_1660),
.Y(n_2311)
);

INVx2_ASAP7_75t_L g2312 ( 
.A(n_1681),
.Y(n_2312)
);

INVx3_ASAP7_75t_L g2313 ( 
.A(n_1681),
.Y(n_2313)
);

NAND2xp5_ASAP7_75t_L g2314 ( 
.A(n_1879),
.B(n_1657),
.Y(n_2314)
);

INVx1_ASAP7_75t_L g2315 ( 
.A(n_1678),
.Y(n_2315)
);

AND2x4_ASAP7_75t_L g2316 ( 
.A(n_1825),
.B(n_1603),
.Y(n_2316)
);

INVx2_ASAP7_75t_L g2317 ( 
.A(n_1688),
.Y(n_2317)
);

NOR2xp33_ASAP7_75t_L g2318 ( 
.A(n_1770),
.B(n_1501),
.Y(n_2318)
);

AND2x2_ASAP7_75t_L g2319 ( 
.A(n_1988),
.B(n_1619),
.Y(n_2319)
);

INVx8_ASAP7_75t_L g2320 ( 
.A(n_1988),
.Y(n_2320)
);

NAND2xp5_ASAP7_75t_L g2321 ( 
.A(n_1884),
.B(n_1505),
.Y(n_2321)
);

INVx3_ASAP7_75t_L g2322 ( 
.A(n_1688),
.Y(n_2322)
);

INVx1_ASAP7_75t_L g2323 ( 
.A(n_1702),
.Y(n_2323)
);

INVx2_ASAP7_75t_L g2324 ( 
.A(n_1688),
.Y(n_2324)
);

NOR2xp33_ASAP7_75t_SL g2325 ( 
.A(n_1864),
.B(n_1504),
.Y(n_2325)
);

INVx2_ASAP7_75t_L g2326 ( 
.A(n_1689),
.Y(n_2326)
);

INVx1_ASAP7_75t_L g2327 ( 
.A(n_1704),
.Y(n_2327)
);

INVx2_ASAP7_75t_L g2328 ( 
.A(n_1689),
.Y(n_2328)
);

INVx4_ASAP7_75t_L g2329 ( 
.A(n_1937),
.Y(n_2329)
);

INVx2_ASAP7_75t_L g2330 ( 
.A(n_1689),
.Y(n_2330)
);

INVx2_ASAP7_75t_L g2331 ( 
.A(n_1713),
.Y(n_2331)
);

NAND2xp5_ASAP7_75t_SL g2332 ( 
.A(n_1885),
.B(n_1381),
.Y(n_2332)
);

INVx2_ASAP7_75t_L g2333 ( 
.A(n_1713),
.Y(n_2333)
);

INVx3_ASAP7_75t_L g2334 ( 
.A(n_1713),
.Y(n_2334)
);

INVx2_ASAP7_75t_L g2335 ( 
.A(n_1718),
.Y(n_2335)
);

INVx1_ASAP7_75t_L g2336 ( 
.A(n_1708),
.Y(n_2336)
);

NAND2xp5_ASAP7_75t_L g2337 ( 
.A(n_1888),
.B(n_1522),
.Y(n_2337)
);

INVx2_ASAP7_75t_SL g2338 ( 
.A(n_1694),
.Y(n_2338)
);

INVx2_ASAP7_75t_SL g2339 ( 
.A(n_1694),
.Y(n_2339)
);

INVx2_ASAP7_75t_L g2340 ( 
.A(n_1718),
.Y(n_2340)
);

INVx1_ASAP7_75t_L g2341 ( 
.A(n_1711),
.Y(n_2341)
);

AND2x6_ASAP7_75t_L g2342 ( 
.A(n_1781),
.B(n_1540),
.Y(n_2342)
);

INVx1_ASAP7_75t_L g2343 ( 
.A(n_1715),
.Y(n_2343)
);

INVx5_ASAP7_75t_L g2344 ( 
.A(n_1757),
.Y(n_2344)
);

INVxp67_ASAP7_75t_SL g2345 ( 
.A(n_1937),
.Y(n_2345)
);

INVx2_ASAP7_75t_L g2346 ( 
.A(n_1718),
.Y(n_2346)
);

INVx2_ASAP7_75t_SL g2347 ( 
.A(n_1720),
.Y(n_2347)
);

INVx2_ASAP7_75t_L g2348 ( 
.A(n_1722),
.Y(n_2348)
);

INVx2_ASAP7_75t_L g2349 ( 
.A(n_1722),
.Y(n_2349)
);

NAND2xp5_ASAP7_75t_L g2350 ( 
.A(n_1762),
.B(n_1578),
.Y(n_2350)
);

NAND2xp5_ASAP7_75t_SL g2351 ( 
.A(n_1770),
.B(n_1381),
.Y(n_2351)
);

INVx2_ASAP7_75t_L g2352 ( 
.A(n_1722),
.Y(n_2352)
);

NOR2xp33_ASAP7_75t_L g2353 ( 
.A(n_1783),
.B(n_1589),
.Y(n_2353)
);

NAND2xp5_ASAP7_75t_L g2354 ( 
.A(n_1763),
.B(n_1764),
.Y(n_2354)
);

INVx1_ASAP7_75t_L g2355 ( 
.A(n_1716),
.Y(n_2355)
);

CKINVDCx5p33_ASAP7_75t_R g2356 ( 
.A(n_1853),
.Y(n_2356)
);

NAND2xp33_ASAP7_75t_SL g2357 ( 
.A(n_1783),
.B(n_1553),
.Y(n_2357)
);

HB1xp67_ASAP7_75t_L g2358 ( 
.A(n_1890),
.Y(n_2358)
);

NAND2xp5_ASAP7_75t_SL g2359 ( 
.A(n_1910),
.B(n_1392),
.Y(n_2359)
);

INVx1_ASAP7_75t_L g2360 ( 
.A(n_1724),
.Y(n_2360)
);

INVxp67_ASAP7_75t_SL g2361 ( 
.A(n_1941),
.Y(n_2361)
);

NAND2xp5_ASAP7_75t_L g2362 ( 
.A(n_1659),
.B(n_1594),
.Y(n_2362)
);

INVx2_ASAP7_75t_L g2363 ( 
.A(n_1729),
.Y(n_2363)
);

INVx2_ASAP7_75t_L g2364 ( 
.A(n_1729),
.Y(n_2364)
);

INVx1_ASAP7_75t_L g2365 ( 
.A(n_1727),
.Y(n_2365)
);

INVx2_ASAP7_75t_L g2366 ( 
.A(n_1729),
.Y(n_2366)
);

INVx1_ASAP7_75t_L g2367 ( 
.A(n_1728),
.Y(n_2367)
);

HB1xp67_ASAP7_75t_L g2368 ( 
.A(n_1890),
.Y(n_2368)
);

INVx2_ASAP7_75t_L g2369 ( 
.A(n_1743),
.Y(n_2369)
);

NAND2xp5_ASAP7_75t_SL g2370 ( 
.A(n_1910),
.B(n_1392),
.Y(n_2370)
);

INVx2_ASAP7_75t_L g2371 ( 
.A(n_1743),
.Y(n_2371)
);

INVx2_ASAP7_75t_L g2372 ( 
.A(n_1743),
.Y(n_2372)
);

INVx3_ASAP7_75t_L g2373 ( 
.A(n_1766),
.Y(n_2373)
);

INVx3_ASAP7_75t_L g2374 ( 
.A(n_1766),
.Y(n_2374)
);

INVx2_ASAP7_75t_L g2375 ( 
.A(n_1766),
.Y(n_2375)
);

AND2x2_ASAP7_75t_L g2376 ( 
.A(n_1940),
.B(n_1619),
.Y(n_2376)
);

AND3x2_ASAP7_75t_L g2377 ( 
.A(n_1990),
.B(n_1473),
.C(n_1602),
.Y(n_2377)
);

AND2x2_ASAP7_75t_L g2378 ( 
.A(n_1940),
.B(n_1625),
.Y(n_2378)
);

NAND2xp5_ASAP7_75t_SL g2379 ( 
.A(n_1791),
.B(n_1633),
.Y(n_2379)
);

INVx1_ASAP7_75t_L g2380 ( 
.A(n_2056),
.Y(n_2380)
);

INVx1_ASAP7_75t_L g2381 ( 
.A(n_2056),
.Y(n_2381)
);

INVx1_ASAP7_75t_L g2382 ( 
.A(n_2062),
.Y(n_2382)
);

NAND2xp5_ASAP7_75t_L g2383 ( 
.A(n_2057),
.B(n_1732),
.Y(n_2383)
);

INVx2_ASAP7_75t_L g2384 ( 
.A(n_2036),
.Y(n_2384)
);

INVx1_ASAP7_75t_L g2385 ( 
.A(n_2062),
.Y(n_2385)
);

NAND2xp5_ASAP7_75t_L g2386 ( 
.A(n_2057),
.B(n_1661),
.Y(n_2386)
);

INVx1_ASAP7_75t_L g2387 ( 
.A(n_2063),
.Y(n_2387)
);

INVx1_ASAP7_75t_L g2388 ( 
.A(n_2063),
.Y(n_2388)
);

NOR2xp67_ASAP7_75t_L g2389 ( 
.A(n_2028),
.B(n_1525),
.Y(n_2389)
);

XOR2xp5_ASAP7_75t_L g2390 ( 
.A(n_2294),
.B(n_1795),
.Y(n_2390)
);

BUFx2_ASAP7_75t_L g2391 ( 
.A(n_2158),
.Y(n_2391)
);

XOR2xp5_ASAP7_75t_L g2392 ( 
.A(n_2294),
.B(n_1813),
.Y(n_2392)
);

INVx1_ASAP7_75t_L g2393 ( 
.A(n_2067),
.Y(n_2393)
);

AND2x2_ASAP7_75t_L g2394 ( 
.A(n_2149),
.B(n_1906),
.Y(n_2394)
);

NAND2xp5_ASAP7_75t_SL g2395 ( 
.A(n_2093),
.B(n_2059),
.Y(n_2395)
);

INVx2_ASAP7_75t_L g2396 ( 
.A(n_2036),
.Y(n_2396)
);

NOR2xp33_ASAP7_75t_L g2397 ( 
.A(n_2093),
.B(n_1746),
.Y(n_2397)
);

INVx1_ASAP7_75t_L g2398 ( 
.A(n_2067),
.Y(n_2398)
);

NAND2xp5_ASAP7_75t_L g2399 ( 
.A(n_2134),
.B(n_2257),
.Y(n_2399)
);

INVx1_ASAP7_75t_L g2400 ( 
.A(n_2069),
.Y(n_2400)
);

INVx1_ASAP7_75t_L g2401 ( 
.A(n_2069),
.Y(n_2401)
);

XOR2xp5_ASAP7_75t_L g2402 ( 
.A(n_2033),
.B(n_1813),
.Y(n_2402)
);

INVx1_ASAP7_75t_L g2403 ( 
.A(n_2071),
.Y(n_2403)
);

NOR2xp33_ASAP7_75t_L g2404 ( 
.A(n_2072),
.B(n_1746),
.Y(n_2404)
);

INVx2_ASAP7_75t_SL g2405 ( 
.A(n_2158),
.Y(n_2405)
);

NAND2x1p5_ASAP7_75t_L g2406 ( 
.A(n_2079),
.B(n_1873),
.Y(n_2406)
);

INVxp33_ASAP7_75t_L g2407 ( 
.A(n_2015),
.Y(n_2407)
);

NOR2xp33_ASAP7_75t_L g2408 ( 
.A(n_2023),
.B(n_1906),
.Y(n_2408)
);

INVx1_ASAP7_75t_L g2409 ( 
.A(n_2071),
.Y(n_2409)
);

INVx2_ASAP7_75t_L g2410 ( 
.A(n_2047),
.Y(n_2410)
);

NAND2xp33_ASAP7_75t_R g2411 ( 
.A(n_2202),
.B(n_2073),
.Y(n_2411)
);

INVx1_ASAP7_75t_L g2412 ( 
.A(n_2074),
.Y(n_2412)
);

AOI21xp5_ASAP7_75t_L g2413 ( 
.A1(n_2350),
.A2(n_1779),
.B(n_1769),
.Y(n_2413)
);

NAND2xp5_ASAP7_75t_L g2414 ( 
.A(n_2134),
.B(n_1785),
.Y(n_2414)
);

INVx1_ASAP7_75t_L g2415 ( 
.A(n_2074),
.Y(n_2415)
);

INVx1_ASAP7_75t_L g2416 ( 
.A(n_2077),
.Y(n_2416)
);

INVx2_ASAP7_75t_L g2417 ( 
.A(n_2047),
.Y(n_2417)
);

AND2x4_ASAP7_75t_L g2418 ( 
.A(n_2035),
.B(n_1874),
.Y(n_2418)
);

INVx1_ASAP7_75t_L g2419 ( 
.A(n_2077),
.Y(n_2419)
);

NAND2xp33_ASAP7_75t_R g2420 ( 
.A(n_2202),
.B(n_1993),
.Y(n_2420)
);

INVx1_ASAP7_75t_L g2421 ( 
.A(n_2085),
.Y(n_2421)
);

HB1xp67_ASAP7_75t_L g2422 ( 
.A(n_2248),
.Y(n_2422)
);

AND2x2_ASAP7_75t_L g2423 ( 
.A(n_2149),
.B(n_1924),
.Y(n_2423)
);

XOR2xp5_ASAP7_75t_L g2424 ( 
.A(n_2033),
.B(n_1993),
.Y(n_2424)
);

INVx1_ASAP7_75t_L g2425 ( 
.A(n_2085),
.Y(n_2425)
);

INVxp33_ASAP7_75t_L g2426 ( 
.A(n_2015),
.Y(n_2426)
);

INVx1_ASAP7_75t_L g2427 ( 
.A(n_2104),
.Y(n_2427)
);

NAND2xp5_ASAP7_75t_SL g2428 ( 
.A(n_2213),
.B(n_1901),
.Y(n_2428)
);

INVx2_ASAP7_75t_L g2429 ( 
.A(n_2048),
.Y(n_2429)
);

INVx1_ASAP7_75t_L g2430 ( 
.A(n_2104),
.Y(n_2430)
);

INVx1_ASAP7_75t_L g2431 ( 
.A(n_2105),
.Y(n_2431)
);

INVx1_ASAP7_75t_L g2432 ( 
.A(n_2105),
.Y(n_2432)
);

INVxp67_ASAP7_75t_SL g2433 ( 
.A(n_2027),
.Y(n_2433)
);

INVx1_ASAP7_75t_L g2434 ( 
.A(n_2107),
.Y(n_2434)
);

INVx1_ASAP7_75t_L g2435 ( 
.A(n_2107),
.Y(n_2435)
);

INVx1_ASAP7_75t_L g2436 ( 
.A(n_2110),
.Y(n_2436)
);

NAND2xp5_ASAP7_75t_L g2437 ( 
.A(n_2257),
.B(n_1792),
.Y(n_2437)
);

INVx1_ASAP7_75t_L g2438 ( 
.A(n_2110),
.Y(n_2438)
);

INVx1_ASAP7_75t_L g2439 ( 
.A(n_2139),
.Y(n_2439)
);

AND2x2_ASAP7_75t_L g2440 ( 
.A(n_2204),
.B(n_1924),
.Y(n_2440)
);

INVx1_ASAP7_75t_L g2441 ( 
.A(n_2139),
.Y(n_2441)
);

CKINVDCx5p33_ASAP7_75t_R g2442 ( 
.A(n_2356),
.Y(n_2442)
);

AOI21xp5_ASAP7_75t_L g2443 ( 
.A1(n_2350),
.A2(n_2020),
.B(n_2017),
.Y(n_2443)
);

BUFx3_ASAP7_75t_L g2444 ( 
.A(n_2248),
.Y(n_2444)
);

AND2x4_ASAP7_75t_L g2445 ( 
.A(n_2035),
.B(n_1881),
.Y(n_2445)
);

INVx4_ASAP7_75t_SL g2446 ( 
.A(n_2079),
.Y(n_2446)
);

XOR2xp5_ASAP7_75t_L g2447 ( 
.A(n_2356),
.B(n_1055),
.Y(n_2447)
);

NOR2xp33_ASAP7_75t_L g2448 ( 
.A(n_2054),
.B(n_1922),
.Y(n_2448)
);

INVx1_ASAP7_75t_L g2449 ( 
.A(n_2142),
.Y(n_2449)
);

AND2x2_ASAP7_75t_L g2450 ( 
.A(n_2204),
.B(n_1638),
.Y(n_2450)
);

INVx1_ASAP7_75t_L g2451 ( 
.A(n_2142),
.Y(n_2451)
);

NOR2xp33_ASAP7_75t_L g2452 ( 
.A(n_2087),
.B(n_1922),
.Y(n_2452)
);

NOR2xp33_ASAP7_75t_SL g2453 ( 
.A(n_2018),
.B(n_1959),
.Y(n_2453)
);

XNOR2xp5_ASAP7_75t_L g2454 ( 
.A(n_2289),
.B(n_1055),
.Y(n_2454)
);

INVx1_ASAP7_75t_L g2455 ( 
.A(n_2120),
.Y(n_2455)
);

NOR2xp33_ASAP7_75t_L g2456 ( 
.A(n_2108),
.B(n_1932),
.Y(n_2456)
);

INVx3_ASAP7_75t_L g2457 ( 
.A(n_2313),
.Y(n_2457)
);

INVx1_ASAP7_75t_L g2458 ( 
.A(n_2120),
.Y(n_2458)
);

AND2x2_ASAP7_75t_L g2459 ( 
.A(n_2070),
.B(n_1625),
.Y(n_2459)
);

INVx1_ASAP7_75t_L g2460 ( 
.A(n_2123),
.Y(n_2460)
);

INVx1_ASAP7_75t_L g2461 ( 
.A(n_2123),
.Y(n_2461)
);

INVx1_ASAP7_75t_L g2462 ( 
.A(n_2128),
.Y(n_2462)
);

INVx1_ASAP7_75t_L g2463 ( 
.A(n_2128),
.Y(n_2463)
);

INVx2_ASAP7_75t_L g2464 ( 
.A(n_2048),
.Y(n_2464)
);

CKINVDCx20_ASAP7_75t_R g2465 ( 
.A(n_2169),
.Y(n_2465)
);

INVx1_ASAP7_75t_L g2466 ( 
.A(n_2129),
.Y(n_2466)
);

AND2x2_ASAP7_75t_L g2467 ( 
.A(n_2070),
.B(n_1932),
.Y(n_2467)
);

CKINVDCx20_ASAP7_75t_R g2468 ( 
.A(n_2169),
.Y(n_2468)
);

INVx1_ASAP7_75t_L g2469 ( 
.A(n_2129),
.Y(n_2469)
);

INVx1_ASAP7_75t_L g2470 ( 
.A(n_2133),
.Y(n_2470)
);

INVx1_ASAP7_75t_L g2471 ( 
.A(n_2133),
.Y(n_2471)
);

INVx4_ASAP7_75t_SL g2472 ( 
.A(n_2079),
.Y(n_2472)
);

INVx1_ASAP7_75t_L g2473 ( 
.A(n_2135),
.Y(n_2473)
);

NOR2x1_ASAP7_75t_L g2474 ( 
.A(n_2028),
.B(n_1791),
.Y(n_2474)
);

INVx1_ASAP7_75t_L g2475 ( 
.A(n_2135),
.Y(n_2475)
);

NOR2xp67_ASAP7_75t_L g2476 ( 
.A(n_2220),
.B(n_1339),
.Y(n_2476)
);

INVx2_ASAP7_75t_L g2477 ( 
.A(n_2050),
.Y(n_2477)
);

NAND2xp33_ASAP7_75t_SL g2478 ( 
.A(n_2080),
.B(n_1823),
.Y(n_2478)
);

INVxp67_ASAP7_75t_L g2479 ( 
.A(n_2065),
.Y(n_2479)
);

BUFx2_ASAP7_75t_L g2480 ( 
.A(n_2238),
.Y(n_2480)
);

INVx2_ASAP7_75t_L g2481 ( 
.A(n_2050),
.Y(n_2481)
);

INVx1_ASAP7_75t_L g2482 ( 
.A(n_2272),
.Y(n_2482)
);

CKINVDCx20_ASAP7_75t_R g2483 ( 
.A(n_2238),
.Y(n_2483)
);

INVx2_ASAP7_75t_SL g2484 ( 
.A(n_2259),
.Y(n_2484)
);

INVx1_ASAP7_75t_L g2485 ( 
.A(n_2272),
.Y(n_2485)
);

CKINVDCx16_ASAP7_75t_R g2486 ( 
.A(n_2325),
.Y(n_2486)
);

INVx1_ASAP7_75t_L g2487 ( 
.A(n_2119),
.Y(n_2487)
);

INVx2_ASAP7_75t_L g2488 ( 
.A(n_2053),
.Y(n_2488)
);

INVx1_ASAP7_75t_L g2489 ( 
.A(n_2119),
.Y(n_2489)
);

INVx1_ASAP7_75t_L g2490 ( 
.A(n_2124),
.Y(n_2490)
);

NAND2xp5_ASAP7_75t_L g2491 ( 
.A(n_2121),
.B(n_1799),
.Y(n_2491)
);

INVx2_ASAP7_75t_L g2492 ( 
.A(n_2053),
.Y(n_2492)
);

CKINVDCx5p33_ASAP7_75t_R g2493 ( 
.A(n_2116),
.Y(n_2493)
);

INVx1_ASAP7_75t_L g2494 ( 
.A(n_2124),
.Y(n_2494)
);

INVx1_ASAP7_75t_L g2495 ( 
.A(n_2125),
.Y(n_2495)
);

INVx1_ASAP7_75t_L g2496 ( 
.A(n_2125),
.Y(n_2496)
);

INVxp33_ASAP7_75t_L g2497 ( 
.A(n_2068),
.Y(n_2497)
);

AND2x2_ASAP7_75t_L g2498 ( 
.A(n_2094),
.B(n_1433),
.Y(n_2498)
);

INVx1_ASAP7_75t_L g2499 ( 
.A(n_2138),
.Y(n_2499)
);

NAND2xp5_ASAP7_75t_L g2500 ( 
.A(n_2121),
.B(n_1801),
.Y(n_2500)
);

INVx1_ASAP7_75t_L g2501 ( 
.A(n_2138),
.Y(n_2501)
);

NOR2xp67_ASAP7_75t_L g2502 ( 
.A(n_2220),
.B(n_1440),
.Y(n_2502)
);

INVx1_ASAP7_75t_L g2503 ( 
.A(n_2261),
.Y(n_2503)
);

NOR2xp33_ASAP7_75t_L g2504 ( 
.A(n_2167),
.B(n_1823),
.Y(n_2504)
);

NAND2xp33_ASAP7_75t_R g2505 ( 
.A(n_2233),
.B(n_1950),
.Y(n_2505)
);

NOR2xp33_ASAP7_75t_L g2506 ( 
.A(n_2184),
.B(n_1858),
.Y(n_2506)
);

INVx1_ASAP7_75t_L g2507 ( 
.A(n_2261),
.Y(n_2507)
);

CKINVDCx20_ASAP7_75t_R g2508 ( 
.A(n_2098),
.Y(n_2508)
);

INVx3_ASAP7_75t_R g2509 ( 
.A(n_2068),
.Y(n_2509)
);

INVx1_ASAP7_75t_L g2510 ( 
.A(n_2268),
.Y(n_2510)
);

INVx1_ASAP7_75t_L g2511 ( 
.A(n_2268),
.Y(n_2511)
);

INVx1_ASAP7_75t_L g2512 ( 
.A(n_2276),
.Y(n_2512)
);

AOI21xp5_ASAP7_75t_L g2513 ( 
.A1(n_2017),
.A2(n_2029),
.B(n_2020),
.Y(n_2513)
);

XNOR2x2_ASAP7_75t_L g2514 ( 
.A(n_2259),
.B(n_563),
.Y(n_2514)
);

INVx2_ASAP7_75t_SL g2515 ( 
.A(n_2358),
.Y(n_2515)
);

INVxp33_ASAP7_75t_SL g2516 ( 
.A(n_2325),
.Y(n_2516)
);

NOR2xp33_ASAP7_75t_L g2517 ( 
.A(n_2283),
.B(n_1926),
.Y(n_2517)
);

INVx2_ASAP7_75t_L g2518 ( 
.A(n_2058),
.Y(n_2518)
);

XOR2xp5_ASAP7_75t_L g2519 ( 
.A(n_2269),
.B(n_1074),
.Y(n_2519)
);

INVxp67_ASAP7_75t_SL g2520 ( 
.A(n_2027),
.Y(n_2520)
);

INVx1_ASAP7_75t_L g2521 ( 
.A(n_2276),
.Y(n_2521)
);

NAND2x1p5_ASAP7_75t_L g2522 ( 
.A(n_2079),
.B(n_1883),
.Y(n_2522)
);

AND2x2_ASAP7_75t_L g2523 ( 
.A(n_2094),
.B(n_1437),
.Y(n_2523)
);

CKINVDCx20_ASAP7_75t_R g2524 ( 
.A(n_2252),
.Y(n_2524)
);

NOR2xp33_ASAP7_75t_L g2525 ( 
.A(n_2283),
.B(n_1926),
.Y(n_2525)
);

INVx1_ASAP7_75t_L g2526 ( 
.A(n_2281),
.Y(n_2526)
);

INVx1_ASAP7_75t_L g2527 ( 
.A(n_2281),
.Y(n_2527)
);

INVx1_ASAP7_75t_L g2528 ( 
.A(n_2284),
.Y(n_2528)
);

XNOR2x2_ASAP7_75t_L g2529 ( 
.A(n_2208),
.B(n_2217),
.Y(n_2529)
);

INVx1_ASAP7_75t_L g2530 ( 
.A(n_2284),
.Y(n_2530)
);

INVx1_ASAP7_75t_L g2531 ( 
.A(n_2288),
.Y(n_2531)
);

INVx3_ASAP7_75t_L g2532 ( 
.A(n_2313),
.Y(n_2532)
);

INVx1_ASAP7_75t_L g2533 ( 
.A(n_2288),
.Y(n_2533)
);

INVxp67_ASAP7_75t_L g2534 ( 
.A(n_2368),
.Y(n_2534)
);

INVx1_ASAP7_75t_L g2535 ( 
.A(n_2291),
.Y(n_2535)
);

NOR2xp33_ASAP7_75t_L g2536 ( 
.A(n_2286),
.B(n_1926),
.Y(n_2536)
);

INVx1_ASAP7_75t_L g2537 ( 
.A(n_2291),
.Y(n_2537)
);

INVx1_ASAP7_75t_L g2538 ( 
.A(n_2315),
.Y(n_2538)
);

INVx1_ASAP7_75t_L g2539 ( 
.A(n_2315),
.Y(n_2539)
);

INVxp67_ASAP7_75t_SL g2540 ( 
.A(n_2027),
.Y(n_2540)
);

INVx1_ASAP7_75t_L g2541 ( 
.A(n_2323),
.Y(n_2541)
);

AND2x2_ASAP7_75t_L g2542 ( 
.A(n_2055),
.B(n_2090),
.Y(n_2542)
);

INVx1_ASAP7_75t_L g2543 ( 
.A(n_2323),
.Y(n_2543)
);

NOR2xp33_ASAP7_75t_L g2544 ( 
.A(n_2286),
.B(n_1886),
.Y(n_2544)
);

AND2x2_ASAP7_75t_L g2545 ( 
.A(n_2055),
.B(n_1461),
.Y(n_2545)
);

INVx1_ASAP7_75t_L g2546 ( 
.A(n_2327),
.Y(n_2546)
);

BUFx3_ASAP7_75t_L g2547 ( 
.A(n_2176),
.Y(n_2547)
);

NOR2xp33_ASAP7_75t_L g2548 ( 
.A(n_2237),
.B(n_1889),
.Y(n_2548)
);

XOR2xp5_ASAP7_75t_L g2549 ( 
.A(n_2293),
.B(n_1074),
.Y(n_2549)
);

NAND2xp33_ASAP7_75t_SL g2550 ( 
.A(n_2080),
.B(n_1495),
.Y(n_2550)
);

INVx1_ASAP7_75t_L g2551 ( 
.A(n_2327),
.Y(n_2551)
);

CKINVDCx5p33_ASAP7_75t_R g2552 ( 
.A(n_2116),
.Y(n_2552)
);

INVx1_ASAP7_75t_L g2553 ( 
.A(n_2336),
.Y(n_2553)
);

INVx1_ASAP7_75t_L g2554 ( 
.A(n_2336),
.Y(n_2554)
);

NAND2xp5_ASAP7_75t_L g2555 ( 
.A(n_2171),
.B(n_1802),
.Y(n_2555)
);

BUFx3_ASAP7_75t_L g2556 ( 
.A(n_2176),
.Y(n_2556)
);

INVx1_ASAP7_75t_L g2557 ( 
.A(n_2341),
.Y(n_2557)
);

NOR2xp33_ASAP7_75t_L g2558 ( 
.A(n_2155),
.B(n_1893),
.Y(n_2558)
);

INVx1_ASAP7_75t_L g2559 ( 
.A(n_2341),
.Y(n_2559)
);

AND2x2_ASAP7_75t_L g2560 ( 
.A(n_2090),
.B(n_1468),
.Y(n_2560)
);

INVx1_ASAP7_75t_L g2561 ( 
.A(n_2343),
.Y(n_2561)
);

AND2x2_ASAP7_75t_L g2562 ( 
.A(n_2060),
.B(n_1468),
.Y(n_2562)
);

NOR2xp33_ASAP7_75t_L g2563 ( 
.A(n_2151),
.B(n_1904),
.Y(n_2563)
);

INVx1_ASAP7_75t_L g2564 ( 
.A(n_2343),
.Y(n_2564)
);

AND2x2_ASAP7_75t_L g2565 ( 
.A(n_2182),
.B(n_1469),
.Y(n_2565)
);

AND2x2_ASAP7_75t_L g2566 ( 
.A(n_2182),
.B(n_2101),
.Y(n_2566)
);

INVx1_ASAP7_75t_L g2567 ( 
.A(n_2355),
.Y(n_2567)
);

INVx1_ASAP7_75t_L g2568 ( 
.A(n_2355),
.Y(n_2568)
);

NAND2xp5_ASAP7_75t_SL g2569 ( 
.A(n_2122),
.B(n_2314),
.Y(n_2569)
);

AND2x2_ASAP7_75t_L g2570 ( 
.A(n_2101),
.B(n_1469),
.Y(n_2570)
);

OR2x2_ASAP7_75t_L g2571 ( 
.A(n_2233),
.B(n_1908),
.Y(n_2571)
);

INVxp67_ASAP7_75t_SL g2572 ( 
.A(n_2027),
.Y(n_2572)
);

INVx2_ASAP7_75t_SL g2573 ( 
.A(n_2131),
.Y(n_2573)
);

INVx1_ASAP7_75t_L g2574 ( 
.A(n_2360),
.Y(n_2574)
);

INVx1_ASAP7_75t_L g2575 ( 
.A(n_2360),
.Y(n_2575)
);

CKINVDCx20_ASAP7_75t_R g2576 ( 
.A(n_2357),
.Y(n_2576)
);

NAND2xp5_ASAP7_75t_SL g2577 ( 
.A(n_2122),
.B(n_1913),
.Y(n_2577)
);

INVx1_ASAP7_75t_L g2578 ( 
.A(n_2365),
.Y(n_2578)
);

INVx1_ASAP7_75t_L g2579 ( 
.A(n_2365),
.Y(n_2579)
);

NAND2xp33_ASAP7_75t_SL g2580 ( 
.A(n_2080),
.B(n_1915),
.Y(n_2580)
);

NOR2xp33_ASAP7_75t_L g2581 ( 
.A(n_2122),
.B(n_1917),
.Y(n_2581)
);

INVx2_ASAP7_75t_L g2582 ( 
.A(n_2058),
.Y(n_2582)
);

INVx1_ASAP7_75t_L g2583 ( 
.A(n_2367),
.Y(n_2583)
);

XNOR2xp5_ASAP7_75t_L g2584 ( 
.A(n_2377),
.B(n_1089),
.Y(n_2584)
);

INVx1_ASAP7_75t_L g2585 ( 
.A(n_2367),
.Y(n_2585)
);

INVx1_ASAP7_75t_L g2586 ( 
.A(n_2255),
.Y(n_2586)
);

CKINVDCx20_ASAP7_75t_R g2587 ( 
.A(n_2130),
.Y(n_2587)
);

AND2x2_ASAP7_75t_L g2588 ( 
.A(n_2173),
.B(n_1481),
.Y(n_2588)
);

INVx2_ASAP7_75t_L g2589 ( 
.A(n_2064),
.Y(n_2589)
);

INVx1_ASAP7_75t_L g2590 ( 
.A(n_2255),
.Y(n_2590)
);

INVx2_ASAP7_75t_SL g2591 ( 
.A(n_2131),
.Y(n_2591)
);

NOR2xp33_ASAP7_75t_L g2592 ( 
.A(n_2314),
.B(n_2280),
.Y(n_2592)
);

XNOR2x2_ASAP7_75t_L g2593 ( 
.A(n_2208),
.B(n_576),
.Y(n_2593)
);

XOR2xp5_ASAP7_75t_L g2594 ( 
.A(n_2061),
.B(n_1089),
.Y(n_2594)
);

NOR2xp33_ASAP7_75t_L g2595 ( 
.A(n_2018),
.B(n_1918),
.Y(n_2595)
);

INVx1_ASAP7_75t_L g2596 ( 
.A(n_2264),
.Y(n_2596)
);

INVx1_ASAP7_75t_L g2597 ( 
.A(n_2264),
.Y(n_2597)
);

INVx1_ASAP7_75t_L g2598 ( 
.A(n_2064),
.Y(n_2598)
);

INVx1_ASAP7_75t_L g2599 ( 
.A(n_2066),
.Y(n_2599)
);

INVx1_ASAP7_75t_L g2600 ( 
.A(n_2066),
.Y(n_2600)
);

XNOR2xp5_ASAP7_75t_SL g2601 ( 
.A(n_2180),
.B(n_1608),
.Y(n_2601)
);

AND2x4_ASAP7_75t_L g2602 ( 
.A(n_2035),
.B(n_2051),
.Y(n_2602)
);

INVx1_ASAP7_75t_L g2603 ( 
.A(n_2075),
.Y(n_2603)
);

INVx1_ASAP7_75t_L g2604 ( 
.A(n_2075),
.Y(n_2604)
);

INVx1_ASAP7_75t_L g2605 ( 
.A(n_2082),
.Y(n_2605)
);

AND2x2_ASAP7_75t_L g2606 ( 
.A(n_2109),
.B(n_1481),
.Y(n_2606)
);

AND2x2_ASAP7_75t_L g2607 ( 
.A(n_2109),
.B(n_1486),
.Y(n_2607)
);

XOR2x2_ASAP7_75t_L g2608 ( 
.A(n_2246),
.B(n_1612),
.Y(n_2608)
);

INVx2_ASAP7_75t_L g2609 ( 
.A(n_2082),
.Y(n_2609)
);

INVx1_ASAP7_75t_L g2610 ( 
.A(n_2088),
.Y(n_2610)
);

OAI21xp5_ASAP7_75t_L g2611 ( 
.A1(n_2043),
.A2(n_1808),
.B(n_1805),
.Y(n_2611)
);

INVx1_ASAP7_75t_L g2612 ( 
.A(n_2088),
.Y(n_2612)
);

INVx1_ASAP7_75t_L g2613 ( 
.A(n_2092),
.Y(n_2613)
);

INVx1_ASAP7_75t_L g2614 ( 
.A(n_2092),
.Y(n_2614)
);

INVx1_ASAP7_75t_L g2615 ( 
.A(n_2096),
.Y(n_2615)
);

NAND2xp5_ASAP7_75t_L g2616 ( 
.A(n_2118),
.B(n_1811),
.Y(n_2616)
);

INVx1_ASAP7_75t_L g2617 ( 
.A(n_2096),
.Y(n_2617)
);

INVx4_ASAP7_75t_L g2618 ( 
.A(n_2299),
.Y(n_2618)
);

CKINVDCx14_ASAP7_75t_R g2619 ( 
.A(n_2160),
.Y(n_2619)
);

INVx1_ASAP7_75t_L g2620 ( 
.A(n_2099),
.Y(n_2620)
);

INVx1_ASAP7_75t_L g2621 ( 
.A(n_2099),
.Y(n_2621)
);

AND2x2_ASAP7_75t_L g2622 ( 
.A(n_2265),
.B(n_1486),
.Y(n_2622)
);

INVx1_ASAP7_75t_L g2623 ( 
.A(n_2102),
.Y(n_2623)
);

AND2x2_ASAP7_75t_SL g2624 ( 
.A(n_2226),
.B(n_1720),
.Y(n_2624)
);

XOR2xp5_ASAP7_75t_L g2625 ( 
.A(n_2197),
.B(n_1094),
.Y(n_2625)
);

INVx1_ASAP7_75t_L g2626 ( 
.A(n_2102),
.Y(n_2626)
);

AND2x4_ASAP7_75t_L g2627 ( 
.A(n_2051),
.B(n_1919),
.Y(n_2627)
);

INVxp33_ASAP7_75t_L g2628 ( 
.A(n_2160),
.Y(n_2628)
);

NAND2xp5_ASAP7_75t_L g2629 ( 
.A(n_2309),
.B(n_1814),
.Y(n_2629)
);

AND2x6_ASAP7_75t_L g2630 ( 
.A(n_2043),
.B(n_1720),
.Y(n_2630)
);

INVx1_ASAP7_75t_L g2631 ( 
.A(n_2103),
.Y(n_2631)
);

INVx1_ASAP7_75t_L g2632 ( 
.A(n_2103),
.Y(n_2632)
);

BUFx5_ASAP7_75t_L g2633 ( 
.A(n_2045),
.Y(n_2633)
);

INVx1_ASAP7_75t_L g2634 ( 
.A(n_2106),
.Y(n_2634)
);

INVx1_ASAP7_75t_L g2635 ( 
.A(n_2106),
.Y(n_2635)
);

AND2x4_ASAP7_75t_L g2636 ( 
.A(n_2051),
.B(n_1920),
.Y(n_2636)
);

AND2x2_ASAP7_75t_L g2637 ( 
.A(n_2265),
.B(n_1730),
.Y(n_2637)
);

INVx1_ASAP7_75t_L g2638 ( 
.A(n_2111),
.Y(n_2638)
);

INVx1_ASAP7_75t_SL g2639 ( 
.A(n_2232),
.Y(n_2639)
);

INVx1_ASAP7_75t_L g2640 ( 
.A(n_2111),
.Y(n_2640)
);

INVx2_ASAP7_75t_SL g2641 ( 
.A(n_2232),
.Y(n_2641)
);

INVx1_ASAP7_75t_L g2642 ( 
.A(n_2114),
.Y(n_2642)
);

NAND2xp33_ASAP7_75t_R g2643 ( 
.A(n_2235),
.B(n_1950),
.Y(n_2643)
);

NOR2xp33_ASAP7_75t_L g2644 ( 
.A(n_2018),
.B(n_1512),
.Y(n_2644)
);

CKINVDCx20_ASAP7_75t_R g2645 ( 
.A(n_2130),
.Y(n_2645)
);

INVx2_ASAP7_75t_L g2646 ( 
.A(n_2114),
.Y(n_2646)
);

INVx1_ASAP7_75t_L g2647 ( 
.A(n_2117),
.Y(n_2647)
);

INVx1_ASAP7_75t_L g2648 ( 
.A(n_2117),
.Y(n_2648)
);

INVx1_ASAP7_75t_L g2649 ( 
.A(n_2147),
.Y(n_2649)
);

NOR2xp33_ASAP7_75t_L g2650 ( 
.A(n_2018),
.B(n_1512),
.Y(n_2650)
);

CKINVDCx20_ASAP7_75t_R g2651 ( 
.A(n_2221),
.Y(n_2651)
);

INVx1_ASAP7_75t_L g2652 ( 
.A(n_2147),
.Y(n_2652)
);

INVx1_ASAP7_75t_L g2653 ( 
.A(n_2156),
.Y(n_2653)
);

AND2x4_ASAP7_75t_L g2654 ( 
.A(n_2176),
.B(n_1730),
.Y(n_2654)
);

INVx1_ASAP7_75t_L g2655 ( 
.A(n_2156),
.Y(n_2655)
);

BUFx6f_ASAP7_75t_L g2656 ( 
.A(n_2311),
.Y(n_2656)
);

NOR2xp33_ASAP7_75t_L g2657 ( 
.A(n_2078),
.B(n_1559),
.Y(n_2657)
);

INVx1_ASAP7_75t_L g2658 ( 
.A(n_2161),
.Y(n_2658)
);

INVx1_ASAP7_75t_L g2659 ( 
.A(n_2161),
.Y(n_2659)
);

INVx1_ASAP7_75t_L g2660 ( 
.A(n_2166),
.Y(n_2660)
);

INVx1_ASAP7_75t_L g2661 ( 
.A(n_2166),
.Y(n_2661)
);

INVx1_ASAP7_75t_L g2662 ( 
.A(n_2267),
.Y(n_2662)
);

INVx1_ASAP7_75t_L g2663 ( 
.A(n_2267),
.Y(n_2663)
);

NOR2xp33_ASAP7_75t_L g2664 ( 
.A(n_2337),
.B(n_1559),
.Y(n_2664)
);

XNOR2x2_ASAP7_75t_SL g2665 ( 
.A(n_2235),
.B(n_1094),
.Y(n_2665)
);

INVx1_ASAP7_75t_L g2666 ( 
.A(n_2183),
.Y(n_2666)
);

NOR2xp33_ASAP7_75t_L g2667 ( 
.A(n_2052),
.B(n_1561),
.Y(n_2667)
);

INVx1_ASAP7_75t_L g2668 ( 
.A(n_2183),
.Y(n_2668)
);

INVx1_ASAP7_75t_L g2669 ( 
.A(n_2185),
.Y(n_2669)
);

INVx1_ASAP7_75t_L g2670 ( 
.A(n_2185),
.Y(n_2670)
);

AND2x4_ASAP7_75t_L g2671 ( 
.A(n_2176),
.B(n_1730),
.Y(n_2671)
);

XOR2xp5_ASAP7_75t_L g2672 ( 
.A(n_2239),
.B(n_1145),
.Y(n_2672)
);

NAND2xp33_ASAP7_75t_R g2673 ( 
.A(n_2251),
.B(n_1735),
.Y(n_2673)
);

INVx1_ASAP7_75t_L g2674 ( 
.A(n_2187),
.Y(n_2674)
);

INVx1_ASAP7_75t_L g2675 ( 
.A(n_2187),
.Y(n_2675)
);

INVx1_ASAP7_75t_L g2676 ( 
.A(n_2191),
.Y(n_2676)
);

INVx1_ASAP7_75t_L g2677 ( 
.A(n_2191),
.Y(n_2677)
);

INVx1_ASAP7_75t_L g2678 ( 
.A(n_2193),
.Y(n_2678)
);

XNOR2xp5_ASAP7_75t_L g2679 ( 
.A(n_2112),
.B(n_1145),
.Y(n_2679)
);

NOR2xp33_ASAP7_75t_L g2680 ( 
.A(n_2052),
.B(n_1561),
.Y(n_2680)
);

INVxp33_ASAP7_75t_SL g2681 ( 
.A(n_2318),
.Y(n_2681)
);

AND2x4_ASAP7_75t_L g2682 ( 
.A(n_2042),
.B(n_1735),
.Y(n_2682)
);

INVx1_ASAP7_75t_L g2683 ( 
.A(n_2193),
.Y(n_2683)
);

INVx1_ASAP7_75t_L g2684 ( 
.A(n_2194),
.Y(n_2684)
);

AND2x2_ASAP7_75t_L g2685 ( 
.A(n_2251),
.B(n_1735),
.Y(n_2685)
);

AND2x2_ASAP7_75t_L g2686 ( 
.A(n_2231),
.B(n_1736),
.Y(n_2686)
);

NOR2xp33_ASAP7_75t_L g2687 ( 
.A(n_2321),
.B(n_1580),
.Y(n_2687)
);

INVx2_ASAP7_75t_L g2688 ( 
.A(n_2081),
.Y(n_2688)
);

NAND2xp33_ASAP7_75t_R g2689 ( 
.A(n_2295),
.B(n_1736),
.Y(n_2689)
);

XNOR2xp5_ASAP7_75t_L g2690 ( 
.A(n_2112),
.B(n_1172),
.Y(n_2690)
);

NOR2xp33_ASAP7_75t_L g2691 ( 
.A(n_2321),
.B(n_1580),
.Y(n_2691)
);

INVx1_ASAP7_75t_L g2692 ( 
.A(n_2194),
.Y(n_2692)
);

CKINVDCx20_ASAP7_75t_R g2693 ( 
.A(n_2221),
.Y(n_2693)
);

INVx1_ASAP7_75t_L g2694 ( 
.A(n_2195),
.Y(n_2694)
);

INVx1_ASAP7_75t_L g2695 ( 
.A(n_2195),
.Y(n_2695)
);

INVx1_ASAP7_75t_L g2696 ( 
.A(n_2199),
.Y(n_2696)
);

NOR2xp67_ASAP7_75t_L g2697 ( 
.A(n_2095),
.B(n_1444),
.Y(n_2697)
);

INVx2_ASAP7_75t_SL g2698 ( 
.A(n_2231),
.Y(n_2698)
);

INVx1_ASAP7_75t_L g2699 ( 
.A(n_2199),
.Y(n_2699)
);

CKINVDCx16_ASAP7_75t_R g2700 ( 
.A(n_2221),
.Y(n_2700)
);

INVx1_ASAP7_75t_L g2701 ( 
.A(n_2200),
.Y(n_2701)
);

INVx1_ASAP7_75t_L g2702 ( 
.A(n_2200),
.Y(n_2702)
);

BUFx3_ASAP7_75t_L g2703 ( 
.A(n_2316),
.Y(n_2703)
);

INVx1_ASAP7_75t_L g2704 ( 
.A(n_2223),
.Y(n_2704)
);

INVx1_ASAP7_75t_L g2705 ( 
.A(n_2223),
.Y(n_2705)
);

XOR2xp5_ASAP7_75t_L g2706 ( 
.A(n_2243),
.B(n_1172),
.Y(n_2706)
);

INVx1_ASAP7_75t_L g2707 ( 
.A(n_2225),
.Y(n_2707)
);

INVxp33_ASAP7_75t_L g2708 ( 
.A(n_2353),
.Y(n_2708)
);

INVxp33_ASAP7_75t_L g2709 ( 
.A(n_2154),
.Y(n_2709)
);

INVx1_ASAP7_75t_L g2710 ( 
.A(n_2225),
.Y(n_2710)
);

INVxp33_ASAP7_75t_L g2711 ( 
.A(n_2163),
.Y(n_2711)
);

CKINVDCx20_ASAP7_75t_R g2712 ( 
.A(n_2221),
.Y(n_2712)
);

AND2x2_ASAP7_75t_L g2713 ( 
.A(n_2376),
.B(n_1736),
.Y(n_2713)
);

AND2x2_ASAP7_75t_L g2714 ( 
.A(n_2376),
.B(n_1749),
.Y(n_2714)
);

INVx1_ASAP7_75t_L g2715 ( 
.A(n_2227),
.Y(n_2715)
);

INVxp33_ASAP7_75t_L g2716 ( 
.A(n_2218),
.Y(n_2716)
);

INVx2_ASAP7_75t_L g2717 ( 
.A(n_2081),
.Y(n_2717)
);

CKINVDCx5p33_ASAP7_75t_R g2718 ( 
.A(n_2249),
.Y(n_2718)
);

INVx1_ASAP7_75t_L g2719 ( 
.A(n_2227),
.Y(n_2719)
);

INVx5_ASAP7_75t_L g2720 ( 
.A(n_2079),
.Y(n_2720)
);

INVx1_ASAP7_75t_L g2721 ( 
.A(n_2230),
.Y(n_2721)
);

INVx1_ASAP7_75t_L g2722 ( 
.A(n_2230),
.Y(n_2722)
);

AOI22xp33_ASAP7_75t_L g2723 ( 
.A1(n_2448),
.A2(n_2089),
.B1(n_2097),
.B2(n_2378),
.Y(n_2723)
);

INVx1_ASAP7_75t_L g2724 ( 
.A(n_2380),
.Y(n_2724)
);

INVx1_ASAP7_75t_SL g2725 ( 
.A(n_2480),
.Y(n_2725)
);

INVx2_ASAP7_75t_L g2726 ( 
.A(n_2384),
.Y(n_2726)
);

AOI22xp5_ASAP7_75t_L g2727 ( 
.A1(n_2448),
.A2(n_2452),
.B1(n_2504),
.B2(n_2428),
.Y(n_2727)
);

AOI22xp5_ASAP7_75t_L g2728 ( 
.A1(n_2452),
.A2(n_2379),
.B1(n_2046),
.B2(n_2083),
.Y(n_2728)
);

NAND2xp33_ASAP7_75t_L g2729 ( 
.A(n_2399),
.B(n_2342),
.Y(n_2729)
);

NAND2xp5_ASAP7_75t_L g2730 ( 
.A(n_2399),
.B(n_2378),
.Y(n_2730)
);

NAND2xp5_ASAP7_75t_SL g2731 ( 
.A(n_2681),
.B(n_2504),
.Y(n_2731)
);

INVx1_ASAP7_75t_L g2732 ( 
.A(n_2381),
.Y(n_2732)
);

INVx2_ASAP7_75t_L g2733 ( 
.A(n_2396),
.Y(n_2733)
);

INVx1_ASAP7_75t_SL g2734 ( 
.A(n_2483),
.Y(n_2734)
);

NAND2xp5_ASAP7_75t_SL g2735 ( 
.A(n_2592),
.B(n_2249),
.Y(n_2735)
);

NOR2xp33_ASAP7_75t_L g2736 ( 
.A(n_2708),
.B(n_1190),
.Y(n_2736)
);

INVx2_ASAP7_75t_L g2737 ( 
.A(n_2410),
.Y(n_2737)
);

NOR3xp33_ASAP7_75t_L g2738 ( 
.A(n_2687),
.B(n_2145),
.C(n_2146),
.Y(n_2738)
);

BUFx3_ASAP7_75t_L g2739 ( 
.A(n_2444),
.Y(n_2739)
);

INVx1_ASAP7_75t_L g2740 ( 
.A(n_2382),
.Y(n_2740)
);

NAND2xp5_ASAP7_75t_L g2741 ( 
.A(n_2592),
.B(n_2089),
.Y(n_2741)
);

NAND2xp33_ASAP7_75t_L g2742 ( 
.A(n_2656),
.B(n_2342),
.Y(n_2742)
);

INVx1_ASAP7_75t_L g2743 ( 
.A(n_2385),
.Y(n_2743)
);

INVx2_ASAP7_75t_L g2744 ( 
.A(n_2417),
.Y(n_2744)
);

INVx1_ASAP7_75t_L g2745 ( 
.A(n_2387),
.Y(n_2745)
);

NAND2xp5_ASAP7_75t_SL g2746 ( 
.A(n_2588),
.B(n_2249),
.Y(n_2746)
);

INVx2_ASAP7_75t_L g2747 ( 
.A(n_2429),
.Y(n_2747)
);

NOR2xp33_ASAP7_75t_L g2748 ( 
.A(n_2408),
.B(n_1190),
.Y(n_2748)
);

INVx2_ASAP7_75t_L g2749 ( 
.A(n_2464),
.Y(n_2749)
);

INVx2_ASAP7_75t_L g2750 ( 
.A(n_2477),
.Y(n_2750)
);

NAND2xp5_ASAP7_75t_SL g2751 ( 
.A(n_2397),
.B(n_2404),
.Y(n_2751)
);

NAND2xp5_ASAP7_75t_L g2752 ( 
.A(n_2383),
.B(n_2089),
.Y(n_2752)
);

INVx2_ASAP7_75t_L g2753 ( 
.A(n_2481),
.Y(n_2753)
);

CKINVDCx5p33_ASAP7_75t_R g2754 ( 
.A(n_2442),
.Y(n_2754)
);

OAI22xp33_ASAP7_75t_L g2755 ( 
.A1(n_2397),
.A2(n_2042),
.B1(n_2100),
.B2(n_2076),
.Y(n_2755)
);

NAND2xp5_ASAP7_75t_L g2756 ( 
.A(n_2544),
.B(n_2041),
.Y(n_2756)
);

NOR2xp33_ASAP7_75t_L g2757 ( 
.A(n_2408),
.B(n_1238),
.Y(n_2757)
);

NAND2xp5_ASAP7_75t_SL g2758 ( 
.A(n_2404),
.B(n_2249),
.Y(n_2758)
);

INVx1_ASAP7_75t_L g2759 ( 
.A(n_2388),
.Y(n_2759)
);

NAND2xp5_ASAP7_75t_SL g2760 ( 
.A(n_2456),
.B(n_2306),
.Y(n_2760)
);

INVx1_ASAP7_75t_L g2761 ( 
.A(n_2393),
.Y(n_2761)
);

INVx2_ASAP7_75t_SL g2762 ( 
.A(n_2484),
.Y(n_2762)
);

INVx1_ASAP7_75t_L g2763 ( 
.A(n_2398),
.Y(n_2763)
);

NAND2xp5_ASAP7_75t_L g2764 ( 
.A(n_2544),
.B(n_2362),
.Y(n_2764)
);

NOR2xp33_ASAP7_75t_L g2765 ( 
.A(n_2506),
.B(n_1238),
.Y(n_2765)
);

AOI22xp5_ASAP7_75t_L g2766 ( 
.A1(n_2506),
.A2(n_2351),
.B1(n_2305),
.B2(n_2319),
.Y(n_2766)
);

OR2x6_ASAP7_75t_L g2767 ( 
.A(n_2405),
.B(n_2299),
.Y(n_2767)
);

INVx2_ASAP7_75t_L g2768 ( 
.A(n_2488),
.Y(n_2768)
);

NAND2xp5_ASAP7_75t_L g2769 ( 
.A(n_2558),
.B(n_2031),
.Y(n_2769)
);

INVx1_ASAP7_75t_L g2770 ( 
.A(n_2400),
.Y(n_2770)
);

NOR2xp33_ASAP7_75t_L g2771 ( 
.A(n_2407),
.B(n_2040),
.Y(n_2771)
);

NAND2xp5_ASAP7_75t_SL g2772 ( 
.A(n_2456),
.B(n_2306),
.Y(n_2772)
);

NAND2xp5_ASAP7_75t_SL g2773 ( 
.A(n_2687),
.B(n_2338),
.Y(n_2773)
);

A2O1A1Ixp33_ASAP7_75t_L g2774 ( 
.A1(n_2517),
.A2(n_2262),
.B(n_2270),
.C(n_2266),
.Y(n_2774)
);

NOR2xp33_ASAP7_75t_L g2775 ( 
.A(n_2426),
.B(n_1669),
.Y(n_2775)
);

NAND3xp33_ASAP7_75t_L g2776 ( 
.A(n_2395),
.B(n_2298),
.C(n_2278),
.Y(n_2776)
);

NOR2xp33_ASAP7_75t_L g2777 ( 
.A(n_2497),
.B(n_2628),
.Y(n_2777)
);

AND3x1_ASAP7_75t_L g2778 ( 
.A(n_2667),
.B(n_2305),
.C(n_2295),
.Y(n_2778)
);

BUFx6f_ASAP7_75t_L g2779 ( 
.A(n_2656),
.Y(n_2779)
);

INVx1_ASAP7_75t_L g2780 ( 
.A(n_2401),
.Y(n_2780)
);

NOR3xp33_ASAP7_75t_L g2781 ( 
.A(n_2691),
.B(n_2332),
.C(n_2132),
.Y(n_2781)
);

INVx1_ASAP7_75t_L g2782 ( 
.A(n_2403),
.Y(n_2782)
);

CKINVDCx5p33_ASAP7_75t_R g2783 ( 
.A(n_2420),
.Y(n_2783)
);

NOR2xp33_ASAP7_75t_L g2784 ( 
.A(n_2691),
.B(n_1669),
.Y(n_2784)
);

NOR2xp33_ASAP7_75t_L g2785 ( 
.A(n_2548),
.B(n_1771),
.Y(n_2785)
);

NOR2xp33_ASAP7_75t_L g2786 ( 
.A(n_2548),
.B(n_1771),
.Y(n_2786)
);

A2O1A1Ixp33_ASAP7_75t_L g2787 ( 
.A1(n_2517),
.A2(n_2262),
.B(n_2270),
.C(n_2266),
.Y(n_2787)
);

NAND2xp5_ASAP7_75t_SL g2788 ( 
.A(n_2698),
.B(n_2338),
.Y(n_2788)
);

BUFx8_ASAP7_75t_L g2789 ( 
.A(n_2391),
.Y(n_2789)
);

NAND2xp5_ASAP7_75t_L g2790 ( 
.A(n_2558),
.B(n_2205),
.Y(n_2790)
);

OAI22xp5_ASAP7_75t_L g2791 ( 
.A1(n_2383),
.A2(n_2198),
.B1(n_2275),
.B2(n_2273),
.Y(n_2791)
);

INVx2_ASAP7_75t_SL g2792 ( 
.A(n_2422),
.Y(n_2792)
);

INVxp67_ASAP7_75t_L g2793 ( 
.A(n_2422),
.Y(n_2793)
);

BUFx6f_ASAP7_75t_SL g2794 ( 
.A(n_2573),
.Y(n_2794)
);

NAND2xp5_ASAP7_75t_L g2795 ( 
.A(n_2563),
.B(n_2525),
.Y(n_2795)
);

INVx2_ASAP7_75t_L g2796 ( 
.A(n_2492),
.Y(n_2796)
);

AOI22xp5_ASAP7_75t_L g2797 ( 
.A1(n_2576),
.A2(n_2319),
.B1(n_2113),
.B2(n_2141),
.Y(n_2797)
);

INVx2_ASAP7_75t_L g2798 ( 
.A(n_2518),
.Y(n_2798)
);

O2A1O1Ixp33_ASAP7_75t_L g2799 ( 
.A1(n_2569),
.A2(n_2137),
.B(n_2256),
.C(n_2359),
.Y(n_2799)
);

INVx1_ASAP7_75t_L g2800 ( 
.A(n_2409),
.Y(n_2800)
);

NAND2xp5_ASAP7_75t_SL g2801 ( 
.A(n_2566),
.B(n_2339),
.Y(n_2801)
);

NAND2xp5_ASAP7_75t_SL g2802 ( 
.A(n_2450),
.B(n_2339),
.Y(n_2802)
);

INVx2_ASAP7_75t_L g2803 ( 
.A(n_2582),
.Y(n_2803)
);

BUFx6f_ASAP7_75t_L g2804 ( 
.A(n_2656),
.Y(n_2804)
);

AOI221xp5_ASAP7_75t_L g2805 ( 
.A1(n_2657),
.A2(n_1892),
.B1(n_776),
.B2(n_829),
.C(n_774),
.Y(n_2805)
);

NAND2xp5_ASAP7_75t_SL g2806 ( 
.A(n_2542),
.B(n_2347),
.Y(n_2806)
);

OAI22xp5_ASAP7_75t_L g2807 ( 
.A1(n_2414),
.A2(n_2274),
.B1(n_2273),
.B2(n_2275),
.Y(n_2807)
);

INVx2_ASAP7_75t_SL g2808 ( 
.A(n_2515),
.Y(n_2808)
);

INVx2_ASAP7_75t_SL g2809 ( 
.A(n_2591),
.Y(n_2809)
);

INVx2_ASAP7_75t_L g2810 ( 
.A(n_2589),
.Y(n_2810)
);

OAI221xp5_ASAP7_75t_L g2811 ( 
.A1(n_2657),
.A2(n_2370),
.B1(n_2100),
.B2(n_2186),
.C(n_2136),
.Y(n_2811)
);

NAND2xp5_ASAP7_75t_L g2812 ( 
.A(n_2563),
.B(n_2076),
.Y(n_2812)
);

NAND2xp5_ASAP7_75t_L g2813 ( 
.A(n_2525),
.B(n_2136),
.Y(n_2813)
);

NAND2xp5_ASAP7_75t_L g2814 ( 
.A(n_2414),
.B(n_2437),
.Y(n_2814)
);

INVx2_ASAP7_75t_L g2815 ( 
.A(n_2609),
.Y(n_2815)
);

INVx1_ASAP7_75t_L g2816 ( 
.A(n_2412),
.Y(n_2816)
);

INVx2_ASAP7_75t_L g2817 ( 
.A(n_2646),
.Y(n_2817)
);

AND2x2_ASAP7_75t_L g2818 ( 
.A(n_2440),
.B(n_1749),
.Y(n_2818)
);

NAND2xp5_ASAP7_75t_L g2819 ( 
.A(n_2536),
.B(n_2302),
.Y(n_2819)
);

INVx1_ASAP7_75t_L g2820 ( 
.A(n_2415),
.Y(n_2820)
);

NAND2xp5_ASAP7_75t_L g2821 ( 
.A(n_2536),
.B(n_2302),
.Y(n_2821)
);

BUFx6f_ASAP7_75t_L g2822 ( 
.A(n_2602),
.Y(n_2822)
);

INVx3_ASAP7_75t_L g2823 ( 
.A(n_2618),
.Y(n_2823)
);

NAND2xp5_ASAP7_75t_L g2824 ( 
.A(n_2437),
.B(n_2491),
.Y(n_2824)
);

NOR2xp33_ASAP7_75t_SL g2825 ( 
.A(n_2618),
.B(n_2014),
.Y(n_2825)
);

INVx2_ASAP7_75t_L g2826 ( 
.A(n_2598),
.Y(n_2826)
);

NAND2xp5_ASAP7_75t_SL g2827 ( 
.A(n_2602),
.B(n_2347),
.Y(n_2827)
);

NAND2xp33_ASAP7_75t_L g2828 ( 
.A(n_2633),
.B(n_2342),
.Y(n_2828)
);

NAND2xp5_ASAP7_75t_L g2829 ( 
.A(n_2629),
.B(n_2186),
.Y(n_2829)
);

NAND3xp33_ASAP7_75t_L g2830 ( 
.A(n_2474),
.B(n_2277),
.C(n_2210),
.Y(n_2830)
);

NOR2xp33_ASAP7_75t_L g2831 ( 
.A(n_2664),
.B(n_1612),
.Y(n_2831)
);

NAND2xp5_ASAP7_75t_L g2832 ( 
.A(n_2629),
.B(n_2189),
.Y(n_2832)
);

INVx1_ASAP7_75t_L g2833 ( 
.A(n_2416),
.Y(n_2833)
);

OAI22xp5_ASAP7_75t_L g2834 ( 
.A1(n_2433),
.A2(n_2274),
.B1(n_2049),
.B2(n_2045),
.Y(n_2834)
);

NAND2xp5_ASAP7_75t_L g2835 ( 
.A(n_2616),
.B(n_2189),
.Y(n_2835)
);

INVx1_ASAP7_75t_L g2836 ( 
.A(n_2419),
.Y(n_2836)
);

NAND2xp5_ASAP7_75t_L g2837 ( 
.A(n_2616),
.B(n_2205),
.Y(n_2837)
);

NOR2xp33_ASAP7_75t_L g2838 ( 
.A(n_2664),
.B(n_1627),
.Y(n_2838)
);

INVx1_ASAP7_75t_L g2839 ( 
.A(n_2421),
.Y(n_2839)
);

AOI22xp33_ASAP7_75t_L g2840 ( 
.A1(n_2529),
.A2(n_2097),
.B1(n_2258),
.B2(n_2342),
.Y(n_2840)
);

NOR2xp33_ASAP7_75t_L g2841 ( 
.A(n_2639),
.B(n_1627),
.Y(n_2841)
);

INVx2_ASAP7_75t_L g2842 ( 
.A(n_2599),
.Y(n_2842)
);

NAND3xp33_ASAP7_75t_L g2843 ( 
.A(n_2581),
.B(n_2277),
.C(n_2140),
.Y(n_2843)
);

OR2x2_ASAP7_75t_L g2844 ( 
.A(n_2639),
.B(n_2258),
.Y(n_2844)
);

NAND2xp5_ASAP7_75t_L g2845 ( 
.A(n_2491),
.B(n_2316),
.Y(n_2845)
);

NOR2xp67_ASAP7_75t_L g2846 ( 
.A(n_2644),
.B(n_1583),
.Y(n_2846)
);

INVx2_ASAP7_75t_L g2847 ( 
.A(n_2600),
.Y(n_2847)
);

NOR3x1_ASAP7_75t_L g2848 ( 
.A(n_2641),
.B(n_1304),
.C(n_1303),
.Y(n_2848)
);

INVx2_ASAP7_75t_L g2849 ( 
.A(n_2603),
.Y(n_2849)
);

INVx2_ASAP7_75t_L g2850 ( 
.A(n_2604),
.Y(n_2850)
);

NOR2xp33_ASAP7_75t_L g2851 ( 
.A(n_2479),
.B(n_1644),
.Y(n_2851)
);

NAND2xp5_ASAP7_75t_L g2852 ( 
.A(n_2500),
.B(n_2316),
.Y(n_2852)
);

OR2x2_ASAP7_75t_L g2853 ( 
.A(n_2394),
.B(n_2316),
.Y(n_2853)
);

INVx2_ASAP7_75t_SL g2854 ( 
.A(n_2571),
.Y(n_2854)
);

NAND2xp33_ASAP7_75t_L g2855 ( 
.A(n_2633),
.B(n_2342),
.Y(n_2855)
);

NAND2xp5_ASAP7_75t_L g2856 ( 
.A(n_2500),
.B(n_2049),
.Y(n_2856)
);

OAI21xp5_ASAP7_75t_L g2857 ( 
.A1(n_2443),
.A2(n_2038),
.B(n_2034),
.Y(n_2857)
);

INVx1_ASAP7_75t_L g2858 ( 
.A(n_2425),
.Y(n_2858)
);

AOI22xp5_ASAP7_75t_L g2859 ( 
.A1(n_2673),
.A2(n_2342),
.B1(n_2097),
.B2(n_2115),
.Y(n_2859)
);

NOR2xp67_ASAP7_75t_L g2860 ( 
.A(n_2644),
.B(n_1582),
.Y(n_2860)
);

BUFx6f_ASAP7_75t_L g2861 ( 
.A(n_2547),
.Y(n_2861)
);

AND2x6_ASAP7_75t_SL g2862 ( 
.A(n_2667),
.B(n_1644),
.Y(n_2862)
);

NOR2xp33_ASAP7_75t_L g2863 ( 
.A(n_2479),
.B(n_1582),
.Y(n_2863)
);

NAND2xp5_ASAP7_75t_SL g2864 ( 
.A(n_2389),
.B(n_2311),
.Y(n_2864)
);

INVx4_ASAP7_75t_L g2865 ( 
.A(n_2720),
.Y(n_2865)
);

A2O1A1Ixp33_ASAP7_75t_L g2866 ( 
.A1(n_2581),
.A2(n_2498),
.B(n_2523),
.C(n_2680),
.Y(n_2866)
);

OR2x6_ASAP7_75t_L g2867 ( 
.A(n_2534),
.B(n_2299),
.Y(n_2867)
);

NAND2xp5_ASAP7_75t_L g2868 ( 
.A(n_2555),
.B(n_2016),
.Y(n_2868)
);

OR2x2_ASAP7_75t_L g2869 ( 
.A(n_2423),
.B(n_2467),
.Y(n_2869)
);

NAND2xp5_ASAP7_75t_SL g2870 ( 
.A(n_2459),
.B(n_2311),
.Y(n_2870)
);

NAND2xp5_ASAP7_75t_SL g2871 ( 
.A(n_2682),
.B(n_2311),
.Y(n_2871)
);

INVx2_ASAP7_75t_L g2872 ( 
.A(n_2605),
.Y(n_2872)
);

INVx2_ASAP7_75t_L g2873 ( 
.A(n_2610),
.Y(n_2873)
);

NAND2xp5_ASAP7_75t_L g2874 ( 
.A(n_2555),
.B(n_2016),
.Y(n_2874)
);

INVx2_ASAP7_75t_L g2875 ( 
.A(n_2612),
.Y(n_2875)
);

INVx2_ASAP7_75t_L g2876 ( 
.A(n_2613),
.Y(n_2876)
);

INVx2_ASAP7_75t_L g2877 ( 
.A(n_2614),
.Y(n_2877)
);

NAND2xp5_ASAP7_75t_SL g2878 ( 
.A(n_2682),
.B(n_2214),
.Y(n_2878)
);

INVx2_ASAP7_75t_SL g2879 ( 
.A(n_2508),
.Y(n_2879)
);

INVx2_ASAP7_75t_L g2880 ( 
.A(n_2615),
.Y(n_2880)
);

NAND2xp5_ASAP7_75t_L g2881 ( 
.A(n_2637),
.B(n_2140),
.Y(n_2881)
);

NAND2xp5_ASAP7_75t_L g2882 ( 
.A(n_2503),
.B(n_2342),
.Y(n_2882)
);

AOI22xp5_ASAP7_75t_L g2883 ( 
.A1(n_2689),
.A2(n_2115),
.B1(n_2320),
.B2(n_2299),
.Y(n_2883)
);

INVx1_ASAP7_75t_L g2884 ( 
.A(n_2427),
.Y(n_2884)
);

NOR2xp33_ASAP7_75t_L g2885 ( 
.A(n_2534),
.B(n_1583),
.Y(n_2885)
);

OAI22xp5_ASAP7_75t_L g2886 ( 
.A1(n_2433),
.A2(n_2019),
.B1(n_2022),
.B2(n_2021),
.Y(n_2886)
);

NOR2xp33_ASAP7_75t_L g2887 ( 
.A(n_2516),
.B(n_1628),
.Y(n_2887)
);

AO22x1_ASAP7_75t_L g2888 ( 
.A1(n_2680),
.A2(n_1706),
.B1(n_1777),
.B2(n_1686),
.Y(n_2888)
);

NAND2xp5_ASAP7_75t_L g2889 ( 
.A(n_2507),
.B(n_2214),
.Y(n_2889)
);

INVx1_ASAP7_75t_SL g2890 ( 
.A(n_2606),
.Y(n_2890)
);

NOR2xp33_ASAP7_75t_L g2891 ( 
.A(n_2619),
.B(n_2594),
.Y(n_2891)
);

O2A1O1Ixp33_ASAP7_75t_L g2892 ( 
.A1(n_2577),
.A2(n_2143),
.B(n_1815),
.C(n_1830),
.Y(n_2892)
);

NOR2xp33_ASAP7_75t_L g2893 ( 
.A(n_2625),
.B(n_1628),
.Y(n_2893)
);

NAND2xp5_ASAP7_75t_L g2894 ( 
.A(n_2386),
.B(n_2019),
.Y(n_2894)
);

AOI22xp33_ASAP7_75t_SL g2895 ( 
.A1(n_2593),
.A2(n_2320),
.B1(n_2299),
.B2(n_1686),
.Y(n_2895)
);

INVx2_ASAP7_75t_SL g2896 ( 
.A(n_2562),
.Y(n_2896)
);

NAND2xp5_ASAP7_75t_SL g2897 ( 
.A(n_2607),
.B(n_2214),
.Y(n_2897)
);

INVx2_ASAP7_75t_L g2898 ( 
.A(n_2617),
.Y(n_2898)
);

AOI221xp5_ASAP7_75t_L g2899 ( 
.A1(n_2549),
.A2(n_582),
.B1(n_595),
.B2(n_606),
.C(n_594),
.Y(n_2899)
);

INVx2_ASAP7_75t_L g2900 ( 
.A(n_2620),
.Y(n_2900)
);

INVx1_ASAP7_75t_L g2901 ( 
.A(n_2430),
.Y(n_2901)
);

INVx2_ASAP7_75t_L g2902 ( 
.A(n_2621),
.Y(n_2902)
);

BUFx6f_ASAP7_75t_L g2903 ( 
.A(n_2556),
.Y(n_2903)
);

AOI22xp5_ASAP7_75t_L g2904 ( 
.A1(n_2565),
.A2(n_2115),
.B1(n_2320),
.B2(n_2263),
.Y(n_2904)
);

NOR2xp33_ASAP7_75t_L g2905 ( 
.A(n_2709),
.B(n_1345),
.Y(n_2905)
);

INVx1_ASAP7_75t_L g2906 ( 
.A(n_2431),
.Y(n_2906)
);

INVx3_ASAP7_75t_L g2907 ( 
.A(n_2457),
.Y(n_2907)
);

AND2x6_ASAP7_75t_SL g2908 ( 
.A(n_2650),
.B(n_1345),
.Y(n_2908)
);

NOR3xp33_ASAP7_75t_L g2909 ( 
.A(n_2478),
.B(n_2215),
.C(n_1616),
.Y(n_2909)
);

INVx1_ASAP7_75t_L g2910 ( 
.A(n_2432),
.Y(n_2910)
);

NOR2xp33_ASAP7_75t_L g2911 ( 
.A(n_2711),
.B(n_2716),
.Y(n_2911)
);

OAI221xp5_ASAP7_75t_L g2912 ( 
.A1(n_2643),
.A2(n_606),
.B1(n_610),
.B2(n_595),
.C(n_594),
.Y(n_2912)
);

O2A1O1Ixp33_ASAP7_75t_L g2913 ( 
.A1(n_2386),
.A2(n_2143),
.B(n_1815),
.C(n_1830),
.Y(n_2913)
);

AND2x2_ASAP7_75t_L g2914 ( 
.A(n_2570),
.B(n_1749),
.Y(n_2914)
);

NAND2xp5_ASAP7_75t_SL g2915 ( 
.A(n_2654),
.B(n_2263),
.Y(n_2915)
);

BUFx5_ASAP7_75t_L g2916 ( 
.A(n_2630),
.Y(n_2916)
);

NAND2xp5_ASAP7_75t_SL g2917 ( 
.A(n_2654),
.B(n_2263),
.Y(n_2917)
);

INVx2_ASAP7_75t_L g2918 ( 
.A(n_2623),
.Y(n_2918)
);

NAND2xp5_ASAP7_75t_L g2919 ( 
.A(n_2510),
.B(n_2320),
.Y(n_2919)
);

INVx1_ASAP7_75t_L g2920 ( 
.A(n_2434),
.Y(n_2920)
);

INVx2_ASAP7_75t_SL g2921 ( 
.A(n_2418),
.Y(n_2921)
);

NAND2xp5_ASAP7_75t_SL g2922 ( 
.A(n_2671),
.B(n_2320),
.Y(n_2922)
);

NAND2xp5_ASAP7_75t_L g2923 ( 
.A(n_2511),
.B(n_2081),
.Y(n_2923)
);

NAND2xp5_ASAP7_75t_SL g2924 ( 
.A(n_2671),
.B(n_2086),
.Y(n_2924)
);

INVx1_ASAP7_75t_L g2925 ( 
.A(n_2435),
.Y(n_2925)
);

NAND2xp5_ASAP7_75t_L g2926 ( 
.A(n_2512),
.B(n_2084),
.Y(n_2926)
);

NAND2xp5_ASAP7_75t_SL g2927 ( 
.A(n_2685),
.B(n_2086),
.Y(n_2927)
);

BUFx5_ASAP7_75t_L g2928 ( 
.A(n_2630),
.Y(n_2928)
);

INVx2_ASAP7_75t_SL g2929 ( 
.A(n_2418),
.Y(n_2929)
);

AO22x1_ASAP7_75t_L g2930 ( 
.A1(n_2718),
.A2(n_1777),
.B1(n_1847),
.B2(n_1706),
.Y(n_2930)
);

NOR2xp67_ASAP7_75t_L g2931 ( 
.A(n_2650),
.B(n_1815),
.Y(n_2931)
);

BUFx2_ASAP7_75t_L g2932 ( 
.A(n_2651),
.Y(n_2932)
);

NAND2xp5_ASAP7_75t_SL g2933 ( 
.A(n_2545),
.B(n_2560),
.Y(n_2933)
);

NAND2xp5_ASAP7_75t_SL g2934 ( 
.A(n_2686),
.B(n_2086),
.Y(n_2934)
);

NAND2xp5_ASAP7_75t_L g2935 ( 
.A(n_2521),
.B(n_2084),
.Y(n_2935)
);

NOR3xp33_ASAP7_75t_L g2936 ( 
.A(n_2486),
.B(n_1830),
.C(n_1940),
.Y(n_2936)
);

NAND2xp5_ASAP7_75t_L g2937 ( 
.A(n_2526),
.B(n_2084),
.Y(n_2937)
);

NOR2xp33_ASAP7_75t_L g2938 ( 
.A(n_2509),
.B(n_1706),
.Y(n_2938)
);

INVx2_ASAP7_75t_L g2939 ( 
.A(n_2626),
.Y(n_2939)
);

INVx2_ASAP7_75t_SL g2940 ( 
.A(n_2445),
.Y(n_2940)
);

INVx2_ASAP7_75t_L g2941 ( 
.A(n_2631),
.Y(n_2941)
);

INVx1_ASAP7_75t_L g2942 ( 
.A(n_2436),
.Y(n_2942)
);

AOI22xp5_ASAP7_75t_L g2943 ( 
.A1(n_2524),
.A2(n_2164),
.B1(n_2188),
.B2(n_2086),
.Y(n_2943)
);

AND2x6_ASAP7_75t_SL g2944 ( 
.A(n_2601),
.B(n_1959),
.Y(n_2944)
);

AO221x1_ASAP7_75t_L g2945 ( 
.A1(n_2665),
.A2(n_2188),
.B1(n_2086),
.B2(n_2148),
.C(n_2181),
.Y(n_2945)
);

NAND2xp5_ASAP7_75t_L g2946 ( 
.A(n_2527),
.B(n_2091),
.Y(n_2946)
);

NAND2xp5_ASAP7_75t_L g2947 ( 
.A(n_2520),
.B(n_2021),
.Y(n_2947)
);

NOR3xp33_ASAP7_75t_L g2948 ( 
.A(n_2700),
.B(n_1963),
.C(n_1085),
.Y(n_2948)
);

INVx1_ASAP7_75t_L g2949 ( 
.A(n_2438),
.Y(n_2949)
);

AND2x2_ASAP7_75t_L g2950 ( 
.A(n_2622),
.B(n_1963),
.Y(n_2950)
);

NAND2xp5_ASAP7_75t_L g2951 ( 
.A(n_2520),
.B(n_2022),
.Y(n_2951)
);

OR2x6_ASAP7_75t_L g2952 ( 
.A(n_2703),
.B(n_2014),
.Y(n_2952)
);

O2A1O1Ixp5_ASAP7_75t_L g2953 ( 
.A1(n_2413),
.A2(n_2354),
.B(n_2361),
.C(n_2345),
.Y(n_2953)
);

NAND2xp5_ASAP7_75t_SL g2954 ( 
.A(n_2595),
.B(n_2188),
.Y(n_2954)
);

BUFx6f_ASAP7_75t_L g2955 ( 
.A(n_2445),
.Y(n_2955)
);

INVx2_ASAP7_75t_L g2956 ( 
.A(n_2632),
.Y(n_2956)
);

HB1xp67_ASAP7_75t_L g2957 ( 
.A(n_2713),
.Y(n_2957)
);

NAND2xp5_ASAP7_75t_SL g2958 ( 
.A(n_2595),
.B(n_2188),
.Y(n_2958)
);

BUFx8_ASAP7_75t_L g2959 ( 
.A(n_2714),
.Y(n_2959)
);

NOR2xp33_ASAP7_75t_R g2960 ( 
.A(n_2411),
.B(n_1777),
.Y(n_2960)
);

INVx2_ASAP7_75t_L g2961 ( 
.A(n_2634),
.Y(n_2961)
);

NAND2xp5_ASAP7_75t_SL g2962 ( 
.A(n_2627),
.B(n_2188),
.Y(n_2962)
);

NAND2xp5_ASAP7_75t_SL g2963 ( 
.A(n_2627),
.B(n_1963),
.Y(n_2963)
);

AOI22xp33_ASAP7_75t_L g2964 ( 
.A1(n_2624),
.A2(n_2164),
.B1(n_2242),
.B2(n_2236),
.Y(n_2964)
);

INVx2_ASAP7_75t_SL g2965 ( 
.A(n_2636),
.Y(n_2965)
);

INVx2_ASAP7_75t_SL g2966 ( 
.A(n_2636),
.Y(n_2966)
);

NAND2xp5_ASAP7_75t_SL g2967 ( 
.A(n_2624),
.B(n_2127),
.Y(n_2967)
);

AOI22xp5_ASAP7_75t_L g2968 ( 
.A1(n_2643),
.A2(n_2164),
.B1(n_2025),
.B2(n_2044),
.Y(n_2968)
);

INVx5_ASAP7_75t_L g2969 ( 
.A(n_2630),
.Y(n_2969)
);

NOR2xp33_ASAP7_75t_L g2970 ( 
.A(n_2672),
.B(n_1847),
.Y(n_2970)
);

NAND2xp5_ASAP7_75t_SL g2971 ( 
.A(n_2528),
.B(n_2127),
.Y(n_2971)
);

NAND2xp5_ASAP7_75t_L g2972 ( 
.A(n_2540),
.B(n_2024),
.Y(n_2972)
);

NAND2xp5_ASAP7_75t_L g2973 ( 
.A(n_2530),
.B(n_2091),
.Y(n_2973)
);

NAND2xp5_ASAP7_75t_SL g2974 ( 
.A(n_2531),
.B(n_2533),
.Y(n_2974)
);

INVxp67_ASAP7_75t_SL g2975 ( 
.A(n_2540),
.Y(n_2975)
);

INVx2_ASAP7_75t_L g2976 ( 
.A(n_2635),
.Y(n_2976)
);

INVx2_ASAP7_75t_SL g2977 ( 
.A(n_2514),
.Y(n_2977)
);

NAND2xp5_ASAP7_75t_SL g2978 ( 
.A(n_2535),
.B(n_2127),
.Y(n_2978)
);

INVxp67_ASAP7_75t_L g2979 ( 
.A(n_2505),
.Y(n_2979)
);

AOI21xp5_ASAP7_75t_L g2980 ( 
.A1(n_2572),
.A2(n_2025),
.B(n_2014),
.Y(n_2980)
);

NAND2xp5_ASAP7_75t_L g2981 ( 
.A(n_2537),
.B(n_2538),
.Y(n_2981)
);

OAI22xp5_ASAP7_75t_L g2982 ( 
.A1(n_2572),
.A2(n_2541),
.B1(n_2546),
.B2(n_2543),
.Y(n_2982)
);

INVx2_ASAP7_75t_L g2983 ( 
.A(n_2638),
.Y(n_2983)
);

AND2x6_ASAP7_75t_SL g2984 ( 
.A(n_2392),
.B(n_1847),
.Y(n_2984)
);

AND2x4_ASAP7_75t_L g2985 ( 
.A(n_2539),
.B(n_2354),
.Y(n_2985)
);

OR2x6_ASAP7_75t_L g2986 ( 
.A(n_2476),
.B(n_2014),
.Y(n_2986)
);

NAND2xp5_ASAP7_75t_L g2987 ( 
.A(n_2551),
.B(n_2091),
.Y(n_2987)
);

NAND2xp5_ASAP7_75t_L g2988 ( 
.A(n_2553),
.B(n_2026),
.Y(n_2988)
);

INVx1_ASAP7_75t_L g2989 ( 
.A(n_2666),
.Y(n_2989)
);

INVx1_ASAP7_75t_L g2990 ( 
.A(n_2668),
.Y(n_2990)
);

NAND2xp5_ASAP7_75t_L g2991 ( 
.A(n_2554),
.B(n_2557),
.Y(n_2991)
);

NAND2xp5_ASAP7_75t_L g2992 ( 
.A(n_2559),
.B(n_2026),
.Y(n_2992)
);

A2O1A1Ixp33_ASAP7_75t_L g2993 ( 
.A1(n_2561),
.A2(n_2025),
.B(n_2044),
.C(n_2014),
.Y(n_2993)
);

OAI22xp33_ASAP7_75t_L g2994 ( 
.A1(n_2453),
.A2(n_2025),
.B1(n_2044),
.B2(n_2242),
.Y(n_2994)
);

NOR2xp33_ASAP7_75t_L g2995 ( 
.A(n_2706),
.B(n_2027),
.Y(n_2995)
);

AOI22xp5_ASAP7_75t_L g2996 ( 
.A1(n_2502),
.A2(n_2044),
.B1(n_2025),
.B2(n_1816),
.Y(n_2996)
);

NAND2xp5_ASAP7_75t_L g2997 ( 
.A(n_2633),
.B(n_2024),
.Y(n_2997)
);

INVx2_ASAP7_75t_SL g2998 ( 
.A(n_2693),
.Y(n_2998)
);

NAND2xp5_ASAP7_75t_L g2999 ( 
.A(n_2633),
.B(n_2026),
.Y(n_2999)
);

NAND2xp5_ASAP7_75t_L g3000 ( 
.A(n_2633),
.B(n_2029),
.Y(n_3000)
);

INVx1_ASAP7_75t_L g3001 ( 
.A(n_2669),
.Y(n_3001)
);

INVx2_ASAP7_75t_SL g3002 ( 
.A(n_2712),
.Y(n_3002)
);

INVx1_ASAP7_75t_L g3003 ( 
.A(n_2670),
.Y(n_3003)
);

AOI22xp5_ASAP7_75t_L g3004 ( 
.A1(n_2550),
.A2(n_2567),
.B1(n_2568),
.B2(n_2564),
.Y(n_3004)
);

INVx4_ASAP7_75t_L g3005 ( 
.A(n_2720),
.Y(n_3005)
);

INVx2_ASAP7_75t_L g3006 ( 
.A(n_2640),
.Y(n_3006)
);

NOR2xp33_ASAP7_75t_L g3007 ( 
.A(n_2519),
.B(n_2260),
.Y(n_3007)
);

OAI21xp33_ASAP7_75t_L g3008 ( 
.A1(n_2574),
.A2(n_612),
.B(n_610),
.Y(n_3008)
);

NAND2xp5_ASAP7_75t_L g3009 ( 
.A(n_2575),
.B(n_2236),
.Y(n_3009)
);

INVx2_ASAP7_75t_SL g3010 ( 
.A(n_2447),
.Y(n_3010)
);

AOI22xp33_ASAP7_75t_L g3011 ( 
.A1(n_2439),
.A2(n_2441),
.B1(n_2451),
.B2(n_2449),
.Y(n_3011)
);

NAND2xp5_ASAP7_75t_SL g3012 ( 
.A(n_2578),
.B(n_2127),
.Y(n_3012)
);

INVx1_ASAP7_75t_L g3013 ( 
.A(n_2674),
.Y(n_3013)
);

INVx2_ASAP7_75t_SL g3014 ( 
.A(n_2454),
.Y(n_3014)
);

NAND3xp33_ASAP7_75t_L g3015 ( 
.A(n_2413),
.B(n_2150),
.C(n_2144),
.Y(n_3015)
);

BUFx3_ASAP7_75t_L g3016 ( 
.A(n_2493),
.Y(n_3016)
);

NAND2xp5_ASAP7_75t_L g3017 ( 
.A(n_2579),
.B(n_2583),
.Y(n_3017)
);

INVx2_ASAP7_75t_L g3018 ( 
.A(n_2642),
.Y(n_3018)
);

AOI221xp5_ASAP7_75t_L g3019 ( 
.A1(n_2585),
.A2(n_620),
.B1(n_622),
.B2(n_613),
.C(n_612),
.Y(n_3019)
);

INVx2_ASAP7_75t_L g3020 ( 
.A(n_2647),
.Y(n_3020)
);

NAND2x1p5_ASAP7_75t_L g3021 ( 
.A(n_2969),
.B(n_2720),
.Y(n_3021)
);

INVx2_ASAP7_75t_L g3022 ( 
.A(n_2826),
.Y(n_3022)
);

AOI21xp5_ASAP7_75t_L g3023 ( 
.A1(n_2828),
.A2(n_2044),
.B(n_2170),
.Y(n_3023)
);

AO21x2_ASAP7_75t_L g3024 ( 
.A1(n_2859),
.A2(n_2611),
.B(n_2443),
.Y(n_3024)
);

AOI21xp5_ASAP7_75t_L g3025 ( 
.A1(n_2855),
.A2(n_2190),
.B(n_2170),
.Y(n_3025)
);

O2A1O1Ixp33_ASAP7_75t_L g3026 ( 
.A1(n_2785),
.A2(n_2453),
.B(n_2652),
.C(n_2649),
.Y(n_3026)
);

NAND2xp5_ASAP7_75t_L g3027 ( 
.A(n_2764),
.B(n_2586),
.Y(n_3027)
);

OR2x2_ASAP7_75t_L g3028 ( 
.A(n_2869),
.B(n_2590),
.Y(n_3028)
);

NAND2xp5_ASAP7_75t_SL g3029 ( 
.A(n_2727),
.B(n_2697),
.Y(n_3029)
);

INVx1_ASAP7_75t_L g3030 ( 
.A(n_2724),
.Y(n_3030)
);

AOI21xp5_ASAP7_75t_L g3031 ( 
.A1(n_2814),
.A2(n_2190),
.B(n_2170),
.Y(n_3031)
);

INVx2_ASAP7_75t_SL g3032 ( 
.A(n_2789),
.Y(n_3032)
);

OAI22xp5_ASAP7_75t_L g3033 ( 
.A1(n_2866),
.A2(n_2455),
.B1(n_2460),
.B2(n_2458),
.Y(n_3033)
);

AND2x2_ASAP7_75t_L g3034 ( 
.A(n_2818),
.B(n_2596),
.Y(n_3034)
);

A2O1A1Ixp33_ASAP7_75t_L g3035 ( 
.A1(n_2765),
.A2(n_2461),
.B(n_2463),
.C(n_2462),
.Y(n_3035)
);

AOI21xp5_ASAP7_75t_L g3036 ( 
.A1(n_2814),
.A2(n_2729),
.B(n_2824),
.Y(n_3036)
);

AOI21xp5_ASAP7_75t_L g3037 ( 
.A1(n_2824),
.A2(n_2190),
.B(n_2170),
.Y(n_3037)
);

OAI21xp5_ASAP7_75t_L g3038 ( 
.A1(n_2795),
.A2(n_2611),
.B(n_2485),
.Y(n_3038)
);

NOR2xp33_ASAP7_75t_L g3039 ( 
.A(n_2731),
.B(n_2390),
.Y(n_3039)
);

INVx2_ASAP7_75t_L g3040 ( 
.A(n_2842),
.Y(n_3040)
);

O2A1O1Ixp33_ASAP7_75t_SL g3041 ( 
.A1(n_2756),
.A2(n_2655),
.B(n_2658),
.C(n_2653),
.Y(n_3041)
);

NAND2xp5_ASAP7_75t_L g3042 ( 
.A(n_2730),
.B(n_2597),
.Y(n_3042)
);

INVxp67_ASAP7_75t_L g3043 ( 
.A(n_2777),
.Y(n_3043)
);

AOI21xp5_ASAP7_75t_L g3044 ( 
.A1(n_2752),
.A2(n_2206),
.B(n_2190),
.Y(n_3044)
);

INVx1_ASAP7_75t_SL g3045 ( 
.A(n_2725),
.Y(n_3045)
);

O2A1O1Ixp33_ASAP7_75t_L g3046 ( 
.A1(n_2786),
.A2(n_2660),
.B(n_2661),
.C(n_2659),
.Y(n_3046)
);

AOI21xp5_ASAP7_75t_L g3047 ( 
.A1(n_2752),
.A2(n_2245),
.B(n_2206),
.Y(n_3047)
);

NAND2x1_ASAP7_75t_L g3048 ( 
.A(n_2865),
.B(n_2206),
.Y(n_3048)
);

NAND2xp5_ASAP7_75t_L g3049 ( 
.A(n_2751),
.B(n_2662),
.Y(n_3049)
);

AND2x2_ASAP7_75t_L g3050 ( 
.A(n_2995),
.B(n_2663),
.Y(n_3050)
);

NAND2xp5_ASAP7_75t_L g3051 ( 
.A(n_2890),
.B(n_2466),
.Y(n_3051)
);

NOR2xp33_ASAP7_75t_L g3052 ( 
.A(n_2748),
.B(n_2584),
.Y(n_3052)
);

OAI22xp5_ASAP7_75t_L g3053 ( 
.A1(n_2728),
.A2(n_2469),
.B1(n_2471),
.B2(n_2470),
.Y(n_3053)
);

INVx4_ASAP7_75t_L g3054 ( 
.A(n_2779),
.Y(n_3054)
);

AO21x1_ASAP7_75t_L g3055 ( 
.A1(n_2735),
.A2(n_2958),
.B(n_2954),
.Y(n_3055)
);

AOI21xp5_ASAP7_75t_L g3056 ( 
.A1(n_2774),
.A2(n_2245),
.B(n_2206),
.Y(n_3056)
);

NAND2xp5_ASAP7_75t_L g3057 ( 
.A(n_2890),
.B(n_2790),
.Y(n_3057)
);

BUFx6f_ASAP7_75t_L g3058 ( 
.A(n_2779),
.Y(n_3058)
);

BUFx6f_ASAP7_75t_L g3059 ( 
.A(n_2779),
.Y(n_3059)
);

AND2x4_ASAP7_75t_L g3060 ( 
.A(n_2822),
.B(n_2446),
.Y(n_3060)
);

AOI21xp5_ASAP7_75t_L g3061 ( 
.A1(n_2787),
.A2(n_2250),
.B(n_2245),
.Y(n_3061)
);

NAND2xp5_ASAP7_75t_SL g3062 ( 
.A(n_2725),
.B(n_2784),
.Y(n_3062)
);

A2O1A1Ixp33_ASAP7_75t_L g3063 ( 
.A1(n_2776),
.A2(n_2473),
.B(n_2475),
.C(n_2482),
.Y(n_3063)
);

AOI21xp5_ASAP7_75t_L g3064 ( 
.A1(n_2980),
.A2(n_2250),
.B(n_2245),
.Y(n_3064)
);

NAND2xp5_ASAP7_75t_L g3065 ( 
.A(n_2812),
.B(n_2633),
.Y(n_3065)
);

INVx2_ASAP7_75t_L g3066 ( 
.A(n_2847),
.Y(n_3066)
);

BUFx3_ASAP7_75t_L g3067 ( 
.A(n_2739),
.Y(n_3067)
);

INVx1_ASAP7_75t_L g3068 ( 
.A(n_2732),
.Y(n_3068)
);

NAND2xp5_ASAP7_75t_L g3069 ( 
.A(n_2829),
.B(n_2832),
.Y(n_3069)
);

NAND2xp5_ASAP7_75t_SL g3070 ( 
.A(n_2757),
.B(n_2608),
.Y(n_3070)
);

NOR3xp33_ASAP7_75t_L g3071 ( 
.A(n_2831),
.B(n_2580),
.C(n_1090),
.Y(n_3071)
);

AOI21xp5_ASAP7_75t_L g3072 ( 
.A1(n_2868),
.A2(n_2329),
.B(n_2250),
.Y(n_3072)
);

INVx3_ASAP7_75t_L g3073 ( 
.A(n_2823),
.Y(n_3073)
);

NAND2xp5_ASAP7_75t_L g3074 ( 
.A(n_2835),
.B(n_2487),
.Y(n_3074)
);

NAND2xp5_ASAP7_75t_L g3075 ( 
.A(n_2837),
.B(n_2489),
.Y(n_3075)
);

INVx3_ASAP7_75t_L g3076 ( 
.A(n_2823),
.Y(n_3076)
);

INVxp67_ASAP7_75t_L g3077 ( 
.A(n_2911),
.Y(n_3077)
);

NAND2xp5_ASAP7_75t_L g3078 ( 
.A(n_2845),
.B(n_2852),
.Y(n_3078)
);

NAND2xp5_ASAP7_75t_L g3079 ( 
.A(n_2975),
.B(n_2490),
.Y(n_3079)
);

NOR2xp33_ASAP7_75t_L g3080 ( 
.A(n_2979),
.B(n_2424),
.Y(n_3080)
);

NAND2xp5_ASAP7_75t_L g3081 ( 
.A(n_2950),
.B(n_2494),
.Y(n_3081)
);

OAI21xp5_ASAP7_75t_L g3082 ( 
.A1(n_2830),
.A2(n_2513),
.B(n_2496),
.Y(n_3082)
);

OAI21xp5_ASAP7_75t_L g3083 ( 
.A1(n_2830),
.A2(n_2843),
.B(n_2776),
.Y(n_3083)
);

INVx3_ASAP7_75t_L g3084 ( 
.A(n_2865),
.Y(n_3084)
);

AOI21xp5_ASAP7_75t_L g3085 ( 
.A1(n_2868),
.A2(n_2329),
.B(n_2250),
.Y(n_3085)
);

NOR2xp67_ASAP7_75t_L g3086 ( 
.A(n_2754),
.B(n_2552),
.Y(n_3086)
);

AOI21xp5_ASAP7_75t_L g3087 ( 
.A1(n_2874),
.A2(n_2329),
.B(n_2513),
.Y(n_3087)
);

OR2x2_ASAP7_75t_L g3088 ( 
.A(n_2734),
.B(n_2402),
.Y(n_3088)
);

O2A1O1Ixp33_ASAP7_75t_L g3089 ( 
.A1(n_2977),
.A2(n_2495),
.B(n_2501),
.C(n_2499),
.Y(n_3089)
);

CKINVDCx10_ASAP7_75t_R g3090 ( 
.A(n_2794),
.Y(n_3090)
);

O2A1O1Ixp33_ASAP7_75t_SL g3091 ( 
.A1(n_2769),
.A2(n_2707),
.B(n_2710),
.C(n_2705),
.Y(n_3091)
);

AND2x2_ASAP7_75t_L g3092 ( 
.A(n_3007),
.B(n_2587),
.Y(n_3092)
);

A2O1A1Ixp33_ASAP7_75t_L g3093 ( 
.A1(n_2799),
.A2(n_2694),
.B(n_2719),
.C(n_2677),
.Y(n_3093)
);

NOR2xp33_ASAP7_75t_L g3094 ( 
.A(n_2736),
.B(n_2679),
.Y(n_3094)
);

NAND2xp5_ASAP7_75t_L g3095 ( 
.A(n_2853),
.B(n_2675),
.Y(n_3095)
);

NOR2xp33_ASAP7_75t_R g3096 ( 
.A(n_2783),
.B(n_2465),
.Y(n_3096)
);

INVx1_ASAP7_75t_SL g3097 ( 
.A(n_2734),
.Y(n_3097)
);

NOR2xp67_ASAP7_75t_L g3098 ( 
.A(n_2808),
.B(n_2762),
.Y(n_3098)
);

AOI21xp5_ASAP7_75t_L g3099 ( 
.A1(n_2874),
.A2(n_2329),
.B(n_2720),
.Y(n_3099)
);

OAI22xp5_ASAP7_75t_L g3100 ( 
.A1(n_2943),
.A2(n_2522),
.B1(n_2406),
.B2(n_2692),
.Y(n_3100)
);

NAND2xp5_ASAP7_75t_L g3101 ( 
.A(n_2766),
.B(n_2676),
.Y(n_3101)
);

NAND2x1_ASAP7_75t_L g3102 ( 
.A(n_3005),
.B(n_2952),
.Y(n_3102)
);

NAND2xp5_ASAP7_75t_SL g3103 ( 
.A(n_2854),
.B(n_2690),
.Y(n_3103)
);

AOI21x1_ASAP7_75t_L g3104 ( 
.A1(n_2758),
.A2(n_2683),
.B(n_2678),
.Y(n_3104)
);

NOR2xp33_ASAP7_75t_L g3105 ( 
.A(n_2838),
.B(n_2887),
.Y(n_3105)
);

AND2x2_ASAP7_75t_SL g3106 ( 
.A(n_2778),
.B(n_2665),
.Y(n_3106)
);

NAND2xp5_ASAP7_75t_L g3107 ( 
.A(n_2957),
.B(n_2684),
.Y(n_3107)
);

INVx1_ASAP7_75t_L g3108 ( 
.A(n_2740),
.Y(n_3108)
);

NAND2xp5_ASAP7_75t_L g3109 ( 
.A(n_2985),
.B(n_2695),
.Y(n_3109)
);

AOI21x1_ASAP7_75t_L g3110 ( 
.A1(n_2813),
.A2(n_2699),
.B(n_2696),
.Y(n_3110)
);

INVx2_ASAP7_75t_L g3111 ( 
.A(n_2849),
.Y(n_3111)
);

AOI22xp5_ASAP7_75t_L g3112 ( 
.A1(n_2775),
.A2(n_2645),
.B1(n_2468),
.B2(n_2630),
.Y(n_3112)
);

INVx3_ASAP7_75t_L g3113 ( 
.A(n_3005),
.Y(n_3113)
);

HB1xp67_ASAP7_75t_L g3114 ( 
.A(n_2792),
.Y(n_3114)
);

NAND2xp5_ASAP7_75t_L g3115 ( 
.A(n_2985),
.B(n_2701),
.Y(n_3115)
);

CKINVDCx5p33_ASAP7_75t_R g3116 ( 
.A(n_2944),
.Y(n_3116)
);

NAND2xp5_ASAP7_75t_L g3117 ( 
.A(n_2914),
.B(n_2702),
.Y(n_3117)
);

NAND2x1p5_ASAP7_75t_L g3118 ( 
.A(n_2969),
.B(n_2804),
.Y(n_3118)
);

OAI21xp5_ASAP7_75t_L g3119 ( 
.A1(n_2843),
.A2(n_2648),
.B(n_2704),
.Y(n_3119)
);

AOI21xp5_ASAP7_75t_L g3120 ( 
.A1(n_2894),
.A2(n_2279),
.B(n_2344),
.Y(n_3120)
);

AND2x2_ASAP7_75t_L g3121 ( 
.A(n_2896),
.B(n_1307),
.Y(n_3121)
);

NOR2xp33_ASAP7_75t_L g3122 ( 
.A(n_2933),
.B(n_2793),
.Y(n_3122)
);

NAND2xp5_ASAP7_75t_L g3123 ( 
.A(n_2881),
.B(n_2715),
.Y(n_3123)
);

INVx2_ASAP7_75t_L g3124 ( 
.A(n_2850),
.Y(n_3124)
);

INVx1_ASAP7_75t_L g3125 ( 
.A(n_2743),
.Y(n_3125)
);

AOI21xp5_ASAP7_75t_L g3126 ( 
.A1(n_2894),
.A2(n_2279),
.B(n_2344),
.Y(n_3126)
);

NAND2xp5_ASAP7_75t_SL g3127 ( 
.A(n_2797),
.B(n_2457),
.Y(n_3127)
);

INVx3_ASAP7_75t_L g3128 ( 
.A(n_2952),
.Y(n_3128)
);

AND2x2_ASAP7_75t_SL g3129 ( 
.A(n_2778),
.B(n_2721),
.Y(n_3129)
);

NAND2xp5_ASAP7_75t_L g3130 ( 
.A(n_2981),
.B(n_2991),
.Y(n_3130)
);

O2A1O1Ixp5_ASAP7_75t_L g3131 ( 
.A1(n_2773),
.A2(n_2722),
.B(n_2150),
.C(n_2152),
.Y(n_3131)
);

O2A1O1Ixp33_ASAP7_75t_L g3132 ( 
.A1(n_2738),
.A2(n_1311),
.B(n_1308),
.C(n_1091),
.Y(n_3132)
);

INVx3_ASAP7_75t_L g3133 ( 
.A(n_2952),
.Y(n_3133)
);

BUFx6f_ASAP7_75t_L g3134 ( 
.A(n_2804),
.Y(n_3134)
);

AOI21xp5_ASAP7_75t_L g3135 ( 
.A1(n_2741),
.A2(n_2279),
.B(n_2344),
.Y(n_3135)
);

AND2x2_ASAP7_75t_L g3136 ( 
.A(n_2844),
.B(n_1084),
.Y(n_3136)
);

A2O1A1Ixp33_ASAP7_75t_L g3137 ( 
.A1(n_2781),
.A2(n_2532),
.B(n_2717),
.C(n_2688),
.Y(n_3137)
);

O2A1O1Ixp5_ASAP7_75t_L g3138 ( 
.A1(n_2746),
.A2(n_2152),
.B(n_2153),
.C(n_2144),
.Y(n_3138)
);

AOI22xp5_ASAP7_75t_L g3139 ( 
.A1(n_2841),
.A2(n_2630),
.B1(n_2037),
.B2(n_2522),
.Y(n_3139)
);

INVx1_ASAP7_75t_L g3140 ( 
.A(n_2745),
.Y(n_3140)
);

NAND2xp5_ASAP7_75t_L g3141 ( 
.A(n_3017),
.B(n_2532),
.Y(n_3141)
);

INVx1_ASAP7_75t_L g3142 ( 
.A(n_2759),
.Y(n_3142)
);

NAND2xp5_ASAP7_75t_L g3143 ( 
.A(n_2741),
.B(n_2406),
.Y(n_3143)
);

NAND2xp5_ASAP7_75t_L g3144 ( 
.A(n_2947),
.B(n_2034),
.Y(n_3144)
);

INVx1_ASAP7_75t_L g3145 ( 
.A(n_2761),
.Y(n_3145)
);

INVx2_ASAP7_75t_L g3146 ( 
.A(n_2872),
.Y(n_3146)
);

NOR2xp33_ASAP7_75t_L g3147 ( 
.A(n_2771),
.B(n_2285),
.Y(n_3147)
);

OAI22xp5_ASAP7_75t_L g3148 ( 
.A1(n_2840),
.A2(n_2271),
.B1(n_2282),
.B2(n_2260),
.Y(n_3148)
);

AOI21xp5_ASAP7_75t_L g3149 ( 
.A1(n_2997),
.A2(n_2279),
.B(n_2344),
.Y(n_3149)
);

OAI22xp5_ASAP7_75t_L g3150 ( 
.A1(n_2723),
.A2(n_3004),
.B1(n_2811),
.B2(n_2968),
.Y(n_3150)
);

NOR3xp33_ASAP7_75t_L g3151 ( 
.A(n_2805),
.B(n_1093),
.C(n_1092),
.Y(n_3151)
);

NAND2xp5_ASAP7_75t_L g3152 ( 
.A(n_2947),
.B(n_2038),
.Y(n_3152)
);

NAND2xp5_ASAP7_75t_SL g3153 ( 
.A(n_2846),
.B(n_2446),
.Y(n_3153)
);

OAI321xp33_ASAP7_75t_L g3154 ( 
.A1(n_2912),
.A2(n_1100),
.A3(n_1097),
.B1(n_1102),
.B2(n_1098),
.C(n_1096),
.Y(n_3154)
);

O2A1O1Ixp33_ASAP7_75t_L g3155 ( 
.A1(n_2802),
.A2(n_1106),
.B(n_1107),
.C(n_1105),
.Y(n_3155)
);

OAI21xp5_ASAP7_75t_L g3156 ( 
.A1(n_3015),
.A2(n_2039),
.B(n_2153),
.Y(n_3156)
);

NAND2xp5_ASAP7_75t_L g3157 ( 
.A(n_2951),
.B(n_2039),
.Y(n_3157)
);

NOR2xp33_ASAP7_75t_L g3158 ( 
.A(n_3010),
.B(n_2285),
.Y(n_3158)
);

NAND2xp5_ASAP7_75t_L g3159 ( 
.A(n_2951),
.B(n_2157),
.Y(n_3159)
);

BUFx2_ASAP7_75t_L g3160 ( 
.A(n_2789),
.Y(n_3160)
);

BUFx4f_ASAP7_75t_L g3161 ( 
.A(n_2804),
.Y(n_3161)
);

OAI22xp5_ASAP7_75t_L g3162 ( 
.A1(n_3011),
.A2(n_2271),
.B1(n_2282),
.B2(n_2260),
.Y(n_3162)
);

INVx2_ASAP7_75t_L g3163 ( 
.A(n_2873),
.Y(n_3163)
);

OAI21xp5_ASAP7_75t_L g3164 ( 
.A1(n_3015),
.A2(n_2159),
.B(n_2157),
.Y(n_3164)
);

NAND2xp5_ASAP7_75t_L g3165 ( 
.A(n_2972),
.B(n_2159),
.Y(n_3165)
);

INVx1_ASAP7_75t_L g3166 ( 
.A(n_2763),
.Y(n_3166)
);

INVx1_ASAP7_75t_L g3167 ( 
.A(n_2770),
.Y(n_3167)
);

AOI21xp5_ASAP7_75t_L g3168 ( 
.A1(n_2997),
.A2(n_2279),
.B(n_2344),
.Y(n_3168)
);

NOR2xp33_ASAP7_75t_L g3169 ( 
.A(n_2879),
.B(n_2290),
.Y(n_3169)
);

AOI21xp5_ASAP7_75t_L g3170 ( 
.A1(n_2972),
.A2(n_2344),
.B(n_2032),
.Y(n_3170)
);

INVx2_ASAP7_75t_L g3171 ( 
.A(n_2875),
.Y(n_3171)
);

NAND2xp5_ASAP7_75t_L g3172 ( 
.A(n_2819),
.B(n_2162),
.Y(n_3172)
);

NOR2xp33_ASAP7_75t_L g3173 ( 
.A(n_3014),
.B(n_2290),
.Y(n_3173)
);

INVx1_ASAP7_75t_L g3174 ( 
.A(n_2780),
.Y(n_3174)
);

INVx1_ASAP7_75t_L g3175 ( 
.A(n_2782),
.Y(n_3175)
);

INVx2_ASAP7_75t_L g3176 ( 
.A(n_2876),
.Y(n_3176)
);

INVx1_ASAP7_75t_L g3177 ( 
.A(n_2800),
.Y(n_3177)
);

OAI21xp5_ASAP7_75t_L g3178 ( 
.A1(n_2791),
.A2(n_2165),
.B(n_2162),
.Y(n_3178)
);

CKINVDCx20_ASAP7_75t_R g3179 ( 
.A(n_3016),
.Y(n_3179)
);

NOR2xp33_ASAP7_75t_SL g3180 ( 
.A(n_2860),
.B(n_2030),
.Y(n_3180)
);

NAND2xp5_ASAP7_75t_L g3181 ( 
.A(n_2821),
.B(n_2760),
.Y(n_3181)
);

NAND2xp33_ASAP7_75t_L g3182 ( 
.A(n_2916),
.B(n_2037),
.Y(n_3182)
);

AND2x2_ASAP7_75t_SL g3183 ( 
.A(n_2742),
.B(n_2165),
.Y(n_3183)
);

CKINVDCx6p67_ASAP7_75t_R g3184 ( 
.A(n_2794),
.Y(n_3184)
);

INVx1_ASAP7_75t_L g3185 ( 
.A(n_2816),
.Y(n_3185)
);

NAND2xp5_ASAP7_75t_L g3186 ( 
.A(n_2772),
.B(n_2168),
.Y(n_3186)
);

AOI21xp5_ASAP7_75t_L g3187 ( 
.A1(n_2994),
.A2(n_2032),
.B(n_2030),
.Y(n_3187)
);

OAI21xp33_ASAP7_75t_L g3188 ( 
.A1(n_2899),
.A2(n_620),
.B(n_613),
.Y(n_3188)
);

A2O1A1Ixp33_ASAP7_75t_L g3189 ( 
.A1(n_2913),
.A2(n_2282),
.B(n_2287),
.C(n_2271),
.Y(n_3189)
);

AOI21xp5_ASAP7_75t_L g3190 ( 
.A1(n_3000),
.A2(n_2292),
.B(n_2287),
.Y(n_3190)
);

INVx1_ASAP7_75t_L g3191 ( 
.A(n_2820),
.Y(n_3191)
);

INVx1_ASAP7_75t_L g3192 ( 
.A(n_2833),
.Y(n_3192)
);

OAI21x1_ASAP7_75t_L g3193 ( 
.A1(n_2857),
.A2(n_2148),
.B(n_2126),
.Y(n_3193)
);

AND2x2_ASAP7_75t_L g3194 ( 
.A(n_2921),
.B(n_1108),
.Y(n_3194)
);

NAND2xp5_ASAP7_75t_L g3195 ( 
.A(n_2856),
.B(n_2168),
.Y(n_3195)
);

AOI22xp5_ASAP7_75t_L g3196 ( 
.A1(n_2851),
.A2(n_1822),
.B1(n_1831),
.B2(n_1818),
.Y(n_3196)
);

NAND2xp5_ASAP7_75t_L g3197 ( 
.A(n_2856),
.B(n_2172),
.Y(n_3197)
);

INVx2_ASAP7_75t_L g3198 ( 
.A(n_2877),
.Y(n_3198)
);

NAND2xp5_ASAP7_75t_L g3199 ( 
.A(n_2836),
.B(n_2172),
.Y(n_3199)
);

OAI21xp5_ASAP7_75t_L g3200 ( 
.A1(n_2882),
.A2(n_2175),
.B(n_2174),
.Y(n_3200)
);

INVx1_ASAP7_75t_L g3201 ( 
.A(n_2839),
.Y(n_3201)
);

INVx4_ASAP7_75t_L g3202 ( 
.A(n_2822),
.Y(n_3202)
);

NAND2xp5_ASAP7_75t_L g3203 ( 
.A(n_2858),
.B(n_2174),
.Y(n_3203)
);

NAND2xp5_ASAP7_75t_L g3204 ( 
.A(n_2884),
.B(n_2175),
.Y(n_3204)
);

AOI21xp5_ASAP7_75t_L g3205 ( 
.A1(n_3000),
.A2(n_2292),
.B(n_2287),
.Y(n_3205)
);

NOR2xp67_ASAP7_75t_L g3206 ( 
.A(n_2998),
.B(n_2177),
.Y(n_3206)
);

INVx3_ASAP7_75t_L g3207 ( 
.A(n_2822),
.Y(n_3207)
);

INVx2_ASAP7_75t_L g3208 ( 
.A(n_2880),
.Y(n_3208)
);

NAND2xp5_ASAP7_75t_L g3209 ( 
.A(n_2901),
.B(n_2177),
.Y(n_3209)
);

NAND2xp5_ASAP7_75t_L g3210 ( 
.A(n_2906),
.B(n_2178),
.Y(n_3210)
);

INVx1_ASAP7_75t_L g3211 ( 
.A(n_2910),
.Y(n_3211)
);

INVx3_ASAP7_75t_L g3212 ( 
.A(n_2969),
.Y(n_3212)
);

OAI21xp5_ASAP7_75t_L g3213 ( 
.A1(n_2964),
.A2(n_2179),
.B(n_2178),
.Y(n_3213)
);

NAND2xp5_ASAP7_75t_L g3214 ( 
.A(n_2920),
.B(n_2179),
.Y(n_3214)
);

INVx1_ASAP7_75t_L g3215 ( 
.A(n_2925),
.Y(n_3215)
);

NOR2xp33_ASAP7_75t_L g3216 ( 
.A(n_2863),
.B(n_2296),
.Y(n_3216)
);

AOI22xp5_ASAP7_75t_L g3217 ( 
.A1(n_2936),
.A2(n_1844),
.B1(n_1848),
.B2(n_1834),
.Y(n_3217)
);

INVx2_ASAP7_75t_L g3218 ( 
.A(n_2898),
.Y(n_3218)
);

AO21x1_ASAP7_75t_L g3219 ( 
.A1(n_2982),
.A2(n_1999),
.B(n_1983),
.Y(n_3219)
);

OAI22xp5_ASAP7_75t_L g3220 ( 
.A1(n_2904),
.A2(n_2300),
.B1(n_2292),
.B2(n_2373),
.Y(n_3220)
);

AOI21xp5_ASAP7_75t_L g3221 ( 
.A1(n_2825),
.A2(n_2791),
.B(n_2993),
.Y(n_3221)
);

OR2x6_ASAP7_75t_L g3222 ( 
.A(n_2930),
.B(n_2192),
.Y(n_3222)
);

NAND2xp5_ASAP7_75t_L g3223 ( 
.A(n_2942),
.B(n_2192),
.Y(n_3223)
);

AOI21xp5_ASAP7_75t_L g3224 ( 
.A1(n_2825),
.A2(n_2300),
.B(n_2297),
.Y(n_3224)
);

AOI21xp5_ASAP7_75t_L g3225 ( 
.A1(n_2999),
.A2(n_2300),
.B(n_2297),
.Y(n_3225)
);

NAND2xp5_ASAP7_75t_L g3226 ( 
.A(n_3057),
.B(n_2929),
.Y(n_3226)
);

AOI22xp5_ASAP7_75t_L g3227 ( 
.A1(n_3052),
.A2(n_2885),
.B1(n_2893),
.B2(n_2948),
.Y(n_3227)
);

NAND3xp33_ASAP7_75t_SL g3228 ( 
.A(n_3071),
.B(n_2960),
.C(n_2895),
.Y(n_3228)
);

AOI21xp5_ASAP7_75t_L g3229 ( 
.A1(n_3023),
.A2(n_3036),
.B(n_3025),
.Y(n_3229)
);

AOI21xp5_ASAP7_75t_L g3230 ( 
.A1(n_3078),
.A2(n_2999),
.B(n_2834),
.Y(n_3230)
);

AOI21xp5_ASAP7_75t_L g3231 ( 
.A1(n_3031),
.A2(n_2834),
.B(n_2807),
.Y(n_3231)
);

AOI22xp5_ASAP7_75t_L g3232 ( 
.A1(n_3106),
.A2(n_3070),
.B1(n_3094),
.B2(n_3029),
.Y(n_3232)
);

NAND2xp5_ASAP7_75t_SL g3233 ( 
.A(n_3062),
.B(n_3130),
.Y(n_3233)
);

INVx1_ASAP7_75t_SL g3234 ( 
.A(n_3045),
.Y(n_3234)
);

INVx2_ASAP7_75t_L g3235 ( 
.A(n_3022),
.Y(n_3235)
);

INVx4_ASAP7_75t_L g3236 ( 
.A(n_3161),
.Y(n_3236)
);

INVx1_ASAP7_75t_L g3237 ( 
.A(n_3030),
.Y(n_3237)
);

NAND2xp5_ASAP7_75t_L g3238 ( 
.A(n_3069),
.B(n_2940),
.Y(n_3238)
);

NOR2xp33_ASAP7_75t_L g3239 ( 
.A(n_3077),
.B(n_2891),
.Y(n_3239)
);

AOI22xp5_ASAP7_75t_L g3240 ( 
.A1(n_3105),
.A2(n_2970),
.B1(n_2801),
.B2(n_3008),
.Y(n_3240)
);

AOI21xp5_ASAP7_75t_L g3241 ( 
.A1(n_3037),
.A2(n_2807),
.B(n_2857),
.Y(n_3241)
);

NOR2xp33_ASAP7_75t_L g3242 ( 
.A(n_3043),
.B(n_3002),
.Y(n_3242)
);

AOI21xp5_ASAP7_75t_L g3243 ( 
.A1(n_3087),
.A2(n_2886),
.B(n_2969),
.Y(n_3243)
);

NAND2xp5_ASAP7_75t_SL g3244 ( 
.A(n_3122),
.B(n_2931),
.Y(n_3244)
);

NAND2xp5_ASAP7_75t_L g3245 ( 
.A(n_3050),
.B(n_2965),
.Y(n_3245)
);

NAND2xp5_ASAP7_75t_SL g3246 ( 
.A(n_3117),
.B(n_2919),
.Y(n_3246)
);

INVx1_ASAP7_75t_L g3247 ( 
.A(n_3068),
.Y(n_3247)
);

NAND2xp5_ASAP7_75t_L g3248 ( 
.A(n_3034),
.B(n_3136),
.Y(n_3248)
);

NAND2xp5_ASAP7_75t_SL g3249 ( 
.A(n_3026),
.B(n_2861),
.Y(n_3249)
);

AOI21xp5_ASAP7_75t_L g3250 ( 
.A1(n_3180),
.A2(n_3085),
.B(n_3072),
.Y(n_3250)
);

AOI21x1_ASAP7_75t_L g3251 ( 
.A1(n_3110),
.A2(n_3221),
.B(n_3061),
.Y(n_3251)
);

AOI21xp5_ASAP7_75t_L g3252 ( 
.A1(n_3180),
.A2(n_2886),
.B(n_2967),
.Y(n_3252)
);

NAND2xp5_ASAP7_75t_L g3253 ( 
.A(n_3027),
.B(n_2966),
.Y(n_3253)
);

NAND2xp5_ASAP7_75t_L g3254 ( 
.A(n_3028),
.B(n_2809),
.Y(n_3254)
);

NAND2xp5_ASAP7_75t_SL g3255 ( 
.A(n_3046),
.B(n_2861),
.Y(n_3255)
);

AOI21xp5_ASAP7_75t_L g3256 ( 
.A1(n_3144),
.A2(n_2883),
.B(n_2953),
.Y(n_3256)
);

INVx1_ASAP7_75t_L g3257 ( 
.A(n_3108),
.Y(n_3257)
);

INVxp67_ASAP7_75t_SL g3258 ( 
.A(n_3051),
.Y(n_3258)
);

INVx2_ASAP7_75t_L g3259 ( 
.A(n_3040),
.Y(n_3259)
);

AOI21xp5_ASAP7_75t_L g3260 ( 
.A1(n_3152),
.A2(n_2982),
.B(n_2909),
.Y(n_3260)
);

AOI21xp5_ASAP7_75t_L g3261 ( 
.A1(n_3157),
.A2(n_2755),
.B(n_2871),
.Y(n_3261)
);

A2O1A1Ixp33_ASAP7_75t_L g3262 ( 
.A1(n_3035),
.A2(n_2892),
.B(n_2897),
.C(n_2806),
.Y(n_3262)
);

NAND2xp5_ASAP7_75t_L g3263 ( 
.A(n_3181),
.B(n_3109),
.Y(n_3263)
);

NOR2xp33_ASAP7_75t_L g3264 ( 
.A(n_3039),
.B(n_2932),
.Y(n_3264)
);

NOR2xp67_ASAP7_75t_SL g3265 ( 
.A(n_3154),
.B(n_3116),
.Y(n_3265)
);

INVx2_ASAP7_75t_L g3266 ( 
.A(n_3066),
.Y(n_3266)
);

O2A1O1Ixp33_ASAP7_75t_SL g3267 ( 
.A1(n_3153),
.A2(n_2864),
.B(n_2870),
.C(n_2922),
.Y(n_3267)
);

NAND2xp5_ASAP7_75t_L g3268 ( 
.A(n_3115),
.B(n_3019),
.Y(n_3268)
);

AOI21xp5_ASAP7_75t_L g3269 ( 
.A1(n_3038),
.A2(n_2978),
.B(n_2971),
.Y(n_3269)
);

NAND2xp5_ASAP7_75t_L g3270 ( 
.A(n_3095),
.B(n_2949),
.Y(n_3270)
);

NAND2xp5_ASAP7_75t_SL g3271 ( 
.A(n_3045),
.B(n_2861),
.Y(n_3271)
);

INVx2_ASAP7_75t_L g3272 ( 
.A(n_3111),
.Y(n_3272)
);

AOI21xp5_ASAP7_75t_L g3273 ( 
.A1(n_3120),
.A2(n_3012),
.B(n_2992),
.Y(n_3273)
);

AND2x4_ASAP7_75t_L g3274 ( 
.A(n_3207),
.B(n_2867),
.Y(n_3274)
);

NAND2xp5_ASAP7_75t_L g3275 ( 
.A(n_3074),
.B(n_2989),
.Y(n_3275)
);

OAI22xp5_ASAP7_75t_L g3276 ( 
.A1(n_3196),
.A2(n_2867),
.B1(n_3001),
.B2(n_2990),
.Y(n_3276)
);

AOI21xp5_ASAP7_75t_L g3277 ( 
.A1(n_3126),
.A2(n_2988),
.B(n_2934),
.Y(n_3277)
);

INVx2_ASAP7_75t_SL g3278 ( 
.A(n_3067),
.Y(n_3278)
);

CKINVDCx8_ASAP7_75t_R g3279 ( 
.A(n_3090),
.Y(n_3279)
);

INVxp67_ASAP7_75t_L g3280 ( 
.A(n_3114),
.Y(n_3280)
);

O2A1O1Ixp5_ASAP7_75t_L g3281 ( 
.A1(n_3150),
.A2(n_2927),
.B(n_2888),
.C(n_2974),
.Y(n_3281)
);

AOI21xp5_ASAP7_75t_L g3282 ( 
.A1(n_3056),
.A2(n_2986),
.B(n_2996),
.Y(n_3282)
);

AND2x2_ASAP7_75t_L g3283 ( 
.A(n_3194),
.B(n_2955),
.Y(n_3283)
);

AOI21xp5_ASAP7_75t_L g3284 ( 
.A1(n_3065),
.A2(n_2986),
.B(n_3009),
.Y(n_3284)
);

OR2x2_ASAP7_75t_L g3285 ( 
.A(n_3097),
.B(n_3088),
.Y(n_3285)
);

AND2x2_ASAP7_75t_L g3286 ( 
.A(n_3097),
.B(n_3121),
.Y(n_3286)
);

AOI21xp5_ASAP7_75t_L g3287 ( 
.A1(n_3044),
.A2(n_2986),
.B(n_2889),
.Y(n_3287)
);

AO21x1_ASAP7_75t_L g3288 ( 
.A1(n_3089),
.A2(n_3033),
.B(n_3053),
.Y(n_3288)
);

AOI21xp5_ASAP7_75t_L g3289 ( 
.A1(n_3047),
.A2(n_2878),
.B(n_2924),
.Y(n_3289)
);

NAND2xp5_ASAP7_75t_SL g3290 ( 
.A(n_3081),
.B(n_2903),
.Y(n_3290)
);

OAI21xp5_ASAP7_75t_L g3291 ( 
.A1(n_3101),
.A2(n_2788),
.B(n_2963),
.Y(n_3291)
);

AND2x2_ASAP7_75t_L g3292 ( 
.A(n_3092),
.B(n_2955),
.Y(n_3292)
);

INVx5_ASAP7_75t_L g3293 ( 
.A(n_3058),
.Y(n_3293)
);

AND2x2_ASAP7_75t_L g3294 ( 
.A(n_3158),
.B(n_2955),
.Y(n_3294)
);

O2A1O1Ixp33_ASAP7_75t_L g3295 ( 
.A1(n_3154),
.A2(n_2938),
.B(n_2962),
.C(n_2827),
.Y(n_3295)
);

INVxp67_ASAP7_75t_SL g3296 ( 
.A(n_3107),
.Y(n_3296)
);

OAI22xp5_ASAP7_75t_L g3297 ( 
.A1(n_3112),
.A2(n_3216),
.B1(n_3139),
.B2(n_3123),
.Y(n_3297)
);

AND2x2_ASAP7_75t_L g3298 ( 
.A(n_3173),
.B(n_2903),
.Y(n_3298)
);

O2A1O1Ixp33_ASAP7_75t_L g3299 ( 
.A1(n_3188),
.A2(n_2915),
.B(n_2917),
.C(n_3003),
.Y(n_3299)
);

NAND2xp5_ASAP7_75t_L g3300 ( 
.A(n_3075),
.B(n_3013),
.Y(n_3300)
);

AOI21xp5_ASAP7_75t_L g3301 ( 
.A1(n_3099),
.A2(n_2945),
.B(n_2926),
.Y(n_3301)
);

INVx2_ASAP7_75t_L g3302 ( 
.A(n_3124),
.Y(n_3302)
);

NAND2xp5_ASAP7_75t_L g3303 ( 
.A(n_3042),
.B(n_2903),
.Y(n_3303)
);

AOI21xp5_ASAP7_75t_L g3304 ( 
.A1(n_3064),
.A2(n_2935),
.B(n_2923),
.Y(n_3304)
);

AND2x2_ASAP7_75t_L g3305 ( 
.A(n_3147),
.B(n_2848),
.Y(n_3305)
);

AOI21xp5_ASAP7_75t_L g3306 ( 
.A1(n_3170),
.A2(n_3187),
.B(n_3168),
.Y(n_3306)
);

NAND2xp5_ASAP7_75t_SL g3307 ( 
.A(n_3206),
.B(n_2959),
.Y(n_3307)
);

NAND2xp5_ASAP7_75t_SL g3308 ( 
.A(n_3049),
.B(n_3169),
.Y(n_3308)
);

NAND2xp5_ASAP7_75t_L g3309 ( 
.A(n_3188),
.B(n_2959),
.Y(n_3309)
);

AOI21xp5_ASAP7_75t_L g3310 ( 
.A1(n_3149),
.A2(n_2946),
.B(n_2937),
.Y(n_3310)
);

INVx2_ASAP7_75t_L g3311 ( 
.A(n_3146),
.Y(n_3311)
);

NOR2xp33_ASAP7_75t_L g3312 ( 
.A(n_3080),
.B(n_2905),
.Y(n_3312)
);

AOI21xp5_ASAP7_75t_L g3313 ( 
.A1(n_3135),
.A2(n_2987),
.B(n_2973),
.Y(n_3313)
);

NOR2x1_ASAP7_75t_L g3314 ( 
.A(n_3086),
.B(n_2867),
.Y(n_3314)
);

NAND2xp5_ASAP7_75t_SL g3315 ( 
.A(n_3163),
.B(n_2900),
.Y(n_3315)
);

NAND2xp5_ASAP7_75t_L g3316 ( 
.A(n_3171),
.B(n_2941),
.Y(n_3316)
);

OAI22xp5_ASAP7_75t_L g3317 ( 
.A1(n_3217),
.A2(n_2767),
.B1(n_2918),
.B2(n_2902),
.Y(n_3317)
);

AND2x4_ASAP7_75t_L g3318 ( 
.A(n_3207),
.B(n_2767),
.Y(n_3318)
);

NAND2xp5_ASAP7_75t_L g3319 ( 
.A(n_3176),
.B(n_2976),
.Y(n_3319)
);

AOI21x1_ASAP7_75t_L g3320 ( 
.A1(n_3104),
.A2(n_2201),
.B(n_2196),
.Y(n_3320)
);

NAND2xp5_ASAP7_75t_SL g3321 ( 
.A(n_3198),
.B(n_2939),
.Y(n_3321)
);

BUFx2_ASAP7_75t_L g3322 ( 
.A(n_3058),
.Y(n_3322)
);

AOI21xp5_ASAP7_75t_L g3323 ( 
.A1(n_3083),
.A2(n_2767),
.B(n_2907),
.Y(n_3323)
);

NAND2xp5_ASAP7_75t_L g3324 ( 
.A(n_3208),
.B(n_3006),
.Y(n_3324)
);

NAND3xp33_ASAP7_75t_L g3325 ( 
.A(n_3151),
.B(n_878),
.C(n_622),
.Y(n_3325)
);

NOR2xp33_ASAP7_75t_L g3326 ( 
.A(n_3103),
.B(n_2862),
.Y(n_3326)
);

INVx2_ASAP7_75t_L g3327 ( 
.A(n_3218),
.Y(n_3327)
);

INVx2_ASAP7_75t_L g3328 ( 
.A(n_3125),
.Y(n_3328)
);

NOR3xp33_ASAP7_75t_L g3329 ( 
.A(n_3182),
.B(n_1111),
.C(n_1109),
.Y(n_3329)
);

OAI22xp5_ASAP7_75t_L g3330 ( 
.A1(n_3129),
.A2(n_2956),
.B1(n_2983),
.B2(n_2961),
.Y(n_3330)
);

NAND2xp5_ASAP7_75t_L g3331 ( 
.A(n_3140),
.B(n_3018),
.Y(n_3331)
);

NOR3xp33_ASAP7_75t_L g3332 ( 
.A(n_3132),
.B(n_1113),
.C(n_1112),
.Y(n_3332)
);

INVx2_ASAP7_75t_L g3333 ( 
.A(n_3142),
.Y(n_3333)
);

CKINVDCx10_ASAP7_75t_R g3334 ( 
.A(n_3096),
.Y(n_3334)
);

AOI21xp5_ASAP7_75t_L g3335 ( 
.A1(n_3091),
.A2(n_2907),
.B(n_3020),
.Y(n_3335)
);

NAND2xp5_ASAP7_75t_L g3336 ( 
.A(n_3145),
.B(n_2726),
.Y(n_3336)
);

OAI21xp5_ASAP7_75t_L g3337 ( 
.A1(n_3127),
.A2(n_2737),
.B(n_2733),
.Y(n_3337)
);

OAI21xp5_ASAP7_75t_L g3338 ( 
.A1(n_3093),
.A2(n_2747),
.B(n_2744),
.Y(n_3338)
);

AOI21xp5_ASAP7_75t_L g3339 ( 
.A1(n_3041),
.A2(n_3224),
.B(n_3189),
.Y(n_3339)
);

NAND2xp5_ASAP7_75t_SL g3340 ( 
.A(n_3098),
.B(n_2916),
.Y(n_3340)
);

O2A1O1Ixp33_ASAP7_75t_L g3341 ( 
.A1(n_3063),
.A2(n_1117),
.B(n_1118),
.C(n_1116),
.Y(n_3341)
);

INVx2_ASAP7_75t_L g3342 ( 
.A(n_3166),
.Y(n_3342)
);

AOI22xp5_ASAP7_75t_L g3343 ( 
.A1(n_3055),
.A2(n_3100),
.B1(n_3143),
.B2(n_3167),
.Y(n_3343)
);

NOR2xp33_ASAP7_75t_L g3344 ( 
.A(n_3179),
.B(n_2908),
.Y(n_3344)
);

INVx1_ASAP7_75t_L g3345 ( 
.A(n_3174),
.Y(n_3345)
);

O2A1O1Ixp33_ASAP7_75t_SL g3346 ( 
.A1(n_3102),
.A2(n_2750),
.B(n_2753),
.C(n_2749),
.Y(n_3346)
);

OAI21x1_ASAP7_75t_L g3347 ( 
.A1(n_3193),
.A2(n_2148),
.B(n_2126),
.Y(n_3347)
);

AO21x1_ASAP7_75t_L g3348 ( 
.A1(n_3220),
.A2(n_2796),
.B(n_2768),
.Y(n_3348)
);

A2O1A1Ixp33_ASAP7_75t_SL g3349 ( 
.A1(n_3082),
.A2(n_2803),
.B(n_2810),
.C(n_2798),
.Y(n_3349)
);

INVx2_ASAP7_75t_L g3350 ( 
.A(n_3175),
.Y(n_3350)
);

NOR2xp33_ASAP7_75t_L g3351 ( 
.A(n_3160),
.B(n_2984),
.Y(n_3351)
);

INVx1_ASAP7_75t_L g3352 ( 
.A(n_3177),
.Y(n_3352)
);

INVx1_ASAP7_75t_L g3353 ( 
.A(n_3185),
.Y(n_3353)
);

INVx1_ASAP7_75t_L g3354 ( 
.A(n_3191),
.Y(n_3354)
);

OAI22xp5_ASAP7_75t_L g3355 ( 
.A1(n_3183),
.A2(n_3079),
.B1(n_3215),
.B2(n_3211),
.Y(n_3355)
);

NOR2xp33_ASAP7_75t_SL g3356 ( 
.A(n_3184),
.B(n_2916),
.Y(n_3356)
);

AOI21xp5_ASAP7_75t_L g3357 ( 
.A1(n_3024),
.A2(n_2928),
.B(n_2916),
.Y(n_3357)
);

O2A1O1Ixp33_ASAP7_75t_L g3358 ( 
.A1(n_3155),
.A2(n_1122),
.B(n_1123),
.C(n_1121),
.Y(n_3358)
);

AOI21xp5_ASAP7_75t_L g3359 ( 
.A1(n_3024),
.A2(n_2928),
.B(n_2916),
.Y(n_3359)
);

INVx3_ASAP7_75t_L g3360 ( 
.A(n_3060),
.Y(n_3360)
);

OAI22xp5_ASAP7_75t_L g3361 ( 
.A1(n_3192),
.A2(n_2817),
.B1(n_2815),
.B2(n_883),
.Y(n_3361)
);

INVx1_ASAP7_75t_SL g3362 ( 
.A(n_3058),
.Y(n_3362)
);

BUFx2_ASAP7_75t_L g3363 ( 
.A(n_3059),
.Y(n_3363)
);

INVx4_ASAP7_75t_L g3364 ( 
.A(n_3161),
.Y(n_3364)
);

INVx2_ASAP7_75t_L g3365 ( 
.A(n_3201),
.Y(n_3365)
);

INVx2_ASAP7_75t_SL g3366 ( 
.A(n_3059),
.Y(n_3366)
);

INVx4_ASAP7_75t_L g3367 ( 
.A(n_3059),
.Y(n_3367)
);

NAND2xp5_ASAP7_75t_L g3368 ( 
.A(n_3141),
.B(n_878),
.Y(n_3368)
);

O2A1O1Ixp33_ASAP7_75t_L g3369 ( 
.A1(n_3137),
.A2(n_1129),
.B(n_1131),
.C(n_1125),
.Y(n_3369)
);

INVx1_ASAP7_75t_L g3370 ( 
.A(n_3199),
.Y(n_3370)
);

AOI21xp5_ASAP7_75t_L g3371 ( 
.A1(n_3082),
.A2(n_2928),
.B(n_2201),
.Y(n_3371)
);

NAND2xp5_ASAP7_75t_L g3372 ( 
.A(n_3172),
.B(n_883),
.Y(n_3372)
);

INVx2_ASAP7_75t_L g3373 ( 
.A(n_3203),
.Y(n_3373)
);

INVx3_ASAP7_75t_L g3374 ( 
.A(n_3060),
.Y(n_3374)
);

AOI21xp5_ASAP7_75t_L g3375 ( 
.A1(n_3195),
.A2(n_2928),
.B(n_2203),
.Y(n_3375)
);

A2O1A1Ixp33_ASAP7_75t_L g3376 ( 
.A1(n_3119),
.A2(n_2301),
.B(n_2303),
.C(n_2296),
.Y(n_3376)
);

NAND2x1p5_ASAP7_75t_L g3377 ( 
.A(n_3128),
.B(n_2126),
.Y(n_3377)
);

NOR2xp33_ASAP7_75t_L g3378 ( 
.A(n_3032),
.B(n_815),
.Y(n_3378)
);

AOI21xp5_ASAP7_75t_L g3379 ( 
.A1(n_3197),
.A2(n_3165),
.B(n_3159),
.Y(n_3379)
);

AOI21xp5_ASAP7_75t_L g3380 ( 
.A1(n_3213),
.A2(n_3156),
.B(n_3190),
.Y(n_3380)
);

NAND2xp5_ASAP7_75t_L g3381 ( 
.A(n_3204),
.B(n_884),
.Y(n_3381)
);

NAND2xp5_ASAP7_75t_L g3382 ( 
.A(n_3209),
.B(n_884),
.Y(n_3382)
);

O2A1O1Ixp33_ASAP7_75t_SL g3383 ( 
.A1(n_3048),
.A2(n_2301),
.B(n_2304),
.C(n_2303),
.Y(n_3383)
);

AOI21xp5_ASAP7_75t_L g3384 ( 
.A1(n_3156),
.A2(n_2928),
.B(n_2203),
.Y(n_3384)
);

OAI22xp5_ASAP7_75t_L g3385 ( 
.A1(n_3128),
.A2(n_887),
.B1(n_889),
.B2(n_885),
.Y(n_3385)
);

NAND2x1p5_ASAP7_75t_L g3386 ( 
.A(n_3133),
.B(n_2181),
.Y(n_3386)
);

NAND2xp5_ASAP7_75t_L g3387 ( 
.A(n_3210),
.B(n_885),
.Y(n_3387)
);

AOI21xp5_ASAP7_75t_L g3388 ( 
.A1(n_3205),
.A2(n_2211),
.B(n_2196),
.Y(n_3388)
);

NAND2xp5_ASAP7_75t_L g3389 ( 
.A(n_3214),
.B(n_887),
.Y(n_3389)
);

OAI22x1_ASAP7_75t_L g3390 ( 
.A1(n_3133),
.A2(n_891),
.B1(n_895),
.B2(n_889),
.Y(n_3390)
);

NAND2xp5_ASAP7_75t_L g3391 ( 
.A(n_3223),
.B(n_891),
.Y(n_3391)
);

INVx2_ASAP7_75t_L g3392 ( 
.A(n_3186),
.Y(n_3392)
);

NAND2xp5_ASAP7_75t_L g3393 ( 
.A(n_3202),
.B(n_3054),
.Y(n_3393)
);

AOI21xp5_ASAP7_75t_L g3394 ( 
.A1(n_3148),
.A2(n_2212),
.B(n_2211),
.Y(n_3394)
);

OAI22xp5_ASAP7_75t_L g3395 ( 
.A1(n_3222),
.A2(n_898),
.B1(n_901),
.B2(n_895),
.Y(n_3395)
);

INVx1_ASAP7_75t_L g3396 ( 
.A(n_3219),
.Y(n_3396)
);

AND2x4_ASAP7_75t_L g3397 ( 
.A(n_3202),
.B(n_2446),
.Y(n_3397)
);

BUFx2_ASAP7_75t_L g3398 ( 
.A(n_3134),
.Y(n_3398)
);

BUFx6f_ASAP7_75t_L g3399 ( 
.A(n_3134),
.Y(n_3399)
);

AOI21xp5_ASAP7_75t_L g3400 ( 
.A1(n_3200),
.A2(n_3178),
.B(n_3225),
.Y(n_3400)
);

INVx3_ASAP7_75t_L g3401 ( 
.A(n_3118),
.Y(n_3401)
);

INVx2_ASAP7_75t_L g3402 ( 
.A(n_3073),
.Y(n_3402)
);

AOI21xp5_ASAP7_75t_L g3403 ( 
.A1(n_3178),
.A2(n_2216),
.B(n_2212),
.Y(n_3403)
);

AOI21xp5_ASAP7_75t_L g3404 ( 
.A1(n_3164),
.A2(n_2222),
.B(n_2216),
.Y(n_3404)
);

AND2x2_ASAP7_75t_L g3405 ( 
.A(n_3134),
.B(n_1132),
.Y(n_3405)
);

AOI21xp5_ASAP7_75t_L g3406 ( 
.A1(n_3164),
.A2(n_2224),
.B(n_2222),
.Y(n_3406)
);

NOR2xp67_ASAP7_75t_L g3407 ( 
.A(n_3054),
.B(n_2224),
.Y(n_3407)
);

NAND2xp5_ASAP7_75t_L g3408 ( 
.A(n_3073),
.B(n_898),
.Y(n_3408)
);

NAND2xp5_ASAP7_75t_L g3409 ( 
.A(n_3076),
.B(n_901),
.Y(n_3409)
);

A2O1A1Ixp33_ASAP7_75t_SL g3410 ( 
.A1(n_3212),
.A2(n_2207),
.B(n_2209),
.C(n_2181),
.Y(n_3410)
);

BUFx8_ASAP7_75t_L g3411 ( 
.A(n_3222),
.Y(n_3411)
);

INVx2_ASAP7_75t_L g3412 ( 
.A(n_3076),
.Y(n_3412)
);

INVx4_ASAP7_75t_L g3413 ( 
.A(n_3118),
.Y(n_3413)
);

INVx5_ASAP7_75t_L g3414 ( 
.A(n_3212),
.Y(n_3414)
);

NAND2xp5_ASAP7_75t_L g3415 ( 
.A(n_3084),
.B(n_903),
.Y(n_3415)
);

NOR2xp33_ASAP7_75t_L g3416 ( 
.A(n_3222),
.B(n_816),
.Y(n_3416)
);

BUFx2_ASAP7_75t_L g3417 ( 
.A(n_3084),
.Y(n_3417)
);

A2O1A1Ixp33_ASAP7_75t_L g3418 ( 
.A1(n_3131),
.A2(n_2307),
.B(n_2308),
.C(n_2304),
.Y(n_3418)
);

AND2x2_ASAP7_75t_L g3419 ( 
.A(n_3113),
.B(n_1134),
.Y(n_3419)
);

BUFx2_ASAP7_75t_L g3420 ( 
.A(n_3113),
.Y(n_3420)
);

AOI21xp5_ASAP7_75t_L g3421 ( 
.A1(n_3162),
.A2(n_2229),
.B(n_2228),
.Y(n_3421)
);

NOR3xp33_ASAP7_75t_L g3422 ( 
.A(n_3138),
.B(n_1138),
.C(n_1135),
.Y(n_3422)
);

NOR2x1_ASAP7_75t_L g3423 ( 
.A(n_3021),
.B(n_2313),
.Y(n_3423)
);

AOI21xp5_ASAP7_75t_L g3424 ( 
.A1(n_3021),
.A2(n_2229),
.B(n_2228),
.Y(n_3424)
);

OAI22xp5_ASAP7_75t_L g3425 ( 
.A1(n_3105),
.A2(n_908),
.B1(n_909),
.B2(n_903),
.Y(n_3425)
);

NOR2xp33_ASAP7_75t_L g3426 ( 
.A(n_3077),
.B(n_817),
.Y(n_3426)
);

OAI22xp5_ASAP7_75t_L g3427 ( 
.A1(n_3105),
.A2(n_909),
.B1(n_916),
.B2(n_908),
.Y(n_3427)
);

NOR2xp33_ASAP7_75t_SL g3428 ( 
.A(n_3105),
.B(n_916),
.Y(n_3428)
);

NAND2xp5_ASAP7_75t_L g3429 ( 
.A(n_3057),
.B(n_919),
.Y(n_3429)
);

INVx2_ASAP7_75t_L g3430 ( 
.A(n_3022),
.Y(n_3430)
);

INVxp67_ASAP7_75t_SL g3431 ( 
.A(n_3258),
.Y(n_3431)
);

INVx1_ASAP7_75t_L g3432 ( 
.A(n_3396),
.Y(n_3432)
);

CKINVDCx14_ASAP7_75t_R g3433 ( 
.A(n_3344),
.Y(n_3433)
);

OA21x2_ASAP7_75t_L g3434 ( 
.A1(n_3339),
.A2(n_2240),
.B(n_2234),
.Y(n_3434)
);

BUFx6f_ASAP7_75t_L g3435 ( 
.A(n_3399),
.Y(n_3435)
);

AO31x2_ASAP7_75t_L g3436 ( 
.A1(n_3348),
.A2(n_2240),
.A3(n_2241),
.B(n_2234),
.Y(n_3436)
);

OAI21x1_ASAP7_75t_L g3437 ( 
.A1(n_3250),
.A2(n_2209),
.B(n_2207),
.Y(n_3437)
);

NAND3x1_ASAP7_75t_L g3438 ( 
.A(n_3232),
.B(n_1140),
.C(n_1139),
.Y(n_3438)
);

AND2x2_ASAP7_75t_L g3439 ( 
.A(n_3286),
.B(n_1147),
.Y(n_3439)
);

OAI21x1_ASAP7_75t_L g3440 ( 
.A1(n_3229),
.A2(n_3251),
.B(n_3306),
.Y(n_3440)
);

CKINVDCx5p33_ASAP7_75t_R g3441 ( 
.A(n_3334),
.Y(n_3441)
);

NAND2xp5_ASAP7_75t_SL g3442 ( 
.A(n_3227),
.B(n_2241),
.Y(n_3442)
);

OR2x2_ASAP7_75t_L g3443 ( 
.A(n_3285),
.B(n_1646),
.Y(n_3443)
);

OAI21x1_ASAP7_75t_L g3444 ( 
.A1(n_3282),
.A2(n_2209),
.B(n_2207),
.Y(n_3444)
);

INVx2_ASAP7_75t_L g3445 ( 
.A(n_3328),
.Y(n_3445)
);

INVx2_ASAP7_75t_L g3446 ( 
.A(n_3333),
.Y(n_3446)
);

AO31x2_ASAP7_75t_L g3447 ( 
.A1(n_3288),
.A2(n_2247),
.A3(n_2253),
.B(n_2244),
.Y(n_3447)
);

INVx1_ASAP7_75t_L g3448 ( 
.A(n_3237),
.Y(n_3448)
);

OAI21x1_ASAP7_75t_L g3449 ( 
.A1(n_3357),
.A2(n_2254),
.B(n_2219),
.Y(n_3449)
);

OAI21xp5_ASAP7_75t_L g3450 ( 
.A1(n_3325),
.A2(n_1153),
.B(n_1152),
.Y(n_3450)
);

AO22x2_ASAP7_75t_L g3451 ( 
.A1(n_3297),
.A2(n_2472),
.B1(n_1157),
.B2(n_1158),
.Y(n_3451)
);

OR2x2_ASAP7_75t_L g3452 ( 
.A(n_3248),
.B(n_1646),
.Y(n_3452)
);

AOI221xp5_ASAP7_75t_SL g3453 ( 
.A1(n_3425),
.A2(n_1162),
.B1(n_1163),
.B2(n_1161),
.C(n_1154),
.Y(n_3453)
);

NAND2xp33_ASAP7_75t_L g3454 ( 
.A(n_3314),
.B(n_919),
.Y(n_3454)
);

INVx5_ASAP7_75t_L g3455 ( 
.A(n_3293),
.Y(n_3455)
);

NAND2xp5_ASAP7_75t_L g3456 ( 
.A(n_3263),
.B(n_818),
.Y(n_3456)
);

OA21x2_ASAP7_75t_L g3457 ( 
.A1(n_3256),
.A2(n_2247),
.B(n_2244),
.Y(n_3457)
);

AND2x2_ASAP7_75t_L g3458 ( 
.A(n_3292),
.B(n_1434),
.Y(n_3458)
);

BUFx6f_ASAP7_75t_L g3459 ( 
.A(n_3399),
.Y(n_3459)
);

AOI21xp5_ASAP7_75t_L g3460 ( 
.A1(n_3230),
.A2(n_2253),
.B(n_2307),
.Y(n_3460)
);

INVx1_ASAP7_75t_L g3461 ( 
.A(n_3247),
.Y(n_3461)
);

OAI21x1_ASAP7_75t_L g3462 ( 
.A1(n_3359),
.A2(n_2254),
.B(n_2219),
.Y(n_3462)
);

INVx1_ASAP7_75t_L g3463 ( 
.A(n_3257),
.Y(n_3463)
);

NAND3xp33_ASAP7_75t_L g3464 ( 
.A(n_3428),
.B(n_934),
.C(n_921),
.Y(n_3464)
);

OAI21xp5_ASAP7_75t_L g3465 ( 
.A1(n_3325),
.A2(n_2308),
.B(n_2001),
.Y(n_3465)
);

OAI21x1_ASAP7_75t_SL g3466 ( 
.A1(n_3291),
.A2(n_3295),
.B(n_3323),
.Y(n_3466)
);

INVx4_ASAP7_75t_L g3467 ( 
.A(n_3293),
.Y(n_3467)
);

AO31x2_ASAP7_75t_L g3468 ( 
.A1(n_3243),
.A2(n_2312),
.A3(n_2317),
.B(n_2310),
.Y(n_3468)
);

OAI21x1_ASAP7_75t_L g3469 ( 
.A1(n_3320),
.A2(n_2254),
.B(n_2219),
.Y(n_3469)
);

OAI21x1_ASAP7_75t_L g3470 ( 
.A1(n_3287),
.A2(n_2334),
.B(n_2322),
.Y(n_3470)
);

BUFx2_ASAP7_75t_SL g3471 ( 
.A(n_3278),
.Y(n_3471)
);

AOI221xp5_ASAP7_75t_SL g3472 ( 
.A1(n_3427),
.A2(n_937),
.B1(n_939),
.B2(n_934),
.C(n_921),
.Y(n_3472)
);

OAI21xp5_ASAP7_75t_L g3473 ( 
.A1(n_3281),
.A2(n_2005),
.B(n_2000),
.Y(n_3473)
);

AOI21xp5_ASAP7_75t_L g3474 ( 
.A1(n_3400),
.A2(n_1854),
.B(n_1852),
.Y(n_3474)
);

OAI21xp5_ASAP7_75t_L g3475 ( 
.A1(n_3232),
.A2(n_3262),
.B(n_3244),
.Y(n_3475)
);

NOR2xp33_ASAP7_75t_L g3476 ( 
.A(n_3239),
.B(n_824),
.Y(n_3476)
);

OAI22xp5_ASAP7_75t_L g3477 ( 
.A1(n_3227),
.A2(n_939),
.B1(n_940),
.B2(n_937),
.Y(n_3477)
);

NAND2xp5_ASAP7_75t_L g3478 ( 
.A(n_3296),
.B(n_825),
.Y(n_3478)
);

INVx1_ASAP7_75t_L g3479 ( 
.A(n_3345),
.Y(n_3479)
);

OAI22xp5_ASAP7_75t_L g3480 ( 
.A1(n_3240),
.A2(n_943),
.B1(n_947),
.B2(n_940),
.Y(n_3480)
);

NAND3xp33_ASAP7_75t_L g3481 ( 
.A(n_3428),
.B(n_947),
.C(n_943),
.Y(n_3481)
);

AOI221x1_ASAP7_75t_L g3482 ( 
.A1(n_3390),
.A2(n_2013),
.B1(n_2010),
.B2(n_2006),
.C(n_1972),
.Y(n_3482)
);

AOI21x1_ASAP7_75t_L g3483 ( 
.A1(n_3249),
.A2(n_2312),
.B(n_2310),
.Y(n_3483)
);

INVx2_ASAP7_75t_L g3484 ( 
.A(n_3342),
.Y(n_3484)
);

INVx1_ASAP7_75t_SL g3485 ( 
.A(n_3234),
.Y(n_3485)
);

OAI21xp5_ASAP7_75t_L g3486 ( 
.A1(n_3284),
.A2(n_1861),
.B(n_1855),
.Y(n_3486)
);

AO21x1_ASAP7_75t_L g3487 ( 
.A1(n_3255),
.A2(n_2324),
.B(n_2317),
.Y(n_3487)
);

AO31x2_ASAP7_75t_L g3488 ( 
.A1(n_3241),
.A2(n_2326),
.A3(n_2328),
.B(n_2324),
.Y(n_3488)
);

AO21x1_ASAP7_75t_L g3489 ( 
.A1(n_3355),
.A2(n_2328),
.B(n_2326),
.Y(n_3489)
);

AOI21xp5_ASAP7_75t_L g3490 ( 
.A1(n_3380),
.A2(n_1869),
.B(n_1867),
.Y(n_3490)
);

OAI21x1_ASAP7_75t_L g3491 ( 
.A1(n_3375),
.A2(n_2334),
.B(n_2322),
.Y(n_3491)
);

OAI21xp5_ASAP7_75t_L g3492 ( 
.A1(n_3260),
.A2(n_1872),
.B(n_2330),
.Y(n_3492)
);

OAI21x1_ASAP7_75t_SL g3493 ( 
.A1(n_3261),
.A2(n_3338),
.B(n_3343),
.Y(n_3493)
);

NAND2xp5_ASAP7_75t_SL g3494 ( 
.A(n_3240),
.B(n_2472),
.Y(n_3494)
);

OAI21x1_ASAP7_75t_L g3495 ( 
.A1(n_3304),
.A2(n_2334),
.B(n_2322),
.Y(n_3495)
);

INVx3_ASAP7_75t_L g3496 ( 
.A(n_3360),
.Y(n_3496)
);

NAND2xp5_ASAP7_75t_L g3497 ( 
.A(n_3233),
.B(n_826),
.Y(n_3497)
);

OAI21x1_ASAP7_75t_L g3498 ( 
.A1(n_3388),
.A2(n_3313),
.B(n_3273),
.Y(n_3498)
);

INVx2_ASAP7_75t_L g3499 ( 
.A(n_3350),
.Y(n_3499)
);

AOI22x1_ASAP7_75t_L g3500 ( 
.A1(n_3335),
.A2(n_950),
.B1(n_948),
.B2(n_828),
.Y(n_3500)
);

AO31x2_ASAP7_75t_L g3501 ( 
.A1(n_3231),
.A2(n_2331),
.A3(n_2333),
.B(n_2330),
.Y(n_3501)
);

NOR2xp33_ASAP7_75t_L g3502 ( 
.A(n_3264),
.B(n_827),
.Y(n_3502)
);

BUFx2_ASAP7_75t_L g3503 ( 
.A(n_3298),
.Y(n_3503)
);

OAI21xp5_ASAP7_75t_L g3504 ( 
.A1(n_3301),
.A2(n_2333),
.B(n_2331),
.Y(n_3504)
);

OAI21x1_ASAP7_75t_L g3505 ( 
.A1(n_3347),
.A2(n_2374),
.B(n_2373),
.Y(n_3505)
);

OR2x6_ASAP7_75t_L g3506 ( 
.A(n_3307),
.B(n_3236),
.Y(n_3506)
);

AND2x2_ASAP7_75t_L g3507 ( 
.A(n_3283),
.B(n_1434),
.Y(n_3507)
);

NAND2xp5_ASAP7_75t_SL g3508 ( 
.A(n_3305),
.B(n_2472),
.Y(n_3508)
);

OAI21x1_ASAP7_75t_L g3509 ( 
.A1(n_3277),
.A2(n_2374),
.B(n_2373),
.Y(n_3509)
);

AND2x2_ASAP7_75t_L g3510 ( 
.A(n_3294),
.B(n_1447),
.Y(n_3510)
);

AO21x2_ASAP7_75t_L g3511 ( 
.A1(n_3371),
.A2(n_2340),
.B(n_2335),
.Y(n_3511)
);

AOI21x1_ASAP7_75t_L g3512 ( 
.A1(n_3289),
.A2(n_2340),
.B(n_2335),
.Y(n_3512)
);

NAND2xp5_ASAP7_75t_L g3513 ( 
.A(n_3238),
.B(n_832),
.Y(n_3513)
);

AND2x4_ASAP7_75t_L g3514 ( 
.A(n_3274),
.B(n_2346),
.Y(n_3514)
);

CKINVDCx14_ASAP7_75t_R g3515 ( 
.A(n_3351),
.Y(n_3515)
);

AND2x4_ASAP7_75t_L g3516 ( 
.A(n_3274),
.B(n_2346),
.Y(n_3516)
);

NAND2xp5_ASAP7_75t_L g3517 ( 
.A(n_3253),
.B(n_834),
.Y(n_3517)
);

AO31x2_ASAP7_75t_L g3518 ( 
.A1(n_3252),
.A2(n_2349),
.A3(n_2352),
.B(n_2348),
.Y(n_3518)
);

INVx4_ASAP7_75t_L g3519 ( 
.A(n_3293),
.Y(n_3519)
);

INVx1_ASAP7_75t_L g3520 ( 
.A(n_3352),
.Y(n_3520)
);

A2O1A1Ixp33_ASAP7_75t_L g3521 ( 
.A1(n_3416),
.A2(n_950),
.B(n_948),
.C(n_845),
.Y(n_3521)
);

OAI21x1_ASAP7_75t_L g3522 ( 
.A1(n_3310),
.A2(n_2374),
.B(n_2349),
.Y(n_3522)
);

INVx8_ASAP7_75t_L g3523 ( 
.A(n_3399),
.Y(n_3523)
);

BUFx4_ASAP7_75t_SL g3524 ( 
.A(n_3322),
.Y(n_3524)
);

INVx1_ASAP7_75t_L g3525 ( 
.A(n_3353),
.Y(n_3525)
);

INVx2_ASAP7_75t_L g3526 ( 
.A(n_3365),
.Y(n_3526)
);

AOI21xp5_ASAP7_75t_L g3527 ( 
.A1(n_3379),
.A2(n_2352),
.B(n_2348),
.Y(n_3527)
);

OA22x2_ASAP7_75t_L g3528 ( 
.A1(n_3309),
.A2(n_846),
.B1(n_847),
.B2(n_840),
.Y(n_3528)
);

INVxp67_ASAP7_75t_SL g3529 ( 
.A(n_3303),
.Y(n_3529)
);

OAI21x1_ASAP7_75t_L g3530 ( 
.A1(n_3403),
.A2(n_2364),
.B(n_2363),
.Y(n_3530)
);

BUFx3_ASAP7_75t_L g3531 ( 
.A(n_3363),
.Y(n_3531)
);

OAI21x1_ASAP7_75t_SL g3532 ( 
.A1(n_3343),
.A2(n_2364),
.B(n_2363),
.Y(n_3532)
);

NAND2xp5_ASAP7_75t_L g3533 ( 
.A(n_3226),
.B(n_848),
.Y(n_3533)
);

INVx2_ASAP7_75t_L g3534 ( 
.A(n_3430),
.Y(n_3534)
);

OAI21x1_ASAP7_75t_L g3535 ( 
.A1(n_3384),
.A2(n_2369),
.B(n_2366),
.Y(n_3535)
);

OAI21x1_ASAP7_75t_L g3536 ( 
.A1(n_3404),
.A2(n_2369),
.B(n_2366),
.Y(n_3536)
);

OAI21xp5_ASAP7_75t_L g3537 ( 
.A1(n_3246),
.A2(n_2372),
.B(n_2371),
.Y(n_3537)
);

O2A1O1Ixp5_ASAP7_75t_L g3538 ( 
.A1(n_3265),
.A2(n_2372),
.B(n_2375),
.C(n_2371),
.Y(n_3538)
);

AOI21xp33_ASAP7_75t_L g3539 ( 
.A1(n_3299),
.A2(n_1970),
.B(n_1968),
.Y(n_3539)
);

AND2x2_ASAP7_75t_L g3540 ( 
.A(n_3234),
.B(n_1447),
.Y(n_3540)
);

AOI21xp5_ASAP7_75t_L g3541 ( 
.A1(n_3269),
.A2(n_2375),
.B(n_1981),
.Y(n_3541)
);

AOI221xp5_ASAP7_75t_L g3542 ( 
.A1(n_3385),
.A2(n_860),
.B1(n_863),
.B2(n_853),
.C(n_849),
.Y(n_3542)
);

NAND2xp5_ASAP7_75t_L g3543 ( 
.A(n_3308),
.B(n_873),
.Y(n_3543)
);

BUFx2_ASAP7_75t_SL g3544 ( 
.A(n_3236),
.Y(n_3544)
);

AOI21xp5_ASAP7_75t_L g3545 ( 
.A1(n_3275),
.A2(n_3300),
.B(n_3346),
.Y(n_3545)
);

NAND2xp5_ASAP7_75t_SL g3546 ( 
.A(n_3312),
.B(n_1599),
.Y(n_3546)
);

NAND2xp5_ASAP7_75t_L g3547 ( 
.A(n_3270),
.B(n_3392),
.Y(n_3547)
);

INVx3_ASAP7_75t_L g3548 ( 
.A(n_3360),
.Y(n_3548)
);

OAI21xp5_ASAP7_75t_L g3549 ( 
.A1(n_3268),
.A2(n_959),
.B(n_874),
.Y(n_3549)
);

OAI21x1_ASAP7_75t_L g3550 ( 
.A1(n_3406),
.A2(n_1833),
.B(n_1828),
.Y(n_3550)
);

OAI22x1_ASAP7_75t_L g3551 ( 
.A1(n_3354),
.A2(n_6),
.B1(n_2),
.B2(n_4),
.Y(n_3551)
);

BUFx6f_ASAP7_75t_L g3552 ( 
.A(n_3364),
.Y(n_3552)
);

CKINVDCx5p33_ASAP7_75t_R g3553 ( 
.A(n_3279),
.Y(n_3553)
);

OAI21x1_ASAP7_75t_L g3554 ( 
.A1(n_3394),
.A2(n_1833),
.B(n_1828),
.Y(n_3554)
);

OAI21xp5_ASAP7_75t_L g3555 ( 
.A1(n_3426),
.A2(n_1662),
.B(n_1828),
.Y(n_3555)
);

AOI21xp5_ASAP7_75t_L g3556 ( 
.A1(n_3267),
.A2(n_1965),
.B(n_1941),
.Y(n_3556)
);

OR2x2_ASAP7_75t_L g3557 ( 
.A(n_3245),
.B(n_3254),
.Y(n_3557)
);

OAI21xp5_ASAP7_75t_L g3558 ( 
.A1(n_3372),
.A2(n_1835),
.B(n_1833),
.Y(n_3558)
);

AOI21xp5_ASAP7_75t_L g3559 ( 
.A1(n_3356),
.A2(n_1965),
.B(n_1941),
.Y(n_3559)
);

OR2x2_ASAP7_75t_L g3560 ( 
.A(n_3235),
.B(n_1599),
.Y(n_3560)
);

NAND2xp5_ASAP7_75t_L g3561 ( 
.A(n_3370),
.B(n_1599),
.Y(n_3561)
);

NAND2xp5_ASAP7_75t_L g3562 ( 
.A(n_3373),
.B(n_1599),
.Y(n_3562)
);

BUFx3_ASAP7_75t_L g3563 ( 
.A(n_3398),
.Y(n_3563)
);

AOI21xp5_ASAP7_75t_L g3564 ( 
.A1(n_3356),
.A2(n_1965),
.B(n_1941),
.Y(n_3564)
);

NAND2xp5_ASAP7_75t_SL g3565 ( 
.A(n_3276),
.B(n_1600),
.Y(n_3565)
);

OAI21x1_ASAP7_75t_L g3566 ( 
.A1(n_3421),
.A2(n_1838),
.B(n_1835),
.Y(n_3566)
);

AOI21xp5_ASAP7_75t_L g3567 ( 
.A1(n_3349),
.A2(n_1974),
.B(n_1965),
.Y(n_3567)
);

OAI22xp5_ASAP7_75t_L g3568 ( 
.A1(n_3242),
.A2(n_1838),
.B1(n_1841),
.B2(n_1835),
.Y(n_3568)
);

INVx2_ASAP7_75t_L g3569 ( 
.A(n_3259),
.Y(n_3569)
);

OAI21xp5_ASAP7_75t_L g3570 ( 
.A1(n_3368),
.A2(n_1841),
.B(n_1838),
.Y(n_3570)
);

INVx1_ASAP7_75t_SL g3571 ( 
.A(n_3271),
.Y(n_3571)
);

NAND2xp5_ASAP7_75t_L g3572 ( 
.A(n_3429),
.B(n_1600),
.Y(n_3572)
);

BUFx2_ASAP7_75t_L g3573 ( 
.A(n_3367),
.Y(n_3573)
);

OA21x2_ASAP7_75t_L g3574 ( 
.A1(n_3418),
.A2(n_1607),
.B(n_1600),
.Y(n_3574)
);

NAND2xp5_ASAP7_75t_L g3575 ( 
.A(n_3266),
.B(n_3272),
.Y(n_3575)
);

NAND2xp5_ASAP7_75t_L g3576 ( 
.A(n_3302),
.B(n_1600),
.Y(n_3576)
);

NAND2xp5_ASAP7_75t_L g3577 ( 
.A(n_3311),
.B(n_1607),
.Y(n_3577)
);

INVx5_ASAP7_75t_L g3578 ( 
.A(n_3364),
.Y(n_3578)
);

OAI21xp5_ASAP7_75t_L g3579 ( 
.A1(n_3381),
.A2(n_1876),
.B(n_1841),
.Y(n_3579)
);

NAND2xp5_ASAP7_75t_L g3580 ( 
.A(n_3327),
.B(n_3331),
.Y(n_3580)
);

OA22x2_ASAP7_75t_L g3581 ( 
.A1(n_3280),
.A2(n_8),
.B1(n_4),
.B2(n_6),
.Y(n_3581)
);

BUFx3_ASAP7_75t_L g3582 ( 
.A(n_3366),
.Y(n_3582)
);

NOR2x1_ASAP7_75t_L g3583 ( 
.A(n_3228),
.B(n_1542),
.Y(n_3583)
);

AOI221xp5_ASAP7_75t_SL g3584 ( 
.A1(n_3395),
.A2(n_1623),
.B1(n_1632),
.B2(n_1611),
.C(n_1607),
.Y(n_3584)
);

OAI22x1_ASAP7_75t_L g3585 ( 
.A1(n_3290),
.A2(n_12),
.B1(n_8),
.B2(n_10),
.Y(n_3585)
);

NAND2xp5_ASAP7_75t_L g3586 ( 
.A(n_3316),
.B(n_1607),
.Y(n_3586)
);

AO21x2_ASAP7_75t_L g3587 ( 
.A1(n_3422),
.A2(n_1975),
.B(n_1974),
.Y(n_3587)
);

BUFx4f_ASAP7_75t_L g3588 ( 
.A(n_3374),
.Y(n_3588)
);

AOI21xp5_ASAP7_75t_SL g3589 ( 
.A1(n_3317),
.A2(n_1975),
.B(n_1974),
.Y(n_3589)
);

AOI21xp5_ASAP7_75t_L g3590 ( 
.A1(n_3383),
.A2(n_1975),
.B(n_1974),
.Y(n_3590)
);

OAI21x1_ASAP7_75t_L g3591 ( 
.A1(n_3424),
.A2(n_1909),
.B(n_1876),
.Y(n_3591)
);

NOR2x1_ASAP7_75t_R g3592 ( 
.A(n_3367),
.B(n_1611),
.Y(n_3592)
);

AOI21xp5_ASAP7_75t_L g3593 ( 
.A1(n_3340),
.A2(n_1978),
.B(n_1975),
.Y(n_3593)
);

INVx1_ASAP7_75t_L g3594 ( 
.A(n_3336),
.Y(n_3594)
);

OR2x2_ASAP7_75t_L g3595 ( 
.A(n_3319),
.B(n_1611),
.Y(n_3595)
);

INVx2_ASAP7_75t_L g3596 ( 
.A(n_3324),
.Y(n_3596)
);

INVx1_ASAP7_75t_L g3597 ( 
.A(n_3337),
.Y(n_3597)
);

INVx1_ASAP7_75t_L g3598 ( 
.A(n_3411),
.Y(n_3598)
);

NAND2xp5_ASAP7_75t_SL g3599 ( 
.A(n_3330),
.B(n_1611),
.Y(n_3599)
);

OAI21x1_ASAP7_75t_L g3600 ( 
.A1(n_3423),
.A2(n_1909),
.B(n_1876),
.Y(n_3600)
);

INVx1_ASAP7_75t_L g3601 ( 
.A(n_3411),
.Y(n_3601)
);

BUFx6f_ASAP7_75t_SL g3602 ( 
.A(n_3397),
.Y(n_3602)
);

AOI21xp5_ASAP7_75t_L g3603 ( 
.A1(n_3410),
.A2(n_1982),
.B(n_1978),
.Y(n_3603)
);

BUFx2_ASAP7_75t_L g3604 ( 
.A(n_3374),
.Y(n_3604)
);

NAND2xp5_ASAP7_75t_L g3605 ( 
.A(n_3382),
.B(n_1623),
.Y(n_3605)
);

NAND2xp5_ASAP7_75t_L g3606 ( 
.A(n_3387),
.B(n_1623),
.Y(n_3606)
);

OAI21x1_ASAP7_75t_L g3607 ( 
.A1(n_3377),
.A2(n_1909),
.B(n_1978),
.Y(n_3607)
);

OAI22xp5_ASAP7_75t_L g3608 ( 
.A1(n_3326),
.A2(n_1982),
.B1(n_1987),
.B2(n_1978),
.Y(n_3608)
);

OAI21x1_ASAP7_75t_L g3609 ( 
.A1(n_3377),
.A2(n_1987),
.B(n_1982),
.Y(n_3609)
);

NAND2xp5_ASAP7_75t_L g3610 ( 
.A(n_3389),
.B(n_1623),
.Y(n_3610)
);

AOI21xp5_ASAP7_75t_L g3611 ( 
.A1(n_3376),
.A2(n_3321),
.B(n_3315),
.Y(n_3611)
);

OAI21x1_ASAP7_75t_L g3612 ( 
.A1(n_3386),
.A2(n_1987),
.B(n_1982),
.Y(n_3612)
);

BUFx2_ASAP7_75t_L g3613 ( 
.A(n_3417),
.Y(n_3613)
);

AOI21xp5_ASAP7_75t_L g3614 ( 
.A1(n_3414),
.A2(n_2002),
.B(n_1987),
.Y(n_3614)
);

OAI21xp5_ASAP7_75t_L g3615 ( 
.A1(n_3391),
.A2(n_3329),
.B(n_3369),
.Y(n_3615)
);

OAI21x1_ASAP7_75t_L g3616 ( 
.A1(n_3386),
.A2(n_2008),
.B(n_2002),
.Y(n_3616)
);

INVx1_ASAP7_75t_L g3617 ( 
.A(n_3402),
.Y(n_3617)
);

NAND2xp5_ASAP7_75t_L g3618 ( 
.A(n_3419),
.B(n_1632),
.Y(n_3618)
);

BUFx2_ASAP7_75t_L g3619 ( 
.A(n_3420),
.Y(n_3619)
);

AOI21xp5_ASAP7_75t_L g3620 ( 
.A1(n_3414),
.A2(n_3318),
.B(n_3407),
.Y(n_3620)
);

OAI21x1_ASAP7_75t_L g3621 ( 
.A1(n_3341),
.A2(n_2008),
.B(n_2002),
.Y(n_3621)
);

AOI21xp33_ASAP7_75t_L g3622 ( 
.A1(n_3361),
.A2(n_1632),
.B(n_2002),
.Y(n_3622)
);

OAI22xp5_ASAP7_75t_L g3623 ( 
.A1(n_3415),
.A2(n_2008),
.B1(n_1663),
.B2(n_1680),
.Y(n_3623)
);

CKINVDCx6p67_ASAP7_75t_R g3624 ( 
.A(n_3362),
.Y(n_3624)
);

OAI21x1_ASAP7_75t_L g3625 ( 
.A1(n_3412),
.A2(n_3401),
.B(n_3358),
.Y(n_3625)
);

AOI21xp5_ASAP7_75t_L g3626 ( 
.A1(n_3414),
.A2(n_2008),
.B(n_1672),
.Y(n_3626)
);

OA21x2_ASAP7_75t_L g3627 ( 
.A1(n_3408),
.A2(n_1632),
.B(n_1620),
.Y(n_3627)
);

OAI21xp33_ASAP7_75t_L g3628 ( 
.A1(n_3332),
.A2(n_1546),
.B(n_1543),
.Y(n_3628)
);

AND2x2_ASAP7_75t_L g3629 ( 
.A(n_3405),
.B(n_3362),
.Y(n_3629)
);

AND2x4_ASAP7_75t_L g3630 ( 
.A(n_3318),
.B(n_303),
.Y(n_3630)
);

AOI21x1_ASAP7_75t_L g3631 ( 
.A1(n_3393),
.A2(n_1399),
.B(n_1354),
.Y(n_3631)
);

NOR2x1_ASAP7_75t_SL g3632 ( 
.A(n_3413),
.B(n_3409),
.Y(n_3632)
);

NAND2xp5_ASAP7_75t_L g3633 ( 
.A(n_3401),
.B(n_12),
.Y(n_3633)
);

NAND2xp5_ASAP7_75t_L g3634 ( 
.A(n_3413),
.B(n_3378),
.Y(n_3634)
);

BUFx6f_ASAP7_75t_L g3635 ( 
.A(n_3397),
.Y(n_3635)
);

AOI21xp5_ASAP7_75t_L g3636 ( 
.A1(n_3229),
.A2(n_1672),
.B(n_1663),
.Y(n_3636)
);

AOI21xp33_ASAP7_75t_L g3637 ( 
.A1(n_3297),
.A2(n_14),
.B(n_15),
.Y(n_3637)
);

AOI21x1_ASAP7_75t_L g3638 ( 
.A1(n_3320),
.A2(n_1399),
.B(n_1354),
.Y(n_3638)
);

INVx1_ASAP7_75t_L g3639 ( 
.A(n_3396),
.Y(n_3639)
);

AOI22xp5_ASAP7_75t_L g3640 ( 
.A1(n_3428),
.A2(n_1560),
.B1(n_1399),
.B2(n_1354),
.Y(n_3640)
);

O2A1O1Ixp5_ASAP7_75t_L g3641 ( 
.A1(n_3288),
.A2(n_1768),
.B(n_1757),
.C(n_17),
.Y(n_3641)
);

OAI21xp5_ASAP7_75t_L g3642 ( 
.A1(n_3325),
.A2(n_1399),
.B(n_1354),
.Y(n_3642)
);

AO31x2_ASAP7_75t_L g3643 ( 
.A1(n_3348),
.A2(n_1757),
.A3(n_1768),
.B(n_1399),
.Y(n_3643)
);

INVx1_ASAP7_75t_SL g3644 ( 
.A(n_3485),
.Y(n_3644)
);

NAND2xp5_ASAP7_75t_L g3645 ( 
.A(n_3529),
.B(n_15),
.Y(n_3645)
);

NAND3xp33_ASAP7_75t_L g3646 ( 
.A(n_3549),
.B(n_1546),
.C(n_1543),
.Y(n_3646)
);

BUFx3_ASAP7_75t_L g3647 ( 
.A(n_3503),
.Y(n_3647)
);

INVx3_ASAP7_75t_L g3648 ( 
.A(n_3445),
.Y(n_3648)
);

INVx1_ASAP7_75t_L g3649 ( 
.A(n_3432),
.Y(n_3649)
);

BUFx2_ASAP7_75t_L g3650 ( 
.A(n_3613),
.Y(n_3650)
);

OR2x2_ASAP7_75t_L g3651 ( 
.A(n_3431),
.B(n_16),
.Y(n_3651)
);

HB1xp67_ASAP7_75t_L g3652 ( 
.A(n_3619),
.Y(n_3652)
);

INVx1_ASAP7_75t_L g3653 ( 
.A(n_3432),
.Y(n_3653)
);

INVx1_ASAP7_75t_L g3654 ( 
.A(n_3639),
.Y(n_3654)
);

AOI21xp5_ASAP7_75t_L g3655 ( 
.A1(n_3545),
.A2(n_3493),
.B(n_3559),
.Y(n_3655)
);

INVx1_ASAP7_75t_SL g3656 ( 
.A(n_3557),
.Y(n_3656)
);

OR2x2_ASAP7_75t_L g3657 ( 
.A(n_3463),
.B(n_18),
.Y(n_3657)
);

AOI22xp33_ASAP7_75t_SL g3658 ( 
.A1(n_3475),
.A2(n_22),
.B1(n_20),
.B2(n_21),
.Y(n_3658)
);

AND2x2_ASAP7_75t_L g3659 ( 
.A(n_3629),
.B(n_20),
.Y(n_3659)
);

BUFx6f_ASAP7_75t_L g3660 ( 
.A(n_3435),
.Y(n_3660)
);

AOI22xp33_ASAP7_75t_L g3661 ( 
.A1(n_3637),
.A2(n_1546),
.B1(n_1543),
.B2(n_1432),
.Y(n_3661)
);

CKINVDCx5p33_ASAP7_75t_R g3662 ( 
.A(n_3441),
.Y(n_3662)
);

NAND2xp5_ASAP7_75t_L g3663 ( 
.A(n_3547),
.B(n_21),
.Y(n_3663)
);

AND2x4_ASAP7_75t_L g3664 ( 
.A(n_3463),
.B(n_3479),
.Y(n_3664)
);

NOR2xp67_ASAP7_75t_L g3665 ( 
.A(n_3443),
.B(n_22),
.Y(n_3665)
);

INVx2_ASAP7_75t_L g3666 ( 
.A(n_3446),
.Y(n_3666)
);

INVx1_ASAP7_75t_L g3667 ( 
.A(n_3479),
.Y(n_3667)
);

OAI21xp33_ASAP7_75t_L g3668 ( 
.A1(n_3476),
.A2(n_1546),
.B(n_1543),
.Y(n_3668)
);

AOI21xp5_ASAP7_75t_L g3669 ( 
.A1(n_3564),
.A2(n_1672),
.B(n_1663),
.Y(n_3669)
);

BUFx3_ASAP7_75t_L g3670 ( 
.A(n_3531),
.Y(n_3670)
);

OAI22xp5_ASAP7_75t_L g3671 ( 
.A1(n_3464),
.A2(n_1443),
.B1(n_1452),
.B2(n_1432),
.Y(n_3671)
);

INVx1_ASAP7_75t_L g3672 ( 
.A(n_3520),
.Y(n_3672)
);

NAND2x1p5_ASAP7_75t_L g3673 ( 
.A(n_3455),
.B(n_1432),
.Y(n_3673)
);

AND2x4_ASAP7_75t_L g3674 ( 
.A(n_3520),
.B(n_3525),
.Y(n_3674)
);

CKINVDCx20_ASAP7_75t_R g3675 ( 
.A(n_3553),
.Y(n_3675)
);

CKINVDCx5p33_ASAP7_75t_R g3676 ( 
.A(n_3524),
.Y(n_3676)
);

AOI21xp5_ASAP7_75t_L g3677 ( 
.A1(n_3589),
.A2(n_1680),
.B(n_1672),
.Y(n_3677)
);

AND2x2_ASAP7_75t_L g3678 ( 
.A(n_3448),
.B(n_23),
.Y(n_3678)
);

INVx1_ASAP7_75t_L g3679 ( 
.A(n_3639),
.Y(n_3679)
);

AOI21xp5_ASAP7_75t_L g3680 ( 
.A1(n_3556),
.A2(n_3486),
.B(n_3466),
.Y(n_3680)
);

AND2x4_ASAP7_75t_L g3681 ( 
.A(n_3525),
.B(n_305),
.Y(n_3681)
);

AND2x2_ASAP7_75t_L g3682 ( 
.A(n_3461),
.B(n_24),
.Y(n_3682)
);

NAND2xp5_ASAP7_75t_L g3683 ( 
.A(n_3594),
.B(n_24),
.Y(n_3683)
);

AOI21xp5_ASAP7_75t_L g3684 ( 
.A1(n_3636),
.A2(n_1682),
.B(n_1680),
.Y(n_3684)
);

AOI21xp5_ASAP7_75t_SL g3685 ( 
.A1(n_3615),
.A2(n_1443),
.B(n_1432),
.Y(n_3685)
);

INVx2_ASAP7_75t_L g3686 ( 
.A(n_3484),
.Y(n_3686)
);

O2A1O1Ixp5_ASAP7_75t_L g3687 ( 
.A1(n_3565),
.A2(n_28),
.B(n_25),
.C(n_26),
.Y(n_3687)
);

AND2x2_ASAP7_75t_L g3688 ( 
.A(n_3510),
.B(n_25),
.Y(n_3688)
);

NOR2xp33_ASAP7_75t_L g3689 ( 
.A(n_3502),
.B(n_26),
.Y(n_3689)
);

AND2x2_ASAP7_75t_L g3690 ( 
.A(n_3458),
.B(n_29),
.Y(n_3690)
);

BUFx2_ASAP7_75t_L g3691 ( 
.A(n_3598),
.Y(n_3691)
);

INVx3_ASAP7_75t_L g3692 ( 
.A(n_3499),
.Y(n_3692)
);

INVx2_ASAP7_75t_L g3693 ( 
.A(n_3526),
.Y(n_3693)
);

AOI21xp5_ASAP7_75t_L g3694 ( 
.A1(n_3641),
.A2(n_1682),
.B(n_1680),
.Y(n_3694)
);

NAND2xp5_ASAP7_75t_L g3695 ( 
.A(n_3594),
.B(n_30),
.Y(n_3695)
);

NOR2xp33_ASAP7_75t_SL g3696 ( 
.A(n_3588),
.B(n_1479),
.Y(n_3696)
);

NAND2xp5_ASAP7_75t_L g3697 ( 
.A(n_3596),
.B(n_30),
.Y(n_3697)
);

BUFx6f_ASAP7_75t_L g3698 ( 
.A(n_3435),
.Y(n_3698)
);

BUFx2_ASAP7_75t_L g3699 ( 
.A(n_3598),
.Y(n_3699)
);

CKINVDCx5p33_ASAP7_75t_R g3700 ( 
.A(n_3515),
.Y(n_3700)
);

AND2x2_ASAP7_75t_L g3701 ( 
.A(n_3571),
.B(n_32),
.Y(n_3701)
);

AOI21xp5_ASAP7_75t_L g3702 ( 
.A1(n_3490),
.A2(n_1683),
.B(n_1682),
.Y(n_3702)
);

NAND2x1p5_ASAP7_75t_L g3703 ( 
.A(n_3455),
.B(n_1443),
.Y(n_3703)
);

NAND2xp5_ASAP7_75t_L g3704 ( 
.A(n_3580),
.B(n_32),
.Y(n_3704)
);

NAND2x1_ASAP7_75t_L g3705 ( 
.A(n_3467),
.B(n_1443),
.Y(n_3705)
);

BUFx6f_ASAP7_75t_L g3706 ( 
.A(n_3435),
.Y(n_3706)
);

BUFx2_ASAP7_75t_L g3707 ( 
.A(n_3601),
.Y(n_3707)
);

INVx1_ASAP7_75t_L g3708 ( 
.A(n_3597),
.Y(n_3708)
);

INVx2_ASAP7_75t_SL g3709 ( 
.A(n_3523),
.Y(n_3709)
);

NAND2xp5_ASAP7_75t_L g3710 ( 
.A(n_3534),
.B(n_3569),
.Y(n_3710)
);

OA21x2_ASAP7_75t_L g3711 ( 
.A1(n_3584),
.A2(n_33),
.B(n_34),
.Y(n_3711)
);

AOI21xp5_ASAP7_75t_L g3712 ( 
.A1(n_3599),
.A2(n_1683),
.B(n_1682),
.Y(n_3712)
);

INVx1_ASAP7_75t_L g3713 ( 
.A(n_3597),
.Y(n_3713)
);

AO21x1_ASAP7_75t_L g3714 ( 
.A1(n_3480),
.A2(n_34),
.B(n_35),
.Y(n_3714)
);

INVx3_ASAP7_75t_L g3715 ( 
.A(n_3459),
.Y(n_3715)
);

AOI21xp5_ASAP7_75t_L g3716 ( 
.A1(n_3474),
.A2(n_3504),
.B(n_3498),
.Y(n_3716)
);

AOI22xp5_ASAP7_75t_L g3717 ( 
.A1(n_3438),
.A2(n_1452),
.B1(n_1464),
.B2(n_1460),
.Y(n_3717)
);

INVx1_ASAP7_75t_L g3718 ( 
.A(n_3617),
.Y(n_3718)
);

AOI21xp5_ASAP7_75t_L g3719 ( 
.A1(n_3555),
.A2(n_1691),
.B(n_1683),
.Y(n_3719)
);

NAND2x1p5_ASAP7_75t_L g3720 ( 
.A(n_3455),
.B(n_1452),
.Y(n_3720)
);

INVx2_ASAP7_75t_L g3721 ( 
.A(n_3617),
.Y(n_3721)
);

OAI21xp33_ASAP7_75t_L g3722 ( 
.A1(n_3477),
.A2(n_1460),
.B(n_1452),
.Y(n_3722)
);

NAND2xp5_ASAP7_75t_L g3723 ( 
.A(n_3439),
.B(n_36),
.Y(n_3723)
);

INVx2_ASAP7_75t_L g3724 ( 
.A(n_3575),
.Y(n_3724)
);

OR2x2_ASAP7_75t_L g3725 ( 
.A(n_3452),
.B(n_37),
.Y(n_3725)
);

BUFx3_ASAP7_75t_L g3726 ( 
.A(n_3563),
.Y(n_3726)
);

INVx1_ASAP7_75t_L g3727 ( 
.A(n_3488),
.Y(n_3727)
);

HB1xp67_ASAP7_75t_L g3728 ( 
.A(n_3604),
.Y(n_3728)
);

OA21x2_ASAP7_75t_L g3729 ( 
.A1(n_3440),
.A2(n_38),
.B(n_41),
.Y(n_3729)
);

AOI21xp5_ASAP7_75t_L g3730 ( 
.A1(n_3590),
.A2(n_1691),
.B(n_1683),
.Y(n_3730)
);

NOR4xp25_ASAP7_75t_L g3731 ( 
.A(n_3481),
.B(n_45),
.C(n_42),
.D(n_43),
.Y(n_3731)
);

AOI21xp5_ASAP7_75t_L g3732 ( 
.A1(n_3588),
.A2(n_1698),
.B(n_1691),
.Y(n_3732)
);

NAND2xp5_ASAP7_75t_L g3733 ( 
.A(n_3540),
.B(n_45),
.Y(n_3733)
);

NAND2xp5_ASAP7_75t_L g3734 ( 
.A(n_3456),
.B(n_46),
.Y(n_3734)
);

BUFx2_ASAP7_75t_L g3735 ( 
.A(n_3601),
.Y(n_3735)
);

NAND2xp5_ASAP7_75t_L g3736 ( 
.A(n_3507),
.B(n_47),
.Y(n_3736)
);

INVx3_ASAP7_75t_L g3737 ( 
.A(n_3459),
.Y(n_3737)
);

INVx2_ASAP7_75t_L g3738 ( 
.A(n_3496),
.Y(n_3738)
);

INVx2_ASAP7_75t_L g3739 ( 
.A(n_3496),
.Y(n_3739)
);

NAND2xp5_ASAP7_75t_L g3740 ( 
.A(n_3478),
.B(n_3533),
.Y(n_3740)
);

INVx1_ASAP7_75t_SL g3741 ( 
.A(n_3471),
.Y(n_3741)
);

BUFx2_ASAP7_75t_L g3742 ( 
.A(n_3573),
.Y(n_3742)
);

INVx1_ASAP7_75t_L g3743 ( 
.A(n_3488),
.Y(n_3743)
);

INVx1_ASAP7_75t_L g3744 ( 
.A(n_3488),
.Y(n_3744)
);

AOI21xp5_ASAP7_75t_L g3745 ( 
.A1(n_3494),
.A2(n_1698),
.B(n_1691),
.Y(n_3745)
);

INVx5_ASAP7_75t_SL g3746 ( 
.A(n_3506),
.Y(n_3746)
);

CKINVDCx5p33_ASAP7_75t_R g3747 ( 
.A(n_3433),
.Y(n_3747)
);

AOI21xp5_ASAP7_75t_L g3748 ( 
.A1(n_3442),
.A2(n_1699),
.B(n_1698),
.Y(n_3748)
);

NAND2xp5_ASAP7_75t_SL g3749 ( 
.A(n_3634),
.B(n_1460),
.Y(n_3749)
);

INVx2_ASAP7_75t_L g3750 ( 
.A(n_3548),
.Y(n_3750)
);

NAND2x1_ASAP7_75t_L g3751 ( 
.A(n_3467),
.B(n_1460),
.Y(n_3751)
);

NOR2xp33_ASAP7_75t_L g3752 ( 
.A(n_3513),
.B(n_3517),
.Y(n_3752)
);

INVx2_ASAP7_75t_L g3753 ( 
.A(n_3548),
.Y(n_3753)
);

NAND2xp5_ASAP7_75t_SL g3754 ( 
.A(n_3583),
.B(n_1464),
.Y(n_3754)
);

BUFx2_ASAP7_75t_L g3755 ( 
.A(n_3624),
.Y(n_3755)
);

INVx3_ASAP7_75t_L g3756 ( 
.A(n_3459),
.Y(n_3756)
);

NAND2xp5_ASAP7_75t_L g3757 ( 
.A(n_3632),
.B(n_47),
.Y(n_3757)
);

OAI21x1_ASAP7_75t_L g3758 ( 
.A1(n_3512),
.A2(n_309),
.B(n_307),
.Y(n_3758)
);

BUFx3_ASAP7_75t_L g3759 ( 
.A(n_3582),
.Y(n_3759)
);

AND2x2_ASAP7_75t_L g3760 ( 
.A(n_3632),
.B(n_49),
.Y(n_3760)
);

CKINVDCx20_ASAP7_75t_R g3761 ( 
.A(n_3552),
.Y(n_3761)
);

INVx2_ASAP7_75t_SL g3762 ( 
.A(n_3523),
.Y(n_3762)
);

AOI22xp5_ASAP7_75t_L g3763 ( 
.A1(n_3454),
.A2(n_1464),
.B1(n_1560),
.B2(n_1620),
.Y(n_3763)
);

NOR2xp33_ASAP7_75t_L g3764 ( 
.A(n_3528),
.B(n_49),
.Y(n_3764)
);

AOI21xp5_ASAP7_75t_L g3765 ( 
.A1(n_3611),
.A2(n_1699),
.B(n_1698),
.Y(n_3765)
);

BUFx8_ASAP7_75t_SL g3766 ( 
.A(n_3602),
.Y(n_3766)
);

OAI22xp5_ASAP7_75t_L g3767 ( 
.A1(n_3521),
.A2(n_1464),
.B1(n_1703),
.B2(n_1699),
.Y(n_3767)
);

NAND2xp5_ASAP7_75t_L g3768 ( 
.A(n_3546),
.B(n_3543),
.Y(n_3768)
);

CKINVDCx20_ASAP7_75t_R g3769 ( 
.A(n_3552),
.Y(n_3769)
);

INVx1_ASAP7_75t_L g3770 ( 
.A(n_3501),
.Y(n_3770)
);

AND2x4_ASAP7_75t_L g3771 ( 
.A(n_3506),
.B(n_310),
.Y(n_3771)
);

INVx1_ASAP7_75t_L g3772 ( 
.A(n_3501),
.Y(n_3772)
);

OR2x6_ASAP7_75t_SL g3773 ( 
.A(n_3633),
.B(n_50),
.Y(n_3773)
);

OAI22xp5_ASAP7_75t_L g3774 ( 
.A1(n_3508),
.A2(n_1703),
.B1(n_1709),
.B2(n_1699),
.Y(n_3774)
);

NAND2xp5_ASAP7_75t_L g3775 ( 
.A(n_3497),
.B(n_51),
.Y(n_3775)
);

BUFx3_ASAP7_75t_L g3776 ( 
.A(n_3552),
.Y(n_3776)
);

AOI21xp5_ASAP7_75t_L g3777 ( 
.A1(n_3628),
.A2(n_1709),
.B(n_1703),
.Y(n_3777)
);

INVx1_ASAP7_75t_L g3778 ( 
.A(n_3501),
.Y(n_3778)
);

INVx1_ASAP7_75t_L g3779 ( 
.A(n_3518),
.Y(n_3779)
);

OR2x2_ASAP7_75t_SL g3780 ( 
.A(n_3572),
.B(n_51),
.Y(n_3780)
);

NAND2xp5_ASAP7_75t_L g3781 ( 
.A(n_3551),
.B(n_54),
.Y(n_3781)
);

INVx1_ASAP7_75t_SL g3782 ( 
.A(n_3630),
.Y(n_3782)
);

BUFx2_ASAP7_75t_L g3783 ( 
.A(n_3519),
.Y(n_3783)
);

INVx1_ASAP7_75t_L g3784 ( 
.A(n_3518),
.Y(n_3784)
);

NAND2xp5_ASAP7_75t_L g3785 ( 
.A(n_3514),
.B(n_54),
.Y(n_3785)
);

OR2x2_ASAP7_75t_SL g3786 ( 
.A(n_3635),
.B(n_55),
.Y(n_3786)
);

INVx2_ASAP7_75t_L g3787 ( 
.A(n_3560),
.Y(n_3787)
);

INVx8_ASAP7_75t_L g3788 ( 
.A(n_3578),
.Y(n_3788)
);

A2O1A1Ixp33_ASAP7_75t_L g3789 ( 
.A1(n_3472),
.A2(n_58),
.B(n_56),
.C(n_57),
.Y(n_3789)
);

INVx2_ASAP7_75t_SL g3790 ( 
.A(n_3635),
.Y(n_3790)
);

OR2x6_ASAP7_75t_L g3791 ( 
.A(n_3544),
.B(n_1703),
.Y(n_3791)
);

OR2x6_ASAP7_75t_L g3792 ( 
.A(n_3620),
.B(n_1925),
.Y(n_3792)
);

BUFx2_ASAP7_75t_L g3793 ( 
.A(n_3519),
.Y(n_3793)
);

AND2x6_ASAP7_75t_L g3794 ( 
.A(n_3630),
.B(n_1709),
.Y(n_3794)
);

INVx6_ASAP7_75t_L g3795 ( 
.A(n_3578),
.Y(n_3795)
);

AOI21xp5_ASAP7_75t_L g3796 ( 
.A1(n_3492),
.A2(n_3451),
.B(n_3434),
.Y(n_3796)
);

HB1xp67_ASAP7_75t_L g3797 ( 
.A(n_3625),
.Y(n_3797)
);

AOI21xp5_ASAP7_75t_L g3798 ( 
.A1(n_3451),
.A2(n_1721),
.B(n_1709),
.Y(n_3798)
);

OR2x6_ASAP7_75t_L g3799 ( 
.A(n_3635),
.B(n_1721),
.Y(n_3799)
);

INVx1_ASAP7_75t_L g3800 ( 
.A(n_3518),
.Y(n_3800)
);

AOI21xp33_ASAP7_75t_L g3801 ( 
.A1(n_3453),
.A2(n_56),
.B(n_57),
.Y(n_3801)
);

CKINVDCx5p33_ASAP7_75t_R g3802 ( 
.A(n_3602),
.Y(n_3802)
);

AND2x2_ASAP7_75t_L g3803 ( 
.A(n_3514),
.B(n_58),
.Y(n_3803)
);

OAI22xp5_ASAP7_75t_L g3804 ( 
.A1(n_3581),
.A2(n_3500),
.B1(n_3578),
.B2(n_3605),
.Y(n_3804)
);

A2O1A1Ixp33_ASAP7_75t_L g3805 ( 
.A1(n_3450),
.A2(n_3542),
.B(n_3642),
.C(n_3610),
.Y(n_3805)
);

AOI22xp33_ASAP7_75t_L g3806 ( 
.A1(n_3585),
.A2(n_1560),
.B1(n_1654),
.B2(n_1620),
.Y(n_3806)
);

NAND2x1p5_ASAP7_75t_L g3807 ( 
.A(n_3516),
.B(n_1721),
.Y(n_3807)
);

INVx2_ASAP7_75t_SL g3808 ( 
.A(n_3516),
.Y(n_3808)
);

AND2x2_ASAP7_75t_L g3809 ( 
.A(n_3595),
.B(n_59),
.Y(n_3809)
);

NOR2xp33_ASAP7_75t_SL g3810 ( 
.A(n_3592),
.B(n_1479),
.Y(n_3810)
);

INVx1_ASAP7_75t_L g3811 ( 
.A(n_3468),
.Y(n_3811)
);

AND3x1_ASAP7_75t_SL g3812 ( 
.A(n_3482),
.B(n_59),
.C(n_61),
.Y(n_3812)
);

OAI22xp5_ASAP7_75t_L g3813 ( 
.A1(n_3500),
.A2(n_1742),
.B1(n_1750),
.B2(n_1721),
.Y(n_3813)
);

INVx1_ASAP7_75t_SL g3814 ( 
.A(n_3606),
.Y(n_3814)
);

INVx1_ASAP7_75t_L g3815 ( 
.A(n_3468),
.Y(n_3815)
);

BUFx6f_ASAP7_75t_L g3816 ( 
.A(n_3609),
.Y(n_3816)
);

BUFx12f_ASAP7_75t_L g3817 ( 
.A(n_3538),
.Y(n_3817)
);

HB1xp67_ASAP7_75t_L g3818 ( 
.A(n_3468),
.Y(n_3818)
);

OAI22x1_ASAP7_75t_L g3819 ( 
.A1(n_3483),
.A2(n_64),
.B1(n_62),
.B2(n_63),
.Y(n_3819)
);

INVx1_ASAP7_75t_L g3820 ( 
.A(n_3561),
.Y(n_3820)
);

AOI22xp33_ASAP7_75t_L g3821 ( 
.A1(n_3579),
.A2(n_1560),
.B1(n_1654),
.B2(n_1620),
.Y(n_3821)
);

INVx1_ASAP7_75t_L g3822 ( 
.A(n_3447),
.Y(n_3822)
);

INVx1_ASAP7_75t_SL g3823 ( 
.A(n_3618),
.Y(n_3823)
);

INVx2_ASAP7_75t_L g3824 ( 
.A(n_3447),
.Y(n_3824)
);

NOR2xp33_ASAP7_75t_L g3825 ( 
.A(n_3562),
.B(n_63),
.Y(n_3825)
);

CKINVDCx5p33_ASAP7_75t_R g3826 ( 
.A(n_3576),
.Y(n_3826)
);

AND2x2_ASAP7_75t_L g3827 ( 
.A(n_3489),
.B(n_64),
.Y(n_3827)
);

INVx1_ASAP7_75t_SL g3828 ( 
.A(n_3577),
.Y(n_3828)
);

INVx1_ASAP7_75t_L g3829 ( 
.A(n_3447),
.Y(n_3829)
);

NAND2xp5_ASAP7_75t_SL g3830 ( 
.A(n_3558),
.B(n_1479),
.Y(n_3830)
);

INVx4_ASAP7_75t_L g3831 ( 
.A(n_3627),
.Y(n_3831)
);

BUFx2_ASAP7_75t_L g3832 ( 
.A(n_3612),
.Y(n_3832)
);

BUFx2_ASAP7_75t_L g3833 ( 
.A(n_3616),
.Y(n_3833)
);

BUFx10_ASAP7_75t_L g3834 ( 
.A(n_3608),
.Y(n_3834)
);

OAI21xp5_ASAP7_75t_L g3835 ( 
.A1(n_3570),
.A2(n_1560),
.B(n_1654),
.Y(n_3835)
);

OAI22xp33_ASAP7_75t_L g3836 ( 
.A1(n_3640),
.A2(n_67),
.B1(n_65),
.B2(n_66),
.Y(n_3836)
);

NAND2xp5_ASAP7_75t_L g3837 ( 
.A(n_3586),
.B(n_65),
.Y(n_3837)
);

NAND2xp5_ASAP7_75t_L g3838 ( 
.A(n_3457),
.B(n_66),
.Y(n_3838)
);

INVxp67_ASAP7_75t_L g3839 ( 
.A(n_3465),
.Y(n_3839)
);

AND2x4_ASAP7_75t_L g3840 ( 
.A(n_3600),
.B(n_311),
.Y(n_3840)
);

OAI22xp5_ASAP7_75t_L g3841 ( 
.A1(n_3568),
.A2(n_1750),
.B1(n_1772),
.B2(n_1742),
.Y(n_3841)
);

NAND2xp5_ASAP7_75t_L g3842 ( 
.A(n_3457),
.B(n_68),
.Y(n_3842)
);

AOI22xp5_ASAP7_75t_L g3843 ( 
.A1(n_3623),
.A2(n_1654),
.B1(n_1479),
.B2(n_1508),
.Y(n_3843)
);

AND2x2_ASAP7_75t_L g3844 ( 
.A(n_3627),
.B(n_69),
.Y(n_3844)
);

OA21x2_ASAP7_75t_L g3845 ( 
.A1(n_3621),
.A2(n_70),
.B(n_71),
.Y(n_3845)
);

AOI22xp5_ASAP7_75t_L g3846 ( 
.A1(n_3487),
.A2(n_1654),
.B1(n_1480),
.B2(n_1524),
.Y(n_3846)
);

NAND2xp5_ASAP7_75t_L g3847 ( 
.A(n_3511),
.B(n_71),
.Y(n_3847)
);

O2A1O1Ixp5_ASAP7_75t_SL g3848 ( 
.A1(n_3539),
.A2(n_74),
.B(n_72),
.C(n_73),
.Y(n_3848)
);

AND2x4_ASAP7_75t_L g3849 ( 
.A(n_3607),
.B(n_313),
.Y(n_3849)
);

AND2x2_ASAP7_75t_L g3850 ( 
.A(n_3473),
.B(n_74),
.Y(n_3850)
);

INVx2_ASAP7_75t_SL g3851 ( 
.A(n_3444),
.Y(n_3851)
);

CKINVDCx20_ASAP7_75t_R g3852 ( 
.A(n_3537),
.Y(n_3852)
);

NOR2xp33_ASAP7_75t_L g3853 ( 
.A(n_3631),
.B(n_75),
.Y(n_3853)
);

INVx2_ASAP7_75t_SL g3854 ( 
.A(n_3535),
.Y(n_3854)
);

CKINVDCx5p33_ASAP7_75t_R g3855 ( 
.A(n_3593),
.Y(n_3855)
);

INVx1_ASAP7_75t_L g3856 ( 
.A(n_3436),
.Y(n_3856)
);

NAND2xp33_ASAP7_75t_L g3857 ( 
.A(n_3614),
.B(n_1742),
.Y(n_3857)
);

AND2x2_ASAP7_75t_L g3858 ( 
.A(n_3436),
.B(n_75),
.Y(n_3858)
);

AND2x2_ASAP7_75t_SL g3859 ( 
.A(n_3574),
.B(n_3434),
.Y(n_3859)
);

A2O1A1Ixp33_ASAP7_75t_L g3860 ( 
.A1(n_3541),
.A2(n_79),
.B(n_76),
.C(n_78),
.Y(n_3860)
);

INVx1_ASAP7_75t_L g3861 ( 
.A(n_3436),
.Y(n_3861)
);

BUFx3_ASAP7_75t_L g3862 ( 
.A(n_3532),
.Y(n_3862)
);

AOI22xp33_ASAP7_75t_L g3863 ( 
.A1(n_3622),
.A2(n_3587),
.B1(n_3527),
.B2(n_3460),
.Y(n_3863)
);

INVx2_ASAP7_75t_SL g3864 ( 
.A(n_3470),
.Y(n_3864)
);

INVx2_ASAP7_75t_L g3865 ( 
.A(n_3449),
.Y(n_3865)
);

NAND2xp5_ASAP7_75t_L g3866 ( 
.A(n_3643),
.B(n_76),
.Y(n_3866)
);

INVx1_ASAP7_75t_L g3867 ( 
.A(n_3664),
.Y(n_3867)
);

INVx1_ASAP7_75t_L g3868 ( 
.A(n_3664),
.Y(n_3868)
);

OAI22xp5_ASAP7_75t_L g3869 ( 
.A1(n_3658),
.A2(n_3574),
.B1(n_3626),
.B2(n_3567),
.Y(n_3869)
);

INVx2_ASAP7_75t_L g3870 ( 
.A(n_3674),
.Y(n_3870)
);

INVx1_ASAP7_75t_L g3871 ( 
.A(n_3674),
.Y(n_3871)
);

CKINVDCx16_ASAP7_75t_R g3872 ( 
.A(n_3761),
.Y(n_3872)
);

BUFx10_ASAP7_75t_L g3873 ( 
.A(n_3676),
.Y(n_3873)
);

OAI21xp5_ASAP7_75t_SL g3874 ( 
.A1(n_3689),
.A2(n_78),
.B(n_79),
.Y(n_3874)
);

AOI22xp33_ASAP7_75t_SL g3875 ( 
.A1(n_3850),
.A2(n_3437),
.B1(n_3591),
.B2(n_3522),
.Y(n_3875)
);

INVxp67_ASAP7_75t_SL g3876 ( 
.A(n_3708),
.Y(n_3876)
);

CKINVDCx5p33_ASAP7_75t_R g3877 ( 
.A(n_3662),
.Y(n_3877)
);

INVx1_ASAP7_75t_L g3878 ( 
.A(n_3667),
.Y(n_3878)
);

INVx6_ASAP7_75t_L g3879 ( 
.A(n_3759),
.Y(n_3879)
);

BUFx3_ASAP7_75t_L g3880 ( 
.A(n_3766),
.Y(n_3880)
);

INVx3_ASAP7_75t_L g3881 ( 
.A(n_3648),
.Y(n_3881)
);

OAI22xp5_ASAP7_75t_L g3882 ( 
.A1(n_3786),
.A2(n_3780),
.B1(n_3781),
.B2(n_3773),
.Y(n_3882)
);

INVx1_ASAP7_75t_L g3883 ( 
.A(n_3672),
.Y(n_3883)
);

CKINVDCx11_ASAP7_75t_R g3884 ( 
.A(n_3675),
.Y(n_3884)
);

CKINVDCx11_ASAP7_75t_R g3885 ( 
.A(n_3769),
.Y(n_3885)
);

INVx1_ASAP7_75t_L g3886 ( 
.A(n_3649),
.Y(n_3886)
);

INVx2_ASAP7_75t_L g3887 ( 
.A(n_3721),
.Y(n_3887)
);

AOI22xp33_ASAP7_75t_L g3888 ( 
.A1(n_3714),
.A2(n_3495),
.B1(n_3509),
.B2(n_3491),
.Y(n_3888)
);

NAND2xp5_ASAP7_75t_L g3889 ( 
.A(n_3656),
.B(n_3643),
.Y(n_3889)
);

NAND2x1p5_ASAP7_75t_L g3890 ( 
.A(n_3742),
.B(n_3462),
.Y(n_3890)
);

OAI22xp5_ASAP7_75t_L g3891 ( 
.A1(n_3789),
.A2(n_3603),
.B1(n_3638),
.B2(n_84),
.Y(n_3891)
);

INVx1_ASAP7_75t_L g3892 ( 
.A(n_3649),
.Y(n_3892)
);

CKINVDCx20_ASAP7_75t_R g3893 ( 
.A(n_3747),
.Y(n_3893)
);

AOI22xp5_ASAP7_75t_L g3894 ( 
.A1(n_3812),
.A2(n_3530),
.B1(n_3536),
.B2(n_3554),
.Y(n_3894)
);

INVx6_ASAP7_75t_L g3895 ( 
.A(n_3660),
.Y(n_3895)
);

AOI22xp33_ASAP7_75t_SL g3896 ( 
.A1(n_3646),
.A2(n_3550),
.B1(n_3566),
.B2(n_3469),
.Y(n_3896)
);

INVx3_ASAP7_75t_L g3897 ( 
.A(n_3648),
.Y(n_3897)
);

INVx1_ASAP7_75t_SL g3898 ( 
.A(n_3650),
.Y(n_3898)
);

NAND2xp33_ASAP7_75t_SL g3899 ( 
.A(n_3700),
.B(n_80),
.Y(n_3899)
);

AOI22xp33_ASAP7_75t_SL g3900 ( 
.A1(n_3852),
.A2(n_3505),
.B1(n_86),
.B2(n_80),
.Y(n_3900)
);

BUFx2_ASAP7_75t_SL g3901 ( 
.A(n_3670),
.Y(n_3901)
);

BUFx2_ASAP7_75t_L g3902 ( 
.A(n_3647),
.Y(n_3902)
);

CKINVDCx5p33_ASAP7_75t_R g3903 ( 
.A(n_3802),
.Y(n_3903)
);

OAI22xp5_ASAP7_75t_L g3904 ( 
.A1(n_3860),
.A2(n_88),
.B1(n_81),
.B2(n_87),
.Y(n_3904)
);

AOI22xp33_ASAP7_75t_L g3905 ( 
.A1(n_3764),
.A2(n_1508),
.B1(n_1524),
.B2(n_1480),
.Y(n_3905)
);

AND2x2_ASAP7_75t_L g3906 ( 
.A(n_3652),
.B(n_3643),
.Y(n_3906)
);

AOI22xp33_ASAP7_75t_L g3907 ( 
.A1(n_3752),
.A2(n_1508),
.B1(n_1524),
.B2(n_1480),
.Y(n_3907)
);

INVx1_ASAP7_75t_L g3908 ( 
.A(n_3653),
.Y(n_3908)
);

INVx3_ASAP7_75t_L g3909 ( 
.A(n_3692),
.Y(n_3909)
);

OAI22xp5_ASAP7_75t_L g3910 ( 
.A1(n_3805),
.A2(n_91),
.B1(n_89),
.B2(n_90),
.Y(n_3910)
);

BUFx3_ASAP7_75t_L g3911 ( 
.A(n_3726),
.Y(n_3911)
);

BUFx10_ASAP7_75t_L g3912 ( 
.A(n_3771),
.Y(n_3912)
);

BUFx6f_ASAP7_75t_L g3913 ( 
.A(n_3660),
.Y(n_3913)
);

OAI22xp5_ASAP7_75t_L g3914 ( 
.A1(n_3839),
.A2(n_92),
.B1(n_89),
.B2(n_91),
.Y(n_3914)
);

CKINVDCx14_ASAP7_75t_R g3915 ( 
.A(n_3755),
.Y(n_3915)
);

INVx2_ASAP7_75t_L g3916 ( 
.A(n_3692),
.Y(n_3916)
);

BUFx8_ASAP7_75t_L g3917 ( 
.A(n_3803),
.Y(n_3917)
);

AOI22xp33_ASAP7_75t_L g3918 ( 
.A1(n_3801),
.A2(n_1508),
.B1(n_1524),
.B2(n_1480),
.Y(n_3918)
);

NAND2xp5_ASAP7_75t_L g3919 ( 
.A(n_3814),
.B(n_93),
.Y(n_3919)
);

BUFx2_ASAP7_75t_SL g3920 ( 
.A(n_3741),
.Y(n_3920)
);

INVx4_ASAP7_75t_L g3921 ( 
.A(n_3788),
.Y(n_3921)
);

INVx2_ASAP7_75t_L g3922 ( 
.A(n_3718),
.Y(n_3922)
);

INVx2_ASAP7_75t_L g3923 ( 
.A(n_3666),
.Y(n_3923)
);

CKINVDCx11_ASAP7_75t_R g3924 ( 
.A(n_3644),
.Y(n_3924)
);

CKINVDCx5p33_ASAP7_75t_R g3925 ( 
.A(n_3776),
.Y(n_3925)
);

INVx3_ASAP7_75t_L g3926 ( 
.A(n_3795),
.Y(n_3926)
);

CKINVDCx11_ASAP7_75t_R g3927 ( 
.A(n_3691),
.Y(n_3927)
);

INVx1_ASAP7_75t_L g3928 ( 
.A(n_3653),
.Y(n_3928)
);

INVx1_ASAP7_75t_L g3929 ( 
.A(n_3654),
.Y(n_3929)
);

INVx4_ASAP7_75t_L g3930 ( 
.A(n_3788),
.Y(n_3930)
);

INVx2_ASAP7_75t_L g3931 ( 
.A(n_3686),
.Y(n_3931)
);

CKINVDCx8_ASAP7_75t_R g3932 ( 
.A(n_3660),
.Y(n_3932)
);

OAI22xp5_ASAP7_75t_L g3933 ( 
.A1(n_3661),
.A2(n_96),
.B1(n_94),
.B2(n_95),
.Y(n_3933)
);

INVx2_ASAP7_75t_L g3934 ( 
.A(n_3693),
.Y(n_3934)
);

INVx2_ASAP7_75t_R g3935 ( 
.A(n_3708),
.Y(n_3935)
);

INVx6_ASAP7_75t_L g3936 ( 
.A(n_3698),
.Y(n_3936)
);

OAI22xp33_ASAP7_75t_R g3937 ( 
.A1(n_3657),
.A2(n_100),
.B1(n_95),
.B2(n_97),
.Y(n_3937)
);

INVx3_ASAP7_75t_L g3938 ( 
.A(n_3795),
.Y(n_3938)
);

INVx2_ASAP7_75t_SL g3939 ( 
.A(n_3698),
.Y(n_3939)
);

INVx1_ASAP7_75t_L g3940 ( 
.A(n_3654),
.Y(n_3940)
);

INVx1_ASAP7_75t_L g3941 ( 
.A(n_3679),
.Y(n_3941)
);

INVx1_ASAP7_75t_SL g3942 ( 
.A(n_3728),
.Y(n_3942)
);

AOI22xp33_ASAP7_75t_L g3943 ( 
.A1(n_3817),
.A2(n_1538),
.B1(n_1750),
.B2(n_1742),
.Y(n_3943)
);

AOI22xp33_ASAP7_75t_L g3944 ( 
.A1(n_3760),
.A2(n_1538),
.B1(n_1925),
.B2(n_1772),
.Y(n_3944)
);

AOI22xp33_ASAP7_75t_SL g3945 ( 
.A1(n_3746),
.A2(n_101),
.B1(n_97),
.B2(n_100),
.Y(n_3945)
);

AOI22xp33_ASAP7_75t_L g3946 ( 
.A1(n_3740),
.A2(n_1538),
.B1(n_1925),
.B2(n_1772),
.Y(n_3946)
);

AOI22xp5_ASAP7_75t_L g3947 ( 
.A1(n_3836),
.A2(n_103),
.B1(n_101),
.B2(n_102),
.Y(n_3947)
);

INVx1_ASAP7_75t_L g3948 ( 
.A(n_3679),
.Y(n_3948)
);

AOI22xp33_ASAP7_75t_L g3949 ( 
.A1(n_3804),
.A2(n_1538),
.B1(n_1772),
.B2(n_1750),
.Y(n_3949)
);

OAI22xp33_ASAP7_75t_L g3950 ( 
.A1(n_3717),
.A2(n_107),
.B1(n_104),
.B2(n_106),
.Y(n_3950)
);

OAI22xp33_ASAP7_75t_L g3951 ( 
.A1(n_3757),
.A2(n_108),
.B1(n_104),
.B2(n_106),
.Y(n_3951)
);

INVx1_ASAP7_75t_L g3952 ( 
.A(n_3713),
.Y(n_3952)
);

OAI22xp33_ASAP7_75t_L g3953 ( 
.A1(n_3782),
.A2(n_111),
.B1(n_109),
.B2(n_110),
.Y(n_3953)
);

AOI22xp33_ASAP7_75t_L g3954 ( 
.A1(n_3768),
.A2(n_1925),
.B1(n_1784),
.B2(n_1787),
.Y(n_3954)
);

INVx4_ASAP7_75t_L g3955 ( 
.A(n_3698),
.Y(n_3955)
);

INVx6_ASAP7_75t_L g3956 ( 
.A(n_3706),
.Y(n_3956)
);

AND2x2_ASAP7_75t_L g3957 ( 
.A(n_3699),
.B(n_109),
.Y(n_3957)
);

OAI22xp33_ASAP7_75t_L g3958 ( 
.A1(n_3826),
.A2(n_115),
.B1(n_112),
.B2(n_114),
.Y(n_3958)
);

AOI22xp33_ASAP7_75t_L g3959 ( 
.A1(n_3771),
.A2(n_1898),
.B1(n_1784),
.B2(n_1787),
.Y(n_3959)
);

AOI22xp33_ASAP7_75t_SL g3960 ( 
.A1(n_3746),
.A2(n_117),
.B1(n_112),
.B2(n_116),
.Y(n_3960)
);

INVx2_ASAP7_75t_L g3961 ( 
.A(n_3724),
.Y(n_3961)
);

INVx3_ASAP7_75t_SL g3962 ( 
.A(n_3709),
.Y(n_3962)
);

AOI22xp33_ASAP7_75t_L g3963 ( 
.A1(n_3668),
.A2(n_1784),
.B1(n_1787),
.B2(n_1780),
.Y(n_3963)
);

AOI22xp33_ASAP7_75t_L g3964 ( 
.A1(n_3862),
.A2(n_1784),
.B1(n_1787),
.B2(n_1780),
.Y(n_3964)
);

CKINVDCx11_ASAP7_75t_R g3965 ( 
.A(n_3707),
.Y(n_3965)
);

NAND2xp5_ASAP7_75t_L g3966 ( 
.A(n_3823),
.B(n_116),
.Y(n_3966)
);

OAI22xp5_ASAP7_75t_L g3967 ( 
.A1(n_3734),
.A2(n_119),
.B1(n_117),
.B2(n_118),
.Y(n_3967)
);

CKINVDCx20_ASAP7_75t_R g3968 ( 
.A(n_3808),
.Y(n_3968)
);

AOI22xp33_ASAP7_75t_L g3969 ( 
.A1(n_3853),
.A2(n_1898),
.B1(n_1794),
.B2(n_1798),
.Y(n_3969)
);

BUFx8_ASAP7_75t_L g3970 ( 
.A(n_3659),
.Y(n_3970)
);

HB1xp67_ASAP7_75t_L g3971 ( 
.A(n_3713),
.Y(n_3971)
);

INVx1_ASAP7_75t_L g3972 ( 
.A(n_3710),
.Y(n_3972)
);

INVx1_ASAP7_75t_L g3973 ( 
.A(n_3787),
.Y(n_3973)
);

INVx1_ASAP7_75t_L g3974 ( 
.A(n_3797),
.Y(n_3974)
);

INVx2_ASAP7_75t_L g3975 ( 
.A(n_3738),
.Y(n_3975)
);

AOI22xp33_ASAP7_75t_SL g3976 ( 
.A1(n_3827),
.A2(n_123),
.B1(n_118),
.B2(n_120),
.Y(n_3976)
);

INVx2_ASAP7_75t_L g3977 ( 
.A(n_3739),
.Y(n_3977)
);

INVx1_ASAP7_75t_L g3978 ( 
.A(n_3820),
.Y(n_3978)
);

INVx2_ASAP7_75t_L g3979 ( 
.A(n_3750),
.Y(n_3979)
);

OAI22xp33_ASAP7_75t_L g3980 ( 
.A1(n_3680),
.A2(n_132),
.B1(n_124),
.B2(n_125),
.Y(n_3980)
);

INVx4_ASAP7_75t_L g3981 ( 
.A(n_3706),
.Y(n_3981)
);

BUFx10_ASAP7_75t_L g3982 ( 
.A(n_3825),
.Y(n_3982)
);

AOI22xp33_ASAP7_75t_L g3983 ( 
.A1(n_3735),
.A2(n_1794),
.B1(n_1798),
.B2(n_1780),
.Y(n_3983)
);

BUFx2_ASAP7_75t_SL g3984 ( 
.A(n_3665),
.Y(n_3984)
);

INVx1_ASAP7_75t_L g3985 ( 
.A(n_3753),
.Y(n_3985)
);

AOI22xp33_ASAP7_75t_SL g3986 ( 
.A1(n_3655),
.A2(n_134),
.B1(n_124),
.B2(n_133),
.Y(n_3986)
);

INVx1_ASAP7_75t_L g3987 ( 
.A(n_3866),
.Y(n_3987)
);

INVx1_ASAP7_75t_L g3988 ( 
.A(n_3858),
.Y(n_3988)
);

BUFx12f_ASAP7_75t_L g3989 ( 
.A(n_3725),
.Y(n_3989)
);

BUFx3_ASAP7_75t_L g3990 ( 
.A(n_3706),
.Y(n_3990)
);

BUFx12f_ASAP7_75t_L g3991 ( 
.A(n_3688),
.Y(n_3991)
);

BUFx3_ASAP7_75t_L g3992 ( 
.A(n_3715),
.Y(n_3992)
);

BUFx3_ASAP7_75t_L g3993 ( 
.A(n_3715),
.Y(n_3993)
);

AND2x2_ASAP7_75t_L g3994 ( 
.A(n_3783),
.B(n_135),
.Y(n_3994)
);

NAND2xp5_ASAP7_75t_L g3995 ( 
.A(n_3828),
.B(n_135),
.Y(n_3995)
);

NAND2xp5_ASAP7_75t_L g3996 ( 
.A(n_3838),
.B(n_136),
.Y(n_3996)
);

INVx1_ASAP7_75t_L g3997 ( 
.A(n_3842),
.Y(n_3997)
);

BUFx4f_ASAP7_75t_SL g3998 ( 
.A(n_3737),
.Y(n_3998)
);

BUFx12f_ASAP7_75t_L g3999 ( 
.A(n_3690),
.Y(n_3999)
);

INVx2_ASAP7_75t_L g4000 ( 
.A(n_3793),
.Y(n_4000)
);

BUFx2_ASAP7_75t_L g4001 ( 
.A(n_3737),
.Y(n_4001)
);

INVx1_ASAP7_75t_L g4002 ( 
.A(n_3778),
.Y(n_4002)
);

CKINVDCx20_ASAP7_75t_R g4003 ( 
.A(n_3790),
.Y(n_4003)
);

INVx1_ASAP7_75t_SL g4004 ( 
.A(n_3651),
.Y(n_4004)
);

BUFx2_ASAP7_75t_L g4005 ( 
.A(n_3756),
.Y(n_4005)
);

AOI22xp33_ASAP7_75t_L g4006 ( 
.A1(n_3681),
.A2(n_1794),
.B1(n_1798),
.B2(n_1780),
.Y(n_4006)
);

INVx2_ASAP7_75t_L g4007 ( 
.A(n_3756),
.Y(n_4007)
);

AND2x2_ASAP7_75t_L g4008 ( 
.A(n_3701),
.B(n_136),
.Y(n_4008)
);

NAND2xp5_ASAP7_75t_L g4009 ( 
.A(n_3645),
.B(n_138),
.Y(n_4009)
);

INVx3_ASAP7_75t_L g4010 ( 
.A(n_3816),
.Y(n_4010)
);

BUFx4f_ASAP7_75t_SL g4011 ( 
.A(n_3762),
.Y(n_4011)
);

CKINVDCx20_ASAP7_75t_R g4012 ( 
.A(n_3733),
.Y(n_4012)
);

INVx2_ASAP7_75t_L g4013 ( 
.A(n_3832),
.Y(n_4013)
);

INVx1_ASAP7_75t_L g4014 ( 
.A(n_3778),
.Y(n_4014)
);

OAI22xp33_ASAP7_75t_L g4015 ( 
.A1(n_3767),
.A2(n_141),
.B1(n_138),
.B2(n_140),
.Y(n_4015)
);

BUFx6f_ASAP7_75t_SL g4016 ( 
.A(n_3681),
.Y(n_4016)
);

INVx2_ASAP7_75t_L g4017 ( 
.A(n_3833),
.Y(n_4017)
);

INVx1_ASAP7_75t_L g4018 ( 
.A(n_3811),
.Y(n_4018)
);

BUFx2_ASAP7_75t_L g4019 ( 
.A(n_3792),
.Y(n_4019)
);

CKINVDCx20_ASAP7_75t_R g4020 ( 
.A(n_3723),
.Y(n_4020)
);

CKINVDCx14_ASAP7_75t_R g4021 ( 
.A(n_3794),
.Y(n_4021)
);

AOI22xp33_ASAP7_75t_SL g4022 ( 
.A1(n_3794),
.A2(n_142),
.B1(n_140),
.B2(n_141),
.Y(n_4022)
);

OAI22xp5_ASAP7_75t_L g4023 ( 
.A1(n_3775),
.A2(n_144),
.B1(n_142),
.B2(n_143),
.Y(n_4023)
);

AOI22xp5_ASAP7_75t_L g4024 ( 
.A1(n_3722),
.A2(n_147),
.B1(n_143),
.B2(n_146),
.Y(n_4024)
);

NAND2xp5_ASAP7_75t_SL g4025 ( 
.A(n_3855),
.B(n_1412),
.Y(n_4025)
);

INVx1_ASAP7_75t_L g4026 ( 
.A(n_3815),
.Y(n_4026)
);

BUFx10_ASAP7_75t_L g4027 ( 
.A(n_3849),
.Y(n_4027)
);

AND2x2_ASAP7_75t_L g4028 ( 
.A(n_3809),
.B(n_147),
.Y(n_4028)
);

CKINVDCx11_ASAP7_75t_R g4029 ( 
.A(n_3834),
.Y(n_4029)
);

AOI22xp33_ASAP7_75t_L g4030 ( 
.A1(n_3749),
.A2(n_1798),
.B1(n_1819),
.B2(n_1794),
.Y(n_4030)
);

AOI22xp33_ASAP7_75t_L g4031 ( 
.A1(n_3736),
.A2(n_1824),
.B1(n_1836),
.B2(n_1819),
.Y(n_4031)
);

INVx2_ASAP7_75t_L g4032 ( 
.A(n_3816),
.Y(n_4032)
);

BUFx12f_ASAP7_75t_L g4033 ( 
.A(n_3678),
.Y(n_4033)
);

INVx1_ASAP7_75t_L g4034 ( 
.A(n_3770),
.Y(n_4034)
);

BUFx6f_ASAP7_75t_SL g4035 ( 
.A(n_3849),
.Y(n_4035)
);

BUFx12f_ASAP7_75t_L g4036 ( 
.A(n_3682),
.Y(n_4036)
);

INVx1_ASAP7_75t_L g4037 ( 
.A(n_3772),
.Y(n_4037)
);

BUFx12f_ASAP7_75t_L g4038 ( 
.A(n_3799),
.Y(n_4038)
);

BUFx2_ASAP7_75t_L g4039 ( 
.A(n_3792),
.Y(n_4039)
);

INVx1_ASAP7_75t_L g4040 ( 
.A(n_3856),
.Y(n_4040)
);

NAND2xp5_ASAP7_75t_L g4041 ( 
.A(n_3997),
.B(n_3844),
.Y(n_4041)
);

BUFx2_ASAP7_75t_L g4042 ( 
.A(n_3926),
.Y(n_4042)
);

HB1xp67_ASAP7_75t_L g4043 ( 
.A(n_3942),
.Y(n_4043)
);

NAND2xp5_ASAP7_75t_L g4044 ( 
.A(n_3987),
.B(n_3847),
.Y(n_4044)
);

CKINVDCx20_ASAP7_75t_R g4045 ( 
.A(n_3884),
.Y(n_4045)
);

AOI21xp5_ASAP7_75t_SL g4046 ( 
.A1(n_3910),
.A2(n_3729),
.B(n_3819),
.Y(n_4046)
);

OR2x2_ASAP7_75t_L g4047 ( 
.A(n_3988),
.B(n_3818),
.Y(n_4047)
);

INVx2_ASAP7_75t_L g4048 ( 
.A(n_3870),
.Y(n_4048)
);

INVx3_ASAP7_75t_SL g4049 ( 
.A(n_3877),
.Y(n_4049)
);

NAND2xp5_ASAP7_75t_L g4050 ( 
.A(n_3972),
.B(n_3663),
.Y(n_4050)
);

OA21x2_ASAP7_75t_L g4051 ( 
.A1(n_3974),
.A2(n_3765),
.B(n_3779),
.Y(n_4051)
);

INVx1_ASAP7_75t_L g4052 ( 
.A(n_3886),
.Y(n_4052)
);

BUFx3_ASAP7_75t_L g4053 ( 
.A(n_3880),
.Y(n_4053)
);

AND2x2_ASAP7_75t_L g4054 ( 
.A(n_3898),
.B(n_3864),
.Y(n_4054)
);

OA21x2_ASAP7_75t_L g4055 ( 
.A1(n_4040),
.A2(n_3779),
.B(n_3856),
.Y(n_4055)
);

OR2x2_ASAP7_75t_L g4056 ( 
.A(n_3942),
.B(n_3822),
.Y(n_4056)
);

OAI22xp5_ASAP7_75t_L g4057 ( 
.A1(n_3874),
.A2(n_3685),
.B1(n_3695),
.B2(n_3683),
.Y(n_4057)
);

INVx1_ASAP7_75t_L g4058 ( 
.A(n_3892),
.Y(n_4058)
);

AND2x2_ASAP7_75t_L g4059 ( 
.A(n_3898),
.B(n_3831),
.Y(n_4059)
);

AND2x2_ASAP7_75t_L g4060 ( 
.A(n_4000),
.B(n_3902),
.Y(n_4060)
);

CKINVDCx5p33_ASAP7_75t_R g4061 ( 
.A(n_3885),
.Y(n_4061)
);

NAND2xp5_ASAP7_75t_L g4062 ( 
.A(n_3978),
.B(n_3704),
.Y(n_4062)
);

INVx3_ASAP7_75t_L g4063 ( 
.A(n_3926),
.Y(n_4063)
);

AOI21x1_ASAP7_75t_SL g4064 ( 
.A1(n_3889),
.A2(n_3785),
.B(n_3697),
.Y(n_4064)
);

OR2x2_ASAP7_75t_L g4065 ( 
.A(n_3867),
.B(n_3829),
.Y(n_4065)
);

NAND2xp5_ASAP7_75t_L g4066 ( 
.A(n_3961),
.B(n_3731),
.Y(n_4066)
);

OAI22xp5_ASAP7_75t_L g4067 ( 
.A1(n_3874),
.A2(n_4024),
.B1(n_3947),
.B2(n_3882),
.Y(n_4067)
);

AOI21x1_ASAP7_75t_SL g4068 ( 
.A1(n_3996),
.A2(n_3837),
.B(n_3840),
.Y(n_4068)
);

AND2x2_ASAP7_75t_L g4069 ( 
.A(n_3868),
.B(n_3831),
.Y(n_4069)
);

AOI21xp5_ASAP7_75t_L g4070 ( 
.A1(n_3910),
.A2(n_3891),
.B(n_3716),
.Y(n_4070)
);

AOI21xp5_ASAP7_75t_SL g4071 ( 
.A1(n_4016),
.A2(n_3729),
.B(n_3711),
.Y(n_4071)
);

INVx2_ASAP7_75t_SL g4072 ( 
.A(n_3879),
.Y(n_4072)
);

NOR2xp67_ASAP7_75t_L g4073 ( 
.A(n_3938),
.B(n_3796),
.Y(n_4073)
);

OR2x2_ASAP7_75t_L g4074 ( 
.A(n_3871),
.B(n_3861),
.Y(n_4074)
);

AOI21xp5_ASAP7_75t_L g4075 ( 
.A1(n_3891),
.A2(n_3719),
.B(n_3830),
.Y(n_4075)
);

OAI22xp5_ASAP7_75t_L g4076 ( 
.A1(n_4024),
.A2(n_3711),
.B1(n_3806),
.B2(n_3798),
.Y(n_4076)
);

AOI21xp5_ASAP7_75t_L g4077 ( 
.A1(n_3904),
.A2(n_3754),
.B(n_3777),
.Y(n_4077)
);

HB1xp67_ASAP7_75t_L g4078 ( 
.A(n_3971),
.Y(n_4078)
);

AOI21x1_ASAP7_75t_SL g4079 ( 
.A1(n_3996),
.A2(n_3840),
.B(n_3834),
.Y(n_4079)
);

OA22x2_ASAP7_75t_L g4080 ( 
.A1(n_3882),
.A2(n_3791),
.B1(n_3774),
.B2(n_3763),
.Y(n_4080)
);

AOI21xp5_ASAP7_75t_L g4081 ( 
.A1(n_3904),
.A2(n_3857),
.B(n_3748),
.Y(n_4081)
);

AOI21xp5_ASAP7_75t_L g4082 ( 
.A1(n_3980),
.A2(n_3677),
.B(n_3694),
.Y(n_4082)
);

INVx1_ASAP7_75t_L g4083 ( 
.A(n_3908),
.Y(n_4083)
);

NAND2x1p5_ASAP7_75t_L g4084 ( 
.A(n_3938),
.B(n_3845),
.Y(n_4084)
);

AND2x2_ASAP7_75t_L g4085 ( 
.A(n_3915),
.B(n_4004),
.Y(n_4085)
);

AND2x2_ASAP7_75t_L g4086 ( 
.A(n_4004),
.B(n_3973),
.Y(n_4086)
);

AOI21xp5_ASAP7_75t_SL g4087 ( 
.A1(n_4016),
.A2(n_3791),
.B(n_3845),
.Y(n_4087)
);

HB1xp67_ASAP7_75t_L g4088 ( 
.A(n_4013),
.Y(n_4088)
);

AOI21xp5_ASAP7_75t_L g4089 ( 
.A1(n_4025),
.A2(n_3702),
.B(n_3712),
.Y(n_4089)
);

INVx2_ASAP7_75t_SL g4090 ( 
.A(n_3879),
.Y(n_4090)
);

HB1xp67_ASAP7_75t_L g4091 ( 
.A(n_4017),
.Y(n_4091)
);

NAND2xp5_ASAP7_75t_L g4092 ( 
.A(n_3985),
.B(n_3863),
.Y(n_4092)
);

BUFx2_ASAP7_75t_L g4093 ( 
.A(n_4001),
.Y(n_4093)
);

AND2x2_ASAP7_75t_L g4094 ( 
.A(n_3920),
.B(n_3851),
.Y(n_4094)
);

INVx2_ASAP7_75t_L g4095 ( 
.A(n_3881),
.Y(n_4095)
);

O2A1O1Ixp33_ASAP7_75t_L g4096 ( 
.A1(n_4023),
.A2(n_3687),
.B(n_3745),
.C(n_3671),
.Y(n_4096)
);

INVx4_ASAP7_75t_L g4097 ( 
.A(n_4011),
.Y(n_4097)
);

AOI21xp5_ASAP7_75t_L g4098 ( 
.A1(n_4015),
.A2(n_3835),
.B(n_3669),
.Y(n_4098)
);

AOI21xp5_ASAP7_75t_SL g4099 ( 
.A1(n_4035),
.A2(n_3703),
.B(n_3673),
.Y(n_4099)
);

INVx3_ASAP7_75t_SL g4100 ( 
.A(n_3903),
.Y(n_4100)
);

OR2x2_ASAP7_75t_L g4101 ( 
.A(n_3922),
.B(n_3861),
.Y(n_4101)
);

INVx2_ASAP7_75t_L g4102 ( 
.A(n_3881),
.Y(n_4102)
);

AOI21xp5_ASAP7_75t_SL g4103 ( 
.A1(n_4035),
.A2(n_3720),
.B(n_3732),
.Y(n_4103)
);

OAI22xp5_ASAP7_75t_L g4104 ( 
.A1(n_3947),
.A2(n_3807),
.B1(n_3846),
.B2(n_3859),
.Y(n_4104)
);

OAI22xp5_ASAP7_75t_L g4105 ( 
.A1(n_3976),
.A2(n_3841),
.B1(n_3800),
.B2(n_3784),
.Y(n_4105)
);

OAI22xp5_ASAP7_75t_L g4106 ( 
.A1(n_3986),
.A2(n_3743),
.B1(n_3744),
.B2(n_3727),
.Y(n_4106)
);

INVx2_ASAP7_75t_L g4107 ( 
.A(n_3897),
.Y(n_4107)
);

INVx2_ASAP7_75t_L g4108 ( 
.A(n_3897),
.Y(n_4108)
);

NAND2xp5_ASAP7_75t_L g4109 ( 
.A(n_3923),
.B(n_3854),
.Y(n_4109)
);

OAI22xp5_ASAP7_75t_L g4110 ( 
.A1(n_4022),
.A2(n_3727),
.B1(n_3730),
.B2(n_3843),
.Y(n_4110)
);

AND2x2_ASAP7_75t_L g4111 ( 
.A(n_3927),
.B(n_3865),
.Y(n_4111)
);

OAI22xp5_ASAP7_75t_L g4112 ( 
.A1(n_3945),
.A2(n_3824),
.B1(n_3799),
.B2(n_3705),
.Y(n_4112)
);

O2A1O1Ixp33_ASAP7_75t_L g4113 ( 
.A1(n_4023),
.A2(n_3967),
.B(n_3951),
.C(n_3914),
.Y(n_4113)
);

NAND2xp5_ASAP7_75t_L g4114 ( 
.A(n_3931),
.B(n_3848),
.Y(n_4114)
);

OAI22xp5_ASAP7_75t_L g4115 ( 
.A1(n_3960),
.A2(n_3751),
.B1(n_3816),
.B2(n_3813),
.Y(n_4115)
);

NAND2xp5_ASAP7_75t_L g4116 ( 
.A(n_3934),
.B(n_3684),
.Y(n_4116)
);

HB1xp67_ASAP7_75t_L g4117 ( 
.A(n_3916),
.Y(n_4117)
);

OAI22xp5_ASAP7_75t_L g4118 ( 
.A1(n_3900),
.A2(n_3821),
.B1(n_3794),
.B2(n_3810),
.Y(n_4118)
);

AOI21xp5_ASAP7_75t_L g4119 ( 
.A1(n_3869),
.A2(n_3696),
.B(n_3758),
.Y(n_4119)
);

CKINVDCx5p33_ASAP7_75t_R g4120 ( 
.A(n_3924),
.Y(n_4120)
);

AND2x2_ASAP7_75t_L g4121 ( 
.A(n_3965),
.B(n_3794),
.Y(n_4121)
);

NAND2x1p5_ASAP7_75t_L g4122 ( 
.A(n_3909),
.B(n_1819),
.Y(n_4122)
);

OAI22xp5_ASAP7_75t_L g4123 ( 
.A1(n_3967),
.A2(n_150),
.B1(n_148),
.B2(n_149),
.Y(n_4123)
);

BUFx2_ASAP7_75t_L g4124 ( 
.A(n_4005),
.Y(n_4124)
);

INVx1_ASAP7_75t_L g4125 ( 
.A(n_3928),
.Y(n_4125)
);

BUFx3_ASAP7_75t_L g4126 ( 
.A(n_3893),
.Y(n_4126)
);

OAI22xp5_ASAP7_75t_L g4127 ( 
.A1(n_3914),
.A2(n_151),
.B1(n_149),
.B2(n_150),
.Y(n_4127)
);

NAND2xp5_ASAP7_75t_L g4128 ( 
.A(n_3975),
.B(n_151),
.Y(n_4128)
);

NAND2xp5_ASAP7_75t_L g4129 ( 
.A(n_3977),
.B(n_154),
.Y(n_4129)
);

BUFx3_ASAP7_75t_L g4130 ( 
.A(n_3873),
.Y(n_4130)
);

CKINVDCx12_ASAP7_75t_R g4131 ( 
.A(n_4008),
.Y(n_4131)
);

OAI22xp5_ASAP7_75t_L g4132 ( 
.A1(n_3958),
.A2(n_157),
.B1(n_154),
.B2(n_156),
.Y(n_4132)
);

AOI21x1_ASAP7_75t_SL g4133 ( 
.A1(n_4009),
.A2(n_3906),
.B(n_3995),
.Y(n_4133)
);

INVx2_ASAP7_75t_L g4134 ( 
.A(n_3909),
.Y(n_4134)
);

AND2x2_ASAP7_75t_L g4135 ( 
.A(n_3901),
.B(n_159),
.Y(n_4135)
);

O2A1O1Ixp33_ASAP7_75t_L g4136 ( 
.A1(n_3953),
.A2(n_164),
.B(n_160),
.C(n_162),
.Y(n_4136)
);

HB1xp67_ASAP7_75t_L g4137 ( 
.A(n_3979),
.Y(n_4137)
);

AND2x2_ASAP7_75t_L g4138 ( 
.A(n_3872),
.B(n_160),
.Y(n_4138)
);

NAND2xp5_ASAP7_75t_L g4139 ( 
.A(n_3887),
.B(n_164),
.Y(n_4139)
);

INVx2_ASAP7_75t_SL g4140 ( 
.A(n_3911),
.Y(n_4140)
);

OA21x2_ASAP7_75t_L g4141 ( 
.A1(n_4002),
.A2(n_165),
.B(n_166),
.Y(n_4141)
);

NAND2xp5_ASAP7_75t_L g4142 ( 
.A(n_3878),
.B(n_166),
.Y(n_4142)
);

HB1xp67_ASAP7_75t_L g4143 ( 
.A(n_3952),
.Y(n_4143)
);

A2O1A1Ixp33_ASAP7_75t_L g4144 ( 
.A1(n_3899),
.A2(n_169),
.B(n_167),
.C(n_168),
.Y(n_4144)
);

INVx1_ASAP7_75t_L g4145 ( 
.A(n_3929),
.Y(n_4145)
);

INVx1_ASAP7_75t_L g4146 ( 
.A(n_3940),
.Y(n_4146)
);

OAI22xp5_ASAP7_75t_L g4147 ( 
.A1(n_3933),
.A2(n_170),
.B1(n_167),
.B2(n_169),
.Y(n_4147)
);

AOI21xp5_ASAP7_75t_SL g4148 ( 
.A1(n_3869),
.A2(n_3930),
.B(n_3921),
.Y(n_4148)
);

BUFx3_ASAP7_75t_L g4149 ( 
.A(n_3873),
.Y(n_4149)
);

AND2x2_ASAP7_75t_L g4150 ( 
.A(n_3962),
.B(n_170),
.Y(n_4150)
);

NAND2xp5_ASAP7_75t_L g4151 ( 
.A(n_3883),
.B(n_171),
.Y(n_4151)
);

NAND2xp5_ASAP7_75t_L g4152 ( 
.A(n_3941),
.B(n_172),
.Y(n_4152)
);

INVx2_ASAP7_75t_L g4153 ( 
.A(n_4007),
.Y(n_4153)
);

AOI21x1_ASAP7_75t_SL g4154 ( 
.A1(n_4009),
.A2(n_172),
.B(n_174),
.Y(n_4154)
);

BUFx2_ASAP7_75t_SL g4155 ( 
.A(n_4003),
.Y(n_4155)
);

OAI22xp5_ASAP7_75t_L g4156 ( 
.A1(n_3933),
.A2(n_178),
.B1(n_176),
.B2(n_177),
.Y(n_4156)
);

INVx1_ASAP7_75t_L g4157 ( 
.A(n_3948),
.Y(n_4157)
);

INVx1_ASAP7_75t_L g4158 ( 
.A(n_3876),
.Y(n_4158)
);

OR2x2_ASAP7_75t_L g4159 ( 
.A(n_3935),
.B(n_177),
.Y(n_4159)
);

O2A1O1Ixp5_ASAP7_75t_L g4160 ( 
.A1(n_3950),
.A2(n_181),
.B(n_179),
.C(n_180),
.Y(n_4160)
);

AOI21x1_ASAP7_75t_SL g4161 ( 
.A1(n_3919),
.A2(n_3966),
.B(n_3994),
.Y(n_4161)
);

NAND2xp5_ASAP7_75t_L g4162 ( 
.A(n_3992),
.B(n_183),
.Y(n_4162)
);

HB1xp67_ASAP7_75t_L g4163 ( 
.A(n_4032),
.Y(n_4163)
);

INVx1_ASAP7_75t_L g4164 ( 
.A(n_4018),
.Y(n_4164)
);

NAND2xp5_ASAP7_75t_L g4165 ( 
.A(n_3993),
.B(n_184),
.Y(n_4165)
);

O2A1O1Ixp5_ASAP7_75t_L g4166 ( 
.A1(n_4010),
.A2(n_186),
.B(n_184),
.C(n_185),
.Y(n_4166)
);

INVx2_ASAP7_75t_L g4167 ( 
.A(n_4010),
.Y(n_4167)
);

A2O1A1Ixp33_ASAP7_75t_L g4168 ( 
.A1(n_3984),
.A2(n_188),
.B(n_185),
.C(n_187),
.Y(n_4168)
);

CKINVDCx6p67_ASAP7_75t_R g4169 ( 
.A(n_4029),
.Y(n_4169)
);

OAI22xp5_ASAP7_75t_L g4170 ( 
.A1(n_3937),
.A2(n_3894),
.B1(n_3949),
.B2(n_4021),
.Y(n_4170)
);

AOI21xp5_ASAP7_75t_L g4171 ( 
.A1(n_3918),
.A2(n_1824),
.B(n_1819),
.Y(n_4171)
);

INVx1_ASAP7_75t_L g4172 ( 
.A(n_4026),
.Y(n_4172)
);

INVx1_ASAP7_75t_L g4173 ( 
.A(n_4034),
.Y(n_4173)
);

INVx1_ASAP7_75t_L g4174 ( 
.A(n_4037),
.Y(n_4174)
);

O2A1O1Ixp33_ASAP7_75t_L g4175 ( 
.A1(n_3905),
.A2(n_192),
.B(n_189),
.C(n_190),
.Y(n_4175)
);

AND2x2_ASAP7_75t_L g4176 ( 
.A(n_3925),
.B(n_189),
.Y(n_4176)
);

BUFx6f_ASAP7_75t_SL g4177 ( 
.A(n_4097),
.Y(n_4177)
);

NAND2xp33_ASAP7_75t_R g4178 ( 
.A(n_4120),
.B(n_3957),
.Y(n_4178)
);

AOI222xp33_ASAP7_75t_L g4179 ( 
.A1(n_4067),
.A2(n_3982),
.B1(n_3989),
.B2(n_4028),
.C1(n_4020),
.C2(n_3970),
.Y(n_4179)
);

CKINVDCx8_ASAP7_75t_R g4180 ( 
.A(n_4155),
.Y(n_4180)
);

NAND2xp5_ASAP7_75t_L g4181 ( 
.A(n_4043),
.B(n_4019),
.Y(n_4181)
);

HB1xp67_ASAP7_75t_L g4182 ( 
.A(n_4078),
.Y(n_4182)
);

NAND2xp33_ASAP7_75t_R g4183 ( 
.A(n_4061),
.B(n_4039),
.Y(n_4183)
);

NAND2xp33_ASAP7_75t_R g4184 ( 
.A(n_4159),
.B(n_190),
.Y(n_4184)
);

NOR3xp33_ASAP7_75t_SL g4185 ( 
.A(n_4067),
.B(n_4014),
.C(n_3930),
.Y(n_4185)
);

CKINVDCx5p33_ASAP7_75t_R g4186 ( 
.A(n_4045),
.Y(n_4186)
);

AOI22xp33_ASAP7_75t_L g4187 ( 
.A1(n_4070),
.A2(n_3982),
.B1(n_4036),
.B2(n_4033),
.Y(n_4187)
);

INVx1_ASAP7_75t_L g4188 ( 
.A(n_4143),
.Y(n_4188)
);

INVx1_ASAP7_75t_L g4189 ( 
.A(n_4164),
.Y(n_4189)
);

OA21x2_ASAP7_75t_L g4190 ( 
.A1(n_4073),
.A2(n_3888),
.B(n_3969),
.Y(n_4190)
);

BUFx3_ASAP7_75t_L g4191 ( 
.A(n_4126),
.Y(n_4191)
);

NAND2xp5_ASAP7_75t_L g4192 ( 
.A(n_4158),
.B(n_3894),
.Y(n_4192)
);

INVx1_ASAP7_75t_L g4193 ( 
.A(n_4172),
.Y(n_4193)
);

BUFx4f_ASAP7_75t_SL g4194 ( 
.A(n_4169),
.Y(n_4194)
);

NAND2xp5_ASAP7_75t_L g4195 ( 
.A(n_4044),
.B(n_3939),
.Y(n_4195)
);

OR2x2_ASAP7_75t_L g4196 ( 
.A(n_4041),
.B(n_4047),
.Y(n_4196)
);

AND2x2_ASAP7_75t_L g4197 ( 
.A(n_4085),
.B(n_3921),
.Y(n_4197)
);

BUFx2_ASAP7_75t_L g4198 ( 
.A(n_4093),
.Y(n_4198)
);

OR2x2_ASAP7_75t_L g4199 ( 
.A(n_4092),
.B(n_3890),
.Y(n_4199)
);

INVx1_ASAP7_75t_L g4200 ( 
.A(n_4173),
.Y(n_4200)
);

NOR2xp33_ASAP7_75t_R g4201 ( 
.A(n_4131),
.B(n_4012),
.Y(n_4201)
);

CKINVDCx5p33_ASAP7_75t_R g4202 ( 
.A(n_4049),
.Y(n_4202)
);

CKINVDCx5p33_ASAP7_75t_R g4203 ( 
.A(n_4100),
.Y(n_4203)
);

INVx2_ASAP7_75t_L g4204 ( 
.A(n_4167),
.Y(n_4204)
);

A2O1A1Ixp33_ASAP7_75t_L g4205 ( 
.A1(n_4113),
.A2(n_4136),
.B(n_4168),
.C(n_4160),
.Y(n_4205)
);

INVx1_ASAP7_75t_L g4206 ( 
.A(n_4174),
.Y(n_4206)
);

HB1xp67_ASAP7_75t_L g4207 ( 
.A(n_4056),
.Y(n_4207)
);

AND2x2_ASAP7_75t_L g4208 ( 
.A(n_4111),
.B(n_4027),
.Y(n_4208)
);

BUFx2_ASAP7_75t_L g4209 ( 
.A(n_4124),
.Y(n_4209)
);

OAI22xp5_ASAP7_75t_L g4210 ( 
.A1(n_4170),
.A2(n_3943),
.B1(n_3968),
.B2(n_3944),
.Y(n_4210)
);

INVx2_ASAP7_75t_L g4211 ( 
.A(n_4069),
.Y(n_4211)
);

OR2x6_ASAP7_75t_L g4212 ( 
.A(n_4148),
.B(n_4038),
.Y(n_4212)
);

INVx2_ASAP7_75t_L g4213 ( 
.A(n_4065),
.Y(n_4213)
);

NAND2xp5_ASAP7_75t_L g4214 ( 
.A(n_4050),
.B(n_4086),
.Y(n_4214)
);

INVx1_ASAP7_75t_L g4215 ( 
.A(n_4052),
.Y(n_4215)
);

HB1xp67_ASAP7_75t_L g4216 ( 
.A(n_4074),
.Y(n_4216)
);

AOI21xp33_ASAP7_75t_L g4217 ( 
.A1(n_4123),
.A2(n_3970),
.B(n_3991),
.Y(n_4217)
);

BUFx2_ASAP7_75t_L g4218 ( 
.A(n_4042),
.Y(n_4218)
);

INVx2_ASAP7_75t_L g4219 ( 
.A(n_4054),
.Y(n_4219)
);

AO31x2_ASAP7_75t_L g4220 ( 
.A1(n_4106),
.A2(n_3955),
.A3(n_3981),
.B(n_3932),
.Y(n_4220)
);

INVx1_ASAP7_75t_L g4221 ( 
.A(n_4058),
.Y(n_4221)
);

INVx1_ASAP7_75t_L g4222 ( 
.A(n_4083),
.Y(n_4222)
);

INVx8_ASAP7_75t_L g4223 ( 
.A(n_4135),
.Y(n_4223)
);

INVx2_ASAP7_75t_L g4224 ( 
.A(n_4095),
.Y(n_4224)
);

OAI22xp5_ASAP7_75t_L g4225 ( 
.A1(n_4170),
.A2(n_3963),
.B1(n_3959),
.B2(n_4006),
.Y(n_4225)
);

NAND2xp5_ASAP7_75t_L g4226 ( 
.A(n_4062),
.B(n_3990),
.Y(n_4226)
);

NAND2xp5_ASAP7_75t_L g4227 ( 
.A(n_4066),
.B(n_4027),
.Y(n_4227)
);

AND2x4_ASAP7_75t_L g4228 ( 
.A(n_4063),
.B(n_3955),
.Y(n_4228)
);

OR2x6_ASAP7_75t_L g4229 ( 
.A(n_4087),
.B(n_3981),
.Y(n_4229)
);

BUFx3_ASAP7_75t_L g4230 ( 
.A(n_4053),
.Y(n_4230)
);

AO31x2_ASAP7_75t_L g4231 ( 
.A1(n_4106),
.A2(n_3998),
.A3(n_3895),
.B(n_3956),
.Y(n_4231)
);

AOI22xp33_ASAP7_75t_L g4232 ( 
.A1(n_4080),
.A2(n_3999),
.B1(n_3912),
.B2(n_3917),
.Y(n_4232)
);

A2O1A1Ixp33_ASAP7_75t_L g4233 ( 
.A1(n_4144),
.A2(n_4031),
.B(n_3964),
.C(n_3907),
.Y(n_4233)
);

AND2x2_ASAP7_75t_L g4234 ( 
.A(n_4060),
.B(n_3912),
.Y(n_4234)
);

AND2x4_ASAP7_75t_L g4235 ( 
.A(n_4063),
.B(n_3913),
.Y(n_4235)
);

AND2x2_ASAP7_75t_L g4236 ( 
.A(n_4059),
.B(n_3895),
.Y(n_4236)
);

AND2x2_ASAP7_75t_L g4237 ( 
.A(n_4094),
.B(n_4088),
.Y(n_4237)
);

OR2x2_ASAP7_75t_L g4238 ( 
.A(n_4137),
.B(n_3913),
.Y(n_4238)
);

INVx1_ASAP7_75t_L g4239 ( 
.A(n_4125),
.Y(n_4239)
);

AND2x2_ASAP7_75t_L g4240 ( 
.A(n_4091),
.B(n_3936),
.Y(n_4240)
);

CKINVDCx16_ASAP7_75t_R g4241 ( 
.A(n_4130),
.Y(n_4241)
);

BUFx8_ASAP7_75t_SL g4242 ( 
.A(n_4149),
.Y(n_4242)
);

BUFx3_ASAP7_75t_L g4243 ( 
.A(n_4140),
.Y(n_4243)
);

INVx2_ASAP7_75t_L g4244 ( 
.A(n_4102),
.Y(n_4244)
);

AND2x2_ASAP7_75t_L g4245 ( 
.A(n_4163),
.B(n_3936),
.Y(n_4245)
);

AND2x2_ASAP7_75t_L g4246 ( 
.A(n_4121),
.B(n_3956),
.Y(n_4246)
);

OAI21xp5_ASAP7_75t_L g4247 ( 
.A1(n_4046),
.A2(n_3946),
.B(n_3875),
.Y(n_4247)
);

INVx1_ASAP7_75t_SL g4248 ( 
.A(n_4150),
.Y(n_4248)
);

INVx2_ASAP7_75t_L g4249 ( 
.A(n_4107),
.Y(n_4249)
);

INVx1_ASAP7_75t_L g4250 ( 
.A(n_4145),
.Y(n_4250)
);

NOR2xp33_ASAP7_75t_R g4251 ( 
.A(n_4097),
.B(n_4072),
.Y(n_4251)
);

AND2x2_ASAP7_75t_L g4252 ( 
.A(n_4048),
.B(n_3913),
.Y(n_4252)
);

AND2x2_ASAP7_75t_L g4253 ( 
.A(n_4108),
.B(n_3896),
.Y(n_4253)
);

INVx2_ASAP7_75t_L g4254 ( 
.A(n_4134),
.Y(n_4254)
);

INVx2_ASAP7_75t_L g4255 ( 
.A(n_4146),
.Y(n_4255)
);

OR2x2_ASAP7_75t_L g4256 ( 
.A(n_4109),
.B(n_3954),
.Y(n_4256)
);

NAND2xp33_ASAP7_75t_SL g4257 ( 
.A(n_4138),
.B(n_4090),
.Y(n_4257)
);

AO31x2_ASAP7_75t_L g4258 ( 
.A1(n_4105),
.A2(n_196),
.A3(n_193),
.B(n_195),
.Y(n_4258)
);

BUFx2_ASAP7_75t_L g4259 ( 
.A(n_4117),
.Y(n_4259)
);

OAI21x1_ASAP7_75t_L g4260 ( 
.A1(n_4084),
.A2(n_3983),
.B(n_4030),
.Y(n_4260)
);

AOI22xp33_ASAP7_75t_L g4261 ( 
.A1(n_4080),
.A2(n_3917),
.B1(n_1836),
.B2(n_1859),
.Y(n_4261)
);

NAND3xp33_ASAP7_75t_SL g4262 ( 
.A(n_4075),
.B(n_195),
.C(n_196),
.Y(n_4262)
);

NAND2xp33_ASAP7_75t_R g4263 ( 
.A(n_4176),
.B(n_197),
.Y(n_4263)
);

NAND3xp33_ASAP7_75t_SL g4264 ( 
.A(n_4115),
.B(n_4057),
.C(n_4119),
.Y(n_4264)
);

NOR2xp33_ASAP7_75t_R g4265 ( 
.A(n_4162),
.B(n_199),
.Y(n_4265)
);

INVx3_ASAP7_75t_L g4266 ( 
.A(n_4153),
.Y(n_4266)
);

INVx1_ASAP7_75t_L g4267 ( 
.A(n_4157),
.Y(n_4267)
);

OAI22xp5_ASAP7_75t_L g4268 ( 
.A1(n_4105),
.A2(n_201),
.B1(n_199),
.B2(n_200),
.Y(n_4268)
);

AND2x4_ASAP7_75t_L g4269 ( 
.A(n_4116),
.B(n_200),
.Y(n_4269)
);

INVx2_ASAP7_75t_L g4270 ( 
.A(n_4101),
.Y(n_4270)
);

AND2x2_ASAP7_75t_SL g4271 ( 
.A(n_4141),
.B(n_205),
.Y(n_4271)
);

CKINVDCx5p33_ASAP7_75t_R g4272 ( 
.A(n_4165),
.Y(n_4272)
);

AND2x2_ASAP7_75t_L g4273 ( 
.A(n_4084),
.B(n_205),
.Y(n_4273)
);

AND2x2_ASAP7_75t_L g4274 ( 
.A(n_4142),
.B(n_4151),
.Y(n_4274)
);

OR2x2_ASAP7_75t_SL g4275 ( 
.A(n_4141),
.B(n_206),
.Y(n_4275)
);

NOR3xp33_ASAP7_75t_SL g4276 ( 
.A(n_4112),
.B(n_206),
.C(n_208),
.Y(n_4276)
);

NOR2x1p5_ASAP7_75t_L g4277 ( 
.A(n_4114),
.B(n_209),
.Y(n_4277)
);

NAND3xp33_ASAP7_75t_SL g4278 ( 
.A(n_4115),
.B(n_210),
.C(n_211),
.Y(n_4278)
);

NAND2xp5_ASAP7_75t_L g4279 ( 
.A(n_4152),
.B(n_4128),
.Y(n_4279)
);

AO21x2_ASAP7_75t_L g4280 ( 
.A1(n_4071),
.A2(n_210),
.B(n_211),
.Y(n_4280)
);

INVx2_ASAP7_75t_L g4281 ( 
.A(n_4055),
.Y(n_4281)
);

AOI22xp33_ASAP7_75t_L g4282 ( 
.A1(n_4123),
.A2(n_1898),
.B1(n_1870),
.B2(n_1863),
.Y(n_4282)
);

INVx1_ASAP7_75t_L g4283 ( 
.A(n_4055),
.Y(n_4283)
);

CKINVDCx11_ASAP7_75t_R g4284 ( 
.A(n_4112),
.Y(n_4284)
);

NOR2xp33_ASAP7_75t_R g4285 ( 
.A(n_4129),
.B(n_212),
.Y(n_4285)
);

AOI22xp33_ASAP7_75t_L g4286 ( 
.A1(n_4118),
.A2(n_1898),
.B1(n_1870),
.B2(n_1863),
.Y(n_4286)
);

AO31x2_ASAP7_75t_L g4287 ( 
.A1(n_4076),
.A2(n_213),
.A3(n_214),
.B(n_215),
.Y(n_4287)
);

XNOR2xp5_ASAP7_75t_L g4288 ( 
.A(n_4057),
.B(n_214),
.Y(n_4288)
);

OAI22xp5_ASAP7_75t_L g4289 ( 
.A1(n_4127),
.A2(n_215),
.B1(n_217),
.B2(n_219),
.Y(n_4289)
);

CKINVDCx5p33_ASAP7_75t_R g4290 ( 
.A(n_4103),
.Y(n_4290)
);

INVx1_ASAP7_75t_L g4291 ( 
.A(n_4139),
.Y(n_4291)
);

OR2x2_ASAP7_75t_L g4292 ( 
.A(n_4051),
.B(n_217),
.Y(n_4292)
);

INVx1_ASAP7_75t_L g4293 ( 
.A(n_4122),
.Y(n_4293)
);

AND2x2_ASAP7_75t_L g4294 ( 
.A(n_4122),
.B(n_219),
.Y(n_4294)
);

AOI22xp5_ASAP7_75t_L g4295 ( 
.A1(n_4118),
.A2(n_221),
.B1(n_222),
.B2(n_224),
.Y(n_4295)
);

AND2x2_ASAP7_75t_L g4296 ( 
.A(n_4099),
.B(n_224),
.Y(n_4296)
);

NAND2xp5_ASAP7_75t_L g4297 ( 
.A(n_4077),
.B(n_225),
.Y(n_4297)
);

INVx2_ASAP7_75t_L g4298 ( 
.A(n_4051),
.Y(n_4298)
);

OA21x2_ASAP7_75t_L g4299 ( 
.A1(n_4082),
.A2(n_225),
.B(n_227),
.Y(n_4299)
);

CKINVDCx20_ASAP7_75t_R g4300 ( 
.A(n_4132),
.Y(n_4300)
);

INVx2_ASAP7_75t_L g4301 ( 
.A(n_4166),
.Y(n_4301)
);

NOR2xp33_ASAP7_75t_R g4302 ( 
.A(n_4161),
.B(n_227),
.Y(n_4302)
);

NOR3xp33_ASAP7_75t_SL g4303 ( 
.A(n_4132),
.B(n_228),
.C(n_229),
.Y(n_4303)
);

INVx1_ASAP7_75t_L g4304 ( 
.A(n_4076),
.Y(n_4304)
);

BUFx3_ASAP7_75t_L g4305 ( 
.A(n_4194),
.Y(n_4305)
);

INVx2_ASAP7_75t_L g4306 ( 
.A(n_4281),
.Y(n_4306)
);

AND2x4_ASAP7_75t_L g4307 ( 
.A(n_4231),
.B(n_4229),
.Y(n_4307)
);

INVx2_ASAP7_75t_L g4308 ( 
.A(n_4298),
.Y(n_4308)
);

AND2x4_ASAP7_75t_L g4309 ( 
.A(n_4231),
.B(n_4089),
.Y(n_4309)
);

BUFx2_ASAP7_75t_L g4310 ( 
.A(n_4212),
.Y(n_4310)
);

OR2x2_ASAP7_75t_L g4311 ( 
.A(n_4304),
.B(n_4110),
.Y(n_4311)
);

INVx2_ASAP7_75t_L g4312 ( 
.A(n_4283),
.Y(n_4312)
);

INVx2_ASAP7_75t_L g4313 ( 
.A(n_4259),
.Y(n_4313)
);

OA21x2_ASAP7_75t_L g4314 ( 
.A1(n_4247),
.A2(n_4081),
.B(n_4098),
.Y(n_4314)
);

INVx2_ASAP7_75t_L g4315 ( 
.A(n_4255),
.Y(n_4315)
);

INVx1_ASAP7_75t_L g4316 ( 
.A(n_4215),
.Y(n_4316)
);

INVx1_ASAP7_75t_SL g4317 ( 
.A(n_4201),
.Y(n_4317)
);

BUFx3_ASAP7_75t_L g4318 ( 
.A(n_4242),
.Y(n_4318)
);

INVx3_ASAP7_75t_L g4319 ( 
.A(n_4229),
.Y(n_4319)
);

INVx3_ASAP7_75t_L g4320 ( 
.A(n_4229),
.Y(n_4320)
);

AND2x2_ASAP7_75t_L g4321 ( 
.A(n_4231),
.B(n_4104),
.Y(n_4321)
);

OA21x2_ASAP7_75t_L g4322 ( 
.A1(n_4247),
.A2(n_4127),
.B(n_4171),
.Y(n_4322)
);

INVx2_ASAP7_75t_L g4323 ( 
.A(n_4266),
.Y(n_4323)
);

INVx2_ASAP7_75t_L g4324 ( 
.A(n_4266),
.Y(n_4324)
);

HB1xp67_ASAP7_75t_L g4325 ( 
.A(n_4182),
.Y(n_4325)
);

INVx1_ASAP7_75t_L g4326 ( 
.A(n_4221),
.Y(n_4326)
);

NAND2xp5_ASAP7_75t_L g4327 ( 
.A(n_4274),
.B(n_4104),
.Y(n_4327)
);

OR2x2_ASAP7_75t_L g4328 ( 
.A(n_4192),
.B(n_4110),
.Y(n_4328)
);

AND2x2_ASAP7_75t_L g4329 ( 
.A(n_4220),
.B(n_4133),
.Y(n_4329)
);

NOR2xp33_ASAP7_75t_L g4330 ( 
.A(n_4177),
.B(n_4147),
.Y(n_4330)
);

INVx1_ASAP7_75t_L g4331 ( 
.A(n_4222),
.Y(n_4331)
);

INVx2_ASAP7_75t_L g4332 ( 
.A(n_4292),
.Y(n_4332)
);

BUFx2_ASAP7_75t_L g4333 ( 
.A(n_4212),
.Y(n_4333)
);

INVx2_ASAP7_75t_L g4334 ( 
.A(n_4280),
.Y(n_4334)
);

INVx2_ASAP7_75t_L g4335 ( 
.A(n_4280),
.Y(n_4335)
);

HB1xp67_ASAP7_75t_L g4336 ( 
.A(n_4198),
.Y(n_4336)
);

OAI21x1_ASAP7_75t_L g4337 ( 
.A1(n_4192),
.A2(n_4064),
.B(n_4079),
.Y(n_4337)
);

OAI21xp5_ASAP7_75t_L g4338 ( 
.A1(n_4264),
.A2(n_4156),
.B(n_4147),
.Y(n_4338)
);

INVx2_ASAP7_75t_L g4339 ( 
.A(n_4224),
.Y(n_4339)
);

OA21x2_ASAP7_75t_L g4340 ( 
.A1(n_4185),
.A2(n_4156),
.B(n_4068),
.Y(n_4340)
);

INVx2_ASAP7_75t_L g4341 ( 
.A(n_4244),
.Y(n_4341)
);

INVx2_ASAP7_75t_L g4342 ( 
.A(n_4249),
.Y(n_4342)
);

INVx2_ASAP7_75t_L g4343 ( 
.A(n_4254),
.Y(n_4343)
);

INVx3_ASAP7_75t_L g4344 ( 
.A(n_4220),
.Y(n_4344)
);

INVx2_ASAP7_75t_L g4345 ( 
.A(n_4204),
.Y(n_4345)
);

A2O1A1Ixp33_ASAP7_75t_L g4346 ( 
.A1(n_4205),
.A2(n_4175),
.B(n_4096),
.C(n_4154),
.Y(n_4346)
);

INVx1_ASAP7_75t_L g4347 ( 
.A(n_4239),
.Y(n_4347)
);

OR2x2_ASAP7_75t_L g4348 ( 
.A(n_4216),
.B(n_228),
.Y(n_4348)
);

AOI22xp33_ASAP7_75t_L g4349 ( 
.A1(n_4284),
.A2(n_229),
.B1(n_231),
.B2(n_233),
.Y(n_4349)
);

AO21x2_ASAP7_75t_L g4350 ( 
.A1(n_4268),
.A2(n_231),
.B(n_234),
.Y(n_4350)
);

OA21x2_ASAP7_75t_L g4351 ( 
.A1(n_4260),
.A2(n_234),
.B(n_235),
.Y(n_4351)
);

INVx2_ASAP7_75t_L g4352 ( 
.A(n_4250),
.Y(n_4352)
);

AOI211xp5_ASAP7_75t_L g4353 ( 
.A1(n_4268),
.A2(n_235),
.B(n_236),
.C(n_237),
.Y(n_4353)
);

NAND2xp5_ASAP7_75t_L g4354 ( 
.A(n_4291),
.B(n_237),
.Y(n_4354)
);

AO21x2_ASAP7_75t_L g4355 ( 
.A1(n_4297),
.A2(n_238),
.B(n_240),
.Y(n_4355)
);

HB1xp67_ASAP7_75t_L g4356 ( 
.A(n_4209),
.Y(n_4356)
);

OR2x6_ASAP7_75t_L g4357 ( 
.A(n_4212),
.B(n_241),
.Y(n_4357)
);

AOI21xp33_ASAP7_75t_L g4358 ( 
.A1(n_4301),
.A2(n_242),
.B(n_244),
.Y(n_4358)
);

HB1xp67_ASAP7_75t_L g4359 ( 
.A(n_4218),
.Y(n_4359)
);

OR2x2_ASAP7_75t_L g4360 ( 
.A(n_4207),
.B(n_244),
.Y(n_4360)
);

OA21x2_ASAP7_75t_L g4361 ( 
.A1(n_4261),
.A2(n_245),
.B(n_246),
.Y(n_4361)
);

BUFx3_ASAP7_75t_L g4362 ( 
.A(n_4180),
.Y(n_4362)
);

OAI22xp5_ASAP7_75t_L g4363 ( 
.A1(n_4232),
.A2(n_245),
.B1(n_246),
.B2(n_247),
.Y(n_4363)
);

AND2x2_ASAP7_75t_L g4364 ( 
.A(n_4220),
.B(n_247),
.Y(n_4364)
);

INVx2_ASAP7_75t_L g4365 ( 
.A(n_4267),
.Y(n_4365)
);

AND2x2_ASAP7_75t_L g4366 ( 
.A(n_4253),
.B(n_248),
.Y(n_4366)
);

AND2x2_ASAP7_75t_L g4367 ( 
.A(n_4228),
.B(n_250),
.Y(n_4367)
);

OAI221xp5_ASAP7_75t_L g4368 ( 
.A1(n_4295),
.A2(n_250),
.B1(n_251),
.B2(n_252),
.C(n_255),
.Y(n_4368)
);

AND2x2_ASAP7_75t_L g4369 ( 
.A(n_4228),
.B(n_252),
.Y(n_4369)
);

INVx1_ASAP7_75t_L g4370 ( 
.A(n_4189),
.Y(n_4370)
);

BUFx2_ASAP7_75t_L g4371 ( 
.A(n_4251),
.Y(n_4371)
);

INVx1_ASAP7_75t_L g4372 ( 
.A(n_4193),
.Y(n_4372)
);

INVx1_ASAP7_75t_L g4373 ( 
.A(n_4200),
.Y(n_4373)
);

AND2x2_ASAP7_75t_L g4374 ( 
.A(n_4237),
.B(n_256),
.Y(n_4374)
);

INVx2_ASAP7_75t_L g4375 ( 
.A(n_4206),
.Y(n_4375)
);

AND2x2_ASAP7_75t_L g4376 ( 
.A(n_4270),
.B(n_256),
.Y(n_4376)
);

INVx1_ASAP7_75t_L g4377 ( 
.A(n_4188),
.Y(n_4377)
);

INVx1_ASAP7_75t_L g4378 ( 
.A(n_4213),
.Y(n_4378)
);

AOI21xp5_ASAP7_75t_SL g4379 ( 
.A1(n_4278),
.A2(n_4299),
.B(n_4262),
.Y(n_4379)
);

OR2x2_ASAP7_75t_L g4380 ( 
.A(n_4196),
.B(n_257),
.Y(n_4380)
);

OR2x2_ASAP7_75t_L g4381 ( 
.A(n_4214),
.B(n_4287),
.Y(n_4381)
);

INVx3_ASAP7_75t_L g4382 ( 
.A(n_4235),
.Y(n_4382)
);

AND2x4_ASAP7_75t_L g4383 ( 
.A(n_4287),
.B(n_4258),
.Y(n_4383)
);

OA21x2_ASAP7_75t_L g4384 ( 
.A1(n_4227),
.A2(n_4276),
.B(n_4217),
.Y(n_4384)
);

INVx2_ASAP7_75t_L g4385 ( 
.A(n_4275),
.Y(n_4385)
);

AND2x2_ASAP7_75t_L g4386 ( 
.A(n_4235),
.B(n_257),
.Y(n_4386)
);

INVx1_ASAP7_75t_L g4387 ( 
.A(n_4271),
.Y(n_4387)
);

AOI22xp33_ASAP7_75t_SL g4388 ( 
.A1(n_4302),
.A2(n_258),
.B1(n_260),
.B2(n_261),
.Y(n_4388)
);

HB1xp67_ASAP7_75t_L g4389 ( 
.A(n_4287),
.Y(n_4389)
);

INVx1_ASAP7_75t_L g4390 ( 
.A(n_4258),
.Y(n_4390)
);

INVx2_ASAP7_75t_L g4391 ( 
.A(n_4238),
.Y(n_4391)
);

AOI221xp5_ASAP7_75t_L g4392 ( 
.A1(n_4288),
.A2(n_261),
.B1(n_262),
.B2(n_263),
.C(n_264),
.Y(n_4392)
);

NOR2xp33_ASAP7_75t_L g4393 ( 
.A(n_4177),
.B(n_262),
.Y(n_4393)
);

AND2x2_ASAP7_75t_L g4394 ( 
.A(n_4211),
.B(n_265),
.Y(n_4394)
);

AND2x2_ASAP7_75t_L g4395 ( 
.A(n_4219),
.B(n_267),
.Y(n_4395)
);

AND2x2_ASAP7_75t_L g4396 ( 
.A(n_4245),
.B(n_4248),
.Y(n_4396)
);

NOR2x1_ASAP7_75t_R g4397 ( 
.A(n_4290),
.B(n_267),
.Y(n_4397)
);

INVx1_ASAP7_75t_L g4398 ( 
.A(n_4258),
.Y(n_4398)
);

INVx2_ASAP7_75t_L g4399 ( 
.A(n_4269),
.Y(n_4399)
);

INVx3_ASAP7_75t_L g4400 ( 
.A(n_4241),
.Y(n_4400)
);

OA21x2_ASAP7_75t_L g4401 ( 
.A1(n_4217),
.A2(n_271),
.B(n_272),
.Y(n_4401)
);

INVx4_ASAP7_75t_L g4402 ( 
.A(n_4296),
.Y(n_4402)
);

AND2x2_ASAP7_75t_L g4403 ( 
.A(n_4248),
.B(n_273),
.Y(n_4403)
);

OR2x2_ASAP7_75t_L g4404 ( 
.A(n_4279),
.B(n_273),
.Y(n_4404)
);

INVx1_ASAP7_75t_L g4405 ( 
.A(n_4299),
.Y(n_4405)
);

HB1xp67_ASAP7_75t_L g4406 ( 
.A(n_4336),
.Y(n_4406)
);

NOR2x1_ASAP7_75t_L g4407 ( 
.A(n_4364),
.B(n_4277),
.Y(n_4407)
);

INVx2_ASAP7_75t_L g4408 ( 
.A(n_4312),
.Y(n_4408)
);

INVx2_ASAP7_75t_L g4409 ( 
.A(n_4312),
.Y(n_4409)
);

AND2x4_ASAP7_75t_L g4410 ( 
.A(n_4400),
.B(n_4197),
.Y(n_4410)
);

INVx1_ASAP7_75t_L g4411 ( 
.A(n_4352),
.Y(n_4411)
);

INVx1_ASAP7_75t_L g4412 ( 
.A(n_4352),
.Y(n_4412)
);

INVx3_ASAP7_75t_L g4413 ( 
.A(n_4400),
.Y(n_4413)
);

INVx1_ASAP7_75t_L g4414 ( 
.A(n_4365),
.Y(n_4414)
);

AND2x2_ASAP7_75t_L g4415 ( 
.A(n_4400),
.B(n_4199),
.Y(n_4415)
);

INVx1_ASAP7_75t_L g4416 ( 
.A(n_4365),
.Y(n_4416)
);

BUFx3_ASAP7_75t_L g4417 ( 
.A(n_4318),
.Y(n_4417)
);

INVx2_ASAP7_75t_L g4418 ( 
.A(n_4308),
.Y(n_4418)
);

NAND2xp5_ASAP7_75t_L g4419 ( 
.A(n_4385),
.B(n_4269),
.Y(n_4419)
);

INVx1_ASAP7_75t_L g4420 ( 
.A(n_4375),
.Y(n_4420)
);

INVx1_ASAP7_75t_L g4421 ( 
.A(n_4375),
.Y(n_4421)
);

AND2x2_ASAP7_75t_L g4422 ( 
.A(n_4310),
.B(n_4236),
.Y(n_4422)
);

INVx2_ASAP7_75t_L g4423 ( 
.A(n_4308),
.Y(n_4423)
);

AND2x4_ASAP7_75t_L g4424 ( 
.A(n_4382),
.B(n_4208),
.Y(n_4424)
);

NAND2xp5_ASAP7_75t_L g4425 ( 
.A(n_4385),
.B(n_4273),
.Y(n_4425)
);

INVx1_ASAP7_75t_L g4426 ( 
.A(n_4316),
.Y(n_4426)
);

INVx2_ASAP7_75t_L g4427 ( 
.A(n_4306),
.Y(n_4427)
);

AND2x2_ASAP7_75t_L g4428 ( 
.A(n_4310),
.B(n_4333),
.Y(n_4428)
);

AND2x2_ASAP7_75t_L g4429 ( 
.A(n_4333),
.B(n_4240),
.Y(n_4429)
);

INVx1_ASAP7_75t_SL g4430 ( 
.A(n_4371),
.Y(n_4430)
);

AND2x2_ASAP7_75t_L g4431 ( 
.A(n_4382),
.B(n_4234),
.Y(n_4431)
);

INVx2_ASAP7_75t_L g4432 ( 
.A(n_4306),
.Y(n_4432)
);

AND2x4_ASAP7_75t_L g4433 ( 
.A(n_4382),
.B(n_4243),
.Y(n_4433)
);

INVx1_ASAP7_75t_SL g4434 ( 
.A(n_4371),
.Y(n_4434)
);

INVx1_ASAP7_75t_L g4435 ( 
.A(n_4316),
.Y(n_4435)
);

NAND2xp5_ASAP7_75t_L g4436 ( 
.A(n_4387),
.B(n_4300),
.Y(n_4436)
);

INVx1_ASAP7_75t_L g4437 ( 
.A(n_4326),
.Y(n_4437)
);

INVx2_ASAP7_75t_L g4438 ( 
.A(n_4396),
.Y(n_4438)
);

AND2x2_ASAP7_75t_L g4439 ( 
.A(n_4321),
.B(n_4252),
.Y(n_4439)
);

HB1xp67_ASAP7_75t_L g4440 ( 
.A(n_4356),
.Y(n_4440)
);

AND2x4_ASAP7_75t_L g4441 ( 
.A(n_4307),
.B(n_4293),
.Y(n_4441)
);

NOR2x1_ASAP7_75t_L g4442 ( 
.A(n_4364),
.B(n_4230),
.Y(n_4442)
);

OR2x2_ASAP7_75t_L g4443 ( 
.A(n_4332),
.B(n_4256),
.Y(n_4443)
);

INVx1_ASAP7_75t_L g4444 ( 
.A(n_4326),
.Y(n_4444)
);

AND2x2_ASAP7_75t_L g4445 ( 
.A(n_4321),
.B(n_4246),
.Y(n_4445)
);

INVx2_ASAP7_75t_L g4446 ( 
.A(n_4396),
.Y(n_4446)
);

INVx1_ASAP7_75t_L g4447 ( 
.A(n_4331),
.Y(n_4447)
);

INVx2_ASAP7_75t_L g4448 ( 
.A(n_4399),
.Y(n_4448)
);

NAND2xp5_ASAP7_75t_L g4449 ( 
.A(n_4387),
.B(n_4179),
.Y(n_4449)
);

INVx1_ASAP7_75t_L g4450 ( 
.A(n_4331),
.Y(n_4450)
);

INVx2_ASAP7_75t_L g4451 ( 
.A(n_4399),
.Y(n_4451)
);

INVx2_ASAP7_75t_L g4452 ( 
.A(n_4359),
.Y(n_4452)
);

AND2x2_ASAP7_75t_L g4453 ( 
.A(n_4307),
.B(n_4187),
.Y(n_4453)
);

NAND2xp5_ASAP7_75t_SL g4454 ( 
.A(n_4402),
.B(n_4179),
.Y(n_4454)
);

INVx1_ASAP7_75t_L g4455 ( 
.A(n_4347),
.Y(n_4455)
);

INVx1_ASAP7_75t_L g4456 ( 
.A(n_4347),
.Y(n_4456)
);

AND2x4_ASAP7_75t_L g4457 ( 
.A(n_4307),
.B(n_4191),
.Y(n_4457)
);

HB1xp67_ASAP7_75t_L g4458 ( 
.A(n_4325),
.Y(n_4458)
);

INVx4_ASAP7_75t_R g4459 ( 
.A(n_4318),
.Y(n_4459)
);

AND2x2_ASAP7_75t_L g4460 ( 
.A(n_4329),
.B(n_4319),
.Y(n_4460)
);

AND2x2_ASAP7_75t_L g4461 ( 
.A(n_4329),
.B(n_4190),
.Y(n_4461)
);

AND2x2_ASAP7_75t_L g4462 ( 
.A(n_4319),
.B(n_4190),
.Y(n_4462)
);

AND2x2_ASAP7_75t_L g4463 ( 
.A(n_4319),
.B(n_4181),
.Y(n_4463)
);

AND2x2_ASAP7_75t_L g4464 ( 
.A(n_4320),
.B(n_4195),
.Y(n_4464)
);

OR2x2_ASAP7_75t_L g4465 ( 
.A(n_4332),
.B(n_4226),
.Y(n_4465)
);

INVx2_ASAP7_75t_L g4466 ( 
.A(n_4323),
.Y(n_4466)
);

INVx1_ASAP7_75t_L g4467 ( 
.A(n_4370),
.Y(n_4467)
);

AOI22xp5_ASAP7_75t_L g4468 ( 
.A1(n_4314),
.A2(n_4295),
.B1(n_4184),
.B2(n_4257),
.Y(n_4468)
);

NOR2xp67_ASAP7_75t_L g4469 ( 
.A(n_4320),
.B(n_4202),
.Y(n_4469)
);

INVx1_ASAP7_75t_L g4470 ( 
.A(n_4370),
.Y(n_4470)
);

AND2x2_ASAP7_75t_L g4471 ( 
.A(n_4320),
.B(n_4314),
.Y(n_4471)
);

OR2x2_ASAP7_75t_L g4472 ( 
.A(n_4390),
.B(n_4223),
.Y(n_4472)
);

AOI221xp5_ASAP7_75t_L g4473 ( 
.A1(n_4454),
.A2(n_4338),
.B1(n_4346),
.B2(n_4379),
.C(n_4383),
.Y(n_4473)
);

AOI22xp33_ASAP7_75t_L g4474 ( 
.A1(n_4449),
.A2(n_4314),
.B1(n_4322),
.B2(n_4384),
.Y(n_4474)
);

OA21x2_ASAP7_75t_L g4475 ( 
.A1(n_4468),
.A2(n_4335),
.B(n_4334),
.Y(n_4475)
);

AO21x2_ASAP7_75t_L g4476 ( 
.A1(n_4461),
.A2(n_4335),
.B(n_4334),
.Y(n_4476)
);

OAI22xp5_ASAP7_75t_L g4477 ( 
.A1(n_4442),
.A2(n_4314),
.B1(n_4328),
.B2(n_4388),
.Y(n_4477)
);

AOI21xp33_ASAP7_75t_L g4478 ( 
.A1(n_4442),
.A2(n_4322),
.B(n_4328),
.Y(n_4478)
);

NAND2xp5_ASAP7_75t_L g4479 ( 
.A(n_4430),
.B(n_4434),
.Y(n_4479)
);

NOR5xp2_ASAP7_75t_SL g4480 ( 
.A(n_4459),
.B(n_4263),
.C(n_4392),
.D(n_4358),
.E(n_4363),
.Y(n_4480)
);

INVx1_ASAP7_75t_SL g4481 ( 
.A(n_4417),
.Y(n_4481)
);

INVx3_ASAP7_75t_L g4482 ( 
.A(n_4417),
.Y(n_4482)
);

AND2x2_ASAP7_75t_L g4483 ( 
.A(n_4422),
.B(n_4402),
.Y(n_4483)
);

INVx1_ASAP7_75t_L g4484 ( 
.A(n_4426),
.Y(n_4484)
);

AND2x2_ASAP7_75t_L g4485 ( 
.A(n_4422),
.B(n_4402),
.Y(n_4485)
);

AOI22xp33_ASAP7_75t_L g4486 ( 
.A1(n_4407),
.A2(n_4322),
.B1(n_4384),
.B2(n_4383),
.Y(n_4486)
);

NAND4xp25_ASAP7_75t_L g4487 ( 
.A(n_4407),
.B(n_4349),
.C(n_4353),
.D(n_4330),
.Y(n_4487)
);

INVx1_ASAP7_75t_L g4488 ( 
.A(n_4426),
.Y(n_4488)
);

NAND3xp33_ASAP7_75t_L g4489 ( 
.A(n_4458),
.B(n_4379),
.C(n_4322),
.Y(n_4489)
);

AOI22xp33_ASAP7_75t_L g4490 ( 
.A1(n_4436),
.A2(n_4384),
.B1(n_4383),
.B2(n_4368),
.Y(n_4490)
);

INVx2_ASAP7_75t_SL g4491 ( 
.A(n_4459),
.Y(n_4491)
);

AOI221xp5_ASAP7_75t_L g4492 ( 
.A1(n_4406),
.A2(n_4383),
.B1(n_4440),
.B2(n_4389),
.C(n_4428),
.Y(n_4492)
);

AND2x4_ASAP7_75t_L g4493 ( 
.A(n_4469),
.B(n_4313),
.Y(n_4493)
);

INVx5_ASAP7_75t_L g4494 ( 
.A(n_4413),
.Y(n_4494)
);

AOI22xp33_ASAP7_75t_L g4495 ( 
.A1(n_4425),
.A2(n_4384),
.B1(n_4327),
.B2(n_4311),
.Y(n_4495)
);

AOI22xp33_ASAP7_75t_L g4496 ( 
.A1(n_4410),
.A2(n_4311),
.B1(n_4355),
.B2(n_4350),
.Y(n_4496)
);

AND2x4_ASAP7_75t_L g4497 ( 
.A(n_4413),
.B(n_4313),
.Y(n_4497)
);

OAI211xp5_ASAP7_75t_L g4498 ( 
.A1(n_4461),
.A2(n_4390),
.B(n_4398),
.C(n_4303),
.Y(n_4498)
);

INVx1_ASAP7_75t_L g4499 ( 
.A(n_4435),
.Y(n_4499)
);

INVx2_ASAP7_75t_L g4500 ( 
.A(n_4413),
.Y(n_4500)
);

OAI211xp5_ASAP7_75t_SL g4501 ( 
.A1(n_4419),
.A2(n_4317),
.B(n_4405),
.C(n_4354),
.Y(n_4501)
);

NOR2xp33_ASAP7_75t_L g4502 ( 
.A(n_4410),
.B(n_4305),
.Y(n_4502)
);

AOI222xp33_ASAP7_75t_L g4503 ( 
.A1(n_4428),
.A2(n_4397),
.B1(n_4398),
.B2(n_4405),
.C1(n_4393),
.C2(n_4366),
.Y(n_4503)
);

INVx1_ASAP7_75t_L g4504 ( 
.A(n_4435),
.Y(n_4504)
);

INVx2_ASAP7_75t_L g4505 ( 
.A(n_4429),
.Y(n_4505)
);

INVx2_ASAP7_75t_L g4506 ( 
.A(n_4429),
.Y(n_4506)
);

AO21x2_ASAP7_75t_L g4507 ( 
.A1(n_4471),
.A2(n_4403),
.B(n_4366),
.Y(n_4507)
);

OAI31xp33_ASAP7_75t_L g4508 ( 
.A1(n_4453),
.A2(n_4381),
.A3(n_4309),
.B(n_4210),
.Y(n_4508)
);

OAI21x1_ASAP7_75t_L g4509 ( 
.A1(n_4460),
.A2(n_4344),
.B(n_4337),
.Y(n_4509)
);

INVx2_ASAP7_75t_L g4510 ( 
.A(n_4433),
.Y(n_4510)
);

INVx2_ASAP7_75t_L g4511 ( 
.A(n_4433),
.Y(n_4511)
);

OAI21xp5_ASAP7_75t_L g4512 ( 
.A1(n_4453),
.A2(n_4337),
.B(n_4340),
.Y(n_4512)
);

AOI21xp5_ASAP7_75t_L g4513 ( 
.A1(n_4410),
.A2(n_4397),
.B(n_4357),
.Y(n_4513)
);

INVx1_ASAP7_75t_L g4514 ( 
.A(n_4505),
.Y(n_4514)
);

AND2x2_ASAP7_75t_L g4515 ( 
.A(n_4482),
.B(n_4445),
.Y(n_4515)
);

NAND2xp5_ASAP7_75t_L g4516 ( 
.A(n_4481),
.B(n_4452),
.Y(n_4516)
);

AOI33xp33_ASAP7_75t_L g4517 ( 
.A1(n_4473),
.A2(n_4452),
.A3(n_4438),
.B1(n_4446),
.B2(n_4448),
.B3(n_4451),
.Y(n_4517)
);

AND2x4_ASAP7_75t_L g4518 ( 
.A(n_4494),
.B(n_4457),
.Y(n_4518)
);

AND2x2_ASAP7_75t_L g4519 ( 
.A(n_4482),
.B(n_4445),
.Y(n_4519)
);

INVx1_ASAP7_75t_L g4520 ( 
.A(n_4505),
.Y(n_4520)
);

AND2x2_ASAP7_75t_L g4521 ( 
.A(n_4491),
.B(n_4433),
.Y(n_4521)
);

AND2x2_ASAP7_75t_L g4522 ( 
.A(n_4483),
.B(n_4431),
.Y(n_4522)
);

AND2x2_ASAP7_75t_SL g4523 ( 
.A(n_4486),
.B(n_4474),
.Y(n_4523)
);

AND2x2_ASAP7_75t_L g4524 ( 
.A(n_4485),
.B(n_4431),
.Y(n_4524)
);

OR2x2_ASAP7_75t_L g4525 ( 
.A(n_4507),
.B(n_4438),
.Y(n_4525)
);

INVx2_ASAP7_75t_L g4526 ( 
.A(n_4494),
.Y(n_4526)
);

INVx2_ASAP7_75t_SL g4527 ( 
.A(n_4494),
.Y(n_4527)
);

NAND2xp5_ASAP7_75t_L g4528 ( 
.A(n_4506),
.B(n_4448),
.Y(n_4528)
);

AND2x4_ASAP7_75t_L g4529 ( 
.A(n_4494),
.B(n_4457),
.Y(n_4529)
);

BUFx2_ASAP7_75t_L g4530 ( 
.A(n_4493),
.Y(n_4530)
);

INVx1_ASAP7_75t_L g4531 ( 
.A(n_4506),
.Y(n_4531)
);

INVx1_ASAP7_75t_L g4532 ( 
.A(n_4484),
.Y(n_4532)
);

AND2x2_ASAP7_75t_L g4533 ( 
.A(n_4493),
.B(n_4457),
.Y(n_4533)
);

INVx2_ASAP7_75t_L g4534 ( 
.A(n_4476),
.Y(n_4534)
);

INVx1_ASAP7_75t_L g4535 ( 
.A(n_4488),
.Y(n_4535)
);

INVx2_ASAP7_75t_L g4536 ( 
.A(n_4476),
.Y(n_4536)
);

HB1xp67_ASAP7_75t_L g4537 ( 
.A(n_4507),
.Y(n_4537)
);

BUFx2_ASAP7_75t_L g4538 ( 
.A(n_4493),
.Y(n_4538)
);

INVx2_ASAP7_75t_L g4539 ( 
.A(n_4497),
.Y(n_4539)
);

AND2x4_ASAP7_75t_L g4540 ( 
.A(n_4497),
.B(n_4446),
.Y(n_4540)
);

INVxp67_ASAP7_75t_L g4541 ( 
.A(n_4530),
.Y(n_4541)
);

INVx1_ASAP7_75t_L g4542 ( 
.A(n_4537),
.Y(n_4542)
);

AND2x2_ASAP7_75t_SL g4543 ( 
.A(n_4523),
.B(n_4486),
.Y(n_4543)
);

INVx1_ASAP7_75t_L g4544 ( 
.A(n_4530),
.Y(n_4544)
);

NOR2xp33_ASAP7_75t_L g4545 ( 
.A(n_4523),
.B(n_4502),
.Y(n_4545)
);

AND2x2_ASAP7_75t_L g4546 ( 
.A(n_4521),
.B(n_4502),
.Y(n_4546)
);

HB1xp67_ASAP7_75t_L g4547 ( 
.A(n_4538),
.Y(n_4547)
);

INVx1_ASAP7_75t_L g4548 ( 
.A(n_4538),
.Y(n_4548)
);

INVx1_ASAP7_75t_L g4549 ( 
.A(n_4525),
.Y(n_4549)
);

NAND2xp5_ASAP7_75t_L g4550 ( 
.A(n_4515),
.B(n_4519),
.Y(n_4550)
);

NAND2xp5_ASAP7_75t_L g4551 ( 
.A(n_4515),
.B(n_4503),
.Y(n_4551)
);

AND2x2_ASAP7_75t_L g4552 ( 
.A(n_4521),
.B(n_4510),
.Y(n_4552)
);

HB1xp67_ASAP7_75t_L g4553 ( 
.A(n_4525),
.Y(n_4553)
);

AND2x2_ASAP7_75t_L g4554 ( 
.A(n_4519),
.B(n_4510),
.Y(n_4554)
);

INVx1_ASAP7_75t_L g4555 ( 
.A(n_4514),
.Y(n_4555)
);

INVxp67_ASAP7_75t_SL g4556 ( 
.A(n_4533),
.Y(n_4556)
);

INVxp67_ASAP7_75t_L g4557 ( 
.A(n_4533),
.Y(n_4557)
);

INVxp67_ASAP7_75t_L g4558 ( 
.A(n_4518),
.Y(n_4558)
);

AOI22xp5_ASAP7_75t_L g4559 ( 
.A1(n_4543),
.A2(n_4523),
.B1(n_4477),
.B2(n_4490),
.Y(n_4559)
);

OR2x2_ASAP7_75t_L g4560 ( 
.A(n_4550),
.B(n_4516),
.Y(n_4560)
);

NAND2xp5_ASAP7_75t_L g4561 ( 
.A(n_4556),
.B(n_4522),
.Y(n_4561)
);

OR2x2_ASAP7_75t_L g4562 ( 
.A(n_4551),
.B(n_4479),
.Y(n_4562)
);

NAND2xp5_ASAP7_75t_L g4563 ( 
.A(n_4552),
.B(n_4522),
.Y(n_4563)
);

OR2x2_ASAP7_75t_L g4564 ( 
.A(n_4557),
.B(n_4451),
.Y(n_4564)
);

NAND2xp5_ASAP7_75t_L g4565 ( 
.A(n_4552),
.B(n_4524),
.Y(n_4565)
);

INVx1_ASAP7_75t_L g4566 ( 
.A(n_4547),
.Y(n_4566)
);

AND2x2_ASAP7_75t_L g4567 ( 
.A(n_4546),
.B(n_4524),
.Y(n_4567)
);

AND2x2_ASAP7_75t_L g4568 ( 
.A(n_4546),
.B(n_4554),
.Y(n_4568)
);

NAND4xp25_ASAP7_75t_L g4569 ( 
.A(n_4545),
.B(n_4474),
.C(n_4508),
.D(n_4495),
.Y(n_4569)
);

INVx2_ASAP7_75t_L g4570 ( 
.A(n_4554),
.Y(n_4570)
);

INVx1_ASAP7_75t_L g4571 ( 
.A(n_4544),
.Y(n_4571)
);

AND2x2_ASAP7_75t_L g4572 ( 
.A(n_4545),
.B(n_4511),
.Y(n_4572)
);

NAND2xp5_ASAP7_75t_L g4573 ( 
.A(n_4543),
.B(n_4511),
.Y(n_4573)
);

NAND2xp5_ASAP7_75t_L g4574 ( 
.A(n_4558),
.B(n_4517),
.Y(n_4574)
);

OR2x2_ASAP7_75t_L g4575 ( 
.A(n_4548),
.B(n_4541),
.Y(n_4575)
);

AND2x2_ASAP7_75t_L g4576 ( 
.A(n_4553),
.B(n_4513),
.Y(n_4576)
);

INVx1_ASAP7_75t_SL g4577 ( 
.A(n_4568),
.Y(n_4577)
);

OAI22xp33_ASAP7_75t_L g4578 ( 
.A1(n_4559),
.A2(n_4489),
.B1(n_4512),
.B2(n_4487),
.Y(n_4578)
);

INVx1_ASAP7_75t_L g4579 ( 
.A(n_4561),
.Y(n_4579)
);

NAND2xp5_ASAP7_75t_SL g4580 ( 
.A(n_4559),
.B(n_4478),
.Y(n_4580)
);

AOI21xp33_ASAP7_75t_SL g4581 ( 
.A1(n_4573),
.A2(n_4475),
.B(n_4490),
.Y(n_4581)
);

HB1xp67_ASAP7_75t_L g4582 ( 
.A(n_4567),
.Y(n_4582)
);

AND2x2_ASAP7_75t_L g4583 ( 
.A(n_4572),
.B(n_4305),
.Y(n_4583)
);

NOR2xp33_ASAP7_75t_L g4584 ( 
.A(n_4569),
.B(n_4562),
.Y(n_4584)
);

INVx1_ASAP7_75t_L g4585 ( 
.A(n_4570),
.Y(n_4585)
);

NOR2xp67_ASAP7_75t_SL g4586 ( 
.A(n_4575),
.B(n_4362),
.Y(n_4586)
);

OR2x2_ASAP7_75t_L g4587 ( 
.A(n_4563),
.B(n_4528),
.Y(n_4587)
);

AOI21xp33_ASAP7_75t_SL g4588 ( 
.A1(n_4565),
.A2(n_4475),
.B(n_4527),
.Y(n_4588)
);

INVxp67_ASAP7_75t_L g4589 ( 
.A(n_4582),
.Y(n_4589)
);

INVx1_ASAP7_75t_L g4590 ( 
.A(n_4577),
.Y(n_4590)
);

BUFx4f_ASAP7_75t_SL g4591 ( 
.A(n_4583),
.Y(n_4591)
);

INVx1_ASAP7_75t_SL g4592 ( 
.A(n_4577),
.Y(n_4592)
);

INVx1_ASAP7_75t_SL g4593 ( 
.A(n_4587),
.Y(n_4593)
);

NAND2xp5_ASAP7_75t_L g4594 ( 
.A(n_4581),
.B(n_4566),
.Y(n_4594)
);

INVx1_ASAP7_75t_L g4595 ( 
.A(n_4585),
.Y(n_4595)
);

INVx2_ASAP7_75t_L g4596 ( 
.A(n_4579),
.Y(n_4596)
);

INVx1_ASAP7_75t_L g4597 ( 
.A(n_4586),
.Y(n_4597)
);

O2A1O1Ixp33_ASAP7_75t_L g4598 ( 
.A1(n_4594),
.A2(n_4580),
.B(n_4578),
.C(n_4588),
.Y(n_4598)
);

AOI22xp5_ASAP7_75t_L g4599 ( 
.A1(n_4592),
.A2(n_4569),
.B1(n_4584),
.B2(n_4495),
.Y(n_4599)
);

INVx1_ASAP7_75t_L g4600 ( 
.A(n_4590),
.Y(n_4600)
);

AND2x4_ASAP7_75t_L g4601 ( 
.A(n_4589),
.B(n_4571),
.Y(n_4601)
);

INVx1_ASAP7_75t_L g4602 ( 
.A(n_4594),
.Y(n_4602)
);

A2O1A1O1Ixp25_ASAP7_75t_L g4603 ( 
.A1(n_4597),
.A2(n_4574),
.B(n_4498),
.C(n_4542),
.D(n_4549),
.Y(n_4603)
);

INVx1_ASAP7_75t_L g4604 ( 
.A(n_4595),
.Y(n_4604)
);

AOI222xp33_ASAP7_75t_L g4605 ( 
.A1(n_4591),
.A2(n_4492),
.B1(n_4576),
.B2(n_4534),
.C1(n_4536),
.C2(n_4501),
.Y(n_4605)
);

NAND2xp5_ASAP7_75t_L g4606 ( 
.A(n_4593),
.B(n_4560),
.Y(n_4606)
);

INVx1_ASAP7_75t_L g4607 ( 
.A(n_4596),
.Y(n_4607)
);

INVx1_ASAP7_75t_L g4608 ( 
.A(n_4590),
.Y(n_4608)
);

OAI21xp33_ASAP7_75t_L g4609 ( 
.A1(n_4597),
.A2(n_4529),
.B(n_4518),
.Y(n_4609)
);

INVx1_ASAP7_75t_L g4610 ( 
.A(n_4606),
.Y(n_4610)
);

NAND2xp33_ASAP7_75t_R g4611 ( 
.A(n_4601),
.B(n_4480),
.Y(n_4611)
);

AOI21xp33_ASAP7_75t_SL g4612 ( 
.A1(n_4598),
.A2(n_4605),
.B(n_4609),
.Y(n_4612)
);

AOI322xp5_ASAP7_75t_L g4613 ( 
.A1(n_4599),
.A2(n_4602),
.A3(n_4603),
.B1(n_4608),
.B2(n_4600),
.C1(n_4607),
.C2(n_4496),
.Y(n_4613)
);

INVx1_ASAP7_75t_L g4614 ( 
.A(n_4604),
.Y(n_4614)
);

INVx1_ASAP7_75t_L g4615 ( 
.A(n_4606),
.Y(n_4615)
);

INVx1_ASAP7_75t_L g4616 ( 
.A(n_4606),
.Y(n_4616)
);

AOI221xp5_ASAP7_75t_L g4617 ( 
.A1(n_4598),
.A2(n_4531),
.B1(n_4514),
.B2(n_4520),
.C(n_4532),
.Y(n_4617)
);

AOI222xp33_ASAP7_75t_L g4618 ( 
.A1(n_4602),
.A2(n_4536),
.B1(n_4534),
.B2(n_4520),
.C1(n_4531),
.C2(n_4555),
.Y(n_4618)
);

NOR2xp33_ASAP7_75t_L g4619 ( 
.A(n_4612),
.B(n_4564),
.Y(n_4619)
);

INVx1_ASAP7_75t_L g4620 ( 
.A(n_4610),
.Y(n_4620)
);

NAND2xp5_ASAP7_75t_L g4621 ( 
.A(n_4617),
.B(n_4527),
.Y(n_4621)
);

INVx1_ASAP7_75t_L g4622 ( 
.A(n_4615),
.Y(n_4622)
);

INVx1_ASAP7_75t_SL g4623 ( 
.A(n_4616),
.Y(n_4623)
);

INVxp67_ASAP7_75t_L g4624 ( 
.A(n_4611),
.Y(n_4624)
);

NOR2xp33_ASAP7_75t_L g4625 ( 
.A(n_4614),
.B(n_4518),
.Y(n_4625)
);

INVx1_ASAP7_75t_L g4626 ( 
.A(n_4618),
.Y(n_4626)
);

OAI221xp5_ASAP7_75t_L g4627 ( 
.A1(n_4619),
.A2(n_4613),
.B1(n_4526),
.B2(n_4475),
.C(n_4536),
.Y(n_4627)
);

NAND4xp25_ASAP7_75t_L g4628 ( 
.A(n_4625),
.B(n_4526),
.C(n_4529),
.D(n_4518),
.Y(n_4628)
);

INVx1_ASAP7_75t_L g4629 ( 
.A(n_4621),
.Y(n_4629)
);

INVx1_ASAP7_75t_L g4630 ( 
.A(n_4626),
.Y(n_4630)
);

NAND2xp5_ASAP7_75t_SL g4631 ( 
.A(n_4623),
.B(n_4529),
.Y(n_4631)
);

AOI221xp5_ASAP7_75t_L g4632 ( 
.A1(n_4624),
.A2(n_4534),
.B1(n_4535),
.B2(n_4532),
.C(n_4529),
.Y(n_4632)
);

NAND4xp25_ASAP7_75t_L g4633 ( 
.A(n_4620),
.B(n_4535),
.C(n_4539),
.D(n_4540),
.Y(n_4633)
);

INVx2_ASAP7_75t_L g4634 ( 
.A(n_4622),
.Y(n_4634)
);

NAND2xp5_ASAP7_75t_L g4635 ( 
.A(n_4625),
.B(n_4539),
.Y(n_4635)
);

NOR3x1_ASAP7_75t_L g4636 ( 
.A(n_4621),
.B(n_4509),
.C(n_4504),
.Y(n_4636)
);

NOR2xp33_ASAP7_75t_L g4637 ( 
.A(n_4625),
.B(n_4539),
.Y(n_4637)
);

OAI211xp5_ASAP7_75t_SL g4638 ( 
.A1(n_4624),
.A2(n_4496),
.B(n_4500),
.C(n_4404),
.Y(n_4638)
);

OA21x2_ASAP7_75t_L g4639 ( 
.A1(n_4626),
.A2(n_4500),
.B(n_4540),
.Y(n_4639)
);

NAND3xp33_ASAP7_75t_L g4640 ( 
.A(n_4625),
.B(n_4540),
.C(n_4499),
.Y(n_4640)
);

NAND4xp25_ASAP7_75t_SL g4641 ( 
.A(n_4623),
.B(n_4471),
.C(n_4460),
.D(n_4462),
.Y(n_4641)
);

AOI211xp5_ASAP7_75t_L g4642 ( 
.A1(n_4627),
.A2(n_4540),
.B(n_4497),
.C(n_4403),
.Y(n_4642)
);

AOI21xp5_ASAP7_75t_L g4643 ( 
.A1(n_4631),
.A2(n_4404),
.B(n_4443),
.Y(n_4643)
);

NAND2xp5_ASAP7_75t_L g4644 ( 
.A(n_4637),
.B(n_4472),
.Y(n_4644)
);

NOR2x1_ASAP7_75t_L g4645 ( 
.A(n_4639),
.B(n_4362),
.Y(n_4645)
);

NOR3xp33_ASAP7_75t_L g4646 ( 
.A(n_4629),
.B(n_4186),
.C(n_4443),
.Y(n_4646)
);

OAI221xp5_ASAP7_75t_L g4647 ( 
.A1(n_4628),
.A2(n_4357),
.B1(n_4472),
.B2(n_4344),
.C(n_4401),
.Y(n_4647)
);

NOR2xp33_ASAP7_75t_L g4648 ( 
.A(n_4638),
.B(n_4203),
.Y(n_4648)
);

OR2x2_ASAP7_75t_L g4649 ( 
.A(n_4641),
.B(n_4465),
.Y(n_4649)
);

NAND2xp5_ASAP7_75t_L g4650 ( 
.A(n_4632),
.B(n_4415),
.Y(n_4650)
);

NAND4xp75_ASAP7_75t_L g4651 ( 
.A(n_4630),
.B(n_4401),
.C(n_4462),
.D(n_4351),
.Y(n_4651)
);

NOR2xp33_ASAP7_75t_L g4652 ( 
.A(n_4635),
.B(n_4415),
.Y(n_4652)
);

NOR2xp33_ASAP7_75t_L g4653 ( 
.A(n_4640),
.B(n_4463),
.Y(n_4653)
);

NAND2xp5_ASAP7_75t_L g4654 ( 
.A(n_4636),
.B(n_4463),
.Y(n_4654)
);

INVx1_ASAP7_75t_L g4655 ( 
.A(n_4633),
.Y(n_4655)
);

NAND2xp5_ASAP7_75t_L g4656 ( 
.A(n_4634),
.B(n_4464),
.Y(n_4656)
);

NAND2xp5_ASAP7_75t_SL g4657 ( 
.A(n_4640),
.B(n_4344),
.Y(n_4657)
);

AND3x1_ASAP7_75t_L g4658 ( 
.A(n_4637),
.B(n_4369),
.C(n_4367),
.Y(n_4658)
);

OAI21xp5_ASAP7_75t_SL g4659 ( 
.A1(n_4638),
.A2(n_4369),
.B(n_4367),
.Y(n_4659)
);

INVx1_ASAP7_75t_L g4660 ( 
.A(n_4635),
.Y(n_4660)
);

NAND2xp5_ASAP7_75t_L g4661 ( 
.A(n_4637),
.B(n_4464),
.Y(n_4661)
);

NAND2xp5_ASAP7_75t_L g4662 ( 
.A(n_4637),
.B(n_4418),
.Y(n_4662)
);

INVxp67_ASAP7_75t_L g4663 ( 
.A(n_4637),
.Y(n_4663)
);

NAND2xp5_ASAP7_75t_L g4664 ( 
.A(n_4637),
.B(n_4418),
.Y(n_4664)
);

O2A1O1Ixp33_ASAP7_75t_L g4665 ( 
.A1(n_4631),
.A2(n_4357),
.B(n_4289),
.C(n_4480),
.Y(n_4665)
);

NAND3xp33_ASAP7_75t_L g4666 ( 
.A(n_4645),
.B(n_4655),
.C(n_4663),
.Y(n_4666)
);

BUFx2_ASAP7_75t_L g4667 ( 
.A(n_4658),
.Y(n_4667)
);

OAI21xp5_ASAP7_75t_SL g4668 ( 
.A1(n_4652),
.A2(n_4386),
.B(n_4309),
.Y(n_4668)
);

INVx1_ASAP7_75t_L g4669 ( 
.A(n_4650),
.Y(n_4669)
);

NOR3xp33_ASAP7_75t_L g4670 ( 
.A(n_4660),
.B(n_4289),
.C(n_4272),
.Y(n_4670)
);

NAND2xp5_ASAP7_75t_L g4671 ( 
.A(n_4642),
.B(n_4659),
.Y(n_4671)
);

NAND5xp2_ASAP7_75t_L g4672 ( 
.A(n_4648),
.B(n_4286),
.C(n_4386),
.D(n_4374),
.E(n_4395),
.Y(n_4672)
);

INVx1_ASAP7_75t_L g4673 ( 
.A(n_4661),
.Y(n_4673)
);

NOR3xp33_ASAP7_75t_L g4674 ( 
.A(n_4646),
.B(n_4656),
.C(n_4644),
.Y(n_4674)
);

NAND4xp75_ASAP7_75t_L g4675 ( 
.A(n_4657),
.B(n_4401),
.C(n_4351),
.D(n_4437),
.Y(n_4675)
);

NOR2xp33_ASAP7_75t_L g4676 ( 
.A(n_4653),
.B(n_4465),
.Y(n_4676)
);

NOR3xp33_ASAP7_75t_L g4677 ( 
.A(n_4654),
.B(n_4664),
.C(n_4662),
.Y(n_4677)
);

NAND2xp5_ASAP7_75t_L g4678 ( 
.A(n_4643),
.B(n_4423),
.Y(n_4678)
);

NOR2xp33_ASAP7_75t_L g4679 ( 
.A(n_4649),
.B(n_4360),
.Y(n_4679)
);

AOI221xp5_ASAP7_75t_L g4680 ( 
.A1(n_4665),
.A2(n_4265),
.B1(n_4427),
.B2(n_4432),
.C(n_4423),
.Y(n_4680)
);

AOI211x1_ASAP7_75t_SL g4681 ( 
.A1(n_4647),
.A2(n_4432),
.B(n_4427),
.C(n_4409),
.Y(n_4681)
);

NAND4xp25_ASAP7_75t_L g4682 ( 
.A(n_4651),
.B(n_4178),
.C(n_4360),
.D(n_4380),
.Y(n_4682)
);

AOI22xp33_ASAP7_75t_SL g4683 ( 
.A1(n_4652),
.A2(n_4401),
.B1(n_4357),
.B2(n_4441),
.Y(n_4683)
);

AND2x2_ASAP7_75t_L g4684 ( 
.A(n_4658),
.B(n_4439),
.Y(n_4684)
);

AOI221xp5_ASAP7_75t_L g4685 ( 
.A1(n_4653),
.A2(n_4470),
.B1(n_4467),
.B2(n_4437),
.C(n_4456),
.Y(n_4685)
);

NAND3xp33_ASAP7_75t_L g4686 ( 
.A(n_4645),
.B(n_4409),
.C(n_4408),
.Y(n_4686)
);

O2A1O1Ixp33_ASAP7_75t_L g4687 ( 
.A1(n_4655),
.A2(n_4408),
.B(n_4467),
.C(n_4470),
.Y(n_4687)
);

A2O1A1Ixp33_ASAP7_75t_L g4688 ( 
.A1(n_4652),
.A2(n_4444),
.B(n_4456),
.C(n_4455),
.Y(n_4688)
);

NOR4xp25_ASAP7_75t_L g4689 ( 
.A(n_4655),
.B(n_4444),
.C(n_4455),
.D(n_4450),
.Y(n_4689)
);

NAND2xp5_ASAP7_75t_SL g4690 ( 
.A(n_4645),
.B(n_4441),
.Y(n_4690)
);

NAND2x1_ASAP7_75t_SL g4691 ( 
.A(n_4645),
.B(n_4447),
.Y(n_4691)
);

NAND3xp33_ASAP7_75t_L g4692 ( 
.A(n_4645),
.B(n_4450),
.C(n_4447),
.Y(n_4692)
);

NAND2xp5_ASAP7_75t_L g4693 ( 
.A(n_4642),
.B(n_4374),
.Y(n_4693)
);

NAND4xp25_ASAP7_75t_L g4694 ( 
.A(n_4666),
.B(n_4380),
.C(n_4348),
.D(n_4395),
.Y(n_4694)
);

NOR2xp33_ASAP7_75t_SL g4695 ( 
.A(n_4667),
.B(n_4424),
.Y(n_4695)
);

NAND5xp2_ASAP7_75t_L g4696 ( 
.A(n_4674),
.B(n_4394),
.C(n_4376),
.D(n_4294),
.E(n_4416),
.Y(n_4696)
);

NOR3xp33_ASAP7_75t_L g4697 ( 
.A(n_4671),
.B(n_4348),
.C(n_4411),
.Y(n_4697)
);

INVx1_ASAP7_75t_L g4698 ( 
.A(n_4684),
.Y(n_4698)
);

NAND2xp5_ASAP7_75t_L g4699 ( 
.A(n_4679),
.B(n_4376),
.Y(n_4699)
);

OAI321xp33_ASAP7_75t_L g4700 ( 
.A1(n_4690),
.A2(n_4420),
.A3(n_4412),
.B1(n_4414),
.B2(n_4416),
.C(n_4421),
.Y(n_4700)
);

NAND3xp33_ASAP7_75t_L g4701 ( 
.A(n_4677),
.B(n_4412),
.C(n_4411),
.Y(n_4701)
);

NOR3xp33_ASAP7_75t_L g4702 ( 
.A(n_4669),
.B(n_4420),
.C(n_4414),
.Y(n_4702)
);

AOI211xp5_ASAP7_75t_L g4703 ( 
.A1(n_4673),
.A2(n_4421),
.B(n_4466),
.C(n_4285),
.Y(n_4703)
);

AOI222xp33_ASAP7_75t_L g4704 ( 
.A1(n_4680),
.A2(n_4466),
.B1(n_4394),
.B2(n_4441),
.C1(n_4309),
.C2(n_4439),
.Y(n_4704)
);

NOR2xp33_ASAP7_75t_L g4705 ( 
.A(n_4693),
.B(n_4424),
.Y(n_4705)
);

NOR5xp2_ASAP7_75t_L g4706 ( 
.A(n_4686),
.B(n_4377),
.C(n_4441),
.D(n_4373),
.E(n_4372),
.Y(n_4706)
);

NOR3xp33_ASAP7_75t_L g4707 ( 
.A(n_4678),
.B(n_4381),
.C(n_4309),
.Y(n_4707)
);

NOR3xp33_ASAP7_75t_L g4708 ( 
.A(n_4676),
.B(n_4377),
.C(n_4424),
.Y(n_4708)
);

NAND3xp33_ASAP7_75t_L g4709 ( 
.A(n_4692),
.B(n_4351),
.C(n_4183),
.Y(n_4709)
);

NOR2x1_ASAP7_75t_L g4710 ( 
.A(n_4682),
.B(n_4355),
.Y(n_4710)
);

NAND2xp5_ASAP7_75t_L g4711 ( 
.A(n_4670),
.B(n_4668),
.Y(n_4711)
);

NAND3xp33_ASAP7_75t_SL g4712 ( 
.A(n_4681),
.B(n_4391),
.C(n_4373),
.Y(n_4712)
);

AOI221xp5_ASAP7_75t_SL g4713 ( 
.A1(n_4687),
.A2(n_4372),
.B1(n_4391),
.B2(n_4315),
.C(n_4323),
.Y(n_4713)
);

NAND2xp5_ASAP7_75t_L g4714 ( 
.A(n_4691),
.B(n_4689),
.Y(n_4714)
);

INVx1_ASAP7_75t_L g4715 ( 
.A(n_4688),
.Y(n_4715)
);

NAND4xp25_ASAP7_75t_SL g4716 ( 
.A(n_4685),
.B(n_4378),
.C(n_4324),
.D(n_4315),
.Y(n_4716)
);

AOI21xp33_ASAP7_75t_L g4717 ( 
.A1(n_4683),
.A2(n_4355),
.B(n_4351),
.Y(n_4717)
);

XNOR2x1_ASAP7_75t_L g4718 ( 
.A(n_4675),
.B(n_274),
.Y(n_4718)
);

XOR2xp5_ASAP7_75t_L g4719 ( 
.A(n_4718),
.B(n_275),
.Y(n_4719)
);

INVx1_ASAP7_75t_SL g4720 ( 
.A(n_4695),
.Y(n_4720)
);

NAND2xp5_ASAP7_75t_L g4721 ( 
.A(n_4703),
.B(n_4672),
.Y(n_4721)
);

AND2x2_ASAP7_75t_L g4722 ( 
.A(n_4705),
.B(n_4697),
.Y(n_4722)
);

INVx2_ASAP7_75t_SL g4723 ( 
.A(n_4698),
.Y(n_4723)
);

AND2x2_ASAP7_75t_L g4724 ( 
.A(n_4708),
.B(n_4378),
.Y(n_4724)
);

AOI211xp5_ASAP7_75t_L g4725 ( 
.A1(n_4711),
.A2(n_4210),
.B(n_277),
.C(n_278),
.Y(n_4725)
);

HB1xp67_ASAP7_75t_L g4726 ( 
.A(n_4714),
.Y(n_4726)
);

NOR2xp33_ASAP7_75t_L g4727 ( 
.A(n_4699),
.B(n_4223),
.Y(n_4727)
);

NOR2xp33_ASAP7_75t_L g4728 ( 
.A(n_4701),
.B(n_4715),
.Y(n_4728)
);

NAND2xp5_ASAP7_75t_L g4729 ( 
.A(n_4702),
.B(n_4223),
.Y(n_4729)
);

NOR3xp33_ASAP7_75t_L g4730 ( 
.A(n_4710),
.B(n_276),
.C(n_278),
.Y(n_4730)
);

AOI211xp5_ASAP7_75t_L g4731 ( 
.A1(n_4717),
.A2(n_280),
.B(n_282),
.C(n_283),
.Y(n_4731)
);

INVx1_ASAP7_75t_L g4732 ( 
.A(n_4712),
.Y(n_4732)
);

INVxp67_ASAP7_75t_SL g4733 ( 
.A(n_4706),
.Y(n_4733)
);

NOR2xp33_ASAP7_75t_R g4734 ( 
.A(n_4716),
.B(n_280),
.Y(n_4734)
);

INVx1_ASAP7_75t_SL g4735 ( 
.A(n_4709),
.Y(n_4735)
);

OAI21xp33_ASAP7_75t_L g4736 ( 
.A1(n_4707),
.A2(n_4324),
.B(n_4339),
.Y(n_4736)
);

INVx2_ASAP7_75t_L g4737 ( 
.A(n_4729),
.Y(n_4737)
);

AND2x4_ASAP7_75t_L g4738 ( 
.A(n_4723),
.B(n_4696),
.Y(n_4738)
);

INVx1_ASAP7_75t_L g4739 ( 
.A(n_4727),
.Y(n_4739)
);

INVx1_ASAP7_75t_L g4740 ( 
.A(n_4719),
.Y(n_4740)
);

AOI22xp5_ASAP7_75t_L g4741 ( 
.A1(n_4720),
.A2(n_4694),
.B1(n_4704),
.B2(n_4713),
.Y(n_4741)
);

OA211x2_ASAP7_75t_L g4742 ( 
.A1(n_4728),
.A2(n_4700),
.B(n_284),
.C(n_285),
.Y(n_4742)
);

NOR2x1_ASAP7_75t_L g4743 ( 
.A(n_4732),
.B(n_4350),
.Y(n_4743)
);

INVx1_ASAP7_75t_L g4744 ( 
.A(n_4724),
.Y(n_4744)
);

XNOR2xp5_ASAP7_75t_L g4745 ( 
.A(n_4731),
.B(n_283),
.Y(n_4745)
);

NOR3xp33_ASAP7_75t_L g4746 ( 
.A(n_4726),
.B(n_285),
.C(n_286),
.Y(n_4746)
);

OR3x2_ASAP7_75t_L g4747 ( 
.A(n_4734),
.B(n_287),
.C(n_288),
.Y(n_4747)
);

NOR2xp33_ASAP7_75t_L g4748 ( 
.A(n_4735),
.B(n_287),
.Y(n_4748)
);

NAND4xp75_ASAP7_75t_L g4749 ( 
.A(n_4722),
.B(n_4340),
.C(n_289),
.D(n_292),
.Y(n_4749)
);

INVxp67_ASAP7_75t_L g4750 ( 
.A(n_4733),
.Y(n_4750)
);

INVx1_ASAP7_75t_L g4751 ( 
.A(n_4730),
.Y(n_4751)
);

AND2x2_ASAP7_75t_L g4752 ( 
.A(n_4725),
.B(n_4339),
.Y(n_4752)
);

NOR3xp33_ASAP7_75t_L g4753 ( 
.A(n_4750),
.B(n_4721),
.C(n_4736),
.Y(n_4753)
);

AND2x2_ASAP7_75t_L g4754 ( 
.A(n_4738),
.B(n_4341),
.Y(n_4754)
);

NOR3x1_ASAP7_75t_L g4755 ( 
.A(n_4751),
.B(n_288),
.C(n_289),
.Y(n_4755)
);

NOR4xp25_ASAP7_75t_L g4756 ( 
.A(n_4744),
.B(n_292),
.C(n_293),
.D(n_295),
.Y(n_4756)
);

NOR3xp33_ASAP7_75t_L g4757 ( 
.A(n_4739),
.B(n_296),
.C(n_298),
.Y(n_4757)
);

NOR2x1_ASAP7_75t_L g4758 ( 
.A(n_4748),
.B(n_4350),
.Y(n_4758)
);

NAND4xp75_ASAP7_75t_L g4759 ( 
.A(n_4742),
.B(n_4340),
.C(n_298),
.D(n_299),
.Y(n_4759)
);

OAI21xp33_ASAP7_75t_L g4760 ( 
.A1(n_4741),
.A2(n_4342),
.B(n_4341),
.Y(n_4760)
);

INVx2_ASAP7_75t_L g4761 ( 
.A(n_4747),
.Y(n_4761)
);

NOR2x1p5_ASAP7_75t_L g4762 ( 
.A(n_4737),
.B(n_296),
.Y(n_4762)
);

NAND3x1_ASAP7_75t_L g4763 ( 
.A(n_4746),
.B(n_4740),
.C(n_4752),
.Y(n_4763)
);

NAND3xp33_ASAP7_75t_L g4764 ( 
.A(n_4745),
.B(n_4340),
.C(n_4345),
.Y(n_4764)
);

NOR3xp33_ASAP7_75t_L g4765 ( 
.A(n_4743),
.B(n_4749),
.C(n_4345),
.Y(n_4765)
);

NOR3xp33_ASAP7_75t_L g4766 ( 
.A(n_4750),
.B(n_4343),
.C(n_4342),
.Y(n_4766)
);

INVx1_ASAP7_75t_L g4767 ( 
.A(n_4748),
.Y(n_4767)
);

AND2x2_ASAP7_75t_L g4768 ( 
.A(n_4750),
.B(n_4343),
.Y(n_4768)
);

OAI21xp5_ASAP7_75t_L g4769 ( 
.A1(n_4750),
.A2(n_4361),
.B(n_4233),
.Y(n_4769)
);

NOR3xp33_ASAP7_75t_L g4770 ( 
.A(n_4750),
.B(n_314),
.C(n_316),
.Y(n_4770)
);

OAI211xp5_ASAP7_75t_SL g4771 ( 
.A1(n_4753),
.A2(n_320),
.B(n_323),
.C(n_324),
.Y(n_4771)
);

AND3x4_ASAP7_75t_L g4772 ( 
.A(n_4765),
.B(n_329),
.C(n_330),
.Y(n_4772)
);

INVx2_ASAP7_75t_L g4773 ( 
.A(n_4755),
.Y(n_4773)
);

INVx1_ASAP7_75t_L g4774 ( 
.A(n_4762),
.Y(n_4774)
);

CKINVDCx5p33_ASAP7_75t_R g4775 ( 
.A(n_4761),
.Y(n_4775)
);

INVx1_ASAP7_75t_L g4776 ( 
.A(n_4768),
.Y(n_4776)
);

BUFx3_ASAP7_75t_L g4777 ( 
.A(n_4754),
.Y(n_4777)
);

CKINVDCx5p33_ASAP7_75t_R g4778 ( 
.A(n_4767),
.Y(n_4778)
);

CKINVDCx5p33_ASAP7_75t_R g4779 ( 
.A(n_4763),
.Y(n_4779)
);

NAND2xp5_ASAP7_75t_SL g4780 ( 
.A(n_4756),
.B(n_4282),
.Y(n_4780)
);

INVx1_ASAP7_75t_SL g4781 ( 
.A(n_4759),
.Y(n_4781)
);

INVx1_ASAP7_75t_SL g4782 ( 
.A(n_4757),
.Y(n_4782)
);

AND3x4_ASAP7_75t_L g4783 ( 
.A(n_4766),
.B(n_4770),
.C(n_4760),
.Y(n_4783)
);

OAI22xp5_ASAP7_75t_SL g4784 ( 
.A1(n_4781),
.A2(n_4769),
.B1(n_4764),
.B2(n_4758),
.Y(n_4784)
);

OAI22xp5_ASAP7_75t_L g4785 ( 
.A1(n_4779),
.A2(n_4361),
.B1(n_4225),
.B2(n_1412),
.Y(n_4785)
);

AND2x2_ASAP7_75t_L g4786 ( 
.A(n_4773),
.B(n_4361),
.Y(n_4786)
);

OAI211xp5_ASAP7_75t_SL g4787 ( 
.A1(n_4782),
.A2(n_331),
.B(n_333),
.C(n_336),
.Y(n_4787)
);

A2O1A1Ixp33_ASAP7_75t_L g4788 ( 
.A1(n_4777),
.A2(n_4225),
.B(n_343),
.C(n_344),
.Y(n_4788)
);

NOR3xp33_ASAP7_75t_L g4789 ( 
.A(n_4776),
.B(n_338),
.C(n_346),
.Y(n_4789)
);

AND2x2_ASAP7_75t_L g4790 ( 
.A(n_4774),
.B(n_4361),
.Y(n_4790)
);

INVx1_ASAP7_75t_L g4791 ( 
.A(n_4784),
.Y(n_4791)
);

INVx1_ASAP7_75t_L g4792 ( 
.A(n_4786),
.Y(n_4792)
);

INVx1_ASAP7_75t_L g4793 ( 
.A(n_4790),
.Y(n_4793)
);

OAI22x1_ASAP7_75t_L g4794 ( 
.A1(n_4789),
.A2(n_4772),
.B1(n_4783),
.B2(n_4775),
.Y(n_4794)
);

AOI22xp5_ASAP7_75t_L g4795 ( 
.A1(n_4787),
.A2(n_4778),
.B1(n_4771),
.B2(n_4780),
.Y(n_4795)
);

INVx1_ASAP7_75t_L g4796 ( 
.A(n_4788),
.Y(n_4796)
);

INVx1_ASAP7_75t_L g4797 ( 
.A(n_4785),
.Y(n_4797)
);

INVx1_ASAP7_75t_L g4798 ( 
.A(n_4793),
.Y(n_4798)
);

NAND2xp5_ASAP7_75t_L g4799 ( 
.A(n_4792),
.B(n_348),
.Y(n_4799)
);

AND3x1_ASAP7_75t_L g4800 ( 
.A(n_4791),
.B(n_350),
.C(n_353),
.Y(n_4800)
);

NOR3x2_ASAP7_75t_L g4801 ( 
.A(n_4794),
.B(n_354),
.C(n_355),
.Y(n_4801)
);

AOI21xp5_ASAP7_75t_L g4802 ( 
.A1(n_4796),
.A2(n_4797),
.B(n_4795),
.Y(n_4802)
);

XNOR2xp5_ASAP7_75t_L g4803 ( 
.A(n_4794),
.B(n_357),
.Y(n_4803)
);

XOR2xp5_ASAP7_75t_L g4804 ( 
.A(n_4803),
.B(n_4802),
.Y(n_4804)
);

OAI22xp5_ASAP7_75t_L g4805 ( 
.A1(n_4798),
.A2(n_1412),
.B1(n_362),
.B2(n_363),
.Y(n_4805)
);

INVx1_ASAP7_75t_L g4806 ( 
.A(n_4800),
.Y(n_4806)
);

OA21x2_ASAP7_75t_L g4807 ( 
.A1(n_4799),
.A2(n_4801),
.B(n_367),
.Y(n_4807)
);

INVx1_ASAP7_75t_L g4808 ( 
.A(n_4803),
.Y(n_4808)
);

AOI22x1_ASAP7_75t_L g4809 ( 
.A1(n_4804),
.A2(n_359),
.B1(n_371),
.B2(n_372),
.Y(n_4809)
);

AOI21xp5_ASAP7_75t_L g4810 ( 
.A1(n_4806),
.A2(n_1412),
.B(n_1863),
.Y(n_4810)
);

INVx2_ASAP7_75t_L g4811 ( 
.A(n_4807),
.Y(n_4811)
);

OAI22xp5_ASAP7_75t_SL g4812 ( 
.A1(n_4808),
.A2(n_4805),
.B1(n_375),
.B2(n_377),
.Y(n_4812)
);

AOI22xp5_ASAP7_75t_L g4813 ( 
.A1(n_4812),
.A2(n_374),
.B1(n_379),
.B2(n_380),
.Y(n_4813)
);

OAI22xp5_ASAP7_75t_L g4814 ( 
.A1(n_4811),
.A2(n_381),
.B1(n_383),
.B2(n_384),
.Y(n_4814)
);

AOI21xp5_ASAP7_75t_L g4815 ( 
.A1(n_4810),
.A2(n_1870),
.B(n_1863),
.Y(n_4815)
);

AOI21x1_ASAP7_75t_L g4816 ( 
.A1(n_4809),
.A2(n_389),
.B(n_390),
.Y(n_4816)
);

AOI21x1_ASAP7_75t_L g4817 ( 
.A1(n_4811),
.A2(n_393),
.B(n_397),
.Y(n_4817)
);

OAI21xp33_ASAP7_75t_L g4818 ( 
.A1(n_4813),
.A2(n_398),
.B(n_399),
.Y(n_4818)
);

OR2x2_ASAP7_75t_L g4819 ( 
.A(n_4815),
.B(n_407),
.Y(n_4819)
);

INVxp33_ASAP7_75t_SL g4820 ( 
.A(n_4814),
.Y(n_4820)
);

OAI21xp5_ASAP7_75t_L g4821 ( 
.A1(n_4816),
.A2(n_409),
.B(n_410),
.Y(n_4821)
);

AOI22xp33_ASAP7_75t_L g4822 ( 
.A1(n_4817),
.A2(n_1870),
.B1(n_1860),
.B2(n_1859),
.Y(n_4822)
);

AOI21xp5_ASAP7_75t_L g4823 ( 
.A1(n_4815),
.A2(n_1860),
.B(n_1859),
.Y(n_4823)
);

INVx3_ASAP7_75t_SL g4824 ( 
.A(n_4816),
.Y(n_4824)
);

AOI21xp5_ASAP7_75t_L g4825 ( 
.A1(n_4815),
.A2(n_1860),
.B(n_1859),
.Y(n_4825)
);

INVx1_ASAP7_75t_L g4826 ( 
.A(n_4816),
.Y(n_4826)
);

AOI21xp5_ASAP7_75t_L g4827 ( 
.A1(n_4815),
.A2(n_1860),
.B(n_1836),
.Y(n_4827)
);

AOI22xp33_ASAP7_75t_L g4828 ( 
.A1(n_4820),
.A2(n_1836),
.B1(n_1824),
.B2(n_1451),
.Y(n_4828)
);

AOI22xp33_ASAP7_75t_L g4829 ( 
.A1(n_4818),
.A2(n_4826),
.B1(n_4824),
.B2(n_4821),
.Y(n_4829)
);

OAI22xp33_ASAP7_75t_L g4830 ( 
.A1(n_4819),
.A2(n_4827),
.B1(n_4825),
.B2(n_4823),
.Y(n_4830)
);

AOI22xp5_ASAP7_75t_L g4831 ( 
.A1(n_4822),
.A2(n_411),
.B1(n_413),
.B2(n_418),
.Y(n_4831)
);

AOI22xp33_ASAP7_75t_L g4832 ( 
.A1(n_4820),
.A2(n_1824),
.B1(n_1451),
.B2(n_1450),
.Y(n_4832)
);

AO22x2_ASAP7_75t_L g4833 ( 
.A1(n_4826),
.A2(n_420),
.B1(n_424),
.B2(n_425),
.Y(n_4833)
);

AOI22xp33_ASAP7_75t_L g4834 ( 
.A1(n_4820),
.A2(n_1451),
.B1(n_1450),
.B2(n_1442),
.Y(n_4834)
);

AOI22xp5_ASAP7_75t_L g4835 ( 
.A1(n_4820),
.A2(n_429),
.B1(n_430),
.B2(n_432),
.Y(n_4835)
);

AOI22xp5_ASAP7_75t_L g4836 ( 
.A1(n_4820),
.A2(n_433),
.B1(n_441),
.B2(n_442),
.Y(n_4836)
);

AO22x2_ASAP7_75t_L g4837 ( 
.A1(n_4826),
.A2(n_443),
.B1(n_446),
.B2(n_447),
.Y(n_4837)
);

NOR2x1_ASAP7_75t_L g4838 ( 
.A(n_4830),
.B(n_1768),
.Y(n_4838)
);

AOI21xp5_ASAP7_75t_L g4839 ( 
.A1(n_4829),
.A2(n_1451),
.B(n_1425),
.Y(n_4839)
);

OAI21x1_ASAP7_75t_L g4840 ( 
.A1(n_4828),
.A2(n_4832),
.B(n_4834),
.Y(n_4840)
);

OAI21xp5_ASAP7_75t_L g4841 ( 
.A1(n_4831),
.A2(n_452),
.B(n_453),
.Y(n_4841)
);

AO21x2_ASAP7_75t_L g4842 ( 
.A1(n_4835),
.A2(n_461),
.B(n_467),
.Y(n_4842)
);

OAI21xp5_ASAP7_75t_L g4843 ( 
.A1(n_4836),
.A2(n_469),
.B(n_470),
.Y(n_4843)
);

OAI21x1_ASAP7_75t_L g4844 ( 
.A1(n_4833),
.A2(n_472),
.B(n_473),
.Y(n_4844)
);

AO221x2_ASAP7_75t_L g4845 ( 
.A1(n_4837),
.A2(n_474),
.B1(n_477),
.B2(n_479),
.C(n_481),
.Y(n_4845)
);

OAI21xp5_ASAP7_75t_SL g4846 ( 
.A1(n_4829),
.A2(n_482),
.B(n_492),
.Y(n_4846)
);

INVxp67_ASAP7_75t_L g4847 ( 
.A(n_4838),
.Y(n_4847)
);

AOI22xp33_ASAP7_75t_L g4848 ( 
.A1(n_4842),
.A2(n_1450),
.B1(n_1442),
.B2(n_1425),
.Y(n_4848)
);

OAI22xp33_ASAP7_75t_L g4849 ( 
.A1(n_4843),
.A2(n_497),
.B1(n_498),
.B2(n_500),
.Y(n_4849)
);

AOI22x1_ASAP7_75t_L g4850 ( 
.A1(n_4839),
.A2(n_502),
.B1(n_506),
.B2(n_509),
.Y(n_4850)
);

AOI221xp5_ASAP7_75t_L g4851 ( 
.A1(n_4847),
.A2(n_4841),
.B1(n_4846),
.B2(n_4844),
.C(n_4840),
.Y(n_4851)
);

AOI21xp5_ASAP7_75t_L g4852 ( 
.A1(n_4851),
.A2(n_4848),
.B(n_4849),
.Y(n_4852)
);

AOI211xp5_ASAP7_75t_L g4853 ( 
.A1(n_4852),
.A2(n_4850),
.B(n_4845),
.C(n_517),
.Y(n_4853)
);


endmodule