module fake_jpeg_3386_n_155 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_39, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_155);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_39;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_155;

wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_73;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_150;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_6),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_37),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_23),
.Y(n_43)
);

BUFx5_ASAP7_75t_L g44 ( 
.A(n_21),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_17),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_11),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_40),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_20),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_14),
.Y(n_49)
);

BUFx5_ASAP7_75t_L g50 ( 
.A(n_39),
.Y(n_50)
);

INVx11_ASAP7_75t_L g51 ( 
.A(n_22),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_24),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_9),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_2),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_7),
.Y(n_55)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_55),
.Y(n_56)
);

INVx2_ASAP7_75t_SL g73 ( 
.A(n_56),
.Y(n_73)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_51),
.Y(n_57)
);

INVx5_ASAP7_75t_L g67 ( 
.A(n_57),
.Y(n_67)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_51),
.Y(n_58)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_58),
.Y(n_72)
);

INVx11_ASAP7_75t_L g59 ( 
.A(n_52),
.Y(n_59)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_59),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_54),
.B(n_41),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_60),
.B(n_49),
.Y(n_65)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_52),
.Y(n_61)
);

BUFx12f_ASAP7_75t_L g69 ( 
.A(n_61),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_53),
.B(n_0),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_SL g68 ( 
.A(n_62),
.B(n_42),
.Y(n_68)
);

AND2x2_ASAP7_75t_L g63 ( 
.A(n_60),
.B(n_52),
.Y(n_63)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_63),
.B(n_71),
.C(n_66),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_56),
.A2(n_55),
.B1(n_43),
.B2(n_54),
.Y(n_64)
);

OAI22xp33_ASAP7_75t_L g76 ( 
.A1(n_64),
.A2(n_59),
.B1(n_50),
.B2(n_44),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_65),
.B(n_46),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_57),
.Y(n_66)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_66),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_68),
.B(n_0),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_58),
.Y(n_71)
);

INVx1_ASAP7_75t_SL g79 ( 
.A(n_71),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_64),
.A2(n_55),
.B1(n_62),
.B2(n_43),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_74),
.A2(n_76),
.B1(n_61),
.B2(n_67),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g91 ( 
.A(n_75),
.B(n_88),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_63),
.B(n_45),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_77),
.B(n_80),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_SL g78 ( 
.A(n_73),
.B(n_47),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_78),
.B(n_84),
.Y(n_97)
);

INVx1_ASAP7_75t_SL g80 ( 
.A(n_73),
.Y(n_80)
);

INVxp67_ASAP7_75t_SL g81 ( 
.A(n_69),
.Y(n_81)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_81),
.Y(n_93)
);

INVx1_ASAP7_75t_SL g82 ( 
.A(n_69),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_82),
.B(n_83),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_72),
.B(n_48),
.Y(n_83)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_69),
.Y(n_86)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_86),
.Y(n_102)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_67),
.Y(n_87)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_87),
.Y(n_104)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_85),
.Y(n_89)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_89),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_80),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_90),
.B(n_92),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_85),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g96 ( 
.A(n_82),
.B(n_1),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_96),
.B(n_101),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_SL g118 ( 
.A1(n_98),
.A2(n_103),
.B(n_3),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_79),
.A2(n_61),
.B1(n_70),
.B2(n_50),
.Y(n_99)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_99),
.Y(n_106)
);

AOI21xp5_ASAP7_75t_L g100 ( 
.A1(n_81),
.A2(n_79),
.B(n_70),
.Y(n_100)
);

AOI21xp5_ASAP7_75t_L g121 ( 
.A1(n_100),
.A2(n_26),
.B(n_35),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_84),
.B(n_19),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_74),
.A2(n_44),
.B1(n_2),
.B2(n_3),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_97),
.B(n_18),
.C(n_36),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_105),
.B(n_110),
.Y(n_130)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_104),
.Y(n_108)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_108),
.Y(n_123)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_95),
.Y(n_109)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_109),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_91),
.B(n_1),
.Y(n_110)
);

CKINVDCx16_ASAP7_75t_R g112 ( 
.A(n_100),
.Y(n_112)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_112),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_94),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_113),
.Y(n_124)
);

XOR2xp5_ASAP7_75t_L g114 ( 
.A(n_101),
.B(n_25),
.Y(n_114)
);

AOI21xp5_ASAP7_75t_L g125 ( 
.A1(n_114),
.A2(n_116),
.B(n_99),
.Y(n_125)
);

XOR2xp5_ASAP7_75t_L g116 ( 
.A(n_98),
.B(n_16),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_102),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_117),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_118),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_103),
.B(n_4),
.Y(n_119)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_119),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_89),
.Y(n_120)
);

AO21x1_ASAP7_75t_L g122 ( 
.A1(n_120),
.A2(n_121),
.B(n_93),
.Y(n_122)
);

AOI21xp5_ASAP7_75t_SL g140 ( 
.A1(n_122),
.A2(n_5),
.B(n_7),
.Y(n_140)
);

XOR2xp5_ASAP7_75t_L g138 ( 
.A(n_125),
.B(n_126),
.Y(n_138)
);

AOI32xp33_ASAP7_75t_L g126 ( 
.A1(n_107),
.A2(n_106),
.A3(n_121),
.B1(n_116),
.B2(n_115),
.Y(n_126)
);

AOI21xp5_ASAP7_75t_L g128 ( 
.A1(n_115),
.A2(n_15),
.B(n_34),
.Y(n_128)
);

OAI21xp33_ASAP7_75t_SL g137 ( 
.A1(n_128),
.A2(n_131),
.B(n_27),
.Y(n_137)
);

O2A1O1Ixp33_ASAP7_75t_L g131 ( 
.A1(n_105),
.A2(n_13),
.B(n_33),
.C(n_32),
.Y(n_131)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_132),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_124),
.B(n_114),
.C(n_111),
.Y(n_136)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_136),
.Y(n_143)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_137),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_134),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_139),
.A2(n_140),
.B1(n_141),
.B2(n_130),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_SL g141 ( 
.A(n_130),
.B(n_127),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_138),
.A2(n_129),
.B1(n_133),
.B2(n_123),
.Y(n_142)
);

XOR2xp5_ASAP7_75t_L g146 ( 
.A(n_142),
.B(n_122),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_144),
.B(n_137),
.C(n_135),
.Y(n_147)
);

XNOR2x1_ASAP7_75t_L g148 ( 
.A(n_146),
.B(n_147),
.Y(n_148)
);

XOR2xp5_ASAP7_75t_L g149 ( 
.A(n_148),
.B(n_143),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_SL g150 ( 
.A1(n_149),
.A2(n_145),
.B(n_142),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_150),
.B(n_131),
.C(n_29),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_151),
.B(n_28),
.C(n_31),
.Y(n_152)
);

AND2x2_ASAP7_75t_L g153 ( 
.A(n_152),
.B(n_12),
.Y(n_153)
);

OAI311xp33_ASAP7_75t_L g154 ( 
.A1(n_153),
.A2(n_30),
.A3(n_38),
.B1(n_10),
.C1(n_8),
.Y(n_154)
);

XOR2xp5_ASAP7_75t_L g155 ( 
.A(n_154),
.B(n_10),
.Y(n_155)
);


endmodule