module real_jpeg_26503_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_68;
wire n_247;
wire n_146;
wire n_83;
wire n_78;
wire n_249;
wire n_215;
wire n_176;
wire n_166;
wire n_221;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_131;
wire n_47;
wire n_163;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_243;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_200;
wire n_48;
wire n_164;
wire n_184;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_13;
wire n_120;
wire n_113;
wire n_155;
wire n_199;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_238;
wire n_67;
wire n_79;
wire n_178;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_44;
wire n_28;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_121;
wire n_234;
wire n_106;
wire n_172;
wire n_160;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_192;
wire n_203;
wire n_100;
wire n_198;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_205;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_228;
wire n_150;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_241;
wire n_103;
wire n_225;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_216;
wire n_244;
wire n_128;
wire n_213;
wire n_167;
wire n_179;
wire n_133;
wire n_202;
wire n_138;
wire n_25;
wire n_217;
wire n_53;
wire n_127;
wire n_210;
wire n_206;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;
wire n_16;

INVx11_ASAP7_75t_SL g63 ( 
.A(n_0),
.Y(n_63)
);

HB1xp67_ASAP7_75t_L g82 ( 
.A(n_1),
.Y(n_82)
);

INVx11_ASAP7_75t_L g103 ( 
.A(n_1),
.Y(n_103)
);

INVx5_ASAP7_75t_L g142 ( 
.A(n_1),
.Y(n_142)
);

BUFx12_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_3),
.A2(n_42),
.B1(n_44),
.B2(n_65),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_3),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_L g77 ( 
.A1(n_3),
.A2(n_61),
.B1(n_62),
.B2(n_65),
.Y(n_77)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_4),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_L g39 ( 
.A1(n_5),
.A2(n_22),
.B1(n_23),
.B2(n_40),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_5),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_5),
.A2(n_40),
.B1(n_42),
.B2(n_44),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_5),
.A2(n_40),
.B1(n_61),
.B2(n_62),
.Y(n_102)
);

BUFx2_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

INVx8_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

INVx11_ASAP7_75t_L g59 ( 
.A(n_8),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_8),
.A2(n_59),
.B1(n_61),
.B2(n_62),
.Y(n_60)
);

AOI21xp33_ASAP7_75t_L g183 ( 
.A1(n_8),
.A2(n_11),
.B(n_62),
.Y(n_183)
);

AOI22xp33_ASAP7_75t_SL g26 ( 
.A1(n_9),
.A2(n_27),
.B1(n_28),
.B2(n_29),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_9),
.Y(n_29)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_9),
.A2(n_22),
.B1(n_23),
.B2(n_29),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_9),
.A2(n_29),
.B1(n_42),
.B2(n_44),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_9),
.A2(n_29),
.B1(n_61),
.B2(n_62),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g41 ( 
.A1(n_10),
.A2(n_42),
.B1(n_43),
.B2(n_44),
.Y(n_41)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_10),
.Y(n_43)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_10),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g31 ( 
.A1(n_11),
.A2(n_27),
.B1(n_28),
.B2(n_32),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_11),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_L g47 ( 
.A1(n_11),
.A2(n_22),
.B1(n_23),
.B2(n_32),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_11),
.A2(n_32),
.B1(n_42),
.B2(n_44),
.Y(n_87)
);

AOI21xp33_ASAP7_75t_SL g124 ( 
.A1(n_11),
.A2(n_22),
.B(n_25),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_11),
.A2(n_32),
.B1(n_61),
.B2(n_62),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_11),
.B(n_21),
.Y(n_155)
);

AOI21xp33_ASAP7_75t_SL g163 ( 
.A1(n_11),
.A2(n_42),
.B(n_50),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_11),
.B(n_41),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_112),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_110),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_SL g14 ( 
.A(n_15),
.B(n_93),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_15),
.B(n_93),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g15 ( 
.A1(n_16),
.A2(n_74),
.B1(n_75),
.B2(n_92),
.Y(n_15)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_16),
.Y(n_92)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_66),
.Y(n_16)
);

AOI22xp5_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_19),
.B1(n_35),
.B2(n_36),
.Y(n_17)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_18),
.A2(n_19),
.B1(n_148),
.B2(n_149),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_18),
.A2(n_19),
.B1(n_226),
.B2(n_227),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_18),
.B(n_224),
.C(n_226),
.Y(n_242)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_19),
.B(n_109),
.C(n_131),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_26),
.B(n_30),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_21),
.B(n_34),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_21),
.B(n_33),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_21),
.A2(n_31),
.B1(n_33),
.B2(n_107),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g21 ( 
.A1(n_22),
.A2(n_23),
.B1(n_24),
.B2(n_25),
.Y(n_21)
);

AOI22xp33_ASAP7_75t_L g49 ( 
.A1(n_22),
.A2(n_23),
.B1(n_43),
.B2(n_50),
.Y(n_49)
);

A2O1A1Ixp33_ASAP7_75t_L g162 ( 
.A1(n_22),
.A2(n_32),
.B(n_51),
.C(n_163),
.Y(n_162)
);

INVx11_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

AOI22xp33_ASAP7_75t_L g34 ( 
.A1(n_24),
.A2(n_25),
.B1(n_27),
.B2(n_28),
.Y(n_34)
);

A2O1A1Ixp33_ASAP7_75t_L g123 ( 
.A1(n_24),
.A2(n_28),
.B(n_32),
.C(n_124),
.Y(n_123)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_26),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_28),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_31),
.B(n_33),
.Y(n_30)
);

CKINVDCx14_ASAP7_75t_R g90 ( 
.A(n_31),
.Y(n_90)
);

A2O1A1Ixp33_ASAP7_75t_L g182 ( 
.A1(n_32),
.A2(n_42),
.B(n_59),
.C(n_183),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_32),
.B(n_197),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_SL g200 ( 
.A(n_32),
.B(n_60),
.Y(n_200)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_L g36 ( 
.A1(n_37),
.A2(n_38),
.B1(n_52),
.B2(n_53),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_38),
.Y(n_37)
);

AOI21xp5_ASAP7_75t_L g38 ( 
.A1(n_39),
.A2(n_41),
.B(n_45),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_41),
.B(n_49),
.Y(n_48)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_41),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_41),
.B(n_48),
.Y(n_228)
);

CKINVDCx16_ASAP7_75t_R g44 ( 
.A(n_42),
.Y(n_44)
);

OAI22xp33_ASAP7_75t_L g57 ( 
.A1(n_42),
.A2(n_44),
.B1(n_58),
.B2(n_59),
.Y(n_57)
);

INVxp67_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

OAI21xp5_ASAP7_75t_L g109 ( 
.A1(n_46),
.A2(n_71),
.B(n_73),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_47),
.B(n_48),
.Y(n_46)
);

CKINVDCx14_ASAP7_75t_R g72 ( 
.A(n_47),
.Y(n_72)
);

INVxp67_ASAP7_75t_L g70 ( 
.A(n_48),
.Y(n_70)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_53),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_SL g53 ( 
.A(n_54),
.B(n_64),
.Y(n_53)
);

INVxp33_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_55),
.B(n_133),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g55 ( 
.A(n_56),
.B(n_60),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_56),
.A2(n_60),
.B1(n_64),
.B2(n_68),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_56),
.B(n_87),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_56),
.A2(n_60),
.B1(n_87),
.B2(n_105),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_57),
.B(n_60),
.Y(n_56)
);

INVx11_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

OAI21xp5_ASAP7_75t_L g84 ( 
.A1(n_60),
.A2(n_68),
.B(n_85),
.Y(n_84)
);

INVxp67_ASAP7_75t_L g139 ( 
.A(n_60),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_SL g195 ( 
.A(n_61),
.B(n_196),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_62),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_62),
.B(n_81),
.Y(n_80)
);

INVx11_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

AOI21xp5_ASAP7_75t_L g97 ( 
.A1(n_66),
.A2(n_67),
.B(n_69),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_67),
.B(n_69),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_69),
.A2(n_106),
.B1(n_119),
.B2(n_120),
.Y(n_118)
);

CKINVDCx16_ASAP7_75t_R g120 ( 
.A(n_69),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_69),
.B(n_153),
.C(n_154),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_69),
.A2(n_120),
.B1(n_170),
.B2(n_172),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_70),
.A2(n_71),
.B1(n_72),
.B2(n_73),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g227 ( 
.A(n_72),
.B(n_228),
.Y(n_227)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

AOI21xp33_ASAP7_75t_L g75 ( 
.A1(n_76),
.A2(n_83),
.B(n_88),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_76),
.B(n_84),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_76),
.A2(n_88),
.B1(n_89),
.B2(n_96),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_76),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_76),
.A2(n_84),
.B1(n_96),
.B2(n_241),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_77),
.B(n_78),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_77),
.A2(n_80),
.B1(n_102),
.B2(n_103),
.Y(n_101)
);

INVxp33_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_79),
.B(n_145),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_80),
.B(n_81),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_80),
.A2(n_103),
.B1(n_126),
.B2(n_127),
.Y(n_125)
);

INVxp67_ASAP7_75t_L g144 ( 
.A(n_80),
.Y(n_144)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

XOR2xp5_ASAP7_75t_L g94 ( 
.A(n_83),
.B(n_95),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_84),
.Y(n_241)
);

INVxp67_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

AOI21xp5_ASAP7_75t_L g137 ( 
.A1(n_86),
.A2(n_138),
.B(n_139),
.Y(n_137)
);

INVxp67_ASAP7_75t_L g133 ( 
.A(n_87),
.Y(n_133)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_91),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_97),
.C(n_98),
.Y(n_93)
);

XOR2xp5_ASAP7_75t_L g248 ( 
.A(n_94),
.B(n_97),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_98),
.A2(n_99),
.B1(n_247),
.B2(n_248),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_99),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_100),
.B(n_106),
.C(n_108),
.Y(n_99)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_100),
.B(n_238),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_101),
.B(n_104),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_101),
.A2(n_104),
.B1(n_177),
.B2(n_222),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_101),
.Y(n_222)
);

OAI21xp5_ASAP7_75t_SL g141 ( 
.A1(n_102),
.A2(n_142),
.B(n_143),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_L g153 ( 
.A1(n_103),
.A2(n_126),
.B(n_143),
.Y(n_153)
);

INVx11_ASAP7_75t_L g198 ( 
.A(n_103),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_104),
.A2(n_175),
.B1(n_176),
.B2(n_177),
.Y(n_174)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_104),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_L g185 ( 
.A1(n_104),
.A2(n_177),
.B1(n_186),
.B2(n_187),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_104),
.B(n_125),
.C(n_187),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_104),
.B(n_168),
.C(n_176),
.Y(n_211)
);

INVxp67_ASAP7_75t_L g138 ( 
.A(n_105),
.Y(n_138)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_106),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_106),
.B(n_120),
.C(n_121),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_106),
.A2(n_108),
.B1(n_109),
.B2(n_119),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_108),
.A2(n_109),
.B1(n_131),
.B2(n_132),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_108),
.B(n_137),
.C(n_161),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_108),
.A2(n_109),
.B1(n_136),
.B2(n_137),
.Y(n_207)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

AOI21xp5_ASAP7_75t_L g112 ( 
.A1(n_113),
.A2(n_244),
.B(n_249),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_SL g113 ( 
.A1(n_114),
.A2(n_232),
.B(n_243),
.Y(n_113)
);

O2A1O1Ixp33_ASAP7_75t_SL g114 ( 
.A1(n_115),
.A2(n_156),
.B(n_216),
.C(n_231),
.Y(n_114)
);

AND2x2_ASAP7_75t_L g115 ( 
.A(n_116),
.B(n_146),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_116),
.B(n_146),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g116 ( 
.A(n_117),
.B(n_128),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_117),
.B(n_129),
.C(n_135),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_SL g117 ( 
.A(n_118),
.B(n_121),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_122),
.B(n_125),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_122),
.A2(n_123),
.B1(n_125),
.B2(n_151),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_123),
.Y(n_122)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_125),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_125),
.A2(n_151),
.B1(n_185),
.B2(n_188),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_125),
.B(n_200),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_125),
.B(n_200),
.Y(n_201)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_127),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_129),
.A2(n_130),
.B1(n_134),
.B2(n_135),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_130),
.Y(n_129)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_135),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_136),
.A2(n_137),
.B1(n_140),
.B2(n_141),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_136),
.A2(n_137),
.B1(n_182),
.B2(n_192),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_136),
.B(n_141),
.Y(n_224)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_SL g181 ( 
.A(n_137),
.B(n_182),
.Y(n_181)
);

CKINVDCx16_ASAP7_75t_R g140 ( 
.A(n_141),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_145),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_150),
.C(n_152),
.Y(n_146)
);

XOR2xp5_ASAP7_75t_L g212 ( 
.A(n_147),
.B(n_213),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_148),
.Y(n_149)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_150),
.B(n_152),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_153),
.A2(n_154),
.B1(n_155),
.B2(n_171),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_153),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_153),
.B(n_195),
.Y(n_194)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_SL g156 ( 
.A(n_157),
.B(n_215),
.Y(n_156)
);

AOI21xp5_ASAP7_75t_L g157 ( 
.A1(n_158),
.A2(n_210),
.B(n_214),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_L g158 ( 
.A1(n_159),
.A2(n_178),
.B(n_209),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_167),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_160),
.B(n_167),
.Y(n_209)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_161),
.B(n_207),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_162),
.A2(n_164),
.B1(n_165),
.B2(n_166),
.Y(n_161)
);

CKINVDCx16_ASAP7_75t_R g166 ( 
.A(n_162),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_164),
.B(n_166),
.Y(n_175)
);

CKINVDCx16_ASAP7_75t_R g164 ( 
.A(n_165),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_168),
.A2(n_169),
.B1(n_173),
.B2(n_174),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_170),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_171),
.B(n_191),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_SL g202 ( 
.A(n_171),
.B(n_191),
.Y(n_202)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_175),
.Y(n_176)
);

AOI21xp5_ASAP7_75t_L g178 ( 
.A1(n_179),
.A2(n_204),
.B(n_208),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_L g179 ( 
.A1(n_180),
.A2(n_189),
.B(n_203),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_184),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_181),
.B(n_184),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_182),
.Y(n_192)
);

CKINVDCx16_ASAP7_75t_R g188 ( 
.A(n_185),
.Y(n_188)
);

CKINVDCx16_ASAP7_75t_R g187 ( 
.A(n_186),
.Y(n_187)
);

AOI21xp5_ASAP7_75t_L g189 ( 
.A1(n_190),
.A2(n_193),
.B(n_202),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_L g193 ( 
.A1(n_194),
.A2(n_199),
.B(n_201),
.Y(n_193)
);

INVx5_ASAP7_75t_SL g197 ( 
.A(n_198),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_205),
.B(n_206),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_205),
.B(n_206),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_211),
.B(n_212),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_211),
.B(n_212),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_217),
.B(n_218),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_SL g231 ( 
.A(n_217),
.B(n_218),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_219),
.A2(n_220),
.B1(n_229),
.B2(n_230),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_221),
.B(n_223),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_221),
.B(n_223),
.C(n_230),
.Y(n_233)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_224),
.B(n_225),
.Y(n_223)
);

CKINVDCx14_ASAP7_75t_R g226 ( 
.A(n_227),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_229),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_233),
.B(n_234),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_SL g243 ( 
.A(n_233),
.B(n_234),
.Y(n_243)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_235),
.B(n_242),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_236),
.A2(n_237),
.B1(n_239),
.B2(n_240),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_236),
.B(n_240),
.C(n_242),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_237),
.Y(n_236)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_245),
.B(n_246),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_SL g249 ( 
.A(n_245),
.B(n_246),
.Y(n_249)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);


endmodule