module fake_jpeg_16385_n_322 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_322);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_322;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_4),
.Y(n_15)
);

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

BUFx6f_ASAP7_75t_SL g17 ( 
.A(n_14),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

INVx11_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_3),
.Y(n_24)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

BUFx10_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_1),
.Y(n_27)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

BUFx10_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_0),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_13),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_18),
.Y(n_32)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_32),
.Y(n_48)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_17),
.Y(n_33)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_33),
.Y(n_45)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_26),
.Y(n_34)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_34),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_18),
.Y(n_35)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_25),
.B(n_1),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_36),
.B(n_37),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_24),
.B(n_30),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_26),
.Y(n_38)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_38),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_26),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_39),
.B(n_40),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g40 ( 
.A(n_20),
.B(n_1),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_SL g41 ( 
.A1(n_33),
.A2(n_17),
.B1(n_25),
.B2(n_28),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_41),
.A2(n_28),
.B1(n_42),
.B2(n_45),
.Y(n_62)
);

INVx5_ASAP7_75t_L g42 ( 
.A(n_33),
.Y(n_42)
);

INVx5_ASAP7_75t_L g78 ( 
.A(n_42),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g43 ( 
.A1(n_36),
.A2(n_17),
.B1(n_25),
.B2(n_28),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_L g63 ( 
.A1(n_43),
.A2(n_54),
.B1(n_22),
.B2(n_20),
.Y(n_63)
);

BUFx2_ASAP7_75t_L g44 ( 
.A(n_32),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_44),
.Y(n_60)
);

INVx8_ASAP7_75t_L g49 ( 
.A(n_32),
.Y(n_49)
);

INVx3_ASAP7_75t_SL g70 ( 
.A(n_49),
.Y(n_70)
);

MAJIxp5_ASAP7_75t_L g52 ( 
.A(n_36),
.B(n_16),
.C(n_29),
.Y(n_52)
);

AND2x2_ASAP7_75t_L g73 ( 
.A(n_52),
.B(n_38),
.Y(n_73)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_32),
.Y(n_53)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_53),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_38),
.A2(n_22),
.B1(n_25),
.B2(n_28),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_37),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_55),
.B(n_40),
.Y(n_67)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_42),
.Y(n_58)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_58),
.Y(n_93)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_51),
.Y(n_59)
);

BUFx2_ASAP7_75t_L g106 ( 
.A(n_59),
.Y(n_106)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_51),
.Y(n_61)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_61),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g105 ( 
.A(n_62),
.B(n_63),
.Y(n_105)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_48),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_64),
.B(n_67),
.Y(n_91)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_46),
.Y(n_65)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_65),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_53),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_66),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_53),
.Y(n_68)
);

INVx11_ASAP7_75t_L g107 ( 
.A(n_68),
.Y(n_107)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_45),
.Y(n_69)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_69),
.Y(n_102)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_45),
.Y(n_71)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_71),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_L g72 ( 
.A1(n_50),
.A2(n_22),
.B1(n_55),
.B2(n_52),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_72),
.A2(n_79),
.B1(n_82),
.B2(n_20),
.Y(n_88)
);

XNOR2x1_ASAP7_75t_SL g109 ( 
.A(n_73),
.B(n_41),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_50),
.B(n_31),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_74),
.B(n_75),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_56),
.B(n_31),
.Y(n_75)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_48),
.Y(n_76)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_76),
.Y(n_104)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_48),
.Y(n_77)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_77),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_46),
.A2(n_22),
.B1(n_31),
.B2(n_30),
.Y(n_79)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_44),
.Y(n_80)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_80),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_56),
.B(n_26),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_81),
.B(n_83),
.Y(n_112)
);

OAI22xp33_ASAP7_75t_L g82 ( 
.A1(n_49),
.A2(n_35),
.B1(n_18),
.B2(n_21),
.Y(n_82)
);

CKINVDCx16_ASAP7_75t_R g83 ( 
.A(n_54),
.Y(n_83)
);

INVx13_ASAP7_75t_L g84 ( 
.A(n_65),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_84),
.B(n_86),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_66),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_88),
.A2(n_57),
.B1(n_23),
.B2(n_71),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_73),
.B(n_52),
.Y(n_89)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_89),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_78),
.A2(n_46),
.B1(n_49),
.B2(n_47),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_90),
.A2(n_100),
.B1(n_70),
.B2(n_47),
.Y(n_118)
);

A2O1A1Ixp33_ASAP7_75t_L g92 ( 
.A1(n_73),
.A2(n_43),
.B(n_30),
.C(n_27),
.Y(n_92)
);

XOR2x1_ASAP7_75t_L g121 ( 
.A(n_92),
.B(n_97),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_59),
.B(n_43),
.Y(n_95)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_95),
.Y(n_123)
);

AOI21xp33_ASAP7_75t_L g97 ( 
.A1(n_62),
.A2(n_24),
.B(n_27),
.Y(n_97)
);

CKINVDCx14_ASAP7_75t_R g98 ( 
.A(n_58),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_98),
.B(n_111),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_61),
.B(n_23),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_L g130 ( 
.A1(n_99),
.A2(n_27),
.B(n_24),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_78),
.A2(n_49),
.B1(n_47),
.B2(n_23),
.Y(n_100)
);

AND2x2_ASAP7_75t_L g117 ( 
.A(n_109),
.B(n_82),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_70),
.B(n_41),
.C(n_39),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_110),
.B(n_34),
.C(n_35),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_68),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_104),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_113),
.B(n_132),
.Y(n_144)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_85),
.Y(n_114)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_114),
.Y(n_146)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_85),
.Y(n_115)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_115),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_SL g162 ( 
.A1(n_117),
.A2(n_128),
.B(n_131),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_118),
.A2(n_122),
.B1(n_57),
.B2(n_99),
.Y(n_147)
);

HB1xp67_ASAP7_75t_L g119 ( 
.A(n_93),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_119),
.B(n_136),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_124),
.B(n_129),
.C(n_93),
.Y(n_142)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_101),
.Y(n_125)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_125),
.Y(n_150)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_94),
.Y(n_126)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_126),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_109),
.A2(n_89),
.B1(n_105),
.B2(n_95),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_127),
.A2(n_91),
.B1(n_87),
.B2(n_96),
.Y(n_152)
);

AND2x2_ASAP7_75t_L g128 ( 
.A(n_110),
.B(n_60),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_112),
.B(n_39),
.C(n_34),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_L g157 ( 
.A1(n_130),
.A2(n_104),
.B(n_111),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_SL g131 ( 
.A1(n_105),
.A2(n_69),
.B(n_16),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_102),
.Y(n_132)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_102),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_133),
.B(n_135),
.Y(n_160)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_101),
.Y(n_134)
);

INVxp67_ASAP7_75t_L g153 ( 
.A(n_134),
.Y(n_153)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_103),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_103),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_96),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_137),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g138 ( 
.A(n_108),
.Y(n_138)
);

INVx3_ASAP7_75t_L g161 ( 
.A(n_138),
.Y(n_161)
);

CKINVDCx14_ASAP7_75t_R g140 ( 
.A(n_139),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_140),
.B(n_142),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_117),
.A2(n_105),
.B1(n_112),
.B2(n_92),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_141),
.A2(n_147),
.B1(n_163),
.B2(n_164),
.Y(n_183)
);

OAI32xp33_ASAP7_75t_L g143 ( 
.A1(n_121),
.A2(n_120),
.A3(n_127),
.B1(n_123),
.B2(n_117),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_143),
.B(n_134),
.Y(n_175)
);

INVx2_ASAP7_75t_SL g145 ( 
.A(n_126),
.Y(n_145)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_145),
.Y(n_177)
);

FAx1_ASAP7_75t_SL g151 ( 
.A(n_121),
.B(n_87),
.CI(n_91),
.CON(n_151),
.SN(n_151)
);

NOR2xp33_ASAP7_75t_SL g191 ( 
.A(n_151),
.B(n_157),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_152),
.B(n_154),
.Y(n_178)
);

INVxp67_ASAP7_75t_L g154 ( 
.A(n_116),
.Y(n_154)
);

BUFx24_ASAP7_75t_SL g155 ( 
.A(n_120),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_155),
.B(n_166),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_L g158 ( 
.A1(n_128),
.A2(n_86),
.B(n_106),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_L g171 ( 
.A1(n_158),
.A2(n_159),
.B(n_129),
.Y(n_171)
);

AOI21xp5_ASAP7_75t_L g159 ( 
.A1(n_131),
.A2(n_94),
.B(n_2),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_123),
.A2(n_107),
.B1(n_77),
.B2(n_76),
.Y(n_163)
);

AOI22xp33_ASAP7_75t_SL g164 ( 
.A1(n_115),
.A2(n_107),
.B1(n_80),
.B2(n_84),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_124),
.A2(n_35),
.B1(n_44),
.B2(n_106),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_165),
.A2(n_167),
.B1(n_170),
.B2(n_161),
.Y(n_185)
);

INVxp67_ASAP7_75t_L g166 ( 
.A(n_125),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_128),
.A2(n_84),
.B1(n_106),
.B2(n_44),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_133),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_168),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_122),
.A2(n_108),
.B1(n_12),
.B2(n_13),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_L g218 ( 
.A(n_171),
.B(n_172),
.Y(n_218)
);

OAI21xp5_ASAP7_75t_L g172 ( 
.A1(n_159),
.A2(n_130),
.B(n_135),
.Y(n_172)
);

INVx1_ASAP7_75t_SL g173 ( 
.A(n_160),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_173),
.B(n_176),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_175),
.A2(n_181),
.B1(n_184),
.B2(n_190),
.Y(n_205)
);

INVxp67_ASAP7_75t_L g176 ( 
.A(n_169),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_152),
.B(n_18),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_179),
.B(n_180),
.Y(n_222)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_145),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_154),
.A2(n_138),
.B1(n_21),
.B2(n_19),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_141),
.A2(n_21),
.B1(n_19),
.B2(n_15),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_185),
.B(n_195),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_143),
.B(n_18),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_186),
.B(n_187),
.Y(n_225)
);

INVxp67_ASAP7_75t_L g187 ( 
.A(n_144),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_157),
.B(n_21),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_188),
.B(n_189),
.Y(n_226)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_145),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_158),
.A2(n_108),
.B1(n_19),
.B2(n_15),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_162),
.A2(n_15),
.B1(n_19),
.B2(n_10),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_192),
.A2(n_200),
.B1(n_170),
.B2(n_149),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_151),
.B(n_15),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_193),
.B(n_194),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_150),
.Y(n_194)
);

INVx1_ASAP7_75t_SL g195 ( 
.A(n_153),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_150),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_196),
.Y(n_204)
);

CKINVDCx16_ASAP7_75t_R g198 ( 
.A(n_148),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_198),
.B(n_201),
.Y(n_215)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_148),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_199),
.Y(n_207)
);

AOI21xp5_ASAP7_75t_L g200 ( 
.A1(n_162),
.A2(n_1),
.B(n_2),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_156),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_146),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_202),
.B(n_16),
.Y(n_228)
);

OAI21xp5_ASAP7_75t_L g203 ( 
.A1(n_142),
.A2(n_2),
.B(n_3),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_203),
.B(n_5),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_174),
.B(n_151),
.C(n_167),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_206),
.B(n_208),
.C(n_220),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_171),
.B(n_165),
.C(n_156),
.Y(n_208)
);

CKINVDCx14_ASAP7_75t_R g245 ( 
.A(n_211),
.Y(n_245)
);

INVxp67_ASAP7_75t_L g212 ( 
.A(n_181),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_212),
.B(n_224),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_183),
.A2(n_166),
.B1(n_153),
.B2(n_161),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_213),
.A2(n_216),
.B1(n_173),
.B2(n_187),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_178),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_216)
);

OAI22x1_ASAP7_75t_L g217 ( 
.A1(n_192),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_217),
.A2(n_212),
.B1(n_224),
.B2(n_200),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_182),
.B(n_202),
.Y(n_219)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_219),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_175),
.B(n_16),
.C(n_29),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_191),
.B(n_16),
.C(n_29),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_221),
.B(n_227),
.C(n_196),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_SL g244 ( 
.A(n_223),
.B(n_203),
.Y(n_244)
);

INVxp67_ASAP7_75t_L g224 ( 
.A(n_190),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_193),
.B(n_16),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_228),
.B(n_189),
.Y(n_240)
);

AND2x2_ASAP7_75t_L g229 ( 
.A(n_218),
.B(n_188),
.Y(n_229)
);

CKINVDCx16_ASAP7_75t_R g252 ( 
.A(n_229),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_230),
.A2(n_234),
.B1(n_235),
.B2(n_241),
.Y(n_256)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_215),
.Y(n_231)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_231),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g232 ( 
.A(n_218),
.B(n_186),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_232),
.B(n_239),
.C(n_249),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_216),
.B(n_182),
.Y(n_233)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_233),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_210),
.A2(n_179),
.B1(n_194),
.B2(n_185),
.Y(n_235)
);

BUFx2_ASAP7_75t_L g238 ( 
.A(n_209),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_238),
.Y(n_257)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_240),
.Y(n_260)
);

OAI21xp5_ASAP7_75t_L g241 ( 
.A1(n_225),
.A2(n_191),
.B(n_172),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_207),
.B(n_176),
.Y(n_242)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_242),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_222),
.B(n_180),
.Y(n_243)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_243),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_SL g264 ( 
.A(n_244),
.B(n_223),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_214),
.Y(n_246)
);

BUFx24_ASAP7_75t_SL g250 ( 
.A(n_246),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_208),
.A2(n_195),
.B1(n_199),
.B2(n_201),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_248),
.A2(n_220),
.B1(n_217),
.B2(n_177),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_206),
.B(n_184),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_236),
.B(n_213),
.C(n_226),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_254),
.B(n_255),
.C(n_261),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_236),
.B(n_221),
.C(n_204),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_SL g281 ( 
.A(n_258),
.B(n_16),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_248),
.B(n_227),
.C(n_177),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_239),
.B(n_205),
.C(n_211),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_262),
.B(n_266),
.C(n_230),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_264),
.B(n_234),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_249),
.B(n_205),
.C(n_197),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_254),
.B(n_247),
.C(n_232),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_267),
.B(n_274),
.C(n_279),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_259),
.B(n_231),
.Y(n_268)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_268),
.Y(n_290)
);

HB1xp67_ASAP7_75t_L g269 ( 
.A(n_265),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_L g289 ( 
.A(n_269),
.B(n_273),
.Y(n_289)
);

XOR2xp5_ASAP7_75t_L g270 ( 
.A(n_253),
.B(n_229),
.Y(n_270)
);

XOR2xp5_ASAP7_75t_L g284 ( 
.A(n_270),
.B(n_278),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_260),
.B(n_241),
.Y(n_271)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_271),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_257),
.B(n_235),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g293 ( 
.A(n_275),
.B(n_11),
.Y(n_293)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_251),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_276),
.A2(n_277),
.B1(n_281),
.B2(n_5),
.Y(n_287)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_263),
.Y(n_277)
);

XOR2xp5_ASAP7_75t_L g278 ( 
.A(n_253),
.B(n_229),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_262),
.B(n_245),
.C(n_237),
.Y(n_279)
);

XOR2xp5_ASAP7_75t_L g280 ( 
.A(n_256),
.B(n_238),
.Y(n_280)
);

XOR2xp5_ASAP7_75t_L g285 ( 
.A(n_280),
.B(n_264),
.Y(n_285)
);

OAI21x1_ASAP7_75t_SL g282 ( 
.A1(n_280),
.A2(n_250),
.B(n_261),
.Y(n_282)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_282),
.Y(n_297)
);

AOI22xp33_ASAP7_75t_SL g283 ( 
.A1(n_270),
.A2(n_252),
.B1(n_255),
.B2(n_266),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_283),
.B(n_293),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_285),
.B(n_11),
.C(n_7),
.Y(n_304)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_287),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_272),
.B(n_29),
.C(n_26),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_288),
.B(n_291),
.C(n_294),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_274),
.B(n_29),
.C(n_26),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_272),
.B(n_29),
.C(n_26),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_SL g295 ( 
.A(n_292),
.B(n_278),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g307 ( 
.A(n_295),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_290),
.B(n_289),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_SL g308 ( 
.A(n_299),
.B(n_300),
.Y(n_308)
);

HB1xp67_ASAP7_75t_L g300 ( 
.A(n_286),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_288),
.B(n_29),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_301),
.B(n_303),
.C(n_304),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_284),
.B(n_10),
.C(n_7),
.Y(n_303)
);

INVx6_ASAP7_75t_L g305 ( 
.A(n_299),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_305),
.B(n_311),
.Y(n_313)
);

XOR2xp5_ASAP7_75t_L g306 ( 
.A(n_298),
.B(n_284),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_306),
.B(n_310),
.C(n_9),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_297),
.B(n_285),
.C(n_283),
.Y(n_310)
);

NAND3xp33_ASAP7_75t_L g311 ( 
.A(n_302),
.B(n_8),
.C(n_9),
.Y(n_311)
);

AOI21xp5_ASAP7_75t_L g312 ( 
.A1(n_308),
.A2(n_296),
.B(n_8),
.Y(n_312)
);

OAI21xp5_ASAP7_75t_L g315 ( 
.A1(n_312),
.A2(n_314),
.B(n_311),
.Y(n_315)
);

AOI21xp5_ASAP7_75t_L g316 ( 
.A1(n_315),
.A2(n_313),
.B(n_306),
.Y(n_316)
);

AO221x1_ASAP7_75t_L g317 ( 
.A1(n_316),
.A2(n_305),
.B1(n_307),
.B2(n_309),
.C(n_12),
.Y(n_317)
);

OR2x2_ASAP7_75t_L g318 ( 
.A(n_317),
.B(n_9),
.Y(n_318)
);

OAI21xp5_ASAP7_75t_SL g319 ( 
.A1(n_318),
.A2(n_11),
.B(n_13),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_319),
.B(n_14),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_320),
.B(n_6),
.Y(n_321)
);

AOI21xp5_ASAP7_75t_L g322 ( 
.A1(n_321),
.A2(n_6),
.B(n_14),
.Y(n_322)
);


endmodule