module fake_jpeg_4658_n_138 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_138);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_138;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_11;
wire n_131;
wire n_56;
wire n_79;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

INVx1_ASAP7_75t_L g11 ( 
.A(n_5),
.Y(n_11)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_10),
.Y(n_12)
);

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_4),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_3),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_1),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_0),
.B(n_10),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

BUFx10_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

BUFx12_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_12),
.B(n_0),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_24),
.B(n_27),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_21),
.Y(n_25)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_25),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_21),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_26),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_12),
.B(n_0),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_28),
.B(n_29),
.Y(n_34)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_19),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_19),
.Y(n_30)
);

INVx5_ASAP7_75t_L g45 ( 
.A(n_30),
.Y(n_45)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_20),
.Y(n_31)
);

CKINVDCx16_ASAP7_75t_R g35 ( 
.A(n_31),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_32),
.Y(n_40)
);

AND2x2_ASAP7_75t_L g37 ( 
.A(n_29),
.B(n_15),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_37),
.B(n_38),
.Y(n_48)
);

AND2x2_ASAP7_75t_L g38 ( 
.A(n_30),
.B(n_15),
.Y(n_38)
);

OAI22xp33_ASAP7_75t_L g41 ( 
.A1(n_32),
.A2(n_22),
.B1(n_16),
.B2(n_13),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_L g49 ( 
.A1(n_41),
.A2(n_14),
.B1(n_11),
.B2(n_18),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_31),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_42),
.B(n_43),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_25),
.Y(n_43)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_27),
.Y(n_44)
);

HB1xp67_ASAP7_75t_L g56 ( 
.A(n_44),
.Y(n_56)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_45),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_46),
.B(n_53),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_42),
.B(n_22),
.Y(n_47)
);

XNOR2xp5_ASAP7_75t_L g67 ( 
.A(n_47),
.B(n_50),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_49),
.A2(n_57),
.B1(n_39),
.B2(n_17),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_35),
.B(n_20),
.Y(n_50)
);

A2O1A1Ixp33_ASAP7_75t_L g51 ( 
.A1(n_34),
.A2(n_17),
.B(n_14),
.C(n_20),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_51),
.B(n_52),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_35),
.B(n_20),
.Y(n_52)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_45),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_54),
.B(n_36),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g57 ( 
.A1(n_37),
.A2(n_32),
.B1(n_18),
.B2(n_11),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_47),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_58),
.B(n_59),
.Y(n_71)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_56),
.Y(n_59)
);

MAJIxp5_ASAP7_75t_L g60 ( 
.A(n_50),
.B(n_33),
.C(n_38),
.Y(n_60)
);

OAI21xp5_ASAP7_75t_SL g79 ( 
.A1(n_60),
.A2(n_63),
.B(n_68),
.Y(n_79)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_55),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_62),
.B(n_64),
.Y(n_76)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_52),
.Y(n_64)
);

OAI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_57),
.A2(n_38),
.B1(n_37),
.B2(n_41),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_65),
.A2(n_70),
.B1(n_20),
.B2(n_16),
.Y(n_81)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_49),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_SL g78 ( 
.A(n_66),
.B(n_16),
.Y(n_78)
);

AO22x1_ASAP7_75t_L g68 ( 
.A1(n_48),
.A2(n_39),
.B1(n_40),
.B2(n_44),
.Y(n_68)
);

AO22x1_ASAP7_75t_L g75 ( 
.A1(n_68),
.A2(n_54),
.B1(n_36),
.B2(n_43),
.Y(n_75)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_69),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_67),
.B(n_48),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_72),
.B(n_77),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_61),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_73),
.B(n_80),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_58),
.A2(n_54),
.B1(n_46),
.B2(n_53),
.Y(n_74)
);

INVxp67_ASAP7_75t_L g83 ( 
.A(n_74),
.Y(n_83)
);

OA21x2_ASAP7_75t_L g88 ( 
.A1(n_75),
.A2(n_23),
.B(n_2),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_67),
.B(n_51),
.Y(n_77)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_78),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_79),
.B(n_26),
.C(n_23),
.Y(n_87)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_59),
.Y(n_80)
);

AO21x1_ASAP7_75t_L g85 ( 
.A1(n_81),
.A2(n_68),
.B(n_62),
.Y(n_85)
);

XOR2xp5_ASAP7_75t_L g84 ( 
.A(n_72),
.B(n_60),
.Y(n_84)
);

XOR2xp5_ASAP7_75t_L g98 ( 
.A(n_84),
.B(n_87),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_85),
.B(n_86),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_SL g86 ( 
.A(n_76),
.B(n_70),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_88),
.A2(n_75),
.B1(n_82),
.B2(n_80),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g91 ( 
.A(n_71),
.Y(n_91)
);

CKINVDCx14_ASAP7_75t_R g96 ( 
.A(n_91),
.Y(n_96)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_74),
.Y(n_92)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_92),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_73),
.B(n_9),
.Y(n_93)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_93),
.Y(n_105)
);

AOI21xp5_ASAP7_75t_L g95 ( 
.A1(n_87),
.A2(n_79),
.B(n_75),
.Y(n_95)
);

NOR3xp33_ASAP7_75t_L g109 ( 
.A(n_95),
.B(n_102),
.C(n_82),
.Y(n_109)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_89),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_97),
.B(n_99),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_94),
.B(n_77),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_100),
.B(n_101),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_88),
.Y(n_101)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_94),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_104),
.A2(n_83),
.B1(n_85),
.B2(n_90),
.Y(n_106)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_106),
.Y(n_121)
);

XOR2xp5_ASAP7_75t_L g107 ( 
.A(n_98),
.B(n_84),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_107),
.B(n_111),
.C(n_103),
.Y(n_116)
);

NAND3xp33_ASAP7_75t_L g108 ( 
.A(n_95),
.B(n_91),
.C(n_88),
.Y(n_108)
);

XNOR2xp5_ASAP7_75t_L g117 ( 
.A(n_108),
.B(n_23),
.Y(n_117)
);

AOI21xp5_ASAP7_75t_L g119 ( 
.A1(n_109),
.A2(n_113),
.B(n_1),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_98),
.B(n_83),
.C(n_23),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_110),
.B(n_96),
.C(n_97),
.Y(n_115)
);

XOR2xp5_ASAP7_75t_L g111 ( 
.A(n_99),
.B(n_102),
.Y(n_111)
);

INVxp67_ASAP7_75t_L g113 ( 
.A(n_100),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_115),
.B(n_116),
.C(n_118),
.Y(n_127)
);

NOR3xp33_ASAP7_75t_L g126 ( 
.A(n_117),
.B(n_119),
.C(n_8),
.Y(n_126)
);

XNOR2xp5_ASAP7_75t_L g118 ( 
.A(n_114),
.B(n_105),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_108),
.B(n_1),
.C(n_3),
.Y(n_120)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_120),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_121),
.A2(n_113),
.B1(n_112),
.B2(n_6),
.Y(n_123)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_123),
.Y(n_128)
);

O2A1O1Ixp33_ASAP7_75t_L g124 ( 
.A1(n_115),
.A2(n_4),
.B(n_5),
.C(n_6),
.Y(n_124)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_124),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_118),
.B(n_4),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_L g129 ( 
.A1(n_125),
.A2(n_126),
.B(n_8),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_129),
.B(n_7),
.Y(n_134)
);

XNOR2xp5_ASAP7_75t_L g130 ( 
.A(n_127),
.B(n_6),
.Y(n_130)
);

XOR2xp5_ASAP7_75t_L g132 ( 
.A(n_130),
.B(n_125),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_132),
.B(n_133),
.Y(n_135)
);

NOR3xp33_ASAP7_75t_SL g133 ( 
.A(n_131),
.B(n_128),
.C(n_122),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_134),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_L g137 ( 
.A1(n_135),
.A2(n_133),
.B(n_130),
.Y(n_137)
);

XOR2xp5_ASAP7_75t_L g138 ( 
.A(n_137),
.B(n_136),
.Y(n_138)
);


endmodule