module fake_netlist_1_11920_n_610 (n_53, n_67, n_45, n_20, n_2, n_38, n_44, n_64, n_54, n_62, n_36, n_47, n_37, n_69, n_34, n_5, n_23, n_8, n_28, n_31, n_22, n_46, n_48, n_58, n_57, n_11, n_25, n_16, n_26, n_13, n_30, n_33, n_50, n_52, n_49, n_59, n_73, n_3, n_18, n_60, n_66, n_32, n_0, n_41, n_1, n_35, n_55, n_65, n_12, n_9, n_70, n_17, n_63, n_14, n_10, n_15, n_56, n_71, n_42, n_24, n_19, n_61, n_21, n_6, n_4, n_74, n_72, n_51, n_29, n_43, n_7, n_68, n_40, n_27, n_39, n_610);
input n_53;
input n_67;
input n_45;
input n_20;
input n_2;
input n_38;
input n_44;
input n_64;
input n_54;
input n_62;
input n_36;
input n_47;
input n_37;
input n_69;
input n_34;
input n_5;
input n_23;
input n_8;
input n_28;
input n_31;
input n_22;
input n_46;
input n_48;
input n_58;
input n_57;
input n_11;
input n_25;
input n_16;
input n_26;
input n_13;
input n_30;
input n_33;
input n_50;
input n_52;
input n_49;
input n_59;
input n_73;
input n_3;
input n_18;
input n_60;
input n_66;
input n_32;
input n_0;
input n_41;
input n_1;
input n_35;
input n_55;
input n_65;
input n_12;
input n_9;
input n_70;
input n_17;
input n_63;
input n_14;
input n_10;
input n_15;
input n_56;
input n_71;
input n_42;
input n_24;
input n_19;
input n_61;
input n_21;
input n_6;
input n_4;
input n_74;
input n_72;
input n_51;
input n_29;
input n_43;
input n_7;
input n_68;
input n_40;
input n_27;
input n_39;
output n_610;
wire n_117;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_154;
wire n_328;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_532;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_586;
wire n_244;
wire n_540;
wire n_563;
wire n_141;
wire n_119;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_593;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_367;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_108;
wire n_91;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_77;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_172;
wire n_329;
wire n_251;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_271;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_446;
wire n_423;
wire n_342;
wire n_420;
wire n_370;
wire n_589;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_357;
wire n_90;
wire n_245;
wire n_260;
wire n_78;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_208;
wire n_200;
wire n_573;
wire n_126;
wire n_178;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_75;
wire n_376;
wire n_552;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_76;
wire n_520;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_438;
wire n_134;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_583;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_84;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_444;
wire n_176;
wire n_521;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_132;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g75 ( .A(n_20), .Y(n_75) );
INVx1_ASAP7_75t_L g76 ( .A(n_53), .Y(n_76) );
BUFx2_ASAP7_75t_SL g77 ( .A(n_18), .Y(n_77) );
INVxp33_ASAP7_75t_L g78 ( .A(n_55), .Y(n_78) );
INVx1_ASAP7_75t_L g79 ( .A(n_4), .Y(n_79) );
INVx1_ASAP7_75t_L g80 ( .A(n_9), .Y(n_80) );
INVx1_ASAP7_75t_L g81 ( .A(n_34), .Y(n_81) );
INVx1_ASAP7_75t_L g82 ( .A(n_59), .Y(n_82) );
INVx1_ASAP7_75t_L g83 ( .A(n_11), .Y(n_83) );
INVx1_ASAP7_75t_L g84 ( .A(n_27), .Y(n_84) );
INVx1_ASAP7_75t_L g85 ( .A(n_58), .Y(n_85) );
INVxp33_ASAP7_75t_SL g86 ( .A(n_19), .Y(n_86) );
INVxp67_ASAP7_75t_SL g87 ( .A(n_11), .Y(n_87) );
NOR2xp67_ASAP7_75t_L g88 ( .A(n_7), .B(n_22), .Y(n_88) );
CKINVDCx5p33_ASAP7_75t_R g89 ( .A(n_15), .Y(n_89) );
INVxp67_ASAP7_75t_L g90 ( .A(n_2), .Y(n_90) );
CKINVDCx5p33_ASAP7_75t_R g91 ( .A(n_56), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_40), .Y(n_92) );
INVx1_ASAP7_75t_L g93 ( .A(n_26), .Y(n_93) );
INVx1_ASAP7_75t_L g94 ( .A(n_15), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_65), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_13), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_39), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_64), .Y(n_98) );
INVxp33_ASAP7_75t_SL g99 ( .A(n_62), .Y(n_99) );
NAND2xp5_ASAP7_75t_L g100 ( .A(n_73), .B(n_71), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_25), .Y(n_101) );
BUFx6f_ASAP7_75t_L g102 ( .A(n_63), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_10), .Y(n_103) );
INVx2_ASAP7_75t_L g104 ( .A(n_41), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_17), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_67), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_52), .Y(n_107) );
INVxp33_ASAP7_75t_SL g108 ( .A(n_70), .Y(n_108) );
INVxp67_ASAP7_75t_SL g109 ( .A(n_45), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_29), .Y(n_110) );
CKINVDCx20_ASAP7_75t_R g111 ( .A(n_22), .Y(n_111) );
CKINVDCx5p33_ASAP7_75t_R g112 ( .A(n_18), .Y(n_112) );
CKINVDCx16_ASAP7_75t_R g113 ( .A(n_25), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_50), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_60), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_43), .Y(n_116) );
INVxp67_ASAP7_75t_SL g117 ( .A(n_54), .Y(n_117) );
INVxp33_ASAP7_75t_SL g118 ( .A(n_30), .Y(n_118) );
INVx4_ASAP7_75t_R g119 ( .A(n_33), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_8), .Y(n_120) );
NOR2xp33_ASAP7_75t_L g121 ( .A(n_86), .B(n_0), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_76), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_76), .Y(n_123) );
CKINVDCx20_ASAP7_75t_R g124 ( .A(n_113), .Y(n_124) );
BUFx6f_ASAP7_75t_L g125 ( .A(n_102), .Y(n_125) );
CKINVDCx5p33_ASAP7_75t_R g126 ( .A(n_89), .Y(n_126) );
INVx2_ASAP7_75t_L g127 ( .A(n_102), .Y(n_127) );
INVx2_ASAP7_75t_L g128 ( .A(n_102), .Y(n_128) );
INVx2_ASAP7_75t_L g129 ( .A(n_102), .Y(n_129) );
NAND2xp5_ASAP7_75t_L g130 ( .A(n_90), .B(n_0), .Y(n_130) );
AND2x4_ASAP7_75t_L g131 ( .A(n_75), .B(n_1), .Y(n_131) );
BUFx6f_ASAP7_75t_L g132 ( .A(n_102), .Y(n_132) );
CKINVDCx20_ASAP7_75t_R g133 ( .A(n_111), .Y(n_133) );
BUFx6f_ASAP7_75t_L g134 ( .A(n_104), .Y(n_134) );
NAND2xp5_ASAP7_75t_L g135 ( .A(n_101), .B(n_1), .Y(n_135) );
CKINVDCx5p33_ASAP7_75t_R g136 ( .A(n_112), .Y(n_136) );
INVx1_ASAP7_75t_L g137 ( .A(n_81), .Y(n_137) );
INVx1_ASAP7_75t_L g138 ( .A(n_81), .Y(n_138) );
AND2x4_ASAP7_75t_L g139 ( .A(n_75), .B(n_2), .Y(n_139) );
CKINVDCx5p33_ASAP7_75t_R g140 ( .A(n_99), .Y(n_140) );
CKINVDCx5p33_ASAP7_75t_R g141 ( .A(n_108), .Y(n_141) );
INVx1_ASAP7_75t_L g142 ( .A(n_82), .Y(n_142) );
INVx1_ASAP7_75t_L g143 ( .A(n_82), .Y(n_143) );
CKINVDCx5p33_ASAP7_75t_R g144 ( .A(n_118), .Y(n_144) );
CKINVDCx20_ASAP7_75t_R g145 ( .A(n_77), .Y(n_145) );
INVx1_ASAP7_75t_L g146 ( .A(n_84), .Y(n_146) );
CKINVDCx20_ASAP7_75t_R g147 ( .A(n_77), .Y(n_147) );
CKINVDCx20_ASAP7_75t_R g148 ( .A(n_79), .Y(n_148) );
CKINVDCx5p33_ASAP7_75t_R g149 ( .A(n_91), .Y(n_149) );
INVx2_ASAP7_75t_L g150 ( .A(n_104), .Y(n_150) );
INVxp67_ASAP7_75t_L g151 ( .A(n_103), .Y(n_151) );
INVx1_ASAP7_75t_L g152 ( .A(n_84), .Y(n_152) );
HB1xp67_ASAP7_75t_L g153 ( .A(n_79), .Y(n_153) );
CKINVDCx20_ASAP7_75t_R g154 ( .A(n_80), .Y(n_154) );
AND2x2_ASAP7_75t_L g155 ( .A(n_78), .B(n_3), .Y(n_155) );
CKINVDCx5p33_ASAP7_75t_R g156 ( .A(n_98), .Y(n_156) );
INVx2_ASAP7_75t_L g157 ( .A(n_85), .Y(n_157) );
NAND2xp5_ASAP7_75t_L g158 ( .A(n_120), .B(n_3), .Y(n_158) );
NAND2xp5_ASAP7_75t_L g159 ( .A(n_85), .B(n_4), .Y(n_159) );
CKINVDCx5p33_ASAP7_75t_R g160 ( .A(n_109), .Y(n_160) );
INVx2_ASAP7_75t_L g161 ( .A(n_125), .Y(n_161) );
INVx2_ASAP7_75t_L g162 ( .A(n_125), .Y(n_162) );
BUFx2_ASAP7_75t_L g163 ( .A(n_126), .Y(n_163) );
BUFx4f_ASAP7_75t_L g164 ( .A(n_131), .Y(n_164) );
NAND2x1p5_ASAP7_75t_L g165 ( .A(n_131), .B(n_97), .Y(n_165) );
NAND2x1p5_ASAP7_75t_L g166 ( .A(n_131), .B(n_97), .Y(n_166) );
OAI221xp5_ASAP7_75t_L g167 ( .A1(n_151), .A2(n_80), .B1(n_94), .B2(n_96), .C(n_83), .Y(n_167) );
BUFx10_ASAP7_75t_L g168 ( .A(n_149), .Y(n_168) );
NAND3x1_ASAP7_75t_L g169 ( .A(n_121), .B(n_83), .C(n_94), .Y(n_169) );
NAND2xp5_ASAP7_75t_L g170 ( .A(n_122), .B(n_110), .Y(n_170) );
HB1xp67_ASAP7_75t_L g171 ( .A(n_136), .Y(n_171) );
NOR2x1_ASAP7_75t_L g172 ( .A(n_130), .B(n_107), .Y(n_172) );
OR2x2_ASAP7_75t_L g173 ( .A(n_153), .B(n_105), .Y(n_173) );
BUFx6f_ASAP7_75t_L g174 ( .A(n_125), .Y(n_174) );
BUFx6f_ASAP7_75t_L g175 ( .A(n_125), .Y(n_175) );
AOI22xp33_ASAP7_75t_L g176 ( .A1(n_131), .A2(n_105), .B1(n_96), .B2(n_87), .Y(n_176) );
INVx2_ASAP7_75t_L g177 ( .A(n_134), .Y(n_177) );
NAND2xp5_ASAP7_75t_SL g178 ( .A(n_156), .B(n_107), .Y(n_178) );
AO22x2_ASAP7_75t_L g179 ( .A1(n_139), .A2(n_106), .B1(n_93), .B2(n_116), .Y(n_179) );
INVx1_ASAP7_75t_L g180 ( .A(n_134), .Y(n_180) );
OAI22x1_ASAP7_75t_L g181 ( .A1(n_139), .A2(n_92), .B1(n_93), .B2(n_95), .Y(n_181) );
INVx1_ASAP7_75t_L g182 ( .A(n_134), .Y(n_182) );
INVx2_ASAP7_75t_L g183 ( .A(n_125), .Y(n_183) );
INVx8_ASAP7_75t_L g184 ( .A(n_139), .Y(n_184) );
BUFx6f_ASAP7_75t_L g185 ( .A(n_125), .Y(n_185) );
INVx2_ASAP7_75t_L g186 ( .A(n_132), .Y(n_186) );
BUFx4f_ASAP7_75t_L g187 ( .A(n_139), .Y(n_187) );
INVx2_ASAP7_75t_L g188 ( .A(n_134), .Y(n_188) );
NAND2x1p5_ASAP7_75t_L g189 ( .A(n_122), .B(n_110), .Y(n_189) );
INVx2_ASAP7_75t_L g190 ( .A(n_134), .Y(n_190) );
AND2x4_ASAP7_75t_L g191 ( .A(n_123), .B(n_88), .Y(n_191) );
INVxp67_ASAP7_75t_SL g192 ( .A(n_155), .Y(n_192) );
AND2x4_ASAP7_75t_L g193 ( .A(n_123), .B(n_137), .Y(n_193) );
INVx3_ASAP7_75t_L g194 ( .A(n_157), .Y(n_194) );
INVx2_ASAP7_75t_L g195 ( .A(n_132), .Y(n_195) );
NOR2xp33_ASAP7_75t_L g196 ( .A(n_140), .B(n_92), .Y(n_196) );
NOR2xp33_ASAP7_75t_L g197 ( .A(n_141), .B(n_95), .Y(n_197) );
BUFx3_ASAP7_75t_L g198 ( .A(n_150), .Y(n_198) );
AND2x4_ASAP7_75t_L g199 ( .A(n_137), .B(n_106), .Y(n_199) );
NAND2xp5_ASAP7_75t_L g200 ( .A(n_138), .B(n_114), .Y(n_200) );
HB1xp67_ASAP7_75t_L g201 ( .A(n_155), .Y(n_201) );
INVx1_ASAP7_75t_L g202 ( .A(n_134), .Y(n_202) );
BUFx4f_ASAP7_75t_L g203 ( .A(n_138), .Y(n_203) );
INVx2_ASAP7_75t_L g204 ( .A(n_132), .Y(n_204) );
INVx1_ASAP7_75t_L g205 ( .A(n_157), .Y(n_205) );
AND2x4_ASAP7_75t_L g206 ( .A(n_142), .B(n_114), .Y(n_206) );
INVx1_ASAP7_75t_L g207 ( .A(n_157), .Y(n_207) );
HB1xp67_ASAP7_75t_L g208 ( .A(n_148), .Y(n_208) );
NAND2xp5_ASAP7_75t_L g209 ( .A(n_142), .B(n_115), .Y(n_209) );
INVx2_ASAP7_75t_L g210 ( .A(n_127), .Y(n_210) );
NAND2xp5_ASAP7_75t_SL g211 ( .A(n_160), .B(n_116), .Y(n_211) );
INVx4_ASAP7_75t_L g212 ( .A(n_132), .Y(n_212) );
INVx2_ASAP7_75t_L g213 ( .A(n_127), .Y(n_213) );
INVx1_ASAP7_75t_L g214 ( .A(n_150), .Y(n_214) );
INVx1_ASAP7_75t_SL g215 ( .A(n_124), .Y(n_215) );
INVx4_ASAP7_75t_L g216 ( .A(n_132), .Y(n_216) );
NOR3xp33_ASAP7_75t_SL g217 ( .A(n_167), .B(n_144), .C(n_158), .Y(n_217) );
AO22x1_ASAP7_75t_L g218 ( .A1(n_172), .A2(n_117), .B1(n_152), .B2(n_146), .Y(n_218) );
INVx1_ASAP7_75t_SL g219 ( .A(n_163), .Y(n_219) );
INVx1_ASAP7_75t_L g220 ( .A(n_205), .Y(n_220) );
NAND2xp5_ASAP7_75t_L g221 ( .A(n_193), .B(n_143), .Y(n_221) );
INVx2_ASAP7_75t_SL g222 ( .A(n_184), .Y(n_222) );
AND2x4_ASAP7_75t_L g223 ( .A(n_192), .B(n_146), .Y(n_223) );
NOR3xp33_ASAP7_75t_SL g224 ( .A(n_196), .B(n_197), .C(n_178), .Y(n_224) );
NOR2xp33_ASAP7_75t_L g225 ( .A(n_201), .B(n_147), .Y(n_225) );
NAND2xp5_ASAP7_75t_L g226 ( .A(n_193), .B(n_152), .Y(n_226) );
AOI22xp5_ASAP7_75t_L g227 ( .A1(n_179), .A2(n_143), .B1(n_159), .B2(n_135), .Y(n_227) );
BUFx3_ASAP7_75t_L g228 ( .A(n_184), .Y(n_228) );
BUFx2_ASAP7_75t_L g229 ( .A(n_163), .Y(n_229) );
INVx2_ASAP7_75t_L g230 ( .A(n_194), .Y(n_230) );
AND2x4_ASAP7_75t_L g231 ( .A(n_172), .B(n_145), .Y(n_231) );
INVx1_ASAP7_75t_L g232 ( .A(n_205), .Y(n_232) );
INVxp67_ASAP7_75t_SL g233 ( .A(n_165), .Y(n_233) );
BUFx12f_ASAP7_75t_SL g234 ( .A(n_199), .Y(n_234) );
NOR2xp33_ASAP7_75t_R g235 ( .A(n_168), .B(n_154), .Y(n_235) );
NAND2xp5_ASAP7_75t_L g236 ( .A(n_193), .B(n_115), .Y(n_236) );
INVx2_ASAP7_75t_L g237 ( .A(n_194), .Y(n_237) );
AND2x2_ASAP7_75t_L g238 ( .A(n_193), .B(n_5), .Y(n_238) );
INVx1_ASAP7_75t_L g239 ( .A(n_207), .Y(n_239) );
BUFx2_ASAP7_75t_L g240 ( .A(n_184), .Y(n_240) );
INVx1_ASAP7_75t_SL g241 ( .A(n_215), .Y(n_241) );
AND2x4_ASAP7_75t_L g242 ( .A(n_176), .B(n_5), .Y(n_242) );
INVx2_ASAP7_75t_L g243 ( .A(n_194), .Y(n_243) );
NAND2xp5_ASAP7_75t_L g244 ( .A(n_203), .B(n_100), .Y(n_244) );
INVx3_ASAP7_75t_L g245 ( .A(n_184), .Y(n_245) );
OAI22xp5_ASAP7_75t_SL g246 ( .A1(n_208), .A2(n_133), .B1(n_129), .B2(n_128), .Y(n_246) );
NAND2xp5_ASAP7_75t_L g247 ( .A(n_203), .B(n_129), .Y(n_247) );
BUFx3_ASAP7_75t_L g248 ( .A(n_184), .Y(n_248) );
NAND2xp5_ASAP7_75t_L g249 ( .A(n_203), .B(n_129), .Y(n_249) );
NAND2xp5_ASAP7_75t_L g250 ( .A(n_199), .B(n_128), .Y(n_250) );
AND2x4_ASAP7_75t_L g251 ( .A(n_211), .B(n_6), .Y(n_251) );
O2A1O1Ixp33_ASAP7_75t_L g252 ( .A1(n_173), .A2(n_127), .B(n_128), .C(n_119), .Y(n_252) );
NOR3xp33_ASAP7_75t_SL g253 ( .A(n_170), .B(n_6), .C(n_7), .Y(n_253) );
INVx1_ASAP7_75t_L g254 ( .A(n_207), .Y(n_254) );
NOR2xp33_ASAP7_75t_R g255 ( .A(n_168), .B(n_36), .Y(n_255) );
INVx2_ASAP7_75t_L g256 ( .A(n_194), .Y(n_256) );
NOR2xp33_ASAP7_75t_L g257 ( .A(n_173), .B(n_37), .Y(n_257) );
NAND2xp5_ASAP7_75t_L g258 ( .A(n_199), .B(n_132), .Y(n_258) );
INVx3_ASAP7_75t_L g259 ( .A(n_198), .Y(n_259) );
INVx3_ASAP7_75t_L g260 ( .A(n_198), .Y(n_260) );
NAND2xp5_ASAP7_75t_L g261 ( .A(n_199), .B(n_8), .Y(n_261) );
OR2x2_ASAP7_75t_L g262 ( .A(n_171), .B(n_9), .Y(n_262) );
AND2x2_ASAP7_75t_L g263 ( .A(n_179), .B(n_10), .Y(n_263) );
NAND2xp5_ASAP7_75t_L g264 ( .A(n_206), .B(n_12), .Y(n_264) );
NAND2xp5_ASAP7_75t_SL g265 ( .A(n_164), .B(n_38), .Y(n_265) );
AND2x4_ASAP7_75t_L g266 ( .A(n_206), .B(n_12), .Y(n_266) );
BUFx6f_ASAP7_75t_L g267 ( .A(n_164), .Y(n_267) );
INVx3_ASAP7_75t_L g268 ( .A(n_198), .Y(n_268) );
INVx5_ASAP7_75t_L g269 ( .A(n_212), .Y(n_269) );
BUFx3_ASAP7_75t_L g270 ( .A(n_165), .Y(n_270) );
INVx1_ASAP7_75t_L g271 ( .A(n_189), .Y(n_271) );
NAND2xp33_ASAP7_75t_SL g272 ( .A(n_181), .B(n_13), .Y(n_272) );
INVx1_ASAP7_75t_L g273 ( .A(n_189), .Y(n_273) );
INVx1_ASAP7_75t_L g274 ( .A(n_189), .Y(n_274) );
INVx4_ASAP7_75t_L g275 ( .A(n_164), .Y(n_275) );
BUFx2_ASAP7_75t_L g276 ( .A(n_234), .Y(n_276) );
INVx1_ASAP7_75t_L g277 ( .A(n_220), .Y(n_277) );
O2A1O1Ixp33_ASAP7_75t_SL g278 ( .A1(n_265), .A2(n_200), .B(n_209), .C(n_214), .Y(n_278) );
O2A1O1Ixp5_ASAP7_75t_L g279 ( .A1(n_218), .A2(n_187), .B(n_206), .C(n_191), .Y(n_279) );
INVx1_ASAP7_75t_SL g280 ( .A(n_219), .Y(n_280) );
BUFx3_ASAP7_75t_L g281 ( .A(n_228), .Y(n_281) );
AOI21xp5_ASAP7_75t_SL g282 ( .A1(n_266), .A2(n_165), .B(n_166), .Y(n_282) );
CKINVDCx20_ASAP7_75t_R g283 ( .A(n_235), .Y(n_283) );
BUFx2_ASAP7_75t_L g284 ( .A(n_234), .Y(n_284) );
INVx2_ASAP7_75t_L g285 ( .A(n_220), .Y(n_285) );
AND2x4_ASAP7_75t_L g286 ( .A(n_270), .B(n_206), .Y(n_286) );
OR2x2_ASAP7_75t_L g287 ( .A(n_229), .B(n_166), .Y(n_287) );
AOI21xp5_ASAP7_75t_L g288 ( .A1(n_221), .A2(n_187), .B(n_166), .Y(n_288) );
INVx1_ASAP7_75t_L g289 ( .A(n_232), .Y(n_289) );
O2A1O1Ixp33_ASAP7_75t_L g290 ( .A1(n_226), .A2(n_236), .B(n_264), .C(n_261), .Y(n_290) );
A2O1A1Ixp33_ASAP7_75t_SL g291 ( .A1(n_257), .A2(n_214), .B(n_177), .C(n_188), .Y(n_291) );
INVx2_ASAP7_75t_L g292 ( .A(n_232), .Y(n_292) );
NAND2xp5_ASAP7_75t_L g293 ( .A(n_223), .B(n_179), .Y(n_293) );
INVx2_ASAP7_75t_L g294 ( .A(n_239), .Y(n_294) );
AO32x2_ASAP7_75t_L g295 ( .A1(n_246), .A2(n_216), .A3(n_212), .B1(n_179), .B2(n_181), .Y(n_295) );
INVx2_ASAP7_75t_L g296 ( .A(n_239), .Y(n_296) );
AO21x2_ASAP7_75t_L g297 ( .A1(n_227), .A2(n_252), .B(n_263), .Y(n_297) );
HB1xp67_ASAP7_75t_L g298 ( .A(n_241), .Y(n_298) );
NAND2xp5_ASAP7_75t_SL g299 ( .A(n_228), .B(n_168), .Y(n_299) );
INVx1_ASAP7_75t_SL g300 ( .A(n_229), .Y(n_300) );
OAI22xp33_ASAP7_75t_L g301 ( .A1(n_227), .A2(n_187), .B1(n_191), .B2(n_168), .Y(n_301) );
A2O1A1Ixp33_ASAP7_75t_L g302 ( .A1(n_254), .A2(n_191), .B(n_202), .C(n_182), .Y(n_302) );
BUFx4f_ASAP7_75t_SL g303 ( .A(n_251), .Y(n_303) );
AOI21xp5_ASAP7_75t_L g304 ( .A1(n_244), .A2(n_202), .B(n_180), .Y(n_304) );
O2A1O1Ixp33_ASAP7_75t_SL g305 ( .A1(n_258), .A2(n_180), .B(n_182), .C(n_177), .Y(n_305) );
INVx1_ASAP7_75t_L g306 ( .A(n_254), .Y(n_306) );
AND2x4_ASAP7_75t_L g307 ( .A(n_270), .B(n_191), .Y(n_307) );
OAI22xp5_ASAP7_75t_L g308 ( .A1(n_233), .A2(n_169), .B1(n_190), .B2(n_188), .Y(n_308) );
INVx1_ASAP7_75t_L g309 ( .A(n_271), .Y(n_309) );
AND2x4_ASAP7_75t_L g310 ( .A(n_270), .B(n_14), .Y(n_310) );
INVx2_ASAP7_75t_L g311 ( .A(n_230), .Y(n_311) );
BUFx2_ASAP7_75t_L g312 ( .A(n_240), .Y(n_312) );
INVx1_ASAP7_75t_L g313 ( .A(n_271), .Y(n_313) );
INVx3_ASAP7_75t_L g314 ( .A(n_228), .Y(n_314) );
AOI22xp5_ASAP7_75t_L g315 ( .A1(n_266), .A2(n_169), .B1(n_212), .B2(n_216), .Y(n_315) );
BUFx2_ASAP7_75t_L g316 ( .A(n_240), .Y(n_316) );
AND2x4_ASAP7_75t_L g317 ( .A(n_248), .B(n_14), .Y(n_317) );
AOI21xp33_ASAP7_75t_L g318 ( .A1(n_222), .A2(n_216), .B(n_212), .Y(n_318) );
INVx1_ASAP7_75t_SL g319 ( .A(n_266), .Y(n_319) );
NOR2xp33_ASAP7_75t_L g320 ( .A(n_231), .B(n_16), .Y(n_320) );
INVx1_ASAP7_75t_L g321 ( .A(n_273), .Y(n_321) );
OAI22xp5_ASAP7_75t_L g322 ( .A1(n_282), .A2(n_266), .B1(n_274), .B2(n_273), .Y(n_322) );
OAI21x1_ASAP7_75t_L g323 ( .A1(n_290), .A2(n_263), .B(n_238), .Y(n_323) );
AOI22xp33_ASAP7_75t_L g324 ( .A1(n_303), .A2(n_242), .B1(n_251), .B2(n_238), .Y(n_324) );
HB1xp67_ASAP7_75t_L g325 ( .A(n_312), .Y(n_325) );
INVx2_ASAP7_75t_L g326 ( .A(n_285), .Y(n_326) );
OAI222xp33_ASAP7_75t_L g327 ( .A1(n_301), .A2(n_242), .B1(n_262), .B2(n_251), .C1(n_274), .C2(n_231), .Y(n_327) );
AOI21xp5_ASAP7_75t_L g328 ( .A1(n_282), .A2(n_250), .B(n_249), .Y(n_328) );
AOI22xp33_ASAP7_75t_L g329 ( .A1(n_320), .A2(n_242), .B1(n_251), .B2(n_223), .Y(n_329) );
INVx2_ASAP7_75t_L g330 ( .A(n_285), .Y(n_330) );
INVx2_ASAP7_75t_L g331 ( .A(n_292), .Y(n_331) );
INVx4_ASAP7_75t_L g332 ( .A(n_310), .Y(n_332) );
AND2x2_ASAP7_75t_L g333 ( .A(n_292), .B(n_223), .Y(n_333) );
AND2x2_ASAP7_75t_L g334 ( .A(n_294), .B(n_223), .Y(n_334) );
OAI221xp5_ASAP7_75t_L g335 ( .A1(n_293), .A2(n_217), .B1(n_224), .B2(n_246), .C(n_262), .Y(n_335) );
INVx1_ASAP7_75t_L g336 ( .A(n_294), .Y(n_336) );
AOI22xp33_ASAP7_75t_SL g337 ( .A1(n_310), .A2(n_242), .B1(n_231), .B2(n_225), .Y(n_337) );
AND2x2_ASAP7_75t_L g338 ( .A(n_296), .B(n_248), .Y(n_338) );
CKINVDCx5p33_ASAP7_75t_R g339 ( .A(n_283), .Y(n_339) );
NOR2xp33_ASAP7_75t_L g340 ( .A(n_287), .B(n_231), .Y(n_340) );
OR2x2_ASAP7_75t_L g341 ( .A(n_300), .B(n_218), .Y(n_341) );
AOI21xp33_ASAP7_75t_L g342 ( .A1(n_297), .A2(n_247), .B(n_267), .Y(n_342) );
AOI22xp33_ASAP7_75t_L g343 ( .A1(n_317), .A2(n_310), .B1(n_296), .B2(n_289), .Y(n_343) );
INVx1_ASAP7_75t_L g344 ( .A(n_277), .Y(n_344) );
OAI21x1_ASAP7_75t_L g345 ( .A1(n_288), .A2(n_190), .B(n_260), .Y(n_345) );
INVx2_ASAP7_75t_L g346 ( .A(n_277), .Y(n_346) );
INVx3_ASAP7_75t_L g347 ( .A(n_286), .Y(n_347) );
AND2x2_ASAP7_75t_L g348 ( .A(n_289), .B(n_248), .Y(n_348) );
OAI22xp5_ASAP7_75t_L g349 ( .A1(n_319), .A2(n_275), .B1(n_222), .B2(n_259), .Y(n_349) );
AND2x4_ASAP7_75t_L g350 ( .A(n_309), .B(n_275), .Y(n_350) );
NAND2x1_ASAP7_75t_L g351 ( .A(n_306), .B(n_310), .Y(n_351) );
OAI22xp33_ASAP7_75t_L g352 ( .A1(n_332), .A2(n_280), .B1(n_298), .B2(n_287), .Y(n_352) );
INVx5_ASAP7_75t_SL g353 ( .A(n_350), .Y(n_353) );
AOI22xp33_ASAP7_75t_L g354 ( .A1(n_337), .A2(n_317), .B1(n_272), .B2(n_308), .Y(n_354) );
INVx1_ASAP7_75t_L g355 ( .A(n_336), .Y(n_355) );
OAI22xp33_ASAP7_75t_L g356 ( .A1(n_332), .A2(n_312), .B1(n_316), .B2(n_315), .Y(n_356) );
AOI221xp5_ASAP7_75t_L g357 ( .A1(n_335), .A2(n_284), .B1(n_276), .B2(n_307), .C(n_279), .Y(n_357) );
AOI22xp33_ASAP7_75t_L g358 ( .A1(n_337), .A2(n_317), .B1(n_307), .B2(n_316), .Y(n_358) );
AOI221xp5_ASAP7_75t_L g359 ( .A1(n_335), .A2(n_284), .B1(n_276), .B2(n_307), .C(n_306), .Y(n_359) );
NAND2xp5_ASAP7_75t_L g360 ( .A(n_340), .B(n_307), .Y(n_360) );
AO21x2_ASAP7_75t_L g361 ( .A1(n_342), .A2(n_291), .B(n_297), .Y(n_361) );
OAI31xp33_ASAP7_75t_L g362 ( .A1(n_327), .A2(n_317), .A3(n_321), .B(n_313), .Y(n_362) );
NAND2xp5_ASAP7_75t_L g363 ( .A(n_340), .B(n_309), .Y(n_363) );
OAI21xp5_ASAP7_75t_SL g364 ( .A1(n_343), .A2(n_286), .B(n_313), .Y(n_364) );
INVx3_ASAP7_75t_L g365 ( .A(n_332), .Y(n_365) );
AND2x2_ASAP7_75t_L g366 ( .A(n_333), .B(n_321), .Y(n_366) );
OR2x2_ASAP7_75t_L g367 ( .A(n_343), .B(n_297), .Y(n_367) );
INVx1_ASAP7_75t_L g368 ( .A(n_336), .Y(n_368) );
AOI22xp33_ASAP7_75t_L g369 ( .A1(n_324), .A2(n_286), .B1(n_275), .B2(n_281), .Y(n_369) );
OAI22xp33_ASAP7_75t_L g370 ( .A1(n_332), .A2(n_286), .B1(n_275), .B2(n_281), .Y(n_370) );
OAI21xp33_ASAP7_75t_L g371 ( .A1(n_329), .A2(n_253), .B(n_302), .Y(n_371) );
OAI22xp5_ASAP7_75t_L g372 ( .A1(n_324), .A2(n_314), .B1(n_311), .B2(n_260), .Y(n_372) );
AND2x4_ASAP7_75t_L g373 ( .A(n_332), .B(n_314), .Y(n_373) );
INVx2_ASAP7_75t_L g374 ( .A(n_326), .Y(n_374) );
AOI222xp33_ASAP7_75t_L g375 ( .A1(n_327), .A2(n_299), .B1(n_314), .B2(n_267), .C1(n_311), .C2(n_230), .Y(n_375) );
NOR2x1_ASAP7_75t_SL g376 ( .A(n_332), .B(n_267), .Y(n_376) );
AND2x2_ASAP7_75t_L g377 ( .A(n_333), .B(n_295), .Y(n_377) );
OR2x2_ASAP7_75t_L g378 ( .A(n_355), .B(n_351), .Y(n_378) );
NOR2x2_ASAP7_75t_L g379 ( .A(n_374), .B(n_339), .Y(n_379) );
OR2x6_ASAP7_75t_L g380 ( .A(n_364), .B(n_351), .Y(n_380) );
OAI33xp33_ASAP7_75t_L g381 ( .A1(n_352), .A2(n_341), .A3(n_322), .B1(n_344), .B2(n_336), .B3(n_349), .Y(n_381) );
NAND2xp5_ASAP7_75t_L g382 ( .A(n_366), .B(n_329), .Y(n_382) );
INVx2_ASAP7_75t_L g383 ( .A(n_374), .Y(n_383) );
OAI221xp5_ASAP7_75t_L g384 ( .A1(n_359), .A2(n_322), .B1(n_351), .B2(n_341), .C(n_325), .Y(n_384) );
AND2x2_ASAP7_75t_L g385 ( .A(n_366), .B(n_346), .Y(n_385) );
INVx1_ASAP7_75t_L g386 ( .A(n_355), .Y(n_386) );
CKINVDCx5p33_ASAP7_75t_R g387 ( .A(n_358), .Y(n_387) );
AND2x2_ASAP7_75t_L g388 ( .A(n_368), .B(n_346), .Y(n_388) );
AND2x4_ASAP7_75t_SL g389 ( .A(n_365), .B(n_350), .Y(n_389) );
OAI332xp33_ASAP7_75t_L g390 ( .A1(n_363), .A2(n_341), .A3(n_344), .B1(n_346), .B2(n_326), .B3(n_330), .C1(n_331), .C2(n_24), .Y(n_390) );
AOI21xp5_ASAP7_75t_L g391 ( .A1(n_374), .A2(n_330), .B(n_331), .Y(n_391) );
INVx2_ASAP7_75t_SL g392 ( .A(n_365), .Y(n_392) );
INVx1_ASAP7_75t_L g393 ( .A(n_368), .Y(n_393) );
BUFx2_ASAP7_75t_L g394 ( .A(n_365), .Y(n_394) );
AND2x2_ASAP7_75t_L g395 ( .A(n_377), .B(n_346), .Y(n_395) );
OAI22xp5_ASAP7_75t_SL g396 ( .A1(n_354), .A2(n_339), .B1(n_325), .B2(n_344), .Y(n_396) );
OAI221xp5_ASAP7_75t_L g397 ( .A1(n_357), .A2(n_342), .B1(n_347), .B2(n_328), .C(n_333), .Y(n_397) );
AO21x2_ASAP7_75t_L g398 ( .A1(n_361), .A2(n_345), .B(n_323), .Y(n_398) );
OAI21xp5_ASAP7_75t_SL g399 ( .A1(n_362), .A2(n_350), .B(n_334), .Y(n_399) );
OR2x2_ASAP7_75t_L g400 ( .A(n_367), .B(n_326), .Y(n_400) );
AOI21xp5_ASAP7_75t_L g401 ( .A1(n_362), .A2(n_326), .B(n_330), .Y(n_401) );
AND2x4_ASAP7_75t_SL g402 ( .A(n_365), .B(n_350), .Y(n_402) );
NOR2xp33_ASAP7_75t_L g403 ( .A(n_360), .B(n_347), .Y(n_403) );
AOI22xp33_ASAP7_75t_L g404 ( .A1(n_371), .A2(n_347), .B1(n_350), .B2(n_334), .Y(n_404) );
INVx2_ASAP7_75t_L g405 ( .A(n_377), .Y(n_405) );
AOI221xp5_ASAP7_75t_L g406 ( .A1(n_364), .A2(n_347), .B1(n_348), .B2(n_328), .C(n_330), .Y(n_406) );
INVx2_ASAP7_75t_L g407 ( .A(n_361), .Y(n_407) );
NOR4xp25_ASAP7_75t_SL g408 ( .A(n_375), .B(n_295), .C(n_278), .D(n_255), .Y(n_408) );
OAI211xp5_ASAP7_75t_L g409 ( .A1(n_375), .A2(n_323), .B(n_331), .C(n_348), .Y(n_409) );
AND2x2_ASAP7_75t_L g410 ( .A(n_405), .B(n_367), .Y(n_410) );
AOI22xp33_ASAP7_75t_L g411 ( .A1(n_396), .A2(n_356), .B1(n_369), .B2(n_353), .Y(n_411) );
INVx2_ASAP7_75t_L g412 ( .A(n_383), .Y(n_412) );
OR2x2_ASAP7_75t_L g413 ( .A(n_405), .B(n_361), .Y(n_413) );
AO31x2_ASAP7_75t_L g414 ( .A1(n_401), .A2(n_372), .A3(n_331), .B(n_376), .Y(n_414) );
NOR2x1_ASAP7_75t_L g415 ( .A(n_378), .B(n_370), .Y(n_415) );
AND2x2_ASAP7_75t_L g416 ( .A(n_395), .B(n_353), .Y(n_416) );
AND2x2_ASAP7_75t_L g417 ( .A(n_395), .B(n_353), .Y(n_417) );
NAND2xp5_ASAP7_75t_L g418 ( .A(n_386), .B(n_323), .Y(n_418) );
NAND2xp5_ASAP7_75t_L g419 ( .A(n_393), .B(n_323), .Y(n_419) );
OAI31xp33_ASAP7_75t_L g420 ( .A1(n_384), .A2(n_338), .A3(n_349), .B(n_373), .Y(n_420) );
OAI22xp5_ASAP7_75t_L g421 ( .A1(n_399), .A2(n_353), .B1(n_373), .B2(n_338), .Y(n_421) );
AOI21xp5_ASAP7_75t_L g422 ( .A1(n_391), .A2(n_345), .B(n_376), .Y(n_422) );
INVx2_ASAP7_75t_SL g423 ( .A(n_389), .Y(n_423) );
INVx1_ASAP7_75t_SL g424 ( .A(n_379), .Y(n_424) );
OAI211xp5_ASAP7_75t_L g425 ( .A1(n_399), .A2(n_338), .B(n_295), .C(n_353), .Y(n_425) );
INVx2_ASAP7_75t_L g426 ( .A(n_383), .Y(n_426) );
OAI22xp5_ASAP7_75t_L g427 ( .A1(n_380), .A2(n_373), .B1(n_295), .B2(n_245), .Y(n_427) );
AND2x2_ASAP7_75t_L g428 ( .A(n_385), .B(n_373), .Y(n_428) );
OR2x2_ASAP7_75t_SL g429 ( .A(n_378), .B(n_295), .Y(n_429) );
OAI33xp33_ASAP7_75t_L g430 ( .A1(n_396), .A2(n_16), .A3(n_17), .B1(n_19), .B2(n_20), .B3(n_21), .Y(n_430) );
INVx2_ASAP7_75t_SL g431 ( .A(n_389), .Y(n_431) );
INVx2_ASAP7_75t_L g432 ( .A(n_407), .Y(n_432) );
OAI21xp5_ASAP7_75t_SL g433 ( .A1(n_409), .A2(n_267), .B(n_245), .Y(n_433) );
INVx1_ASAP7_75t_L g434 ( .A(n_393), .Y(n_434) );
NOR2xp33_ASAP7_75t_SL g435 ( .A(n_380), .B(n_267), .Y(n_435) );
NAND2xp5_ASAP7_75t_L g436 ( .A(n_388), .B(n_345), .Y(n_436) );
INVx2_ASAP7_75t_L g437 ( .A(n_407), .Y(n_437) );
AND2x4_ASAP7_75t_L g438 ( .A(n_380), .B(n_345), .Y(n_438) );
OAI221xp5_ASAP7_75t_L g439 ( .A1(n_404), .A2(n_260), .B1(n_268), .B2(n_259), .C(n_304), .Y(n_439) );
AND2x2_ASAP7_75t_L g440 ( .A(n_385), .B(n_21), .Y(n_440) );
NOR2x1_ASAP7_75t_L g441 ( .A(n_394), .B(n_268), .Y(n_441) );
HB1xp67_ASAP7_75t_L g442 ( .A(n_388), .Y(n_442) );
INVx3_ASAP7_75t_L g443 ( .A(n_380), .Y(n_443) );
AND2x4_ASAP7_75t_L g444 ( .A(n_380), .B(n_68), .Y(n_444) );
NAND2xp5_ASAP7_75t_L g445 ( .A(n_400), .B(n_237), .Y(n_445) );
AOI31xp33_ASAP7_75t_L g446 ( .A1(n_381), .A2(n_305), .A3(n_318), .B(n_23), .Y(n_446) );
AND2x2_ASAP7_75t_L g447 ( .A(n_400), .B(n_23), .Y(n_447) );
NAND2xp5_ASAP7_75t_L g448 ( .A(n_382), .B(n_237), .Y(n_448) );
AND2x2_ASAP7_75t_L g449 ( .A(n_394), .B(n_24), .Y(n_449) );
INVx2_ASAP7_75t_L g450 ( .A(n_398), .Y(n_450) );
AND2x4_ASAP7_75t_L g451 ( .A(n_398), .B(n_28), .Y(n_451) );
INVx1_ASAP7_75t_L g452 ( .A(n_398), .Y(n_452) );
AND2x2_ASAP7_75t_L g453 ( .A(n_392), .B(n_243), .Y(n_453) );
OAI33xp33_ASAP7_75t_L g454 ( .A1(n_387), .A2(n_162), .A3(n_161), .B1(n_183), .B2(n_186), .B3(n_195), .Y(n_454) );
AND2x2_ASAP7_75t_L g455 ( .A(n_392), .B(n_243), .Y(n_455) );
INVx2_ASAP7_75t_L g456 ( .A(n_397), .Y(n_456) );
NAND2xp5_ASAP7_75t_L g457 ( .A(n_442), .B(n_390), .Y(n_457) );
AND2x2_ASAP7_75t_L g458 ( .A(n_410), .B(n_406), .Y(n_458) );
AND2x2_ASAP7_75t_L g459 ( .A(n_410), .B(n_402), .Y(n_459) );
NOR2xp33_ASAP7_75t_L g460 ( .A(n_424), .B(n_387), .Y(n_460) );
OR2x2_ASAP7_75t_L g461 ( .A(n_418), .B(n_402), .Y(n_461) );
AND2x4_ASAP7_75t_L g462 ( .A(n_443), .B(n_403), .Y(n_462) );
AND2x2_ASAP7_75t_L g463 ( .A(n_434), .B(n_408), .Y(n_463) );
OR2x2_ASAP7_75t_L g464 ( .A(n_418), .B(n_210), .Y(n_464) );
AND2x2_ASAP7_75t_L g465 ( .A(n_434), .B(n_31), .Y(n_465) );
INVx2_ASAP7_75t_L g466 ( .A(n_432), .Y(n_466) );
AND2x2_ASAP7_75t_L g467 ( .A(n_443), .B(n_32), .Y(n_467) );
NAND2xp5_ASAP7_75t_L g468 ( .A(n_440), .B(n_256), .Y(n_468) );
NAND3xp33_ASAP7_75t_L g469 ( .A(n_452), .B(n_174), .C(n_175), .Y(n_469) );
AND2x4_ASAP7_75t_L g470 ( .A(n_443), .B(n_35), .Y(n_470) );
INVx1_ASAP7_75t_L g471 ( .A(n_432), .Y(n_471) );
OR2x2_ASAP7_75t_L g472 ( .A(n_419), .B(n_213), .Y(n_472) );
INVx1_ASAP7_75t_L g473 ( .A(n_432), .Y(n_473) );
AND2x2_ASAP7_75t_L g474 ( .A(n_443), .B(n_42), .Y(n_474) );
NAND2xp5_ASAP7_75t_L g475 ( .A(n_440), .B(n_256), .Y(n_475) );
INVx2_ASAP7_75t_L g476 ( .A(n_437), .Y(n_476) );
AND2x2_ASAP7_75t_L g477 ( .A(n_428), .B(n_44), .Y(n_477) );
NAND2xp5_ASAP7_75t_SL g478 ( .A(n_424), .B(n_268), .Y(n_478) );
NAND2xp5_ASAP7_75t_L g479 ( .A(n_447), .B(n_259), .Y(n_479) );
INVx1_ASAP7_75t_SL g480 ( .A(n_449), .Y(n_480) );
INVx1_ASAP7_75t_L g481 ( .A(n_437), .Y(n_481) );
INVxp67_ASAP7_75t_SL g482 ( .A(n_412), .Y(n_482) );
NOR2x1_ASAP7_75t_L g483 ( .A(n_444), .B(n_216), .Y(n_483) );
INVx1_ASAP7_75t_L g484 ( .A(n_437), .Y(n_484) );
AND2x4_ASAP7_75t_L g485 ( .A(n_438), .B(n_46), .Y(n_485) );
NAND2xp5_ASAP7_75t_L g486 ( .A(n_447), .B(n_210), .Y(n_486) );
INVx3_ASAP7_75t_L g487 ( .A(n_451), .Y(n_487) );
BUFx2_ASAP7_75t_L g488 ( .A(n_412), .Y(n_488) );
OR2x2_ASAP7_75t_L g489 ( .A(n_419), .B(n_429), .Y(n_489) );
CKINVDCx16_ASAP7_75t_R g490 ( .A(n_423), .Y(n_490) );
INVx1_ASAP7_75t_L g491 ( .A(n_412), .Y(n_491) );
BUFx2_ASAP7_75t_L g492 ( .A(n_426), .Y(n_492) );
OR2x2_ASAP7_75t_L g493 ( .A(n_429), .B(n_213), .Y(n_493) );
NAND2xp5_ASAP7_75t_L g494 ( .A(n_449), .B(n_47), .Y(n_494) );
INVx2_ASAP7_75t_L g495 ( .A(n_426), .Y(n_495) );
INVx2_ASAP7_75t_L g496 ( .A(n_426), .Y(n_496) );
AND2x2_ASAP7_75t_L g497 ( .A(n_452), .B(n_48), .Y(n_497) );
NAND2xp5_ASAP7_75t_L g498 ( .A(n_416), .B(n_49), .Y(n_498) );
INVx1_ASAP7_75t_L g499 ( .A(n_445), .Y(n_499) );
NOR3xp33_ASAP7_75t_SL g500 ( .A(n_430), .B(n_51), .C(n_57), .Y(n_500) );
NOR2xp33_ASAP7_75t_L g501 ( .A(n_423), .B(n_61), .Y(n_501) );
NAND4xp25_ASAP7_75t_SL g502 ( .A(n_425), .B(n_66), .C(n_69), .D(n_72), .Y(n_502) );
INVx1_ASAP7_75t_L g503 ( .A(n_413), .Y(n_503) );
HB1xp67_ASAP7_75t_L g504 ( .A(n_431), .Y(n_504) );
INVxp67_ASAP7_75t_L g505 ( .A(n_416), .Y(n_505) );
NAND2xp5_ASAP7_75t_SL g506 ( .A(n_444), .B(n_269), .Y(n_506) );
NAND2xp5_ASAP7_75t_SL g507 ( .A(n_490), .B(n_444), .Y(n_507) );
NOR2xp67_ASAP7_75t_L g508 ( .A(n_502), .B(n_433), .Y(n_508) );
OAI22xp5_ASAP7_75t_L g509 ( .A1(n_457), .A2(n_411), .B1(n_421), .B2(n_425), .Y(n_509) );
OAI22xp5_ASAP7_75t_L g510 ( .A1(n_500), .A2(n_421), .B1(n_444), .B2(n_427), .Y(n_510) );
NOR3xp33_ASAP7_75t_L g511 ( .A(n_478), .B(n_430), .C(n_446), .Y(n_511) );
AOI22xp33_ASAP7_75t_L g512 ( .A1(n_462), .A2(n_427), .B1(n_438), .B2(n_456), .Y(n_512) );
AOI21xp33_ASAP7_75t_L g513 ( .A1(n_493), .A2(n_446), .B(n_450), .Y(n_513) );
NOR2x1_ASAP7_75t_L g514 ( .A(n_483), .B(n_441), .Y(n_514) );
OAI21xp5_ASAP7_75t_L g515 ( .A1(n_506), .A2(n_441), .B(n_422), .Y(n_515) );
AOI22xp5_ASAP7_75t_L g516 ( .A1(n_460), .A2(n_435), .B1(n_415), .B2(n_417), .Y(n_516) );
O2A1O1Ixp33_ASAP7_75t_L g517 ( .A1(n_493), .A2(n_420), .B(n_448), .C(n_451), .Y(n_517) );
NAND4xp75_ASAP7_75t_L g518 ( .A(n_463), .B(n_417), .C(n_422), .D(n_450), .Y(n_518) );
AOI22xp5_ASAP7_75t_L g519 ( .A1(n_462), .A2(n_438), .B1(n_451), .B2(n_454), .Y(n_519) );
AND2x2_ASAP7_75t_L g520 ( .A(n_505), .B(n_436), .Y(n_520) );
NAND2x1p5_ASAP7_75t_L g521 ( .A(n_485), .B(n_455), .Y(n_521) );
OAI321xp33_ASAP7_75t_L g522 ( .A1(n_463), .A2(n_439), .A3(n_448), .B1(n_445), .B2(n_455), .C(n_453), .Y(n_522) );
NAND2xp5_ASAP7_75t_L g523 ( .A(n_503), .B(n_414), .Y(n_523) );
AOI22xp5_ASAP7_75t_L g524 ( .A1(n_462), .A2(n_453), .B1(n_439), .B2(n_245), .Y(n_524) );
NAND2xp5_ASAP7_75t_L g525 ( .A(n_489), .B(n_414), .Y(n_525) );
AOI21xp33_ASAP7_75t_SL g526 ( .A1(n_504), .A2(n_74), .B(n_414), .Y(n_526) );
NAND2xp5_ASAP7_75t_L g527 ( .A(n_499), .B(n_414), .Y(n_527) );
AOI22xp5_ASAP7_75t_L g528 ( .A1(n_458), .A2(n_414), .B1(n_162), .B2(n_186), .Y(n_528) );
OAI22xp5_ASAP7_75t_L g529 ( .A1(n_480), .A2(n_414), .B1(n_269), .B2(n_161), .Y(n_529) );
INVx1_ASAP7_75t_L g530 ( .A(n_489), .Y(n_530) );
A2O1A1Ixp33_ASAP7_75t_L g531 ( .A1(n_501), .A2(n_161), .B(n_162), .C(n_204), .Y(n_531) );
AND2x2_ASAP7_75t_L g532 ( .A(n_459), .B(n_186), .Y(n_532) );
AOI322xp5_ASAP7_75t_L g533 ( .A1(n_458), .A2(n_183), .A3(n_195), .B1(n_204), .B2(n_185), .C1(n_175), .C2(n_174), .Y(n_533) );
INVx1_ASAP7_75t_L g534 ( .A(n_488), .Y(n_534) );
OAI221xp5_ASAP7_75t_SL g535 ( .A1(n_461), .A2(n_183), .B1(n_195), .B2(n_204), .C(n_185), .Y(n_535) );
AOI221xp5_ASAP7_75t_L g536 ( .A1(n_486), .A2(n_475), .B1(n_468), .B2(n_479), .C(n_481), .Y(n_536) );
AOI222xp33_ASAP7_75t_L g537 ( .A1(n_477), .A2(n_174), .B1(n_175), .B2(n_185), .C1(n_269), .C2(n_459), .Y(n_537) );
NAND3xp33_ASAP7_75t_L g538 ( .A(n_467), .B(n_174), .C(n_175), .Y(n_538) );
INVxp67_ASAP7_75t_L g539 ( .A(n_477), .Y(n_539) );
OR2x2_ASAP7_75t_L g540 ( .A(n_461), .B(n_174), .Y(n_540) );
AOI22xp5_ASAP7_75t_L g541 ( .A1(n_485), .A2(n_174), .B1(n_175), .B2(n_185), .Y(n_541) );
INVx1_ASAP7_75t_L g542 ( .A(n_488), .Y(n_542) );
INVx2_ASAP7_75t_L g543 ( .A(n_492), .Y(n_543) );
AOI311xp33_ASAP7_75t_L g544 ( .A1(n_471), .A2(n_175), .A3(n_185), .B(n_269), .C(n_484), .Y(n_544) );
AOI321xp33_ASAP7_75t_SL g545 ( .A1(n_487), .A2(n_185), .A3(n_269), .B1(n_485), .B2(n_470), .C(n_494), .Y(n_545) );
INVx1_ASAP7_75t_L g546 ( .A(n_491), .Y(n_546) );
AOI221xp5_ASAP7_75t_L g547 ( .A1(n_471), .A2(n_269), .B1(n_481), .B2(n_484), .C(n_473), .Y(n_547) );
OAI21x1_ASAP7_75t_SL g548 ( .A1(n_510), .A2(n_496), .B(n_495), .Y(n_548) );
NOR3x1_ASAP7_75t_L g549 ( .A(n_509), .B(n_498), .C(n_469), .Y(n_549) );
INVx3_ASAP7_75t_L g550 ( .A(n_521), .Y(n_550) );
NAND3xp33_ASAP7_75t_SL g551 ( .A(n_511), .B(n_474), .C(n_467), .Y(n_551) );
INVx1_ASAP7_75t_L g552 ( .A(n_546), .Y(n_552) );
AOI221xp5_ASAP7_75t_L g553 ( .A1(n_530), .A2(n_465), .B1(n_473), .B2(n_487), .C(n_491), .Y(n_553) );
HB1xp67_ASAP7_75t_L g554 ( .A(n_534), .Y(n_554) );
INVx2_ASAP7_75t_L g555 ( .A(n_542), .Y(n_555) );
AND2x2_ASAP7_75t_L g556 ( .A(n_520), .B(n_487), .Y(n_556) );
OR2x2_ASAP7_75t_L g557 ( .A(n_525), .B(n_482), .Y(n_557) );
NAND2xp5_ASAP7_75t_SL g558 ( .A(n_508), .B(n_470), .Y(n_558) );
NOR3xp33_ASAP7_75t_SL g559 ( .A(n_522), .B(n_497), .C(n_472), .Y(n_559) );
AND2x2_ASAP7_75t_L g560 ( .A(n_525), .B(n_466), .Y(n_560) );
INVx1_ASAP7_75t_L g561 ( .A(n_543), .Y(n_561) );
NAND2xp33_ASAP7_75t_L g562 ( .A(n_521), .B(n_497), .Y(n_562) );
AND2x2_ASAP7_75t_L g563 ( .A(n_512), .B(n_476), .Y(n_563) );
INVx1_ASAP7_75t_L g564 ( .A(n_527), .Y(n_564) );
INVx1_ASAP7_75t_L g565 ( .A(n_523), .Y(n_565) );
INVx2_ASAP7_75t_L g566 ( .A(n_523), .Y(n_566) );
INVxp67_ASAP7_75t_SL g567 ( .A(n_538), .Y(n_567) );
XOR2x2_ASAP7_75t_L g568 ( .A(n_507), .B(n_464), .Y(n_568) );
NAND2xp5_ASAP7_75t_L g569 ( .A(n_536), .B(n_476), .Y(n_569) );
NOR2xp33_ASAP7_75t_L g570 ( .A(n_539), .B(n_464), .Y(n_570) );
NAND2xp33_ASAP7_75t_SL g571 ( .A(n_545), .B(n_496), .Y(n_571) );
NAND2xp5_ASAP7_75t_L g572 ( .A(n_516), .B(n_517), .Y(n_572) );
NOR2xp33_ASAP7_75t_L g573 ( .A(n_518), .B(n_472), .Y(n_573) );
OAI21xp33_ASAP7_75t_SL g574 ( .A1(n_558), .A2(n_519), .B(n_515), .Y(n_574) );
INVx1_ASAP7_75t_L g575 ( .A(n_554), .Y(n_575) );
AOI22xp5_ASAP7_75t_L g576 ( .A1(n_551), .A2(n_524), .B1(n_532), .B2(n_537), .Y(n_576) );
A2O1A1Ixp33_ASAP7_75t_L g577 ( .A1(n_559), .A2(n_526), .B(n_513), .C(n_514), .Y(n_577) );
NOR2xp33_ASAP7_75t_L g578 ( .A(n_572), .B(n_540), .Y(n_578) );
AOI21xp33_ASAP7_75t_L g579 ( .A1(n_573), .A2(n_529), .B(n_528), .Y(n_579) );
OAI221xp5_ASAP7_75t_L g580 ( .A1(n_571), .A2(n_544), .B1(n_547), .B2(n_541), .C(n_535), .Y(n_580) );
NOR3xp33_ASAP7_75t_L g581 ( .A(n_571), .B(n_531), .C(n_495), .Y(n_581) );
AOI22xp5_ASAP7_75t_L g582 ( .A1(n_568), .A2(n_533), .B1(n_562), .B2(n_563), .Y(n_582) );
AOI21xp5_ASAP7_75t_SL g583 ( .A1(n_567), .A2(n_553), .B(n_562), .Y(n_583) );
OAI21xp5_ASAP7_75t_L g584 ( .A1(n_569), .A2(n_568), .B(n_550), .Y(n_584) );
OAI31xp33_ASAP7_75t_L g585 ( .A1(n_550), .A2(n_563), .A3(n_564), .B(n_570), .Y(n_585) );
NAND2xp5_ASAP7_75t_SL g586 ( .A(n_548), .B(n_550), .Y(n_586) );
INVx2_ASAP7_75t_SL g587 ( .A(n_557), .Y(n_587) );
AND2x2_ASAP7_75t_L g588 ( .A(n_560), .B(n_556), .Y(n_588) );
AOI22xp33_ASAP7_75t_L g589 ( .A1(n_548), .A2(n_564), .B1(n_565), .B2(n_556), .Y(n_589) );
INVx2_ASAP7_75t_L g590 ( .A(n_557), .Y(n_590) );
NAND2xp5_ASAP7_75t_SL g591 ( .A(n_584), .B(n_566), .Y(n_591) );
INVx5_ASAP7_75t_L g592 ( .A(n_587), .Y(n_592) );
AOI22xp33_ASAP7_75t_L g593 ( .A1(n_581), .A2(n_555), .B1(n_552), .B2(n_561), .Y(n_593) );
AOI221xp5_ASAP7_75t_L g594 ( .A1(n_583), .A2(n_585), .B1(n_589), .B2(n_574), .C(n_575), .Y(n_594) );
AOI222xp33_ASAP7_75t_L g595 ( .A1(n_586), .A2(n_549), .B1(n_555), .B2(n_577), .C1(n_590), .C2(n_580), .Y(n_595) );
NAND2xp5_ASAP7_75t_L g596 ( .A(n_590), .B(n_588), .Y(n_596) );
OAI22xp5_ASAP7_75t_SL g597 ( .A1(n_576), .A2(n_583), .B1(n_577), .B2(n_586), .Y(n_597) );
NAND3xp33_ASAP7_75t_SL g598 ( .A(n_579), .B(n_577), .C(n_584), .Y(n_598) );
NAND2xp5_ASAP7_75t_L g599 ( .A(n_578), .B(n_587), .Y(n_599) );
OAI221xp5_ASAP7_75t_SL g600 ( .A1(n_574), .A2(n_585), .B1(n_583), .B2(n_582), .C(n_577), .Y(n_600) );
CKINVDCx5p33_ASAP7_75t_R g601 ( .A(n_598), .Y(n_601) );
XOR2xp5_ASAP7_75t_L g602 ( .A(n_597), .B(n_599), .Y(n_602) );
OAI211xp5_ASAP7_75t_L g603 ( .A1(n_595), .A2(n_600), .B(n_594), .C(n_591), .Y(n_603) );
NAND3x1_ASAP7_75t_L g604 ( .A(n_603), .B(n_596), .C(n_592), .Y(n_604) );
INVx1_ASAP7_75t_L g605 ( .A(n_601), .Y(n_605) );
AND2x4_ASAP7_75t_L g606 ( .A(n_605), .B(n_592), .Y(n_606) );
INVx1_ASAP7_75t_L g607 ( .A(n_604), .Y(n_607) );
AND2x4_ASAP7_75t_L g608 ( .A(n_606), .B(n_592), .Y(n_608) );
AOI22xp5_ASAP7_75t_L g609 ( .A1(n_608), .A2(n_606), .B1(n_602), .B2(n_607), .Y(n_609) );
AOI21xp5_ASAP7_75t_L g610 ( .A1(n_609), .A2(n_608), .B(n_593), .Y(n_610) );
endmodule