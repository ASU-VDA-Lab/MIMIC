module fake_jpeg_10896_n_589 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_589);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_589;

wire n_529;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_547;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_582;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_387;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_539;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_442;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_570;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_419;
wire n_378;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx3_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

INVx3_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

BUFx8_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_16),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

INVxp67_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_5),
.Y(n_26)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_15),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_16),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_8),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_3),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_6),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_8),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_13),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_6),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_2),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_10),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_4),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_14),
.Y(n_42)
);

BUFx5_ASAP7_75t_L g43 ( 
.A(n_1),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_9),
.Y(n_44)
);

BUFx24_ASAP7_75t_L g45 ( 
.A(n_17),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_13),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_17),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_9),
.Y(n_48)
);

BUFx8_ASAP7_75t_L g49 ( 
.A(n_17),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_9),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_5),
.Y(n_51)
);

BUFx8_ASAP7_75t_L g52 ( 
.A(n_0),
.Y(n_52)
);

BUFx2_ASAP7_75t_L g53 ( 
.A(n_14),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_11),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_1),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_11),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_15),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_42),
.B(n_47),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_58),
.B(n_78),
.Y(n_135)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_35),
.Y(n_59)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_59),
.Y(n_137)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_35),
.Y(n_60)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_60),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_29),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_61),
.Y(n_127)
);

OR2x2_ASAP7_75t_L g62 ( 
.A(n_47),
.B(n_16),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_62),
.B(n_71),
.Y(n_125)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_21),
.Y(n_63)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_63),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_29),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_64),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_31),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_65),
.Y(n_145)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_31),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g172 ( 
.A(n_66),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_33),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g173 ( 
.A(n_67),
.Y(n_173)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_33),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g192 ( 
.A(n_68),
.Y(n_192)
);

BUFx2_ASAP7_75t_L g69 ( 
.A(n_45),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g142 ( 
.A(n_69),
.Y(n_142)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_49),
.Y(n_70)
);

INVx3_ASAP7_75t_L g131 ( 
.A(n_70),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_45),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_44),
.Y(n_72)
);

INVx6_ASAP7_75t_L g129 ( 
.A(n_72),
.Y(n_129)
);

INVx13_ASAP7_75t_L g73 ( 
.A(n_45),
.Y(n_73)
);

INVx13_ASAP7_75t_L g153 ( 
.A(n_73),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_45),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_74),
.B(n_93),
.Y(n_140)
);

HB1xp67_ASAP7_75t_L g75 ( 
.A(n_24),
.Y(n_75)
);

CKINVDCx16_ASAP7_75t_R g183 ( 
.A(n_75),
.Y(n_183)
);

BUFx12f_ASAP7_75t_L g76 ( 
.A(n_49),
.Y(n_76)
);

BUFx3_ASAP7_75t_L g146 ( 
.A(n_76),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_44),
.Y(n_77)
);

INVx6_ASAP7_75t_L g148 ( 
.A(n_77),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_42),
.B(n_15),
.Y(n_78)
);

INVx11_ASAP7_75t_L g79 ( 
.A(n_20),
.Y(n_79)
);

INVx11_ASAP7_75t_L g143 ( 
.A(n_79),
.Y(n_143)
);

BUFx4f_ASAP7_75t_SL g80 ( 
.A(n_25),
.Y(n_80)
);

INVxp67_ASAP7_75t_SL g124 ( 
.A(n_80),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_32),
.B(n_14),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_81),
.B(n_88),
.Y(n_138)
);

BUFx3_ASAP7_75t_L g82 ( 
.A(n_25),
.Y(n_82)
);

BUFx12f_ASAP7_75t_L g128 ( 
.A(n_82),
.Y(n_128)
);

BUFx6f_ASAP7_75t_SL g83 ( 
.A(n_20),
.Y(n_83)
);

INVx11_ASAP7_75t_L g188 ( 
.A(n_83),
.Y(n_188)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_54),
.Y(n_84)
);

INVx6_ASAP7_75t_L g154 ( 
.A(n_84),
.Y(n_154)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_21),
.Y(n_85)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_85),
.Y(n_149)
);

BUFx3_ASAP7_75t_L g86 ( 
.A(n_28),
.Y(n_86)
);

BUFx3_ASAP7_75t_L g155 ( 
.A(n_86),
.Y(n_155)
);

INVx2_ASAP7_75t_SL g87 ( 
.A(n_28),
.Y(n_87)
);

INVx4_ASAP7_75t_SL g132 ( 
.A(n_87),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_32),
.B(n_0),
.Y(n_88)
);

BUFx12_ASAP7_75t_L g89 ( 
.A(n_49),
.Y(n_89)
);

BUFx12_ASAP7_75t_L g130 ( 
.A(n_89),
.Y(n_130)
);

BUFx3_ASAP7_75t_L g90 ( 
.A(n_43),
.Y(n_90)
);

INVx5_ASAP7_75t_L g161 ( 
.A(n_90),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_54),
.Y(n_91)
);

INVx6_ASAP7_75t_L g166 ( 
.A(n_91),
.Y(n_166)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_49),
.Y(n_92)
);

INVx3_ASAP7_75t_L g177 ( 
.A(n_92),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_53),
.Y(n_93)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_23),
.Y(n_94)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_94),
.Y(n_165)
);

BUFx5_ASAP7_75t_L g95 ( 
.A(n_43),
.Y(n_95)
);

BUFx2_ASAP7_75t_L g197 ( 
.A(n_95),
.Y(n_197)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_56),
.Y(n_96)
);

INVx8_ASAP7_75t_L g167 ( 
.A(n_96),
.Y(n_167)
);

INVx5_ASAP7_75t_L g97 ( 
.A(n_32),
.Y(n_97)
);

INVx4_ASAP7_75t_L g144 ( 
.A(n_97),
.Y(n_144)
);

INVx11_ASAP7_75t_L g98 ( 
.A(n_20),
.Y(n_98)
);

INVx11_ASAP7_75t_L g189 ( 
.A(n_98),
.Y(n_189)
);

BUFx12f_ASAP7_75t_L g99 ( 
.A(n_20),
.Y(n_99)
);

INVx4_ASAP7_75t_L g171 ( 
.A(n_99),
.Y(n_171)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_40),
.Y(n_100)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_100),
.Y(n_152)
);

AND2x2_ASAP7_75t_L g101 ( 
.A(n_27),
.B(n_0),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_101),
.B(n_105),
.Y(n_141)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_32),
.Y(n_102)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_102),
.Y(n_123)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_23),
.Y(n_103)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_103),
.Y(n_182)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_18),
.Y(n_104)
);

INVx3_ASAP7_75t_L g134 ( 
.A(n_104),
.Y(n_134)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_30),
.Y(n_105)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_40),
.Y(n_106)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_106),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_53),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_107),
.B(n_111),
.Y(n_159)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_18),
.Y(n_108)
);

INVx4_ASAP7_75t_L g181 ( 
.A(n_108),
.Y(n_181)
);

INVx8_ASAP7_75t_L g109 ( 
.A(n_56),
.Y(n_109)
);

INVx3_ASAP7_75t_SL g169 ( 
.A(n_109),
.Y(n_169)
);

INVx5_ASAP7_75t_L g110 ( 
.A(n_19),
.Y(n_110)
);

INVx4_ASAP7_75t_L g186 ( 
.A(n_110),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_53),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_57),
.Y(n_112)
);

INVx8_ASAP7_75t_L g187 ( 
.A(n_112),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_27),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_113),
.B(n_114),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_22),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_57),
.Y(n_115)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_115),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_22),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_116),
.B(n_50),
.Y(n_178)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_19),
.Y(n_117)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_117),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_57),
.Y(n_118)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_118),
.Y(n_174)
);

BUFx5_ASAP7_75t_L g119 ( 
.A(n_52),
.Y(n_119)
);

BUFx10_ASAP7_75t_L g193 ( 
.A(n_119),
.Y(n_193)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_38),
.Y(n_120)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_120),
.Y(n_175)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_38),
.Y(n_121)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_121),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_62),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_SL g208 ( 
.A(n_122),
.B(n_133),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_SL g133 ( 
.A(n_101),
.B(n_26),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_70),
.B(n_34),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_139),
.B(n_150),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_104),
.B(n_26),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_108),
.B(n_55),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_151),
.B(n_184),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_66),
.A2(n_55),
.B1(n_51),
.B2(n_34),
.Y(n_156)
);

OAI22xp33_ASAP7_75t_SL g229 ( 
.A1(n_156),
.A2(n_180),
.B1(n_96),
.B2(n_91),
.Y(n_229)
);

AOI21xp33_ASAP7_75t_SL g158 ( 
.A1(n_79),
.A2(n_24),
.B(n_52),
.Y(n_158)
);

OR2x2_ASAP7_75t_SL g212 ( 
.A(n_158),
.B(n_73),
.Y(n_212)
);

AOI22xp33_ASAP7_75t_L g160 ( 
.A1(n_112),
.A2(n_30),
.B1(n_36),
.B2(n_46),
.Y(n_160)
);

OA22x2_ASAP7_75t_L g244 ( 
.A1(n_160),
.A2(n_77),
.B1(n_67),
.B2(n_65),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_98),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_SL g253 ( 
.A(n_162),
.B(n_168),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_89),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_178),
.B(n_196),
.Y(n_203)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_102),
.Y(n_179)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_179),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_115),
.A2(n_37),
.B1(n_51),
.B2(n_41),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_110),
.B(n_41),
.Y(n_184)
);

CKINVDCx12_ASAP7_75t_R g185 ( 
.A(n_89),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_185),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_SL g190 ( 
.A(n_80),
.B(n_37),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_SL g263 ( 
.A(n_190),
.B(n_194),
.Y(n_263)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_118),
.Y(n_191)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_191),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_SL g194 ( 
.A(n_80),
.B(n_48),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_87),
.B(n_48),
.C(n_46),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_195),
.B(n_69),
.C(n_124),
.Y(n_206)
);

OR2x2_ASAP7_75t_L g196 ( 
.A(n_92),
.B(n_36),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_141),
.B(n_1),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_198),
.B(n_236),
.Y(n_276)
);

BUFx6f_ASAP7_75t_L g199 ( 
.A(n_127),
.Y(n_199)
);

BUFx6f_ASAP7_75t_L g298 ( 
.A(n_199),
.Y(n_298)
);

AND2x2_ASAP7_75t_SL g202 ( 
.A(n_137),
.B(n_99),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_202),
.B(n_206),
.C(n_210),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_125),
.B(n_97),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_SL g290 ( 
.A(n_204),
.B(n_205),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_138),
.B(n_121),
.Y(n_205)
);

AOI22xp33_ASAP7_75t_SL g207 ( 
.A1(n_124),
.A2(n_76),
.B1(n_99),
.B2(n_109),
.Y(n_207)
);

INVxp67_ASAP7_75t_L g291 ( 
.A(n_207),
.Y(n_291)
);

AND2x2_ASAP7_75t_L g209 ( 
.A(n_132),
.B(n_76),
.Y(n_209)
);

INVx1_ASAP7_75t_SL g275 ( 
.A(n_209),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_126),
.B(n_120),
.C(n_64),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_135),
.B(n_50),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_211),
.B(n_226),
.Y(n_268)
);

NOR2x1_ASAP7_75t_L g285 ( 
.A(n_212),
.B(n_264),
.Y(n_285)
);

INVx6_ASAP7_75t_L g213 ( 
.A(n_129),
.Y(n_213)
);

INVx4_ASAP7_75t_L g280 ( 
.A(n_213),
.Y(n_280)
);

BUFx2_ASAP7_75t_L g214 ( 
.A(n_171),
.Y(n_214)
);

BUFx3_ASAP7_75t_L g277 ( 
.A(n_214),
.Y(n_277)
);

INVx13_ASAP7_75t_L g215 ( 
.A(n_153),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_215),
.Y(n_295)
);

AOI22xp33_ASAP7_75t_SL g217 ( 
.A1(n_197),
.A2(n_82),
.B1(n_86),
.B2(n_90),
.Y(n_217)
);

AOI22xp33_ASAP7_75t_SL g283 ( 
.A1(n_217),
.A2(n_248),
.B1(n_254),
.B2(n_262),
.Y(n_283)
);

AND2x2_ASAP7_75t_L g220 ( 
.A(n_132),
.B(n_119),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_220),
.B(n_234),
.C(n_193),
.Y(n_281)
);

BUFx6f_ASAP7_75t_SL g221 ( 
.A(n_143),
.Y(n_221)
);

INVx4_ASAP7_75t_L g293 ( 
.A(n_221),
.Y(n_293)
);

INVx8_ASAP7_75t_L g222 ( 
.A(n_127),
.Y(n_222)
);

INVx3_ASAP7_75t_L g271 ( 
.A(n_222),
.Y(n_271)
);

INVx3_ASAP7_75t_L g223 ( 
.A(n_142),
.Y(n_223)
);

INVx4_ASAP7_75t_L g316 ( 
.A(n_223),
.Y(n_316)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_163),
.Y(n_224)
);

INVx2_ASAP7_75t_L g297 ( 
.A(n_224),
.Y(n_297)
);

INVx2_ASAP7_75t_SL g225 ( 
.A(n_142),
.Y(n_225)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_225),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_140),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_149),
.B(n_165),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_227),
.B(n_228),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_159),
.B(n_39),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_SL g304 ( 
.A1(n_229),
.A2(n_148),
.B1(n_234),
.B2(n_173),
.Y(n_304)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_174),
.Y(n_230)
);

INVx2_ASAP7_75t_L g299 ( 
.A(n_230),
.Y(n_299)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_175),
.Y(n_231)
);

INVx2_ASAP7_75t_L g313 ( 
.A(n_231),
.Y(n_313)
);

CKINVDCx16_ASAP7_75t_R g232 ( 
.A(n_143),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_232),
.B(n_241),
.Y(n_273)
);

BUFx3_ASAP7_75t_L g233 ( 
.A(n_146),
.Y(n_233)
);

INVx3_ASAP7_75t_L g287 ( 
.A(n_233),
.Y(n_287)
);

AND2x2_ASAP7_75t_SL g234 ( 
.A(n_147),
.B(n_95),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_182),
.Y(n_235)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_235),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_196),
.B(n_1),
.Y(n_236)
);

BUFx6f_ASAP7_75t_L g237 ( 
.A(n_136),
.Y(n_237)
);

INVx3_ASAP7_75t_L g302 ( 
.A(n_237),
.Y(n_302)
);

BUFx3_ASAP7_75t_L g238 ( 
.A(n_146),
.Y(n_238)
);

INVx3_ASAP7_75t_L g308 ( 
.A(n_238),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_152),
.B(n_2),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_239),
.B(n_246),
.Y(n_307)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_176),
.Y(n_240)
);

INVx2_ASAP7_75t_L g315 ( 
.A(n_240),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_183),
.B(n_39),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_170),
.B(n_157),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_242),
.B(n_250),
.Y(n_279)
);

BUFx6f_ASAP7_75t_L g243 ( 
.A(n_136),
.Y(n_243)
);

INVx3_ASAP7_75t_L g311 ( 
.A(n_243),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_L g300 ( 
.A1(n_244),
.A2(n_148),
.B1(n_166),
.B2(n_154),
.Y(n_300)
);

INVx4_ASAP7_75t_L g245 ( 
.A(n_144),
.Y(n_245)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_245),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_164),
.B(n_2),
.Y(n_246)
);

BUFx6f_ASAP7_75t_L g247 ( 
.A(n_145),
.Y(n_247)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_247),
.Y(n_305)
);

AOI22xp33_ASAP7_75t_SL g248 ( 
.A1(n_197),
.A2(n_84),
.B1(n_72),
.B2(n_68),
.Y(n_248)
);

INVx3_ASAP7_75t_L g249 ( 
.A(n_144),
.Y(n_249)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_249),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_131),
.B(n_61),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_188),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_251),
.B(n_252),
.Y(n_286)
);

INVx6_ASAP7_75t_L g252 ( 
.A(n_129),
.Y(n_252)
);

BUFx6f_ASAP7_75t_L g254 ( 
.A(n_145),
.Y(n_254)
);

INVx5_ASAP7_75t_L g255 ( 
.A(n_171),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_255),
.B(n_256),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_SL g256 ( 
.A(n_177),
.B(n_2),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_123),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_257),
.B(n_265),
.Y(n_296)
);

INVx3_ASAP7_75t_L g258 ( 
.A(n_123),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g306 ( 
.A(n_258),
.Y(n_306)
);

AOI22xp33_ASAP7_75t_L g259 ( 
.A1(n_160),
.A2(n_52),
.B1(n_4),
.B2(n_5),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_L g269 ( 
.A1(n_259),
.A2(n_261),
.B1(n_169),
.B2(n_188),
.Y(n_269)
);

INVx11_ASAP7_75t_L g260 ( 
.A(n_189),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_260),
.Y(n_310)
);

AOI22xp33_ASAP7_75t_L g261 ( 
.A1(n_167),
.A2(n_52),
.B1(n_7),
.B2(n_8),
.Y(n_261)
);

AOI22xp33_ASAP7_75t_SL g262 ( 
.A1(n_169),
.A2(n_3),
.B1(n_7),
.B2(n_8),
.Y(n_262)
);

CKINVDCx9p33_ASAP7_75t_R g264 ( 
.A(n_153),
.Y(n_264)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_172),
.Y(n_265)
);

BUFx3_ASAP7_75t_L g266 ( 
.A(n_128),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_266),
.B(n_128),
.Y(n_314)
);

AND2x2_ASAP7_75t_L g348 ( 
.A(n_269),
.B(n_281),
.Y(n_348)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_212),
.A2(n_172),
.B1(n_166),
.B2(n_154),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g326 ( 
.A1(n_272),
.A2(n_309),
.B1(n_321),
.B2(n_202),
.Y(n_326)
);

AND2x2_ASAP7_75t_SL g284 ( 
.A(n_206),
.B(n_193),
.Y(n_284)
);

AND2x2_ASAP7_75t_L g361 ( 
.A(n_284),
.B(n_238),
.Y(n_361)
);

AOI22xp33_ASAP7_75t_SL g288 ( 
.A1(n_236),
.A2(n_193),
.B1(n_161),
.B2(n_155),
.Y(n_288)
);

INVxp67_ASAP7_75t_L g354 ( 
.A(n_288),
.Y(n_354)
);

OAI21xp5_ASAP7_75t_L g292 ( 
.A1(n_203),
.A2(n_155),
.B(n_134),
.Y(n_292)
);

AOI21xp5_ASAP7_75t_L g332 ( 
.A1(n_292),
.A2(n_294),
.B(n_303),
.Y(n_332)
);

AOI21xp5_ASAP7_75t_L g294 ( 
.A1(n_220),
.A2(n_189),
.B(n_161),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_L g323 ( 
.A1(n_300),
.A2(n_304),
.B1(n_222),
.B2(n_213),
.Y(n_323)
);

NOR2x1_ASAP7_75t_L g301 ( 
.A(n_208),
.B(n_181),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_SL g333 ( 
.A(n_301),
.B(n_317),
.Y(n_333)
);

AOI21xp5_ASAP7_75t_L g303 ( 
.A1(n_220),
.A2(n_209),
.B(n_253),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_SL g309 ( 
.A1(n_200),
.A2(n_192),
.B1(n_173),
.B2(n_167),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_239),
.B(n_187),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_312),
.B(n_319),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_314),
.B(n_264),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_263),
.B(n_181),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_246),
.B(n_187),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_201),
.B(n_134),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_SL g342 ( 
.A(n_320),
.B(n_214),
.Y(n_342)
);

OAI22xp5_ASAP7_75t_L g321 ( 
.A1(n_244),
.A2(n_192),
.B1(n_186),
.B2(n_128),
.Y(n_321)
);

AOI21xp5_ASAP7_75t_L g322 ( 
.A1(n_209),
.A2(n_186),
.B(n_130),
.Y(n_322)
);

OAI21xp5_ASAP7_75t_SL g353 ( 
.A1(n_322),
.A2(n_225),
.B(n_130),
.Y(n_353)
);

AOI22xp5_ASAP7_75t_L g387 ( 
.A1(n_323),
.A2(n_324),
.B1(n_338),
.B2(n_306),
.Y(n_387)
);

OAI22xp5_ASAP7_75t_L g324 ( 
.A1(n_304),
.A2(n_244),
.B1(n_210),
.B2(n_198),
.Y(n_324)
);

AND2x6_ASAP7_75t_L g325 ( 
.A(n_284),
.B(n_218),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_SL g395 ( 
.A(n_325),
.B(n_345),
.Y(n_395)
);

OAI22xp5_ASAP7_75t_L g376 ( 
.A1(n_326),
.A2(n_328),
.B1(n_329),
.B2(n_339),
.Y(n_376)
);

AOI22xp5_ASAP7_75t_L g328 ( 
.A1(n_272),
.A2(n_244),
.B1(n_234),
.B2(n_202),
.Y(n_328)
);

AOI22xp5_ASAP7_75t_L g329 ( 
.A1(n_284),
.A2(n_265),
.B1(n_252),
.B2(n_240),
.Y(n_329)
);

INVx3_ASAP7_75t_L g330 ( 
.A(n_271),
.Y(n_330)
);

INVx2_ASAP7_75t_L g377 ( 
.A(n_330),
.Y(n_377)
);

INVxp67_ASAP7_75t_L g393 ( 
.A(n_331),
.Y(n_393)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_301),
.B(n_218),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g381 ( 
.A(n_334),
.B(n_342),
.Y(n_381)
);

INVx6_ASAP7_75t_L g335 ( 
.A(n_298),
.Y(n_335)
);

HB1xp67_ASAP7_75t_L g366 ( 
.A(n_335),
.Y(n_366)
);

A2O1A1Ixp33_ASAP7_75t_L g336 ( 
.A1(n_278),
.A2(n_215),
.B(n_216),
.C(n_219),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_336),
.B(n_355),
.Y(n_371)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_274),
.Y(n_337)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_337),
.Y(n_368)
);

OAI22xp5_ASAP7_75t_SL g338 ( 
.A1(n_300),
.A2(n_231),
.B1(n_230),
.B2(n_224),
.Y(n_338)
);

AOI22xp5_ASAP7_75t_L g339 ( 
.A1(n_309),
.A2(n_258),
.B1(n_199),
.B2(n_243),
.Y(n_339)
);

BUFx12_ASAP7_75t_L g340 ( 
.A(n_295),
.Y(n_340)
);

CKINVDCx20_ASAP7_75t_R g389 ( 
.A(n_340),
.Y(n_389)
);

INVx3_ASAP7_75t_L g341 ( 
.A(n_271),
.Y(n_341)
);

INVx1_ASAP7_75t_SL g402 ( 
.A(n_341),
.Y(n_402)
);

XOR2xp5_ASAP7_75t_L g343 ( 
.A(n_307),
.B(n_260),
.Y(n_343)
);

XNOR2xp5_ASAP7_75t_L g370 ( 
.A(n_343),
.B(n_358),
.Y(n_370)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_274),
.Y(n_344)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_344),
.Y(n_378)
);

AND2x6_ASAP7_75t_L g345 ( 
.A(n_290),
.B(n_221),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_296),
.Y(n_346)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_346),
.Y(n_382)
);

INVx5_ASAP7_75t_L g347 ( 
.A(n_280),
.Y(n_347)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_347),
.Y(n_390)
);

INVx3_ASAP7_75t_L g349 ( 
.A(n_280),
.Y(n_349)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_349),
.Y(n_394)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_297),
.Y(n_350)
);

AOI22xp33_ASAP7_75t_SL g391 ( 
.A1(n_350),
.A2(n_351),
.B1(n_363),
.B2(n_365),
.Y(n_391)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_297),
.Y(n_351)
);

NOR2xp33_ASAP7_75t_L g352 ( 
.A(n_268),
.B(n_279),
.Y(n_352)
);

CKINVDCx16_ASAP7_75t_R g374 ( 
.A(n_352),
.Y(n_374)
);

OAI21xp5_ASAP7_75t_SL g388 ( 
.A1(n_353),
.A2(n_356),
.B(n_359),
.Y(n_388)
);

AND2x6_ASAP7_75t_L g355 ( 
.A(n_285),
.B(n_130),
.Y(n_355)
);

NAND2x1_ASAP7_75t_L g356 ( 
.A(n_285),
.B(n_245),
.Y(n_356)
);

OAI22xp33_ASAP7_75t_SL g357 ( 
.A1(n_283),
.A2(n_249),
.B1(n_254),
.B2(n_247),
.Y(n_357)
);

AOI22xp5_ASAP7_75t_SL g375 ( 
.A1(n_357),
.A2(n_291),
.B1(n_275),
.B2(n_310),
.Y(n_375)
);

MAJIxp5_ASAP7_75t_L g358 ( 
.A(n_278),
.B(n_223),
.C(n_237),
.Y(n_358)
);

OR2x2_ASAP7_75t_L g359 ( 
.A(n_281),
.B(n_255),
.Y(n_359)
);

AND2x6_ASAP7_75t_L g360 ( 
.A(n_292),
.B(n_266),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_360),
.B(n_362),
.Y(n_372)
);

XOR2xp5_ASAP7_75t_L g386 ( 
.A(n_361),
.B(n_318),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g362 ( 
.A(n_307),
.B(n_319),
.Y(n_362)
);

INVx13_ASAP7_75t_L g363 ( 
.A(n_295),
.Y(n_363)
);

AND2x2_ASAP7_75t_L g364 ( 
.A(n_275),
.B(n_233),
.Y(n_364)
);

OAI21xp5_ASAP7_75t_L g385 ( 
.A1(n_364),
.A2(n_294),
.B(n_306),
.Y(n_385)
);

INVx5_ASAP7_75t_L g365 ( 
.A(n_302),
.Y(n_365)
);

OAI22xp5_ASAP7_75t_SL g367 ( 
.A1(n_326),
.A2(n_312),
.B1(n_289),
.B2(n_291),
.Y(n_367)
);

AOI22xp5_ASAP7_75t_L g406 ( 
.A1(n_367),
.A2(n_383),
.B1(n_401),
.B2(n_403),
.Y(n_406)
);

BUFx24_ASAP7_75t_SL g369 ( 
.A(n_333),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_L g407 ( 
.A(n_369),
.B(n_364),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_362),
.B(n_286),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_373),
.B(n_379),
.Y(n_413)
);

OAI22xp5_ASAP7_75t_L g404 ( 
.A1(n_375),
.A2(n_329),
.B1(n_353),
.B2(n_339),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_327),
.B(n_276),
.Y(n_379)
);

AOI21xp5_ASAP7_75t_L g380 ( 
.A1(n_354),
.A2(n_322),
.B(n_303),
.Y(n_380)
);

AOI21xp5_ASAP7_75t_L g433 ( 
.A1(n_380),
.A2(n_399),
.B(n_385),
.Y(n_433)
);

OAI22xp5_ASAP7_75t_SL g383 ( 
.A1(n_328),
.A2(n_270),
.B1(n_273),
.B2(n_276),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_343),
.B(n_310),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_384),
.B(n_398),
.Y(n_428)
);

AND2x2_ASAP7_75t_L g425 ( 
.A(n_385),
.B(n_387),
.Y(n_425)
);

INVxp67_ASAP7_75t_L g414 ( 
.A(n_386),
.Y(n_414)
);

OAI21xp5_ASAP7_75t_L g392 ( 
.A1(n_356),
.A2(n_267),
.B(n_318),
.Y(n_392)
);

AO21x1_ASAP7_75t_L g429 ( 
.A1(n_392),
.A2(n_396),
.B(n_397),
.Y(n_429)
);

OAI21xp5_ASAP7_75t_L g396 ( 
.A1(n_332),
.A2(n_267),
.B(n_282),
.Y(n_396)
);

OAI21xp5_ASAP7_75t_L g397 ( 
.A1(n_332),
.A2(n_282),
.B(n_287),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_358),
.B(n_336),
.Y(n_398)
);

OAI21xp5_ASAP7_75t_L g399 ( 
.A1(n_354),
.A2(n_287),
.B(n_308),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_348),
.B(n_305),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_400),
.B(n_349),
.Y(n_430)
);

OAI22xp5_ASAP7_75t_SL g401 ( 
.A1(n_359),
.A2(n_305),
.B1(n_311),
.B2(n_302),
.Y(n_401)
);

OAI22xp5_ASAP7_75t_SL g403 ( 
.A1(n_348),
.A2(n_311),
.B1(n_298),
.B2(n_313),
.Y(n_403)
);

AOI22xp5_ASAP7_75t_L g440 ( 
.A1(n_404),
.A2(n_410),
.B1(n_423),
.B2(n_431),
.Y(n_440)
);

CKINVDCx20_ASAP7_75t_R g405 ( 
.A(n_366),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_405),
.B(n_422),
.Y(n_443)
);

INVxp67_ASAP7_75t_L g450 ( 
.A(n_407),
.Y(n_450)
);

NOR2xp33_ASAP7_75t_SL g408 ( 
.A(n_381),
.B(n_361),
.Y(n_408)
);

NOR2xp33_ASAP7_75t_SL g452 ( 
.A(n_408),
.B(n_416),
.Y(n_452)
);

MAJIxp5_ASAP7_75t_L g409 ( 
.A(n_370),
.B(n_361),
.C(n_348),
.Y(n_409)
);

MAJIxp5_ASAP7_75t_L g445 ( 
.A(n_409),
.B(n_412),
.C(n_432),
.Y(n_445)
);

OAI22xp5_ASAP7_75t_SL g410 ( 
.A1(n_387),
.A2(n_345),
.B1(n_325),
.B2(n_360),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_368),
.Y(n_411)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_411),
.Y(n_444)
);

XOR2xp5_ASAP7_75t_L g412 ( 
.A(n_370),
.B(n_364),
.Y(n_412)
);

AOI22xp5_ASAP7_75t_L g415 ( 
.A1(n_376),
.A2(n_338),
.B1(n_355),
.B2(n_330),
.Y(n_415)
);

OAI22xp5_ASAP7_75t_L g442 ( 
.A1(n_415),
.A2(n_375),
.B1(n_396),
.B2(n_395),
.Y(n_442)
);

NOR2xp33_ASAP7_75t_L g416 ( 
.A(n_389),
.B(n_341),
.Y(n_416)
);

NOR2xp33_ASAP7_75t_L g417 ( 
.A(n_389),
.B(n_382),
.Y(n_417)
);

CKINVDCx14_ASAP7_75t_R g460 ( 
.A(n_417),
.Y(n_460)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_368),
.Y(n_418)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_418),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_SL g419 ( 
.A(n_373),
.B(n_340),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_SL g441 ( 
.A(n_419),
.B(n_420),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_SL g420 ( 
.A(n_379),
.B(n_340),
.Y(n_420)
);

NOR2xp33_ASAP7_75t_L g421 ( 
.A(n_382),
.B(n_365),
.Y(n_421)
);

NOR3xp33_ASAP7_75t_L g449 ( 
.A(n_421),
.B(n_390),
.C(n_394),
.Y(n_449)
);

CKINVDCx20_ASAP7_75t_R g422 ( 
.A(n_381),
.Y(n_422)
);

OAI22xp5_ASAP7_75t_L g423 ( 
.A1(n_372),
.A2(n_395),
.B1(n_371),
.B2(n_400),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_378),
.Y(n_424)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_424),
.Y(n_461)
);

CKINVDCx20_ASAP7_75t_R g426 ( 
.A(n_401),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g446 ( 
.A(n_426),
.B(n_436),
.Y(n_446)
);

NOR2xp33_ASAP7_75t_L g427 ( 
.A(n_383),
.B(n_316),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_SL g453 ( 
.A(n_427),
.B(n_374),
.Y(n_453)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_430),
.Y(n_463)
);

OAI22xp5_ASAP7_75t_L g431 ( 
.A1(n_372),
.A2(n_335),
.B1(n_363),
.B2(n_347),
.Y(n_431)
);

MAJIxp5_ASAP7_75t_L g432 ( 
.A(n_398),
.B(n_384),
.C(n_386),
.Y(n_432)
);

OAI21xp5_ASAP7_75t_L g439 ( 
.A1(n_433),
.A2(n_388),
.B(n_380),
.Y(n_439)
);

XOR2xp5_ASAP7_75t_L g434 ( 
.A(n_388),
.B(n_316),
.Y(n_434)
);

MAJIxp5_ASAP7_75t_L g454 ( 
.A(n_434),
.B(n_412),
.C(n_409),
.Y(n_454)
);

NAND4xp25_ASAP7_75t_SL g435 ( 
.A(n_371),
.B(n_277),
.C(n_308),
.D(n_293),
.Y(n_435)
);

CKINVDCx20_ASAP7_75t_R g456 ( 
.A(n_435),
.Y(n_456)
);

CKINVDCx20_ASAP7_75t_R g436 ( 
.A(n_378),
.Y(n_436)
);

CKINVDCx20_ASAP7_75t_R g437 ( 
.A(n_374),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_L g455 ( 
.A(n_437),
.B(n_438),
.Y(n_455)
);

INVxp67_ASAP7_75t_L g438 ( 
.A(n_392),
.Y(n_438)
);

OAI21xp5_ASAP7_75t_L g493 ( 
.A1(n_439),
.A2(n_435),
.B(n_411),
.Y(n_493)
);

AOI22xp5_ASAP7_75t_L g485 ( 
.A1(n_442),
.A2(n_466),
.B1(n_404),
.B2(n_425),
.Y(n_485)
);

AOI22xp5_ASAP7_75t_L g447 ( 
.A1(n_431),
.A2(n_376),
.B1(n_367),
.B2(n_403),
.Y(n_447)
);

OAI22xp5_ASAP7_75t_SL g484 ( 
.A1(n_447),
.A2(n_448),
.B1(n_429),
.B2(n_428),
.Y(n_484)
);

AOI22xp5_ASAP7_75t_L g448 ( 
.A1(n_426),
.A2(n_397),
.B1(n_399),
.B2(n_393),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_L g481 ( 
.A(n_449),
.B(n_451),
.Y(n_481)
);

OA22x2_ASAP7_75t_L g451 ( 
.A1(n_406),
.A2(n_377),
.B1(n_402),
.B2(n_394),
.Y(n_451)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_453),
.Y(n_471)
);

MAJx2_ASAP7_75t_L g495 ( 
.A(n_454),
.B(n_299),
.C(n_293),
.Y(n_495)
);

CKINVDCx20_ASAP7_75t_R g458 ( 
.A(n_417),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_L g490 ( 
.A(n_458),
.B(n_459),
.Y(n_490)
);

CKINVDCx20_ASAP7_75t_R g459 ( 
.A(n_416),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_SL g462 ( 
.A(n_422),
.B(n_390),
.Y(n_462)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_462),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_L g464 ( 
.A(n_420),
.B(n_377),
.Y(n_464)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_464),
.Y(n_474)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_419),
.Y(n_465)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_465),
.Y(n_491)
);

OAI22xp5_ASAP7_75t_L g466 ( 
.A1(n_415),
.A2(n_391),
.B1(n_402),
.B2(n_277),
.Y(n_466)
);

XOR2xp5_ASAP7_75t_L g467 ( 
.A(n_432),
.B(n_315),
.Y(n_467)
);

XOR2xp5_ASAP7_75t_L g488 ( 
.A(n_467),
.B(n_425),
.Y(n_488)
);

CKINVDCx16_ASAP7_75t_R g468 ( 
.A(n_430),
.Y(n_468)
);

NOR2xp33_ASAP7_75t_L g475 ( 
.A(n_468),
.B(n_437),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_413),
.B(n_315),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_469),
.Y(n_470)
);

MAJIxp5_ASAP7_75t_SL g473 ( 
.A(n_439),
.B(n_425),
.C(n_408),
.Y(n_473)
);

OAI21xp5_ASAP7_75t_SL g500 ( 
.A1(n_473),
.A2(n_483),
.B(n_460),
.Y(n_500)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_475),
.Y(n_496)
);

INVx2_ASAP7_75t_L g476 ( 
.A(n_465),
.Y(n_476)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_476),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_SL g477 ( 
.A(n_450),
.B(n_413),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_SL g511 ( 
.A(n_477),
.B(n_482),
.Y(n_511)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_464),
.Y(n_478)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_478),
.Y(n_508)
);

OAI22x1_ASAP7_75t_L g479 ( 
.A1(n_448),
.A2(n_406),
.B1(n_429),
.B2(n_433),
.Y(n_479)
);

OAI22xp5_ASAP7_75t_L g505 ( 
.A1(n_479),
.A2(n_456),
.B1(n_446),
.B2(n_441),
.Y(n_505)
);

MAJIxp5_ASAP7_75t_L g480 ( 
.A(n_445),
.B(n_414),
.C(n_434),
.Y(n_480)
);

MAJIxp5_ASAP7_75t_L g498 ( 
.A(n_480),
.B(n_487),
.C(n_489),
.Y(n_498)
);

NOR2xp33_ASAP7_75t_L g482 ( 
.A(n_453),
.B(n_421),
.Y(n_482)
);

AOI21xp33_ASAP7_75t_L g483 ( 
.A1(n_455),
.A2(n_428),
.B(n_423),
.Y(n_483)
);

AOI22xp5_ASAP7_75t_L g507 ( 
.A1(n_484),
.A2(n_466),
.B1(n_463),
.B2(n_468),
.Y(n_507)
);

OAI22xp5_ASAP7_75t_SL g501 ( 
.A1(n_485),
.A2(n_440),
.B1(n_447),
.B2(n_446),
.Y(n_501)
);

OAI22xp5_ASAP7_75t_L g486 ( 
.A1(n_440),
.A2(n_429),
.B1(n_436),
.B2(n_405),
.Y(n_486)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_486),
.Y(n_515)
);

MAJIxp5_ASAP7_75t_L g487 ( 
.A(n_445),
.B(n_454),
.C(n_467),
.Y(n_487)
);

XNOR2xp5_ASAP7_75t_L g497 ( 
.A(n_488),
.B(n_495),
.Y(n_497)
);

MAJIxp5_ASAP7_75t_L g489 ( 
.A(n_443),
.B(n_410),
.C(n_424),
.Y(n_489)
);

NOR2xp33_ASAP7_75t_L g492 ( 
.A(n_458),
.B(n_418),
.Y(n_492)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_492),
.Y(n_517)
);

XOR2xp5_ASAP7_75t_L g514 ( 
.A(n_493),
.B(n_461),
.Y(n_514)
);

XNOR2xp5_ASAP7_75t_SL g494 ( 
.A(n_441),
.B(n_313),
.Y(n_494)
);

XNOR2xp5_ASAP7_75t_SL g512 ( 
.A(n_494),
.B(n_461),
.Y(n_512)
);

MAJIxp5_ASAP7_75t_L g499 ( 
.A(n_487),
.B(n_443),
.C(n_459),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_499),
.B(n_502),
.Y(n_530)
);

INVxp67_ASAP7_75t_L g526 ( 
.A(n_500),
.Y(n_526)
);

AOI22xp5_ASAP7_75t_L g519 ( 
.A1(n_501),
.A2(n_505),
.B1(n_509),
.B2(n_491),
.Y(n_519)
);

MAJIxp5_ASAP7_75t_L g502 ( 
.A(n_480),
.B(n_455),
.C(n_462),
.Y(n_502)
);

CKINVDCx16_ASAP7_75t_R g503 ( 
.A(n_490),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_L g531 ( 
.A(n_503),
.B(n_504),
.Y(n_531)
);

MAJIxp5_ASAP7_75t_L g504 ( 
.A(n_488),
.B(n_442),
.C(n_451),
.Y(n_504)
);

OAI22xp5_ASAP7_75t_SL g522 ( 
.A1(n_507),
.A2(n_516),
.B1(n_476),
.B2(n_472),
.Y(n_522)
);

OAI22xp5_ASAP7_75t_SL g509 ( 
.A1(n_485),
.A2(n_456),
.B1(n_463),
.B2(n_452),
.Y(n_509)
);

XNOR2xp5_ASAP7_75t_L g510 ( 
.A(n_495),
.B(n_469),
.Y(n_510)
);

XNOR2xp5_ASAP7_75t_L g521 ( 
.A(n_510),
.B(n_514),
.Y(n_521)
);

XNOR2x1_ASAP7_75t_L g523 ( 
.A(n_512),
.B(n_513),
.Y(n_523)
);

XNOR2xp5_ASAP7_75t_SL g513 ( 
.A(n_479),
.B(n_452),
.Y(n_513)
);

AOI22xp5_ASAP7_75t_L g516 ( 
.A1(n_484),
.A2(n_451),
.B1(n_457),
.B2(n_444),
.Y(n_516)
);

MAJIxp5_ASAP7_75t_L g518 ( 
.A(n_489),
.B(n_451),
.C(n_457),
.Y(n_518)
);

NOR2xp33_ASAP7_75t_L g532 ( 
.A(n_518),
.B(n_490),
.Y(n_532)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_519),
.Y(n_543)
);

XOR2xp5_ASAP7_75t_L g520 ( 
.A(n_497),
.B(n_493),
.Y(n_520)
);

XOR2xp5_ASAP7_75t_L g540 ( 
.A(n_520),
.B(n_536),
.Y(n_540)
);

AOI22xp5_ASAP7_75t_L g538 ( 
.A1(n_522),
.A2(n_501),
.B1(n_508),
.B2(n_518),
.Y(n_538)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_509),
.Y(n_524)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_524),
.Y(n_546)
);

CKINVDCx20_ASAP7_75t_R g525 ( 
.A(n_511),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_L g541 ( 
.A(n_525),
.B(n_528),
.Y(n_541)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_517),
.Y(n_527)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_527),
.Y(n_549)
);

XNOR2xp5_ASAP7_75t_L g528 ( 
.A(n_498),
.B(n_473),
.Y(n_528)
);

BUFx5_ASAP7_75t_L g529 ( 
.A(n_496),
.Y(n_529)
);

NOR2xp33_ASAP7_75t_L g545 ( 
.A(n_529),
.B(n_532),
.Y(n_545)
);

NOR2xp33_ASAP7_75t_L g533 ( 
.A(n_499),
.B(n_471),
.Y(n_533)
);

NOR2xp33_ASAP7_75t_L g550 ( 
.A(n_533),
.B(n_534),
.Y(n_550)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_506),
.Y(n_534)
);

NOR2xp33_ASAP7_75t_L g535 ( 
.A(n_502),
.B(n_481),
.Y(n_535)
);

NOR2xp33_ASAP7_75t_L g551 ( 
.A(n_535),
.B(n_510),
.Y(n_551)
);

XOR2xp5_ASAP7_75t_L g536 ( 
.A(n_497),
.B(n_481),
.Y(n_536)
);

AOI21xp5_ASAP7_75t_L g537 ( 
.A1(n_526),
.A2(n_515),
.B(n_514),
.Y(n_537)
);

AOI21xp5_ASAP7_75t_L g553 ( 
.A1(n_537),
.A2(n_542),
.B(n_544),
.Y(n_553)
);

XOR2xp5_ASAP7_75t_L g561 ( 
.A(n_538),
.B(n_539),
.Y(n_561)
);

AOI22xp5_ASAP7_75t_L g539 ( 
.A1(n_526),
.A2(n_504),
.B1(n_478),
.B2(n_474),
.Y(n_539)
);

MAJIxp5_ASAP7_75t_L g542 ( 
.A(n_530),
.B(n_498),
.C(n_513),
.Y(n_542)
);

OAI21xp5_ASAP7_75t_L g544 ( 
.A1(n_531),
.A2(n_507),
.B(n_470),
.Y(n_544)
);

AND2x2_ASAP7_75t_L g547 ( 
.A(n_519),
.B(n_516),
.Y(n_547)
);

XOR2xp5_ASAP7_75t_L g563 ( 
.A(n_547),
.B(n_538),
.Y(n_563)
);

OAI21xp5_ASAP7_75t_SL g548 ( 
.A1(n_528),
.A2(n_470),
.B(n_512),
.Y(n_548)
);

AOI21xp5_ASAP7_75t_SL g554 ( 
.A1(n_548),
.A2(n_537),
.B(n_544),
.Y(n_554)
);

NOR2xp33_ASAP7_75t_SL g558 ( 
.A(n_551),
.B(n_444),
.Y(n_558)
);

OAI21xp5_ASAP7_75t_SL g552 ( 
.A1(n_541),
.A2(n_529),
.B(n_536),
.Y(n_552)
);

AOI21xp5_ASAP7_75t_L g564 ( 
.A1(n_552),
.A2(n_557),
.B(n_560),
.Y(n_564)
);

INVxp67_ASAP7_75t_L g571 ( 
.A(n_554),
.Y(n_571)
);

MAJIxp5_ASAP7_75t_L g555 ( 
.A(n_542),
.B(n_521),
.C(n_520),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_L g570 ( 
.A(n_555),
.B(n_556),
.Y(n_570)
);

NOR2xp33_ASAP7_75t_L g556 ( 
.A(n_549),
.B(n_521),
.Y(n_556)
);

MAJIxp5_ASAP7_75t_L g557 ( 
.A(n_540),
.B(n_523),
.C(n_494),
.Y(n_557)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_558),
.Y(n_567)
);

NOR2xp33_ASAP7_75t_L g559 ( 
.A(n_543),
.B(n_299),
.Y(n_559)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_559),
.Y(n_568)
);

NOR2xp33_ASAP7_75t_L g560 ( 
.A(n_539),
.B(n_523),
.Y(n_560)
);

AOI22xp5_ASAP7_75t_L g562 ( 
.A1(n_546),
.A2(n_3),
.B1(n_7),
.B2(n_10),
.Y(n_562)
);

MAJIxp5_ASAP7_75t_L g565 ( 
.A(n_562),
.B(n_545),
.C(n_550),
.Y(n_565)
);

MAJIxp5_ASAP7_75t_L g572 ( 
.A(n_563),
.B(n_547),
.C(n_11),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_L g573 ( 
.A(n_565),
.B(n_561),
.Y(n_573)
);

AOI21xp5_ASAP7_75t_L g566 ( 
.A1(n_553),
.A2(n_548),
.B(n_540),
.Y(n_566)
);

AOI21x1_ASAP7_75t_L g577 ( 
.A1(n_566),
.A2(n_557),
.B(n_554),
.Y(n_577)
);

OA21x2_ASAP7_75t_SL g569 ( 
.A1(n_555),
.A2(n_547),
.B(n_10),
.Y(n_569)
);

CKINVDCx20_ASAP7_75t_R g578 ( 
.A(n_569),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_SL g576 ( 
.A(n_572),
.B(n_3),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_L g579 ( 
.A(n_573),
.B(n_574),
.Y(n_579)
);

CKINVDCx16_ASAP7_75t_R g574 ( 
.A(n_570),
.Y(n_574)
);

MAJIxp5_ASAP7_75t_L g575 ( 
.A(n_564),
.B(n_563),
.C(n_561),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_L g581 ( 
.A(n_575),
.B(n_576),
.Y(n_581)
);

AOI21xp5_ASAP7_75t_SL g580 ( 
.A1(n_577),
.A2(n_571),
.B(n_567),
.Y(n_580)
);

OAI21xp5_ASAP7_75t_L g583 ( 
.A1(n_580),
.A2(n_571),
.B(n_575),
.Y(n_583)
);

NOR2xp33_ASAP7_75t_L g582 ( 
.A(n_578),
.B(n_572),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_L g584 ( 
.A(n_582),
.B(n_568),
.Y(n_584)
);

OAI21xp33_ASAP7_75t_L g585 ( 
.A1(n_583),
.A2(n_584),
.B(n_579),
.Y(n_585)
);

OR2x2_ASAP7_75t_L g586 ( 
.A(n_585),
.B(n_581),
.Y(n_586)
);

OAI31xp33_ASAP7_75t_L g587 ( 
.A1(n_586),
.A2(n_12),
.A3(n_13),
.B(n_585),
.Y(n_587)
);

XNOR2xp5_ASAP7_75t_L g588 ( 
.A(n_587),
.B(n_12),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_SL g589 ( 
.A(n_588),
.B(n_12),
.Y(n_589)
);


endmodule