module fake_netlist_1_12642_n_719 (n_44, n_81, n_69, n_22, n_57, n_88, n_52, n_26, n_50, n_33, n_73, n_49, n_80, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_87, n_74, n_7, n_29, n_45, n_85, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_91, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_84, n_55, n_12, n_86, n_75, n_72, n_43, n_76, n_89, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_83, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_82, n_15, n_61, n_21, n_51, n_39, n_719);
input n_44;
input n_81;
input n_69;
input n_22;
input n_57;
input n_88;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_80;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_87;
input n_74;
input n_7;
input n_29;
input n_45;
input n_85;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_84;
input n_55;
input n_12;
input n_86;
input n_75;
input n_72;
input n_43;
input n_76;
input n_89;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_83;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_82;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_719;
wire n_117;
wire n_663;
wire n_707;
wire n_361;
wire n_513;
wire n_185;
wire n_705;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_701;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_672;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_715;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_702;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_563;
wire n_540;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_697;
wire n_554;
wire n_712;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_711;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_708;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_696;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_243;
wire n_235;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_338;
wire n_519;
wire n_699;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_689;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_704;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_710;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_706;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_357;
wire n_653;
wire n_716;
wire n_260;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_718;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_717;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_684;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_597;
wire n_498;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_714;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_618;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_688;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_266;
wire n_683;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_695;
wire n_469;
wire n_585;
wire n_713;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_709;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_132;
wire n_99;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
BUFx6f_ASAP7_75t_L g92 ( .A(n_69), .Y(n_92) );
INVx1_ASAP7_75t_L g93 ( .A(n_12), .Y(n_93) );
INVx1_ASAP7_75t_L g94 ( .A(n_33), .Y(n_94) );
BUFx6f_ASAP7_75t_L g95 ( .A(n_15), .Y(n_95) );
INVxp67_ASAP7_75t_SL g96 ( .A(n_79), .Y(n_96) );
BUFx6f_ASAP7_75t_L g97 ( .A(n_26), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_86), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_68), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_88), .Y(n_100) );
INVx2_ASAP7_75t_L g101 ( .A(n_41), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_82), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_67), .Y(n_103) );
CKINVDCx5p33_ASAP7_75t_R g104 ( .A(n_13), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_59), .Y(n_105) );
CKINVDCx16_ASAP7_75t_R g106 ( .A(n_37), .Y(n_106) );
CKINVDCx5p33_ASAP7_75t_R g107 ( .A(n_28), .Y(n_107) );
INVxp33_ASAP7_75t_L g108 ( .A(n_85), .Y(n_108) );
INVx1_ASAP7_75t_SL g109 ( .A(n_60), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_52), .Y(n_110) );
INVx2_ASAP7_75t_L g111 ( .A(n_42), .Y(n_111) );
CKINVDCx5p33_ASAP7_75t_R g112 ( .A(n_17), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_6), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_17), .Y(n_114) );
CKINVDCx5p33_ASAP7_75t_R g115 ( .A(n_2), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_54), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_65), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_62), .Y(n_118) );
CKINVDCx16_ASAP7_75t_R g119 ( .A(n_5), .Y(n_119) );
CKINVDCx14_ASAP7_75t_R g120 ( .A(n_5), .Y(n_120) );
INVx1_ASAP7_75t_SL g121 ( .A(n_83), .Y(n_121) );
CKINVDCx5p33_ASAP7_75t_R g122 ( .A(n_40), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_31), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_47), .Y(n_124) );
INVx1_ASAP7_75t_L g125 ( .A(n_35), .Y(n_125) );
INVx1_ASAP7_75t_L g126 ( .A(n_66), .Y(n_126) );
BUFx2_ASAP7_75t_L g127 ( .A(n_7), .Y(n_127) );
INVx1_ASAP7_75t_L g128 ( .A(n_36), .Y(n_128) );
HB1xp67_ASAP7_75t_L g129 ( .A(n_4), .Y(n_129) );
CKINVDCx20_ASAP7_75t_R g130 ( .A(n_55), .Y(n_130) );
INVxp67_ASAP7_75t_L g131 ( .A(n_29), .Y(n_131) );
INVx3_ASAP7_75t_L g132 ( .A(n_95), .Y(n_132) );
AND2x4_ASAP7_75t_L g133 ( .A(n_101), .B(n_0), .Y(n_133) );
INVx1_ASAP7_75t_L g134 ( .A(n_102), .Y(n_134) );
INVx1_ASAP7_75t_L g135 ( .A(n_102), .Y(n_135) );
OA21x2_ASAP7_75t_L g136 ( .A1(n_103), .A2(n_0), .B(n_1), .Y(n_136) );
INVx2_ASAP7_75t_L g137 ( .A(n_92), .Y(n_137) );
INVx1_ASAP7_75t_L g138 ( .A(n_103), .Y(n_138) );
INVx1_ASAP7_75t_L g139 ( .A(n_105), .Y(n_139) );
NOR2x1_ASAP7_75t_L g140 ( .A(n_94), .B(n_1), .Y(n_140) );
INVx1_ASAP7_75t_L g141 ( .A(n_105), .Y(n_141) );
AND2x4_ASAP7_75t_L g142 ( .A(n_101), .B(n_2), .Y(n_142) );
INVx2_ASAP7_75t_L g143 ( .A(n_92), .Y(n_143) );
HB1xp67_ASAP7_75t_L g144 ( .A(n_127), .Y(n_144) );
INVx3_ASAP7_75t_L g145 ( .A(n_95), .Y(n_145) );
INVx3_ASAP7_75t_L g146 ( .A(n_95), .Y(n_146) );
INVx5_ASAP7_75t_L g147 ( .A(n_92), .Y(n_147) );
INVx3_ASAP7_75t_L g148 ( .A(n_95), .Y(n_148) );
INVx1_ASAP7_75t_L g149 ( .A(n_128), .Y(n_149) );
INVx1_ASAP7_75t_L g150 ( .A(n_128), .Y(n_150) );
INVxp67_ASAP7_75t_L g151 ( .A(n_127), .Y(n_151) );
HB1xp67_ASAP7_75t_L g152 ( .A(n_120), .Y(n_152) );
INVx1_ASAP7_75t_L g153 ( .A(n_133), .Y(n_153) );
OR2x2_ASAP7_75t_L g154 ( .A(n_144), .B(n_119), .Y(n_154) );
INVx4_ASAP7_75t_L g155 ( .A(n_133), .Y(n_155) );
NAND2xp5_ASAP7_75t_L g156 ( .A(n_151), .B(n_106), .Y(n_156) );
AOI22xp33_ASAP7_75t_L g157 ( .A1(n_133), .A2(n_93), .B1(n_114), .B2(n_113), .Y(n_157) );
INVx2_ASAP7_75t_L g158 ( .A(n_132), .Y(n_158) );
INVx4_ASAP7_75t_L g159 ( .A(n_133), .Y(n_159) );
INVx2_ASAP7_75t_L g160 ( .A(n_132), .Y(n_160) );
INVx1_ASAP7_75t_L g161 ( .A(n_133), .Y(n_161) );
BUFx6f_ASAP7_75t_L g162 ( .A(n_147), .Y(n_162) );
INVx1_ASAP7_75t_L g163 ( .A(n_133), .Y(n_163) );
INVx2_ASAP7_75t_L g164 ( .A(n_147), .Y(n_164) );
AND2x2_ASAP7_75t_L g165 ( .A(n_151), .B(n_129), .Y(n_165) );
NAND2xp5_ASAP7_75t_L g166 ( .A(n_152), .B(n_108), .Y(n_166) );
INVx2_ASAP7_75t_L g167 ( .A(n_147), .Y(n_167) );
NAND2xp5_ASAP7_75t_L g168 ( .A(n_152), .B(n_104), .Y(n_168) );
INVx1_ASAP7_75t_L g169 ( .A(n_142), .Y(n_169) );
INVx1_ASAP7_75t_L g170 ( .A(n_142), .Y(n_170) );
NAND2xp5_ASAP7_75t_SL g171 ( .A(n_138), .B(n_107), .Y(n_171) );
NAND2xp5_ASAP7_75t_L g172 ( .A(n_144), .B(n_104), .Y(n_172) );
NOR2xp33_ASAP7_75t_L g173 ( .A(n_134), .B(n_131), .Y(n_173) );
INVx1_ASAP7_75t_L g174 ( .A(n_142), .Y(n_174) );
BUFx6f_ASAP7_75t_L g175 ( .A(n_147), .Y(n_175) );
INVx2_ASAP7_75t_L g176 ( .A(n_132), .Y(n_176) );
NAND3xp33_ASAP7_75t_L g177 ( .A(n_142), .B(n_112), .C(n_115), .Y(n_177) );
INVx1_ASAP7_75t_L g178 ( .A(n_142), .Y(n_178) );
INVx2_ASAP7_75t_SL g179 ( .A(n_138), .Y(n_179) );
AOI22xp33_ASAP7_75t_L g180 ( .A1(n_142), .A2(n_93), .B1(n_95), .B2(n_115), .Y(n_180) );
AO22x1_ASAP7_75t_L g181 ( .A1(n_140), .A2(n_141), .B1(n_139), .B2(n_138), .Y(n_181) );
OR2x6_ASAP7_75t_L g182 ( .A(n_140), .B(n_98), .Y(n_182) );
BUFx3_ASAP7_75t_L g183 ( .A(n_147), .Y(n_183) );
INVx1_ASAP7_75t_L g184 ( .A(n_136), .Y(n_184) );
NAND2xp5_ASAP7_75t_L g185 ( .A(n_179), .B(n_134), .Y(n_185) );
OAI22xp5_ASAP7_75t_SL g186 ( .A1(n_154), .A2(n_130), .B1(n_112), .B2(n_136), .Y(n_186) );
INVx1_ASAP7_75t_L g187 ( .A(n_153), .Y(n_187) );
INVx2_ASAP7_75t_SL g188 ( .A(n_155), .Y(n_188) );
AOI21xp5_ASAP7_75t_L g189 ( .A1(n_179), .A2(n_139), .B(n_141), .Y(n_189) );
NOR2xp33_ASAP7_75t_L g190 ( .A(n_166), .B(n_135), .Y(n_190) );
AOI22xp33_ASAP7_75t_L g191 ( .A1(n_155), .A2(n_136), .B1(n_139), .B2(n_141), .Y(n_191) );
OAI22xp5_ASAP7_75t_L g192 ( .A1(n_180), .A2(n_130), .B1(n_149), .B2(n_135), .Y(n_192) );
NAND2xp5_ASAP7_75t_L g193 ( .A(n_156), .B(n_149), .Y(n_193) );
NOR2xp33_ASAP7_75t_L g194 ( .A(n_168), .B(n_150), .Y(n_194) );
HB1xp67_ASAP7_75t_L g195 ( .A(n_154), .Y(n_195) );
OAI221xp5_ASAP7_75t_L g196 ( .A1(n_157), .A2(n_150), .B1(n_136), .B2(n_96), .C(n_100), .Y(n_196) );
NAND2xp5_ASAP7_75t_L g197 ( .A(n_173), .B(n_107), .Y(n_197) );
OR2x6_ASAP7_75t_L g198 ( .A(n_182), .B(n_136), .Y(n_198) );
NAND2xp5_ASAP7_75t_L g199 ( .A(n_155), .B(n_122), .Y(n_199) );
INVx8_ASAP7_75t_L g200 ( .A(n_182), .Y(n_200) );
NAND3xp33_ASAP7_75t_SL g201 ( .A(n_172), .B(n_122), .C(n_109), .Y(n_201) );
NAND2xp5_ASAP7_75t_L g202 ( .A(n_155), .B(n_121), .Y(n_202) );
INVx2_ASAP7_75t_L g203 ( .A(n_184), .Y(n_203) );
AOI22xp33_ASAP7_75t_L g204 ( .A1(n_159), .A2(n_136), .B1(n_99), .B2(n_110), .Y(n_204) );
INVx1_ASAP7_75t_L g205 ( .A(n_153), .Y(n_205) );
NAND2xp5_ASAP7_75t_SL g206 ( .A(n_159), .B(n_116), .Y(n_206) );
INVx1_ASAP7_75t_L g207 ( .A(n_161), .Y(n_207) );
OAI22xp5_ASAP7_75t_L g208 ( .A1(n_177), .A2(n_125), .B1(n_117), .B2(n_118), .Y(n_208) );
BUFx3_ASAP7_75t_L g209 ( .A(n_161), .Y(n_209) );
NAND2xp5_ASAP7_75t_L g210 ( .A(n_159), .B(n_123), .Y(n_210) );
NAND2xp5_ASAP7_75t_L g211 ( .A(n_159), .B(n_124), .Y(n_211) );
NOR2xp67_ASAP7_75t_L g212 ( .A(n_165), .B(n_3), .Y(n_212) );
NAND2xp5_ASAP7_75t_SL g213 ( .A(n_184), .B(n_126), .Y(n_213) );
NAND2xp5_ASAP7_75t_SL g214 ( .A(n_163), .B(n_111), .Y(n_214) );
NAND2xp5_ASAP7_75t_L g215 ( .A(n_171), .B(n_111), .Y(n_215) );
AOI22xp33_ASAP7_75t_L g216 ( .A1(n_182), .A2(n_148), .B1(n_132), .B2(n_146), .Y(n_216) );
INVxp67_ASAP7_75t_L g217 ( .A(n_165), .Y(n_217) );
NAND2xp5_ASAP7_75t_L g218 ( .A(n_163), .B(n_147), .Y(n_218) );
NAND2xp5_ASAP7_75t_L g219 ( .A(n_169), .B(n_147), .Y(n_219) );
NAND2xp5_ASAP7_75t_L g220 ( .A(n_169), .B(n_147), .Y(n_220) );
INVx4_ASAP7_75t_L g221 ( .A(n_183), .Y(n_221) );
INVx2_ASAP7_75t_SL g222 ( .A(n_170), .Y(n_222) );
NAND2xp33_ASAP7_75t_L g223 ( .A(n_170), .B(n_92), .Y(n_223) );
NAND2xp5_ASAP7_75t_L g224 ( .A(n_174), .B(n_147), .Y(n_224) );
NAND2xp5_ASAP7_75t_L g225 ( .A(n_174), .B(n_178), .Y(n_225) );
AOI22xp5_ASAP7_75t_L g226 ( .A1(n_182), .A2(n_148), .B1(n_146), .B2(n_145), .Y(n_226) );
NAND2xp5_ASAP7_75t_L g227 ( .A(n_190), .B(n_182), .Y(n_227) );
NAND2xp5_ASAP7_75t_L g228 ( .A(n_194), .B(n_181), .Y(n_228) );
NOR2xp67_ASAP7_75t_L g229 ( .A(n_195), .B(n_178), .Y(n_229) );
NAND2xp5_ASAP7_75t_L g230 ( .A(n_193), .B(n_217), .Y(n_230) );
A2O1A1Ixp33_ASAP7_75t_L g231 ( .A1(n_222), .A2(n_181), .B(n_137), .C(n_143), .Y(n_231) );
AOI21xp5_ASAP7_75t_L g232 ( .A1(n_213), .A2(n_167), .B(n_164), .Y(n_232) );
AOI21xp5_ASAP7_75t_L g233 ( .A1(n_213), .A2(n_167), .B(n_164), .Y(n_233) );
AOI21xp5_ASAP7_75t_L g234 ( .A1(n_203), .A2(n_167), .B(n_164), .Y(n_234) );
NAND2xp5_ASAP7_75t_SL g235 ( .A(n_192), .B(n_92), .Y(n_235) );
AOI22xp5_ASAP7_75t_L g236 ( .A1(n_186), .A2(n_97), .B1(n_148), .B2(n_146), .Y(n_236) );
AOI33xp33_ASAP7_75t_L g237 ( .A1(n_216), .A2(n_137), .A3(n_143), .B1(n_158), .B2(n_160), .B3(n_176), .Y(n_237) );
OAI22xp5_ASAP7_75t_L g238 ( .A1(n_200), .A2(n_148), .B1(n_132), .B2(n_145), .Y(n_238) );
INVx3_ASAP7_75t_L g239 ( .A(n_209), .Y(n_239) );
INVx1_ASAP7_75t_SL g240 ( .A(n_199), .Y(n_240) );
NAND2xp5_ASAP7_75t_L g241 ( .A(n_212), .B(n_145), .Y(n_241) );
OAI21x1_ASAP7_75t_L g242 ( .A1(n_203), .A2(n_148), .B(n_145), .Y(n_242) );
AOI21xp5_ASAP7_75t_L g243 ( .A1(n_189), .A2(n_158), .B(n_176), .Y(n_243) );
INVx3_ASAP7_75t_SL g244 ( .A(n_200), .Y(n_244) );
NOR2xp33_ASAP7_75t_L g245 ( .A(n_197), .B(n_3), .Y(n_245) );
NAND2xp5_ASAP7_75t_SL g246 ( .A(n_222), .B(n_97), .Y(n_246) );
INVx3_ASAP7_75t_L g247 ( .A(n_209), .Y(n_247) );
NAND2xp5_ASAP7_75t_SL g248 ( .A(n_200), .B(n_97), .Y(n_248) );
NAND2xp5_ASAP7_75t_L g249 ( .A(n_200), .B(n_187), .Y(n_249) );
NAND2xp5_ASAP7_75t_SL g250 ( .A(n_188), .B(n_97), .Y(n_250) );
AOI21xp5_ASAP7_75t_L g251 ( .A1(n_185), .A2(n_160), .B(n_183), .Y(n_251) );
NOR2xp33_ASAP7_75t_L g252 ( .A(n_201), .B(n_4), .Y(n_252) );
INVx3_ASAP7_75t_L g253 ( .A(n_221), .Y(n_253) );
BUFx4f_ASAP7_75t_L g254 ( .A(n_198), .Y(n_254) );
A2O1A1Ixp33_ASAP7_75t_L g255 ( .A1(n_205), .A2(n_137), .B(n_143), .C(n_145), .Y(n_255) );
INVxp67_ASAP7_75t_L g256 ( .A(n_188), .Y(n_256) );
AND2x4_ASAP7_75t_L g257 ( .A(n_207), .B(n_6), .Y(n_257) );
AOI21xp5_ASAP7_75t_L g258 ( .A1(n_206), .A2(n_183), .B(n_175), .Y(n_258) );
AOI21xp5_ASAP7_75t_L g259 ( .A1(n_206), .A2(n_175), .B(n_162), .Y(n_259) );
INVx3_ASAP7_75t_L g260 ( .A(n_221), .Y(n_260) );
NAND2xp5_ASAP7_75t_L g261 ( .A(n_230), .B(n_225), .Y(n_261) );
OAI22xp5_ASAP7_75t_L g262 ( .A1(n_254), .A2(n_198), .B1(n_196), .B2(n_204), .Y(n_262) );
NAND2xp5_ASAP7_75t_L g263 ( .A(n_227), .B(n_208), .Y(n_263) );
A2O1A1Ixp33_ASAP7_75t_L g264 ( .A1(n_245), .A2(n_226), .B(n_210), .C(n_211), .Y(n_264) );
NAND2xp5_ASAP7_75t_L g265 ( .A(n_229), .B(n_202), .Y(n_265) );
AOI22xp5_ASAP7_75t_L g266 ( .A1(n_257), .A2(n_236), .B1(n_228), .B2(n_254), .Y(n_266) );
INVx1_ASAP7_75t_L g267 ( .A(n_237), .Y(n_267) );
OAI21x1_ASAP7_75t_L g268 ( .A1(n_242), .A2(n_191), .B(n_214), .Y(n_268) );
AND2x2_ASAP7_75t_L g269 ( .A(n_244), .B(n_198), .Y(n_269) );
AOI21xp5_ASAP7_75t_L g270 ( .A1(n_243), .A2(n_224), .B(n_218), .Y(n_270) );
INVx1_ASAP7_75t_L g271 ( .A(n_239), .Y(n_271) );
BUFx3_ASAP7_75t_L g272 ( .A(n_244), .Y(n_272) );
OAI21x1_ASAP7_75t_L g273 ( .A1(n_232), .A2(n_214), .B(n_219), .Y(n_273) );
OAI21x1_ASAP7_75t_SL g274 ( .A1(n_249), .A2(n_215), .B(n_220), .Y(n_274) );
HB1xp67_ASAP7_75t_L g275 ( .A(n_257), .Y(n_275) );
NAND2xp5_ASAP7_75t_SL g276 ( .A(n_240), .B(n_221), .Y(n_276) );
NAND2xp5_ASAP7_75t_L g277 ( .A(n_245), .B(n_198), .Y(n_277) );
OAI21x1_ASAP7_75t_L g278 ( .A1(n_233), .A2(n_143), .B(n_137), .Y(n_278) );
NAND2xp5_ASAP7_75t_SL g279 ( .A(n_239), .B(n_97), .Y(n_279) );
AO21x1_ASAP7_75t_L g280 ( .A1(n_235), .A2(n_223), .B(n_146), .Y(n_280) );
AOI21xp5_ASAP7_75t_L g281 ( .A1(n_251), .A2(n_223), .B(n_175), .Y(n_281) );
NOR2xp33_ASAP7_75t_L g282 ( .A(n_247), .B(n_7), .Y(n_282) );
INVx1_ASAP7_75t_SL g283 ( .A(n_247), .Y(n_283) );
OAI21x1_ASAP7_75t_L g284 ( .A1(n_259), .A2(n_146), .B(n_51), .Y(n_284) );
INVx1_ASAP7_75t_L g285 ( .A(n_267), .Y(n_285) );
INVx1_ASAP7_75t_L g286 ( .A(n_267), .Y(n_286) );
OAI21xp5_ASAP7_75t_L g287 ( .A1(n_264), .A2(n_231), .B(n_234), .Y(n_287) );
BUFx6f_ASAP7_75t_L g288 ( .A(n_284), .Y(n_288) );
OA21x2_ASAP7_75t_L g289 ( .A1(n_284), .A2(n_255), .B(n_241), .Y(n_289) );
INVx3_ASAP7_75t_L g290 ( .A(n_272), .Y(n_290) );
INVx1_ASAP7_75t_L g291 ( .A(n_261), .Y(n_291) );
AOI221xp5_ASAP7_75t_L g292 ( .A1(n_263), .A2(n_252), .B1(n_238), .B2(n_248), .C(n_256), .Y(n_292) );
OAI21x1_ASAP7_75t_L g293 ( .A1(n_278), .A2(n_246), .B(n_250), .Y(n_293) );
OAI21xp5_ASAP7_75t_L g294 ( .A1(n_268), .A2(n_252), .B(n_258), .Y(n_294) );
NAND2xp5_ASAP7_75t_L g295 ( .A(n_266), .B(n_253), .Y(n_295) );
AOI21xp5_ASAP7_75t_L g296 ( .A1(n_270), .A2(n_256), .B(n_260), .Y(n_296) );
INVx1_ASAP7_75t_L g297 ( .A(n_274), .Y(n_297) );
BUFx6f_ASAP7_75t_L g298 ( .A(n_278), .Y(n_298) );
INVx2_ASAP7_75t_SL g299 ( .A(n_272), .Y(n_299) );
INVx2_ASAP7_75t_L g300 ( .A(n_273), .Y(n_300) );
XNOR2xp5_ASAP7_75t_L g301 ( .A(n_275), .B(n_253), .Y(n_301) );
INVx2_ASAP7_75t_L g302 ( .A(n_273), .Y(n_302) );
BUFx12f_ASAP7_75t_L g303 ( .A(n_269), .Y(n_303) );
OAI21x1_ASAP7_75t_SL g304 ( .A1(n_274), .A2(n_260), .B(n_9), .Y(n_304) );
INVx1_ASAP7_75t_L g305 ( .A(n_271), .Y(n_305) );
OA21x2_ASAP7_75t_L g306 ( .A1(n_268), .A2(n_50), .B(n_91), .Y(n_306) );
OAI21x1_ASAP7_75t_L g307 ( .A1(n_281), .A2(n_49), .B(n_90), .Y(n_307) );
INVx1_ASAP7_75t_L g308 ( .A(n_305), .Y(n_308) );
INVx1_ASAP7_75t_L g309 ( .A(n_305), .Y(n_309) );
INVx1_ASAP7_75t_L g310 ( .A(n_297), .Y(n_310) );
BUFx3_ASAP7_75t_L g311 ( .A(n_303), .Y(n_311) );
INVx1_ASAP7_75t_L g312 ( .A(n_297), .Y(n_312) );
INVx2_ASAP7_75t_L g313 ( .A(n_300), .Y(n_313) );
OA21x2_ASAP7_75t_L g314 ( .A1(n_294), .A2(n_277), .B(n_280), .Y(n_314) );
AND2x4_ASAP7_75t_L g315 ( .A(n_295), .B(n_271), .Y(n_315) );
INVx1_ASAP7_75t_SL g316 ( .A(n_290), .Y(n_316) );
INVx2_ASAP7_75t_L g317 ( .A(n_300), .Y(n_317) );
INVx1_ASAP7_75t_L g318 ( .A(n_304), .Y(n_318) );
AOI22xp33_ASAP7_75t_L g319 ( .A1(n_291), .A2(n_262), .B1(n_266), .B2(n_265), .Y(n_319) );
AOI21x1_ASAP7_75t_L g320 ( .A1(n_304), .A2(n_262), .B(n_279), .Y(n_320) );
INVx1_ASAP7_75t_L g321 ( .A(n_285), .Y(n_321) );
NOR2xp33_ASAP7_75t_L g322 ( .A(n_291), .B(n_269), .Y(n_322) );
INVx2_ASAP7_75t_L g323 ( .A(n_300), .Y(n_323) );
OAI21xp5_ASAP7_75t_L g324 ( .A1(n_287), .A2(n_282), .B(n_276), .Y(n_324) );
OAI21xp5_ASAP7_75t_L g325 ( .A1(n_287), .A2(n_283), .B(n_280), .Y(n_325) );
AND2x2_ASAP7_75t_L g326 ( .A(n_285), .B(n_283), .Y(n_326) );
OR2x2_ASAP7_75t_L g327 ( .A(n_295), .B(n_8), .Y(n_327) );
INVx2_ASAP7_75t_L g328 ( .A(n_302), .Y(n_328) );
INVx3_ASAP7_75t_L g329 ( .A(n_290), .Y(n_329) );
HB1xp67_ASAP7_75t_L g330 ( .A(n_299), .Y(n_330) );
INVx1_ASAP7_75t_L g331 ( .A(n_286), .Y(n_331) );
INVx1_ASAP7_75t_L g332 ( .A(n_286), .Y(n_332) );
INVx1_ASAP7_75t_L g333 ( .A(n_302), .Y(n_333) );
AND2x2_ASAP7_75t_L g334 ( .A(n_290), .B(n_8), .Y(n_334) );
INVx1_ASAP7_75t_L g335 ( .A(n_302), .Y(n_335) );
AND2x4_ASAP7_75t_L g336 ( .A(n_294), .B(n_53), .Y(n_336) );
INVx1_ASAP7_75t_L g337 ( .A(n_306), .Y(n_337) );
OAI21xp5_ASAP7_75t_L g338 ( .A1(n_296), .A2(n_9), .B(n_10), .Y(n_338) );
AND2x4_ASAP7_75t_L g339 ( .A(n_290), .B(n_56), .Y(n_339) );
INVx1_ASAP7_75t_L g340 ( .A(n_306), .Y(n_340) );
INVx1_ASAP7_75t_L g341 ( .A(n_310), .Y(n_341) );
BUFx6f_ASAP7_75t_L g342 ( .A(n_320), .Y(n_342) );
AND2x2_ASAP7_75t_L g343 ( .A(n_308), .B(n_298), .Y(n_343) );
AO21x2_ASAP7_75t_L g344 ( .A1(n_325), .A2(n_296), .B(n_307), .Y(n_344) );
NOR2xp33_ASAP7_75t_L g345 ( .A(n_322), .B(n_299), .Y(n_345) );
INVxp67_ASAP7_75t_L g346 ( .A(n_330), .Y(n_346) );
INVx1_ASAP7_75t_L g347 ( .A(n_310), .Y(n_347) );
INVx2_ASAP7_75t_L g348 ( .A(n_313), .Y(n_348) );
OR2x2_ASAP7_75t_L g349 ( .A(n_312), .B(n_301), .Y(n_349) );
INVx3_ASAP7_75t_L g350 ( .A(n_336), .Y(n_350) );
INVxp67_ASAP7_75t_SL g351 ( .A(n_327), .Y(n_351) );
NAND2x1p5_ASAP7_75t_SL g352 ( .A(n_334), .B(n_289), .Y(n_352) );
INVx2_ASAP7_75t_L g353 ( .A(n_313), .Y(n_353) );
INVx1_ASAP7_75t_L g354 ( .A(n_312), .Y(n_354) );
AND2x2_ASAP7_75t_L g355 ( .A(n_308), .B(n_298), .Y(n_355) );
INVx1_ASAP7_75t_L g356 ( .A(n_309), .Y(n_356) );
INVx1_ASAP7_75t_L g357 ( .A(n_309), .Y(n_357) );
AND2x2_ASAP7_75t_L g358 ( .A(n_315), .B(n_298), .Y(n_358) );
OR2x6_ASAP7_75t_L g359 ( .A(n_318), .B(n_288), .Y(n_359) );
INVx1_ASAP7_75t_L g360 ( .A(n_333), .Y(n_360) );
INVx2_ASAP7_75t_L g361 ( .A(n_313), .Y(n_361) );
HB1xp67_ASAP7_75t_L g362 ( .A(n_334), .Y(n_362) );
NAND2xp5_ASAP7_75t_L g363 ( .A(n_321), .B(n_301), .Y(n_363) );
INVx1_ASAP7_75t_L g364 ( .A(n_333), .Y(n_364) );
AND2x2_ASAP7_75t_L g365 ( .A(n_315), .B(n_298), .Y(n_365) );
INVx2_ASAP7_75t_L g366 ( .A(n_317), .Y(n_366) );
INVx1_ASAP7_75t_L g367 ( .A(n_335), .Y(n_367) );
INVx1_ASAP7_75t_L g368 ( .A(n_335), .Y(n_368) );
HB1xp67_ASAP7_75t_L g369 ( .A(n_311), .Y(n_369) );
HB1xp67_ASAP7_75t_L g370 ( .A(n_311), .Y(n_370) );
OAI31xp33_ASAP7_75t_L g371 ( .A1(n_311), .A2(n_303), .A3(n_292), .B(n_12), .Y(n_371) );
INVx3_ASAP7_75t_L g372 ( .A(n_336), .Y(n_372) );
OR2x2_ASAP7_75t_L g373 ( .A(n_327), .B(n_298), .Y(n_373) );
NOR2xp33_ASAP7_75t_L g374 ( .A(n_321), .B(n_303), .Y(n_374) );
INVx3_ASAP7_75t_L g375 ( .A(n_336), .Y(n_375) );
INVx3_ASAP7_75t_L g376 ( .A(n_336), .Y(n_376) );
INVx2_ASAP7_75t_SL g377 ( .A(n_329), .Y(n_377) );
HB1xp67_ASAP7_75t_L g378 ( .A(n_316), .Y(n_378) );
INVx1_ASAP7_75t_L g379 ( .A(n_331), .Y(n_379) );
NOR2xp33_ASAP7_75t_L g380 ( .A(n_331), .B(n_10), .Y(n_380) );
NAND2xp5_ASAP7_75t_L g381 ( .A(n_332), .B(n_292), .Y(n_381) );
HB1xp67_ASAP7_75t_L g382 ( .A(n_316), .Y(n_382) );
INVx2_ASAP7_75t_L g383 ( .A(n_317), .Y(n_383) );
HB1xp67_ASAP7_75t_L g384 ( .A(n_329), .Y(n_384) );
BUFx2_ASAP7_75t_L g385 ( .A(n_317), .Y(n_385) );
INVx3_ASAP7_75t_L g386 ( .A(n_323), .Y(n_386) );
AND2x2_ASAP7_75t_L g387 ( .A(n_315), .B(n_298), .Y(n_387) );
INVx2_ASAP7_75t_L g388 ( .A(n_323), .Y(n_388) );
INVx5_ASAP7_75t_SL g389 ( .A(n_339), .Y(n_389) );
BUFx6f_ASAP7_75t_L g390 ( .A(n_320), .Y(n_390) );
AOI22xp5_ASAP7_75t_L g391 ( .A1(n_319), .A2(n_289), .B1(n_306), .B2(n_288), .Y(n_391) );
INVx2_ASAP7_75t_L g392 ( .A(n_323), .Y(n_392) );
AND2x2_ASAP7_75t_L g393 ( .A(n_315), .B(n_288), .Y(n_393) );
INVx4_ASAP7_75t_L g394 ( .A(n_339), .Y(n_394) );
NOR2x1_ASAP7_75t_L g395 ( .A(n_318), .B(n_306), .Y(n_395) );
INVx2_ASAP7_75t_L g396 ( .A(n_328), .Y(n_396) );
NAND2xp5_ASAP7_75t_L g397 ( .A(n_332), .B(n_289), .Y(n_397) );
NAND2xp5_ASAP7_75t_L g398 ( .A(n_351), .B(n_326), .Y(n_398) );
AND2x2_ASAP7_75t_L g399 ( .A(n_343), .B(n_314), .Y(n_399) );
AND2x2_ASAP7_75t_L g400 ( .A(n_343), .B(n_314), .Y(n_400) );
OR2x2_ASAP7_75t_L g401 ( .A(n_373), .B(n_328), .Y(n_401) );
AND2x2_ASAP7_75t_L g402 ( .A(n_355), .B(n_314), .Y(n_402) );
INVx1_ASAP7_75t_L g403 ( .A(n_356), .Y(n_403) );
INVx2_ASAP7_75t_L g404 ( .A(n_385), .Y(n_404) );
BUFx2_ASAP7_75t_L g405 ( .A(n_394), .Y(n_405) );
OR2x2_ASAP7_75t_L g406 ( .A(n_373), .B(n_328), .Y(n_406) );
INVx1_ASAP7_75t_L g407 ( .A(n_341), .Y(n_407) );
INVxp67_ASAP7_75t_L g408 ( .A(n_369), .Y(n_408) );
HB1xp67_ASAP7_75t_L g409 ( .A(n_370), .Y(n_409) );
NAND2xp5_ASAP7_75t_L g410 ( .A(n_363), .B(n_326), .Y(n_410) );
NAND2xp5_ASAP7_75t_L g411 ( .A(n_357), .B(n_338), .Y(n_411) );
INVxp67_ASAP7_75t_L g412 ( .A(n_345), .Y(n_412) );
AND2x2_ASAP7_75t_L g413 ( .A(n_355), .B(n_314), .Y(n_413) );
INVx4_ASAP7_75t_L g414 ( .A(n_394), .Y(n_414) );
INVx2_ASAP7_75t_L g415 ( .A(n_385), .Y(n_415) );
AND2x2_ASAP7_75t_L g416 ( .A(n_358), .B(n_314), .Y(n_416) );
INVx1_ASAP7_75t_L g417 ( .A(n_341), .Y(n_417) );
INVx1_ASAP7_75t_L g418 ( .A(n_347), .Y(n_418) );
HB1xp67_ASAP7_75t_L g419 ( .A(n_346), .Y(n_419) );
INVx2_ASAP7_75t_L g420 ( .A(n_348), .Y(n_420) );
AND2x2_ASAP7_75t_L g421 ( .A(n_358), .B(n_337), .Y(n_421) );
INVx1_ASAP7_75t_L g422 ( .A(n_347), .Y(n_422) );
INVx2_ASAP7_75t_L g423 ( .A(n_348), .Y(n_423) );
HB1xp67_ASAP7_75t_L g424 ( .A(n_362), .Y(n_424) );
AND2x2_ASAP7_75t_L g425 ( .A(n_365), .B(n_337), .Y(n_425) );
INVx1_ASAP7_75t_L g426 ( .A(n_354), .Y(n_426) );
AND2x2_ASAP7_75t_L g427 ( .A(n_365), .B(n_340), .Y(n_427) );
AND2x2_ASAP7_75t_L g428 ( .A(n_387), .B(n_340), .Y(n_428) );
NAND2xp5_ASAP7_75t_L g429 ( .A(n_357), .B(n_329), .Y(n_429) );
NOR2xp33_ASAP7_75t_L g430 ( .A(n_349), .B(n_11), .Y(n_430) );
INVx1_ASAP7_75t_L g431 ( .A(n_354), .Y(n_431) );
NAND2xp5_ASAP7_75t_L g432 ( .A(n_379), .B(n_329), .Y(n_432) );
INVx2_ASAP7_75t_SL g433 ( .A(n_394), .Y(n_433) );
NOR2xp33_ASAP7_75t_L g434 ( .A(n_349), .B(n_11), .Y(n_434) );
INVx1_ASAP7_75t_L g435 ( .A(n_379), .Y(n_435) );
INVx1_ASAP7_75t_L g436 ( .A(n_360), .Y(n_436) );
INVx2_ASAP7_75t_L g437 ( .A(n_348), .Y(n_437) );
INVx1_ASAP7_75t_L g438 ( .A(n_360), .Y(n_438) );
NAND2xp5_ASAP7_75t_L g439 ( .A(n_381), .B(n_324), .Y(n_439) );
HB1xp67_ASAP7_75t_L g440 ( .A(n_378), .Y(n_440) );
OR2x2_ASAP7_75t_L g441 ( .A(n_364), .B(n_325), .Y(n_441) );
INVx1_ASAP7_75t_L g442 ( .A(n_367), .Y(n_442) );
NAND2xp5_ASAP7_75t_L g443 ( .A(n_374), .B(n_324), .Y(n_443) );
AND2x2_ASAP7_75t_L g444 ( .A(n_387), .B(n_288), .Y(n_444) );
NAND2xp5_ASAP7_75t_L g445 ( .A(n_380), .B(n_339), .Y(n_445) );
INVx1_ASAP7_75t_L g446 ( .A(n_367), .Y(n_446) );
INVx2_ASAP7_75t_L g447 ( .A(n_361), .Y(n_447) );
INVx1_ASAP7_75t_L g448 ( .A(n_368), .Y(n_448) );
BUFx3_ASAP7_75t_L g449 ( .A(n_377), .Y(n_449) );
AND2x2_ASAP7_75t_L g450 ( .A(n_393), .B(n_288), .Y(n_450) );
INVx2_ASAP7_75t_L g451 ( .A(n_361), .Y(n_451) );
OR2x2_ASAP7_75t_L g452 ( .A(n_368), .B(n_339), .Y(n_452) );
AND2x2_ASAP7_75t_L g453 ( .A(n_393), .B(n_288), .Y(n_453) );
AND2x2_ASAP7_75t_L g454 ( .A(n_386), .B(n_306), .Y(n_454) );
INVx2_ASAP7_75t_L g455 ( .A(n_361), .Y(n_455) );
AND2x2_ASAP7_75t_L g456 ( .A(n_386), .B(n_350), .Y(n_456) );
INVx1_ASAP7_75t_L g457 ( .A(n_366), .Y(n_457) );
AND2x4_ASAP7_75t_L g458 ( .A(n_350), .B(n_307), .Y(n_458) );
BUFx2_ASAP7_75t_L g459 ( .A(n_382), .Y(n_459) );
AND2x2_ASAP7_75t_L g460 ( .A(n_386), .B(n_289), .Y(n_460) );
NAND2xp5_ASAP7_75t_L g461 ( .A(n_389), .B(n_14), .Y(n_461) );
INVx2_ASAP7_75t_L g462 ( .A(n_366), .Y(n_462) );
OR2x2_ASAP7_75t_L g463 ( .A(n_397), .B(n_289), .Y(n_463) );
AND2x2_ASAP7_75t_L g464 ( .A(n_386), .B(n_307), .Y(n_464) );
OR2x2_ASAP7_75t_L g465 ( .A(n_366), .B(n_14), .Y(n_465) );
INVx1_ASAP7_75t_L g466 ( .A(n_383), .Y(n_466) );
INVx2_ASAP7_75t_L g467 ( .A(n_383), .Y(n_467) );
INVx1_ASAP7_75t_L g468 ( .A(n_383), .Y(n_468) );
HB1xp67_ASAP7_75t_L g469 ( .A(n_384), .Y(n_469) );
INVx2_ASAP7_75t_L g470 ( .A(n_388), .Y(n_470) );
NAND2xp5_ASAP7_75t_L g471 ( .A(n_389), .B(n_16), .Y(n_471) );
AND2x2_ASAP7_75t_L g472 ( .A(n_350), .B(n_16), .Y(n_472) );
INVx1_ASAP7_75t_L g473 ( .A(n_388), .Y(n_473) );
AND2x2_ASAP7_75t_L g474 ( .A(n_350), .B(n_18), .Y(n_474) );
NAND3xp33_ASAP7_75t_L g475 ( .A(n_371), .B(n_19), .C(n_175), .Y(n_475) );
AND2x2_ASAP7_75t_L g476 ( .A(n_416), .B(n_376), .Y(n_476) );
NAND2xp5_ASAP7_75t_L g477 ( .A(n_424), .B(n_396), .Y(n_477) );
INVxp67_ASAP7_75t_L g478 ( .A(n_409), .Y(n_478) );
NAND2xp5_ASAP7_75t_L g479 ( .A(n_410), .B(n_396), .Y(n_479) );
AND2x2_ASAP7_75t_L g480 ( .A(n_416), .B(n_376), .Y(n_480) );
BUFx2_ASAP7_75t_SL g481 ( .A(n_414), .Y(n_481) );
AND2x2_ASAP7_75t_L g482 ( .A(n_399), .B(n_376), .Y(n_482) );
AND2x2_ASAP7_75t_L g483 ( .A(n_399), .B(n_376), .Y(n_483) );
INVxp67_ASAP7_75t_L g484 ( .A(n_440), .Y(n_484) );
OR2x2_ASAP7_75t_L g485 ( .A(n_398), .B(n_396), .Y(n_485) );
INVx1_ASAP7_75t_SL g486 ( .A(n_419), .Y(n_486) );
INVx2_ASAP7_75t_L g487 ( .A(n_420), .Y(n_487) );
INVx1_ASAP7_75t_L g488 ( .A(n_407), .Y(n_488) );
AND2x2_ASAP7_75t_L g489 ( .A(n_400), .B(n_375), .Y(n_489) );
AND2x2_ASAP7_75t_L g490 ( .A(n_400), .B(n_375), .Y(n_490) );
OAI21xp5_ASAP7_75t_L g491 ( .A1(n_430), .A2(n_391), .B(n_395), .Y(n_491) );
INVx1_ASAP7_75t_L g492 ( .A(n_417), .Y(n_492) );
INVx1_ASAP7_75t_L g493 ( .A(n_417), .Y(n_493) );
INVx1_ASAP7_75t_L g494 ( .A(n_418), .Y(n_494) );
OR2x2_ASAP7_75t_L g495 ( .A(n_408), .B(n_388), .Y(n_495) );
INVx1_ASAP7_75t_L g496 ( .A(n_418), .Y(n_496) );
OR2x2_ASAP7_75t_L g497 ( .A(n_459), .B(n_392), .Y(n_497) );
INVx2_ASAP7_75t_L g498 ( .A(n_420), .Y(n_498) );
INVxp67_ASAP7_75t_L g499 ( .A(n_459), .Y(n_499) );
INVx1_ASAP7_75t_L g500 ( .A(n_422), .Y(n_500) );
AND2x2_ASAP7_75t_L g501 ( .A(n_402), .B(n_372), .Y(n_501) );
AND2x2_ASAP7_75t_L g502 ( .A(n_402), .B(n_372), .Y(n_502) );
INVx1_ASAP7_75t_L g503 ( .A(n_422), .Y(n_503) );
NAND2xp5_ASAP7_75t_L g504 ( .A(n_439), .B(n_392), .Y(n_504) );
OR2x2_ASAP7_75t_L g505 ( .A(n_401), .B(n_392), .Y(n_505) );
OR2x2_ASAP7_75t_L g506 ( .A(n_401), .B(n_353), .Y(n_506) );
OR2x2_ASAP7_75t_L g507 ( .A(n_406), .B(n_353), .Y(n_507) );
INVx1_ASAP7_75t_L g508 ( .A(n_426), .Y(n_508) );
INVx2_ASAP7_75t_L g509 ( .A(n_423), .Y(n_509) );
INVx1_ASAP7_75t_L g510 ( .A(n_426), .Y(n_510) );
INVx2_ASAP7_75t_L g511 ( .A(n_423), .Y(n_511) );
NAND2xp5_ASAP7_75t_L g512 ( .A(n_403), .B(n_372), .Y(n_512) );
AND2x2_ASAP7_75t_L g513 ( .A(n_413), .B(n_375), .Y(n_513) );
AND2x2_ASAP7_75t_L g514 ( .A(n_413), .B(n_375), .Y(n_514) );
AND2x2_ASAP7_75t_SL g515 ( .A(n_405), .B(n_342), .Y(n_515) );
INVx2_ASAP7_75t_L g516 ( .A(n_437), .Y(n_516) );
AND2x2_ASAP7_75t_L g517 ( .A(n_421), .B(n_359), .Y(n_517) );
AND2x4_ASAP7_75t_L g518 ( .A(n_405), .B(n_359), .Y(n_518) );
INVx2_ASAP7_75t_L g519 ( .A(n_437), .Y(n_519) );
NAND2xp5_ASAP7_75t_L g520 ( .A(n_435), .B(n_377), .Y(n_520) );
AND2x2_ASAP7_75t_L g521 ( .A(n_421), .B(n_425), .Y(n_521) );
OR2x2_ASAP7_75t_L g522 ( .A(n_469), .B(n_352), .Y(n_522) );
AND2x2_ASAP7_75t_L g523 ( .A(n_425), .B(n_359), .Y(n_523) );
INVx1_ASAP7_75t_L g524 ( .A(n_431), .Y(n_524) );
AND2x2_ASAP7_75t_L g525 ( .A(n_427), .B(n_359), .Y(n_525) );
NAND2xp5_ASAP7_75t_L g526 ( .A(n_431), .B(n_352), .Y(n_526) );
OAI22xp5_ASAP7_75t_L g527 ( .A1(n_445), .A2(n_359), .B1(n_391), .B2(n_395), .Y(n_527) );
NAND2x1_ASAP7_75t_L g528 ( .A(n_414), .B(n_390), .Y(n_528) );
AND2x2_ASAP7_75t_L g529 ( .A(n_427), .B(n_344), .Y(n_529) );
INVx1_ASAP7_75t_L g530 ( .A(n_438), .Y(n_530) );
INVx1_ASAP7_75t_L g531 ( .A(n_438), .Y(n_531) );
NAND2xp5_ASAP7_75t_L g532 ( .A(n_436), .B(n_344), .Y(n_532) );
INVx2_ASAP7_75t_L g533 ( .A(n_447), .Y(n_533) );
BUFx3_ASAP7_75t_L g534 ( .A(n_449), .Y(n_534) );
NAND2xp5_ASAP7_75t_L g535 ( .A(n_442), .B(n_390), .Y(n_535) );
OR2x2_ASAP7_75t_L g536 ( .A(n_428), .B(n_390), .Y(n_536) );
AND2x2_ASAP7_75t_L g537 ( .A(n_444), .B(n_390), .Y(n_537) );
INVx2_ASAP7_75t_L g538 ( .A(n_447), .Y(n_538) );
INVx1_ASAP7_75t_L g539 ( .A(n_446), .Y(n_539) );
INVx2_ASAP7_75t_L g540 ( .A(n_451), .Y(n_540) );
AND2x2_ASAP7_75t_L g541 ( .A(n_444), .B(n_390), .Y(n_541) );
OR2x2_ASAP7_75t_L g542 ( .A(n_452), .B(n_390), .Y(n_542) );
INVx2_ASAP7_75t_L g543 ( .A(n_451), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g544 ( .A(n_448), .B(n_342), .Y(n_544) );
INVx2_ASAP7_75t_L g545 ( .A(n_455), .Y(n_545) );
AND2x2_ASAP7_75t_L g546 ( .A(n_450), .B(n_342), .Y(n_546) );
AND2x2_ASAP7_75t_L g547 ( .A(n_450), .B(n_342), .Y(n_547) );
AND2x2_ASAP7_75t_L g548 ( .A(n_453), .B(n_342), .Y(n_548) );
AND2x2_ASAP7_75t_L g549 ( .A(n_453), .B(n_342), .Y(n_549) );
OR2x2_ASAP7_75t_L g550 ( .A(n_441), .B(n_19), .Y(n_550) );
INVx2_ASAP7_75t_L g551 ( .A(n_455), .Y(n_551) );
INVx1_ASAP7_75t_L g552 ( .A(n_429), .Y(n_552) );
OR2x2_ASAP7_75t_L g553 ( .A(n_452), .B(n_20), .Y(n_553) );
AND2x2_ASAP7_75t_L g554 ( .A(n_456), .B(n_293), .Y(n_554) );
INVx3_ASAP7_75t_L g555 ( .A(n_414), .Y(n_555) );
INVx1_ASAP7_75t_L g556 ( .A(n_432), .Y(n_556) );
INVx2_ASAP7_75t_L g557 ( .A(n_462), .Y(n_557) );
OR2x2_ASAP7_75t_L g558 ( .A(n_404), .B(n_415), .Y(n_558) );
OR2x2_ASAP7_75t_L g559 ( .A(n_404), .B(n_21), .Y(n_559) );
INVx1_ASAP7_75t_L g560 ( .A(n_465), .Y(n_560) );
INVx1_ASAP7_75t_L g561 ( .A(n_465), .Y(n_561) );
AND2x2_ASAP7_75t_L g562 ( .A(n_456), .B(n_293), .Y(n_562) );
INVx1_ASAP7_75t_L g563 ( .A(n_472), .Y(n_563) );
OR2x2_ASAP7_75t_L g564 ( .A(n_521), .B(n_441), .Y(n_564) );
AND2x2_ASAP7_75t_L g565 ( .A(n_521), .B(n_412), .Y(n_565) );
AND2x2_ASAP7_75t_L g566 ( .A(n_517), .B(n_433), .Y(n_566) );
INVx2_ASAP7_75t_L g567 ( .A(n_497), .Y(n_567) );
AND2x2_ASAP7_75t_L g568 ( .A(n_517), .B(n_433), .Y(n_568) );
INVx1_ASAP7_75t_L g569 ( .A(n_539), .Y(n_569) );
OR2x2_ASAP7_75t_L g570 ( .A(n_485), .B(n_415), .Y(n_570) );
AOI21x1_ASAP7_75t_L g571 ( .A1(n_528), .A2(n_472), .B(n_474), .Y(n_571) );
INVx1_ASAP7_75t_L g572 ( .A(n_488), .Y(n_572) );
OR2x2_ASAP7_75t_L g573 ( .A(n_477), .B(n_457), .Y(n_573) );
INVx1_ASAP7_75t_L g574 ( .A(n_492), .Y(n_574) );
AND2x2_ASAP7_75t_L g575 ( .A(n_523), .B(n_449), .Y(n_575) );
OAI21xp5_ASAP7_75t_L g576 ( .A1(n_550), .A2(n_434), .B(n_475), .Y(n_576) );
AND2x2_ASAP7_75t_L g577 ( .A(n_523), .B(n_460), .Y(n_577) );
INVx1_ASAP7_75t_L g578 ( .A(n_493), .Y(n_578) );
INVx1_ASAP7_75t_L g579 ( .A(n_494), .Y(n_579) );
INVx1_ASAP7_75t_SL g580 ( .A(n_481), .Y(n_580) );
AND2x4_ASAP7_75t_L g581 ( .A(n_534), .B(n_458), .Y(n_581) );
OR2x2_ASAP7_75t_L g582 ( .A(n_506), .B(n_457), .Y(n_582) );
NAND2xp5_ASAP7_75t_L g583 ( .A(n_552), .B(n_411), .Y(n_583) );
NAND3xp33_ASAP7_75t_L g584 ( .A(n_491), .B(n_443), .C(n_461), .Y(n_584) );
INVx1_ASAP7_75t_L g585 ( .A(n_496), .Y(n_585) );
BUFx2_ASAP7_75t_L g586 ( .A(n_534), .Y(n_586) );
AOI32xp33_ASAP7_75t_L g587 ( .A1(n_486), .A2(n_474), .A3(n_471), .B1(n_458), .B2(n_464), .Y(n_587) );
INVx1_ASAP7_75t_L g588 ( .A(n_500), .Y(n_588) );
OA21x2_ASAP7_75t_L g589 ( .A1(n_532), .A2(n_473), .B(n_468), .Y(n_589) );
NAND2xp5_ASAP7_75t_L g590 ( .A(n_556), .B(n_473), .Y(n_590) );
INVx1_ASAP7_75t_L g591 ( .A(n_503), .Y(n_591) );
INVx1_ASAP7_75t_L g592 ( .A(n_508), .Y(n_592) );
AND2x2_ASAP7_75t_L g593 ( .A(n_525), .B(n_460), .Y(n_593) );
NAND2xp5_ASAP7_75t_L g594 ( .A(n_529), .B(n_468), .Y(n_594) );
OR2x2_ASAP7_75t_L g595 ( .A(n_507), .B(n_466), .Y(n_595) );
AOI22xp5_ASAP7_75t_L g596 ( .A1(n_563), .A2(n_458), .B1(n_466), .B2(n_464), .Y(n_596) );
OA21x2_ASAP7_75t_SL g597 ( .A1(n_518), .A2(n_454), .B(n_463), .Y(n_597) );
OR2x2_ASAP7_75t_L g598 ( .A(n_505), .B(n_470), .Y(n_598) );
AND2x2_ASAP7_75t_L g599 ( .A(n_525), .B(n_470), .Y(n_599) );
INVxp67_ASAP7_75t_L g600 ( .A(n_522), .Y(n_600) );
HB1xp67_ASAP7_75t_L g601 ( .A(n_499), .Y(n_601) );
AND2x2_ASAP7_75t_L g602 ( .A(n_478), .B(n_462), .Y(n_602) );
INVx1_ASAP7_75t_L g603 ( .A(n_510), .Y(n_603) );
AND2x2_ASAP7_75t_L g604 ( .A(n_482), .B(n_483), .Y(n_604) );
AND2x2_ASAP7_75t_L g605 ( .A(n_482), .B(n_467), .Y(n_605) );
INVx1_ASAP7_75t_L g606 ( .A(n_524), .Y(n_606) );
INVx1_ASAP7_75t_L g607 ( .A(n_530), .Y(n_607) );
AND2x2_ASAP7_75t_L g608 ( .A(n_483), .B(n_489), .Y(n_608) );
NAND2xp5_ASAP7_75t_L g609 ( .A(n_529), .B(n_467), .Y(n_609) );
NAND2xp5_ASAP7_75t_L g610 ( .A(n_504), .B(n_463), .Y(n_610) );
AND2x2_ASAP7_75t_L g611 ( .A(n_489), .B(n_454), .Y(n_611) );
INVx1_ASAP7_75t_L g612 ( .A(n_531), .Y(n_612) );
INVx1_ASAP7_75t_L g613 ( .A(n_495), .Y(n_613) );
INVx1_ASAP7_75t_SL g614 ( .A(n_515), .Y(n_614) );
AND2x2_ASAP7_75t_L g615 ( .A(n_490), .B(n_22), .Y(n_615) );
NAND2xp5_ASAP7_75t_L g616 ( .A(n_479), .B(n_293), .Y(n_616) );
INVx1_ASAP7_75t_L g617 ( .A(n_558), .Y(n_617) );
OAI211xp5_ASAP7_75t_SL g618 ( .A1(n_484), .A2(n_23), .B(n_24), .C(n_25), .Y(n_618) );
INVxp67_ASAP7_75t_L g619 ( .A(n_526), .Y(n_619) );
NAND2x1p5_ASAP7_75t_L g620 ( .A(n_555), .B(n_27), .Y(n_620) );
NAND2xp5_ASAP7_75t_SL g621 ( .A(n_515), .B(n_30), .Y(n_621) );
NAND2x1p5_ASAP7_75t_L g622 ( .A(n_553), .B(n_32), .Y(n_622) );
HB1xp67_ASAP7_75t_L g623 ( .A(n_487), .Y(n_623) );
INVx2_ASAP7_75t_L g624 ( .A(n_487), .Y(n_624) );
INVx1_ASAP7_75t_L g625 ( .A(n_520), .Y(n_625) );
BUFx3_ASAP7_75t_L g626 ( .A(n_518), .Y(n_626) );
AND2x2_ASAP7_75t_L g627 ( .A(n_501), .B(n_34), .Y(n_627) );
INVx1_ASAP7_75t_L g628 ( .A(n_512), .Y(n_628) );
NAND2xp5_ASAP7_75t_L g629 ( .A(n_560), .B(n_38), .Y(n_629) );
INVxp33_ASAP7_75t_L g630 ( .A(n_586), .Y(n_630) );
AND2x2_ASAP7_75t_L g631 ( .A(n_604), .B(n_501), .Y(n_631) );
AOI22xp33_ASAP7_75t_L g632 ( .A1(n_584), .A2(n_527), .B1(n_518), .B2(n_514), .Y(n_632) );
INVx1_ASAP7_75t_L g633 ( .A(n_590), .Y(n_633) );
OAI22xp5_ASAP7_75t_L g634 ( .A1(n_580), .A2(n_550), .B1(n_536), .B2(n_514), .Y(n_634) );
HB1xp67_ASAP7_75t_L g635 ( .A(n_623), .Y(n_635) );
AND2x2_ASAP7_75t_L g636 ( .A(n_608), .B(n_502), .Y(n_636) );
AND2x4_ASAP7_75t_SL g637 ( .A(n_566), .B(n_476), .Y(n_637) );
AND2x2_ASAP7_75t_L g638 ( .A(n_577), .B(n_502), .Y(n_638) );
NAND3xp33_ASAP7_75t_SL g639 ( .A(n_580), .B(n_559), .C(n_561), .Y(n_639) );
OAI21xp33_ASAP7_75t_SL g640 ( .A1(n_597), .A2(n_476), .B(n_480), .Y(n_640) );
INVxp33_ASAP7_75t_L g641 ( .A(n_620), .Y(n_641) );
AND2x2_ASAP7_75t_L g642 ( .A(n_593), .B(n_513), .Y(n_642) );
AOI21xp5_ASAP7_75t_L g643 ( .A1(n_621), .A2(n_535), .B(n_544), .Y(n_643) );
INVx1_ASAP7_75t_L g644 ( .A(n_564), .Y(n_644) );
A2O1A1Ixp33_ASAP7_75t_L g645 ( .A1(n_587), .A2(n_480), .B(n_513), .C(n_541), .Y(n_645) );
OAI22xp5_ASAP7_75t_L g646 ( .A1(n_614), .A2(n_542), .B1(n_537), .B2(n_541), .Y(n_646) );
AOI21xp5_ASAP7_75t_L g647 ( .A1(n_620), .A2(n_543), .B(n_557), .Y(n_647) );
AOI32xp33_ASAP7_75t_L g648 ( .A1(n_614), .A2(n_537), .A3(n_546), .B1(n_549), .B2(n_548), .Y(n_648) );
INVx1_ASAP7_75t_L g649 ( .A(n_601), .Y(n_649) );
AOI32xp33_ASAP7_75t_L g650 ( .A1(n_565), .A2(n_546), .A3(n_547), .B1(n_549), .B2(n_548), .Y(n_650) );
AOI21xp33_ASAP7_75t_SL g651 ( .A1(n_576), .A2(n_547), .B(n_562), .Y(n_651) );
OAI21xp33_ASAP7_75t_L g652 ( .A1(n_619), .A2(n_562), .B(n_554), .Y(n_652) );
INVxp67_ASAP7_75t_L g653 ( .A(n_601), .Y(n_653) );
NAND2xp5_ASAP7_75t_L g654 ( .A(n_628), .B(n_551), .Y(n_654) );
OAI31xp33_ASAP7_75t_L g655 ( .A1(n_600), .A2(n_545), .A3(n_543), .B(n_540), .Y(n_655) );
INVx1_ASAP7_75t_L g656 ( .A(n_569), .Y(n_656) );
AND2x2_ASAP7_75t_L g657 ( .A(n_599), .B(n_540), .Y(n_657) );
INVx1_ASAP7_75t_L g658 ( .A(n_573), .Y(n_658) );
AOI21xp5_ASAP7_75t_L g659 ( .A1(n_618), .A2(n_538), .B(n_533), .Y(n_659) );
NAND2xp5_ASAP7_75t_L g660 ( .A(n_583), .B(n_519), .Y(n_660) );
NAND2xp5_ASAP7_75t_L g661 ( .A(n_583), .B(n_516), .Y(n_661) );
AOI221xp5_ASAP7_75t_L g662 ( .A1(n_600), .A2(n_511), .B1(n_509), .B2(n_498), .C(n_45), .Y(n_662) );
AOI22xp5_ASAP7_75t_L g663 ( .A1(n_625), .A2(n_596), .B1(n_581), .B2(n_568), .Y(n_663) );
NOR4xp25_ASAP7_75t_L g664 ( .A(n_617), .B(n_509), .C(n_43), .D(n_44), .Y(n_664) );
INVx1_ASAP7_75t_L g665 ( .A(n_572), .Y(n_665) );
OAI21xp5_ASAP7_75t_L g666 ( .A1(n_571), .A2(n_39), .B(n_46), .Y(n_666) );
NOR4xp25_ASAP7_75t_L g667 ( .A(n_613), .B(n_48), .C(n_57), .D(n_58), .Y(n_667) );
OAI21xp33_ASAP7_75t_L g668 ( .A1(n_640), .A2(n_594), .B(n_610), .Y(n_668) );
AOI311xp33_ASAP7_75t_L g669 ( .A1(n_645), .A2(n_579), .A3(n_574), .B(n_612), .C(n_578), .Y(n_669) );
AOI221xp5_ASAP7_75t_L g670 ( .A1(n_651), .A2(n_594), .B1(n_602), .B2(n_588), .C(n_591), .Y(n_670) );
INVx1_ASAP7_75t_L g671 ( .A(n_633), .Y(n_671) );
OAI221xp5_ASAP7_75t_L g672 ( .A1(n_632), .A2(n_626), .B1(n_622), .B2(n_609), .C(n_603), .Y(n_672) );
AOI222xp33_ASAP7_75t_L g673 ( .A1(n_653), .A2(n_609), .B1(n_585), .B2(n_606), .C1(n_607), .C2(n_592), .Y(n_673) );
AOI221xp5_ASAP7_75t_L g674 ( .A1(n_634), .A2(n_611), .B1(n_567), .B2(n_605), .C(n_581), .Y(n_674) );
AOI22xp5_ASAP7_75t_L g675 ( .A1(n_663), .A2(n_575), .B1(n_615), .B2(n_627), .Y(n_675) );
NAND2xp5_ASAP7_75t_L g676 ( .A(n_649), .B(n_589), .Y(n_676) );
AOI221xp5_ASAP7_75t_L g677 ( .A1(n_652), .A2(n_650), .B1(n_648), .B2(n_630), .C(n_646), .Y(n_677) );
AOI22xp5_ASAP7_75t_L g678 ( .A1(n_658), .A2(n_589), .B1(n_570), .B2(n_622), .Y(n_678) );
OAI22xp33_ASAP7_75t_L g679 ( .A1(n_641), .A2(n_595), .B1(n_582), .B2(n_598), .Y(n_679) );
NAND2xp33_ASAP7_75t_SL g680 ( .A(n_635), .B(n_629), .Y(n_680) );
AOI221xp5_ASAP7_75t_L g681 ( .A1(n_644), .A2(n_616), .B1(n_629), .B2(n_624), .C(n_64), .Y(n_681) );
AOI22xp5_ASAP7_75t_L g682 ( .A1(n_639), .A2(n_616), .B1(n_61), .B2(n_63), .Y(n_682) );
OAI22xp5_ASAP7_75t_L g683 ( .A1(n_637), .A2(n_70), .B1(n_71), .B2(n_72), .Y(n_683) );
NAND4xp25_ASAP7_75t_L g684 ( .A(n_662), .B(n_73), .C(n_74), .D(n_75), .Y(n_684) );
AOI21xp5_ASAP7_75t_L g685 ( .A1(n_647), .A2(n_76), .B(n_77), .Y(n_685) );
AOI22xp5_ASAP7_75t_L g686 ( .A1(n_639), .A2(n_78), .B1(n_80), .B2(n_81), .Y(n_686) );
NOR4xp25_ASAP7_75t_L g687 ( .A(n_662), .B(n_84), .C(n_87), .D(n_89), .Y(n_687) );
OAI221xp5_ASAP7_75t_SL g688 ( .A1(n_655), .A2(n_162), .B1(n_175), .B2(n_664), .C(n_659), .Y(n_688) );
OAI21xp33_ASAP7_75t_SL g689 ( .A1(n_631), .A2(n_162), .B(n_175), .Y(n_689) );
AOI221x1_ASAP7_75t_L g690 ( .A1(n_659), .A2(n_162), .B1(n_666), .B2(n_647), .C(n_656), .Y(n_690) );
NAND4xp25_ASAP7_75t_L g691 ( .A(n_643), .B(n_162), .C(n_660), .D(n_661), .Y(n_691) );
AND2x4_ASAP7_75t_L g692 ( .A(n_665), .B(n_636), .Y(n_692) );
NOR3xp33_ASAP7_75t_L g693 ( .A(n_643), .B(n_654), .C(n_667), .Y(n_693) );
NAND4xp75_ASAP7_75t_L g694 ( .A(n_638), .B(n_640), .C(n_576), .D(n_659), .Y(n_694) );
OAI31xp33_ASAP7_75t_L g695 ( .A1(n_642), .A2(n_645), .A3(n_580), .B(n_630), .Y(n_695) );
OAI21xp5_ASAP7_75t_SL g696 ( .A1(n_657), .A2(n_641), .B(n_580), .Y(n_696) );
INVx1_ASAP7_75t_L g697 ( .A(n_671), .Y(n_697) );
NAND2xp5_ASAP7_75t_L g698 ( .A(n_673), .B(n_693), .Y(n_698) );
NAND4xp25_ASAP7_75t_L g699 ( .A(n_688), .B(n_695), .C(n_690), .D(n_691), .Y(n_699) );
NAND3xp33_ASAP7_75t_L g700 ( .A(n_669), .B(n_677), .C(n_668), .Y(n_700) );
AOI22xp5_ASAP7_75t_L g701 ( .A1(n_694), .A2(n_696), .B1(n_672), .B2(n_674), .Y(n_701) );
AOI21xp5_ASAP7_75t_L g702 ( .A1(n_689), .A2(n_680), .B(n_687), .Y(n_702) );
CKINVDCx5p33_ASAP7_75t_R g703 ( .A(n_698), .Y(n_703) );
NAND3x1_ASAP7_75t_L g704 ( .A(n_701), .B(n_678), .C(n_682), .Y(n_704) );
NAND4xp25_ASAP7_75t_L g705 ( .A(n_700), .B(n_684), .C(n_681), .D(n_686), .Y(n_705) );
OAI22xp5_ASAP7_75t_L g706 ( .A1(n_702), .A2(n_675), .B1(n_670), .B2(n_679), .Y(n_706) );
HB1xp67_ASAP7_75t_L g707 ( .A(n_703), .Y(n_707) );
INVx2_ASAP7_75t_L g708 ( .A(n_704), .Y(n_708) );
NAND2xp5_ASAP7_75t_L g709 ( .A(n_706), .B(n_697), .Y(n_709) );
INVx1_ASAP7_75t_L g710 ( .A(n_707), .Y(n_710) );
INVx3_ASAP7_75t_L g711 ( .A(n_708), .Y(n_711) );
HB1xp67_ASAP7_75t_L g712 ( .A(n_710), .Y(n_712) );
INVx2_ASAP7_75t_L g713 ( .A(n_710), .Y(n_713) );
OAI22x1_ASAP7_75t_L g714 ( .A1(n_713), .A2(n_711), .B1(n_709), .B2(n_699), .Y(n_714) );
OAI21xp5_ASAP7_75t_L g715 ( .A1(n_712), .A2(n_711), .B(n_705), .Y(n_715) );
OAI21xp5_ASAP7_75t_L g716 ( .A1(n_715), .A2(n_711), .B(n_685), .Y(n_716) );
XNOR2x1_ASAP7_75t_L g717 ( .A(n_716), .B(n_714), .Y(n_717) );
OAI21xp5_ASAP7_75t_L g718 ( .A1(n_717), .A2(n_711), .B(n_676), .Y(n_718) );
OAI21xp5_ASAP7_75t_L g719 ( .A1(n_718), .A2(n_692), .B(n_683), .Y(n_719) );
endmodule